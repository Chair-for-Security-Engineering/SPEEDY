module SPEEDY_Rounds5_0 ( Ciphertext, Key, Plaintext );
  input [191:0] Ciphertext;
  input [191:0] Key;
  output [191:0] Plaintext;
  wire   n1, n2, n7, n10, n14, n16, n17, n19, n21, n22, n24, n26, n27, n29,
         n30, n31, n32, n33, n39, n40, n42, n44, n46, n48, n49, n50, n55, n57,
         n59, n60, n61, n63, n64, n65, n66, n67, n70, n73, n75, n77, n78, n79,
         n80, n81, n83, n84, n85, n87, n89, n91, n92, n93, n97, n98, n99, n100,
         n101, n103, n105, n106, n107, n109, n110, n111, n112, n114, n115,
         n118, n120, n124, n125, n127, n129, n130, n131, n132, n133, n137,
         n138, n139, n141, n144, n146, n147, n148, n149, n152, n153, n157,
         n159, n161, n162, n163, n169, n170, n171, n172, n173, n177, n178,
         n179, n180, n185, n187, n188, n189, n191, n193, n195, n197, n200,
         n201, n202, n204, n205, n208, n209, n211, n212, n213, n214, n215,
         n216, n217, n219, n222, n223, n224, n227, n231, n233, n238, n240,
         n242, n243, n244, n245, n246, n247, n248, n254, n255, n256, n258,
         n260, n261, n262, n263, n264, n266, n269, n270, n271, n273, n274,
         n275, n277, n279, n281, n282, n283, n284, n286, n287, n288, n291,
         n292, n295, n296, n298, n299, n300, n301, n302, n304, n305, n306,
         n307, n309, n312, n313, n314, n315, n317, n318, n320, n321, n322,
         n323, n324, n327, n328, n331, n333, n337, n339, n342, n344, n345,
         n348, n349, n351, n352, n353, n354, n356, n357, n358, n359, n362,
         n364, n365, n367, n372, n375, n376, n377, n381, n382, n383, n386,
         n387, n391, n392, n393, n399, n400, n401, n402, n403, n404, n406,
         n408, n409, n411, n412, n414, n416, n419, n423, n424, n426, n429,
         n430, n431, n432, n433, n434, n435, n436, n439, n440, n442, n445,
         n447, n449, n454, n455, n457, n461, n462, n463, n466, n467, n469,
         n470, n472, n473, n476, n478, n482, n483, n484, n485, n486, n489,
         n490, n491, n493, n495, n496, n499, n502, n504, n506, n507, n508,
         n517, n518, n521, n522, n523, n524, n525, n527, n531, n532, n533,
         n535, n536, n537, n540, n541, n543, n544, n545, n548, n550, n551,
         n555, n559, n560, n562, n565, n567, n569, n571, n574, n576, n577,
         n578, n579, n580, n582, n586, n588, n590, n591, n592, n594, n595,
         n596, n597, n599, n600, n601, n602, n603, n604, n605, n608, n609,
         n610, n611, n614, n616, n617, n618, n620, n622, n623, n624, n625,
         n627, n628, n630, n635, n637, n638, n639, n641, n645, n647, n648,
         n651, n652, n653, n656, n657, n658, n660, n664, n665, n666, n667,
         n670, n671, n672, n673, n674, n677, n678, n680, n682, n684, n685,
         n686, n687, n688, n689, n695, n696, n697, n699, n701, n703, n707,
         n708, n709, n710, n711, n715, n717, n718, n721, n724, n725, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n746, n747, n748, n750, n752,
         n753, n754, n755, n756, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n813, n814, n815, n816, n817, n818, n819, n820,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n833,
         n834, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n853, n854, n856, n857, n858, n859,
         n861, n863, n865, n866, n868, n869, n870, n872, n873, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n886, n887, n888,
         n889, n891, n892, n893, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n908, n909, n910, n911, n913, n914, n915,
         n916, n917, n918, n920, n921, n922, n925, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n940, n941, n942, n943,
         n944, n946, n948, n949, n951, n952, n953, n955, n957, n959, n960,
         n961, n963, n964, n965, n967, n968, n970, n971, n972, n973, n974,
         n976, n978, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1015, n1017, n1018, n1019, n1020, n1021, n1023, n1024,
         n1025, n1031, n1032, n1033, n1034, n1035, n1036, n1038, n1039, n1041,
         n1042, n1045, n1048, n1050, n1051, n1052, n1053, n1056, n1057, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1077, n1078, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1089, n1093, n1094, n1095, n1096, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1106, n1110, n1111, n1112, n1113,
         n1115, n1116, n1117, n1119, n1121, n1122, n1124, n1128, n1129, n1132,
         n1133, n1135, n1136, n1138, n1139, n1140, n1141, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1157,
         n1158, n1160, n1161, n1162, n1163, n1164, n1165, n1167, n1170, n1171,
         n1172, n1174, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1187, n1188, n1189, n1190, n1192, n1193, n1196, n1197, n1198,
         n1200, n1203, n1205, n1208, n1209, n1212, n1213, n1214, n1217, n1218,
         n1219, n1221, n1224, n1225, n1226, n1227, n1230, n1232, n1233, n1235,
         n1237, n1238, n1239, n1243, n1244, n1248, n1252, n1253, n1254, n1255,
         n1256, n1257, n1259, n1260, n1261, n1262, n1263, n1265, n1266, n1267,
         n1268, n1269, n1270, n1272, n1273, n1274, n1275, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1301, n1303, n1304, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1341, n1342, n1343, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1358, n1359, n1360, n1362, n1363, n1364, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1447, n1448, n1449, n1450, n1452, n1453,
         n1455, n1456, n1457, n1458, n1459, n1461, n1462, n1463, n1464, n1465,
         n1466, n1468, n1469, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1479, n1480, n1481, n1482, n1483, n1484, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1497, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1509, n1510, n1511, n1512,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1527, n1528, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1561, n1562, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1585, n1586, n1587, n1590, n1591,
         n1592, n1593, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1663, n1664, n1666, n1667, n1669,
         n1670, n1671, n1672, n1673, n1674, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1704, n1705, n1706, n1708, n1709, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1721, n1723, n1724, n1725, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1765, n1766, n1767, n1769, n1770, n1771, n1772,
         n1773, n1775, n1776, n1777, n1779, n1780, n1781, n1782, n1783, n1785,
         n1786, n1787, n1788, n1789, n1790, n1792, n1793, n1794, n1795, n1796,
         n1798, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1852, n1853, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1865, n1866, n1867,
         n1868, n1869, n1871, n1872, n1875, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1915, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1938, n1939, n1940, n1941, n1942, n1943, n1945, n1946, n1947, n1948,
         n1951, n1952, n1953, n1955, n1956, n1957, n1958, n1959, n1960, n1962,
         n1963, n1967, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1979,
         n1981, n1982, n1983, n1985, n1986, n1987, n1988, n1989, n1990, n1993,
         n1994, n1995, n1996, n1998, n1999, n2000, n2001, n2002, n2004, n2005,
         n2006, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2017, n2018,
         n2019, n2020, n2021, n2023, n2024, n2025, n2026, n2028, n2029, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2046, n2047, n2049, n2051, n2052, n2053, n2056, n2057, n2059,
         n2060, n2061, n2062, n2063, n2064, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2078, n2079, n2081, n2082,
         n2083, n2086, n2087, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2100, n2101, n2102, n2103, n2104, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2140, n2141, n2142,
         n2143, n2144, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2157, n2158, n2159, n2160, n2161, n2162, n2164, n2166, n2167,
         n2168, n2169, n2170, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2182, n2183, n2184, n2185, n2187, n2191, n2192, n2193,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2210, n2212, n2213, n2215, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2230, n2232, n2233, n2234, n2235,
         n2236, n2240, n2241, n2242, n2245, n2246, n2247, n2250, n2252, n2253,
         n2255, n2256, n2257, n2258, n2259, n2260, n2262, n2263, n2264, n2265,
         n2266, n2267, n2269, n2271, n2273, n2274, n2275, n2276, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2301, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2312,
         n2313, n2314, n2315, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2348, n2349, n2350, n2351, n2352, n2354, n2355, n2356,
         n2357, n2361, n2362, n2364, n2365, n2367, n2369, n2370, n2371, n2372,
         n2373, n2374, n2376, n2378, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2406, n2407,
         n2408, n2409, n2410, n2412, n2413, n2416, n2417, n2418, n2419, n2420,
         n2422, n2425, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2448, n2450, n2451, n2452, n2453, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2472, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2489, n2490, n2491, n2493, n2494,
         n2495, n2496, n2499, n2500, n2501, n2502, n2504, n2505, n2506, n2507,
         n2508, n2510, n2511, n2512, n2513, n2514, n2516, n2519, n2522, n2524,
         n2530, n2531, n2532, n2533, n2535, n2538, n2540, n2541, n2542, n2543,
         n2544, n2546, n2547, n2548, n2550, n2551, n2553, n2557, n2560, n2561,
         n2562, n2564, n2565, n2567, n2568, n2569, n2570, n2571, n2572, n2574,
         n2576, n2578, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2607, n2608, n2609, n2610,
         n2612, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2625, n2626, n2628, n2629, n2630, n2631, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2644, n2645, n2646,
         n2647, n2650, n2651, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2674, n2675, n2676, n2677, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2697, n2698, n2699, n2700, n2701, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2712, n2713, n2714, n2715, n2716, n2717, n2719,
         n2721, n2722, n2723, n2724, n2726, n2727, n2729, n2730, n2731, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2769, n2770, n2771, n2772, n2775, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2800, n2801,
         n2803, n2804, n2805, n2806, n2807, n2810, n2811, n2812, n2814, n2816,
         n2817, n2820, n2821, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2840,
         n2841, n2842, n2843, n2846, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2870, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2889, n2890, n2891,
         n2892, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2911, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2928,
         n2929, n2930, n2933, n2934, n2935, n2937, n2939, n2940, n2941, n2942,
         n2944, n2947, n2948, n2950, n2951, n2952, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2965, n2968, n2970, n2971,
         n2973, n2974, n2975, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2987, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3001, n3003, n3004, n3005, n3006, n3007, n3009, n3010,
         n3011, n3012, n3013, n3015, n3018, n3019, n3021, n3022, n3023, n3025,
         n3026, n3027, n3029, n3030, n3031, n3032, n3033, n3035, n3036, n3037,
         n3038, n3039, n3042, n3043, n3044, n3046, n3047, n3048, n3049, n3050,
         n3052, n3053, n3054, n3055, n3057, n3059, n3060, n3061, n3064, n3065,
         n3069, n3070, n3071, n3072, n3073, n3076, n3077, n3078, n3080, n3081,
         n3082, n3085, n3086, n3087, n3090, n3091, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3101, n3102, n3103, n3104, n3105, n3108, n3109,
         n3111, n3112, n3113, n3116, n3117, n3118, n3119, n3122, n3123, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3139, n3140, n3142, n3145, n3148, n3149, n3150, n3151, n3154, n3155,
         n3156, n3159, n3161, n3162, n3163, n3164, n3165, n3167, n3168, n3169,
         n3171, n3172, n3173, n3174, n3175, n3177, n3178, n3180, n3181, n3182,
         n3183, n3184, n3185, n3187, n3188, n3190, n3191, n3193, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3227, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3274,
         n3275, n3277, n3279, n3281, n3282, n3284, n3285, n3287, n3288, n3289,
         n3290, n3291, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3310, n3311,
         n3313, n3314, n3315, n3316, n3317, n3318, n3320, n3322, n3323, n3324,
         n3325, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3338, n3339, n3340, n3341, n3344, n3345, n3346, n3347, n3348, n3350,
         n3351, n3352, n3353, n3354, n3356, n3357, n3358, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3379, n3380, n3381, n3382, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3402, n3403, n3404, n3405, n3406, n3407, n3409,
         n3410, n3412, n3413, n3414, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3440, n3441, n3442, n3443,
         n3444, n3445, n3448, n3449, n3450, n3451, n3452, n3453, n3455, n3457,
         n3458, n3459, n3460, n3461, n3462, n3464, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3482, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3495, n3497, n3499, n3500, n3501, n3503, n3504, n3505,
         n3507, n3510, n3511, n3512, n3513, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3540, n3541, n3543,
         n3544, n3545, n3547, n3548, n3549, n3550, n3551, n3553, n3555, n3556,
         n3559, n3560, n3561, n3562, n3563, n3564, n3566, n3567, n3568, n3570,
         n3571, n3572, n3573, n3574, n3575, n3578, n3579, n3580, n3581, n3582,
         n3583, n3585, n3588, n3589, n3590, n3591, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3602, n3603, n3604, n3605, n3606, n3607,
         n3609, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3625, n3626, n3628, n3630, n3631, n3633, n3634,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3656, n3657, n3658, n3659,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3677, n3678, n3679, n3680, n3681,
         n3684, n3685, n3686, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3705, n3706, n3707,
         n3708, n3710, n3713, n3715, n3716, n3717, n3718, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3728, n3729, n3730, n3732, n3733, n3734,
         n3735, n3737, n3738, n3739, n3741, n3743, n3745, n3746, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3775, n3776, n3777, n3780, n3781, n3782, n3785, n3786, n3787, n3789,
         n3790, n3793, n3794, n3797, n3798, n3799, n3800, n3804, n3806, n3807,
         n3808, n3809, n3811, n3813, n3814, n3815, n3816, n3817, n3818, n3820,
         n3821, n3822, n3823, n3824, n3825, n3827, n3828, n3829, n3830, n3831,
         n3835, n3836, n3837, n3838, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3849, n3852, n3853, n3854, n3855, n3856, n3857, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3868, n3869, n3870, n3871,
         n3875, n3878, n3879, n3881, n3884, n3885, n3887, n3888, n3889, n3890,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3907, n3908, n3910, n3911, n3913, n3914, n3916, n3917,
         n3918, n3919, n3920, n3921, n3923, n3925, n3927, n3928, n3929, n3930,
         n3932, n3933, n3934, n3935, n3937, n3938, n3939, n3940, n3941, n3942,
         n3944, n3945, n3946, n3947, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3969, n3970, n3971, n3975, n3976, n3979, n3980, n3981, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3999, n4001, n4002, n4003, n4005, n4006, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4017, n4018, n4019, n4020,
         n4021, n4023, n4024, n4025, n4027, n4029, n4030, n4031, n4033, n4034,
         n4035, n4036, n4037, n4038, n4041, n4042, n4043, n4046, n4047, n4048,
         n4049, n4051, n4052, n4054, n4055, n4056, n4057, n4059, n4061, n4062,
         n4063, n4064, n4065, n4068, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4090, n4091, n4092, n4093, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4109, n4111, n4112,
         n4115, n4116, n4117, n4118, n4119, n4121, n4123, n4124, n4125, n4126,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4156, n4157, n4158, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4178, n4181, n4182, n4183, n4184, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4224, n4226, n4227, n4228, n4229, n4231, n4232,
         n4233, n4234, n4237, n4238, n4239, n4240, n4241, n4243, n4244, n4245,
         n4248, n4249, n4250, n4252, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4268, n4269, n4270,
         n4271, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4304,
         n4305, n4308, n4310, n4311, n4312, n4313, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4326, n4327, n4328, n4329,
         n4331, n4332, n4333, n4334, n4335, n4336, n4339, n4340, n4341, n4342,
         n4343, n4344, n4346, n4347, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4361, n4362, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4373, n4374, n4375, n4376, n4378, n4380,
         n4383, n4386, n4387, n4388, n4389, n4391, n4392, n4393, n4394, n4395,
         n4396, n4398, n4399, n4403, n4404, n4405, n4409, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4420, n4422, n4424, n4425, n4428, n4430,
         n4431, n4433, n4436, n4437, n4439, n4440, n4441, n4442, n4443, n4444,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4457,
         n4459, n4460, n4463, n4464, n4465, n4466, n4467, n4468, n4470, n4473,
         n4476, n4477, n4479, n4480, n4481, n4482, n4483, n4485, n4487, n4488,
         n4489, n4491, n4493, n4495, n4496, n4497, n4499, n4503, n4504, n4506,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4519, n4521, n4522,
         n4525, n4526, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4537,
         n4538, n4539, n4540, n4541, n4543, n4544, n4546, n4547, n4548, n4549,
         n4551, n4556, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4579, n4580, n4581, n4584, n4585, n4587, n4588, n4589, n4591,
         n4592, n4594, n4595, n4598, n4601, n4602, n4604, n4606, n4607, n4609,
         n4611, n4613, n4614, n4615, n4616, n4617, n4619, n4620, n4621, n4622,
         n4623, n4624, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4654, n4655, n4657,
         n4658, n4659, n4660, n4661, n4663, n4664, n4666, n4667, n4669, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4695, n4696, n4697, n4699, n4700, n4701, n4703, n4706, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4721, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4740, n4743, n4744, n4745, n4746, n4747, n4748, n4751, n4754,
         n4756, n4757, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4769,
         n4771, n4773, n4774, n4775, n4776, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4787, n4789, n4790, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4805, n4806, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4819, n4821, n4822,
         n4824, n4825, n4826, n4827, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4838, n4839, n4840, n4842, n4844, n4845, n4846, n4847, n4848,
         n4850, n4851, n4852, n4853, n4854, n4855, n4858, n4859, n4860, n4863,
         n4864, n4865, n4867, n4868, n4869, n4870, n4871, n4873, n4874, n4876,
         n4879, n4880, n4881, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4897, n4898, n4899, n4900, n4901,
         n4903, n4904, n4907, n4908, n4911, n4914, n4915, n4917, n4918, n4919,
         n4921, n4922, n4924, n4926, n4928, n4929, n4930, n4933, n4934, n4936,
         n4937, n4938, n4940, n4941, n4943, n4945, n4947, n4949, n4950, n4951,
         n4952, n4953, n4955, n4956, n4958, n4960, n4961, n4962, n4963, n4964,
         n4967, n4968, n4969, n4971, n4972, n4973, n4977, n4978, n4980, n4981,
         n4982, n4984, n4985, n4986, n4988, n4989, n4990, n4991, n4993, n4995,
         n4996, n4998, n4999, n5000, n5001, n5003, n5004, n5005, n5008, n5009,
         n5011, n5013, n5017, n5019, n5020, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5033, n5037, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5048, n5049, n5050, n5051, n5053, n5054, n5055,
         n5056, n5057, n5059, n5060, n5061, n5062, n5063, n5065, n5068, n5069,
         n5070, n5072, n5073, n5075, n5076, n5078, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5098, n5099, n5100, n5101, n5103, n5104, n5105, n5107, n5108,
         n5109, n5110, n5112, n5113, n5114, n5115, n5117, n5118, n5119, n5120,
         n5122, n5123, n5124, n5125, n5126, n5127, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5152, n5153, n5154, n5155,
         n5156, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5169, n5170, n5171, n5172, n5173, n5175, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5192, n5193, n5194, n5195, n5196, n5198, n5199, n5200, n5202, n5203,
         n5204, n5205, n5206, n5208, n5209, n5210, n5211, n5212, n5214, n5215,
         n5216, n5217, n5218, n5219, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5231, n5232, n5233, n5234, n5235, n5236, n5238, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5250, n5251, n5252, n5253,
         n5254, n5255, n5258, n5259, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5271, n5272, n5273, n5275, n5276, n5277, n5278, n5279,
         n5280, n5282, n5283, n5284, n5285, n5287, n5289, n5290, n5291, n5292,
         n5293, n5294, n5296, n5297, n5298, n5299, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5315, n5316,
         n5317, n5318, n5319, n5322, n5323, n5324, n5326, n5327, n5328, n5330,
         n5332, n5333, n5334, n5335, n5336, n5337, n5339, n5340, n5341, n5342,
         n5343, n5345, n5346, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5362, n5363, n5364, n5365,
         n5367, n5368, n5369, n5371, n5373, n5374, n5376, n5377, n5382, n5383,
         n5384, n5385, n5386, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5414, n5415, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5481, n5482, n5483, n5484,
         n5487, n5488, n5489, n5490, n5491, n5493, n5494, n5495, n5496, n5497,
         n5498, n5502, n5505, n5506, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5527, n5528, n5529, n5531, n5532, n5533, n5534, n5536,
         n5537, n5541, n5543, n5544, n5545, n5547, n5548, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5560, n5561, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5591, n5593, n5594, n5595, n5596, n5597, n5599, n5600,
         n5602, n5603, n5604, n5607, n5609, n5610, n5611, n5612, n5614, n5615,
         n5619, n5620, n5621, n5622, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5649, n5650, n5651, n5652, n5653,
         n5654, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5672, n5673, n5674, n5675,
         n5676, n5678, n5679, n5680, n5681, n5682, n5684, n5685, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5696, n5697, n5698, n5699, n5700,
         n5701, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5740, n5741, n5742, n5743, n5744,
         n5745, n5747, n5748, n5749, n5752, n5754, n5755, n5757, n5758, n5760,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5785, n5786, n5787, n5788, n5790, n5791, n5792, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5805, n5806, n5807,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5818, n5819,
         n5822, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5833, n5834,
         n5836, n5837, n5838, n5839, n5841, n5842, n5846, n5847, n5848, n5849,
         n5851, n5853, n5854, n5855, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5883, n5884, n5885, n5886,
         n5887, n5889, n5890, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5902, n5903, n5906, n5907, n5908, n5909, n5910, n5911,
         n5913, n5914, n5917, n5919, n5920, n5922, n5923, n5924, n5927, n5928,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5957, n5958, n5959, n5960,
         n5961, n5963, n5964, n5965, n5966, n5968, n5969, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5995,
         n5996, n5997, n5999, n6000, n6001, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6024, n6025, n6026, n6027, n6028, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6040, n6041, n6043,
         n6045, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6065, n6067,
         n6068, n6070, n6071, n6072, n6073, n6075, n6076, n6077, n6078, n6080,
         n6081, n6082, n6083, n6084, n6085, n6087, n6088, n6089, n6090, n6091,
         n6092, n6095, n6096, n6097, n6098, n6100, n6101, n6102, n6103, n6105,
         n6106, n6107, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6148, n6149,
         n6150, n6151, n6152, n6153, n6157, n6159, n6160, n6161, n6162, n6164,
         n6166, n6167, n6168, n6170, n6171, n6173, n6174, n6177, n6178, n6179,
         n6180, n6181, n6184, n6187, n6188, n6191, n6192, n6194, n6195, n6197,
         n6198, n6199, n6200, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6235, n6236, n6237, n6238, n6241, n6243, n6244, n6245,
         n6247, n6248, n6250, n6251, n6252, n6253, n6255, n6256, n6257, n6259,
         n6260, n6262, n6268, n6269, n6270, n6271, n6273, n6274, n6275, n6276,
         n6277, n6280, n6281, n6282, n6283, n6284, n6285, n6288, n6289, n6290,
         n6291, n6293, n6294, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6311, n6312, n6313,
         n6314, n6316, n6317, n6318, n6319, n6321, n6322, n6323, n6324, n6326,
         n6329, n6330, n6331, n6332, n6333, n6336, n6337, n6338, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6403, n6404, n6405, n6406, n6407, n6408,
         n6410, n6411, n6412, n6414, n6415, n6416, n6417, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6431, n6432, n6435,
         n6437, n6438, n6439, n6440, n6441, n6442, n6444, n6445, n6447, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6462, n6463,
         n6464, n6465, n6467, n6469, n6473, n6474, n6475, n6481, n6482, n6483,
         n6484, n6486, n6489, n6490, n6491, n6493, n6494, n6495, n6496, n6497,
         n6498, n6500, n6501, n6502, n6504, n6505, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6519, n6520, n6522,
         n6523, n6524, n6526, n6527, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6544, n6545,
         n6546, n6547, n6548, n6549, n6551, n6552, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6570, n6571, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6592, n6593, n6595, n6596, n6597, n6598, n6599, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6615, n6616, n6617, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6632, n6633, n6635, n6636, n6638, n6639,
         n6640, n6641, n6643, n6644, n6645, n6647, n6649, n6651, n6654, n6655,
         n6656, n6657, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6669, n6670, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6682, n6684, n6685, n6686, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6698, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6711, n6713, n6714, n6715, n6716, n6717, n6718,
         n6720, n6721, n6722, n6723, n6725, n6726, n6727, n6728, n6730, n6731,
         n6732, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6742, n6743,
         n6744, n6745, n6747, n6748, n6749, n6750, n6751, n6752, n6754, n6755,
         n6756, n6758, n6759, n6760, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6784, n6785, n6786, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6799, n6800, n6801, n6803, n6804,
         n6805, n6807, n6808, n6809, n6810, n6812, n6813, n6815, n6816, n6817,
         n6818, n6820, n6822, n6823, n6824, n6825, n6826, n6827, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6838, n6839, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6852, n6853,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6865,
         n6866, n6867, n6868, n6869, n6871, n6872, n6873, n6874, n6875, n6876,
         n6878, n6879, n6880, n6881, n6883, n6885, n6886, n6888, n6889, n6890,
         n6891, n6892, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6906, n6907, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6917, n6918, n6919, n6920, n6922, n6923, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6940, n6941, n6943, n6944, n6946, n6947, n6949, n6950,
         n6952, n6953, n6954, n6955, n6956, n6957, n6959, n6960, n6961, n6963,
         n6965, n6967, n6968, n6969, n6971, n6973, n6974, n6975, n6977, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6987, n6988, n6989, n6990,
         n6991, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7001, n7002,
         n7004, n7005, n7006, n7007, n7008, n7009, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7040, n7041, n7042, n7043, n7047, n7048, n7049, n7050, n7051,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7067, n7068, n7069, n7070, n7071, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7084, n7086, n7087, n7092,
         n7093, n7094, n7095, n7096, n7098, n7099, n7100, n7102, n7103, n7104,
         n7105, n7106, n7109, n7110, n7111, n7112, n7113, n7115, n7116, n7117,
         n7118, n7120, n7123, n7125, n7127, n7129, n7130, n7132, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7159, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7171, n7172, n7173,
         n7174, n7175, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7190, n7191, n7192, n7194, n7195, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7211, n7212, n7213, n7214, n7215, n7216, n7218, n7219, n7220, n7222,
         n7225, n7226, n7228, n7229, n7230, n7231, n7232, n7234, n7235, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7249, n7252, n7253, n7254, n7256, n7257, n7258, n7259, n7260, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7277, n7280, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7292, n7293, n7295, n7296, n7297, n7298, n7299, n7300, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7311, n7313, n7314,
         n7315, n7317, n7318, n7320, n7321, n7322, n7323, n7324, n7326, n7327,
         n7328, n7331, n7332, n7333, n7335, n7336, n7337, n7338, n7340, n7341,
         n7342, n7343, n7345, n7346, n7347, n7348, n7349, n7350, n7352, n7354,
         n7355, n7356, n7358, n7359, n7360, n7361, n7362, n7363, n7365, n7366,
         n7367, n7370, n7371, n7373, n7374, n7375, n7376, n7377, n7380, n7381,
         n7383, n7385, n7386, n7388, n7389, n7390, n7392, n7394, n7395, n7396,
         n7397, n7398, n7400, n7401, n7402, n7403, n7404, n7405, n7408, n7410,
         n7414, n7415, n7417, n7418, n7420, n7421, n7423, n7424, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7441, n7442, n7444, n7445, n7446, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7456, n7459, n7461, n7462, n7463, n7464,
         n7465, n7466, n7468, n7469, n7474, n7475, n7477, n7481, n7483, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7494, n7495, n7496,
         n7499, n7500, n7501, n7502, n7504, n7506, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7522, n7525,
         n7527, n7528, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7544, n7546, n7548, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7571, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7593, n7594, n7595, n7596, n7598, n7600, n7601, n7602,
         n7603, n7604, n7605, n7607, n7608, n7610, n7612, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7622, n7626, n7627, n7628, n7629, n7630,
         n7632, n7633, n7634, n7635, n7637, n7639, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7660, n7661, n7662, n7663, n7666, n7668,
         n7672, n7673, n7674, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7702, n7703, n7705, n7708, n7710,
         n7711, n7713, n7714, n7715, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7727, n7728, n7729, n7730, n7731, n7732, n7735, n7736,
         n7737, n7738, n7741, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7752, n7753, n7754, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7771, n7772,
         n7773, n7774, n7775, n7776, n7778, n7779, n7782, n7784, n7785, n7786,
         n7787, n7788, n7789, n7791, n7794, n7795, n7797, n7799, n7800, n7801,
         n7802, n7803, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7816, n7817, n7818, n7819, n7821, n7823, n7824, n7826,
         n7827, n7828, n7829, n7830, n7831, n7834, n7835, n7836, n7838, n7839,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7896, n7902, n7903, n7904, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7923, n7924, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7935, n7937, n7941, n7942, n7943, n7944, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7969, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7993,
         n7995, n7996, n7997, n7998, n7999, n8000, n8002, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8012, n8014, n8015, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8035, n8036, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8068, n8069, n8070, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8080, n8081, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8093, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8108, n8109, n8110, n8111,
         n8113, n8114, n8115, n8116, n8117, n8119, n8120, n8121, n8122, n8123,
         n8125, n8126, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8141, n8142, n8143, n8144, n8146, n8147, n8148,
         n8149, n8150, n8152, n8153, n8155, n8156, n8157, n8158, n8159, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8173, n8174, n8175, n8177, n8178, n8179, n8180, n8181, n8182, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8208, n8209, n8211, n8212, n8213, n8214, n8215, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8236, n8237, n8238, n8239, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8254,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8266,
         n8267, n8268, n8269, n8270, n8271, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8285, n8287, n8288, n8289, n8290,
         n8292, n8293, n8294, n8295, n8296, n8298, n8299, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8311, n8312, n8314, n8315,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8335, n8336, n8337,
         n8338, n8340, n8341, n8342, n8343, n8344, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8359, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8371, n8372, n8373,
         n8374, n8375, n8377, n8378, n8380, n8381, n8384, n8385, n8386, n8387,
         n8389, n8391, n8392, n8394, n8395, n8396, n8397, n8398, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8408, n8409, n8410, n8411, n8412,
         n8413, n8415, n8416, n8417, n8418, n8419, n8420, n8422, n8423, n8424,
         n8425, n8426, n8427, n8429, n8430, n8431, n8432, n8433, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8452, n8453, n8454, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8483, n8484, n8485, n8486, n8487, n8489, n8492, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8502, n8505, n8506, n8507, n8508, n8509,
         n8511, n8513, n8514, n8516, n8517, n8518, n8520, n8521, n8522, n8523,
         n8525, n8526, n8527, n8528, n8529, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8556, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8567, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8578, n8579, n8581, n8582, n8583, n8584,
         n8586, n8587, n8588, n8589, n8590, n8591, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8606, n8608,
         n8609, n8612, n8613, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8628, n8629, n8630, n8631, n8632,
         n8633, n8636, n8637, n8639, n8640, n8642, n8643, n8645, n8646, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8662, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8678, n8679, n8680, n8683,
         n8684, n8685, n8687, n8688, n8689, n8690, n8691, n8692, n8694, n8695,
         n8696, n8697, n8699, n8700, n8701, n8702, n8703, n8704, n8706, n8707,
         n8708, n8710, n8711, n8713, n8714, n8715, n8716, n8719, n8720, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8744, n8745, n8746, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8756, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8769, n8770, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8784, n8785, n8786, n8788, n8789, n8790, n8791, n8792, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8810, n8811, n8812, n8813, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8832, n8833, n8835, n8836, n8837, n8839, n8840, n8841, n8842,
         n8843, n8844, n8846, n8847, n8848, n8850, n8851, n8852, n8853, n8854,
         n8856, n8858, n8859, n8860, n8861, n8862, n8864, n8865, n8866, n8868,
         n8869, n8870, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8882, n8884, n8885, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8895, n8896, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8911, n8912, n8913, n8914, n8915, n8917,
         n8918, n8919, n8921, n8922, n8923, n8924, n8929, n8931, n8932, n8933,
         n8934, n8936, n8937, n8938, n8940, n8941, n8942, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8968,
         n8969, n8973, n8974, n8975, n8976, n8977, n8979, n8981, n8982, n8983,
         n8984, n8985, n8986, n8989, n8990, n8992, n8994, n8995, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9005, n9007, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9017, n9018, n9019, n9022, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9034, n9035, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9049, n9050, n9051, n9052, n9055, n9056, n9057, n9058, n9059, n9060,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9071, n9072,
         n9075, n9076, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9105, n9106, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9166, n9167, n9168, n9169, n9170, n9173, n9175, n9176, n9177, n9178,
         n9179, n9180, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9205, n9207, n9208, n9209, n9211, n9212, n9214, n9215, n9216, n9217,
         n9219, n9221, n9222, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9236, n9238, n9240, n9241, n9242, n9243,
         n9244, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9263, n9264, n9265,
         n9266, n9267, n9269, n9273, n9274, n9277, n9278, n9279, n9280, n9281,
         n9283, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9301, n9302, n9304, n9306,
         n9307, n9311, n9314, n9315, n9316, n9317, n9318, n9319, n9321, n9322,
         n9323, n9324, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9334,
         n9335, n9337, n9338, n9339, n9340, n9342, n9343, n9344, n9345, n9346,
         n9350, n9351, n9353, n9354, n9355, n9356, n9357, n9358, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9424, n9426, n9427, n9428, n9429,
         n9430, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9440, n9442,
         n9443, n9444, n9445, n9446, n9447, n9449, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9459, n9460, n9461, n9462, n9463, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9499,
         n9500, n9501, n9503, n9504, n9505, n9506, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9517, n9519, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9538, n9539, n9540, n9541, n9542, n9543, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9579, n9580,
         n9581, n9582, n9583, n9584, n9586, n9587, n9588, n9589, n9590, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9605, n9606, n9607, n9608, n9609, n9610, n9613, n9615, n9616, n9617,
         n9618, n9619, n9621, n9622, n9627, n9628, n9629, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9641, n9642, n9643, n9646, n9648,
         n9649, n9650, n9652, n9653, n9654, n9655, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9671, n9672, n9673, n9674,
         n9675, n9677, n9679, n9682, n9683, n9685, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9695, n9696, n9697, n9698, n9700, n9701, n9702,
         n9703, n9704, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9729, n9730, n9731, n9736, n9737, n9739, n9740, n9742,
         n9743, n9744, n9745, n9746, n9748, n9749, n9751, n9752, n9753, n9755,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9775, n9776, n9777, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9801,
         n9802, n9803, n9804, n9805, n9806, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9836, n9837, n9839, n9842, n9843, n9845, n9847, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9858, n9860, n9861, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9878, n9880, n9882, n9883, n9884, n9885, n9886, n9888, n9889,
         n9890, n9891, n9892, n9894, n9896, n9898, n9899, n9904, n9907, n9908,
         n9909, n9910, n9912, n9913, n9914, n9915, n9917, n9918, n9920, n9922,
         n9924, n9925, n9926, n9928, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9940, n9941, n9943, n9945, n9946, n9947, n9948,
         n9953, n9954, n9956, n9959, n9962, n9963, n9967, n9968, n9969, n9971,
         n9972, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9983, n9984,
         n9986, n9987, n9988, n9989, n9991, n9992, n9993, n9995, n9997, n9998,
         n10000, n10001, n10003, n10004, n10005, n10008, n10010, n10013,
         n10015, n10016, n10017, n10019, n10021, n10022, n10023, n10024,
         n10025, n10027, n10030, n10031, n10032, n10033, n10035, n10036,
         n10038, n10040, n10041, n10043, n10044, n10045, n10046, n10047,
         n10049, n10052, n10053, n10055, n10056, n10057, n10058, n10060,
         n10061, n10062, n10063, n10064, n10065, n10067, n10068, n10069,
         n10070, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10084, n10085, n10086, n10087, n10088,
         n10090, n10091, n10095, n10096, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10110,
         n10111, n10112, n10113, n10115, n10116, n10117, n10118, n10119,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10131, n10132, n10133, n10134, n10137, n10138, n10139,
         n10140, n10141, n10145, n10148, n10150, n10151, n10152, n10153,
         n10155, n10156, n10157, n10159, n10160, n10165, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10183, n10184, n10185, n10187, n10190,
         n10191, n10192, n10193, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10205, n10206, n10210, n10211,
         n10214, n10217, n10218, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10232, n10233, n10235, n10236, n10237,
         n10239, n10240, n10241, n10243, n10244, n10245, n10247, n10248,
         n10250, n10251, n10252, n10253, n10254, n10255, n10258, n10263,
         n10264, n10265, n10267, n10268, n10269, n10270, n10271, n10273,
         n10274, n10275, n10277, n10278, n10279, n10282, n10283, n10284,
         n10285, n10286, n10288, n10289, n10291, n10292, n10293, n10294,
         n10295, n10298, n10299, n10300, n10302, n10303, n10304, n10305,
         n10307, n10309, n10310, n10311, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10324, n10325, n10327,
         n10328, n10329, n10333, n10334, n10335, n10337, n10339, n10340,
         n10341, n10344, n10345, n10346, n10347, n10348, n10349, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10360,
         n10361, n10362, n10363, n10364, n10366, n10367, n10368, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10381, n10383, n10389, n10390, n10391, n10393, n10394,
         n10395, n10397, n10398, n10399, n10401, n10402, n10403, n10404,
         n10405, n10406, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10419, n10420, n10422, n10425,
         n10426, n10427, n10428, n10430, n10431, n10434, n10436, n10437,
         n10441, n10442, n10443, n10445, n10446, n10447, n10448, n10449,
         n10450, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10461, n10463, n10464, n10466, n10469, n10470, n10472,
         n10473, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10490,
         n10492, n10493, n10494, n10495, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10510, n10512, n10513, n10515, n10517, n10519, n10521, n10522,
         n10523, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10535, n10536, n10537, n10538, n10539, n10540,
         n10542, n10543, n10544, n10545, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10562, n10563, n10566, n10567,
         n10569, n10571, n10572, n10573, n10574, n10575, n10577, n10578,
         n10579, n10580, n10583, n10584, n10585, n10587, n10590, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10606, n10608, n10611, n10613, n10615, n10617,
         n10618, n10619, n10620, n10621, n10622, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10634, n10635,
         n10636, n10637, n10639, n10640, n10641, n10642, n10643, n10645,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10656, n10658, n10660, n10661, n10662, n10663, n10664, n10665,
         n10668, n10669, n10670, n10671, n10673, n10675, n10676, n10677,
         n10678, n10680, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10694, n10698, n10699, n10700,
         n10703, n10705, n10706, n10707, n10708, n10709, n10711, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10721, n10722,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10780, n10781, n10782,
         n10783, n10784, n10786, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10798, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10815, n10816, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10847,
         n10848, n10849, n10852, n10853, n10855, n10858, n10859, n10860,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10882, n10883, n10884, n10885, n10887, n10888,
         n10889, n10891, n10893, n10894, n10896, n10897, n10898, n10899,
         n10900, n10902, n10904, n10906, n10907, n10908, n10909, n10910,
         n10911, n10914, n10915, n10917, n10918, n10919, n10920, n10922,
         n10923, n10924, n10925, n10926, n10927, n10930, n10932, n10933,
         n10936, n10937, n10938, n10939, n10941, n10942, n10944, n10945,
         n10946, n10947, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10975, n10976, n10977, n10978, n10979, n10981,
         n10983, n10984, n10985, n10986, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11101, n11102, n11104, n11105, n11106,
         n11108, n11110, n11111, n11113, n11114, n11118, n11119, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11142, n11143, n11144, n11145, n11147,
         n11149, n11150, n11153, n11154, n11155, n11156, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11169, n11170, n11171, n11172, n11174, n11175, n11176, n11177,
         n11178, n11179, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11200, n11201, n11202, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11229, n11230, n11231,
         n11232, n11233, n11234, n11236, n11237, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11252, n11254, n11255, n11256, n11260, n11261, n11262,
         n11263, n11264, n11265, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11278, n11279, n11280,
         n11281, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11304, n11305, n11307,
         n11309, n11310, n11311, n11312, n11314, n11316, n11317, n11318,
         n11319, n11321, n11322, n11323, n11324, n11325, n11327, n11328,
         n11329, n11333, n11336, n11337, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11372, n11373, n11374, n11375, n11378, n11380, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11390, n11391, n11393,
         n11394, n11395, n11396, n11397, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11409, n11410, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11423, n11424, n11425,
         n11426, n11427, n11429, n11430, n11433, n11434, n11435, n11436,
         n11437, n11439, n11440, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11452, n11455, n11456, n11457, n11458,
         n11459, n11460, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11483, n11484, n11485,
         n11486, n11487, n11488, n11490, n11492, n11493, n11494, n11495,
         n11497, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11513, n11514, n11515,
         n11516, n11517, n11519, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11534,
         n11536, n11537, n11538, n11539, n11542, n11543, n11544, n11545,
         n11546, n11548, n11549, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11561, n11562, n11563, n11564, n11565,
         n11566, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11577, n11578, n11579, n11580, n11581, n11582, n11586,
         n11587, n11588, n11589, n11590, n11592, n11593, n11594, n11595,
         n11599, n11600, n11601, n11605, n11606, n11607, n11608, n11609,
         n11610, n11612, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11627, n11628,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11649, n11650, n11652, n11654, n11655, n11656, n11657,
         n11658, n11659, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11675,
         n11676, n11677, n11678, n11679, n11680, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11691, n11692, n11693,
         n11698, n11699, n11700, n11701, n11702, n11704, n11705, n11708,
         n11709, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11725, n11726, n11727, n11728, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11741,
         n11742, n11743, n11744, n11746, n11747, n11748, n11749, n11750,
         n11751, n11753, n11754, n11755, n11756, n11757, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11792, n11793,
         n11794, n11795, n11797, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11828, n11829, n11830, n11831,
         n11832, n11833, n11835, n11836, n11837, n11838, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11863, n11864, n11866, n11867, n11868, n11869,
         n11870, n11871, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11890, n11891, n11892, n11893, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11903, n11904, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11945, n11946, n11947, n11948, n11949, n11950,
         n11954, n11955, n11956, n11957, n11959, n11961, n11962, n11963,
         n11965, n11967, n11968, n11970, n11971, n11973, n11975, n11977,
         n11978, n11980, n11981, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11992, n11993, n11994, n11995, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12033,
         n12034, n12036, n12037, n12038, n12039, n12040, n12042, n12043,
         n12044, n12045, n12049, n12050, n12051, n12052, n12055, n12056,
         n12057, n12058, n12060, n12062, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12076,
         n12077, n12078, n12080, n12081, n12082, n12084, n12085, n12086,
         n12087, n12088, n12089, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12114,
         n12116, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12127, n12128, n12129, n12130, n12131, n12133, n12134, n12135,
         n12137, n12140, n12141, n12142, n12143, n12145, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12194, n12195, n12196, n12197, n12198,
         n12199, n12201, n12203, n12205, n12206, n12208, n12209, n12210,
         n12212, n12214, n12215, n12216, n12220, n12221, n12225, n12226,
         n12227, n12229, n12230, n12231, n12232, n12234, n12235, n12236,
         n12237, n12239, n12240, n12243, n12244, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12257, n12258, n12260,
         n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
         n12271, n12272, n12273, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12304, n12307,
         n12310, n12312, n12313, n12314, n12315, n12317, n12318, n12320,
         n12321, n12322, n12323, n12325, n12327, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12384,
         n12386, n12387, n12389, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12419, n12420, n12421, n12422, n12423,
         n12424, n12426, n12428, n12430, n12431, n12432, n12433, n12434,
         n12436, n12439, n12440, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12464, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12477, n12478, n12479, n12480, n12482,
         n12483, n12484, n12486, n12487, n12489, n12491, n12492, n12493,
         n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501,
         n12502, n12503, n12504, n12505, n12506, n12507, n12509, n12511,
         n12512, n12513, n12514, n12515, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12539,
         n12540, n12541, n12542, n12543, n12545, n12546, n12547, n12548,
         n12549, n12550, n12552, n12553, n12554, n12555, n12556, n12557,
         n12558, n12559, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12595, n12596, n12597, n12598, n12599,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12614, n12615, n12616, n12618,
         n12619, n12620, n12624, n12625, n12626, n12629, n12630, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12665, n12666, n12667,
         n12668, n12669, n12673, n12674, n12675, n12676, n12677, n12679,
         n12680, n12681, n12682, n12685, n12686, n12687, n12688, n12689,
         n12690, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12714, n12715,
         n12716, n12717, n12720, n12722, n12723, n12725, n12727, n12728,
         n12729, n12730, n12731, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12779, n12780, n12781, n12782,
         n12783, n12785, n12786, n12787, n12788, n12789, n12791, n12794,
         n12797, n12798, n12799, n12800, n12803, n12804, n12805, n12806,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12838, n12840, n12841, n12842, n12843, n12844,
         n12845, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12868, n12869, n12871, n12872, n12874,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12887, n12889, n12890, n12891, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12907, n12908, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12927, n12929, n12930, n12932,
         n12933, n12935, n12936, n12937, n12938, n12940, n12941, n12942,
         n12943, n12944, n12945, n12947, n12948, n12952, n12953, n12954,
         n12955, n12956, n12957, n12959, n12960, n12961, n12962, n12963,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12995, n12996, n12997, n12998, n12999,
         n13000, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13018, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13052,
         n13053, n13054, n13055, n13056, n13057, n13059, n13060, n13061,
         n13062, n13064, n13067, n13068, n13069, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13102, n13103, n13104, n13105, n13107, n13108, n13109,
         n13112, n13114, n13115, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13131,
         n13132, n13133, n13135, n13136, n13137, n13138, n13139, n13141,
         n13142, n13143, n13144, n13145, n13147, n13148, n13149, n13151,
         n13152, n13153, n13155, n13156, n13159, n13162, n13163, n13164,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13187, n13188, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13213, n13214, n13215, n13216, n13218, n13219,
         n13220, n13221, n13225, n13228, n13229, n13230, n13232, n13233,
         n13234, n13235, n13237, n13238, n13239, n13240, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13251, n13254,
         n13255, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13270, n13272, n13274, n13276,
         n13277, n13278, n13280, n13281, n13283, n13284, n13285, n13286,
         n13288, n13289, n13290, n13291, n13292, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13319, n13320, n13321,
         n13322, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13338, n13339,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13350,
         n13352, n13353, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13372, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13452, n13453, n13454, n13456, n13457, n13458,
         n13459, n13460, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13475, n13476,
         n13478, n13479, n13480, n13481, n13482, n13483, n13485, n13486,
         n13487, n13489, n13490, n13492, n13493, n13496, n13497, n13498,
         n13500, n13501, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13522, n13524, n13525, n13526,
         n13527, n13528, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13541, n13544, n13545, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13557,
         n13558, n13559, n13561, n13562, n13563, n13564, n13565, n13566,
         n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
         n13575, n13576, n13578, n13579, n13580, n13581, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13599, n13600, n13601, n13603,
         n13605, n13607, n13608, n13609, n13610, n13613, n13614, n13615,
         n13616, n13618, n13619, n13620, n13621, n13622, n13623, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13638, n13639, n13640, n13642, n13643, n13645, n13647,
         n13650, n13651, n13652, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13666, n13667,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13712,
         n13713, n13714, n13716, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13737, n13739, n13740, n13742, n13743,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13755, n13756, n13757, n13759, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13778, n13780, n13781, n13782,
         n13783, n13785, n13786, n13787, n13788, n13790, n13792, n13793,
         n13794, n13795, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13817, n13818, n13819, n13821,
         n13822, n13823, n13824, n13825, n13826, n13828, n13830, n13831,
         n13832, n13833, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13850,
         n13851, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13862, n13863, n13864, n13865, n13866, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13877, n13878,
         n13879, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13909, n13911, n13912, n13914, n13915,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13925,
         n13926, n13928, n13929, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13942, n13943, n13944,
         n13945, n13947, n13949, n13950, n13952, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13978, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13992, n13994, n13996, n13997,
         n13998, n13999, n14002, n14003, n14004, n14005, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14036, n14037, n14038, n14039, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14049, n14050, n14051, n14052,
         n14054, n14055, n14056, n14058, n14059, n14060, n14061, n14062,
         n14063, n14064, n14065, n14067, n14068, n14069, n14070, n14072,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14095, n14096, n14097, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14114, n14115, n14118, n14119,
         n14120, n14121, n14122, n14127, n14128, n14129, n14131, n14132,
         n14133, n14134, n14135, n14136, n14138, n14139, n14141, n14142,
         n14143, n14144, n14145, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14174, n14176, n14177, n14178,
         n14180, n14181, n14183, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14196, n14199, n14200,
         n14201, n14202, n14203, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14235, n14236, n14238,
         n14240, n14241, n14242, n14243, n14245, n14246, n14247, n14249,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14298, n14299, n14300, n14301,
         n14302, n14303, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14319,
         n14320, n14322, n14323, n14324, n14325, n14326, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14339, n14341, n14342, n14343, n14344, n14345, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14356, n14357, n14358,
         n14359, n14360, n14361, n14363, n14364, n14365, n14366, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14382, n14383, n14384, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14407, n14408, n14409, n14411, n14412, n14414, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14454, n14456, n14457, n14458, n14459, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14477, n14478, n14480,
         n14481, n14482, n14484, n14485, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14508,
         n14510, n14512, n14513, n14514, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14541, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14555, n14556,
         n14558, n14560, n14561, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14573, n14574, n14575, n14576,
         n14577, n14578, n14580, n14581, n14582, n14583, n14584, n14586,
         n14587, n14588, n14589, n14590, n14593, n14594, n14595, n14596,
         n14597, n14600, n14601, n14602, n14603, n14604, n14605, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14626, n14627, n14628, n14629, n14630, n14633, n14635,
         n14636, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14650, n14651, n14654, n14655,
         n14656, n14657, n14658, n14659, n14661, n14662, n14663, n14665,
         n14666, n14667, n14668, n14669, n14671, n14672, n14674, n14675,
         n14676, n14677, n14678, n14679, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14728, n14729, n14730, n14731, n14732, n14733, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14778, n14779, n14780,
         n14782, n14783, n14784, n14785, n14786, n14787, n14789, n14792,
         n14793, n14794, n14796, n14797, n14798, n14800, n14801, n14803,
         n14804, n14806, n14807, n14808, n14809, n14810, n14811, n14813,
         n14814, n14815, n14816, n14818, n14819, n14820, n14824, n14825,
         n14826, n14827, n14828, n14831, n14833, n14834, n14836, n14837,
         n14839, n14840, n14841, n14842, n14843, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14884, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14899, n14900, n14901, n14903,
         n14904, n14905, n14906, n14908, n14909, n14910, n14911, n14913,
         n14914, n14915, n14916, n14918, n14919, n14920, n14921, n14922,
         n14924, n14925, n14927, n14929, n14930, n14931, n14934, n14935,
         n14936, n14937, n14938, n14940, n14941, n14943, n14944, n14945,
         n14946, n14947, n14948, n14950, n14951, n14952, n14953, n14954,
         n14955, n14958, n14960, n14961, n14962, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14973, n14974, n14975,
         n14977, n14978, n14980, n14981, n14982, n14985, n14986, n14987,
         n14988, n14990, n14991, n14993, n14994, n14997, n14999, n15000,
         n15001, n15002, n15003, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15015, n15016, n15017, n15018, n15020,
         n15021, n15022, n15023, n15025, n15026, n15028, n15029, n15030,
         n15031, n15032, n15033, n15034, n15036, n15038, n15039, n15040,
         n15041, n15043, n15044, n15045, n15046, n15047, n15051, n15053,
         n15054, n15055, n15056, n15058, n15059, n15060, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15078, n15079, n15081, n15082,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15099, n15100,
         n15101, n15102, n15105, n15108, n15109, n15110, n15111, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15122, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
         n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15152,
         n15153, n15154, n15155, n15156, n15157, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15170, n15171,
         n15173, n15174, n15175, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
         n15207, n15208, n15209, n15211, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15222, n15223, n15225, n15227,
         n15229, n15232, n15233, n15234, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15249,
         n15250, n15252, n15254, n15256, n15257, n15258, n15260, n15261,
         n15262, n15265, n15266, n15267, n15269, n15271, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15313, n15314, n15315, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15328, n15329,
         n15330, n15332, n15333, n15334, n15336, n15337, n15338, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15348, n15349,
         n15351, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15365, n15366, n15367, n15369,
         n15370, n15371, n15372, n15374, n15376, n15377, n15378, n15379,
         n15380, n15381, n15383, n15385, n15386, n15387, n15393, n15394,
         n15395, n15397, n15398, n15399, n15401, n15402, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15432, n15433, n15434, n15435, n15436, n15439, n15440,
         n15441, n15442, n15444, n15445, n15446, n15447, n15449, n15450,
         n15452, n15453, n15454, n15457, n15458, n15459, n15460, n15461,
         n15462, n15464, n15466, n15467, n15469, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15480, n15481, n15482,
         n15483, n15484, n15485, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15500,
         n15501, n15502, n15503, n15505, n15507, n15508, n15509, n15510,
         n15511, n15512, n15513, n15514, n15515, n15516, n15519, n15520,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15544, n15545, n15546, n15547, n15548, n15549,
         n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15560, n15561, n15562, n15563, n15564, n15566, n15567,
         n15568, n15569, n15571, n15572, n15573, n15574, n15575, n15576,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15599, n15601, n15602, n15603,
         n15605, n15606, n15609, n15610, n15611, n15612, n15613, n15614,
         n15615, n15616, n15617, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15642,
         n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
         n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
         n15661, n15662, n15663, n15664, n15665, n15666, n15669, n15670,
         n15671, n15672, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15689, n15690, n15692, n15693, n15695, n15697, n15698, n15699,
         n15700, n15701, n15703, n15704, n15705, n15706, n15707, n15708,
         n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,
         n15717, n15718, n15719, n15720, n15722, n15723, n15724, n15725,
         n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
         n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
         n15742, n15743, n15745, n15746, n15747, n15748, n15749, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15761, n15762,
         n15763, n15765, n15766, n15768, n15769, n15770, n15771, n15772,
         n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780,
         n15781, n15782, n15783, n15784, n15785, n15786, n15788, n15789,
         n15790, n15791, n15792, n15793, n15794, n15795, n15797, n15798,
         n15799, n15800, n15801, n15802, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15813, n15814, n15815, n15816,
         n15817, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15828, n15829, n15830, n15831, n15832, n15834, n15835,
         n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15844,
         n15845, n15846, n15847, n15848, n15849, n15850, n15853, n15854,
         n15856, n15857, n15858, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15869, n15870, n15871, n15872, n15873, n15875,
         n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
         n15885, n15886, n15888, n15889, n15890, n15892, n15893, n15894,
         n15896, n15897, n15898, n15899, n15902, n15903, n15904, n15906,
         n15907, n15908, n15909, n15912, n15913, n15914, n15915, n15916,
         n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15937, n15938, n15940, n15941, n15942,
         n15943, n15944, n15945, n15946, n15947, n15949, n15950, n15951,
         n15953, n15955, n15957, n15958, n15960, n15961, n15962, n15963,
         n15964, n15966, n15967, n15968, n15969, n15970, n15971, n15972,
         n15974, n15975, n15976, n15978, n15979, n15981, n15982, n15983,
         n15984, n15985, n15986, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15998, n15999, n16001, n16002,
         n16004, n16006, n16007, n16008, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16020, n16021, n16024,
         n16025, n16026, n16027, n16028, n16030, n16032, n16034, n16035,
         n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043,
         n16045, n16046, n16047, n16048, n16049, n16050, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16062,
         n16063, n16065, n16066, n16068, n16069, n16071, n16072, n16073,
         n16074, n16076, n16077, n16079, n16080, n16081, n16082, n16083,
         n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
         n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16101,
         n16102, n16103, n16106, n16107, n16108, n16109, n16110, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16122, n16123, n16125, n16126, n16127, n16128, n16132, n16133,
         n16134, n16135, n16136, n16138, n16139, n16140, n16142, n16143,
         n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
         n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159,
         n16160, n16161, n16162, n16163, n16164, n16168, n16171, n16172,
         n16173, n16174, n16175, n16176, n16177, n16179, n16181, n16182,
         n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190,
         n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198,
         n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206,
         n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16215,
         n16217, n16218, n16219, n16220, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16260, n16261, n16262, n16263, n16264, n16266, n16267, n16268,
         n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16278,
         n16279, n16280, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16346, n16347, n16349, n16353, n16354, n16355, n16357, n16358,
         n16360, n16361, n16363, n16365, n16366, n16367, n16368, n16369,
         n16370, n16372, n16373, n16375, n16376, n16377, n16378, n16379,
         n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387,
         n16388, n16389, n16391, n16392, n16393, n16394, n16395, n16396,
         n16397, n16398, n16400, n16401, n16402, n16403, n16404, n16406,
         n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415,
         n16416, n16418, n16419, n16420, n16421, n16422, n16423, n16425,
         n16426, n16427, n16428, n16430, n16431, n16432, n16434, n16435,
         n16436, n16437, n16438, n16439, n16440, n16442, n16443, n16444,
         n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452,
         n16453, n16455, n16456, n16457, n16458, n16459, n16460, n16461,
         n16462, n16464, n16465, n16466, n16467, n16468, n16469, n16470,
         n16471, n16472, n16473, n16474, n16475, n16476, n16480, n16481,
         n16483, n16484, n16485, n16486, n16487, n16489, n16490, n16491,
         n16492, n16493, n16494, n16496, n16497, n16500, n16501, n16502,
         n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510,
         n16511, n16513, n16514, n16515, n16516, n16517, n16518, n16519,
         n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527,
         n16528, n16529, n16530, n16531, n16532, n16533, n16535, n16536,
         n16538, n16539, n16540, n16542, n16543, n16545, n16546, n16547,
         n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555,
         n16556, n16557, n16558, n16559, n16561, n16562, n16563, n16564,
         n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16573,
         n16574, n16576, n16578, n16579, n16580, n16581, n16582, n16583,
         n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591,
         n16592, n16593, n16594, n16595, n16596, n16597, n16599, n16601,
         n16603, n16604, n16605, n16606, n16607, n16608, n16610, n16611,
         n16612, n16613, n16614, n16616, n16617, n16618, n16619, n16620,
         n16621, n16622, n16624, n16625, n16626, n16627, n16628, n16629,
         n16630, n16631, n16632, n16633, n16634, n16635, n16637, n16638,
         n16639, n16641, n16642, n16643, n16644, n16645, n16646, n16647,
         n16648, n16649, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16688, n16689, n16690,
         n16691, n16692, n16694, n16695, n16696, n16698, n16700, n16701,
         n16702, n16703, n16705, n16706, n16707, n16708, n16709, n16710,
         n16711, n16712, n16713, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16738, n16739, n16740, n16741, n16742, n16744, n16745, n16746,
         n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754,
         n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762,
         n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771,
         n16772, n16773, n16775, n16776, n16777, n16778, n16779, n16780,
         n16782, n16783, n16786, n16787, n16788, n16789, n16790, n16791,
         n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799,
         n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16808,
         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
         n16819, n16820, n16821, n16823, n16824, n16827, n16828, n16829,
         n16830, n16831, n16832, n16833, n16835, n16836, n16837, n16838,
         n16840, n16842, n16843, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16856, n16857, n16858,
         n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866,
         n16867, n16868, n16869, n16870, n16872, n16873, n16876, n16877,
         n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885,
         n16886, n16887, n16888, n16890, n16891, n16892, n16893, n16894,
         n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902,
         n16903, n16904, n16906, n16907, n16908, n16909, n16910, n16911,
         n16912, n16914, n16915, n16916, n16917, n16919, n16920, n16921,
         n16922, n16925, n16929, n16930, n16932, n16933, n16935, n16936,
         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
         n16945, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16968, n16969, n16970,
         n16971, n16972, n16974, n16976, n16978, n16979, n16980, n16981,
         n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989,
         n16990, n16991, n16992, n16993, n16994, n16995, n16997, n16998,
         n17000, n17002, n17003, n17004, n17005, n17006, n17008, n17009,
         n17010, n17012, n17013, n17015, n17016, n17017, n17018, n17019,
         n17020, n17023, n17024, n17025, n17026, n17027, n17028, n17029,
         n17030, n17032, n17033, n17034, n17035, n17036, n17037, n17038,
         n17039, n17040, n17041, n17042, n17043, n17046, n17047, n17048,
         n17051, n17053, n17054, n17055, n17056, n17057, n17058, n17059,
         n17060, n17061, n17063, n17064, n17069, n17070, n17071, n17072,
         n17073, n17076, n17077, n17078, n17079, n17080, n17081, n17082,
         n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090,
         n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098,
         n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
         n17108, n17109, n17110, n17111, n17112, n17114, n17115, n17116,
         n17117, n17118, n17119, n17120, n17122, n17124, n17125, n17126,
         n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134,
         n17135, n17137, n17138, n17139, n17140, n17141, n17143, n17144,
         n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154,
         n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162,
         n17163, n17164, n17165, n17166, n17168, n17170, n17171, n17172,
         n17173, n17174, n17175, n17176, n17177, n17180, n17181, n17182,
         n17183, n17184, n17185, n17186, n17189, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17215, n17216, n17217, n17218,
         n17219, n17220, n17221, n17223, n17224, n17225, n17226, n17227,
         n17228, n17230, n17231, n17232, n17233, n17234, n17235, n17236,
         n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244,
         n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252,
         n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261,
         n17263, n17264, n17265, n17266, n17267, n17268, n17270, n17271,
         n17272, n17273, n17274, n17275, n17277, n17278, n17279, n17280,
         n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,
         n17289, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17311, n17312, n17315, n17316, n17317, n17318,
         n17319, n17320, n17321, n17322, n17324, n17326, n17328, n17329,
         n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340,
         n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348,
         n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356,
         n17357, n17359, n17360, n17361, n17362, n17363, n17364, n17365,
         n17366, n17367, n17368, n17370, n17371, n17372, n17373, n17374,
         n17375, n17376, n17377, n17378, n17379, n17380, n17382, n17383,
         n17384, n17385, n17387, n17389, n17390, n17391, n17392, n17394,
         n17395, n17396, n17397, n17398, n17400, n17401, n17402, n17403,
         n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411,
         n17412, n17413, n17414, n17415, n17416, n17418, n17419, n17420,
         n17422, n17423, n17425, n17426, n17427, n17428, n17429, n17430,
         n17431, n17432, n17433, n17434, n17436, n17437, n17438, n17439,
         n17441, n17442, n17444, n17446, n17447, n17448, n17450, n17451,
         n17452, n17453, n17455, n17457, n17458, n17459, n17460, n17462,
         n17463, n17464, n17466, n17467, n17468, n17470, n17471, n17472,
         n17473, n17474, n17476, n17477, n17478, n17479, n17481, n17482,
         n17483, n17484, n17486, n17487, n17488, n17489, n17490, n17491,
         n17492, n17494, n17495, n17496, n17497, n17498, n17499, n17500,
         n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508,
         n17509, n17510, n17511, n17512, n17513, n17514, n17516, n17517,
         n17518, n17520, n17521, n17522, n17523, n17524, n17525, n17526,
         n17527, n17528, n17529, n17530, n17532, n17533, n17536, n17537,
         n17538, n17540, n17542, n17543, n17544, n17545, n17546, n17547,
         n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555,
         n17556, n17557, n17558, n17559, n17560, n17562, n17563, n17564,
         n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574,
         n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17583,
         n17584, n17586, n17589, n17590, n17591, n17592, n17594, n17595,
         n17596, n17597, n17598, n17599, n17601, n17602, n17603, n17604,
         n17605, n17606, n17607, n17608, n17610, n17611, n17612, n17613,
         n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
         n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630,
         n17631, n17632, n17633, n17634, n17635, n17637, n17638, n17639,
         n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647,
         n17648, n17649, n17650, n17651, n17652, n17654, n17655, n17656,
         n17657, n17660, n17661, n17663, n17664, n17665, n17666, n17667,
         n17668, n17670, n17671, n17672, n17673, n17675, n17677, n17678,
         n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686,
         n17687, n17688, n17689, n17691, n17692, n17693, n17697, n17700,
         n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708,
         n17710, n17711, n17712, n17713, n17714, n17715, n17717, n17718,
         n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726,
         n17727, n17728, n17729, n17731, n17733, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17743, n17744, n17745, n17746,
         n17747, n17750, n17751, n17752, n17753, n17754, n17755, n17756,
         n17757, n17758, n17759, n17761, n17762, n17763, n17764, n17765,
         n17766, n17768, n17769, n17770, n17771, n17772, n17773, n17774,
         n17775, n17776, n17777, n17778, n17780, n17781, n17783, n17784,
         n17785, n17786, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17798, n17799, n17800, n17801, n17802,
         n17803, n17805, n17806, n17808, n17809, n17810, n17813, n17815,
         n17816, n17817, n17818, n17821, n17824, n17827, n17828, n17829,
         n17831, n17833, n17834, n17835, n17836, n17837, n17838, n17840,
         n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848,
         n17849, n17850, n17851, n17852, n17853, n17855, n17856, n17857,
         n17859, n17860, n17861, n17862, n17863, n17865, n17866, n17867,
         n17868, n17869, n17870, n17872, n17873, n17874, n17875, n17876,
         n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885,
         n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893,
         n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902,
         n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17911,
         n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919,
         n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17928,
         n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,
         n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944,
         n17945, n17947, n17948, n17949, n17950, n17951, n17952, n17954,
         n17955, n17957, n17958, n17959, n17960, n17961, n17962, n17963,
         n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971,
         n17972, n17975, n17977, n17978, n17979, n17980, n17981, n17982,
         n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17991,
         n17992, n17993, n17994, n17996, n17997, n17998, n17999, n18000,
         n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008,
         n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016,
         n18018, n18019, n18020, n18021, n18022, n18023, n18027, n18028,
         n18029, n18031, n18032, n18033, n18034, n18035, n18036, n18037,
         n18038, n18039, n18041, n18042, n18043, n18045, n18046, n18047,
         n18048, n18049, n18050, n18051, n18053, n18054, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18065, n18066,
         n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18075,
         n18076, n18077, n18078, n18079, n18080, n18081, n18083, n18084,
         n18085, n18086, n18087, n18088, n18089, n18091, n18092, n18093,
         n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102,
         n18103, n18104, n18106, n18107, n18108, n18109, n18111, n18112,
         n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120,
         n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,
         n18129, n18130, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18142, n18143, n18144, n18145, n18146, n18147,
         n18148, n18149, n18150, n18151, n18153, n18154, n18155, n18156,
         n18158, n18159, n18160, n18162, n18167, n18169, n18170, n18172,
         n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180,
         n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188,
         n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196,
         n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205,
         n18206, n18207, n18208, n18209, n18211, n18213, n18214, n18215,
         n18216, n18218, n18219, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18246, n18247, n18248, n18249, n18250,
         n18251, n18252, n18254, n18255, n18256, n18257, n18258, n18259,
         n18260, n18261, n18262, n18263, n18264, n18265, n18268, n18269,
         n18270, n18271, n18273, n18276, n18277, n18278, n18281, n18282,
         n18283, n18284, n18285, n18286, n18287, n18288, n18290, n18291,
         n18292, n18293, n18294, n18295, n18296, n18297, n18299, n18300,
         n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308,
         n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317,
         n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325,
         n18326, n18327, n18328, n18330, n18331, n18333, n18334, n18335,
         n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343,
         n18344, n18348, n18349, n18351, n18352, n18354, n18355, n18356,
         n18357, n18358, n18361, n18362, n18363, n18364, n18365, n18366,
         n18368, n18370, n18371, n18372, n18373, n18374, n18375, n18376,
         n18377, n18379, n18380, n18381, n18382, n18383, n18385, n18386,
         n18387, n18388, n18389, n18390, n18391, n18393, n18394, n18395,
         n18396, n18397, n18398, n18399, n18401, n18402, n18405, n18406,
         n18407, n18408, n18410, n18411, n18413, n18414, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18430, n18431, n18432, n18433, n18434,
         n18435, n18440, n18441, n18442, n18443, n18444, n18446, n18447,
         n18448, n18450, n18451, n18452, n18453, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18505, n18506,
         n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514,
         n18515, n18516, n18518, n18519, n18520, n18521, n18522, n18523,
         n18524, n18525, n18526, n18528, n18529, n18530, n18531, n18532,
         n18533, n18534, n18536, n18537, n18538, n18539, n18540, n18541,
         n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549,
         n18550, n18551, n18553, n18554, n18555, n18557, n18558, n18559,
         n18560, n18561, n18562, n18564, n18565, n18566, n18568, n18569,
         n18570, n18571, n18573, n18574, n18575, n18576, n18578, n18579,
         n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18589,
         n18590, n18592, n18593, n18594, n18595, n18596, n18597, n18598,
         n18599, n18600, n18601, n18602, n18603, n18605, n18606, n18607,
         n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615,
         n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623,
         n18624, n18625, n18629, n18630, n18631, n18632, n18633, n18634,
         n18635, n18637, n18638, n18639, n18640, n18641, n18642, n18644,
         n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652,
         n18655, n18656, n18658, n18659, n18660, n18661, n18662, n18664,
         n18665, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18685, n18686, n18687, n18688, n18690, n18691,
         n18693, n18695, n18696, n18698, n18699, n18700, n18701, n18702,
         n18704, n18705, n18706, n18707, n18708, n18709, n18711, n18712,
         n18713, n18714, n18715, n18716, n18717, n18720, n18721, n18722,
         n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730,
         n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
         n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747,
         n18748, n18750, n18751, n18752, n18753, n18754, n18755, n18756,
         n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764,
         n18765, n18766, n18767, n18769, n18770, n18771, n18773, n18774,
         n18775, n18776, n18777, n18779, n18780, n18781, n18782, n18783,
         n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18792,
         n18793, n18794, n18796, n18797, n18799, n18800, n18801, n18802,
         n18803, n18804, n18806, n18807, n18808, n18809, n18810, n18811,
         n18812, n18813, n18814, n18815, n18816, n18817, n18819, n18820,
         n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18829,
         n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837,
         n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18846,
         n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854,
         n18855, n18856, n18857, n18858, n18859, n18861, n18862, n18863,
         n18864, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882,
         n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890,
         n18891, n18892, n18895, n18896, n18897, n18898, n18899, n18900,
         n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908,
         n18909, n18910, n18911, n18914, n18915, n18916, n18917, n18918,
         n18919, n18920, n18922, n18923, n18924, n18925, n18926, n18927,
         n18929, n18930, n18931, n18932, n18933, n18935, n18936, n18937,
         n18938, n18939, n18941, n18943, n18944, n18945, n18946, n18947,
         n18950, n18951, n18954, n18955, n18956, n18957, n18958, n18959,
         n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967,
         n18968, n18969, n18971, n18972, n18973, n18974, n18975, n18976,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18986,
         n18987, n18989, n18990, n18991, n18992, n18993, n18995, n18996,
         n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004,
         n19005, n19006, n19007, n19008, n19009, n19010, n19012, n19013,
         n19015, n19017, n19018, n19019, n19020, n19021, n19022, n19023,
         n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031,
         n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039,
         n19040, n19041, n19042, n19043, n19044, n19045, n19047, n19048,
         n19049, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19062, n19064, n19065, n19066, n19067,
         n19068, n19069, n19070, n19071, n19072, n19073, n19075, n19076,
         n19077, n19078, n19079, n19080, n19081, n19083, n19085, n19087,
         n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095,
         n19096, n19098, n19100, n19101, n19102, n19103, n19105, n19106,
         n19107, n19108, n19109, n19110, n19112, n19113, n19114, n19118,
         n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126,
         n19127, n19129, n19130, n19131, n19132, n19133, n19134, n19137,
         n19138, n19139, n19140, n19142, n19144, n19145, n19146, n19147,
         n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155,
         n19156, n19158, n19159, n19160, n19161, n19163, n19165, n19167,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19181, n19183, n19184, n19185, n19186, n19187,
         n19188, n19189, n19190, n19191, n19192, n19193, n19195, n19196,
         n19197, n19198, n19200, n19201, n19202, n19203, n19204, n19206,
         n19207, n19208, n19209, n19210, n19212, n19214, n19215, n19216,
         n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224,
         n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232,
         n19233, n19237, n19238, n19240, n19241, n19242, n19243, n19245,
         n19246, n19248, n19249, n19250, n19252, n19253, n19254, n19255,
         n19256, n19258, n19260, n19261, n19262, n19263, n19265, n19266,
         n19268, n19269, n19270, n19271, n19273, n19274, n19275, n19276,
         n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19285,
         n19287, n19289, n19290, n19291, n19292, n19294, n19295, n19296,
         n19297, n19299, n19300, n19301, n19302, n19303, n19305, n19306,
         n19307, n19309, n19311, n19312, n19313, n19314, n19316, n19317,
         n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326,
         n19328, n19329, n19330, n19331, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19346,
         n19347, n19348, n19349, n19351, n19352, n19353, n19354, n19356,
         n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364,
         n19365, n19367, n19368, n19369, n19371, n19372, n19373, n19374,
         n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19383,
         n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19392,
         n19393, n19395, n19396, n19397, n19400, n19401, n19402, n19403,
         n19404, n19407, n19409, n19410, n19411, n19412, n19413, n19416,
         n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19426,
         n19428, n19430, n19431, n19432, n19433, n19434, n19435, n19437,
         n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445,
         n19446, n19448, n19449, n19450, n19451, n19452, n19453, n19454,
         n19455, n19456, n19457, n19458, n19460, n19461, n19462, n19464,
         n19465, n19466, n19467, n19471, n19473, n19474, n19475, n19476,
         n19477, n19478, n19479, n19481, n19482, n19483, n19484, n19485,
         n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493,
         n19494, n19496, n19497, n19499, n19500, n19501, n19502, n19503,
         n19504, n19505, n19507, n19509, n19510, n19511, n19512, n19514,
         n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522,
         n19523, n19524, n19525, n19526, n19527, n19529, n19530, n19531,
         n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539,
         n19540, n19541, n19543, n19544, n19545, n19546, n19547, n19548,
         n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556,
         n19557, n19558, n19559, n19560, n19562, n19563, n19564, n19565,
         n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573,
         n19574, n19575, n19577, n19578, n19581, n19584, n19587, n19588,
         n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19597,
         n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605,
         n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613,
         n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621,
         n19622, n19624, n19625, n19626, n19627, n19628, n19629, n19630,
         n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638,
         n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646,
         n19647, n19648, n19649, n19652, n19653, n19654, n19656, n19658,
         n19661, n19662, n19663, n19664, n19665, n19666, n19670, n19671,
         n19672, n19674, n19675, n19676, n19677, n19678, n19679, n19680,
         n19681, n19682, n19683, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706,
         n19707, n19708, n19709, n19711, n19712, n19713, n19714, n19715,
         n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723,
         n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19735,
         n19736, n19737, n19738, n19739, n19740, n19742, n19743, n19746,
         n19747, n19748, n19750, n19751, n19752, n19753, n19754, n19755,
         n19756, n19757, n19758, n19759, n19760, n19761, n19763, n19764,
         n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772,
         n19773, n19774, n19775, n19777, n19778, n19780, n19781, n19782,
         n19783, n19785, n19786, n19787, n19788, n19789, n19790, n19791,
         n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19800,
         n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808,
         n19809, n19810, n19811, n19813, n19814, n19816, n19817, n19818,
         n19819, n19821, n19822, n19823, n19824, n19825, n19826, n19827,
         n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835,
         n19836, n19838, n19841, n19843, n19844, n19845, n19847, n19848,
         n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856,
         n19857, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19870, n19871, n19872, n19873, n19874,
         n19876, n19878, n19879, n19882, n19883, n19884, n19885, n19886,
         n19887, n19888, n19889, n19890, n19891, n19893, n19894, n19896,
         n19897, n19899, n19900, n19902, n19903, n19904, n19905, n19907,
         n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915,
         n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19924,
         n19925, n19926, n19927, n19928, n19929, n19931, n19932, n19933,
         n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942,
         n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950,
         n19951, n19952, n19953, n19954, n19955, n19956, n19958, n19959,
         n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967,
         n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975,
         n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983,
         n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991,
         n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999,
         n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007,
         n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015,
         n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023,
         n20024, n20025, n20026, n20028, n20029, n20031, n20032, n20034,
         n20037, n20038, n20039, n20040, n20041, n20042, n20044, n20045,
         n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053,
         n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061,
         n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069,
         n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077,
         n20078, n20079, n20080, n20081, n20083, n20084, n20085, n20086,
         n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094,
         n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102,
         n20103, n20105, n20106, n20107, n20108, n20109, n20110, n20111,
         n20112, n20113, n20114, n20115, n20116, n20118, n20121, n20122,
         n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130,
         n20131, n20132, n20134, n20136, n20137, n20138, n20139, n20140,
         n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148,
         n20151, n20152, n20153, n20155, n20156, n20157, n20158, n20159,
         n20160, n20161, n20162, n20163, n20165, n20166, n20167, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20190, n20191, n20193, n20194, n20195,
         n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205,
         n20206, n20207, n20208, n20209, n20211, n20212, n20213, n20214,
         n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222,
         n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230,
         n20232, n20234, n20235, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20248, n20249, n20250,
         n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258,
         n20259, n20260, n20261, n20262, n20263, n20264, n20266, n20268,
         n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276,
         n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284,
         n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292,
         n20293, n20294, n20297, n20298, n20299, n20300, n20301, n20302,
         n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310,
         n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318,
         n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326,
         n20328, n20329, n20330, n20331, n20332, n20334, n20335, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20347, n20348, n20349, n20351, n20352, n20353, n20354, n20355,
         n20356, n20357, n20360, n20361, n20362, n20363, n20364, n20365,
         n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374,
         n20375, n20376, n20378, n20380, n20381, n20382, n20383, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20399, n20400, n20401, n20402,
         n20403, n20404, n20406, n20407, n20408, n20409, n20410, n20411,
         n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419,
         n20421, n20423, n20425, n20426, n20427, n20428, n20429, n20430,
         n20431, n20432, n20433, n20435, n20436, n20437, n20438, n20439,
         n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448,
         n20449, n20451, n20452, n20455, n20456, n20457, n20458, n20460,
         n20461, n20462, n20464, n20466, n20468, n20469, n20470, n20471,
         n20472, n20473, n20474, n20476, n20477, n20478, n20479, n20480,
         n20481, n20484, n20485, n20486, n20487, n20488, n20489, n20491,
         n20492, n20493, n20495, n20496, n20497, n20498, n20501, n20502,
         n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511,
         n20512, n20513, n20514, n20516, n20517, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20533, n20534, n20535, n20538, n20539, n20540,
         n20541, n20544, n20545, n20546, n20547, n20548, n20549, n20550,
         n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20559,
         n20560, n20561, n20562, n20563, n20565, n20566, n20567, n20568,
         n20569, n20570, n20571, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20584, n20585, n20586,
         n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594,
         n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602,
         n20603, n20605, n20606, n20607, n20608, n20609, n20610, n20611,
         n20613, n20614, n20615, n20616, n20617, n20619, n20620, n20621,
         n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629,
         n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637,
         n20638, n20639, n20642, n20643, n20645, n20646, n20648, n20649,
         n20650, n20652, n20653, n20654, n20655, n20656, n20657, n20658,
         n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666,
         n20667, n20668, n20669, n20670, n20671, n20673, n20674, n20675,
         n20676, n20678, n20679, n20680, n20682, n20683, n20684, n20685,
         n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693,
         n20694, n20695, n20696, n20699, n20700, n20701, n20703, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20719, n20720, n20721, n20722,
         n20723, n20724, n20725, n20726, n20728, n20730, n20731, n20733,
         n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741,
         n20742, n20743, n20745, n20747, n20749, n20750, n20751, n20752,
         n20753, n20754, n20755, n20756, n20757, n20758, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20769, n20770,
         n20771, n20772, n20773, n20774, n20776, n20777, n20778, n20779,
         n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787,
         n20788, n20789, n20790, n20791, n20792, n20793, n20796, n20797,
         n20798, n20799, n20800, n20802, n20803, n20806, n20807, n20808,
         n20809, n20810, n20811, n20812, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20826,
         n20828, n20830, n20831, n20832, n20834, n20835, n20836, n20837,
         n20838, n20839, n20841, n20842, n20844, n20845, n20846, n20847,
         n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855,
         n20856, n20857, n20859, n20860, n20861, n20862, n20863, n20864,
         n20865, n20867, n20869, n20870, n20871, n20872, n20874, n20875,
         n20876, n20878, n20879, n20881, n20882, n20883, n20886, n20887,
         n20888, n20889, n20891, n20892, n20893, n20894, n20895, n20896,
         n20897, n20898, n20899, n20900, n20901, n20902, n20904, n20905,
         n20907, n20908, n20909, n20911, n20912, n20913, n20915, n20916,
         n20917, n20918, n20919, n20921, n20922, n20923, n20925, n20926,
         n20927, n20929, n20930, n20931, n20932, n20933, n20934, n20935,
         n20936, n20937, n20938, n20940, n20941, n20942, n20944, n20945,
         n20946, n20947, n20948, n20950, n20951, n20953, n20954, n20955,
         n20956, n20957, n20958, n20960, n20962, n20963, n20964, n20965,
         n20966, n20968, n20969, n20970, n20971, n20972, n20974, n20975,
         n20978, n20979, n20980, n20982, n20983, n20984, n20985, n20987,
         n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20996,
         n20998, n20999, n21000, n21001, n21005, n21006, n21008, n21009,
         n21010, n21011, n21014, n21016, n21017, n21018, n21019, n21020,
         n21021, n21022, n21023, n21024, n21025, n21027, n21028, n21029,
         n21030, n21032, n21033, n21034, n21035, n21036, n21037, n21039,
         n21040, n21041, n21042, n21044, n21046, n21050, n21051, n21052,
         n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062,
         n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070,
         n21071, n21073, n21074, n21079, n21081, n21082, n21083, n21084,
         n21085, n21086, n21087, n21088, n21090, n21092, n21094, n21095,
         n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21104,
         n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112,
         n21113, n21114, n21115, n21117, n21118, n21119, n21120, n21121,
         n21122, n21124, n21125, n21126, n21127, n21128, n21129, n21130,
         n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138,
         n21139, n21140, n21141, n21142, n21143, n21146, n21147, n21148,
         n21150, n21151, n21152, n21153, n21154, n21156, n21157, n21158,
         n21159, n21160, n21161, n21162, n21163, n21165, n21166, n21167,
         n21168, n21169, n21170, n21171, n21172, n21173, n21176, n21177,
         n21178, n21179, n21181, n21183, n21184, n21185, n21186, n21187,
         n21188, n21189, n21190, n21191, n21193, n21194, n21196, n21198,
         n21199, n21200, n21203, n21204, n21205, n21206, n21207, n21209,
         n21210, n21211, n21212, n21214, n21215, n21216, n21217, n21218,
         n21219, n21220, n21222, n21223, n21225, n21226, n21227, n21228,
         n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236,
         n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244,
         n21245, n21246, n21248, n21249, n21251, n21252, n21253, n21254,
         n21255, n21257, n21258, n21259, n21260, n21261, n21262, n21263,
         n21264, n21265, n21266, n21268, n21269, n21270, n21271, n21272,
         n21273, n21274, n21275, n21276, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21303, n21304, n21305, n21307,
         n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315,
         n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21324,
         n21325, n21326, n21328, n21329, n21330, n21331, n21332, n21333,
         n21334, n21335, n21336, n21339, n21340, n21341, n21342, n21343,
         n21344, n21345, n21346, n21347, n21348, n21349, n21351, n21352,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21379, n21380, n21381, n21382, n21383, n21384, n21385, n21386,
         n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394,
         n21395, n21397, n21398, n21399, n21400, n21401, n21402, n21403,
         n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411,
         n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419,
         n21420, n21421, n21422, n21424, n21425, n21426, n21427, n21428,
         n21429, n21430, n21431, n21432, n21433, n21434, n21436, n21437,
         n21438, n21439, n21440, n21441, n21442, n21443, n21445, n21446,
         n21447, n21448, n21449, n21450, n21451, n21452, n21453, n21454,
         n21455, n21456, n21457, n21459, n21460, n21461, n21462, n21463,
         n21464, n21465, n21466, n21467, n21468, n21469, n21470, n21471,
         n21473, n21474, n21475, n21476, n21477, n21478, n21479, n21480,
         n21481, n21482, n21483, n21484, n21485, n21486, n21487, n21488,
         n21489, n21490, n21491, n21492, n21493, n21494, n21495, n21496,
         n21497, n21498, n21499, n21501, n21502, n21503, n21504, n21506,
         n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21516,
         n21517, n21518, n21519, n21520, n21521, n21522, n21525, n21526,
         n21527, n21528, n21529, n21530, n21531, n21532, n21535, n21536,
         n21537, n21538, n21541, n21542, n21543, n21544, n21545, n21546,
         n21547, n21548, n21549, n21550, n21551, n21552, n21555, n21556,
         n21557, n21558, n21559, n21560, n21561, n21562, n21563, n21564,
         n21565, n21566, n21567, n21568, n21569, n21570, n21572, n21573,
         n21574, n21575, n21576, n21577, n21578, n21579, n21580, n21581,
         n21582, n21584, n21585, n21586, n21588, n21589, n21590, n21591,
         n21592, n21593, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21604, n21605, n21606, n21607, n21608, n21609, n21610,
         n21611, n21612, n21613, n21614, n21615, n21616, n21617, n21620,
         n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628,
         n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21638,
         n21639, n21640, n21641, n21642, n21643, n21644, n21645, n21649,
         n21650, n21651, n21653, n21655, n21656, n21657, n21659, n21660,
         n21661, n21662, n21663, n21664, n21665, n21666, n21667, n21668,
         n21669, n21671, n21672, n21673, n21674, n21675, n21676, n21677,
         n21678, n21679, n21680, n21681, n21682, n21683, n21684, n21685,
         n21686, n21687, n21688, n21689, n21690, n21691, n21692, n21693,
         n21694, n21695, n21696, n21697, n21699, n21700, n21701, n21702,
         n21703, n21704, n21705, n21706, n21707, n21708, n21709, n21710,
         n21711, n21712, n21713, n21714, n21715, n21716, n21717, n21718,
         n21719, n21720, n21721, n21722, n21723, n21724, n21725, n21726,
         n21727, n21728, n21729, n21730, n21731, n21732, n21733, n21734,
         n21735, n21736, n21737, n21738, n21740, n21741, n21742, n21743,
         n21744, n21745, n21746, n21747, n21748, n21749, n21750, n21751,
         n21752, n21753, n21754, n21755, n21756, n21757, n21758, n21759,
         n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767,
         n21768, n21769, n21771, n21773, n21774, n21775, n21776, n21777,
         n21778, n21779, n21780, n21781, n21784, n21785, n21786, n21787,
         n21788, n21789, n21790, n21791, n21792, n21793, n21794, n21795,
         n21796, n21798, n21799, n21800, n21801, n21802, n21803, n21804,
         n21805, n21806, n21807, n21808, n21809, n21810, n21811, n21812,
         n21813, n21814, n21816, n21817, n21819, n21820, n21821, n21822,
         n21823, n21824, n21825, n21826, n21828, n21829, n21830, n21831,
         n21832, n21833, n21834, n21835, n21837, n21838, n21839, n21840,
         n21841, n21842, n21843, n21844, n21847, n21848, n21849, n21850,
         n21851, n21852, n21854, n21855, n21856, n21857, n21859, n21860,
         n21861, n21862, n21863, n21864, n21865, n21866, n21867, n21868,
         n21869, n21870, n21875, n21876, n21877, n21878, n21879, n21880,
         n21881, n21883, n21884, n21885, n21886, n21887, n21888, n21890,
         n21891, n21892, n21893, n21894, n21895, n21896, n21897, n21899,
         n21900, n21903, n21904, n21905, n21906, n21908, n21909, n21910,
         n21911, n21912, n21913, n21914, n21915, n21916, n21917, n21918,
         n21919, n21920, n21921, n21922, n21923, n21924, n21925, n21927,
         n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935,
         n21937, n21938, n21939, n21940, n21941, n21942, n21943, n21944,
         n21945, n21946, n21947, n21948, n21949, n21950, n21951, n21952,
         n21953, n21954, n21955, n21956, n21957, n21958, n21959, n21960,
         n21961, n21962, n21963, n21964, n21965, n21966, n21967, n21968,
         n21969, n21970, n21971, n21972, n21973, n21974, n21975, n21976,
         n21977, n21978, n21980, n21982, n21983, n21984, n21985, n21986,
         n21987, n21988, n21989, n21990, n21991, n21992, n21993, n21994,
         n21996, n21997, n21998, n21999, n22000, n22002, n22003, n22004,
         n22005, n22006, n22007, n22008, n22009, n22010, n22011, n22012,
         n22014, n22015, n22016, n22017, n22018, n22019, n22020, n22021,
         n22022, n22023, n22024, n22025, n22026, n22027, n22029, n22030,
         n22032, n22033, n22034, n22035, n22036, n22038, n22039, n22040,
         n22041, n22042, n22043, n22044, n22045, n22047, n22048, n22050,
         n22051, n22053, n22056, n22057, n22058, n22059, n22060, n22061,
         n22062, n22063, n22064, n22065, n22066, n22067, n22068, n22069,
         n22070, n22071, n22072, n22073, n22074, n22078, n22079, n22080,
         n22081, n22082, n22083, n22084, n22085, n22086, n22087, n22088,
         n22089, n22091, n22092, n22093, n22094, n22095, n22097, n22098,
         n22099, n22100, n22101, n22102, n22103, n22104, n22105, n22106,
         n22107, n22108, n22109, n22110, n22111, n22112, n22113, n22114,
         n22115, n22116, n22117, n22118, n22119, n22120, n22121, n22122,
         n22123, n22124, n22126, n22127, n22128, n22129, n22130, n22131,
         n22139, n22141, n22142, n22143, n22144, n22145, n22146, n22148,
         n22150, n22152, n22153, n22154, n22155, n22156, n22157, n22158,
         n22159, n22160, n22161, n22162, n22163, n22164, n22166, n22168,
         n22169, n22170, n22171, n22172, n22173, n22174, n22176, n22177,
         n22180, n22181, n22182, n22184, n22185, n22186, n22187, n22188,
         n22189, n22190, n22191, n22195, n22197, n22198, n22199, n22200,
         n22201, n22202, n22203, n22204, n22205, n22206, n22207, n22208,
         n22209, n22210, n22211, n22212, n22213, n22214, n22215, n22217,
         n22219, n22220, n22221, n22222, n22223, n22224, n22225, n22226,
         n22227, n22228, n22229, n22230, n22231, n22232, n22233, n22234,
         n22235, n22236, n22237, n22239, n22241, n22242, n22243, n22244,
         n22246, n22247, n22248, n22249, n22250, n22252, n22253, n22254,
         n22255, n22256, n22257, n22258, n22259, n22260, n22262, n22263,
         n22264, n22265, n22266, n22267, n22268, n22269, n22271, n22273,
         n22274, n22276, n22277, n22278, n22279, n22280, n22281, n22282,
         n22283, n22284, n22285, n22286, n22287, n22288, n22289, n22290,
         n22291, n22292, n22293, n22294, n22295, n22296, n22297, n22299,
         n22301, n22302, n22303, n22304, n22305, n22307, n22308, n22310,
         n22311, n22312, n22313, n22314, n22315, n22316, n22317, n22318,
         n22319, n22320, n22321, n22322, n22323, n22325, n22326, n22329,
         n22330, n22331, n22332, n22333, n22334, n22336, n22337, n22338,
         n22339, n22340, n22342, n22343, n22344, n22345, n22346, n22348,
         n22349, n22350, n22351, n22352, n22353, n22355, n22357, n22359,
         n22360, n22361, n22362, n22363, n22364, n22365, n22367, n22370,
         n22372, n22373, n22374, n22376, n22377, n22378, n22379, n22380,
         n22381, n22382, n22383, n22384, n22385, n22386, n22387, n22388,
         n22389, n22390, n22391, n22394, n22395, n22396, n22397, n22398,
         n22401, n22402, n22404, n22406, n22408, n22409, n22410, n22411,
         n22412, n22413, n22414, n22415, n22416, n22417, n22418, n22419,
         n22421, n22422, n22423, n22424, n22426, n22427, n22428, n22429,
         n22430, n22431, n22432, n22433, n22434, n22435, n22436, n22439,
         n22440, n22442, n22443, n22444, n22446, n22447, n22448, n22450,
         n22451, n22452, n22453, n22454, n22455, n22456, n22457, n22458,
         n22459, n22461, n22462, n22463, n22464, n22466, n22468, n22469,
         n22470, n22471, n22472, n22473, n22474, n22476, n22477, n22478,
         n22479, n22480, n22481, n22482, n22483, n22484, n22485, n22486,
         n22487, n22488, n22489, n22491, n22494, n22495, n22496, n22497,
         n22498, n22499, n22500, n22502, n22503, n22504, n22505, n22506,
         n22508, n22509, n22510, n22512, n22513, n22514, n22515, n22516,
         n22518, n22519, n22520, n22521, n22523, n22524, n22525, n22526,
         n22527, n22528, n22530, n22531, n22533, n22534, n22535, n22536,
         n22537, n22538, n22539, n22540, n22541, n22542, n22544, n22545,
         n22546, n22547, n22549, n22550, n22551, n22552, n22553, n22554,
         n22555, n22556, n22557, n22558, n22559, n22560, n22561, n22564,
         n22565, n22566, n22569, n22570, n22571, n22572, n22573, n22574,
         n22576, n22577, n22578, n22579, n22580, n22581, n22583, n22584,
         n22586, n22587, n22588, n22589, n22591, n22592, n22593, n22594,
         n22595, n22596, n22597, n22598, n22599, n22601, n22602, n22603,
         n22604, n22605, n22606, n22607, n22608, n22609, n22613, n22614,
         n22617, n22618, n22619, n22620, n22621, n22622, n22625, n22626,
         n22627, n22628, n22629, n22630, n22632, n22633, n22635, n22637,
         n22638, n22639, n22640, n22641, n22642, n22643, n22645, n22646,
         n22647, n22648, n22650, n22651, n22652, n22653, n22654, n22656,
         n22657, n22658, n22659, n22660, n22661, n22662, n22664, n22666,
         n22667, n22668, n22669, n22670, n22671, n22673, n22674, n22675,
         n22676, n22677, n22678, n22679, n22680, n22681, n22682, n22683,
         n22684, n22689, n22690, n22691, n22693, n22694, n22695, n22696,
         n22697, n22698, n22699, n22700, n22701, n22702, n22703, n22704,
         n22705, n22706, n22707, n22708, n22709, n22710, n22711, n22712,
         n22713, n22714, n22715, n22716, n22717, n22718, n22719, n22720,
         n22721, n22723, n22724, n22725, n22726, n22727, n22728, n22731,
         n22732, n22733, n22734, n22735, n22736, n22737, n22738, n22739,
         n22741, n22742, n22743, n22744, n22745, n22746, n22747, n22748,
         n22749, n22750, n22751, n22752, n22753, n22755, n22756, n22757,
         n22758, n22759, n22760, n22761, n22762, n22763, n22764, n22765,
         n22767, n22768, n22769, n22772, n22773, n22775, n22776, n22777,
         n22778, n22779, n22780, n22781, n22782, n22783, n22785, n22786,
         n22787, n22788, n22790, n22792, n22794, n22795, n22796, n22797,
         n22798, n22799, n22800, n22801, n22802, n22803, n22804, n22805,
         n22806, n22807, n22809, n22810, n22811, n22812, n22813, n22814,
         n22815, n22817, n22818, n22819, n22820, n22821, n22822, n22823,
         n22824, n22825, n22831, n22832, n22835, n22836, n22837, n22838,
         n22839, n22840, n22841, n22842, n22844, n22845, n22846, n22847,
         n22848, n22850, n22851, n22852, n22853, n22855, n22856, n22857,
         n22858, n22859, n22860, n22861, n22863, n22864, n22865, n22866,
         n22867, n22868, n22869, n22870, n22871, n22872, n22873, n22874,
         n22875, n22876, n22877, n22878, n22879, n22880, n22881, n22882,
         n22883, n22884, n22885, n22886, n22887, n22889, n22890, n22891,
         n22892, n22893, n22894, n22895, n22896, n22897, n22898, n22899,
         n22900, n22902, n22903, n22905, n22907, n22908, n22909, n22910,
         n22911, n22912, n22913, n22915, n22916, n22918, n22919, n22921,
         n22922, n22923, n22925, n22926, n22927, n22928, n22929, n22930,
         n22931, n22932, n22933, n22934, n22935, n22936, n22937, n22939,
         n22940, n22941, n22942, n22943, n22944, n22945, n22947, n22948,
         n22949, n22950, n22951, n22952, n22953, n22954, n22956, n22957,
         n22958, n22959, n22961, n22962, n22963, n22964, n22965, n22966,
         n22967, n22968, n22969, n22971, n22972, n22973, n22975, n22976,
         n22977, n22978, n22979, n22980, n22981, n22983, n22985, n22986,
         n22988, n22989, n22990, n22991, n22992, n22993, n22994, n22995,
         n22996, n22997, n22998, n22999, n23000, n23002, n23003, n23004,
         n23005, n23006, n23007, n23008, n23013, n23014, n23015, n23016,
         n23017, n23018, n23019, n23020, n23021, n23022, n23024, n23025,
         n23027, n23028, n23030, n23032, n23033, n23035, n23036, n23037,
         n23039, n23040, n23041, n23042, n23044, n23046, n23047, n23048,
         n23049, n23050, n23051, n23052, n23053, n23054, n23055, n23056,
         n23058, n23059, n23061, n23062, n23063, n23064, n23065, n23067,
         n23068, n23069, n23070, n23071, n23072, n23073, n23074, n23076,
         n23077, n23078, n23080, n23083, n23084, n23085, n23086, n23087,
         n23088, n23089, n23090, n23092, n23093, n23094, n23095, n23096,
         n23097, n23098, n23099, n23101, n23102, n23104, n23106, n23107,
         n23108, n23110, n23111, n23112, n23113, n23114, n23115, n23116,
         n23117, n23118, n23119, n23120, n23121, n23122, n23123, n23124,
         n23125, n23126, n23127, n23128, n23129, n23130, n23131, n23132,
         n23133, n23134, n23135, n23136, n23137, n23138, n23139, n23140,
         n23141, n23143, n23144, n23145, n23146, n23147, n23148, n23149,
         n23150, n23151, n23152, n23153, n23154, n23155, n23156, n23157,
         n23158, n23159, n23160, n23162, n23163, n23164, n23165, n23166,
         n23167, n23168, n23169, n23170, n23173, n23174, n23175, n23176,
         n23177, n23178, n23179, n23180, n23181, n23182, n23184, n23185,
         n23186, n23187, n23188, n23191, n23192, n23193, n23194, n23195,
         n23196, n23197, n23199, n23200, n23204, n23206, n23207, n23208,
         n23209, n23210, n23211, n23212, n23213, n23215, n23216, n23217,
         n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225,
         n23226, n23227, n23229, n23230, n23231, n23232, n23236, n23237,
         n23238, n23239, n23241, n23242, n23243, n23245, n23246, n23247,
         n23248, n23249, n23250, n23251, n23252, n23253, n23254, n23256,
         n23257, n23258, n23259, n23260, n23261, n23263, n23264, n23266,
         n23267, n23269, n23270, n23271, n23272, n23273, n23274, n23275,
         n23276, n23277, n23278, n23279, n23280, n23281, n23282, n23283,
         n23284, n23285, n23286, n23287, n23288, n23289, n23290, n23292,
         n23294, n23295, n23297, n23298, n23299, n23300, n23301, n23302,
         n23303, n23305, n23306, n23307, n23309, n23311, n23312, n23313,
         n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23323,
         n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331,
         n23332, n23333, n23334, n23335, n23337, n23339, n23340, n23341,
         n23342, n23343, n23344, n23345, n23346, n23347, n23348, n23349,
         n23350, n23351, n23352, n23353, n23354, n23355, n23356, n23357,
         n23360, n23361, n23362, n23363, n23364, n23365, n23366, n23367,
         n23368, n23369, n23370, n23371, n23372, n23373, n23375, n23376,
         n23377, n23380, n23381, n23383, n23385, n23386, n23387, n23388,
         n23389, n23390, n23394, n23395, n23396, n23397, n23398, n23399,
         n23400, n23401, n23402, n23403, n23405, n23406, n23407, n23408,
         n23409, n23410, n23411, n23412, n23414, n23415, n23416, n23417,
         n23418, n23419, n23420, n23421, n23422, n23424, n23425, n23426,
         n23427, n23429, n23430, n23432, n23434, n23435, n23436, n23437,
         n23439, n23440, n23442, n23443, n23445, n23446, n23447, n23448,
         n23449, n23451, n23452, n23453, n23454, n23455, n23456, n23457,
         n23458, n23459, n23461, n23463, n23464, n23465, n23466, n23467,
         n23468, n23469, n23470, n23471, n23472, n23474, n23475, n23476,
         n23477, n23478, n23479, n23480, n23481, n23482, n23484, n23485,
         n23486, n23487, n23488, n23489, n23490, n23491, n23492, n23493,
         n23495, n23496, n23497, n23498, n23500, n23501, n23502, n23503,
         n23504, n23505, n23506, n23507, n23508, n23509, n23510, n23514,
         n23515, n23516, n23517, n23518, n23519, n23520, n23522, n23525,
         n23526, n23528, n23529, n23531, n23532, n23533, n23534, n23535,
         n23537, n23538, n23540, n23541, n23542, n23544, n23545, n23546,
         n23547, n23548, n23549, n23550, n23551, n23552, n23553, n23554,
         n23555, n23556, n23557, n23558, n23559, n23561, n23562, n23563,
         n23564, n23565, n23566, n23567, n23568, n23569, n23571, n23572,
         n23573, n23574, n23575, n23576, n23577, n23578, n23579, n23580,
         n23581, n23582, n23583, n23584, n23585, n23586, n23587, n23588,
         n23589, n23590, n23591, n23592, n23594, n23595, n23596, n23597,
         n23598, n23599, n23600, n23601, n23602, n23603, n23604, n23606,
         n23608, n23610, n23611, n23612, n23613, n23614, n23616, n23617,
         n23618, n23619, n23620, n23622, n23623, n23624, n23625, n23626,
         n23627, n23628, n23629, n23630, n23631, n23633, n23634, n23635,
         n23636, n23637, n23638, n23639, n23640, n23641, n23642, n23643,
         n23644, n23645, n23646, n23647, n23648, n23649, n23650, n23651,
         n23652, n23654, n23655, n23656, n23658, n23659, n23661, n23663,
         n23665, n23666, n23667, n23668, n23669, n23670, n23674, n23676,
         n23677, n23678, n23679, n23680, n23681, n23682, n23683, n23685,
         n23687, n23688, n23689, n23690, n23692, n23693, n23695, n23696,
         n23697, n23698, n23699, n23700, n23701, n23702, n23703, n23704,
         n23705, n23706, n23707, n23708, n23709, n23711, n23712, n23713,
         n23714, n23716, n23717, n23718, n23719, n23720, n23721, n23722,
         n23723, n23724, n23726, n23727, n23730, n23731, n23732, n23733,
         n23734, n23735, n23736, n23737, n23738, n23739, n23740, n23741,
         n23742, n23743, n23744, n23745, n23746, n23747, n23748, n23749,
         n23750, n23752, n23753, n23754, n23756, n23757, n23758, n23759,
         n23760, n23761, n23762, n23763, n23764, n23765, n23766, n23767,
         n23768, n23769, n23770, n23771, n23772, n23773, n23774, n23775,
         n23777, n23778, n23779, n23780, n23781, n23782, n23783, n23784,
         n23785, n23786, n23787, n23789, n23790, n23791, n23792, n23793,
         n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801,
         n23802, n23804, n23805, n23807, n23808, n23809, n23810, n23811,
         n23812, n23813, n23814, n23816, n23817, n23818, n23819, n23821,
         n23822, n23823, n23824, n23825, n23826, n23827, n23828, n23829,
         n23830, n23831, n23832, n23833, n23834, n23835, n23836, n23837,
         n23838, n23839, n23840, n23841, n23842, n23845, n23849, n23850,
         n23851, n23852, n23853, n23855, n23856, n23857, n23858, n23859,
         n23860, n23861, n23862, n23863, n23865, n23866, n23869, n23870,
         n23871, n23872, n23873, n23874, n23875, n23876, n23877, n23878,
         n23879, n23880, n23881, n23882, n23883, n23884, n23885, n23886,
         n23887, n23888, n23890, n23891, n23892, n23893, n23894, n23895,
         n23897, n23898, n23899, n23900, n23901, n23902, n23903, n23904,
         n23905, n23906, n23907, n23908, n23909, n23910, n23912, n23914,
         n23915, n23916, n23917, n23918, n23919, n23920, n23921, n23922,
         n23924, n23925, n23926, n23927, n23928, n23929, n23930, n23931,
         n23932, n23933, n23934, n23935, n23936, n23937, n23938, n23939,
         n23940, n23941, n23942, n23943, n23944, n23945, n23947, n23949,
         n23950, n23952, n23953, n23954, n23955, n23956, n23957, n23962,
         n23964, n23965, n23967, n23968, n23969, n23970, n23971, n23972,
         n23973, n23974, n23975, n23976, n23977, n23979, n23980, n23982,
         n23983, n23984, n23985, n23986, n23987, n23988, n23989, n23990,
         n23991, n23992, n23993, n23994, n23995, n23996, n23997, n23998,
         n23999, n24000, n24001, n24002, n24003, n24004, n24005, n24006,
         n24007, n24008, n24009, n24010, n24011, n24012, n24013, n24014,
         n24017, n24018, n24019, n24020, n24021, n24022, n24023, n24024,
         n24025, n24027, n24028, n24030, n24031, n24032, n24033, n24034,
         n24035, n24036, n24037, n24038, n24039, n24040, n24041, n24043,
         n24044, n24046, n24047, n24048, n24049, n24050, n24051, n24052,
         n24053, n24054, n24055, n24056, n24057, n24058, n24059, n24060,
         n24061, n24062, n24063, n24064, n24065, n24066, n24067, n24068,
         n24069, n24071, n24072, n24073, n24074, n24075, n24076, n24077,
         n24078, n24079, n24080, n24081, n24083, n24084, n24085, n24086,
         n24087, n24088, n24089, n24090, n24091, n24092, n24093, n24094,
         n24095, n24096, n24097, n24098, n24099, n24100, n24101, n24102,
         n24103, n24105, n24108, n24109, n24110, n24111, n24112, n24113,
         n24114, n24115, n24117, n24118, n24120, n24121, n24122, n24123,
         n24124, n24126, n24128, n24129, n24130, n24132, n24133, n24134,
         n24135, n24136, n24138, n24139, n24140, n24141, n24142, n24144,
         n24145, n24146, n24147, n24148, n24150, n24151, n24152, n24153,
         n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161,
         n24162, n24163, n24164, n24165, n24166, n24167, n24169, n24170,
         n24171, n24172, n24173, n24174, n24176, n24177, n24178, n24179,
         n24180, n24181, n24182, n24183, n24184, n24185, n24188, n24189,
         n24190, n24191, n24192, n24193, n24194, n24195, n24196, n24197,
         n24198, n24199, n24200, n24201, n24202, n24203, n24204, n24205,
         n24206, n24207, n24208, n24209, n24210, n24211, n24212, n24213,
         n24214, n24215, n24216, n24217, n24219, n24221, n24222, n24223,
         n24224, n24225, n24226, n24227, n24228, n24229, n24230, n24231,
         n24232, n24233, n24234, n24235, n24236, n24238, n24239, n24240,
         n24241, n24243, n24244, n24246, n24247, n24248, n24249, n24250,
         n24251, n24252, n24254, n24255, n24256, n24257, n24258, n24259,
         n24261, n24262, n24263, n24264, n24265, n24266, n24267, n24270,
         n24271, n24272, n24273, n24274, n24275, n24276, n24277, n24278,
         n24279, n24282, n24283, n24284, n24286, n24287, n24290, n24291,
         n24292, n24293, n24294, n24295, n24296, n24297, n24298, n24299,
         n24300, n24301, n24302, n24304, n24305, n24306, n24309, n24310,
         n24311, n24312, n24313, n24314, n24315, n24316, n24317, n24318,
         n24319, n24320, n24321, n24322, n24323, n24324, n24325, n24326,
         n24327, n24328, n24329, n24330, n24331, n24332, n24333, n24334,
         n24335, n24336, n24337, n24338, n24339, n24340, n24341, n24342,
         n24343, n24344, n24345, n24346, n24347, n24348, n24349, n24350,
         n24351, n24352, n24353, n24354, n24355, n24356, n24357, n24358,
         n24359, n24360, n24361, n24362, n24363, n24364, n24365, n24366,
         n24367, n24368, n24370, n24371, n24373, n24374, n24375, n24376,
         n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385,
         n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393,
         n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401,
         n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409,
         n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24418,
         n24419, n24420, n24421, n24422, n24424, n24425, n24427, n24428,
         n24429, n24430, n24431, n24432, n24434, n24435, n24436, n24437,
         n24438, n24439, n24440, n24441, n24442, n24444, n24447, n24448,
         n24449, n24450, n24451, n24452, n24453, n24454, n24455, n24457,
         n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465,
         n24466, n24467, n24468, n24470, n24471, n24472, n24473, n24475,
         n24476, n24477, n24479, n24480, n24481, n24482, n24483, n24485,
         n24486, n24488, n24489, n24490, n24491, n24492, n24493, n24494,
         n24496, n24497, n24498, n24499, n24501, n24502, n24503, n24504,
         n24505, n24506, n24508, n24509, n24510, n24511, n24512, n24513,
         n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521,
         n24522, n24523, n24524, n24526, n24527, n24529, n24530, n24533,
         n24534, n24535, n24536, n24537, n24538, n24539, n24540, n24541,
         n24543, n24544, n24545, n24547, n24548, n24549, n24550, n24551,
         n24552, n24553, n24555, n24556, n24557, n24558, n24559, n24560,
         n24561, n24562, n24563, n24564, n24566, n24568, n24569, n24570,
         n24571, n24574, n24575, n24576, n24577, n24578, n24579, n24580,
         n24581, n24582, n24583, n24584, n24585, n24586, n24589, n24591,
         n24592, n24593, n24594, n24595, n24596, n24597, n24598, n24599,
         n24600, n24603, n24606, n24607, n24608, n24609, n24610, n24611,
         n24612, n24613, n24614, n24615, n24617, n24618, n24621, n24622,
         n24623, n24624, n24625, n24626, n24627, n24628, n24629, n24630,
         n24631, n24632, n24633, n24634, n24635, n24636, n24637, n24638,
         n24639, n24640, n24641, n24643, n24644, n24645, n24646, n24647,
         n24648, n24649, n24650, n24651, n24653, n24654, n24656, n24658,
         n24659, n24660, n24661, n24662, n24663, n24664, n24666, n24667,
         n24668, n24669, n24670, n24671, n24672, n24673, n24674, n24675,
         n24676, n24677, n24679, n24680, n24681, n24682, n24683, n24684,
         n24685, n24686, n24688, n24689, n24690, n24691, n24692, n24694,
         n24696, n24697, n24698, n24699, n24700, n24701, n24702, n24703,
         n24704, n24706, n24708, n24710, n24711, n24712, n24713, n24714,
         n24715, n24716, n24717, n24719, n24720, n24721, n24722, n24723,
         n24724, n24725, n24726, n24728, n24729, n24730, n24731, n24732,
         n24733, n24734, n24735, n24737, n24739, n24742, n24743, n24744,
         n24745, n24746, n24748, n24749, n24750, n24751, n24752, n24753,
         n24755, n24756, n24757, n24758, n24759, n24760, n24762, n24764,
         n24765, n24766, n24767, n24768, n24770, n24774, n24775, n24776,
         n24777, n24779, n24780, n24781, n24782, n24784, n24785, n24786,
         n24787, n24788, n24790, n24791, n24792, n24794, n24796, n24797,
         n24798, n24799, n24801, n24802, n24803, n24804, n24805, n24806,
         n24807, n24808, n24809, n24810, n24811, n24812, n24813, n24815,
         n24816, n24817, n24818, n24820, n24821, n24822, n24823, n24824,
         n24825, n24826, n24827, n24828, n24829, n24830, n24831, n24834,
         n24835, n24836, n24837, n24838, n24839, n24840, n24842, n24844,
         n24848, n24849, n24850, n24851, n24852, n24853, n24854, n24855,
         n24856, n24858, n24859, n24860, n24861, n24862, n24863, n24864,
         n24865, n24866, n24867, n24868, n24869, n24870, n24871, n24872,
         n24873, n24874, n24875, n24877, n24878, n24879, n24880, n24881,
         n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889,
         n24890, n24891, n24893, n24894, n24895, n24896, n24897, n24898,
         n24900, n24901, n24902, n24903, n24904, n24906, n24908, n24909,
         n24911, n24912, n24913, n24915, n24916, n24917, n24918, n24919,
         n24920, n24921, n24922, n24923, n24924, n24925, n24926, n24927,
         n24928, n24929, n24930, n24931, n24932, n24933, n24934, n24935,
         n24940, n24941, n24942, n24943, n24944, n24945, n24946, n24947,
         n24948, n24949, n24950, n24951, n24952, n24953, n24954, n24956,
         n24957, n24958, n24959, n24960, n24961, n24962, n24963, n24964,
         n24965, n24966, n24967, n24968, n24969, n24970, n24973, n24974,
         n24975, n24976, n24977, n24978, n24979, n24980, n24981, n24982,
         n24983, n24984, n24985, n24987, n24988, n24989, n24990, n24991,
         n24992, n24993, n24994, n24996, n24997, n24999, n25000, n25001,
         n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009,
         n25010, n25011, n25012, n25013, n25014, n25016, n25017, n25018,
         n25020, n25021, n25022, n25023, n25025, n25026, n25027, n25029,
         n25030, n25031, n25032, n25033, n25034, n25035, n25036, n25037,
         n25038, n25039, n25040, n25041, n25042, n25043, n25044, n25046,
         n25047, n25048, n25050, n25051, n25052, n25053, n25054, n25055,
         n25056, n25058, n25059, n25060, n25061, n25062, n25063, n25064,
         n25065, n25066, n25067, n25068, n25069, n25070, n25071, n25072,
         n25073, n25074, n25075, n25076, n25077, n25078, n25080, n25081,
         n25082, n25083, n25085, n25086, n25087, n25088, n25089, n25090,
         n25091, n25092, n25093, n25094, n25095, n25096, n25098, n25099,
         n25100, n25101, n25103, n25104, n25106, n25107, n25109, n25110,
         n25111, n25112, n25113, n25115, n25116, n25117, n25118, n25119,
         n25120, n25121, n25124, n25125, n25126, n25127, n25128, n25129,
         n25130, n25131, n25132, n25134, n25136, n25137, n25138, n25139,
         n25140, n25141, n25142, n25144, n25145, n25146, n25147, n25148,
         n25149, n25150, n25151, n25152, n25154, n25155, n25156, n25157,
         n25158, n25159, n25160, n25161, n25162, n25163, n25164, n25165,
         n25166, n25167, n25168, n25169, n25170, n25171, n25172, n25173,
         n25174, n25175, n25176, n25177, n25179, n25180, n25181, n25182,
         n25183, n25184, n25185, n25186, n25187, n25188, n25190, n25191,
         n25192, n25193, n25194, n25196, n25197, n25198, n25199, n25200,
         n25201, n25202, n25203, n25204, n25205, n25206, n25208, n25209,
         n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25218,
         n25219, n25220, n25221, n25222, n25224, n25225, n25227, n25229,
         n25230, n25231, n25232, n25233, n25235, n25236, n25237, n25238,
         n25239, n25240, n25241, n25242, n25243, n25244, n25245, n25246,
         n25247, n25248, n25249, n25250, n25251, n25252, n25253, n25254,
         n25256, n25257, n25258, n25259, n25261, n25262, n25263, n25264,
         n25265, n25266, n25267, n25268, n25269, n25270, n25272, n25273,
         n25274, n25275, n25277, n25279, n25280, n25281, n25282, n25283,
         n25284, n25285, n25286, n25287, n25288, n25290, n25292, n25293,
         n25294, n25296, n25297, n25298, n25299, n25300, n25301, n25302,
         n25304, n25305, n25306, n25307, n25308, n25309, n25310, n25311,
         n25312, n25313, n25314, n25315, n25316, n25317, n25318, n25320,
         n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329,
         n25331, n25332, n25333, n25334, n25336, n25337, n25338, n25339,
         n25340, n25341, n25342, n25343, n25344, n25345, n25346, n25347,
         n25348, n25349, n25350, n25351, n25352, n25353, n25354, n25355,
         n25356, n25357, n25358, n25359, n25360, n25361, n25362, n25363,
         n25364, n25365, n25366, n25367, n25368, n25370, n25371, n25372,
         n25373, n25374, n25375, n25376, n25377, n25378, n25381, n25383,
         n25384, n25385, n25386, n25387, n25388, n25389, n25390, n25391,
         n25392, n25393, n25394, n25395, n25396, n25397, n25398, n25399,
         n25401, n25402, n25403, n25404, n25405, n25407, n25409, n25410,
         n25411, n25412, n25413, n25414, n25415, n25416, n25417, n25418,
         n25419, n25420, n25421, n25422, n25423, n25424, n25426, n25427,
         n25428, n25429, n25430, n25432, n25433, n25434, n25435, n25437,
         n25438, n25439, n25440, n25442, n25443, n25444, n25445, n25446,
         n25447, n25448, n25449, n25450, n25451, n25452, n25453, n25454,
         n25455, n25456, n25457, n25458, n25459, n25461, n25462, n25465,
         n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473,
         n25474, n25475, n25476, n25477, n25479, n25480, n25481, n25482,
         n25483, n25484, n25486, n25487, n25488, n25489, n25490, n25491,
         n25492, n25493, n25494, n25495, n25497, n25499, n25500, n25501,
         n25502, n25503, n25504, n25506, n25507, n25508, n25509, n25510,
         n25511, n25512, n25513, n25514, n25515, n25516, n25517, n25518,
         n25519, n25522, n25524, n25525, n25526, n25527, n25528, n25529,
         n25530, n25531, n25532, n25533, n25534, n25535, n25537, n25538,
         n25541, n25542, n25545, n25546, n25547, n25548, n25549, n25550,
         n25551, n25553, n25555, n25556, n25557, n25558, n25559, n25561,
         n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569,
         n25570, n25571, n25572, n25574, n25575, n25576, n25578, n25579,
         n25580, n25582, n25584, n25585, n25586, n25589, n25590, n25591,
         n25592, n25594, n25595, n25596, n25598, n25599, n25600, n25601,
         n25602, n25603, n25604, n25605, n25606, n25608, n25609, n25610,
         n25611, n25612, n25616, n25617, n25618, n25619, n25620, n25621,
         n25622, n25623, n25624, n25625, n25626, n25627, n25628, n25629,
         n25630, n25631, n25632, n25633, n25634, n25635, n25636, n25637,
         n25638, n25639, n25640, n25641, n25642, n25643, n25644, n25645,
         n25646, n25647, n25648, n25649, n25650, n25651, n25652, n25653,
         n25654, n25657, n25658, n25659, n25660, n25661, n25663, n25664,
         n25665, n25666, n25667, n25668, n25669, n25670, n25671, n25672,
         n25675, n25676, n25677, n25679, n25680, n25681, n25682, n25683,
         n25684, n25685, n25686, n25687, n25688, n25689, n25690, n25691,
         n25692, n25693, n25694, n25695, n25696, n25697, n25698, n25700,
         n25701, n25702, n25703, n25704, n25705, n25706, n25707, n25708,
         n25709, n25710, n25711, n25712, n25713, n25714, n25715, n25716,
         n25717, n25718, n25719, n25720, n25721, n25722, n25724, n25725,
         n25728, n25729, n25730, n25731, n25732, n25733, n25734, n25735,
         n25736, n25737, n25738, n25739, n25740, n25741, n25742, n25743,
         n25744, n25745, n25746, n25747, n25749, n25751, n25752, n25753,
         n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25762,
         n25763, n25764, n25765, n25766, n25767, n25769, n25770, n25771,
         n25772, n25773, n25774, n25775, n25776, n25777, n25779, n25781,
         n25783, n25784, n25785, n25786, n25787, n25788, n25789, n25790,
         n25791, n25792, n25793, n25794, n25795, n25797, n25798, n25800,
         n25801, n25803, n25804, n25805, n25806, n25807, n25809, n25810,
         n25811, n25812, n25813, n25814, n25815, n25816, n25817, n25818,
         n25819, n25820, n25821, n25822, n25823, n25824, n25825, n25826,
         n25828, n25830, n25831, n25833, n25835, n25836, n25837, n25838,
         n25839, n25840, n25841, n25842, n25843, n25844, n25845, n25847,
         n25848, n25849, n25850, n25851, n25852, n25853, n25854, n25855,
         n25856, n25857, n25858, n25859, n25860, n25861, n25862, n25863,
         n25864, n25865, n25866, n25867, n25868, n25869, n25870, n25872,
         n25873, n25874, n25876, n25877, n25878, n25879, n25881, n25882,
         n25884, n25885, n25886, n25887, n25888, n25891, n25893, n25894,
         n25895, n25896, n25897, n25898, n25899, n25900, n25903, n25904,
         n25905, n25906, n25907, n25909, n25910, n25911, n25912, n25913,
         n25914, n25915, n25918, n25919, n25920, n25921, n25922, n25923,
         n25924, n25925, n25926, n25927, n25928, n25929, n25930, n25931,
         n25932, n25933, n25934, n25935, n25936, n25937, n25938, n25939,
         n25940, n25942, n25943, n25944, n25946, n25947, n25948, n25949,
         n25951, n25952, n25953, n25954, n25955, n25956, n25957, n25958,
         n25959, n25960, n25961, n25962, n25963, n25964, n25965, n25966,
         n25967, n25968, n25969, n25970, n25972, n25973, n25975, n25976,
         n25978, n25979, n25980, n25982, n25983, n25984, n25986, n25987,
         n25988, n25989, n25990, n25991, n25992, n25993, n25994, n25995,
         n25996, n25997, n25998, n25999, n26000, n26002, n26003, n26004,
         n26006, n26007, n26008, n26009, n26010, n26011, n26012, n26014,
         n26015, n26016, n26017, n26019, n26020, n26021, n26022, n26023,
         n26024, n26025, n26026, n26027, n26028, n26029, n26030, n26031,
         n26032, n26034, n26035, n26036, n26037, n26038, n26039, n26040,
         n26041, n26043, n26044, n26045, n26046, n26047, n26048, n26049,
         n26050, n26052, n26053, n26054, n26056, n26057, n26058, n26059,
         n26060, n26061, n26062, n26063, n26064, n26065, n26066, n26067,
         n26069, n26070, n26071, n26072, n26074, n26075, n26076, n26077,
         n26078, n26079, n26080, n26081, n26084, n26085, n26086, n26087,
         n26088, n26089, n26090, n26091, n26092, n26093, n26094, n26095,
         n26096, n26097, n26098, n26099, n26100, n26101, n26102, n26103,
         n26104, n26105, n26107, n26108, n26109, n26110, n26111, n26112,
         n26113, n26114, n26117, n26118, n26119, n26120, n26121, n26122,
         n26124, n26125, n26126, n26127, n26128, n26129, n26130, n26131,
         n26132, n26133, n26134, n26135, n26138, n26139, n26141, n26142,
         n26143, n26144, n26145, n26146, n26147, n26148, n26150, n26151,
         n26153, n26154, n26155, n26156, n26158, n26159, n26160, n26161,
         n26162, n26163, n26165, n26166, n26167, n26168, n26169, n26170,
         n26171, n26172, n26173, n26174, n26175, n26176, n26178, n26179,
         n26180, n26181, n26182, n26183, n26184, n26185, n26186, n26187,
         n26189, n26190, n26191, n26192, n26194, n26196, n26198, n26200,
         n26201, n26202, n26204, n26205, n26206, n26208, n26209, n26210,
         n26211, n26212, n26213, n26214, n26216, n26217, n26218, n26219,
         n26220, n26221, n26222, n26223, n26224, n26226, n26227, n26228,
         n26229, n26231, n26232, n26234, n26235, n26236, n26237, n26238,
         n26239, n26240, n26241, n26242, n26243, n26245, n26246, n26247,
         n26248, n26250, n26251, n26252, n26253, n26254, n26255, n26256,
         n26257, n26258, n26260, n26262, n26263, n26264, n26265, n26266,
         n26267, n26268, n26269, n26270, n26271, n26272, n26273, n26274,
         n26275, n26276, n26277, n26278, n26279, n26280, n26281, n26282,
         n26283, n26284, n26285, n26286, n26287, n26288, n26289, n26292,
         n26293, n26294, n26296, n26297, n26298, n26299, n26300, n26301,
         n26302, n26303, n26304, n26305, n26306, n26307, n26308, n26310,
         n26311, n26312, n26313, n26314, n26315, n26316, n26317, n26318,
         n26319, n26320, n26321, n26322, n26323, n26324, n26325, n26326,
         n26327, n26328, n26329, n26330, n26331, n26332, n26333, n26334,
         n26335, n26336, n26337, n26338, n26339, n26340, n26341, n26342,
         n26343, n26344, n26345, n26346, n26347, n26348, n26349, n26350,
         n26351, n26352, n26353, n26354, n26355, n26356, n26357, n26358,
         n26359, n26360, n26361, n26362, n26363, n26364, n26365, n26366,
         n26367, n26368, n26369, n26370, n26371, n26372, n26373, n26374,
         n26375, n26376, n26377, n26378, n26379, n26380, n26381, n26383,
         n26384, n26385, n26386, n26387, n26388, n26389, n26390, n26391,
         n26393, n26394, n26395, n26396, n26397, n26398, n26399, n26400,
         n26401, n26402, n26403, n26404, n26405, n26406, n26407, n26408,
         n26409, n26410, n26411, n26412, n26413, n26414, n26415, n26416,
         n26417, n26418, n26419, n26420, n26421, n26422, n26423, n26424,
         n26425, n26426, n26427, n26428, n26429, n26430, n26431, n26432,
         n26433, n26434, n26435, n26436, n26437, n26438, n26439, n26440,
         n26441, n26444, n26445, n26446, n26447, n26448, n26449, n26450,
         n26451, n26452, n26453, n26454, n26455, n26456, n26457, n26458,
         n26459, n26460, n26461, n26462, n26463, n26464, n26465, n26467,
         n26468, n26469, n26470, n26471, n26472, n26473, n26475, n26476,
         n26477, n26479, n26480, n26481, n26482, n26483, n26484, n26485,
         n26487, n26488, n26489, n26490, n26491, n26492, n26493, n26494,
         n26495, n26496, n26497, n26498, n26499, n26500, n26501, n26502,
         n26503, n26504, n26505, n26506, n26507, n26508, n26509, n26510,
         n26511, n26512, n26514, n26515, n26516, n26517, n26518, n26519,
         n26520, n26521, n26522, n26523, n26524, n26525, n26526, n26527,
         n26528, n26529, n26530, n26531, n26532, n26533, n26534, n26535,
         n26536, n26537, n26538, n26539, n26540, n26541, n26542, n26543,
         n26544, n26546, n26547, n26548, n26549, n26550, n26551, n26552,
         n26553, n26554, n26555, n26556, n26557, n26558, n26559, n26560,
         n26561, n26562, n26563, n26564, n26565, n26566, n26567, n26568,
         n26569, n26570, n26571, n26572, n26573, n26574, n26575, n26576,
         n26577, n26578, n26579, n26580, n26581, n26582, n26583, n26585,
         n26586, n26587, n26588, n26589, n26591, n26592, n26593, n26594,
         n26595, n26596, n26597, n26598, n26599, n26600, n26601, n26602,
         n26603, n26604, n26605, n26606, n26607, n26608, n26609, n26610,
         n26611, n26612, n26613, n26614, n26615, n26616, n26618, n26619,
         n26620, n26621, n26622, n26623, n26624, n26625, n26626, n26627,
         n26628, n26629, n26630, n26631, n26632, n26633, n26634, n26635,
         n26636, n26637, n26638, n26639, n26640, n26641, n26642, n26643,
         n26644, n26645, n26646, n26647, n26648, n26649, n26650, n26651,
         n26652, n26653, n26654, n26655, n26656, n26657, n26658, n26660,
         n26661, n26662, n26663, n26664, n26665, n26666, n26667, n26668,
         n26669, n26670, n26671, n26672, n26673, n26674, n26675, n26676,
         n26677, n26678, n26679, n26680, n26682, n26683, n26684, n26685,
         n26686, n26687, n26688, n26689, n26690, n26691, n26692, n26693,
         n26694, n26695, n26696, n26698, n26699, n26700, n26701, n26702,
         n26703, n26704, n26705, n26706, n26707, n26708, n26709, n26710,
         n26711, n26712, n26713, n26714, n26715, n26716, n26717, n26718,
         n26719, n26720, n26721, n26723, n26724, n26725, n26726, n26728,
         n26730, n26732, n26733, n26734, n26735, n26736, n26737, n26738,
         n26739, n26740, n26741, n26742, n26743, n26744, n26745, n26746,
         n26747, n26749, n26750, n26752, n26753, n26754, n26755, n26756,
         n26757, n26758, n26759, n26760, n26761, n26762, n26763, n26764,
         n26765, n26766, n26767, n26768, n26769, n26770, n26771, n26772,
         n26773, n26776, n26777, n26778, n26779, n26780, n26781, n26782,
         n26783, n26784, n26785, n26786, n26787, n26788, n26789, n26790,
         n26791, n26792, n26793, n26794, n26795, n26796, n26797, n26798,
         n26799, n26800, n26801, n26802, n26804, n26805, n26806, n26807,
         n26808, n26809, n26810, n26811, n26812, n26813, n26814, n26815,
         n26816, n26817, n26818, n26819, n26820, n26821, n26822, n26823,
         n26824, n26825, n26826, n26827, n26828, n26830, n26831, n26832,
         n26833, n26834, n26835, n26836, n26837, n26838, n26839, n26840,
         n26841, n26842, n26843, n26844, n26845, n26846, n26847, n26848,
         n26849, n26850, n26851, n26852, n26853, n26854, n26856, n26857,
         n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865,
         n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873,
         n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881,
         n26882, n26883, n26884, n26885, n26886, n26887, n26888, n26889,
         n26890, n26891, n26892, n26893, n26895, n26896, n26897, n26898,
         n26900, n26901, n26903, n26905, n26906, n26907, n26910, n26911,
         n26912, n26913, n26914, n26916, n26918, n26919, n26920, n26921,
         n26922, n26923, n26924, n26925, n26926, n26927, n26928, n26929,
         n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937,
         n26938, n26940, n26941, n26942, n26944, n26945, n26946, n26948,
         n26949, n26950, n26951, n26952, n26953, n26954, n26955, n26956,
         n26957, n26958, n26959, n26960, n26961, n26963, n26964, n26965,
         n26966, n26967, n26968, n26969, n26970, n26971, n26972, n26973,
         n26974, n26975, n26976, n26977, n26978, n26979, n26980, n26981,
         n26982, n26983, n26985, n26986, n26987, n26988, n26989, n26990,
         n26991, n26992, n26993, n26994, n26997, n26998, n26999, n27000,
         n27001, n27003, n27004, n27005, n27006, n27007, n27008, n27010,
         n27011, n27013, n27014, n27015, n27016, n27017, n27018, n27020,
         n27021, n27022, n27023, n27024, n27025, n27026, n27027, n27028,
         n27029, n27030, n27031, n27032, n27033, n27035, n27036, n27037,
         n27038, n27039, n27040, n27042, n27043, n27044, n27045, n27047,
         n27048, n27049, n27050, n27051, n27052, n27053, n27054, n27056,
         n27057, n27058, n27059, n27060, n27061, n27062, n27063, n27064,
         n27065, n27066, n27067, n27068, n27069, n27071, n27072, n27073,
         n27074, n27075, n27076, n27077, n27078, n27079, n27080, n27081,
         n27082, n27083, n27084, n27085, n27087, n27088, n27090, n27091,
         n27092, n27093, n27094, n27095, n27096, n27097, n27098, n27099,
         n27100, n27101, n27102, n27103, n27104, n27105, n27106, n27107,
         n27108, n27109, n27111, n27112, n27113, n27114, n27115, n27117,
         n27118, n27120, n27121, n27122, n27123, n27124, n27125, n27126,
         n27127, n27128, n27129, n27130, n27131, n27132, n27133, n27134,
         n27135, n27136, n27137, n27138, n27139, n27140, n27141, n27142,
         n27143, n27144, n27145, n27146, n27147, n27149, n27150, n27151,
         n27152, n27153, n27154, n27155, n27156, n27157, n27158, n27159,
         n27160, n27161, n27162, n27163, n27164, n27165, n27166, n27168,
         n27169, n27170, n27171, n27172, n27173, n27174, n27175, n27176,
         n27177, n27178, n27179, n27180, n27181, n27182, n27183, n27184,
         n27185, n27187, n27188, n27189, n27190, n27191, n27192, n27193,
         n27194, n27195, n27196, n27197, n27198, n27199, n27200, n27201,
         n27202, n27203, n27204, n27205, n27206, n27207, n27208, n27209,
         n27210, n27211, n27212, n27213, n27214, n27215, n27216, n27217,
         n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225,
         n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233,
         n27234, n27235, n27236, n27238, n27239, n27240, n27241, n27242,
         n27243, n27244, n27245, n27246, n27247, n27248, n27249, n27250,
         n27251, n27254, n27255, n27256, n27258, n27259, n27260, n27261,
         n27262, n27263, n27264, n27265, n27266, n27267, n27268, n27269,
         n27270, n27271, n27272, n27273, n27274, n27275, n27276, n27277,
         n27278, n27279, n27280, n27282, n27283, n27284, n27285, n27286,
         n27287, n27288, n27289, n27290, n27291, n27292, n27293, n27295,
         n27296, n27298, n27299, n27300, n27301, n27302, n27303, n27304,
         n27305, n27306, n27307, n27308, n27309, n27310, n27311, n27312,
         n27313, n27314, n27315, n27316, n27317, n27318, n27320, n27321,
         n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329,
         n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337,
         n27338, n27339, n27340, n27341, n27342, n27343, n27344, n27345,
         n27346, n27347, n27348, n27349, n27350, n27351, n27352, n27353,
         n27354, n27355, n27356, n27357, n27358, n27360, n27361, n27362,
         n27363, n27365, n27366, n27367, n27368, n27369, n27370, n27371,
         n27372, n27373, n27374, n27375, n27376, n27377, n27378, n27379,
         n27380, n27381, n27382, n27383, n27384, n27385, n27386, n27387,
         n27388, n27389, n27390, n27391, n27392, n27393, n27394, n27395,
         n27396, n27397, n27398, n27399, n27400, n27401, n27402, n27403,
         n27404, n27405, n27406, n27407, n27408, n27409, n27410, n27411,
         n27412, n27413, n27414, n27415, n27416, n27417, n27418, n27419,
         n27421, n27422, n27423, n27424, n27425, n27426, n27427, n27428,
         n27429, n27430, n27431, n27432, n27433, n27434, n27435, n27436,
         n27437, n27438, n27439, n27440, n27441, n27442, n27443, n27444,
         n27445, n27446, n27447, n27448, n27449, n27450, n27451, n27452,
         n27453, n27454, n27455, n27457, n27458, n27459, n27460, n27464,
         n27465, n27466, n27467, n27469, n27470, n27471, n27472, n27473,
         n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481,
         n27482, n27483, n27484, n27485, n27486, n27487, n27488, n27489,
         n27491, n27492, n27493, n27494, n27495, n27496, n27497, n27498,
         n27499, n27500, n27501, n27502, n27503, n27504, n27505, n27506,
         n27507, n27508, n27509, n27510, n27511, n27512, n27513, n27514,
         n27515, n27516, n27517, n27518, n27519, n27520, n27521, n27522,
         n27523, n27524, n27525, n27526, n27527, n27528, n27529, n27530,
         n27531, n27532, n27533, n27534, n27535, n27536, n27537, n27538,
         n27539, n27540, n27541, n27542, n27543, n27544, n27545, n27546,
         n27547, n27548, n27549, n27550, n27551, n27552, n27553, n27554,
         n27555, n27556, n27557, n27558, n27559, n27560, n27561, n27562,
         n27563, n27564, n27565, n27566, n27567, n27568, n27569, n27570,
         n27571, n27572, n27573, n27574, n27575, n27576, n27577, n27578,
         n27579, n27580, n27581, n27582, n27583, n27584, n27585, n27586,
         n27587, n27588, n27589, n27590, n27591, n27592, n27593, n27594,
         n27595, n27596, n27597, n27598, n27599, n27600, n27601, n27602,
         n27603, n27604, n27605, n27606, n27607, n27608, n27609, n27610,
         n27611, n27612, n27613, n27614, n27615, n27616, n27617, n27618,
         n27619, n27620, n27621, n27622, n27623, n27624, n27625, n27626,
         n27627, n27628, n27629, n27630, n27631, n27632, n27633, n27634,
         n27635, n27637, n27638, n27639, n27640, n27641, n27642, n27643,
         n27644, n27646, n27647, n27648, n27649, n27650, n27651, n27653,
         n27654, n27655, n27656, n27657, n27658, n27660, n27661, n27662,
         n27663, n27664, n27665, n27666, n27668, n27669, n27670, n27671,
         n27672, n27673, n27674, n27675, n27676, n27677, n27678, n27679,
         n27680, n27681, n27682, n27683, n27684, n27685, n27686, n27687,
         n27689, n27690, n27691, n27692, n27693, n27694, n27695, n27696,
         n27697, n27698, n27699, n27700, n27701, n27702, n27703, n27704,
         n27705, n27706, n27708, n27709, n27710, n27712, n27713, n27714,
         n27715, n27716, n27717, n27718, n27719, n27720, n27721, n27722,
         n27724, n27725, n27727, n27728, n27729, n27730, n27731, n27732,
         n27733, n27734, n27735, n27736, n27737, n27738, n27739, n27740,
         n27741, n27742, n27743, n27744, n27746, n27748, n27749, n27750,
         n27751, n27752, n27753, n27754, n27756, n27757, n27758, n27759,
         n27761, n27762, n27763, n27764, n27765, n27766, n27767, n27768,
         n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27777,
         n27778, n27779, n27780, n27781, n27782, n27783, n27784, n27785,
         n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793,
         n27794, n27795, n27796, n27797, n27798, n27799, n27800, n27801,
         n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809,
         n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817,
         n27818, n27819, n27820, n27821, n27822, n27823, n27824, n27825,
         n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833,
         n27834, n27836, n27837, n27838, n27839, n27840, n27841, n27842,
         n27843, n27844, n27845, n27846, n27847, n27849, n27850, n27851,
         n27852, n27853, n27854, n27855, n27856, n27857, n27858, n27859,
         n27860, n27861, n27862, n27863, n27864, n27865, n27866, n27868,
         n27869, n27870, n27871, n27872, n27873, n27874, n27875, n27876,
         n27877, n27878, n27879, n27880, n27882, n27883, n27884, n27885,
         n27886, n27887, n27888, n27889, n27890, n27891, n27892, n27893,
         n27894, n27895, n27896, n27897, n27898, n27899, n27900, n27902,
         n27903, n27904, n27905, n27906, n27907, n27908, n27909, n27910,
         n27911, n27912, n27913, n27914, n27915, n27916, n27917, n27918,
         n27919, n27920, n27921, n27922, n27923, n27924, n27925, n27926,
         n27927, n27928, n27929, n27930, n27931, n27932, n27933, n27934,
         n27935, n27936, n27937, n27938, n27939, n27940, n27941, n27943,
         n27944, n27945, n27946, n27948, n27949, n27950, n27951, n27954,
         n27955, n27956, n27957, n27958, n27959, n27960, n27961, n27962,
         n27963, n27964, n27965, n27966, n27967, n27968, n27969, n27970,
         n27971, n27972, n27973, n27974, n27975, n27976, n27977, n27978,
         n27979, n27980, n27981, n27982, n27983, n27984, n27985, n27988,
         n27989, n27990, n27991, n27992, n27993, n27994, n27995, n27996,
         n27997, n27998, n28000, n28001, n28002, n28003, n28004, n28005,
         n28006, n28007, n28008, n28011, n28012, n28013, n28014, n28015,
         n28016, n28017, n28018, n28020, n28021, n28022, n28023, n28024,
         n28025, n28026, n28027, n28028, n28029, n28030, n28031, n28032,
         n28033, n28034, n28035, n28036, n28037, n28038, n28039, n28040,
         n28042, n28043, n28044, n28045, n28046, n28047, n28048, n28049,
         n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057,
         n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28065,
         n28066, n28067, n28068, n28069, n28070, n28071, n28072, n28073,
         n28074, n28075, n28076, n28077, n28078, n28079, n28080, n28081,
         n28082, n28083, n28084, n28085, n28086, n28087, n28088, n28090,
         n28091, n28092, n28093, n28094, n28095, n28096, n28097, n28098,
         n28099, n28100, n28101, n28102, n28103, n28104, n28105, n28106,
         n28107, n28108, n28109, n28110, n28111, n28112, n28113, n28114,
         n28115, n28116, n28117, n28118, n28119, n28120, n28121, n28122,
         n28123, n28124, n28125, n28126, n28127, n28128, n28129, n28130,
         n28131, n28132, n28133, n28134, n28135, n28136, n28137, n28138,
         n28139, n28140, n28141, n28142, n28143, n28144, n28145, n28146,
         n28147, n28148, n28149, n28150, n28151, n28155, n28156, n28157,
         n28158, n28159, n28160, n28161, n28162, n28163, n28164, n28165,
         n28166, n28167, n28168, n28169, n28170, n28171, n28172, n28173,
         n28174, n28175, n28176, n28177, n28178, n28180, n28182, n28183,
         n28184, n28185, n28186, n28187, n28188, n28189, n28190, n28191,
         n28192, n28193, n28194, n28195, n28196, n28197, n28198, n28199,
         n28200, n28201, n28202, n28204, n28205, n28206, n28207, n28208,
         n28209, n28210, n28211, n28212, n28213, n28214, n28216, n28217,
         n28218, n28219, n28220, n28221, n28222, n28223, n28224, n28225,
         n28226, n28227, n28228, n28229, n28230, n28231, n28232, n28233,
         n28234, n28235, n28236, n28237, n28238, n28239, n28240, n28241,
         n28242, n28243, n28244, n28245, n28246, n28247, n28248, n28250,
         n28252, n28253, n28254, n28255, n28256, n28257, n28258, n28259,
         n28260, n28261, n28262, n28264, n28265, n28266, n28267, n28268,
         n28269, n28270, n28271, n28272, n28273, n28274, n28275, n28276,
         n28277, n28278, n28279, n28280, n28281, n28282, n28283, n28284,
         n28285, n28286, n28287, n28288, n28289, n28290, n28291, n28293,
         n28294, n28295, n28296, n28297, n28298, n28299, n28300, n28301,
         n28302, n28303, n28304, n28305, n28306, n28307, n28308, n28309,
         n28310, n28311, n28312, n28313, n28314, n28315, n28316, n28317,
         n28318, n28319, n28320, n28321, n28322, n28323, n28324, n28325,
         n28326, n28327, n28328, n28329, n28330, n28331, n28332, n28333,
         n28334, n28335, n28336, n28337, n28338, n28339, n28340, n28341,
         n28342, n28343, n28344, n28345, n28346, n28347, n28348, n28349,
         n28350, n28351, n28352, n28353, n28354, n28355, n28356, n28357,
         n28359, n28360, n28361, n28362, n28363, n28364, n28366, n28367,
         n28368, n28369, n28370, n28371, n28372, n28374, n28375, n28376,
         n28377, n28378, n28379, n28380, n28381, n28382, n28383, n28384,
         n28386, n28387, n28388, n28390, n28391, n28393, n28394, n28395,
         n28396, n28397, n28398, n28399, n28400, n28401, n28402, n28403,
         n28405, n28406, n28407, n28409, n28410, n28411, n28412, n28413,
         n28414, n28415, n28416, n28417, n28418, n28419, n28420, n28421,
         n28422, n28423, n28424, n28425, n28426, n28427, n28428, n28429,
         n28430, n28432, n28433, n28434, n28435, n28436, n28437, n28438,
         n28440, n28441, n28442, n28444, n28445, n28446, n28447, n28448,
         n28449, n28450, n28451, n28452, n28453, n28454, n28455, n28456,
         n28457, n28458, n28459, n28460, n28461, n28462, n28463, n28464,
         n28465, n28466, n28467, n28468, n28469, n28470, n28471, n28472,
         n28473, n28474, n28475, n28476, n28477, n28478, n28479, n28480,
         n28481, n28483, n28484, n28485, n28486, n28487, n28488, n28489,
         n28490, n28491, n28492, n28494, n28495, n28496, n28497, n28498,
         n28499, n28500, n28501, n28502, n28503, n28504, n28505, n28506,
         n28507, n28508, n28509, n28510, n28511, n28512, n28513, n28514,
         n28515, n28516, n28517, n28518, n28519, n28520, n28521, n28522,
         n28523, n28524, n28525, n28526, n28527, n28528, n28529, n28531,
         n28532, n28533, n28534, n28535, n28536, n28537, n28538, n28539,
         n28540, n28541, n28542, n28543, n28544, n28545, n28546, n28547,
         n28548, n28549, n28550, n28551, n28552, n28553, n28554, n28555,
         n28556, n28557, n28558, n28559, n28560, n28562, n28563, n28564,
         n28565, n28570, n28571, n28572, n28574, n28575, n28576, n28577,
         n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585,
         n28586, n28587, n28588, n28589, n28590, n28591, n28592, n28593,
         n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28602,
         n28603, n28604, n28605, n28606, n28607, n28608, n28609, n28610,
         n28611, n28612, n28613, n28614, n28615, n28616, n28617, n28618,
         n28619, n28620, n28621, n28622, n28623, n28624, n28625, n28626,
         n28627, n28628, n28629, n28630, n28631, n28632, n28633, n28634,
         n28635, n28636, n28638, n28639, n28640, n28642, n28643, n28644,
         n28645, n28646, n28647, n28648, n28649, n28650, n28651, n28652,
         n28653, n28654, n28655, n28656, n28657, n28658, n28659, n28660,
         n28661, n28662, n28663, n28664, n28665, n28666, n28667, n28668,
         n28669, n28670, n28671, n28672, n28673, n28674, n28675, n28676,
         n28677, n28678, n28679, n28681, n28682, n28683, n28684, n28685,
         n28686, n28687, n28688, n28689, n28690, n28691, n28692, n28693,
         n28694, n28695, n28696, n28697, n28698, n28699, n28701, n28702,
         n28703, n28704, n28705, n28706, n28707, n28710, n28711, n28712,
         n28713, n28714, n28715, n28716, n28717, n28720, n28721, n28722,
         n28723, n28725, n28726, n28727, n28728, n28730, n28731, n28732,
         n28733, n28734, n28735, n28736, n28737, n28738, n28739, n28740,
         n28743, n28744, n28745, n28746, n28748, n28749, n28750, n28751,
         n28752, n28753, n28754, n28755, n28756, n28757, n28758, n28760,
         n28761, n28762, n28763, n28764, n28768, n28769, n28770, n28771,
         n28772, n28773, n28774, n28775, n28776, n28777, n28778, n28779,
         n28780, n28781, n28782, n28783, n28784, n28785, n28786, n28787,
         n28788, n28789, n28790, n28791, n28792, n28793, n28794, n28795,
         n28796, n28797, n28798, n28799, n28800, n28801, n28802, n28803,
         n28804, n28805, n28806, n28807, n28808, n28809, n28810, n28811,
         n28812, n28813, n28814, n28815, n28816, n28817, n28818, n28819,
         n28820, n28821, n28823, n28824, n28825, n28826, n28827, n28828,
         n28829, n28830, n28831, n28832, n28833, n28834, n28835, n28836,
         n28837, n28838, n28839, n28840, n28841, n28842, n28843, n28844,
         n28845, n28846, n28847, n28848, n28850, n28851, n28852, n28853,
         n28854, n28855, n28856, n28857, n28858, n28859, n28860, n28861,
         n28862, n28863, n28864, n28865, n28866, n28867, n28868, n28869,
         n28870, n28871, n28872, n28873, n28874, n28875, n28876, n28877,
         n28878, n28879, n28880, n28881, n28882, n28883, n28884, n28885,
         n28886, n28887, n28888, n28889, n28890, n28891, n28892, n28893,
         n28894, n28895, n28896, n28897, n28898, n28899, n28900, n28901,
         n28902, n28903, n28904, n28905, n28907, n28908, n28909, n28911,
         n28912, n28913, n28914, n28915, n28916, n28917, n28918, n28919,
         n28920, n28921, n28922, n28923, n28924, n28925, n28926, n28927,
         n28928, n28929, n28930, n28931, n28932, n28933, n28934, n28935,
         n28937, n28938, n28939, n28940, n28941, n28942, n28943, n28944,
         n28945, n28947, n28948, n28949, n28950, n28951, n28952, n28953,
         n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961,
         n28962, n28964, n28965, n28966, n28969, n28970, n28971, n28972,
         n28973, n28974, n28975, n28976, n28977, n28978, n28979, n28980,
         n28981, n28982, n28983, n28984, n28985, n28986, n28987, n28988,
         n28989, n28990, n28991, n28992, n28993, n28994, n28995, n28996,
         n28997, n28999, n29000, n29001, n29002, n29003, n29004, n29007,
         n29008, n29009, n29010, n29011, n29012, n29013, n29014, n29015,
         n29016, n29017, n29018, n29019, n29020, n29021, n29022, n29024,
         n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033,
         n29034, n29035, n29036, n29037, n29038, n29039, n29040, n29041,
         n29043, n29045, n29047, n29050, n29051, n29052, n29053, n29054,
         n29055, n29056, n29057, n29058, n29059, n29060, n29061, n29062,
         n29063, n29064, n29065, n29066, n29067, n29068, n29069, n29070,
         n29071, n29072, n29073, n29074, n29075, n29076, n29077, n29078,
         n29079, n29080, n29083, n29084, n29085, n29086, n29087, n29088,
         n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29098,
         n29099, n29100, n29102, n29103, n29104, n29105, n29106, n29107,
         n29108, n29109, n29110, n29111, n29112, n29113, n29114, n29115,
         n29116, n29117, n29118, n29119, n29120, n29121, n29122, n29123,
         n29124, n29125, n29127, n29128, n29129, n29130, n29131, n29132,
         n29133, n29134, n29135, n29136, n29137, n29138, n29139, n29140,
         n29141, n29142, n29143, n29144, n29145, n29146, n29147, n29148,
         n29149, n29150, n29151, n29152, n29153, n29154, n29155, n29156,
         n29158, n29159, n29160, n29161, n29162, n29163, n29164, n29165,
         n29166, n29167, n29168, n29169, n29170, n29171, n29172, n29173,
         n29174, n29175, n29176, n29177, n29178, n29179, n29180, n29181,
         n29182, n29183, n29184, n29185, n29187, n29188, n29189, n29190,
         n29191, n29192, n29193, n29194, n29195, n29196, n29197, n29198,
         n29199, n29200, n29201, n29202, n29203, n29204, n29205, n29206,
         n29207, n29208, n29209, n29210, n29211, n29212, n29213, n29215,
         n29218, n29219, n29220, n29221, n29222, n29223, n29224, n29225,
         n29227, n29228, n29229, n29230, n29231, n29232, n29233, n29234,
         n29235, n29236, n29237, n29238, n29239, n29240, n29241, n29242,
         n29243, n29244, n29245, n29246, n29247, n29248, n29249, n29250,
         n29251, n29252, n29254, n29255, n29256, n29257, n29258, n29259,
         n29260, n29262, n29263, n29264, n29265, n29266, n29267, n29268,
         n29269, n29271, n29272, n29273, n29274, n29275, n29276, n29277,
         n29278, n29279, n29280, n29281, n29282, n29283, n29284, n29285,
         n29286, n29287, n29288, n29289, n29290, n29291, n29292, n29293,
         n29294, n29295, n29296, n29297, n29298, n29300, n29301, n29302,
         n29303, n29304, n29306, n29307, n29308, n29309, n29310, n29311,
         n29312, n29313, n29314, n29315, n29316, n29317, n29318, n29319,
         n29320, n29321, n29322, n29323, n29324, n29325, n29327, n29328,
         n29329, n29330, n29331, n29332, n29333, n29334, n29335, n29336,
         n29337, n29338, n29339, n29340, n29341, n29342, n29343, n29344,
         n29345, n29346, n29347, n29350, n29351, n29352, n29353, n29354,
         n29355, n29356, n29357, n29358, n29359, n29361, n29362, n29363,
         n29364, n29365, n29366, n29367, n29368, n29369, n29370, n29371,
         n29372, n29373, n29374, n29375, n29376, n29377, n29378, n29379,
         n29380, n29381, n29382, n29383, n29384, n29385, n29386, n29387,
         n29388, n29389, n29390, n29391, n29392, n29393, n29394, n29395,
         n29396, n29397, n29398, n29399, n29400, n29401, n29402, n29403,
         n29404, n29405, n29406, n29407, n29408, n29409, n29410, n29411,
         n29412, n29413, n29414, n29415, n29416, n29417, n29418, n29420,
         n29421, n29422, n29423, n29424, n29425, n29426, n29427, n29428,
         n29430, n29431, n29432, n29433, n29434, n29435, n29436, n29437,
         n29438, n29439, n29440, n29441, n29442, n29443, n29444, n29445,
         n29446, n29447, n29448, n29449, n29450, n29451, n29452, n29453,
         n29455, n29456, n29457, n29458, n29459, n29460, n29461, n29462,
         n29463, n29464, n29465, n29466, n29467, n29469, n29470, n29471,
         n29472, n29473, n29474, n29475, n29476, n29477, n29478, n29480,
         n29481, n29482, n29483, n29484, n29485, n29486, n29487, n29488,
         n29489, n29490, n29491, n29492, n29493, n29494, n29495, n29496,
         n29497, n29498, n29499, n29500, n29501, n29502, n29503, n29505,
         n29506, n29507, n29508, n29509, n29510, n29511, n29512, n29513,
         n29514, n29515, n29516, n29517, n29519, n29520, n29521, n29522,
         n29523, n29524, n29525, n29526, n29527, n29528, n29529, n29530,
         n29531, n29532, n29533, n29534, n29535, n29538, n29539, n29540,
         n29541, n29542, n29543, n29544, n29545, n29546, n29547, n29548,
         n29549, n29550, n29551, n29552, n29553, n29554, n29555, n29557,
         n29558, n29559, n29560, n29561, n29562, n29564, n29565, n29566,
         n29567, n29568, n29569, n29570, n29571, n29572, n29573, n29574,
         n29575, n29576, n29577, n29578, n29579, n29580, n29583, n29584,
         n29585, n29586, n29587, n29588, n29589, n29590, n29591, n29592,
         n29593, n29594, n29595, n29596, n29597, n29598, n29600, n29601,
         n29602, n29603, n29604, n29605, n29607, n29608, n29609, n29610,
         n29611, n29612, n29613, n29614, n29615, n29616, n29617, n29618,
         n29619, n29620, n29621, n29622, n29623, n29624, n29625, n29626,
         n29627, n29628, n29629, n29630, n29631, n29632, n29633, n29634,
         n29635, n29636, n29638, n29639, n29640, n29641, n29642, n29643,
         n29644, n29645, n29646, n29647, n29648, n29649, n29651, n29652,
         n29653, n29654, n29655, n29656, n29657, n29658, n29659, n29660,
         n29661, n29662, n29663, n29664, n29665, n29666, n29667, n29668,
         n29669, n29670, n29671, n29672, n29673, n29674, n29675, n29676,
         n29677, n29678, n29679, n29680, n29681, n29682, n29683, n29684,
         n29685, n29686, n29687, n29688, n29689, n29690, n29691, n29692,
         n29694, n29695, n29696, n29697, n29698, n29699, n29700, n29701,
         n29702, n29703, n29704, n29705, n29706, n29707, n29708, n29709,
         n29710, n29711, n29712, n29713, n29714, n29716, n29717, n29718,
         n29719, n29720, n29721, n29722, n29723, n29724, n29725, n29726,
         n29727, n29728, n29729, n29730, n29731, n29732, n29733, n29734,
         n29735, n29736, n29737, n29738, n29739, n29740, n29742, n29743,
         n29744, n29745, n29746, n29747, n29748, n29749, n29750, n29751,
         n29752, n29753, n29754, n29756, n29757, n29759, n29760, n29761,
         n29763, n29764, n29765, n29766, n29767, n29768, n29769, n29770,
         n29771, n29772, n29773, n29774, n29775, n29776, n29777, n29778,
         n29779, n29780, n29781, n29782, n29783, n29784, n29785, n29786,
         n29787, n29789, n29790, n29791, n29792, n29793, n29794, n29795,
         n29797, n29798, n29800, n29801, n29802, n29803, n29804, n29805,
         n29806, n29807, n29808, n29809, n29810, n29811, n29812, n29813,
         n29814, n29815, n29816, n29817, n29818, n29819, n29820, n29821,
         n29822, n29823, n29824, n29825, n29826, n29827, n29828, n29829,
         n29830, n29832, n29833, n29834, n29835, n29836, n29837, n29838,
         n29839, n29840, n29841, n29842, n29843, n29844, n29845, n29846,
         n29847, n29848, n29849, n29850, n29851, n29852, n29853, n29854,
         n29855, n29856, n29857, n29858, n29859, n29860, n29861, n29862,
         n29863, n29864, n29865, n29868, n29869, n29871, n29872, n29873,
         n29874, n29875, n29876, n29877, n29878, n29879, n29881, n29882,
         n29883, n29884, n29885, n29886, n29887, n29888, n29889, n29890,
         n29891, n29892, n29893, n29894, n29895, n29896, n29898, n29899,
         n29900, n29901, n29902, n29903, n29904, n29905, n29906, n29907,
         n29908, n29909, n29910, n29911, n29912, n29913, n29914, n29915,
         n29916, n29917, n29918, n29919, n29920, n29921, n29922, n29923,
         n29924, n29925, n29927, n29928, n29929, n29930, n29931, n29932,
         n29933, n29934, n29935, n29936, n29937, n29938, n29939, n29940,
         n29941, n29942, n29943, n29944, n29945, n29946, n29948, n29949,
         n29950, n29951, n29952, n29953, n29954, n29955, n29956, n29957,
         n29959, n29960, n29961, n29962, n29963, n29964, n29965, n29966,
         n29967, n29968, n29969, n29970, n29971, n29972, n29973, n29974,
         n29976, n29977, n29978, n29979, n29980, n29981, n29982, n29983,
         n29984, n29985, n29986, n29987, n29988, n29989, n29990, n29991,
         n29992, n29993, n29994, n29995, n29996, n29997, n29998, n29999,
         n30000, n30001, n30002, n30003, n30004, n30005, n30006, n30007,
         n30008, n30009, n30010, n30011, n30012, n30013, n30014, n30016,
         n30017, n30018, n30019, n30020, n30021, n30022, n30023, n30024,
         n30025, n30026, n30027, n30028, n30029, n30030, n30031, n30032,
         n30033, n30034, n30035, n30036, n30037, n30038, n30039, n30040,
         n30041, n30042, n30043, n30044, n30045, n30046, n30047, n30048,
         n30049, n30050, n30051, n30052, n30053, n30054, n30055, n30056,
         n30057, n30058, n30059, n30061, n30062, n30063, n30064, n30065,
         n30066, n30067, n30068, n30069, n30070, n30071, n30072, n30073,
         n30074, n30075, n30076, n30077, n30078, n30079, n30080, n30081,
         n30082, n30084, n30085, n30086, n30087, n30088, n30089, n30090,
         n30091, n30092, n30093, n30094, n30096, n30097, n30098, n30099,
         n30101, n30102, n30103, n30104, n30105, n30106, n30107, n30108,
         n30109, n30110, n30111, n30112, n30113, n30114, n30115, n30116,
         n30117, n30118, n30119, n30120, n30121, n30122, n30123, n30124,
         n30125, n30126, n30127, n30128, n30129, n30130, n30131, n30132,
         n30133, n30134, n30135, n30136, n30137, n30138, n30139, n30140,
         n30141, n30142, n30143, n30144, n30145, n30146, n30147, n30148,
         n30149, n30150, n30151, n30152, n30153, n30154, n30155, n30156,
         n30157, n30158, n30159, n30160, n30161, n30162, n30163, n30164,
         n30165, n30166, n30167, n30168, n30169, n30170, n30172, n30173,
         n30174, n30175, n30176, n30177, n30178, n30179, n30180, n30181,
         n30182, n30183, n30184, n30185, n30187, n30188, n30189, n30190,
         n30192, n30193, n30194, n30195, n30196, n30197, n30198, n30199,
         n30200, n30201, n30205, n30206, n30207, n30209, n30210, n30211,
         n30212, n30213, n30214, n30215, n30216, n30217, n30218, n30219,
         n30220, n30221, n30222, n30223, n30224, n30225, n30226, n30227,
         n30228, n30229, n30230, n30231, n30232, n30233, n30234, n30235,
         n30236, n30237, n30238, n30239, n30240, n30241, n30242, n30243,
         n30244, n30245, n30246, n30247, n30248, n30250, n30251, n30252,
         n30253, n30254, n30255, n30258, n30259, n30260, n30261, n30262,
         n30263, n30264, n30265, n30266, n30267, n30268, n30269, n30271,
         n30273, n30274, n30275, n30276, n30277, n30278, n30279, n30280,
         n30281, n30282, n30283, n30284, n30285, n30286, n30288, n30291,
         n30292, n30293, n30294, n30295, n30296, n30297, n30298, n30299,
         n30300, n30301, n30302, n30303, n30304, n30305, n30306, n30307,
         n30308, n30309, n30310, n30311, n30312, n30313, n30314, n30316,
         n30317, n30318, n30319, n30320, n30321, n30322, n30323, n30324,
         n30325, n30326, n30327, n30328, n30329, n30330, n30331, n30332,
         n30333, n30334, n30335, n30336, n30337, n30338, n30339, n30340,
         n30341, n30342, n30343, n30344, n30345, n30347, n30348, n30349,
         n30350, n30351, n30352, n30354, n30355, n30356, n30358, n30359,
         n30360, n30361, n30362, n30363, n30364, n30365, n30367, n30368,
         n30369, n30370, n30371, n30372, n30373, n30374, n30375, n30376,
         n30377, n30378, n30379, n30380, n30381, n30382, n30383, n30384,
         n30385, n30386, n30387, n30388, n30389, n30390, n30391, n30392,
         n30393, n30394, n30395, n30396, n30397, n30398, n30399, n30400,
         n30401, n30402, n30403, n30404, n30405, n30406, n30407, n30408,
         n30409, n30410, n30411, n30412, n30413, n30414, n30415, n30416,
         n30417, n30418, n30419, n30421, n30422, n30423, n30424, n30425,
         n30427, n30429, n30430, n30431, n30432, n30433, n30434, n30435,
         n30436, n30437, n30438, n30439, n30440, n30441, n30442, n30443,
         n30444, n30445, n30446, n30447, n30448, n30449, n30450, n30451,
         n30452, n30454, n30455, n30456, n30457, n30458, n30459, n30460,
         n30461, n30462, n30463, n30465, n30466, n30467, n30468, n30469,
         n30470, n30471, n30472, n30473, n30474, n30475, n30476, n30477,
         n30478, n30479, n30480, n30481, n30482, n30483, n30484, n30486,
         n30487, n30488, n30489, n30490, n30491, n30492, n30493, n30494,
         n30495, n30496, n30497, n30498, n30499, n30500, n30501, n30502,
         n30504, n30505, n30506, n30507, n30508, n30509, n30510, n30511,
         n30513, n30514, n30517, n30518, n30519, n30520, n30521, n30522,
         n30523, n30524, n30525, n30526, n30527, n30528, n30529, n30530,
         n30531, n30532, n30533, n30534, n30535, n30536, n30537, n30538,
         n30540, n30541, n30543, n30544, n30545, n30546, n30547, n30548,
         n30549, n30550, n30551, n30552, n30553, n30554, n30555, n30556,
         n30557, n30558, n30559, n30560, n30561, n30562, n30563, n30564,
         n30565, n30566, n30567, n30568, n30569, n30570, n30571, n30573,
         n30574, n30575, n30576, n30577, n30578, n30579, n30580, n30581,
         n30582, n30583, n30584, n30585, n30586, n30587, n30588, n30589,
         n30590, n30591, n30592, n30593, n30594, n30595, n30596, n30597,
         n30598, n30599, n30601, n30602, n30603, n30604, n30606, n30607,
         n30608, n30609, n30610, n30613, n30614, n30616, n30617, n30618,
         n30619, n30620, n30621, n30622, n30623, n30624, n30625, n30626,
         n30627, n30628, n30629, n30630, n30631, n30632, n30633, n30634,
         n30635, n30636, n30637, n30638, n30639, n30640, n30641, n30642,
         n30643, n30645, n30646, n30647, n30648, n30649, n30650, n30651,
         n30653, n30654, n30655, n30656, n30657, n30658, n30659, n30660,
         n30661, n30662, n30663, n30664, n30665, n30666, n30667, n30668,
         n30669, n30670, n30671, n30672, n30673, n30675, n30676, n30677,
         n30678, n30679, n30680, n30681, n30682, n30683, n30684, n30685,
         n30686, n30687, n30688, n30689, n30691, n30692, n30693, n30695,
         n30696, n30697, n30698, n30699, n30700, n30701, n30702, n30703,
         n30704, n30705, n30706, n30707, n30708, n30709, n30710, n30711,
         n30712, n30713, n30714, n30715, n30716, n30717, n30718, n30719,
         n30720, n30721, n30722, n30723, n30724, n30725, n30726, n30727,
         n30728, n30729, n30730, n30731, n30733, n30735, n30736, n30737,
         n30738, n30739, n30740, n30741, n30742, n30743, n30744, n30745,
         n30746, n30747, n30748, n30749, n30750, n30751, n30752, n30753,
         n30754, n30755, n30757, n30758, n30759, n30760, n30761, n30762,
         n30763, n30764, n30765, n30766, n30767, n30768, n30769, n30770,
         n30771, n30772, n30773, n30774, n30775, n30776, n30777, n30778,
         n30779, n30780, n30781, n30782, n30783, n30784, n30785, n30786,
         n30787, n30788, n30789, n30790, n30791, n30792, n30793, n30794,
         n30795, n30796, n30797, n30798, n30799, n30801, n30802, n30803,
         n30804, n30805, n30806, n30807, n30808, n30809, n30810, n30811,
         n30812, n30813, n30814, n30815, n30816, n30817, n30818, n30819,
         n30820, n30822, n30823, n30824, n30825, n30826, n30827, n30828,
         n30829, n30830, n30831, n30832, n30833, n30834, n30835, n30836,
         n30837, n30838, n30839, n30840, n30841, n30842, n30843, n30844,
         n30845, n30846, n30848, n30849, n30850, n30851, n30852, n30853,
         n30854, n30855, n30856, n30857, n30858, n30859, n30860, n30861,
         n30862, n30863, n30864, n30865, n30866, n30867, n30869, n30870,
         n30871, n30873, n30874, n30875, n30876, n30877, n30878, n30881,
         n30882, n30883, n30884, n30885, n30886, n30887, n30888, n30889,
         n30890, n30891, n30892, n30893, n30894, n30895, n30896, n30897,
         n30898, n30899, n30900, n30901, n30903, n30904, n30906, n30907,
         n30908, n30909, n30910, n30911, n30912, n30913, n30914, n30915,
         n30916, n30917, n30918, n30919, n30920, n30921, n30922, n30924,
         n30925, n30926, n30927, n30928, n30929, n30930, n30931, n30932,
         n30933, n30934, n30935, n30936, n30937, n30938, n30939, n30940,
         n30941, n30943, n30944, n30945, n30946, n30947, n30948, n30949,
         n30950, n30951, n30952, n30953, n30954, n30955, n30956, n30957,
         n30958, n30959, n30960, n30961, n30962, n30963, n30964, n30965,
         n30967, n30968, n30969, n30970, n30971, n30972, n30973, n30974,
         n30975, n30976, n30977, n30979, n30980, n30981, n30982, n30983,
         n30984, n30985, n30986, n30987, n30988, n30989, n30990, n30992,
         n30993, n30994, n30995, n30996, n30998, n30999, n31000, n31001,
         n31002, n31003, n31004, n31005, n31006, n31007, n31008, n31009,
         n31010, n31011, n31012, n31013, n31014, n31015, n31016, n31017,
         n31018, n31019, n31020, n31022, n31023, n31024, n31025, n31026,
         n31027, n31028, n31029, n31030, n31031, n31032, n31033, n31034,
         n31035, n31036, n31037, n31038, n31039, n31040, n31041, n31042,
         n31043, n31044, n31045, n31046, n31047, n31048, n31049, n31050,
         n31051, n31052, n31053, n31054, n31055, n31056, n31057, n31058,
         n31059, n31060, n31061, n31062, n31063, n31065, n31066, n31068,
         n31069, n31070, n31071, n31072, n31073, n31074, n31075, n31076,
         n31077, n31079, n31080, n31081, n31082, n31083, n31084, n31085,
         n31086, n31088, n31089, n31090, n31091, n31092, n31093, n31094,
         n31095, n31096, n31097, n31098, n31099, n31100, n31101, n31102,
         n31104, n31105, n31106, n31107, n31108, n31109, n31110, n31111,
         n31112, n31113, n31114, n31115, n31116, n31117, n31118, n31119,
         n31120, n31121, n31122, n31123, n31124, n31125, n31126, n31127,
         n31128, n31129, n31131, n31132, n31133, n31134, n31135, n31136,
         n31137, n31138, n31139, n31140, n31141, n31142, n31143, n31144,
         n31145, n31146, n31147, n31148, n31149, n31150, n31151, n31152,
         n31153, n31154, n31155, n31156, n31159, n31160, n31161, n31162,
         n31163, n31164, n31165, n31166, n31167, n31168, n31169, n31170,
         n31171, n31173, n31174, n31175, n31176, n31177, n31178, n31179,
         n31182, n31183, n31184, n31185, n31187, n31188, n31189, n31190,
         n31191, n31192, n31193, n31194, n31195, n31196, n31197, n31198,
         n31199, n31200, n31201, n31202, n31203, n31204, n31205, n31206,
         n31207, n31208, n31209, n31210, n31211, n31212, n31213, n31214,
         n31215, n31216, n31217, n31218, n31219, n31220, n31221, n31222,
         n31223, n31224, n31225, n31226, n31227, n31228, n31229, n31230,
         n31231, n31232, n31233, n31234, n31236, n31237, n31238, n31239,
         n31240, n31241, n31242, n31243, n31244, n31245, n31246, n31247,
         n31248, n31249, n31250, n31251, n31252, n31253, n31254, n31255,
         n31256, n31257, n31258, n31259, n31260, n31261, n31262, n31263,
         n31264, n31265, n31266, n31267, n31268, n31269, n31270, n31271,
         n31272, n31273, n31274, n31275, n31276, n31277, n31278, n31279,
         n31280, n31281, n31282, n31284, n31285, n31286, n31287, n31288,
         n31289, n31290, n31291, n31292, n31293, n31294, n31296, n31297,
         n31298, n31299, n31300, n31301, n31302, n31303, n31305, n31306,
         n31307, n31308, n31309, n31310, n31311, n31312, n31313, n31314,
         n31315, n31316, n31317, n31318, n31319, n31320, n31321, n31322,
         n31323, n31324, n31325, n31326, n31327, n31329, n31330, n31331,
         n31332, n31333, n31334, n31335, n31336, n31338, n31339, n31340,
         n31341, n31342, n31344, n31345, n31346, n31347, n31348, n31349,
         n31350, n31351, n31354, n31355, n31356, n31357, n31358, n31359,
         n31360, n31361, n31362, n31365, n31366, n31367, n31368, n31369,
         n31370, n31371, n31372, n31373, n31374, n31375, n31376, n31377,
         n31378, n31379, n31380, n31381, n31382, n31383, n31384, n31385,
         n31386, n31387, n31388, n31389, n31390, n31391, n31392, n31393,
         n31394, n31395, n31397, n31398, n31399, n31401, n31403, n31404,
         n31405, n31406, n31407, n31408, n31409, n31410, n31411, n31412,
         n31413, n31414, n31417, n31418, n31419, n31420, n31421, n31422,
         n31423, n31424, n31425, n31426, n31427, n31428, n31429, n31430,
         n31431, n31432, n31433, n31434, n31435, n31436, n31437, n31438,
         n31439, n31440, n31442, n31444, n31445, n31446, n31447, n31448,
         n31449, n31450, n31452, n31453, n31454, n31455, n31456, n31458,
         n31459, n31460, n31461, n31463, n31464, n31465, n31466, n31468,
         n31469, n31470, n31472, n31473, n31474, n31475, n31476, n31477,
         n31479, n31480, n31481, n31482, n31483, n31484, n31485, n31486,
         n31487, n31489, n31490, n31491, n31492, n31493, n31494, n31495,
         n31496, n31497, n31498, n31499, n31502, n31503, n31504, n31505,
         n31506, n31507, n31508, n31509, n31510, n31511, n31512, n31513,
         n31514, n31515, n31516, n31517, n31518, n31519, n31520, n31521,
         n31522, n31523, n31524, n31525, n31526, n31528, n31529, n31530,
         n31531, n31532, n31533, n31534, n31535, n31536, n31537, n31538,
         n31539, n31540, n31541, n31542, n31543, n31544, n31545, n31546,
         n31547, n31548, n31549, n31550, n31551, n31552, n31553, n31554,
         n31555, n31556, n31558, n31559, n31560, n31561, n31562, n31563,
         n31565, n31566, n31568, n31569, n31570, n31571, n31572, n31573,
         n31574, n31575, n31576, n31577, n31579, n31581, n31582, n31583,
         n31584, n31585, n31587, n31588, n31589, n31590, n31591, n31592,
         n31593, n31594, n31595, n31597, n31598, n31599, n31600, n31601,
         n31602, n31603, n31604, n31605, n31606, n31607, n31608, n31609,
         n31610, n31611, n31612, n31613, n31614, n31615, n31616, n31617,
         n31618, n31619, n31622, n31623, n31624, n31625, n31626, n31627,
         n31628, n31629, n31630, n31632, n31633, n31634, n31635, n31637,
         n31638, n31639, n31640, n31641, n31642, n31643, n31644, n31645,
         n31646, n31647, n31648, n31649, n31650, n31651, n31653, n31654,
         n31655, n31656, n31657, n31658, n31659, n31660, n31661, n31663,
         n31664, n31665, n31666, n31667, n31668, n31669, n31670, n31671,
         n31672, n31673, n31674, n31675, n31676, n31677, n31678, n31679,
         n31680, n31681, n31682, n31683, n31684, n31685, n31686, n31687,
         n31688, n31689, n31690, n31691, n31692, n31693, n31694, n31695,
         n31696, n31697, n31698, n31699, n31700, n31701, n31702, n31703,
         n31704, n31705, n31706, n31707, n31708, n31709, n31710, n31711,
         n31712, n31713, n31714, n31715, n31716, n31718, n31719, n31720,
         n31721, n31722, n31724, n31725, n31727, n31728, n31729, n31730,
         n31731, n31732, n31734, n31735, n31736, n31737, n31738, n31739,
         n31740, n31741, n31742, n31743, n31744, n31745, n31746, n31747,
         n31748, n31749, n31750, n31751, n31752, n31753, n31754, n31755,
         n31756, n31757, n31758, n31759, n31760, n31761, n31762, n31763,
         n31764, n31765, n31766, n31767, n31768, n31769, n31770, n31771,
         n31772, n31773, n31774, n31775, n31776, n31777, n31778, n31779,
         n31780, n31781, n31782, n31783, n31784, n31785, n31786, n31787,
         n31788, n31789, n31791, n31792, n31793, n31794, n31795, n31796,
         n31797, n31798, n31799, n31800, n31801, n31802, n31803, n31804,
         n31805, n31806, n31808, n31809, n31810, n31811, n31812, n31813,
         n31814, n31815, n31816, n31817, n31818, n31819, n31820, n31821,
         n31823, n31824, n31825, n31826, n31827, n31828, n31830, n31831,
         n31832, n31833, n31834, n31835, n31836, n31837, n31838, n31839,
         n31840, n31841, n31842, n31843, n31844, n31845, n31846, n31847,
         n31848, n31849, n31850, n31851, n31852, n31853, n31854, n31855,
         n31856, n31857, n31858, n31859, n31860, n31861, n31862, n31863,
         n31864, n31865, n31866, n31867, n31868, n31869, n31870, n31871,
         n31872, n31873, n31874, n31875, n31876, n31877, n31878, n31879,
         n31880, n31881, n31882, n31883, n31884, n31885, n31886, n31887,
         n31888, n31889, n31890, n31892, n31893, n31894, n31895, n31896,
         n31897, n31898, n31899, n31900, n31901, n31902, n31905, n31906,
         n31907, n31908, n31909, n31910, n31911, n31912, n31913, n31914,
         n31915, n31916, n31917, n31918, n31919, n31920, n31921, n31922,
         n31923, n31924, n31925, n31926, n31927, n31928, n31929, n31930,
         n31931, n31932, n31933, n31935, n31936, n31937, n31938, n31939,
         n31940, n31941, n31943, n31944, n31945, n31946, n31947, n31948,
         n31950, n31951, n31952, n31953, n31954, n31955, n31956, n31957,
         n31958, n31959, n31960, n31961, n31962, n31964, n31965, n31966,
         n31967, n31968, n31969, n31970, n31971, n31972, n31973, n31974,
         n31975, n31976, n31977, n31978, n31979, n31980, n31981, n31982,
         n31983, n31984, n31985, n31986, n31987, n31988, n31989, n31990,
         n31991, n31992, n31993, n31994, n31995, n31996, n31997, n31998,
         n31999, n32000, n32001, n32002, n32003, n32004, n32005, n32006,
         n32007, n32008, n32009, n32010, n32011, n32012, n32013, n32014,
         n32015, n32016, n32017, n32018, n32019, n32020, n32021, n32022,
         n32023, n32024, n32025, n32026, n32027, n32028, n32029, n32030,
         n32031, n32032, n32033, n32034, n32035, n32036, n32037, n32038,
         n32039, n32040, n32041, n32042, n32043, n32044, n32045, n32046,
         n32047, n32048, n32049, n32051, n32052, n32053, n32054, n32055,
         n32056, n32057, n32058, n32059, n32060, n32061, n32062, n32063,
         n32064, n32065, n32066, n32067, n32068, n32069, n32070, n32071,
         n32072, n32073, n32074, n32075, n32076, n32077, n32078, n32079,
         n32080, n32081, n32082, n32083, n32084, n32085, n32086, n32087,
         n32088, n32089, n32090, n32091, n32092, n32093, n32094, n32095,
         n32096, n32097, n32098, n32099, n32100, n32101, n32102, n32103,
         n32104, n32105, n32106, n32107, n32108, n32109, n32110, n32111,
         n32112, n32113, n32114, n32115, n32116, n32117, n32118, n32119,
         n32120, n32121, n32122, n32123, n32124, n32125, n32126, n32127,
         n32128, n32129, n32130, n32132, n32133, n32134, n32135, n32136,
         n32137, n32138, n32139, n32140, n32141, n32142, n32143, n32144,
         n32145, n32148, n32149, n32150, n32153, n32154, n32155, n32156,
         n32157, n32158, n32159, n32160, n32161, n32162, n32163, n32164,
         n32165, n32166, n32167, n32168, n32169, n32170, n32171, n32172,
         n32173, n32174, n32175, n32176, n32177, n32178, n32179, n32180,
         n32181, n32182, n32183, n32184, n32185, n32186, n32187, n32188,
         n32189, n32190, n32191, n32192, n32193, n32194, n32196, n32199,
         n32200, n32201, n32202, n32203, n32204, n32205, n32206, n32207,
         n32208, n32210, n32211, n32212, n32213, n32214, n32215, n32216,
         n32217, n32218, n32219, n32220, n32221, n32222, n32223, n32224,
         n32226, n32227, n32228, n32229, n32230, n32231, n32232, n32233,
         n32234, n32235, n32236, n32237, n32238, n32239, n32241, n32242,
         n32243, n32244, n32246, n32247, n32248, n32249, n32250, n32251,
         n32252, n32253, n32255, n32256, n32257, n32258, n32259, n32260,
         n32261, n32262, n32263, n32264, n32265, n32266, n32267, n32268,
         n32269, n32270, n32271, n32272, n32273, n32274, n32275, n32276,
         n32278, n32279, n32280, n32281, n32282, n32283, n32284, n32285,
         n32286, n32287, n32288, n32289, n32290, n32291, n32292, n32293,
         n32294, n32295, n32296, n32297, n32298, n32299, n32300, n32301,
         n32302, n32303, n32304, n32305, n32306, n32307, n32308, n32309,
         n32310, n32311, n32312, n32313, n32314, n32315, n32316, n32317,
         n32318, n32319, n32320, n32321, n32322, n32323, n32324, n32325,
         n32326, n32327, n32328, n32329, n32330, n32331, n32332, n32333,
         n32334, n32335, n32336, n32337, n32338, n32339, n32340, n32341,
         n32342, n32343, n32344, n32345, n32346, n32348, n32349, n32350,
         n32351, n32352, n32353, n32354, n32355, n32356, n32357, n32358,
         n32359, n32360, n32361, n32363, n32364, n32365, n32366, n32367,
         n32368, n32369, n32370, n32371, n32372, n32373, n32374, n32375,
         n32376, n32377, n32378, n32379, n32380, n32381, n32382, n32383,
         n32384, n32385, n32386, n32387, n32388, n32389, n32390, n32391,
         n32392, n32393, n32394, n32395, n32396, n32397, n32398, n32399,
         n32400, n32401, n32402, n32403, n32405, n32406, n32407, n32408,
         n32409, n32410, n32411, n32412, n32413, n32414, n32415, n32416,
         n32417, n32418, n32420, n32421, n32422, n32423, n32424, n32425,
         n32426, n32427, n32428, n32429, n32430, n32431, n32432, n32435,
         n32436, n32437, n32438, n32439, n32440, n32441, n32442, n32443,
         n32444, n32445, n32446, n32447, n32448, n32449, n32450, n32451,
         n32452, n32453, n32454, n32455, n32456, n32457, n32458, n32459,
         n32460, n32461, n32462, n32463, n32464, n32465, n32466, n32467,
         n32468, n32469, n32470, n32471, n32472, n32473, n32474, n32475,
         n32476, n32479, n32481, n32482, n32483, n32484, n32485, n32486,
         n32487, n32488, n32489, n32490, n32491, n32492, n32493, n32494,
         n32495, n32496, n32497, n32498, n32499, n32500, n32501, n32502,
         n32503, n32504, n32505, n32506, n32507, n32508, n32509, n32510,
         n32511, n32512, n32513, n32514, n32515, n32516, n32517, n32519,
         n32520, n32521, n32522, n32523, n32524, n32525, n32526, n32527,
         n32528, n32529, n32530, n32531, n32532, n32533, n32534, n32535,
         n32536, n32537, n32538, n32539, n32540, n32541, n32542, n32543,
         n32544, n32545, n32546, n32547, n32548, n32549, n32550, n32551,
         n32552, n32553, n32554, n32556, n32557, n32558, n32559, n32560,
         n32561, n32562, n32563, n32564, n32565, n32566, n32567, n32568,
         n32569, n32570, n32571, n32572, n32573, n32574, n32575, n32576,
         n32577, n32578, n32579, n32580, n32581, n32582, n32583, n32584,
         n32585, n32586, n32587, n32588, n32589, n32590, n32591, n32592,
         n32593, n32594, n32595, n32596, n32598, n32599, n32600, n32601,
         n32602, n32604, n32605, n32606, n32608, n32609, n32610, n32611,
         n32612, n32613, n32614, n32615, n32616, n32617, n32618, n32619,
         n32620, n32621, n32622, n32623, n32624, n32625, n32626, n32627,
         n32628, n32629, n32630, n32631, n32632, n32633, n32634, n32635,
         n32636, n32637, n32638, n32639, n32640, n32641, n32642, n32643,
         n32644, n32645, n32646, n32648, n32649, n32650, n32653, n32654,
         n32655, n32657, n32658, n32659, n32660, n32661, n32662, n32663,
         n32664, n32665, n32666, n32667, n32668, n32669, n32670, n32671,
         n32672, n32673, n32674, n32675, n32676, n32677, n32678, n32679,
         n32680, n32681, n32682, n32684, n32685, n32686, n32687, n32688,
         n32689, n32690, n32691, n32692, n32694, n32695, n32696, n32697,
         n32699, n32700, n32702, n32703, n32704, n32706, n32707, n32708,
         n32709, n32710, n32711, n32712, n32713, n32714, n32715, n32716,
         n32717, n32718, n32719, n32720, n32721, n32722, n32723, n32724,
         n32725, n32726, n32728, n32729, n32730, n32731, n32732, n32733,
         n32734, n32735, n32736, n32737, n32738, n32739, n32740, n32741,
         n32742, n32743, n32744, n32745, n32746, n32747, n32748, n32749,
         n32750, n32751, n32752, n32753, n32754, n32755, n32756, n32757,
         n32758, n32760, n32763, n32764, n32765, n32766, n32767, n32768,
         n32769, n32770, n32771, n32772, n32773, n32774, n32775, n32776,
         n32777, n32778, n32779, n32780, n32781, n32782, n32784, n32785,
         n32786, n32787, n32788, n32789, n32790, n32791, n32792, n32793,
         n32794, n32795, n32796, n32797, n32798, n32799, n32800, n32801,
         n32802, n32803, n32804, n32805, n32806, n32807, n32808, n32809,
         n32810, n32811, n32812, n32813, n32814, n32815, n32816, n32819,
         n32820, n32821, n32822, n32823, n32824, n32827, n32828, n32829,
         n32831, n32832, n32833, n32834, n32835, n32836, n32837, n32838,
         n32839, n32840, n32841, n32842, n32843, n32844, n32845, n32846,
         n32847, n32848, n32849, n32850, n32851, n32852, n32853, n32854,
         n32855, n32856, n32857, n32858, n32859, n32860, n32861, n32862,
         n32864, n32865, n32867, n32868, n32869, n32870, n32871, n32872,
         n32875, n32878, n32879, n32880, n32882, n32883, n32884, n32885,
         n32886, n32887, n32889, n32890, n32891, n32892, n32893, n32895,
         n32896, n32897, n32898, n32899, n32900, n32901, n32902, n32903,
         n32904, n32905, n32906, n32907, n32908, n32910, n32911, n32912,
         n32913, n32914, n32915, n32916, n32917, n32918, n32919, n32920,
         n32921, n32922, n32923, n32924, n32925, n32926, n32927, n32928,
         n32929, n32930, n32931, n32932, n32933, n32934, n32936, n32937,
         n32938, n32939, n32940, n32941, n32942, n32943, n32944, n32945,
         n32946, n32947, n32948, n32949, n32950, n32951, n32952, n32953,
         n32955, n32956, n32958, n32959, n32961, n32963, n32964, n32965,
         n32966, n32967, n32968, n32969, n32970, n32971, n32972, n32973,
         n32974, n32975, n32976, n32977, n32978, n32979, n32981, n32982,
         n32984, n32985, n32986, n32987, n32988, n32989, n32990, n32991,
         n32992, n32993, n32994, n32995, n32996, n32997, n32998, n32999,
         n33000, n33001, n33002, n33003, n33004, n33005, n33006, n33007,
         n33010, n33011, n33012, n33013, n33014, n33015, n33016, n33017,
         n33018, n33019, n33021, n33022, n33023, n33024, n33025, n33026,
         n33027, n33028, n33029, n33030, n33031, n33032, n33033, n33034,
         n33035, n33036, n33037, n33038, n33039, n33040, n33041, n33042,
         n33043, n33044, n33045, n33046, n33047, n33048, n33049, n33050,
         n33051, n33052, n33053, n33054, n33055, n33056, n33057, n33058,
         n33059, n33060, n33061, n33062, n33063, n33064, n33065, n33067,
         n33068, n33069, n33070, n33071, n33072, n33073, n33074, n33075,
         n33076, n33077, n33079, n33081, n33083, n33084, n33085, n33086,
         n33087, n33088, n33089, n33092, n33094, n33095, n33096, n33097,
         n33098, n33099, n33100, n33101, n33103, n33104, n33105, n33107,
         n33108, n33109, n33110, n33111, n33112, n33115, n33116, n33117,
         n33118, n33119, n33121, n33122, n33124, n33125, n33126, n33127,
         n33128, n33129, n33130, n33131, n33132, n33133, n33134, n33135,
         n33136, n33137, n33138, n33139, n33140, n33141, n33142, n33143,
         n33144, n33145, n33146, n33147, n33148, n33149, n33150, n33151,
         n33152, n33153, n33154, n33155, n33156, n33157, n33158, n33159,
         n33160, n33161, n33162, n33163, n33164, n33165, n33166, n33167,
         n33168, n33169, n33170, n33171, n33172, n33173, n33174, n33175,
         n33176, n33177, n33178, n33179, n33180, n33181, n33182, n33183,
         n33184, n33185, n33186, n33187, n33188, n33189, n33190, n33191,
         n33192, n33193, n33194, n33195, n33196, n33197, n33198, n33199,
         n33200, n33201, n33202, n33203, n33204, n33205, n33206, n33207,
         n33208, n33209, n33210, n33212, n33213, n33214, n33215, n33216,
         n33219, n33220, n33221, n33222, n33223, n33224, n33226, n33227,
         n33228, n33229, n33230, n33231, n33232, n33233, n33234, n33235,
         n33236, n33237, n33238, n33239, n33240, n33242, n33243, n33244,
         n33245, n33246, n33247, n33248, n33249, n33250, n33251, n33252,
         n33253, n33254, n33255, n33256, n33257, n33258, n33259, n33260,
         n33261, n33262, n33263, n33264, n33265, n33266, n33267, n33268,
         n33269, n33270, n33271, n33272, n33273, n33274, n33275, n33276,
         n33277, n33278, n33279, n33280, n33281, n33282, n33283, n33284,
         n33285, n33286, n33287, n33288, n33289, n33291, n33292, n33293,
         n33294, n33295, n33296, n33297, n33298, n33299, n33300, n33301,
         n33302, n33303, n33304, n33305, n33306, n33307, n33308, n33309,
         n33310, n33311, n33312, n33314, n33315, n33316, n33317, n33319,
         n33320, n33321, n33322, n33323, n33324, n33326, n33327, n33328,
         n33329, n33330, n33332, n33333, n33334, n33335, n33336, n33337,
         n33338, n33339, n33341, n33342, n33344, n33345, n33347, n33348,
         n33349, n33350, n33351, n33352, n33353, n33354, n33355, n33356,
         n33357, n33358, n33359, n33360, n33361, n33362, n33364, n33367,
         n33368, n33369, n33370, n33371, n33372, n33374, n33375, n33376,
         n33377, n33378, n33379, n33380, n33381, n33384, n33385, n33386,
         n33387, n33388, n33389, n33390, n33391, n33393, n33394, n33395,
         n33396, n33397, n33398, n33399, n33400, n33401, n33402, n33403,
         n33404, n33405, n33406, n33407, n33408, n33409, n33410, n33411,
         n33412, n33413, n33414, n33415, n33417, n33418, n33419, n33420,
         n33421, n33422, n33423, n33424, n33425, n33426, n33427, n33428,
         n33429, n33430, n33431, n33432, n33433, n33434, n33435, n33436,
         n33437, n33438, n33439, n33440, n33441, n33442, n33443, n33445,
         n33446, n33447, n33448, n33449, n33450, n33451, n33453, n33454,
         n33455, n33456, n33457, n33458, n33459, n33460, n33462, n33463,
         n33464, n33465, n33466, n33467, n33468, n33469, n33470, n33471,
         n33474, n33475, n33476, n33477, n33478, n33479, n33480, n33481,
         n33482, n33483, n33484, n33485, n33486, n33487, n33488, n33489,
         n33490, n33492, n33493, n33494, n33495, n33496, n33497, n33498,
         n33499, n33500, n33501, n33502, n33503, n33504, n33505, n33506,
         n33507, n33508, n33509, n33510, n33511, n33512, n33513, n33514,
         n33515, n33517, n33518, n33519, n33520, n33521, n33522, n33523,
         n33524, n33525, n33526, n33527, n33528, n33529, n33530, n33531,
         n33532, n33533, n33534, n33535, n33536, n33537, n33538, n33539,
         n33540, n33541, n33542, n33543, n33544, n33545, n33546, n33547,
         n33548, n33549, n33550, n33551, n33552, n33553, n33554, n33555,
         n33556, n33557, n33558, n33559, n33560, n33561, n33562, n33563,
         n33564, n33565, n33566, n33567, n33568, n33570, n33571, n33573,
         n33574, n33575, n33576, n33577, n33578, n33579, n33580, n33581,
         n33582, n33583, n33584, n33585, n33587, n33588, n33589, n33590,
         n33592, n33593, n33594, n33595, n33596, n33597, n33598, n33599,
         n33600, n33601, n33602, n33603, n33606, n33607, n33608, n33609,
         n33610, n33611, n33612, n33613, n33614, n33615, n33616, n33617,
         n33618, n33619, n33620, n33621, n33622, n33623, n33624, n33625,
         n33626, n33627, n33628, n33629, n33630, n33631, n33632, n33633,
         n33634, n33635, n33637, n33638, n33639, n33640, n33641, n33642,
         n33643, n33644, n33645, n33647, n33648, n33649, n33650, n33651,
         n33652, n33653, n33654, n33655, n33656, n33657, n33658, n33660,
         n33661, n33662, n33663, n33664, n33666, n33668, n33669, n33670,
         n33672, n33673, n33674, n33675, n33676, n33677, n33678, n33679,
         n33680, n33681, n33682, n33683, n33684, n33685, n33686, n33687,
         n33689, n33690, n33691, n33692, n33693, n33694, n33695, n33696,
         n33697, n33698, n33699, n33700, n33701, n33702, n33703, n33704,
         n33705, n33706, n33707, n33708, n33709, n33710, n33713, n33714,
         n33715, n33716, n33717, n33718, n33719, n33720, n33721, n33722,
         n33723, n33724, n33725, n33726, n33728, n33729, n33730, n33731,
         n33732, n33733, n33734, n33735, n33736, n33737, n33738, n33739,
         n33740, n33741, n33742, n33743, n33744, n33745, n33746, n33747,
         n33748, n33749, n33750, n33751, n33752, n33753, n33754, n33756,
         n33757, n33758, n33759, n33760, n33761, n33762, n33763, n33764,
         n33765, n33766, n33767, n33770, n33771, n33773, n33774, n33775,
         n33776, n33777, n33778, n33779, n33780, n33781, n33782, n33783,
         n33784, n33785, n33786, n33787, n33788, n33789, n33790, n33791,
         n33793, n33794, n33795, n33796, n33797, n33798, n33799, n33800,
         n33801, n33802, n33803, n33804, n33807, n33808, n33809, n33810,
         n33811, n33812, n33813, n33814, n33815, n33816, n33817, n33818,
         n33819, n33820, n33821, n33823, n33824, n33825, n33826, n33827,
         n33828, n33829, n33830, n33831, n33832, n33833, n33834, n33835,
         n33836, n33837, n33838, n33839, n33840, n33841, n33842, n33843,
         n33844, n33845, n33846, n33847, n33848, n33849, n33850, n33851,
         n33852, n33853, n33854, n33855, n33856, n33857, n33858, n33859,
         n33860, n33861, n33862, n33863, n33864, n33865, n33866, n33867,
         n33868, n33869, n33870, n33871, n33872, n33873, n33874, n33876,
         n33877, n33878, n33879, n33880, n33881, n33882, n33883, n33884,
         n33885, n33886, n33887, n33888, n33889, n33890, n33891, n33892,
         n33893, n33894, n33895, n33896, n33897, n33898, n33899, n33900,
         n33901, n33902, n33903, n33904, n33905, n33906, n33907, n33908,
         n33909, n33911, n33912, n33914, n33915, n33916, n33917, n33918,
         n33919, n33920, n33921, n33922, n33923, n33924, n33925, n33926,
         n33927, n33928, n33929, n33930, n33931, n33932, n33933, n33935,
         n33936, n33937, n33938, n33939, n33940, n33941, n33942, n33943,
         n33944, n33945, n33946, n33947, n33948, n33949, n33950, n33951,
         n33952, n33953, n33954, n33955, n33956, n33957, n33960, n33961,
         n33962, n33963, n33964, n33965, n33966, n33967, n33968, n33969,
         n33970, n33971, n33972, n33973, n33974, n33975, n33976, n33977,
         n33978, n33979, n33980, n33981, n33982, n33983, n33984, n33985,
         n33986, n33987, n33988, n33989, n33990, n33991, n33992, n33993,
         n33994, n33995, n33996, n33997, n33998, n33999, n34000, n34001,
         n34002, n34003, n34004, n34005, n34006, n34007, n34008, n34009,
         n34011, n34014, n34015, n34016, n34017, n34018, n34019, n34020,
         n34021, n34022, n34023, n34024, n34025, n34026, n34027, n34028,
         n34029, n34030, n34031, n34032, n34033, n34034, n34035, n34036,
         n34037, n34039, n34040, n34041, n34042, n34043, n34044, n34045,
         n34046, n34047, n34048, n34049, n34050, n34051, n34052, n34053,
         n34054, n34055, n34056, n34057, n34059, n34060, n34061, n34062,
         n34063, n34064, n34065, n34066, n34067, n34068, n34069, n34070,
         n34071, n34072, n34073, n34074, n34075, n34076, n34077, n34078,
         n34079, n34080, n34081, n34082, n34083, n34084, n34085, n34086,
         n34087, n34088, n34089, n34090, n34091, n34092, n34093, n34094,
         n34095, n34096, n34097, n34098, n34099, n34100, n34101, n34102,
         n34103, n34104, n34105, n34106, n34107, n34108, n34109, n34110,
         n34111, n34112, n34113, n34114, n34115, n34116, n34117, n34118,
         n34119, n34120, n34121, n34122, n34123, n34124, n34125, n34126,
         n34127, n34128, n34129, n34130, n34131, n34132, n34133, n34134,
         n34135, n34136, n34137, n34138, n34139, n34140, n34142, n34143,
         n34144, n34146, n34147, n34148, n34149, n34150, n34151, n34152,
         n34153, n34154, n34155, n34156, n34157, n34158, n34159, n34160,
         n34161, n34162, n34163, n34164, n34165, n34166, n34167, n34168,
         n34169, n34170, n34171, n34172, n34173, n34174, n34175, n34176,
         n34178, n34179, n34180, n34181, n34182, n34183, n34184, n34185,
         n34186, n34187, n34188, n34189, n34190, n34191, n34192, n34193,
         n34194, n34195, n34196, n34197, n34198, n34200, n34201, n34202,
         n34203, n34204, n34205, n34206, n34207, n34208, n34209, n34210,
         n34211, n34213, n34214, n34215, n34216, n34217, n34218, n34219,
         n34220, n34221, n34222, n34224, n34225, n34226, n34227, n34228,
         n34232, n34233, n34234, n34235, n34236, n34237, n34238, n34239,
         n34240, n34241, n34242, n34243, n34244, n34246, n34247, n34248,
         n34249, n34250, n34251, n34252, n34253, n34254, n34255, n34257,
         n34258, n34259, n34260, n34261, n34262, n34263, n34264, n34265,
         n34266, n34268, n34269, n34270, n34271, n34272, n34273, n34274,
         n34275, n34276, n34277, n34278, n34280, n34281, n34282, n34283,
         n34284, n34285, n34286, n34287, n34288, n34289, n34290, n34291,
         n34292, n34293, n34294, n34295, n34298, n34300, n34302, n34303,
         n34304, n34305, n34306, n34307, n34308, n34309, n34310, n34311,
         n34312, n34313, n34314, n34315, n34316, n34317, n34318, n34319,
         n34320, n34321, n34322, n34323, n34324, n34325, n34326, n34327,
         n34329, n34330, n34331, n34332, n34333, n34334, n34335, n34336,
         n34337, n34338, n34340, n34341, n34342, n34343, n34344, n34345,
         n34346, n34347, n34348, n34349, n34350, n34351, n34352, n34353,
         n34355, n34356, n34357, n34358, n34359, n34360, n34361, n34362,
         n34363, n34364, n34365, n34366, n34368, n34369, n34370, n34371,
         n34372, n34373, n34374, n34375, n34376, n34377, n34378, n34379,
         n34380, n34381, n34382, n34383, n34384, n34385, n34386, n34387,
         n34388, n34389, n34390, n34391, n34392, n34393, n34394, n34395,
         n34397, n34398, n34399, n34400, n34402, n34403, n34404, n34405,
         n34406, n34407, n34408, n34409, n34410, n34412, n34413, n34414,
         n34415, n34416, n34417, n34418, n34419, n34420, n34421, n34422,
         n34423, n34424, n34425, n34426, n34427, n34428, n34429, n34430,
         n34431, n34432, n34433, n34434, n34435, n34436, n34437, n34438,
         n34439, n34440, n34441, n34442, n34443, n34444, n34445, n34446,
         n34447, n34448, n34450, n34451, n34452, n34453, n34454, n34455,
         n34456, n34457, n34458, n34459, n34460, n34461, n34462, n34463,
         n34464, n34465, n34466, n34467, n34468, n34469, n34470, n34471,
         n34472, n34474, n34475, n34476, n34477, n34478, n34479, n34480,
         n34481, n34482, n34483, n34484, n34485, n34486, n34487, n34488,
         n34490, n34491, n34492, n34493, n34494, n34495, n34496, n34497,
         n34498, n34499, n34500, n34501, n34502, n34503, n34504, n34505,
         n34506, n34507, n34508, n34509, n34510, n34511, n34512, n34513,
         n34514, n34515, n34516, n34517, n34518, n34519, n34520, n34521,
         n34522, n34523, n34524, n34525, n34526, n34527, n34528, n34529,
         n34530, n34531, n34532, n34533, n34534, n34535, n34536, n34537,
         n34538, n34539, n34540, n34541, n34542, n34543, n34544, n34545,
         n34546, n34547, n34548, n34549, n34550, n34551, n34552, n34553,
         n34554, n34555, n34557, n34558, n34559, n34560, n34561, n34562,
         n34563, n34564, n34565, n34566, n34567, n34568, n34569, n34570,
         n34571, n34572, n34573, n34574, n34575, n34577, n34578, n34579,
         n34581, n34582, n34583, n34585, n34586, n34587, n34588, n34589,
         n34590, n34591, n34592, n34593, n34594, n34595, n34596, n34597,
         n34598, n34599, n34600, n34601, n34602, n34603, n34604, n34606,
         n34607, n34608, n34609, n34610, n34611, n34612, n34613, n34614,
         n34615, n34616, n34618, n34619, n34620, n34621, n34622, n34623,
         n34624, n34625, n34626, n34627, n34628, n34630, n34631, n34632,
         n34633, n34634, n34635, n34636, n34637, n34638, n34639, n34640,
         n34641, n34642, n34643, n34644, n34645, n34646, n34647, n34649,
         n34650, n34651, n34652, n34653, n34654, n34655, n34656, n34657,
         n34658, n34660, n34661, n34662, n34663, n34664, n34665, n34666,
         n34667, n34668, n34669, n34670, n34671, n34672, n34673, n34674,
         n34675, n34676, n34677, n34679, n34680, n34681, n34682, n34683,
         n34684, n34685, n34687, n34688, n34689, n34691, n34694, n34695,
         n34696, n34697, n34698, n34699, n34700, n34701, n34702, n34703,
         n34704, n34705, n34706, n34707, n34708, n34709, n34710, n34711,
         n34713, n34714, n34715, n34716, n34717, n34718, n34719, n34720,
         n34721, n34722, n34723, n34724, n34725, n34726, n34727, n34730,
         n34731, n34732, n34733, n34734, n34735, n34736, n34737, n34738,
         n34739, n34740, n34741, n34742, n34743, n34744, n34745, n34746,
         n34747, n34748, n34749, n34750, n34751, n34752, n34753, n34754,
         n34755, n34758, n34759, n34760, n34761, n34763, n34764, n34765,
         n34766, n34767, n34768, n34769, n34770, n34771, n34773, n34774,
         n34775, n34776, n34777, n34778, n34779, n34780, n34781, n34783,
         n34784, n34785, n34786, n34787, n34789, n34790, n34791, n34792,
         n34793, n34795, n34796, n34797, n34798, n34799, n34800, n34801,
         n34802, n34804, n34805, n34806, n34807, n34808, n34809, n34810,
         n34811, n34815, n34816, n34817, n34818, n34819, n34820, n34821,
         n34822, n34823, n34825, n34826, n34827, n34828, n34829, n34830,
         n34832, n34833, n34834, n34835, n34836, n34837, n34838, n34839,
         n34840, n34841, n34842, n34843, n34844, n34845, n34846, n34847,
         n34848, n34849, n34850, n34851, n34852, n34853, n34854, n34855,
         n34856, n34857, n34858, n34859, n34860, n34861, n34862, n34863,
         n34864, n34865, n34866, n34868, n34869, n34870, n34871, n34872,
         n34873, n34874, n34875, n34876, n34877, n34878, n34879, n34881,
         n34882, n34883, n34884, n34885, n34886, n34887, n34888, n34889,
         n34890, n34891, n34892, n34893, n34894, n34895, n34896, n34897,
         n34898, n34899, n34902, n34903, n34904, n34906, n34907, n34908,
         n34909, n34910, n34911, n34912, n34913, n34914, n34915, n34916,
         n34917, n34918, n34919, n34920, n34921, n34923, n34924, n34925,
         n34926, n34927, n34928, n34929, n34930, n34931, n34932, n34933,
         n34934, n34935, n34936, n34937, n34938, n34940, n34941, n34942,
         n34946, n34947, n34948, n34949, n34950, n34951, n34952, n34953,
         n34956, n34957, n34958, n34959, n34960, n34961, n34962, n34963,
         n34964, n34965, n34966, n34967, n34968, n34969, n34970, n34971,
         n34972, n34973, n34974, n34976, n34977, n34978, n34979, n34980,
         n34981, n34982, n34983, n34984, n34986, n34988, n34989, n34990,
         n34991, n34992, n34993, n34994, n34995, n34996, n34997, n34998,
         n34999, n35001, n35002, n35003, n35004, n35005, n35006, n35007,
         n35008, n35011, n35013, n35014, n35015, n35016, n35017, n35018,
         n35019, n35020, n35021, n35022, n35023, n35024, n35025, n35026,
         n35027, n35029, n35030, n35031, n35032, n35033, n35034, n35035,
         n35036, n35037, n35038, n35039, n35041, n35042, n35044, n35045,
         n35046, n35047, n35048, n35049, n35050, n35051, n35052, n35053,
         n35054, n35055, n35056, n35057, n35059, n35061, n35062, n35063,
         n35064, n35065, n35066, n35067, n35068, n35070, n35071, n35072,
         n35073, n35075, n35076, n35077, n35078, n35079, n35080, n35081,
         n35082, n35083, n35084, n35085, n35086, n35087, n35089, n35091,
         n35092, n35093, n35094, n35095, n35096, n35097, n35098, n35099,
         n35100, n35101, n35102, n35103, n35104, n35105, n35108, n35109,
         n35110, n35111, n35112, n35113, n35114, n35115, n35116, n35117,
         n35118, n35119, n35120, n35121, n35122, n35124, n35125, n35126,
         n35128, n35130, n35131, n35132, n35133, n35134, n35135, n35136,
         n35137, n35138, n35139, n35140, n35141, n35142, n35143, n35144,
         n35145, n35146, n35147, n35148, n35149, n35150, n35151, n35152,
         n35153, n35154, n35159, n35160, n35161, n35162, n35163, n35164,
         n35165, n35167, n35170, n35171, n35173, n35174, n35176, n35177,
         n35178, n35179, n35180, n35181, n35182, n35183, n35184, n35185,
         n35186, n35187, n35188, n35189, n35190, n35191, n35192, n35194,
         n35195, n35196, n35197, n35198, n35199, n35200, n35201, n35202,
         n35203, n35204, n35205, n35206, n35207, n35208, n35209, n35210,
         n35211, n35212, n35213, n35214, n35215, n35217, n35218, n35219,
         n35220, n35222, n35224, n35225, n35226, n35228, n35229, n35230,
         n35231, n35232, n35233, n35234, n35235, n35236, n35238, n35240,
         n35241, n35242, n35243, n35244, n35245, n35246, n35247, n35248,
         n35249, n35250, n35251, n35252, n35254, n35255, n35256, n35257,
         n35258, n35259, n35260, n35261, n35262, n35263, n35264, n35265,
         n35266, n35267, n35268, n35269, n35270, n35271, n35272, n35273,
         n35274, n35275, n35276, n35277, n35278, n35279, n35280, n35281,
         n35282, n35283, n35284, n35285, n35286, n35287, n35288, n35289,
         n35290, n35291, n35292, n35294, n35295, n35296, n35297, n35298,
         n35299, n35300, n35301, n35302, n35303, n35304, n35305, n35306,
         n35307, n35308, n35309, n35310, n35311, n35312, n35313, n35314,
         n35315, n35316, n35317, n35318, n35319, n35320, n35321, n35322,
         n35323, n35324, n35325, n35326, n35327, n35328, n35329, n35330,
         n35331, n35333, n35334, n35335, n35336, n35337, n35338, n35339,
         n35340, n35341, n35343, n35344, n35345, n35346, n35348, n35349,
         n35350, n35351, n35352, n35353, n35354, n35355, n35357, n35358,
         n35360, n35361, n35362, n35363, n35364, n35365, n35366, n35367,
         n35368, n35369, n35370, n35371, n35372, n35373, n35374, n35375,
         n35376, n35377, n35378, n35379, n35380, n35381, n35382, n35383,
         n35384, n35385, n35386, n35387, n35388, n35389, n35390, n35391,
         n35392, n35393, n35394, n35395, n35396, n35397, n35398, n35399,
         n35400, n35401, n35402, n35403, n35404, n35405, n35407, n35408,
         n35409, n35410, n35411, n35412, n35413, n35414, n35415, n35416,
         n35417, n35418, n35419, n35420, n35421, n35422, n35423, n35424,
         n35425, n35426, n35427, n35428, n35429, n35430, n35431, n35432,
         n35433, n35434, n35435, n35436, n35437, n35438, n35439, n35440,
         n35441, n35443, n35444, n35445, n35446, n35447, n35449, n35450,
         n35451, n35452, n35453, n35454, n35455, n35456, n35457, n35458,
         n35459, n35460, n35461, n35463, n35464, n35465, n35466, n35467,
         n35468, n35469, n35470, n35472, n35473, n35476, n35478, n35480,
         n35482, n35483, n35484, n35485, n35486, n35487, n35488, n35489,
         n35490, n35491, n35492, n35493, n35494, n35495, n35496, n35497,
         n35499, n35500, n35501, n35502, n35503, n35504, n35505, n35506,
         n35507, n35508, n35509, n35510, n35511, n35512, n35513, n35514,
         n35515, n35516, n35517, n35518, n35519, n35520, n35521, n35522,
         n35523, n35524, n35525, n35526, n35528, n35529, n35530, n35532,
         n35533, n35534, n35535, n35536, n35537, n35538, n35540, n35541,
         n35543, n35544, n35546, n35547, n35548, n35549, n35550, n35551,
         n35552, n35554, n35555, n35556, n35557, n35558, n35559, n35560,
         n35561, n35562, n35563, n35564, n35565, n35566, n35567, n35568,
         n35569, n35570, n35571, n35572, n35573, n35574, n35575, n35576,
         n35577, n35578, n35579, n35580, n35581, n35582, n35583, n35584,
         n35585, n35588, n35589, n35590, n35591, n35592, n35593, n35594,
         n35595, n35598, n35599, n35600, n35602, n35603, n35604, n35605,
         n35606, n35607, n35608, n35609, n35611, n35612, n35613, n35614,
         n35615, n35617, n35618, n35619, n35620, n35621, n35622, n35623,
         n35624, n35625, n35626, n35627, n35628, n35629, n35630, n35631,
         n35632, n35633, n35634, n35635, n35637, n35638, n35639, n35641,
         n35642, n35643, n35644, n35645, n35646, n35647, n35648, n35649,
         n35650, n35651, n35652, n35653, n35654, n35655, n35656, n35657,
         n35658, n35659, n35660, n35661, n35662, n35663, n35664, n35665,
         n35666, n35667, n35668, n35669, n35670, n35673, n35674, n35675,
         n35677, n35678, n35679, n35680, n35681, n35682, n35683, n35684,
         n35685, n35686, n35687, n35688, n35689, n35690, n35691, n35692,
         n35694, n35695, n35696, n35697, n35698, n35699, n35700, n35701,
         n35702, n35703, n35704, n35705, n35706, n35707, n35708, n35709,
         n35710, n35711, n35712, n35713, n35714, n35715, n35717, n35718,
         n35719, n35721, n35722, n35723, n35724, n35725, n35726, n35728,
         n35729, n35730, n35731, n35732, n35733, n35734, n35735, n35737,
         n35738, n35739, n35740, n35741, n35743, n35744, n35745, n35746,
         n35747, n35748, n35749, n35750, n35751, n35752, n35753, n35754,
         n35755, n35756, n35758, n35759, n35760, n35761, n35762, n35763,
         n35764, n35765, n35766, n35767, n35768, n35769, n35770, n35771,
         n35772, n35773, n35774, n35775, n35776, n35777, n35778, n35779,
         n35780, n35781, n35782, n35783, n35785, n35786, n35787, n35788,
         n35789, n35790, n35791, n35792, n35793, n35794, n35795, n35796,
         n35797, n35798, n35799, n35800, n35801, n35802, n35803, n35804,
         n35805, n35806, n35807, n35808, n35809, n35810, n35811, n35813,
         n35815, n35816, n35817, n35818, n35819, n35820, n35821, n35822,
         n35823, n35824, n35826, n35827, n35828, n35830, n35832, n35833,
         n35834, n35835, n35836, n35837, n35838, n35839, n35840, n35841,
         n35842, n35844, n35845, n35846, n35847, n35848, n35849, n35850,
         n35851, n35852, n35854, n35855, n35856, n35857, n35858, n35859,
         n35860, n35861, n35862, n35863, n35864, n35865, n35866, n35867,
         n35868, n35869, n35870, n35871, n35873, n35874, n35876, n35877,
         n35878, n35879, n35880, n35881, n35882, n35883, n35884, n35885,
         n35886, n35887, n35888, n35889, n35890, n35892, n35894, n35895,
         n35896, n35897, n35898, n35899, n35900, n35901, n35902, n35903,
         n35905, n35906, n35907, n35908, n35909, n35910, n35911, n35912,
         n35913, n35914, n35915, n35916, n35917, n35918, n35919, n35920,
         n35921, n35922, n35923, n35924, n35925, n35926, n35927, n35928,
         n35929, n35930, n35931, n35932, n35933, n35934, n35935, n35936,
         n35937, n35938, n35939, n35940, n35941, n35942, n35943, n35944,
         n35945, n35946, n35947, n35948, n35949, n35950, n35951, n35952,
         n35953, n35954, n35955, n35956, n35957, n35958, n35959, n35960,
         n35961, n35962, n35963, n35964, n35965, n35966, n35967, n35968,
         n35969, n35970, n35971, n35972, n35973, n35974, n35975, n35976,
         n35977, n35978, n35979, n35980, n35981, n35982, n35983, n35984,
         n35985, n35986, n35987, n35988, n35989, n35990, n35991, n35992,
         n35993, n35994, n35995, n35996, n35997, n35999, n36000, n36001,
         n36002, n36003, n36004, n36005, n36006, n36007, n36008, n36009,
         n36010, n36011, n36012, n36013, n36014, n36015, n36016, n36017,
         n36018, n36019, n36020, n36021, n36022, n36024, n36025, n36026,
         n36027, n36028, n36029, n36030, n36031, n36032, n36034, n36035,
         n36036, n36037, n36038, n36039, n36040, n36041, n36042, n36043,
         n36044, n36045, n36046, n36047, n36048, n36049, n36050, n36051,
         n36052, n36053, n36054, n36055, n36056, n36057, n36058, n36059,
         n36060, n36061, n36062, n36063, n36065, n36066, n36067, n36068,
         n36069, n36070, n36071, n36072, n36074, n36075, n36076, n36077,
         n36079, n36080, n36081, n36082, n36083, n36084, n36086, n36087,
         n36088, n36089, n36090, n36091, n36092, n36093, n36094, n36095,
         n36096, n36097, n36098, n36099, n36100, n36101, n36102, n36103,
         n36104, n36105, n36106, n36107, n36108, n36109, n36110, n36111,
         n36112, n36113, n36114, n36115, n36116, n36117, n36118, n36119,
         n36120, n36121, n36122, n36123, n36124, n36125, n36127, n36129,
         n36130, n36131, n36132, n36133, n36134, n36135, n36136, n36137,
         n36138, n36139, n36140, n36141, n36142, n36144, n36145, n36146,
         n36147, n36148, n36149, n36150, n36151, n36152, n36153, n36154,
         n36155, n36156, n36157, n36158, n36159, n36160, n36161, n36162,
         n36163, n36164, n36165, n36166, n36167, n36168, n36169, n36170,
         n36171, n36172, n36173, n36174, n36175, n36176, n36177, n36178,
         n36179, n36180, n36181, n36182, n36183, n36184, n36185, n36186,
         n36187, n36188, n36189, n36190, n36191, n36192, n36193, n36194,
         n36195, n36196, n36197, n36198, n36199, n36200, n36201, n36202,
         n36203, n36204, n36205, n36206, n36207, n36209, n36210, n36211,
         n36212, n36213, n36215, n36216, n36217, n36218, n36219, n36220,
         n36221, n36223, n36224, n36225, n36226, n36227, n36228, n36229,
         n36231, n36232, n36233, n36234, n36235, n36237, n36238, n36239,
         n36240, n36241, n36242, n36243, n36244, n36245, n36246, n36247,
         n36248, n36249, n36252, n36253, n36255, n36256, n36257, n36258,
         n36259, n36260, n36261, n36262, n36263, n36264, n36265, n36266,
         n36267, n36268, n36269, n36271, n36272, n36273, n36274, n36275,
         n36276, n36277, n36278, n36279, n36280, n36281, n36282, n36283,
         n36284, n36285, n36287, n36288, n36289, n36290, n36291, n36292,
         n36293, n36294, n36295, n36297, n36298, n36299, n36300, n36301,
         n36302, n36303, n36304, n36305, n36306, n36307, n36308, n36309,
         n36310, n36311, n36312, n36313, n36315, n36317, n36318, n36319,
         n36320, n36321, n36322, n36323, n36324, n36325, n36326, n36327,
         n36328, n36329, n36331, n36332, n36333, n36334, n36335, n36336,
         n36337, n36338, n36339, n36340, n36341, n36342, n36343, n36344,
         n36345, n36346, n36347, n36348, n36349, n36350, n36351, n36352,
         n36353, n36354, n36356, n36357, n36358, n36359, n36360, n36361,
         n36362, n36363, n36364, n36365, n36366, n36368, n36369, n36370,
         n36371, n36372, n36373, n36374, n36375, n36377, n36378, n36379,
         n36380, n36381, n36384, n36385, n36386, n36389, n36390, n36391,
         n36393, n36394, n36395, n36396, n36398, n36399, n36401, n36402,
         n36403, n36404, n36405, n36406, n36407, n36408, n36409, n36410,
         n36411, n36412, n36413, n36414, n36415, n36416, n36417, n36418,
         n36419, n36420, n36421, n36422, n36423, n36424, n36425, n36427,
         n36428, n36429, n36430, n36431, n36432, n36433, n36434, n36435,
         n36436, n36437, n36438, n36439, n36440, n36441, n36442, n36443,
         n36444, n36445, n36446, n36447, n36448, n36449, n36450, n36451,
         n36452, n36453, n36454, n36455, n36456, n36458, n36459, n36460,
         n36461, n36462, n36463, n36464, n36465, n36466, n36467, n36468,
         n36469, n36470, n36471, n36472, n36473, n36474, n36475, n36476,
         n36477, n36478, n36480, n36481, n36482, n36483, n36484, n36485,
         n36486, n36487, n36488, n36489, n36490, n36491, n36492, n36493,
         n36494, n36495, n36496, n36497, n36498, n36499, n36500, n36501,
         n36503, n36504, n36505, n36506, n36507, n36508, n36509, n36510,
         n36511, n36512, n36513, n36514, n36515, n36517, n36518, n36519,
         n36520, n36522, n36523, n36524, n36525, n36526, n36527, n36528,
         n36529, n36530, n36531, n36532, n36533, n36534, n36535, n36536,
         n36537, n36538, n36539, n36540, n36541, n36542, n36543, n36544,
         n36545, n36546, n36547, n36548, n36549, n36550, n36551, n36552,
         n36553, n36554, n36555, n36556, n36557, n36558, n36559, n36560,
         n36561, n36563, n36564, n36565, n36566, n36567, n36568, n36569,
         n36570, n36572, n36573, n36574, n36575, n36576, n36577, n36578,
         n36579, n36580, n36582, n36583, n36584, n36585, n36586, n36587,
         n36588, n36589, n36590, n36591, n36592, n36593, n36594, n36595,
         n36596, n36597, n36598, n36599, n36600, n36601, n36602, n36604,
         n36605, n36606, n36607, n36608, n36609, n36610, n36611, n36612,
         n36613, n36614, n36615, n36616, n36617, n36618, n36619, n36620,
         n36621, n36622, n36623, n36624, n36625, n36626, n36627, n36628,
         n36629, n36630, n36631, n36632, n36633, n36634, n36635, n36636,
         n36637, n36638, n36639, n36640, n36641, n36642, n36643, n36644,
         n36645, n36646, n36647, n36648, n36649, n36650, n36651, n36652,
         n36653, n36654, n36656, n36657, n36658, n36659, n36660, n36661,
         n36662, n36663, n36664, n36665, n36666, n36667, n36669, n36670,
         n36671, n36672, n36673, n36674, n36675, n36676, n36677, n36678,
         n36679, n36680, n36681, n36682, n36683, n36685, n36686, n36687,
         n36688, n36689, n36690, n36691, n36692, n36693, n36694, n36695,
         n36696, n36697, n36698, n36699, n36700, n36701, n36703, n36705,
         n36706, n36707, n36708, n36709, n36710, n36711, n36712, n36713,
         n36715, n36716, n36717, n36718, n36719, n36720, n36721, n36722,
         n36723, n36724, n36725, n36726, n36727, n36728, n36729, n36730,
         n36731, n36732, n36733, n36734, n36735, n36736, n36737, n36738,
         n36739, n36740, n36741, n36742, n36743, n36744, n36745, n36746,
         n36747, n36748, n36749, n36750, n36751, n36752, n36753, n36754,
         n36755, n36756, n36758, n36759, n36760, n36761, n36763, n36764,
         n36765, n36766, n36767, n36768, n36769, n36770, n36771, n36772,
         n36773, n36774, n36775, n36776, n36777, n36778, n36779, n36780,
         n36781, n36782, n36783, n36785, n36786, n36787, n36788, n36789,
         n36790, n36791, n36792, n36793, n36794, n36796, n36798, n36799,
         n36800, n36801, n36803, n36804, n36805, n36806, n36808, n36809,
         n36810, n36811, n36812, n36813, n36814, n36815, n36816, n36817,
         n36818, n36819, n36820, n36821, n36822, n36823, n36824, n36825,
         n36826, n36827, n36828, n36829, n36830, n36831, n36832, n36833,
         n36834, n36835, n36837, n36838, n36841, n36842, n36843, n36844,
         n36846, n36847, n36848, n36850, n36851, n36852, n36853, n36854,
         n36855, n36856, n36857, n36858, n36859, n36860, n36861, n36862,
         n36863, n36864, n36865, n36866, n36867, n36868, n36869, n36870,
         n36871, n36872, n36873, n36874, n36875, n36876, n36878, n36879,
         n36880, n36881, n36882, n36883, n36884, n36886, n36888, n36889,
         n36890, n36891, n36892, n36893, n36894, n36895, n36897, n36898,
         n36899, n36900, n36901, n36902, n36903, n36904, n36905, n36906,
         n36907, n36908, n36909, n36910, n36911, n36912, n36913, n36914,
         n36915, n36916, n36917, n36918, n36919, n36920, n36921, n36922,
         n36923, n36924, n36926, n36927, n36928, n36929, n36930, n36931,
         n36932, n36933, n36934, n36935, n36936, n36937, n36938, n36939,
         n36940, n36941, n36942, n36943, n36944, n36945, n36946, n36947,
         n36948, n36949, n36950, n36951, n36952, n36953, n36954, n36955,
         n36956, n36957, n36958, n36959, n36960, n36961, n36962, n36963,
         n36964, n36965, n36966, n36967, n36968, n36969, n36970, n36971,
         n36972, n36973, n36974, n36975, n36976, n36978, n36979, n36980,
         n36981, n36982, n36983, n36984, n36986, n36987, n36988, n36989,
         n36990, n36991, n36992, n36993, n36994, n36995, n36996, n36997,
         n36998, n36999, n37000, n37001, n37002, n37003, n37004, n37005,
         n37006, n37007, n37008, n37009, n37010, n37011, n37012, n37013,
         n37014, n37015, n37016, n37017, n37018, n37019, n37020, n37021,
         n37022, n37023, n37024, n37025, n37026, n37027, n37028, n37029,
         n37030, n37031, n37032, n37033, n37034, n37035, n37036, n37037,
         n37038, n37039, n37040, n37041, n37042, n37043, n37044, n37045,
         n37046, n37047, n37048, n37049, n37050, n37051, n37052, n37053,
         n37054, n37055, n37056, n37057, n37058, n37059, n37060, n37061,
         n37062, n37064, n37065, n37067, n37068, n37069, n37070, n37072,
         n37073, n37074, n37075, n37076, n37077, n37078, n37079, n37080,
         n37081, n37082, n37083, n37084, n37085, n37086, n37087, n37090,
         n37091, n37092, n37093, n37094, n37095, n37096, n37097, n37098,
         n37099, n37100, n37101, n37102, n37104, n37105, n37106, n37107,
         n37108, n37109, n37110, n37111, n37112, n37113, n37114, n37115,
         n37116, n37117, n37118, n37119, n37120, n37121, n37123, n37125,
         n37126, n37127, n37128, n37129, n37130, n37131, n37132, n37133,
         n37134, n37135, n37136, n37137, n37138, n37139, n37140, n37141,
         n37142, n37143, n37144, n37145, n37146, n37147, n37148, n37149,
         n37150, n37151, n37152, n37153, n37154, n37155, n37156, n37157,
         n37158, n37159, n37160, n37161, n37162, n37163, n37164, n37165,
         n37166, n37167, n37168, n37169, n37170, n37171, n37172, n37173,
         n37174, n37175, n37176, n37177, n37178, n37179, n37180, n37181,
         n37182, n37183, n37184, n37185, n37187, n37188, n37189, n37190,
         n37191, n37192, n37193, n37194, n37196, n37197, n37198, n37199,
         n37200, n37203, n37204, n37205, n37206, n37207, n37208, n37209,
         n37210, n37211, n37212, n37214, n37216, n37217, n37218, n37219,
         n37220, n37221, n37222, n37223, n37224, n37225, n37227, n37228,
         n37229, n37230, n37231, n37232, n37233, n37234, n37235, n37236,
         n37237, n37238, n37239, n37240, n37242, n37243, n37244, n37245,
         n37246, n37247, n37248, n37249, n37252, n37253, n37254, n37255,
         n37256, n37257, n37258, n37259, n37260, n37261, n37262, n37263,
         n37264, n37265, n37266, n37267, n37268, n37269, n37270, n37271,
         n37272, n37273, n37274, n37276, n37277, n37278, n37279, n37280,
         n37281, n37282, n37283, n37284, n37285, n37286, n37287, n37288,
         n37289, n37290, n37291, n37292, n37293, n37294, n37295, n37296,
         n37297, n37298, n37299, n37300, n37301, n37302, n37303, n37304,
         n37305, n37306, n37307, n37308, n37309, n37310, n37311, n37312,
         n37313, n37314, n37315, n37316, n37317, n37319, n37321, n37322,
         n37323, n37324, n37325, n37326, n37327, n37328, n37329, n37330,
         n37331, n37332, n37333, n37334, n37335, n37336, n37337, n37338,
         n37339, n37340, n37341, n37342, n37343, n37344, n37345, n37346,
         n37347, n37348, n37349, n37350, n37351, n37352, n37354, n37355,
         n37356, n37357, n37358, n37359, n37360, n37361, n37363, n37364,
         n37365, n37366, n37367, n37368, n37369, n37370, n37371, n37373,
         n37374, n37375, n37376, n37378, n37379, n37380, n37381, n37382,
         n37383, n37384, n37385, n37386, n37387, n37388, n37389, n37390,
         n37391, n37392, n37393, n37394, n37395, n37396, n37397, n37398,
         n37399, n37400, n37401, n37402, n37403, n37404, n37405, n37406,
         n37407, n37408, n37409, n37410, n37411, n37412, n37413, n37414,
         n37415, n37416, n37418, n37419, n37420, n37421, n37422, n37423,
         n37424, n37425, n37426, n37427, n37428, n37429, n37430, n37431,
         n37432, n37433, n37434, n37435, n37436, n37437, n37439, n37440,
         n37441, n37442, n37443, n37444, n37445, n37446, n37447, n37448,
         n37449, n37451, n37452, n37453, n37454, n37455, n37456, n37457,
         n37458, n37459, n37460, n37461, n37462, n37463, n37464, n37465,
         n37466, n37467, n37468, n37469, n37470, n37471, n37472, n37473,
         n37474, n37475, n37476, n37477, n37478, n37479, n37480, n37481,
         n37482, n37483, n37484, n37485, n37486, n37487, n37488, n37489,
         n37490, n37491, n37492, n37493, n37494, n37495, n37496, n37497,
         n37498, n37499, n37500, n37501, n37502, n37503, n37504, n37505,
         n37506, n37507, n37508, n37509, n37510, n37511, n37512, n37513,
         n37514, n37515, n37516, n37517, n37518, n37519, n37520, n37521,
         n37522, n37523, n37524, n37525, n37526, n37527, n37528, n37529,
         n37530, n37531, n37532, n37533, n37534, n37535, n37536, n37537,
         n37538, n37539, n37541, n37542, n37543, n37544, n37545, n37546,
         n37547, n37549, n37550, n37552, n37553, n37554, n37555, n37556,
         n37557, n37558, n37559, n37560, n37561, n37562, n37563, n37564,
         n37565, n37566, n37567, n37568, n37569, n37570, n37571, n37572,
         n37573, n37574, n37575, n37576, n37577, n37578, n37579, n37580,
         n37581, n37582, n37583, n37584, n37585, n37586, n37587, n37588,
         n37590, n37592, n37593, n37594, n37595, n37596, n37597, n37598,
         n37600, n37601, n37602, n37603, n37604, n37605, n37606, n37607,
         n37608, n37609, n37610, n37611, n37612, n37613, n37614, n37615,
         n37616, n37617, n37618, n37619, n37620, n37621, n37622, n37623,
         n37624, n37625, n37626, n37627, n37628, n37629, n37630, n37631,
         n37632, n37633, n37634, n37635, n37636, n37637, n37638, n37639,
         n37640, n37641, n37642, n37643, n37644, n37645, n37646, n37647,
         n37648, n37649, n37650, n37651, n37652, n37653, n37654, n37655,
         n37656, n37657, n37659, n37660, n37661, n37662, n37663, n37664,
         n37665, n37666, n37667, n37668, n37669, n37670, n37671, n37673,
         n37674, n37675, n37676, n37677, n37678, n37679, n37680, n37681,
         n37682, n37683, n37684, n37685, n37686, n37687, n37688, n37689,
         n37690, n37691, n37692, n37693, n37694, n37695, n37696, n37697,
         n37698, n37699, n37701, n37702, n37703, n37704, n37705, n37706,
         n37708, n37709, n37710, n37711, n37712, n37713, n37714, n37715,
         n37716, n37717, n37718, n37719, n37720, n37721, n37722, n37723,
         n37724, n37725, n37726, n37727, n37729, n37730, n37731, n37732,
         n37733, n37734, n37735, n37736, n37737, n37738, n37739, n37740,
         n37741, n37742, n37743, n37744, n37745, n37746, n37747, n37748,
         n37749, n37750, n37751, n37752, n37753, n37754, n37755, n37757,
         n37758, n37759, n37760, n37761, n37762, n37763, n37764, n37765,
         n37766, n37767, n37768, n37769, n37770, n37772, n37773, n37774,
         n37775, n37777, n37778, n37779, n37780, n37781, n37782, n37783,
         n37785, n37786, n37787, n37788, n37789, n37790, n37791, n37792,
         n37793, n37794, n37795, n37796, n37797, n37798, n37799, n37800,
         n37801, n37802, n37803, n37804, n37805, n37806, n37807, n37808,
         n37809, n37810, n37811, n37812, n37813, n37814, n37816, n37817,
         n37818, n37819, n37820, n37821, n37822, n37823, n37824, n37825,
         n37827, n37828, n37829, n37830, n37831, n37832, n37833, n37834,
         n37835, n37836, n37837, n37838, n37839, n37840, n37842, n37843,
         n37844, n37845, n37846, n37847, n37848, n37849, n37850, n37851,
         n37852, n37853, n37854, n37855, n37856, n37857, n37858, n37859,
         n37860, n37861, n37862, n37863, n37864, n37865, n37866, n37867,
         n37868, n37869, n37870, n37871, n37872, n37873, n37874, n37875,
         n37876, n37877, n37878, n37879, n37880, n37881, n37882, n37883,
         n37884, n37885, n37886, n37887, n37888, n37889, n37890, n37891,
         n37892, n37893, n37894, n37895, n37896, n37897, n37898, n37899,
         n37900, n37901, n37902, n37904, n37906, n37907, n37908, n37909,
         n37910, n37911, n37912, n37913, n37914, n37915, n37916, n37917,
         n37919, n37920, n37921, n37922, n37923, n37924, n37926, n37927,
         n37928, n37930, n37931, n37933, n37934, n37935, n37936, n37937,
         n37938, n37939, n37940, n37941, n37942, n37943, n37944, n37945,
         n37946, n37947, n37948, n37949, n37950, n37951, n37952, n37953,
         n37954, n37955, n37956, n37957, n37958, n37959, n37960, n37961,
         n37962, n37963, n37964, n37965, n37966, n37967, n37969, n37970,
         n37971, n37972, n37973, n37974, n37975, n37978, n37979, n37980,
         n37981, n37982, n37983, n37984, n37985, n37986, n37987, n37988,
         n37989, n37990, n37991, n37992, n37993, n37994, n37995, n37996,
         n37997, n37998, n37999, n38000, n38001, n38002, n38003, n38004,
         n38005, n38006, n38007, n38008, n38009, n38010, n38011, n38012,
         n38013, n38014, n38015, n38017, n38018, n38020, n38021, n38022,
         n38023, n38024, n38025, n38026, n38027, n38028, n38029, n38030,
         n38031, n38032, n38033, n38034, n38035, n38036, n38037, n38038,
         n38039, n38040, n38041, n38042, n38043, n38044, n38045, n38046,
         n38047, n38048, n38049, n38050, n38051, n38055, n38056, n38057,
         n38058, n38059, n38060, n38061, n38062, n38063, n38064, n38065,
         n38066, n38067, n38068, n38069, n38070, n38071, n38072, n38073,
         n38074, n38075, n38076, n38077, n38078, n38079, n38080, n38081,
         n38083, n38084, n38085, n38086, n38087, n38088, n38089, n38090,
         n38091, n38092, n38093, n38094, n38095, n38096, n38097, n38098,
         n38099, n38100, n38101, n38102, n38103, n38104, n38105, n38106,
         n38107, n38108, n38109, n38110, n38111, n38112, n38113, n38114,
         n38115, n38116, n38117, n38118, n38119, n38120, n38121, n38122,
         n38123, n38124, n38125, n38126, n38127, n38128, n38129, n38130,
         n38131, n38132, n38133, n38134, n38135, n38136, n38137, n38138,
         n38139, n38140, n38142, n38144, n38145, n38146, n38147, n38148,
         n38149, n38150, n38151, n38152, n38153, n38154, n38155, n38156,
         n38158, n38159, n38160, n38161, n38162, n38163, n38164, n38165,
         n38166, n38167, n38168, n38169, n38170, n38171, n38172, n38173,
         n38174, n38175, n38176, n38177, n38178, n38179, n38180, n38181,
         n38182, n38183, n38184, n38185, n38186, n38187, n38188, n38189,
         n38190, n38191, n38192, n38193, n38194, n38196, n38197, n38198,
         n38199, n38200, n38201, n38203, n38204, n38205, n38206, n38207,
         n38208, n38209, n38210, n38211, n38212, n38213, n38214, n38215,
         n38216, n38217, n38218, n38219, n38220, n38221, n38222, n38223,
         n38224, n38225, n38226, n38227, n38228, n38229, n38230, n38231,
         n38232, n38233, n38234, n38235, n38236, n38237, n38238, n38239,
         n38240, n38241, n38242, n38243, n38244, n38245, n38246, n38247,
         n38248, n38249, n38250, n38251, n38252, n38253, n38254, n38255,
         n38257, n38258, n38259, n38260, n38262, n38263, n38264, n38265,
         n38266, n38267, n38269, n38270, n38271, n38272, n38273, n38274,
         n38275, n38276, n38277, n38278, n38279, n38280, n38281, n38282,
         n38283, n38284, n38285, n38286, n38287, n38288, n38289, n38290,
         n38291, n38292, n38293, n38294, n38295, n38297, n38298, n38299,
         n38300, n38301, n38302, n38303, n38304, n38305, n38306, n38307,
         n38308, n38309, n38310, n38311, n38312, n38313, n38314, n38315,
         n38316, n38317, n38318, n38319, n38320, n38321, n38322, n38323,
         n38324, n38325, n38326, n38327, n38328, n38329, n38330, n38331,
         n38332, n38333, n38334, n38335, n38336, n38337, n38338, n38339,
         n38340, n38341, n38342, n38343, n38344, n38345, n38346, n38347,
         n38348, n38349, n38350, n38351, n38352, n38353, n38354, n38355,
         n38357, n38358, n38359, n38360, n38361, n38362, n38363, n38364,
         n38365, n38366, n38367, n38368, n38369, n38370, n38371, n38372,
         n38373, n38374, n38375, n38376, n38377, n38378, n38379, n38380,
         n38381, n38382, n38383, n38384, n38385, n38386, n38387, n38388,
         n38389, n38390, n38391, n38392, n38393, n38394, n38395, n38397,
         n38398, n38399, n38400, n38401, n38402, n38403, n38404, n38405,
         n38406, n38407, n38408, n38409, n38410, n38411, n38412, n38413,
         n38414, n38415, n38416, n38417, n38418, n38419, n38420, n38421,
         n38422, n38423, n38424, n38425, n38426, n38428, n38429, n38430,
         n38431, n38432, n38433, n38434, n38435, n38436, n38437, n38438,
         n38439, n38440, n38441, n38442, n38443, n38444, n38445, n38446,
         n38447, n38448, n38449, n38450, n38451, n38452, n38453, n38454,
         n38455, n38456, n38457, n38458, n38459, n38460, n38461, n38462,
         n38463, n38464, n38465, n38466, n38467, n38468, n38469, n38470,
         n38471, n38472, n38473, n38474, n38475, n38476, n38477, n38478,
         n38479, n38480, n38481, n38482, n38483, n38484, n38485, n38486,
         n38487, n38488, n38489, n38490, n38491, n38493, n38494, n38495,
         n38496, n38497, n38498, n38499, n38500, n38501, n38502, n38503,
         n38504, n38505, n38506, n38507, n38509, n38510, n38511, n38512,
         n38513, n38514, n38516, n38517, n38518, n38519, n38520, n38521,
         n38522, n38523, n38524, n38525, n38526, n38527, n38529, n38530,
         n38531, n38532, n38533, n38534, n38535, n38536, n38537, n38538,
         n38540, n38541, n38542, n38543, n38544, n38545, n38546, n38547,
         n38548, n38549, n38550, n38551, n38552, n38553, n38554, n38555,
         n38556, n38557, n38558, n38559, n38560, n38561, n38562, n38563,
         n38564, n38565, n38566, n38567, n38568, n38569, n38570, n38571,
         n38572, n38573, n38574, n38575, n38576, n38577, n38578, n38579,
         n38580, n38581, n38582, n38583, n38584, n38585, n38586, n38587,
         n38588, n38589, n38590, n38591, n38592, n38593, n38595, n38596,
         n38597, n38598, n38599, n38600, n38601, n38602, n38603, n38604,
         n38605, n38606, n38607, n38608, n38609, n38610, n38611, n38612,
         n38613, n38614, n38615, n38616, n38617, n38618, n38619, n38620,
         n38621, n38622, n38623, n38624, n38625, n38626, n38627, n38628,
         n38629, n38630, n38631, n38632, n38633, n38634, n38635, n38636,
         n38637, n38638, n38639, n38640, n38641, n38642, n38643, n38644,
         n38645, n38646, n38647, n38648, n38649, n38650, n38651, n38652,
         n38653, n38654, n38655, n38656, n38658, n38659, n38660, n38661,
         n38662, n38663, n38664, n38665, n38666, n38667, n38668, n38669,
         n38670, n38671, n38672, n38674, n38675, n38676, n38677, n38678,
         n38679, n38680, n38681, n38682, n38683, n38684, n38685, n38686,
         n38689, n38690, n38691, n38692, n38693, n38695, n38696, n38697,
         n38698, n38699, n38700, n38701, n38702, n38703, n38704, n38705,
         n38706, n38707, n38708, n38709, n38710, n38711, n38713, n38714,
         n38715, n38716, n38718, n38720, n38721, n38722, n38723, n38724,
         n38725, n38726, n38727, n38728, n38729, n38731, n38732, n38733,
         n38734, n38735, n38736, n38737, n38738, n38739, n38740, n38741,
         n38742, n38743, n38744, n38745, n38746, n38747, n38748, n38749,
         n38750, n38752, n38753, n38754, n38755, n38756, n38757, n38758,
         n38759, n38760, n38761, n38762, n38763, n38764, n38765, n38766,
         n38767, n38768, n38769, n38770, n38771, n38772, n38773, n38774,
         n38775, n38776, n38777, n38778, n38779, n38780, n38781, n38782,
         n38784, n38785, n38786, n38787, n38788, n38789, n38790, n38791,
         n38792, n38793, n38794, n38795, n38796, n38797, n38798, n38799,
         n38800, n38801, n38802, n38803, n38804, n38805, n38806, n38807,
         n38808, n38809, n38810, n38811, n38812, n38813, n38814, n38815,
         n38816, n38817, n38818, n38819, n38820, n38821, n38823, n38824,
         n38825, n38826, n38828, n38829, n38830, n38831, n38832, n38833,
         n38834, n38835, n38836, n38837, n38838, n38839, n38840, n38841,
         n38842, n38843, n38844, n38845, n38846, n38847, n38848, n38849,
         n38850, n38851, n38852, n38853, n38854, n38855, n38856, n38857,
         n38858, n38859, n38860, n38861, n38862, n38863, n38864, n38865,
         n38866, n38867, n38868, n38869, n38870, n38871, n38872, n38873,
         n38874, n38877, n38878, n38880, n38881, n38882, n38883, n38884,
         n38885, n38886, n38887, n38888, n38889, n38890, n38891, n38892,
         n38893, n38894, n38895, n38896, n38897, n38898, n38899, n38900,
         n38901, n38902, n38903, n38904, n38905, n38906, n38907, n38908,
         n38909, n38910, n38911, n38912, n38913, n38914, n38915, n38916,
         n38917, n38918, n38919, n38920, n38921, n38922, n38923, n38924,
         n38925, n38926, n38927, n38928, n38929, n38930, n38931, n38932,
         n38933, n38934, n38935, n38936, n38938, n38939, n38940, n38941,
         n38942, n38943, n38944, n38945, n38946, n38947, n38948, n38949,
         n38950, n38951, n38952, n38953, n38954, n38955, n38956, n38957,
         n38958, n38959, n38960, n38961, n38962, n38963, n38964, n38966,
         n38967, n38968, n38969, n38970, n38971, n38972, n38973, n38974,
         n38975, n38976, n38977, n38978, n38979, n38980, n38981, n38982,
         n38983, n38984, n38985, n38986, n38987, n38988, n38989, n38990,
         n38991, n38992, n38993, n38994, n38995, n38996, n38997, n38998,
         n38999, n39000, n39001, n39002, n39003, n39004, n39005, n39006,
         n39007, n39008, n39009, n39010, n39011, n39012, n39013, n39014,
         n39015, n39016, n39017, n39018, n39019, n39021, n39022, n39023,
         n39025, n39026, n39028, n39029, n39030, n39032, n39033, n39034,
         n39035, n39036, n39037, n39038, n39039, n39040, n39041, n39042,
         n39043, n39044, n39045, n39046, n39047, n39048, n39049, n39050,
         n39051, n39052, n39053, n39054, n39055, n39056, n39057, n39058,
         n39059, n39060, n39062, n39063, n39064, n39065, n39066, n39067,
         n39068, n39069, n39070, n39071, n39072, n39073, n39074, n39076,
         n39077, n39078, n39079, n39080, n39081, n39082, n39083, n39084,
         n39086, n39087, n39088, n39089, n39090, n39091, n39092, n39093,
         n39094, n39095, n39096, n39097, n39098, n39099, n39100, n39101,
         n39102, n39103, n39104, n39106, n39107, n39109, n39110, n39111,
         n39112, n39113, n39114, n39115, n39116, n39117, n39118, n39119,
         n39120, n39123, n39124, n39125, n39126, n39127, n39128, n39129,
         n39130, n39131, n39132, n39133, n39134, n39135, n39136, n39137,
         n39139, n39140, n39141, n39142, n39143, n39144, n39145, n39146,
         n39147, n39148, n39149, n39150, n39151, n39152, n39153, n39156,
         n39158, n39159, n39160, n39161, n39162, n39163, n39164, n39165,
         n39166, n39167, n39168, n39169, n39170, n39171, n39172, n39173,
         n39175, n39176, n39177, n39178, n39179, n39180, n39181, n39182,
         n39183, n39184, n39185, n39186, n39187, n39188, n39189, n39190,
         n39191, n39192, n39193, n39194, n39195, n39196, n39197, n39198,
         n39199, n39200, n39201, n39202, n39203, n39204, n39205, n39206,
         n39207, n39208, n39209, n39210, n39211, n39212, n39213, n39214,
         n39215, n39216, n39217, n39218, n39219, n39220, n39221, n39222,
         n39223, n39224, n39225, n39226, n39227, n39228, n39230, n39231,
         n39232, n39233, n39234, n39235, n39237, n39238, n39239, n39240,
         n39241, n39242, n39243, n39244, n39245, n39246, n39247, n39248,
         n39249, n39250, n39251, n39252, n39253, n39254, n39255, n39256,
         n39257, n39258, n39259, n39260, n39261, n39262, n39263, n39264,
         n39265, n39267, n39268, n39269, n39270, n39271, n39272, n39273,
         n39274, n39275, n39276, n39277, n39278, n39279, n39280, n39281,
         n39282, n39283, n39284, n39285, n39286, n39287, n39288, n39289,
         n39290, n39291, n39292, n39293, n39294, n39295, n39296, n39297,
         n39298, n39299, n39300, n39301, n39302, n39303, n39304, n39305,
         n39306, n39307, n39308, n39309, n39310, n39311, n39312, n39313,
         n39314, n39315, n39317, n39318, n39319, n39320, n39321, n39322,
         n39323, n39324, n39325, n39326, n39327, n39328, n39329, n39330,
         n39331, n39332, n39333, n39334, n39335, n39336, n39337, n39338,
         n39339, n39341, n39342, n39343, n39344, n39345, n39346, n39347,
         n39348, n39349, n39350, n39351, n39352, n39353, n39354, n39357,
         n39358, n39359, n39360, n39361, n39362, n39363, n39364, n39365,
         n39366, n39367, n39368, n39369, n39371, n39372, n39373, n39374,
         n39375, n39376, n39377, n39378, n39379, n39380, n39382, n39383,
         n39384, n39385, n39386, n39387, n39388, n39389, n39390, n39391,
         n39392, n39393, n39394, n39395, n39396, n39397, n39398, n39399,
         n39400, n39401, n39402, n39403, n39404, n39405, n39406, n39407,
         n39408, n39409, n39410, n39411, n39412, n39413, n39414, n39415,
         n39416, n39417, n39418, n39419, n39420, n39421, n39423, n39424,
         n39425, n39426, n39427, n39428, n39429, n39430, n39431, n39432,
         n39433, n39434, n39435, n39436, n39437, n39438, n39439, n39441,
         n39442, n39443, n39444, n39445, n39446, n39447, n39448, n39449,
         n39450, n39451, n39452, n39453, n39454, n39455, n39456, n39457,
         n39458, n39459, n39460, n39461, n39462, n39463, n39464, n39465,
         n39466, n39467, n39468, n39469, n39470, n39471, n39472, n39473,
         n39475, n39476, n39477, n39478, n39479, n39480, n39481, n39482,
         n39485, n39486, n39487, n39488, n39489, n39490, n39491, n39492,
         n39493, n39494, n39495, n39496, n39497, n39498, n39501, n39502,
         n39503, n39504, n39505, n39506, n39507, n39508, n39509, n39510,
         n39511, n39512, n39513, n39514, n39515, n39516, n39517, n39520,
         n39521, n39522, n39523, n39524, n39525, n39526, n39527, n39528,
         n39529, n39530, n39531, n39532, n39533, n39534, n39535, n39536,
         n39537, n39538, n39539, n39540, n39541, n39542, n39543, n39544,
         n39545, n39547, n39549, n39550, n39551, n39552, n39553, n39554,
         n39555, n39556, n39557, n39558, n39559, n39560, n39561, n39562,
         n39563, n39564, n39565, n39566, n39567, n39568, n39569, n39570,
         n39571, n39572, n39573, n39574, n39575, n39576, n39577, n39578,
         n39579, n39581, n39582, n39583, n39584, n39585, n39586, n39587,
         n39589, n39590, n39591, n39592, n39593, n39594, n39595, n39596,
         n39597, n39598, n39599, n39600, n39601, n39602, n39603, n39604,
         n39605, n39606, n39607, n39608, n39609, n39610, n39611, n39612,
         n39613, n39614, n39615, n39616, n39617, n39618, n39619, n39621,
         n39622, n39623, n39624, n39625, n39626, n39627, n39628, n39629,
         n39630, n39631, n39632, n39633, n39634, n39635, n39636, n39637,
         n39638, n39639, n39640, n39642, n39643, n39644, n39645, n39646,
         n39647, n39648, n39649, n39650, n39651, n39652, n39653, n39655,
         n39656, n39657, n39658, n39659, n39660, n39661, n39663, n39664,
         n39665, n39666, n39667, n39668, n39669, n39670, n39671, n39672,
         n39673, n39674, n39675, n39676, n39677, n39678, n39680, n39681,
         n39682, n39683, n39684, n39685, n39687, n39688, n39689, n39690,
         n39691, n39692, n39694, n39695, n39696, n39697, n39698, n39699,
         n39700, n39702, n39703, n39704, n39705, n39706, n39707, n39708,
         n39709, n39710, n39711, n39712, n39713, n39714, n39715, n39716,
         n39719, n39720, n39721, n39722, n39723, n39724, n39725, n39726,
         n39727, n39728, n39729, n39730, n39731, n39732, n39733, n39734,
         n39735, n39736, n39737, n39738, n39739, n39740, n39741, n39742,
         n39743, n39744, n39745, n39746, n39747, n39749, n39750, n39751,
         n39752, n39753, n39755, n39756, n39757, n39758, n39759, n39760,
         n39761, n39762, n39763, n39764, n39765, n39766, n39767, n39768,
         n39769, n39770, n39771, n39772, n39773, n39774, n39775, n39776,
         n39779, n39781, n39782, n39783, n39784, n39785, n39786, n39787,
         n39788, n39789, n39791, n39792, n39793, n39794, n39795, n39796,
         n39797, n39798, n39799, n39800, n39801, n39802, n39803, n39804,
         n39805, n39806, n39808, n39809, n39810, n39811, n39812, n39813,
         n39814, n39815, n39816, n39817, n39818, n39819, n39820, n39821,
         n39822, n39823, n39824, n39826, n39827, n39828, n39829, n39830,
         n39831, n39832, n39833, n39834, n39835, n39836, n39837, n39838,
         n39839, n39841, n39842, n39843, n39844, n39845, n39846, n39847,
         n39848, n39849, n39850, n39851, n39852, n39853, n39854, n39856,
         n39857, n39858, n39859, n39860, n39861, n39862, n39863, n39864,
         n39865, n39866, n39867, n39868, n39869, n39870, n39871, n39872,
         n39873, n39874, n39875, n39876, n39877, n39878, n39879, n39880,
         n39881, n39882, n39883, n39885, n39886, n39887, n39888, n39890,
         n39891, n39893, n39894, n39895, n39896, n39897, n39898, n39899,
         n39900, n39901, n39902, n39903, n39904, n39905, n39906, n39907,
         n39908, n39909, n39910, n39911, n39912, n39914, n39915, n39916,
         n39917, n39918, n39919, n39920, n39921, n39922, n39923, n39924,
         n39926, n39928, n39929, n39930, n39931, n39932, n39933, n39934,
         n39935, n39936, n39937, n39938, n39939, n39940, n39941, n39942,
         n39943, n39944, n39945, n39946, n39947, n39948, n39949, n39950,
         n39951, n39952, n39953, n39954, n39955, n39956, n39957, n39958,
         n39959, n39960, n39961, n39962, n39964, n39965, n39966, n39967,
         n39968, n39970, n39971, n39972, n39973, n39974, n39975, n39976,
         n39977, n39978, n39979, n39980, n39981, n39982, n39983, n39984,
         n39985, n39986, n39987, n39988, n39990, n39992, n39993, n39994,
         n39995, n39997, n39998, n39999, n40000, n40001, n40002, n40003,
         n40004, n40006, n40007, n40008, n40009, n40012, n40015, n40016,
         n40017, n40018, n40019, n40020, n40021, n40022, n40023, n40024,
         n40025, n40026, n40027, n40028, n40029, n40030, n40031, n40032,
         n40033, n40034, n40035, n40036, n40037, n40038, n40039, n40040,
         n40041, n40042, n40043, n40044, n40046, n40047, n40048, n40049,
         n40050, n40051, n40052, n40053, n40054, n40055, n40056, n40057,
         n40058, n40059, n40060, n40061, n40062, n40063, n40064, n40065,
         n40066, n40067, n40068, n40069, n40070, n40072, n40074, n40075,
         n40076, n40077, n40078, n40079, n40080, n40081, n40082, n40084,
         n40085, n40086, n40087, n40088, n40089, n40090, n40091, n40092,
         n40093, n40094, n40095, n40096, n40097, n40098, n40099, n40100,
         n40101, n40102, n40103, n40104, n40105, n40106, n40107, n40108,
         n40110, n40111, n40112, n40114, n40115, n40116, n40117, n40118,
         n40119, n40120, n40121, n40123, n40124, n40125, n40126, n40127,
         n40128, n40129, n40130, n40131, n40132, n40133, n40134, n40135,
         n40136, n40137, n40138, n40139, n40140, n40142, n40143, n40145,
         n40146, n40147, n40148, n40149, n40150, n40151, n40154, n40155,
         n40158, n40159, n40162, n40163, n40165, n40166, n40167, n40168,
         n40169, n40170, n40171, n40172, n40173, n40174, n40175, n40176,
         n40177, n40179, n40180, n40181, n40182, n40183, n40184, n40185,
         n40186, n40187, n40189, n40190, n40192, n40193, n40194, n40196,
         n40197, n40198, n40199, n40200, n40201, n40202, n40203, n40204,
         n40205, n40206, n40207, n40208, n40209, n40210, n40211, n40212,
         n40213, n40215, n40216, n40217, n40218, n40219, n40220, n40221,
         n40222, n40223, n40224, n40225, n40226, n40227, n40228, n40229,
         n40230, n40231, n40232, n40233, n40234, n40235, n40236, n40237,
         n40238, n40239, n40240, n40241, n40242, n40243, n40244, n40245,
         n40246, n40247, n40248, n40249, n40250, n40251, n40252, n40253,
         n40254, n40255, n40256, n40257, n40258, n40260, n40263, n40264,
         n40265, n40266, n40267, n40268, n40269, n40270, n40271, n40272,
         n40273, n40274, n40275, n40276, n40277, n40278, n40279, n40280,
         n40281, n40283, n40284, n40286, n40287, n40288, n40289, n40291,
         n40292, n40293, n40294, n40295, n40296, n40297, n40298, n40299,
         n40300, n40301, n40302, n40303, n40304, n40306, n40307, n40308,
         n40309, n40310, n40311, n40312, n40313, n40314, n40315, n40316,
         n40317, n40318, n40319, n40320, n40322, n40323, n40324, n40325,
         n40326, n40327, n40328, n40329, n40330, n40331, n40332, n40333,
         n40334, n40335, n40336, n40337, n40338, n40339, n40340, n40341,
         n40342, n40343, n40344, n40345, n40346, n40347, n40348, n40349,
         n40350, n40352, n40353, n40354, n40355, n40356, n40357, n40358,
         n40359, n40360, n40361, n40362, n40363, n40364, n40365, n40366,
         n40367, n40368, n40369, n40370, n40371, n40372, n40373, n40374,
         n40375, n40376, n40377, n40378, n40379, n40380, n40381, n40382,
         n40383, n40384, n40385, n40386, n40387, n40388, n40389, n40390,
         n40391, n40392, n40393, n40394, n40395, n40396, n40397, n40398,
         n40400, n40401, n40402, n40403, n40404, n40405, n40406, n40408,
         n40409, n40410, n40411, n40412, n40413, n40414, n40415, n40416,
         n40417, n40420, n40421, n40422, n40423, n40424, n40425, n40427,
         n40428, n40429, n40430, n40431, n40432, n40433, n40434, n40435,
         n40437, n40438, n40439, n40441, n40443, n40444, n40445, n40446,
         n40447, n40448, n40449, n40450, n40451, n40452, n40453, n40454,
         n40456, n40457, n40458, n40459, n40460, n40461, n40462, n40463,
         n40464, n40465, n40466, n40468, n40469, n40470, n40471, n40472,
         n40473, n40474, n40475, n40476, n40477, n40478, n40479, n40481,
         n40482, n40484, n40485, n40486, n40487, n40488, n40489, n40490,
         n40491, n40492, n40493, n40494, n40495, n40497, n40498, n40499,
         n40500, n40501, n40502, n40503, n40507, n40508, n40509, n40511,
         n40512, n40513, n40514, n40515, n40516, n40517, n40518, n40519,
         n40520, n40521, n40522, n40523, n40524, n40525, n40526, n40527,
         n40528, n40529, n40530, n40531, n40532, n40533, n40534, n40535,
         n40536, n40537, n40538, n40539, n40540, n40541, n40542, n40543,
         n40544, n40545, n40546, n40547, n40548, n40549, n40550, n40551,
         n40552, n40553, n40554, n40556, n40557, n40558, n40559, n40560,
         n40561, n40563, n40564, n40565, n40568, n40569, n40570, n40571,
         n40572, n40573, n40575, n40576, n40577, n40578, n40579, n40580,
         n40581, n40582, n40583, n40584, n40585, n40586, n40587, n40588,
         n40589, n40590, n40591, n40592, n40593, n40595, n40596, n40597,
         n40598, n40599, n40600, n40601, n40602, n40603, n40604, n40605,
         n40606, n40607, n40608, n40609, n40611, n40612, n40613, n40614,
         n40615, n40616, n40617, n40618, n40619, n40622, n40623, n40625,
         n40626, n40627, n40628, n40629, n40631, n40633, n40634, n40635,
         n40636, n40638, n40639, n40641, n40642, n40643, n40644, n40645,
         n40646, n40647, n40648, n40649, n40650, n40651, n40653, n40654,
         n40655, n40656, n40657, n40658, n40659, n40661, n40662, n40663,
         n40664, n40665, n40666, n40667, n40668, n40669, n40670, n40671,
         n40673, n40674, n40675, n40676, n40677, n40678, n40680, n40682,
         n40683, n40685, n40686, n40687, n40688, n40689, n40690, n40691,
         n40692, n40693, n40694, n40695, n40696, n40697, n40698, n40699,
         n40700, n40701, n40702, n40703, n40704, n40705, n40706, n40707,
         n40708, n40709, n40710, n40711, n40712, n40713, n40714, n40716,
         n40717, n40718, n40720, n40721, n40722, n40723, n40724, n40726,
         n40727, n40728, n40729, n40731, n40732, n40733, n40734, n40737,
         n40738, n40741, n40742, n40744, n40745, n40746, n40747, n40748,
         n40749, n40750, n40751, n40752, n40753, n40754, n40755, n40756,
         n40758, n40759, n40760, n40761, n40763, n40764, n40765, n40766,
         n40767, n40768, n40769, n40770, n40771, n40772, n40773, n40774,
         n40775, n40776, n40777, n40778, n40779, n40780, n40781, n40782,
         n40783, n40784, n40785, n40786, n40787, n40788, n40789, n40790,
         n40791, n40792, n40794, n40797, n40798, n40799, n40800, n40801,
         n40802, n40803, n40804, n40805, n40806, n40807, n40808, n40810,
         n40812, n40813, n40814, n40815, n40817, n40818, n40819, n40820,
         n40821, n40822, n40823, n40824, n40825, n40826, n40829, n40830,
         n40831, n40832, n40833, n40834, n40835, n40836, n40837, n40839,
         n40840, n40841, n40842, n40843, n40844, n40845, n40846, n40847,
         n40848, n40849, n40850, n40851, n40852, n40853, n40854, n40855,
         n40856, n40857, n40858, n40860, n40862, n40863, n40864, n40865,
         n40866, n40867, n40868, n40869, n40870, n40872, n40873, n40874,
         n40875, n40876, n40877, n40878, n40879, n40880, n40881, n40882,
         n40883, n40884, n40885, n40886, n40887, n40888, n40889, n40890,
         n40891, n40893, n40894, n40895, n40896, n40897, n40898, n40899,
         n40900, n40901, n40902, n40903, n40904, n40905, n40906, n40908,
         n40909, n40910, n40911, n40912, n40913, n40914, n40915, n40916,
         n40917, n40918, n40919, n40920, n40921, n40922, n40923, n40924,
         n40925, n40928, n40929, n40930, n40931, n40932, n40933, n40934,
         n40935, n40936, n40937, n40938, n40939, n40941, n40942, n40943,
         n40944, n40946, n40947, n40948, n40949, n40951, n40952, n40954,
         n40955, n40956, n40957, n40958, n40959, n40960, n40961, n40962,
         n40963, n40964, n40965, n40966, n40967, n40968, n40969, n40970,
         n40971, n40972, n40973, n40974, n40975, n40976, n40977, n40979,
         n40980, n40982, n40983, n40984, n40985, n40986, n40987, n40989,
         n40990, n40991, n40992, n40993, n40994, n40995, n40996, n40997,
         n40998, n40999, n41000, n41001, n41002, n41003, n41004, n41006,
         n41007, n41009, n41012, n41013, n41014, n41015, n41016, n41017,
         n41019, n41020, n41021, n41022, n41023, n41024, n41025, n41026,
         n41027, n41028, n41029, n41030, n41031, n41032, n41033, n41034,
         n41035, n41036, n41037, n41038, n41039, n41040, n41041, n41042,
         n41043, n41044, n41045, n41046, n41047, n41048, n41049, n41051,
         n41052, n41053, n41054, n41055, n41056, n41057, n41058, n41059,
         n41060, n41061, n41062, n41063, n41064, n41065, n41066, n41067,
         n41069, n41072, n41073, n41074, n41075, n41076, n41077, n41078,
         n41079, n41080, n41081, n41082, n41083, n41084, n41085, n41086,
         n41087, n41088, n41089, n41090, n41091, n41092, n41093, n41094,
         n41096, n41097, n41098, n41099, n41100, n41101, n41102, n41103,
         n41105, n41106, n41107, n41108, n41109, n41110, n41111, n41112,
         n41113, n41115, n41116, n41117, n41118, n41119, n41120, n41121,
         n41122, n41123, n41124, n41125, n41126, n41127, n41128, n41129,
         n41131, n41132, n41133, n41134, n41135, n41136, n41137, n41138,
         n41139, n41140, n41141, n41142, n41144, n41145, n41146, n41147,
         n41148, n41149, n41150, n41152, n41153, n41154, n41155, n41156,
         n41157, n41158, n41159, n41160, n41161, n41162, n41163, n41164,
         n41165, n41166, n41167, n41168, n41169, n41170, n41171, n41172,
         n41173, n41174, n41175, n41176, n41177, n41178, n41179, n41180,
         n41181, n41182, n41183, n41184, n41185, n41186, n41187, n41188,
         n41189, n41190, n41191, n41192, n41193, n41194, n41195, n41197,
         n41198, n41199, n41200, n41204, n41205, n41206, n41207, n41208,
         n41209, n41210, n41211, n41212, n41213, n41214, n41215, n41216,
         n41217, n41219, n41220, n41222, n41223, n41224, n41225, n41226,
         n41228, n41229, n41230, n41231, n41232, n41234, n41235, n41236,
         n41237, n41238, n41239, n41240, n41241, n41242, n41243, n41244,
         n41245, n41246, n41247, n41248, n41249, n41250, n41251, n41252,
         n41253, n41254, n41255, n41256, n41257, n41258, n41259, n41260,
         n41261, n41262, n41263, n41264, n41267, n41269, n41270, n41271,
         n41272, n41273, n41274, n41275, n41276, n41277, n41278, n41279,
         n41280, n41281, n41282, n41283, n41285, n41286, n41287, n41288,
         n41289, n41290, n41291, n41292, n41293, n41294, n41295, n41296,
         n41297, n41298, n41299, n41300, n41301, n41302, n41303, n41304,
         n41305, n41306, n41307, n41308, n41310, n41311, n41312, n41313,
         n41314, n41316, n41318, n41319, n41320, n41321, n41322, n41323,
         n41324, n41325, n41326, n41327, n41328, n41329, n41330, n41331,
         n41333, n41334, n41335, n41336, n41337, n41338, n41339, n41340,
         n41341, n41342, n41343, n41344, n41345, n41346, n41347, n41348,
         n41349, n41350, n41351, n41352, n41353, n41354, n41355, n41356,
         n41357, n41358, n41359, n41360, n41361, n41362, n41363, n41364,
         n41365, n41366, n41367, n41368, n41369, n41370, n41371, n41372,
         n41374, n41375, n41376, n41377, n41378, n41379, n41380, n41381,
         n41382, n41383, n41384, n41385, n41386, n41387, n41388, n41389,
         n41390, n41391, n41392, n41393, n41394, n41395, n41396, n41397,
         n41399, n41400, n41401, n41402, n41403, n41404, n41405, n41408,
         n41409, n41410, n41411, n41412, n41413, n41414, n41415, n41417,
         n41418, n41419, n41420, n41422, n41423, n41424, n41425, n41426,
         n41427, n41428, n41429, n41430, n41431, n41432, n41433, n41434,
         n41435, n41436, n41437, n41438, n41439, n41440, n41441, n41442,
         n41443, n41444, n41445, n41446, n41447, n41448, n41449, n41450,
         n41451, n41452, n41453, n41454, n41455, n41456, n41457, n41458,
         n41459, n41460, n41461, n41462, n41463, n41464, n41465, n41466,
         n41467, n41469, n41470, n41471, n41472, n41473, n41474, n41476,
         n41477, n41478, n41479, n41480, n41481, n41482, n41483, n41484,
         n41485, n41486, n41487, n41488, n41489, n41490, n41491, n41492,
         n41494, n41495, n41496, n41497, n41498, n41499, n41500, n41501,
         n41503, n41504, n41505, n41506, n41507, n41509, n41510, n41511,
         n41512, n41513, n41514, n41515, n41516, n41517, n41518, n41519,
         n41520, n41521, n41522, n41523, n41524, n41525, n41526, n41527,
         n41528, n41529, n41530, n41531, n41532, n41533, n41534, n41535,
         n41536, n41537, n41538, n41539, n41540, n41541, n41542, n41543,
         n41544, n41545, n41546, n41547, n41548, n41549, n41550, n41551,
         n41553, n41554, n41555, n41556, n41557, n41558, n41559, n41560,
         n41561, n41562, n41563, n41564, n41565, n41566, n41567, n41568,
         n41570, n41571, n41574, n41575, n41576, n41577, n41579, n41581,
         n41582, n41583, n41584, n41585, n41587, n41588, n41589, n41591,
         n41592, n41593, n41594, n41595, n41596, n41597, n41598, n41599,
         n41600, n41601, n41602, n41603, n41604, n41605, n41606, n41607,
         n41610, n41611, n41612, n41613, n41614, n41615, n41616, n41617,
         n41619, n41620, n41621, n41622, n41624, n41625, n41626, n41627,
         n41628, n41629, n41630, n41631, n41632, n41633, n41634, n41635,
         n41636, n41637, n41638, n41639, n41640, n41641, n41642, n41643,
         n41644, n41645, n41646, n41647, n41648, n41649, n41650, n41651,
         n41652, n41653, n41654, n41655, n41656, n41657, n41658, n41659,
         n41660, n41661, n41662, n41663, n41665, n41666, n41668, n41669,
         n41670, n41672, n41673, n41674, n41675, n41676, n41677, n41678,
         n41679, n41680, n41682, n41683, n41684, n41685, n41686, n41688,
         n41689, n41690, n41691, n41692, n41693, n41694, n41695, n41696,
         n41697, n41698, n41699, n41700, n41701, n41702, n41703, n41704,
         n41705, n41706, n41707, n41708, n41710, n41711, n41712, n41713,
         n41714, n41715, n41716, n41717, n41718, n41719, n41720, n41721,
         n41722, n41724, n41725, n41726, n41727, n41728, n41729, n41730,
         n41732, n41733, n41734, n41735, n41736, n41737, n41738, n41739,
         n41740, n41741, n41742, n41743, n41744, n41745, n41747, n41748,
         n41749, n41751, n41752, n41753, n41754, n41755, n41756, n41757,
         n41758, n41759, n41762, n41764, n41765, n41766, n41767, n41768,
         n41769, n41770, n41772, n41773, n41775, n41777, n41778, n41779,
         n41780, n41781, n41782, n41783, n41784, n41785, n41786, n41787,
         n41788, n41789, n41790, n41791, n41792, n41793, n41794, n41795,
         n41796, n41797, n41798, n41799, n41800, n41801, n41802, n41803,
         n41804, n41805, n41806, n41807, n41808, n41809, n41810, n41811,
         n41812, n41813, n41814, n41816, n41817, n41818, n41819, n41820,
         n41821, n41822, n41823, n41824, n41825, n41827, n41828, n41830,
         n41831, n41832, n41833, n41834, n41835, n41836, n41837, n41838,
         n41839, n41840, n41842, n41843, n41844, n41845, n41846, n41847,
         n41849, n41850, n41851, n41852, n41853, n41854, n41855, n41856,
         n41857, n41858, n41859, n41861, n41862, n41863, n41865, n41866,
         n41867, n41868, n41869, n41870, n41871, n41872, n41873, n41874,
         n41875, n41876, n41877, n41879, n41880, n41881, n41882, n41883,
         n41884, n41885, n41886, n41887, n41888, n41889, n41890, n41891,
         n41892, n41893, n41894, n41895, n41896, n41897, n41898, n41899,
         n41900, n41901, n41902, n41903, n41904, n41906, n41907, n41908,
         n41909, n41910, n41911, n41912, n41914, n41915, n41916, n41918,
         n41919, n41920, n41921, n41922, n41923, n41924, n41925, n41926,
         n41928, n41929, n41930, n41931, n41932, n41933, n41934, n41935,
         n41936, n41937, n41938, n41940, n41941, n41942, n41943, n41944,
         n41945, n41946, n41947, n41948, n41949, n41950, n41951, n41952,
         n41953, n41954, n41955, n41956, n41958, n41959, n41961, n41962,
         n41963, n41964, n41965, n41966, n41967, n41968, n41969, n41970,
         n41971, n41972, n41973, n41974, n41975, n41976, n41977, n41979,
         n41980, n41981, n41982, n41983, n41984, n41985, n41986, n41987,
         n41988, n41989, n41990, n41991, n41995, n41996, n41997, n41998,
         n41999, n42001, n42003, n42004, n42006, n42007, n42008, n42009,
         n42010, n42011, n42012, n42013, n42014, n42015, n42016, n42017,
         n42018, n42019, n42020, n42021, n42022, n42023, n42024, n42025,
         n42026, n42027, n42028, n42029, n42030, n42031, n42032, n42033,
         n42034, n42035, n42036, n42037, n42038, n42040, n42041, n42042,
         n42043, n42044, n42045, n42046, n42049, n42050, n42051, n42053,
         n42054, n42055, n42056, n42057, n42058, n42059, n42060, n42061,
         n42062, n42063, n42064, n42065, n42066, n42067, n42068, n42069,
         n42070, n42071, n42072, n42073, n42074, n42075, n42076, n42077,
         n42078, n42079, n42080, n42081, n42082, n42084, n42085, n42086,
         n42087, n42088, n42089, n42090, n42091, n42092, n42093, n42094,
         n42095, n42096, n42097, n42098, n42099, n42100, n42101, n42102,
         n42103, n42104, n42105, n42107, n42108, n42110, n42111, n42112,
         n42113, n42115, n42117, n42118, n42119, n42120, n42121, n42122,
         n42123, n42124, n42125, n42126, n42127, n42128, n42129, n42130,
         n42131, n42132, n42133, n42135, n42136, n42137, n42138, n42139,
         n42140, n42141, n42142, n42143, n42146, n42147, n42148, n42149,
         n42150, n42151, n42152, n42153, n42154, n42155, n42156, n42157,
         n42158, n42159, n42160, n42161, n42162, n42163, n42164, n42165,
         n42166, n42167, n42168, n42169, n42170, n42171, n42172, n42174,
         n42175, n42176, n42177, n42178, n42179, n42180, n42181, n42184,
         n42185, n42186, n42187, n42188, n42189, n42190, n42191, n42194,
         n42195, n42196, n42197, n42198, n42199, n42200, n42201, n42202,
         n42203, n42204, n42205, n42207, n42208, n42209, n42210, n42211,
         n42213, n42214, n42215, n42216, n42217, n42218, n42219, n42220,
         n42221, n42222, n42223, n42224, n42225, n42226, n42227, n42228,
         n42230, n42231, n42232, n42233, n42234, n42235, n42236, n42237,
         n42238, n42239, n42240, n42242, n42243, n42244, n42245, n42247,
         n42248, n42249, n42251, n42252, n42253, n42254, n42255, n42256,
         n42257, n42258, n42259, n42260, n42261, n42262, n42263, n42264,
         n42265, n42266, n42267, n42268, n42269, n42270, n42271, n42273,
         n42275, n42276, n42277, n42278, n42279, n42280, n42281, n42282,
         n42283, n42284, n42285, n42286, n42287, n42288, n42289, n42290,
         n42291, n42292, n42293, n42294, n42295, n42296, n42298, n42299,
         n42300, n42301, n42302, n42303, n42304, n42305, n42306, n42307,
         n42308, n42309, n42310, n42311, n42312, n42313, n42314, n42316,
         n42317, n42318, n42319, n42320, n42321, n42322, n42323, n42324,
         n42325, n42326, n42327, n42328, n42329, n42330, n42331, n42332,
         n42333, n42334, n42336, n42337, n42338, n42339, n42340, n42341,
         n42342, n42343, n42344, n42345, n42346, n42347, n42348, n42349,
         n42350, n42351, n42352, n42353, n42354, n42355, n42356, n42357,
         n42358, n42359, n42360, n42361, n42362, n42363, n42364, n42365,
         n42366, n42367, n42368, n42369, n42370, n42371, n42372, n42373,
         n42374, n42375, n42376, n42377, n42378, n42379, n42380, n42381,
         n42382, n42383, n42384, n42385, n42386, n42387, n42388, n42389,
         n42390, n42391, n42392, n42393, n42394, n42395, n42396, n42397,
         n42398, n42399, n42400, n42401, n42402, n42403, n42404, n42405,
         n42406, n42407, n42408, n42409, n42410, n42411, n42412, n42413,
         n42414, n42415, n42416, n42417, n42418, n42419, n42420, n42421,
         n42422, n42423, n42424, n42425, n42426, n42427, n42428, n42429,
         n42430, n42431, n42432, n42433, n42434, n42435, n42436, n42437,
         n42438, n42439, n42441, n42442, n42443, n42444, n42446, n42447,
         n42448, n42449, n42450, n42451, n42452, n42453, n42454, n42455,
         n42457, n42458, n42460, n42461, n42463, n42464, n42465, n42466,
         n42467, n42468, n42470, n42471, n42472, n42473, n42474, n42475,
         n42476, n42477, n42478, n42479, n42480, n42481, n42482, n42483,
         n42484, n42485, n42486, n42487, n42488, n42489, n42490, n42491,
         n42492, n42493, n42494, n42495, n42496, n42497, n42498, n42499,
         n42500, n42501, n42502, n42503, n42504, n42505, n42506, n42507,
         n42508, n42509, n42510, n42511, n42512, n42513, n42514, n42515,
         n42516, n42517, n42518, n42519, n42520, n42521, n42522, n42523,
         n42524, n42526, n42527, n42528, n42529, n42530, n42531, n42532,
         n42533, n42534, n42535, n42536, n42537, n42538, n42539, n42540,
         n42541, n42542, n42543, n42544, n42545, n42546, n42548, n42549,
         n42550, n42551, n42552, n42553, n42554, n42555, n42556, n42557,
         n42558, n42559, n42560, n42562, n42563, n42564, n42565, n42566,
         n42567, n42568, n42569, n42571, n42572, n42573, n42574, n42575,
         n42576, n42577, n42578, n42579, n42580, n42581, n42583, n42584,
         n42585, n42586, n42587, n42588, n42589, n42590, n42591, n42592,
         n42593, n42594, n42595, n42596, n42597, n42598, n42599, n42600,
         n42601, n42602, n42604, n42605, n42606, n42607, n42608, n42609,
         n42610, n42611, n42612, n42613, n42614, n42615, n42617, n42618,
         n42619, n42620, n42621, n42622, n42623, n42624, n42625, n42626,
         n42627, n42628, n42629, n42630, n42631, n42633, n42634, n42635,
         n42636, n42638, n42639, n42640, n42641, n42642, n42643, n42644,
         n42645, n42646, n42648, n42650, n42651, n42652, n42653, n42654,
         n42655, n42656, n42657, n42658, n42659, n42660, n42661, n42662,
         n42663, n42664, n42665, n42666, n42667, n42668, n42669, n42670,
         n42671, n42672, n42673, n42674, n42675, n42676, n42677, n42678,
         n42679, n42680, n42681, n42682, n42683, n42684, n42685, n42686,
         n42687, n42688, n42689, n42690, n42691, n42692, n42693, n42694,
         n42695, n42696, n42697, n42698, n42699, n42700, n42701, n42702,
         n42703, n42704, n42705, n42707, n42708, n42709, n42710, n42711,
         n42712, n42713, n42714, n42715, n42716, n42717, n42718, n42719,
         n42720, n42721, n42723, n42724, n42725, n42726, n42730, n42731,
         n42732, n42733, n42734, n42735, n42736, n42737, n42738, n42739,
         n42740, n42741, n42742, n42743, n42744, n42745, n42746, n42747,
         n42748, n42749, n42750, n42751, n42752, n42753, n42754, n42755,
         n42756, n42757, n42758, n42759, n42760, n42761, n42762, n42763,
         n42764, n42765, n42766, n42767, n42768, n42769, n42770, n42771,
         n42772, n42775, n42776, n42777, n42778, n42779, n42780, n42781,
         n42782, n42783, n42784, n42785, n42786, n42787, n42788, n42789,
         n42790, n42792, n42794, n42796, n42797, n42798, n42799, n42800,
         n42801, n42802, n42803, n42804, n42805, n42806, n42807, n42808,
         n42809, n42810, n42812, n42813, n42814, n42815, n42816, n42819,
         n42821, n42822, n42823, n42824, n42825, n42826, n42827, n42829,
         n42830, n42831, n42832, n42833, n42834, n42835, n42836, n42837,
         n42838, n42839, n42840, n42841, n42842, n42843, n42844, n42845,
         n42846, n42847, n42848, n42849, n42850, n42852, n42853, n42854,
         n42855, n42856, n42857, n42858, n42860, n42861, n42863, n42864,
         n42865, n42866, n42867, n42868, n42869, n42870, n42871, n42872,
         n42873, n42874, n42875, n42876, n42877, n42878, n42879, n42881,
         n42882, n42883, n42884, n42885, n42887, n42888, n42889, n42890,
         n42891, n42892, n42893, n42894, n42895, n42896, n42898, n42899,
         n42900, n42901, n42902, n42903, n42904, n42905, n42907, n42908,
         n42909, n42910, n42911, n42912, n42913, n42914, n42915, n42916,
         n42917, n42918, n42919, n42920, n42921, n42922, n42923, n42924,
         n42925, n42926, n42927, n42928, n42929, n42930, n42931, n42932,
         n42934, n42935, n42936, n42937, n42938, n42939, n42940, n42941,
         n42942, n42943, n42944, n42945, n42946, n42947, n42948, n42949,
         n42950, n42951, n42952, n42953, n42954, n42955, n42956, n42957,
         n42958, n42959, n42960, n42962, n42963, n42964, n42965, n42966,
         n42967, n42968, n42969, n42970, n42971, n42972, n42973, n42974,
         n42975, n42976, n42978, n42979, n42980, n42982, n42983, n42984,
         n42985, n42986, n42987, n42988, n42989, n42990, n42991, n42993,
         n42994, n42995, n42996, n42997, n42998, n42999, n43000, n43001,
         n43002, n43003, n43004, n43005, n43006, n43007, n43008, n43009,
         n43010, n43011, n43012, n43013, n43014, n43015, n43016, n43017,
         n43018, n43019, n43020, n43021, n43022, n43023, n43024, n43025,
         n43026, n43027, n43028, n43029, n43030, n43031, n43032, n43034,
         n43035, n43036, n43037, n43038, n43039, n43040, n43041, n43042,
         n43043, n43044, n43045, n43048, n43049, n43050, n43051, n43052,
         n43053, n43054, n43055, n43056, n43057, n43058, n43059, n43060,
         n43061, n43062, n43063, n43064, n43065, n43066, n43067, n43068,
         n43069, n43070, n43072, n43074, n43076, n43077, n43078, n43079,
         n43080, n43081, n43082, n43084, n43085, n43086, n43087, n43088,
         n43089, n43090, n43091, n43092, n43093, n43094, n43096, n43097,
         n43098, n43099, n43100, n43101, n43102, n43104, n43105, n43106,
         n43107, n43108, n43109, n43110, n43111, n43112, n43113, n43114,
         n43115, n43116, n43117, n43118, n43119, n43120, n43121, n43122,
         n43123, n43124, n43125, n43126, n43127, n43128, n43129, n43130,
         n43131, n43132, n43133, n43134, n43135, n43136, n43137, n43138,
         n43139, n43140, n43141, n43142, n43143, n43144, n43145, n43146,
         n43147, n43148, n43149, n43150, n43151, n43153, n43154, n43155,
         n43156, n43157, n43158, n43159, n43161, n43162, n43163, n43164,
         n43165, n43166, n43167, n43168, n43169, n43170, n43172, n43173,
         n43175, n43176, n43177, n43178, n43180, n43181, n43182, n43183,
         n43184, n43185, n43187, n43188, n43189, n43190, n43191, n43192,
         n43193, n43194, n43195, n43196, n43197, n43198, n43199, n43200,
         n43202, n43203, n43205, n43206, n43207, n43208, n43209, n43210,
         n43212, n43213, n43214, n43215, n43217, n43218, n43219, n43220,
         n43222, n43223, n43224, n43225, n43226, n43227, n43228, n43229,
         n43230, n43231, n43232, n43233, n43234, n43235, n43236, n43237,
         n43240, n43241, n43242, n43243, n43244, n43245, n43246, n43247,
         n43248, n43249, n43250, n43251, n43252, n43253, n43254, n43255,
         n43256, n43257, n43258, n43259, n43260, n43261, n43262, n43263,
         n43264, n43265, n43266, n43268, n43269, n43270, n43271, n43272,
         n43273, n43275, n43276, n43277, n43278, n43279, n43280, n43281,
         n43282, n43283, n43284, n43285, n43286, n43288, n43289, n43290,
         n43291, n43292, n43294, n43295, n43296, n43297, n43298, n43299,
         n43300, n43301, n43302, n43303, n43304, n43305, n43306, n43307,
         n43308, n43309, n43310, n43311, n43312, n43313, n43314, n43315,
         n43316, n43317, n43318, n43319, n43320, n43321, n43322, n43323,
         n43324, n43325, n43326, n43327, n43328, n43329, n43330, n43331,
         n43332, n43333, n43334, n43335, n43336, n43337, n43338, n43339,
         n43341, n43342, n43343, n43344, n43345, n43346, n43347, n43348,
         n43349, n43350, n43351, n43352, n43353, n43354, n43355, n43356,
         n43357, n43358, n43359, n43360, n43361, n43362, n43363, n43364,
         n43365, n43366, n43368, n43369, n43370, n43371, n43372, n43373,
         n43374, n43375, n43376, n43377, n43378, n43379, n43380, n43381,
         n43382, n43383, n43384, n43386, n43387, n43389, n43390, n43391,
         n43392, n43393, n43394, n43395, n43396, n43398, n43399, n43400,
         n43401, n43402, n43403, n43404, n43405, n43406, n43407, n43408,
         n43409, n43410, n43412, n43413, n43414, n43415, n43416, n43417,
         n43418, n43421, n43422, n43423, n43424, n43425, n43426, n43427,
         n43428, n43429, n43430, n43431, n43432, n43433, n43434, n43435,
         n43436, n43437, n43438, n43439, n43440, n43441, n43443, n43444,
         n43445, n43446, n43447, n43448, n43449, n43450, n43451, n43452,
         n43453, n43454, n43455, n43456, n43457, n43458, n43459, n43460,
         n43462, n43463, n43464, n43465, n43466, n43467, n43468, n43469,
         n43470, n43471, n43472, n43473, n43474, n43475, n43476, n43477,
         n43478, n43479, n43480, n43481, n43482, n43483, n43484, n43485,
         n43486, n43487, n43489, n43490, n43491, n43492, n43493, n43494,
         n43495, n43496, n43497, n43498, n43499, n43502, n43504, n43505,
         n43506, n43507, n43508, n43509, n43510, n43511, n43513, n43514,
         n43515, n43516, n43517, n43518, n43521, n43523, n43525, n43526,
         n43527, n43528, n43530, n43531, n43532, n43533, n43534, n43535,
         n43536, n43537, n43538, n43539, n43540, n43541, n43542, n43543,
         n43544, n43545, n43546, n43547, n43548, n43549, n43550, n43551,
         n43552, n43553, n43554, n43555, n43556, n43557, n43558, n43559,
         n43560, n43561, n43563, n43564, n43565, n43566, n43567, n43568,
         n43569, n43570, n43571, n43572, n43573, n43574, n43575, n43576,
         n43577, n43578, n43579, n43580, n43581, n43582, n43583, n43584,
         n43585, n43586, n43587, n43588, n43589, n43590, n43591, n43592,
         n43593, n43594, n43595, n43596, n43597, n43598, n43599, n43600,
         n43601, n43602, n43603, n43605, n43606, n43607, n43608, n43609,
         n43610, n43611, n43612, n43614, n43615, n43616, n43617, n43618,
         n43620, n43621, n43622, n43623, n43624, n43625, n43626, n43627,
         n43629, n43630, n43631, n43633, n43634, n43635, n43636, n43637,
         n43638, n43639, n43640, n43641, n43642, n43643, n43644, n43645,
         n43646, n43647, n43648, n43649, n43651, n43652, n43653, n43654,
         n43655, n43656, n43657, n43658, n43659, n43661, n43662, n43663,
         n43664, n43665, n43666, n43667, n43668, n43669, n43670, n43671,
         n43672, n43673, n43674, n43675, n43676, n43677, n43678, n43679,
         n43680, n43681, n43682, n43683, n43684, n43686, n43687, n43688,
         n43689, n43690, n43691, n43692, n43693, n43694, n43695, n43696,
         n43697, n43698, n43699, n43700, n43701, n43702, n43703, n43704,
         n43705, n43708, n43709, n43710, n43711, n43712, n43713, n43714,
         n43715, n43716, n43717, n43718, n43719, n43720, n43721, n43722,
         n43723, n43724, n43725, n43726, n43727, n43728, n43729, n43730,
         n43731, n43732, n43733, n43734, n43735, n43736, n43737, n43738,
         n43741, n43742, n43743, n43745, n43746, n43747, n43748, n43749,
         n43750, n43751, n43752, n43753, n43754, n43756, n43757, n43758,
         n43759, n43760, n43761, n43762, n43763, n43764, n43766, n43768,
         n43769, n43770, n43771, n43772, n43773, n43774, n43775, n43776,
         n43777, n43778, n43779, n43780, n43781, n43782, n43783, n43784,
         n43785, n43786, n43787, n43788, n43789, n43790, n43791, n43792,
         n43793, n43794, n43795, n43796, n43797, n43798, n43799, n43800,
         n43801, n43802, n43803, n43804, n43805, n43806, n43807, n43808,
         n43809, n43810, n43811, n43814, n43815, n43816, n43817, n43818,
         n43819, n43820, n43821, n43822, n43823, n43825, n43826, n43827,
         n43828, n43829, n43830, n43831, n43833, n43834, n43836, n43837,
         n43839, n43840, n43841, n43842, n43843, n43844, n43845, n43846,
         n43847, n43848, n43849, n43850, n43851, n43852, n43853, n43854,
         n43855, n43856, n43857, n43858, n43859, n43860, n43861, n43862,
         n43863, n43864, n43865, n43866, n43867, n43868, n43869, n43870,
         n43871, n43872, n43873, n43874, n43875, n43877, n43878, n43880,
         n43881, n43882, n43883, n43884, n43885, n43886, n43887, n43889,
         n43890, n43891, n43892, n43893, n43894, n43895, n43896, n43897,
         n43898, n43899, n43900, n43901, n43902, n43903, n43904, n43905,
         n43906, n43907, n43908, n43909, n43910, n43911, n43912, n43913,
         n43914, n43915, n43916, n43917, n43918, n43919, n43920, n43921,
         n43922, n43923, n43924, n43925, n43926, n43927, n43928, n43929,
         n43930, n43931, n43932, n43933, n43934, n43935, n43936, n43937,
         n43938, n43939, n43940, n43941, n43942, n43944, n43945, n43946,
         n43947, n43948, n43949, n43950, n43951, n43953, n43954, n43955,
         n43956, n43957, n43958, n43959, n43960, n43961, n43962, n43963,
         n43964, n43965, n43966, n43967, n43968, n43969, n43970, n43971,
         n43972, n43973, n43974, n43975, n43976, n43977, n43978, n43979,
         n43980, n43981, n43982, n43983, n43984, n43985, n43986, n43987,
         n43988, n43989, n43990, n43991, n43992, n43993, n43994, n43995,
         n43996, n43997, n43998, n44000, n44001, n44002, n44003, n44004,
         n44005, n44006, n44007, n44008, n44009, n44011, n44013, n44014,
         n44015, n44016, n44017, n44018, n44020, n44021, n44022, n44023,
         n44024, n44025, n44026, n44027, n44028, n44029, n44030, n44031,
         n44032, n44033, n44034, n44035, n44036, n44037, n44038, n44039,
         n44040, n44041, n44042, n44043, n44044, n44045, n44046, n44047,
         n44048, n44049, n44050, n44051, n44052, n44053, n44054, n44055,
         n44056, n44057, n44058, n44059, n44060, n44061, n44062, n44063,
         n44064, n44065, n44066, n44067, n44068, n44069, n44070, n44071,
         n44072, n44073, n44074, n44075, n44076, n44077, n44078, n44079,
         n44080, n44081, n44082, n44083, n44084, n44085, n44086, n44087,
         n44088, n44089, n44090, n44091, n44092, n44093, n44094, n44095,
         n44096, n44097, n44098, n44099, n44100, n44101, n44102, n44103,
         n44104, n44105, n44107, n44108, n44109, n44110, n44111, n44112,
         n44113, n44114, n44115, n44116, n44117, n44118, n44119, n44120,
         n44121, n44122, n44123, n44124, n44125, n44126, n44127, n44128,
         n44129, n44130, n44131, n44132, n44133, n44134, n44135, n44137,
         n44138, n44139, n44140, n44141, n44142, n44143, n44144, n44145,
         n44147, n44148, n44149, n44150, n44151, n44152, n44153, n44154,
         n44155, n44156, n44157, n44158, n44159, n44160, n44161, n44162,
         n44163, n44164, n44165, n44166, n44167, n44168, n44169, n44170,
         n44171, n44172, n44173, n44174, n44175, n44176, n44177, n44178,
         n44179, n44180, n44181, n44182, n44183, n44184, n44185, n44186,
         n44187, n44188, n44190, n44191, n44192, n44193, n44194, n44195,
         n44196, n44197, n44198, n44199, n44200, n44201, n44202, n44203,
         n44204, n44205, n44206, n44207, n44208, n44211, n44212, n44213,
         n44214, n44215, n44216, n44217, n44218, n44219, n44220, n44222,
         n44223, n44224, n44225, n44226, n44227, n44228, n44229, n44230,
         n44231, n44232, n44233, n44234, n44235, n44236, n44237, n44238,
         n44239, n44240, n44241, n44242, n44243, n44244, n44245, n44246,
         n44247, n44248, n44249, n44250, n44252, n44253, n44254, n44255,
         n44256, n44257, n44258, n44260, n44261, n44262, n44263, n44264,
         n44265, n44266, n44267, n44268, n44269, n44270, n44271, n44272,
         n44273, n44274, n44275, n44276, n44277, n44278, n44279, n44281,
         n44282, n44283, n44284, n44285, n44286, n44287, n44289, n44290,
         n44291, n44292, n44293, n44294, n44296, n44297, n44298, n44299,
         n44300, n44301, n44302, n44303, n44304, n44307, n44309, n44310,
         n44311, n44312, n44313, n44314, n44315, n44316, n44317, n44318,
         n44319, n44321, n44322, n44323, n44324, n44325, n44326, n44328,
         n44329, n44330, n44331, n44332, n44333, n44334, n44336, n44337,
         n44338, n44339, n44340, n44341, n44342, n44343, n44344, n44345,
         n44346, n44347, n44348, n44350, n44351, n44352, n44353, n44354,
         n44355, n44356, n44357, n44358, n44359, n44360, n44362, n44363,
         n44364, n44365, n44366, n44367, n44368, n44369, n44370, n44371,
         n44372, n44373, n44374, n44375, n44376, n44377, n44378, n44379,
         n44380, n44381, n44382, n44383, n44384, n44385, n44386, n44387,
         n44388, n44389, n44390, n44391, n44392, n44393, n44394, n44395,
         n44397, n44398, n44399, n44400, n44401, n44402, n44403, n44404,
         n44405, n44406, n44407, n44408, n44409, n44410, n44411, n44412,
         n44413, n44414, n44415, n44416, n44417, n44418, n44419, n44420,
         n44421, n44422, n44424, n44425, n44426, n44427, n44428, n44429,
         n44430, n44431, n44432, n44433, n44434, n44435, n44436, n44437,
         n44438, n44439, n44440, n44441, n44442, n44443, n44444, n44445,
         n44446, n44447, n44448, n44450, n44451, n44452, n44453, n44454,
         n44455, n44456, n44457, n44458, n44459, n44460, n44461, n44462,
         n44463, n44464, n44465, n44466, n44467, n44468, n44469, n44470,
         n44471, n44472, n44473, n44474, n44475, n44476, n44477, n44478,
         n44479, n44480, n44483, n44484, n44485, n44486, n44487, n44488,
         n44489, n44490, n44491, n44492, n44493, n44494, n44495, n44496,
         n44497, n44498, n44499, n44501, n44502, n44503, n44504, n44505,
         n44506, n44507, n44508, n44509, n44510, n44511, n44512, n44513,
         n44514, n44515, n44516, n44517, n44518, n44519, n44520, n44523,
         n44524, n44526, n44527, n44528, n44529, n44530, n44531, n44532,
         n44533, n44534, n44535, n44536, n44537, n44538, n44539, n44540,
         n44541, n44542, n44543, n44544, n44545, n44546, n44547, n44548,
         n44549, n44550, n44551, n44552, n44553, n44554, n44556, n44557,
         n44558, n44559, n44560, n44562, n44563, n44564, n44565, n44566,
         n44567, n44568, n44569, n44570, n44572, n44573, n44575, n44576,
         n44577, n44578, n44579, n44580, n44581, n44582, n44583, n44584,
         n44585, n44586, n44587, n44588, n44589, n44590, n44591, n44592,
         n44593, n44594, n44595, n44596, n44597, n44598, n44599, n44600,
         n44601, n44602, n44603, n44604, n44606, n44607, n44608, n44609,
         n44610, n44611, n44612, n44613, n44614, n44615, n44616, n44617,
         n44618, n44619, n44620, n44621, n44622, n44623, n44624, n44625,
         n44626, n44627, n44628, n44629, n44630, n44631, n44632, n44633,
         n44634, n44635, n44636, n44637, n44638, n44639, n44640, n44641,
         n44642, n44643, n44645, n44646, n44647, n44649, n44651, n44652,
         n44653, n44654, n44655, n44657, n44658, n44660, n44661, n44662,
         n44663, n44664, n44665, n44666, n44667, n44668, n44669, n44670,
         n44671, n44672, n44674, n44675, n44677, n44678, n44679, n44680,
         n44681, n44682, n44683, n44684, n44685, n44686, n44687, n44688,
         n44689, n44690, n44692, n44694, n44698, n44699, n44700, n44702,
         n44703, n44704, n44705, n44706, n44707, n44708, n44709, n44710,
         n44711, n44713, n44714, n44715, n44716, n44717, n44718, n44719,
         n44720, n44721, n44722, n44723, n44724, n44725, n44726, n44727,
         n44728, n44729, n44730, n44731, n44732, n44733, n44734, n44735,
         n44736, n44738, n44739, n44740, n44741, n44742, n44743, n44744,
         n44745, n44746, n44747, n44748, n44749, n44750, n44751, n44752,
         n44753, n44754, n44755, n44757, n44758, n44759, n44760, n44761,
         n44762, n44763, n44764, n44766, n44767, n44768, n44769, n44770,
         n44771, n44773, n44774, n44775, n44776, n44777, n44778, n44779,
         n44780, n44781, n44782, n44783, n44784, n44785, n44786, n44787,
         n44788, n44789, n44790, n44791, n44792, n44793, n44794, n44795,
         n44796, n44797, n44798, n44800, n44802, n44803, n44804, n44805,
         n44806, n44807, n44808, n44809, n44810, n44811, n44812, n44813,
         n44814, n44815, n44816, n44817, n44819, n44820, n44821, n44822,
         n44823, n44824, n44825, n44826, n44827, n44828, n44829, n44830,
         n44831, n44832, n44833, n44834, n44835, n44836, n44837, n44838,
         n44839, n44840, n44841, n44842, n44843, n44844, n44845, n44846,
         n44847, n44848, n44849, n44850, n44851, n44852, n44853, n44854,
         n44856, n44857, n44858, n44859, n44860, n44861, n44862, n44863,
         n44864, n44865, n44866, n44868, n44871, n44872, n44874, n44876,
         n44877, n44878, n44879, n44880, n44881, n44883, n44885, n44886,
         n44887, n44888, n44889, n44890, n44891, n44892, n44893, n44894,
         n44895, n44896, n44897, n44898, n44899, n44900, n44901, n44902,
         n44903, n44904, n44905, n44906, n44907, n44908, n44909, n44910,
         n44911, n44912, n44913, n44914, n44915, n44916, n44917, n44918,
         n44919, n44920, n44921, n44922, n44923, n44924, n44925, n44926,
         n44927, n44928, n44929, n44930, n44931, n44932, n44933, n44934,
         n44935, n44936, n44937, n44938, n44939, n44940, n44941, n44942,
         n44943, n44944, n44945, n44946, n44947, n44948, n44949, n44950,
         n44951, n44952, n44953, n44954, n44955, n44956, n44957, n44959,
         n44960, n44961, n44962, n44963, n44964, n44965, n44966, n44967,
         n44968, n44969, n44970, n44971, n44972, n44973, n44974, n44976,
         n44977, n44978, n44979, n44980, n44981, n44982, n44983, n44984,
         n44985, n44986, n44987, n44988, n44989, n44990, n44991, n44992,
         n44993, n44994, n44995, n44996, n44997, n44998, n44999, n45000,
         n45001, n45002, n45003, n45004, n45006, n45007, n45008, n45009,
         n45010, n45011, n45012, n45013, n45014, n45015, n45016, n45017,
         n45018, n45019, n45020, n45021, n45022, n45024, n45025, n45026,
         n45027, n45028, n45029, n45030, n45031, n45032, n45033, n45035,
         n45036, n45037, n45038, n45039, n45040, n45041, n45042, n45043,
         n45044, n45045, n45046, n45047, n45048, n45049, n45050, n45051,
         n45052, n45053, n45054, n45055, n45057, n45058, n45059, n45060,
         n45061, n45062, n45063, n45064, n45065, n45066, n45067, n45068,
         n45069, n45070, n45071, n45074, n45075, n45076, n45077, n45078,
         n45079, n45080, n45081, n45082, n45083, n45084, n45085, n45086,
         n45087, n45088, n45089, n45090, n45091, n45092, n45093, n45094,
         n45095, n45096, n45097, n45098, n45099, n45100, n45101, n45102,
         n45103, n45104, n45105, n45106, n45107, n45108, n45110, n45111,
         n45112, n45113, n45114, n45115, n45116, n45117, n45119, n45120,
         n45121, n45122, n45123, n45124, n45125, n45126, n45127, n45128,
         n45129, n45130, n45131, n45132, n45133, n45134, n45135, n45136,
         n45137, n45138, n45139, n45140, n45141, n45142, n45143, n45144,
         n45145, n45146, n45147, n45148, n45149, n45150, n45151, n45152,
         n45153, n45154, n45155, n45156, n45157, n45158, n45159, n45160,
         n45161, n45162, n45163, n45164, n45165, n45166, n45167, n45170,
         n45171, n45172, n45173, n45174, n45175, n45176, n45177, n45178,
         n45179, n45181, n45182, n45183, n45184, n45185, n45186, n45187,
         n45188, n45189, n45190, n45191, n45192, n45193, n45194, n45195,
         n45196, n45197, n45198, n45199, n45200, n45201, n45202, n45203,
         n45204, n45205, n45206, n45207, n45208, n45209, n45210, n45211,
         n45212, n45213, n45214, n45215, n45216, n45218, n45219, n45220,
         n45221, n45222, n45223, n45224, n45225, n45226, n45227, n45229,
         n45231, n45233, n45234, n45235, n45236, n45237, n45238, n45239,
         n45240, n45241, n45242, n45243, n45244, n45245, n45246, n45247,
         n45249, n45250, n45251, n45252, n45253, n45254, n45255, n45256,
         n45257, n45258, n45259, n45260, n45261, n45262, n45263, n45264,
         n45265, n45267, n45269, n45270, n45271, n45274, n45275, n45276,
         n45277, n45278, n45279, n45280, n45281, n45282, n45284, n45285,
         n45286, n45287, n45288, n45289, n45290, n45291, n45293, n45294,
         n45295, n45296, n45297, n45298, n45299, n45300, n45301, n45302,
         n45303, n45304, n45306, n45308, n45309, n45310, n45311, n45312,
         n45313, n45314, n45315, n45316, n45317, n45318, n45319, n45320,
         n45321, n45322, n45323, n45324, n45325, n45326, n45327, n45328,
         n45329, n45330, n45331, n45332, n45333, n45334, n45335, n45336,
         n45337, n45338, n45339, n45340, n45341, n45342, n45343, n45344,
         n45345, n45346, n45347, n45348, n45349, n45350, n45351, n45352,
         n45353, n45354, n45355, n45356, n45357, n45358, n45359, n45360,
         n45361, n45362, n45363, n45364, n45365, n45366, n45367, n45368,
         n45370, n45371, n45372, n45373, n45375, n45376, n45377, n45378,
         n45379, n45380, n45381, n45382, n45383, n45385, n45386, n45387,
         n45388, n45389, n45390, n45391, n45392, n45393, n45394, n45395,
         n45396, n45397, n45398, n45399, n45400, n45401, n45402, n45403,
         n45404, n45405, n45406, n45407, n45408, n45409, n45411, n45412,
         n45413, n45414, n45416, n45417, n45418, n45419, n45420, n45421,
         n45422, n45423, n45424, n45425, n45426, n45427, n45428, n45429,
         n45430, n45431, n45432, n45433, n45434, n45435, n45436, n45437,
         n45438, n45439, n45440, n45442, n45443, n45444, n45445, n45446,
         n45447, n45448, n45449, n45450, n45451, n45452, n45453, n45454,
         n45455, n45456, n45457, n45458, n45459, n45461, n45462, n45463,
         n45464, n45465, n45466, n45467, n45468, n45469, n45470, n45471,
         n45472, n45473, n45474, n45475, n45476, n45477, n45479, n45480,
         n45481, n45482, n45483, n45484, n45485, n45486, n45487, n45488,
         n45489, n45490, n45491, n45492, n45493, n45494, n45495, n45498,
         n45499, n45500, n45501, n45503, n45504, n45505, n45506, n45507,
         n45508, n45509, n45510, n45511, n45512, n45513, n45515, n45516,
         n45517, n45518, n45519, n45520, n45521, n45522, n45523, n45524,
         n45525, n45526, n45527, n45528, n45529, n45530, n45531, n45532,
         n45533, n45534, n45535, n45536, n45537, n45538, n45539, n45540,
         n45541, n45543, n45544, n45545, n45546, n45547, n45549, n45550,
         n45551, n45552, n45553, n45554, n45555, n45556, n45557, n45558,
         n45559, n45561, n45562, n45563, n45565, n45566, n45567, n45568,
         n45569, n45570, n45571, n45572, n45573, n45574, n45576, n45577,
         n45578, n45579, n45580, n45581, n45582, n45584, n45586, n45587,
         n45588, n45589, n45590, n45591, n45592, n45594, n45595, n45596,
         n45597, n45599, n45601, n45602, n45603, n45604, n45606, n45607,
         n45608, n45609, n45610, n45611, n45612, n45613, n45614, n45617,
         n45618, n45619, n45620, n45621, n45622, n45623, n45624, n45627,
         n45628, n45629, n45630, n45631, n45632, n45633, n45634, n45635,
         n45636, n45637, n45638, n45639, n45640, n45641, n45642, n45643,
         n45644, n45645, n45646, n45647, n45648, n45650, n45651, n45652,
         n45653, n45654, n45655, n45656, n45657, n45658, n45659, n45660,
         n45661, n45662, n45663, n45664, n45665, n45666, n45667, n45668,
         n45669, n45670, n45672, n45673, n45674, n45675, n45676, n45677,
         n45678, n45679, n45680, n45681, n45682, n45683, n45684, n45685,
         n45686, n45687, n45689, n45690, n45691, n45692, n45694, n45695,
         n45696, n45697, n45698, n45699, n45700, n45701, n45702, n45703,
         n45704, n45705, n45706, n45708, n45709, n45710, n45711, n45712,
         n45713, n45714, n45715, n45716, n45717, n45718, n45719, n45720,
         n45721, n45722, n45723, n45724, n45725, n45726, n45727, n45728,
         n45729, n45730, n45731, n45733, n45734, n45736, n45737, n45739,
         n45740, n45741, n45744, n45745, n45746, n45747, n45748, n45749,
         n45750, n45751, n45752, n45754, n45755, n45756, n45757, n45758,
         n45759, n45760, n45761, n45762, n45763, n45764, n45765, n45766,
         n45767, n45768, n45769, n45770, n45771, n45772, n45773, n45774,
         n45775, n45776, n45777, n45779, n45780, n45781, n45782, n45783,
         n45784, n45785, n45786, n45787, n45788, n45790, n45791, n45792,
         n45793, n45794, n45796, n45798, n45799, n45800, n45801, n45802,
         n45803, n45804, n45805, n45806, n45807, n45808, n45809, n45810,
         n45811, n45812, n45813, n45815, n45816, n45817, n45818, n45819,
         n45820, n45821, n45822, n45823, n45826, n45827, n45828, n45829,
         n45830, n45831, n45832, n45833, n45834, n45835, n45836, n45837,
         n45838, n45839, n45840, n45841, n45842, n45843, n45844, n45845,
         n45846, n45847, n45848, n45849, n45850, n45852, n45853, n45854,
         n45855, n45856, n45857, n45858, n45859, n45860, n45861, n45862,
         n45865, n45866, n45867, n45868, n45869, n45870, n45871, n45872,
         n45873, n45874, n45875, n45876, n45877, n45878, n45879, n45880,
         n45881, n45882, n45883, n45884, n45885, n45887, n45888, n45889,
         n45891, n45892, n45894, n45895, n45896, n45897, n45898, n45899,
         n45900, n45901, n45902, n45903, n45904, n45905, n45906, n45907,
         n45908, n45910, n45911, n45912, n45913, n45914, n45916, n45920,
         n45921, n45922, n45923, n45924, n45925, n45926, n45927, n45929,
         n45930, n45931, n45932, n45933, n45934, n45935, n45936, n45937,
         n45939, n45940, n45941, n45942, n45943, n45944, n45945, n45946,
         n45947, n45948, n45949, n45950, n45951, n45952, n45953, n45954,
         n45955, n45957, n45958, n45959, n45960, n45961, n45962, n45964,
         n45965, n45966, n45967, n45968, n45969, n45970, n45971, n45972,
         n45974, n45975, n45976, n45977, n45978, n45979, n45980, n45982,
         n45983, n45984, n45985, n45986, n45987, n45988, n45989, n45990,
         n45991, n45992, n45993, n45994, n45995, n45997, n45998, n45999,
         n46000, n46001, n46002, n46003, n46004, n46005, n46006, n46007,
         n46008, n46009, n46010, n46011, n46012, n46013, n46014, n46015,
         n46016, n46017, n46018, n46019, n46020, n46022, n46023, n46024,
         n46025, n46026, n46027, n46028, n46029, n46030, n46031, n46032,
         n46033, n46034, n46035, n46036, n46037, n46038, n46039, n46040,
         n46041, n46042, n46044, n46045, n46046, n46047, n46048, n46049,
         n46050, n46052, n46053, n46054, n46055, n46056, n46057, n46058,
         n46059, n46060, n46061, n46062, n46063, n46064, n46066, n46067,
         n46068, n46069, n46070, n46072, n46073, n46074, n46075, n46076,
         n46077, n46078, n46079, n46080, n46081, n46082, n46083, n46084,
         n46085, n46086, n46087, n46088, n46089, n46090, n46091, n46092,
         n46093, n46094, n46095, n46096, n46097, n46098, n46099, n46100,
         n46101, n46102, n46103, n46104, n46105, n46106, n46107, n46108,
         n46109, n46111, n46112, n46113, n46114, n46115, n46116, n46117,
         n46118, n46120, n46121, n46122, n46123, n46124, n46125, n46126,
         n46127, n46128, n46129, n46130, n46131, n46132, n46133, n46135,
         n46136, n46137, n46140, n46141, n46142, n46143, n46144, n46145,
         n46146, n46147, n46148, n46149, n46150, n46151, n46152, n46153,
         n46154, n46155, n46156, n46157, n46159, n46160, n46161, n46162,
         n46163, n46164, n46165, n46166, n46167, n46168, n46169, n46170,
         n46171, n46172, n46173, n46174, n46175, n46176, n46177, n46178,
         n46180, n46181, n46182, n46183, n46184, n46185, n46186, n46187,
         n46188, n46189, n46190, n46191, n46192, n46193, n46194, n46195,
         n46196, n46197, n46198, n46199, n46200, n46201, n46202, n46203,
         n46204, n46206, n46207, n46208, n46209, n46210, n46211, n46212,
         n46213, n46214, n46215, n46216, n46217, n46218, n46219, n46220,
         n46221, n46222, n46223, n46224, n46225, n46226, n46227, n46228,
         n46229, n46230, n46231, n46232, n46233, n46234, n46235, n46236,
         n46237, n46238, n46239, n46240, n46241, n46243, n46244, n46245,
         n46246, n46247, n46248, n46249, n46250, n46251, n46252, n46253,
         n46254, n46255, n46256, n46257, n46258, n46259, n46260, n46261,
         n46262, n46263, n46264, n46265, n46266, n46267, n46268, n46269,
         n46270, n46271, n46272, n46273, n46274, n46275, n46276, n46277,
         n46278, n46279, n46280, n46281, n46282, n46283, n46284, n46285,
         n46286, n46287, n46288, n46289, n46290, n46291, n46292, n46293,
         n46296, n46297, n46298, n46299, n46300, n46301, n46302, n46303,
         n46304, n46305, n46306, n46307, n46308, n46309, n46310, n46311,
         n46312, n46314, n46315, n46316, n46317, n46318, n46319, n46321,
         n46322, n46323, n46324, n46325, n46326, n46327, n46328, n46329,
         n46330, n46331, n46332, n46333, n46336, n46337, n46338, n46339,
         n46340, n46341, n46342, n46343, n46344, n46345, n46346, n46347,
         n46348, n46349, n46350, n46351, n46352, n46353, n46354, n46355,
         n46356, n46357, n46358, n46359, n46360, n46361, n46362, n46363,
         n46364, n46365, n46366, n46367, n46368, n46369, n46370, n46371,
         n46372, n46373, n46374, n46375, n46376, n46377, n46378, n46379,
         n46380, n46381, n46382, n46383, n46384, n46385, n46386, n46387,
         n46388, n46389, n46390, n46391, n46392, n46393, n46394, n46395,
         n46396, n46397, n46398, n46399, n46400, n46401, n46402, n46403,
         n46404, n46405, n46406, n46407, n46408, n46409, n46410, n46412,
         n46413, n46414, n46415, n46416, n46417, n46418, n46421, n46422,
         n46423, n46424, n46425, n46426, n46427, n46428, n46429, n46430,
         n46431, n46432, n46433, n46434, n46436, n46437, n46438, n46439,
         n46440, n46441, n46442, n46443, n46444, n46445, n46446, n46447,
         n46448, n46449, n46450, n46451, n46452, n46453, n46454, n46455,
         n46456, n46457, n46458, n46460, n46461, n46462, n46463, n46464,
         n46465, n46466, n46467, n46468, n46469, n46470, n46471, n46472,
         n46473, n46474, n46475, n46476, n46477, n46481, n46482, n46483,
         n46484, n46486, n46487, n46488, n46489, n46490, n46491, n46492,
         n46493, n46494, n46495, n46496, n46497, n46498, n46499, n46500,
         n46501, n46502, n46503, n46504, n46505, n46506, n46507, n46508,
         n46509, n46510, n46511, n46513, n46514, n46515, n46516, n46517,
         n46518, n46519, n46520, n46521, n46522, n46523, n46524, n46525,
         n46526, n46527, n46528, n46529, n46531, n46532, n46533, n46534,
         n46535, n46536, n46537, n46538, n46539, n46540, n46543, n46544,
         n46545, n46546, n46547, n46549, n46550, n46551, n46552, n46553,
         n46554, n46555, n46556, n46557, n46558, n46559, n46560, n46561,
         n46562, n46563, n46564, n46565, n46566, n46568, n46570, n46571,
         n46572, n46573, n46576, n46577, n46578, n46579, n46580, n46581,
         n46582, n46583, n46584, n46585, n46586, n46587, n46588, n46589,
         n46590, n46591, n46592, n46593, n46594, n46595, n46596, n46597,
         n46598, n46599, n46601, n46602, n46603, n46604, n46605, n46606,
         n46607, n46608, n46609, n46610, n46611, n46612, n46613, n46614,
         n46615, n46616, n46617, n46618, n46619, n46620, n46621, n46622,
         n46623, n46624, n46625, n46626, n46628, n46629, n46630, n46631,
         n46632, n46633, n46634, n46635, n46636, n46637, n46638, n46639,
         n46640, n46641, n46642, n46643, n46644, n46645, n46646, n46647,
         n46648, n46649, n46650, n46651, n46652, n46653, n46654, n46655,
         n46656, n46657, n46658, n46659, n46660, n46661, n46662, n46663,
         n46665, n46666, n46668, n46669, n46670, n46671, n46672, n46673,
         n46674, n46676, n46677, n46679, n46680, n46681, n46682, n46683,
         n46684, n46685, n46686, n46687, n46688, n46689, n46690, n46691,
         n46692, n46693, n46694, n46695, n46696, n46697, n46698, n46699,
         n46700, n46701, n46702, n46703, n46704, n46705, n46706, n46707,
         n46708, n46709, n46710, n46711, n46712, n46713, n46714, n46715,
         n46716, n46717, n46718, n46719, n46720, n46721, n46722, n46723,
         n46725, n46726, n46727, n46728, n46729, n46730, n46731, n46732,
         n46733, n46735, n46736, n46737, n46738, n46739, n46740, n46741,
         n46742, n46744, n46745, n46746, n46747, n46748, n46749, n46751,
         n46752, n46753, n46754, n46755, n46756, n46757, n46758, n46759,
         n46760, n46761, n46762, n46763, n46764, n46765, n46767, n46770,
         n46771, n46773, n46777, n46778, n46782, n46783, n46784, n46785,
         n46786, n46787, n46788, n46789, n46790, n46792, n46793, n46794,
         n46796, n46797, n46798, n46799, n46800, n46801, n46802, n46803,
         n46804, n46805, n46806, n46807, n46809, n46810, n46812, n46813,
         n46814, n46815, n46816, n46817, n46818, n46819, n46820, n46821,
         n46822, n46823, n46824, n46825, n46826, n46827, n46828, n46829,
         n46830, n46831, n46833, n46835, n46836, n46837, n46838, n46839,
         n46840, n46841, n46842, n46843, n46844, n46845, n46846, n46847,
         n46848, n46849, n46850, n46851, n46852, n46853, n46854, n46855,
         n46856, n46858, n46859, n46860, n46861, n46862, n46863, n46864,
         n46865, n46866, n46867, n46868, n46869, n46870, n46871, n46872,
         n46873, n46874, n46875, n46876, n46877, n46878, n46879, n46880,
         n46882, n46883, n46884, n46885, n46886, n46887, n46889, n46890,
         n46891, n46892, n46893, n46894, n46896, n46897, n46898, n46899,
         n46900, n46901, n46902, n46903, n46904, n46905, n46906, n46907,
         n46908, n46910, n46911, n46912, n46913, n46914, n46915, n46916,
         n46918, n46919, n46920, n46921, n46922, n46923, n46924, n46925,
         n46926, n46927, n46928, n46929, n46930, n46931, n46932, n46933,
         n46934, n46935, n46936, n46937, n46940, n46941, n46942, n46943,
         n46944, n46945, n46946, n46947, n46948, n46949, n46950, n46951,
         n46952, n46957, n46958, n46959, n46960, n46961, n46962, n46963,
         n46964, n46965, n46967, n46968, n46969, n46971, n46972, n46973,
         n46974, n46975, n46976, n46977, n46978, n46979, n46980, n46981,
         n46982, n46983, n46984, n46985, n46986, n46987, n46988, n46989,
         n46990, n46991, n46992, n46993, n46994, n46995, n46996, n46997,
         n46998, n46999, n47000, n47001, n47002, n47003, n47004, n47005,
         n47006, n47007, n47008, n47009, n47010, n47011, n47012, n47013,
         n47014, n47015, n47016, n47017, n47018, n47019, n47020, n47021,
         n47022, n47023, n47024, n47025, n47026, n47027, n47028, n47029,
         n47030, n47031, n47032, n47033, n47034, n47035, n47036, n47037,
         n47039, n47040, n47041, n47042, n47044, n47045, n47046, n47047,
         n47049, n47051, n47052, n47053, n47054, n47055, n47056, n47057,
         n47058, n47059, n47060, n47061, n47062, n47063, n47064, n47068,
         n47069, n47070, n47071, n47072, n47073, n47074, n47075, n47077,
         n47078, n47079, n47080, n47081, n47082, n47083, n47084, n47085,
         n47086, n47087, n47088, n47089, n47090, n47091, n47092, n47093,
         n47094, n47095, n47096, n47097, n47098, n47099, n47100, n47101,
         n47102, n47104, n47105, n47106, n47107, n47108, n47110, n47111,
         n47112, n47113, n47115, n47116, n47117, n47118, n47119, n47120,
         n47121, n47122, n47123, n47124, n47125, n47126, n47127, n47128,
         n47129, n47130, n47131, n47132, n47133, n47135, n47136, n47137,
         n47139, n47140, n47141, n47142, n47143, n47144, n47145, n47146,
         n47148, n47149, n47150, n47151, n47152, n47153, n47154, n47155,
         n47156, n47157, n47158, n47159, n47160, n47161, n47163, n47164,
         n47165, n47166, n47167, n47168, n47169, n47170, n47171, n47172,
         n47173, n47174, n47175, n47176, n47177, n47178, n47179, n47180,
         n47181, n47182, n47183, n47184, n47185, n47186, n47187, n47188,
         n47189, n47190, n47192, n47193, n47194, n47195, n47196, n47197,
         n47199, n47200, n47201, n47202, n47203, n47204, n47206, n47207,
         n47208, n47209, n47210, n47211, n47213, n47214, n47215, n47216,
         n47217, n47218, n47219, n47221, n47222, n47223, n47224, n47226,
         n47227, n47228, n47229, n47230, n47231, n47232, n47233, n47236,
         n47237, n47238, n47239, n47240, n47241, n47243, n47244, n47245,
         n47246, n47247, n47248, n47249, n47250, n47251, n47252, n47253,
         n47254, n47255, n47256, n47257, n47259, n47260, n47261, n47262,
         n47263, n47264, n47265, n47266, n47267, n47268, n47269, n47270,
         n47271, n47272, n47273, n47274, n47275, n47276, n47277, n47278,
         n47279, n47280, n47281, n47282, n47283, n47284, n47285, n47286,
         n47287, n47288, n47289, n47290, n47291, n47292, n47293, n47294,
         n47295, n47296, n47297, n47298, n47299, n47300, n47301, n47302,
         n47303, n47304, n47305, n47306, n47307, n47308, n47309, n47310,
         n47311, n47312, n47313, n47314, n47315, n47316, n47317, n47318,
         n47319, n47321, n47322, n47323, n47324, n47325, n47326, n47327,
         n47328, n47329, n47331, n47332, n47333, n47334, n47335, n47336,
         n47337, n47338, n47339, n47340, n47341, n47342, n47343, n47344,
         n47345, n47346, n47347, n47348, n47349, n47350, n47351, n47352,
         n47353, n47354, n47355, n47356, n47357, n47358, n47359, n47360,
         n47361, n47362, n47363, n47364, n47365, n47366, n47367, n47368,
         n47369, n47370, n47371, n47372, n47373, n47375, n47376, n47377,
         n47378, n47379, n47380, n47381, n47382, n47383, n47384, n47385,
         n47386, n47387, n47388, n47389, n47390, n47391, n47392, n47393,
         n47394, n47395, n47396, n47397, n47398, n47399, n47400, n47401,
         n47403, n47404, n47405, n47406, n47407, n47408, n47409, n47411,
         n47413, n47414, n47415, n47416, n47417, n47418, n47419, n47420,
         n47421, n47422, n47423, n47424, n47425, n47426, n47427, n47428,
         n47429, n47430, n47431, n47432, n47433, n47434, n47435, n47436,
         n47437, n47439, n47441, n47442, n47443, n47444, n47445, n47446,
         n47447, n47448, n47449, n47450, n47451, n47452, n47453, n47454,
         n47455, n47456, n47457, n47458, n47460, n47461, n47462, n47463,
         n47464, n47465, n47466, n47467, n47468, n47469, n47470, n47471,
         n47472, n47473, n47474, n47475, n47476, n47477, n47478, n47479,
         n47480, n47481, n47482, n47483, n47484, n47485, n47486, n47487,
         n47488, n47489, n47490, n47491, n47492, n47493, n47494, n47495,
         n47496, n47497, n47498, n47499, n47500, n47501, n47502, n47503,
         n47504, n47505, n47506, n47508, n47509, n47510, n47511, n47512,
         n47513, n47515, n47516, n47517, n47518, n47519, n47520, n47521,
         n47522, n47523, n47524, n47525, n47526, n47527, n47529, n47530,
         n47531, n47532, n47533, n47534, n47535, n47536, n47537, n47538,
         n47539, n47540, n47541, n47542, n47543, n47544, n47545, n47546,
         n47547, n47548, n47549, n47550, n47551, n47552, n47553, n47554,
         n47555, n47557, n47558, n47559, n47560, n47561, n47562, n47563,
         n47564, n47565, n47566, n47568, n47570, n47571, n47572, n47573,
         n47574, n47575, n47576, n47577, n47578, n47579, n47580, n47581,
         n47582, n47583, n47584, n47585, n47586, n47587, n47588, n47589,
         n47590, n47591, n47592, n47593, n47594, n47595, n47596, n47597,
         n47598, n47599, n47600, n47601, n47602, n47603, n47604, n47605,
         n47606, n47607, n47608, n47609, n47610, n47611, n47612, n47613,
         n47615, n47616, n47617, n47618, n47619, n47620, n47621, n47622,
         n47623, n47624, n47625, n47626, n47627, n47628, n47629, n47631,
         n47632, n47633, n47634, n47635, n47636, n47637, n47638, n47639,
         n47640, n47641, n47642, n47643, n47644, n47645, n47646, n47647,
         n47648, n47649, n47650, n47651, n47652, n47653, n47654, n47655,
         n47656, n47657, n47659, n47660, n47661, n47662, n47663, n47664,
         n47665, n47666, n47667, n47668, n47669, n47670, n47671, n47672,
         n47673, n47674, n47675, n47676, n47677, n47680, n47681, n47682,
         n47683, n47685, n47686, n47687, n47688, n47689, n47690, n47691,
         n47692, n47693, n47694, n47695, n47696, n47697, n47698, n47699,
         n47700, n47701, n47702, n47703, n47704, n47705, n47706, n47707,
         n47708, n47709, n47710, n47711, n47712, n47713, n47714, n47716,
         n47717, n47718, n47719, n47720, n47721, n47722, n47723, n47724,
         n47725, n47726, n47727, n47728, n47729, n47730, n47731, n47732,
         n47733, n47734, n47735, n47736, n47737, n47738, n47739, n47740,
         n47741, n47743, n47744, n47745, n47746, n47747, n47748, n47749,
         n47750, n47752, n47753, n47754, n47755, n47756, n47757, n47759,
         n47760, n47761, n47762, n47763, n47765, n47766, n47768, n47769,
         n47770, n47771, n47772, n47773, n47774, n47775, n47776, n47777,
         n47778, n47779, n47780, n47783, n47785, n47786, n47787, n47788,
         n47789, n47790, n47792, n47793, n47794, n47796, n47797, n47798,
         n47799, n47800, n47801, n47802, n47803, n47804, n47805, n47806,
         n47807, n47808, n47809, n47810, n47811, n47812, n47813, n47814,
         n47815, n47816, n47817, n47818, n47819, n47820, n47821, n47823,
         n47824, n47825, n47826, n47827, n47828, n47830, n47831, n47832,
         n47833, n47834, n47837, n47838, n47839, n47840, n47841, n47843,
         n47844, n47845, n47846, n47847, n47848, n47850, n47851, n47852,
         n47853, n47855, n47856, n47857, n47858, n47860, n47861, n47862,
         n47863, n47864, n47865, n47866, n47867, n47868, n47869, n47870,
         n47871, n47872, n47873, n47874, n47875, n47876, n47877, n47878,
         n47879, n47880, n47881, n47882, n47883, n47884, n47885, n47886,
         n47887, n47888, n47889, n47890, n47891, n47892, n47894, n47895,
         n47896, n47897, n47898, n47899, n47900, n47901, n47902, n47903,
         n47904, n47905, n47906, n47907, n47908, n47909, n47910, n47911,
         n47912, n47913, n47914, n47915, n47916, n47917, n47918, n47919,
         n47920, n47921, n47922, n47923, n47924, n47925, n47926, n47927,
         n47928, n47929, n47930, n47931, n47932, n47933, n47934, n47935,
         n47936, n47937, n47938, n47939, n47940, n47941, n47942, n47943,
         n47944, n47945, n47946, n47947, n47948, n47949, n47950, n47951,
         n47952, n47954, n47955, n47956, n47957, n47958, n47959, n47961,
         n47962, n47963, n47964, n47965, n47966, n47967, n47968, n47969,
         n47970, n47971, n47972, n47975, n47976, n47977, n47978, n47979,
         n47980, n47981, n47982, n47983, n47984, n47985, n47986, n47987,
         n47988, n47989, n47990, n47991, n47992, n47993, n47994, n47995,
         n47996, n47997, n47998, n47999, n48000, n48001, n48002, n48003,
         n48004, n48005, n48006, n48007, n48008, n48009, n48010, n48011,
         n48012, n48014, n48015, n48016, n48017, n48018, n48019, n48020,
         n48021, n48022, n48023, n48024, n48025, n48026, n48027, n48028,
         n48029, n48030, n48031, n48033, n48034, n48035, n48036, n48037,
         n48038, n48039, n48040, n48041, n48044, n48045, n48046, n48048,
         n48049, n48050, n48051, n48053, n48054, n48055, n48056, n48057,
         n48058, n48059, n48060, n48061, n48063, n48064, n48065, n48066,
         n48067, n48068, n48069, n48070, n48071, n48072, n48073, n48074,
         n48075, n48076, n48077, n48078, n48079, n48080, n48081, n48082,
         n48084, n48085, n48086, n48087, n48088, n48089, n48090, n48091,
         n48092, n48093, n48094, n48095, n48096, n48097, n48098, n48099,
         n48100, n48101, n48102, n48103, n48104, n48105, n48107, n48108,
         n48109, n48110, n48111, n48112, n48113, n48114, n48115, n48118,
         n48119, n48120, n48121, n48122, n48123, n48124, n48125, n48126,
         n48128, n48129, n48130, n48131, n48132, n48133, n48134, n48135,
         n48136, n48137, n48138, n48139, n48140, n48141, n48142, n48144,
         n48145, n48146, n48147, n48148, n48149, n48150, n48151, n48152,
         n48153, n48154, n48155, n48156, n48157, n48158, n48159, n48160,
         n48161, n48162, n48163, n48164, n48165, n48166, n48167, n48168,
         n48169, n48170, n48171, n48173, n48174, n48175, n48176, n48177,
         n48178, n48179, n48180, n48182, n48183, n48184, n48185, n48186,
         n48189, n48191, n48192, n48193, n48194, n48196, n48197, n48198,
         n48199, n48200, n48201, n48202, n48203, n48204, n48205, n48206,
         n48208, n48209, n48210, n48211, n48212, n48213, n48214, n48215,
         n48216, n48218, n48219, n48220, n48221, n48222, n48223, n48224,
         n48225, n48226, n48227, n48228, n48229, n48231, n48232, n48233,
         n48234, n48236, n48237, n48238, n48239, n48240, n48241, n48242,
         n48243, n48244, n48246, n48247, n48248, n48249, n48250, n48251,
         n48252, n48253, n48254, n48258, n48259, n48260, n48261, n48262,
         n48265, n48266, n48267, n48268, n48269, n48270, n48272, n48273,
         n48274, n48275, n48276, n48277, n48278, n48279, n48280, n48281,
         n48282, n48283, n48286, n48287, n48288, n48289, n48290, n48292,
         n48293, n48294, n48295, n48298, n48299, n48300, n48301, n48302,
         n48303, n48305, n48307, n48308, n48309, n48310, n48311, n48312,
         n48313, n48314, n48315, n48316, n48317, n48318, n48319, n48320,
         n48321, n48322, n48323, n48324, n48325, n48327, n48329, n48330,
         n48332, n48333, n48334, n48336, n48337, n48338, n48339, n48340,
         n48341, n48342, n48345, n48346, n48347, n48348, n48349, n48350,
         n48352, n48353, n48354, n48355, n48356, n48358, n48359, n48360,
         n48362, n48363, n48364, n48365, n48366, n48367, n48368, n48369,
         n48370, n48371, n48372, n48373, n48374, n48375, n48376, n48377,
         n48378, n48379, n48380, n48381, n48382, n48383, n48385, n48386,
         n48387, n48388, n48389, n48390, n48391, n48392, n48393, n48394,
         n48395, n48396, n48397, n48398, n48399, n48401, n48402, n48404,
         n48407, n48410, n48411, n48412, n48413, n48414, n48415, n48416,
         n48417, n48418, n48419, n48420, n48421, n48422, n48423, n48424,
         n48425, n48426, n48427, n48428, n48429, n48430, n48431, n48432,
         n48433, n48434, n48435, n48436, n48437, n48438, n48439, n48440,
         n48441, n48442, n48443, n48444, n48445, n48446, n48447, n48448,
         n48449, n48450, n48451, n48452, n48453, n48454, n48455, n48456,
         n48457, n48458, n48459, n48460, n48461, n48462, n48463, n48464,
         n48465, n48466, n48467, n48468, n48469, n48470, n48471, n48472,
         n48473, n48474, n48475, n48477, n48478, n48479, n48480, n48481,
         n48482, n48483, n48484, n48485, n48486, n48487, n48488, n48489,
         n48490, n48491, n48492, n48493, n48494, n48495, n48496, n48497,
         n48498, n48499, n48500, n48501, n48503, n48504, n48506, n48507,
         n48508, n48510, n48511, n48512, n48513, n48514, n48515, n48516,
         n48517, n48518, n48519, n48520, n48521, n48522, n48523, n48524,
         n48526, n48527, n48528, n48529, n48530, n48533, n48534, n48535,
         n48536, n48537, n48538, n48539, n48540, n48541, n48542, n48543,
         n48544, n48545, n48546, n48547, n48548, n48549, n48551, n48552,
         n48553, n48554, n48555, n48556, n48557, n48558, n48559, n48560,
         n48561, n48562, n48563, n48564, n48565, n48566, n48567, n48568,
         n48569, n48570, n48571, n48572, n48573, n48574, n48575, n48576,
         n48577, n48578, n48579, n48580, n48581, n48582, n48583, n48584,
         n48585, n48586, n48587, n48588, n48589, n48590, n48591, n48592,
         n48593, n48594, n48595, n48596, n48597, n48599, n48600, n48601,
         n48602, n48603, n48604, n48605, n48606, n48607, n48608, n48609,
         n48610, n48612, n48613, n48614, n48615, n48616, n48617, n48618,
         n48619, n48620, n48621, n48622, n48623, n48624, n48625, n48626,
         n48627, n48628, n48629, n48630, n48631, n48632, n48633, n48634,
         n48635, n48636, n48637, n48638, n48639, n48640, n48641, n48642,
         n48644, n48645, n48646, n48647, n48648, n48649, n48650, n48651,
         n48652, n48653, n48654, n48656, n48657, n48658, n48659, n48660,
         n48661, n48662, n48663, n48664, n48665, n48666, n48667, n48668,
         n48669, n48670, n48671, n48672, n48673, n48675, n48676, n48677,
         n48678, n48679, n48680, n48681, n48682, n48683, n48684, n48685,
         n48686, n48687, n48688, n48689, n48690, n48691, n48692, n48693,
         n48694, n48695, n48697, n48698, n48699, n48701, n48702, n48703,
         n48704, n48705, n48706, n48707, n48709, n48710, n48711, n48712,
         n48713, n48714, n48715, n48716, n48717, n48718, n48719, n48720,
         n48721, n48722, n48723, n48724, n48725, n48726, n48727, n48728,
         n48729, n48730, n48731, n48732, n48733, n48734, n48735, n48736,
         n48737, n48738, n48739, n48740, n48741, n48742, n48744, n48745,
         n48746, n48747, n48748, n48749, n48750, n48751, n48752, n48753,
         n48754, n48755, n48756, n48757, n48758, n48759, n48760, n48761,
         n48762, n48763, n48764, n48766, n48767, n48768, n48769, n48770,
         n48771, n48772, n48773, n48774, n48775, n48776, n48778, n48779,
         n48780, n48781, n48783, n48784, n48785, n48786, n48787, n48788,
         n48790, n48791, n48792, n48793, n48794, n48795, n48796, n48797,
         n48798, n48799, n48800, n48801, n48802, n48803, n48804, n48805,
         n48806, n48807, n48808, n48809, n48810, n48811, n48812, n48813,
         n48814, n48816, n48818, n48819, n48820, n48821, n48822, n48823,
         n48824, n48825, n48826, n48827, n48828, n48829, n48830, n48831,
         n48832, n48833, n48834, n48836, n48837, n48838, n48839, n48840,
         n48841, n48842, n48843, n48844, n48845, n48846, n48847, n48848,
         n48850, n48851, n48852, n48853, n48854, n48855, n48856, n48857,
         n48858, n48859, n48860, n48862, n48863, n48864, n48865, n48866,
         n48867, n48868, n48869, n48870, n48871, n48872, n48873, n48874,
         n48875, n48876, n48877, n48878, n48879, n48880, n48881, n48882,
         n48883, n48884, n48885, n48886, n48887, n48888, n48889, n48890,
         n48891, n48892, n48893, n48894, n48895, n48896, n48897, n48898,
         n48900, n48901, n48902, n48903, n48904, n48906, n48907, n48908,
         n48909, n48910, n48911, n48912, n48913, n48914, n48915, n48916,
         n48917, n48918, n48919, n48920, n48921, n48922, n48923, n48924,
         n48925, n48926, n48927, n48928, n48929, n48930, n48931, n48932,
         n48933, n48934, n48935, n48936, n48937, n48938, n48939, n48942,
         n48943, n48944, n48945, n48946, n48947, n48948, n48949, n48950,
         n48951, n48952, n48953, n48954, n48955, n48956, n48957, n48958,
         n48959, n48960, n48961, n48962, n48963, n48964, n48965, n48966,
         n48967, n48968, n48969, n48970, n48971, n48972, n48973, n48974,
         n48975, n48976, n48977, n48978, n48979, n48980, n48981, n48983,
         n48984, n48985, n48986, n48987, n48989, n48990, n48991, n48992,
         n48994, n48995, n48996, n48997, n48998, n48999, n49000, n49001,
         n49002, n49003, n49004, n49005, n49006, n49007, n49008, n49009,
         n49010, n49011, n49012, n49013, n49014, n49016, n49017, n49018,
         n49019, n49020, n49021, n49023, n49024, n49025, n49026, n49027,
         n49028, n49029, n49030, n49031, n49032, n49033, n49034, n49035,
         n49036, n49037, n49038, n49039, n49041, n49042, n49043, n49044,
         n49045, n49046, n49047, n49048, n49049, n49050, n49051, n49052,
         n49053, n49054, n49055, n49056, n49057, n49058, n49059, n49060,
         n49061, n49062, n49063, n49064, n49065, n49066, n49067, n49068,
         n49069, n49071, n49072, n49073, n49074, n49075, n49076, n49077,
         n49078, n49079, n49080, n49081, n49082, n49083, n49084, n49085,
         n49086, n49087, n49088, n49089, n49090, n49091, n49092, n49093,
         n49094, n49095, n49096, n49097, n49098, n49099, n49100, n49101,
         n49102, n49103, n49104, n49105, n49106, n49107, n49108, n49109,
         n49110, n49111, n49112, n49113, n49114, n49115, n49116, n49117,
         n49118, n49119, n49120, n49121, n49122, n49123, n49124, n49125,
         n49126, n49127, n49128, n49129, n49130, n49131, n49132, n49133,
         n49134, n49135, n49136, n49137, n49138, n49139, n49140, n49141,
         n49142, n49144, n49145, n49146, n49147, n49149, n49150, n49151,
         n49152, n49153, n49154, n49155, n49156, n49157, n49158, n49159,
         n49160, n49161, n49162, n49163, n49164, n49165, n49166, n49167,
         n49168, n49169, n49170, n49171, n49172, n49173, n49174, n49175,
         n49176, n49177, n49178, n49179, n49180, n49181, n49182, n49183,
         n49184, n49185, n49186, n49187, n49188, n49189, n49190, n49191,
         n49192, n49193, n49194, n49195, n49196, n49197, n49198, n49199,
         n49200, n49201, n49202, n49203, n49205, n49206, n49207, n49209,
         n49210, n49211, n49213, n49214, n49215, n49216, n49217, n49218,
         n49219, n49220, n49221, n49222, n49223, n49224, n49225, n49226,
         n49227, n49228, n49229, n49231, n49232, n49233, n49234, n49235,
         n49236, n49237, n49238, n49239, n49240, n49241, n49243, n49244,
         n49245, n49247, n49248, n49249, n49250, n49251, n49252, n49253,
         n49254, n49255, n49256, n49257, n49258, n49259, n49260, n49261,
         n49262, n49263, n49264, n49265, n49266, n49267, n49268, n49269,
         n49270, n49271, n49272, n49273, n49274, n49275, n49276, n49277,
         n49278, n49280, n49281, n49282, n49283, n49284, n49286, n49287,
         n49288, n49289, n49290, n49291, n49292, n49293, n49294, n49295,
         n49296, n49298, n49299, n49300, n49301, n49302, n49303, n49304,
         n49305, n49306, n49307, n49308, n49309, n49310, n49311, n49312,
         n49313, n49314, n49315, n49316, n49317, n49318, n49319, n49320,
         n49321, n49322, n49323, n49324, n49325, n49326, n49327, n49328,
         n49329, n49330, n49331, n49332, n49333, n49334, n49335, n49336,
         n49337, n49338, n49339, n49340, n49341, n49342, n49343, n49344,
         n49345, n49346, n49347, n49348, n49349, n49350, n49351, n49352,
         n49353, n49354, n49355, n49356, n49357, n49358, n49359, n49360,
         n49361, n49362, n49363, n49364, n49365, n49366, n49367, n49368,
         n49369, n49370, n49371, n49372, n49373, n49374, n49375, n49376,
         n49377, n49378, n49379, n49380, n49382, n49383, n49384, n49385,
         n49386, n49387, n49388, n49389, n49390, n49391, n49393, n49394,
         n49395, n49396, n49397, n49398, n49399, n49400, n49401, n49402,
         n49403, n49404, n49405, n49406, n49407, n49408, n49409, n49410,
         n49411, n49412, n49413, n49414, n49415, n49416, n49419, n49420,
         n49421, n49422, n49425, n49426, n49427, n49428, n49429, n49430,
         n49431, n49432, n49433, n49434, n49435, n49436, n49437, n49438,
         n49439, n49440, n49441, n49442, n49443, n49444, n49445, n49446,
         n49447, n49448, n49449, n49450, n49451, n49452, n49453, n49454,
         n49455, n49456, n49458, n49459, n49460, n49461, n49462, n49463,
         n49464, n49465, n49466, n49467, n49469, n49470, n49471, n49472,
         n49473, n49475, n49476, n49477, n49478, n49482, n49483, n49484,
         n49485, n49486, n49487, n49488, n49489, n49490, n49491, n49492,
         n49493, n49494, n49495, n49496, n49498, n49499, n49500, n49501,
         n49502, n49503, n49504, n49505, n49506, n49507, n49508, n49510,
         n49511, n49512, n49513, n49514, n49515, n49516, n49520, n49521,
         n49522, n49523, n49524, n49525, n49526, n49527, n49528, n49529,
         n49530, n49531, n49532, n49533, n49534, n49535, n49536, n49538,
         n49539, n49540, n49541, n49542, n49543, n49544, n49545, n49546,
         n49547, n49548, n49549, n49550, n49551, n49552, n49553, n49554,
         n49555, n49556, n49557, n49558, n49559, n49560, n49561, n49562,
         n49563, n49564, n49565, n49566, n49567, n49568, n49569, n49570,
         n49571, n49572, n49573, n49574, n49575, n49576, n49578, n49579,
         n49580, n49581, n49582, n49583, n49584, n49585, n49586, n49587,
         n49588, n49589, n49590, n49591, n49593, n49594, n49595, n49597,
         n49598, n49599, n49600, n49601, n49602, n49603, n49604, n49605,
         n49606, n49607, n49608, n49609, n49610, n49612, n49613, n49614,
         n49617, n49618, n49619, n49620, n49621, n49622, n49623, n49624,
         n49625, n49626, n49627, n49628, n49629, n49630, n49631, n49632,
         n49633, n49634, n49635, n49637, n49638, n49639, n49640, n49641,
         n49642, n49643, n49644, n49645, n49646, n49647, n49648, n49649,
         n49650, n49651, n49652, n49653, n49654, n49655, n49656, n49657,
         n49658, n49659, n49661, n49662, n49664, n49665, n49666, n49667,
         n49668, n49669, n49670, n49671, n49673, n49674, n49675, n49676,
         n49677, n49678, n49679, n49681, n49682, n49684, n49685, n49686,
         n49687, n49688, n49689, n49691, n49692, n49693, n49694, n49695,
         n49696, n49697, n49698, n49699, n49700, n49701, n49702, n49703,
         n49704, n49705, n49706, n49707, n49708, n49709, n49710, n49711,
         n49712, n49713, n49714, n49715, n49716, n49717, n49718, n49719,
         n49720, n49721, n49722, n49723, n49724, n49725, n49726, n49727,
         n49728, n49729, n49730, n49731, n49732, n49733, n49734, n49735,
         n49736, n49737, n49738, n49739, n49740, n49741, n49742, n49743,
         n49744, n49745, n49748, n49749, n49750, n49751, n49752, n49753,
         n49754, n49755, n49756, n49757, n49758, n49759, n49760, n49761,
         n49762, n49763, n49764, n49765, n49766, n49767, n49768, n49769,
         n49770, n49771, n49772, n49774, n49775, n49776, n49777, n49778,
         n49779, n49780, n49781, n49782, n49783, n49784, n49785, n49787,
         n49788, n49789, n49790, n49791, n49792, n49793, n49794, n49795,
         n49796, n49797, n49798, n49799, n49802, n49803, n49804, n49805,
         n49806, n49807, n49808, n49809, n49810, n49811, n49813, n49814,
         n49815, n49816, n49817, n49818, n49819, n49820, n49821, n49822,
         n49823, n49824, n49825, n49827, n49828, n49829, n49830, n49831,
         n49832, n49833, n49834, n49835, n49836, n49838, n49839, n49840,
         n49841, n49842, n49843, n49844, n49845, n49846, n49847, n49848,
         n49849, n49850, n49851, n49852, n49853, n49854, n49855, n49856,
         n49857, n49858, n49859, n49860, n49861, n49862, n49863, n49864,
         n49865, n49866, n49867, n49868, n49869, n49870, n49871, n49873,
         n49874, n49875, n49876, n49877, n49878, n49879, n49881, n49882,
         n49883, n49884, n49885, n49886, n49887, n49888, n49889, n49890,
         n49891, n49893, n49894, n49895, n49897, n49898, n49899, n49900,
         n49901, n49902, n49903, n49904, n49905, n49906, n49907, n49908,
         n49909, n49910, n49911, n49912, n49913, n49914, n49915, n49916,
         n49917, n49918, n49919, n49920, n49921, n49922, n49923, n49924,
         n49926, n49927, n49928, n49929, n49930, n49931, n49932, n49933,
         n49934, n49935, n49936, n49937, n49938, n49939, n49940, n49941,
         n49942, n49943, n49944, n49945, n49946, n49947, n49948, n49949,
         n49950, n49951, n49952, n49953, n49954, n49955, n49956, n49957,
         n49958, n49959, n49960, n49961, n49962, n49963, n49964, n49965,
         n49966, n49967, n49968, n49969, n49970, n49971, n49972, n49973,
         n49976, n49977, n49978, n49979, n49980, n49981, n49982, n49983,
         n49985, n49986, n49989, n49990, n49991, n49993, n49994, n49996,
         n49997, n49998, n49999, n50000, n50001, n50002, n50004, n50005,
         n50006, n50007, n50009, n50010, n50011, n50012, n50013, n50014,
         n50015, n50016, n50017, n50018, n50019, n50020, n50021, n50022,
         n50023, n50025, n50026, n50027, n50028, n50030, n50031, n50032,
         n50033, n50034, n50035, n50036, n50037, n50038, n50039, n50040,
         n50041, n50042, n50043, n50044, n50045, n50046, n50047, n50048,
         n50049, n50050, n50051, n50052, n50053, n50054, n50055, n50056,
         n50057, n50058, n50059, n50060, n50062, n50063, n50064, n50065,
         n50066, n50067, n50068, n50069, n50070, n50071, n50072, n50073,
         n50074, n50075, n50076, n50077, n50078, n50079, n50080, n50081,
         n50082, n50083, n50084, n50086, n50087, n50088, n50090, n50091,
         n50092, n50093, n50094, n50095, n50096, n50097, n50098, n50099,
         n50100, n50101, n50102, n50103, n50104, n50105, n50107, n50108,
         n50109, n50110, n50111, n50112, n50113, n50114, n50115, n50117,
         n50119, n50120, n50121, n50122, n50123, n50124, n50125, n50126,
         n50127, n50128, n50129, n50130, n50131, n50132, n50133, n50134,
         n50136, n50137, n50138, n50139, n50140, n50141, n50142, n50143,
         n50144, n50145, n50146, n50147, n50148, n50149, n50150, n50151,
         n50152, n50153, n50154, n50155, n50157, n50159, n50160, n50161,
         n50162, n50163, n50164, n50165, n50166, n50167, n50168, n50169,
         n50170, n50171, n50172, n50173, n50174, n50175, n50176, n50177,
         n50178, n50179, n50180, n50181, n50182, n50183, n50184, n50185,
         n50186, n50187, n50188, n50189, n50190, n50191, n50192, n50193,
         n50194, n50195, n50196, n50197, n50198, n50199, n50200, n50201,
         n50202, n50203, n50204, n50205, n50206, n50207, n50208, n50209,
         n50210, n50211, n50212, n50213, n50214, n50215, n50216, n50218,
         n50219, n50220, n50221, n50222, n50223, n50225, n50227, n50228,
         n50229, n50230, n50231, n50232, n50233, n50234, n50235, n50236,
         n50237, n50238, n50239, n50240, n50241, n50242, n50243, n50244,
         n50245, n50246, n50247, n50248, n50249, n50250, n50251, n50252,
         n50253, n50254, n50255, n50257, n50258, n50259, n50260, n50261,
         n50262, n50263, n50264, n50265, n50266, n50267, n50268, n50269,
         n50270, n50271, n50272, n50273, n50274, n50275, n50276, n50277,
         n50278, n50280, n50281, n50282, n50283, n50284, n50285, n50286,
         n50287, n50288, n50289, n50290, n50291, n50292, n50293, n50294,
         n50295, n50296, n50297, n50298, n50300, n50301, n50302, n50303,
         n50304, n50305, n50306, n50307, n50308, n50309, n50310, n50312,
         n50313, n50314, n50315, n50316, n50317, n50318, n50319, n50320,
         n50321, n50322, n50323, n50324, n50325, n50326, n50328, n50329,
         n50330, n50331, n50332, n50333, n50334, n50336, n50337, n50338,
         n50339, n50340, n50341, n50342, n50343, n50345, n50346, n50348,
         n50349, n50350, n50351, n50352, n50353, n50354, n50355, n50357,
         n50358, n50359, n50360, n50361, n50362, n50363, n50364, n50365,
         n50366, n50367, n50369, n50370, n50371, n50372, n50373, n50374,
         n50375, n50376, n50378, n50379, n50380, n50381, n50382, n50383,
         n50384, n50385, n50386, n50387, n50388, n50389, n50390, n50391,
         n50392, n50393, n50394, n50395, n50396, n50397, n50398, n50399,
         n50400, n50401, n50402, n50403, n50404, n50405, n50406, n50407,
         n50408, n50409, n50410, n50411, n50412, n50413, n50414, n50415,
         n50416, n50417, n50418, n50419, n50420, n50421, n50422, n50423,
         n50424, n50425, n50426, n50427, n50428, n50429, n50430, n50431,
         n50433, n50434, n50435, n50436, n50437, n50438, n50439, n50440,
         n50441, n50442, n50443, n50444, n50446, n50447, n50448, n50449,
         n50450, n50451, n50452, n50453, n50454, n50455, n50456, n50457,
         n50458, n50459, n50460, n50461, n50462, n50463, n50464, n50465,
         n50466, n50467, n50468, n50469, n50470, n50471, n50472, n50473,
         n50474, n50475, n50476, n50477, n50478, n50480, n50482, n50484,
         n50485, n50486, n50487, n50488, n50489, n50490, n50491, n50492,
         n50493, n50494, n50495, n50496, n50497, n50498, n50499, n50500,
         n50501, n50502, n50503, n50504, n50505, n50506, n50507, n50508,
         n50509, n50510, n50511, n50512, n50513, n50514, n50515, n50516,
         n50517, n50518, n50519, n50520, n50521, n50522, n50523, n50524,
         n50525, n50526, n50527, n50528, n50529, n50530, n50531, n50532,
         n50533, n50534, n50535, n50536, n50537, n50538, n50539, n50540,
         n50541, n50543, n50544, n50545, n50546, n50547, n50548, n50549,
         n50550, n50551, n50552, n50553, n50554, n50555, n50556, n50557,
         n50558, n50559, n50560, n50561, n50562, n50563, n50564, n50565,
         n50566, n50567, n50568, n50569, n50570, n50571, n50572, n50573,
         n50574, n50575, n50576, n50577, n50578, n50579, n50580, n50581,
         n50582, n50583, n50584, n50585, n50586, n50587, n50588, n50589,
         n50590, n50591, n50592, n50593, n50594, n50595, n50596, n50597,
         n50598, n50599, n50600, n50601, n50602, n50603, n50604, n50606,
         n50607, n50608, n50609, n50610, n50611, n50612, n50613, n50614,
         n50615, n50616, n50617, n50618, n50619, n50620, n50621, n50622,
         n50623, n50624, n50625, n50626, n50627, n50628, n50629, n50630,
         n50631, n50632, n50633, n50634, n50635, n50636, n50637, n50638,
         n50639, n50640, n50641, n50642, n50643, n50644, n50646, n50648,
         n50649, n50650, n50651, n50652, n50653, n50654, n50655, n50656,
         n50657, n50658, n50660, n50661, n50662, n50663, n50664, n50665,
         n50666, n50667, n50668, n50669, n50670, n50671, n50672, n50673,
         n50674, n50675, n50676, n50678, n50679, n50680, n50681, n50682,
         n50683, n50684, n50685, n50686, n50687, n50688, n50689, n50690,
         n50691, n50692, n50693, n50694, n50695, n50696, n50697, n50698,
         n50699, n50700, n50701, n50702, n50703, n50704, n50705, n50706,
         n50707, n50708, n50709, n50710, n50711, n50712, n50713, n50714,
         n50715, n50716, n50717, n50718, n50719, n50720, n50721, n50722,
         n50723, n50724, n50725, n50726, n50727, n50728, n50729, n50730,
         n50731, n50732, n50733, n50734, n50735, n50736, n50737, n50738,
         n50739, n50740, n50741, n50742, n50743, n50745, n50746, n50747,
         n50748, n50749, n50750, n50751, n50752, n50754, n50755, n50756,
         n50757, n50758, n50759, n50760, n50761, n50762, n50763, n50764,
         n50765, n50766, n50767, n50768, n50769, n50770, n50771, n50772,
         n50773, n50775, n50776, n50777, n50778, n50779, n50780, n50781,
         n50782, n50783, n50784, n50785, n50786, n50787, n50788, n50789,
         n50790, n50791, n50792, n50793, n50794, n50795, n50796, n50797,
         n50798, n50799, n50800, n50801, n50802, n50803, n50804, n50806,
         n50807, n50808, n50809, n50810, n50811, n50814, n50816, n50817,
         n50818, n50820, n50821, n50822, n50823, n50824, n50825, n50826,
         n50828, n50829, n50830, n50831, n50832, n50833, n50834, n50835,
         n50836, n50837, n50838, n50839, n50840, n50841, n50842, n50843,
         n50844, n50845, n50846, n50847, n50848, n50849, n50850, n50851,
         n50852, n50853, n50855, n50856, n50857, n50858, n50859, n50860,
         n50861, n50862, n50863, n50864, n50865, n50866, n50867, n50868,
         n50869, n50870, n50871, n50872, n50873, n50874, n50875, n50876,
         n50878, n50879, n50880, n50882, n50883, n50884, n50885, n50886,
         n50887, n50888, n50889, n50890, n50892, n50893, n50894, n50895,
         n50896, n50898, n50899, n50900, n50901, n50902, n50903, n50904,
         n50905, n50906, n50907, n50908, n50909, n50910, n50911, n50912,
         n50913, n50914, n50915, n50916, n50917, n50918, n50919, n50920,
         n50921, n50923, n50924, n50925, n50926, n50927, n50929, n50930,
         n50931, n50932, n50933, n50934, n50935, n50936, n50937, n50938,
         n50939, n50940, n50941, n50942, n50943, n50944, n50945, n50946,
         n50947, n50948, n50949, n50951, n50952, n50953, n50954, n50955,
         n50956, n50957, n50958, n50959, n50960, n50961, n50962, n50963,
         n50964, n50965, n50966, n50967, n50968, n50969, n50970, n50971,
         n50972, n50973, n50974, n50975, n50976, n50977, n50978, n50979,
         n50980, n50981, n50982, n50983, n50984, n50985, n50986, n50987,
         n50988, n50989, n50990, n50991, n50992, n50993, n50994, n50995,
         n50997, n50998, n50999, n51000, n51001, n51002, n51003, n51004,
         n51005, n51006, n51007, n51008, n51009, n51010, n51011, n51012,
         n51013, n51015, n51016, n51017, n51018, n51019, n51020, n51021,
         n51022, n51023, n51024, n51025, n51026, n51027, n51028, n51029,
         n51030, n51031, n51032, n51033, n51034, n51035, n51036, n51037,
         n51038, n51039, n51040, n51041, n51042, n51043, n51044, n51045,
         n51046, n51047, n51048, n51049, n51050, n51051, n51052, n51053,
         n51054, n51056, n51057, n51058, n51059, n51060, n51061, n51062,
         n51063, n51064, n51065, n51066, n51067, n51068, n51069, n51070,
         n51071, n51072, n51073, n51074, n51075, n51076, n51077, n51078,
         n51080, n51081, n51082, n51083, n51084, n51085, n51086, n51087,
         n51088, n51089, n51090, n51091, n51092, n51093, n51094, n51095,
         n51096, n51097, n51099, n51100, n51101, n51102, n51103, n51104,
         n51105, n51106, n51107, n51110, n51112, n51113, n51114, n51115,
         n51116, n51119, n51120, n51121, n51122, n51123, n51124, n51125,
         n51126, n51127, n51128, n51129, n51130, n51131, n51132, n51133,
         n51134, n51135, n51136, n51137, n51138, n51139, n51140, n51141,
         n51142, n51143, n51144, n51145, n51146, n51147, n51148, n51149,
         n51150, n51151, n51152, n51153, n51154, n51155, n51156, n51158,
         n51159, n51160, n51161, n51162, n51163, n51164, n51165, n51166,
         n51167, n51168, n51169, n51170, n51171, n51172, n51173, n51174,
         n51175, n51176, n51177, n51178, n51179, n51180, n51181, n51185,
         n51186, n51187, n51188, n51189, n51190, n51191, n51192, n51193,
         n51194, n51195, n51196, n51197, n51198, n51199, n51200, n51201,
         n51202, n51203, n51204, n51205, n51206, n51207, n51208, n51209,
         n51210, n51211, n51213, n51214, n51215, n51216, n51217, n51218,
         n51219, n51220, n51221, n51222, n51223, n51224, n51225, n51226,
         n51227, n51228, n51229, n51230, n51231, n51232, n51233, n51234,
         n51235, n51236, n51237, n51238, n51239, n51240, n51241, n51242,
         n51243, n51244, n51245, n51246, n51247, n51248, n51249, n51250,
         n51251, n51252, n51253, n51254, n51256, n51257, n51258, n51259,
         n51260, n51261, n51262, n51263, n51264, n51265, n51266, n51267,
         n51268, n51269, n51270, n51271, n51273, n51274, n51275, n51276,
         n51277, n51278, n51279, n51280, n51281, n51282, n51283, n51284,
         n51285, n51286, n51287, n51288, n51289, n51290, n51291, n51292,
         n51293, n51294, n51295, n51296, n51297, n51298, n51299, n51300,
         n51301, n51302, n51303, n51304, n51305, n51306, n51307, n51308,
         n51309, n51310, n51311, n51312, n51313, n51314, n51315, n51316,
         n51317, n51318, n51319, n51320, n51321, n51322, n51323, n51324,
         n51325, n51326, n51327, n51328, n51329, n51330, n51331, n51332,
         n51333, n51334, n51335, n51337, n51338, n51339, n51340, n51341,
         n51342, n51343, n51344, n51345, n51346, n51347, n51348, n51349,
         n51350, n51351, n51352, n51353, n51354, n51355, n51356, n51357,
         n51358, n51360, n51361, n51362, n51363, n51364, n51365, n51366,
         n51367, n51368, n51369, n51370, n51371, n51372, n51373, n51374,
         n51375, n51376, n51377, n51379, n51380, n51381, n51382, n51383,
         n51384, n51385, n51386, n51387, n51388, n51389, n51390, n51391,
         n51392, n51393, n51394, n51395, n51396, n51397, n51398, n51399,
         n51400, n51402, n51403, n51404, n51405, n51406, n51407, n51408,
         n51409, n51410, n51411, n51412, n51413, n51414, n51415, n51416,
         n51417, n51418, n51419, n51420, n51421, n51422, n51423, n51424,
         n51425, n51426, n51428, n51429, n51430, n51431, n51432, n51433,
         n51434, n51435, n51437, n51438, n51439, n51440, n51441, n51442,
         n51443, n51444, n51445, n51446, n51447, n51448, n51449, n51450,
         n51451, n51452, n51453, n51454, n51455, n51456, n51457, n51458,
         n51459, n51460, n51461, n51462, n51463, n51465, n51466, n51467,
         n51468, n51469, n51470, n51472, n51473, n51474, n51475, n51476,
         n51477, n51478, n51479, n51480, n51481, n51482, n51483, n51484,
         n51485, n51486, n51487, n51488, n51489, n51490, n51491, n51492,
         n51493, n51494, n51495, n51496, n51497, n51498, n51499, n51500,
         n51501, n51502, n51503, n51504, n51505, n51506, n51507, n51508,
         n51509, n51510, n51511, n51512, n51513, n51514, n51515, n51516,
         n51517, n51518, n51519, n51520, n51521, n51522, n51523, n51524,
         n51525, n51526, n51527, n51528, n51529, n51530, n51531, n51532,
         n51533, n51534, n51535, n51536, n51537, n51538, n51539, n51540,
         n51541, n51542, n51543, n51544, n51545, n51546, n51547, n51548,
         n51549, n51550, n51551, n51552, n51553, n51554, n51555, n51556,
         n51557, n51558, n51559, n51560, n51561, n51562, n51563, n51565,
         n51567, n51568, n51569, n51570, n51572, n51573, n51574, n51575,
         n51576, n51577, n51578, n51579, n51580, n51581, n51582, n51583,
         n51584, n51585, n51586, n51587, n51588, n51589, n51590, n51591,
         n51592, n51593, n51594, n51595, n51596, n51597, n51598, n51599,
         n51600, n51601, n51602, n51604, n51605, n51606, n51607, n51608,
         n51609, n51610, n51611, n51612, n51613, n51614, n51615, n51616,
         n51617, n51618, n51619, n51620, n51621, n51622, n51623, n51624,
         n51625, n51626, n51627, n51628, n51629, n51630, n51631, n51632,
         n51633, n51635, n51636, n51637, n51638, n51639, n51640, n51641,
         n51642, n51643, n51644, n51645, n51646, n51647, n51648, n51649,
         n51650, n51651, n51652, n51653, n51654, n51655, n51656, n51657,
         n51658, n51659, n51660, n51661, n51662, n51663, n51664, n51665,
         n51666, n51667, n51668, n51669, n51670, n51671, n51672, n51673,
         n51674, n51675, n51676, n51677, n51678, n51679, n51680, n51681,
         n51682, n51683, n51684, n51685, n51686, n51687, n51688, n51689,
         n51690, n51691, n51692, n51693, n51694, n51695, n51696, n51697,
         n51699, n51700, n51701, n51702, n51703, n51704, n51705, n51706,
         n51707, n51709, n51710, n51711, n51712, n51713, n51714, n51715,
         n51716, n51717, n51718, n51719, n51720, n51721, n51722, n51723,
         n51724, n51725, n51726, n51727, n51729, n51730, n51731, n51732,
         n51733, n51734, n51735, n51736, n51737, n51738, n51740, n51741,
         n51742, n51743, n51744, n51745, n51746, n51748, n51749, n51750,
         n51751, n51752, n51753, n51754, n51755, n51756, n51757, n51758,
         n51759, n51760, n51761, n51762, n51763, n51764, n51765, n51766,
         n51767, n51768, n51769, n51770, n51771, n51772, n51775, n51776,
         n51777, n51779, n51780, n51781, n51782, n51783, n51786, n51788,
         n51789, n51790, n51792, n51793, n51794, n51795, n51796, n51797,
         n51798, n51799, n51800, n51801, n51802, n51803, n51804, n51805,
         n51806, n51807, n51808, n51809, n51810, n51812, n51813, n51814,
         n51815, n51816, n51817, n51818, n51819, n51820, n51821, n51823,
         n51824, n51825, n51826, n51827, n51828, n51829, n51830, n51831,
         n51832, n51833, n51834, n51835, n51837, n51838, n51839, n51840,
         n51841, n51842, n51843, n51844, n51845, n51846, n51847, n51848,
         n51849, n51850, n51851, n51852, n51853, n51855, n51858, n51859,
         n51860, n51861, n51862, n51863, n51864, n51865, n51866, n51867,
         n51868, n51869, n51870, n51871, n51872, n51873, n51874, n51875,
         n51876, n51877, n51878, n51879, n51880, n51881, n51882, n51884,
         n51886, n51887, n51888, n51889, n51890, n51891, n51892, n51893,
         n51894, n51895, n51897, n51898, n51899, n51900, n51901, n51902,
         n51903, n51904, n51905, n51906, n51907, n51908, n51909, n51910,
         n51911, n51912, n51913, n51914, n51915, n51916, n51917, n51918,
         n51919, n51920, n51921, n51922, n51924, n51925, n51926, n51927,
         n51928, n51929, n51930, n51931, n51932, n51933, n51934, n51935,
         n51936, n51937, n51939, n51940, n51941, n51942, n51943, n51944,
         n51945, n51946, n51947, n51948, n51949, n51950, n51951, n51952,
         n51953, n51954, n51955, n51956, n51957, n51958, n51959, n51960,
         n51961, n51962, n51963, n51964, n51965, n51966, n51967, n51968,
         n51969, n51970, n51971, n51972, n51973, n51974, n51975, n51976,
         n51977, n51978, n51979, n51980, n51981, n51982, n51983, n51984,
         n51985, n51986, n51987, n51988, n51989, n51990, n51991, n51992,
         n51993, n51994, n51995, n51996, n51997, n51998, n51999, n52000,
         n52001, n52002, n52003, n52004, n52005, n52006, n52007, n52008,
         n52009, n52010, n52011, n52012, n52013, n52014, n52015, n52016,
         n52017, n52018, n52019, n52020, n52021, n52022, n52023, n52024,
         n52025, n52026, n52028, n52029, n52030, n52031, n52032, n52033,
         n52034, n52035, n52036, n52037, n52038, n52039, n52040, n52041,
         n52042, n52043, n52044, n52045, n52046, n52047, n52048, n52049,
         n52050, n52051, n52052, n52053, n52054, n52055, n52058, n52059,
         n52060, n52061, n52062, n52063, n52064, n52065, n52066, n52067,
         n52068, n52069, n52070, n52071, n52072, n52073, n52075, n52076,
         n52077, n52078, n52079, n52080, n52081, n52082, n52083, n52084,
         n52085, n52086, n52087, n52088, n52089, n52090, n52091, n52092,
         n52093, n52094, n52095, n52096, n52097, n52098, n52099, n52100,
         n52101, n52102, n52103, n52104, n52105, n52106, n52107, n52108,
         n52109, n52110, n52111, n52112, n52113, n52114, n52115, n52116,
         n52117, n52118, n52119, n52120, n52121, n52122, n52123, n52124,
         n52125, n52126, n52127, n52129, n52130, n52131, n52133, n52134,
         n52135, n52136, n52137, n52138, n52139, n52140, n52141, n52142,
         n52143, n52144, n52145, n52146, n52147, n52148, n52149, n52150,
         n52151, n52152, n52153, n52154, n52155, n52156, n52157, n52159,
         n52160, n52161, n52162, n52164, n52165, n52166, n52167, n52168,
         n52169, n52170, n52171, n52172, n52173, n52174, n52175, n52176,
         n52177, n52178, n52179, n52180, n52181, n52182, n52183, n52184,
         n52185, n52186, n52187, n52188, n52189, n52190, n52192, n52193,
         n52195, n52196, n52197, n52198, n52199, n52200, n52201, n52202,
         n52203, n52204, n52205, n52206, n52207, n52208, n52209, n52210,
         n52211, n52212, n52213, n52216, n52217, n52218, n52219, n52220,
         n52222, n52223, n52224, n52225, n52226, n52227, n52228, n52229,
         n52230, n52231, n52232, n52233, n52234, n52235, n52236, n52237,
         n52238, n52239, n52240, n52241, n52245, n52246, n52247, n52248,
         n52249, n52250, n52251, n52252, n52253, n52254, n52255, n52256,
         n52257, n52258, n52259, n52261, n52262, n52263, n52264, n52265,
         n52266, n52267, n52268, n52269, n52270, n52271, n52272, n52273,
         n52275, n52276, n52277, n52278, n52279, n52280, n52281, n52282,
         n52283, n52284, n52285, n52287, n52288, n52289, n52291, n52292,
         n52293, n52294, n52295, n52296, n52297, n52298, n52299, n52300,
         n52301, n52302, n52303, n52304, n52305, n52307, n52309, n52310,
         n52311, n52312, n52313, n52314, n52315, n52317, n52319, n52320,
         n52321, n52322, n52323, n52325, n52326, n52327, n52328, n52329,
         n52330, n52331, n52332, n52333, n52334, n52335, n52336, n52337,
         n52338, n52339, n52340, n52341, n52342, n52343, n52344, n52345,
         n52346, n52348, n52349, n52350, n52351, n52352, n52353, n52354,
         n52355, n52356, n52357, n52358, n52360, n52361, n52362, n52363,
         n52364, n52365, n52366, n52367, n52368, n52369, n52370, n52371,
         n52372, n52373, n52374, n52375, n52376, n52377, n52378, n52379,
         n52380, n52381, n52382, n52383, n52384, n52385, n52386, n52387,
         n52388, n52389, n52390, n52393, n52394, n52396, n52397, n52398,
         n52399, n52400, n52401, n52402, n52403, n52404, n52405, n52406,
         n52407, n52408, n52409, n52410, n52411, n52412, n52413, n52414,
         n52415, n52416, n52417, n52418, n52419, n52420, n52421, n52422,
         n52423, n52424, n52425, n52426, n52427, n52428, n52429, n52430,
         n52431, n52432, n52433, n52434, n52435, n52436, n52437, n52438,
         n52439, n52440, n52441, n52442, n52443, n52444, n52445, n52446,
         n52447, n52448, n52449, n52450, n52451, n52452, n52453, n52454,
         n52455, n52456, n52457, n52458, n52459, n52460, n52461, n52462,
         n52463, n52464, n52465, n52466, n52467, n52468, n52469, n52470,
         n52471, n52472, n52473, n52475, n52476, n52477, n52478, n52479,
         n52480, n52482, n52483, n52484, n52485, n52486, n52487, n52488,
         n52489, n52490, n52491, n52492, n52493, n52494, n52495, n52496,
         n52497, n52498, n52499, n52500, n52501, n52502, n52503, n52504,
         n52505, n52506, n52507, n52508, n52509, n52510, n52511, n52512,
         n52513, n52514, n52515, n52516, n52517, n52518, n52519, n52520,
         n52521, n52522, n52523, n52524, n52525, n52526, n52527, n52529,
         n52530, n52531, n52532, n52533, n52534, n52535, n52536, n52537,
         n52538, n52539, n52540, n52541, n52543, n52544, n52545, n52546,
         n52547, n52548, n52549, n52550, n52551, n52552, n52553, n52554,
         n52555, n52556, n52557, n52558, n52559, n52560, n52561, n52562,
         n52563, n52564, n52565, n52566, n52567, n52568, n52569, n52570,
         n52572, n52573, n52574, n52575, n52576, n52577, n52578, n52579,
         n52580, n52581, n52582, n52583, n52584, n52585, n52586, n52587,
         n52588, n52589, n52590, n52591, n52592, n52593, n52594, n52595,
         n52596, n52597, n52598, n52599, n52600, n52601, n52602, n52603,
         n52604, n52605, n52606, n52607, n52608, n52609, n52610, n52611,
         n52612, n52613, n52614, n52615, n52616, n52617, n52618, n52619,
         n52620, n52621, n52622, n52623, n52624, n52625, n52626, n52627,
         n52628, n52629, n52630, n52631, n52632, n52633, n52634, n52635,
         n52636, n52637, n52638, n52639, n52640, n52641, n52642, n52643,
         n52645, n52646, n52647, n52648, n52649, n52650, n52651, n52652,
         n52653, n52654, n52655, n52656, n52657, n52658, n52659, n52661,
         n52662, n52665, n52667, n52668, n52669, n52670, n52671, n52672,
         n52673, n52674, n52675, n52676, n52677, n52678, n52679, n52680,
         n52681, n52682, n52683, n52685, n52686, n52687, n52688, n52689,
         n52690, n52691, n52692, n52694, n52695, n52696, n52697, n52698,
         n52699, n52700, n52701, n52702, n52703, n52704, n52705, n52706,
         n52707, n52708, n52709, n52710, n52712, n52713, n52714, n52715,
         n52716, n52717, n52719, n52720, n52721, n52723, n52725, n52726,
         n52727, n52728, n52729, n52730, n52731, n52732, n52733, n52734,
         n52735, n52737, n52738, n52739, n52743, n52744, n52745, n52746,
         n52747, n52748, n52749, n52750, n52751, n52752, n52753, n52754,
         n52755, n52756, n52757, n52758, n52759, n52760, n52761, n52762,
         n52763, n52765, n52766, n52767, n52768, n52769, n52770, n52771,
         n52772, n52774, n52775, n52776, n52778, n52779, n52780, n52781,
         n52782, n52783, n52784, n52786, n52787, n52788, n52789, n52790,
         n52792, n52794, n52795, n52796, n52797, n52798, n52799, n52800,
         n52801, n52802, n52803, n52804, n52805, n52806, n52807, n52808,
         n52809, n52810, n52811, n52812, n52813, n52814, n52815, n52816,
         n52817, n52818, n52819, n52820, n52821, n52822, n52823, n52824,
         n52825, n52826, n52827, n52828, n52829, n52830, n52831, n52832,
         n52833, n52834, n52835, n52836, n52837, n52838, n52839, n52840,
         n52841, n52842, n52843, n52844, n52845, n52846, n52847, n52848,
         n52849, n52850, n52851, n52852, n52853, n52854, n52855, n52856,
         n52857, n52858, n52859, n52860, n52861, n52862, n52863, n52864,
         n52865, n52866, n52868, n52869, n52870, n52871, n52872, n52873,
         n52874, n52876, n52878, n52879, n52880, n52881, n52882, n52883,
         n52884, n52885, n52886, n52887, n52888, n52889, n52890, n52892,
         n52893, n52894, n52895, n52896, n52897, n52898, n52899, n52900,
         n52901, n52903, n52904, n52905, n52906, n52907, n52908, n52909,
         n52910, n52911, n52912, n52913, n52914, n52916, n52917, n52918,
         n52919, n52920, n52921, n52922, n52923, n52924, n52925, n52926,
         n52927, n52928, n52929, n52930, n52931, n52932, n52933, n52935,
         n52937, n52938, n52940, n52943, n52944, n52945, n52946, n52948,
         n52949, n52950, n52951, n52952, n52953, n52954, n52955, n52957,
         n52958, n52959, n52961, n52962, n52963, n52964, n52965, n52966,
         n52967, n52968, n52969, n52970, n52972, n52973, n52974, n52975,
         n52976, n52977, n52978, n52979, n52980, n52982, n52983, n52984,
         n52985, n52986, n52987, n52988, n52989, n52990, n52992, n52993,
         n52994, n52995, n52996, n52997, n52998, n52999, n53000, n53001,
         n53002, n53003, n53004, n53005, n53006, n53007, n53008, n53009,
         n53010, n53011, n53012, n53013, n53014, n53015, n53016, n53017,
         n53018, n53019, n53020, n53021, n53022, n53023, n53024, n53025,
         n53026, n53027, n53029, n53030, n53031, n53032, n53033, n53034,
         n53035, n53036, n53037, n53038, n53039, n53040, n53041, n53042,
         n53043, n53044, n53045, n53046, n53047, n53048, n53049, n53050,
         n53051, n53052, n53053, n53054, n53055, n53056, n53057, n53058,
         n53059, n53060, n53061, n53062, n53063, n53064, n53066, n53067,
         n53068, n53070, n53071, n53072, n53073, n53074, n53075, n53076,
         n53077, n53078, n53079, n53080, n53081, n53082, n53083, n53084,
         n53085, n53086, n53087, n53088, n53089, n53090, n53091, n53092,
         n53093, n53094, n53095, n53096, n53097, n53098, n53099, n53100,
         n53101, n53102, n53103, n53104, n53105, n53106, n53107, n53108,
         n53109, n53110, n53111, n53112, n53113, n53114, n53115, n53116,
         n53117, n53118, n53119, n53120, n53121, n53122, n53123, n53124,
         n53126, n53127, n53128, n53129, n53130, n53131, n53132, n53133,
         n53135, n53136, n53137, n53138, n53139, n53140, n53141, n53142,
         n53143, n53144, n53145, n53146, n53147, n53148, n53149, n53150,
         n53153, n53154, n53155, n53156, n53157, n53158, n53159, n53160,
         n53161, n53162, n53163, n53164, n53165, n53166, n53167, n53168,
         n53169, n53170, n53171, n53172, n53173, n53174, n53175, n53176,
         n53177, n53178, n53179, n53180, n53181, n53182, n53183, n53184,
         n53185, n53186, n53187, n53188, n53189, n53190, n53192, n53193,
         n53194, n53195, n53196, n53197, n53198, n53199, n53200, n53201,
         n53202, n53203, n53204, n53205, n53206, n53207, n53208, n53209,
         n53212, n53213, n53214, n53215, n53216, n53218, n53219, n53220,
         n53221, n53222, n53223, n53224, n53225, n53226, n53227, n53228,
         n53229, n53230, n53231, n53232, n53233, n53234, n53235, n53236,
         n53237, n53238, n53239, n53240, n53241, n53242, n53243, n53244,
         n53246, n53247, n53248, n53249, n53250, n53251, n53252, n53253,
         n53254, n53255, n53257, n53258, n53259, n53260, n53261, n53262,
         n53264, n53265, n53266, n53267, n53268, n53269, n53270, n53271,
         n53272, n53273, n53274, n53275, n53276, n53277, n53278, n53279,
         n53280, n53281, n53282, n53283, n53284, n53285, n53286, n53287,
         n53288, n53289, n53291, n53292, n53293, n53294, n53295, n53296,
         n53297, n53298, n53300, n53301, n53302, n53303, n53304, n53305,
         n53306, n53307, n53308, n53309, n53310, n53311, n53312, n53313,
         n53314, n53315, n53316, n53317, n53318, n53319, n53320, n53321,
         n53322, n53323, n53324, n53325, n53326, n53327, n53328, n53329,
         n53331, n53332, n53333, n53334, n53335, n53336, n53337, n53338,
         n53339, n53340, n53341, n53342, n53344, n53345, n53346, n53347,
         n53348, n53349, n53350, n53351, n53352, n53353, n53354, n53355,
         n53356, n53357, n53358, n53359, n53361, n53362, n53363, n53364,
         n53365, n53366, n53368, n53369, n53370, n53371, n53372, n53373,
         n53374, n53375, n53376, n53377, n53378, n53379, n53380, n53381,
         n53382, n53383, n53384, n53385, n53386, n53387, n53388, n53389,
         n53390, n53391, n53392, n53393, n53394, n53395, n53396, n53397,
         n53398, n53399, n53400, n53402, n53403, n53404, n53405, n53406,
         n53407, n53408, n53409, n53410, n53411, n53412, n53413, n53414,
         n53415, n53416, n53417, n53418, n53419, n53420, n53421, n53422,
         n53423, n53424, n53425, n53426, n53427, n53428, n53429, n53430,
         n53431, n53432, n53433, n53434, n53435, n53436, n53437, n53438,
         n53439, n53440, n53441, n53442, n53443, n53444, n53445, n53446,
         n53447, n53448, n53449, n53450, n53451, n53452, n53454, n53455,
         n53456, n53457, n53458, n53459, n53460, n53461, n53462, n53463,
         n53464, n53465, n53466, n53467, n53468, n53469, n53470, n53471,
         n53472, n53473, n53474, n53475, n53476, n53477, n53478, n53479,
         n53480, n53481, n53482, n53483, n53484, n53485, n53486, n53487,
         n53489, n53490, n53491, n53492, n53493, n53494, n53495, n53496,
         n53497, n53498, n53499, n53500, n53501, n53502, n53503, n53504,
         n53505, n53506, n53507, n53508, n53509, n53510, n53511, n53512,
         n53513, n53514, n53515, n53516, n53517, n53518, n53519, n53520,
         n53521, n53522, n53523, n53524, n53525, n53526, n53527, n53528,
         n53529, n53530, n53531, n53532, n53533, n53534, n53535, n53536,
         n53537, n53538, n53539, n53540, n53541, n53542, n53543, n53544,
         n53545, n53546, n53547, n53548, n53549, n53551, n53552, n53554,
         n53555, n53556, n53557, n53558, n53559, n53560, n53561, n53562,
         n53563, n53564, n53565, n53566, n53567, n53568, n53569, n53570,
         n53572, n53575, n53576, n53577, n53578, n53580, n53581, n53582,
         n53583, n53584, n53585, n53586, n53587, n53588, n53589, n53590,
         n53591, n53592, n53593, n53594, n53595, n53596, n53597, n53598,
         n53600, n53601, n53602, n53603, n53604, n53605, n53606, n53607,
         n53608, n53609, n53610, n53611, n53612, n53613, n53614, n53615,
         n53616, n53617, n53618, n53619, n53620, n53621, n53622, n53623,
         n53624, n53625, n53626, n53627, n53628, n53629, n53630, n53631,
         n53632, n53633, n53634, n53635, n53636, n53637, n53638, n53639,
         n53640, n53641, n53642, n53643, n53644, n53645, n53646, n53647,
         n53648, n53649, n53650, n53651, n53652, n53653, n53654, n53655,
         n53656, n53657, n53658, n53659, n53660, n53661, n53662, n53663,
         n53664, n53665, n53666, n53667, n53668, n53669, n53670, n53671,
         n53672, n53673, n53674, n53675, n53676, n53677, n53678, n53679,
         n53680, n53682, n53683, n53684, n53685, n53687, n53688, n53689,
         n53690, n53691, n53692, n53693, n53694, n53695, n53696, n53697,
         n53698, n53699, n53700, n53701, n53702, n53703, n53704, n53705,
         n53706, n53707, n53708, n53709, n53711, n53712, n53713, n53714,
         n53715, n53716, n53717, n53718, n53719, n53720, n53721, n53723,
         n53724, n53725, n53726, n53727, n53728, n53729, n53730, n53731,
         n53732, n53733, n53734, n53735, n53736, n53737, n53738, n53739,
         n53740, n53741, n53742, n53743, n53744, n53745, n53746, n53747,
         n53748, n53749, n53750, n53751, n53752, n53753, n53754, n53755,
         n53756, n53757, n53758, n53759, n53761, n53762, n53763, n53764,
         n53765, n53766, n53767, n53768, n53770, n53771, n53772, n53773,
         n53774, n53775, n53776, n53777, n53778, n53779, n53780, n53781,
         n53782, n53783, n53784, n53785, n53786, n53787, n53789, n53790,
         n53791, n53792, n53793, n53794, n53795, n53796, n53797, n53798,
         n53799, n53800, n53801, n53802, n53803, n53804, n53805, n53807,
         n53808, n53809, n53810, n53811, n53812, n53813, n53814, n53815,
         n53816, n53817, n53818, n53819, n53820, n53821, n53822, n53823,
         n53824, n53825, n53826, n53827, n53828, n53829, n53830, n53831,
         n53832, n53833, n53834, n53835, n53836, n53837, n53841, n53843,
         n53844, n53845, n53847, n53848, n53849, n53850, n53851, n53852,
         n53853, n53854, n53855, n53856, n53857, n53858, n53859, n53860,
         n53861, n53862, n53863, n53864, n53865, n53867, n53868, n53869,
         n53870, n53871, n53872, n53873, n53875, n53876, n53877, n53878,
         n53879, n53880, n53881, n53882, n53883, n53884, n53885, n53886,
         n53887, n53888, n53889, n53890, n53891, n53892, n53893, n53894,
         n53895, n53896, n53897, n53899, n53900, n53901, n53902, n53903,
         n53904, n53905, n53906, n53907, n53908, n53909, n53910, n53911,
         n53912, n53913, n53914, n53915, n53916, n53917, n53918, n53919,
         n53920, n53921, n53922, n53923, n53924, n53925, n53926, n53927,
         n53928, n53929, n53930, n53931, n53932, n53933, n53935, n53936,
         n53937, n53938, n53939, n53940, n53941, n53942, n53943, n53944,
         n53945, n53946, n53947, n53948, n53949, n53950, n53951, n53952,
         n53953, n53955, n53956, n53957, n53958, n53959, n53960, n53961,
         n53962, n53964, n53965, n53966, n53967, n53968, n53969, n53970,
         n53971, n53972, n53973, n53974, n53975, n53976, n53977, n53979,
         n53980, n53981, n53982, n53983, n53984, n53985, n53986, n53987,
         n53988, n53989, n53991, n53992, n53993, n53994, n53995, n53996,
         n53997, n53998, n53999, n54000, n54001, n54002, n54003, n54004,
         n54006, n54007, n54009, n54010, n54012, n54013, n54014, n54015,
         n54016, n54017, n54018, n54019, n54020, n54021, n54022, n54023,
         n54024, n54025, n54026, n54027, n54028, n54029, n54030, n54031,
         n54032, n54033, n54034, n54035, n54036, n54037, n54039, n54041,
         n54043, n54044, n54045, n54046, n54047, n54048, n54049, n54050,
         n54051, n54052, n54053, n54054, n54055, n54056, n54057, n54058,
         n54059, n54060, n54061, n54062, n54063, n54064, n54065, n54066,
         n54067, n54068, n54069, n54070, n54071, n54072, n54073, n54074,
         n54075, n54077, n54079, n54081, n54082, n54083, n54084, n54085,
         n54086, n54087, n54088, n54089, n54090, n54091, n54092, n54093,
         n54094, n54095, n54096, n54097, n54098, n54100, n54102, n54103,
         n54104, n54105, n54106, n54107, n54108, n54109, n54110, n54111,
         n54112, n54113, n54115, n54116, n54117, n54118, n54119, n54120,
         n54121, n54122, n54123, n54124, n54125, n54126, n54127, n54128,
         n54130, n54131, n54132, n54133, n54134, n54135, n54136, n54137,
         n54138, n54139, n54140, n54141, n54143, n54144, n54145, n54146,
         n54147, n54148, n54149, n54150, n54151, n54152, n54153, n54155,
         n54156, n54157, n54158, n54159, n54160, n54161, n54162, n54165,
         n54166, n54167, n54168, n54169, n54170, n54171, n54172, n54173,
         n54174, n54175, n54176, n54177, n54178, n54179, n54180, n54181,
         n54182, n54183, n54184, n54185, n54186, n54187, n54188, n54189,
         n54190, n54191, n54192, n54193, n54194, n54195, n54196, n54197,
         n54198, n54199, n54200, n54201, n54202, n54203, n54204, n54205,
         n54207, n54208, n54209, n54210, n54211, n54212, n54213, n54214,
         n54215, n54216, n54217, n54218, n54219, n54221, n54222, n54223,
         n54224, n54225, n54226, n54227, n54228, n54229, n54230, n54231,
         n54232, n54233, n54234, n54235, n54236, n54237, n54238, n54239,
         n54240, n54241, n54242, n54243, n54244, n54245, n54246, n54247,
         n54248, n54249, n54250, n54251, n54252, n54253, n54254, n54255,
         n54256, n54257, n54258, n54259, n54260, n54261, n54262, n54263,
         n54264, n54265, n54266, n54267, n54268, n54269, n54270, n54271,
         n54272, n54273, n54274, n54275, n54276, n54277, n54278, n54280,
         n54281, n54282, n54284, n54285, n54286, n54287, n54288, n54289,
         n54291, n54292, n54294, n54295, n54296, n54297, n54298, n54299,
         n54300, n54302, n54303, n54304, n54305, n54307, n54308, n54309,
         n54310, n54311, n54312, n54314, n54316, n54317, n54318, n54319,
         n54320, n54321, n54322, n54323, n54324, n54325, n54326, n54327,
         n54328, n54330, n54331, n54332, n54333, n54334, n54335, n54336,
         n54337, n54338, n54340, n54341, n54342, n54343, n54344, n54345,
         n54346, n54347, n54348, n54349, n54350, n54351, n54352, n54353,
         n54354, n54355, n54356, n54357, n54358, n54359, n54360, n54361,
         n54362, n54363, n54364, n54365, n54366, n54367, n54368, n54369,
         n54370, n54371, n54372, n54373, n54374, n54375, n54376, n54377,
         n54378, n54379, n54380, n54381, n54382, n54383, n54384, n54385,
         n54386, n54387, n54388, n54390, n54391, n54392, n54393, n54394,
         n54395, n54396, n54397, n54399, n54400, n54401, n54402, n54403,
         n54404, n54405, n54406, n54407, n54408, n54409, n54410, n54411,
         n54412, n54413, n54414, n54415, n54417, n54418, n54419, n54420,
         n54421, n54422, n54423, n54424, n54425, n54426, n54427, n54428,
         n54429, n54430, n54431, n54432, n54433, n54434, n54435, n54436,
         n54437, n54438, n54439, n54440, n54441, n54442, n54443, n54444,
         n54445, n54446, n54447, n54448, n54450, n54451, n54452, n54453,
         n54454, n54455, n54456, n54457, n54459, n54460, n54461, n54462,
         n54463, n54464, n54465, n54466, n54467, n54468, n54469, n54470,
         n54471, n54472, n54473, n54474, n54475, n54476, n54477, n54478,
         n54479, n54480, n54481, n54482, n54483, n54484, n54485, n54486,
         n54487, n54488, n54489, n54490, n54492, n54493, n54494, n54495,
         n54496, n54498, n54499, n54500, n54501, n54502, n54503, n54504,
         n54505, n54506, n54507, n54508, n54510, n54511, n54512, n54513,
         n54514, n54515, n54517, n54520, n54522, n54523, n54524, n54525,
         n54526, n54527, n54528, n54529, n54530, n54531, n54532, n54533,
         n54534, n54535, n54536, n54537, n54538, n54539, n54540, n54541,
         n54542, n54543, n54544, n54545, n54546, n54547, n54548, n54549,
         n54550, n54551, n54552, n54553, n54554, n54555, n54556, n54558,
         n54559, n54560, n54561, n54562, n54563, n54564, n54565, n54566,
         n54567, n54568, n54569, n54570, n54571, n54572, n54573, n54574,
         n54575, n54576, n54577, n54578, n54579, n54580, n54581, n54582,
         n54583, n54584, n54585, n54587, n54588, n54589, n54590, n54591,
         n54592, n54593, n54594, n54595, n54596, n54597, n54598, n54599,
         n54600, n54601, n54602, n54603, n54604, n54605, n54606, n54607,
         n54608, n54609, n54610, n54611, n54612, n54613, n54614, n54615,
         n54616, n54617, n54618, n54619, n54620, n54621, n54622, n54623,
         n54624, n54625, n54626, n54627, n54628, n54629, n54630, n54631,
         n54632, n54633, n54634, n54635, n54636, n54637, n54638, n54639,
         n54640, n54641, n54643, n54645, n54646, n54647, n54648, n54649,
         n54650, n54651, n54652, n54653, n54654, n54655, n54656, n54657,
         n54658, n54659, n54660, n54661, n54662, n54664, n54665, n54666,
         n54667, n54668, n54669, n54670, n54671, n54672, n54673, n54674,
         n54675, n54676, n54677, n54678, n54679, n54680, n54681, n54682,
         n54683, n54684, n54685, n54686, n54687, n54688, n54689, n54690,
         n54691, n54692, n54693, n54694, n54695, n54696, n54697, n54698,
         n54699, n54700, n54701, n54702, n54703, n54704, n54705, n54706,
         n54707, n54708, n54709, n54710, n54711, n54712, n54713, n54714,
         n54715, n54716, n54717, n54718, n54719, n54720, n54721, n54722,
         n54723, n54724, n54725, n54726, n54727, n54728, n54729, n54730,
         n54731, n54732, n54733, n54734, n54735, n54736, n54737, n54738,
         n54739, n54740, n54741, n54742, n54743, n54744, n54745, n54746,
         n54747, n54748, n54749, n54750, n54751, n54752, n54753, n54754,
         n54755, n54756, n54757, n54758, n54759, n54761, n54762, n54763,
         n54764, n54766, n54767, n54768, n54769, n54770, n54771, n54772,
         n54773, n54774, n54775, n54776, n54777, n54778, n54779, n54780,
         n54781, n54782, n54783, n54784, n54785, n54786, n54787, n54788,
         n54789, n54790, n54791, n54792, n54793, n54794, n54796, n54797,
         n54798, n54799, n54801, n54802, n54803, n54804, n54805, n54806,
         n54807, n54809, n54810, n54811, n54813, n54814, n54815, n54816,
         n54817, n54818, n54819, n54821, n54822, n54823, n54824, n54825,
         n54826, n54827, n54829, n54830, n54831, n54832, n54835, n54838,
         n54839, n54840, n54841, n54842, n54843, n54844, n54845, n54846,
         n54847, n54848, n54849, n54852, n54853, n54854, n54855, n54857,
         n54858, n54859, n54860, n54861, n54862, n54863, n54866, n54867,
         n54868, n54869, n54870, n54871, n54872, n54873, n54874, n54875,
         n54876, n54877, n54879, n54880, n54881, n54882, n54883, n54884,
         n54885, n54886, n54887, n54888, n54890, n54891, n54892, n54893,
         n54894, n54895, n54896, n54898, n54899, n54900, n54901, n54902,
         n54903, n54904, n54905, n54906, n54907, n54908, n54909, n54911,
         n54912, n54913, n54914, n54915, n54916, n54917, n54918, n54919,
         n54920, n54921, n54922, n54923, n54925, n54926, n54927, n54928,
         n54929, n54930, n54931, n54932, n54933, n54934, n54935, n54936,
         n54938, n54939, n54941, n54942, n54943, n54944, n54945, n54948,
         n54949, n54950, n54951, n54952, n54953, n54954, n54955, n54956,
         n54957, n54958, n54959, n54960, n54961, n54963, n54964, n54965,
         n54966, n54967, n54968, n54970, n54971, n54972, n54973, n54974,
         n54975, n54976, n54977, n54978, n54979, n54980, n54981, n54982,
         n54983, n54984, n54987, n54989, n54990, n54991, n54992, n54993,
         n54994, n54995, n54996, n54997, n54998, n54999, n55000, n55001,
         n55002, n55003, n55004, n55005, n55006, n55007, n55008, n55009,
         n55011, n55012, n55013, n55014, n55015, n55016, n55017, n55018,
         n55019, n55020, n55021, n55022, n55023, n55024, n55025, n55026,
         n55027, n55029, n55030, n55031, n55032, n55033, n55034, n55035,
         n55036, n55037, n55038, n55039, n55040, n55041, n55042, n55043,
         n55044, n55045, n55046, n55047, n55048, n55049, n55050, n55051,
         n55052, n55053, n55054, n55056, n55057, n55058, n55059, n55060,
         n55061, n55062, n55063, n55064, n55065, n55066, n55067, n55068,
         n55069, n55070, n55071, n55074, n55075, n55076, n55077, n55078,
         n55079, n55080, n55081, n55082, n55084, n55085, n55086, n55087,
         n55088, n55089, n55090, n55092, n55094, n55095, n55096, n55097,
         n55098, n55099, n55101, n55102, n55103, n55104, n55105, n55106,
         n55107, n55108, n55110, n55111, n55112, n55113, n55114, n55115,
         n55116, n55117, n55118, n55119, n55120, n55121, n55122, n55123,
         n55124, n55125, n55126, n55127, n55128, n55129, n55130, n55131,
         n55132, n55133, n55134, n55135, n55136, n55137, n55138, n55139,
         n55140, n55141, n55142, n55143, n55144, n55145, n55146, n55147,
         n55148, n55149, n55150, n55151, n55152, n55153, n55154, n55155,
         n55156, n55157, n55158, n55159, n55160, n55161, n55162, n55163,
         n55164, n55165, n55166, n55167, n55168, n55169, n55170, n55171,
         n55172, n55173, n55174, n55175, n55176, n55177, n55178, n55179,
         n55180, n55181, n55182, n55183, n55184, n55185, n55186, n55187,
         n55189, n55190, n55191, n55192, n55193, n55195, n55196, n55197,
         n55198, n55199, n55200, n55201, n55202, n55203, n55204, n55205,
         n55206, n55207, n55208, n55209, n55210, n55211, n55212, n55214,
         n55215, n55216, n55217, n55218, n55219, n55221, n55222, n55223,
         n55224, n55225, n55226, n55227, n55228, n55229, n55230, n55231,
         n55232, n55233, n55234, n55235, n55236, n55237, n55238, n55239,
         n55240, n55241, n55242, n55244, n55245, n55246, n55247, n55248,
         n55249, n55250, n55252, n55253, n55254, n55255, n55256, n55257,
         n55258, n55259, n55260, n55261, n55262, n55263, n55264, n55265,
         n55266, n55267, n55268, n55269, n55270, n55271, n55272, n55273,
         n55275, n55276, n55277, n55278, n55279, n55280, n55281, n55282,
         n55283, n55284, n55285, n55286, n55287, n55288, n55289, n55290,
         n55291, n55292, n55293, n55294, n55295, n55296, n55297, n55298,
         n55299, n55300, n55301, n55302, n55303, n55304, n55305, n55306,
         n55307, n55308, n55309, n55310, n55311, n55312, n55315, n55316,
         n55317, n55318, n55319, n55320, n55321, n55322, n55323, n55324,
         n55326, n55327, n55329, n55331, n55332, n55333, n55334, n55335,
         n55336, n55337, n55338, n55339, n55340, n55341, n55342, n55343,
         n55345, n55346, n55347, n55349, n55350, n55351, n55352, n55353,
         n55354, n55355, n55356, n55358, n55359, n55360, n55361, n55362,
         n55363, n55364, n55365, n55366, n55367, n55368, n55369, n55370,
         n55371, n55372, n55373, n55374, n55375, n55376, n55377, n55378,
         n55379, n55380, n55381, n55382, n55383, n55384, n55385, n55386,
         n55387, n55388, n55389, n55391, n55392, n55394, n55395, n55396,
         n55397, n55398, n55399, n55400, n55401, n55402, n55403, n55404,
         n55406, n55407, n55408, n55410, n55411, n55412, n55413, n55414,
         n55415, n55416, n55417, n55418, n55419, n55420, n55421, n55423,
         n55424, n55425, n55426, n55427, n55428, n55429, n55430, n55431,
         n55432, n55433, n55434, n55435, n55436, n55437, n55438, n55439,
         n55440, n55441, n55442, n55443, n55444, n55445, n55446, n55447,
         n55448, n55449, n55450, n55451, n55452, n55453, n55454, n55455,
         n55456, n55457, n55458, n55459, n55460, n55461, n55462, n55463,
         n55465, n55466, n55468, n55469, n55470, n55471, n55472, n55473,
         n55474, n55475, n55476, n55477, n55478, n55479, n55480, n55481,
         n55483, n55484, n55485, n55486, n55487, n55488, n55489, n55491,
         n55492, n55493, n55494, n55495, n55496, n55497, n55498, n55499,
         n55500, n55501, n55502, n55503, n55504, n55505, n55506, n55507,
         n55508, n55509, n55510, n55511, n55512, n55513, n55514, n55515,
         n55516, n55518, n55519, n55520, n55521, n55522, n55523, n55524,
         n55525, n55526, n55527, n55528, n55529, n55530, n55531, n55532,
         n55533, n55534, n55535, n55537, n55538, n55539, n55540, n55541,
         n55542, n55543, n55544, n55545, n55546, n55547, n55548, n55549,
         n55550, n55551, n55552, n55553, n55554, n55555, n55556, n55557,
         n55558, n55559, n55560, n55561, n55562, n55563, n55564, n55565,
         n55566, n55567, n55568, n55569, n55570, n55571, n55572, n55573,
         n55574, n55575, n55576, n55577, n55578, n55579, n55580, n55581,
         n55582, n55583, n55584, n55585, n55586, n55587, n55588, n55589,
         n55590, n55591, n55592, n55593, n55594, n55595, n55596, n55597,
         n55598, n55599, n55600, n55601, n55602, n55603, n55604, n55607,
         n55608, n55609, n55610, n55611, n55612, n55613, n55614, n55615,
         n55616, n55617, n55618, n55619, n55620, n55621, n55622, n55623,
         n55624, n55625, n55626, n55627, n55628, n55629, n55630, n55631,
         n55632, n55633, n55634, n55635, n55636, n55637, n55638, n55639,
         n55640, n55641, n55642, n55643, n55644, n55645, n55646, n55647,
         n55648, n55649, n55650, n55651, n55652, n55653, n55654, n55655,
         n55656, n55657, n55658, n55659, n55660, n55661, n55662, n55663,
         n55664, n55665, n55666, n55667, n55668, n55669, n55670, n55671,
         n55672, n55673, n55674, n55675, n55676, n55677, n55678, n55679,
         n55680, n55681, n55682, n55683, n55684, n55685, n55686, n55687,
         n55688, n55689, n55690, n55691, n55692, n55693, n55694, n55695,
         n55696, n55697, n55698, n55699, n55700, n55701, n55702, n55703,
         n55704, n55705, n55706, n55707, n55708, n55709, n55710, n55711,
         n55712, n55713, n55714, n55715, n55716, n55717, n55718, n55719,
         n55720, n55721, n55722, n55724, n55725, n55726, n55727, n55728,
         n55729, n55730, n55731, n55732, n55733, n55734, n55735, n55737,
         n55738, n55739, n55740, n55741, n55742, n55744, n55746, n55747,
         n55748, n55749, n55750, n55751, n55752, n55753, n55754, n55755,
         n55756, n55757, n55758, n55759, n55760, n55761, n55762, n55763,
         n55764, n55765, n55766, n55767, n55768, n55769, n55770, n55771,
         n55772, n55773, n55774, n55775, n55776, n55777, n55778, n55779,
         n55780, n55781, n55782, n55783, n55784, n55786, n55788, n55789,
         n55790, n55791, n55792, n55793, n55794, n55795, n55796, n55797,
         n55799, n55800, n55801, n55802, n55803, n55804, n55805, n55806,
         n55807, n55808, n55809, n55810, n55811, n55812, n55813, n55814,
         n55815, n55816, n55817, n55818, n55819, n55820, n55821, n55822,
         n55824, n55825, n55826, n55827, n55828, n55829, n55831, n55832,
         n55833, n55834, n55835, n55836, n55837, n55838, n55839, n55840,
         n55842, n55843, n55844, n55845, n55846, n55847, n55850, n55851,
         n55852, n55853, n55854, n55855, n55856, n55857, n55858, n55859,
         n55860, n55861, n55862, n55863, n55864, n55865, n55866, n55867,
         n55868, n55869, n55870, n55871, n55872, n55873, n55874, n55875,
         n55876, n55877, n55878, n55879, n55880, n55881, n55882, n55883,
         n55884, n55885, n55886, n55887, n55888, n55889, n55890, n55891,
         n55892, n55893, n55894, n55895, n55896, n55897, n55898, n55899,
         n55900, n55901, n55902, n55903, n55904, n55905, n55906, n55908,
         n55909, n55910, n55911, n55912, n55913, n55914, n55915, n55916,
         n55917, n55918, n55919, n55920, n55921, n55922, n55923, n55924,
         n55925, n55926, n55927, n55928, n55930, n55931, n55932, n55933,
         n55934, n55935, n55936, n55937, n55938, n55939, n55940, n55941,
         n55942, n55944, n55947, n55948, n55949, n55950, n55951, n55952,
         n55953, n55955, n55956, n55957, n55958, n55961, n55962, n55964,
         n55965, n55966, n55967, n55968, n55969, n55970, n55971, n55972,
         n55973, n55974, n55975, n55976, n55977, n55978, n55979, n55980,
         n55981, n55982, n55983, n55984, n55985, n55986, n55987, n55988,
         n55989, n55990, n55991, n55992, n55993, n55994, n55995, n55996,
         n55997, n55998, n55999, n56000, n56001, n56002, n56003, n56004,
         n56005, n56006, n56007, n56008, n56009, n56010, n56011, n56012,
         n56013, n56014, n56015, n56017, n56018, n56019, n56020, n56023,
         n56024, n56025, n56026, n56027, n56028, n56029, n56030, n56031,
         n56032, n56033, n56034, n56035, n56036, n56037, n56038, n56039,
         n56040, n56041, n56042, n56043, n56044, n56045, n56046, n56047,
         n56048, n56049, n56050, n56051, n56052, n56053, n56054, n56055,
         n56056, n56057, n56058, n56059, n56060, n56061, n56062, n56063,
         n56064, n56065, n56066, n56067, n56068, n56069, n56070, n56071,
         n56072, n56073, n56074, n56075, n56076, n56077, n56078, n56079,
         n56080, n56081, n56082, n56083, n56084, n56085, n56087, n56088,
         n56089, n56090, n56091, n56092, n56093, n56094, n56095, n56096,
         n56097, n56098, n56099, n56100, n56101, n56102, n56103, n56104,
         n56105, n56106, n56107, n56108, n56110, n56111, n56112, n56113,
         n56114, n56115, n56117, n56118, n56119, n56120, n56121, n56122,
         n56123, n56124, n56125, n56126, n56127, n56128, n56129, n56130,
         n56131, n56132, n56133, n56134, n56135, n56136, n56137, n56138,
         n56139, n56140, n56141, n56142, n56143, n56144, n56145, n56146,
         n56147, n56148, n56149, n56150, n56151, n56152, n56153, n56154,
         n56155, n56157, n56158, n56159, n56160, n56161, n56162, n56163,
         n56164, n56165, n56166, n56167, n56168, n56169, n56170, n56171,
         n56172, n56173, n56174, n56175, n56176, n56177, n56178, n56179,
         n56180, n56181, n56182, n56183, n56184, n56185, n56186, n56187,
         n56188, n56189, n56190, n56191, n56192, n56194, n56195, n56196,
         n56197, n56198, n56199, n56200, n56201, n56202, n56203, n56204,
         n56205, n56206, n56207, n56208, n56209, n56210, n56211, n56212,
         n56213, n56214, n56215, n56216, n56217, n56218, n56219, n56220,
         n56221, n56222, n56223, n56224, n56225, n56226, n56227, n56228,
         n56229, n56230, n56231, n56232, n56233, n56234, n56235, n56236,
         n56237, n56238, n56239, n56240, n56241, n56242, n56243, n56244,
         n56245, n56246, n56247, n56248, n56249, n56250, n56251, n56252,
         n56253, n56254, n56255, n56256, n56257, n56258, n56259, n56260,
         n56261, n56263, n56264, n56265, n56266, n56267, n56268, n56269,
         n56270, n56271, n56272, n56273, n56274, n56275, n56276, n56277,
         n56278, n56279, n56280, n56281, n56282, n56283, n56284, n56285,
         n56286, n56287, n56288, n56289, n56290, n56291, n56292, n56293,
         n56294, n56295, n56296, n56297, n56298, n56299, n56300, n56301,
         n56302, n56303, n56304, n56305, n56306, n56307, n56308, n56309,
         n56311, n56312, n56313, n56314, n56315, n56316, n56317, n56318,
         n56319, n56320, n56321, n56322, n56323, n56324, n56325, n56326,
         n56327, n56328, n56329, n56330, n56331, n56332, n56333, n56334,
         n56335, n56336, n56338, n56339, n56340, n56341, n56342, n56343,
         n56344, n56346, n56347, n56348, n56349, n56350, n56351, n56352,
         n56353, n56355, n56356, n56357, n56358, n56359, n56360, n56361,
         n56362, n56363, n56364, n56365, n56367, n56368, n56369, n56370,
         n56371, n56372, n56373, n56374, n56375, n56377, n56379, n56380,
         n56381, n56382, n56383, n56384, n56385, n56386, n56387, n56388,
         n56389, n56390, n56391, n56392, n56393, n56394, n56396, n56397,
         n56398, n56399, n56401, n56402, n56403, n56404, n56405, n56406,
         n56407, n56408, n56409, n56411, n56412, n56413, n56414, n56415,
         n56417, n56418, n56419, n56420, n56421, n56422, n56423, n56424,
         n56425, n56426, n56428, n56430, n56431, n56432, n56433, n56434,
         n56435, n56436, n56437, n56438, n56439, n56440, n56441, n56443,
         n56444, n56445, n56446, n56448, n56451, n56452, n56453, n56454,
         n56455, n56456, n56457, n56458, n56459, n56460, n56461, n56462,
         n56463, n56464, n56465, n56466, n56467, n56468, n56469, n56470,
         n56472, n56473, n56474, n56475, n56476, n56477, n56478, n56479,
         n56480, n56481, n56482, n56483, n56484, n56485, n56486, n56487,
         n56488, n56489, n56490, n56491, n56492, n56493, n56494, n56495,
         n56496, n56497, n56498, n56499, n56500, n56501, n56502, n56503,
         n56504, n56505, n56506, n56507, n56508, n56509, n56510, n56511,
         n56512, n56513, n56514, n56516, n56517, n56518, n56519, n56520,
         n56521, n56522, n56523, n56524, n56525, n56526, n56529, n56530,
         n56531, n56532, n56533, n56534, n56536, n56537, n56538, n56539,
         n56540, n56541, n56542, n56543, n56544, n56545, n56546, n56547,
         n56548, n56549, n56550, n56551, n56552, n56553, n56554, n56555,
         n56556, n56557, n56558, n56559, n56560, n56562, n56563, n56564,
         n56565, n56566, n56567, n56568, n56569, n56570, n56571, n56572,
         n56573, n56574, n56575, n56579, n56580, n56581, n56582, n56583,
         n56584, n56585, n56586, n56587, n56588, n56590, n56591, n56592,
         n56593, n56594, n56595, n56596, n56597, n56598, n56599, n56600,
         n56601, n56602, n56604, n56605, n56606, n56607, n56608, n56609,
         n56610, n56611, n56612, n56613, n56614, n56615, n56616, n56619,
         n56620, n56621, n56622, n56623, n56624, n56626, n56627, n56628,
         n56629, n56630, n56631, n56632, n56633, n56634, n56635, n56636,
         n56637, n56638, n56639, n56640, n56641, n56642, n56644, n56645,
         n56646, n56647, n56648, n56649, n56651, n56652, n56653, n56654,
         n56658, n56659, n56660, n56661, n56662, n56663, n56664, n56665,
         n56666, n56667, n56668, n56669, n56670, n56672, n56673, n56674,
         n56676, n56677, n56678, n56679, n56680, n56681, n56682, n56683,
         n56684, n56685, n56686, n56687, n56688, n56689, n56690, n56691,
         n56692, n56693, n56694, n56695, n56696, n56697, n56698, n56699,
         n56700, n56701, n56702, n56703, n56704, n56705, n56706, n56707,
         n56708, n56710, n56711, n56712, n56713, n56714, n56716, n56717,
         n56718, n56719, n56721, n56722, n56723, n56724, n56725, n56726,
         n56727, n56728, n56729, n56730, n56731, n56732, n56733, n56734,
         n56735, n56736, n56737, n56738, n56739, n56740, n56741, n56742,
         n56743, n56744, n56745, n56746, n56747, n56749, n56751, n56752,
         n56753, n56754, n56755, n56756, n56757, n56758, n56759, n56760,
         n56761, n56762, n56763, n56764, n56765, n56766, n56767, n56768,
         n56769, n56770, n56771, n56772, n56773, n56774, n56775, n56776,
         n56777, n56778, n56779, n56780, n56781, n56782, n56783, n56784,
         n56785, n56786, n56787, n56788, n56789, n56790, n56791, n56792,
         n56793, n56795, n56796, n56797, n56799, n56800, n56802, n56803,
         n56804, n56805, n56806, n56807, n56808, n56809, n56810, n56812,
         n56813, n56814, n56815, n56816, n56817, n56818, n56819, n56820,
         n56821, n56822, n56823, n56824, n56825, n56826, n56827, n56829,
         n56830, n56831, n56832, n56833, n56834, n56836, n56837, n56838,
         n56839, n56840, n56841, n56842, n56843, n56844, n56845, n56846,
         n56848, n56849, n56850, n56851, n56852, n56853, n56854, n56855,
         n56856, n56857, n56858, n56859, n56860, n56861, n56862, n56863,
         n56864, n56865, n56866, n56867, n56868, n56869, n56870, n56871,
         n56872, n56873, n56874, n56875, n56876, n56877, n56879, n56880,
         n56881, n56882, n56883, n56884, n56885, n56886, n56887, n56888,
         n56889, n56890, n56891, n56892, n56893, n56894, n56895, n56896,
         n56897, n56899, n56900, n56901, n56902, n56903, n56904, n56905,
         n56906, n56907, n56908, n56909, n56910, n56911, n56913, n56914,
         n56915, n56916, n56917, n56918, n56919, n56921, n56922, n56923,
         n56924, n56925, n56926, n56928, n56929, n56930, n56931, n56933,
         n56935, n56936, n56937, n56939, n56940, n56941, n56942, n56943,
         n56944, n56945, n56946, n56947, n56948, n56949, n56950, n56952,
         n56953, n56954, n56955, n56956, n56957, n56958, n56959, n56960,
         n56961, n56962, n56963, n56964, n56965, n56966, n56967, n56968,
         n56970, n56971, n56972, n56973, n56974, n56975, n56976, n56977,
         n56978, n56979, n56980, n56981, n56982, n56983, n56984, n56985,
         n56986, n56987, n56988, n56989, n56990, n56991, n56992, n56993,
         n56995, n56996, n56997, n56998, n56999, n57000, n57001, n57002,
         n57004, n57005, n57006, n57007, n57008, n57009, n57010, n57011,
         n57012, n57013, n57014, n57015, n57017, n57018, n57019, n57020,
         n57022, n57023, n57024, n57025, n57026, n57027, n57029, n57030,
         n57031, n57032, n57034, n57035, n57036, n57037, n57038, n57039,
         n57040, n57041, n57042, n57043, n57044, n57046, n57047, n57048,
         n57049, n57050, n57051, n57052, n57053, n57054, n57055, n57056,
         n57057, n57058, n57060, n57061, n57062, n57063, n57064, n57065,
         n57066, n57067, n57068, n57069, n57070, n57072, n57073, n57074,
         n57075, n57076, n57078, n57079, n57081, n57083, n57084, n57086,
         n57087, n57088, n57089, n57090, n57091, n57092, n57093, n57094,
         n57095, n57096, n57097, n57098, n57099, n57101, n57102, n57104,
         n57105, n57106, n57107, n57108, n57109, n57110, n57111, n57112,
         n57113, n57114, n57115, n57116, n57119, n57120, n57121, n57122,
         n57123, n57124, n57125, n57126, n57127, n57128, n57129, n57130,
         n57131, n57132, n57133, n57134, n57135, n57136, n57137, n57138,
         n57140, n57142, n57143, n57144, n57146, n57148, n57149, n57150,
         n57153, n57154, n57155, n57156, n57157, n57158, n57159, n57160,
         n57161, n57162, n57164, n57165, n57166, n57167, n57168, n57169,
         n57171, n57172, n57173, n57174, n57175, n57177, n57178, n57179,
         n57182, n57183, n57184, n57185, n57186, n57187, n57191, n57192,
         n57193, n57194, n57195, n57196, n57197, n57198, n57199, n57200,
         n57201, n57202, n57203, n57204, n57205, n57207, n57208, n57209,
         n57210, n57211, n57212, n57213, n57214, n57216, n57217, n57218,
         n57219, n57220, n57221, n57222, n57223, n57224, n57225, n57226,
         n57227, n57228, n57229, n57230, n57231, n57232, n57233, n57234,
         n57235, n57236, n57237, n57238, n57239, n57240, n57241, n57243,
         n57244, n57245, n57247, n57248, n57249, n57250, n57251, n57252,
         n57253, n57254, n57255, n57256, n57257, n57258, n57259, n57260,
         n57261, n57262, n57263, n57264, n57265, n57266, n57267, n57268,
         n57269, n57270, n57271, n57272, n57273, n57274, n57275, n57276,
         n57277, n57278, n57279, n57280, n57281, n57282, n57283, n57285,
         n57287, n57288, n57289, n57290, n57291, n57292, n57293, n57294,
         n57295, n57296, n57297, n57298, n57299, n57300, n57301, n57302,
         n57303, n57304, n57305, n57306, n57309, n57310, n57311, n57312,
         n57313, n57314, n57315, n57316, n57317, n57318, n57319, n57320,
         n57321, n57322, n57323, n57324, n57325, n57326, n57327, n57328,
         n57329, n57330, n57331, n57332, n57333, n57334, n57335, n57336,
         n57337, n57338, n57339, n57340, n57341, n57342, n57344, n57345,
         n57346, n57347, n57348, n57349, n57350, n57351, n57352, n57353,
         n57354, n57355, n57356, n57357, n57358, n57359, n57360, n57361,
         n57363, n57364, n57365, n57366, n57367, n57368, n57369, n57370,
         n57371, n57372, n57373, n57375, n57376, n57377, n57378, n57379,
         n57380, n57381, n57382, n57383, n57385, n57387, n57388, n57389,
         n57390, n57391, n57392, n57393, n57394, n57395, n57396, n57397,
         n57398, n57399, n57400, n57401, n57402, n57403, n57404, n57405,
         n57406, n57407, n57408, n57409, n57410, n57411, n57412, n57413,
         n57414, n57415, n57416, n57417, n57419, n57420, n57421, n57423,
         n57424, n57425, n57426, n57427, n57428, n57429, n57430, n57431,
         n57432, n57433, n57434, n57435, n57436, n57437, n57438, n57439,
         n57440, n57441, n57442, n57443, n57444, n57445, n57446, n57447,
         n57448, n57450, n57451, n57452, n57453, n57454, n57455, n57456,
         n57458, n57459, n57461, n57462, n57463, n57465, n57466, n57467,
         n57468, n57470, n57471, n57473, n57474, n57476, n57477, n57479,
         n57480, n57481, n57482, n57483, n57485, n57486, n57487, n57488,
         n57489, n57490, n57492, n57494, n57495, n57496, n57497, n57499,
         n57501, n57502, n57507, n57508, n57509, n57510, n57514, n57515,
         n57517, n57519, n57521, n57522, n57523, n57525, n57526, n57528,
         n57529, n57530, n57531, n57532, n57534, n57535, n57536, n57537,
         n57538, n57541, n57542, n57543, n57544, n57545, n57546, n57547,
         n57549, n57550, n57551, n57553, n57555, n57557, n57558, n57559,
         n57563, n57564, n57566, n57568, n57569, n57570, n57571, n57572,
         n57573, n57574, n57576, n57577, n57580, n57582, n57586, n57587,
         n57589, n57590, n57591, n57592, n57593, n57595, n57596, n57597,
         n57598, n57599, n57600, n57603, n57605, n57606, n57607, n57608,
         n57609, n57610, n57611, n57612, n57613, n57614, n57615, n57616,
         n57617, n57618, n57619, n57620, n57621, n57622, n57623, n57624,
         n57625, n57626, n57628, n57629, n57630, n57631, n57632, n57633,
         n57634, n57635, n57636, n57637, n57638, n57639, n57640, n57641,
         n57644, n57647, n57648, n57649, n57651, n57652, n57654, n57655,
         n57656, n57657, n57658, n57660, n57664, n57665, n57666, n57667,
         n57668, n57669, n57670, n57672, n57673, n57674, n57675, n57676,
         n57677, n57678, n57679, n57680, n57681, n57682, n57683, n57684,
         n57685, n57686, n57687, n57688, n57689, n57690, n57691, n57692,
         n57693, n57694, n57695, n57696, n57697, n57698, n57699, n57700,
         n57701, n57704, n57705, n57706, n57707, n57708, n57709, n57710,
         n57711, n57714, n57716, n57717, n57719, n57720, n57721, n57722,
         n57723, n57727, n57728, n57729, n57730, n57731, n57732, n57733,
         n57734, n57735, n57738, n57739, n57740, n57742, n57744, n57746,
         n57747, n57748, n57749, n57750, n57751, n57752, n57753, n57754,
         n57755, n57756, n57757, n57758, n57759, n57760, n57762, n57764,
         n57766, n57768, n57769, n57772, n57773, n57774, n57775, n57776,
         n57777, n57778, n57780, n57781, n57782, n57783, n57784, n57785,
         n57786, n57788, n57789, n57790, n57791, n57792, n57796, n57799,
         n57802, n57803, n57805, n57806, n57808, n57809, n57810, n57812,
         n57815, n57816, n57819, n57820, n57821, n57822, n57824, n57826,
         n57827, n57828, n57829, n57830, n57831, n57832, n57836, n57837,
         n57838, n57839, n57842, n57844, n57845, n57846, n57847, n57848,
         n57851, n57852, n57854, n57856, n57857, n57860, n57861, n57862,
         n57863, n57864, n57865, n57866, n57868, n57869, n57870, n57871,
         n57872, n57873, n57874, n57875, n57876, n57878, n57881, n57882,
         n57883, n57884, n57885, n57886, n57888, n57889, n57890, n57892,
         n57893, n57894, n57896, n57898, n57899, n57900, n57901, n57907,
         n57908, n57909, n57910, n57911, n57912, n57914, n57915, n57918,
         n57919, n57920, n57921, n57922, n57924, n57925, n57926, n57927,
         n57930, n57931, n57932, n57935, n57936, n57937, n57938, n57939,
         n57940, n57941, n57944, n57945, n57947, n57948, n57949, n57950,
         n57951, n57952, n57953, n57954, n57955, n57956, n57957, n57958,
         n57960, n57962, n57963, n57964, n57965, n57966, n57967, n57970,
         n57971, n57972, n57973, n57974, n57975, n57976, n57978, n57979,
         n57983, n57984, n57985, n57986, n57987, n57988, n57989, n57990,
         n57991, n57992, n57993, n57995, n57996, n57997, n57998, n57999,
         n58000, n58001, n58002, n58004, n58005, n58006, n58009, n58013,
         n58014, n58016, n58017, n58018, n58019, n58020, n58022, n58024,
         n58025, n58026, n58027, n58029, n58030, n58031, n58032, n58033,
         n58035, n58036, n58037, n58039, n58040, n58042, n58043, n58045,
         n58046, n58047, n58048, n58050, n58051, n58052, n58053, n58055,
         n58058, n58059, n58060, n58061, n58062, n58064, n58065, n58068,
         n58069, n58073, n58074, n58075, n58076, n58077, n58078, n58079,
         n58080, n58081, n58082, n58083, n58084, n58085, n58086, n58088,
         n58089, n58090, n58091, n58092, n58094, n58095, n58096, n58097,
         n58098, n58099, n58102, n58103, n58104, n58105, n58107, n58108,
         n58109, n58111, n58112, n58113, n58115, n58116, n58117, n58119,
         n58122, n58123, n58124, n58125, n58127, n58128, n58129, n58130,
         n58131, n58132, n58133, n58134, n58135, n58136, n58137, n58139,
         n58140, n58145, n58146, n58147, n58148, n58150, n58151, n58152,
         n58153, n58154, n58155, n58156, n58157, n58158, n58160, n58161,
         n58162, n58163, n58164, n58168, n58169, n58171, n58172, n58174,
         n58175, n58176, n58177, n58178, n58179, n58180, n58184, n58185,
         n58186, n58187, n58189, n58191, n58192, n58193, n58195, n58198,
         n58199, n58201, n58203, n58204, n58205, n58206, n58207, n58208,
         n58209, n58210, n58211, n58212, n58213, n58214, n58215, n58218,
         n58220, n58221, n58222, n58223, n58225, n58226, n58227, n58229,
         n58231, n58232, n58233, n58234, n58235, n58236, n58237, n58238,
         n58240, n58241, n58243, n58244, n58245, n58246, n58247, n58248,
         n58249, n58250, n58252, n58254, n58255, n58257, n58258, n58259,
         n58261, n58262, n58264, n58265, n58267, n58269, n58271, n58272,
         n58273, n58274, n58275, n58277, n58279, n58280, n58281, n58282,
         n58283, n58284, n58285, n58286, n58288, n58289, n58290, n58292,
         n58293, n58294, n58296, n58297, n58298, n58299, n58300, n58301,
         n58302, n58303, n58304, n58305, n58306, n58307, n58309, n58310,
         n58312, n58313, n58316, n58318, n58320, n58321, n58322, n58323,
         n58324, n58325, n58326, n58327, n58328, n58330, n58332, n58333,
         n58335, n58336, n58338, n58339, n58340, n58341, n58343, n58346,
         n58347, n58348, n58349, n58351, n58352, n58353, n58354, n58355,
         n58357, n58364, n58365, n58366, n58367, n58368, n58369, n58370,
         n58371, n58372, n58373, n58375, n58377, n58378, n58379, n58380,
         n58382, n58384, n58385, n58386, n58387, n58388, n58390, n58392,
         n58393, n58394, n58395, n58396, n58398, n58399, n58400, n58401,
         n58402, n58404, n58406, n58407, n58408, n58409, n58414, n58415,
         n58416, n58417, n58418, n58419, n58420, n58421, n58422, n58423,
         n58424, n58426, n58427, n58428, n58429, n58430, n58431, n58432,
         n58433, n58434, n58435, n58437, n58440, n58442, n58443, n58444,
         n58445, n58446, n58447, n58448, n58449, n58450, n58451, n58453,
         n58455, n58456, n58457, n58460, n58461, n58462, n58463, n58466,
         n58467, n58468, n58470, n58472, n58473, n58474, n58475, n58476,
         n58477, n58479, n58480, n58481, n58483, n58484, n58485, n58486,
         n58488, n58489, n58490, n58491, n58492, n58498, n58499, n58500,
         n58502, n58503, n58504, n58505, n58506, n58510, n58511, n58513,
         n58514, n58517, n58518, n58519, n58520, n58521, n58522, n58524,
         n58525, n58526, n58527, n58528, n58529, n58530, n58531, n58532,
         n58533, n58534, n58535, n58537, n58538, n58540, n58541, n58544,
         n58546, n58548, n58549, n58550, n58551, n58552, n58553, n58555,
         n58557, n58559, n58560, n58561, n58562, n58563, n58564, n58565,
         n58567, n58568, n58570, n58571, n58572, n58573, n58574, n58575,
         n58577, n58578, n58580, n58581, n58582, n58583, n58584, n58585,
         n58586, n58587, n58588, n58589, n58591, n58594, n58596, n58598,
         n58599, n58601, n58603, n58604, n58606, n58608, n58609, n58610,
         n58612, n58613, n58615, n58616, n58617, n58618, n58619, n58620,
         n58621, n58624, n58625, n58626, n58628, n58629, n58630, n58633,
         n58634, n58635, n58636, n58637, n58639, n58640, n58641, n58644,
         n58645, n58646, n58647, n58648, n58649, n58650, n58651, n58653,
         n58654, n58655, n58656, n58657, n58660, n58661, n58663, n58664,
         n58665, n58666, n58667, n58668, n58669, n58672, n58674, n58675,
         n58676, n58678, n58680, n58681, n58683, n58684, n58685, n58687,
         n58688, n58689, n58690, n58691, n58692, n58693, n58694, n58695,
         n58696, n58697, n58700, n58701, n58702, n58703, n58704, n58705,
         n58708, n58710, n58713, n58715, n58716, n58717, n58718, n58720,
         n58721, n58722, n58723, n58725, n58727, n58728, n58729, n58730,
         n58731, n58732, n58734, n58735, n58736, n58738, n58740, n58743,
         n58744, n58745, n58747, n58748, n58749, n58750, n58751, n58753,
         n58754, n58755, n58756, n58757, n58759, n58760, n58762, n58763,
         n58764, n58765, n58766, n58767, n58768, n58769, n58770, n58771,
         n58772, n58775, n58776, n58777, n58780, n58781, n58782, n58783,
         n58784, n58785, n58787, n58789, n58790, n58791, n58792, n58793,
         n58794, n58795, n58796, n58797, n58798, n58799, n58800, n58801,
         n58802, n58806, n58807, n58808, n58809, n58810, n58811, n58812,
         n58813, n58814, n58815, n58816, n58817, n58818, n58819, n58822,
         n58823, n58824, n58825, n58826, n58827, n58828, n58829, n58830,
         n58831, n58832, n58834, n58835, n58836, n58837, n58838, n58839,
         n58840, n58841, n58842, n58843, n58844, n58845, n58846, n58850,
         n58851, n58852, n58853, n58855, n58856, n58858, n58859, n58860,
         n58861, n58862, n58863, n58864, n58867, n58868, n58869, n58871,
         n58872, n58873, n58874, n58876, n58878, n58879, n58880, n58881,
         n58882, n58883, n58884, n58885, n58886, n58888, n58889, n58891,
         n58892, n58895, n58896, n58897, n58898, n58900, n58904, n58905,
         n58907, n58908, n58909, n58910, n58912, n58913, n58914, n58916,
         n58917, n58918, n58920, n58921, n58922, n58923, n58924, n58925,
         n58926, n58927, n58928, n58929, n58931, n58932, n58933, n58934,
         n58937, n58938, n58939, n58940, n58941, n58942, n58943, n58944,
         n58945, n58946, n58947, n58949, n58954, n58955, n58957, n58958,
         n58959, n58961, n58962, n58963, n58964, n58965, n58967, n58968,
         n58969, n58970, n58971, n58972, n58974, n58975, n58976, n58977,
         n58978, n58980, n58981, n58983, n58984, n58985, n58987, n58988,
         n58989, n58990, n58991, n58994, n58995, n58996, n58997, n58998,
         n58999, n59000, n59001, n59003, n59004, n59005, n59006, n59008,
         n59009, n59011, n59012, n59013, n59014, n59015, n59016, n59017,
         n59018, n59019, n59020, n59021, n59023, n59024, n59026, n59028,
         n59029, n59030, n59032, n59034, n59035, n59036, n59037, n59038,
         n59039, n59040, n59041, n59043, n59044, n59045, n59046, n59048,
         n59049, n59051, n59052, n59053, n59056, n59057, n59058, n59059,
         n59062, n59063, n59064, n59065, n59066, n59067, n59068, n59069,
         n59071, n59072, n59074, n59075, n59076, n59078, n59079, n59080,
         n59081, n59082, n59083, n59084, n59085, n59086, n59087, n59088,
         n59089, n59090, n59091, n59093, n59094, n59095, n59096, n59097,
         n59098, n59099, n59100, n59101, n59102, n59103, n59104, n59105,
         n59106, n59107, n59108, n59109, n59110, n59113, n59115, n59116,
         n59117, n59119, n59120, n59121, n59122, n59123, n59125, n59126,
         n59127, n59128, n59129, n59130, n59131, n59134, n59135, n59136,
         n59137, n59138, n59139, n59140, n59141, n59142, n59143, n59146,
         n59147, n59149, n59150, n59151, n59153, n59154, n59155, n59156,
         n59157, n59158, n59159, n59160, n59163, n59165, n59166, n59167,
         n59168, n59169, n59172, n59173, n59174, n59175, n59176, n59177,
         n59179, n59180, n59181, n59183, n59184, n59185, n59186, n59188,
         n59190, n59192, n59193, n59195, n59196, n59197, n59198, n59199,
         n59200, n59202, n59203, n59205, n59206, n59207, n59208, n59209,
         n59210, n59211, n59212, n59214, n59215, n59216, n59217, n59218,
         n59221, n59222, n59224, n59225, n59226, n59227, n59228, n59229,
         n59230, n59231, n59232, n59233, n59236, n59237, n59238, n59239,
         n59240, n59241, n59244, n59245, n59248, n59249, n59250, n59252,
         n59255, n59256, n59257, n59258, n59259, n59260, n59261, n59262,
         n59263, n59264, n59266, n59267, n59268, n59269, n59270, n59271,
         n59272, n59273, n59274, n59275, n59276, n59277, n59279, n59280,
         n59281, n59282, n59284, n59285, n59286, n59287, n59288, n59289,
         n59291, n59292, n59293, n59294, n59296, n59297, n59298, n59299,
         n59300, n59301, n59302, n59303, n59305, n59306, n59307, n59309,
         n59310, n59311, n59312, n59315, n59316, n59317, n59319, n59320,
         n59321, n59322, n59323, n59324, n59325, n59326, n59328, n59329,
         n59330, n59331, n59332, n59333, n59334, n59335, n59336, n59337,
         n59340, n59341, n59342, n59343, n59344, n59345, n59346, n59347,
         n59348, n59351, n59354, n59355, n59356, n59358, n59360, n59361,
         n59362, n59363, n59364, n59365, n59366, n59369, n59370, n59372,
         n59373, n59374, n59375, n59376, n59377, n59378, n59379, n59381,
         n59382, n59383, n59384, n59387, n59388, n59389, n59390, n59391,
         n59392, n59393, n59394, n59395, n59396, n59397, n59398, n59399,
         n59400, n59402, n59403, n59404, n59406, n59407, n59408, n59409,
         n59412, n59415, n59416, n59417, n59418, n59419, n59420, n59421,
         n59422, n59424, n59425, n59426, n59427, n59428, n59429, n59431,
         n59432, n59435, n59437, n59439, n59440, n59442, n59443, n59444,
         n59445, n59446, n59447, n59449, n59451, n59452, n59453, n59454,
         n59455, n59458, n59460, n59461, n59462, n59463, n59464, n59465,
         n59467, n59468, n59469, n59470, n59471, n59472, n59473, n59474,
         n59475, n59476, n59477, n59479, n59481, n59482, n59483, n59485,
         n59486, n59487, n59488, n59490, n59491, n59492, n59493, n59495,
         n59496, n59497, n59499, n59501, n59505, n59506, n59507, n59508,
         n59510, n59514, n59515, n59516, n59517, n59518, n59521, n59522,
         n59523, n59528, n59530, n59531, n59532, n59533, n59534, n59536,
         n59537, n59538, n59539, n59541, n59542, n59543, n59544, n59545,
         n59546, n59547, n59550, n59551, n59552, n59553, n59554, n59555,
         n59557, n59558, n59559, n59560, n59561, n59562, n59563, n59565,
         n59566, n59567, n59568, n59569, n59570, n59571, n59572, n59574,
         n59575, n59576, n59577, n59581, n59582, n59583, n59585, n59586,
         n59587, n59588, n59589, n59590, n59591, n59593, n59594, n59597,
         n59599, n59601, n59602, n59603, n59604, n59607, n59608, n59609,
         n59610, n59611, n59613, n59614, n59615, n59616, n59617, n59618,
         n59619, n59620, n59621, n59622, n59625, n59626, n59627, n59628,
         n59629, n59630, n59631, n59632, n59633, n59634, n59637, n59638,
         n59639, n59640, n59641, n59642, n59644, n59645, n59646, n59647,
         n59648, n59649, n59650, n59651, n59652, n59655, n59657, n59658,
         n59660, n59661, n59662, n59663, n59664, n59665, n59667, n59668,
         n59669, n59670, n59671, n59672, n59673, n59674, n59675, n59676,
         n59678, n59679, n59680, n59681, n59682, n59684, n59685, n59686,
         n59687, n59688, n59689, n59690, n59691, n59692, n59694, n59695,
         n59696, n59697, n59698, n59699, n59700, n59701, n59703, n59705,
         n59706, n59707, n59708, n59709, n59710, n59711, n59713, n59714,
         n59715, n59716, n59717, n59718, n59719, n59720, n59721, n59722,
         n59723, n59724, n59728, n59730, n59731, n59732, n59733, n59734,
         n59735, n59736, n59737, n59739, n59741, n59744, n59746, n59747,
         n59749, n59750, n59751, n59752, n59753, n59754, n59755, n59758,
         n59759, n59760, n59763, n59764, n59765, n59767, n59769, n59770,
         n59771, n59772, n59773, n59775, n59776, n59777, n59779, n59780,
         n59781, n59782, n59783, n59785, n59786, n59787, n59788, n59789,
         n59790, n59791, n59792, n59794, n59795, n59797, n59798, n59799,
         n59801, n59802, n59803, n59804, n59805, n59806, n59808, n59809,
         n59810, n59811, n59812, n59813, n59815, n59817, n59818, n59820,
         n59821, n59822, n59823, n59824, n59825, n59826, n59827, n59828,
         n59829, n59831, n59832, n59833, n59834, n59835, n59836, n59838,
         n59841, n59842, n59843, n59844, n59845, n59847, n59848, n59849,
         n59851, n59852, n59853, n59854, n59855, n59856, n59858, n59859,
         n59860, n59861, n59862, n59863, n59866, n59867, n59868, n59871,
         n59872, n59873, n59874, n59875, n59876, n59877, n59878, n59879,
         n59880, n59881, n59882, n59883, n59884, n59885, n59887, n59888,
         n59889, n59890, n59891, n59892, n59893, n59894, n59895, n59896,
         n59898, n59899, n59900, n59903, n59904, n59905, n59907, n59909,
         n59910, n59911, n59912, n59913, n59914, n59915, n59916, n59918,
         n59920, n59922, n59923, n59924, n59925, n59926, n59927, n59928,
         n59929, n59930, n59931, n59932, n59933, n59934, n59935, n59936,
         n59937, n59938, n59939, n59940, n59941, n59942, n59943, n59944,
         n59945, n59946, n59947, n59948, n59949, n59950, n59951, n59952,
         n59954, n59956, n59957, n59958, n59959, n59961, n59962, n59963,
         n59964, n59965, n59966, n59967, n59968, n59969, n59970, n59972,
         n59973, n59974, n59975, n59976, n59977, n59979, n59980, n59981,
         n59982, n59983, n59984, n59985, n59987, n59988, n59989, n59990,
         n59991, n59992, n59993, n59994, n59998, n60000, n60001, n60002,
         n60003, n60004, n60005, n60006, n60008, n60009, n60010, n60011,
         n60012, n60013, n60014, n60018, n60019, n60020, n60021, n60022,
         n60023, n60024, n60026, n60028, n60030, n60031, n60032, n60033,
         n60034, n60037, n60038, n60039, n60041, n60042, n60043, n60045,
         n60046, n60049, n60050, n60052, n60054, n60055, n60056, n60058,
         n60059, n60062, n60063, n60064, n60065, n60066, n60069, n60070,
         n60071, n60072, n60073, n60074, n60075, n60076, n60077, n60078,
         n60079, n60081, n60082, n60083, n60084, n60085, n60086, n60087,
         n60088, n60091, n60092, n60093, n60094, n60095, n60097, n60099,
         n60100, n60101, n60102, n60103, n60104, n60105, n60106, n60107,
         n60108, n60109, n60110, n60111, n60112, n60113, n60114, n60115,
         n60116, n60118, n60119, n60121, n60122, n60123, n60124, n60125,
         n60126, n60127, n60128, n60129, n60130, n60131, n60132, n60133,
         n60134, n60135, n60138, n60139, n60140, n60141, n60142, n60143,
         n60144, n60145, n60146, n60147, n60148, n60149, n60151, n60152,
         n60153, n60154, n60155, n60156, n60157, n60159, n60161, n60162,
         n60163, n60164, n60165, n60166, n60167, n60168, n60169, n60170,
         n60171, n60172, n60173, n60174, n60175, n60176, n60179, n60180,
         n60181, n60183, n60185, n60186, n60187, n60188, n60189, n60191,
         n60194, n60195, n60196, n60198, n60199, n60200, n60201, n60202,
         n60203, n60204, n60206, n60207, n60209, n60210, n60212, n60213,
         n60214, n60215, n60216, n60218, n60219, n60220, n60221, n60222,
         n60223, n60224, n60225, n60226, n60227, n60228, n60229, n60230,
         n60232, n60233, n60234, n60236, n60237, n60238, n60239, n60240,
         n60241, n60242, n60243, n60245, n60247, n60248, n60249, n60250,
         n60251, n60252, n60256, n60257, n60258, n60259, n60261, n60262,
         n60264, n60265, n60267, n60268, n60270, n60272, n60274, n60275,
         n60276, n60278, n60279, n60280, n60282, n60283, n60284, n60285,
         n60287, n60289, n60290, n60291, n60292, n60293, n60294, n60295,
         n60297, n60298, n60300, n60301, n60302, n60303, n60305, n60306,
         n60308, n60309, n60310, n60311, n60312, n60313, n60314, n60315,
         n60316, n60318, n60319, n60321, n60323, n60324, n60325, n60326,
         n60327, n60328, n60329, n60333, n60334, n60335, n60336, n60337,
         n60338, n60339, n60342, n60343, n60344, n60345, n60347, n60348,
         n60349, n60350, n60351, n60353, n60355, n60356, n60358, n60360,
         n60361, n60362, n60363, n60364, n60365, n60366, n60367, n60368,
         n60370, n60372, n60373, n60374, n60375, n60376, n60377, n60378,
         n60380, n60381, n60382, n60383, n60384, n60386, n60387, n60388,
         n60390, n60391, n60392, n60393, n60394, n60395, n60397, n60398,
         n60399, n60400, n60401, n60404, n60405, n60407, n60408, n60409,
         n60410, n60411, n60413, n60415, n60416, n60417, n60419, n60420,
         n60421, n60422, n60423, n60425, n60426, n60428, n60429, n60430,
         n60431, n60432, n60433, n60434, n60435, n60437, n60439, n60440,
         n60441, n60444, n60447, n60448, n60449, n60450, n60451, n60452,
         n60453, n60455, n60456, n60457, n60458, n60459, n60461, n60462,
         n60464, n60465, n60466, n60467, n60469, n60470, n60471, n60472,
         n60473, n60474, n60475, n60476, n60479, n60480, n60482, n60483,
         n60484, n60485, n60486, n60487, n60488, n60489, n60490, n60492,
         n60493, n60494, n60495, n60496, n60497, n60498, n60499, n60500,
         n60501, n60502, n60503, n60504, n60505, n60507, n60508, n60509,
         n60510, n60511, n60513, n60514, n60515, n60516, n60517, n60518,
         n60519, n60520, n60522, n60523, n60524, n60525, n60526, n60527,
         n60528, n60529, n60530, n60531, n60532, n60533, n60534, n60537,
         n60538, n60539, n60540, n60541, n60542, n60543, n60544, n60545,
         n60546, n60547, n60548, n60549, n60550, n60551, n60552, n60553,
         n60554, n60555, n60556, n60557, n60559, n60560, n60561, n60562,
         n60563, n60564, n60565, n60567, n60568, n60570, n60571, n60572,
         n60573, n60574, n60575, n60576, n60577, n60578, n60579, n60580,
         n60581, n60582, n60583, n60584, n60585, n60587, n60590, n60591,
         n60592, n60593, n60594, n60595, n60597, n60599, n60600, n60601,
         n60602, n60603, n60604, n60606, n60608, n60609, n60610, n60612,
         n60614, n60615, n60616, n60617, n60619, n60620, n60621, n60622,
         n60624, n60625, n60626, n60627, n60628, n60629, n60630, n60631,
         n60632, n60633, n60634, n60635, n60636, n60637, n60639, n60641,
         n60642, n60643, n60644, n60645, n60647, n60648, n60649, n60650,
         n60651, n60652, n60653, n60654, n60655, n60656, n60657, n60659,
         n60661, n60662, n60663, n60665, n60666, n60667, n60668, n60669,
         n60670, n60672, n60674, n60675, n60676, n60677, n60681, n60682,
         n60683, n60684, n60685, n60686, n60687, n60688, n60690, n60691,
         n60692, n60693, n60694, n60695, n60696, n60697, n60699, n60700,
         n60701, n60702, n60706, n60707, n60708, n60709, n60710, n60711,
         n60713, n60714, n60715, n60716, n60717, n60718, n60719, n60720,
         n60721, n60722, n60723, n60724, n60725, n60726, n60727, n60728,
         n60730, n60731, n60732, n60734, n60735, n60736, n60737, n60738,
         n60740, n60741, n60742, n60743, n60744, n60746, n60749, n60750,
         n60751, n60752, n60753, n60754, n60755, n60756, n60757, n60758,
         n60759, n60760, n60761, n60762, n60763, n60764, n60765, n60766,
         n60767, n60768, n60770, n60771, n60772, n60774, n60776, n60777,
         n60778, n60779, n60780, n60781, n60782, n60783, n60784, n60786,
         n60788, n60789, n60792, n60793, n60794, n60795, n60796, n60797,
         n60798, n60799, n60801, n60803, n60804, n60805, n60807, n60808,
         n60809, n60810, n60811, n60812, n60813, n60814, n60815, n60816,
         n60817, n60818, n60819, n60820, n60821, n60822, n60823, n60824,
         n60825, n60826, n60828, n60829, n60830, n60831, n60832, n60833,
         n60835, n60836, n60837, n60838, n60839, n60840, n60841, n60842,
         n60843, n60844, n60845, n60846, n60848, n60849, n60850, n60851,
         n60853, n60854, n60855, n60856, n60857, n60858, n60859, n60860,
         n60861, n60862, n60863, n60865, n60866, n60867, n60868, n60869,
         n60870, n60871, n60872, n60874, n60875, n60876, n60877, n60878,
         n60879, n60880, n60881, n60882, n60883, n60884, n60885, n60886,
         n60887, n60888, n60889, n60890, n60891, n60892, n60893, n60894,
         n60895, n60897, n60898, n60899, n60900, n60901, n60902, n60903,
         n60904, n60906, n60908, n60909, n60910, n60911, n60912, n60913,
         n60914, n60915, n60916, n60918, n60919, n60921, n60922, n60923,
         n60925, n60926, n60927, n60928, n60929, n60930, n60931, n60932,
         n60934, n60935, n60937, n60939, n60940, n60941, n60942, n60943,
         n60945, n60946, n60947, n60948, n60949, n60950, n60951, n60952,
         n60953, n60954, n60955, n60956, n60957, n60958, n60959, n60960,
         n60961, n60962, n60963, n60964, n60966, n60967, n60968, n60969,
         n60970, n60971, n60973, n60974, n60975, n60977, n60979, n60980,
         n60981, n60982, n60983, n60984, n60985, n60987, n60988, n60989,
         n60990, n60992, n60993, n60994, n60996, n60997, n60998, n60999,
         n61000, n61001, n61004, n61005, n61006, n61007, n61008, n61009,
         n61010, n61011, n61012, n61013, n61014, n61016, n61017, n61018,
         n61020, n61021, n61022, n61023, n61025, n61026, n61027, n61028,
         n61030, n61032, n61033, n61034, n61035, n61037, n61039, n61041,
         n61042, n61043, n61044, n61045, n61046, n61047, n61048, n61049,
         n61050, n61052, n61053, n61054, n61055, n61057, n61058, n61061,
         n61064, n61065, n61066, n61067, n61069, n61070, n61071, n61072,
         n61074, n61075, n61076, n61077, n61078, n61079, n61081, n61082,
         n61083, n61086, n61087, n61088, n61089, n61090, n61091, n61092,
         n61094, n61095, n61096, n61099, n61100, n61101, n61102, n61103,
         n61104, n61105, n61106, n61107, n61108, n61109, n61110, n61111,
         n61112, n61115, n61116, n61117, n61119, n61120, n61121, n61122,
         n61123, n61124, n61125, n61126, n61127, n61128, n61129, n61130,
         n61131, n61132, n61133, n61134, n61135, n61136, n61137, n61138,
         n61139, n61140, n61142, n61143, n61144, n61145, n61146, n61147,
         n61149, n61150, n61151, n61152, n61153, n61155, n61156, n61157,
         n61158, n61159, n61160, n61162, n61164, n61165, n61166, n61167,
         n61168, n61169, n61170, n61171, n61173, n61174, n61175, n61176,
         n61177, n61178, n61179, n61180, n61181, n61182, n61183, n61184,
         n61186, n61187, n61191, n61192, n61193, n61194, n61195, n61196,
         n61197, n61198, n61202, n61203, n61204, n61205, n61207, n61208,
         n61209, n61210, n61211, n61212, n61213, n61215, n61216, n61218,
         n61219, n61220, n61221, n61222, n61223, n61225, n61226, n61228,
         n61229, n61231, n61232, n61233, n61234, n61235, n61236, n61237,
         n61238, n61239, n61240, n61241, n61242, n61243, n61244, n61246,
         n61247, n61248, n61249, n61250, n61251, n61252, n61253, n61255,
         n61256, n61257, n61258, n61260, n61261, n61262, n61263, n61264,
         n61265, n61267, n61270, n61272, n61273, n61277, n61278, n61279,
         n61280, n61281, n61282, n61283, n61284, n61285, n61286, n61287,
         n61288, n61289, n61290, n61291, n61292, n61293, n61294, n61295,
         n61297, n61298, n61299, n61300, n61304, n61305, n61306, n61307,
         n61308, n61309, n61310, n61311, n61312, n61313, n61314, n61315,
         n61316, n61317, n61318, n61319, n61320, n61321, n61324, n61325,
         n61326, n61327, n61330, n61331, n61332, n61333, n61334, n61335,
         n61337, n61338, n61340, n61341, n61343, n61344, n61346, n61347,
         n61348, n61349, n61350, n61352, n61354, n61355, n61356, n61358,
         n61359, n61360, n61361, n61362, n61363, n61364, n61365, n61366,
         n61368, n61371, n61372, n61373, n61374, n61375, n61376, n61380,
         n61382, n61383, n61384, n61385, n61386, n61387, n61388, n61389,
         n61390, n61391, n61392, n61394, n61395, n61397, n61398, n61399,
         n61400, n61401, n61402, n61403, n61405, n61407, n61409, n61410,
         n61411, n61412, n61413, n61414, n61415, n61416, n61417, n61418,
         n61419, n61420, n61421, n61422, n61423, n61424, n61426, n61429,
         n61432, n61433, n61434, n61435, n61436, n61438, n61439, n61440,
         n61441, n61442, n61443, n61444, n61445, n61446, n61447, n61449,
         n61450, n61452, n61455, n61457, n61458, n61461, n61462, n61463,
         n61464, n61465, n61467, n61468, n61469, n61470, n61472, n61473,
         n61474, n61475, n61476, n61477, n61478, n61479, n61483, n61484,
         n61487, n61488, n61489, n61490, n61491, n61492, n61494, n61496,
         n61497, n61498, n61499, n61500, n61501, n61502, n61503, n61506,
         n61507, n61508, n61509, n61510, n61511, n61512, n61513, n61516,
         n61517, n61518, n61519, n61520, n61521, n61522, n61523, n61524,
         n61525, n61526, n61527, n61528, n61529, n61530, n61531, n61532,
         n61533, n61534, n61535, n61536, n61537, n61538, n61539, n61540,
         n61541, n61543, n61544, n61545, n61546, n61547, n61548, n61549,
         n61550, n61551, n61552, n61553, n61554, n61555, n61556, n61557,
         n61558, n61559, n61560, n61561, n61563, n61564, n61565, n61566,
         n61567, n61569, n61571, n61572, n61573, n61574, n61575, n61576,
         n61577, n61578, n61579, n61581, n61582, n61583, n61584, n61590,
         n61591, n61592, n61593, n61594, n61595, n61596, n61597, n61598,
         n61599, n61601, n61602, n61603, n61604, n61605, n61606, n61608,
         n61609, n61610, n61611, n61612, n61613, n61614, n61617, n61618,
         n61619, n61620, n61622, n61623, n61624, n61625, n61626, n61627,
         n61628, n61629, n61630, n61631, n61632, n61633, n61634, n61636,
         n61638, n61640, n61641, n61642, n61643, n61644, n61646, n61647,
         n61648, n61649, n61650, n61651, n61652, n61653, n61654, n61655,
         n61656, n61657, n61658, n61659, n61660, n61661, n61662, n61663,
         n61664, n61665, n61666, n61667, n61668, n61669, n61670, n61671,
         n61672, n61673, n61674, n61675, n61676, n61677, n61678, n61679,
         n61680, n61681, n61682, n61683, n61684, n61685, n61686, n61687,
         n61688, n61690, n61691, n61693, n61694, n61695, n61696, n61697,
         n61698, n61699, n61700, n61701, n61702, n61703, n61704, n61705,
         n61706, n61707, n61708, n61709, n61710, n61711, n61712, n61713,
         n61714, n61715, n61716, n61717, n61718, n61719, n61720, n61721,
         n61722, n61723, n61724, n61725, n61726, n61727, n61728, n61729,
         n61730, n61731, n61732, n61733, n61734, n61735, n61736, n61737,
         n61738, n61739, n61740, n61741, n61742, n61743, n61744, n61745,
         n61746, n61747, n61748, n61749, n61750, n61751, n61752, n61753,
         n61754, n61755, n61756, n61757, n61758, n61759, n61760, n61761,
         n61762, n61763, n61764, n61765, n61766, n61767, n61768, n61769,
         n61770, n61771, n61772, n61773, n61774, n61775, n61776, n61777,
         n61778, n61779, n61780, n61781, n61782, n61783, n61784, n61785,
         n61786, n61787, n61788, n61789, n61790, n61791, n61792, n61793,
         n61794, n61795, n61796, n61797, n61798, n61799, n61800, n61801,
         n61802, n61803, n61804, n61805, n61806, n61807, n61808, n61809,
         n61810, n61811, n61812, n61813, n61814, n61815, n61816, n61817,
         n61818, n61819, n61820, n61821, n61822, n61823, n61824, n61825,
         n61826, n61827, n61828, n61829, n61830, n61831, n61832, n61833,
         n61834, n61835, n61836, n61837, n61838, n61839, n61840, n61841,
         n61842, n61843, n61844, n61845, n61846, n61847, n61848, n61849,
         n61850, n61851, n61852, n61853, n61854, n61855, n61856, n61857,
         n61858, n61859, n61860, n61861, n61862, n61863, n61864, n61865,
         n61866, n61867, n61868, n61869, n61870, n61871, n61872, n61873,
         n61874, n61875, n61876, n61877, n61878, n61879, n61880, n61881,
         n61882, n61883, n61884, n61885, n61886, n61887, n61888, n61889,
         n61890, n61891, n61892, n61893, n61894, n61895, n61896, n61897,
         n61898, n61899, n61900, n61901, n61902, n61903, n61904, n61905,
         n61906, n61907, n61908, n61909, n61910, n61911, n61912, n61913,
         n61914, n61915, n61916, n61917, n61918, n61919, n61920, n61921,
         n61922, n61923, n61924, n61925, n61926, n61927, n61928, n61929,
         n61930, n61931, n61932, n61933, n61934, n61935, n61936, n61937,
         n61938, n61939, n61940, n61941, n61942, n61943, n61944, n61945,
         n61946, n61947, n61948, n61949, n61950, n61951, n61952, n61953,
         n61954, n61955, n61956, n61957, n61958, n61959, n61960, n61961,
         n61962, n61963, n61964, n61965, n61966, n61967, n61968, n61969,
         n61970, n61971, n61972, n61973, n61974, n61975, n61976, n61977,
         n61978, n61979, n61980, n61981, n61982, n61983, n61984, n61985,
         n61986, n61987, n61988, n61989, n61990, n61991, n61992, n61993,
         n61994, n61995, n61996, n61997, n61998, n61999, n62000, n62001,
         n62002, n62003, n62004, n62005, n62006, n62007, n62008, n62009,
         n62010, n62011, n62012, n62013, n62014, n62015, n62016, n62017,
         n62018, n62019, n62020, n62021, n62022, n62023, n62024, n62025,
         n62026, n62027, n62028, n62029, n62030, n62031, n62032, n62033,
         n62034, n62035, n62036, n62037, n62038, n62039, n62040, n62041,
         n62042, n62043, n62044, n62045, n62046, n62047, n62048, n62049,
         n62050, n62051, n62052, n62053, n62054, n62055, n62056, n62057,
         n62058, n62059, n62060, n62061, n62062, n62063, n62064, n62065,
         n62066, n62067, n62068, n62069, n62070, n62071, n62072, n62073,
         n62074, n62075, n62076, n62077, n62078, n62079, n62080, n62081,
         n62082, n62083, n62084, n62085, n62086, n62087, n62088, n62089,
         n62090, n62091, n62092, n62093, n62094, n62095, n62096, n62097,
         n62098, n62099, n62100, n62101, n62102, n62103, n62104, n62105,
         n62106, n62107, n62108, n62109, n62110, n62111, n62112, n62113,
         n62114, n62115, n62116, n62117, n62118, n62119, n62120, n62121,
         n62122, n62123, n62124, n62125, n62126, n62127, n62128, n62129,
         n62130, n62131, n62132, n62133, n62134, n62135, n62136, n62137,
         n62138, n62139, n62140, n62141, n62142, n62143, n62144, n62145,
         n62146, n62147, n62148, n62149, n62150, n62151, n62152, n62153,
         n62154, n62155, n62156, n62157, n62158, n62159, n62160, n62161,
         n62162, n62163, n62164, n62165, n62166, n62167, n62168, n62169,
         n62170, n62171, n62172, n62173, n62174, n62175, n62176, n62177,
         n62178, n62179, n62180, n62181, n62183, n62184, n62185, n62186,
         n62187, n62188, n62189, n62190, n62191, n62192, n62193, n62194,
         n62195, n62196, n62197, n62198, n62199, n62200, n62201, n62202,
         n62203, n62204, n62205, n62206, n62207, n62208, n62209, n62210,
         n62211, n62212, n62213, n62214, n62215, n62216, n62217, n62218,
         n62219, n62220, n62221, n62222, n62223, n62224, n62225, n62226,
         n62227, n62228, n62229, n62230, n62231, n62232, n62233, n62234,
         n62235, n62236, n62237, n62238, n62239, n62240, n62241, n62242,
         n62243, n62244, n62245, n62246, n62247, n62248, n62249, n62250,
         n62251, n62252, n62253, n62254, n62255, n62256, n62257, n62258,
         n62259, n62260, n62261, n62262, n62263, n62264, n62265, n62266,
         n62267, n62268, n62269, n62270, n62271, n62272, n62273, n62274,
         n62275, n62276, n62277, n62278, n62279, n62280, n62281, n62282,
         n62283, n62284, n62285, n62286, n62287, n62288, n62289, n62290,
         n62291, n62292, n62293, n62294, n62295, n62296, n62297, n62298,
         n62299, n62300, n62301, n62302, n62303, n62304, n62305, n62306,
         n62307, n62308, n62309, n62310, n62311, n62312, n62313, n62314,
         n62315, n62316, n62317, n62318, n62319, n62320, n62321, n62322,
         n62323, n62324, n62325, n62326, n62327, n62328, n62329, n62330,
         n62331, n62332, n62333, n62334, n62335, n62336, n62337, n62338,
         n62339, n62340, n62341, n62342, n62343, n62344, n62345, n62346,
         n62347, n62348, n62349, n62350, n62351, n62352, n62353, n62354,
         n62355, n62356, n62357, n62358, n62359, n62360, n62361, n62362,
         n62363, n62364, n62365, n62366, n62367, n62368, n62369, n62370,
         n62371, n62372, n62373, n62374, n62375, n62376, n62377, n62378,
         n62379, n62380, n62381, n62382, n62383, n62384, n62385, n62386,
         n62387, n62388, n62389, n62390, n62391, n62392, n62393, n62394,
         n62395, n62396, n62398, n62399, n62400, n62401, n62402, n62403,
         n62404, n62405, n62406, n62407, n62408, n62409, n62410, n62411,
         n62412, n62413, n62414, n62415, n62416, n62417, n62418, n62419,
         n62420, n62421, n62422, n62423, n62424, n62425, n62426, n62427,
         n62428, n62429, n62430, n62431, n62432, n62433, n62434, n62435,
         n62436, n62437, n62438, n62439, n62440, n62441, n62442, n62443,
         n62444, n62445, n62446, n62447, n62448, n62449, n62450, n62451,
         n62452, n62455, n62456, n62457, n62458, n62459, n62460, n62461,
         n62462, n62463, n62464, n62465, n62466, n62467, n62468, n62469,
         n62470, n62471, n62472, n62473, n62474, n62475, n62476, n62477,
         n62479, n62480, n62481, n62482, n62483, n62484, n62485, n62486,
         n62487, n62488, n62489, n62490, n62491, n62492, n62493, n62494,
         n62495, n62496, n62497, n62498, n62499, n62500, n62501, n62502,
         n62503, n62504, n62505, n62506, n62507, n62508, n62509, n62510,
         n62511, n62512, n62513, n62514, n62515, n62516, n62517, n62518,
         n62519, n62520, n62521, n62522, n62523, n62524, n62525, n62526,
         n62527, n62528, n62529, n62530, n62531, n62532, n62533, n62534,
         n62535, n62536, n62537, n62538, n62539, n62540, n62541, n62542,
         n62543, n62544, n62545, n62546, n62547, n62548, n62549, n62550,
         n62551, n62552, n62553, n62554, n62555, n62556, n62557, n62558,
         n62559, n62560, n62561, n62562, n62563, n62564, n62565, n62566,
         n62567, n62568, n62569, n62570, n62571, n62572, n62573, n62574,
         n62575, n62576, n62577, n62578, n62579, n62580, n62581, n62582,
         n62583, n62584, n62585, n62586, n62587, n62588, n62589, n62590,
         n62591, n62592, n62593, n62594, n62595, n62596, n62597, n62598,
         n62599, n62600, n62601, n62602, n62603, n62604, n62605, n62606,
         n62607, n62608, n62609, n62610, n62611, n62612, n62613, n62614,
         n62615, n62616, n62617, n62618, n62619, n62620, n62621, n62622,
         n62623, n62624, n62625, n62626, n62627, n62628, n62629, n62630,
         n62631, n62632, n62633, n62634, n62635, n62636, n62637, n62638,
         n62639, n62640, n62641, n62642, n62643, n62644, n62645, n62646,
         n62647, n62648, n62649, n62650, n62651, n62652, n62653, n62654,
         n62655, n62656, n62657, n62658, n62659, n62660, n62661, n62662,
         n62663, n62664, n62665, n62666, n62667, n62668, n62669, n62670,
         n62671, n62672, n62673, n62674, n62675, n62676, n62677, n62678,
         n62679, n62680, n62681, n62682, n62683, n62684, n62685, n62686,
         n62687, n62688, n62689, n62690, n62691, n62692, n62693, n62694,
         n62695, n62696, n62697, n62698, n62699, n62700, n62701, n62702,
         n62703, n62704, n62705, n62706, n62707, n62708, n62709, n62710,
         n62711, n62712, n62713, n62714, n62715, n62716, n62717, n62718,
         n62719, n62720, n62721, n62722, n62723, n62724, n62725, n62726,
         n62727, n62729, n62730, n62731, n62732, n62733, n62734, n62735,
         n62736, n62737, n62738, n62739, n62740, n62741, n62742, n62743,
         n62744, n62745, n62746, n62747, n62748, n62749, n62750, n62751,
         n62752, n62753, n62754, n62755, n62756, n62757, n62758, n62759,
         n62760, n62761, n62762, n62763, n62764, n62765, n62766, n62767,
         n62768, n62769, n62770, n62771, n62772, n62773, n62774, n62775,
         n62776, n62777, n62778, n62779, n62780, n62781, n62782, n62783,
         n62784, n62785, n62786, n62787, n62788, n62789, n62790, n62791,
         n62792, n62793, n62794, n62795, n62796, n62797, n62798, n62799,
         n62800, n62801, n62802, n62803, n62804, n62805, n62806, n62807,
         n62808, n62809, n62810, n62811, n62812, n62813, n62814, n62815,
         n62817, n62818, n62819, n62820, n62821, n62822, n62823, n62824,
         n62825, n62826, n62827, n62828, n62829, n62830, n62831, n62832,
         n62833, n62834, n62835, n62836, n62837, n62838, n62839, n62840,
         n62841, n62842, n62843, n62844, n62845, n62846, n62847, n62848,
         n62849, n62850, n62851, n62852, n62853, n62854, n62855, n62856,
         n62857, n62858, n62859, n62860, n62861, n62862, n62863, n62864,
         n62865, n62866, n62867, n62868, n62869, n62870, n62871, n62872,
         n62873, n62874, n62875, n62876, n62877, n62878, n62879, n62880,
         n62881, n62882, n62883, n62884, n62885, n62886, n62887, n62888,
         n62889, n62890, n62891, n62892, n62893, n62894, n62895, n62896,
         n62897, n62898, n62899, n62900, n62901, n62902, n62903, n62904,
         n62905, n62906, n62907, n62908, n62909, n62910, n62911, n62912,
         n62913, n62914, n62915, n62916, n62917, n62918, n62919, n62920,
         n62921, n62922, n62923, n62924, n62925, n62926, n62927, n62928,
         n62929, n62930, n62931, n62932, n62933, n62934, n62935, n62936,
         n62937, n62938, n62939, n62940, n62941, n62942, n62943, n62944,
         n62945, n62946, n62947, n62948, n62949, n62950, n62951, n62952,
         n62953, n62954, n62955, n62956, n62957, n62958, n62959, n62960,
         n62961, n62962, n62963, n62964, n62965, n62966, n62967, n62968,
         n62969, n62970, n62971, n62972, n62973, n62974, n62975, n62976,
         n62977, n62978, n62979, n62980, n62981, n62982, n62983, n62984,
         n62985, n62986, n62987, n62988, n62989, n62990, n62991, n62992,
         n62993, n62994, n62995, n62996, n62997, n62998, n62999, n63000,
         n63001, n63002, n63003, n63004, n63005, n63006, n63007, n63008,
         n63009, n63010, n63011, n63012, n63013, n63014, n63015, n63016,
         n63017, n63018, n63019, n63020, n63021, n63022, n63023, n63024,
         n63025, n63026, n63027, n63028, n63029, n63030, n63031, n63032,
         n63033, n63034, n63035, n63036, n63037, n63038, n63039, n63040,
         n63041, n63042, n63043, n63044, n63045, n63046, n63047, n63048,
         n63049, n63050, n63051, n63052, n63053, n63054, n63055, n63056,
         n63057, n63058, n63059, n63060, n63061, n63062, n63063, n63064,
         n63065, n63066, n63067, n63068, n63069, n63070, n63071, n63072,
         n63073, n63074, n63075, n63076, n63077, n63078, n63079, n63080,
         n63081, n63082, n63083, n63084, n63085, n63086, n63087, n63088,
         n63089, n63090, n63091, n63092, n63093, n63094, n63095, n63096,
         n63097, n63098, n63099, n63100, n63101, n63102, n63103, n63104,
         n63105, n63106, n63107, n63108, n63109, n63110, n63111, n63112,
         n63113, n63114, n63115, n63116, n63117, n63118, n63119, n63120,
         n63121, n63122, n63123, n63124, n63125, n63126, n63127, n63128,
         n63129, n63130, n63131, n63132, n63133, n63134, n63135, n63136,
         n63137, n63138, n63139, n63140, n63141, n63142, n63144, n63145,
         n63146, n63147, n63148, n63149, n63150, n63151, n63152, n63153,
         n63154, n63155, n63156, n63157, n63158, n63159, n63160, n63161,
         n63162, n63163, n63164, n63165, n63166, n63167, n63168, n63169,
         n63170, n63171, n63172, n63173, n63174, n63175, n63176, n63177,
         n63178, n63179, n63180, n63181, n63182, n63183, n63184, n63185,
         n63186, n63187, n63188, n63189, n63190, n63191, n63192, n63193,
         n63194, n63195, n63196, n63197, n63198, n63199, n63200, n63201,
         n63202, n63203, n63204, n63205, n63206, n63207, n63208, n63209,
         n63210, n63211, n63212, n63213, n63214, n63215, n63216, n63217,
         n63218, n63219, n63220, n63221, n63222, n63223, n63224, n63225,
         n63226, n63227, n63228, n63229, n63230, n63231, n63232, n63233,
         n63234, n63235, n63236, n63237, n63238, n63239, n63240, n63241,
         n63242, n63243, n63244, n63245, n63246, n63247, n63248, n63249,
         n63250, n63251, n63252, n63253, n63254, n63255, n63256, n63257,
         n63258, n63259, n63260, n63261, n63262, n63263, n63264, n63265,
         n63266, n63267, n63268, n63269, n63270, n63271, n63272, n63273,
         n63274, n63275, n63276, n63277, n63278, n63279, n63280, n63281,
         n63282, n63283, n63284, n63285, n63286, n63287, n63288, n63289,
         n63290, n63291, n63292, n63293, n63294, n63295, n63296, n63297,
         n63298, n63299, n63300, n63301, n63302, n63303, n63304, n63305,
         n63306, n63307, n63308, n63309, n63310, n63311, n63312, n63313,
         n63314, n63315, n63316, n63317, n63318, n63319, n63320, n63321,
         n63322, n63323, n63324, n63325, n63326, n63327, n63328, n63329,
         n63330, n63331, n63332, n63333, n63334, n63335, n63336, n63337,
         n63338, n63339, n63340, n63341, n63342, n63343, n63344, n63345,
         n63346, n63347, n63348, n63349, n63350, n63351, n63352, n63353,
         n63354, n63355, n63356, n63357, n63358, n63359, n63360, n63361,
         n63362, n63363, n63364, n63365, n63366, n63367, n63368, n63369,
         n63370, n63371, n63372, n63373, n63374, n63375, n63376, n63377,
         n63378, n63379, n63380, n63381, n63382, n63383, n63384, n63385,
         n63386, n63387, n63388, n63389, n63390, n63391, n63392, n63393,
         n63394, n63395, n63396, n63397, n63398, n63399, n63400, n63401,
         n63402, n63403, n63404, n63405, n63406, n63407, n63409, n63410,
         n63411, n63412, n63413, n63414, n63415, n63416, n63417, n63418,
         n63419, n63420, n63421, n63422, n63423, n63424, n63425, n63426,
         n63427, n63428, n63429, n63430, n63431, n63432, n63433, n63435,
         n63436, n63437, n63438, n63439, n63440, n63441, n63442, n63443,
         n63444, n63445, n63446, n63447, n63448, n63449, n63450, n63451,
         n63452, n63453, n63454, n63455, n63456, n63457, n63458, n63459,
         n63460, n63461, n63462, n63463, n63464, n63465, n63466, n63467,
         n63468, n63469, n63470, n63471, n63472, n63473, n63474, n63475,
         n63476, n63477, n63478, n63479, n63480, n63481, n63482, n63483,
         n63484, n63485, n63486, n63487, n63488, n63489, n63490, n63491,
         n63492, n63493, n63494, n63495, n63496, n63497, n63498, n63499,
         n63500, n63501, n63502, n63503, n63504, n63505, n63506, n63507,
         n63508, n63509, n63510, n63511, n63512, n63513, n63514, n63515,
         n63516, n63517, n63518, n63519, n63520, n63521, n63522, n63523,
         n63524, n63525, n63526, n63527, n63528, n63529, n63530, n63531,
         n63532, n63533, n63534, n63535, n63536, n63537, n63538, n63539,
         n63540, n63541, n63542, n63543, n63544, n63545, n63546, n63547,
         n63548, n63549, n63550, n63551, n63552, n63553, n63554, n63555,
         n63556, n63557, n63558, n63559, n63560, n63562, n63563, n63564,
         n63565, n63566, n63567, n63568, n63569, n63570, n63571, n63572,
         n63573, n63574, n63575, n63576, n63577, n63578, n63579, n63580,
         n63581, n63582, n63583, n63584, n63585, n63586, n63587, n63588,
         n63589, n63590, n63591, n63592, n63593, n63594, n63595, n63596,
         n63597, n63598, n63599, n63600, n63601, n63602, n63603, n63604,
         n63605, n63606, n63607, n63608, n63609, n63610, n63611, n63612,
         n63613, n63614, n63615, n63616, n63617, n63618, n63619, n63620,
         n63621, n63622, n63623, n63624, n63625, n63626, n63627, n63628,
         n63629, n63630, n63631, n63632, n63633, n63634, n63635, n63636,
         n63637, n63638, n63639, n63640, n63641, n63642, n63643, n63644,
         n63645, n63646, n63647, n63648, n63649, n63650, n63651, n63652,
         n63653, n63654, n63655, n63656, n63657, n63658, n63659, n63660,
         n63661, n63662, n63663, n63664, n63665, n63666, n63667, n63668,
         n63669, n63670, n63671, n63672, n63673, n63674, n63675, n63676,
         n63677, n63678, n63679, n63680, n63681, n63682, n63683, n63684,
         n63685, n63686, n63687, n63688, n63689, n63690, n63691, n63692,
         n63693, n63694, n63695, n63696, n63697, n63698, n63699, n63700,
         n63701, n63702, n63703, n63704, n63705, n63706, n63707, n63708,
         n63709, n63710, n63711, n63712, n63713, n63714, n63715, n63716,
         n63717, n63718, n63719, n63720, n63721, n63722, n63723, n63724,
         n63725, n63726, n63727, n63728, n63729, n63730, n63731, n63732,
         n63733, n63734, n63735, n63736, n63737, n63738, n63739, n63740,
         n63741, n63742, n63743, n63744, n63745, n63746, n63747, n63748,
         n63749, n63750, n63751, n63752, n63753, n63754, n63755, n63756,
         n63757, n63758, n63759, n63760, n63761, n63762, n63763, n63764,
         n63765, n63766, n63767, n63768, n63769, n63770, n63771, n63772,
         n63773, n63774, n63775, n63776, n63777, n63778, n63779, n63780,
         n63781, n63782, n63783, n63784, n63785, n63786, n63787, n63788,
         n63789, n63790, n63791, n63792, n63793, n63794, n63795, n63796,
         n63797, n63798, n63799, n63800, n63801, n63802, n63803, n63804,
         n63805, n63806, n63807, n63808, n63809, n63810, n63811, n63812,
         n63813, n63814, n63815, n63816, n63817, n63818, n63819, n63820,
         n63821, n63822, n63823, n63824, n63825, n63826, n63827, n63828,
         n63829, n63830, n63831, n63832, n63833, n63834, n63835, n63836,
         n63837, n63838, n63839, n63840, n63841, n63842, n63843, n63844,
         n63845, n63846, n63848, n63849, n63850, n63851, n63852, n63853,
         n63854, n63855, n63856, n63857, n63858, n63859, n63860, n63861,
         n63862, n63863, n63864, n63865, n63866, n63867, n63868, n63869,
         n63870, n63871, n63872, n63873, n63874, n63875, n63876, n63877,
         n63878, n63879, n63880, n63881, n63882, n63883, n63884, n63885,
         n63886, n63887, n63888, n63889, n63890, n63891, n63892, n63893,
         n63894, n63895, n63896, n63897, n63898, n63899, n63900, n63901,
         n63902, n63903, n63904, n63905, n63906, n63907, n63908, n63909,
         n63910, n63911, n63912, n63913, n63914, n63915, n63916, n63917,
         n63918, n63919, n63920, n63921, n63922, n63923, n63924, n63925,
         n63926, n63927, n63928, n63929, n63930, n63931, n63932, n63933,
         n63934, n63935, n63936, n63937, n63938, n63939, n63940, n63941,
         n63942, n63943, n63944, n63945, n63946, n63947, n63948, n63949,
         n63950, n63951, n63952, n63953, n63954, n63955, n63956, n63957,
         n63958, n63959, n63960, n63961, n63962, n63963, n63964, n63965,
         n63966, n63967, n63968, n63969, n63970, n63971, n63972, n63973,
         n63974, n63975, n63976, n63977, n63978, n63979, n63980, n63981,
         n63982, n63983, n63984, n63985, n63986, n63987, n63988, n63989,
         n63990, n63991, n63992, n63993, n63994, n63995, n63996, n63997,
         n63998, n63999, n64000, n64001, n64002, n64003, n64004, n64005,
         n64006, n64007, n64008, n64009, n64010, n64011, n64012, n64013,
         n64014, n64015, n64016, n64017, n64018, n64019, n64020, n64021,
         n64022, n64023, n64024, n64025, n64026, n64027, n64028, n64029,
         n64030, n64031, n64032, n64033, n64034, n64035, n64036, n64037,
         n64038, n64039, n64040, n64041, n64042, n64043, n64044, n64045,
         n64046, n64047, n64048, n64049, n64050, n64051, n64052, n64053,
         n64054, n64055, n64056, n64057, n64058, n64059, n64060, n64061,
         n64062, n64063, n64064, n64065, n64066, n64067, n64068, n64069,
         n64070, n64071, n64072, n64073, n64074, n64075, n64076, n64077,
         n64078, n64079, n64080, n64081, n64082, n64083, n64084, n64085,
         n64086, n64087, n64088, n64089, n64090, n64091, n64092, n64093,
         n64094, n64095, n64096, n64097, n64098, n64099, n64100, n64101,
         n64102, n64103, n64104, n64105, n64106, n64107, n64108, n64109,
         n64110, n64111, n64112, n64113, n64114, n64115, n64116, n64117,
         n64118, n64119, n64120, n64121, n64122, n64123, n64124, n64125,
         n64126, n64127, n64128, n64129, n64130, n64131, n64132, n64133,
         n64134, n64135, n64136, n64137, n64138, n64139, n64140, n64141,
         n64142, n64143, n64144, n64145, n64146, n64147, n64148, n64149,
         n64150, n64151, n64152, n64153, n64154, n64155, n64156, n64157,
         n64158, n64159, n64160, n64161, n64162, n64163, n64164, n64165,
         n64166, n64167, n64168, n64169, n64170, n64171, n64172, n64173,
         n64174, n64175, n64176, n64177, n64178, n64179, n64180, n64181,
         n64182, n64183, n64184, n64185, n64186, n64187, n64188, n64189,
         n64190, n64191, n64192, n64193, n64194, n64195, n64196, n64197,
         n64198, n64199, n64200, n64201, n64202, n64203, n64204, n64205,
         n64206, n64207, n64208, n64209, n64210, n64211, n64212, n64213,
         n64214, n64215, n64216, n64217, n64218, n64219, n64220, n64221,
         n64222, n64223, n64224, n64225, n64226, n64227, n64228, n64229,
         n64230, n64231, n64232, n64233, n64234, n64235, n64236, n64237,
         n64238, n64239, n64240, n64241, n64242, n64243, n64244, n64245,
         n64246, n64247, n64248, n64249, n64250, n64251, n64252, n64253,
         n64254, n64255, n64256, n64257, n64258, n64259, n64260, n64261,
         n64262, n64263, n64264, n64265, n64266, n64267, n64268, n64269,
         n64270, n64271, n64272, n64273, n64274, n64275, n64276, n64277,
         n64278, n64279, n64280, n64281, n64282, n64283, n64284, n64285,
         n64286, n64287, n64288, n64289, n64290, n64291, n64292, n64293,
         n64294, n64295, n64296, n64297, n64298, n64299, n64300, n64301,
         n64302, n64303, n64304, n64305, n64306, n64307, n64308, n64309,
         n64310, n64311, n64312, n64313, n64314, n64315, n64316, n64317,
         n64318, n64319, n64320, n64321, n64322, n64323, n64324, n64325,
         n64326, n64327, n64328, n64329, n64330, n64332, n64333, n64334,
         n64335, n64336, n64337, n64338, n64339, n64340, n64341, n64342,
         n64343, n64344, n64345, n64346, n64347, n64348, n64349, n64350,
         n64351, n64352, n64353, n64354, n64355, n64356, n64357, n64358,
         n64359, n64360, n64361, n64362, n64363, n64364, n64365, n64366,
         n64367, n64368, n64369, n64370, n64371, n64372, n64373, n64374,
         n64375, n64376, n64377, n64378, n64379, n64380, n64381, n64382,
         n64383, n64384, n64385, n64386, n64387, n64388, n64389, n64390,
         n64391, n64392, n64393, n64394, n64395, n64396, n64397, n64398,
         n64399, n64400, n64401, n64402, n64403, n64404, n64405, n64406,
         n64407, n64408, n64409, n64410, n64411, n64412, n64413, n64414,
         n64415, n64416, n64417, n64418, n64419, n64420, n64421, n64422,
         n64423, n64424, n64425, n64426, n64427, n64428, n64429, n64430,
         n64431, n64432, n64433, n64434, n64435, n64436, n64437, n64438,
         n64439, n64440, n64441, n64442, n64443, n64444, n64445, n64446,
         n64447, n64448, n64449, n64450, n64451, n64452, n64453, n64454,
         n64455, n64456, n64457, n64458, n64459, n64460, n64461, n64462,
         n64463, n64464, n64465, n64466, n64468, n64469, n64470, n64471,
         n64472, n64473, n64474, n64475, n64476, n64477, n64478, n64479,
         n64480, n64481, n64482, n64483, n64484, n64485, n64486, n64487,
         n64488, n64489, n64490, n64491, n64492, n64493, n64494, n64495,
         n64496, n64497, n64498, n64499, n64500, n64501, n64502, n64503,
         n64504, n64505, n64506, n64507, n64508, n64509, n64510, n64511,
         n64512, n64513, n64514, n64515, n64516, n64517, n64518, n64519,
         n64520, n64521, n64522, n64523, n64524, n64525, n64526, n64527,
         n64528, n64529, n64530, n64531, n64532, n64533, n64534, n64535,
         n64536, n64537, n64538, n64539, n64540, n64541, n64542, n64543,
         n64544, n64545, n64546, n64547, n64548, n64549, n64550, n64551,
         n64552, n64553, n64554, n64555, n64556, n64557, n64558, n64559,
         n64560, n64561, n64562, n64563, n64564, n64565, n64566, n64567,
         n64568, n64569, n64570, n64571, n64572, n64573, n64574, n64575,
         n64576, n64577, n64578, n64579, n64580, n64581, n64582, n64583,
         n64584, n64585, n64586, n64587, n64588, n64589, n64590, n64591,
         n64592, n64593, n64594, n64595, n64596, n64597, n64598, n64599,
         n64600, n64601, n64602, n64603, n64604, n64605, n64606, n64607,
         n64608, n64609, n64610, n64611, n64612, n64613, n64614, n64615,
         n64616, n64617, n64618, n64619, n64620, n64621, n64622, n64623,
         n64624, n64625, n64626, n64627, n64628, n64629, n64630, n64631,
         n64632, n64634, n64635, n64636, n64637, n64638, n64639, n64640,
         n64641, n64642, n64643, n64644, n64645, n64646, n64647, n64649,
         n64650, n64651, n64652, n64653, n64654, n64655, n64656, n64657,
         n64658, n64659, n64660, n64661, n64662, n64663, n64664, n64665,
         n64666, n64667, n64668, n64669, n64670, n64671, n64672, n64673,
         n64674, n64675, n64676, n64677, n64678, n64679, n64680, n64681,
         n64682, n64683, n64684, n64685, n64686, n64687, n64688, n64689,
         n64690, n64691, n64692, n64693, n64694, n64695, n64696, n64697,
         n64698, n64699, n64700, n64701, n64702, n64703, n64704, n64705,
         n64706, n64707, n64708, n64709, n64710, n64711, n64712, n64713,
         n64714, n64715, n64716, n64717, n64718, n64719, n64720, n64721,
         n64722, n64723, n64724, n64725, n64726, n64727, n64728, n64729,
         n64730, n64731, n64732, n64733, n64734, n64735, n64736, n64737,
         n64738, n64739, n64740, n64741, n64742, n64743, n64744, n64745,
         n64746, n64747, n64748, n64749, n64750, n64751, n64752, n64753,
         n64754, n64755, n64756, n64757, n64758, n64759, n64760, n64761,
         n64762, n64763, n64764, n64765, n64766, n64767, n64768, n64769,
         n64770, n64771, n64772, n64773, n64774, n64775, n64776, n64777,
         n64778, n64779, n64780, n64781, n64782, n64783, n64784, n64785,
         n64786, n64787, n64788, n64789, n64790, n64791, n64792, n64793,
         n64794, n64795, n64796, n64797, n64798, n64799, n64800, n64801,
         n64802, n64803, n64804, n64805, n64806, n64807, n64808, n64809,
         n64810, n64811, n64812, n64813, n64814, n64815, n64816, n64817,
         n64818, n64819, n64820, n64821, n64822, n64823, n64824, n64825,
         n64826, n64827, n64828, n64829, n64830, n64831, n64832, n64833,
         n64834, n64835, n64836, n64837, n64838, n64839, n64840, n64841,
         n64842, n64843, n64844, n64845, n64846, n64847, n64848, n64849,
         n64850, n64851, n64852, n64853, n64854, n64855, n64856, n64857,
         n64858, n64859, n64860, n64861, n64862, n64863, n64864, n64865,
         n64867, n64868, n64869, n64870, n64871, n64872, n64873, n64874,
         n64875, n64876, n64877, n64878, n64879, n64880, n64881, n64882,
         n64883, n64884, n64885, n64886, n64887, n64888, n64889, n64890,
         n64891, n64892, n64893, n64894, n64895, n64896, n64897, n64898,
         n64899, n64900, n64901, n64902, n64903, n64904, n64905, n64906,
         n64907, n64908, n64909, n64910, n64911, n64912, n64913, n64914,
         n64915, n64916, n64917, n64918, n64919, n64920, n64921, n64922,
         n64923, n64924, n64925, n64926, n64927, n64928, n64929, n64930,
         n64931, n64932, n64933, n64934, n64935, n64936, n64937, n64938,
         n64939, n64940, n64941, n64942, n64943, n64944, n64945, n64946,
         n64947, n64948, n64949, n64950, n64951, n64952, n64953, n64954,
         n64955, n64956, n64957, n64958, n64959, n64960, n64961, n64962,
         n64963, n64964, n64965, n64966, n64967, n64968, n64969, n64970,
         n64971, n64972, n64973, n64974, n64975, n64976, n64977, n64978,
         n64979, n64980, n64981, n64982, n64983, n64984, n64985, n64986,
         n64987, n64988, n64989, n64990, n64991, n64992, n64993, n64994,
         n64995, n64996, n64997, n64998, n64999, n65000, n65001, n65002,
         n65003, n65004, n65005, n65006, n65007, n65008, n65009, n65010,
         n65011, n65012, n65013, n65014, n65015, n65016, n65017, n65018,
         n65019, n65020, n65021, n65022, n65023, n65024, n65025, n65026,
         n65027, n65028, n65029, n65030, n65031, n65032, n65033, n65034,
         n65035, n65036, n65037, n65038, n65039, n65040, n65041, n65042,
         n65043, n65044, n65045, n65046, n65047, n65048, n65049, n65050,
         n65051, n65052, n65053, n65054, n65055, n65056, n65057, n65058,
         n65059, n65060, n65061, n65062, n65063, n65064, n65065, n65066,
         n65067, n65068, n65069, n65070, n65071, n65072, n65073, n65074,
         n65075, n65076, n65077, n65078, n65079, n65080, n65081, n65082,
         n65083, n65084, n65085, n65086, n65087, n65088, n65089, n65090,
         n65091, n65092, n65093, n65094, n65095, n65096, n65097, n65098,
         n65099, n65100, n65101, n65102, n65103, n65104, n65105, n65106,
         n65107, n65108, n65109, n65110, n65111, n65112, n65113, n65114,
         n65115, n65116, n65117, n65118, n65119, n65120, n65121, n65122,
         n65123, n65124, n65125, n65126, n65127, n65128, n65129, n65130,
         n65131, n65132, n65133, n65134, n65135, n65136, n65137, n65138,
         n65139, n65140, n65141, n65142, n65143, n65144, n65145, n65146,
         n65147, n65148, n65149, n65150, n65151, n65152, n65153, n65154,
         n65155, n65156, n65157, n65158, n65159, n65160, n65161, n65162,
         n65163, n65164, n65165, n65166, n65167, n65168, n65169, n65170,
         n65171, n65172, n65173, n65174, n65175, n65176, n65177, n65178,
         n65179, n65180, n65181, n65182, n65183, n65184, n65185, n65186,
         n65187, n65188, n65189, n65190, n65191, n65192, n65193, n65194,
         n65195, n65196, n65197, n65198, n65199, n65201, n65202, n65203,
         n65204, n65205, n65206, n65207, n65208, n65209, n65210, n65211,
         n65212, n65213, n65214, n65215, n65216, n65217, n65218, n65219,
         n65220, n65221, n65222, n65224, n65225, n65226, n65227, n65228,
         n65229, n65230, n65231, n65232, n65233, n65234, n65235, n65236,
         n65237, n65238, n65239, n65240, n65241, n65242, n65243, n65244,
         n65245, n65246, n65247, n65248, n65249, n65250, n65251, n65252,
         n65253, n65254, n65255, n65256, n65257, n65258, n65259, n65260,
         n65261, n65262, n65263, n65264, n65265, n65266, n65267, n65268,
         n65269, n65270, n65271, n65272, n65273, n65274, n65275, n65276,
         n65277, n65278, n65279, n65280, n65281, n65282, n65283;

  INV_X1 U2 ( .I(n53102), .ZN(n53103) );
  INV_X1 U3 ( .I(n53174), .ZN(n53175) );
  INV_X1 U4 ( .I(n55052), .ZN(n55053) );
  INV_X1 U5 ( .I(n55534), .ZN(n55535) );
  INV_X1 U6 ( .I(n56949), .ZN(n56950) );
  INV_X1 U7 ( .I(n54734), .ZN(n54735) );
  INV_X1 U8 ( .I(n55765), .ZN(n55766) );
  NOR2_X1 U13 ( .A1(n21119), .A2(n21115), .ZN(n21114) );
  INV_X1 U18 ( .I(n55179), .ZN(n524) );
  NAND2_X1 U20 ( .A1(n54510), .A2(n54549), .ZN(n677) );
  AOI21_X1 U22 ( .A1(n53165), .A2(n61690), .B(n544), .ZN(n780) );
  NOR4_X1 U24 ( .A1(n51562), .A2(n51561), .A3(n51563), .A4(n56790), .ZN(n5896)
         );
  NOR2_X1 U25 ( .A1(n53466), .A2(n53506), .ZN(n5966) );
  AOI21_X1 U26 ( .A1(n55048), .A2(n55094), .B(n9068), .ZN(n8409) );
  OAI22_X1 U27 ( .A1(n15922), .A2(n53106), .B1(n53105), .B2(n53108), .ZN(
        n53123) );
  NAND2_X1 U28 ( .A1(n17959), .A2(n57997), .ZN(n54867) );
  INV_X1 U29 ( .I(n12156), .ZN(n544) );
  AND2_X1 U32 ( .A1(n53274), .A2(n53267), .Z(n1163) );
  NAND2_X1 U37 ( .A1(n6559), .A2(n6561), .ZN(n5114) );
  NAND2_X1 U39 ( .A1(n19222), .A2(n54530), .ZN(n54527) );
  INV_X1 U43 ( .I(n53329), .ZN(n213) );
  NOR2_X1 U44 ( .A1(n23448), .A2(n54723), .ZN(n54672) );
  NAND3_X1 U47 ( .A1(n54280), .A2(n54268), .A3(n19404), .ZN(n54234) );
  AOI21_X1 U48 ( .A1(n22516), .A2(n14778), .B(n4996), .ZN(n57087) );
  NOR2_X1 U50 ( .A1(n54010), .A2(n54001), .ZN(n53952) );
  NOR2_X1 U55 ( .A1(n54914), .A2(n17959), .ZN(n12690) );
  NOR2_X1 U66 ( .A1(n53148), .A2(n23856), .ZN(n3195) );
  NAND2_X1 U84 ( .A1(n19735), .A2(n53294), .ZN(n53280) );
  NAND2_X1 U97 ( .A1(n53324), .A2(n12923), .ZN(n53315) );
  NAND3_X1 U100 ( .A1(n12827), .A2(n53294), .A3(n4283), .ZN(n53274) );
  OR2_X1 U104 ( .A1(n16489), .A2(n7240), .Z(n15972) );
  INV_X1 U108 ( .I(n24535), .ZN(n53046) );
  NAND2_X1 U112 ( .A1(n55885), .A2(n55893), .ZN(n55870) );
  OR2_X1 U116 ( .A1(n56290), .A2(n22430), .Z(n1187) );
  NAND2_X1 U117 ( .A1(n56168), .A2(n56182), .ZN(n56173) );
  NOR2_X1 U123 ( .A1(n4336), .A2(n54913), .ZN(n2053) );
  INV_X2 U134 ( .I(n23956), .ZN(n22889) );
  NAND2_X1 U135 ( .A1(n24063), .A2(n14428), .ZN(n55341) );
  INV_X1 U154 ( .I(n56191), .ZN(n56171) );
  INV_X1 U158 ( .I(n59180), .ZN(n56313) );
  INV_X1 U163 ( .I(n24117), .ZN(n17799) );
  NOR2_X1 U167 ( .A1(n53699), .A2(n53672), .ZN(n53649) );
  NAND2_X1 U170 ( .A1(n56047), .A2(n56108), .ZN(n56072) );
  NOR2_X1 U182 ( .A1(n23956), .A2(n61361), .ZN(n12575) );
  NAND2_X1 U184 ( .A1(n53808), .A2(n53809), .ZN(n53789) );
  BUF_X2 U190 ( .I(n54902), .Z(n14635) );
  INV_X1 U193 ( .I(n18119), .ZN(n1582) );
  NOR2_X1 U199 ( .A1(n60115), .A2(n1450), .ZN(n15405) );
  OR2_X1 U200 ( .A1(n15245), .A2(n55387), .Z(n4955) );
  INV_X1 U204 ( .I(n53355), .ZN(n11963) );
  INV_X1 U208 ( .I(n24063), .ZN(n55364) );
  NOR2_X1 U209 ( .A1(n23318), .A2(n1591), .ZN(n56349) );
  BUF_X2 U212 ( .I(n8905), .Z(n2049) );
  INV_X2 U219 ( .I(n55768), .ZN(n55812) );
  INV_X2 U223 ( .I(n55868), .ZN(n55885) );
  INV_X2 U226 ( .I(n53729), .ZN(n25011) );
  INV_X1 U229 ( .I(n54257), .ZN(n54277) );
  INV_X2 U235 ( .I(n8905), .ZN(n1919) );
  BUF_X2 U237 ( .I(n25676), .Z(n25675) );
  INV_X2 U238 ( .I(n22362), .ZN(n9068) );
  BUF_X4 U250 ( .I(n53326), .Z(n17012) );
  INV_X2 U252 ( .I(n53146), .ZN(n53129) );
  AND2_X1 U254 ( .A1(n8397), .A2(n55011), .Z(n1162) );
  BUF_X4 U268 ( .I(n53243), .Z(n1232) );
  NAND2_X1 U275 ( .A1(n54683), .A2(n58283), .ZN(n8327) );
  AOI21_X1 U276 ( .A1(n56363), .A2(n13575), .B(n59827), .ZN(n18008) );
  OR2_X1 U291 ( .A1(n60181), .A2(n1260), .Z(n1182) );
  OR2_X1 U292 ( .A1(n56591), .A2(n20737), .Z(n16163) );
  AOI21_X1 U302 ( .A1(n7159), .A2(n12917), .B(n53548), .ZN(n10837) );
  AOI21_X1 U303 ( .A1(n53606), .A2(n53603), .B(n53605), .ZN(n12000) );
  AOI21_X1 U304 ( .A1(n58477), .A2(n13575), .B(n56364), .ZN(n5884) );
  AOI21_X1 U305 ( .A1(n52667), .A2(n21225), .B(n57058), .ZN(n21236) );
  INV_X1 U308 ( .I(n11521), .ZN(n55665) );
  AOI21_X1 U315 ( .A1(n54636), .A2(n54635), .B(n1373), .ZN(n3944) );
  NOR2_X1 U318 ( .A1(n1151), .A2(n4181), .ZN(n25107) );
  NAND2_X1 U323 ( .A1(n50933), .A2(n50951), .ZN(n75) );
  NOR2_X1 U324 ( .A1(n65011), .A2(n55414), .ZN(n54984) );
  OR2_X1 U327 ( .A1(n56433), .A2(n55986), .Z(n50899) );
  NAND3_X1 U330 ( .A1(n54779), .A2(n54780), .A3(n2200), .ZN(n2468) );
  NAND2_X1 U332 ( .A1(n52668), .A2(n57067), .ZN(n52667) );
  NOR2_X1 U345 ( .A1(n56268), .A2(n14324), .ZN(n55666) );
  NAND2_X1 U350 ( .A1(n54605), .A2(n60439), .ZN(n54779) );
  AND2_X1 U356 ( .A1(n55262), .A2(n63194), .Z(n1143) );
  NAND2_X1 U372 ( .A1(n1613), .A2(n54997), .ZN(n52946) );
  NOR4_X1 U378 ( .A1(n55470), .A2(n61282), .A3(n2180), .A4(n57901), .ZN(n55479) );
  NAND2_X1 U382 ( .A1(n55472), .A2(n55728), .ZN(n15315) );
  NAND2_X1 U387 ( .A1(n55438), .A2(n16073), .ZN(n55436) );
  INV_X1 U389 ( .I(n53877), .ZN(n53015) );
  NAND3_X1 U390 ( .A1(n54983), .A2(n55416), .A3(n52572), .ZN(n52574) );
  NAND3_X1 U391 ( .A1(n23157), .A2(n23974), .A3(n52840), .ZN(n53194) );
  OAI21_X1 U392 ( .A1(n53227), .A2(n53455), .B(n53580), .ZN(n53228) );
  INV_X1 U395 ( .I(n55679), .ZN(n55294) );
  NAND2_X1 U402 ( .A1(n51890), .A2(n56250), .ZN(n51185) );
  NAND2_X1 U409 ( .A1(n16948), .A2(n55412), .ZN(n55256) );
  INV_X2 U411 ( .I(n19167), .ZN(n1613) );
  INV_X2 U414 ( .I(n55442), .ZN(n55438) );
  OR2_X1 U425 ( .A1(n57026), .A2(n53212), .Z(n1151) );
  NOR2_X1 U427 ( .A1(n12574), .A2(n13232), .ZN(n53209) );
  INV_X1 U441 ( .I(n57026), .ZN(n23102) );
  NAND2_X1 U462 ( .A1(n24647), .A2(n52270), .ZN(n56598) );
  INV_X1 U463 ( .I(n61736), .ZN(n9089) );
  NAND3_X1 U465 ( .A1(n23025), .A2(n23476), .A3(n60002), .ZN(n53449) );
  INV_X2 U473 ( .I(n5227), .ZN(n15761) );
  INV_X1 U499 ( .I(n53858), .ZN(n22885) );
  INV_X2 U516 ( .I(n23873), .ZN(n12282) );
  NAND2_X1 U518 ( .A1(n54860), .A2(n18230), .ZN(n17937) );
  CLKBUF_X4 U520 ( .I(n6115), .Z(n3376) );
  INV_X1 U524 ( .I(n1459), .ZN(n53547) );
  BUF_X2 U530 ( .I(n14332), .Z(n12818) );
  INV_X2 U531 ( .I(n19811), .ZN(n23873) );
  INV_X2 U533 ( .I(n55444), .ZN(n5907) );
  INV_X1 U554 ( .I(n24787), .ZN(n13155) );
  INV_X1 U555 ( .I(n50633), .ZN(n531) );
  INV_X1 U561 ( .I(n50614), .ZN(n20008) );
  INV_X1 U571 ( .I(n19519), .ZN(n51615) );
  INV_X1 U572 ( .I(n25969), .ZN(n26201) );
  BUF_X2 U575 ( .I(n49727), .Z(n51522) );
  INV_X1 U576 ( .I(n23422), .ZN(n1465) );
  BUF_X2 U580 ( .I(n12379), .Z(n16969) );
  INV_X1 U581 ( .I(n56008), .ZN(n50718) );
  INV_X2 U585 ( .I(n2256), .ZN(n15487) );
  BUF_X2 U593 ( .I(n52596), .Z(n1625) );
  INV_X1 U602 ( .I(n24061), .ZN(n1901) );
  BUF_X2 U603 ( .I(n52201), .Z(n19530) );
  BUF_X2 U608 ( .I(n10825), .Z(n10398) );
  INV_X1 U611 ( .I(n26028), .ZN(n4245) );
  BUF_X2 U614 ( .I(n51510), .Z(n24758) );
  BUF_X2 U618 ( .I(n51810), .Z(n23422) );
  INV_X1 U620 ( .I(n52446), .ZN(n7744) );
  NAND3_X1 U630 ( .A1(n1096), .A2(n49894), .A3(n10263), .ZN(n25818) );
  NOR2_X1 U632 ( .A1(n16571), .A2(n11002), .ZN(n11001) );
  NAND3_X1 U633 ( .A1(n49728), .A2(n50400), .A3(n1381), .ZN(n49035) );
  NOR2_X1 U646 ( .A1(n12844), .A2(n26098), .ZN(n12843) );
  INV_X1 U648 ( .I(n49795), .ZN(n48433) );
  NOR3_X1 U650 ( .A1(n48928), .A2(n48927), .A3(n48926), .ZN(n48935) );
  AOI22_X1 U652 ( .A1(n49304), .A2(n49303), .B1(n24236), .B2(n24235), .ZN(
        n23659) );
  NOR3_X1 U659 ( .A1(n15131), .A2(n50120), .A3(n15130), .ZN(n15128) );
  NAND2_X1 U661 ( .A1(n49655), .A2(n3055), .ZN(n15005) );
  AOI21_X1 U663 ( .A1(n13692), .A2(n19107), .B(n48927), .ZN(n48373) );
  NOR2_X1 U672 ( .A1(n48716), .A2(n22867), .ZN(n50120) );
  NOR2_X1 U678 ( .A1(n48413), .A2(n1630), .ZN(n48417) );
  NAND3_X1 U685 ( .A1(n3347), .A2(n49581), .A3(n1637), .ZN(n48939) );
  NOR2_X1 U686 ( .A1(n9534), .A2(n15154), .ZN(n14858) );
  NOR2_X1 U687 ( .A1(n42), .A2(n15961), .ZN(n49569) );
  NAND2_X1 U690 ( .A1(n21189), .A2(n1377), .ZN(n10264) );
  INV_X1 U692 ( .I(n12595), .ZN(n48065) );
  NOR2_X1 U694 ( .A1(n13684), .A2(n50340), .ZN(n50261) );
  AND2_X1 U695 ( .A1(n49312), .A2(n1638), .Z(n1117) );
  NAND2_X1 U704 ( .A1(n25781), .A2(n19437), .ZN(n5763) );
  AOI21_X1 U705 ( .A1(n50275), .A2(n826), .B(n15967), .ZN(n14036) );
  OAI22_X1 U711 ( .A1(n50212), .A2(n47996), .B1(n7588), .B2(n50222), .ZN(
        n47997) );
  INV_X2 U716 ( .I(n18469), .ZN(n48811) );
  NAND2_X1 U723 ( .A1(n13684), .A2(n50340), .ZN(n49934) );
  INV_X1 U733 ( .I(n49049), .ZN(n49056) );
  NAND2_X1 U737 ( .A1(n49014), .A2(n49005), .ZN(n48453) );
  NAND2_X1 U746 ( .A1(n6716), .A2(n10563), .ZN(n49011) );
  NAND3_X1 U759 ( .A1(n46368), .A2(n4647), .A3(n5544), .ZN(n6894) );
  NAND2_X1 U760 ( .A1(n3461), .A2(n6977), .ZN(n467) );
  NOR2_X1 U764 ( .A1(n25018), .A2(n19589), .ZN(n47971) );
  NAND2_X1 U771 ( .A1(n48950), .A2(n22869), .ZN(n4310) );
  NAND2_X1 U772 ( .A1(n49029), .A2(n1381), .ZN(n6804) );
  NAND3_X1 U776 ( .A1(n48803), .A2(n18469), .A3(n6633), .ZN(n14097) );
  OAI21_X1 U779 ( .A1(n1291), .A2(n15793), .B(n50330), .ZN(n50332) );
  NOR2_X1 U780 ( .A1(n60719), .A2(n1205), .ZN(n6184) );
  NAND4_X1 U781 ( .A1(n47976), .A2(n49772), .A3(n48949), .A4(n22869), .ZN(
        n46090) );
  NAND3_X1 U782 ( .A1(n49408), .A2(n7086), .A3(n49272), .ZN(n46370) );
  INV_X1 U801 ( .I(n46850), .ZN(n50376) );
  NOR2_X1 U802 ( .A1(n1474), .A2(n2810), .ZN(n48073) );
  NAND2_X1 U805 ( .A1(n1643), .A2(n7952), .ZN(n21537) );
  NOR2_X1 U810 ( .A1(n13550), .A2(n57194), .ZN(n48774) );
  NAND2_X1 U821 ( .A1(n50331), .A2(n50257), .ZN(n50330) );
  NAND2_X1 U833 ( .A1(n50426), .A2(n23063), .ZN(n49253) );
  NOR2_X1 U841 ( .A1(n1382), .A2(n9983), .ZN(n49530) );
  NOR2_X1 U843 ( .A1(n19705), .A2(n7115), .ZN(n48819) );
  NOR2_X1 U852 ( .A1(n565), .A2(n3031), .ZN(n9379) );
  NAND2_X1 U857 ( .A1(n17874), .A2(n49600), .ZN(n48314) );
  NOR2_X1 U861 ( .A1(n50399), .A2(n25944), .ZN(n15167) );
  INV_X4 U878 ( .I(n20138), .ZN(n24374) );
  NAND2_X1 U888 ( .A1(n50378), .A2(n46850), .ZN(n50092) );
  INV_X2 U913 ( .I(n8044), .ZN(n19705) );
  INV_X2 U925 ( .I(n21870), .ZN(n13024) );
  INV_X1 U926 ( .I(n11246), .ZN(n17683) );
  INV_X2 U939 ( .I(n17379), .ZN(n48064) );
  INV_X1 U979 ( .I(n48701), .ZN(n49484) );
  INV_X2 U980 ( .I(n49637), .ZN(n1641) );
  NAND2_X1 U991 ( .A1(n48852), .A2(n49493), .ZN(n48701) );
  NAND2_X1 U1002 ( .A1(n4870), .A2(n46761), .ZN(n49888) );
  NAND2_X1 U1005 ( .A1(n22780), .A2(n49500), .ZN(n1631) );
  INV_X2 U1006 ( .I(n21320), .ZN(n47970) );
  AOI22_X1 U1028 ( .A1(n2151), .A2(n46023), .B1(n2150), .B2(n45634), .ZN(
        n26174) );
  NAND2_X1 U1032 ( .A1(n47841), .A2(n47840), .ZN(n87) );
  NOR2_X1 U1039 ( .A1(n11526), .A2(n16245), .ZN(n20274) );
  NAND2_X1 U1040 ( .A1(n48114), .A2(n13267), .ZN(n49859) );
  NAND2_X1 U1046 ( .A1(n2069), .A2(n20917), .ZN(n44074) );
  AND2_X1 U1064 ( .A1(n47574), .A2(n47573), .Z(n1071) );
  INV_X1 U1067 ( .I(n47297), .ZN(n1661) );
  NAND4_X1 U1073 ( .A1(n19740), .A2(n19739), .A3(n47244), .A4(n22303), .ZN(
        n19738) );
  NAND3_X1 U1080 ( .A1(n46048), .A2(n59861), .A3(n6497), .ZN(n6432) );
  NAND2_X1 U1081 ( .A1(n18227), .A2(n47407), .ZN(n43827) );
  NOR2_X1 U1085 ( .A1(n20624), .A2(n48640), .ZN(n12995) );
  INV_X1 U1089 ( .I(n46020), .ZN(n45601) );
  NAND2_X1 U1090 ( .A1(n64766), .A2(n48146), .ZN(n21819) );
  NAND2_X1 U1091 ( .A1(n43191), .A2(n47821), .ZN(n13971) );
  AOI22_X1 U1092 ( .A1(n47743), .A2(n59008), .B1(n63647), .B2(n47729), .ZN(
        n45914) );
  NAND3_X1 U1093 ( .A1(n17670), .A2(n24893), .A3(n47407), .ZN(n47408) );
  NOR2_X1 U1110 ( .A1(n47683), .A2(n45267), .ZN(n47420) );
  NAND2_X1 U1115 ( .A1(n23113), .A2(n1328), .ZN(n6660) );
  INV_X1 U1116 ( .I(n47217), .ZN(n537) );
  NAND4_X1 U1129 ( .A1(n3220), .A2(n48189), .A3(n2403), .A4(n23813), .ZN(n3219) );
  NOR3_X1 U1166 ( .A1(n47806), .A2(n47700), .A3(n11492), .ZN(n47808) );
  NAND3_X1 U1167 ( .A1(n12850), .A2(n1480), .A3(n23035), .ZN(n47511) );
  NOR2_X1 U1168 ( .A1(n47746), .A2(n62788), .ZN(n46737) );
  NAND2_X1 U1169 ( .A1(n6188), .A2(n6192), .ZN(n6187) );
  NOR2_X1 U1175 ( .A1(n7930), .A2(n47700), .ZN(n223) );
  AND2_X1 U1177 ( .A1(n47231), .A2(n10193), .Z(n6494) );
  INV_X1 U1181 ( .I(n22736), .ZN(n47371) );
  BUF_X2 U1184 ( .I(n45432), .Z(n47367) );
  NAND3_X1 U1193 ( .A1(n9368), .A2(n18570), .A3(n48199), .ZN(n47199) );
  INV_X1 U1194 ( .I(n3770), .ZN(n31) );
  NAND3_X1 U1197 ( .A1(n46025), .A2(n47298), .A3(n344), .ZN(n2149) );
  INV_X2 U1198 ( .I(n44065), .ZN(n45517) );
  INV_X1 U1200 ( .I(n46976), .ZN(n1655) );
  NOR2_X1 U1209 ( .A1(n47605), .A2(n61025), .ZN(n3770) );
  INV_X1 U1215 ( .I(n45075), .ZN(n46927) );
  INV_X1 U1227 ( .I(n3686), .ZN(n20140) );
  NAND2_X1 U1234 ( .A1(n23969), .A2(n23167), .ZN(n47896) );
  BUF_X2 U1236 ( .I(n13719), .Z(n47902) );
  NAND2_X1 U1245 ( .A1(n24545), .A2(n7816), .ZN(n48467) );
  INV_X1 U1246 ( .I(n22684), .ZN(n47531) );
  INV_X2 U1257 ( .I(n45591), .ZN(n47894) );
  INV_X1 U1268 ( .I(n8733), .ZN(n19921) );
  INV_X1 U1269 ( .I(n45889), .ZN(n47121) );
  NOR2_X1 U1272 ( .A1(n48135), .A2(n20996), .ZN(n7816) );
  INV_X2 U1273 ( .I(n1212), .ZN(n48518) );
  NOR2_X1 U1274 ( .A1(n47534), .A2(n24801), .ZN(n47016) );
  NOR2_X1 U1288 ( .A1(n45201), .A2(n47811), .ZN(n45202) );
  INV_X2 U1291 ( .I(n25007), .ZN(n47868) );
  INV_X2 U1292 ( .I(n45432), .ZN(n21451) );
  INV_X1 U1310 ( .I(n25148), .ZN(n48596) );
  CLKBUF_X4 U1316 ( .I(n46561), .Z(n1212) );
  INV_X2 U1328 ( .I(n43595), .ZN(n47881) );
  INV_X1 U1339 ( .I(n16557), .ZN(n115) );
  INV_X1 U1340 ( .I(n13853), .ZN(n44606) );
  INV_X1 U1342 ( .I(n46395), .ZN(n387) );
  INV_X1 U1345 ( .I(n15561), .ZN(n19766) );
  INV_X1 U1346 ( .I(n44386), .ZN(n8813) );
  INV_X1 U1348 ( .I(n12265), .ZN(n1671) );
  INV_X1 U1349 ( .I(n673), .ZN(n46436) );
  INV_X1 U1352 ( .I(n5989), .ZN(n5990) );
  INV_X1 U1360 ( .I(n8187), .ZN(n26167) );
  BUF_X2 U1373 ( .I(n43944), .Z(n46164) );
  INV_X1 U1375 ( .I(n9242), .ZN(n44895) );
  INV_X1 U1376 ( .I(n18728), .ZN(n132) );
  INV_X1 U1387 ( .I(n24278), .ZN(n1489) );
  INV_X1 U1406 ( .I(n23256), .ZN(n578) );
  INV_X2 U1407 ( .I(n24262), .ZN(n5360) );
  INV_X1 U1412 ( .I(n6564), .ZN(n11111) );
  INV_X1 U1414 ( .I(n44022), .ZN(n46211) );
  INV_X1 U1416 ( .I(n60556), .ZN(n1898) );
  INV_X2 U1418 ( .I(n20754), .ZN(n24262) );
  NOR2_X1 U1441 ( .A1(n20987), .A2(n43983), .ZN(n20173) );
  NOR2_X1 U1447 ( .A1(n41589), .A2(n401), .ZN(n7374) );
  OAI21_X1 U1455 ( .A1(n403), .A2(n402), .B(n7451), .ZN(n401) );
  NAND2_X1 U1464 ( .A1(n42343), .A2(n64346), .ZN(n9697) );
  NAND2_X1 U1468 ( .A1(n43608), .A2(n8171), .ZN(n19939) );
  AOI21_X1 U1469 ( .A1(n16156), .A2(n43475), .B(n43456), .ZN(n16746) );
  NAND2_X1 U1470 ( .A1(n20632), .A2(n1713), .ZN(n42679) );
  OAI21_X1 U1472 ( .A1(n40880), .A2(n39431), .B(n40882), .ZN(n39432) );
  OR2_X1 U1478 ( .A1(n5398), .A2(n62600), .Z(n16135) );
  NAND2_X1 U1482 ( .A1(n43917), .A2(n61743), .ZN(n43489) );
  OAI22_X1 U1487 ( .A1(n23819), .A2(n41644), .B1(n15091), .B2(n23811), .ZN(
        n42117) );
  INV_X1 U1488 ( .I(n2197), .ZN(n39880) );
  NOR2_X1 U1489 ( .A1(n24386), .A2(n1335), .ZN(n43366) );
  INV_X1 U1493 ( .I(n25672), .ZN(n170) );
  INV_X1 U1497 ( .I(n43012), .ZN(n41682) );
  OR2_X1 U1499 ( .A1(n43339), .A2(n23561), .Z(n993) );
  NOR2_X1 U1500 ( .A1(n42386), .A2(n42694), .ZN(n41971) );
  AND4_X1 U1501 ( .A1(n5341), .A2(n43573), .A3(n43572), .A4(n1397), .Z(n1025)
         );
  OAI21_X1 U1502 ( .A1(n41956), .A2(n5972), .B(n600), .ZN(n17303) );
  OAI21_X1 U1503 ( .A1(n12313), .A2(n42066), .B(n13751), .ZN(n20040) );
  OAI21_X1 U1505 ( .A1(n11229), .A2(n4106), .B(n1708), .ZN(n43603) );
  NAND2_X1 U1506 ( .A1(n42628), .A2(n577), .ZN(n660) );
  INV_X1 U1508 ( .I(n43872), .ZN(n402) );
  NOR2_X1 U1510 ( .A1(n8687), .A2(n41325), .ZN(n15878) );
  NOR2_X1 U1511 ( .A1(n42653), .A2(n1715), .ZN(n42745) );
  OAI21_X1 U1514 ( .A1(n42423), .A2(n43282), .B(n43107), .ZN(n6534) );
  INV_X1 U1516 ( .I(n43338), .ZN(n42590) );
  NAND2_X1 U1520 ( .A1(n22282), .A2(n41695), .ZN(n42736) );
  NAND2_X1 U1536 ( .A1(n22716), .A2(n23314), .ZN(n3204) );
  NAND2_X1 U1553 ( .A1(n601), .A2(n5972), .ZN(n600) );
  AND2_X1 U1554 ( .A1(n4322), .A2(n22939), .Z(n995) );
  NAND3_X1 U1567 ( .A1(n24981), .A2(n42998), .A3(n8343), .ZN(n39861) );
  NAND2_X1 U1568 ( .A1(n42653), .A2(n1335), .ZN(n42734) );
  NAND2_X1 U1576 ( .A1(n42140), .A2(n10004), .ZN(n42659) );
  INV_X1 U1582 ( .I(n18724), .ZN(n19742) );
  INV_X1 U1586 ( .I(n24386), .ZN(n42653) );
  INV_X1 U1587 ( .I(n24024), .ZN(n41695) );
  INV_X1 U1591 ( .I(n43416), .ZN(n601) );
  NOR2_X1 U1596 ( .A1(n43582), .A2(n43572), .ZN(n12154) );
  INV_X1 U1603 ( .I(n41757), .ZN(n42965) );
  NOR2_X1 U1606 ( .A1(n42985), .A2(n14409), .ZN(n43957) );
  INV_X1 U1613 ( .I(n8247), .ZN(n42369) );
  NAND2_X1 U1632 ( .A1(n19591), .A2(n43289), .ZN(n43111) );
  NAND3_X1 U1634 ( .A1(n21073), .A2(n43487), .A3(n43486), .ZN(n43914) );
  CLKBUF_X4 U1638 ( .I(n39841), .Z(n4659) );
  NAND2_X1 U1650 ( .A1(n12312), .A2(n43464), .ZN(n42065) );
  NOR2_X1 U1652 ( .A1(n42872), .A2(n43816), .ZN(n16545) );
  NAND2_X1 U1682 ( .A1(n8139), .A2(n5787), .ZN(n43869) );
  BUF_X2 U1687 ( .I(n41254), .Z(n43889) );
  NOR2_X1 U1695 ( .A1(n20922), .A2(n1301), .ZN(n5369) );
  INV_X1 U1702 ( .I(n5262), .ZN(n42001) );
  NAND2_X1 U1705 ( .A1(n43910), .A2(n43490), .ZN(n43776) );
  NOR2_X1 U1720 ( .A1(n25534), .A2(n42080), .ZN(n42396) );
  INV_X2 U1721 ( .I(n42993), .ZN(n11476) );
  INV_X2 U1727 ( .I(n41254), .ZN(n43897) );
  INV_X2 U1735 ( .I(n2879), .ZN(n42838) );
  NAND2_X1 U1736 ( .A1(n59898), .A2(n42600), .ZN(n42032) );
  NAND2_X1 U1739 ( .A1(n1301), .A2(n41614), .ZN(n42357) );
  INV_X2 U1740 ( .I(n20586), .ZN(n42585) );
  INV_X1 U1748 ( .I(n42027), .ZN(n42022) );
  OR2_X1 U1756 ( .A1(n26247), .A2(n20047), .Z(n25924) );
  INV_X2 U1768 ( .I(n42695), .ZN(n41970) );
  OAI21_X1 U1780 ( .A1(n13091), .A2(n41916), .B(n42242), .ZN(n13090) );
  NOR2_X1 U1783 ( .A1(n41080), .A2(n24862), .ZN(n15072) );
  NOR2_X1 U1788 ( .A1(n984), .A2(n40852), .ZN(n41080) );
  INV_X1 U1793 ( .I(n37996), .ZN(n40334) );
  NAND2_X1 U1797 ( .A1(n40471), .A2(n40470), .ZN(n40476) );
  NAND3_X1 U1803 ( .A1(n701), .A2(n40489), .A3(n40490), .ZN(n40497) );
  OAI21_X1 U1805 ( .A1(n40766), .A2(n40402), .B(n41423), .ZN(n11196) );
  AND2_X1 U1808 ( .A1(n42266), .A2(n40804), .Z(n5516) );
  NOR3_X1 U1815 ( .A1(n61264), .A2(n9980), .A3(n19438), .ZN(n42485) );
  OR2_X1 U1816 ( .A1(n6412), .A2(n42277), .Z(n999) );
  OR2_X1 U1820 ( .A1(n40107), .A2(n23711), .Z(n994) );
  NAND2_X1 U1822 ( .A1(n13034), .A2(n41255), .ZN(n41925) );
  NOR2_X1 U1823 ( .A1(n7696), .A2(n20047), .ZN(n7695) );
  NAND3_X1 U1830 ( .A1(n40049), .A2(n16962), .A3(n40103), .ZN(n25069) );
  NAND4_X1 U1836 ( .A1(n3536), .A2(n42300), .A3(n41269), .A4(n988), .ZN(n3535)
         );
  NAND2_X1 U1837 ( .A1(n40029), .A2(n14014), .ZN(n14013) );
  INV_X1 U1846 ( .I(n23399), .ZN(n40034) );
  INV_X1 U1866 ( .I(n3946), .ZN(n14815) );
  INV_X1 U1870 ( .I(n3505), .ZN(n40057) );
  INV_X1 U1877 ( .I(n8536), .ZN(n41194) );
  NOR2_X1 U1880 ( .A1(n41800), .A2(n41944), .ZN(n41802) );
  NAND3_X1 U1883 ( .A1(n42465), .A2(n24633), .A3(n23399), .ZN(n14524) );
  NAND2_X1 U1887 ( .A1(n9198), .A2(n40946), .ZN(n18610) );
  INV_X1 U1891 ( .I(n40614), .ZN(n39057) );
  INV_X1 U1895 ( .I(n40571), .ZN(n39486) );
  INV_X1 U1918 ( .I(n42277), .ZN(n41928) );
  NAND2_X1 U1925 ( .A1(n23610), .A2(n40708), .ZN(n11631) );
  NAND2_X1 U1935 ( .A1(n287), .A2(n25247), .ZN(n40791) );
  CLKBUF_X2 U1939 ( .I(n41182), .Z(n9915) );
  NOR2_X1 U1944 ( .A1(n60928), .A2(n12523), .ZN(n41014) );
  NAND2_X1 U1947 ( .A1(n40645), .A2(n7011), .ZN(n40648) );
  INV_X1 U1953 ( .I(n39007), .ZN(n41411) );
  NOR2_X1 U1957 ( .A1(n41212), .A2(n13050), .ZN(n40401) );
  INV_X1 U1966 ( .I(n37926), .ZN(n40465) );
  NAND2_X1 U1968 ( .A1(n38264), .A2(n41270), .ZN(n12264) );
  NAND2_X1 U1969 ( .A1(n40257), .A2(n37926), .ZN(n40932) );
  OAI21_X1 U1973 ( .A1(n41379), .A2(n41384), .B(n41122), .ZN(n2338) );
  NOR2_X1 U1978 ( .A1(n41874), .A2(n40842), .ZN(n40841) );
  INV_X1 U1989 ( .I(n41019), .ZN(n23355) );
  INV_X2 U2001 ( .I(n41182), .ZN(n11787) );
  NOR2_X1 U2006 ( .A1(n10954), .A2(n40994), .ZN(n40143) );
  NAND2_X1 U2007 ( .A1(n41950), .A2(n20348), .ZN(n13756) );
  NAND2_X1 U2033 ( .A1(n21255), .A2(n36648), .ZN(n40232) );
  INV_X2 U2052 ( .I(n36648), .ZN(n11126) );
  BUF_X2 U2063 ( .I(n40970), .Z(n18704) );
  BUF_X2 U2074 ( .I(n65271), .Z(n6058) );
  INV_X2 U2084 ( .I(n41383), .ZN(n41385) );
  INV_X2 U2094 ( .I(n19990), .ZN(n20046) );
  INV_X2 U2099 ( .I(n13434), .ZN(n41383) );
  INV_X2 U2100 ( .I(n8908), .ZN(n14165) );
  INV_X2 U2101 ( .I(n961), .ZN(n41444) );
  INV_X1 U2103 ( .I(n38861), .ZN(n1751) );
  INV_X1 U2107 ( .I(n17078), .ZN(n13696) );
  INV_X1 U2108 ( .I(n25376), .ZN(n38500) );
  INV_X1 U2110 ( .I(n65210), .ZN(n38308) );
  INV_X1 U2114 ( .I(n12880), .ZN(n15699) );
  INV_X1 U2117 ( .I(n13664), .ZN(n39358) );
  NAND2_X1 U2121 ( .A1(n8232), .A2(n8231), .ZN(n39372) );
  INV_X1 U2129 ( .I(n37556), .ZN(n8984) );
  INV_X1 U2130 ( .I(n39732), .ZN(n39460) );
  INV_X1 U2140 ( .I(n61949), .ZN(n628) );
  INV_X1 U2142 ( .I(n11829), .ZN(n38973) );
  BUF_X2 U2150 ( .I(n22452), .Z(n19381) );
  BUF_X2 U2154 ( .I(n23922), .Z(n12356) );
  INV_X1 U2156 ( .I(n51946), .ZN(n1902) );
  INV_X1 U2160 ( .I(n55034), .ZN(n18699) );
  INV_X1 U2161 ( .I(n56335), .ZN(n189) );
  BUF_X2 U2169 ( .I(n20470), .Z(n20234) );
  INV_X1 U2172 ( .I(n55792), .ZN(n22202) );
  NAND2_X1 U2173 ( .A1(n466), .A2(n1761), .ZN(n11210) );
  INV_X1 U2174 ( .I(n37967), .ZN(n1761) );
  NOR2_X1 U2182 ( .A1(n34377), .A2(n10087), .ZN(n490) );
  NOR2_X1 U2192 ( .A1(n36095), .A2(n36094), .ZN(n36103) );
  NAND3_X1 U2193 ( .A1(n19509), .A2(n60659), .A3(n25571), .ZN(n917) );
  NOR2_X1 U2202 ( .A1(n36786), .A2(n5978), .ZN(n5977) );
  OAI21_X1 U2206 ( .A1(n16127), .A2(n36665), .B(n63697), .ZN(n17664) );
  NAND2_X1 U2210 ( .A1(n36701), .A2(n36700), .ZN(n622) );
  NAND3_X1 U2220 ( .A1(n3692), .A2(n18583), .A3(n23357), .ZN(n22301) );
  NOR2_X1 U2222 ( .A1(n26052), .A2(n34841), .ZN(n11178) );
  NAND2_X1 U2226 ( .A1(n36009), .A2(n61747), .ZN(n7967) );
  NAND3_X1 U2228 ( .A1(n36507), .A2(n36586), .A3(n36506), .ZN(n8242) );
  NOR4_X1 U2233 ( .A1(n37271), .A2(n37270), .A3(n22733), .A4(n37268), .ZN(
        n37274) );
  NAND2_X1 U2235 ( .A1(n37420), .A2(n22595), .ZN(n16355) );
  NOR2_X1 U2238 ( .A1(n9633), .A2(n1419), .ZN(n35162) );
  INV_X1 U2241 ( .I(n17595), .ZN(n17720) );
  NOR2_X1 U2253 ( .A1(n23766), .A2(n18205), .ZN(n36698) );
  NOR2_X1 U2255 ( .A1(n37363), .A2(n2594), .ZN(n36586) );
  NAND2_X1 U2261 ( .A1(n3691), .A2(n37212), .ZN(n36978) );
  NAND2_X1 U2271 ( .A1(n8356), .A2(n36553), .ZN(n36372) );
  NAND2_X1 U2272 ( .A1(n36185), .A2(n36196), .ZN(n36111) );
  INV_X1 U2277 ( .I(n35888), .ZN(n31786) );
  NAND2_X1 U2285 ( .A1(n13297), .A2(n34872), .ZN(n7805) );
  NOR2_X1 U2329 ( .A1(n4263), .A2(n35361), .ZN(n36415) );
  NAND2_X1 U2332 ( .A1(n35885), .A2(n35883), .ZN(n34878) );
  NAND2_X1 U2336 ( .A1(n1776), .A2(n2362), .ZN(n12967) );
  NAND3_X1 U2346 ( .A1(n20431), .A2(n3590), .A3(n8487), .ZN(n484) );
  NAND2_X1 U2349 ( .A1(n22503), .A2(n23801), .ZN(n19893) );
  INV_X1 U2352 ( .I(n14915), .ZN(n37028) );
  OAI21_X1 U2357 ( .A1(n36437), .A2(n1419), .B(n36436), .ZN(n36438) );
  NOR2_X1 U2368 ( .A1(n22169), .A2(n3458), .ZN(n25163) );
  AND2_X1 U2373 ( .A1(n5205), .A2(n19473), .Z(n8438) );
  BUF_X2 U2407 ( .I(n33933), .Z(n37084) );
  NOR2_X1 U2408 ( .A1(n36852), .A2(n26213), .ZN(n36665) );
  NAND2_X1 U2409 ( .A1(n15171), .A2(n36926), .ZN(n14753) );
  NOR2_X1 U2416 ( .A1(n36170), .A2(n3458), .ZN(n2761) );
  NAND2_X1 U2418 ( .A1(n15743), .A2(n37184), .ZN(n37010) );
  CLKBUF_X4 U2429 ( .I(n34288), .Z(n8177) );
  CLKBUF_X8 U2430 ( .I(n32940), .Z(n8356) );
  BUF_X2 U2463 ( .I(n37358), .Z(n19573) );
  INV_X2 U2480 ( .I(n34469), .ZN(n24198) );
  NAND2_X1 U2482 ( .A1(n33813), .A2(n33812), .ZN(n33819) );
  NOR3_X1 U2487 ( .A1(n33759), .A2(n34798), .A3(n33468), .ZN(n15571) );
  NAND3_X1 U2504 ( .A1(n33595), .A2(n33600), .A3(n9679), .ZN(n33308) );
  OR2_X1 U2516 ( .A1(n35748), .A2(n61496), .Z(n15838) );
  NAND2_X1 U2517 ( .A1(n16614), .A2(n8780), .ZN(n32802) );
  NOR2_X1 U2532 ( .A1(n64958), .A2(n1345), .ZN(n14092) );
  INV_X1 U2533 ( .I(n35222), .ZN(n16506) );
  AND2_X1 U2534 ( .A1(n34193), .A2(n58447), .Z(n16066) );
  AOI21_X1 U2537 ( .A1(n34247), .A2(n15184), .B(n34246), .ZN(n15185) );
  OAI21_X1 U2540 ( .A1(n6527), .A2(n35628), .B(n35205), .ZN(n35209) );
  NOR2_X1 U2541 ( .A1(n34382), .A2(n1805), .ZN(n13735) );
  INV_X1 U2543 ( .I(n33337), .ZN(n2) );
  OAI21_X1 U2544 ( .A1(n2346), .A2(n64234), .B(n34188), .ZN(n19780) );
  INV_X1 U2550 ( .I(n34113), .ZN(n34118) );
  NAND2_X1 U2574 ( .A1(n61699), .A2(n33319), .ZN(n35630) );
  NAND2_X1 U2583 ( .A1(n33513), .A2(n25404), .ZN(n34964) );
  AND2_X1 U2585 ( .A1(n34221), .A2(n35799), .Z(n910) );
  NAND2_X1 U2595 ( .A1(n33433), .A2(n34587), .ZN(n11401) );
  NAND3_X1 U2598 ( .A1(n34142), .A2(n57898), .A3(n19663), .ZN(n19662) );
  AND2_X1 U2627 ( .A1(n35713), .A2(n17304), .Z(n16240) );
  INV_X1 U2629 ( .I(n33513), .ZN(n34542) );
  NAND2_X1 U2633 ( .A1(n35218), .A2(n17400), .ZN(n35663) );
  NAND2_X1 U2634 ( .A1(n14247), .A2(n65189), .ZN(n35020) );
  NAND2_X1 U2642 ( .A1(n34993), .A2(n12953), .ZN(n34994) );
  NAND2_X1 U2643 ( .A1(n31976), .A2(n35301), .ZN(n34748) );
  BUF_X2 U2644 ( .I(n31659), .Z(n33406) );
  CLKBUF_X2 U2645 ( .I(n3082), .Z(n8694) );
  INV_X1 U2650 ( .I(n34953), .ZN(n34569) );
  AND4_X1 U2657 ( .A1(n18300), .A2(n23834), .A3(n551), .A4(n34993), .Z(n903)
         );
  NAND2_X1 U2661 ( .A1(n4097), .A2(n19119), .ZN(n322) );
  INV_X1 U2691 ( .I(n17255), .ZN(n33550) );
  INV_X1 U2694 ( .I(n11182), .ZN(n35279) );
  NAND2_X1 U2703 ( .A1(n13487), .A2(n24089), .ZN(n17304) );
  NAND2_X1 U2704 ( .A1(n35735), .A2(n18651), .ZN(n34414) );
  CLKBUF_X2 U2710 ( .I(n34035), .Z(n2635) );
  INV_X1 U2715 ( .I(n64603), .ZN(n33961) );
  NAND2_X1 U2719 ( .A1(n31767), .A2(n32892), .ZN(n32889) );
  NOR2_X1 U2721 ( .A1(n32914), .A2(n33503), .ZN(n30960) );
  OAI21_X1 U2723 ( .A1(n60669), .A2(n10504), .B(n35765), .ZN(n18395) );
  INV_X2 U2727 ( .I(n34783), .ZN(n33776) );
  INV_X1 U2730 ( .I(n31842), .ZN(n16481) );
  INV_X1 U2731 ( .I(n34161), .ZN(n34002) );
  NAND2_X1 U2744 ( .A1(n16402), .A2(n1546), .ZN(n34438) );
  INV_X2 U2745 ( .I(n12658), .ZN(n35218) );
  BUF_X2 U2746 ( .I(n32529), .Z(n33568) );
  INV_X4 U2747 ( .I(n1547), .ZN(n34658) );
  NOR2_X1 U2750 ( .A1(n34530), .A2(n34961), .ZN(n33503) );
  INV_X1 U2752 ( .I(n59138), .ZN(n33621) );
  INV_X2 U2754 ( .I(n25844), .ZN(n35709) );
  INV_X1 U2767 ( .I(n1542), .ZN(n5085) );
  INV_X1 U2771 ( .I(n34331), .ZN(n35774) );
  INV_X1 U2776 ( .I(n227), .ZN(n31659) );
  INV_X2 U2777 ( .I(n8456), .ZN(n32846) );
  INV_X2 U2780 ( .I(n2923), .ZN(n5604) );
  INV_X1 U2785 ( .I(n24831), .ZN(n665) );
  INV_X1 U2789 ( .I(n15464), .ZN(n33186) );
  INV_X1 U2793 ( .I(n14665), .ZN(n32085) );
  INV_X1 U2794 ( .I(n18964), .ZN(n24666) );
  INV_X1 U2796 ( .I(n5436), .ZN(n5437) );
  INV_X1 U2798 ( .I(n31344), .ZN(n33891) );
  INV_X1 U2800 ( .I(n32335), .ZN(n32590) );
  INV_X1 U2803 ( .I(n14563), .ZN(n19069) );
  BUF_X2 U2824 ( .I(n33856), .Z(n23869) );
  BUF_X2 U2828 ( .I(n15732), .Z(n15733) );
  INV_X1 U2838 ( .I(n31599), .ZN(n32035) );
  OAI21_X1 U2852 ( .A1(n30818), .A2(n30822), .B(n29932), .ZN(n29836) );
  AOI21_X1 U2853 ( .A1(n30891), .A2(n603), .B(n3486), .ZN(n29723) );
  AOI21_X1 U2859 ( .A1(n28290), .A2(n11568), .B(n11566), .ZN(n28298) );
  NOR2_X1 U2860 ( .A1(n29279), .A2(n8752), .ZN(n22099) );
  NOR3_X1 U2863 ( .A1(n17786), .A2(n17785), .A3(n17784), .ZN(n17783) );
  NAND3_X1 U2865 ( .A1(n30776), .A2(n20551), .A3(n62202), .ZN(n20695) );
  OAI21_X1 U2866 ( .A1(n2253), .A2(n100), .B(n16631), .ZN(n2296) );
  INV_X1 U2870 ( .I(n33185), .ZN(n1985) );
  NAND2_X1 U2872 ( .A1(n31168), .A2(n327), .ZN(n31169) );
  INV_X1 U2873 ( .I(n28579), .ZN(n124) );
  NAND2_X1 U2882 ( .A1(n30162), .A2(n60111), .ZN(n17490) );
  OAI21_X1 U2884 ( .A1(n29902), .A2(n29569), .B(n29905), .ZN(n11816) );
  AOI21_X1 U2892 ( .A1(n29808), .A2(n16219), .B(n1350), .ZN(n9002) );
  NAND4_X1 U2894 ( .A1(n30884), .A2(n30885), .A3(n31241), .A4(n23008), .ZN(
        n20077) );
  CLKBUF_X2 U2902 ( .I(Key[34]), .Z(n53685) );
  OAI21_X1 U2908 ( .A1(n27354), .A2(n22838), .B(n22837), .ZN(n27363) );
  NAND2_X1 U2909 ( .A1(n30223), .A2(n770), .ZN(n29808) );
  NAND2_X1 U2912 ( .A1(n17281), .A2(n17483), .ZN(n17481) );
  NOR2_X1 U2914 ( .A1(n29564), .A2(n11263), .ZN(n28958) );
  AOI22_X1 U2916 ( .A1(n29262), .A2(n1317), .B1(n29268), .B2(n8218), .ZN(
        n29263) );
  NAND4_X1 U2919 ( .A1(n59658), .A2(n24852), .A3(n10068), .A4(n2795), .ZN(
        n5985) );
  AOI22_X1 U2921 ( .A1(n14350), .A2(n12376), .B1(n19572), .B2(n30385), .ZN(
        n29498) );
  AND2_X1 U2928 ( .A1(n19363), .A2(n23705), .Z(n770) );
  NAND2_X1 U2929 ( .A1(n30455), .A2(n20859), .ZN(n30451) );
  NOR2_X1 U2940 ( .A1(n23055), .A2(n21532), .ZN(n30212) );
  CLKBUF_X2 U2946 ( .I(n21512), .Z(n3426) );
  BUF_X2 U2948 ( .I(n46180), .Z(n1190) );
  NAND2_X1 U2956 ( .A1(n31053), .A2(n579), .ZN(n30687) );
  NAND3_X1 U2958 ( .A1(n12165), .A2(n30050), .A3(n12164), .ZN(n12163) );
  NAND3_X1 U2960 ( .A1(n29959), .A2(n18472), .A3(n30767), .ZN(n26439) );
  NAND2_X1 U2961 ( .A1(n1859), .A2(n1253), .ZN(n30443) );
  NAND3_X1 U2962 ( .A1(n30369), .A2(n30375), .A3(n1437), .ZN(n5859) );
  NAND4_X1 U2965 ( .A1(n31243), .A2(n9654), .A3(n19255), .A4(n1435), .ZN(
        n24238) );
  NAND2_X1 U2970 ( .A1(n24504), .A2(n22411), .ZN(n596) );
  OR2_X1 U2983 ( .A1(n30845), .A2(n8470), .Z(n30214) );
  NAND2_X1 U2986 ( .A1(n28933), .A2(n29209), .ZN(n30684) );
  NOR2_X1 U2992 ( .A1(n10629), .A2(n5631), .ZN(n30099) );
  NAND2_X1 U2998 ( .A1(n30334), .A2(n23140), .ZN(n29943) );
  INV_X2 U3013 ( .I(n7426), .ZN(n1278) );
  NOR2_X1 U3018 ( .A1(n22374), .A2(n26740), .ZN(n30239) );
  NAND2_X1 U3026 ( .A1(n17745), .A2(n29747), .ZN(n30780) );
  NAND2_X1 U3028 ( .A1(n30455), .A2(n18402), .ZN(n30360) );
  NOR2_X1 U3030 ( .A1(n30695), .A2(n31055), .ZN(n29034) );
  AND2_X1 U3034 ( .A1(n24564), .A2(n20391), .Z(n759) );
  INV_X1 U3040 ( .I(n27789), .ZN(n1849) );
  NAND2_X1 U3042 ( .A1(n23988), .A2(n13731), .ZN(n30303) );
  NOR2_X1 U3044 ( .A1(n2269), .A2(n61622), .ZN(n2369) );
  AOI21_X1 U3045 ( .A1(n11909), .A2(n12893), .B(n603), .ZN(n5692) );
  NOR2_X1 U3049 ( .A1(n30376), .A2(n23004), .ZN(n20606) );
  INV_X1 U3089 ( .I(n30087), .ZN(n30085) );
  INV_X2 U3093 ( .I(n31074), .ZN(n25384) );
  BUF_X2 U3097 ( .I(n4921), .Z(n9434) );
  NAND2_X1 U3099 ( .A1(n29202), .A2(n12130), .ZN(n30224) );
  NOR2_X1 U3106 ( .A1(n13320), .A2(n15533), .ZN(n28762) );
  CLKBUF_X2 U3107 ( .I(Key[72]), .Z(n54517) );
  NOR2_X1 U3115 ( .A1(n14200), .A2(n29913), .ZN(n17719) );
  INV_X1 U3117 ( .I(n29889), .ZN(n603) );
  INV_X2 U3120 ( .I(n9153), .ZN(n31085) );
  INV_X1 U3130 ( .I(n30255), .ZN(n9047) );
  INV_X1 U3137 ( .I(n15791), .ZN(n29521) );
  INV_X2 U3146 ( .I(n24196), .ZN(n30211) );
  BUF_X2 U3151 ( .I(Key[20]), .Z(n51019) );
  NAND2_X1 U3163 ( .A1(n21832), .A2(n15689), .ZN(n24448) );
  OAI21_X1 U3164 ( .A1(n15196), .A2(n15195), .B(n29173), .ZN(n29201) );
  OAI21_X1 U3176 ( .A1(n29116), .A2(n2142), .B(n29115), .ZN(n29200) );
  NOR2_X1 U3178 ( .A1(n28213), .A2(n28214), .ZN(n13623) );
  NOR4_X1 U3180 ( .A1(n26313), .A2(n26637), .A3(n2704), .A4(n26312), .ZN(
        n26314) );
  NAND2_X1 U3184 ( .A1(n26266), .A2(n11134), .ZN(n11133) );
  NAND3_X1 U3185 ( .A1(n29329), .A2(n29328), .A3(n29330), .ZN(n29331) );
  AND2_X1 U3188 ( .A1(n28370), .A2(n26331), .Z(n15904) );
  NAND3_X1 U3190 ( .A1(n27217), .A2(n29295), .A3(n1360), .ZN(n27225) );
  NAND4_X1 U3193 ( .A1(n27694), .A2(n27695), .A3(n27696), .A4(n27697), .ZN(
        n27706) );
  NAND2_X1 U3195 ( .A1(n11374), .A2(n29652), .ZN(n10917) );
  AOI21_X1 U3196 ( .A1(n29653), .A2(n29652), .B(n29668), .ZN(n29655) );
  NOR2_X1 U3199 ( .A1(n29129), .A2(n8436), .ZN(n27969) );
  OAI22_X1 U3200 ( .A1(n62406), .A2(n8436), .B1(n8613), .B2(n10399), .ZN(
        n15211) );
  NAND2_X1 U3201 ( .A1(n11605), .A2(n29166), .ZN(n14227) );
  NOR3_X2 U3202 ( .A1(n27147), .A2(n27146), .A3(n27145), .ZN(n4706) );
  NAND2_X1 U3213 ( .A1(n1931), .A2(n27970), .ZN(n13805) );
  NAND2_X1 U3215 ( .A1(n23665), .A2(n2513), .ZN(n28218) );
  NOR2_X1 U3217 ( .A1(n61643), .A2(n28035), .ZN(n28037) );
  OAI21_X1 U3218 ( .A1(n27115), .A2(n11267), .B(n57318), .ZN(n14222) );
  NAND2_X1 U3222 ( .A1(n27405), .A2(n3087), .ZN(n27270) );
  NAND3_X1 U3226 ( .A1(n28225), .A2(n19170), .A3(n23166), .ZN(n14149) );
  NOR3_X1 U3227 ( .A1(n26635), .A2(n22902), .A3(n10321), .ZN(n26636) );
  INV_X1 U3231 ( .I(n8436), .ZN(n22929) );
  INV_X1 U3238 ( .I(n28230), .ZN(n28031) );
  NOR2_X1 U3245 ( .A1(n28472), .A2(n28630), .ZN(n29713) );
  INV_X1 U3248 ( .I(n28396), .ZN(n28416) );
  INV_X1 U3251 ( .I(n7775), .ZN(n26580) );
  NAND2_X1 U3252 ( .A1(n28072), .A2(n23586), .ZN(n26524) );
  NAND2_X1 U3256 ( .A1(n26654), .A2(n21132), .ZN(n27579) );
  NAND2_X1 U3258 ( .A1(n29381), .A2(n29652), .ZN(n27338) );
  INV_X1 U3259 ( .I(n29128), .ZN(n26732) );
  INV_X1 U3260 ( .I(n26034), .ZN(n5306) );
  INV_X1 U3262 ( .I(n21132), .ZN(n27577) );
  INV_X1 U3263 ( .I(n27410), .ZN(n1880) );
  INV_X1 U3264 ( .I(n8113), .ZN(n10805) );
  NAND2_X1 U3266 ( .A1(n20782), .A2(n21068), .ZN(n91) );
  NAND2_X1 U3267 ( .A1(n8113), .A2(n58601), .ZN(n29669) );
  NAND2_X1 U3277 ( .A1(n29682), .A2(n25341), .ZN(n27678) );
  NAND2_X1 U3282 ( .A1(n28030), .A2(n28033), .ZN(n27094) );
  INV_X1 U3287 ( .I(n29697), .ZN(n29682) );
  INV_X1 U3296 ( .I(n11514), .ZN(n29161) );
  INV_X1 U3305 ( .I(n20581), .ZN(n28640) );
  INV_X1 U3307 ( .I(n7371), .ZN(n29146) );
  INV_X1 U3308 ( .I(n20070), .ZN(n1566) );
  NAND2_X1 U3314 ( .A1(n23876), .A2(n28271), .ZN(n28027) );
  NAND2_X1 U3320 ( .A1(n16446), .A2(n9940), .ZN(n28384) );
  NOR2_X1 U3326 ( .A1(n28033), .A2(n27051), .ZN(n26577) );
  NAND3_X1 U3327 ( .A1(n28804), .A2(n18515), .A3(n28813), .ZN(n27323) );
  INV_X1 U3329 ( .I(n1321), .ZN(n28254) );
  INV_X1 U3330 ( .I(n856), .ZN(n12030) );
  INV_X1 U3331 ( .I(n27381), .ZN(n28245) );
  OAI21_X1 U3333 ( .A1(n22810), .A2(n19522), .B(n10914), .ZN(n27430) );
  NOR2_X1 U3336 ( .A1(n27622), .A2(n10914), .ZN(n26599) );
  OAI21_X1 U3339 ( .A1(n27232), .A2(n14633), .B(n27470), .ZN(n20510) );
  INV_X1 U3341 ( .I(n29673), .ZN(n29375) );
  NOR2_X1 U3342 ( .A1(n26260), .A2(n64155), .ZN(n26517) );
  NAND2_X1 U3343 ( .A1(n24498), .A2(n28076), .ZN(n16903) );
  INV_X1 U3348 ( .I(n26945), .ZN(n28831) );
  INV_X1 U3352 ( .I(n7760), .ZN(n26043) );
  INV_X1 U3356 ( .I(n26270), .ZN(n28076) );
  INV_X2 U3362 ( .I(n28187), .ZN(n29691) );
  INV_X1 U3364 ( .I(n26192), .ZN(n19972) );
  INV_X1 U3365 ( .I(n2066), .ZN(n28873) );
  INV_X1 U3368 ( .I(n27051), .ZN(n28030) );
  NOR2_X1 U3373 ( .A1(n28588), .A2(n28595), .ZN(n28846) );
  NOR2_X1 U3382 ( .A1(n1894), .A2(n1447), .ZN(n28351) );
  NAND2_X1 U3394 ( .A1(n1360), .A2(n27494), .ZN(n26969) );
  NOR2_X1 U3396 ( .A1(n19452), .A2(n10403), .ZN(n27498) );
  INV_X1 U3408 ( .I(n28221), .ZN(n27996) );
  INV_X2 U3416 ( .I(n27292), .ZN(n29144) );
  INV_X1 U3419 ( .I(n27478), .ZN(n27228) );
  BUF_X2 U3427 ( .I(n27366), .Z(n23170) );
  BUF_X2 U3428 ( .I(n26691), .Z(n23504) );
  NAND2_X1 U3429 ( .A1(n19619), .A2(n19883), .ZN(n19566) );
  INV_X1 U3430 ( .I(n24039), .ZN(n26344) );
  INV_X1 U3431 ( .I(n26279), .ZN(n27135) );
  INV_X2 U3434 ( .I(n14903), .ZN(n27533) );
  INV_X2 U3438 ( .I(n26691), .ZN(n10403) );
  BUF_X2 U3442 ( .I(Key[145]), .Z(n56155) );
  NAND3_X2 U3448 ( .A1(n32968), .A2(n32969), .A3(n32967), .ZN(n32970) );
  NAND2_X2 U3449 ( .A1(n18831), .A2(n3399), .ZN(n3398) );
  INV_X4 U3457 ( .I(n23914), .ZN(n34253) );
  INV_X2 U3460 ( .I(n42395), .ZN(n42403) );
  NOR2_X2 U3461 ( .A1(n14260), .A2(n64651), .ZN(n44451) );
  BUF_X2 U3462 ( .I(n30535), .Z(n33143) );
  BUF_X2 U3468 ( .I(n15410), .Z(n20948) );
  BUF_X2 U3470 ( .I(n25690), .Z(n9660) );
  INV_X2 U3472 ( .I(n13950), .ZN(n35318) );
  INV_X2 U3485 ( .I(n14242), .ZN(n306) );
  INV_X2 U3491 ( .I(n11590), .ZN(n41379) );
  NAND2_X2 U3494 ( .A1(n42509), .A2(n42508), .ZN(n2800) );
  NAND2_X2 U3502 ( .A1(n37931), .A2(n3306), .ZN(n41511) );
  NOR2_X2 U3531 ( .A1(n55101), .A2(n54960), .ZN(n55097) );
  OAI21_X2 U3532 ( .A1(n2658), .A2(n27932), .B(n2657), .ZN(n2656) );
  NOR2_X2 U3534 ( .A1(n26842), .A2(n30122), .ZN(n26846) );
  BUF_X4 U3535 ( .I(n40979), .Z(n42347) );
  AOI21_X1 U3543 ( .A1(n42967), .A2(n18721), .B(n17152), .ZN(n17151) );
  NAND2_X2 U3547 ( .A1(n43460), .A2(n12312), .ZN(n42962) );
  NOR3_X2 U3555 ( .A1(n54485), .A2(n54484), .A3(n54483), .ZN(n54486) );
  NOR2_X2 U3557 ( .A1(n60433), .A2(n54565), .ZN(n54572) );
  NAND2_X2 U3559 ( .A1(n15071), .A2(n35974), .ZN(n19699) );
  NOR2_X2 U3561 ( .A1(n45991), .A2(n59802), .ZN(n1663) );
  NAND2_X2 U3567 ( .A1(n21102), .A2(n45807), .ZN(n19652) );
  INV_X4 U3571 ( .I(n36746), .ZN(n36338) );
  NAND2_X2 U3578 ( .A1(n22464), .A2(n4428), .ZN(n16227) );
  NAND2_X2 U3579 ( .A1(n14240), .A2(n40277), .ZN(n5537) );
  NAND2_X2 U3580 ( .A1(n7952), .A2(n8251), .ZN(n15436) );
  INV_X2 U3587 ( .I(n8293), .ZN(n15731) );
  NAND2_X2 U3593 ( .A1(n47515), .A2(n10333), .ZN(n47512) );
  NAND3_X2 U3603 ( .A1(n41079), .A2(n9790), .A3(n40854), .ZN(n40849) );
  OAI21_X1 U3606 ( .A1(n43581), .A2(n5398), .B(n11018), .ZN(n2625) );
  AOI21_X2 U3615 ( .A1(n48125), .A2(n48124), .B(n22712), .ZN(n22711) );
  NOR2_X2 U3620 ( .A1(n5531), .A2(n57199), .ZN(n41017) );
  INV_X4 U3627 ( .I(n39427), .ZN(n2735) );
  INV_X4 U3635 ( .I(n36838), .ZN(n36852) );
  NOR3_X2 U3637 ( .A1(n41157), .A2(n15943), .A3(n41156), .ZN(n5212) );
  NAND2_X2 U3649 ( .A1(n10140), .A2(n31189), .ZN(n31571) );
  OAI21_X2 U3653 ( .A1(n27897), .A2(n17274), .B(n1889), .ZN(n28644) );
  NAND4_X2 U3656 ( .A1(n45691), .A2(n45692), .A3(n45690), .A4(n45689), .ZN(
        n45698) );
  BUF_X4 U3668 ( .I(n34350), .Z(n4591) );
  NAND2_X2 U3677 ( .A1(n49224), .A2(n5946), .ZN(n49152) );
  INV_X4 U3689 ( .I(n61164), .ZN(n43912) );
  INV_X4 U3697 ( .I(n18385), .ZN(n8474) );
  NOR2_X2 U3704 ( .A1(n5004), .A2(n5003), .ZN(n13459) );
  INV_X2 U3707 ( .I(n38781), .ZN(n24663) );
  NAND2_X2 U3709 ( .A1(n22794), .A2(n18335), .ZN(n56572) );
  NOR2_X2 U3714 ( .A1(n21388), .A2(n13081), .ZN(n18989) );
  NAND2_X2 U3715 ( .A1(n18989), .A2(n34305), .ZN(n34775) );
  NOR2_X2 U3719 ( .A1(n18335), .A2(n25134), .ZN(n56282) );
  AOI21_X2 U3723 ( .A1(n33952), .A2(n33953), .B(n20066), .ZN(n20065) );
  INV_X4 U3725 ( .I(n617), .ZN(n49382) );
  BUF_X4 U3729 ( .I(n33872), .Z(n8329) );
  NOR3_X2 U3732 ( .A1(n6407), .A2(n19529), .A3(n28848), .ZN(n4832) );
  NAND2_X2 U3734 ( .A1(n19948), .A2(n35148), .ZN(n35355) );
  INV_X4 U3735 ( .I(n42387), .ZN(n41972) );
  NOR2_X2 U3737 ( .A1(n24644), .A2(n3566), .ZN(n42262) );
  NAND2_X2 U3743 ( .A1(n11150), .A2(n23278), .ZN(n47622) );
  INV_X4 U3748 ( .I(n30492), .ZN(n25527) );
  NAND2_X2 U3749 ( .A1(n14446), .A2(n26041), .ZN(n54047) );
  AOI22_X2 U3755 ( .A1(n22127), .A2(n21023), .B1(n16062), .B2(n30073), .ZN(
        n22126) );
  BUF_X4 U3758 ( .I(n42225), .Z(n5980) );
  NAND3_X2 U3801 ( .A1(n5063), .A2(n5062), .A3(n5061), .ZN(n5060) );
  NAND3_X2 U3808 ( .A1(n40291), .A2(n60153), .A3(n321), .ZN(n40230) );
  OAI21_X2 U3810 ( .A1(n6937), .A2(n11497), .B(n41615), .ZN(n14240) );
  AOI22_X2 U3811 ( .A1(n34276), .A2(n34786), .B1(n34277), .B2(n62373), .ZN(
        n34285) );
  BUF_X4 U3816 ( .I(n41987), .Z(n22999) );
  OAI21_X2 U3823 ( .A1(n59376), .A2(n3306), .B(n3304), .ZN(n40249) );
  NAND3_X2 U3845 ( .A1(n17306), .A2(n27284), .A3(n28560), .ZN(n17305) );
  BUF_X4 U3851 ( .I(n24170), .Z(n24169) );
  INV_X4 U3864 ( .I(n33898), .ZN(n33204) );
  INV_X2 U3866 ( .I(n21036), .ZN(n40038) );
  INV_X2 U3868 ( .I(n34378), .ZN(n36520) );
  NAND3_X1 U3886 ( .A1(n55101), .A2(n62822), .A3(n591), .ZN(n3371) );
  NAND2_X1 U3888 ( .A1(n63039), .A2(n59180), .ZN(n56311) );
  INV_X1 U3889 ( .I(n61914), .ZN(n1598) );
  NAND2_X1 U3892 ( .A1(n9067), .A2(n55102), .ZN(n3369) );
  NOR2_X1 U3893 ( .A1(n55014), .A2(n1960), .ZN(n1959) );
  NAND2_X1 U3894 ( .A1(n9102), .A2(n55068), .ZN(n10773) );
  NOR2_X1 U3897 ( .A1(n34355), .A2(n34350), .ZN(n21196) );
  OR2_X1 U3901 ( .A1(n54006), .A2(n2851), .Z(n21121) );
  NOR2_X1 U3905 ( .A1(n9067), .A2(n54960), .ZN(n3372) );
  NOR2_X1 U3906 ( .A1(n9097), .A2(n55075), .ZN(n9093) );
  OAI21_X1 U3907 ( .A1(n55077), .A2(n55089), .B(n62822), .ZN(n9094) );
  INV_X1 U3915 ( .I(n41925), .ZN(n10201) );
  INV_X1 U3918 ( .I(n53437), .ZN(n12956) );
  OAI21_X1 U3922 ( .A1(n10773), .A2(n55057), .B(n55074), .ZN(n10772) );
  OAI21_X1 U3927 ( .A1(n11521), .A2(n61321), .B(n13022), .ZN(n13021) );
  NAND2_X1 U3929 ( .A1(n54192), .A2(n54197), .ZN(n54193) );
  NAND2_X1 U3934 ( .A1(n21590), .A2(n3525), .ZN(n53142) );
  NAND4_X1 U3943 ( .A1(n10774), .A2(n10772), .A3(n55059), .A4(n55058), .ZN(
        n9831) );
  NAND2_X1 U3950 ( .A1(n53522), .A2(n53529), .ZN(n14022) );
  NAND2_X1 U3953 ( .A1(n53355), .A2(n52762), .ZN(n53347) );
  NAND2_X1 U3957 ( .A1(n53492), .A2(n9595), .ZN(n53517) );
  NAND2_X1 U3958 ( .A1(n54614), .A2(n54430), .ZN(n4241) );
  NAND2_X1 U3961 ( .A1(n5193), .A2(n5172), .ZN(n56162) );
  INV_X1 U3964 ( .I(n2866), .ZN(n15937) );
  OAI21_X1 U3965 ( .A1(n2866), .A2(n63022), .B(n63020), .ZN(n2865) );
  NAND2_X1 U3966 ( .A1(n22749), .A2(n4319), .ZN(n13333) );
  BUF_X4 U3969 ( .I(n48536), .Z(n22464) );
  OAI21_X1 U3972 ( .A1(n55097), .A2(n11548), .B(n4985), .ZN(n55058) );
  AOI22_X1 U3973 ( .A1(n55095), .A2(n4985), .B1(n11548), .B2(n25220), .ZN(
        n55085) );
  NAND2_X1 U3982 ( .A1(n37354), .A2(n23226), .ZN(n18123) );
  INV_X1 U3983 ( .I(n53797), .ZN(n53825) );
  INV_X1 U3987 ( .I(n13503), .ZN(n53775) );
  NAND2_X1 U3988 ( .A1(n46910), .A2(n179), .ZN(n16879) );
  AND2_X1 U3989 ( .A1(n20615), .A2(n53673), .Z(n1181) );
  NOR2_X1 U3990 ( .A1(n25220), .A2(n15520), .ZN(n55042) );
  INV_X1 U3997 ( .I(n53676), .ZN(n53702) );
  NAND2_X1 U3998 ( .A1(n19475), .A2(n53676), .ZN(n53687) );
  AOI22_X1 U4004 ( .A1(n54672), .A2(n54755), .B1(n54671), .B2(n54759), .ZN(
        n18564) );
  NAND2_X1 U4014 ( .A1(n56695), .A2(n23785), .ZN(n56696) );
  NAND2_X1 U4016 ( .A1(n56759), .A2(n51565), .ZN(n5892) );
  NAND3_X1 U4023 ( .A1(n20458), .A2(n49065), .A3(n8298), .ZN(n49839) );
  OAI22_X1 U4029 ( .A1(n58232), .A2(n46958), .B1(n58244), .B2(n59406), .ZN(
        n46957) );
  AND2_X1 U4030 ( .A1(n7138), .A2(n1367), .Z(n1170) );
  NOR2_X1 U4042 ( .A1(n28225), .A2(n23170), .ZN(n431) );
  NAND2_X1 U4047 ( .A1(n54978), .A2(n24075), .ZN(n527) );
  INV_X1 U4052 ( .I(n42508), .ZN(n41276) );
  NAND2_X1 U4059 ( .A1(n53789), .A2(n53776), .ZN(n53047) );
  NOR2_X1 U4069 ( .A1(n39136), .A2(n39123), .ZN(n40957) );
  NAND2_X1 U4072 ( .A1(n53598), .A2(n53196), .ZN(n52843) );
  OAI21_X1 U4089 ( .A1(n55308), .A2(n54999), .B(n52118), .ZN(n25718) );
  NAND3_X1 U4095 ( .A1(n49108), .A2(n49109), .A3(n2514), .ZN(n22313) );
  NAND2_X1 U4097 ( .A1(n56174), .A2(n5193), .ZN(n17408) );
  OAI22_X1 U4100 ( .A1(n60105), .A2(n58763), .B1(n20630), .B2(n10869), .ZN(
        n53538) );
  NAND2_X1 U4101 ( .A1(n53535), .A2(n10869), .ZN(n17107) );
  AND2_X1 U4103 ( .A1(n22708), .A2(n10869), .Z(n1180) );
  INV_X2 U4108 ( .I(n57400), .ZN(n1477) );
  NAND2_X1 U4112 ( .A1(n54901), .A2(n2348), .ZN(n54928) );
  NAND3_X1 U4116 ( .A1(n54824), .A2(n5711), .A3(n1607), .ZN(n54336) );
  NOR2_X1 U4117 ( .A1(n41140), .A2(n43578), .ZN(n6971) );
  NOR2_X1 U4130 ( .A1(n15761), .A2(n54437), .ZN(n11463) );
  AOI21_X1 U4131 ( .A1(n56774), .A2(n56808), .B(n56785), .ZN(n13589) );
  AOI21_X1 U4139 ( .A1(n23595), .A2(n53080), .B(n53094), .ZN(n53058) );
  NAND3_X1 U4141 ( .A1(n54391), .A2(n54392), .A3(n54390), .ZN(n6557) );
  NAND3_X1 U4146 ( .A1(n47407), .A2(n18227), .A3(n47858), .ZN(n47867) );
  NOR3_X2 U4147 ( .A1(n17356), .A2(n17355), .A3(n17354), .ZN(n18251) );
  NOR3_X1 U4155 ( .A1(n53220), .A2(n57019), .A3(n57024), .ZN(n53221) );
  NAND2_X1 U4167 ( .A1(n1280), .A2(n54272), .ZN(n54209) );
  OAI21_X1 U4174 ( .A1(n39430), .A2(n6534), .B(n6533), .ZN(n6532) );
  AND2_X1 U4185 ( .A1(n15304), .A2(n52235), .Z(n1152) );
  BUF_X2 U4194 ( .I(n4336), .Z(n4152) );
  NAND2_X1 U4198 ( .A1(n1335), .A2(n43357), .ZN(n12196) );
  OAI22_X1 U4199 ( .A1(n14224), .A2(n55307), .B1(n55309), .B2(n55308), .ZN(
        n55315) );
  INV_X1 U4204 ( .I(n47798), .ZN(n8572) );
  NOR4_X1 U4206 ( .A1(n2531), .A2(n55175), .A3(n16978), .A4(n58813), .ZN(n2530) );
  INV_X4 U4216 ( .I(n8135), .ZN(n47208) );
  NAND2_X1 U4217 ( .A1(n20788), .A2(n48212), .ZN(n14690) );
  NOR2_X1 U4223 ( .A1(n34358), .A2(n34727), .ZN(n34250) );
  NAND2_X2 U4229 ( .A1(n20388), .A2(n20387), .ZN(n32318) );
  AOI21_X1 U4232 ( .A1(n56989), .A2(n52269), .B(n5081), .ZN(n52275) );
  NAND2_X1 U4235 ( .A1(n6061), .A2(n22669), .ZN(n53931) );
  NAND3_X1 U4240 ( .A1(n4830), .A2(n20891), .A3(n60553), .ZN(n55969) );
  NAND2_X1 U4241 ( .A1(n31270), .A2(n31264), .ZN(n31284) );
  OAI22_X1 U4242 ( .A1(n53924), .A2(n54001), .B1(n53902), .B2(n23292), .ZN(
        n21119) );
  NOR2_X1 U4243 ( .A1(n23292), .A2(n6061), .ZN(n53984) );
  NAND2_X1 U4244 ( .A1(n64970), .A2(n4830), .ZN(n55965) );
  OAI21_X1 U4245 ( .A1(n2719), .A2(n36584), .B(n36580), .ZN(n2715) );
  NOR2_X1 U4252 ( .A1(n1714), .A2(n61745), .ZN(n5949) );
  NOR3_X1 U4256 ( .A1(n1456), .A2(n12074), .A3(n1613), .ZN(n8744) );
  AND2_X1 U4257 ( .A1(n55337), .A2(n55345), .Z(n15864) );
  NAND2_X1 U4260 ( .A1(n12962), .A2(n61745), .ZN(n41579) );
  INV_X1 U4261 ( .I(n65022), .ZN(n10) );
  NAND2_X1 U4263 ( .A1(n53509), .A2(n53511), .ZN(n299) );
  NOR3_X2 U4265 ( .A1(n29388), .A2(n29390), .A3(n29389), .ZN(n29391) );
  NAND2_X1 U4267 ( .A1(n42676), .A2(n42838), .ZN(n41729) );
  OAI21_X1 U4273 ( .A1(n13072), .A2(n65275), .B(n1647), .ZN(n11809) );
  NAND2_X1 U4279 ( .A1(n5318), .A2(n13218), .ZN(n5056) );
  NOR2_X1 U4280 ( .A1(n53439), .A2(n53435), .ZN(n12785) );
  OAI22_X1 U4281 ( .A1(n53434), .A2(n53435), .B1(n53439), .B2(n3127), .ZN(
        n23507) );
  INV_X1 U4282 ( .I(n53439), .ZN(n53442) );
  INV_X1 U4298 ( .I(n14332), .ZN(n52237) );
  INV_X2 U4299 ( .I(n54411), .ZN(n1367) );
  INV_X1 U4326 ( .I(n53104), .ZN(n53105) );
  NOR2_X1 U4334 ( .A1(n1438), .A2(n14174), .ZN(n22156) );
  NAND2_X1 U4342 ( .A1(n56539), .A2(n52704), .ZN(n56532) );
  NOR2_X2 U4347 ( .A1(n22431), .A2(n61223), .ZN(n35182) );
  INV_X1 U4354 ( .I(n12049), .ZN(n10739) );
  NAND3_X1 U4357 ( .A1(n54346), .A2(n54348), .A3(n4564), .ZN(n6676) );
  NAND3_X1 U4358 ( .A1(n54345), .A2(n54348), .A3(n54344), .ZN(n6673) );
  CLKBUF_X2 U4364 ( .I(n41506), .Z(n4945) );
  NOR3_X1 U4370 ( .A1(n27678), .A2(n1889), .A3(n29695), .ZN(n27682) );
  INV_X1 U4372 ( .I(n1889), .ZN(n28186) );
  NOR2_X1 U4374 ( .A1(n27678), .A2(n1889), .ZN(n26910) );
  NAND2_X1 U4378 ( .A1(n30441), .A2(n24298), .ZN(n28095) );
  NAND3_X1 U4404 ( .A1(n47087), .A2(n5090), .A3(n14518), .ZN(n48466) );
  OAI21_X1 U4405 ( .A1(n5081), .A2(n52881), .B(n56985), .ZN(n52887) );
  NAND4_X1 U4427 ( .A1(n14438), .A2(n49859), .A3(n49864), .A4(n14436), .ZN(
        n14435) );
  INV_X1 U4428 ( .I(n39317), .ZN(n40294) );
  NAND2_X1 U4432 ( .A1(n12974), .A2(n55722), .ZN(n13025) );
  INV_X4 U4440 ( .I(n1270), .ZN(n42804) );
  NAND2_X2 U4446 ( .A1(n12116), .A2(n19231), .ZN(n35604) );
  NAND2_X1 U4461 ( .A1(n56117), .A2(n56120), .ZN(n7) );
  NOR3_X2 U4464 ( .A1(n25546), .A2(n25548), .A3(n25547), .ZN(n10631) );
  NAND2_X2 U4467 ( .A1(n9548), .A2(n20929), .ZN(n5124) );
  XOR2_X1 U4471 ( .A1(n14901), .A2(n10), .Z(n45425) );
  NAND2_X1 U4477 ( .A1(n35198), .A2(n9329), .ZN(n33324) );
  NOR2_X2 U4478 ( .A1(n22701), .A2(n35629), .ZN(n35198) );
  NAND2_X2 U4482 ( .A1(n1866), .A2(n29905), .ZN(n30857) );
  XOR2_X1 U4483 ( .A1(n61666), .A2(n16), .Z(n15746) );
  XOR2_X1 U4484 ( .A1(n45336), .A2(n25836), .Z(n16) );
  XOR2_X1 U4490 ( .A1(n17), .A2(n46126), .Z(n10116) );
  XOR2_X1 U4491 ( .A1(n46296), .A2(n46123), .Z(n17) );
  XOR2_X1 U4495 ( .A1(n51136), .A2(n50868), .Z(n9632) );
  XOR2_X1 U4498 ( .A1(n20072), .A2(n31342), .Z(n4692) );
  NOR2_X2 U4513 ( .A1(n21717), .A2(n22523), .ZN(n41037) );
  NOR2_X1 U4521 ( .A1(n53947), .A2(n12915), .ZN(n24) );
  XOR2_X1 U4527 ( .A1(n26), .A2(n25316), .Z(n8833) );
  XOR2_X1 U4528 ( .A1(n51050), .A2(n52025), .Z(n26) );
  XOR2_X1 U4529 ( .A1(n27), .A2(n22376), .Z(n43821) );
  INV_X1 U4534 ( .I(n35630), .ZN(n35632) );
  BUF_X2 U4535 ( .I(n15271), .Z(n3478) );
  NAND2_X2 U4555 ( .A1(n33642), .A2(n33117), .ZN(n4266) );
  INV_X2 U4562 ( .I(n3673), .ZN(n25519) );
  XOR2_X1 U4563 ( .A1(n10311), .A2(n39), .Z(n3673) );
  OR2_X1 U4570 ( .A1(n3077), .A2(n54079), .Z(n1148) );
  NAND3_X1 U4573 ( .A1(n59698), .A2(n47663), .A3(n15157), .ZN(n47666) );
  NAND2_X2 U4587 ( .A1(n3667), .A2(n40713), .ZN(n41454) );
  XOR2_X1 U4589 ( .A1(n33032), .A2(n46), .Z(n32488) );
  XOR2_X1 U4590 ( .A1(n33232), .A2(n32479), .Z(n46) );
  XOR2_X1 U4593 ( .A1(n48), .A2(n15462), .Z(n15459) );
  XOR2_X1 U4594 ( .A1(n51846), .A2(n15461), .Z(n48) );
  XOR2_X1 U4596 ( .A1(n49), .A2(n19514), .Z(n32657) );
  XOR2_X1 U4597 ( .A1(n32655), .A2(n33243), .Z(n49) );
  NAND2_X2 U4602 ( .A1(n17401), .A2(n17400), .ZN(n35662) );
  NAND2_X1 U4603 ( .A1(n50), .A2(n43951), .ZN(n11406) );
  NAND3_X2 U4605 ( .A1(n14968), .A2(n18515), .A3(n27442), .ZN(n29369) );
  XOR2_X1 U4618 ( .A1(n57), .A2(n57321), .Z(n12658) );
  XOR2_X1 U4621 ( .A1(n59), .A2(n61667), .Z(n2798) );
  XOR2_X1 U4622 ( .A1(n5027), .A2(n44587), .Z(n59) );
  XOR2_X1 U4624 ( .A1(n60), .A2(n51685), .Z(n6447) );
  XOR2_X1 U4627 ( .A1(n14251), .A2(n44849), .Z(n61) );
  NOR2_X2 U4637 ( .A1(n33103), .A2(n16856), .ZN(n33563) );
  NOR3_X2 U4640 ( .A1(n17788), .A2(n17789), .A3(n17790), .ZN(n67) );
  AND3_X1 U4647 ( .A1(n45501), .A2(n45500), .A3(n45499), .Z(n19686) );
  OAI22_X2 U4649 ( .A1(n36594), .A2(n36593), .B1(n36592), .B2(n36591), .ZN(
        n36602) );
  OAI22_X1 U4652 ( .A1(n56889), .A2(n56888), .B1(n60708), .B2(n56887), .ZN(
        n56900) );
  BUF_X4 U4658 ( .I(n22098), .Z(n19681) );
  INV_X4 U4660 ( .I(n24782), .ZN(n24007) );
  NAND2_X2 U4666 ( .A1(n43656), .A2(n6221), .ZN(n6995) );
  NOR3_X2 U4667 ( .A1(n9081), .A2(n7923), .A3(n7924), .ZN(n43656) );
  XOR2_X1 U4673 ( .A1(n8950), .A2(n33160), .Z(n79) );
  XOR2_X1 U4674 ( .A1(n80), .A2(n7698), .Z(n45341) );
  XOR2_X1 U4675 ( .A1(n10282), .A2(n44826), .Z(n80) );
  OAI21_X1 U4677 ( .A1(n41954), .A2(n41949), .B(n60143), .ZN(n41301) );
  NOR2_X2 U4678 ( .A1(n38273), .A2(n22290), .ZN(n41954) );
  NOR2_X2 U4679 ( .A1(n12912), .A2(n12914), .ZN(n81) );
  AOI22_X1 U4690 ( .A1(n48410), .A2(n62054), .B1(n12845), .B2(n12842), .ZN(
        n12841) );
  AOI22_X1 U4701 ( .A1(n55062), .A2(n55079), .B1(n55064), .B2(n55063), .ZN(n83) );
  XOR2_X1 U4705 ( .A1(n3914), .A2(n3913), .Z(n84) );
  OR2_X1 U4707 ( .A1(n11179), .A2(n61475), .Z(n42054) );
  XOR2_X1 U4708 ( .A1(n85), .A2(n3449), .Z(n20301) );
  XOR2_X1 U4709 ( .A1(n24449), .A2(n44293), .Z(n85) );
  AOI21_X1 U4710 ( .A1(n36820), .A2(n36819), .B(n15200), .ZN(n8098) );
  INV_X2 U4714 ( .I(n22523), .ZN(n1400) );
  NAND2_X1 U4719 ( .A1(n55972), .A2(n55975), .ZN(n55979) );
  NOR2_X2 U4720 ( .A1(n19461), .A2(n10525), .ZN(n30237) );
  AOI21_X2 U4728 ( .A1(n42117), .A2(n58210), .B(n1007), .ZN(n13926) );
  NAND2_X2 U4729 ( .A1(n27387), .A2(n28243), .ZN(n26268) );
  BUF_X2 U4749 ( .I(n15632), .Z(n101) );
  XOR2_X1 U4750 ( .A1(n63892), .A2(n887), .Z(n8423) );
  XOR2_X1 U4751 ( .A1(n23491), .A2(n32101), .Z(n887) );
  XOR2_X1 U4755 ( .A1(n38470), .A2(n37552), .Z(n103) );
  BUF_X2 U4757 ( .I(n38812), .Z(n23583) );
  NAND2_X2 U4759 ( .A1(n15156), .A2(n24837), .ZN(n26286) );
  XOR2_X1 U4760 ( .A1(n2147), .A2(n15087), .Z(n2842) );
  AND2_X1 U4771 ( .A1(n2124), .A2(n1226), .Z(n9198) );
  NAND2_X2 U4774 ( .A1(n25698), .A2(n12164), .ZN(n30254) );
  NOR2_X2 U4783 ( .A1(n54634), .A2(n54860), .ZN(n6580) );
  AND2_X1 U4788 ( .A1(n14530), .A2(n21792), .Z(n47247) );
  XOR2_X1 U4791 ( .A1(n106), .A2(n44626), .Z(n7140) );
  NAND2_X2 U4793 ( .A1(n12051), .A2(n10734), .ZN(n29490) );
  XOR2_X1 U4794 ( .A1(n107), .A2(n54870), .Z(Plaintext[84]) );
  XOR2_X1 U4798 ( .A1(n59218), .A2(n45423), .Z(n45003) );
  OR2_X2 U4803 ( .A1(n32400), .A2(n34359), .Z(n34725) );
  XOR2_X1 U4804 ( .A1(n9358), .A2(n9356), .Z(n32400) );
  NAND2_X2 U4805 ( .A1(n1356), .A2(n8113), .ZN(n29653) );
  BUF_X2 U4812 ( .I(n32513), .Z(n111) );
  XOR2_X1 U4815 ( .A1(n32524), .A2(n24434), .Z(n112) );
  XOR2_X1 U4818 ( .A1(n31827), .A2(n33906), .Z(n31828) );
  XOR2_X1 U4821 ( .A1(n115), .A2(n11102), .Z(n114) );
  INV_X2 U4822 ( .I(n49088), .ZN(n45389) );
  OAI21_X1 U4823 ( .A1(n28121), .A2(n29626), .B(n26948), .ZN(n26949) );
  NOR2_X2 U4827 ( .A1(n57198), .A2(n43464), .ZN(n43478) );
  NOR2_X2 U4841 ( .A1(n24199), .A2(n19590), .ZN(n31101) );
  NAND3_X2 U4843 ( .A1(n18232), .A2(n15802), .A3(n18237), .ZN(n32733) );
  INV_X2 U4851 ( .I(n22477), .ZN(n25428) );
  NOR2_X2 U4852 ( .A1(n3478), .A2(n21159), .ZN(n29063) );
  NOR2_X2 U4855 ( .A1(n1534), .A2(n34161), .ZN(n11874) );
  AOI21_X1 U4859 ( .A1(n26348), .A2(n26349), .B(n28346), .ZN(n26350) );
  BUF_X2 U4864 ( .I(n20882), .Z(n129) );
  XOR2_X1 U4867 ( .A1(n14900), .A2(n132), .Z(n45054) );
  XOR2_X1 U4868 ( .A1(n45326), .A2(n46620), .Z(n14900) );
  BUF_X2 U4871 ( .I(n23699), .Z(n22410) );
  NAND2_X1 U4872 ( .A1(n133), .A2(n22629), .ZN(n22628) );
  NOR2_X2 U4877 ( .A1(n1500), .A2(n4313), .ZN(n40886) );
  INV_X2 U4883 ( .I(n20634), .ZN(n5081) );
  XOR2_X1 U4894 ( .A1(n18478), .A2(n20593), .Z(n2000) );
  NAND2_X1 U4897 ( .A1(n56382), .A2(n137), .ZN(n21857) );
  NAND2_X2 U4916 ( .A1(n11942), .A2(n11949), .ZN(n13392) );
  INV_X4 U4921 ( .I(n21467), .ZN(n21468) );
  XOR2_X1 U4926 ( .A1(n144), .A2(n32028), .Z(n8264) );
  AND2_X1 U4935 ( .A1(n21067), .A2(n21279), .Z(n7574) );
  OAI21_X1 U4945 ( .A1(n7916), .A2(n29302), .B(n10324), .ZN(n7915) );
  AND2_X1 U4951 ( .A1(n22139), .A2(n14729), .Z(n29222) );
  NAND2_X1 U4957 ( .A1(n16810), .A2(n153), .ZN(n17306) );
  NAND2_X1 U4958 ( .A1(n27280), .A2(n28547), .ZN(n153) );
  BUF_X2 U4961 ( .I(n28552), .Z(n19328) );
  NAND2_X1 U4967 ( .A1(n7027), .A2(n53449), .ZN(n53450) );
  NAND2_X2 U4970 ( .A1(n32695), .A2(n33654), .ZN(n33391) );
  INV_X4 U4971 ( .I(n30441), .ZN(n24299) );
  NOR2_X2 U4980 ( .A1(n10699), .A2(n14954), .ZN(n34652) );
  NOR3_X2 U4982 ( .A1(n13983), .A2(n159), .A3(n1530), .ZN(n5185) );
  NOR2_X2 U4994 ( .A1(n10748), .A2(n26089), .ZN(n5008) );
  AND2_X1 U4995 ( .A1(n26450), .A2(n26449), .Z(n215) );
  XOR2_X1 U4997 ( .A1(n50529), .A2(n50530), .Z(n50531) );
  NOR2_X2 U5003 ( .A1(n23757), .A2(n22601), .ZN(n32900) );
  NAND2_X1 U5004 ( .A1(n6726), .A2(n367), .ZN(n856) );
  XNOR2_X1 U5026 ( .A1(n24757), .A2(n5778), .ZN(n1620) );
  NOR3_X1 U5032 ( .A1(n17726), .A2(n27117), .A3(n4488), .ZN(n17725) );
  INV_X4 U5033 ( .I(n25124), .ZN(n1781) );
  XOR2_X1 U5034 ( .A1(n169), .A2(n4273), .Z(n44509) );
  XOR2_X1 U5035 ( .A1(n44505), .A2(n25612), .Z(n169) );
  NOR3_X2 U5038 ( .A1(n171), .A2(n2446), .A3(n170), .ZN(n21212) );
  NOR2_X1 U5039 ( .A1(n2451), .A2(n42736), .ZN(n171) );
  NOR2_X2 U5041 ( .A1(n12979), .A2(n18736), .ZN(n29863) );
  OR2_X1 U5045 ( .A1(n15805), .A2(n35994), .Z(n37043) );
  INV_X4 U5048 ( .I(n1335), .ZN(n6426) );
  NOR2_X2 U5051 ( .A1(n40994), .A2(n40996), .ZN(n40211) );
  NOR4_X2 U5057 ( .A1(n14679), .A2(n26341), .A3(n27601), .A4(n26340), .ZN(
        n14678) );
  NAND2_X2 U5060 ( .A1(n24351), .A2(n36796), .ZN(n36812) );
  BUF_X2 U5061 ( .I(n25689), .Z(n178) );
  AOI22_X1 U5064 ( .A1(n38036), .A2(n38037), .B1(n40991), .B2(n40997), .ZN(
        n38038) );
  XOR2_X1 U5065 ( .A1(n31611), .A2(n31612), .Z(n31619) );
  XOR2_X1 U5066 ( .A1(n9040), .A2(n61497), .Z(n31611) );
  AND2_X1 U5073 ( .A1(n48802), .A2(n17087), .Z(n17086) );
  NAND2_X2 U5074 ( .A1(n6411), .A2(n16590), .ZN(n48802) );
  BUF_X2 U5079 ( .I(n28410), .Z(n180) );
  AOI22_X2 U5080 ( .A1(n36975), .A2(n37233), .B1(n37168), .B2(n37249), .ZN(
        n37451) );
  NAND2_X2 U5081 ( .A1(n9344), .A2(n28313), .ZN(n9251) );
  NAND4_X1 U5090 ( .A1(n61854), .A2(n574), .A3(n34132), .A4(n34144), .ZN(
        n32819) );
  INV_X2 U5110 ( .I(n1203), .ZN(n47180) );
  OAI21_X1 U5116 ( .A1(n288), .A2(n54444), .B(n54446), .ZN(n15026) );
  INV_X4 U5123 ( .I(n28588), .ZN(n29642) );
  NAND2_X1 U5126 ( .A1(n23474), .A2(n27483), .ZN(n15999) );
  NOR3_X1 U5128 ( .A1(n19197), .A2(n54312), .A3(n21296), .ZN(n26155) );
  BUF_X4 U5134 ( .I(Key[79]), .Z(n54708) );
  NAND3_X1 U5135 ( .A1(n54983), .A2(n55412), .A3(n54980), .ZN(n52908) );
  NOR2_X1 U5139 ( .A1(n19871), .A2(n27725), .ZN(n27730) );
  INV_X4 U5140 ( .I(n36338), .ZN(n20720) );
  NAND2_X2 U5143 ( .A1(n9200), .A2(n9185), .ZN(n42593) );
  OR2_X2 U5153 ( .A1(n41019), .A2(n14721), .Z(n40605) );
  NOR2_X2 U5154 ( .A1(n21516), .A2(n46558), .ZN(n5838) );
  AND2_X1 U5159 ( .A1(n56362), .A2(n56554), .Z(n21842) );
  OR2_X1 U5163 ( .A1(n46883), .A2(n9730), .Z(n22246) );
  NAND2_X1 U5170 ( .A1(n29550), .A2(n30786), .ZN(n202) );
  NOR2_X2 U5172 ( .A1(n35144), .A2(n8608), .ZN(n35977) );
  BUF_X2 U5173 ( .I(n38871), .Z(n204) );
  NAND4_X1 U5179 ( .A1(n6558), .A2(n11248), .A3(n6557), .A4(n11249), .ZN(n6556) );
  XOR2_X1 U5186 ( .A1(n208), .A2(n14432), .Z(n6063) );
  NAND2_X2 U5202 ( .A1(n32775), .A2(n21058), .ZN(n5233) );
  INV_X4 U5207 ( .I(n26092), .ZN(n24837) );
  NAND2_X2 U5212 ( .A1(n211), .A2(n28460), .ZN(n28441) );
  NOR3_X2 U5217 ( .A1(n5153), .A2(n29295), .A3(n25532), .ZN(n26959) );
  OAI21_X2 U5228 ( .A1(n45235), .A2(n45234), .B(n59966), .ZN(n25781) );
  NOR2_X1 U5233 ( .A1(n5145), .A2(n59695), .ZN(n5465) );
  XOR2_X1 U5237 ( .A1(n33866), .A2(n64968), .Z(n32676) );
  NAND3_X2 U5239 ( .A1(n20934), .A2(n36750), .A3(n36751), .ZN(n15578) );
  BUF_X2 U5258 ( .I(n31905), .Z(n21059) );
  NAND2_X2 U5266 ( .A1(n9200), .A2(n23003), .ZN(n13825) );
  NAND2_X2 U5268 ( .A1(n54195), .A2(n54196), .ZN(n54203) );
  NOR2_X2 U5269 ( .A1(n18859), .A2(n2984), .ZN(n54195) );
  NAND3_X2 U5285 ( .A1(n52728), .A2(n52727), .A3(n52726), .ZN(n19181) );
  XOR2_X1 U5289 ( .A1(n65273), .A2(n19984), .Z(n2289) );
  NAND2_X2 U5295 ( .A1(n12082), .A2(n25118), .ZN(n40469) );
  OAI22_X1 U5300 ( .A1(n33097), .A2(n16939), .B1(n32802), .B2(n33561), .ZN(
        n32530) );
  NAND2_X2 U5301 ( .A1(n42324), .A2(n23425), .ZN(n42317) );
  BUF_X4 U5305 ( .I(Key[84]), .Z(n54870) );
  BUF_X4 U5306 ( .I(n47911), .Z(n49538) );
  NOR3_X1 U5307 ( .A1(n35906), .A2(n60659), .A3(n35485), .ZN(n3103) );
  NAND2_X2 U5312 ( .A1(n15713), .A2(n57192), .ZN(n52845) );
  INV_X4 U5316 ( .I(n1445), .ZN(n29292) );
  OAI21_X1 U5320 ( .A1(n61683), .A2(n64978), .B(n53836), .ZN(n51858) );
  NAND3_X2 U5334 ( .A1(n3743), .A2(n911), .A3(n31359), .ZN(n37036) );
  XOR2_X1 U5336 ( .A1(n31479), .A2(n240), .Z(n20194) );
  XOR2_X1 U5337 ( .A1(n28796), .A2(n57227), .Z(n240) );
  XOR2_X1 U5345 ( .A1(n23804), .A2(n44817), .Z(n25694) );
  XOR2_X1 U5348 ( .A1(n10746), .A2(n1670), .Z(n45293) );
  INV_X2 U5350 ( .I(n38146), .ZN(n46683) );
  BUF_X4 U5352 ( .I(Key[160]), .Z(n56508) );
  NOR2_X2 U5357 ( .A1(n49363), .A2(n17558), .ZN(n52157) );
  INV_X2 U5360 ( .I(n14538), .ZN(n246) );
  NAND3_X2 U5362 ( .A1(n42607), .A2(n61372), .A3(n5126), .ZN(n42595) );
  AND2_X1 U5381 ( .A1(n33562), .A2(n33563), .Z(n33565) );
  AOI22_X1 U5383 ( .A1(n56197), .A2(n56198), .B1(n56195), .B2(n56196), .ZN(
        n56199) );
  XOR2_X1 U5386 ( .A1(n5449), .A2(n5448), .Z(n5451) );
  NAND2_X1 U5388 ( .A1(n6194), .A2(n45202), .ZN(n6188) );
  NOR2_X2 U5389 ( .A1(n6015), .A2(n49529), .ZN(n3472) );
  NOR2_X1 U5397 ( .A1(n9470), .A2(n9471), .ZN(n9469) );
  NAND2_X2 U5401 ( .A1(n2124), .A2(n40949), .ZN(n38049) );
  INV_X2 U5408 ( .I(n25659), .ZN(n33729) );
  XOR2_X1 U5412 ( .A1(n254), .A2(n15354), .Z(n4890) );
  XOR2_X1 U5414 ( .A1(n4055), .A2(n255), .Z(n4054) );
  XOR2_X1 U5415 ( .A1(n51120), .A2(n51126), .Z(n255) );
  NOR2_X2 U5416 ( .A1(n32885), .A2(n7323), .ZN(n34164) );
  NAND4_X1 U5427 ( .A1(n55048), .A2(n55047), .A3(n55065), .A4(n55046), .ZN(
        n55049) );
  INV_X2 U5429 ( .I(n31114), .ZN(n19697) );
  XOR2_X1 U5437 ( .A1(n5989), .A2(n46697), .Z(n8737) );
  NAND2_X2 U5443 ( .A1(n24250), .A2(n43225), .ZN(n43000) );
  NOR2_X1 U5446 ( .A1(n21837), .A2(n13143), .ZN(n21635) );
  BUF_X2 U5453 ( .I(n11977), .Z(n264) );
  AND3_X1 U5459 ( .A1(n2885), .A2(n12393), .A3(n57211), .Z(n19185) );
  NAND3_X1 U5460 ( .A1(n55104), .A2(n55103), .A3(n4416), .ZN(n392) );
  NOR3_X2 U5462 ( .A1(n14699), .A2(n42889), .A3(n61709), .ZN(n14698) );
  XOR2_X1 U5468 ( .A1(n269), .A2(n12020), .Z(n11985) );
  BUF_X4 U5472 ( .I(n18053), .Z(n4263) );
  BUF_X4 U5473 ( .I(n839), .Z(n10531) );
  AND2_X1 U5476 ( .A1(n33539), .A2(n14330), .Z(n21651) );
  AOI22_X2 U5477 ( .A1(n29382), .A2(n29383), .B1(n5659), .B2(n29381), .ZN(
        n29386) );
  NAND4_X2 U5478 ( .A1(n29387), .A2(n10603), .A3(n29386), .A4(n29385), .ZN(
        n29388) );
  XOR2_X1 U5482 ( .A1(n14945), .A2(n24212), .Z(n10864) );
  NOR2_X2 U5487 ( .A1(n13671), .A2(n22486), .ZN(n54929) );
  NAND2_X2 U5490 ( .A1(n24367), .A2(n15728), .ZN(n8212) );
  NAND2_X2 U5491 ( .A1(n13838), .A2(n1293), .ZN(n24367) );
  NAND2_X1 U5493 ( .A1(n274), .A2(n53971), .ZN(n53935) );
  OAI21_X1 U5494 ( .A1(n53933), .A2(n54006), .B(n53932), .ZN(n274) );
  XOR2_X1 U5502 ( .A1(n275), .A2(n54936), .Z(Plaintext[89]) );
  NAND2_X1 U5507 ( .A1(n27016), .A2(n29113), .ZN(n8806) );
  INV_X4 U5508 ( .I(n23209), .ZN(n27138) );
  BUF_X2 U5511 ( .I(n41430), .Z(n277) );
  BUF_X2 U5514 ( .I(n43915), .Z(n279) );
  XOR2_X1 U5517 ( .A1(n63263), .A2(n8550), .Z(n8551) );
  INV_X2 U5519 ( .I(n281), .ZN(n54459) );
  NOR2_X2 U5520 ( .A1(n55017), .A2(n12127), .ZN(n281) );
  NOR3_X1 U5523 ( .A1(n29298), .A2(n283), .A3(n282), .ZN(n29301) );
  NOR2_X1 U5524 ( .A1(n29296), .A2(n29295), .ZN(n282) );
  NOR2_X1 U5525 ( .A1(n29294), .A2(n29293), .ZN(n283) );
  XOR2_X1 U5526 ( .A1(n43786), .A2(n43782), .Z(n284) );
  NOR2_X2 U5527 ( .A1(n33004), .A2(n32457), .ZN(n20068) );
  NOR2_X2 U5534 ( .A1(n22071), .A2(n54813), .ZN(n5318) );
  AND3_X1 U5537 ( .A1(n42638), .A2(n20888), .A3(n43184), .Z(n19421) );
  XOR2_X1 U5540 ( .A1(n52373), .A2(n51319), .Z(n52629) );
  NAND2_X2 U5541 ( .A1(n8675), .A2(n24566), .ZN(n52373) );
  OR2_X1 U5542 ( .A1(n11463), .A2(n54827), .Z(n288) );
  NOR2_X1 U5547 ( .A1(n5114), .A2(n5113), .ZN(n5112) );
  XOR2_X1 U5553 ( .A1(n24621), .A2(n24040), .Z(n1998) );
  XOR2_X1 U5555 ( .A1(n5676), .A2(n53705), .Z(n292) );
  BUF_X2 U5559 ( .I(n1447), .Z(n296) );
  INV_X2 U5562 ( .I(n34019), .ZN(n1538) );
  XOR2_X1 U5565 ( .A1(n25136), .A2(n18830), .Z(n298) );
  NAND4_X2 U5566 ( .A1(n29263), .A2(n29265), .A3(n29573), .A4(n29264), .ZN(
        n29271) );
  NOR2_X1 U5571 ( .A1(n300), .A2(n299), .ZN(n23639) );
  INV_X1 U5572 ( .I(n53510), .ZN(n300) );
  NOR2_X1 U5575 ( .A1(n14322), .A2(n13426), .ZN(n13425) );
  XOR2_X1 U5584 ( .A1(n33044), .A2(n29259), .Z(n304) );
  NAND3_X1 U5585 ( .A1(n20319), .A2(n1457), .A3(n6351), .ZN(n17106) );
  NAND2_X2 U5586 ( .A1(n23857), .A2(n20349), .ZN(n20319) );
  XOR2_X1 U5587 ( .A1(n2345), .A2(n305), .Z(n21356) );
  XOR2_X1 U5590 ( .A1(n18547), .A2(n15726), .Z(n10884) );
  OAI22_X1 U5599 ( .A1(n22818), .A2(n21390), .B1(n55160), .B2(n55161), .ZN(
        n55174) );
  INV_X4 U5600 ( .I(n15806), .ZN(n47244) );
  XOR2_X1 U5609 ( .A1(n309), .A2(n9194), .Z(n9193) );
  XOR2_X1 U5610 ( .A1(n10896), .A2(n12869), .Z(n309) );
  INV_X1 U5615 ( .I(n23941), .ZN(n55475) );
  NAND2_X2 U5619 ( .A1(n5192), .A2(n30492), .ZN(n6714) );
  NOR3_X2 U5621 ( .A1(n21111), .A2(n21110), .A3(n21109), .ZN(n21108) );
  INV_X2 U5623 ( .I(n312), .ZN(n19609) );
  XOR2_X1 U5625 ( .A1(Ciphertext[175]), .A2(Key[158]), .Z(n23699) );
  OAI21_X1 U5628 ( .A1(n26723), .A2(n26724), .B(n313), .ZN(n26725) );
  NOR2_X1 U5629 ( .A1(n18200), .A2(n16654), .ZN(n313) );
  NAND2_X1 U5631 ( .A1(n11048), .A2(n42431), .ZN(n314) );
  INV_X2 U5634 ( .I(n315), .ZN(n18231) );
  XOR2_X1 U5636 ( .A1(n3753), .A2(n915), .Z(n3751) );
  XOR2_X1 U5637 ( .A1(n3752), .A2(n13115), .Z(n3753) );
  BUF_X4 U5643 ( .I(n36022), .Z(n23626) );
  AOI21_X1 U5652 ( .A1(n53418), .A2(n53419), .B(n53417), .ZN(n53424) );
  NOR2_X1 U5655 ( .A1(n21922), .A2(n25789), .ZN(n16716) );
  NAND2_X2 U5656 ( .A1(n7020), .A2(n53462), .ZN(n21922) );
  NAND2_X2 U5657 ( .A1(n3732), .A2(n14473), .ZN(n47361) );
  AOI21_X1 U5659 ( .A1(n1809), .A2(n33953), .B(n322), .ZN(n21259) );
  AND2_X1 U5661 ( .A1(n46790), .A2(n23185), .Z(n323) );
  OAI22_X2 U5668 ( .A1(n20491), .A2(n31263), .B1(n59755), .B2(n31262), .ZN(
        n31265) );
  NOR2_X1 U5675 ( .A1(n6313), .A2(n5945), .ZN(n5946) );
  AOI22_X1 U5678 ( .A1(n56989), .A2(n56993), .B1(n56612), .B2(n51437), .ZN(
        n51438) );
  NAND2_X2 U5688 ( .A1(n18609), .A2(n1384), .ZN(n48716) );
  NAND3_X2 U5690 ( .A1(n49533), .A2(n49532), .A3(n9983), .ZN(n48904) );
  OAI21_X1 U5692 ( .A1(n40712), .A2(n64366), .B(n333), .ZN(n40714) );
  AOI22_X1 U5693 ( .A1(n3042), .A2(n20994), .B1(n4819), .B2(n41453), .ZN(n333)
         );
  NOR2_X2 U5705 ( .A1(n21033), .A2(n24988), .ZN(n24501) );
  XOR2_X1 U5720 ( .A1(n345), .A2(n26467), .Z(n27433) );
  XOR2_X1 U5721 ( .A1(n56030), .A2(n4921), .Z(n345) );
  NOR2_X2 U5744 ( .A1(n5153), .A2(n26446), .ZN(n29306) );
  XOR2_X1 U5751 ( .A1(n349), .A2(n13642), .Z(n13640) );
  NAND2_X1 U5757 ( .A1(n10741), .A2(n9198), .ZN(n351) );
  AOI21_X1 U5758 ( .A1(n46094), .A2(n48601), .B(n352), .ZN(n46100) );
  NAND2_X2 U5763 ( .A1(n28594), .A2(n28593), .ZN(n29639) );
  XOR2_X1 U5764 ( .A1(n22919), .A2(n26850), .Z(n28594) );
  INV_X2 U5765 ( .I(n353), .ZN(n2614) );
  BUF_X2 U5767 ( .I(n15487), .Z(n354) );
  NOR3_X2 U5770 ( .A1(n356), .A2(n13806), .A3(n13803), .ZN(n14522) );
  INV_X4 U5772 ( .I(n56268), .ZN(n55659) );
  XOR2_X1 U5786 ( .A1(n24858), .A2(n12122), .Z(n365) );
  OAI22_X1 U5791 ( .A1(n35707), .A2(n24089), .B1(n35708), .B2(n1343), .ZN(
        n35721) );
  NOR2_X2 U5794 ( .A1(n36979), .A2(n23742), .ZN(n36610) );
  NAND2_X2 U5801 ( .A1(n3772), .A2(n22756), .ZN(n49451) );
  INV_X2 U5804 ( .I(n367), .ZN(n6727) );
  XOR2_X1 U5805 ( .A1(Ciphertext[177]), .A2(Key[172]), .Z(n367) );
  BUF_X4 U5808 ( .I(n12110), .Z(n10829) );
  INV_X2 U5809 ( .I(n33650), .ZN(n33649) );
  NAND3_X1 U5814 ( .A1(n47906), .A2(n7298), .A3(n61628), .ZN(n45587) );
  INV_X2 U5815 ( .I(n47905), .ZN(n7298) );
  NAND2_X2 U5816 ( .A1(n47570), .A2(n47901), .ZN(n47905) );
  XOR2_X1 U5829 ( .A1(n39247), .A2(n8720), .Z(n8719) );
  XOR2_X1 U5833 ( .A1(n46581), .A2(n1036), .Z(n6057) );
  BUF_X4 U5838 ( .I(Key[175]), .Z(n56849) );
  NAND3_X1 U5843 ( .A1(n56379), .A2(n56547), .A3(n56545), .ZN(n375) );
  NAND2_X2 U5844 ( .A1(n34490), .A2(n35883), .ZN(n35171) );
  NOR2_X2 U5849 ( .A1(n30159), .A2(n25157), .ZN(n17872) );
  NOR2_X2 U5850 ( .A1(n27334), .A2(n27335), .ZN(n30159) );
  NAND2_X2 U5858 ( .A1(n57537), .A2(n29053), .ZN(n30046) );
  AOI22_X1 U5859 ( .A1(n39962), .A2(n39961), .B1(n1272), .B2(n12615), .ZN(
        n39966) );
  OAI22_X1 U5861 ( .A1(n45926), .A2(n45925), .B1(n45924), .B2(n24374), .ZN(
        n381) );
  OAI22_X1 U5862 ( .A1(n382), .A2(n56937), .B1(n56939), .B2(n56963), .ZN(
        n56948) );
  XOR2_X1 U5864 ( .A1(n9005), .A2(n11575), .Z(n383) );
  INV_X2 U5866 ( .I(n21665), .ZN(n43288) );
  NAND4_X2 U5867 ( .A1(n18526), .A2(n23550), .A3(n25626), .A4(n39322), .ZN(
        n21665) );
  NOR2_X2 U5871 ( .A1(n22220), .A2(n28028), .ZN(n28079) );
  XOR2_X1 U5875 ( .A1(n386), .A2(n15862), .Z(n10859) );
  XOR2_X1 U5876 ( .A1(n387), .A2(n20223), .Z(n386) );
  NOR2_X2 U5880 ( .A1(n18909), .A2(n18907), .ZN(n33388) );
  NOR2_X2 U5882 ( .A1(n7972), .A2(n18600), .ZN(n50002) );
  NAND2_X1 U5885 ( .A1(n40226), .A2(n40140), .ZN(n25627) );
  INV_X4 U5896 ( .I(n27966), .ZN(n18423) );
  BUF_X2 U5901 ( .I(n22741), .Z(n15649) );
  NOR2_X1 U5902 ( .A1(n6660), .A2(n6661), .ZN(n6659) );
  INV_X2 U5922 ( .I(n399), .ZN(n6129) );
  NAND2_X2 U5924 ( .A1(n41340), .A2(n41559), .ZN(n43252) );
  XOR2_X1 U5926 ( .A1(n39369), .A2(n37102), .Z(n25641) );
  XOR2_X1 U5929 ( .A1(n31754), .A2(n61883), .Z(n400) );
  NAND2_X2 U5933 ( .A1(n2009), .A2(n17962), .ZN(n20758) );
  OAI21_X1 U5934 ( .A1(n25469), .A2(n59199), .B(n62921), .ZN(n404) );
  NOR2_X2 U5943 ( .A1(n42643), .A2(n16568), .ZN(n20208) );
  NOR2_X1 U5948 ( .A1(n49793), .A2(n23802), .ZN(n49796) );
  NAND2_X2 U5949 ( .A1(n49114), .A2(n1642), .ZN(n49793) );
  NOR2_X1 U5952 ( .A1(n408), .A2(n20264), .ZN(n20263) );
  NOR2_X1 U5953 ( .A1(n19855), .A2(n19856), .ZN(n408) );
  NAND2_X2 U5954 ( .A1(n409), .A2(n49645), .ZN(n11215) );
  NOR2_X2 U5971 ( .A1(n53867), .A2(n52783), .ZN(n4118) );
  XOR2_X1 U5974 ( .A1(n416), .A2(n2565), .Z(n517) );
  XOR2_X1 U5980 ( .A1(n25686), .A2(n8187), .Z(n20854) );
  XOR2_X1 U5981 ( .A1(n419), .A2(n43941), .Z(n8187) );
  INV_X1 U5984 ( .I(n49132), .ZN(n24135) );
  OR3_X1 U5985 ( .A1(n49132), .A2(n50360), .A3(n60209), .Z(n49205) );
  NAND2_X2 U5990 ( .A1(n22273), .A2(n27429), .ZN(n26470) );
  INV_X4 U5992 ( .I(n41568), .ZN(n24715) );
  NOR2_X1 U5994 ( .A1(n14614), .A2(n34657), .ZN(n14613) );
  XOR2_X1 U6002 ( .A1(n1672), .A2(n12265), .Z(n11736) );
  NOR3_X2 U6004 ( .A1(n424), .A2(n4903), .A3(n423), .ZN(n15247) );
  NOR2_X1 U6005 ( .A1(n35440), .A2(n1530), .ZN(n423) );
  NAND2_X1 U6009 ( .A1(n41543), .A2(n41544), .ZN(n426) );
  BUF_X2 U6018 ( .I(n42598), .Z(n429) );
  NAND2_X1 U6021 ( .A1(n22995), .A2(n22996), .ZN(n40048) );
  OR2_X2 U6022 ( .A1(n14354), .A2(n54272), .Z(n54285) );
  NOR2_X1 U6023 ( .A1(n432), .A2(n431), .ZN(n873) );
  NOR3_X2 U6025 ( .A1(n1890), .A2(n22159), .A3(n20734), .ZN(n28005) );
  NAND3_X1 U6026 ( .A1(n41944), .A2(n20227), .A3(n60021), .ZN(n41304) );
  XOR2_X1 U6028 ( .A1(n16691), .A2(n16508), .Z(n11471) );
  BUF_X2 U6029 ( .I(n29644), .Z(n434) );
  OR2_X1 U6031 ( .A1(n43656), .A2(n6221), .Z(n20685) );
  BUF_X2 U6040 ( .I(n22082), .Z(n436) );
  NOR2_X2 U6043 ( .A1(n34771), .A2(n60416), .ZN(n32946) );
  NOR2_X2 U6046 ( .A1(n24039), .A2(n24701), .ZN(n25993) );
  XOR2_X1 U6049 ( .A1(n439), .A2(n23267), .Z(n46576) );
  XOR2_X1 U6050 ( .A1(n46573), .A2(n46572), .Z(n439) );
  NAND2_X1 U6056 ( .A1(n20979), .A2(n49118), .ZN(n49119) );
  XOR2_X1 U6061 ( .A1(n442), .A2(n61654), .Z(n12887) );
  XOR2_X1 U6062 ( .A1(n12889), .A2(n23356), .Z(n442) );
  NOR2_X2 U6068 ( .A1(n28049), .A2(n15156), .ZN(n27126) );
  NAND3_X2 U6071 ( .A1(n35270), .A2(n36824), .A3(n35269), .ZN(n23782) );
  INV_X2 U6075 ( .I(n30705), .ZN(n13531) );
  AND2_X1 U6083 ( .A1(n40559), .A2(n42247), .Z(n449) );
  INV_X4 U6089 ( .I(n28633), .ZN(n28472) );
  XOR2_X1 U6094 ( .A1(n454), .A2(n3449), .Z(n9009) );
  NAND2_X2 U6096 ( .A1(n60054), .A2(n21906), .ZN(n34680) );
  NAND2_X2 U6110 ( .A1(n21605), .A2(n36796), .ZN(n36301) );
  INV_X4 U6111 ( .I(n27690), .ZN(n28471) );
  NAND3_X2 U6115 ( .A1(n16726), .A2(n16723), .A3(n34332), .ZN(n16722) );
  BUF_X2 U6127 ( .I(n9411), .Z(n463) );
  NAND2_X2 U6128 ( .A1(n11987), .A2(n60284), .ZN(n28904) );
  NOR2_X2 U6131 ( .A1(n3993), .A2(n2795), .ZN(n2794) );
  XOR2_X1 U6137 ( .A1(n46657), .A2(n46232), .Z(n7069) );
  XOR2_X1 U6138 ( .A1(n24733), .A2(n19268), .Z(n46657) );
  AND3_X1 U6145 ( .A1(n27289), .A2(n27288), .A3(n13761), .Z(n9583) );
  NOR2_X2 U6147 ( .A1(n34614), .A2(n34613), .ZN(n24273) );
  OAI21_X2 U6155 ( .A1(n4628), .A2(n4627), .B(n34604), .ZN(n31535) );
  NOR2_X2 U6159 ( .A1(n15666), .A2(n1267), .ZN(n46916) );
  NAND2_X2 U6162 ( .A1(n13084), .A2(n13083), .ZN(n31193) );
  BUF_X4 U6172 ( .I(n36567), .Z(n24102) );
  XOR2_X1 U6175 ( .A1(n11499), .A2(n478), .Z(n9770) );
  XOR2_X1 U6176 ( .A1(n46666), .A2(n61669), .Z(n478) );
  XOR2_X1 U6177 ( .A1(n32642), .A2(n54143), .Z(n33048) );
  NAND3_X2 U6178 ( .A1(n29420), .A2(n18160), .A3(n18159), .ZN(n32642) );
  XOR2_X1 U6182 ( .A1(n482), .A2(n22219), .Z(n15847) );
  XOR2_X1 U6183 ( .A1(n50541), .A2(n50540), .Z(n482) );
  XOR2_X1 U6184 ( .A1(n30974), .A2(n483), .Z(n31199) );
  XOR2_X1 U6185 ( .A1(n8590), .A2(n13990), .Z(n483) );
  NAND2_X1 U6189 ( .A1(n20870), .A2(n53403), .ZN(n486) );
  XOR2_X1 U6190 ( .A1(n32642), .A2(n19285), .Z(n13638) );
  NOR2_X2 U6192 ( .A1(n43851), .A2(n23730), .ZN(n22109) );
  NOR3_X2 U6194 ( .A1(n490), .A2(n34379), .A3(n489), .ZN(n34380) );
  NOR2_X1 U6195 ( .A1(n60980), .A2(n37365), .ZN(n489) );
  OR2_X2 U6196 ( .A1(n25598), .A2(n48074), .Z(n11246) );
  NAND2_X2 U6197 ( .A1(n60929), .A2(n13984), .ZN(n9144) );
  NAND2_X2 U6201 ( .A1(n15184), .A2(n32922), .ZN(n34720) );
  NOR2_X1 U6206 ( .A1(n63799), .A2(n910), .ZN(n34225) );
  NAND2_X2 U6208 ( .A1(n4186), .A2(n27414), .ZN(n18375) );
  AOI21_X2 U6209 ( .A1(n37895), .A2(n41912), .B(n42242), .ZN(n40788) );
  NOR2_X1 U6211 ( .A1(n48329), .A2(n2758), .ZN(n2076) );
  BUF_X4 U6215 ( .I(n26670), .Z(n22273) );
  NOR3_X2 U6224 ( .A1(n61844), .A2(n17338), .A3(n17337), .ZN(n17625) );
  NAND4_X1 U6228 ( .A1(n48799), .A2(n47990), .A3(n46965), .A4(n48802), .ZN(
        n499) );
  NOR3_X2 U6240 ( .A1(n18372), .A2(n49569), .A3(n18371), .ZN(n17969) );
  NOR2_X2 U6243 ( .A1(n30058), .A2(n27363), .ZN(n10023) );
  INV_X2 U6245 ( .I(n36434), .ZN(n36437) );
  NAND2_X2 U6246 ( .A1(n1742), .A2(n7237), .ZN(n12152) );
  INV_X2 U6248 ( .I(n9885), .ZN(n6781) );
  NAND2_X2 U6251 ( .A1(n47406), .A2(n47857), .ZN(n10947) );
  AOI21_X2 U6256 ( .A1(n19221), .A2(n5960), .B(n5958), .ZN(n14283) );
  NAND4_X2 U6259 ( .A1(n3407), .A2(n29140), .A3(n3406), .A4(n3405), .ZN(n3404)
         );
  INV_X2 U6262 ( .I(n506), .ZN(n51945) );
  XNOR2_X1 U6263 ( .A1(n50948), .A2(n52358), .ZN(n506) );
  OR2_X2 U6271 ( .A1(n2922), .A2(n2923), .Z(n11182) );
  XOR2_X1 U6272 ( .A1(n23040), .A2(n3863), .Z(n51952) );
  XOR2_X1 U6275 ( .A1(n31884), .A2(n876), .Z(n2991) );
  XOR2_X1 U6276 ( .A1(n31480), .A2(n13367), .Z(n13366) );
  NOR2_X2 U6278 ( .A1(n28746), .A2(n28745), .ZN(n29102) );
  AOI21_X2 U6291 ( .A1(n52863), .A2(n507), .B(n57060), .ZN(n52662) );
  AND2_X1 U6295 ( .A1(n5889), .A2(n56234), .Z(n5887) );
  XOR2_X1 U6304 ( .A1(n15711), .A2(n21098), .Z(n37894) );
  OR2_X2 U6323 ( .A1(n35292), .A2(n523), .Z(n2900) );
  OAI22_X1 U6324 ( .A1(n35284), .A2(n35699), .B1(n35285), .B2(n904), .ZN(n523)
         );
  INV_X2 U6325 ( .I(n25037), .ZN(n32199) );
  NAND3_X2 U6326 ( .A1(n25035), .A2(n25038), .A3(n30624), .ZN(n25037) );
  NOR2_X1 U6333 ( .A1(n527), .A2(n55244), .ZN(n7408) );
  INV_X2 U6348 ( .I(n532), .ZN(n2766) );
  XOR2_X1 U6349 ( .A1(n2769), .A2(n44931), .Z(n532) );
  NOR2_X2 U6350 ( .A1(n1416), .A2(n21921), .ZN(n37393) );
  XOR2_X1 U6356 ( .A1(n38526), .A2(n12356), .Z(n5660) );
  BUF_X2 U6363 ( .I(n52568), .Z(n535) );
  NAND2_X2 U6370 ( .A1(n9675), .A2(n1781), .ZN(n35440) );
  AND2_X1 U6371 ( .A1(n54254), .A2(n14354), .Z(n15923) );
  BUF_X2 U6374 ( .I(n5944), .Z(n540) );
  INV_X2 U6379 ( .I(n21014), .ZN(n2351) );
  NOR2_X2 U6381 ( .A1(n543), .A2(n8311), .ZN(n7767) );
  BUF_X2 U6384 ( .I(n32527), .Z(n33697) );
  OR2_X2 U6389 ( .A1(n41568), .A2(n41699), .Z(n16204) );
  NOR2_X2 U6397 ( .A1(n18975), .A2(n24394), .ZN(n48273) );
  XOR2_X1 U6400 ( .A1(n17766), .A2(n61655), .Z(n14638) );
  OR2_X1 U6401 ( .A1(n63085), .A2(n33613), .Z(n7120) );
  XOR2_X1 U6425 ( .A1(n2425), .A2(n1680), .Z(n3036) );
  XOR2_X1 U6426 ( .A1(n49961), .A2(n49960), .Z(n49962) );
  NAND2_X1 U6429 ( .A1(n31834), .A2(n16481), .ZN(n559) );
  NAND2_X2 U6433 ( .A1(n15689), .A2(n1562), .ZN(n13817) );
  XOR2_X1 U6434 ( .A1(n37625), .A2(n57221), .Z(n39688) );
  NOR2_X2 U6435 ( .A1(n14683), .A2(n14684), .ZN(n37625) );
  XOR2_X1 U6436 ( .A1(n9811), .A2(n562), .Z(n39694) );
  XOR2_X1 U6437 ( .A1(n39692), .A2(n39691), .Z(n562) );
  NAND2_X2 U6440 ( .A1(n43249), .A2(n43248), .ZN(n12262) );
  XOR2_X1 U6443 ( .A1(n1327), .A2(n1473), .Z(n565) );
  XOR2_X1 U6447 ( .A1(n23655), .A2(n567), .Z(n37865) );
  XOR2_X1 U6448 ( .A1(n38972), .A2(n49426), .Z(n567) );
  XOR2_X1 U6452 ( .A1(n569), .A2(n52900), .Z(Plaintext[0]) );
  NAND2_X2 U6456 ( .A1(n10251), .A2(n157), .ZN(n33650) );
  NAND2_X1 U6462 ( .A1(n5620), .A2(n52880), .ZN(n5619) );
  NAND2_X1 U6463 ( .A1(n33649), .A2(n12768), .ZN(n574) );
  INV_X1 U6470 ( .I(n19080), .ZN(n53080) );
  AND2_X1 U6471 ( .A1(n52878), .A2(n19080), .Z(n52879) );
  AOI21_X1 U6477 ( .A1(n27355), .A2(n65186), .B(n16218), .ZN(n19920) );
  BUF_X2 U6478 ( .I(n30159), .Z(n579) );
  XOR2_X1 U6480 ( .A1(n580), .A2(n50599), .Z(n3866) );
  XOR2_X1 U6481 ( .A1(n22256), .A2(n51522), .Z(n580) );
  XOR2_X1 U6486 ( .A1(n3477), .A2(n3259), .Z(n3258) );
  XOR2_X1 U6487 ( .A1(n2897), .A2(n3353), .Z(n3477) );
  XOR2_X1 U6490 ( .A1(n582), .A2(n9707), .Z(n15687) );
  XOR2_X1 U6491 ( .A1(n2391), .A2(n32715), .Z(n582) );
  XOR2_X1 U6497 ( .A1(n50952), .A2(n2070), .Z(n10497) );
  NOR2_X2 U6505 ( .A1(n23955), .A2(n20747), .ZN(n14350) );
  NAND4_X1 U6510 ( .A1(n55039), .A2(n55038), .A3(n55037), .A4(n55064), .ZN(
        n23688) );
  NOR3_X2 U6514 ( .A1(n26396), .A2(n26395), .A3(n26394), .ZN(n26403) );
  XOR2_X1 U6516 ( .A1(n36104), .A2(n21366), .Z(n590) );
  BUF_X2 U6518 ( .I(n22362), .Z(n591) );
  BUF_X4 U6526 ( .I(Key[130]), .Z(n55810) );
  INV_X2 U6527 ( .I(n14007), .ZN(n15474) );
  NAND2_X2 U6528 ( .A1(n4526), .A2(n49005), .ZN(n14007) );
  XOR2_X1 U6530 ( .A1(n44143), .A2(n1052), .Z(n6056) );
  NAND4_X1 U6534 ( .A1(n34810), .A2(n34811), .A3(n35946), .A4(n34817), .ZN(
        n595) );
  OR2_X1 U6536 ( .A1(n56257), .A2(n51888), .Z(n19905) );
  OAI22_X1 U6544 ( .A1(n5594), .A2(n596), .B1(n31080), .B2(n31079), .ZN(n14422) );
  BUF_X2 U6545 ( .I(n3617), .Z(n597) );
  NAND2_X2 U6548 ( .A1(n27352), .A2(n27353), .ZN(n31055) );
  AOI21_X2 U6550 ( .A1(n52252), .A2(n52251), .B(n52250), .ZN(n52261) );
  NOR2_X2 U6557 ( .A1(n35505), .A2(n14753), .ZN(n36922) );
  BUF_X2 U6560 ( .I(n33258), .Z(n602) );
  AND2_X1 U6565 ( .A1(n56962), .A2(n25022), .Z(n16168) );
  AOI21_X1 U6566 ( .A1(n55076), .A2(n55089), .B(n55056), .ZN(n55032) );
  NAND2_X2 U6568 ( .A1(n55088), .A2(n25171), .ZN(n9102) );
  XOR2_X1 U6570 ( .A1(n2191), .A2(n39628), .Z(n604) );
  XOR2_X1 U6571 ( .A1(n605), .A2(n46636), .Z(n6098) );
  INV_X2 U6580 ( .I(n609), .ZN(n26126) );
  XOR2_X1 U6581 ( .A1(Key[121]), .A2(Ciphertext[156]), .Z(n609) );
  NAND2_X2 U6583 ( .A1(n29315), .A2(n29314), .ZN(n24088) );
  XOR2_X1 U6586 ( .A1(n610), .A2(n53308), .Z(Plaintext[17]) );
  NAND4_X2 U6588 ( .A1(n611), .A2(n39891), .A3(n39890), .A4(n39893), .ZN(
        n39897) );
  OAI21_X2 U6589 ( .A1(n57327), .A2(n39888), .B(n40093), .ZN(n611) );
  NOR3_X2 U6590 ( .A1(n12783), .A2(n12782), .A3(n12785), .ZN(n7228) );
  NOR2_X2 U6595 ( .A1(n57039), .A2(n52786), .ZN(n53436) );
  NOR2_X2 U6598 ( .A1(n60417), .A2(n17967), .ZN(n47858) );
  XOR2_X1 U6600 ( .A1(n616), .A2(n836), .Z(n29311) );
  XOR2_X1 U6601 ( .A1(n52317), .A2(n53833), .Z(n616) );
  NAND3_X2 U6603 ( .A1(n43834), .A2(n43833), .A3(n9726), .ZN(n618) );
  BUF_X2 U6605 ( .I(n56155), .Z(n620) );
  NOR3_X1 U6609 ( .A1(n36703), .A2(n623), .A3(n622), .ZN(n36715) );
  INV_X2 U6614 ( .I(n56482), .ZN(n19731) );
  NAND2_X2 U6615 ( .A1(n9311), .A2(n17795), .ZN(n56482) );
  XOR2_X1 U6622 ( .A1(n24145), .A2(n25822), .Z(n31773) );
  NOR3_X2 U6623 ( .A1(n56380), .A2(n56383), .A3(n56387), .ZN(n624) );
  INV_X2 U6625 ( .I(n28318), .ZN(n28051) );
  XOR2_X1 U6627 ( .A1(n38158), .A2(n4922), .Z(n625) );
  NAND3_X2 U6631 ( .A1(n4396), .A2(n52710), .A3(n52709), .ZN(n627) );
  AND2_X1 U6633 ( .A1(n13489), .A2(n14943), .Z(n7260) );
  XOR2_X1 U6634 ( .A1(n12129), .A2(n628), .Z(n11508) );
  XOR2_X1 U6635 ( .A1(n630), .A2(n61671), .Z(n2025) );
  NOR2_X1 U6644 ( .A1(n14422), .A2(n14421), .ZN(n4973) );
  INV_X2 U6646 ( .I(n43513), .ZN(n13678) );
  NAND2_X2 U6648 ( .A1(n15498), .A2(n57075), .ZN(n18219) );
  OR2_X1 U6655 ( .A1(n34117), .A2(n2695), .Z(n2562) );
  XOR2_X1 U6658 ( .A1(n10409), .A2(n21006), .Z(n9714) );
  NAND2_X2 U6661 ( .A1(n5179), .A2(n1352), .ZN(n5688) );
  INV_X2 U6662 ( .I(n602), .ZN(n31486) );
  XOR2_X1 U6663 ( .A1(n638), .A2(n18013), .Z(n35025) );
  NAND2_X2 U6668 ( .A1(n57211), .A2(n24864), .ZN(n35398) );
  NOR2_X2 U6669 ( .A1(n4789), .A2(n43155), .ZN(n43170) );
  XOR2_X1 U6670 ( .A1(Ciphertext[83]), .A2(Key[90]), .Z(n6886) );
  NAND4_X1 U6671 ( .A1(n54248), .A2(n54245), .A3(n54246), .A4(n54247), .ZN(
        n54250) );
  BUF_X4 U6675 ( .I(n48082), .Z(n23617) );
  INV_X2 U6690 ( .I(n12269), .ZN(n13359) );
  NOR2_X1 U6694 ( .A1(n15238), .A2(n645), .ZN(n56465) );
  NOR2_X2 U6699 ( .A1(n11814), .A2(n11815), .ZN(n16490) );
  INV_X2 U6700 ( .I(n647), .ZN(n25141) );
  NAND2_X2 U6704 ( .A1(n41610), .A2(n1699), .ZN(n5364) );
  INV_X2 U6705 ( .I(n648), .ZN(n6306) );
  AND2_X1 U6708 ( .A1(n15738), .A2(n25052), .Z(n30757) );
  XOR2_X1 U6710 ( .A1(n651), .A2(n19237), .Z(n3018) );
  NOR2_X2 U6726 ( .A1(n1233), .A2(n55102), .ZN(n55075) );
  NAND3_X2 U6727 ( .A1(n1959), .A2(n1162), .A3(n54994), .ZN(n55102) );
  AND2_X1 U6728 ( .A1(n3505), .A2(n23711), .Z(n21928) );
  INV_X2 U6729 ( .I(n29340), .ZN(n10828) );
  XOR2_X1 U6731 ( .A1(n16959), .A2(n32201), .Z(n32203) );
  XOR2_X1 U6735 ( .A1(n656), .A2(n15016), .Z(n16835) );
  INV_X2 U6753 ( .I(n54823), .ZN(n14501) );
  NAND2_X2 U6759 ( .A1(n61733), .A2(n14729), .ZN(n30725) );
  INV_X4 U6760 ( .I(n23588), .ZN(n47329) );
  NOR2_X2 U6763 ( .A1(n54549), .A2(n54523), .ZN(n54580) );
  XOR2_X1 U6764 ( .A1(n7999), .A2(n46236), .Z(n13853) );
  XOR2_X1 U6766 ( .A1(n64039), .A2(n44854), .Z(n45035) );
  XOR2_X1 U6768 ( .A1(n666), .A2(n665), .Z(n24830) );
  INV_X2 U6773 ( .I(n35254), .ZN(n1794) );
  INV_X4 U6774 ( .I(n18452), .ZN(n2457) );
  INV_X2 U6775 ( .I(n667), .ZN(n18230) );
  NAND2_X2 U6778 ( .A1(n364), .A2(n59798), .ZN(n22796) );
  NAND2_X2 U6786 ( .A1(n49107), .A2(n49106), .ZN(n49794) );
  XOR2_X1 U6791 ( .A1(n670), .A2(n54556), .Z(Plaintext[75]) );
  OAI21_X1 U6792 ( .A1(n54554), .A2(n54555), .B(n54553), .ZN(n670) );
  BUF_X2 U6798 ( .I(n5054), .Z(n674) );
  NAND2_X2 U6802 ( .A1(n18425), .A2(n22572), .ZN(n54531) );
  NOR3_X2 U6804 ( .A1(n39917), .A2(n39916), .A3(n39915), .ZN(n39918) );
  OAI22_X2 U6807 ( .A1(n7697), .A2(n22760), .B1(n55018), .B2(n55020), .ZN(
        n4984) );
  XOR2_X1 U6810 ( .A1(n52473), .A2(n13687), .Z(n52499) );
  INV_X2 U6811 ( .I(n686), .ZN(n17464) );
  BUF_X4 U6813 ( .I(n55356), .Z(n14428) );
  NOR2_X2 U6820 ( .A1(n26052), .A2(n58580), .ZN(n36081) );
  NOR2_X2 U6821 ( .A1(n36081), .A2(n63430), .ZN(n36780) );
  XOR2_X1 U6823 ( .A1(n45004), .A2(n18727), .Z(n688) );
  NAND3_X2 U6825 ( .A1(n5407), .A2(n29110), .A3(n29109), .ZN(n689) );
  XOR2_X1 U6830 ( .A1(n24803), .A2(n765), .Z(n49708) );
  XOR2_X1 U6843 ( .A1(n18584), .A2(n46354), .Z(n16624) );
  XOR2_X1 U6845 ( .A1(n46292), .A2(n8481), .Z(n46547) );
  NAND2_X2 U6853 ( .A1(n37355), .A2(n4541), .ZN(n37105) );
  BUF_X2 U6854 ( .I(n16379), .Z(n696) );
  AOI22_X1 U6862 ( .A1(n699), .A2(n1311), .B1(n34107), .B2(n35182), .ZN(n23681) );
  INV_X2 U6870 ( .I(n6439), .ZN(n10737) );
  NAND3_X2 U6871 ( .A1(n18380), .A2(n35215), .A3(n57986), .ZN(n33823) );
  NAND2_X1 U6875 ( .A1(n40059), .A2(n13875), .ZN(n25852) );
  XOR2_X1 U6890 ( .A1(n32557), .A2(n808), .Z(n710) );
  NOR3_X2 U6891 ( .A1(n711), .A2(n55446), .A3(n61691), .ZN(n21275) );
  NAND2_X2 U6893 ( .A1(n40145), .A2(n39324), .ZN(n3356) );
  XOR2_X1 U6904 ( .A1(n715), .A2(n19991), .Z(n20048) );
  XOR2_X1 U6907 ( .A1(Ciphertext[172]), .A2(Key[41]), .Z(n4604) );
  NOR2_X1 U6912 ( .A1(n41375), .A2(n61417), .ZN(n2341) );
  INV_X2 U6913 ( .I(n16461), .ZN(n41375) );
  NAND2_X2 U6914 ( .A1(n41385), .A2(n39994), .ZN(n16461) );
  NAND2_X2 U6915 ( .A1(n23015), .A2(n27343), .ZN(n25157) );
  NAND2_X2 U6919 ( .A1(n717), .A2(n23295), .ZN(n53911) );
  BUF_X2 U6923 ( .I(n11360), .Z(n718) );
  NAND2_X1 U6925 ( .A1(n49810), .A2(n49811), .ZN(n49814) );
  NAND2_X2 U6934 ( .A1(n30688), .A2(n29029), .ZN(n27362) );
  INV_X4 U6939 ( .I(n12779), .ZN(n25148) );
  NAND3_X2 U6941 ( .A1(n35238), .A2(n58285), .A3(n8223), .ZN(n37398) );
  XOR2_X1 U6944 ( .A1(n725), .A2(n25530), .Z(n46421) );
  XOR2_X1 U6945 ( .A1(n10139), .A2(n57892), .Z(n725) );
  BUF_X2 U6948 ( .I(n33035), .Z(n727) );
  XOR2_X1 U6950 ( .A1(n17238), .A2(n728), .Z(n11500) );
  XOR2_X1 U6951 ( .A1(n18098), .A2(n46655), .Z(n728) );
  XOR2_X1 U6952 ( .A1(n729), .A2(n44608), .Z(n44805) );
  XOR2_X1 U6953 ( .A1(n64373), .A2(n15354), .Z(n729) );
  NAND2_X1 U6958 ( .A1(n26446), .A2(n1575), .ZN(n29296) );
  NAND2_X1 U6959 ( .A1(n24431), .A2(n28510), .ZN(n28516) );
  NAND2_X1 U6962 ( .A1(n9671), .A2(n27568), .ZN(n13379) );
  NOR2_X1 U6963 ( .A1(n28589), .A2(n29641), .ZN(n28593) );
  INV_X1 U6966 ( .I(n27583), .ZN(n1572) );
  INV_X1 U6968 ( .I(n26994), .ZN(n14968) );
  NAND3_X1 U6970 ( .A1(n1880), .A2(n29128), .A3(n29127), .ZN(n13561) );
  INV_X1 U6971 ( .I(n27204), .ZN(n27530) );
  NOR2_X1 U6977 ( .A1(n62714), .A2(n29141), .ZN(n17451) );
  NOR2_X1 U6978 ( .A1(n13482), .A2(n28664), .ZN(n27694) );
  AOI21_X1 U6979 ( .A1(n29129), .A2(n8436), .B(n8613), .ZN(n14918) );
  NOR2_X1 U6982 ( .A1(n26654), .A2(n26360), .ZN(n27569) );
  NAND3_X1 U6983 ( .A1(n20678), .A2(n19423), .A3(n28813), .ZN(n26990) );
  NAND2_X1 U6984 ( .A1(n26912), .A2(n25341), .ZN(n27892) );
  NAND2_X1 U6987 ( .A1(n26265), .A2(n26528), .ZN(n14797) );
  NAND2_X1 U6990 ( .A1(n5070), .A2(n9411), .ZN(n29530) );
  NOR2_X1 U6998 ( .A1(n23317), .A2(n1438), .ZN(n30284) );
  NAND2_X1 U7000 ( .A1(n5243), .A2(n23446), .ZN(n29500) );
  AOI21_X1 U7003 ( .A1(n15116), .A2(n29123), .B(n3087), .ZN(n15115) );
  NOR2_X1 U7004 ( .A1(n31272), .A2(n31159), .ZN(n6319) );
  NAND3_X1 U7005 ( .A1(n20025), .A2(n28989), .A3(n23315), .ZN(n5422) );
  NAND2_X1 U7006 ( .A1(n30695), .A2(n31051), .ZN(n30170) );
  NOR3_X1 U7010 ( .A1(n24896), .A2(n28696), .A3(n29820), .ZN(n29998) );
  OAI21_X1 U7014 ( .A1(n28989), .A2(n13175), .B(n30021), .ZN(n27736) );
  AOI21_X1 U7022 ( .A1(n27308), .A2(n3052), .B(n1859), .ZN(n1925) );
  NOR2_X1 U7027 ( .A1(n14216), .A2(n30003), .ZN(n13215) );
  NOR2_X1 U7028 ( .A1(n5866), .A2(n22742), .ZN(n5983) );
  NAND2_X1 U7030 ( .A1(n29434), .A2(n28957), .ZN(n29447) );
  INV_X1 U7034 ( .I(n24292), .ZN(n31682) );
  INV_X1 U7035 ( .I(n5435), .ZN(n1822) );
  NAND2_X1 U7037 ( .A1(n57342), .A2(n35709), .ZN(n11618) );
  NOR2_X1 U7038 ( .A1(n35799), .A2(n7272), .ZN(n34222) );
  INV_X1 U7042 ( .I(n34618), .ZN(n1810) );
  INV_X1 U7046 ( .I(n35802), .ZN(n1805) );
  NAND2_X1 U7047 ( .A1(n11477), .A2(n8694), .ZN(n34554) );
  NOR2_X1 U7048 ( .A1(n34798), .A2(n61748), .ZN(n33762) );
  NAND2_X1 U7049 ( .A1(n11182), .A2(n35272), .ZN(n34387) );
  NOR2_X1 U7053 ( .A1(n7883), .A2(n34970), .ZN(n34538) );
  NOR2_X1 U7054 ( .A1(n34972), .A2(n34970), .ZN(n20895) );
  NOR2_X1 U7059 ( .A1(n34714), .A2(n22633), .ZN(n35304) );
  OR2_X1 U7069 ( .A1(n25396), .A2(n21921), .Z(n35925) );
  INV_X1 U7088 ( .I(n22113), .ZN(n1790) );
  OAI21_X1 U7093 ( .A1(n35913), .A2(n6540), .B(n17660), .ZN(n11612) );
  NAND2_X1 U7098 ( .A1(n22659), .A2(n21536), .ZN(n2279) );
  NAND3_X1 U7099 ( .A1(n37357), .A2(n1524), .A3(n36288), .ZN(n18776) );
  INV_X1 U7106 ( .I(n53090), .ZN(n10499) );
  INV_X1 U7111 ( .I(n54168), .ZN(n19545) );
  INV_X1 U7113 ( .I(n16558), .ZN(n15458) );
  NAND2_X1 U7118 ( .A1(n40952), .A2(n40944), .ZN(n10735) );
  NAND2_X1 U7120 ( .A1(n1274), .A2(n42211), .ZN(n38136) );
  OAI21_X1 U7124 ( .A1(n41430), .A2(n41433), .B(n22638), .ZN(n41436) );
  NOR2_X1 U7125 ( .A1(n6412), .A2(n22776), .ZN(n40818) );
  AND2_X1 U7131 ( .A1(n42264), .A2(n42263), .Z(n992) );
  INV_X1 U7139 ( .I(n40645), .ZN(n18836) );
  NOR3_X1 U7140 ( .A1(n23108), .A2(n61950), .A3(n61013), .ZN(n15340) );
  NOR3_X1 U7143 ( .A1(n38045), .A2(n39104), .A3(n40203), .ZN(n15482) );
  NOR2_X1 U7149 ( .A1(n42653), .A2(n6900), .ZN(n6899) );
  NOR2_X1 U7151 ( .A1(n42598), .A2(n42605), .ZN(n41544) );
  INV_X1 U7152 ( .I(n5488), .ZN(n40626) );
  NOR2_X1 U7153 ( .A1(n8536), .A2(n62175), .ZN(n9590) );
  NAND3_X1 U7161 ( .A1(n40794), .A2(n41262), .A3(n11316), .ZN(n11260) );
  OR2_X1 U7164 ( .A1(n42393), .A2(n19517), .Z(n1042) );
  INV_X1 U7167 ( .I(n40417), .ZN(n39981) );
  AOI22_X1 U7169 ( .A1(n40077), .A2(n40076), .B1(n2159), .B2(n40078), .ZN(
        n40079) );
  NOR2_X1 U7174 ( .A1(n11196), .A2(n6879), .ZN(n6878) );
  NOR2_X1 U7178 ( .A1(n42327), .A2(n42324), .ZN(n43017) );
  NOR2_X1 U7179 ( .A1(n12312), .A2(n26020), .ZN(n42413) );
  NOR2_X1 U7188 ( .A1(n6995), .A2(n41254), .ZN(n43247) );
  NOR2_X1 U7190 ( .A1(n1715), .A2(n14920), .ZN(n2450) );
  NOR2_X1 U7193 ( .A1(n43297), .A2(n17176), .ZN(n43950) );
  INV_X1 U7200 ( .I(n56915), .ZN(n15564) );
  NOR3_X1 U7203 ( .A1(n19271), .A2(n42760), .A3(n8937), .ZN(n8936) );
  OAI21_X1 U7204 ( .A1(n43111), .A2(n43282), .B(n43290), .ZN(n6533) );
  INV_X1 U7209 ( .I(n24037), .ZN(n11925) );
  INV_X1 U7210 ( .I(n57096), .ZN(n13281) );
  NOR3_X1 U7214 ( .A1(n16941), .A2(n20841), .A3(n43950), .ZN(n16548) );
  INV_X1 U7215 ( .I(n43953), .ZN(n43301) );
  AOI21_X1 U7218 ( .A1(n14183), .A2(n8213), .B(n41716), .ZN(n41718) );
  INV_X1 U7224 ( .I(n21253), .ZN(n23497) );
  AOI21_X1 U7225 ( .A1(n23643), .A2(n15697), .B(n18196), .ZN(n9512) );
  INV_X1 U7226 ( .I(n44224), .ZN(n46451) );
  NOR2_X1 U7233 ( .A1(n47481), .A2(n6957), .ZN(n48658) );
  NOR2_X1 U7235 ( .A1(n14323), .A2(n23180), .ZN(n47385) );
  NAND2_X1 U7237 ( .A1(n22772), .A2(n47275), .ZN(n47582) );
  NOR2_X1 U7251 ( .A1(n47259), .A2(n24558), .ZN(n44483) );
  NAND2_X1 U7261 ( .A1(n23802), .A2(n47943), .ZN(n47944) );
  NAND3_X1 U7264 ( .A1(n50363), .A2(n20894), .A3(n26208), .ZN(n16540) );
  AND2_X1 U7266 ( .A1(n46957), .A2(n1328), .Z(n1081) );
  INV_X1 U7267 ( .I(n45304), .ZN(n45464) );
  OAI21_X1 U7272 ( .A1(n50143), .A2(n14617), .B(n50062), .ZN(n50064) );
  NAND2_X1 U7277 ( .A1(n406), .A2(n49195), .ZN(n49191) );
  NOR2_X1 U7291 ( .A1(n4297), .A2(n49780), .ZN(n4296) );
  NOR3_X1 U7293 ( .A1(n9324), .A2(n48019), .A3(n48275), .ZN(n9323) );
  NOR2_X1 U7296 ( .A1(n25091), .A2(n2810), .ZN(n49048) );
  INV_X1 U7303 ( .I(n54249), .ZN(n11409) );
  NOR3_X1 U7306 ( .A1(n49830), .A2(n49829), .A3(n49828), .ZN(n49841) );
  INV_X1 U7308 ( .I(n15487), .ZN(n9545) );
  NOR2_X1 U7313 ( .A1(n55265), .A2(n55270), .ZN(n5276) );
  NOR2_X1 U7315 ( .A1(n25160), .A2(n53214), .ZN(n57022) );
  INV_X1 U7316 ( .I(n54998), .ZN(n55306) );
  NAND2_X1 U7317 ( .A1(n64255), .A2(n5276), .ZN(n5275) );
  NAND2_X1 U7318 ( .A1(n10523), .A2(n14457), .ZN(n4125) );
  NOR2_X1 U7319 ( .A1(n52699), .A2(n16329), .ZN(n57010) );
  NAND3_X1 U7320 ( .A1(n55473), .A2(n14352), .A3(n55281), .ZN(n55282) );
  NAND2_X1 U7322 ( .A1(n55323), .A2(n55438), .ZN(n55308) );
  NAND2_X1 U7325 ( .A1(n10040), .A2(n56268), .ZN(n55927) );
  INV_X1 U7330 ( .I(n54431), .ZN(n54780) );
  OAI22_X1 U7332 ( .A1(n55703), .A2(n18597), .B1(n1369), .B2(n62263), .ZN(
        n55708) );
  NOR2_X1 U7333 ( .A1(n24455), .A2(n15730), .ZN(n55975) );
  AOI21_X1 U7341 ( .A1(n54963), .A2(n54964), .B(n9106), .ZN(n9105) );
  NAND4_X1 U7342 ( .A1(n4241), .A2(n54780), .A3(n54779), .A4(n22231), .ZN(
        n4240) );
  NAND2_X1 U7353 ( .A1(n55820), .A2(n55813), .ZN(n55831) );
  INV_X1 U7354 ( .I(n53738), .ZN(n21973) );
  OAI21_X1 U7356 ( .A1(n55082), .A2(n25170), .B(n15520), .ZN(n8408) );
  NAND3_X1 U7360 ( .A1(n53047), .A2(n53798), .A3(n53046), .ZN(n17640) );
  NAND3_X1 U7363 ( .A1(n55780), .A2(n14890), .A3(n24958), .ZN(n55803) );
  NAND4_X1 U7366 ( .A1(n5614), .A2(n53167), .A3(n3525), .A4(n15415), .ZN(
        n53168) );
  NOR2_X1 U7371 ( .A1(n11548), .A2(n55101), .ZN(n10775) );
  NAND3_X1 U7375 ( .A1(n54912), .A2(n54929), .A3(n54911), .ZN(n2051) );
  OAI21_X1 U7381 ( .A1(n13240), .A2(n13239), .B(n53280), .ZN(n53283) );
  AOI21_X1 U7383 ( .A1(n56326), .A2(n56325), .B(n56340), .ZN(n56333) );
  OAI21_X1 U7384 ( .A1(n55074), .A2(n55089), .B(n10775), .ZN(n10774) );
  INV_X1 U7385 ( .I(n51019), .ZN(n53328) );
  INV_X1 U7386 ( .I(n54917), .ZN(n54918) );
  XNOR2_X1 U7388 ( .A1(n31135), .A2(n31630), .ZN(n730) );
  XOR2_X1 U7392 ( .A1(n51928), .A2(n38401), .Z(n733) );
  OR2_X1 U7393 ( .A1(n39124), .A2(n64571), .Z(n734) );
  XNOR2_X1 U7394 ( .A1(n23069), .A2(n52420), .ZN(n735) );
  OR2_X1 U7395 ( .A1(n54904), .A2(n2329), .Z(n736) );
  OR2_X1 U7396 ( .A1(n48730), .A2(n24692), .Z(n737) );
  XNOR2_X1 U7397 ( .A1(n1819), .A2(n65197), .ZN(n738) );
  OR2_X1 U7398 ( .A1(n17379), .A2(n24788), .Z(n739) );
  XNOR2_X1 U7401 ( .A1(n11529), .A2(n6701), .ZN(n742) );
  XNOR2_X1 U7402 ( .A1(n7811), .A2(n24744), .ZN(n743) );
  XNOR2_X1 U7403 ( .A1(n9602), .A2(n20194), .ZN(n744) );
  XNOR2_X1 U7404 ( .A1(n25376), .A2(n37745), .ZN(n746) );
  AND2_X1 U7405 ( .A1(n24879), .A2(n24877), .Z(n747) );
  XNOR2_X1 U7406 ( .A1(n52154), .A2(n52321), .ZN(n748) );
  XNOR2_X1 U7408 ( .A1(n64360), .A2(n32636), .ZN(n750) );
  XNOR2_X1 U7410 ( .A1(n31018), .A2(n61610), .ZN(n752) );
  NOR2_X1 U7413 ( .A1(n28469), .A2(n4848), .ZN(n1971) );
  XNOR2_X1 U7414 ( .A1(n50126), .A2(n50724), .ZN(n756) );
  XNOR2_X1 U7416 ( .A1(n8559), .A2(n58926), .ZN(n758) );
  AND2_X1 U7417 ( .A1(n42660), .A2(n42659), .Z(n760) );
  AND2_X1 U7418 ( .A1(n4497), .A2(n29509), .Z(n761) );
  OR2_X1 U7419 ( .A1(n18223), .A2(n6215), .Z(n762) );
  XNOR2_X1 U7420 ( .A1(n32414), .A2(n23090), .ZN(n763) );
  XNOR2_X1 U7422 ( .A1(n49693), .A2(n49692), .ZN(n765) );
  XNOR2_X1 U7423 ( .A1(n46124), .A2(n44960), .ZN(n766) );
  XNOR2_X1 U7424 ( .A1(n62616), .A2(n55833), .ZN(n767) );
  XNOR2_X1 U7427 ( .A1(n39721), .A2(n18829), .ZN(n768) );
  XNOR2_X1 U7428 ( .A1(n19860), .A2(n24043), .ZN(n769) );
  AND2_X1 U7429 ( .A1(n49728), .A2(n63084), .Z(n771) );
  XNOR2_X1 U7430 ( .A1(n10430), .A2(n11220), .ZN(n772) );
  XNOR2_X1 U7431 ( .A1(n32524), .A2(n32523), .ZN(n773) );
  XNOR2_X1 U7432 ( .A1(Ciphertext[105]), .A2(Ciphertext[102]), .ZN(n774) );
  XNOR2_X1 U7433 ( .A1(n38629), .A2(n39183), .ZN(n776) );
  XNOR2_X1 U7437 ( .A1(n50514), .A2(n53174), .ZN(n778) );
  XNOR2_X1 U7438 ( .A1(n45847), .A2(n53102), .ZN(n779) );
  XNOR2_X1 U7439 ( .A1(n51002), .A2(n51001), .ZN(n781) );
  XNOR2_X1 U7440 ( .A1(n50070), .A2(n50069), .ZN(n782) );
  XNOR2_X1 U7441 ( .A1(n51132), .A2(n47937), .ZN(n783) );
  XNOR2_X1 U7442 ( .A1(n38994), .A2(n15630), .ZN(n784) );
  XNOR2_X1 U7443 ( .A1(n51512), .A2(n56165), .ZN(n785) );
  XNOR2_X1 U7446 ( .A1(n39471), .A2(n39470), .ZN(n788) );
  XNOR2_X1 U7447 ( .A1(n50526), .A2(n36658), .ZN(n789) );
  XNOR2_X1 U7448 ( .A1(n51188), .A2(n38964), .ZN(n790) );
  XNOR2_X1 U7450 ( .A1(n37638), .A2(n24109), .ZN(n792) );
  XNOR2_X1 U7451 ( .A1(n39724), .A2(n27793), .ZN(n793) );
  XNOR2_X1 U7452 ( .A1(n46124), .A2(n56771), .ZN(n794) );
  XNOR2_X1 U7453 ( .A1(n45820), .A2(n45819), .ZN(n796) );
  XNOR2_X1 U7454 ( .A1(n51323), .A2(n44333), .ZN(n797) );
  XNOR2_X1 U7455 ( .A1(n46324), .A2(n46323), .ZN(n799) );
  XNOR2_X1 U7456 ( .A1(n46170), .A2(n38086), .ZN(n800) );
  XNOR2_X1 U7457 ( .A1(n51523), .A2(n44463), .ZN(n801) );
  XNOR2_X1 U7458 ( .A1(n45352), .A2(n45351), .ZN(n802) );
  XNOR2_X1 U7459 ( .A1(n52330), .A2(n52329), .ZN(n803) );
  XOR2_X1 U7460 ( .A1(n52050), .A2(n50777), .Z(n804) );
  XNOR2_X1 U7461 ( .A1(n51169), .A2(n45471), .ZN(n805) );
  XNOR2_X1 U7463 ( .A1(n38575), .A2(n37671), .ZN(n806) );
  XNOR2_X1 U7464 ( .A1(n31489), .A2(n32267), .ZN(n807) );
  XNOR2_X1 U7465 ( .A1(n32561), .A2(n32560), .ZN(n808) );
  XNOR2_X1 U7467 ( .A1(n52530), .A2(n15652), .ZN(n810) );
  XNOR2_X1 U7468 ( .A1(n11111), .A2(n816), .ZN(n811) );
  XNOR2_X1 U7472 ( .A1(n49669), .A2(n38655), .ZN(n813) );
  XOR2_X1 U7473 ( .A1(Ciphertext[70]), .A2(Key[95]), .Z(n814) );
  INV_X1 U7475 ( .I(n11977), .ZN(n11975) );
  XNOR2_X1 U7476 ( .A1(n44746), .A2(n44745), .ZN(n816) );
  XNOR2_X1 U7477 ( .A1(n37349), .A2(n52614), .ZN(n817) );
  XNOR2_X1 U7479 ( .A1(n51596), .A2(n36218), .ZN(n819) );
  XNOR2_X1 U7484 ( .A1(n51614), .A2(n51613), .ZN(n824) );
  XNOR2_X1 U7487 ( .A1(n52320), .A2(n52319), .ZN(n827) );
  XNOR2_X1 U7488 ( .A1(n40459), .A2(n37348), .ZN(n828) );
  XNOR2_X1 U7489 ( .A1(n45416), .A2(n31696), .ZN(n829) );
  INV_X1 U7492 ( .I(n902), .ZN(n35023) );
  OR2_X1 U7493 ( .A1(n27525), .A2(n27204), .Z(n830) );
  XNOR2_X1 U7496 ( .A1(n51817), .A2(n51816), .ZN(n834) );
  XNOR2_X1 U7499 ( .A1(Ciphertext[156]), .A2(Ciphertext[159]), .ZN(n836) );
  XOR2_X1 U7500 ( .A1(Ciphertext[50]), .A2(Key[147]), .Z(n837) );
  AND2_X2 U7504 ( .A1(n10661), .A2(n10602), .Z(n839) );
  BUF_X2 U7505 ( .I(n13204), .Z(n13163) );
  XNOR2_X1 U7506 ( .A1(n44023), .A2(n32097), .ZN(n840) );
  XOR2_X1 U7507 ( .A1(n44949), .A2(n31635), .Z(n841) );
  OR2_X1 U7508 ( .A1(n13817), .A2(n23734), .Z(n842) );
  XNOR2_X1 U7510 ( .A1(n31381), .A2(n44622), .ZN(n843) );
  XNOR2_X1 U7512 ( .A1(n44087), .A2(n31484), .ZN(n844) );
  XOR2_X1 U7513 ( .A1(n30908), .A2(n18467), .Z(n845) );
  OR2_X2 U7514 ( .A1(n28920), .A2(n30292), .Z(n846) );
  OR2_X2 U7515 ( .A1(n27705), .A2(n27706), .Z(n847) );
  XNOR2_X1 U7516 ( .A1(n49967), .A2(n49966), .ZN(n848) );
  XNOR2_X1 U7523 ( .A1(n33164), .A2(n32175), .ZN(n853) );
  XNOR2_X1 U7524 ( .A1(Ciphertext[174]), .A2(Ciphertext[177]), .ZN(n854) );
  XNOR2_X1 U7526 ( .A1(n62323), .A2(n31437), .ZN(n857) );
  INV_X1 U7529 ( .I(n8518), .ZN(n26460) );
  INV_X1 U7533 ( .I(n19144), .ZN(n25966) );
  AND3_X2 U7534 ( .A1(n22959), .A2(n49107), .A3(n49106), .Z(n858) );
  XNOR2_X1 U7536 ( .A1(n51120), .A2(n51032), .ZN(n859) );
  INV_X1 U7537 ( .I(n56229), .ZN(n16753) );
  XNOR2_X1 U7539 ( .A1(n61178), .A2(n51135), .ZN(n861) );
  XNOR2_X1 U7546 ( .A1(n17441), .A2(n63002), .ZN(n865) );
  XNOR2_X1 U7547 ( .A1(n535), .A2(n52567), .ZN(n866) );
  XNOR2_X1 U7549 ( .A1(n19785), .A2(n51592), .ZN(n868) );
  INV_X1 U7550 ( .I(n5056), .ZN(n54444) );
  XNOR2_X1 U7553 ( .A1(n51968), .A2(n39559), .ZN(n870) );
  INV_X4 U7554 ( .I(n3697), .ZN(n27374) );
  XNOR2_X1 U7558 ( .A1(n13181), .A2(n31814), .ZN(n876) );
  XOR2_X1 U7559 ( .A1(n31854), .A2(n31853), .Z(n877) );
  XNOR2_X1 U7560 ( .A1(n30913), .A2(n25886), .ZN(n878) );
  XNOR2_X1 U7562 ( .A1(n17112), .A2(n752), .ZN(n880) );
  XNOR2_X1 U7565 ( .A1(n5009), .A2(n31109), .ZN(n882) );
  AND2_X1 U7566 ( .A1(n12174), .A2(n2370), .Z(n883) );
  INV_X4 U7571 ( .I(n2614), .ZN(n13487) );
  BUF_X2 U7572 ( .I(n5604), .Z(n11186) );
  INV_X2 U7573 ( .I(n30945), .ZN(n33857) );
  XNOR2_X1 U7574 ( .A1(n31930), .A2(n31929), .ZN(n886) );
  INV_X2 U7576 ( .I(n6530), .ZN(n6529) );
  XNOR2_X1 U7577 ( .A1(n33190), .A2(n25843), .ZN(n888) );
  XOR2_X1 U7578 ( .A1(n12976), .A2(n12977), .Z(n889) );
  AND2_X1 U7581 ( .A1(n3903), .A2(n35848), .Z(n891) );
  XNOR2_X1 U7584 ( .A1(n13962), .A2(n5436), .ZN(n893) );
  AND2_X1 U7586 ( .A1(n23117), .A2(n34620), .Z(n896) );
  INV_X2 U7587 ( .I(n34720), .ZN(n15181) );
  XNOR2_X1 U7590 ( .A1(n33172), .A2(n24666), .ZN(n898) );
  XOR2_X1 U7592 ( .A1(n7884), .A2(n25338), .Z(n900) );
  INV_X4 U7594 ( .I(n15144), .ZN(n15756) );
  XOR2_X1 U7596 ( .A1(n25325), .A2(n30988), .Z(n901) );
  OR2_X2 U7598 ( .A1(n13195), .A2(n8514), .Z(n904) );
  AND2_X1 U7600 ( .A1(n18834), .A2(n24983), .Z(n906) );
  INV_X2 U7609 ( .I(n19606), .ZN(n9956) );
  INV_X4 U7614 ( .I(n36256), .ZN(n19231) );
  AND2_X1 U7615 ( .A1(n15085), .A2(n1424), .Z(n914) );
  INV_X2 U7617 ( .I(n38988), .ZN(n4762) );
  XNOR2_X1 U7618 ( .A1(n10402), .A2(n52082), .ZN(n915) );
  XNOR2_X1 U7619 ( .A1(n39275), .A2(n50793), .ZN(n916) );
  INV_X4 U7620 ( .I(n25366), .ZN(n36026) );
  XOR2_X1 U7623 ( .A1(n1762), .A2(n15309), .Z(n920) );
  XNOR2_X1 U7626 ( .A1(n1200), .A2(n805), .ZN(n922) );
  XNOR2_X1 U7629 ( .A1(n36637), .A2(n36636), .ZN(n925) );
  XNOR2_X1 U7631 ( .A1(n23583), .A2(n11751), .ZN(n927) );
  XNOR2_X1 U7633 ( .A1(n38973), .A2(n36018), .ZN(n929) );
  OR2_X1 U7635 ( .A1(n7380), .A2(n36152), .Z(n931) );
  AND3_X2 U7637 ( .A1(n1418), .A2(n35344), .A3(n2418), .Z(n933) );
  XNOR2_X1 U7638 ( .A1(n26021), .A2(n2114), .ZN(n934) );
  XNOR2_X1 U7639 ( .A1(n39710), .A2(n38386), .ZN(n935) );
  XNOR2_X1 U7640 ( .A1(n38786), .A2(n38785), .ZN(n936) );
  XOR2_X1 U7641 ( .A1(n39692), .A2(n38985), .Z(n937) );
  XNOR2_X1 U7645 ( .A1(n38308), .A2(n38371), .ZN(n940) );
  XNOR2_X1 U7647 ( .A1(n58203), .A2(n16312), .ZN(n942) );
  XNOR2_X1 U7648 ( .A1(n38376), .A2(n38375), .ZN(n944) );
  XNOR2_X1 U7650 ( .A1(n39358), .A2(n19217), .ZN(n946) );
  AND2_X1 U7651 ( .A1(n35972), .A2(n35973), .Z(n949) );
  XNOR2_X1 U7653 ( .A1(n37807), .A2(n38821), .ZN(n951) );
  INV_X1 U7655 ( .I(n9255), .ZN(n39190) );
  XNOR2_X1 U7657 ( .A1(n37525), .A2(n37898), .ZN(n953) );
  XNOR2_X1 U7659 ( .A1(n2191), .A2(n6847), .ZN(n955) );
  XNOR2_X1 U7661 ( .A1(n39003), .A2(n39004), .ZN(n957) );
  XNOR2_X1 U7664 ( .A1(n39768), .A2(n24860), .ZN(n959) );
  XNOR2_X1 U7665 ( .A1(n23493), .A2(n37769), .ZN(n960) );
  XNOR2_X1 U7669 ( .A1(n38151), .A2(n768), .ZN(n963) );
  XNOR2_X1 U7670 ( .A1(n37309), .A2(n7212), .ZN(n964) );
  AND2_X1 U7676 ( .A1(n40203), .A2(n40943), .Z(n967) );
  NAND2_X1 U7677 ( .A1(n42284), .A2(n15645), .ZN(n42277) );
  XNOR2_X1 U7678 ( .A1(n38117), .A2(n38116), .ZN(n968) );
  BUF_X4 U7679 ( .I(n38338), .Z(n42427) );
  AND2_X1 U7686 ( .A1(n10735), .A2(n10341), .Z(n973) );
  AND2_X1 U7687 ( .A1(n40722), .A2(n40723), .Z(n974) );
  INV_X4 U7693 ( .I(n41043), .ZN(n3619) );
  INV_X2 U7695 ( .I(n11278), .ZN(n17752) );
  XNOR2_X1 U7697 ( .A1(n37800), .A2(n38219), .ZN(n980) );
  XNOR2_X1 U7698 ( .A1(n21609), .A2(n36243), .ZN(n981) );
  OR2_X1 U7701 ( .A1(n2081), .A2(n40441), .Z(n985) );
  INV_X4 U7703 ( .I(n11818), .ZN(n43601) );
  NAND2_X1 U7706 ( .A1(n24250), .A2(n4659), .ZN(n986) );
  INV_X4 U7708 ( .I(n61475), .ZN(n20601) );
  AND2_X1 U7711 ( .A1(n3535), .A2(n42298), .Z(n987) );
  BUF_X4 U7715 ( .I(n24243), .Z(n9200) );
  INV_X2 U7718 ( .I(n42583), .ZN(n42155) );
  XOR2_X1 U7719 ( .A1(n5639), .A2(n5638), .Z(n990) );
  AND2_X1 U7722 ( .A1(n41836), .A2(n57545), .Z(n991) );
  AND2_X1 U7727 ( .A1(n43715), .A2(n13207), .Z(n1000) );
  XNOR2_X1 U7730 ( .A1(n65082), .A2(n45280), .ZN(n1003) );
  AND2_X1 U7731 ( .A1(n40558), .A2(n41137), .Z(n1004) );
  OR2_X1 U7732 ( .A1(n43342), .A2(n41624), .Z(n1005) );
  XNOR2_X1 U7738 ( .A1(n42179), .A2(n42178), .ZN(n1011) );
  XNOR2_X1 U7741 ( .A1(n18133), .A2(n1003), .ZN(n1013) );
  NOR3_X1 U7747 ( .A1(n43189), .A2(n43188), .A3(n43513), .ZN(n1017) );
  XNOR2_X1 U7749 ( .A1(n23818), .A2(n45408), .ZN(n1018) );
  INV_X2 U7750 ( .I(n41118), .ZN(n39999) );
  XOR2_X1 U7751 ( .A1(n23953), .A2(n46117), .Z(n1019) );
  XNOR2_X1 U7753 ( .A1(n44954), .A2(n44953), .ZN(n1021) );
  XNOR2_X1 U7755 ( .A1(n44806), .A2(n4703), .ZN(n1023) );
  INV_X1 U7762 ( .I(n23314), .ZN(n21800) );
  NOR2_X2 U7767 ( .A1(n1494), .A2(n11609), .ZN(n11608) );
  AND2_X1 U7769 ( .A1(n6899), .A2(n62237), .Z(n1031) );
  XNOR2_X1 U7771 ( .A1(n46519), .A2(n20626), .ZN(n1033) );
  OAI21_X2 U7773 ( .A1(n43777), .A2(n43776), .B(n12091), .ZN(n6233) );
  NOR2_X2 U7774 ( .A1(n16244), .A2(n21517), .ZN(n21516) );
  AND2_X1 U7775 ( .A1(n9063), .A2(n2588), .Z(n1034) );
  XNOR2_X1 U7777 ( .A1(n44089), .A2(n44090), .ZN(n1036) );
  XNOR2_X1 U7779 ( .A1(n45044), .A2(n45043), .ZN(n1038) );
  XOR2_X1 U7780 ( .A1(n5767), .A2(n45333), .Z(n1039) );
  XNOR2_X1 U7782 ( .A1(n44269), .A2(n18900), .ZN(n1041) );
  XOR2_X1 U7786 ( .A1(n45875), .A2(n23566), .Z(n1045) );
  XNOR2_X1 U7790 ( .A1(n2506), .A2(n2504), .ZN(n1050) );
  INV_X4 U7791 ( .I(n2766), .ZN(n44065) );
  XNOR2_X1 U7793 ( .A1(n64013), .A2(n44081), .ZN(n1052) );
  INV_X1 U7795 ( .I(n6563), .ZN(n24576) );
  XNOR2_X1 U7797 ( .A1(n21596), .A2(n6567), .ZN(n1056) );
  INV_X1 U7798 ( .I(n8639), .ZN(n48606) );
  INV_X1 U7799 ( .I(n11416), .ZN(n44577) );
  XNOR2_X1 U7801 ( .A1(n46298), .A2(n24278), .ZN(n1057) );
  OR2_X1 U7806 ( .A1(n41541), .A2(n8799), .Z(n1061) );
  INV_X4 U7808 ( .I(n17464), .ZN(n25896) );
  XNOR2_X1 U7809 ( .A1(n24133), .A2(n44755), .ZN(n1062) );
  XNOR2_X1 U7810 ( .A1(n45099), .A2(n22199), .ZN(n1063) );
  INV_X1 U7812 ( .I(n47653), .ZN(n47830) );
  AND2_X1 U7816 ( .A1(n48582), .A2(n178), .Z(n1065) );
  OR2_X2 U7822 ( .A1(n25444), .A2(n44779), .Z(n1070) );
  OR2_X1 U7824 ( .A1(n45225), .A2(n47605), .Z(n1073) );
  NAND2_X1 U7825 ( .A1(n18570), .A2(n16798), .ZN(n1074) );
  AND2_X1 U7827 ( .A1(n48463), .A2(n14521), .Z(n1075) );
  XNOR2_X1 U7830 ( .A1(n20301), .A2(n1214), .ZN(n1077) );
  INV_X2 U7832 ( .I(n47429), .ZN(n45794) );
  OR2_X2 U7833 ( .A1(n24047), .A2(n21653), .Z(n1078) );
  AND2_X2 U7845 ( .A1(n13719), .A2(n1669), .Z(n1085) );
  AND2_X1 U7849 ( .A1(n47646), .A2(n49687), .Z(n1089) );
  INV_X4 U7853 ( .I(n48729), .ZN(n49929) );
  INV_X4 U7859 ( .I(n48742), .ZN(n13614) );
  INV_X2 U7861 ( .I(n22805), .ZN(n25680) );
  OR2_X1 U7862 ( .A1(n49889), .A2(n10264), .Z(n1096) );
  INV_X4 U7865 ( .I(n49013), .ZN(n25459) );
  AND2_X1 U7866 ( .A1(n24305), .A2(n24304), .Z(n1099) );
  OR2_X1 U7868 ( .A1(n47969), .A2(n47357), .Z(n1101) );
  XNOR2_X1 U7869 ( .A1(n50611), .A2(n3741), .ZN(n1102) );
  AND2_X1 U7871 ( .A1(n22508), .A2(n2179), .Z(n1103) );
  NAND2_X1 U7873 ( .A1(n49466), .A2(n6313), .ZN(n49752) );
  XNOR2_X1 U7875 ( .A1(n18307), .A2(n17234), .ZN(n1106) );
  OR2_X1 U7883 ( .A1(n58636), .A2(n45182), .Z(n1112) );
  AND2_X1 U7884 ( .A1(n18769), .A2(n49539), .Z(n1113) );
  XNOR2_X1 U7889 ( .A1(n51931), .A2(n52092), .ZN(n1116) );
  XNOR2_X1 U7892 ( .A1(n52406), .A2(n52054), .ZN(n1119) );
  INV_X1 U7895 ( .I(n23796), .ZN(n15718) );
  XNOR2_X1 U7896 ( .A1(n51539), .A2(n51538), .ZN(n1122) );
  XNOR2_X1 U7898 ( .A1(n51198), .A2(n1461), .ZN(n1124) );
  INV_X2 U7903 ( .I(n53615), .ZN(n4226) );
  XNOR2_X1 U7905 ( .A1(n51376), .A2(n51377), .ZN(n1128) );
  INV_X4 U7906 ( .I(n56544), .ZN(n52706) );
  XNOR2_X1 U7907 ( .A1(n51772), .A2(n51771), .ZN(n1129) );
  XNOR2_X1 U7909 ( .A1(n8615), .A2(n23032), .ZN(n1132) );
  XOR2_X1 U7912 ( .A1(n13922), .A2(n51417), .Z(n1133) );
  XNOR2_X1 U7913 ( .A1(n50954), .A2(n50953), .ZN(n1135) );
  INV_X1 U7914 ( .I(n55691), .ZN(n20849) );
  AND2_X1 U7923 ( .A1(n25173), .A2(n64808), .Z(n1138) );
  AND2_X2 U7925 ( .A1(n26097), .A2(n2198), .Z(n1139) );
  XNOR2_X1 U7927 ( .A1(n51334), .A2(n52549), .ZN(n1140) );
  OR2_X1 U7928 ( .A1(n53909), .A2(n5025), .Z(n1141) );
  XNOR2_X1 U7932 ( .A1(n52417), .A2(n8821), .ZN(n1144) );
  AND2_X1 U7933 ( .A1(n53378), .A2(n2001), .Z(n1145) );
  BUF_X2 U7936 ( .I(n52380), .Z(n54939) );
  NOR3_X1 U7937 ( .A1(n55471), .A2(n55470), .A3(n55469), .ZN(n1147) );
  OR2_X1 U7939 ( .A1(n8375), .A2(n54470), .Z(n1149) );
  AND2_X1 U7940 ( .A1(n51890), .A2(n56402), .Z(n1150) );
  BUF_X2 U7944 ( .I(n56323), .Z(n12058) );
  INV_X2 U7949 ( .I(n53598), .ZN(n19068) );
  AND2_X1 U7955 ( .A1(n55341), .A2(n55362), .Z(n1165) );
  OR2_X1 U7957 ( .A1(n8325), .A2(n9550), .Z(n1167) );
  BUF_X4 U7960 ( .I(n54191), .Z(n18859) );
  BUF_X2 U7963 ( .I(n25510), .Z(n22401) );
  AND2_X1 U7964 ( .A1(n4336), .A2(n54929), .Z(n1172) );
  AND2_X1 U7966 ( .A1(n54530), .A2(n54558), .Z(n1174) );
  NOR2_X1 U7968 ( .A1(n53184), .A2(n13370), .ZN(n1176) );
  AND2_X1 U7971 ( .A1(n53264), .A2(n53303), .Z(n1178) );
  AND2_X1 U7974 ( .A1(n55347), .A2(n15703), .Z(n1183) );
  INV_X2 U7975 ( .I(n56282), .ZN(n18255) );
  OR2_X1 U7976 ( .A1(n56062), .A2(n56061), .Z(n1184) );
  XNOR2_X1 U7978 ( .A1(n11355), .A2(n20087), .ZN(n1188) );
  AND2_X1 U7979 ( .A1(n20025), .A2(n58696), .Z(n20026) );
  NAND2_X1 U7982 ( .A1(n8437), .A2(n28216), .ZN(n12085) );
  NOR2_X2 U7983 ( .A1(n9144), .A2(n40091), .ZN(n39894) );
  INV_X1 U7995 ( .I(n44227), .ZN(n6006) );
  INV_X2 U7996 ( .I(n44227), .ZN(n43980) );
  NOR3_X1 U8003 ( .A1(n27069), .A2(n27068), .A3(n27067), .ZN(n30024) );
  BUF_X2 U8004 ( .I(n43468), .Z(n1193) );
  NAND2_X1 U8009 ( .A1(n14214), .A2(n42019), .ZN(n43393) );
  NAND3_X2 U8015 ( .A1(n5460), .A2(n16531), .A3(n16530), .ZN(n4839) );
  INV_X1 U8017 ( .I(n51621), .ZN(n7539) );
  NOR3_X2 U8020 ( .A1(n18235), .A2(n15964), .A3(n18233), .ZN(n18232) );
  NAND3_X2 U8023 ( .A1(n38137), .A2(n15797), .A3(n20075), .ZN(n20086) );
  INV_X1 U8029 ( .I(n13364), .ZN(n15736) );
  OAI21_X2 U8038 ( .A1(n33672), .A2(n17283), .B(n12822), .ZN(n12821) );
  NOR2_X2 U8047 ( .A1(n30893), .A2(n20076), .ZN(n30894) );
  NAND4_X2 U8048 ( .A1(n20080), .A2(n31260), .A3(n20078), .A4(n20077), .ZN(
        n20076) );
  AOI21_X2 U8052 ( .A1(n12067), .A2(n31956), .B(n19108), .ZN(n12066) );
  NOR2_X1 U8053 ( .A1(n7092), .A2(n36013), .ZN(n36676) );
  INV_X1 U8055 ( .I(n54021), .ZN(n51870) );
  BUF_X2 U8056 ( .I(n54021), .Z(n11207) );
  NAND3_X1 U8057 ( .A1(n1990), .A2(n33185), .A3(n31169), .ZN(n1983) );
  NOR2_X1 U8065 ( .A1(n19300), .A2(n736), .ZN(n22865) );
  NAND2_X1 U8066 ( .A1(n54890), .A2(n19300), .ZN(n2205) );
  NAND2_X1 U8075 ( .A1(n7932), .A2(n23645), .ZN(n33759) );
  AOI22_X1 U8100 ( .A1(n39881), .A2(n39882), .B1(n5171), .B2(n42006), .ZN(
        n39883) );
  NAND3_X2 U8101 ( .A1(n20476), .A2(n26869), .A3(n26868), .ZN(n26876) );
  NAND2_X1 U8104 ( .A1(n15731), .A2(n60075), .ZN(n42286) );
  INV_X4 U8108 ( .I(n41082), .ZN(n41073) );
  NAND4_X2 U8111 ( .A1(n40343), .A2(n40342), .A3(n40341), .A4(n40340), .ZN(
        n40344) );
  NOR2_X1 U8119 ( .A1(n8029), .A2(n34657), .ZN(n34172) );
  NOR2_X1 U8124 ( .A1(n64416), .A2(n60467), .ZN(n49977) );
  NOR3_X1 U8126 ( .A1(n50340), .A2(n64416), .A3(n50257), .ZN(n21226) );
  OAI22_X1 U8131 ( .A1(n12993), .A2(n48520), .B1(n48519), .B2(n12968), .ZN(
        n48522) );
  NOR2_X1 U8132 ( .A1(n23316), .A2(n12968), .ZN(n48165) );
  INV_X1 U8135 ( .I(n22071), .ZN(n15023) );
  NAND4_X2 U8138 ( .A1(n10307), .A2(n39326), .A3(n39327), .A4(n3466), .ZN(
        n9828) );
  NOR2_X2 U8141 ( .A1(n47601), .A2(n47600), .ZN(n47646) );
  OR2_X2 U8142 ( .A1(n25755), .A2(n1557), .Z(n16907) );
  INV_X1 U8151 ( .I(n18624), .ZN(n3476) );
  INV_X1 U8152 ( .I(n63001), .ZN(n52471) );
  INV_X1 U8155 ( .I(n24753), .ZN(n25177) );
  BUF_X4 U8158 ( .I(n49748), .Z(n16595) );
  NAND2_X1 U8162 ( .A1(n46020), .A2(n46019), .ZN(n24214) );
  NAND4_X2 U8165 ( .A1(n27820), .A2(n27819), .A3(n27818), .A4(n27817), .ZN(
        n27826) );
  NOR2_X2 U8166 ( .A1(n28475), .A2(n27811), .ZN(n27818) );
  OAI21_X2 U8172 ( .A1(n41234), .A2(n1303), .B(n39052), .ZN(n14288) );
  NAND3_X2 U8179 ( .A1(n12996), .A2(n12991), .A3(n12989), .ZN(n12988) );
  NAND4_X1 U8183 ( .A1(n28255), .A2(n28257), .A3(n28256), .A4(n29166), .ZN(
        n28262) );
  NAND3_X1 U8185 ( .A1(n14469), .A2(n54955), .A3(n54611), .ZN(n52386) );
  BUF_X2 U8191 ( .I(n38907), .Z(n24276) );
  NOR2_X1 U8192 ( .A1(n27936), .A2(n10187), .ZN(n27413) );
  NAND4_X1 U8199 ( .A1(n2864), .A2(n54779), .A3(n22231), .A4(n58994), .ZN(
        n54617) );
  NAND2_X1 U8200 ( .A1(n54785), .A2(n54950), .ZN(n2467) );
  NAND2_X1 U8201 ( .A1(n54950), .A2(n1139), .ZN(n2201) );
  NAND2_X1 U8202 ( .A1(n6135), .A2(n2851), .ZN(n53946) );
  BUF_X4 U8207 ( .I(n21713), .Z(n20025) );
  OAI21_X2 U8208 ( .A1(n50270), .A2(n15194), .B(n14254), .ZN(n50282) );
  INV_X1 U8210 ( .I(n36202), .ZN(n36716) );
  NOR2_X1 U8217 ( .A1(n30706), .A2(n24056), .ZN(n15626) );
  NAND4_X2 U8218 ( .A1(n61778), .A2(n2314), .A3(n13965), .A4(n2313), .ZN(n2312) );
  BUF_X4 U8219 ( .I(n9153), .Z(n5267) );
  NAND2_X1 U8221 ( .A1(n59008), .A2(n10053), .ZN(n45908) );
  NAND2_X1 U8231 ( .A1(n42592), .A2(n2884), .ZN(n15307) );
  OAI21_X2 U8233 ( .A1(n60034), .A2(n17488), .B(n36040), .ZN(n4690) );
  NOR2_X1 U8242 ( .A1(n29432), .A2(n28959), .ZN(n29440) );
  INV_X2 U8247 ( .I(n24188), .ZN(n40239) );
  INV_X4 U8248 ( .I(n4899), .ZN(n7854) );
  NAND2_X2 U8250 ( .A1(n25452), .A2(n25454), .ZN(n25449) );
  NAND2_X1 U8252 ( .A1(n56341), .A2(n56352), .ZN(n56328) );
  NAND2_X1 U8256 ( .A1(n33970), .A2(n10358), .ZN(n9542) );
  INV_X2 U8258 ( .I(n55387), .ZN(n55362) );
  NOR2_X1 U8264 ( .A1(n61717), .A2(n412), .ZN(n45941) );
  NAND4_X2 U8274 ( .A1(n22931), .A2(n3681), .A3(n50420), .A4(n48288), .ZN(
        n3680) );
  NOR2_X1 U8281 ( .A1(n63261), .A2(n50004), .ZN(n3461) );
  OAI22_X1 U8285 ( .A1(n35749), .A2(n6051), .B1(n6206), .B2(n61496), .ZN(
        n35746) );
  INV_X1 U8287 ( .I(n38516), .ZN(n25139) );
  INV_X4 U8292 ( .I(n25742), .ZN(n40315) );
  NOR2_X1 U8297 ( .A1(n10193), .A2(n64250), .ZN(n46050) );
  BUF_X4 U8308 ( .I(n8745), .Z(n1225) );
  AOI21_X1 U8310 ( .A1(n48639), .A2(n48630), .B(n48500), .ZN(n48501) );
  NAND3_X2 U8319 ( .A1(n4885), .A2(n8362), .A3(n29362), .ZN(n29363) );
  AND2_X2 U8324 ( .A1(n11188), .A2(n11187), .Z(n5774) );
  NAND2_X1 U8327 ( .A1(n21808), .A2(n21806), .ZN(n1227) );
  BUF_X2 U8328 ( .I(n36178), .Z(n3458) );
  NOR3_X2 U8331 ( .A1(n5860), .A2(n4868), .A3(n57329), .ZN(n5858) );
  INV_X4 U8343 ( .I(n29801), .ZN(n25241) );
  NAND3_X2 U8348 ( .A1(n6858), .A2(n6860), .A3(n762), .ZN(n6024) );
  NOR2_X1 U8352 ( .A1(n9216), .A2(n9215), .ZN(n40074) );
  NOR2_X2 U8355 ( .A1(n25564), .A2(n25565), .ZN(n37818) );
  NAND3_X2 U8356 ( .A1(n21914), .A2(n31309), .A3(n21911), .ZN(n25564) );
  INV_X1 U8359 ( .I(n20351), .ZN(n6225) );
  NAND2_X1 U8366 ( .A1(n591), .A2(n54960), .ZN(n9097) );
  NOR3_X2 U8367 ( .A1(n6825), .A2(n28234), .A3(n15845), .ZN(n6824) );
  BUF_X4 U8369 ( .I(n34342), .Z(n17538) );
  NAND4_X2 U8370 ( .A1(n26419), .A2(n26420), .A3(n26418), .A4(n26417), .ZN(
        n10124) );
  INV_X2 U8377 ( .I(n53901), .ZN(n54012) );
  NAND2_X1 U8381 ( .A1(n3693), .A2(n37211), .ZN(n3692) );
  INV_X4 U8382 ( .I(n1226), .ZN(n40944) );
  BUF_X4 U8391 ( .I(n4898), .Z(n1233) );
  INV_X1 U8392 ( .I(n31719), .ZN(n24664) );
  NAND2_X1 U8400 ( .A1(n49377), .A2(n3472), .ZN(n3497) );
  NAND2_X1 U8401 ( .A1(n7358), .A2(n3472), .ZN(n49536) );
  OR2_X2 U8413 ( .A1(n19491), .A2(n14848), .Z(n54771) );
  INV_X1 U8415 ( .I(n56408), .ZN(n14601) );
  NAND3_X1 U8416 ( .A1(n56408), .A2(n14307), .A3(n56585), .ZN(n51890) );
  NAND2_X1 U8417 ( .A1(n7680), .A2(n8905), .ZN(n2866) );
  BUF_X2 U8420 ( .I(n23587), .Z(n5118) );
  NAND3_X1 U8424 ( .A1(n61971), .A2(n56815), .A3(n56808), .ZN(n51565) );
  BUF_X2 U8428 ( .I(n14108), .Z(n11577) );
  INV_X2 U8430 ( .I(n2583), .ZN(n16529) );
  BUF_X2 U8431 ( .I(n12049), .Z(n2066) );
  NAND4_X1 U8433 ( .A1(n33819), .A2(n33818), .A3(n24497), .A4(n24496), .ZN(
        n1243) );
  NAND4_X1 U8434 ( .A1(n33819), .A2(n33818), .A3(n24497), .A4(n24496), .ZN(
        n1244) );
  BUF_X2 U8435 ( .I(n33930), .Z(n37940) );
  OAI21_X1 U8440 ( .A1(n24215), .A2(n26065), .B(n50769), .ZN(n8274) );
  NAND2_X1 U8442 ( .A1(n2062), .A2(n51606), .ZN(n54437) );
  BUF_X4 U8463 ( .I(n41675), .Z(n1252) );
  NAND2_X1 U8466 ( .A1(n55342), .A2(n55341), .ZN(n55343) );
  INV_X1 U8472 ( .I(n54243), .ZN(n54264) );
  NAND2_X1 U8475 ( .A1(n55820), .A2(n24958), .ZN(n55819) );
  CLKBUF_X2 U8477 ( .I(n54199), .Z(n9968) );
  CLKBUF_X2 U8483 ( .I(n23116), .Z(n3525) );
  NOR3_X1 U8485 ( .A1(n6465), .A2(n6463), .A3(n54327), .ZN(n6218) );
  NAND2_X1 U8487 ( .A1(n8061), .A2(n8060), .ZN(n8059) );
  NAND2_X1 U8488 ( .A1(n51894), .A2(n24403), .ZN(n4748) );
  NOR2_X1 U8489 ( .A1(n53221), .A2(n61686), .ZN(n12630) );
  AOI22_X1 U8492 ( .A1(n55968), .A2(n55967), .B1(n61182), .B2(n55965), .ZN(
        n6011) );
  OAI21_X1 U8494 ( .A1(n54593), .A2(n7788), .B(n7786), .ZN(n7785) );
  NAND3_X1 U8495 ( .A1(n15929), .A2(n53870), .A3(n63679), .ZN(n13661) );
  NAND4_X1 U8498 ( .A1(n51892), .A2(n11524), .A3(n55927), .A4(n22977), .ZN(
        n51894) );
  OR2_X1 U8499 ( .A1(n55719), .A2(n55908), .Z(n24866) );
  NOR2_X1 U8501 ( .A1(n55679), .A2(n55677), .ZN(n55972) );
  NAND2_X1 U8507 ( .A1(n23110), .A2(n59858), .ZN(n56999) );
  INV_X1 U8509 ( .I(n61572), .ZN(n53231) );
  INV_X1 U8511 ( .I(n53586), .ZN(n1605) );
  INV_X1 U8520 ( .I(n55415), .ZN(n55406) );
  BUF_X2 U8524 ( .I(n50461), .Z(n53859) );
  BUF_X2 U8528 ( .I(n57408), .Z(n26009) );
  OAI21_X1 U8534 ( .A1(n48325), .A2(n5636), .B(n49003), .ZN(n5635) );
  INV_X1 U8539 ( .I(n49951), .ZN(n23459) );
  INV_X1 U8540 ( .I(n9306), .ZN(n13692) );
  NAND3_X1 U8546 ( .A1(n49135), .A2(n60209), .A3(n24134), .ZN(n48266) );
  INV_X1 U8548 ( .I(n4109), .ZN(n50023) );
  INV_X1 U8549 ( .I(n50092), .ZN(n1627) );
  NAND2_X1 U8556 ( .A1(n45231), .A2(n49739), .ZN(n48395) );
  NAND3_X1 U8558 ( .A1(n3239), .A2(n24613), .A3(n57610), .ZN(n3238) );
  NOR3_X1 U8562 ( .A1(n47924), .A2(n12580), .A3(n23707), .ZN(n9925) );
  INV_X1 U8564 ( .I(n22788), .ZN(n48019) );
  NOR3_X1 U8567 ( .A1(n50427), .A2(n78), .A3(n50426), .ZN(n48754) );
  INV_X1 U8569 ( .I(n48431), .ZN(n48801) );
  NAND2_X1 U8570 ( .A1(n78), .A2(n45442), .ZN(n2755) );
  INV_X2 U8572 ( .I(n49529), .ZN(n49543) );
  NOR2_X1 U8577 ( .A1(n49720), .A2(n50096), .ZN(n3030) );
  BUF_X4 U8584 ( .I(n47646), .Z(n49674) );
  NAND2_X1 U8592 ( .A1(n63144), .A2(n59861), .ZN(n11468) );
  AOI22_X1 U8593 ( .A1(n42617), .A2(n23361), .B1(n41979), .B2(n25281), .ZN(
        n25284) );
  NAND2_X1 U8595 ( .A1(n9099), .A2(n48478), .ZN(n7953) );
  OAI21_X1 U8599 ( .A1(n45641), .A2(n45640), .B(n46024), .ZN(n45648) );
  INV_X1 U8600 ( .I(n45654), .ZN(n20861) );
  NAND2_X1 U8601 ( .A1(n45519), .A2(n47468), .ZN(n45744) );
  OAI21_X1 U8602 ( .A1(n47824), .A2(n1295), .B(n47823), .ZN(n12205) );
  NAND2_X1 U8609 ( .A1(n15749), .A2(n9045), .ZN(n9100) );
  INV_X1 U8610 ( .I(n8696), .ZN(n44133) );
  AND3_X1 U8614 ( .A1(n2634), .A2(n59071), .A3(n48481), .Z(n3220) );
  BUF_X1 U8615 ( .I(n2179), .Z(n2178) );
  INV_X2 U8627 ( .I(n21356), .ZN(n1265) );
  INV_X1 U8629 ( .I(n45225), .ZN(n47824) );
  INV_X4 U8639 ( .I(n2686), .ZN(n1268) );
  CLKBUF_X2 U8640 ( .I(n24037), .Z(n11515) );
  AOI22_X1 U8647 ( .A1(n43921), .A2(n43920), .B1(n43918), .B2(n43919), .ZN(
        n43932) );
  NOR2_X1 U8653 ( .A1(n42425), .A2(n7349), .ZN(n40880) );
  NAND3_X1 U8654 ( .A1(n43198), .A2(n43197), .A3(n43516), .ZN(n18673) );
  OAI21_X1 U8656 ( .A1(n15695), .A2(n16864), .B(n279), .ZN(n43918) );
  OR2_X1 U8657 ( .A1(n20067), .A2(n43282), .Z(n4971) );
  OAI22_X1 U8659 ( .A1(n18201), .A2(n13105), .B1(n43607), .B2(n41624), .ZN(
        n41625) );
  NOR3_X1 U8662 ( .A1(n43100), .A2(n24250), .A3(n4659), .ZN(n9447) );
  NOR2_X1 U8665 ( .A1(n42411), .A2(n42965), .ZN(n15120) );
  NAND2_X1 U8667 ( .A1(n43326), .A2(n2496), .ZN(n42196) );
  INV_X1 U8668 ( .I(n42422), .ZN(n21408) );
  NOR2_X1 U8670 ( .A1(n15878), .A2(n41792), .ZN(n41793) );
  INV_X1 U8671 ( .I(n42775), .ZN(n18958) );
  NOR3_X1 U8672 ( .A1(n1392), .A2(n42407), .A3(n21055), .ZN(n3804) );
  INV_X1 U8675 ( .I(n42062), .ZN(n43540) );
  NAND2_X1 U8681 ( .A1(n21851), .A2(n8290), .ZN(n13621) );
  NOR2_X1 U8685 ( .A1(n10617), .A2(n42553), .ZN(n42112) );
  NAND2_X1 U8689 ( .A1(n16982), .A2(n22606), .ZN(n43121) );
  NAND3_X1 U8700 ( .A1(n63464), .A2(n40716), .A3(n60810), .ZN(n38839) );
  AOI21_X1 U8708 ( .A1(n973), .A2(n38045), .B(n967), .ZN(n38048) );
  INV_X1 U8713 ( .I(n5642), .ZN(n20645) );
  OAI22_X1 U8720 ( .A1(n39813), .A2(n64308), .B1(n14985), .B2(n39812), .ZN(
        n24270) );
  AOI21_X1 U8721 ( .A1(n1518), .A2(n40239), .B(n40069), .ZN(n36653) );
  NAND2_X1 U8728 ( .A1(n40696), .A2(n1219), .ZN(n40699) );
  INV_X1 U8729 ( .I(n37532), .ZN(n7649) );
  NAND3_X1 U8730 ( .A1(n4150), .A2(n40064), .A3(n65128), .ZN(n39928) );
  NOR2_X1 U8732 ( .A1(n39066), .A2(n7011), .ZN(n7962) );
  NAND2_X1 U8736 ( .A1(n40661), .A2(n41182), .ZN(n9393) );
  INV_X1 U8742 ( .I(n21791), .ZN(n13050) );
  INV_X1 U8749 ( .I(n40994), .ZN(n40215) );
  BUF_X2 U8752 ( .I(n40666), .Z(n23616) );
  INV_X2 U8753 ( .I(n41474), .ZN(n25131) );
  INV_X2 U8760 ( .I(n25884), .ZN(n41474) );
  INV_X1 U8764 ( .I(n37649), .ZN(n1758) );
  BUF_X1 U8765 ( .I(n37301), .Z(n4422) );
  INV_X1 U8768 ( .I(n13809), .ZN(n13115) );
  NAND2_X2 U8776 ( .A1(n4743), .A2(n11983), .ZN(n38777) );
  NOR4_X1 U8779 ( .A1(n4834), .A2(n37003), .A3(n62734), .A4(n61574), .ZN(
        n34883) );
  OAI21_X1 U8788 ( .A1(n21649), .A2(n33608), .B(n36190), .ZN(n17390) );
  NAND2_X1 U8793 ( .A1(n8363), .A2(n1782), .ZN(n35556) );
  OR2_X1 U8801 ( .A1(n32076), .A2(n37184), .Z(n37007) );
  NAND2_X2 U8804 ( .A1(n1903), .A2(n10067), .ZN(n6612) );
  NOR2_X1 U8811 ( .A1(n4512), .A2(n6540), .ZN(n36825) );
  NOR2_X1 U8815 ( .A1(n7933), .A2(n59379), .ZN(n35958) );
  NAND2_X1 U8825 ( .A1(n9178), .A2(n35886), .ZN(n35888) );
  BUF_X2 U8826 ( .I(n33785), .Z(n36422) );
  BUF_X4 U8827 ( .I(n36960), .Z(n1786) );
  OAI21_X1 U8832 ( .A1(n35631), .A2(n35611), .B(n35202), .ZN(n19198) );
  NOR2_X1 U8833 ( .A1(n35015), .A2(n35014), .ZN(n35016) );
  NOR2_X1 U8834 ( .A1(n35035), .A2(n34635), .ZN(n34651) );
  OAI21_X1 U8841 ( .A1(n14092), .A2(n32965), .B(n5529), .ZN(n32968) );
  OAI21_X1 U8843 ( .A1(n35199), .A2(n35200), .B(n35198), .ZN(n8977) );
  NAND2_X2 U8845 ( .A1(n20068), .A2(n33406), .ZN(n33404) );
  NAND2_X1 U8850 ( .A1(n21699), .A2(n5250), .ZN(n33639) );
  NAND3_X1 U8852 ( .A1(n34040), .A2(n2635), .A3(n33978), .ZN(n31536) );
  INV_X1 U8863 ( .I(n35770), .ZN(n1423) );
  INV_X1 U8868 ( .I(n34566), .ZN(n8552) );
  INV_X1 U8872 ( .I(n32955), .ZN(n34797) );
  INV_X1 U8876 ( .I(n22082), .ZN(n34535) );
  OR2_X1 U8881 ( .A1(n32295), .A2(n21725), .Z(n34953) );
  CLKBUF_X2 U8885 ( .I(n22082), .Z(n19246) );
  BUF_X4 U8888 ( .I(n22699), .Z(n11930) );
  NOR2_X2 U8891 ( .A1(n21413), .A2(n29510), .ZN(n21227) );
  INV_X1 U8892 ( .I(n32266), .ZN(n31487) );
  AOI21_X1 U8898 ( .A1(n61007), .A2(n30591), .B(n4082), .ZN(n27731) );
  CLKBUF_X4 U8899 ( .I(n32183), .Z(n24008) );
  AOI21_X1 U8901 ( .A1(n3899), .A2(n3897), .B(n30647), .ZN(n30336) );
  OAI21_X1 U8906 ( .A1(n30220), .A2(n1869), .B(n22416), .ZN(n2224) );
  INV_X2 U8919 ( .I(n6714), .ZN(n28903) );
  OAI21_X1 U8921 ( .A1(n30546), .A2(n30545), .B(n30544), .ZN(n6818) );
  NOR2_X1 U8924 ( .A1(n8521), .A2(n29235), .ZN(n29832) );
  NAND2_X1 U8928 ( .A1(n30251), .A2(n30046), .ZN(n12162) );
  NAND2_X1 U8931 ( .A1(n30392), .A2(n10068), .ZN(n29499) );
  NOR3_X1 U8932 ( .A1(n29266), .A2(n11205), .A3(n846), .ZN(n9688) );
  NAND3_X1 U8935 ( .A1(n25698), .A2(n11656), .A3(n16631), .ZN(n14109) );
  INV_X2 U8939 ( .I(n25512), .ZN(n1847) );
  NOR2_X1 U8940 ( .A1(n14641), .A2(n14217), .ZN(n14216) );
  NAND2_X1 U8943 ( .A1(n31279), .A2(n31270), .ZN(n31272) );
  NAND2_X1 U8959 ( .A1(n30585), .A2(n1437), .ZN(n29481) );
  NAND2_X1 U8969 ( .A1(n30609), .A2(n30347), .ZN(n22555) );
  BUF_X2 U8970 ( .I(n26740), .Z(n30679) );
  BUF_X2 U8975 ( .I(n30255), .Z(n11656) );
  NOR2_X1 U8977 ( .A1(n14222), .A2(n17725), .ZN(n14221) );
  BUF_X2 U8978 ( .I(n10052), .Z(n4257) );
  BUF_X2 U8979 ( .I(n29576), .Z(n23988) );
  INV_X2 U8992 ( .I(n26268), .ZN(n21151) );
  INV_X1 U8996 ( .I(n26809), .ZN(n29139) );
  NOR2_X1 U8997 ( .A1(n12589), .A2(n28168), .ZN(n29602) );
  INV_X1 U9000 ( .I(n21589), .ZN(n18534) );
  CLKBUF_X2 U9002 ( .I(n16667), .Z(n10419) );
  NAND3_X1 U9005 ( .A1(n1320), .A2(n597), .A3(n6522), .ZN(n27396) );
  INV_X1 U9007 ( .I(n12033), .ZN(n14176) );
  INV_X1 U9017 ( .I(n9940), .ZN(n16667) );
  NOR2_X1 U9019 ( .A1(n27204), .A2(n12221), .ZN(n28339) );
  NAND2_X1 U9022 ( .A1(n29384), .A2(n15893), .ZN(n10603) );
  NAND2_X1 U9024 ( .A1(n5306), .A2(n29171), .ZN(n29166) );
  NAND2_X1 U9026 ( .A1(n23578), .A2(n28128), .ZN(n29287) );
  INV_X1 U9032 ( .I(n5627), .ZN(n29115) );
  INV_X1 U9033 ( .I(n28070), .ZN(n22095) );
  BUF_X1 U9037 ( .I(n27582), .Z(n7477) );
  INV_X2 U9042 ( .I(n26824), .ZN(n27655) );
  NOR2_X1 U9044 ( .A1(n28873), .A2(n29663), .ZN(n27337) );
  INV_X2 U9048 ( .I(n28223), .ZN(n1322) );
  BUF_X2 U9051 ( .I(n39555), .Z(n15707) );
  CLKBUF_X2 U9052 ( .I(n27583), .Z(n22541) );
  BUF_X1 U9054 ( .I(n28376), .Z(n22902) );
  INV_X2 U9056 ( .I(n814), .ZN(n1321) );
  INV_X2 U9057 ( .I(n26531), .ZN(n1279) );
  BUF_X2 U9059 ( .I(n27787), .Z(n15712) );
  INV_X1 U9061 ( .I(n23306), .ZN(n50661) );
  BUF_X2 U9062 ( .I(n26360), .Z(n21132) );
  CLKBUF_X2 U9064 ( .I(n28040), .Z(n23943) );
  CLKBUF_X2 U9067 ( .I(Key[16]), .Z(n53284) );
  BUF_X2 U9069 ( .I(Key[62]), .Z(n54231) );
  CLKBUF_X2 U9070 ( .I(Key[56]), .Z(n54153) );
  BUF_X2 U9071 ( .I(Key[17]), .Z(n53308) );
  BUF_X2 U9076 ( .I(Key[2]), .Z(n53076) );
  CLKBUF_X2 U9077 ( .I(Key[86]), .Z(n54896) );
  CLKBUF_X2 U9080 ( .I(Key[93]), .Z(n4561) );
  CLKBUF_X2 U9081 ( .I(Key[29]), .Z(n53530) );
  BUF_X2 U9082 ( .I(Key[177]), .Z(n52734) );
  AOI22_X1 U9089 ( .A1(n53925), .A2(n53952), .B1(n54013), .B2(n54006), .ZN(
        n53944) );
  NAND2_X1 U9090 ( .A1(n14778), .A2(n61687), .ZN(n57101) );
  AOI21_X1 U9092 ( .A1(n52227), .A2(n53148), .B(n52228), .ZN(n3541) );
  NOR2_X1 U9093 ( .A1(n54192), .A2(n54207), .ZN(n54159) );
  INV_X1 U9096 ( .I(n53148), .ZN(n23153) );
  INV_X1 U9100 ( .I(n20525), .ZN(n53114) );
  NAND2_X1 U9101 ( .A1(n1255), .A2(n62800), .ZN(n56822) );
  INV_X1 U9102 ( .I(n15293), .ZN(n18178) );
  AOI21_X1 U9103 ( .A1(n55629), .A2(n19020), .B(n55641), .ZN(n55649) );
  INV_X1 U9105 ( .I(n11144), .ZN(n56336) );
  BUF_X4 U9107 ( .I(n54238), .Z(n1280) );
  NAND2_X1 U9108 ( .A1(n55752), .A2(n55821), .ZN(n55757) );
  INV_X2 U9109 ( .I(n52248), .ZN(n56942) );
  INV_X1 U9111 ( .I(n53727), .ZN(n14845) );
  NOR2_X1 U9116 ( .A1(n12250), .A2(n23323), .ZN(n25525) );
  NAND2_X1 U9117 ( .A1(n12252), .A2(n12251), .ZN(n12250) );
  OAI21_X1 U9118 ( .A1(n52946), .A2(n61081), .B(n17138), .ZN(n54683) );
  NOR2_X1 U9119 ( .A1(n7268), .A2(n15508), .ZN(n7060) );
  NAND2_X1 U9123 ( .A1(n56234), .A2(n12468), .ZN(n52691) );
  NAND2_X1 U9124 ( .A1(n55284), .A2(n15315), .ZN(n15314) );
  INV_X1 U9126 ( .I(n19971), .ZN(n55488) );
  NAND2_X1 U9127 ( .A1(n53231), .A2(n21561), .ZN(n12252) );
  NOR2_X1 U9129 ( .A1(n13794), .A2(n13793), .ZN(n13792) );
  NOR2_X1 U9131 ( .A1(n20740), .A2(n17499), .ZN(n7347) );
  INV_X1 U9132 ( .I(n54956), .ZN(n19499) );
  NOR2_X1 U9133 ( .A1(n52124), .A2(n19644), .ZN(n9489) );
  INV_X1 U9135 ( .I(n55976), .ZN(n14139) );
  NAND2_X1 U9136 ( .A1(n11989), .A2(n56282), .ZN(n56394) );
  INV_X1 U9139 ( .I(n52844), .ZN(n53382) );
  INV_X2 U9144 ( .I(n55966), .ZN(n55974) );
  INV_X1 U9146 ( .I(n52820), .ZN(n57042) );
  NAND2_X1 U9150 ( .A1(n65282), .A2(n53858), .ZN(n22884) );
  NOR2_X1 U9151 ( .A1(n53428), .A2(n53860), .ZN(n53620) );
  NOR2_X1 U9153 ( .A1(n55415), .A2(n55404), .ZN(n8395) );
  AND2_X1 U9154 ( .A1(n56627), .A2(n56631), .Z(n51110) );
  INV_X1 U9157 ( .I(n13774), .ZN(n25232) );
  INV_X1 U9163 ( .I(n51973), .ZN(n25098) );
  INV_X1 U9164 ( .I(n25568), .ZN(n51553) );
  INV_X1 U9166 ( .I(n18485), .ZN(n51757) );
  INV_X2 U9173 ( .I(n52627), .ZN(n1289) );
  NOR2_X1 U9176 ( .A1(n49011), .A2(n5629), .ZN(n44410) );
  NAND3_X1 U9177 ( .A1(n6897), .A2(n49260), .A3(n6896), .ZN(n6895) );
  NAND3_X1 U9180 ( .A1(n23650), .A2(n49722), .A3(n1627), .ZN(n25605) );
  AOI21_X1 U9186 ( .A1(n49450), .A2(n49846), .B(n49843), .ZN(n14860) );
  NAND2_X1 U9193 ( .A1(n13537), .A2(n50216), .ZN(n5188) );
  INV_X1 U9194 ( .I(n48972), .ZN(n15154) );
  NOR2_X1 U9197 ( .A1(n62413), .A2(n49345), .ZN(n50011) );
  INV_X1 U9198 ( .I(n48418), .ZN(n26104) );
  NAND3_X1 U9200 ( .A1(n50402), .A2(n50404), .A3(n50403), .ZN(n7156) );
  OAI21_X1 U9202 ( .A1(n3238), .A2(n16595), .B(n3236), .ZN(n3235) );
  NAND2_X1 U9206 ( .A1(n19523), .A2(n19379), .ZN(n19172) );
  NAND2_X1 U9208 ( .A1(n9594), .A2(n49493), .ZN(n4719) );
  INV_X2 U9209 ( .I(n16985), .ZN(n1633) );
  NAND2_X1 U9211 ( .A1(n15021), .A2(n6130), .ZN(n15635) );
  CLKBUF_X2 U9213 ( .I(n49529), .Z(n9983) );
  NOR2_X1 U9216 ( .A1(n20004), .A2(n49177), .ZN(n11794) );
  INV_X1 U9218 ( .I(n14516), .ZN(n16107) );
  BUF_X2 U9219 ( .I(n45160), .Z(n49698) );
  INV_X2 U9220 ( .I(n49166), .ZN(n49170) );
  NAND2_X1 U9221 ( .A1(n49748), .A2(n49739), .ZN(n49222) );
  NAND2_X1 U9223 ( .A1(n49673), .A2(n48711), .ZN(n49092) );
  BUF_X4 U9225 ( .I(n46047), .Z(n49767) );
  NOR2_X1 U9242 ( .A1(n47691), .A2(n57852), .ZN(n15553) );
  INV_X1 U9244 ( .I(n24820), .ZN(n1651) );
  NAND2_X1 U9247 ( .A1(n47209), .A2(n47208), .ZN(n8134) );
  NOR3_X1 U9248 ( .A1(n508), .A2(n23643), .A3(n24359), .ZN(n44645) );
  NAND2_X1 U9250 ( .A1(n47210), .A2(n15749), .ZN(n8136) );
  NAND2_X1 U9258 ( .A1(n17573), .A2(n48234), .ZN(n48535) );
  INV_X1 U9267 ( .I(n47487), .ZN(n48660) );
  NOR2_X1 U9271 ( .A1(n13746), .A2(n45992), .ZN(n47243) );
  AND2_X1 U9272 ( .A1(n46986), .A2(n2828), .Z(n2827) );
  NOR2_X1 U9273 ( .A1(n47435), .A2(n24252), .ZN(n47732) );
  INV_X2 U9275 ( .I(n5803), .ZN(n1293) );
  NAND2_X1 U9284 ( .A1(n21650), .A2(n13870), .ZN(n13869) );
  INV_X1 U9288 ( .I(n25926), .ZN(n46212) );
  CLKBUF_X2 U9289 ( .I(n8481), .Z(n8480) );
  BUF_X2 U9290 ( .I(n12608), .Z(n12607) );
  INV_X1 U9294 ( .I(n41708), .ZN(n9031) );
  NAND2_X1 U9301 ( .A1(n43118), .A2(n21408), .ZN(n3007) );
  OAI22_X1 U9302 ( .A1(n26187), .A2(n4659), .B1(n8678), .B2(n43225), .ZN(
        n26186) );
  NAND2_X1 U9304 ( .A1(n43282), .A2(n23700), .ZN(n43283) );
  NAND3_X1 U9306 ( .A1(n41727), .A2(n41726), .A3(n41725), .ZN(n41728) );
  NAND3_X1 U9309 ( .A1(n9440), .A2(n43250), .A3(n760), .ZN(n2011) );
  OAI22_X1 U9311 ( .A1(n43953), .A2(n11986), .B1(n16890), .B2(n16911), .ZN(
        n43954) );
  NOR2_X1 U9312 ( .A1(n42339), .A2(n1391), .ZN(n11018) );
  OR2_X1 U9315 ( .A1(n16377), .A2(n19454), .Z(n11366) );
  INV_X2 U9331 ( .I(n6995), .ZN(n1333) );
  NOR2_X1 U9344 ( .A1(n21073), .A2(n43778), .ZN(n42062) );
  NAND2_X1 U9345 ( .A1(n11476), .A2(n42008), .ZN(n15674) );
  BUF_X2 U9361 ( .I(n5971), .Z(n22087) );
  NOR2_X1 U9362 ( .A1(n19241), .A2(n25534), .ZN(n41693) );
  BUF_X4 U9378 ( .I(n42356), .Z(n1301) );
  OAI21_X1 U9383 ( .A1(n3976), .A2(n38344), .B(n42275), .ZN(n11082) );
  AND2_X1 U9384 ( .A1(n14916), .A2(n41312), .Z(n7356) );
  NAND4_X1 U9389 ( .A1(n3109), .A2(n22593), .A3(n40206), .A4(n40207), .ZN(
        n40208) );
  NOR3_X1 U9391 ( .A1(n11096), .A2(n9894), .A3(n17095), .ZN(n3976) );
  NOR3_X1 U9405 ( .A1(n41168), .A2(n7963), .A3(n7962), .ZN(n11385) );
  NAND3_X1 U9407 ( .A1(n40271), .A2(n20047), .A3(n25921), .ZN(n8441) );
  INV_X1 U9411 ( .I(n40500), .ZN(n3612) );
  INV_X1 U9412 ( .I(n40301), .ZN(n40139) );
  INV_X2 U9415 ( .I(n971), .ZN(n1732) );
  INV_X1 U9418 ( .I(n38496), .ZN(n21736) );
  NAND2_X1 U9419 ( .A1(n41401), .A2(n14165), .ZN(n41410) );
  NAND3_X1 U9420 ( .A1(n40523), .A2(n40614), .A3(n23787), .ZN(n40622) );
  INV_X1 U9423 ( .I(n40314), .ZN(n41817) );
  NAND2_X1 U9428 ( .A1(n17450), .A2(n60957), .ZN(n2004) );
  INV_X1 U9430 ( .I(n40413), .ZN(n40753) );
  OR2_X1 U9439 ( .A1(n40995), .A2(n40994), .Z(n6766) );
  NOR2_X1 U9444 ( .A1(n21207), .A2(n42432), .ZN(n4150) );
  INV_X2 U9445 ( .I(n42479), .ZN(n1515) );
  INV_X2 U9453 ( .I(n40644), .ZN(n7011) );
  INV_X2 U9455 ( .I(n11437), .ZN(n1307) );
  INV_X1 U9456 ( .I(n39710), .ZN(n39534) );
  NOR2_X1 U9460 ( .A1(n36902), .A2(n36901), .ZN(n37649) );
  INV_X1 U9462 ( .I(n38469), .ZN(n24533) );
  BUF_X2 U9467 ( .I(n20042), .Z(n20041) );
  NAND3_X1 U9471 ( .A1(n25591), .A2(n35365), .A3(n35364), .ZN(n25590) );
  NAND3_X1 U9476 ( .A1(n35555), .A2(n35556), .A3(n36487), .ZN(n16605) );
  INV_X1 U9478 ( .I(n37092), .ZN(n36642) );
  NOR2_X1 U9479 ( .A1(n4834), .A2(n37007), .ZN(n23750) );
  NAND3_X1 U9485 ( .A1(n10087), .A2(n2592), .A3(n11077), .ZN(n36523) );
  OAI21_X1 U9486 ( .A1(n37370), .A2(n37371), .B(n61704), .ZN(n14341) );
  NAND4_X1 U9487 ( .A1(n24118), .A2(n35900), .A3(n23584), .A4(n35901), .ZN(
        n14925) );
  NAND4_X1 U9499 ( .A1(n1777), .A2(n15171), .A3(n2792), .A4(n34927), .ZN(n2791) );
  OAI21_X1 U9501 ( .A1(n34470), .A2(n59229), .B(n2775), .ZN(n34471) );
  INV_X1 U9502 ( .I(n37408), .ZN(n35918) );
  NOR2_X1 U9503 ( .A1(n61574), .A2(n8010), .ZN(n35877) );
  NOR2_X1 U9506 ( .A1(n36835), .A2(n6984), .ZN(n35914) );
  AOI22_X1 U9508 ( .A1(n11027), .A2(n9041), .B1(n22559), .B2(n36262), .ZN(
        n11031) );
  OAI21_X1 U9513 ( .A1(n25396), .A2(n25964), .B(n1416), .ZN(n36865) );
  OAI21_X1 U9514 ( .A1(n7488), .A2(n24118), .B(n23584), .ZN(n35174) );
  NAND2_X1 U9516 ( .A1(n13983), .A2(n12652), .ZN(n35437) );
  NAND2_X1 U9518 ( .A1(n36427), .A2(n36422), .ZN(n36179) );
  NOR2_X1 U9524 ( .A1(n1785), .A2(n64405), .ZN(n36379) );
  NAND2_X2 U9534 ( .A1(n21780), .A2(n21781), .ZN(n35990) );
  NOR2_X1 U9539 ( .A1(n2399), .A2(n2398), .ZN(n2397) );
  OR2_X1 U9550 ( .A1(n17148), .A2(n35305), .Z(n21485) );
  NAND4_X1 U9555 ( .A1(n34334), .A2(n35775), .A3(n35770), .A4(n32132), .ZN(
        n32135) );
  NAND3_X1 U9568 ( .A1(n11477), .A2(n8694), .A3(n65189), .ZN(n34555) );
  NOR3_X1 U9571 ( .A1(n60819), .A2(n1541), .A3(n34414), .ZN(n12937) );
  INV_X1 U9572 ( .I(n7661), .ZN(n33774) );
  NOR2_X1 U9574 ( .A1(n8051), .A2(n35762), .ZN(n16203) );
  NAND3_X1 U9581 ( .A1(n24077), .A2(n2208), .A3(n35026), .ZN(n34557) );
  OAI21_X1 U9582 ( .A1(n18077), .A2(n1345), .B(n1545), .ZN(n12167) );
  INV_X1 U9583 ( .I(n35786), .ZN(n34334) );
  INV_X1 U9584 ( .I(n32796), .ZN(n20524) );
  CLKBUF_X2 U9589 ( .I(n24331), .Z(n11659) );
  INV_X1 U9596 ( .I(n14111), .ZN(n14112) );
  BUF_X2 U9598 ( .I(n32017), .Z(n35301) );
  INV_X1 U9599 ( .I(n34317), .ZN(n21487) );
  INV_X1 U9601 ( .I(n23714), .ZN(n12013) );
  CLKBUF_X2 U9602 ( .I(n23491), .Z(n2259) );
  INV_X2 U9603 ( .I(n22652), .ZN(n33838) );
  BUF_X1 U9604 ( .I(n60466), .Z(n4663) );
  BUF_X2 U9605 ( .I(n22751), .Z(n9609) );
  INV_X1 U9610 ( .I(n20719), .ZN(n1833) );
  NAND3_X1 U9614 ( .A1(n30390), .A2(n5343), .A3(n29499), .ZN(n27639) );
  NAND2_X1 U9616 ( .A1(n12161), .A2(n4889), .ZN(n2021) );
  NAND3_X1 U9618 ( .A1(n3987), .A2(n3986), .A3(n3984), .ZN(n3983) );
  AOI22_X1 U9621 ( .A1(n3992), .A2(n12743), .B1(n22322), .B2(n3991), .ZN(n3990) );
  AND2_X1 U9622 ( .A1(n61849), .A2(n30888), .Z(n5799) );
  NOR2_X1 U9624 ( .A1(n30049), .A2(n30250), .ZN(n2280) );
  NOR2_X1 U9625 ( .A1(n29421), .A2(n30455), .ZN(n29425) );
  NOR2_X1 U9629 ( .A1(n10151), .A2(n29481), .ZN(n30591) );
  NAND3_X1 U9631 ( .A1(n31030), .A2(n12871), .A3(n31031), .ZN(n3992) );
  NAND2_X1 U9639 ( .A1(n24949), .A2(n29506), .ZN(n28704) );
  OAI22_X1 U9640 ( .A1(n29041), .A2(n29221), .B1(n30288), .B2(n30284), .ZN(
        n17337) );
  NAND2_X1 U9643 ( .A1(n30449), .A2(n30455), .ZN(n18635) );
  OAI21_X1 U9644 ( .A1(n18326), .A2(n30251), .B(n1349), .ZN(n18325) );
  NAND2_X1 U9647 ( .A1(n22748), .A2(n13176), .ZN(n30028) );
  INV_X1 U9652 ( .I(n30250), .ZN(n1841) );
  NAND2_X1 U9653 ( .A1(n30170), .A2(n58999), .ZN(n13481) );
  NOR2_X1 U9655 ( .A1(n1856), .A2(n10734), .ZN(n30384) );
  AND2_X1 U9656 ( .A1(n13766), .A2(n58747), .Z(n13765) );
  OAI21_X1 U9659 ( .A1(n28904), .A2(n30487), .B(n28905), .ZN(n5864) );
  NAND3_X1 U9660 ( .A1(n1436), .A2(n19255), .A3(n58621), .ZN(n31259) );
  AND2_X1 U9664 ( .A1(n30324), .A2(n2119), .Z(n2118) );
  NOR2_X1 U9665 ( .A1(n30331), .A2(n60202), .ZN(n3902) );
  NAND3_X1 U9666 ( .A1(n3426), .A2(n1869), .A3(n16808), .ZN(n9001) );
  NOR2_X1 U9668 ( .A1(n22230), .A2(n61421), .ZN(n29838) );
  NAND2_X1 U9672 ( .A1(n29959), .A2(n29747), .ZN(n30788) );
  NAND2_X1 U9675 ( .A1(n29440), .A2(n25096), .ZN(n31124) );
  NAND2_X1 U9677 ( .A1(n17872), .A2(n60111), .ZN(n31046) );
  INV_X2 U9685 ( .I(n58710), .ZN(n9250) );
  INV_X2 U9687 ( .I(n23569), .ZN(n24728) );
  CLKBUF_X2 U9688 ( .I(n21832), .Z(n10129) );
  INV_X2 U9692 ( .I(n6349), .ZN(n22322) );
  NAND2_X1 U9693 ( .A1(n30338), .A2(n30347), .ZN(n30614) );
  BUF_X2 U9695 ( .I(n22374), .Z(n18198) );
  INV_X1 U9696 ( .I(n30224), .ZN(n1555) );
  NAND2_X1 U9702 ( .A1(n15689), .A2(n29580), .ZN(n29267) );
  INV_X2 U9705 ( .I(n30580), .ZN(n12051) );
  INV_X4 U9706 ( .I(n847), .ZN(n1316) );
  INV_X4 U9711 ( .I(n28426), .ZN(n1317) );
  INV_X2 U9714 ( .I(n15533), .ZN(n29244) );
  OAI21_X1 U9718 ( .A1(n27164), .A2(n9088), .B(n19113), .ZN(n27240) );
  NAND3_X1 U9721 ( .A1(n28874), .A2(n28871), .A3(n5659), .ZN(n10920) );
  NAND2_X1 U9726 ( .A1(n2513), .A2(n3910), .ZN(n29113) );
  INV_X1 U9727 ( .I(n26524), .ZN(n4059) );
  AND2_X1 U9728 ( .A1(n28231), .A2(n14583), .Z(n14581) );
  NAND2_X1 U9733 ( .A1(n27693), .A2(n29600), .ZN(n27695) );
  INV_X1 U9735 ( .I(n31318), .ZN(n31397) );
  NOR2_X1 U9737 ( .A1(n16525), .A2(n28494), .ZN(n26398) );
  NAND2_X1 U9738 ( .A1(n28510), .A2(n7110), .ZN(n26423) );
  NAND2_X1 U9739 ( .A1(n29134), .A2(n7371), .ZN(n26809) );
  INV_X1 U9744 ( .I(n27037), .ZN(n28238) );
  NOR2_X1 U9747 ( .A1(n29144), .A2(n16654), .ZN(n27296) );
  AND2_X1 U9748 ( .A1(n29127), .A2(n57954), .Z(n11510) );
  NAND3_X1 U9751 ( .A1(n8518), .A2(n64445), .A3(n8359), .ZN(n12033) );
  INV_X1 U9757 ( .I(n29156), .ZN(n29149) );
  INV_X1 U9759 ( .I(n28300), .ZN(n28310) );
  INV_X1 U9760 ( .I(n28616), .ZN(n10085) );
  INV_X1 U9763 ( .I(n27414), .ZN(n29163) );
  NOR2_X1 U9764 ( .A1(n29141), .A2(n29145), .ZN(n2662) );
  INV_X1 U9765 ( .I(n20734), .ZN(n28397) );
  NOR2_X1 U9766 ( .A1(n29671), .A2(n28873), .ZN(n29384) );
  AND2_X1 U9767 ( .A1(n28066), .A2(n28072), .Z(n26529) );
  INV_X2 U9770 ( .I(n60505), .ZN(n27387) );
  INV_X2 U9771 ( .I(n20240), .ZN(n1363) );
  INV_X2 U9772 ( .I(n19279), .ZN(n1362) );
  BUF_X2 U9773 ( .I(n30355), .Z(n15710) );
  BUF_X2 U9774 ( .I(n26334), .Z(n27171) );
  NAND2_X1 U9775 ( .A1(n25202), .A2(n26720), .ZN(n12707) );
  INV_X1 U9778 ( .I(n53375), .ZN(n1448) );
  INV_X1 U9779 ( .I(n28303), .ZN(n20437) );
  INV_X1 U9780 ( .I(n53284), .ZN(n1574) );
  CLKBUF_X2 U9781 ( .I(Key[54]), .Z(n54126) );
  CLKBUF_X2 U9784 ( .I(Key[7]), .Z(n50817) );
  CLKBUF_X2 U9785 ( .I(Key[74]), .Z(n54536) );
  CLKBUF_X2 U9786 ( .I(Key[23]), .Z(n53375) );
  CLKBUF_X2 U9787 ( .I(Key[159]), .Z(n56495) );
  AOI21_X1 U9789 ( .A1(n56319), .A2(n11921), .B(n11920), .ZN(n11919) );
  INV_X1 U9791 ( .I(n2746), .ZN(n53668) );
  CLKBUF_X2 U9794 ( .I(n2851), .Z(n9715) );
  NAND2_X1 U9795 ( .A1(n56851), .A2(n60708), .ZN(n52731) );
  OAI22_X1 U9796 ( .A1(n56822), .A2(n12454), .B1(n56895), .B2(n22667), .ZN(
        n17361) );
  OAI21_X1 U9798 ( .A1(n53800), .A2(n53820), .B(n53807), .ZN(n26218) );
  OAI21_X1 U9799 ( .A1(n53346), .A2(n53347), .B(n53345), .ZN(n53364) );
  AND3_X1 U9802 ( .A1(n17961), .A2(n56145), .A3(n56191), .Z(n51259) );
  NAND2_X1 U9804 ( .A1(n11622), .A2(n1367), .ZN(n6091) );
  NAND2_X1 U9806 ( .A1(n56942), .A2(n56958), .ZN(n21370) );
  BUF_X4 U9807 ( .I(n52041), .Z(n55893) );
  NOR2_X1 U9824 ( .A1(n24957), .A2(n55669), .ZN(n24960) );
  NOR2_X1 U9828 ( .A1(n55488), .A2(n55296), .ZN(n9913) );
  NOR2_X1 U9831 ( .A1(n23025), .A2(n58300), .ZN(n7332) );
  NAND2_X1 U9834 ( .A1(n56273), .A2(n58050), .ZN(n23845) );
  NOR3_X1 U9835 ( .A1(n56999), .A2(n5684), .A3(n20921), .ZN(n24424) );
  NAND2_X1 U9842 ( .A1(n17601), .A2(n55906), .ZN(n17027) );
  AOI21_X1 U9843 ( .A1(n11524), .A2(n22977), .B(n11177), .ZN(n11176) );
  OR2_X1 U9846 ( .A1(n12692), .A2(n1373), .Z(n15822) );
  INV_X2 U9847 ( .I(n22804), .ZN(n1369) );
  INV_X1 U9848 ( .I(n55404), .ZN(n54786) );
  INV_X1 U9849 ( .I(n55905), .ZN(n1595) );
  INV_X1 U9851 ( .I(n3567), .ZN(n55681) );
  INV_X1 U9854 ( .I(n55685), .ZN(n1609) );
  NAND2_X1 U9855 ( .A1(n13232), .A2(n1287), .ZN(n52820) );
  INV_X4 U9858 ( .I(n52126), .ZN(n1324) );
  INV_X4 U9861 ( .I(n54640), .ZN(n1373) );
  INV_X2 U9862 ( .I(n26228), .ZN(n1326) );
  BUF_X2 U9865 ( .I(n23852), .Z(n16691) );
  INV_X1 U9866 ( .I(n52604), .ZN(n2060) );
  NOR2_X1 U9868 ( .A1(n1624), .A2(n49978), .ZN(n49982) );
  OAI22_X1 U9872 ( .A1(n14860), .A2(n49849), .B1(n49452), .B2(n49451), .ZN(
        n14859) );
  NOR2_X1 U9875 ( .A1(n50284), .A2(n48721), .ZN(n15130) );
  AOI21_X1 U9879 ( .A1(n48958), .A2(n49260), .B(n47058), .ZN(n12675) );
  NAND2_X1 U9882 ( .A1(n49390), .A2(n49393), .ZN(n48873) );
  NAND3_X1 U9883 ( .A1(n48853), .A2(n59838), .A3(n49491), .ZN(n6119) );
  NOR2_X1 U9885 ( .A1(n49278), .A2(n16411), .ZN(n11415) );
  NOR2_X1 U9887 ( .A1(n49111), .A2(n59493), .ZN(n49113) );
  NAND2_X1 U9888 ( .A1(n44409), .A2(n48323), .ZN(n14401) );
  NAND2_X1 U9896 ( .A1(n16411), .A2(n49287), .ZN(n48919) );
  AOI21_X1 U9898 ( .A1(n12701), .A2(n48391), .B(n6704), .ZN(n6118) );
  NAND2_X1 U9901 ( .A1(n60520), .A2(n61867), .ZN(n15357) );
  NAND3_X1 U9902 ( .A1(n12580), .A2(n61355), .A3(n50093), .ZN(n12629) );
  NAND2_X1 U9904 ( .A1(n50094), .A2(n50376), .ZN(n50095) );
  OAI22_X1 U9909 ( .A1(n11246), .A2(n13554), .B1(n48682), .B2(n2810), .ZN(
        n6227) );
  NOR2_X1 U9917 ( .A1(n50218), .A2(n14335), .ZN(n14516) );
  AOI21_X1 U9924 ( .A1(n58244), .A2(n64960), .B(n46949), .ZN(n6662) );
  NOR2_X1 U9926 ( .A1(n48242), .A2(n47487), .ZN(n16416) );
  NAND2_X1 U9928 ( .A1(n46814), .A2(n2955), .ZN(n11692) );
  OAI21_X1 U9931 ( .A1(n46760), .A2(n46759), .B(n46814), .ZN(n46761) );
  NAND3_X1 U9932 ( .A1(n45525), .A2(n45744), .A3(n45524), .ZN(n26045) );
  OAI21_X1 U9933 ( .A1(n57234), .A2(n58244), .B(n45506), .ZN(n45507) );
  OR2_X1 U9935 ( .A1(n47898), .A2(n45941), .Z(n4352) );
  NAND3_X1 U9936 ( .A1(n43751), .A2(n47735), .A3(n11821), .ZN(n43754) );
  NOR2_X1 U9941 ( .A1(n1263), .A2(n47422), .ZN(n46845) );
  OAI22_X1 U9942 ( .A1(n48250), .A2(n17153), .B1(n48249), .B2(n1476), .ZN(
        n3358) );
  NAND2_X1 U9945 ( .A1(n48246), .A2(n47481), .ZN(n48247) );
  OAI21_X1 U9946 ( .A1(n47243), .A2(n47244), .B(n47615), .ZN(n8649) );
  INV_X1 U9947 ( .I(n11087), .ZN(n46760) );
  NAND2_X1 U9950 ( .A1(n64791), .A2(n7834), .ZN(n21855) );
  NOR2_X1 U9952 ( .A1(n7335), .A2(n64791), .ZN(n48646) );
  INV_X1 U9956 ( .I(n48571), .ZN(n1650) );
  INV_X1 U9958 ( .I(n15748), .ZN(n47377) );
  OAI21_X1 U9960 ( .A1(n60839), .A2(n47487), .B(n48654), .ZN(n17805) );
  NAND3_X1 U9962 ( .A1(n48624), .A2(n48623), .A3(n48620), .ZN(n46364) );
  CLKBUF_X2 U9967 ( .I(n47036), .Z(n23903) );
  INV_X4 U9973 ( .I(n23407), .ZN(n1328) );
  INV_X4 U9975 ( .I(n20344), .ZN(n48148) );
  BUF_X2 U9978 ( .I(n14782), .Z(n13069) );
  INV_X1 U9979 ( .I(n23118), .ZN(n45852) );
  BUF_X2 U9980 ( .I(n44162), .Z(n25872) );
  INV_X2 U9987 ( .I(n5431), .ZN(n1330) );
  BUF_X2 U9991 ( .I(n46446), .Z(n22207) );
  NOR3_X1 U10003 ( .A1(n43954), .A2(n43949), .A3(n25670), .ZN(n11405) );
  NOR2_X1 U10004 ( .A1(n42847), .A2(n15007), .ZN(n15063) );
  NAND2_X1 U10006 ( .A1(n1687), .A2(n12677), .ZN(n43296) );
  NAND3_X1 U10008 ( .A1(n43283), .A2(n18172), .A3(n2735), .ZN(n43284) );
  NAND3_X1 U10010 ( .A1(n18723), .A2(n1299), .A3(n16890), .ZN(n43298) );
  NAND2_X1 U10017 ( .A1(n23838), .A2(n1491), .ZN(n6901) );
  OAI22_X1 U10019 ( .A1(n43737), .A2(n43738), .B1(n43736), .B2(n43735), .ZN(
        n16607) );
  NAND2_X1 U10024 ( .A1(n15252), .A2(n61739), .ZN(n12775) );
  NOR2_X1 U10034 ( .A1(n42915), .A2(n10415), .ZN(n13162) );
  NAND3_X1 U10035 ( .A1(n7451), .A2(n11606), .A3(n1709), .ZN(n3956) );
  NOR3_X1 U10036 ( .A1(n8687), .A2(n43272), .A3(n43270), .ZN(n4328) );
  NAND2_X1 U10037 ( .A1(n43889), .A2(n11635), .ZN(n43142) );
  OR2_X1 U10040 ( .A1(n20650), .A2(n59682), .Z(n42099) );
  INV_X4 U10044 ( .I(n42894), .ZN(n11179) );
  NAND3_X1 U10045 ( .A1(n62546), .A2(n3674), .A3(n59309), .ZN(n42932) );
  BUF_X2 U10050 ( .I(n15029), .Z(n3674) );
  INV_X4 U10067 ( .I(n18126), .ZN(n1335) );
  BUF_X4 U10068 ( .I(n19537), .Z(n5939) );
  INV_X2 U10071 ( .I(n9135), .ZN(n11609) );
  NAND2_X1 U10084 ( .A1(n15008), .A2(n15072), .ZN(n41634) );
  AOI21_X1 U10087 ( .A1(n40053), .A2(n40107), .B(n7695), .ZN(n40059) );
  NOR2_X1 U10092 ( .A1(n40267), .A2(n40329), .ZN(n8442) );
  NAND3_X1 U10093 ( .A1(n42200), .A2(n60947), .A3(n41870), .ZN(n42205) );
  OAI21_X1 U10094 ( .A1(n40209), .A2(n11494), .B(n40208), .ZN(n26159) );
  OAI21_X1 U10098 ( .A1(n41241), .A2(n39857), .B(n41405), .ZN(n39858) );
  OAI21_X1 U10100 ( .A1(n25627), .A2(n39323), .B(n57955), .ZN(n18526) );
  OAI21_X1 U10109 ( .A1(n18421), .A2(n40441), .B(n18420), .ZN(n18413) );
  NOR2_X1 U10111 ( .A1(n38679), .A2(n40636), .ZN(n38680) );
  NAND3_X1 U10112 ( .A1(n12057), .A2(n5642), .A3(n287), .ZN(n42254) );
  NAND2_X1 U10115 ( .A1(n41462), .A2(n41155), .ZN(n18594) );
  NOR2_X1 U10119 ( .A1(n41054), .A2(n11895), .ZN(n40848) );
  NAND3_X1 U10124 ( .A1(n8440), .A2(n25511), .A3(n40106), .ZN(n8439) );
  NAND2_X1 U10125 ( .A1(n41013), .A2(n1511), .ZN(n41026) );
  OAI21_X1 U10126 ( .A1(n16962), .A2(n12284), .B(n40057), .ZN(n12286) );
  NOR2_X1 U10130 ( .A1(n61394), .A2(n41951), .ZN(n5788) );
  NOR2_X1 U10136 ( .A1(n3245), .A2(n64793), .ZN(n15496) );
  INV_X1 U10139 ( .I(n40217), .ZN(n38040) );
  NAND2_X1 U10142 ( .A1(n19438), .A2(n60971), .ZN(n19726) );
  NOR2_X1 U10143 ( .A1(n41183), .A2(n1404), .ZN(n11194) );
  NAND2_X1 U10144 ( .A1(n36996), .A2(n40146), .ZN(n6751) );
  NAND2_X1 U10147 ( .A1(n40272), .A2(n57536), .ZN(n40271) );
  INV_X1 U10148 ( .I(n39821), .ZN(n1724) );
  CLKBUF_X2 U10149 ( .I(n42465), .Z(n9798) );
  AND2_X1 U10150 ( .A1(n39973), .A2(n41079), .Z(n16159) );
  NOR2_X1 U10151 ( .A1(n41444), .A2(n40695), .ZN(n15440) );
  NAND2_X1 U10154 ( .A1(n39905), .A2(n41306), .ZN(n41308) );
  OR2_X1 U10157 ( .A1(n41077), .A2(n64475), .Z(n3282) );
  INV_X1 U10159 ( .I(n23711), .ZN(n1736) );
  OAI21_X1 U10160 ( .A1(n14132), .A2(n40592), .B(n7907), .ZN(n4359) );
  INV_X1 U10166 ( .I(n64242), .ZN(n21255) );
  INV_X1 U10167 ( .I(n41870), .ZN(n42202) );
  NOR2_X1 U10169 ( .A1(n41877), .A2(n41054), .ZN(n41061) );
  CLKBUF_X2 U10172 ( .I(n41158), .Z(n22380) );
  OR2_X1 U10182 ( .A1(n25976), .A2(n40697), .Z(n15441) );
  CLKBUF_X2 U10187 ( .I(n22653), .Z(n11459) );
  OR2_X2 U10188 ( .A1(n25884), .A2(n25132), .Z(n40417) );
  BUF_X2 U10195 ( .I(n21289), .Z(n16476) );
  INV_X1 U10202 ( .I(n24533), .ZN(n1759) );
  BUF_X2 U10205 ( .I(n15247), .Z(n15246) );
  INV_X1 U10211 ( .I(n36878), .ZN(n4831) );
  AOI22_X1 U10214 ( .A1(n12831), .A2(n36415), .B1(n22474), .B2(n36411), .ZN(
        n13929) );
  AND3_X1 U10215 ( .A1(n34881), .A2(n37003), .A3(n37326), .Z(n8680) );
  OAI21_X1 U10227 ( .A1(n35877), .A2(n2942), .B(n37009), .ZN(n16530) );
  AOI21_X1 U10229 ( .A1(n37291), .A2(n37290), .B(n37289), .ZN(n37850) );
  OAI21_X1 U10233 ( .A1(n24370), .A2(n37084), .B(n13666), .ZN(n37092) );
  AOI22_X1 U10234 ( .A1(n34362), .A2(n34837), .B1(n18984), .B2(n34361), .ZN(
        n16735) );
  NOR2_X1 U10238 ( .A1(n36173), .A2(n36427), .ZN(n36123) );
  OR2_X1 U10245 ( .A1(n3458), .A2(n2059), .Z(n6883) );
  NAND2_X1 U10250 ( .A1(n25125), .A2(n36262), .ZN(n11029) );
  NAND2_X1 U10251 ( .A1(n36584), .A2(n798), .ZN(n11143) );
  NAND2_X1 U10255 ( .A1(n58220), .A2(n8177), .ZN(n34289) );
  NOR2_X1 U10262 ( .A1(n1414), .A2(n4304), .ZN(n2775) );
  OR3_X1 U10265 ( .A1(n19368), .A2(n37125), .A3(n57860), .Z(n20382) );
  OR2_X2 U10266 ( .A1(n9178), .A2(n35173), .Z(n7802) );
  NAND2_X1 U10267 ( .A1(n1416), .A2(n25396), .ZN(n35930) );
  NOR2_X1 U10270 ( .A1(n37209), .A2(n23357), .ZN(n36618) );
  NOR2_X1 U10275 ( .A1(n12141), .A2(n36777), .ZN(n36766) );
  NAND2_X1 U10278 ( .A1(n36171), .A2(n36427), .ZN(n33786) );
  NAND2_X1 U10280 ( .A1(n25964), .A2(n1416), .ZN(n37390) );
  NAND2_X1 U10281 ( .A1(n26147), .A2(n10717), .ZN(n36763) );
  BUF_X2 U10283 ( .I(n35990), .Z(n22892) );
  INV_X1 U10284 ( .I(n33933), .ZN(n1783) );
  NOR2_X1 U10287 ( .A1(n24180), .A2(n11319), .ZN(n6054) );
  BUF_X2 U10290 ( .I(n36451), .Z(n23257) );
  OR2_X1 U10293 ( .A1(n24805), .A2(n8049), .Z(n8050) );
  NOR2_X1 U10296 ( .A1(n36740), .A2(n36749), .ZN(n36344) );
  NAND2_X2 U10298 ( .A1(n24506), .A2(n34419), .ZN(n37351) );
  NAND3_X1 U10299 ( .A1(n16203), .A2(n11980), .A3(n35321), .ZN(n13952) );
  AOI21_X1 U10303 ( .A1(n22026), .A2(n33764), .B(n13894), .ZN(n13893) );
  NAND2_X1 U10306 ( .A1(n33765), .A2(n13895), .ZN(n13894) );
  NAND2_X1 U10307 ( .A1(n1532), .A2(n18300), .ZN(n3513) );
  NAND2_X1 U10315 ( .A1(n14811), .A2(n64954), .ZN(n34551) );
  NAND3_X1 U10318 ( .A1(n34998), .A2(n34797), .A3(n14112), .ZN(n33765) );
  AND2_X1 U10320 ( .A1(n34250), .A2(n32424), .Z(n32428) );
  NAND3_X1 U10321 ( .A1(n35219), .A2(n24614), .A3(n6842), .ZN(n4162) );
  NAND4_X1 U10324 ( .A1(n34555), .A2(n64708), .A3(n34557), .A4(n64499), .ZN(
        n10944) );
  NOR2_X1 U10325 ( .A1(n34559), .A2(n64708), .ZN(n10138) );
  NAND3_X1 U10326 ( .A1(n57628), .A2(n35304), .A3(n1801), .ZN(n18370) );
  NAND2_X1 U10331 ( .A1(n19435), .A2(n34146), .ZN(n12588) );
  AND2_X1 U10336 ( .A1(n34003), .A2(n34002), .Z(n34660) );
  OR2_X1 U10346 ( .A1(n21096), .A2(n65205), .Z(n6520) );
  INV_X4 U10347 ( .I(n35756), .ZN(n1533) );
  INV_X1 U10349 ( .I(n35305), .ZN(n1801) );
  NAND2_X1 U10359 ( .A1(n2618), .A2(n1430), .ZN(n33777) );
  INV_X1 U10364 ( .I(n58447), .ZN(n1539) );
  NOR2_X1 U10370 ( .A1(n24083), .A2(n1429), .ZN(n34687) );
  NOR4_X1 U10374 ( .A1(n16402), .A2(n35318), .A3(n35755), .A4(n1546), .ZN(
        n5772) );
  INV_X2 U10376 ( .I(n35318), .ZN(n8051) );
  INV_X1 U10387 ( .I(n24829), .ZN(n33233) );
  INV_X1 U10388 ( .I(n9108), .ZN(n8622) );
  INV_X1 U10390 ( .I(n17624), .ZN(n1828) );
  CLKBUF_X2 U10391 ( .I(n10599), .Z(n16706) );
  INV_X2 U10398 ( .I(n26216), .ZN(n1347) );
  INV_X1 U10400 ( .I(n19622), .ZN(n19514) );
  NAND2_X1 U10404 ( .A1(n30838), .A2(n29526), .ZN(n29527) );
  NAND2_X1 U10405 ( .A1(n2794), .A2(n26587), .ZN(n2875) );
  NAND3_X1 U10408 ( .A1(n13175), .A2(n21478), .A3(n30027), .ZN(n5424) );
  AOI21_X1 U10409 ( .A1(n2285), .A2(n2284), .B(n1841), .ZN(n2283) );
  NOR2_X1 U10411 ( .A1(n29911), .A2(n17719), .ZN(n17718) );
  NAND3_X1 U10415 ( .A1(n6796), .A2(n6794), .A3(n6793), .ZN(n17186) );
  NAND3_X1 U10417 ( .A1(n30258), .A2(n2369), .A3(n16630), .ZN(n29925) );
  NOR2_X1 U10418 ( .A1(n20538), .A2(n30630), .ZN(n24328) );
  NAND2_X1 U10421 ( .A1(n21588), .A2(n3849), .ZN(n21677) );
  INV_X1 U10422 ( .I(n30231), .ZN(n1837) );
  NAND2_X1 U10425 ( .A1(n29215), .A2(n30264), .ZN(n6758) );
  AOI21_X1 U10429 ( .A1(n16949), .A2(n6795), .B(n29998), .ZN(n6794) );
  AOI21_X1 U10434 ( .A1(n2519), .A2(n30211), .B(n30222), .ZN(n2443) );
  NOR2_X1 U10445 ( .A1(n2965), .A2(n24206), .ZN(n30768) );
  NAND2_X1 U10448 ( .A1(n30360), .A2(n18322), .ZN(n30449) );
  OAI21_X1 U10449 ( .A1(n30215), .A2(n30212), .B(n16808), .ZN(n2441) );
  AOI21_X1 U10450 ( .A1(n1555), .A2(n3426), .B(n63691), .ZN(n2445) );
  NAND2_X1 U10454 ( .A1(n759), .A2(n19701), .ZN(n30634) );
  INV_X1 U10455 ( .I(n22322), .ZN(n12743) );
  NAND2_X1 U10459 ( .A1(n29736), .A2(n5631), .ZN(n28689) );
  NAND2_X1 U10464 ( .A1(n30242), .A2(n30677), .ZN(n30244) );
  NAND3_X1 U10467 ( .A1(n30195), .A2(n5631), .A3(n30197), .ZN(n11033) );
  NAND2_X1 U10473 ( .A1(n58448), .A2(n60170), .ZN(n3168) );
  INV_X1 U10474 ( .I(n5242), .ZN(n26585) );
  NAND2_X1 U10475 ( .A1(n4270), .A2(n29506), .ZN(n27635) );
  NOR2_X1 U10476 ( .A1(n11425), .A2(n1558), .ZN(n30454) );
  NAND2_X1 U10479 ( .A1(n12632), .A2(n29455), .ZN(n5910) );
  NOR2_X1 U10480 ( .A1(n30786), .A2(n29747), .ZN(n29965) );
  NAND2_X1 U10485 ( .A1(n30677), .A2(n22374), .ZN(n6615) );
  NOR2_X1 U10486 ( .A1(n13943), .A2(n30526), .ZN(n30123) );
  NAND2_X1 U10491 ( .A1(n28546), .A2(n29586), .ZN(n29079) );
  NAND2_X1 U10492 ( .A1(n60162), .A2(n4999), .ZN(n15269) );
  NAND2_X1 U10497 ( .A1(n30319), .A2(n24896), .ZN(n29274) );
  NOR2_X1 U10505 ( .A1(n2140), .A2(n2138), .ZN(n2137) );
  NOR2_X1 U10509 ( .A1(n9833), .A2(n14922), .ZN(n15772) );
  NAND2_X1 U10515 ( .A1(n27377), .A2(n2141), .ZN(n2140) );
  NAND2_X1 U10518 ( .A1(n28103), .A2(n28105), .ZN(n27193) );
  NOR2_X1 U10519 ( .A1(n28421), .A2(n19227), .ZN(n16859) );
  NOR2_X1 U10521 ( .A1(n27379), .A2(n2142), .ZN(n2141) );
  NOR2_X1 U10522 ( .A1(n762), .A2(n27051), .ZN(n26575) );
  NAND2_X1 U10528 ( .A1(n14450), .A2(n12109), .ZN(n28556) );
  AOI21_X1 U10529 ( .A1(n11138), .A2(n11137), .B(n11136), .ZN(n11135) );
  OAI21_X1 U10532 ( .A1(n28397), .A2(n28414), .B(n28417), .ZN(n8338) );
  OAI22_X1 U10533 ( .A1(n29108), .A2(n27998), .B1(n27368), .B2(n27367), .ZN(
        n2136) );
  NOR2_X1 U10534 ( .A1(n27556), .A2(n22902), .ZN(n26629) );
  NAND3_X1 U10541 ( .A1(n62406), .A2(n8478), .A3(n17046), .ZN(n13919) );
  NOR2_X1 U10544 ( .A1(n27851), .A2(n27717), .ZN(n16419) );
  INV_X1 U10546 ( .I(n19643), .ZN(n27345) );
  NAND2_X1 U10551 ( .A1(n28238), .A2(n60505), .ZN(n26525) );
  NAND2_X1 U10553 ( .A1(n7371), .A2(n16654), .ZN(n27301) );
  INV_X1 U10558 ( .I(n6522), .ZN(n29151) );
  NOR2_X1 U10559 ( .A1(n24734), .A2(n24735), .ZN(n26682) );
  NAND2_X1 U10560 ( .A1(n17274), .A2(n29697), .ZN(n28652) );
  NAND2_X1 U10561 ( .A1(n27538), .A2(n27232), .ZN(n27460) );
  NAND2_X1 U10562 ( .A1(n29119), .A2(n8478), .ZN(n15114) );
  NOR2_X1 U10565 ( .A1(n23225), .A2(n26660), .ZN(n13376) );
  AOI22_X1 U10566 ( .A1(n3825), .A2(n6522), .B1(n29152), .B2(n29153), .ZN(
        n3824) );
  INV_X1 U10569 ( .I(n27847), .ZN(n26421) );
  NAND2_X1 U10570 ( .A1(n26527), .A2(n60505), .ZN(n11134) );
  INV_X1 U10571 ( .I(n28250), .ZN(n28071) );
  NOR2_X1 U10573 ( .A1(n22144), .A2(n26969), .ZN(n27214) );
  BUF_X2 U10574 ( .I(n28300), .Z(n22706) );
  NAND3_X1 U10579 ( .A1(n29107), .A2(n60171), .A3(n63850), .ZN(n27375) );
  AOI21_X1 U10581 ( .A1(n28219), .A2(n28226), .B(n27996), .ZN(n27018) );
  BUF_X2 U10585 ( .I(n23328), .Z(n23324) );
  INV_X2 U10587 ( .I(n21720), .ZN(n29156) );
  NAND2_X1 U10588 ( .A1(n28378), .A2(n469), .ZN(n23252) );
  NAND2_X1 U10590 ( .A1(n19972), .A2(n10236), .ZN(n28161) );
  AND2_X1 U10591 ( .A1(n26347), .A2(n25993), .Z(n3317) );
  INV_X1 U10592 ( .I(n7538), .ZN(n5292) );
  NAND2_X1 U10594 ( .A1(n22735), .A2(n23191), .ZN(n26327) );
  NAND2_X1 U10595 ( .A1(n21086), .A2(n10187), .ZN(n11573) );
  INV_X1 U10596 ( .I(n1570), .ZN(n7772) );
  NOR2_X1 U10598 ( .A1(n27810), .A2(n22648), .ZN(n20561) );
  INV_X1 U10599 ( .I(n11850), .ZN(n27618) );
  NAND2_X1 U10600 ( .A1(n14102), .A2(n28223), .ZN(n24190) );
  INV_X1 U10601 ( .I(n27821), .ZN(n29704) );
  INV_X2 U10602 ( .I(n26653), .ZN(n1354) );
  INV_X1 U10606 ( .I(n25222), .ZN(n25221) );
  CLKBUF_X2 U10607 ( .I(n23352), .Z(n10914) );
  BUF_X1 U10610 ( .I(n28187), .Z(n10473) );
  INV_X1 U10611 ( .I(n2276), .ZN(n27369) );
  INV_X2 U10613 ( .I(n13763), .ZN(n1359) );
  NOR2_X1 U10616 ( .A1(n28223), .A2(n23166), .ZN(n27014) );
  NAND2_X1 U10617 ( .A1(n7760), .A2(n27846), .ZN(n27850) );
  CLKBUF_X2 U10618 ( .I(n15790), .Z(n4715) );
  CLKBUF_X2 U10621 ( .I(n26373), .Z(n26742) );
  BUF_X2 U10622 ( .I(n20814), .Z(n51881) );
  INV_X1 U10626 ( .I(n23754), .ZN(n1449) );
  CLKBUF_X2 U10628 ( .I(Key[161]), .Z(n23968) );
  CLKBUF_X2 U10630 ( .I(Key[67]), .Z(n54376) );
  CLKBUF_X2 U10631 ( .I(Key[37]), .Z(n53748) );
  CLKBUF_X2 U10633 ( .I(Key[30]), .Z(n53641) );
  CLKBUF_X2 U10634 ( .I(Key[106]), .Z(n51946) );
  CLKBUF_X2 U10635 ( .I(Key[18]), .Z(n53318) );
  CLKBUF_X2 U10636 ( .I(Key[108]), .Z(n55335) );
  CLKBUF_X2 U10637 ( .I(Key[104]), .Z(n55196) );
  INV_X2 U10638 ( .I(n15789), .ZN(n1364) );
  CLKBUF_X2 U10640 ( .I(Key[105]), .Z(n24046) );
  CLKBUF_X2 U10642 ( .I(Key[80]), .Z(n54716) );
  NAND3_X1 U10646 ( .A1(n6665), .A2(n19020), .A3(n10988), .ZN(n6664) );
  NAND2_X1 U10647 ( .A1(n2837), .A2(n2831), .ZN(n2830) );
  NOR2_X1 U10650 ( .A1(n61253), .A2(n6080), .ZN(n6075) );
  NAND2_X1 U10651 ( .A1(n1577), .A2(n17286), .ZN(n20636) );
  NAND2_X1 U10652 ( .A1(n61727), .A2(n57320), .ZN(n56331) );
  NAND2_X1 U10654 ( .A1(n53814), .A2(n26218), .ZN(n53822) );
  INV_X1 U10655 ( .I(n53365), .ZN(n11962) );
  OAI21_X1 U10657 ( .A1(n53675), .A2(n53700), .B(n53666), .ZN(n2836) );
  INV_X1 U10658 ( .I(n53346), .ZN(n53331) );
  NOR2_X1 U10659 ( .A1(n518), .A2(n1574), .ZN(n11346) );
  NAND2_X1 U10660 ( .A1(n53664), .A2(n53692), .ZN(n2835) );
  AND3_X1 U10661 ( .A1(n518), .A2(n1574), .A3(n53302), .Z(n16057) );
  OAI21_X1 U10663 ( .A1(n20587), .A2(n56502), .B(n15238), .ZN(n15240) );
  AOI21_X1 U10664 ( .A1(n56736), .A2(n56707), .B(n6954), .ZN(n56690) );
  NAND2_X1 U10665 ( .A1(n54194), .A2(n54196), .ZN(n13712) );
  NAND2_X1 U10666 ( .A1(n54928), .A2(n13671), .ZN(n2491) );
  AOI21_X1 U10668 ( .A1(n10736), .A2(n55822), .B(n22860), .ZN(n55824) );
  NAND2_X1 U10671 ( .A1(n54175), .A2(n54207), .ZN(n54176) );
  NAND2_X1 U10673 ( .A1(n6168), .A2(n53998), .ZN(n53960) );
  INV_X4 U10676 ( .I(n17012), .ZN(n1450) );
  INV_X2 U10677 ( .I(n1256), .ZN(n54281) );
  AND2_X1 U10678 ( .A1(n56182), .A2(n56190), .Z(n56192) );
  NOR2_X1 U10680 ( .A1(n54960), .A2(n5051), .ZN(n8410) );
  BUF_X2 U10683 ( .I(n55387), .Z(n9777) );
  BUF_X4 U10685 ( .I(n55818), .Z(n24958) );
  NAND2_X1 U10689 ( .A1(n52048), .A2(n11010), .ZN(n51963) );
  NAND2_X1 U10690 ( .A1(n65283), .A2(n18548), .ZN(n51966) );
  NOR2_X1 U10696 ( .A1(n52943), .A2(n63194), .ZN(n8055) );
  NAND2_X1 U10703 ( .A1(n51258), .A2(n16753), .ZN(n22618) );
  NAND2_X1 U10704 ( .A1(n56259), .A2(n56582), .ZN(n22293) );
  NAND2_X1 U10705 ( .A1(n23845), .A2(n11521), .ZN(n11680) );
  OAI21_X1 U10706 ( .A1(n7332), .A2(n53586), .B(n53590), .ZN(n13473) );
  NAND3_X1 U10708 ( .A1(n56997), .A2(n61572), .A3(n64424), .ZN(n20361) );
  NAND2_X1 U10711 ( .A1(n22804), .A2(n12026), .ZN(n51257) );
  NOR2_X1 U10714 ( .A1(n57040), .A2(n23563), .ZN(n19615) );
  NAND2_X1 U10715 ( .A1(n1453), .A2(n2959), .ZN(n54106) );
  INV_X1 U10716 ( .I(n16748), .ZN(n20613) );
  NAND2_X1 U10717 ( .A1(n20921), .A2(n53241), .ZN(n20342) );
  NAND3_X1 U10718 ( .A1(n1605), .A2(n53580), .A3(n53455), .ZN(n53458) );
  AND2_X1 U10720 ( .A1(n187), .A2(n56563), .Z(n23376) );
  OR2_X1 U10722 ( .A1(n53384), .A2(n52756), .Z(n12290) );
  NAND3_X1 U10723 ( .A1(n4184), .A2(n12818), .A3(n53212), .ZN(n50739) );
  NOR2_X1 U10728 ( .A1(n52222), .A2(n22977), .ZN(n8595) );
  NAND2_X1 U10729 ( .A1(n56267), .A2(n56268), .ZN(n11683) );
  NAND2_X1 U10731 ( .A1(n54980), .A2(n197), .ZN(n52909) );
  AOI21_X1 U10732 ( .A1(n55678), .A2(n4194), .B(n4830), .ZN(n4195) );
  NOR2_X1 U10735 ( .A1(n24870), .A2(n21169), .ZN(n11237) );
  INV_X2 U10737 ( .I(n818), .ZN(n1368) );
  BUF_X2 U10738 ( .I(n61902), .Z(n52892) );
  CLKBUF_X2 U10739 ( .I(n55497), .Z(n10414) );
  OR2_X1 U10741 ( .A1(n54659), .A2(n54657), .Z(n15782) );
  NOR2_X1 U10742 ( .A1(n12573), .A2(n15718), .ZN(n6952) );
  NOR2_X1 U10743 ( .A1(n54321), .A2(n23736), .ZN(n54320) );
  BUF_X1 U10746 ( .I(n54046), .Z(n5025) );
  CLKBUF_X2 U10748 ( .I(n19555), .Z(n22708) );
  BUF_X2 U10749 ( .I(n54112), .Z(n10425) );
  CLKBUF_X2 U10755 ( .I(n53036), .Z(n9613) );
  CLKBUF_X4 U10756 ( .I(n55671), .Z(n20891) );
  CLKBUF_X2 U10760 ( .I(n53226), .Z(n23476) );
  INV_X2 U10762 ( .I(n54659), .ZN(n1371) );
  CLKBUF_X4 U10766 ( .I(n54689), .Z(n15040) );
  INV_X1 U10768 ( .I(n16508), .ZN(n8975) );
  INV_X1 U10769 ( .I(n5603), .ZN(n51391) );
  OAI21_X1 U10776 ( .A1(n47453), .A2(n25193), .B(n52445), .ZN(n9552) );
  NAND2_X1 U10777 ( .A1(n12604), .A2(n48827), .ZN(n12601) );
  INV_X1 U10778 ( .I(n20593), .ZN(n14966) );
  OAI21_X1 U10786 ( .A1(n48417), .A2(n23156), .B(n7652), .ZN(n48827) );
  NAND2_X1 U10792 ( .A1(n8435), .A2(n8433), .ZN(n8432) );
  NAND2_X1 U10794 ( .A1(n50358), .A2(n48265), .ZN(n48267) );
  INV_X1 U10797 ( .I(n50259), .ZN(n1624) );
  NOR3_X1 U10798 ( .A1(n8724), .A2(n4362), .A3(n8725), .ZN(n4614) );
  OAI22_X1 U10799 ( .A1(n50420), .A2(n22805), .B1(n48289), .B2(n48757), .ZN(
        n3678) );
  NOR2_X1 U10800 ( .A1(n49999), .A2(n49998), .ZN(n16676) );
  NOR2_X1 U10802 ( .A1(n49048), .A2(n16024), .ZN(n20642) );
  NAND3_X1 U10803 ( .A1(n48841), .A2(n16829), .A3(n48843), .ZN(n48002) );
  NAND2_X1 U10804 ( .A1(n49275), .A2(n16986), .ZN(n48776) );
  AOI21_X1 U10820 ( .A1(n48690), .A2(n1474), .B(n17683), .ZN(n6277) );
  AOI21_X1 U10821 ( .A1(n3885), .A2(n14007), .B(n48325), .ZN(n2758) );
  NOR3_X1 U10822 ( .A1(n1261), .A2(n13038), .A3(n62606), .ZN(n14209) );
  NAND2_X1 U10823 ( .A1(n49804), .A2(n858), .ZN(n11219) );
  OAI21_X1 U10824 ( .A1(n49788), .A2(n20708), .B(n7146), .ZN(n49805) );
  NOR2_X1 U10826 ( .A1(n49612), .A2(n49320), .ZN(n7005) );
  INV_X1 U10827 ( .I(n49463), .ZN(n5568) );
  NOR2_X1 U10828 ( .A1(n44667), .A2(n48340), .ZN(n44668) );
  INV_X1 U10833 ( .I(n48419), .ZN(n47966) );
  AND2_X1 U10834 ( .A1(n18007), .A2(n20971), .Z(n10346) );
  NAND2_X1 U10839 ( .A1(n50216), .A2(n7824), .ZN(n25081) );
  INV_X1 U10840 ( .I(n49919), .ZN(n1629) );
  NAND2_X1 U10841 ( .A1(n47796), .A2(n49642), .ZN(n14310) );
  OAI21_X1 U10843 ( .A1(n18844), .A2(n49918), .B(n3065), .ZN(n2983) );
  NOR2_X1 U10846 ( .A1(n49526), .A2(n406), .ZN(n16484) );
  NAND2_X1 U10847 ( .A1(n23141), .A2(n49767), .ZN(n48948) );
  NOR2_X1 U10849 ( .A1(n58645), .A2(n49677), .ZN(n2582) );
  NOR2_X1 U10852 ( .A1(n62744), .A2(n48845), .ZN(n18433) );
  OAI21_X1 U10855 ( .A1(n1471), .A2(n18609), .B(n21092), .ZN(n14831) );
  AND2_X2 U10865 ( .A1(n24332), .A2(n48868), .Z(n7078) );
  NAND2_X1 U10872 ( .A1(n19634), .A2(n60622), .ZN(n8895) );
  INV_X4 U10875 ( .I(n49940), .ZN(n1379) );
  NOR2_X1 U10880 ( .A1(n46074), .A2(n6656), .ZN(n6655) );
  OAI21_X1 U10890 ( .A1(n8573), .A2(n47811), .B(n8571), .ZN(n25899) );
  OAI21_X1 U10892 ( .A1(n45806), .A2(n23850), .B(n23099), .ZN(n13722) );
  NAND2_X1 U10898 ( .A1(n1103), .A2(n47809), .ZN(n5311) );
  OAI21_X1 U10900 ( .A1(n8572), .A2(n45203), .B(n47811), .ZN(n8571) );
  OAI21_X1 U10905 ( .A1(n47536), .A2(n5771), .B(n8820), .ZN(n47537) );
  AND2_X1 U10908 ( .A1(n22093), .A2(n62247), .Z(n16053) );
  INV_X1 U10909 ( .I(n3358), .ZN(n3357) );
  NOR2_X1 U10915 ( .A1(n9794), .A2(n9793), .ZN(n47129) );
  NAND2_X1 U10918 ( .A1(n48152), .A2(n46752), .ZN(n25414) );
  OAI21_X1 U10927 ( .A1(n47691), .A2(n1263), .B(n13497), .ZN(n13496) );
  OAI21_X1 U10929 ( .A1(n59269), .A2(n47128), .B(n1650), .ZN(n9793) );
  NAND2_X1 U10934 ( .A1(n23903), .A2(n45785), .ZN(n44702) );
  NAND2_X1 U10935 ( .A1(n4655), .A2(n178), .ZN(n46482) );
  NAND2_X1 U10936 ( .A1(n60839), .A2(n47000), .ZN(n47484) );
  NAND2_X1 U10937 ( .A1(n8649), .A2(n58155), .ZN(n8645) );
  NAND2_X1 U10938 ( .A1(n48640), .A2(n21855), .ZN(n7051) );
  NAND2_X1 U10940 ( .A1(n47772), .A2(n13566), .ZN(n44554) );
  NAND2_X1 U10944 ( .A1(n47123), .A2(n47119), .ZN(n46762) );
  INV_X1 U10945 ( .I(n8758), .ZN(n13587) );
  AND2_X1 U10947 ( .A1(n47721), .A2(n47720), .Z(n47722) );
  NOR2_X1 U10949 ( .A1(n47250), .A2(n46893), .ZN(n12723) );
  NAND2_X1 U10956 ( .A1(n25026), .A2(n47874), .ZN(n47360) );
  AND2_X1 U10958 ( .A1(n47905), .A2(n23969), .Z(n16143) );
  NOR2_X1 U10961 ( .A1(n47717), .A2(n47883), .ZN(n11896) );
  NAND3_X1 U10962 ( .A1(n47882), .A2(n12647), .A3(n47880), .ZN(n9454) );
  NOR2_X1 U10966 ( .A1(n2955), .A2(n23850), .ZN(n14786) );
  NOR2_X1 U10968 ( .A1(n2223), .A2(n47592), .ZN(n47279) );
  NAND2_X1 U10979 ( .A1(n13356), .A2(n47576), .ZN(n45193) );
  AND2_X1 U10981 ( .A1(n47470), .A2(n1660), .Z(n2826) );
  INV_X1 U10982 ( .I(n7579), .ZN(n14121) );
  NOR2_X1 U10983 ( .A1(n25006), .A2(n11627), .ZN(n47870) );
  CLKBUF_X2 U10984 ( .I(n3733), .Z(n3732) );
  NOR2_X1 U10986 ( .A1(n1267), .A2(n46906), .ZN(n44196) );
  INV_X1 U10988 ( .I(n47880), .ZN(n14474) );
  INV_X1 U10989 ( .I(n14289), .ZN(n11901) );
  INV_X1 U10991 ( .I(n46905), .ZN(n6892) );
  OR2_X1 U10992 ( .A1(n59695), .A2(n23405), .Z(n8224) );
  NAND2_X1 U10994 ( .A1(n6645), .A2(n1482), .ZN(n46942) );
  INV_X1 U10995 ( .I(n47860), .ZN(n25006) );
  INV_X1 U11004 ( .I(n10055), .ZN(n1660) );
  BUF_X2 U11009 ( .I(n47252), .Z(n9730) );
  NOR2_X1 U11010 ( .A1(n48654), .A2(n3365), .ZN(n17318) );
  INV_X4 U11018 ( .I(n6082), .ZN(n1388) );
  BUF_X2 U11021 ( .I(n44181), .Z(n46913) );
  INV_X1 U11022 ( .I(n15266), .ZN(n46407) );
  NOR2_X1 U11023 ( .A1(n10077), .A2(n23006), .ZN(n25494) );
  INV_X1 U11025 ( .I(n19411), .ZN(n14806) );
  INV_X1 U11026 ( .I(n10099), .ZN(n25693) );
  CLKBUF_X2 U11029 ( .I(n44819), .Z(n10099) );
  INV_X2 U11031 ( .I(n26167), .ZN(n8620) );
  INV_X1 U11037 ( .I(n1682), .ZN(n10745) );
  CLKBUF_X2 U11040 ( .I(n16909), .Z(n20772) );
  INV_X1 U11041 ( .I(n24030), .ZN(n7552) );
  INV_X1 U11043 ( .I(n44091), .ZN(n1682) );
  AOI21_X1 U11047 ( .A1(n42623), .A2(n22088), .B(n43681), .ZN(n44091) );
  INV_X1 U11051 ( .I(n44329), .ZN(n46236) );
  AOI22_X1 U11063 ( .A1(n43207), .A2(n22109), .B1(n43060), .B2(n43203), .ZN(
        n43063) );
  AND4_X1 U11065 ( .A1(n43292), .A2(n16659), .A3(n20639), .A4(n11366), .Z(
        n43110) );
  NAND2_X1 U11066 ( .A1(n11405), .A2(n11404), .ZN(n21758) );
  OAI21_X1 U11069 ( .A1(n42543), .A2(n41576), .B(n13099), .ZN(n5930) );
  NOR2_X1 U11072 ( .A1(n42847), .A2(n43742), .ZN(n15657) );
  NAND4_X1 U11074 ( .A1(n15334), .A2(n18154), .A3(n18725), .A4(n7144), .ZN(
        n18153) );
  NAND3_X1 U11075 ( .A1(n43581), .A2(n43583), .A3(n43582), .ZN(n2689) );
  NAND2_X1 U11080 ( .A1(n6563), .A2(n43104), .ZN(n43292) );
  NAND2_X1 U11083 ( .A1(n16940), .A2(n43298), .ZN(n16550) );
  INV_X1 U11087 ( .I(n42011), .ZN(n6111) );
  AND2_X1 U11089 ( .A1(n42927), .A2(n12961), .Z(n15493) );
  AND3_X1 U11091 ( .A1(n43052), .A2(n60843), .A3(n43868), .Z(n43054) );
  NOR2_X1 U11092 ( .A1(n41777), .A2(n42887), .ZN(n24100) );
  OR2_X1 U11094 ( .A1(n57410), .A2(n42973), .Z(n42974) );
  OAI22_X1 U11098 ( .A1(n41696), .A2(n23838), .B1(n59067), .B2(n43359), .ZN(
        n12195) );
  OR2_X1 U11106 ( .A1(n42369), .A2(n43439), .Z(n24996) );
  AOI21_X1 U11107 ( .A1(n3956), .A2(n7720), .B(n61198), .ZN(n3955) );
  INV_X1 U11111 ( .I(n43915), .ZN(n1933) );
  OAI22_X1 U11113 ( .A1(n43346), .A2(n60843), .B1(n43351), .B2(n41594), .ZN(
        n41595) );
  NAND3_X1 U11117 ( .A1(n1333), .A2(n43897), .A3(n3696), .ZN(n43662) );
  NAND2_X1 U11120 ( .A1(n43868), .A2(n7950), .ZN(n6734) );
  INV_X1 U11122 ( .I(n21950), .ZN(n11361) );
  AOI21_X1 U11124 ( .A1(n42737), .A2(n42736), .B(n43364), .ZN(n42738) );
  AND2_X1 U11131 ( .A1(n6563), .A2(n20844), .Z(n8468) );
  INV_X1 U11134 ( .I(n42543), .ZN(n42930) );
  NAND2_X1 U11136 ( .A1(n43156), .A2(n11179), .ZN(n42565) );
  NOR3_X1 U11137 ( .A1(n41714), .A2(n10617), .A3(n41715), .ZN(n16139) );
  INV_X1 U11140 ( .I(n43577), .ZN(n43575) );
  NAND2_X1 U11144 ( .A1(n42395), .A2(n42394), .ZN(n18343) );
  NOR3_X2 U11153 ( .A1(n24715), .A2(n43380), .A3(n41698), .ZN(n42629) );
  NAND3_X1 U11157 ( .A1(n43695), .A2(n16527), .A3(n43698), .ZN(n16998) );
  NOR2_X1 U11158 ( .A1(n43582), .A2(n6865), .ZN(n43574) );
  NAND2_X1 U11159 ( .A1(n1697), .A2(n1500), .ZN(n40283) );
  NAND2_X1 U11163 ( .A1(n12064), .A2(n64156), .ZN(n15637) );
  AOI21_X1 U11164 ( .A1(n42849), .A2(n41561), .B(n41562), .ZN(n3633) );
  NOR2_X1 U11165 ( .A1(n14051), .A2(n3674), .ZN(n13075) );
  NOR2_X1 U11166 ( .A1(n5787), .A2(n8139), .ZN(n38349) );
  AOI21_X1 U11170 ( .A1(n10827), .A2(n1502), .B(n42865), .ZN(n41507) );
  NAND2_X1 U11172 ( .A1(n24179), .A2(n20844), .ZN(n43105) );
  AND2_X1 U11173 ( .A1(n42669), .A2(n10865), .Z(n11881) );
  INV_X1 U11182 ( .I(n42129), .ZN(n42661) );
  NOR2_X1 U11183 ( .A1(n43270), .A2(n2330), .ZN(n13596) );
  INV_X1 U11186 ( .I(n42717), .ZN(n1696) );
  INV_X4 U11188 ( .I(n42080), .ZN(n1392) );
  INV_X1 U11191 ( .I(n6297), .ZN(n15792) );
  NAND2_X1 U11193 ( .A1(n42354), .A2(n20922), .ZN(n41611) );
  INV_X2 U11194 ( .I(n42377), .ZN(n1394) );
  INV_X1 U11197 ( .I(n43717), .ZN(n8690) );
  INV_X1 U11199 ( .I(n19358), .ZN(n1702) );
  INV_X4 U11206 ( .I(n1701), .ZN(n1398) );
  AOI21_X1 U11208 ( .A1(n41250), .A2(n14816), .B(n14813), .ZN(n41252) );
  NAND3_X1 U11215 ( .A1(n7845), .A2(n11631), .A3(n18594), .ZN(n2877) );
  NAND2_X1 U11222 ( .A1(n14814), .A2(n999), .ZN(n14813) );
  INV_X1 U11223 ( .I(n40862), .ZN(n18028) );
  OAI21_X1 U11229 ( .A1(n61708), .A2(n1515), .B(n40350), .ZN(n11101) );
  NOR3_X1 U11232 ( .A1(n5788), .A2(n41800), .A3(n61435), .ZN(n5792) );
  OR3_X1 U11233 ( .A1(n40066), .A2(n64242), .A3(n60113), .Z(n36652) );
  NAND2_X1 U11241 ( .A1(n41447), .A2(n357), .ZN(n41448) );
  OAI22_X1 U11244 ( .A1(n42260), .A2(n40577), .B1(n42262), .B2(n41906), .ZN(
        n15397) );
  NOR2_X1 U11247 ( .A1(n41155), .A2(n1516), .ZN(n13737) );
  INV_X1 U11248 ( .I(n42303), .ZN(n42306) );
  AND4_X1 U11252 ( .A1(n39161), .A2(n39160), .A3(n65206), .A4(n39159), .Z(
        n39162) );
  NAND2_X1 U11253 ( .A1(n20984), .A2(n41155), .ZN(n5675) );
  NOR2_X1 U11254 ( .A1(n41065), .A2(n41876), .ZN(n3048) );
  NAND3_X1 U11261 ( .A1(n13310), .A2(n38496), .A3(n41031), .ZN(n13309) );
  NAND3_X1 U11263 ( .A1(n13307), .A2(n13308), .A3(n38498), .ZN(n8485) );
  INV_X1 U11269 ( .I(n42523), .ZN(n1506) );
  AND3_X1 U11272 ( .A1(n22713), .A2(n8017), .A3(n10481), .Z(n14820) );
  NOR2_X1 U11273 ( .A1(n40507), .A2(n19458), .ZN(n41013) );
  INV_X1 U11274 ( .I(n60652), .ZN(n41002) );
  NOR3_X1 U11275 ( .A1(n60166), .A2(n39118), .A3(n24743), .ZN(n7646) );
  NAND2_X1 U11276 ( .A1(n40217), .A2(n12409), .ZN(n37062) );
  NOR2_X1 U11277 ( .A1(n61986), .A2(n6625), .ZN(n36996) );
  NAND2_X1 U11278 ( .A1(n39118), .A2(n7649), .ZN(n7648) );
  NOR2_X1 U11279 ( .A1(n39418), .A2(n1518), .ZN(n11132) );
  NAND3_X1 U11280 ( .A1(n40123), .A2(n39408), .A3(n42495), .ZN(n39409) );
  NAND2_X1 U11284 ( .A1(n10954), .A2(n3356), .ZN(n6767) );
  NOR2_X1 U11289 ( .A1(n11787), .A2(n41186), .ZN(n7327) );
  NAND2_X1 U11291 ( .A1(n39869), .A2(n38938), .ZN(n12943) );
  NAND2_X1 U11292 ( .A1(n25976), .A2(n15440), .ZN(n15439) );
  INV_X1 U11293 ( .I(n40379), .ZN(n41427) );
  AOI22_X1 U11294 ( .A1(n60166), .A2(n40607), .B1(n41017), .B2(n1512), .ZN(
        n38426) );
  OR2_X1 U11295 ( .A1(n40217), .A2(n62681), .Z(n5394) );
  NAND3_X1 U11297 ( .A1(n40273), .A2(n40328), .A3(n25229), .ZN(n21924) );
  OAI21_X1 U11299 ( .A1(n40541), .A2(n10587), .B(n40648), .ZN(n38406) );
  AOI21_X1 U11300 ( .A1(n61746), .A2(n41806), .B(n42452), .ZN(n6199) );
  INV_X1 U11301 ( .I(n41280), .ZN(n41269) );
  NAND2_X1 U11304 ( .A1(n39104), .A2(n23986), .ZN(n40202) );
  NAND2_X1 U11307 ( .A1(n62291), .A2(n40064), .ZN(n41813) );
  INV_X1 U11308 ( .I(n42465), .ZN(n21865) );
  NAND4_X1 U11309 ( .A1(n40196), .A2(n40200), .A3(n22593), .A4(n40199), .ZN(
        n37416) );
  INV_X1 U11312 ( .I(n11765), .ZN(n25606) );
  NOR2_X1 U11314 ( .A1(n57208), .A2(n40314), .ZN(n15542) );
  INV_X1 U11315 ( .I(n17930), .ZN(n42436) );
  INV_X1 U11318 ( .I(n10883), .ZN(n41478) );
  INV_X1 U11327 ( .I(n21506), .ZN(n39982) );
  CLKBUF_X2 U11331 ( .I(n40934), .Z(n7201) );
  INV_X1 U11334 ( .I(n13985), .ZN(n40316) );
  NAND2_X1 U11335 ( .A1(n8026), .A2(n709), .ZN(n5709) );
  INV_X1 U11338 ( .I(n40956), .ZN(n1740) );
  OR2_X2 U11341 ( .A1(n19010), .A2(n61653), .Z(n16601) );
  CLKBUF_X2 U11347 ( .I(n17382), .Z(n20984) );
  BUF_X2 U11350 ( .I(n26182), .Z(n10294) );
  BUF_X2 U11352 ( .I(n15590), .Z(n11472) );
  INV_X2 U11354 ( .I(n25141), .ZN(n1408) );
  INV_X2 U11357 ( .I(n5271), .ZN(n1409) );
  INV_X2 U11359 ( .I(n22307), .ZN(n1410) );
  INV_X1 U11360 ( .I(n920), .ZN(n10145) );
  INV_X2 U11361 ( .I(n7619), .ZN(n2741) );
  INV_X1 U11363 ( .I(n38386), .ZN(n14751) );
  BUF_X2 U11365 ( .I(n38004), .Z(n23695) );
  INV_X2 U11374 ( .I(n4919), .ZN(n1411) );
  INV_X2 U11375 ( .I(n14755), .ZN(n1412) );
  INV_X1 U11384 ( .I(n37851), .ZN(n6490) );
  BUF_X2 U11385 ( .I(n22949), .Z(n37525) );
  NAND2_X1 U11387 ( .A1(n36694), .A2(n36693), .ZN(n21941) );
  AND2_X1 U11389 ( .A1(n34291), .A2(n37432), .Z(n25212) );
  NOR2_X1 U11390 ( .A1(n933), .A2(n36720), .ZN(n34807) );
  INV_X1 U11391 ( .I(n36694), .ZN(n6132) );
  NOR2_X1 U11394 ( .A1(n933), .A2(n21544), .ZN(n21543) );
  NAND2_X1 U11395 ( .A1(n36409), .A2(n36402), .ZN(n8765) );
  AOI21_X1 U11396 ( .A1(n14264), .A2(n36109), .B(n22474), .ZN(n35115) );
  OAI21_X1 U11399 ( .A1(n36617), .A2(n36618), .B(n7759), .ZN(n36619) );
  INV_X1 U11406 ( .I(n37331), .ZN(n34882) );
  NOR2_X1 U11416 ( .A1(n36447), .A2(n20728), .ZN(n21457) );
  NAND2_X1 U11417 ( .A1(n18352), .A2(n64093), .ZN(n36503) );
  NOR2_X1 U11426 ( .A1(n36773), .A2(n14951), .ZN(n19188) );
  OAI21_X1 U11428 ( .A1(n9933), .A2(n9932), .B(n15754), .ZN(n16635) );
  NOR2_X1 U11429 ( .A1(n37405), .A2(n6540), .ZN(n8976) );
  NOR2_X1 U11433 ( .A1(n36776), .A2(n10718), .ZN(n2807) );
  NOR2_X1 U11437 ( .A1(n37248), .A2(n12458), .ZN(n12457) );
  NAND2_X1 U11439 ( .A1(n2592), .A2(n9783), .ZN(n2591) );
  OR2_X1 U11441 ( .A1(n24660), .A2(n24659), .Z(n37189) );
  NAND3_X1 U11443 ( .A1(n1903), .A2(n1311), .A3(n948), .ZN(n35179) );
  INV_X4 U11444 ( .I(n23226), .ZN(n1524) );
  NAND3_X1 U11446 ( .A1(n35918), .A2(n36325), .A3(n37400), .ZN(n35924) );
  NAND2_X1 U11450 ( .A1(n36576), .A2(n36570), .ZN(n20167) );
  OAI22_X1 U11453 ( .A1(n12031), .A2(n3622), .B1(n36763), .B2(n34004), .ZN(
        n34005) );
  AOI21_X1 U11454 ( .A1(n36301), .A2(n36300), .B(n36808), .ZN(n34579) );
  INV_X2 U11455 ( .I(n12301), .ZN(n4834) );
  AOI21_X1 U11465 ( .A1(n33787), .A2(n36170), .B(n22155), .ZN(n33788) );
  OR3_X1 U11468 ( .A1(n36622), .A2(n36621), .A3(n1527), .Z(n11601) );
  OAI21_X1 U11472 ( .A1(n34923), .A2(n34924), .B(n18509), .ZN(n11832) );
  NAND3_X1 U11473 ( .A1(n36152), .A2(n33526), .A3(n1767), .ZN(n2299) );
  NAND2_X1 U11474 ( .A1(n10165), .A2(n36777), .ZN(n10718) );
  INV_X1 U11475 ( .I(n37314), .ZN(n35083) );
  NAND3_X1 U11476 ( .A1(n37446), .A2(n36969), .A3(n37455), .ZN(n35854) );
  BUF_X4 U11478 ( .I(n32076), .Z(n37333) );
  NAND2_X1 U11481 ( .A1(n35416), .A2(n14952), .ZN(n14951) );
  NOR3_X1 U11482 ( .A1(n36627), .A2(n35447), .A3(n1527), .ZN(n7723) );
  NAND2_X1 U11484 ( .A1(n6606), .A2(n35964), .ZN(n15070) );
  BUF_X4 U11492 ( .I(n37288), .Z(n23226) );
  NAND3_X1 U11495 ( .A1(n10485), .A2(n36742), .A3(n36748), .ZN(n2020) );
  NOR2_X1 U11498 ( .A1(n36740), .A2(n12863), .ZN(n35062) );
  NAND2_X1 U11499 ( .A1(n36170), .A2(n25163), .ZN(n3459) );
  NOR2_X1 U11501 ( .A1(n36605), .A2(n62672), .ZN(n37047) );
  NAND2_X1 U11503 ( .A1(n12652), .A2(n1338), .ZN(n36622) );
  NOR2_X1 U11505 ( .A1(n34855), .A2(n12141), .ZN(n36048) );
  NOR2_X1 U11506 ( .A1(n35903), .A2(n21010), .ZN(n19509) );
  NAND2_X1 U11516 ( .A1(n11272), .A2(n36459), .ZN(n12351) );
  NOR2_X1 U11517 ( .A1(n36774), .A2(n2002), .ZN(n10061) );
  OR2_X1 U11518 ( .A1(n12883), .A2(n9013), .Z(n12882) );
  NOR2_X1 U11520 ( .A1(n36921), .A2(n4304), .ZN(n19764) );
  OAI21_X1 U11525 ( .A1(n36841), .A2(n26213), .B(n61747), .ZN(n4852) );
  INV_X1 U11530 ( .I(n2158), .ZN(n6491) );
  NAND3_X1 U11531 ( .A1(n1415), .A2(n22431), .A3(n3856), .ZN(n11028) );
  NOR2_X1 U11532 ( .A1(n1777), .A2(n34927), .ZN(n35509) );
  NAND2_X1 U11539 ( .A1(n36742), .A2(n20812), .ZN(n35860) );
  NAND3_X1 U11541 ( .A1(n36422), .A2(n36170), .A3(n1227), .ZN(n36177) );
  CLKBUF_X2 U11543 ( .I(n15743), .Z(n10226) );
  NAND2_X1 U11545 ( .A1(n36574), .A2(n64181), .ZN(n36557) );
  OAI21_X1 U11548 ( .A1(n1339), .A2(n36553), .B(n19364), .ZN(n36096) );
  INV_X1 U11549 ( .I(n13210), .ZN(n36459) );
  NOR2_X1 U11553 ( .A1(n35427), .A2(n36944), .ZN(n36952) );
  INV_X4 U11554 ( .I(n2900), .ZN(n1416) );
  INV_X4 U11558 ( .I(n26243), .ZN(n1418) );
  AOI21_X1 U11570 ( .A1(n12982), .A2(n3513), .B(n34065), .ZN(n3512) );
  INV_X4 U11571 ( .I(n24864), .ZN(n1422) );
  OR2_X2 U11574 ( .A1(n15287), .A2(n15284), .Z(n35178) );
  NAND2_X1 U11578 ( .A1(n13770), .A2(n5772), .ZN(n35315) );
  OAI21_X1 U11579 ( .A1(n34652), .A2(n32883), .B(n24664), .ZN(n3132) );
  NAND3_X1 U11585 ( .A1(n20313), .A2(n20314), .A3(n19805), .ZN(n20312) );
  INV_X1 U11590 ( .I(n35782), .ZN(n19997) );
  OAI22_X1 U11591 ( .A1(n17048), .A2(n32890), .B1(n1539), .B2(n2393), .ZN(
        n2392) );
  AND2_X1 U11592 ( .A1(n7345), .A2(n1546), .Z(n10809) );
  NAND2_X1 U11597 ( .A1(n32831), .A2(n18390), .ZN(n2393) );
  AND3_X1 U11605 ( .A1(n20569), .A2(n22598), .A3(n7183), .Z(n32824) );
  NOR3_X1 U11606 ( .A1(n14953), .A2(n34172), .A3(n34660), .ZN(n16989) );
  OAI21_X1 U11607 ( .A1(n1796), .A2(n63085), .B(n33616), .ZN(n20325) );
  OR2_X1 U11610 ( .A1(n35686), .A2(n23313), .Z(n3981) );
  AOI22_X1 U11616 ( .A1(n34041), .A2(n34040), .B1(n34607), .B2(n34039), .ZN(
        n34049) );
  OAI21_X1 U11618 ( .A1(n35819), .A2(n35820), .B(n35818), .ZN(n3487) );
  NOR2_X1 U11619 ( .A1(n33477), .A2(n64958), .ZN(n2306) );
  NAND2_X1 U11621 ( .A1(n33520), .A2(n35021), .ZN(n14045) );
  INV_X1 U11623 ( .I(n34251), .ZN(n34360) );
  INV_X1 U11624 ( .I(n33690), .ZN(n33559) );
  NAND2_X1 U11625 ( .A1(n33975), .A2(n34040), .ZN(n31024) );
  NAND2_X1 U11626 ( .A1(n33621), .A2(n33620), .ZN(n4879) );
  NOR2_X1 U11627 ( .A1(n22428), .A2(n9329), .ZN(n33549) );
  AND2_X1 U11630 ( .A1(n11709), .A2(n7155), .Z(n32296) );
  OR2_X1 U11638 ( .A1(n33419), .A2(n14320), .Z(n14319) );
  NOR2_X1 U11639 ( .A1(n1798), .A2(n33984), .ZN(n4627) );
  NOR2_X1 U11644 ( .A1(n57166), .A2(n34953), .ZN(n12406) );
  AND2_X1 U11647 ( .A1(n34982), .A2(n2322), .Z(n34983) );
  NAND2_X1 U11648 ( .A1(n34002), .A2(n60628), .ZN(n31469) );
  INV_X1 U11649 ( .I(n34550), .ZN(n16580) );
  NAND2_X1 U11652 ( .A1(n10769), .A2(n11659), .ZN(n32132) );
  AOI21_X1 U11654 ( .A1(n22342), .A2(n33478), .B(n5529), .ZN(n33480) );
  INV_X1 U11655 ( .I(n35235), .ZN(n33216) );
  NAND2_X1 U11656 ( .A1(n22909), .A2(n62683), .ZN(n8879) );
  AND2_X1 U11657 ( .A1(n5386), .A2(n32892), .Z(n21431) );
  NOR2_X1 U11659 ( .A1(n32990), .A2(n33548), .ZN(n33543) );
  NAND2_X1 U11661 ( .A1(n1538), .A2(n2208), .ZN(n2210) );
  INV_X1 U11662 ( .I(n13141), .ZN(n17041) );
  INV_X2 U11663 ( .I(n34603), .ZN(n1798) );
  NAND2_X1 U11664 ( .A1(n3489), .A2(n3488), .ZN(n35818) );
  OAI22_X1 U11665 ( .A1(n1537), .A2(n18077), .B1(n34956), .B2(n57166), .ZN(
        n7727) );
  NAND2_X1 U11668 ( .A1(n32870), .A2(n33950), .ZN(n21217) );
  NOR2_X1 U11672 ( .A1(n35799), .A2(n35806), .ZN(n24956) );
  NAND2_X1 U11673 ( .A1(n1813), .A2(n34056), .ZN(n34051) );
  NAND2_X1 U11677 ( .A1(n35821), .A2(n35817), .ZN(n34239) );
  NAND2_X1 U11686 ( .A1(n9030), .A2(n60835), .ZN(n33584) );
  INV_X1 U11691 ( .I(n904), .ZN(n35702) );
  AND2_X1 U11694 ( .A1(n34989), .A2(n34069), .Z(n2273) );
  NAND2_X1 U11695 ( .A1(n34670), .A2(n64358), .ZN(n3745) );
  INV_X4 U11699 ( .I(n34993), .ZN(n1424) );
  INV_X1 U11700 ( .I(n35620), .ZN(n35206) );
  NOR2_X1 U11706 ( .A1(n15756), .A2(n35031), .ZN(n23014) );
  INV_X4 U11710 ( .I(n24935), .ZN(n35816) );
  INV_X1 U11712 ( .I(n15807), .ZN(n35203) );
  INV_X1 U11714 ( .I(n34521), .ZN(n15786) );
  CLKBUF_X2 U11716 ( .I(n22236), .Z(n10337) );
  INV_X2 U11721 ( .I(n25465), .ZN(n1429) );
  INV_X1 U11727 ( .I(n11506), .ZN(n9528) );
  INV_X2 U11729 ( .I(n17299), .ZN(n1550) );
  NAND2_X2 U11736 ( .A1(n8586), .A2(n1836), .ZN(n13963) );
  NOR2_X1 U11737 ( .A1(n13842), .A2(n12897), .ZN(n8461) );
  NOR2_X1 U11751 ( .A1(n2224), .A2(n2445), .ZN(n2444) );
  OAI21_X1 U11755 ( .A1(n24158), .A2(n24159), .B(n24157), .ZN(n31873) );
  NAND2_X2 U11757 ( .A1(n13215), .A2(n13216), .ZN(n32283) );
  AOI22_X1 U11760 ( .A1(n30220), .A2(n7040), .B1(n30219), .B2(n1555), .ZN(
        n30221) );
  NOR2_X1 U11761 ( .A1(n29489), .A2(n15774), .ZN(n17789) );
  OAI22_X1 U11765 ( .A1(n31223), .A2(n7426), .B1(n10923), .B2(n30665), .ZN(
        n10922) );
  OAI22_X1 U11766 ( .A1(n29421), .A2(n15433), .B1(n28289), .B2(n30363), .ZN(
        n11566) );
  NAND2_X1 U11774 ( .A1(n1837), .A2(n1862), .ZN(n14336) );
  INV_X1 U11775 ( .I(n28102), .ZN(n14668) );
  NAND3_X1 U11777 ( .A1(n29400), .A2(n29886), .A3(n29396), .ZN(n1988) );
  NOR2_X1 U11781 ( .A1(n2439), .A2(n2437), .ZN(n2436) );
  NOR2_X1 U11783 ( .A1(n29426), .A2(n20859), .ZN(n28705) );
  NAND2_X1 U11788 ( .A1(n2441), .A2(n2440), .ZN(n2439) );
  INV_X1 U11789 ( .I(n31191), .ZN(n30867) );
  NAND3_X1 U11791 ( .A1(n29574), .A2(n30301), .A3(n29573), .ZN(n15686) );
  NAND2_X1 U11792 ( .A1(n3797), .A2(n29779), .ZN(n27792) );
  OAI22_X1 U11793 ( .A1(n16060), .A2(n30173), .B1(n31054), .B2(n23144), .ZN(
        n27365) );
  OAI21_X1 U11795 ( .A1(n19754), .A2(n4414), .B(n327), .ZN(n4725) );
  NOR2_X1 U11797 ( .A1(n30574), .A2(n15774), .ZN(n17785) );
  NAND4_X1 U11799 ( .A1(n19885), .A2(n26238), .A3(n28980), .A4(n28979), .ZN(
        n19297) );
  OAI21_X1 U11802 ( .A1(n30096), .A2(n22799), .B(n11033), .ZN(n11032) );
  NAND3_X1 U11804 ( .A1(n4764), .A2(n30634), .A3(n30633), .ZN(n5742) );
  NOR2_X1 U11805 ( .A1(n30678), .A2(n30685), .ZN(n4736) );
  NAND2_X1 U11806 ( .A1(n30731), .A2(n30285), .ZN(n7548) );
  INV_X1 U11808 ( .I(n14701), .ZN(n14851) );
  OAI21_X1 U11812 ( .A1(n1553), .A2(n29274), .B(n61052), .ZN(n4101) );
  AOI21_X1 U11814 ( .A1(n30538), .A2(n1277), .B(n24299), .ZN(n29977) );
  AND3_X1 U11819 ( .A1(n60170), .A2(n4999), .A3(n875), .Z(n13182) );
  NAND2_X1 U11824 ( .A1(n1351), .A2(n30123), .ZN(n30120) );
  INV_X1 U11825 ( .I(n30676), .ZN(n30238) );
  NAND2_X1 U11826 ( .A1(n3426), .A2(n9000), .ZN(n8999) );
  NAND3_X1 U11831 ( .A1(n9979), .A2(n20391), .A3(n30740), .ZN(n30741) );
  NAND3_X1 U11833 ( .A1(n28681), .A2(n24564), .A3(n30747), .ZN(n11967) );
  INV_X1 U11836 ( .I(n29248), .ZN(n3797) );
  AOI21_X1 U11838 ( .A1(n28689), .A2(n26308), .B(n57436), .ZN(n11175) );
  NAND2_X1 U11845 ( .A1(n23349), .A2(n30680), .ZN(n15135) );
  NAND2_X1 U11847 ( .A1(n20069), .A2(n31280), .ZN(n4414) );
  NAND2_X1 U11848 ( .A1(n1554), .A2(n30085), .ZN(n2733) );
  NAND2_X1 U11850 ( .A1(n29904), .A2(n18005), .ZN(n30865) );
  NOR2_X1 U11851 ( .A1(n29267), .A2(n1562), .ZN(n29262) );
  NAND2_X1 U11854 ( .A1(n17745), .A2(n29959), .ZN(n29960) );
  NOR3_X1 U11857 ( .A1(n30680), .A2(n19461), .A3(n18198), .ZN(n13844) );
  OAI21_X1 U11859 ( .A1(n60162), .A2(n30455), .B(n20859), .ZN(n28706) );
  NOR2_X1 U11863 ( .A1(n1278), .A2(n25052), .ZN(n10925) );
  NAND2_X1 U11865 ( .A1(n30480), .A2(n9392), .ZN(n30488) );
  NOR2_X1 U11868 ( .A1(n1352), .A2(n60284), .ZN(n4787) );
  NOR3_X1 U11869 ( .A1(n22504), .A2(n8168), .A3(n8166), .ZN(n30350) );
  INV_X1 U11870 ( .I(n30002), .ZN(n30745) );
  AOI21_X1 U11876 ( .A1(n21832), .A2(n1562), .B(n13731), .ZN(n30299) );
  INV_X1 U11877 ( .I(n31284), .ZN(n1857) );
  INV_X1 U11879 ( .I(n30048), .ZN(n30047) );
  NOR2_X1 U11882 ( .A1(n22014), .A2(n11656), .ZN(n30051) );
  NOR2_X1 U11883 ( .A1(n65), .A2(n1868), .ZN(n30385) );
  INV_X1 U11886 ( .I(n25013), .ZN(n30877) );
  BUF_X4 U11889 ( .I(n29862), .Z(n17413) );
  INV_X2 U11890 ( .I(n30395), .ZN(n1557) );
  BUF_X4 U11896 ( .I(n15772), .Z(n1868) );
  BUF_X4 U11897 ( .I(n58273), .Z(n1432) );
  CLKBUF_X2 U11900 ( .I(n30419), .Z(n22878) );
  INV_X2 U11901 ( .I(n28792), .ZN(n30526) );
  NOR2_X1 U11902 ( .A1(n28059), .A2(n16382), .ZN(n18867) );
  NAND2_X1 U11904 ( .A1(n13027), .A2(n28649), .ZN(n26114) );
  INV_X4 U11905 ( .I(n31242), .ZN(n1435) );
  NOR2_X1 U11914 ( .A1(n13028), .A2(n28654), .ZN(n13027) );
  OR2_X1 U11915 ( .A1(n19963), .A2(n19964), .Z(n24264) );
  INV_X1 U11916 ( .I(n4544), .ZN(n43880) );
  OAI21_X1 U11917 ( .A1(n12183), .A2(n27421), .B(n28254), .ZN(n12182) );
  NOR2_X1 U11920 ( .A1(n13918), .A2(n13917), .ZN(n19124) );
  NAND2_X1 U11921 ( .A1(n8806), .A2(n10404), .ZN(n9775) );
  AOI21_X1 U11924 ( .A1(n19170), .A2(n2136), .B(n2135), .ZN(n2134) );
  AOI21_X1 U11925 ( .A1(n29112), .A2(n29113), .B(n29111), .ZN(n29114) );
  OAI22_X1 U11926 ( .A1(n29137), .A2(n18377), .B1(n24941), .B2(n60841), .ZN(
        n8471) );
  NAND2_X1 U11930 ( .A1(n20608), .A2(n18037), .ZN(n18036) );
  OAI22_X1 U11931 ( .A1(n23937), .A2(n28648), .B1(n16185), .B2(n1889), .ZN(
        n27677) );
  NOR2_X1 U11932 ( .A1(n27018), .A2(n4986), .ZN(n21714) );
  NAND2_X1 U11933 ( .A1(n13919), .A2(n12085), .ZN(n13918) );
  INV_X1 U11935 ( .I(n7024), .ZN(n17235) );
  OR2_X1 U11939 ( .A1(n27893), .A2(n27892), .Z(n27894) );
  OAI21_X1 U11940 ( .A1(n27979), .A2(n27978), .B(n27977), .ZN(n18532) );
  AOI21_X1 U11943 ( .A1(n27182), .A2(n1354), .B(n27181), .ZN(n28103) );
  NAND3_X1 U11944 ( .A1(n27604), .A2(n27175), .A3(n14028), .ZN(n9470) );
  NAND2_X1 U11947 ( .A1(n93), .A2(n4059), .ZN(n28252) );
  NAND3_X1 U11949 ( .A1(n3469), .A2(n2661), .A3(n27934), .ZN(n2660) );
  INV_X1 U11953 ( .I(n29302), .ZN(n27496) );
  NOR2_X1 U11954 ( .A1(n7748), .A2(n26618), .ZN(n26664) );
  AOI21_X1 U11958 ( .A1(n28653), .A2(n28652), .B(n28651), .ZN(n28654) );
  NOR2_X1 U11960 ( .A1(n29146), .A2(n6913), .ZN(n3409) );
  NAND2_X1 U11961 ( .A1(n28798), .A2(n17522), .ZN(n28803) );
  INV_X1 U11962 ( .I(n24441), .ZN(n26739) );
  NAND2_X1 U11963 ( .A1(n26514), .A2(n28406), .ZN(n11075) );
  NAND2_X1 U11965 ( .A1(n27137), .A2(n11637), .ZN(n28325) );
  NOR3_X1 U11966 ( .A1(n29695), .A2(n10473), .A3(n491), .ZN(n20464) );
  OAI21_X1 U11969 ( .A1(n20609), .A2(n18038), .B(n28622), .ZN(n18037) );
  NAND2_X1 U11970 ( .A1(n29642), .A2(n1358), .ZN(n29634) );
  AND2_X1 U11971 ( .A1(n29302), .A2(n63883), .Z(n11162) );
  OAI21_X1 U11972 ( .A1(n27373), .A2(n29112), .B(n27375), .ZN(n2135) );
  NAND2_X1 U11973 ( .A1(n26990), .A2(n27323), .ZN(n6773) );
  NAND3_X1 U11975 ( .A1(n3470), .A2(n17047), .A3(n7371), .ZN(n3469) );
  NOR2_X1 U11977 ( .A1(n27716), .A2(n1570), .ZN(n27719) );
  NOR2_X1 U11979 ( .A1(n7499), .A2(n1320), .ZN(n27264) );
  NAND2_X1 U11980 ( .A1(n62083), .A2(n64174), .ZN(n28367) );
  AND3_X1 U11981 ( .A1(n28238), .A2(n28239), .A3(n28237), .Z(n28248) );
  AOI22_X1 U11986 ( .A1(n27929), .A2(n27928), .B1(n16654), .B2(n27927), .ZN(
        n17249) );
  NOR2_X1 U11987 ( .A1(n17451), .A2(n29147), .ZN(n17248) );
  INV_X1 U11988 ( .I(n8202), .ZN(n1877) );
  NAND2_X1 U11991 ( .A1(n1891), .A2(n8202), .ZN(n7630) );
  NAND2_X1 U11993 ( .A1(n28639), .A2(n27675), .ZN(n3749) );
  AND2_X1 U11994 ( .A1(n26660), .A2(n26665), .Z(n13382) );
  INV_X1 U11997 ( .I(n26964), .ZN(n1882) );
  NOR2_X1 U12001 ( .A1(n26043), .A2(n27846), .ZN(n20148) );
  INV_X1 U12002 ( .I(n27360), .ZN(n1884) );
  INV_X1 U12003 ( .I(n28308), .ZN(n1879) );
  NAND2_X1 U12005 ( .A1(n28162), .A2(n10236), .ZN(n29320) );
  NAND2_X1 U12006 ( .A1(n29694), .A2(n20581), .ZN(n13071) );
  NOR2_X1 U12007 ( .A1(n1279), .A2(n22604), .ZN(n4488) );
  NAND2_X1 U12008 ( .A1(n20665), .A2(n22514), .ZN(n26929) );
  NOR2_X1 U12010 ( .A1(n11573), .A2(n29168), .ZN(n11572) );
  AOI21_X1 U12011 ( .A1(n61177), .A2(n15650), .B(n60355), .ZN(n27095) );
  NAND2_X1 U12013 ( .A1(n29107), .A2(n60171), .ZN(n23466) );
  NAND2_X1 U12014 ( .A1(n29105), .A2(n63850), .ZN(n27017) );
  NOR2_X1 U12016 ( .A1(n266), .A2(n24940), .ZN(n27929) );
  OAI21_X1 U12018 ( .A1(n20561), .A2(n28622), .B(n29712), .ZN(n28467) );
  NAND2_X1 U12019 ( .A1(n29171), .A2(n11514), .ZN(n27287) );
  NAND2_X1 U12020 ( .A1(n28008), .A2(n3256), .ZN(n3255) );
  INV_X1 U12022 ( .I(n29168), .ZN(n27285) );
  NAND2_X1 U12023 ( .A1(n17747), .A2(n29142), .ZN(n29143) );
  INV_X1 U12024 ( .I(n27123), .ZN(n27022) );
  OAI21_X1 U12026 ( .A1(n28379), .A2(n13704), .B(n7129), .ZN(n27556) );
  INV_X1 U12027 ( .I(n28027), .ZN(n27959) );
  NOR2_X1 U12028 ( .A1(n28549), .A2(n28557), .ZN(n12109) );
  NOR2_X1 U12031 ( .A1(n1279), .A2(n64174), .ZN(n28370) );
  NOR2_X1 U12033 ( .A1(n26043), .A2(n28510), .ZN(n27847) );
  NOR2_X1 U12034 ( .A1(n29141), .A2(n17747), .ZN(n27933) );
  AND2_X1 U12036 ( .A1(n26613), .A2(n26612), .Z(n14134) );
  NOR2_X1 U12037 ( .A1(n29621), .A2(n22720), .ZN(n28835) );
  INV_X1 U12038 ( .I(n28551), .ZN(n1564) );
  BUF_X2 U12039 ( .I(n20860), .Z(n8296) );
  NAND2_X1 U12041 ( .A1(n7452), .A2(n61021), .ZN(n28013) );
  NAND2_X1 U12045 ( .A1(n12072), .A2(n21086), .ZN(n4187) );
  CLKBUF_X2 U12047 ( .I(n23549), .Z(n22720) );
  INV_X1 U12048 ( .I(n28342), .ZN(n18931) );
  NAND2_X1 U12049 ( .A1(n1322), .A2(n23170), .ZN(n28226) );
  BUF_X2 U12050 ( .I(n23814), .Z(n10544) );
  OR2_X1 U12055 ( .A1(n28312), .A2(n28299), .Z(n27169) );
  NAND2_X1 U12058 ( .A1(n5306), .A2(n28259), .ZN(n27941) );
  CLKBUF_X2 U12059 ( .I(n28311), .Z(n23840) );
  BUF_X2 U12064 ( .I(n23608), .Z(n21068) );
  INV_X1 U12065 ( .I(n27569), .ZN(n1885) );
  BUF_X2 U12068 ( .I(n28054), .Z(n7438) );
  BUF_X2 U12069 ( .I(n26945), .Z(n29628) );
  CLKBUF_X2 U12070 ( .I(n23917), .Z(n10321) );
  INV_X1 U12074 ( .I(n12739), .ZN(n29617) );
  INV_X1 U12078 ( .I(n28260), .ZN(n13194) );
  CLKBUF_X2 U12079 ( .I(n28221), .Z(n24060) );
  INV_X2 U12081 ( .I(n23917), .ZN(n7886) );
  INV_X4 U12083 ( .I(n17747), .ZN(n24940) );
  INV_X4 U12087 ( .I(n29690), .ZN(n28639) );
  INV_X1 U12091 ( .I(n3482), .ZN(n2067) );
  BUF_X2 U12092 ( .I(n23158), .Z(n22765) );
  INV_X2 U12096 ( .I(n5935), .ZN(n1445) );
  INV_X2 U12098 ( .I(n51492), .ZN(n56762) );
  CLKBUF_X2 U12103 ( .I(Key[47]), .Z(n24535) );
  CLKBUF_X2 U12104 ( .I(Key[26]), .Z(n53487) );
  CLKBUF_X2 U12105 ( .I(Key[128]), .Z(n55777) );
  CLKBUF_X4 U12108 ( .I(Key[114]), .Z(n55516) );
  BUF_X2 U12109 ( .I(Key[162]), .Z(n50494) );
  CLKBUF_X2 U12111 ( .I(Key[0]), .Z(n52900) );
  CLKBUF_X2 U12112 ( .I(Key[143]), .Z(n56124) );
  CLKBUF_X2 U12116 ( .I(Key[96]), .Z(n55118) );
  CLKBUF_X2 U12119 ( .I(Key[140]), .Z(n56040) );
  NAND3_X1 U12120 ( .A1(n6664), .A2(n55609), .A3(n55608), .ZN(n6663) );
  NOR3_X1 U12121 ( .A1(n1183), .A2(n9405), .A3(n9404), .ZN(n9403) );
  NAND2_X1 U12123 ( .A1(n16592), .A2(n20376), .ZN(n14842) );
  NOR2_X1 U12125 ( .A1(n2832), .A2(n2830), .ZN(n2829) );
  AOI21_X1 U12127 ( .A1(n56324), .A2(n56312), .B(n9114), .ZN(n9113) );
  OAI21_X1 U12128 ( .A1(n56314), .A2(n9116), .B(n61727), .ZN(n9115) );
  OAI21_X1 U12133 ( .A1(n53331), .A2(n60517), .B(n11962), .ZN(n16780) );
  NAND4_X1 U12134 ( .A1(n53822), .A2(n53045), .A3(n53046), .A4(n53800), .ZN(
        n17641) );
  NOR3_X1 U12136 ( .A1(n53172), .A2(n53171), .A3(n53173), .ZN(n10060) );
  OAI21_X1 U12137 ( .A1(n7566), .A2(n7565), .B(n56961), .ZN(n56974) );
  NAND2_X1 U12139 ( .A1(n53720), .A2(n53737), .ZN(n53754) );
  NAND3_X1 U12140 ( .A1(n12432), .A2(n55832), .A3(n55814), .ZN(n12431) );
  OAI21_X1 U12141 ( .A1(n55824), .A2(n55825), .B(n60855), .ZN(n12430) );
  NOR2_X1 U12142 ( .A1(n56960), .A2(n56959), .ZN(n7566) );
  NAND2_X1 U12143 ( .A1(n1161), .A2(n53505), .ZN(n53523) );
  NAND2_X1 U12144 ( .A1(n57156), .A2(n57124), .ZN(n57114) );
  NOR3_X1 U12145 ( .A1(n53252), .A2(n53253), .A3(n1164), .ZN(n19670) );
  OAI22_X1 U12146 ( .A1(n54203), .A2(n54188), .B1(n54175), .B2(n54118), .ZN(
        n2957) );
  NAND2_X1 U12147 ( .A1(n53645), .A2(n2746), .ZN(n2744) );
  OAI21_X1 U12148 ( .A1(n53149), .A2(n53148), .B(n3284), .ZN(n53150) );
  NOR2_X1 U12150 ( .A1(n11328), .A2(n61971), .ZN(n11327) );
  NAND4_X1 U12153 ( .A1(n54736), .A2(n23448), .A3(n54704), .A4(n54703), .ZN(
        n54705) );
  NAND2_X1 U12154 ( .A1(n19073), .A2(n1585), .ZN(n19072) );
  OR2_X1 U12155 ( .A1(n20957), .A2(n25393), .Z(n56343) );
  NOR3_X1 U12157 ( .A1(n55596), .A2(n55595), .A3(n19183), .ZN(n55599) );
  INV_X1 U12158 ( .I(n17893), .ZN(n15239) );
  NOR2_X1 U12160 ( .A1(n55226), .A2(n1587), .ZN(n7241) );
  NOR2_X1 U12163 ( .A1(n53966), .A2(n6135), .ZN(n53925) );
  OAI21_X1 U12164 ( .A1(n56157), .A2(n56158), .B(n56184), .ZN(n12532) );
  NAND2_X1 U12165 ( .A1(n1586), .A2(n20985), .ZN(n54427) );
  NAND2_X1 U12166 ( .A1(n56959), .A2(n1583), .ZN(n56908) );
  NAND2_X1 U12168 ( .A1(n23631), .A2(n1583), .ZN(n18111) );
  OAI21_X1 U12169 ( .A1(n62699), .A2(n55166), .B(n55163), .ZN(n55122) );
  AND2_X1 U12171 ( .A1(n55643), .A2(n55639), .Z(n19120) );
  NOR2_X1 U12172 ( .A1(n25172), .A2(n54582), .ZN(n14491) );
  INV_X1 U12173 ( .I(n56176), .ZN(n11274) );
  NOR2_X1 U12176 ( .A1(n5476), .A2(n4688), .ZN(n11325) );
  NOR3_X1 U12178 ( .A1(n55786), .A2(n55820), .A3(n60855), .ZN(n11684) );
  NOR2_X1 U12179 ( .A1(n54409), .A2(n6091), .ZN(n54388) );
  INV_X1 U12181 ( .I(n2784), .ZN(n55141) );
  NOR2_X1 U12182 ( .A1(n20735), .A2(n26135), .ZN(n3448) );
  CLKBUF_X2 U12185 ( .I(n53740), .Z(n7240) );
  BUF_X2 U12188 ( .I(n56344), .Z(n22891) );
  NAND2_X1 U12191 ( .A1(n11622), .A2(n11556), .ZN(n54395) );
  NOR2_X1 U12193 ( .A1(n55147), .A2(n62699), .ZN(n55142) );
  NAND3_X1 U12194 ( .A1(n22197), .A2(n18499), .A3(n50463), .ZN(n9617) );
  AOI21_X1 U12203 ( .A1(n17838), .A2(n51966), .B(n17836), .ZN(n17835) );
  NAND2_X1 U12204 ( .A1(n53912), .A2(n5025), .ZN(n10245) );
  OAI21_X1 U12209 ( .A1(n11680), .A2(n11679), .B(n60370), .ZN(n5041) );
  NOR2_X1 U12213 ( .A1(n11804), .A2(n12469), .ZN(n11803) );
  NAND2_X1 U12214 ( .A1(n14377), .A2(n54102), .ZN(n10529) );
  NAND2_X1 U12215 ( .A1(n13473), .A2(n22542), .ZN(n9839) );
  NOR2_X1 U12216 ( .A1(n54106), .A2(n54105), .ZN(n2987) );
  INV_X1 U12217 ( .I(n53911), .ZN(n53912) );
  OAI21_X1 U12218 ( .A1(n53619), .A2(n15362), .B(n53431), .ZN(n53432) );
  AOI21_X1 U12221 ( .A1(n20016), .A2(n51882), .B(n55718), .ZN(n20015) );
  NAND2_X1 U12223 ( .A1(n55718), .A2(n23919), .ZN(n4374) );
  OAI21_X1 U12228 ( .A1(n20613), .A2(n54107), .B(n9137), .ZN(n11939) );
  NAND3_X1 U12229 ( .A1(n57239), .A2(n56369), .A3(n56370), .ZN(n5886) );
  OAI21_X1 U12230 ( .A1(n24463), .A2(n24466), .B(n55453), .ZN(n23454) );
  NOR2_X1 U12233 ( .A1(n53533), .A2(n20630), .ZN(n17259) );
  OAI21_X1 U12236 ( .A1(n53231), .A2(n59858), .B(n20342), .ZN(n20341) );
  AOI21_X1 U12237 ( .A1(n53219), .A2(n1151), .B(n53218), .ZN(n6953) );
  NAND2_X1 U12238 ( .A1(n51253), .A2(n56394), .ZN(n12534) );
  NAND2_X1 U12239 ( .A1(n19971), .A2(n55685), .ZN(n11164) );
  OAI21_X1 U12240 ( .A1(n57191), .A2(n57691), .B(n24321), .ZN(n5420) );
  AOI21_X1 U12242 ( .A1(n16115), .A2(n1369), .B(n50880), .ZN(n51258) );
  OAI21_X1 U12246 ( .A1(n54984), .A2(n10551), .B(n63708), .ZN(n11549) );
  NOR2_X1 U12247 ( .A1(n1598), .A2(n1286), .ZN(n9407) );
  AOI21_X1 U12249 ( .A1(n11118), .A2(n56565), .B(n56397), .ZN(n7762) );
  OAI22_X1 U12250 ( .A1(n56278), .A2(n51264), .B1(n56568), .B2(n56565), .ZN(
        n7766) );
  NAND2_X1 U12251 ( .A1(n18294), .A2(n19971), .ZN(n11010) );
  NOR2_X1 U12252 ( .A1(n18323), .A2(n56563), .ZN(n6944) );
  INV_X1 U12257 ( .I(n4319), .ZN(n54607) );
  AND2_X1 U12259 ( .A1(n61914), .A2(n51453), .Z(n21070) );
  NAND2_X1 U12260 ( .A1(n8513), .A2(n2180), .ZN(n52923) );
  NAND2_X1 U12262 ( .A1(n53384), .A2(n23974), .ZN(n53197) );
  OAI21_X1 U12263 ( .A1(n1608), .A2(n54082), .B(n3664), .ZN(n54083) );
  OR2_X1 U12268 ( .A1(n23401), .A2(n53198), .Z(n52848) );
  NOR2_X1 U12269 ( .A1(n55922), .A2(n24404), .ZN(n11717) );
  AND3_X1 U12272 ( .A1(n53223), .A2(n64521), .A3(n58300), .Z(n53224) );
  AOI21_X1 U12276 ( .A1(n53449), .A2(n57183), .B(n53572), .ZN(n53225) );
  OAI22_X1 U12279 ( .A1(n4195), .A2(n58626), .B1(n4194), .B2(n55679), .ZN(
        n55682) );
  NOR2_X1 U12281 ( .A1(n54320), .A2(n64307), .ZN(n5735) );
  AOI21_X1 U12282 ( .A1(n18195), .A2(n56397), .B(n11989), .ZN(n7765) );
  AOI21_X1 U12283 ( .A1(n53209), .A2(n3127), .B(n23563), .ZN(n12788) );
  OR2_X1 U12285 ( .A1(n23095), .A2(n23334), .Z(n51345) );
  NAND2_X1 U12291 ( .A1(n56227), .A2(n56226), .ZN(n56425) );
  NAND2_X1 U12292 ( .A1(n14142), .A2(n55677), .ZN(n4836) );
  NAND2_X1 U12296 ( .A1(n54596), .A2(n54088), .ZN(n7788) );
  INV_X4 U12303 ( .I(n26089), .ZN(n23025) );
  INV_X1 U12306 ( .I(n13025), .ZN(n10949) );
  INV_X4 U12307 ( .I(n55440), .ZN(n14226) );
  INV_X2 U12313 ( .I(n9159), .ZN(n1459) );
  INV_X1 U12325 ( .I(n9876), .ZN(n12094) );
  INV_X1 U12326 ( .I(n25794), .ZN(n11480) );
  CLKBUF_X2 U12327 ( .I(n51508), .Z(n20723) );
  BUF_X2 U12329 ( .I(n51690), .Z(n22845) );
  INV_X1 U12332 ( .I(n49353), .ZN(n10157) );
  NAND2_X1 U12333 ( .A1(n47557), .A2(n24804), .ZN(n13095) );
  OAI21_X1 U12336 ( .A1(n49185), .A2(n49406), .B(n49410), .ZN(n49186) );
  OAI21_X1 U12341 ( .A1(n3846), .A2(n49195), .B(n3844), .ZN(n47557) );
  BUF_X2 U12344 ( .I(n52176), .Z(n13325) );
  NAND3_X1 U12345 ( .A1(n50268), .A2(n49946), .A3(n61083), .ZN(n25541) );
  OAI22_X1 U12347 ( .A1(n12752), .A2(n12753), .B1(n48846), .B2(n48845), .ZN(
        n12751) );
  INV_X1 U12350 ( .I(n13317), .ZN(n15526) );
  NAND2_X1 U12352 ( .A1(n6679), .A2(n48327), .ZN(n48329) );
  NAND2_X1 U12358 ( .A1(n49342), .A2(n49341), .ZN(n49354) );
  OAI21_X1 U12359 ( .A1(n49805), .A2(n49804), .B(n11219), .ZN(n11218) );
  INV_X1 U12367 ( .I(n8433), .ZN(n48066) );
  AOI21_X1 U12368 ( .A1(n48308), .A2(n59086), .B(n48307), .ZN(n48311) );
  AOI21_X1 U12370 ( .A1(n48745), .A2(n50267), .B(n50268), .ZN(n10714) );
  AOI21_X1 U12372 ( .A1(n61375), .A2(n16543), .B(n49986), .ZN(n49206) );
  NOR2_X1 U12373 ( .A1(n24770), .A2(n49977), .ZN(n15301) );
  NOR3_X1 U12374 ( .A1(n57290), .A2(n49223), .A3(n49227), .ZN(n24267) );
  NOR2_X1 U12376 ( .A1(n50001), .A2(n16676), .ZN(n16675) );
  AOI21_X1 U12380 ( .A1(n49038), .A2(n46852), .B(n46851), .ZN(n46853) );
  NAND2_X1 U12382 ( .A1(n1631), .A2(n49498), .ZN(n16089) );
  NAND2_X1 U12384 ( .A1(n57267), .A2(n1261), .ZN(n48846) );
  AND2_X1 U12388 ( .A1(n50428), .A2(n25680), .Z(n3679) );
  AOI21_X1 U12392 ( .A1(n49520), .A2(n11781), .B(n57267), .ZN(n18431) );
  NOR2_X1 U12396 ( .A1(n7866), .A2(n50240), .ZN(n47759) );
  INV_X1 U12399 ( .I(n48412), .ZN(n48820) );
  OAI21_X1 U12400 ( .A1(n48418), .A2(n11058), .B(n48065), .ZN(n11057) );
  NAND2_X1 U12401 ( .A1(n5568), .A2(n48395), .ZN(n5567) );
  NAND2_X1 U12402 ( .A1(n19042), .A2(n49484), .ZN(n7746) );
  AOI21_X1 U12403 ( .A1(n47966), .A2(n13120), .B(n47965), .ZN(n3703) );
  OAI21_X1 U12406 ( .A1(n7866), .A2(n1632), .B(n4109), .ZN(n50442) );
  AOI22_X1 U12407 ( .A1(n7866), .A2(n16211), .B1(n25744), .B2(n50443), .ZN(
        n50450) );
  INV_X1 U12408 ( .I(n26102), .ZN(n49781) );
  NOR2_X1 U12412 ( .A1(n25459), .A2(n49017), .ZN(n15472) );
  OR2_X1 U12415 ( .A1(n1644), .A2(n48688), .Z(n4412) );
  INV_X1 U12418 ( .I(n49511), .ZN(n16483) );
  OAI21_X1 U12422 ( .A1(n48323), .A2(n49014), .B(n48031), .ZN(n7015) );
  INV_X1 U12423 ( .I(n49356), .ZN(n49436) );
  OAI21_X1 U12424 ( .A1(n49762), .A2(n48897), .B(n19302), .ZN(n4598) );
  NAND2_X1 U12429 ( .A1(n49064), .A2(n49063), .ZN(n49067) );
  AOI21_X1 U12430 ( .A1(n57949), .A2(n4815), .B(n7078), .ZN(n48874) );
  AOI22_X1 U12431 ( .A1(n49926), .A2(n60772), .B1(n1636), .B2(n61835), .ZN(
        n6213) );
  INV_X1 U12435 ( .I(n50441), .ZN(n50232) );
  AND2_X1 U12436 ( .A1(n50401), .A2(n50081), .Z(n50076) );
  NAND2_X1 U12439 ( .A1(n49331), .A2(n15753), .ZN(n49326) );
  NOR2_X1 U12440 ( .A1(n15167), .A2(n50400), .ZN(n15166) );
  NOR2_X1 U12443 ( .A1(n22867), .A2(n19775), .ZN(n22489) );
  NAND2_X1 U12450 ( .A1(n49419), .A2(n1381), .ZN(n50075) );
  AOI21_X1 U12453 ( .A1(n25473), .A2(n62975), .B(n2477), .ZN(n48376) );
  NOR2_X1 U12454 ( .A1(n50375), .A2(n3031), .ZN(n46851) );
  OAI21_X1 U12455 ( .A1(n48680), .A2(n15737), .B(n48678), .ZN(n17165) );
  INV_X1 U12458 ( .I(n49077), .ZN(n49064) );
  NAND2_X1 U12459 ( .A1(n21367), .A2(n23912), .ZN(n49267) );
  INV_X1 U12460 ( .I(n2477), .ZN(n48983) );
  INV_X1 U12463 ( .I(n14809), .ZN(n49924) );
  NAND2_X1 U12465 ( .A1(n19866), .A2(n15319), .ZN(n49552) );
  NOR2_X1 U12466 ( .A1(n5146), .A2(n49222), .ZN(n49463) );
  AND3_X1 U12469 ( .A1(n17906), .A2(n49372), .A3(n57473), .Z(n25263) );
  NOR2_X1 U12471 ( .A1(n50307), .A2(n50309), .ZN(n49650) );
  NAND2_X1 U12477 ( .A1(n49177), .A2(n12003), .ZN(n5545) );
  NOR2_X1 U12479 ( .A1(n10961), .A2(n49637), .ZN(n10960) );
  BUF_X4 U12480 ( .I(n23247), .Z(n8129) );
  AOI21_X1 U12482 ( .A1(n49686), .A2(n49371), .B(n49687), .ZN(n5497) );
  NOR2_X1 U12484 ( .A1(n23650), .A2(n50376), .ZN(n14065) );
  NOR2_X1 U12485 ( .A1(n14314), .A2(n14315), .ZN(n49900) );
  BUF_X4 U12489 ( .I(n8024), .Z(n1643) );
  NAND2_X1 U12493 ( .A1(n49767), .A2(n49777), .ZN(n4098) );
  BUF_X4 U12498 ( .I(n48141), .Z(n50340) );
  NOR2_X1 U12499 ( .A1(n8695), .A2(n1651), .ZN(n14185) );
  NAND2_X1 U12506 ( .A1(n6283), .A2(n22910), .ZN(n6282) );
  INV_X4 U12507 ( .I(n49720), .ZN(n1473) );
  NAND2_X1 U12516 ( .A1(n46816), .A2(n21304), .ZN(n14789) );
  NOR2_X1 U12517 ( .A1(n58809), .A2(n16416), .ZN(n16415) );
  NAND4_X1 U12518 ( .A1(n62290), .A2(n48101), .A3(n48104), .A4(n23850), .ZN(
        n3093) );
  NAND2_X1 U12526 ( .A1(n1112), .A2(n8923), .ZN(n45188) );
  NAND3_X1 U12528 ( .A1(n46096), .A2(n24801), .A3(n5771), .ZN(n8695) );
  NAND3_X1 U12530 ( .A1(n47396), .A2(n47867), .A3(n47869), .ZN(n47404) );
  NAND3_X1 U12531 ( .A1(n47869), .A2(n70), .A3(n24893), .ZN(n10590) );
  NAND2_X1 U12537 ( .A1(n46267), .A2(n47502), .ZN(n12823) );
  OR2_X1 U12538 ( .A1(n44702), .A2(n45781), .Z(n11444) );
  OAI21_X1 U12552 ( .A1(n8271), .A2(n8270), .B(n46063), .ZN(n21557) );
  NAND2_X1 U12558 ( .A1(n46482), .A2(n23018), .ZN(n12767) );
  AOI21_X1 U12560 ( .A1(n45946), .A2(n47574), .B(n18002), .ZN(n18001) );
  OAI22_X1 U12568 ( .A1(n10250), .A2(n48566), .B1(n13348), .B2(n48565), .ZN(
        n48568) );
  AOI21_X1 U12569 ( .A1(n47637), .A2(n47879), .B(n47636), .ZN(n15030) );
  NOR2_X1 U12570 ( .A1(n8224), .A2(n24114), .ZN(n9743) );
  NAND3_X1 U12572 ( .A1(n48582), .A2(n48581), .A3(n13587), .ZN(n13585) );
  NAND2_X1 U12578 ( .A1(n62748), .A2(n1652), .ZN(n2313) );
  OAI21_X1 U12579 ( .A1(n48651), .A2(n22605), .B(n12620), .ZN(n12619) );
  AOI21_X1 U12580 ( .A1(n46817), .A2(n14786), .B(n46758), .ZN(n14785) );
  OAI21_X1 U12581 ( .A1(n48657), .A2(n48658), .B(n48661), .ZN(n48663) );
  AOI21_X1 U12583 ( .A1(n11896), .A2(n5940), .B(n11901), .ZN(n11900) );
  NOR3_X1 U12584 ( .A1(n9453), .A2(n47361), .A3(n47360), .ZN(n9449) );
  AND3_X1 U12585 ( .A1(n46907), .A2(n1388), .A3(n18361), .Z(n46908) );
  NAND2_X1 U12586 ( .A1(n46980), .A2(n10055), .ZN(n45518) );
  OAI22_X1 U12588 ( .A1(n47857), .A2(n45447), .B1(n25006), .B2(n20912), .ZN(
        n3615) );
  NAND2_X1 U12591 ( .A1(n47800), .A2(n1385), .ZN(n6191) );
  NAND3_X1 U12592 ( .A1(n12723), .A2(n21793), .A3(n47259), .ZN(n12722) );
  NOR2_X1 U12593 ( .A1(n1266), .A2(n47407), .ZN(n13822) );
  NAND2_X1 U12595 ( .A1(n24291), .A2(n45194), .ZN(n18002) );
  NAND3_X1 U12596 ( .A1(n45810), .A2(n47141), .A3(n21451), .ZN(n10676) );
  NAND4_X1 U12597 ( .A1(n6081), .A2(n46913), .A3(n44660), .A4(n23990), .ZN(
        n44207) );
  NOR2_X1 U12599 ( .A1(n12025), .A2(n47690), .ZN(n12024) );
  NAND2_X1 U12602 ( .A1(n45957), .A2(n18951), .ZN(n3181) );
  NOR3_X1 U12608 ( .A1(n61216), .A2(n47422), .A3(n46843), .ZN(n46757) );
  NAND3_X1 U12610 ( .A1(n47373), .A2(n1654), .A3(n23934), .ZN(n14571) );
  AND2_X1 U12615 ( .A1(n23167), .A2(n177), .Z(n16276) );
  INV_X1 U12617 ( .I(n48224), .ZN(n11744) );
  NAND3_X1 U12619 ( .A1(n47517), .A2(n1086), .A3(n47516), .ZN(n10031) );
  NAND2_X1 U12629 ( .A1(n61720), .A2(n47682), .ZN(n13497) );
  NOR2_X1 U12630 ( .A1(n47798), .A2(n23180), .ZN(n18992) );
  NAND2_X1 U12633 ( .A1(n64766), .A2(n60138), .ZN(n21397) );
  AOI21_X1 U12634 ( .A1(n1080), .A2(n13258), .B(n23407), .ZN(n4261) );
  NAND3_X1 U12635 ( .A1(n22905), .A2(n45538), .A3(n1294), .ZN(n11062) );
  OR2_X1 U12639 ( .A1(n47845), .A2(n47844), .Z(n42617) );
  NOR2_X1 U12641 ( .A1(n47377), .A2(n65161), .ZN(n12498) );
  AND2_X1 U12642 ( .A1(n14474), .A2(n47718), .Z(n11908) );
  OAI21_X1 U12643 ( .A1(n8758), .A2(n23542), .B(n9851), .ZN(n21547) );
  OR2_X1 U12646 ( .A1(n47468), .A2(n4380), .Z(n9199) );
  AND3_X1 U12648 ( .A1(n16882), .A2(n48660), .A3(n47488), .Z(n25729) );
  NOR2_X1 U12649 ( .A1(n22468), .A2(n7541), .ZN(n11214) );
  OAI21_X1 U12652 ( .A1(n47559), .A2(n22537), .B(n47664), .ZN(n14456) );
  NAND2_X1 U12654 ( .A1(n47473), .A2(n1660), .ZN(n9176) );
  NOR2_X1 U12657 ( .A1(n48530), .A2(n21177), .ZN(n15163) );
  INV_X4 U12659 ( .I(n1388), .ZN(n15666) );
  NAND2_X1 U12660 ( .A1(n57677), .A2(n47482), .ZN(n19039) );
  OR2_X1 U12661 ( .A1(n45651), .A2(n64888), .Z(n45485) );
  INV_X1 U12665 ( .I(n3562), .ZN(n47237) );
  NAND2_X1 U12666 ( .A1(n47575), .A2(n1085), .ZN(n24291) );
  INV_X1 U12667 ( .I(n47494), .ZN(n11786) );
  INV_X1 U12672 ( .I(n48661), .ZN(n1476) );
  INV_X1 U12673 ( .I(n45536), .ZN(n44699) );
  INV_X1 U12675 ( .I(n47316), .ZN(n46923) );
  NOR2_X1 U12686 ( .A1(n23934), .A2(n21495), .ZN(n20112) );
  AND2_X1 U12687 ( .A1(n47270), .A2(n548), .Z(n47271) );
  OAI21_X1 U12689 ( .A1(n47736), .A2(n45908), .B(n47432), .ZN(n43749) );
  INV_X4 U12701 ( .I(n6938), .ZN(n1664) );
  INV_X2 U12702 ( .I(n16757), .ZN(n46244) );
  CLKBUF_X2 U12703 ( .I(n47472), .Z(n10055) );
  INV_X4 U12706 ( .I(n19935), .ZN(n47534) );
  BUF_X2 U12709 ( .I(n47011), .Z(n20090) );
  INV_X2 U12712 ( .I(n6055), .ZN(n1487) );
  INV_X1 U12716 ( .I(n44955), .ZN(n1673) );
  INV_X1 U12718 ( .I(n44479), .ZN(n1674) );
  BUF_X4 U12722 ( .I(n46442), .Z(n22376) );
  INV_X1 U12723 ( .I(n23641), .ZN(n14461) );
  BUF_X2 U12728 ( .I(n62518), .Z(n17902) );
  BUF_X2 U12729 ( .I(n46305), .Z(n22639) );
  INV_X1 U12737 ( .I(n16519), .ZN(n46428) );
  INV_X2 U12741 ( .I(n9378), .ZN(n1684) );
  NAND2_X1 U12748 ( .A1(n43203), .A2(n43202), .ZN(n19486) );
  NAND2_X1 U12751 ( .A1(n2689), .A2(n43584), .ZN(n2292) );
  AOI21_X1 U12753 ( .A1(n43575), .A2(n43574), .B(n5339), .ZN(n2688) );
  NOR2_X1 U12754 ( .A1(n9445), .A2(n9447), .ZN(n19342) );
  NOR2_X1 U12755 ( .A1(n37534), .A2(n15307), .ZN(n22318) );
  NOR2_X1 U12758 ( .A1(n42742), .A2(n42738), .ZN(n12666) );
  NAND2_X1 U12759 ( .A1(n7576), .A2(n986), .ZN(n9445) );
  AND2_X1 U12760 ( .A1(n43843), .A2(n11750), .Z(n11749) );
  OAI21_X1 U12762 ( .A1(n18021), .A2(n18022), .B(n8290), .ZN(n15174) );
  INV_X1 U12767 ( .I(n40912), .ZN(n4531) );
  NAND2_X1 U12771 ( .A1(n42864), .A2(n9080), .ZN(n8080) );
  NAND2_X1 U12773 ( .A1(n39014), .A2(n39013), .ZN(n13262) );
  NOR2_X1 U12775 ( .A1(n42843), .A2(n8290), .ZN(n15175) );
  NOR2_X1 U12776 ( .A1(n9034), .A2(n1695), .ZN(n3806) );
  NOR2_X1 U12778 ( .A1(n13621), .A2(n13882), .ZN(n15064) );
  NAND2_X1 U12780 ( .A1(n43840), .A2(n19487), .ZN(n11750) );
  AND4_X1 U12784 ( .A1(n43703), .A2(n43702), .A3(n20242), .A4(n16527), .Z(
        n43704) );
  NOR2_X1 U12785 ( .A1(n42565), .A2(n23434), .ZN(n13528) );
  NAND3_X1 U12786 ( .A1(n11362), .A2(n15020), .A3(n43116), .ZN(n11365) );
  AOI21_X1 U12787 ( .A1(n43359), .A2(n13453), .B(n42732), .ZN(n13452) );
  NAND2_X1 U12791 ( .A1(n16890), .A2(n63455), .ZN(n18154) );
  NAND3_X1 U12792 ( .A1(n43955), .A2(n19742), .A3(n63455), .ZN(n11404) );
  AOI21_X1 U12793 ( .A1(n5801), .A2(n1709), .B(n11607), .ZN(n5800) );
  NAND3_X1 U12794 ( .A1(n43251), .A2(n43252), .A3(n43253), .ZN(n15813) );
  NOR3_X1 U12795 ( .A1(n43776), .A2(n43922), .A3(n43489), .ZN(n6072) );
  INV_X1 U12796 ( .I(n24518), .ZN(n41546) );
  NOR2_X1 U12801 ( .A1(n25600), .A2(n43948), .ZN(n43304) );
  AOI21_X1 U12802 ( .A1(n14408), .A2(n19742), .B(n43947), .ZN(n16940) );
  NAND2_X1 U12804 ( .A1(n3730), .A2(n39797), .ZN(n2854) );
  NOR2_X1 U12808 ( .A1(n9446), .A2(n7577), .ZN(n7576) );
  NAND3_X1 U12809 ( .A1(n3953), .A2(n6734), .A3(n7996), .ZN(n3952) );
  NOR2_X1 U12811 ( .A1(n8907), .A2(n8906), .ZN(n15490) );
  NAND2_X1 U12813 ( .A1(n15445), .A2(n9365), .ZN(n16341) );
  NAND3_X1 U12817 ( .A1(n20685), .A2(n3696), .A3(n60593), .ZN(n43653) );
  NOR2_X1 U12818 ( .A1(n21950), .A2(n10111), .ZN(n8469) );
  NAND2_X1 U12820 ( .A1(n41321), .A2(n2856), .ZN(n2855) );
  NOR2_X1 U12821 ( .A1(n63747), .A2(n14051), .ZN(n8906) );
  NAND2_X1 U12823 ( .A1(n19346), .A2(n6007), .ZN(n20294) );
  AOI21_X1 U12825 ( .A1(n43476), .A2(n13751), .B(n43475), .ZN(n43477) );
  NOR2_X1 U12826 ( .A1(n43712), .A2(n43992), .ZN(n20320) );
  NAND2_X1 U12827 ( .A1(n40899), .A2(n1699), .ZN(n40900) );
  AOI21_X1 U12829 ( .A1(n43607), .A2(n43606), .B(n12970), .ZN(n12969) );
  NAND2_X1 U12834 ( .A1(n41693), .A2(n42395), .ZN(n8429) );
  NAND2_X1 U12835 ( .A1(n16649), .A2(n43102), .ZN(n9446) );
  NOR2_X1 U12837 ( .A1(n43564), .A2(n62997), .ZN(n13201) );
  NAND3_X1 U12838 ( .A1(n1333), .A2(n2797), .A3(n43897), .ZN(n43899) );
  AND3_X1 U12840 ( .A1(n46331), .A2(n42642), .A3(n43189), .Z(n41765) );
  NOR2_X1 U12841 ( .A1(n43507), .A2(n43502), .ZN(n43190) );
  AOI21_X1 U12842 ( .A1(n15792), .A2(n61745), .B(n14051), .ZN(n3965) );
  CLKBUF_X2 U12843 ( .I(n42422), .Z(n11362) );
  NAND2_X1 U12844 ( .A1(n43325), .A2(n43326), .ZN(n15032) );
  AND2_X1 U12845 ( .A1(n42780), .A2(n9792), .Z(n7637) );
  AND3_X1 U12849 ( .A1(n43875), .A2(n11608), .A3(n7950), .Z(n5827) );
  NOR2_X1 U12850 ( .A1(n1692), .A2(n64323), .ZN(n7514) );
  NOR2_X1 U12854 ( .A1(n39878), .A2(n43102), .ZN(n42011) );
  NAND3_X1 U12855 ( .A1(n1297), .A2(n61171), .A3(n41584), .ZN(n41585) );
  NOR2_X1 U12856 ( .A1(n43540), .A2(n279), .ZN(n24216) );
  INV_X1 U12862 ( .I(n8687), .ZN(n41790) );
  NOR2_X1 U12863 ( .A1(n57177), .A2(n43130), .ZN(n39802) );
  NAND2_X1 U12865 ( .A1(n12124), .A2(n1392), .ZN(n11817) );
  OAI21_X1 U12866 ( .A1(n43655), .A2(n20183), .B(n64323), .ZN(n3485) );
  NAND2_X1 U12868 ( .A1(n1697), .A2(n20922), .ZN(n40280) );
  NOR2_X1 U12870 ( .A1(n42865), .A2(n4575), .ZN(n4574) );
  INV_X1 U12871 ( .I(n10617), .ZN(n42924) );
  NOR2_X1 U12874 ( .A1(n4789), .A2(n43165), .ZN(n43168) );
  NAND2_X1 U12875 ( .A1(n1705), .A2(n4274), .ZN(n4277) );
  NAND2_X1 U12878 ( .A1(n1700), .A2(n42386), .ZN(n42379) );
  NAND2_X1 U12879 ( .A1(n43335), .A2(n63293), .ZN(n12759) );
  NAND2_X1 U12881 ( .A1(n43140), .A2(n20183), .ZN(n4765) );
  INV_X1 U12882 ( .I(n15502), .ZN(n43207) );
  OAI21_X1 U12883 ( .A1(n42734), .A2(n1715), .B(n41550), .ZN(n13454) );
  OAI22_X1 U12890 ( .A1(n21325), .A2(n21326), .B1(n42138), .B2(n9914), .ZN(
        n3634) );
  NAND2_X1 U12892 ( .A1(n63205), .A2(n13596), .ZN(n13595) );
  INV_X1 U12897 ( .I(n13854), .ZN(n16740) );
  NAND2_X1 U12899 ( .A1(n13478), .A2(n43460), .ZN(n13476) );
  OR3_X1 U12905 ( .A1(n1708), .A2(n62299), .A3(n43601), .Z(n40601) );
  INV_X1 U12906 ( .I(n8537), .ZN(n41661) );
  NAND2_X1 U12908 ( .A1(n20452), .A2(n23434), .ZN(n20451) );
  NAND2_X1 U12909 ( .A1(n63205), .A2(n63529), .ZN(n15218) );
  NAND2_X1 U12910 ( .A1(n24002), .A2(n11747), .ZN(n11746) );
  NAND2_X1 U12911 ( .A1(n43039), .A2(n61171), .ZN(n39015) );
  NOR2_X1 U12916 ( .A1(n18051), .A2(n19517), .ZN(n12124) );
  NAND2_X1 U12917 ( .A1(n43268), .A2(n65217), .ZN(n4335) );
  OR2_X1 U12918 ( .A1(n25440), .A2(n43272), .Z(n2856) );
  NAND2_X1 U12921 ( .A1(n20942), .A2(n24360), .ZN(n15089) );
  NOR2_X1 U12922 ( .A1(n8351), .A2(n1714), .ZN(n8350) );
  NAND2_X1 U12927 ( .A1(n43923), .A2(n21073), .ZN(n1941) );
  NAND2_X1 U12935 ( .A1(n1270), .A2(n61186), .ZN(n42808) );
  NAND2_X1 U12938 ( .A1(n44226), .A2(n6007), .ZN(n43988) );
  NAND2_X1 U12939 ( .A1(n43980), .A2(n6007), .ZN(n44228) );
  INV_X4 U12942 ( .I(n23709), .ZN(n43150) );
  AND2_X1 U12944 ( .A1(n3302), .A2(n43124), .Z(n3327) );
  OR2_X1 U12946 ( .A1(n43225), .A2(n24250), .Z(n19365) );
  INV_X1 U12948 ( .I(n43978), .ZN(n1719) );
  CLKBUF_X4 U12950 ( .I(n42313), .Z(n16880) );
  CLKBUF_X4 U12955 ( .I(n42313), .Z(n44226) );
  OAI21_X1 U12957 ( .A1(n3564), .A2(n42261), .B(n3563), .ZN(n43978) );
  AOI22_X1 U12958 ( .A1(n7929), .A2(n61394), .B1(n41302), .B2(n42237), .ZN(
        n7924) );
  NAND2_X1 U12961 ( .A1(n2877), .A2(n41149), .ZN(n18593) );
  NAND2_X1 U12962 ( .A1(n41952), .A2(n41953), .ZN(n16773) );
  OAI21_X1 U12965 ( .A1(n38275), .A2(n41941), .B(n61394), .ZN(n7749) );
  CLKBUF_X2 U12966 ( .I(n9135), .Z(n8139) );
  AOI21_X1 U12972 ( .A1(n9526), .A2(n9527), .B(n59280), .ZN(n12036) );
  OAI21_X1 U12973 ( .A1(n15776), .A2(n38135), .B(n16297), .ZN(n20075) );
  OAI22_X1 U12976 ( .A1(n41448), .A2(n25430), .B1(n64773), .B2(n41446), .ZN(
        n41450) );
  OAI21_X1 U12979 ( .A1(n41827), .A2(n10479), .B(n4763), .ZN(n41828) );
  NOR2_X1 U12981 ( .A1(n7647), .A2(n7646), .ZN(n7645) );
  OAI21_X1 U12982 ( .A1(n42480), .A2(n42477), .B(n18278), .ZN(n40037) );
  NAND2_X1 U12984 ( .A1(n40069), .A2(n1721), .ZN(n11129) );
  AOI21_X1 U12986 ( .A1(n41803), .A2(n1727), .B(n7337), .ZN(n17076) );
  NOR2_X1 U12992 ( .A1(n6347), .A2(n6346), .ZN(n21165) );
  AND2_X1 U12995 ( .A1(n41461), .A2(n41460), .Z(n3666) );
  OAI21_X1 U12997 ( .A1(n42279), .A2(n58262), .B(n40817), .ZN(n40822) );
  AND2_X1 U13002 ( .A1(n1725), .A2(n59577), .Z(n9527) );
  OAI21_X1 U13007 ( .A1(n40699), .A2(n60653), .B(n41436), .ZN(n17833) );
  AOI21_X1 U13008 ( .A1(n10133), .A2(n41179), .B(n41178), .ZN(n41180) );
  NOR2_X1 U13009 ( .A1(n22943), .A2(n21865), .ZN(n41843) );
  AOI22_X1 U13011 ( .A1(n13309), .A2(n39099), .B1(n13311), .B2(n20726), .ZN(
        n13304) );
  NOR2_X1 U13013 ( .A1(n57545), .A2(n59976), .ZN(n2586) );
  NAND2_X1 U13014 ( .A1(n60509), .A2(n9716), .ZN(n42268) );
  INV_X1 U13018 ( .I(n64773), .ZN(n39844) );
  NAND3_X1 U13019 ( .A1(n41446), .A2(n64773), .A3(n41437), .ZN(n12191) );
  NAND2_X1 U13020 ( .A1(n1723), .A2(n22638), .ZN(n11646) );
  NAND2_X1 U13021 ( .A1(n41458), .A2(n41457), .ZN(n14950) );
  NOR2_X1 U13023 ( .A1(n61435), .A2(n42230), .ZN(n7926) );
  OAI22_X1 U13025 ( .A1(n42269), .A2(n10670), .B1(n42260), .B2(n10668), .ZN(
        n41099) );
  NAND3_X1 U13026 ( .A1(n39039), .A2(n40670), .A3(n39038), .ZN(n39045) );
  AOI21_X1 U13027 ( .A1(n41016), .A2(n1275), .B(n7648), .ZN(n7647) );
  INV_X1 U13028 ( .I(n41248), .ZN(n3457) );
  NAND2_X1 U13029 ( .A1(n40848), .A2(n41885), .ZN(n40862) );
  OAI21_X1 U13030 ( .A1(n41867), .A2(n42520), .B(n41868), .ZN(n25219) );
  NAND2_X1 U13037 ( .A1(n41437), .A2(n23967), .ZN(n10877) );
  OAI22_X1 U13039 ( .A1(n40990), .A2(n12409), .B1(n3356), .B2(n40995), .ZN(
        n10800) );
  NAND2_X1 U13041 ( .A1(n1219), .A2(n41447), .ZN(n6993) );
  AOI21_X1 U13042 ( .A1(n42455), .A2(n16226), .B(n42450), .ZN(n8069) );
  NOR2_X1 U13043 ( .A1(n38045), .A2(n39104), .ZN(n23551) );
  INV_X1 U13046 ( .I(n41155), .ZN(n39019) );
  AOI22_X1 U13048 ( .A1(n15345), .A2(n41235), .B1(n41405), .B2(n1303), .ZN(
        n8917) );
  AOI21_X1 U13050 ( .A1(n40649), .A2(n40648), .B(n22005), .ZN(n22004) );
  NAND2_X1 U13051 ( .A1(n11895), .A2(n57258), .ZN(n12453) );
  AOI21_X1 U13054 ( .A1(n63174), .A2(n1404), .B(n11194), .ZN(n11193) );
  OAI21_X1 U13055 ( .A1(n40998), .A2(n12409), .B(n40211), .ZN(n38036) );
  NAND3_X1 U13056 ( .A1(n25138), .A2(n25140), .A3(n40523), .ZN(n20394) );
  NOR2_X1 U13057 ( .A1(n40657), .A2(n7327), .ZN(n7326) );
  NAND2_X1 U13058 ( .A1(n41192), .A2(n38675), .ZN(n22727) );
  NOR2_X1 U13059 ( .A1(n1745), .A2(n1730), .ZN(n6801) );
  NOR2_X1 U13060 ( .A1(n39959), .A2(n40568), .ZN(n16925) );
  NAND2_X1 U13061 ( .A1(n40990), .A2(n18706), .ZN(n39329) );
  OAI21_X1 U13066 ( .A1(n41311), .A2(n1746), .B(n10593), .ZN(n14916) );
  NAND2_X1 U13067 ( .A1(n2341), .A2(n1731), .ZN(n2340) );
  AND2_X1 U13068 ( .A1(n3946), .A2(n16680), .Z(n11096) );
  NOR2_X1 U13069 ( .A1(n41446), .A2(n277), .ZN(n8246) );
  OAI22_X1 U13070 ( .A1(n5938), .A2(n40403), .B1(n40771), .B2(n58794), .ZN(
        n38933) );
  OAI21_X1 U13073 ( .A1(n40609), .A2(n37530), .B(n58851), .ZN(n25285) );
  NOR2_X1 U13074 ( .A1(n64242), .A2(n6576), .ZN(n39417) );
  NAND2_X1 U13076 ( .A1(n41199), .A2(n40732), .ZN(n9776) );
  NAND2_X1 U13077 ( .A1(n39158), .A2(n40924), .ZN(n11042) );
  AND2_X1 U13078 ( .A1(n40313), .A2(n40314), .Z(n15671) );
  NOR2_X1 U13079 ( .A1(n41276), .A2(n41852), .ZN(n42303) );
  INV_X2 U13081 ( .I(n11084), .ZN(n6689) );
  NAND2_X1 U13082 ( .A1(n41152), .A2(n60139), .ZN(n38843) );
  NAND2_X1 U13083 ( .A1(n63435), .A2(n42237), .ZN(n12733) );
  NAND2_X1 U13084 ( .A1(n3306), .A2(n4968), .ZN(n37927) );
  NOR2_X1 U13087 ( .A1(n40379), .A2(n41435), .ZN(n8245) );
  NOR2_X1 U13089 ( .A1(n19343), .A2(n40568), .ZN(n4134) );
  NOR3_X1 U13090 ( .A1(n11819), .A2(n39957), .A3(n40443), .ZN(n4140) );
  NAND2_X1 U13091 ( .A1(n61417), .A2(n61638), .ZN(n2336) );
  NAND2_X1 U13092 ( .A1(n57207), .A2(n41852), .ZN(n15367) );
  AOI21_X1 U13093 ( .A1(n38197), .A2(n38196), .B(n61916), .ZN(n5814) );
  NAND3_X1 U13094 ( .A1(n18241), .A2(n22913), .A3(n1747), .ZN(n17965) );
  OR2_X1 U13096 ( .A1(n40356), .A2(n664), .Z(n16226) );
  NOR2_X1 U13097 ( .A1(n41039), .A2(n1747), .ZN(n6346) );
  NAND2_X1 U13098 ( .A1(n41944), .A2(n7519), .ZN(n5797) );
  NAND3_X1 U13101 ( .A1(n41898), .A2(n25837), .A3(n42267), .ZN(n41092) );
  NAND2_X1 U13102 ( .A1(n20190), .A2(n42230), .ZN(n9526) );
  NAND4_X1 U13103 ( .A1(n13984), .A2(n42488), .A3(n40123), .A4(n40091), .ZN(
        n40127) );
  NAND2_X1 U13104 ( .A1(n1732), .A2(n62106), .ZN(n2560) );
  OAI21_X1 U13108 ( .A1(n22617), .A2(n22913), .B(n1747), .ZN(n13139) );
  NOR2_X1 U13109 ( .A1(n22617), .A2(n38496), .ZN(n13136) );
  NOR2_X1 U13110 ( .A1(n61658), .A2(n10954), .ZN(n10956) );
  NAND2_X1 U13111 ( .A1(n41186), .A2(n10126), .ZN(n39037) );
  OAI21_X1 U13113 ( .A1(n10452), .A2(n41168), .B(n24781), .ZN(n41159) );
  NAND2_X1 U13114 ( .A1(n41452), .A2(n41451), .ZN(n41458) );
  NAND2_X1 U13116 ( .A1(n41405), .A2(n41237), .ZN(n15343) );
  NOR2_X1 U13117 ( .A1(n41399), .A2(n41412), .ZN(n15341) );
  NAND2_X1 U13118 ( .A1(n14306), .A2(n1275), .ZN(n16468) );
  NAND2_X1 U13120 ( .A1(n58851), .A2(n14306), .ZN(n17768) );
  NAND2_X1 U13123 ( .A1(n40142), .A2(n40210), .ZN(n18713) );
  NOR2_X1 U13124 ( .A1(n41152), .A2(n60139), .ZN(n3042) );
  NAND2_X1 U13125 ( .A1(n40526), .A2(n1740), .ZN(n15426) );
  NAND2_X1 U13127 ( .A1(n1963), .A2(n10554), .ZN(n41825) );
  AND2_X1 U13132 ( .A1(n40443), .A2(n41103), .Z(n5241) );
  NAND2_X1 U13134 ( .A1(n1748), .A2(n971), .ZN(n41111) );
  INV_X1 U13137 ( .I(n40074), .ZN(n40066) );
  INV_X1 U13138 ( .I(n61950), .ZN(n41236) );
  NAND2_X1 U13143 ( .A1(n40732), .A2(n40628), .ZN(n17581) );
  AND2_X1 U13144 ( .A1(n41810), .A2(n664), .Z(n41812) );
  NAND2_X1 U13148 ( .A1(n11677), .A2(n16158), .ZN(n41896) );
  INV_X1 U13149 ( .I(n41428), .ZN(n11718) );
  NAND2_X1 U13150 ( .A1(n18706), .A2(n23752), .ZN(n6752) );
  INV_X1 U13151 ( .I(n40737), .ZN(n41408) );
  NAND2_X1 U13155 ( .A1(n41805), .A2(n24066), .ZN(n6260) );
  BUF_X2 U13159 ( .I(n40928), .Z(n22809) );
  INV_X1 U13163 ( .I(n17915), .ZN(n40556) );
  INV_X2 U13176 ( .I(n6291), .ZN(n41160) );
  INV_X1 U13180 ( .I(n1749), .ZN(n15672) );
  BUF_X2 U13185 ( .I(n17078), .Z(n13695) );
  BUF_X2 U13188 ( .I(n22047), .Z(n7619) );
  INV_X1 U13195 ( .I(n37673), .ZN(n38386) );
  INV_X2 U13204 ( .I(n24274), .ZN(n1520) );
  INV_X2 U13207 ( .I(n20446), .ZN(n1522) );
  BUF_X2 U13209 ( .I(n37873), .Z(n23931) );
  INV_X1 U13212 ( .I(n21239), .ZN(n9371) );
  AND2_X1 U13213 ( .A1(n11072), .A2(n11493), .Z(n14241) );
  CLKBUF_X2 U13215 ( .I(n25155), .Z(n10402) );
  BUF_X2 U13219 ( .I(n38702), .Z(n23199) );
  OAI21_X1 U13221 ( .A1(n36614), .A2(n60431), .B(n18672), .ZN(n18671) );
  AOI22_X1 U13222 ( .A1(n36112), .A2(n36114), .B1(n36111), .B2(n8765), .ZN(
        n8764) );
  NAND2_X1 U13233 ( .A1(n18207), .A2(n36710), .ZN(n36713) );
  NOR2_X1 U13244 ( .A1(n16353), .A2(n35942), .ZN(n8174) );
  NAND2_X1 U13246 ( .A1(n6123), .A2(n37189), .ZN(n6122) );
  AND2_X1 U13247 ( .A1(n19158), .A2(n24010), .Z(n22836) );
  NAND2_X1 U13250 ( .A1(n36872), .A2(n2918), .ZN(n8858) );
  OAI22_X1 U13254 ( .A1(n35607), .A2(n1766), .B1(n9087), .B2(n36201), .ZN(
        n9086) );
  NAND3_X1 U13257 ( .A1(n36826), .A2(n6984), .A3(n36831), .ZN(n11304) );
  AOI21_X1 U13258 ( .A1(n36263), .A2(n11054), .B(n8535), .ZN(n8534) );
  NAND2_X1 U13265 ( .A1(n36582), .A2(n1767), .ZN(n3651) );
  NAND2_X1 U13266 ( .A1(n3649), .A2(n3789), .ZN(n3648) );
  NOR2_X1 U13271 ( .A1(n23146), .A2(n61747), .ZN(n6807) );
  NOR2_X1 U13272 ( .A1(n37339), .A2(n37327), .ZN(n37331) );
  NOR2_X1 U13275 ( .A1(n35984), .A2(n19354), .ZN(n10965) );
  INV_X1 U13276 ( .I(n35147), .ZN(n19948) );
  AOI21_X1 U13278 ( .A1(n20147), .A2(n36698), .B(n35350), .ZN(n34202) );
  AND3_X1 U13283 ( .A1(n35509), .A2(n35508), .A3(n11778), .Z(n11777) );
  NOR2_X1 U13284 ( .A1(n11832), .A2(n23601), .ZN(n10115) );
  INV_X1 U13291 ( .I(n36866), .ZN(n37391) );
  NAND2_X1 U13293 ( .A1(n58743), .A2(n21467), .ZN(n9087) );
  AOI22_X1 U13300 ( .A1(n25343), .A2(n37028), .B1(n22524), .B2(n37029), .ZN(
        n25342) );
  NOR2_X1 U13302 ( .A1(n37333), .A2(n37326), .ZN(n37005) );
  NAND2_X1 U13303 ( .A1(n36848), .A2(n63697), .ZN(n4853) );
  NAND2_X1 U13304 ( .A1(n35181), .A2(n25584), .ZN(n35606) );
  NAND2_X1 U13310 ( .A1(n34874), .A2(n34875), .ZN(n19816) );
  AND2_X1 U13311 ( .A1(n1790), .A2(n64087), .Z(n16263) );
  NOR2_X1 U13314 ( .A1(n61831), .A2(n23778), .ZN(n35105) );
  INV_X1 U13317 ( .I(n16885), .ZN(n10765) );
  OAI22_X1 U13328 ( .A1(n36486), .A2(n36485), .B1(n1782), .B2(n8363), .ZN(
        n36491) );
  NOR3_X1 U13331 ( .A1(n37340), .A2(n37329), .A3(n62734), .ZN(n37330) );
  OAI22_X1 U13333 ( .A1(n36302), .A2(n36303), .B1(n12393), .B2(n36301), .ZN(
        n36317) );
  NAND2_X1 U13334 ( .A1(n61770), .A2(n11028), .ZN(n7254) );
  NOR2_X1 U13335 ( .A1(n8608), .A2(n35353), .ZN(n9932) );
  NAND2_X1 U13337 ( .A1(n10127), .A2(n9041), .ZN(n8085) );
  NAND3_X1 U13341 ( .A1(n34844), .A2(n34845), .A3(n34843), .ZN(n37489) );
  AND2_X1 U13342 ( .A1(n5185), .A2(n63643), .Z(n14172) );
  NAND2_X1 U13344 ( .A1(n36428), .A2(n33789), .ZN(n36432) );
  NOR3_X1 U13345 ( .A1(n35966), .A2(n15432), .A3(n6606), .ZN(n35547) );
  NAND2_X1 U13346 ( .A1(n15038), .A2(n36442), .ZN(n15036) );
  AOI22_X1 U13348 ( .A1(n36869), .A2(n37390), .B1(n60507), .B2(n1413), .ZN(
        n8861) );
  NAND2_X1 U13354 ( .A1(n35966), .A2(n35965), .ZN(n35967) );
  NAND2_X1 U13356 ( .A1(n36451), .A2(n15034), .ZN(n35589) );
  NAND2_X1 U13358 ( .A1(n36920), .A2(n1414), .ZN(n23452) );
  INV_X1 U13359 ( .I(n35426), .ZN(n23944) );
  NOR2_X1 U13361 ( .A1(n798), .A2(n2362), .ZN(n2094) );
  NOR2_X1 U13362 ( .A1(n36378), .A2(n1785), .ZN(n36381) );
  NAND3_X1 U13363 ( .A1(n36130), .A2(n36305), .A3(n36796), .ZN(n36132) );
  INV_X1 U13371 ( .I(n36835), .ZN(n1771) );
  NAND2_X1 U13374 ( .A1(n36939), .A2(n59842), .ZN(n36942) );
  AOI21_X1 U13375 ( .A1(n36938), .A2(n36937), .B(n14629), .ZN(n6167) );
  NAND2_X1 U13380 ( .A1(n35423), .A2(n36743), .ZN(n25154) );
  AND2_X1 U13381 ( .A1(n36852), .A2(n7092), .Z(n16127) );
  OR2_X1 U13383 ( .A1(n10753), .A2(n1777), .Z(n11837) );
  NOR2_X1 U13385 ( .A1(n34863), .A2(n37030), .ZN(n35489) );
  NAND3_X1 U13386 ( .A1(n20020), .A2(n36926), .A3(n36920), .ZN(n34929) );
  AND3_X1 U13387 ( .A1(n34860), .A2(n21010), .A3(n34859), .Z(n34861) );
  NAND3_X1 U13388 ( .A1(n36463), .A2(n36584), .A3(n11272), .ZN(n11273) );
  AND2_X1 U13390 ( .A1(n37945), .A2(n37090), .Z(n22935) );
  NAND2_X1 U13393 ( .A1(n36803), .A2(n57211), .ZN(n34577) );
  NOR2_X1 U13394 ( .A1(n5483), .A2(n63643), .ZN(n12653) );
  INV_X1 U13403 ( .I(n35423), .ZN(n35066) );
  INV_X1 U13405 ( .I(n22295), .ZN(n36430) );
  AOI21_X1 U13407 ( .A1(n36889), .A2(n1421), .B(n36944), .ZN(n34910) );
  NAND2_X1 U13409 ( .A1(n35910), .A2(n21010), .ZN(n3589) );
  BUF_X4 U13410 ( .I(n18348), .Z(n1782) );
  NAND2_X1 U13411 ( .A1(n7028), .A2(n20060), .ZN(n12899) );
  OAI21_X1 U13412 ( .A1(n8356), .A2(n11721), .B(n24102), .ZN(n11720) );
  NOR2_X1 U13413 ( .A1(n36226), .A2(n23257), .ZN(n15009) );
  OR2_X1 U13420 ( .A1(n8474), .A2(n1787), .Z(n35387) );
  BUF_X4 U13427 ( .I(n22254), .Z(n7933) );
  BUF_X4 U13434 ( .I(n37397), .Z(n6540) );
  NAND3_X1 U13441 ( .A1(n36554), .A2(n36553), .A3(n36574), .ZN(n7821) );
  NAND2_X1 U13446 ( .A1(n17892), .A2(n3233), .ZN(n13210) );
  INV_X2 U13449 ( .I(n12110), .ZN(n19539) );
  NOR2_X1 U13452 ( .A1(n8141), .A2(n3551), .ZN(n3550) );
  AOI22_X1 U13453 ( .A1(n32464), .A2(n33621), .B1(n32463), .B2(n32462), .ZN(
        n32465) );
  NAND3_X1 U13465 ( .A1(n35291), .A2(n35290), .A3(n35289), .ZN(n35292) );
  NAND2_X1 U13466 ( .A1(n25100), .A2(n35686), .ZN(n15294) );
  NAND2_X1 U13470 ( .A1(n31514), .A2(n33963), .ZN(n31541) );
  NAND2_X1 U13472 ( .A1(n33430), .A2(n64499), .ZN(n21475) );
  AOI21_X1 U13473 ( .A1(n33571), .A2(n19095), .B(n15614), .ZN(n15613) );
  NAND3_X1 U13477 ( .A1(n33350), .A2(n33349), .A3(n14011), .ZN(n33351) );
  NOR2_X1 U13480 ( .A1(n20325), .A2(n18568), .ZN(n16799) );
  AOI21_X1 U13482 ( .A1(n33404), .A2(n3524), .B(n8142), .ZN(n8141) );
  AOI22_X1 U13483 ( .A1(n33565), .A2(n33564), .B1(n16957), .B2(n33570), .ZN(
        n15612) );
  NAND2_X1 U13486 ( .A1(n11477), .A2(n2206), .ZN(n33430) );
  OAI21_X1 U13487 ( .A1(n64499), .A2(n20439), .B(n21474), .ZN(n21473) );
  AOI21_X1 U13488 ( .A1(n4643), .A2(n10267), .B(n33564), .ZN(n15614) );
  NAND3_X1 U13493 ( .A1(n31536), .A2(n14319), .A3(n31529), .ZN(n18932) );
  AOI21_X1 U13496 ( .A1(n2079), .A2(n34080), .B(n24737), .ZN(n25196) );
  AOI21_X1 U13498 ( .A1(n11433), .A2(n34589), .B(n34595), .ZN(n9812) );
  NAND2_X1 U13500 ( .A1(n35279), .A2(n35802), .ZN(n35281) );
  NAND2_X1 U13503 ( .A1(n9126), .A2(n5477), .ZN(n9125) );
  NAND2_X1 U13506 ( .A1(n11024), .A2(n33348), .ZN(n14011) );
  NOR2_X1 U13508 ( .A1(n18788), .A2(n3487), .ZN(n35824) );
  NAND3_X1 U13513 ( .A1(n17341), .A2(n17342), .A3(n12877), .ZN(n32836) );
  NAND2_X1 U13515 ( .A1(n4879), .A2(n9085), .ZN(n18089) );
  NAND3_X1 U13517 ( .A1(n19570), .A2(n34423), .A3(n35769), .ZN(n5583) );
  OR2_X1 U13520 ( .A1(n1795), .A2(n5410), .Z(n16145) );
  OAI21_X1 U13521 ( .A1(n34333), .A2(n64984), .B(n5874), .ZN(n13851) );
  AND3_X1 U13522 ( .A1(n33987), .A2(n5389), .A3(n11064), .Z(n5388) );
  NAND2_X1 U13529 ( .A1(n12412), .A2(n34155), .ZN(n32842) );
  NAND2_X1 U13534 ( .A1(n13470), .A2(n19457), .ZN(n13469) );
  OAI21_X1 U13536 ( .A1(n34118), .A2(n31727), .B(n59769), .ZN(n31730) );
  NAND2_X1 U13541 ( .A1(n35023), .A2(n11477), .ZN(n16579) );
  INV_X1 U13542 ( .I(n8009), .ZN(n33924) );
  INV_X1 U13543 ( .I(n33960), .ZN(n34079) );
  INV_X1 U13544 ( .I(n64407), .ZN(n21181) );
  NAND2_X1 U13547 ( .A1(n34497), .A2(n5519), .ZN(n5518) );
  NOR3_X1 U13550 ( .A1(n14980), .A2(n33944), .A3(n59769), .ZN(n32865) );
  INV_X1 U13551 ( .I(n2899), .ZN(n2908) );
  AOI21_X1 U13552 ( .A1(n33576), .A2(n33820), .B(n12506), .ZN(n33578) );
  NOR2_X1 U13553 ( .A1(n20835), .A2(n34595), .ZN(n5159) );
  NAND2_X1 U13555 ( .A1(n34196), .A2(n34201), .ZN(n2401) );
  NAND2_X1 U13561 ( .A1(n11709), .A2(n1425), .ZN(n21813) );
  OAI21_X1 U13562 ( .A1(n34601), .A2(n20946), .B(n1798), .ZN(n19603) );
  AND4_X1 U13563 ( .A1(n34134), .A2(n34142), .A3(n33654), .A4(n19416), .Z(
        n31718) );
  NAND3_X1 U13565 ( .A1(n32426), .A2(n32427), .A3(n34731), .ZN(n21455) );
  NAND3_X1 U13571 ( .A1(n34523), .A2(n34051), .A3(n64358), .ZN(n34052) );
  NAND2_X1 U13573 ( .A1(n3174), .A2(n3173), .ZN(n35686) );
  NAND2_X1 U13575 ( .A1(n35778), .A2(n35775), .ZN(n35787) );
  NAND2_X1 U13578 ( .A1(n34186), .A2(n63116), .ZN(n10852) );
  NOR2_X1 U13579 ( .A1(n35280), .A2(n11186), .ZN(n21764) );
  OAI21_X1 U13583 ( .A1(n35646), .A2(n35645), .B(n35650), .ZN(n3442) );
  NOR2_X1 U13586 ( .A1(n25509), .A2(n33004), .ZN(n32452) );
  NAND3_X1 U13589 ( .A1(n33614), .A2(n3549), .A3(n33613), .ZN(n33615) );
  NAND3_X1 U13590 ( .A1(n34795), .A2(n33468), .A3(n14112), .ZN(n15573) );
  NAND3_X1 U13592 ( .A1(n445), .A2(n32684), .A3(n33542), .ZN(n32685) );
  NAND2_X1 U13594 ( .A1(n33397), .A2(n34128), .ZN(n33399) );
  OAI21_X1 U13598 ( .A1(n33963), .A2(n64603), .B(n1810), .ZN(n6344) );
  NOR2_X1 U13601 ( .A1(n31767), .A2(n32891), .ZN(n21432) );
  NOR2_X1 U13604 ( .A1(n63375), .A2(n24614), .ZN(n4881) );
  AOI21_X1 U13605 ( .A1(n7342), .A2(n57546), .B(n35206), .ZN(n35208) );
  NAND2_X1 U13606 ( .A1(n33814), .A2(n16243), .ZN(n24496) );
  NAND2_X1 U13607 ( .A1(n18277), .A2(n32834), .ZN(n5732) );
  INV_X1 U13609 ( .I(n34669), .ZN(n34517) );
  AOI22_X1 U13610 ( .A1(n35287), .A2(n35705), .B1(n35750), .B2(n19265), .ZN(
        n35290) );
  AND2_X1 U13611 ( .A1(n34550), .A2(n34019), .Z(n11083) );
  NAND2_X1 U13612 ( .A1(n60604), .A2(n34725), .ZN(n16819) );
  AND2_X1 U13614 ( .A1(n34026), .A2(n1427), .Z(n9813) );
  AND2_X1 U13616 ( .A1(n18301), .A2(n34989), .Z(n34066) );
  NOR2_X1 U13620 ( .A1(n62683), .A2(n9030), .ZN(n9029) );
  NAND2_X1 U13621 ( .A1(n32945), .A2(n21388), .ZN(n34758) );
  NAND2_X1 U13623 ( .A1(n57166), .A2(n1345), .ZN(n33477) );
  OAI21_X1 U13626 ( .A1(n1424), .A2(n2322), .B(n18300), .ZN(n24875) );
  NAND2_X1 U13627 ( .A1(n33521), .A2(n20785), .ZN(n14046) );
  NOR2_X1 U13628 ( .A1(n8694), .A2(n18136), .ZN(n4700) );
  INV_X1 U13631 ( .I(n25617), .ZN(n33397) );
  INV_X1 U13638 ( .I(n33598), .ZN(n5357) );
  NAND2_X1 U13639 ( .A1(n60926), .A2(n8552), .ZN(n12404) );
  NAND2_X1 U13640 ( .A1(n33560), .A2(n59681), .ZN(n4643) );
  AOI22_X1 U13646 ( .A1(n33752), .A2(n32965), .B1(n20660), .B2(n33756), .ZN(
        n14535) );
  NOR2_X1 U13647 ( .A1(n33601), .A2(n12121), .ZN(n12120) );
  INV_X1 U13648 ( .I(n12413), .ZN(n34157) );
  NAND2_X1 U13649 ( .A1(n12338), .A2(n60054), .ZN(n12340) );
  NOR2_X1 U13652 ( .A1(n34069), .A2(n15085), .ZN(n2765) );
  INV_X1 U13656 ( .I(n34414), .ZN(n18835) );
  NAND2_X1 U13657 ( .A1(n61496), .A2(n34415), .ZN(n34417) );
  INV_X1 U13661 ( .I(n34989), .ZN(n34981) );
  NAND2_X1 U13663 ( .A1(n33775), .A2(n34784), .ZN(n11445) );
  INV_X1 U13665 ( .I(n33801), .ZN(n35658) );
  INV_X1 U13669 ( .I(n5123), .ZN(n35042) );
  OAI22_X1 U13671 ( .A1(n31358), .A2(n3467), .B1(n64358), .B2(n8304), .ZN(
        n30896) );
  INV_X1 U13672 ( .I(n33775), .ZN(n34776) );
  NAND2_X1 U13673 ( .A1(n35656), .A2(n60835), .ZN(n15330) );
  NAND2_X1 U13674 ( .A1(n34198), .A2(n33993), .ZN(n13141) );
  NOR2_X1 U13679 ( .A1(n4097), .A2(n34113), .ZN(n34115) );
  INV_X2 U13680 ( .I(n34427), .ZN(n35777) );
  NOR2_X1 U13690 ( .A1(n16301), .A2(n4496), .ZN(n4355) );
  NOR2_X1 U13692 ( .A1(n33432), .A2(n34589), .ZN(n11402) );
  BUF_X2 U13694 ( .I(n8051), .Z(n8049) );
  INV_X2 U13695 ( .I(n34726), .ZN(n1536) );
  BUF_X2 U13696 ( .I(n34136), .Z(n19416) );
  INV_X4 U13698 ( .I(n5412), .ZN(n34161) );
  NAND2_X1 U13700 ( .A1(n23812), .A2(n15318), .ZN(n10656) );
  NOR2_X1 U13703 ( .A1(n34725), .A2(n23914), .ZN(n9389) );
  NOR2_X1 U13709 ( .A1(n35247), .A2(n62995), .ZN(n15329) );
  NAND2_X1 U13711 ( .A1(n63773), .A2(n35241), .ZN(n35647) );
  CLKBUF_X2 U13713 ( .I(n32868), .Z(n19119) );
  NAND3_X1 U13715 ( .A1(n24286), .A2(n6979), .A3(n57986), .ZN(n6982) );
  INV_X1 U13716 ( .I(n63421), .ZN(n1927) );
  CLKBUF_X2 U13720 ( .I(n1817), .Z(n10566) );
  OR2_X2 U13723 ( .A1(n25659), .A2(n30944), .Z(n33509) );
  INV_X4 U13724 ( .I(n9524), .ZN(n1542) );
  BUF_X2 U13725 ( .I(n33893), .Z(n35283) );
  BUF_X4 U13728 ( .I(n32262), .Z(n1545) );
  INV_X4 U13729 ( .I(n23689), .ZN(n1546) );
  BUF_X2 U13731 ( .I(n35001), .Z(n14111) );
  INV_X1 U13732 ( .I(n22744), .ZN(n24794) );
  INV_X1 U13734 ( .I(n32230), .ZN(n5089) );
  INV_X1 U13736 ( .I(n1819), .ZN(n6457) );
  CLKBUF_X2 U13741 ( .I(n21034), .Z(n8774) );
  INV_X1 U13748 ( .I(n20573), .ZN(n19057) );
  BUF_X2 U13753 ( .I(n30848), .Z(n33164) );
  INV_X1 U13754 ( .I(n33857), .ZN(n3070) );
  NAND2_X1 U13755 ( .A1(n25553), .A2(n3297), .ZN(n3296) );
  INV_X1 U13757 ( .I(n3523), .ZN(n11232) );
  INV_X1 U13759 ( .I(n21128), .ZN(n33896) );
  NOR2_X1 U13763 ( .A1(n3298), .A2(n1899), .ZN(n3297) );
  INV_X1 U13764 ( .I(n24868), .ZN(n5876) );
  BUF_X2 U13765 ( .I(n14565), .Z(n14563) );
  INV_X1 U13766 ( .I(n31943), .ZN(n32655) );
  INV_X1 U13767 ( .I(n14565), .ZN(n6445) );
  BUF_X2 U13768 ( .I(n18547), .Z(n15102) );
  NAND2_X1 U13770 ( .A1(n18765), .A2(n18761), .ZN(n26652) );
  BUF_X4 U13772 ( .I(n30894), .Z(n15725) );
  NOR2_X1 U13774 ( .A1(n25553), .A2(n55150), .ZN(n3301) );
  NAND2_X2 U13777 ( .A1(n22126), .A2(n26372), .ZN(n32483) );
  NOR2_X1 U13780 ( .A1(n14701), .A2(n7981), .ZN(n29465) );
  INV_X1 U13781 ( .I(n3607), .ZN(n6231) );
  AOI21_X1 U13786 ( .A1(n2873), .A2(n4062), .B(n14452), .ZN(n2872) );
  NAND2_X1 U13789 ( .A1(n3816), .A2(n3815), .ZN(n3811) );
  NOR2_X1 U13791 ( .A1(n28985), .A2(n25898), .ZN(n5494) );
  AOI21_X1 U13792 ( .A1(n21659), .A2(n30023), .B(n29725), .ZN(n5425) );
  NOR2_X1 U13795 ( .A1(n30232), .A2(n14336), .ZN(n30235) );
  OAI21_X1 U13798 ( .A1(n13691), .A2(n17413), .B(n12979), .ZN(n13690) );
  NAND2_X1 U13805 ( .A1(n6038), .A2(n30676), .ZN(n18236) );
  AOI22_X1 U13809 ( .A1(n21604), .A2(n11425), .B1(n28706), .B2(n30456), .ZN(
        n6229) );
  NAND3_X1 U13810 ( .A1(n2267), .A2(n30055), .A3(n11656), .ZN(n2282) );
  NAND2_X1 U13812 ( .A1(n30388), .A2(n30387), .ZN(n19515) );
  NAND2_X1 U13815 ( .A1(n5100), .A2(n61162), .ZN(n23679) );
  NAND2_X1 U13816 ( .A1(n5910), .A2(n9891), .ZN(n9890) );
  NAND2_X1 U13818 ( .A1(n30442), .A2(n29983), .ZN(n3815) );
  NAND2_X1 U13821 ( .A1(n3180), .A2(n28704), .ZN(n6179) );
  NOR2_X1 U13822 ( .A1(n27072), .A2(n30028), .ZN(n27738) );
  NAND2_X1 U13824 ( .A1(n4084), .A2(n4083), .ZN(n4082) );
  AOI22_X1 U13826 ( .A1(n20188), .A2(n20187), .B1(n30587), .B2(n59810), .ZN(
        n20186) );
  NOR2_X1 U13829 ( .A1(n4037), .A2(n29511), .ZN(n14452) );
  NAND2_X1 U13830 ( .A1(n28098), .A2(n29449), .ZN(n28102) );
  OAI21_X1 U13832 ( .A1(n30549), .A2(n1839), .B(n30548), .ZN(n6817) );
  NOR2_X1 U13837 ( .A1(n29453), .A2(n28736), .ZN(n28995) );
  NAND2_X1 U13839 ( .A1(n4442), .A2(n24949), .ZN(n5984) );
  INV_X1 U13842 ( .I(n29957), .ZN(n30790) );
  NAND2_X1 U13843 ( .A1(n3993), .A2(n30392), .ZN(n6180) );
  AND2_X1 U13844 ( .A1(n31220), .A2(n1278), .Z(n31222) );
  NAND2_X1 U13846 ( .A1(n22164), .A2(n23370), .ZN(n8335) );
  OAI21_X1 U13847 ( .A1(n1868), .A2(n10427), .B(n10426), .ZN(n30576) );
  NAND2_X1 U13848 ( .A1(n1843), .A2(n30588), .ZN(n24913) );
  INV_X1 U13849 ( .I(n30586), .ZN(n30587) );
  OAI22_X1 U13850 ( .A1(n14641), .A2(n18880), .B1(n30745), .B2(n30740), .ZN(
        n7037) );
  NOR2_X1 U13851 ( .A1(n28925), .A2(n28924), .ZN(n9689) );
  OR3_X1 U13857 ( .A1(n1849), .A2(n29787), .A3(n28943), .Z(n7450) );
  NAND2_X1 U13858 ( .A1(n1844), .A2(n58765), .ZN(n3265) );
  NAND3_X1 U13859 ( .A1(n31102), .A2(n31114), .A3(n1856), .ZN(n10731) );
  NOR2_X1 U13861 ( .A1(n31246), .A2(n11378), .ZN(n31249) );
  NAND2_X1 U13862 ( .A1(n30260), .A2(n30048), .ZN(n2285) );
  OAI21_X1 U13863 ( .A1(n28583), .A2(n31086), .B(n5760), .ZN(n28585) );
  NAND2_X1 U13865 ( .A1(n28422), .A2(n8218), .ZN(n8091) );
  NAND2_X1 U13867 ( .A1(n22627), .A2(n1843), .ZN(n4083) );
  NAND2_X1 U13868 ( .A1(n1861), .A2(n20606), .ZN(n4084) );
  NAND3_X1 U13869 ( .A1(n28778), .A2(n28777), .A3(n19461), .ZN(n28783) );
  NOR2_X1 U13870 ( .A1(n30335), .A2(n3898), .ZN(n3897) );
  NAND2_X1 U13872 ( .A1(n3993), .A2(n11106), .ZN(n2873) );
  OAI21_X1 U13878 ( .A1(n25182), .A2(n13844), .B(n23349), .ZN(n13843) );
  NAND4_X1 U13879 ( .A1(n30750), .A2(n1875), .A3(n23799), .A4(n19929), .ZN(
        n30016) );
  OAI21_X1 U13884 ( .A1(n29451), .A2(n29460), .B(n14868), .ZN(n23176) );
  NAND2_X1 U13887 ( .A1(n3486), .A2(n30885), .ZN(n29400) );
  OR2_X1 U13889 ( .A1(n29793), .A2(n30085), .Z(n3243) );
  OAI21_X1 U13892 ( .A1(n10925), .A2(n31217), .B(n30669), .ZN(n10924) );
  AOI21_X1 U13893 ( .A1(n30386), .A2(n31114), .B(n30385), .ZN(n30388) );
  NAND2_X1 U13896 ( .A1(n20918), .A2(n1858), .ZN(n22837) );
  NOR2_X1 U13897 ( .A1(n29798), .A2(n9197), .ZN(n7737) );
  NOR2_X1 U13898 ( .A1(n12300), .A2(n29538), .ZN(n5865) );
  NOR2_X1 U13899 ( .A1(n16961), .A2(n29992), .ZN(n6795) );
  NOR2_X1 U13900 ( .A1(n30391), .A2(n30392), .ZN(n2796) );
  INV_X1 U13902 ( .I(n29882), .ZN(n29881) );
  NAND2_X1 U13905 ( .A1(n30480), .A2(n25848), .ZN(n11988) );
  NAND2_X1 U13909 ( .A1(n1317), .A2(n11205), .ZN(n11204) );
  NOR2_X1 U13912 ( .A1(n31041), .A2(n30108), .ZN(n30151) );
  INV_X1 U13913 ( .I(n29798), .ZN(n21062) );
  AOI21_X1 U13914 ( .A1(n8336), .A2(n27915), .B(n23370), .ZN(n9287) );
  NOR2_X1 U13915 ( .A1(n64565), .A2(n64940), .ZN(n29522) );
  NOR2_X1 U13916 ( .A1(n29739), .A2(n22796), .ZN(n30093) );
  AND2_X1 U13918 ( .A1(n29490), .A2(n10427), .Z(n15774) );
  OAI21_X1 U13919 ( .A1(n9250), .A2(n58237), .B(n29248), .ZN(n28940) );
  AOI21_X1 U13920 ( .A1(n29248), .A2(n7943), .B(n28937), .ZN(n28941) );
  OAI21_X1 U13923 ( .A1(n1351), .A2(n60214), .B(n22873), .ZN(n8961) );
  AND2_X1 U13924 ( .A1(n30840), .A2(n30223), .Z(n17856) );
  NAND2_X1 U13925 ( .A1(n21876), .A2(n16223), .ZN(n30094) );
  NAND2_X1 U13927 ( .A1(n30352), .A2(n30618), .ZN(n28563) );
  NOR2_X1 U13929 ( .A1(n29001), .A2(n63417), .ZN(n14701) );
  NAND2_X1 U13930 ( .A1(n1868), .A2(n57437), .ZN(n10426) );
  NOR2_X1 U13934 ( .A1(n27900), .A2(n29905), .ZN(n31184) );
  NAND2_X1 U13935 ( .A1(n29457), .A2(n29452), .ZN(n8802) );
  NOR2_X1 U13936 ( .A1(n27789), .A2(n9475), .ZN(n7947) );
  NOR2_X1 U13937 ( .A1(n28762), .A2(n7943), .ZN(n14602) );
  INV_X1 U13939 ( .I(n6615), .ZN(n8946) );
  AND3_X1 U13941 ( .A1(n31161), .A2(n31269), .A3(n22934), .Z(n31162) );
  NAND2_X1 U13942 ( .A1(n20179), .A2(n24206), .ZN(n30779) );
  NAND2_X1 U13943 ( .A1(n31246), .A2(n1435), .ZN(n29890) );
  NAND2_X1 U13945 ( .A1(n6349), .A2(n1315), .ZN(n3989) );
  NAND2_X1 U13949 ( .A1(n30778), .A2(n29959), .ZN(n30785) );
  NAND2_X1 U13952 ( .A1(n28584), .A2(n5267), .ZN(n24502) );
  NAND2_X1 U13953 ( .A1(n29820), .A2(n29993), .ZN(n3723) );
  NAND2_X1 U13955 ( .A1(n30415), .A2(n3085), .ZN(n8642) );
  AOI21_X1 U13956 ( .A1(n10345), .A2(n24896), .B(n29824), .ZN(n4100) );
  AOI21_X1 U13960 ( .A1(n30585), .A2(n22627), .B(n18810), .ZN(n20188) );
  NAND2_X1 U13961 ( .A1(n29458), .A2(n1867), .ZN(n5909) );
  NAND3_X1 U13962 ( .A1(n30214), .A2(n22596), .A3(n16920), .ZN(n8998) );
  OAI21_X1 U13964 ( .A1(n17412), .A2(n64940), .B(n64565), .ZN(n29519) );
  NOR2_X1 U13966 ( .A1(n1432), .A2(n31208), .ZN(n25513) );
  NAND2_X1 U13967 ( .A1(n58644), .A2(n31208), .ZN(n6428) );
  INV_X1 U13968 ( .I(n63417), .ZN(n28098) );
  AND2_X1 U13969 ( .A1(n30271), .A2(n29220), .Z(n28774) );
  NAND2_X1 U13971 ( .A1(n17872), .A2(n58999), .ZN(n9785) );
  NAND2_X1 U13973 ( .A1(n30002), .A2(n22745), .ZN(n28679) );
  AOI21_X1 U13974 ( .A1(n30736), .A2(n31208), .B(n20172), .ZN(n30737) );
  CLKBUF_X2 U13975 ( .I(n1865), .Z(n4444) );
  OR2_X1 U13976 ( .A1(n13280), .A2(n24564), .Z(n30744) );
  NOR2_X1 U13979 ( .A1(n30396), .A2(n22742), .ZN(n6586) );
  NOR2_X1 U13980 ( .A1(n9250), .A2(n7943), .ZN(n7946) );
  NAND2_X1 U13981 ( .A1(n18736), .A2(n17414), .ZN(n13517) );
  CLKBUF_X2 U13984 ( .I(n1862), .Z(n19218) );
  AND2_X1 U13985 ( .A1(n2351), .A2(n30195), .Z(n16223) );
  BUF_X4 U13991 ( .I(n29209), .Z(n19461) );
  CLKBUF_X2 U13997 ( .I(n24335), .Z(n18472) );
  INV_X1 U13999 ( .I(n29846), .ZN(n1867) );
  NAND2_X1 U14002 ( .A1(n5932), .A2(n24263), .ZN(n5931) );
  NOR2_X1 U14004 ( .A1(n23008), .A2(n31254), .ZN(n30886) );
  NOR2_X1 U14005 ( .A1(n23224), .A2(n61421), .ZN(n7403) );
  BUF_X4 U14007 ( .I(n19363), .Z(n21532) );
  CLKBUF_X2 U14008 ( .I(n28080), .Z(n20988) );
  INV_X2 U14010 ( .I(n29432), .ZN(n27150) );
  BUF_X4 U14011 ( .I(n31276), .Z(n6316) );
  NAND2_X1 U14012 ( .A1(n24088), .A2(n24264), .ZN(n5932) );
  INV_X1 U14015 ( .I(n29244), .ZN(n13336) );
  OAI22_X1 U14016 ( .A1(n23419), .A2(n23779), .B1(n23418), .B2(n28271), .ZN(
        n18500) );
  AOI21_X1 U14027 ( .A1(n18914), .A2(n22643), .B(n11051), .ZN(n26473) );
  AOI21_X1 U14031 ( .A1(n26685), .A2(n28348), .B(n26684), .ZN(n26686) );
  AOI21_X1 U14046 ( .A1(n12641), .A2(n12639), .B(n29617), .ZN(n12638) );
  AOI21_X1 U14048 ( .A1(n7371), .A2(n7023), .B(n5468), .ZN(n5467) );
  AOI21_X1 U14049 ( .A1(n27839), .A2(n27841), .B(n27664), .ZN(n17603) );
  OAI21_X1 U14050 ( .A1(n8807), .A2(n28305), .B(n27173), .ZN(n9472) );
  NOR2_X1 U14061 ( .A1(n14533), .A2(n22991), .ZN(n10446) );
  OAI21_X1 U14065 ( .A1(n26540), .A2(n1895), .B(n10946), .ZN(n26300) );
  NOR2_X1 U14066 ( .A1(n11073), .A2(n11773), .ZN(n11759) );
  INV_X1 U14068 ( .I(n10419), .ZN(n7109) );
  OR2_X1 U14069 ( .A1(n27113), .A2(n10946), .Z(n17726) );
  OAI21_X1 U14070 ( .A1(n18534), .A2(n27973), .B(n27390), .ZN(n18533) );
  AOI21_X1 U14071 ( .A1(n11075), .A2(n14780), .B(n1877), .ZN(n7585) );
  NOR2_X1 U14073 ( .A1(n4718), .A2(n4717), .ZN(n12641) );
  AOI21_X1 U14074 ( .A1(n28419), .A2(n11226), .B(n7630), .ZN(n28420) );
  OAI22_X1 U14077 ( .A1(n27496), .A2(n27497), .B1(n59552), .B2(n29297), .ZN(
        n7917) );
  NAND3_X1 U14079 ( .A1(n27064), .A2(n27062), .A3(n27063), .ZN(n27069) );
  NAND2_X1 U14080 ( .A1(n264), .A2(n29609), .ZN(n14938) );
  NOR2_X1 U14084 ( .A1(n3428), .A2(n28650), .ZN(n13028) );
  OAI21_X1 U14088 ( .A1(n18848), .A2(n16515), .B(n26421), .ZN(n16516) );
  AOI21_X1 U14089 ( .A1(n27941), .A2(n1878), .B(n11605), .ZN(n11658) );
  OAI21_X1 U14091 ( .A1(n14134), .A2(n26531), .B(n22110), .ZN(n14133) );
  OR2_X1 U14092 ( .A1(n12422), .A2(n10946), .Z(n12421) );
  AOI21_X1 U14093 ( .A1(n28218), .A2(n3904), .B(n2112), .ZN(n2111) );
  NOR2_X1 U14095 ( .A1(n9468), .A2(n1879), .ZN(n9467) );
  OAI21_X1 U14098 ( .A1(n3200), .A2(n26796), .B(n26795), .ZN(n3199) );
  NAND2_X1 U14099 ( .A1(n522), .A2(n12109), .ZN(n26779) );
  NOR2_X1 U14101 ( .A1(n16793), .A2(n16255), .ZN(n16790) );
  AOI21_X1 U14105 ( .A1(n28029), .A2(n6222), .B(n15978), .ZN(n6822) );
  AOI21_X1 U14107 ( .A1(n27600), .A2(n27073), .B(n1879), .ZN(n12275) );
  AOI21_X1 U14108 ( .A1(n27935), .A2(n29172), .B(n1878), .ZN(n14256) );
  OAI21_X1 U14110 ( .A1(n17248), .A2(n17247), .B(n27934), .ZN(n5468) );
  AOI21_X1 U14112 ( .A1(n3749), .A2(n10598), .B(n29697), .ZN(n20098) );
  NAND2_X1 U14113 ( .A1(n26764), .A2(n64809), .ZN(n27247) );
  INV_X1 U14116 ( .I(n28339), .ZN(n27197) );
  OAI21_X1 U14119 ( .A1(n18200), .A2(n17489), .B(n29146), .ZN(n5471) );
  NAND3_X1 U14121 ( .A1(n29302), .A2(n10324), .A3(n1360), .ZN(n22629) );
  AOI21_X1 U14122 ( .A1(n1440), .A2(n26654), .B(n62784), .ZN(n12929) );
  NOR2_X1 U14124 ( .A1(n57872), .A2(n27022), .ZN(n28043) );
  NOR2_X1 U14125 ( .A1(n18224), .A2(n15650), .ZN(n21300) );
  AND3_X1 U14126 ( .A1(n28231), .A2(n61177), .A3(n9661), .Z(n15978) );
  NAND2_X1 U14127 ( .A1(n6345), .A2(n29643), .ZN(n6408) );
  NAND2_X1 U14128 ( .A1(n59935), .A2(n29642), .ZN(n19550) );
  OR2_X1 U14130 ( .A1(n26935), .A2(n27548), .Z(n16255) );
  NOR2_X1 U14131 ( .A1(n27962), .A2(n7452), .ZN(n10224) );
  AND2_X1 U14133 ( .A1(n16707), .A2(n1355), .Z(n2343) );
  NOR2_X1 U14134 ( .A1(n26794), .A2(n27877), .ZN(n3200) );
  AOI21_X1 U14135 ( .A1(n26804), .A2(n26805), .B(n27255), .ZN(n3202) );
  AOI22_X1 U14137 ( .A1(n22110), .A2(n26322), .B1(n15715), .B2(n28366), .ZN(
        n21042) );
  AND2_X1 U14139 ( .A1(n27179), .A2(n26640), .Z(n8807) );
  NOR2_X1 U14140 ( .A1(n13764), .A2(n29172), .ZN(n13762) );
  OAI21_X1 U14142 ( .A1(n3255), .A2(n28396), .B(n3254), .ZN(n3253) );
  OAI22_X1 U14143 ( .A1(n14227), .A2(n29169), .B1(n29168), .B2(n5306), .ZN(
        n15197) );
  OAI22_X1 U14144 ( .A1(n3332), .A2(n22159), .B1(n3331), .B2(n8202), .ZN(n3330) );
  NAND2_X1 U14145 ( .A1(n22397), .A2(n28397), .ZN(n28006) );
  NOR2_X1 U14147 ( .A1(n29146), .A2(n16654), .ZN(n3414) );
  INV_X1 U14149 ( .I(n27073), .ZN(n27601) );
  OAI22_X1 U14150 ( .A1(n8791), .A2(n28027), .B1(n61035), .B2(n28026), .ZN(
        n22220) );
  NAND3_X1 U14151 ( .A1(n27928), .A2(n27296), .A3(n17747), .ZN(n2661) );
  OR3_X1 U14153 ( .A1(n28342), .A2(n27206), .A3(n28346), .Z(n26595) );
  NAND2_X1 U14154 ( .A1(n26834), .A2(n7110), .ZN(n16515) );
  NAND2_X1 U14156 ( .A1(n29642), .A2(n29641), .ZN(n6603) );
  NAND2_X1 U14157 ( .A1(n29320), .A2(n29321), .ZN(n19963) );
  NAND3_X1 U14158 ( .A1(n29296), .A2(n27495), .A3(n5206), .ZN(n7916) );
  AOI21_X1 U14159 ( .A1(n13376), .A2(n13375), .B(n1885), .ZN(n13374) );
  NAND2_X1 U14162 ( .A1(n28418), .A2(n1891), .ZN(n3293) );
  AOI21_X1 U14164 ( .A1(n28460), .A2(n13007), .B(n28617), .ZN(n13006) );
  INV_X1 U14165 ( .I(n28646), .ZN(n18825) );
  AOI21_X1 U14166 ( .A1(n7220), .A2(n28411), .B(n180), .ZN(n28412) );
  NOR2_X1 U14167 ( .A1(n11052), .A2(n26599), .ZN(n10574) );
  OAI22_X1 U14168 ( .A1(n15763), .A2(n1883), .B1(n27249), .B2(n1443), .ZN(
        n2919) );
  NOR2_X1 U14169 ( .A1(n17619), .A2(n6759), .ZN(n17881) );
  OAI21_X1 U14170 ( .A1(n27807), .A2(n29709), .B(n28623), .ZN(n18035) );
  NOR2_X1 U14172 ( .A1(n13764), .A2(n64012), .ZN(n4821) );
  OAI22_X1 U14175 ( .A1(n28847), .A2(n6515), .B1(n6514), .B2(n6345), .ZN(
        n26854) );
  INV_X1 U14177 ( .I(n11073), .ZN(n27163) );
  AND2_X1 U14178 ( .A1(n20629), .A2(n28622), .Z(n20628) );
  NAND2_X1 U14179 ( .A1(n12072), .A2(n62005), .ZN(n29164) );
  OR3_X1 U14181 ( .A1(n20508), .A2(n27537), .A3(n23474), .Z(n27475) );
  AND2_X1 U14183 ( .A1(n20240), .A2(n10728), .Z(n20214) );
  NAND2_X1 U14184 ( .A1(n26610), .A2(n26540), .ZN(n28359) );
  INV_X1 U14186 ( .I(n22110), .ZN(n15651) );
  AOI22_X1 U14188 ( .A1(n3384), .A2(n28270), .B1(n64374), .B2(n28275), .ZN(
        n8791) );
  NAND3_X1 U14191 ( .A1(n28036), .A2(n10537), .A3(n60355), .ZN(n26571) );
  NAND2_X1 U14193 ( .A1(n1893), .A2(n3117), .ZN(n3332) );
  AND2_X1 U14194 ( .A1(n27849), .A2(n8948), .Z(n8888) );
  NAND2_X1 U14195 ( .A1(n1279), .A2(n22110), .ZN(n21184) );
  INV_X1 U14199 ( .I(n28174), .ZN(n29600) );
  AOI21_X1 U14200 ( .A1(n18931), .A2(n1894), .B(n27526), .ZN(n27207) );
  AND3_X1 U14201 ( .A1(n15477), .A2(n18751), .A3(n1230), .Z(n15534) );
  NAND2_X1 U14203 ( .A1(n27056), .A2(n26577), .ZN(n28232) );
  NAND2_X1 U14204 ( .A1(n23170), .A2(n3865), .ZN(n27373) );
  AND2_X1 U14205 ( .A1(n15477), .A2(n2705), .Z(n2704) );
  AOI21_X1 U14207 ( .A1(n28281), .A2(n60993), .B(n28280), .ZN(n28282) );
  NAND2_X1 U14209 ( .A1(n27174), .A2(n60818), .ZN(n27597) );
  AND2_X1 U14210 ( .A1(n17489), .A2(n6913), .Z(n26718) );
  AOI22_X1 U14211 ( .A1(n7477), .A2(n26660), .B1(n4324), .B2(n26618), .ZN(
        n26620) );
  INV_X2 U14212 ( .I(n8948), .ZN(n27853) );
  OAI22_X1 U14213 ( .A1(n20034), .A2(n29287), .B1(n29285), .B2(n29286), .ZN(
        n29288) );
  NAND2_X1 U14214 ( .A1(n8948), .A2(n7110), .ZN(n24441) );
  INV_X1 U14215 ( .I(n27849), .ZN(n27716) );
  NOR2_X1 U14216 ( .A1(n7499), .A2(n29153), .ZN(n27391) );
  NOR2_X1 U14217 ( .A1(n29141), .A2(n7371), .ZN(n3412) );
  NOR2_X1 U14218 ( .A1(n27136), .A2(n27135), .ZN(n11637) );
  NAND2_X1 U14221 ( .A1(n28543), .A2(n7354), .ZN(n26804) );
  AND2_X1 U14224 ( .A1(n22482), .A2(n24373), .Z(n3825) );
  NOR2_X1 U14225 ( .A1(n1322), .A2(n28221), .ZN(n3865) );
  NAND2_X1 U14226 ( .A1(n28804), .A2(n19423), .ZN(n6775) );
  BUF_X4 U14227 ( .I(n4848), .Z(n1970) );
  NAND2_X1 U14232 ( .A1(n2902), .A2(n26344), .ZN(n16266) );
  INV_X1 U14233 ( .I(n27179), .ZN(n27606) );
  INV_X1 U14236 ( .I(n28381), .ZN(n13702) );
  INV_X1 U14238 ( .I(n23805), .ZN(n10728) );
  INV_X2 U14239 ( .I(n24233), .ZN(n10324) );
  INV_X1 U14240 ( .I(n27543), .ZN(n27464) );
  CLKBUF_X2 U14241 ( .I(n1321), .Z(n17909) );
  INV_X1 U14244 ( .I(n62663), .ZN(n3384) );
  INV_X1 U14246 ( .I(n29145), .ZN(n2657) );
  AOI21_X1 U14247 ( .A1(n29618), .A2(n29617), .B(n29616), .ZN(n14937) );
  NAND2_X1 U14249 ( .A1(n23166), .A2(n1322), .ZN(n5430) );
  INV_X2 U14250 ( .I(n29127), .ZN(n1565) );
  NAND2_X1 U14254 ( .A1(n27056), .A2(n28036), .ZN(n28233) );
  BUF_X2 U14256 ( .I(n29636), .Z(n23386) );
  CLKBUF_X2 U14260 ( .I(n15758), .Z(n22952) );
  CLKBUF_X2 U14266 ( .I(n25785), .Z(n27232) );
  INV_X1 U14271 ( .I(n28674), .ZN(n29618) );
  INV_X2 U14272 ( .I(n29603), .ZN(n1567) );
  CLKBUF_X2 U14276 ( .I(n27494), .Z(n7538) );
  INV_X1 U14281 ( .I(n56065), .ZN(n1897) );
  BUF_X2 U14284 ( .I(n26275), .Z(n27051) );
  BUF_X2 U14286 ( .I(n27279), .Z(n23555) );
  BUF_X2 U14287 ( .I(n26407), .Z(n27283) );
  BUF_X2 U14289 ( .I(n26279), .Z(n26558) );
  CLKBUF_X2 U14290 ( .I(n27185), .Z(n23383) );
  BUF_X4 U14292 ( .I(n21959), .Z(n23942) );
  INV_X1 U14293 ( .I(n55150), .ZN(n1899) );
  CLKBUF_X2 U14300 ( .I(Key[163]), .Z(n56683) );
  CLKBUF_X2 U14301 ( .I(Key[190]), .Z(n57142) );
  CLKBUF_X2 U14302 ( .I(Key[101]), .Z(n23999) );
  CLKBUF_X4 U14303 ( .I(Key[124]), .Z(n55638) );
  CLKBUF_X4 U14310 ( .I(Key[172]), .Z(n24109) );
  CLKBUF_X2 U14312 ( .I(Key[36]), .Z(n53713) );
  CLKBUF_X4 U14313 ( .I(Key[8]), .Z(n53138) );
  CLKBUF_X2 U14314 ( .I(Key[38]), .Z(n50831) );
  CLKBUF_X4 U14318 ( .I(Key[158]), .Z(n56475) );
  CLKBUF_X2 U14319 ( .I(Key[24]), .Z(n23926) );
  NAND2_X1 U14320 ( .A1(n9402), .A2(n9403), .ZN(n9401) );
  NAND2_X1 U14323 ( .A1(n14842), .A2(n14840), .ZN(n14839) );
  NAND3_X1 U14328 ( .A1(n54263), .A2(n54262), .A3(n22641), .ZN(n22640) );
  NAND2_X1 U14329 ( .A1(n17641), .A2(n17640), .ZN(n17639) );
  NAND3_X1 U14332 ( .A1(n21744), .A2(n21750), .A3(n19153), .ZN(n19152) );
  AND2_X1 U14333 ( .A1(n15361), .A2(n53374), .Z(n19836) );
  NOR2_X1 U14334 ( .A1(n21748), .A2(n21745), .ZN(n21744) );
  INV_X1 U14335 ( .I(n53251), .ZN(n19671) );
  NAND4_X1 U14336 ( .A1(n55579), .A2(n55577), .A3(n55578), .A4(n8949), .ZN(
        n55581) );
  NAND3_X1 U14337 ( .A1(n17844), .A2(n17843), .A3(n17842), .ZN(n17841) );
  NAND2_X1 U14340 ( .A1(n12530), .A2(n12529), .ZN(n12528) );
  NAND2_X1 U14342 ( .A1(n12045), .A2(n1187), .ZN(n56294) );
  NAND3_X1 U14345 ( .A1(n9115), .A2(n56316), .A3(n9113), .ZN(n56317) );
  AOI21_X1 U14347 ( .A1(n23403), .A2(n2205), .B(n2204), .ZN(n2203) );
  INV_X1 U14349 ( .I(n53283), .ZN(n13238) );
  NOR2_X1 U14350 ( .A1(n2568), .A2(n5650), .ZN(n5647) );
  NOR2_X1 U14353 ( .A1(n11144), .A2(n12045), .ZN(n14383) );
  NAND2_X1 U14357 ( .A1(n60496), .A2(n53274), .ZN(n53286) );
  NAND2_X1 U14358 ( .A1(n53529), .A2(n53461), .ZN(n5965) );
  NAND3_X1 U14361 ( .A1(n56321), .A2(n11917), .A3(n11916), .ZN(n11915) );
  NAND2_X1 U14362 ( .A1(n15617), .A2(n56183), .ZN(n56201) );
  NAND2_X1 U14364 ( .A1(n54894), .A2(n54895), .ZN(n2204) );
  INV_X1 U14365 ( .I(n23594), .ZN(n5621) );
  NAND3_X1 U14366 ( .A1(n5553), .A2(n55604), .A3(n10381), .ZN(n6665) );
  NOR2_X1 U14367 ( .A1(n21847), .A2(n56823), .ZN(n17363) );
  NOR2_X1 U14370 ( .A1(n12532), .A2(n12526), .ZN(n12531) );
  INV_X1 U14371 ( .I(n56159), .ZN(n12530) );
  AOI21_X1 U14373 ( .A1(n52043), .A2(n21129), .B(n7054), .ZN(n17843) );
  AOI21_X1 U14375 ( .A1(n53810), .A2(n53794), .B(n21746), .ZN(n21745) );
  NAND2_X1 U14376 ( .A1(n2838), .A2(n2836), .ZN(n2832) );
  NAND2_X1 U14377 ( .A1(n19952), .A2(n19951), .ZN(n17842) );
  INV_X1 U14378 ( .I(n2619), .ZN(n2834) );
  NOR2_X1 U14379 ( .A1(n53818), .A2(n19154), .ZN(n19153) );
  NAND2_X1 U14380 ( .A1(n56852), .A2(n22365), .ZN(n22364) );
  OAI21_X1 U14381 ( .A1(n57114), .A2(n57115), .B(n18807), .ZN(n18806) );
  NAND2_X1 U14386 ( .A1(n8827), .A2(n56700), .ZN(n7462) );
  OAI21_X1 U14387 ( .A1(n1172), .A2(n63020), .B(n2865), .ZN(n54934) );
  OAI21_X1 U14388 ( .A1(n19578), .A2(n19577), .B(n518), .ZN(n6946) );
  NOR2_X1 U14390 ( .A1(n56701), .A2(n23785), .ZN(n7464) );
  NAND3_X1 U14393 ( .A1(n19033), .A2(n19032), .A3(n55836), .ZN(n19031) );
  OAI21_X1 U14397 ( .A1(n19036), .A2(n55852), .B(n55870), .ZN(n19035) );
  NAND2_X1 U14398 ( .A1(n9117), .A2(n1582), .ZN(n9116) );
  INV_X1 U14401 ( .I(n55630), .ZN(n10835) );
  NAND3_X1 U14402 ( .A1(n9560), .A2(n56699), .A3(n8618), .ZN(n8826) );
  NAND2_X1 U14404 ( .A1(n3370), .A2(n3369), .ZN(n55103) );
  NAND3_X1 U14405 ( .A1(n55142), .A2(n55141), .A3(n55168), .ZN(n7874) );
  OAI21_X1 U14406 ( .A1(n53471), .A2(n6032), .B(n53513), .ZN(n53472) );
  NAND2_X1 U14407 ( .A1(n10832), .A2(n52224), .ZN(n10081) );
  NOR2_X1 U14408 ( .A1(n55134), .A2(n7988), .ZN(n7987) );
  INV_X1 U14409 ( .I(n8618), .ZN(n8617) );
  NOR2_X1 U14410 ( .A1(n4989), .A2(n54421), .ZN(n23285) );
  INV_X1 U14411 ( .I(n9410), .ZN(n9114) );
  NAND2_X1 U14412 ( .A1(n54722), .A2(n4316), .ZN(n54725) );
  AND2_X1 U14413 ( .A1(n2240), .A2(n11346), .Z(n13237) );
  OAI22_X1 U14414 ( .A1(n21897), .A2(n1165), .B1(n55383), .B2(n22423), .ZN(
        n55331) );
  NAND3_X1 U14415 ( .A1(n20605), .A2(n20300), .A3(n25115), .ZN(n53744) );
  OAI21_X1 U14416 ( .A1(n15240), .A2(n56472), .B(n15239), .ZN(n13076) );
  AOI21_X1 U14418 ( .A1(n55596), .A2(n24297), .B(n55599), .ZN(n55600) );
  NAND3_X1 U14420 ( .A1(n53790), .A2(n53808), .A3(n53809), .ZN(n53773) );
  NAND2_X1 U14422 ( .A1(n20415), .A2(n20416), .ZN(n7054) );
  NOR2_X1 U14423 ( .A1(n4061), .A2(n12915), .ZN(n54013) );
  INV_X1 U14426 ( .I(n54209), .ZN(n54256) );
  NAND2_X1 U14427 ( .A1(n53264), .A2(n62996), .ZN(n53268) );
  NAND2_X1 U14428 ( .A1(n52650), .A2(n62699), .ZN(n52652) );
  INV_X1 U14429 ( .I(n53280), .ZN(n53255) );
  NAND2_X1 U14430 ( .A1(n56928), .A2(n56903), .ZN(n12398) );
  NAND4_X1 U14431 ( .A1(n11685), .A2(n4661), .A3(n55803), .A4(n55761), .ZN(
        n55762) );
  NAND3_X1 U14432 ( .A1(n53996), .A2(n53995), .A3(n54012), .ZN(n54004) );
  INV_X1 U14433 ( .I(n13492), .ZN(n4538) );
  NAND2_X1 U14434 ( .A1(n53996), .A2(n53995), .ZN(n53993) );
  NOR2_X1 U14436 ( .A1(n21121), .A2(n53926), .ZN(n21120) );
  NAND2_X1 U14438 ( .A1(n54387), .A2(n6560), .ZN(n5113) );
  INV_X1 U14441 ( .I(n53463), .ZN(n5964) );
  INV_X1 U14443 ( .I(n19076), .ZN(n11782) );
  INV_X1 U14445 ( .I(n21514), .ZN(n12395) );
  NOR2_X1 U14446 ( .A1(n56350), .A2(n18254), .ZN(n11921) );
  AND2_X1 U14447 ( .A1(n54866), .A2(n7680), .Z(n18740) );
  OAI22_X1 U14448 ( .A1(n53095), .A2(n23212), .B1(n53096), .B2(n12855), .ZN(
        n22912) );
  NAND2_X1 U14449 ( .A1(n12915), .A2(n53992), .ZN(n53937) );
  INV_X1 U14451 ( .I(n53966), .ZN(n53933) );
  NOR2_X1 U14452 ( .A1(n54202), .A2(n54201), .ZN(n13707) );
  INV_X1 U14453 ( .I(n7632), .ZN(n55210) );
  INV_X1 U14454 ( .I(n56814), .ZN(n13591) );
  NAND2_X1 U14457 ( .A1(n53927), .A2(n6168), .ZN(n4061) );
  INV_X1 U14460 ( .I(n56696), .ZN(n56700) );
  INV_X1 U14461 ( .I(n54388), .ZN(n6560) );
  AOI21_X1 U14462 ( .A1(n56192), .A2(n17408), .B(n56191), .ZN(n56197) );
  NOR2_X1 U14464 ( .A1(n54718), .A2(n23448), .ZN(n54668) );
  INV_X1 U14465 ( .I(n57144), .ZN(n4996) );
  INV_X1 U14466 ( .I(n55381), .ZN(n18135) );
  NOR2_X1 U14468 ( .A1(n2039), .A2(n2038), .ZN(n12212) );
  NOR2_X1 U14469 ( .A1(n54580), .A2(n14491), .ZN(n14490) );
  AOI21_X1 U14473 ( .A1(n55786), .A2(n21403), .B(n55829), .ZN(n10247) );
  NAND2_X1 U14474 ( .A1(n11684), .A2(n55760), .ZN(n4661) );
  INV_X1 U14475 ( .I(n3613), .ZN(n56297) );
  INV_X1 U14476 ( .I(n15765), .ZN(n4464) );
  AND2_X1 U14477 ( .A1(n19827), .A2(n61964), .Z(n16217) );
  AND2_X1 U14479 ( .A1(n56961), .A2(n56953), .Z(n14713) );
  NOR2_X1 U14480 ( .A1(n54388), .A2(n11276), .ZN(n54370) );
  NAND2_X1 U14482 ( .A1(n10310), .A2(n55145), .ZN(n7984) );
  NAND2_X1 U14483 ( .A1(n51879), .A2(n51878), .ZN(n17436) );
  NOR3_X1 U14485 ( .A1(n55119), .A2(n62699), .A3(n55168), .ZN(n52651) );
  AND3_X1 U14486 ( .A1(n54891), .A2(n54913), .A3(n22864), .Z(n23403) );
  OAI22_X1 U14487 ( .A1(n53675), .A2(n53695), .B1(n53658), .B2(n53694), .ZN(
        n53646) );
  INV_X1 U14488 ( .I(n56160), .ZN(n12529) );
  INV_X1 U14489 ( .I(n53644), .ZN(n2745) );
  NAND2_X1 U14490 ( .A1(n56192), .A2(n11274), .ZN(n12525) );
  OAI21_X1 U14491 ( .A1(n11325), .A2(n11324), .B(n1170), .ZN(n54371) );
  INV_X1 U14493 ( .I(n9338), .ZN(n9481) );
  NAND3_X1 U14494 ( .A1(n53305), .A2(n19735), .A3(n53294), .ZN(n9480) );
  OR3_X1 U14499 ( .A1(n55820), .A2(n55813), .A3(n55812), .Z(n55814) );
  OR2_X1 U14500 ( .A1(n53083), .A2(n52896), .Z(n52880) );
  INV_X1 U14501 ( .I(n8222), .ZN(n9112) );
  INV_X1 U14502 ( .I(n53160), .ZN(n12155) );
  NAND2_X1 U14504 ( .A1(n6511), .A2(n54877), .ZN(n2475) );
  NAND2_X1 U14505 ( .A1(n55780), .A2(n55820), .ZN(n4977) );
  INV_X1 U14507 ( .I(n15846), .ZN(n55236) );
  INV_X1 U14508 ( .I(n54541), .ZN(n19222) );
  INV_X1 U14509 ( .I(n54395), .ZN(n11324) );
  NOR2_X1 U14510 ( .A1(n5476), .A2(n54392), .ZN(n54369) );
  INV_X1 U14513 ( .I(n56072), .ZN(n56058) );
  INV_X1 U14514 ( .I(n54564), .ZN(n6354) );
  INV_X1 U14516 ( .I(n52301), .ZN(n10833) );
  INV_X1 U14518 ( .I(n54549), .ZN(n6356) );
  NAND2_X1 U14525 ( .A1(n20525), .A2(n53107), .ZN(n23830) );
  AND2_X1 U14526 ( .A1(n63020), .A2(n7680), .Z(n7956) );
  CLKBUF_X2 U14527 ( .I(n55594), .Z(n19183) );
  NOR2_X1 U14528 ( .A1(n2041), .A2(n3285), .ZN(n2039) );
  AND2_X1 U14530 ( .A1(n55503), .A2(n55594), .Z(n15933) );
  INV_X1 U14532 ( .I(n55803), .ZN(n55804) );
  OR2_X1 U14538 ( .A1(n10310), .A2(n7890), .Z(n55134) );
  AND2_X1 U14540 ( .A1(n2049), .A2(n20752), .Z(n54846) );
  AOI21_X1 U14541 ( .A1(n53781), .A2(n58825), .B(n53042), .ZN(n19693) );
  INV_X1 U14546 ( .I(n55038), .ZN(n8412) );
  INV_X1 U14548 ( .I(n56477), .ZN(n56479) );
  NAND2_X1 U14549 ( .A1(n22430), .A2(n20957), .ZN(n56304) );
  INV_X1 U14550 ( .I(n271), .ZN(n11249) );
  CLKBUF_X2 U14551 ( .I(n5193), .Z(n23258) );
  INV_X1 U14554 ( .I(n56816), .ZN(n56766) );
  INV_X2 U14558 ( .I(n25988), .ZN(n3021) );
  CLKBUF_X2 U14560 ( .I(n54901), .Z(n20752) );
  INV_X1 U14561 ( .I(n9424), .ZN(n55363) );
  NOR2_X1 U14563 ( .A1(n9617), .A2(n20560), .ZN(n20559) );
  AND2_X1 U14565 ( .A1(n56182), .A2(n56144), .Z(n15872) );
  AND2_X1 U14566 ( .A1(n1591), .A2(n22430), .Z(n56314) );
  INV_X2 U14570 ( .I(n54383), .ZN(n1586) );
  NAND2_X1 U14575 ( .A1(n1919), .A2(n63020), .ZN(n2493) );
  AND2_X1 U14585 ( .A1(n25268), .A2(n1459), .Z(n15941) );
  CLKBUF_X2 U14591 ( .I(n53998), .Z(n7492) );
  INV_X1 U14595 ( .I(n52223), .ZN(n3307) );
  AND2_X1 U14596 ( .A1(n54876), .A2(n54875), .Z(n54877) );
  AOI21_X1 U14604 ( .A1(n12789), .A2(n12788), .B(n12787), .ZN(n12786) );
  NAND2_X1 U14609 ( .A1(n56260), .A2(n22292), .ZN(n56261) );
  NAND2_X1 U14616 ( .A1(n10845), .A2(n10844), .ZN(n10843) );
  NAND2_X1 U14617 ( .A1(n53022), .A2(n65282), .ZN(n22197) );
  INV_X1 U14622 ( .I(n5041), .ZN(n5040) );
  AOI21_X1 U14627 ( .A1(n10529), .A2(n17375), .B(n17374), .ZN(n14376) );
  INV_X1 U14628 ( .I(n14377), .ZN(n14375) );
  INV_X1 U14629 ( .I(n15509), .ZN(n7061) );
  NAND2_X1 U14630 ( .A1(n18387), .A2(n6391), .ZN(n6390) );
  NAND2_X1 U14632 ( .A1(n5330), .A2(n56359), .ZN(n56236) );
  AOI21_X1 U14633 ( .A1(n12440), .A2(n53197), .B(n12439), .ZN(n52755) );
  OAI21_X1 U14637 ( .A1(n16754), .A2(n9056), .B(n16752), .ZN(n17205) );
  NOR2_X1 U14638 ( .A1(n5886), .A2(n7213), .ZN(n5885) );
  NOR2_X1 U14639 ( .A1(n1176), .A2(n7481), .ZN(n19477) );
  NAND2_X1 U14644 ( .A1(n17376), .A2(n12917), .ZN(n17375) );
  NAND2_X1 U14648 ( .A1(n5419), .A2(n5199), .ZN(n5198) );
  NAND2_X1 U14649 ( .A1(n11939), .A2(n15929), .ZN(n10845) );
  NAND2_X1 U14650 ( .A1(n56280), .A2(n56279), .ZN(n56281) );
  INV_X1 U14657 ( .I(n5278), .ZN(n1957) );
  NAND2_X1 U14660 ( .A1(n51893), .A2(n3616), .ZN(n13859) );
  OAI21_X1 U14662 ( .A1(n10838), .A2(n10837), .B(n10938), .ZN(n10836) );
  INV_X1 U14665 ( .I(n4182), .ZN(n14712) );
  AOI22_X1 U14668 ( .A1(n52486), .A2(n52485), .B1(n52484), .B2(n52483), .ZN(
        n8326) );
  AOI22_X1 U14669 ( .A1(n52234), .A2(n21726), .B1(n52233), .B2(n57036), .ZN(
        n52240) );
  NAND2_X1 U14672 ( .A1(n4375), .A2(n4374), .ZN(n24867) );
  NAND2_X1 U14677 ( .A1(n17329), .A2(n52892), .ZN(n17328) );
  NOR2_X1 U14679 ( .A1(n18927), .A2(n18926), .ZN(n18925) );
  NAND2_X1 U14680 ( .A1(n24311), .A2(n24312), .ZN(n20589) );
  NAND2_X1 U14682 ( .A1(n25499), .A2(n57239), .ZN(n24177) );
  INV_X1 U14686 ( .I(n56127), .ZN(n16330) );
  INV_X1 U14687 ( .I(n20015), .ZN(n20014) );
  AOI21_X1 U14688 ( .A1(n52905), .A2(n54990), .B(n52904), .ZN(n52917) );
  OAI21_X1 U14690 ( .A1(n14804), .A2(n14803), .B(n56229), .ZN(n16642) );
  OAI22_X1 U14694 ( .A1(n56207), .A2(n56638), .B1(n56208), .B2(n56206), .ZN(
        n25410) );
  NAND2_X1 U14695 ( .A1(n53458), .A2(n53457), .ZN(n19353) );
  NAND2_X1 U14697 ( .A1(n65101), .A2(n21248), .ZN(n7555) );
  AOI21_X1 U14699 ( .A1(n17107), .A2(n17106), .B(n1455), .ZN(n14322) );
  NOR2_X1 U14700 ( .A1(n3884), .A2(n54596), .ZN(n6442) );
  NOR2_X1 U14701 ( .A1(n21617), .A2(n15761), .ZN(n18927) );
  OAI21_X1 U14710 ( .A1(n19615), .A2(n19614), .B(n15975), .ZN(n13248) );
  AOI21_X1 U14711 ( .A1(n12290), .A2(n53382), .B(n12289), .ZN(n50672) );
  NAND2_X1 U14712 ( .A1(n52279), .A2(n23526), .ZN(n14577) );
  NAND2_X1 U14713 ( .A1(n57043), .A2(n57042), .ZN(n57044) );
  NOR2_X1 U14714 ( .A1(n54781), .A2(n59879), .ZN(n8903) );
  OAI21_X1 U14720 ( .A1(n51898), .A2(n51897), .B(n51900), .ZN(n24219) );
  NOR2_X1 U14722 ( .A1(n53538), .A2(n19485), .ZN(n19484) );
  NOR2_X1 U14723 ( .A1(n53224), .A2(n53225), .ZN(n53229) );
  OAI21_X1 U14725 ( .A1(n55667), .A2(n55666), .B(n9649), .ZN(n18851) );
  NAND2_X1 U14728 ( .A1(n8448), .A2(n3127), .ZN(n8447) );
  AND2_X1 U14732 ( .A1(n51456), .A2(n56211), .Z(n56413) );
  NOR2_X1 U14733 ( .A1(n20756), .A2(n1458), .ZN(n17838) );
  NOR2_X1 U14735 ( .A1(n57053), .A2(n23248), .ZN(n13422) );
  NOR2_X1 U14737 ( .A1(n7764), .A2(n18255), .ZN(n7763) );
  OAI21_X1 U14738 ( .A1(n25215), .A2(n54961), .B(n2679), .ZN(n54964) );
  INV_X1 U14740 ( .I(n5420), .ZN(n5419) );
  OAI22_X1 U14741 ( .A1(n869), .A2(n14469), .B1(n52382), .B2(n54944), .ZN(
        n7801) );
  INV_X1 U14742 ( .I(n54993), .ZN(n1960) );
  AOI21_X1 U14743 ( .A1(n52744), .A2(n53397), .B(n1180), .ZN(n52748) );
  NAND3_X1 U14744 ( .A1(n57239), .A2(n56554), .A3(n13067), .ZN(n51558) );
  AOI21_X1 U14745 ( .A1(n4126), .A2(n4124), .B(n4121), .ZN(n6462) );
  NAND3_X1 U14747 ( .A1(n52387), .A2(n52386), .A3(n52385), .ZN(n52388) );
  NOR2_X1 U14748 ( .A1(n24142), .A2(n55913), .ZN(n24141) );
  NAND2_X1 U14754 ( .A1(n55977), .A2(n55979), .ZN(n6009) );
  NAND2_X1 U14757 ( .A1(n6464), .A2(n3884), .ZN(n6463) );
  NOR2_X1 U14760 ( .A1(n12535), .A2(n12534), .ZN(n51254) );
  OAI21_X1 U14762 ( .A1(n6395), .A2(n23376), .B(n11121), .ZN(n4740) );
  NOR2_X1 U14763 ( .A1(n17260), .A2(n17259), .ZN(n17258) );
  NAND2_X1 U14764 ( .A1(n52790), .A2(n53436), .ZN(n4116) );
  OAI21_X1 U14765 ( .A1(n11990), .A2(n18269), .B(n56398), .ZN(n18387) );
  INV_X1 U14766 ( .I(n24729), .ZN(n25499) );
  NAND2_X1 U14767 ( .A1(n4255), .A2(n1145), .ZN(n4254) );
  NAND2_X1 U14768 ( .A1(n53546), .A2(n11938), .ZN(n10844) );
  INV_X1 U14771 ( .I(n55717), .ZN(n4375) );
  NAND2_X1 U14772 ( .A1(n24904), .A2(n24903), .ZN(n9266) );
  AOI22_X1 U14774 ( .A1(n64187), .A2(n19356), .B1(n56253), .B2(n56254), .ZN(
        n56260) );
  NAND3_X1 U14776 ( .A1(n16866), .A2(n19401), .A3(n16865), .ZN(n19400) );
  OAI22_X1 U14777 ( .A1(n56627), .A2(n21069), .B1(n56620), .B2(n59449), .ZN(
        n8830) );
  OAI21_X1 U14779 ( .A1(n1147), .A2(n6531), .B(n14351), .ZN(n55483) );
  INV_X1 U14781 ( .I(n18790), .ZN(n55260) );
  OAI21_X1 U14782 ( .A1(n4025), .A2(n21453), .B(n6943), .ZN(n4021) );
  OAI21_X1 U14784 ( .A1(n15180), .A2(n15179), .B(n56564), .ZN(n55944) );
  NOR2_X1 U14785 ( .A1(n53549), .A2(n53547), .ZN(n10839) );
  NAND2_X1 U14786 ( .A1(n9263), .A2(n55974), .ZN(n55449) );
  NAND2_X1 U14787 ( .A1(n51253), .A2(n23377), .ZN(n6395) );
  NAND2_X1 U14788 ( .A1(n57022), .A2(n12818), .ZN(n17553) );
  NOR2_X1 U14789 ( .A1(n21728), .A2(n21582), .ZN(n21727) );
  NAND2_X1 U14790 ( .A1(n51252), .A2(n56396), .ZN(n12535) );
  INV_X1 U14792 ( .I(n55978), .ZN(n6010) );
  NAND2_X1 U14794 ( .A1(n55430), .A2(n10949), .ZN(n50951) );
  NOR2_X1 U14797 ( .A1(n54995), .A2(n7583), .ZN(n54645) );
  NAND2_X1 U14799 ( .A1(n52390), .A2(n52931), .ZN(n7896) );
  INV_X1 U14803 ( .I(n21582), .ZN(n21726) );
  NAND2_X1 U14804 ( .A1(n55666), .A2(n8595), .ZN(n9649) );
  NOR2_X1 U14809 ( .A1(n58326), .A2(n21235), .ZN(n25435) );
  NAND2_X1 U14812 ( .A1(n53403), .A2(n53402), .ZN(n53404) );
  NAND2_X1 U14813 ( .A1(n57041), .A2(n57040), .ZN(n57043) );
  NAND2_X1 U14814 ( .A1(n16644), .A2(n23095), .ZN(n14756) );
  OR3_X1 U14815 ( .A1(n52708), .A2(n56381), .A3(n52707), .Z(n52709) );
  NAND2_X1 U14816 ( .A1(n54643), .A2(n54854), .ZN(n3945) );
  NAND2_X1 U14818 ( .A1(n53238), .A2(n59858), .ZN(n52265) );
  NAND2_X1 U14819 ( .A1(n52133), .A2(n19030), .ZN(n21270) );
  OR3_X1 U14820 ( .A1(n12074), .A2(n54843), .A3(n5279), .Z(n54649) );
  NOR2_X1 U14821 ( .A1(n50546), .A2(n1283), .ZN(n23323) );
  NOR2_X1 U14823 ( .A1(n24674), .A2(n24675), .ZN(n24673) );
  NOR2_X1 U14824 ( .A1(n53438), .A2(n833), .ZN(n13402) );
  INV_X1 U14825 ( .I(n11121), .ZN(n12555) );
  AND2_X1 U14826 ( .A1(n21081), .A2(n16753), .Z(n16752) );
  INV_X1 U14827 ( .I(n16043), .ZN(n13143) );
  INV_X1 U14829 ( .I(n54296), .ZN(n2679) );
  NAND2_X1 U14830 ( .A1(n7765), .A2(n11121), .ZN(n7764) );
  AND3_X1 U14831 ( .A1(n55298), .A2(n55304), .A3(n52918), .Z(n15947) );
  AOI21_X1 U14832 ( .A1(n53606), .A2(n53194), .B(n64910), .ZN(n53195) );
  AOI21_X1 U14835 ( .A1(n11524), .A2(n56265), .B(n13020), .ZN(n13018) );
  INV_X1 U14836 ( .I(n5049), .ZN(n22258) );
  NAND2_X1 U14838 ( .A1(n8446), .A2(n57037), .ZN(n8445) );
  OR2_X1 U14839 ( .A1(n54500), .A2(n24509), .Z(n53841) );
  INV_X1 U14844 ( .I(n54084), .ZN(n54081) );
  NOR2_X1 U14847 ( .A1(n52827), .A2(n12818), .ZN(n19320) );
  OAI21_X1 U14848 ( .A1(n5736), .A2(n54471), .B(n5735), .ZN(n6220) );
  OAI21_X1 U14850 ( .A1(n23526), .A2(n59461), .B(n12468), .ZN(n56560) );
  NAND2_X1 U14851 ( .A1(n57225), .A2(n20653), .ZN(n9866) );
  AOI21_X1 U14858 ( .A1(n53208), .A2(n53445), .B(n53207), .ZN(n12787) );
  NOR2_X1 U14859 ( .A1(n2997), .A2(n1453), .ZN(n9124) );
  OR2_X1 U14861 ( .A1(n55496), .A2(n17979), .Z(n15993) );
  NAND3_X1 U14862 ( .A1(n5057), .A2(n5056), .A3(n54096), .ZN(n18929) );
  NAND2_X1 U14863 ( .A1(n24696), .A2(n13067), .ZN(n26156) );
  NAND2_X1 U14864 ( .A1(n15822), .A2(n4125), .ZN(n4124) );
  NAND2_X1 U14866 ( .A1(n54981), .A2(n54980), .ZN(n8397) );
  NOR2_X1 U14867 ( .A1(n4123), .A2(n62944), .ZN(n4121) );
  OR2_X1 U14873 ( .A1(n16487), .A2(n54110), .Z(n53875) );
  INV_X1 U14874 ( .I(n56636), .ZN(n56219) );
  NOR2_X1 U14875 ( .A1(n56225), .A2(n56430), .ZN(n16754) );
  INV_X1 U14876 ( .I(n57012), .ZN(n24534) );
  OAI22_X1 U14877 ( .A1(n57404), .A2(n4783), .B1(n21877), .B2(n54943), .ZN(
        n54941) );
  NAND2_X1 U14880 ( .A1(n23482), .A2(n54028), .ZN(n53882) );
  NOR2_X1 U14881 ( .A1(n53205), .A2(n3127), .ZN(n50804) );
  OR2_X1 U14882 ( .A1(n55442), .A2(n14225), .Z(n52954) );
  OAI22_X1 U14884 ( .A1(n56228), .A2(n21081), .B1(n56227), .B2(n56226), .ZN(
        n14803) );
  NOR2_X1 U14885 ( .A1(n52951), .A2(n55442), .ZN(n16384) );
  INV_X1 U14887 ( .I(n57029), .ZN(n57034) );
  NOR2_X1 U14891 ( .A1(n19644), .A2(n15485), .ZN(n15484) );
  NOR2_X1 U14892 ( .A1(n55941), .A2(n56567), .ZN(n15180) );
  NAND2_X1 U14895 ( .A1(n61902), .A2(n56985), .ZN(n23625) );
  INV_X1 U14896 ( .I(n54022), .ZN(n54352) );
  NOR2_X1 U14898 ( .A1(n22749), .A2(n54945), .ZN(n2864) );
  NOR2_X1 U14899 ( .A1(n56268), .A2(n24944), .ZN(n14541) );
  NAND2_X1 U14900 ( .A1(n56393), .A2(n11119), .ZN(n11118) );
  NAND2_X1 U14902 ( .A1(n55976), .A2(n3567), .ZN(n52009) );
  INV_X1 U14905 ( .I(n54611), .ZN(n13112) );
  NAND2_X1 U14906 ( .A1(n1370), .A2(n55926), .ZN(n5495) );
  INV_X1 U14907 ( .I(n54452), .ZN(n4126) );
  NAND2_X1 U14908 ( .A1(n54350), .A2(n54349), .ZN(n11394) );
  NOR2_X1 U14911 ( .A1(n5737), .A2(n54599), .ZN(n5736) );
  AND2_X1 U14912 ( .A1(n59831), .A2(n23704), .Z(n17374) );
  AOI21_X1 U14914 ( .A1(n55415), .A2(n55249), .B(n24676), .ZN(n24674) );
  NAND2_X1 U14916 ( .A1(n12282), .A2(n59827), .ZN(n56553) );
  INV_X1 U14917 ( .I(n2903), .ZN(n52881) );
  OAI21_X1 U14918 ( .A1(n818), .A2(n54594), .B(n54473), .ZN(n54474) );
  NOR2_X1 U14919 ( .A1(n51707), .A2(n54471), .ZN(n7791) );
  NAND2_X1 U14920 ( .A1(n54469), .A2(n7787), .ZN(n7786) );
  OR2_X1 U14921 ( .A1(n52816), .A2(n52820), .Z(n52817) );
  NAND2_X1 U14922 ( .A1(n20850), .A2(n55914), .ZN(n9490) );
  NOR2_X1 U14923 ( .A1(n17601), .A2(n52126), .ZN(n17607) );
  OAI21_X1 U14928 ( .A1(n14879), .A2(n55709), .B(n62261), .ZN(n55712) );
  NAND3_X1 U14933 ( .A1(n53580), .A2(n57183), .A3(n21082), .ZN(n53582) );
  NOR2_X1 U14934 ( .A1(n59081), .A2(n54613), .ZN(n4239) );
  OR2_X1 U14935 ( .A1(n53031), .A2(n21697), .Z(n16175) );
  NOR2_X1 U14936 ( .A1(n55427), .A2(n55426), .ZN(n8968) );
  OAI22_X1 U14937 ( .A1(n52737), .A2(n4184), .B1(n25160), .B2(n1372), .ZN(
        n13723) );
  INV_X1 U14938 ( .I(n55452), .ZN(n55453) );
  AOI21_X1 U14939 ( .A1(n55418), .A2(n65011), .B(n61065), .ZN(n15681) );
  OR2_X1 U14940 ( .A1(n56627), .A2(n9388), .Z(n56419) );
  INV_X1 U14944 ( .I(n2201), .ZN(n2200) );
  AND2_X1 U14947 ( .A1(n54470), .A2(n54594), .Z(n22337) );
  INV_X1 U14948 ( .I(n21235), .ZN(n25437) );
  NOR2_X1 U14949 ( .A1(n52673), .A2(n57068), .ZN(n10191) );
  OR2_X1 U14951 ( .A1(n56393), .A2(n56567), .Z(n56278) );
  INV_X1 U14953 ( .I(n55437), .ZN(n14225) );
  INV_X1 U14955 ( .I(n55407), .ZN(n52548) );
  AND2_X1 U14956 ( .A1(n13940), .A2(n53547), .Z(n5656) );
  INV_X1 U14957 ( .I(n54108), .ZN(n53872) );
  OR2_X1 U14958 ( .A1(n54594), .A2(n23736), .Z(n54324) );
  INV_X1 U14961 ( .I(n6211), .ZN(n5737) );
  AND3_X1 U14963 ( .A1(n56412), .A2(n23952), .A3(n57691), .Z(n16046) );
  NAND2_X1 U14964 ( .A1(n52668), .A2(n57061), .ZN(n52669) );
  NAND2_X1 U14966 ( .A1(n56393), .A2(n10183), .ZN(n12553) );
  AND2_X1 U14972 ( .A1(n52946), .A2(n55265), .Z(n8060) );
  INV_X2 U14974 ( .I(n54825), .ZN(n54446) );
  AND2_X1 U14975 ( .A1(n54823), .A2(n15040), .Z(n20095) );
  NOR2_X1 U14978 ( .A1(n56268), .A2(n23447), .ZN(n11523) );
  AND2_X1 U14979 ( .A1(n18597), .A2(n56434), .Z(n16115) );
  INV_X2 U14980 ( .I(n17499), .ZN(n55022) );
  NAND2_X1 U14984 ( .A1(n58626), .A2(n4194), .ZN(n22381) );
  NAND2_X1 U14986 ( .A1(n22760), .A2(n17936), .ZN(n54849) );
  AND2_X1 U14987 ( .A1(n56403), .A2(n56585), .Z(n16160) );
  AND2_X1 U14992 ( .A1(n54088), .A2(n54594), .Z(n7787) );
  OR2_X1 U14996 ( .A1(n54605), .A2(n26095), .Z(n54613) );
  NAND2_X1 U15001 ( .A1(n2062), .A2(n54651), .ZN(n54652) );
  NAND2_X1 U15003 ( .A1(n7148), .A2(n61472), .ZN(n4123) );
  OR2_X1 U15006 ( .A1(n16629), .A2(n56435), .Z(n56226) );
  BUF_X2 U15009 ( .I(n52117), .Z(n55433) );
  INV_X2 U15013 ( .I(n1287), .ZN(n12574) );
  CLKBUF_X2 U15016 ( .I(n54347), .Z(n4564) );
  CLKBUF_X2 U15017 ( .I(n25252), .Z(n23952) );
  INV_X1 U15021 ( .I(n17555), .ZN(n21706) );
  INV_X2 U15023 ( .I(n25168), .ZN(n55936) );
  CLKBUF_X2 U15026 ( .I(n55909), .Z(n23360) );
  AND2_X2 U15031 ( .A1(n6115), .A2(n6116), .Z(n25215) );
  INV_X2 U15036 ( .I(n25948), .ZN(n53383) );
  AND2_X1 U15037 ( .A1(n55306), .A2(n55440), .Z(n16073) );
  INV_X4 U15039 ( .I(n15931), .ZN(n19434) );
  INV_X2 U15042 ( .I(n53031), .ZN(n1611) );
  CLKBUF_X4 U15057 ( .I(n55494), .Z(n18109) );
  BUF_X2 U15061 ( .I(n54615), .Z(n2199) );
  BUF_X2 U15063 ( .I(n50594), .Z(n52857) );
  INV_X1 U15064 ( .I(n54615), .ZN(n2198) );
  CLKBUF_X2 U15067 ( .I(n54998), .Z(n23275) );
  INV_X1 U15069 ( .I(n24284), .ZN(n12598) );
  INV_X2 U15070 ( .I(n24226), .ZN(n56435) );
  BUF_X2 U15071 ( .I(n55676), .Z(n15730) );
  BUF_X4 U15074 ( .I(n51676), .Z(n54594) );
  INV_X1 U15078 ( .I(n23032), .ZN(n22660) );
  INV_X1 U15079 ( .I(n22241), .ZN(n21260) );
  INV_X1 U15083 ( .I(n50644), .ZN(n8856) );
  BUF_X2 U15084 ( .I(n13156), .Z(n10896) );
  BUF_X2 U15085 ( .I(n25395), .Z(n2167) );
  INV_X1 U15087 ( .I(n51003), .ZN(n9298) );
  INV_X1 U15088 ( .I(n51975), .ZN(n9192) );
  INV_X1 U15092 ( .I(n50948), .ZN(n8477) );
  INV_X1 U15093 ( .I(n24776), .ZN(n3863) );
  INV_X1 U15094 ( .I(n16095), .ZN(n8792) );
  CLKBUF_X2 U15096 ( .I(n51987), .Z(n23885) );
  INV_X1 U15097 ( .I(n52637), .ZN(n10252) );
  INV_X1 U15098 ( .I(n51318), .ZN(n12566) );
  INV_X1 U15099 ( .I(n24650), .ZN(n52202) );
  CLKBUF_X2 U15100 ( .I(n10476), .Z(n7070) );
  INV_X1 U15101 ( .I(n52147), .ZN(n2184) );
  CLKBUF_X2 U15102 ( .I(n52541), .Z(n22530) );
  INV_X1 U15103 ( .I(n2933), .ZN(n16960) );
  INV_X1 U15106 ( .I(n12119), .ZN(n52414) );
  INV_X1 U15109 ( .I(n6363), .ZN(n1975) );
  INV_X1 U15110 ( .I(n24739), .ZN(n51043) );
  INV_X2 U15114 ( .I(n25542), .ZN(n1618) );
  INV_X1 U15115 ( .I(n19888), .ZN(n14993) );
  INV_X1 U15121 ( .I(n18644), .ZN(n19688) );
  INV_X1 U15124 ( .I(n50979), .ZN(n10724) );
  INV_X1 U15126 ( .I(n51502), .ZN(n9868) );
  CLKBUF_X2 U15128 ( .I(n21794), .Z(n21097) );
  INV_X1 U15138 ( .I(n17127), .ZN(n6383) );
  INV_X1 U15144 ( .I(n48946), .ZN(n24397) );
  INV_X1 U15145 ( .I(n22153), .ZN(n13885) );
  INV_X1 U15147 ( .I(n52331), .ZN(n20780) );
  INV_X1 U15149 ( .I(n51583), .ZN(n5143) );
  BUF_X2 U15151 ( .I(n2222), .Z(n9506) );
  CLKBUF_X2 U15152 ( .I(n51144), .Z(n23288) );
  INV_X1 U15154 ( .I(n12765), .ZN(n12007) );
  CLKBUF_X2 U15157 ( .I(n51629), .Z(n22305) );
  INV_X1 U15159 ( .I(n2603), .ZN(n15653) );
  CLKBUF_X2 U15162 ( .I(n18486), .Z(n18485) );
  INV_X1 U15163 ( .I(n24074), .ZN(n50670) );
  OAI21_X1 U15164 ( .A1(n13317), .A2(n49198), .B(n49525), .ZN(n49199) );
  NAND2_X1 U15168 ( .A1(n49506), .A2(n49507), .ZN(n5764) );
  CLKBUF_X2 U15171 ( .I(n52453), .Z(n23697) );
  NAND2_X1 U15172 ( .A1(n13886), .A2(n49871), .ZN(n51956) );
  NAND2_X1 U15177 ( .A1(n14779), .A2(n3695), .ZN(n49523) );
  NAND3_X1 U15178 ( .A1(n48939), .A2(n48938), .A3(n49436), .ZN(n8714) );
  OAI21_X1 U15184 ( .A1(n47762), .A2(n8726), .B(n4614), .ZN(n8723) );
  INV_X1 U15188 ( .I(n9156), .ZN(n9155) );
  NAND2_X1 U15189 ( .A1(n23614), .A2(n46778), .ZN(n19782) );
  NOR2_X1 U15190 ( .A1(n4826), .A2(n4825), .ZN(n47071) );
  CLKBUF_X2 U15194 ( .I(n52360), .Z(n4846) );
  INV_X1 U15197 ( .I(n25535), .ZN(n5765) );
  NAND2_X1 U15199 ( .A1(n18430), .A2(n15526), .ZN(n18271) );
  NAND3_X1 U15201 ( .A1(n10486), .A2(n25549), .A3(n56905), .ZN(n12764) );
  NAND2_X1 U15206 ( .A1(n2246), .A2(n2245), .ZN(n11004) );
  AOI21_X1 U15211 ( .A1(n48744), .A2(n10715), .B(n10714), .ZN(n48746) );
  NAND2_X1 U15212 ( .A1(n4300), .A2(n4299), .ZN(n4298) );
  OAI21_X1 U15213 ( .A1(n49945), .A2(n50277), .B(n62244), .ZN(n49953) );
  INV_X1 U15217 ( .I(n11218), .ZN(n11217) );
  INV_X1 U15218 ( .I(n11615), .ZN(n12330) );
  NAND2_X1 U15220 ( .A1(n12367), .A2(n12370), .ZN(n5579) );
  AOI21_X1 U15221 ( .A1(n48290), .A2(n3679), .B(n3678), .ZN(n3677) );
  INV_X1 U15222 ( .I(n12924), .ZN(n50274) );
  NOR2_X1 U15224 ( .A1(n48898), .A2(n6931), .ZN(n4579) );
  INV_X1 U15227 ( .I(n18083), .ZN(n8621) );
  NAND2_X1 U15229 ( .A1(n46084), .A2(n46083), .ZN(n4011) );
  AOI21_X1 U15237 ( .A1(n3919), .A2(n48075), .B(n3918), .ZN(n3917) );
  INV_X1 U15243 ( .I(n48311), .ZN(n9380) );
  OAI21_X1 U15244 ( .A1(n15068), .A2(n48065), .B(n11057), .ZN(n15067) );
  INV_X1 U15245 ( .I(n5697), .ZN(n5696) );
  NOR2_X1 U15246 ( .A1(n18184), .A2(n48771), .ZN(n9824) );
  AOI21_X1 U15247 ( .A1(n10334), .A2(n19219), .B(n19144), .ZN(n16233) );
  AOI21_X1 U15249 ( .A1(n22867), .A2(n57193), .B(n22489), .ZN(n22488) );
  NAND2_X1 U15252 ( .A1(n3845), .A2(n49195), .ZN(n3844) );
  INV_X1 U15254 ( .I(n48989), .ZN(n2647) );
  INV_X1 U15255 ( .I(n47558), .ZN(n13096) );
  NAND2_X1 U15257 ( .A1(n24267), .A2(n24266), .ZN(n10825) );
  INV_X1 U15258 ( .I(n49354), .ZN(n17017) );
  NAND2_X1 U15259 ( .A1(n1104), .A2(n17165), .ZN(n24917) );
  NOR2_X1 U15260 ( .A1(n6610), .A2(n3885), .ZN(n5637) );
  NOR2_X1 U15263 ( .A1(n48003), .A2(n12335), .ZN(n12334) );
  NAND2_X1 U15264 ( .A1(n11887), .A2(n49391), .ZN(n11886) );
  NOR2_X1 U15268 ( .A1(n4503), .A2(n49095), .ZN(n48017) );
  OAI22_X1 U15270 ( .A1(n50449), .A2(n50448), .B1(n50447), .B2(n8878), .ZN(
        n25274) );
  NAND2_X1 U15271 ( .A1(n48820), .A2(n48821), .ZN(n5700) );
  NAND2_X1 U15274 ( .A1(n48073), .A2(n4412), .ZN(n48075) );
  NAND3_X1 U15275 ( .A1(n48862), .A2(n20686), .A3(n16188), .ZN(n48866) );
  OAI22_X1 U15277 ( .A1(n48321), .A2(n7015), .B1(n48324), .B2(n7014), .ZN(
        n7013) );
  INV_X1 U15278 ( .I(n49272), .ZN(n5714) );
  OAI21_X1 U15280 ( .A1(n11290), .A2(n11289), .B(n23156), .ZN(n7652) );
  OAI21_X1 U15281 ( .A1(n49703), .A2(n19302), .B(n4598), .ZN(n49766) );
  NOR2_X1 U15282 ( .A1(n49711), .A2(n14097), .ZN(n46964) );
  INV_X1 U15283 ( .I(n48061), .ZN(n15068) );
  AOI21_X1 U15286 ( .A1(n9535), .A2(n49455), .B(n49454), .ZN(n9534) );
  NAND2_X1 U15287 ( .A1(n49724), .A2(n9409), .ZN(n9408) );
  NOR2_X1 U15290 ( .A1(n14072), .A2(n49843), .ZN(n14070) );
  NAND2_X1 U15291 ( .A1(n48706), .A2(n48705), .ZN(n25039) );
  NAND2_X1 U15295 ( .A1(n49219), .A2(n49220), .ZN(n13972) );
  NOR2_X1 U15297 ( .A1(n49103), .A2(n18081), .ZN(n18080) );
  AOI22_X1 U15298 ( .A1(n49228), .A2(n49229), .B1(n13121), .B2(n49739), .ZN(
        n24266) );
  NOR2_X1 U15300 ( .A1(n49700), .A2(n48680), .ZN(n6931) );
  AOI21_X1 U15302 ( .A1(n49105), .A2(n49104), .B(n18079), .ZN(n18078) );
  NOR2_X1 U15303 ( .A1(n6930), .A2(n6929), .ZN(n4580) );
  INV_X1 U15304 ( .I(n48367), .ZN(n48368) );
  OAI21_X1 U15306 ( .A1(n48794), .A2(n48429), .B(n48810), .ZN(n10906) );
  NAND2_X1 U15307 ( .A1(n48890), .A2(n49703), .ZN(n15625) );
  NOR2_X1 U15310 ( .A1(n23373), .A2(n47995), .ZN(n48000) );
  NOR2_X1 U15311 ( .A1(n9306), .A2(n48925), .ZN(n9696) );
  NAND2_X1 U15313 ( .A1(n17883), .A2(n24768), .ZN(n15302) );
  INV_X1 U15316 ( .I(n16730), .ZN(n49298) );
  NAND2_X1 U15321 ( .A1(n49815), .A2(n22264), .ZN(n8896) );
  NOR2_X1 U15322 ( .A1(n17125), .A2(n49452), .ZN(n17122) );
  NOR2_X1 U15328 ( .A1(n3701), .A2(n47968), .ZN(n3700) );
  INV_X1 U15330 ( .I(n48004), .ZN(n3845) );
  NAND2_X1 U15331 ( .A1(n17682), .A2(n17684), .ZN(n17681) );
  OAI21_X1 U15342 ( .A1(n11351), .A2(n48454), .B(n9853), .ZN(n48456) );
  OAI21_X1 U15343 ( .A1(n48776), .A2(n48775), .B(n48774), .ZN(n3595) );
  INV_X1 U15348 ( .I(n48354), .ZN(n49765) );
  INV_X1 U15352 ( .I(n8878), .ZN(n50446) );
  OAI22_X1 U15353 ( .A1(n47944), .A2(n15220), .B1(n63605), .B2(n49115), .ZN(
        n47945) );
  NOR2_X1 U15354 ( .A1(n50444), .A2(n7867), .ZN(n50022) );
  OAI22_X1 U15355 ( .A1(n48872), .A2(n48871), .B1(n48874), .B2(n48873), .ZN(
        n22320) );
  INV_X1 U15357 ( .I(n49288), .ZN(n7214) );
  NAND2_X1 U15358 ( .A1(n20663), .A2(n20662), .ZN(n20661) );
  OAI21_X1 U15361 ( .A1(n4204), .A2(n149), .B(n47976), .ZN(n4203) );
  NOR2_X1 U15363 ( .A1(n5713), .A2(n49410), .ZN(n49269) );
  NOR2_X1 U15365 ( .A1(n7454), .A2(n48059), .ZN(n48984) );
  INV_X1 U15366 ( .I(n49453), .ZN(n9535) );
  OAI21_X1 U15368 ( .A1(n21269), .A2(n11705), .B(n49069), .ZN(n20237) );
  NAND2_X1 U15369 ( .A1(n49388), .A2(n49387), .ZN(n14032) );
  NAND2_X1 U15372 ( .A1(n49047), .A2(n64167), .ZN(n12370) );
  OAI21_X1 U15374 ( .A1(n49562), .A2(n49563), .B(n63493), .ZN(n17968) );
  NAND2_X1 U15375 ( .A1(n9367), .A2(n49488), .ZN(n48394) );
  NAND2_X1 U15376 ( .A1(n49385), .A2(n49386), .ZN(n14033) );
  OAI21_X1 U15377 ( .A1(n49326), .A2(n49327), .B(n7078), .ZN(n49335) );
  INV_X1 U15379 ( .I(n49073), .ZN(n48305) );
  NOR2_X1 U15381 ( .A1(n49552), .A2(n25128), .ZN(n18371) );
  NAND3_X1 U15382 ( .A1(n12496), .A2(n49316), .A3(n11172), .ZN(n47447) );
  INV_X1 U15383 ( .I(n49839), .ZN(n26189) );
  NAND2_X1 U15384 ( .A1(n49360), .A2(n3351), .ZN(n3350) );
  AND2_X1 U15386 ( .A1(n50269), .A2(n61170), .Z(n25831) );
  NAND2_X1 U15387 ( .A1(n7078), .A2(n15753), .ZN(n11892) );
  NAND2_X1 U15388 ( .A1(n47935), .A2(n14065), .ZN(n15603) );
  OAI22_X1 U15390 ( .A1(n48072), .A2(n49060), .B1(n48071), .B2(n1474), .ZN(
        n3918) );
  NOR2_X1 U15391 ( .A1(n50276), .A2(n62244), .ZN(n50278) );
  AND2_X1 U15393 ( .A1(n11184), .A2(n6323), .Z(n3919) );
  NOR2_X1 U15399 ( .A1(n47926), .A2(n49723), .ZN(n15602) );
  NOR2_X1 U15402 ( .A1(n48923), .A2(n16084), .ZN(n48369) );
  NOR2_X1 U15403 ( .A1(n25263), .A2(n24622), .ZN(n6367) );
  NOR2_X1 U15406 ( .A1(n48453), .A2(n48323), .ZN(n47052) );
  NAND2_X1 U15409 ( .A1(n17126), .A2(n3646), .ZN(n17125) );
  NAND2_X1 U15410 ( .A1(n3646), .A2(n61070), .ZN(n17124) );
  NAND2_X1 U15412 ( .A1(n45613), .A2(n49846), .ZN(n17516) );
  NAND2_X1 U15417 ( .A1(n17335), .A2(n5591), .ZN(n49302) );
  NAND2_X1 U15419 ( .A1(n49697), .A2(n48349), .ZN(n6929) );
  AOI21_X1 U15422 ( .A1(n49740), .A2(n49741), .B(n10831), .ZN(n49745) );
  OAI21_X1 U15423 ( .A1(n1638), .A2(n49315), .B(n17874), .ZN(n9443) );
  NAND2_X1 U15424 ( .A1(n49495), .A2(n64335), .ZN(n9292) );
  NAND2_X1 U15425 ( .A1(n3646), .A2(n49849), .ZN(n14072) );
  NAND2_X1 U15426 ( .A1(n47766), .A2(n7866), .ZN(n8726) );
  NAND4_X1 U15427 ( .A1(n49062), .A2(n17816), .A3(n49077), .A4(n49835), .ZN(
        n45700) );
  NAND3_X1 U15428 ( .A1(n49936), .A2(n50348), .A3(n49934), .ZN(n48142) );
  NAND2_X1 U15429 ( .A1(n49191), .A2(n49510), .ZN(n49194) );
  NAND2_X1 U15432 ( .A1(n15213), .A2(n49172), .ZN(n49173) );
  NOR2_X1 U15434 ( .A1(n10760), .A2(n49606), .ZN(n15848) );
  NOR2_X1 U15435 ( .A1(n48996), .A2(n11820), .ZN(n48706) );
  NAND2_X1 U15437 ( .A1(n49467), .A2(n59966), .ZN(n13121) );
  NAND2_X1 U15440 ( .A1(n48426), .A2(n48427), .ZN(n18239) );
  NOR2_X1 U15442 ( .A1(n26102), .A2(n49767), .ZN(n49784) );
  INV_X1 U15445 ( .I(n20204), .ZN(n49244) );
  INV_X1 U15447 ( .I(n49009), .ZN(n15475) );
  NAND2_X1 U15448 ( .A1(n48407), .A2(n26102), .ZN(n4297) );
  NAND2_X1 U15449 ( .A1(n50093), .A2(n50092), .ZN(n4192) );
  INV_X1 U15450 ( .I(n49018), .ZN(n6716) );
  AOI21_X1 U15451 ( .A1(n15906), .A2(n22926), .B(n61355), .ZN(n49620) );
  OAI21_X1 U15452 ( .A1(n49009), .A2(n49008), .B(n49007), .ZN(n11639) );
  NOR2_X1 U15453 ( .A1(n49767), .A2(n21737), .ZN(n21943) );
  NOR2_X1 U15454 ( .A1(n18625), .A2(n61016), .ZN(n3699) );
  INV_X1 U15455 ( .I(n17793), .ZN(n3701) );
  NAND2_X1 U15456 ( .A1(n63664), .A2(n49711), .ZN(n17090) );
  NOR2_X1 U15460 ( .A1(n19706), .A2(n19705), .ZN(n19704) );
  AND3_X1 U15462 ( .A1(n49266), .A2(n49410), .A3(n49177), .Z(n48964) );
  NAND2_X1 U15463 ( .A1(n12616), .A2(n62033), .ZN(n8711) );
  OR2_X1 U15466 ( .A1(n48039), .A2(n48323), .Z(n6610) );
  AOI21_X1 U15467 ( .A1(n48860), .A2(n9354), .B(n9353), .ZN(n48862) );
  NAND2_X1 U15469 ( .A1(n23500), .A2(n48863), .ZN(n20686) );
  AOI21_X1 U15472 ( .A1(n49138), .A2(n49999), .B(n61375), .ZN(n49139) );
  NOR2_X1 U15478 ( .A1(n1472), .A2(n48453), .ZN(n11351) );
  OAI21_X1 U15480 ( .A1(n49886), .A2(n18608), .B(n57265), .ZN(n13149) );
  INV_X1 U15481 ( .I(n12496), .ZN(n48308) );
  NAND2_X1 U15483 ( .A1(n50291), .A2(n57182), .ZN(n10263) );
  NOR2_X1 U15489 ( .A1(n49767), .A2(n4207), .ZN(n4206) );
  AOI21_X1 U15490 ( .A1(n2868), .A2(n49642), .B(n3065), .ZN(n19520) );
  AOI21_X1 U15491 ( .A1(n48008), .A2(n20971), .B(n49682), .ZN(n4503) );
  AND2_X1 U15492 ( .A1(n48947), .A2(n12845), .Z(n16294) );
  NOR2_X1 U15493 ( .A1(n48948), .A2(n4310), .ZN(n4733) );
  INV_X1 U15496 ( .I(n2983), .ZN(n2982) );
  NAND2_X1 U15501 ( .A1(n15634), .A2(n502), .ZN(n24691) );
  NAND2_X1 U15502 ( .A1(n49919), .A2(n2981), .ZN(n2980) );
  NAND2_X1 U15503 ( .A1(n49643), .A2(n19523), .ZN(n9241) );
  NOR2_X1 U15505 ( .A1(n22869), .A2(n4258), .ZN(n12842) );
  INV_X1 U15506 ( .I(n4418), .ZN(n4417) );
  NOR2_X1 U15507 ( .A1(n48020), .A2(n48832), .ZN(n9324) );
  NAND2_X1 U15508 ( .A1(n19866), .A2(n49170), .ZN(n13633) );
  INV_X1 U15510 ( .I(n46729), .ZN(n50412) );
  INV_X1 U15511 ( .I(n18565), .ZN(n3351) );
  AND2_X1 U15512 ( .A1(n5283), .A2(n15386), .Z(n15906) );
  INV_X1 U15515 ( .I(n4436), .ZN(n44794) );
  INV_X1 U15517 ( .I(n4258), .ZN(n48407) );
  INV_X1 U15518 ( .I(n49641), .ZN(n2868) );
  NAND2_X1 U15519 ( .A1(n48579), .A2(n21537), .ZN(n9500) );
  NAND2_X1 U15520 ( .A1(n49388), .A2(n49382), .ZN(n49336) );
  INV_X1 U15522 ( .I(n10716), .ZN(n15967) );
  OR2_X1 U15523 ( .A1(n23738), .A2(n49006), .Z(n48321) );
  NAND2_X1 U15524 ( .A1(n48707), .A2(n20911), .ZN(n48710) );
  INV_X1 U15526 ( .I(n63943), .ZN(n48675) );
  NAND2_X1 U15528 ( .A1(n49356), .A2(n50044), .ZN(n8457) );
  NAND2_X1 U15529 ( .A1(n12966), .A2(n63943), .ZN(n48673) );
  NOR2_X1 U15534 ( .A1(n18769), .A2(n49430), .ZN(n11002) );
  OAI21_X1 U15538 ( .A1(n3772), .A2(n58269), .B(n58206), .ZN(n45607) );
  NAND2_X1 U15539 ( .A1(n49091), .A2(n16922), .ZN(n2629) );
  NAND2_X1 U15540 ( .A1(n60719), .A2(n49739), .ZN(n49740) );
  NOR2_X1 U15541 ( .A1(n6203), .A2(n5345), .ZN(n23721) );
  INV_X1 U15543 ( .I(n49699), .ZN(n6930) );
  INV_X1 U15550 ( .I(n48822), .ZN(n48821) );
  OR2_X1 U15551 ( .A1(n49846), .A2(n49845), .Z(n49857) );
  NAND3_X1 U15553 ( .A1(n49116), .A2(n47947), .A3(n13878), .ZN(n47349) );
  NAND2_X1 U15555 ( .A1(n4017), .A2(n21550), .ZN(n4827) );
  INV_X1 U15556 ( .I(n49152), .ZN(n49227) );
  AOI21_X1 U15557 ( .A1(n49222), .A2(n10831), .B(n49221), .ZN(n49223) );
  NOR2_X1 U15559 ( .A1(n2262), .A2(n7587), .ZN(n12474) );
  INV_X1 U15560 ( .I(n48774), .ZN(n48924) );
  INV_X1 U15561 ( .I(n49307), .ZN(n48996) );
  NAND2_X1 U15562 ( .A1(n2543), .A2(n49684), .ZN(n2542) );
  INV_X2 U15566 ( .I(n13878), .ZN(n49804) );
  OR4_X1 U15567 ( .A1(n63084), .A2(n50079), .A3(n50403), .A4(n1381), .Z(n49422) );
  NOR2_X1 U15568 ( .A1(n49655), .A2(n14047), .ZN(n49656) );
  AND2_X1 U15570 ( .A1(n50410), .A2(n50411), .Z(n15837) );
  NAND2_X1 U15572 ( .A1(n50310), .A2(n50313), .ZN(n8740) );
  NAND2_X1 U15573 ( .A1(n48268), .A2(n50000), .ZN(n4391) );
  NAND2_X1 U15574 ( .A1(n4098), .A2(n21550), .ZN(n46087) );
  NAND3_X1 U15576 ( .A1(n19998), .A2(n8129), .A3(n59086), .ZN(n47446) );
  NAND2_X1 U15579 ( .A1(n49406), .A2(n10874), .ZN(n2382) );
  INV_X1 U15580 ( .I(n49608), .ZN(n48704) );
  NAND2_X1 U15584 ( .A1(n5497), .A2(n49372), .ZN(n4452) );
  NAND2_X1 U15585 ( .A1(n49373), .A2(n2582), .ZN(n2581) );
  NOR2_X1 U15589 ( .A1(n48073), .A2(n19294), .ZN(n12368) );
  NOR2_X1 U15590 ( .A1(n21334), .A2(n20458), .ZN(n21333) );
  INV_X1 U15592 ( .I(n49561), .ZN(n48279) );
  INV_X4 U15593 ( .I(n20811), .ZN(n48688) );
  AOI21_X1 U15596 ( .A1(n47449), .A2(n7990), .B(n1468), .ZN(n45703) );
  INV_X1 U15597 ( .I(n48897), .ZN(n49760) );
  NAND2_X1 U15604 ( .A1(n49631), .A2(n16197), .ZN(n15356) );
  INV_X1 U15606 ( .I(n12966), .ZN(n48938) );
  AND2_X1 U15607 ( .A1(n49055), .A2(n3971), .Z(n47922) );
  AND2_X1 U15608 ( .A1(n49277), .A2(n49281), .Z(n16862) );
  INV_X1 U15613 ( .I(n49922), .ZN(n2981) );
  NAND3_X1 U15615 ( .A1(n24362), .A2(n60772), .A3(n49635), .ZN(n49633) );
  OR2_X1 U15616 ( .A1(n49496), .A2(n22780), .Z(n5591) );
  NAND2_X1 U15621 ( .A1(n50394), .A2(n4172), .ZN(n50403) );
  INV_X1 U15623 ( .I(n49642), .ZN(n48726) );
  INV_X1 U15625 ( .I(n49752), .ZN(n6203) );
  NAND2_X1 U15627 ( .A1(n50143), .A2(n50307), .ZN(n25113) );
  NAND3_X1 U15628 ( .A1(n16197), .A2(n60772), .A3(n47334), .ZN(n47335) );
  AOI21_X1 U15630 ( .A1(n50220), .A2(n14931), .B(n14516), .ZN(n8355) );
  NOR2_X1 U15631 ( .A1(n14931), .A2(n7586), .ZN(n49338) );
  INV_X1 U15632 ( .I(n50222), .ZN(n50208) );
  NAND2_X1 U15633 ( .A1(n8129), .A2(n25032), .ZN(n20864) );
  NOR2_X1 U15635 ( .A1(n9409), .A2(n50376), .ZN(n50380) );
  NOR2_X1 U15636 ( .A1(n24583), .A2(n1473), .ZN(n24582) );
  OR2_X1 U15637 ( .A1(n64341), .A2(n12701), .Z(n48697) );
  INV_X1 U15638 ( .I(n21367), .ZN(n6897) );
  NOR2_X1 U15639 ( .A1(n49410), .A2(n5545), .ZN(n5544) );
  NOR2_X1 U15640 ( .A1(n49090), .A2(n49677), .ZN(n5429) );
  INV_X1 U15641 ( .I(n15635), .ZN(n15634) );
  NAND2_X1 U15642 ( .A1(n19003), .A2(n49610), .ZN(n10760) );
  INV_X1 U15643 ( .I(n3281), .ZN(n25744) );
  INV_X1 U15644 ( .I(n50267), .ZN(n15194) );
  NAND2_X1 U15645 ( .A1(n49674), .A2(n17906), .ZN(n49366) );
  NOR2_X1 U15646 ( .A1(n1382), .A2(n7358), .ZN(n2245) );
  AOI21_X1 U15648 ( .A1(n1384), .A2(n21092), .B(n1471), .ZN(n46778) );
  NAND2_X1 U15650 ( .A1(n49926), .A2(n48727), .ZN(n48730) );
  AND2_X1 U15651 ( .A1(n50374), .A2(n23650), .Z(n12626) );
  NAND2_X1 U15652 ( .A1(n19705), .A2(n1640), .ZN(n11289) );
  INV_X1 U15653 ( .I(n49885), .ZN(n49889) );
  INV_X2 U15658 ( .I(n50238), .ZN(n1632) );
  NAND2_X1 U15659 ( .A1(n50044), .A2(n50041), .ZN(n50047) );
  INV_X1 U15663 ( .I(n49150), .ZN(n3239) );
  AND2_X1 U15665 ( .A1(n19773), .A2(n50044), .Z(n16256) );
  NOR2_X1 U15667 ( .A1(n49655), .A2(n50296), .ZN(n18158) );
  INV_X1 U15668 ( .I(n50117), .ZN(n49887) );
  NAND2_X1 U15670 ( .A1(n17885), .A2(n23299), .ZN(n50240) );
  OR2_X1 U15672 ( .A1(n3335), .A2(n19773), .Z(n14168) );
  CLKBUF_X2 U15673 ( .I(n22959), .Z(n10015) );
  AND2_X1 U15674 ( .A1(n19144), .A2(n19634), .Z(n16211) );
  OR2_X1 U15677 ( .A1(n57194), .A2(n49276), .Z(n16084) );
  BUF_X4 U15679 ( .I(n23839), .Z(n18882) );
  NAND2_X1 U15681 ( .A1(n22571), .A2(n49166), .ZN(n15349) );
  NOR2_X1 U15682 ( .A1(n49377), .A2(n49538), .ZN(n23576) );
  INV_X1 U15690 ( .I(n10030), .ZN(n3237) );
  CLKBUF_X2 U15692 ( .I(n50331), .Z(n4594) );
  BUF_X4 U15694 ( .I(n49630), .Z(n3658) );
  NAND2_X1 U15695 ( .A1(n25944), .A2(n50394), .ZN(n8995) );
  CLKBUF_X2 U15699 ( .I(n48411), .Z(n7115) );
  BUF_X2 U15712 ( .I(n11795), .Z(n11314) );
  CLKBUF_X2 U15714 ( .I(n49043), .Z(n12579) );
  OR2_X1 U15718 ( .A1(n49459), .A2(n6314), .Z(n16381) );
  INV_X1 U15728 ( .I(n11490), .ZN(n13396) );
  NOR2_X1 U15731 ( .A1(n25457), .A2(n16200), .ZN(n48818) );
  INV_X1 U15734 ( .I(n46047), .ZN(n4271) );
  NAND2_X1 U15736 ( .A1(n16415), .A2(n3249), .ZN(n16414) );
  NAND2_X1 U15737 ( .A1(n15265), .A2(n25899), .ZN(n6732) );
  NAND2_X1 U15741 ( .A1(n47117), .A2(n47116), .ZN(n3096) );
  NAND2_X1 U15746 ( .A1(n14775), .A2(n47372), .ZN(n9816) );
  OAI21_X1 U15750 ( .A1(n6289), .A2(n45777), .B(n45776), .ZN(n6288) );
  NAND2_X1 U15751 ( .A1(n24952), .A2(n24708), .ZN(n23620) );
  NAND2_X1 U15762 ( .A1(n21556), .A2(n21557), .ZN(n21555) );
  NOR2_X1 U15764 ( .A1(n17209), .A2(n17207), .ZN(n17206) );
  NOR2_X1 U15768 ( .A1(n26175), .A2(n44945), .ZN(n25361) );
  NOR2_X1 U15774 ( .A1(n47662), .A2(n47661), .ZN(n24395) );
  AOI21_X1 U15780 ( .A1(n4380), .A2(n46990), .B(n20655), .ZN(n20654) );
  AOI22_X1 U15787 ( .A1(n46924), .A2(n3203), .B1(n46922), .B2(n46923), .ZN(
        n46934) );
  OAI22_X1 U15788 ( .A1(n13821), .A2(n25006), .B1(n47401), .B2(n18227), .ZN(
        n13828) );
  NAND2_X1 U15792 ( .A1(n14691), .A2(n14690), .ZN(n14689) );
  NAND2_X1 U15793 ( .A1(n45974), .A2(n24208), .ZN(n10530) );
  NOR2_X1 U15795 ( .A1(n9934), .A2(n46266), .ZN(n9740) );
  INV_X1 U15797 ( .I(n45771), .ZN(n6280) );
  NOR2_X1 U15798 ( .A1(n48634), .A2(n48633), .ZN(n48638) );
  INV_X1 U15799 ( .I(n45763), .ZN(n6283) );
  INV_X1 U15800 ( .I(n17081), .ZN(n17080) );
  NOR2_X1 U15803 ( .A1(n13933), .A2(n13932), .ZN(n13931) );
  INV_X1 U15805 ( .I(n45773), .ZN(n6289) );
  NAND2_X1 U15807 ( .A1(n17771), .A2(n47111), .ZN(n17770) );
  NAND2_X1 U15811 ( .A1(n45667), .A2(n26240), .ZN(n25003) );
  OAI21_X1 U15812 ( .A1(n4773), .A2(n15835), .B(n48594), .ZN(n12329) );
  OAI21_X1 U15813 ( .A1(n46067), .A2(n60504), .B(n46066), .ZN(n21556) );
  NAND2_X1 U15817 ( .A1(n47203), .A2(n12487), .ZN(n12486) );
  NAND2_X1 U15821 ( .A1(n16703), .A2(n48247), .ZN(n3360) );
  NAND2_X1 U15823 ( .A1(n14695), .A2(n1074), .ZN(n14694) );
  AOI21_X1 U15824 ( .A1(n6786), .A2(n64960), .B(n6657), .ZN(n6656) );
  NAND2_X1 U15826 ( .A1(n11294), .A2(n11295), .ZN(n11292) );
  NAND2_X1 U15833 ( .A1(n47363), .A2(n47366), .ZN(n25033) );
  INV_X1 U15837 ( .I(n47413), .ZN(n13498) );
  NAND2_X1 U15839 ( .A1(n48582), .A2(n11025), .ZN(n46477) );
  NAND2_X1 U15842 ( .A1(n46809), .A2(n2955), .ZN(n14787) );
  OAI21_X1 U15844 ( .A1(n47379), .A2(n12498), .B(n47378), .ZN(n10508) );
  NAND2_X1 U15846 ( .A1(n48094), .A2(n62755), .ZN(n11097) );
  NOR2_X1 U15847 ( .A1(n47638), .A2(n15030), .ZN(n47639) );
  NAND2_X1 U15848 ( .A1(n7367), .A2(n47718), .ZN(n43599) );
  NOR2_X1 U15849 ( .A1(n11900), .A2(n11899), .ZN(n11898) );
  INV_X1 U15850 ( .I(n47365), .ZN(n11897) );
  NOR2_X1 U15851 ( .A1(n11908), .A2(n11904), .ZN(n11903) );
  AND3_X1 U15853 ( .A1(n45535), .A2(n45534), .A3(n45533), .Z(n45543) );
  AOI21_X1 U15854 ( .A1(n17083), .A2(n8507), .B(n17082), .ZN(n17081) );
  INV_X1 U15855 ( .I(n12619), .ZN(n12618) );
  OAI21_X1 U15857 ( .A1(n1476), .A2(n13433), .B(n13432), .ZN(n13933) );
  NAND2_X1 U15858 ( .A1(n45083), .A2(n45082), .ZN(n24452) );
  NAND2_X1 U15862 ( .A1(n14575), .A2(n47139), .ZN(n14574) );
  OAI21_X1 U15864 ( .A1(n16702), .A2(n209), .B(n13759), .ZN(n3468) );
  NOR2_X1 U15865 ( .A1(n45695), .A2(n14911), .ZN(n45697) );
  AOI21_X1 U15867 ( .A1(n46784), .A2(n10250), .B(n46783), .ZN(n46785) );
  AND2_X1 U15870 ( .A1(n47202), .A2(n18787), .Z(n12483) );
  AOI21_X1 U15871 ( .A1(n46845), .A2(n47682), .B(n20568), .ZN(n20567) );
  INV_X1 U15872 ( .I(n47112), .ZN(n47111) );
  NAND2_X1 U15876 ( .A1(n15417), .A2(n45455), .ZN(n2756) );
  AOI22_X1 U15878 ( .A1(n12069), .A2(n20005), .B1(n12024), .B2(n47418), .ZN(
        n12076) );
  OAI21_X1 U15880 ( .A1(n11627), .A2(n20912), .B(n13822), .ZN(n13821) );
  NAND2_X1 U15887 ( .A1(n20831), .A2(n20830), .ZN(n46067) );
  OAI21_X1 U15890 ( .A1(n14569), .A2(n47373), .B(n7218), .ZN(n14568) );
  NAND2_X1 U15891 ( .A1(n47105), .A2(n47104), .ZN(n10437) );
  OR2_X1 U15892 ( .A1(n10450), .A2(n13413), .Z(n15424) );
  NOR2_X1 U15894 ( .A1(n4214), .A2(n3640), .ZN(n16224) );
  NAND3_X1 U15896 ( .A1(n47313), .A2(n47307), .A3(n59687), .ZN(n46920) );
  INV_X1 U15897 ( .I(n3181), .ZN(n46924) );
  NAND2_X1 U15898 ( .A1(n47120), .A2(n60651), .ZN(n10328) );
  NAND2_X1 U15899 ( .A1(n17210), .A2(n12722), .ZN(n17209) );
  NOR2_X1 U15901 ( .A1(n47485), .A2(n47484), .ZN(n13041) );
  OAI21_X1 U15903 ( .A1(n22243), .A2(n47824), .B(n47609), .ZN(n45974) );
  INV_X1 U15904 ( .I(n45971), .ZN(n24208) );
  OAI21_X1 U15908 ( .A1(n47667), .A2(n47668), .B(n21951), .ZN(n19605) );
  NOR2_X1 U15911 ( .A1(n9199), .A2(n2827), .ZN(n20655) );
  NAND2_X1 U15912 ( .A1(n1086), .A2(n11296), .ZN(n11295) );
  OAI22_X1 U15913 ( .A1(n12709), .A2(n12708), .B1(n47001), .B2(n47484), .ZN(
        n25791) );
  NAND3_X1 U15914 ( .A1(n45952), .A2(n12114), .A3(n3181), .ZN(n20268) );
  INV_X1 U15916 ( .I(n46481), .ZN(n5202) );
  NOR2_X1 U15917 ( .A1(n3615), .A2(n45448), .ZN(n3599) );
  AND3_X1 U15921 ( .A1(n47673), .A2(n47672), .A3(n47853), .Z(n47677) );
  NOR2_X1 U15922 ( .A1(n47566), .A2(n24380), .ZN(n18107) );
  OAI22_X1 U15923 ( .A1(n45979), .A2(n47281), .B1(n47275), .B2(n47593), .ZN(
        n45677) );
  NAND2_X1 U15925 ( .A1(n18787), .A2(n63913), .ZN(n7504) );
  NAND2_X1 U15929 ( .A1(n1080), .A2(n45503), .ZN(n6657) );
  NAND2_X1 U15930 ( .A1(n18981), .A2(n18980), .ZN(n18979) );
  OAI21_X1 U15931 ( .A1(n24313), .A2(n57731), .B(n1070), .ZN(n17023) );
  NAND2_X1 U15932 ( .A1(n49863), .A2(n49862), .ZN(n14438) );
  AND2_X1 U15933 ( .A1(n7222), .A2(n47297), .Z(n7077) );
  INV_X1 U15936 ( .I(n48098), .ZN(n48099) );
  INV_X1 U15937 ( .I(n10463), .ZN(n44400) );
  NAND2_X1 U15939 ( .A1(n47492), .A2(n48667), .ZN(n14695) );
  INV_X1 U15941 ( .I(n1064), .ZN(n47047) );
  AOI22_X1 U15942 ( .A1(n14456), .A2(n14741), .B1(n47831), .B2(n14454), .ZN(
        n24380) );
  INV_X1 U15943 ( .I(n44674), .ZN(n47046) );
  NAND2_X1 U15944 ( .A1(n21548), .A2(n21547), .ZN(n48486) );
  NOR2_X1 U15945 ( .A1(n47044), .A2(n61980), .ZN(n17809) );
  INV_X1 U15946 ( .I(n47145), .ZN(n14567) );
  NAND2_X1 U15947 ( .A1(n47396), .A2(n45906), .ZN(n14030) );
  NOR2_X1 U15948 ( .A1(n23865), .A2(n48654), .ZN(n4623) );
  NAND2_X1 U15949 ( .A1(n8224), .A2(n47839), .ZN(n11928) );
  INV_X1 U15953 ( .I(n48535), .ZN(n13267) );
  NOR2_X1 U15954 ( .A1(n48558), .A2(n48557), .ZN(n48570) );
  AOI21_X1 U15955 ( .A1(n48110), .A2(n48111), .B(n48109), .ZN(n14437) );
  NOR2_X1 U15956 ( .A1(n18498), .A2(n16533), .ZN(n14693) );
  INV_X1 U15958 ( .I(n11297), .ZN(n11296) );
  NOR2_X1 U15959 ( .A1(n44771), .A2(n16077), .ZN(n16413) );
  NOR2_X1 U15961 ( .A1(n1328), .A2(n46950), .ZN(n5979) );
  INV_X1 U15962 ( .I(n44771), .ZN(n46108) );
  NAND2_X1 U15963 ( .A1(n18974), .A2(n18973), .ZN(n18981) );
  OAI22_X1 U15965 ( .A1(n47294), .A2(n47295), .B1(n3641), .B2(n47296), .ZN(
        n7222) );
  NAND2_X1 U15966 ( .A1(n46760), .A2(n65062), .ZN(n3094) );
  NAND2_X1 U15968 ( .A1(n20140), .A2(n62230), .ZN(n21638) );
  INV_X1 U15971 ( .I(n16438), .ZN(n7218) );
  NOR2_X1 U15973 ( .A1(n48113), .A2(n57728), .ZN(n15164) );
  NOR2_X1 U15974 ( .A1(n59687), .A2(n5297), .ZN(n46926) );
  NAND2_X1 U15975 ( .A1(n47469), .A2(n46977), .ZN(n9173) );
  OAI21_X1 U15976 ( .A1(n15419), .A2(n15418), .B(n18980), .ZN(n15417) );
  INV_X1 U15978 ( .I(n47671), .ZN(n47672) );
  INV_X1 U15979 ( .I(n46050), .ZN(n6431) );
  AND3_X1 U15981 ( .A1(n47228), .A2(n47229), .A3(n18196), .Z(n46056) );
  NAND2_X1 U15982 ( .A1(n48102), .A2(n20140), .ZN(n45804) );
  INV_X1 U15983 ( .I(n4261), .ZN(n4260) );
  NOR2_X1 U15984 ( .A1(n23361), .A2(n2916), .ZN(n2915) );
  NAND2_X1 U15985 ( .A1(n45488), .A2(n45485), .ZN(n19229) );
  NAND2_X1 U15987 ( .A1(n47441), .A2(n47442), .ZN(n8130) );
  AOI21_X1 U15988 ( .A1(n46925), .A2(n47307), .B(n6935), .ZN(n45083) );
  NOR2_X1 U15990 ( .A1(n10978), .A2(n10977), .ZN(n10975) );
  INV_X1 U15991 ( .I(n45182), .ZN(n7367) );
  NAND2_X1 U15992 ( .A1(n21200), .A2(n47690), .ZN(n21199) );
  NOR2_X1 U15995 ( .A1(n45539), .A2(n11062), .ZN(n45540) );
  NAND2_X1 U15997 ( .A1(n6599), .A2(n59892), .ZN(n45767) );
  NAND2_X1 U15998 ( .A1(n48660), .A2(n48650), .ZN(n13432) );
  NAND2_X1 U15999 ( .A1(n16068), .A2(n1475), .ZN(n13965) );
  OAI21_X1 U16002 ( .A1(n8508), .A2(n23263), .B(n48641), .ZN(n8507) );
  OR2_X1 U16003 ( .A1(n1263), .A2(n47425), .Z(n10763) );
  AOI21_X1 U16004 ( .A1(n45960), .A2(n45966), .B(n3510), .ZN(n22243) );
  NAND2_X1 U16006 ( .A1(n6903), .A2(n48224), .ZN(n46361) );
  NAND2_X1 U16008 ( .A1(n7318), .A2(n8666), .ZN(n47004) );
  AND2_X1 U16009 ( .A1(n47620), .A2(n47619), .Z(n47629) );
  AND3_X1 U16011 ( .A1(n46264), .A2(n46263), .A3(n61146), .Z(n46266) );
  NOR2_X1 U16019 ( .A1(n47807), .A2(n47809), .ZN(n5309) );
  NOR2_X1 U16020 ( .A1(n18992), .A2(n8574), .ZN(n8573) );
  AND3_X1 U16021 ( .A1(n47625), .A2(n62739), .A3(n15360), .Z(n16036) );
  NAND3_X1 U16022 ( .A1(n11744), .A2(n48619), .A3(n22635), .ZN(n11743) );
  AOI21_X1 U16023 ( .A1(n43828), .A2(n6730), .B(n47674), .ZN(n4091) );
  OAI21_X1 U16024 ( .A1(n45206), .A2(n47616), .B(n45205), .ZN(n19737) );
  NAND2_X1 U16026 ( .A1(n61601), .A2(n22239), .ZN(n45578) );
  OAI21_X1 U16027 ( .A1(n48165), .A2(n12990), .B(n48507), .ZN(n12989) );
  OAI21_X1 U16028 ( .A1(n6933), .A2(n7799), .B(n46921), .ZN(n46922) );
  OR2_X1 U16029 ( .A1(n46985), .A2(n19989), .Z(n19988) );
  NAND2_X1 U16031 ( .A1(n45670), .A2(n46882), .ZN(n13446) );
  NAND3_X1 U16032 ( .A1(n47727), .A2(n47880), .A3(n47878), .ZN(n9332) );
  NAND2_X1 U16033 ( .A1(n47399), .A2(n45446), .ZN(n3614) );
  NOR2_X1 U16034 ( .A1(n2169), .A2(n20162), .ZN(n47485) );
  INV_X1 U16035 ( .I(n46069), .ZN(n6788) );
  NAND2_X1 U16038 ( .A1(n47226), .A2(n24340), .ZN(n3081) );
  AOI22_X1 U16039 ( .A1(n46804), .A2(n2499), .B1(n9045), .B2(n48464), .ZN(
        n46805) );
  NAND2_X1 U16040 ( .A1(n46749), .A2(n47381), .ZN(n14575) );
  INV_X1 U16042 ( .I(n45670), .ZN(n46887) );
  NAND2_X1 U16043 ( .A1(n15994), .A2(n44703), .ZN(n18319) );
  NAND2_X1 U16044 ( .A1(n46806), .A2(n46807), .ZN(n24430) );
  OAI21_X1 U16045 ( .A1(n47176), .A2(n47544), .B(n22704), .ZN(n24988) );
  NAND2_X1 U16046 ( .A1(n18321), .A2(n44705), .ZN(n44572) );
  INV_X1 U16047 ( .I(n8643), .ZN(n8648) );
  NAND2_X1 U16048 ( .A1(n8651), .A2(n47237), .ZN(n8646) );
  AOI21_X1 U16049 ( .A1(n45007), .A2(n45006), .B(n7296), .ZN(n14417) );
  AOI21_X1 U16052 ( .A1(n47984), .A2(n47985), .B(n18196), .ZN(n47988) );
  NAND2_X1 U16053 ( .A1(n45445), .A2(n13782), .ZN(n3598) );
  AOI21_X1 U16054 ( .A1(n16074), .A2(n47037), .B(n21712), .ZN(n10463) );
  NAND2_X1 U16055 ( .A1(n45456), .A2(n15421), .ZN(n15420) );
  NAND2_X1 U16058 ( .A1(n11214), .A2(n45985), .ZN(n14414) );
  NAND2_X1 U16059 ( .A1(n47201), .A2(n48191), .ZN(n12487) );
  NAND2_X1 U16060 ( .A1(n5934), .A2(n46894), .ZN(n17210) );
  INV_X1 U16066 ( .I(n48639), .ZN(n8508) );
  AOI22_X1 U16067 ( .A1(n1086), .A2(n47516), .B1(n11786), .B2(n47495), .ZN(
        n47496) );
  INV_X1 U16068 ( .I(n46942), .ZN(n46940) );
  AND2_X1 U16069 ( .A1(n1082), .A2(n48659), .Z(n16190) );
  NAND2_X1 U16070 ( .A1(n3080), .A2(n12249), .ZN(n47226) );
  NAND2_X1 U16071 ( .A1(n63953), .A2(n45493), .ZN(n44343) );
  NAND2_X1 U16073 ( .A1(n48662), .A2(n209), .ZN(n13433) );
  NOR2_X1 U16074 ( .A1(n1667), .A2(n2170), .ZN(n2169) );
  NOR2_X1 U16075 ( .A1(n45536), .A2(n21712), .ZN(n15994) );
  NAND2_X1 U16076 ( .A1(n48588), .A2(n8758), .ZN(n48589) );
  AOI21_X1 U16077 ( .A1(n25026), .A2(n47874), .B(n12647), .ZN(n8924) );
  NOR2_X1 U16081 ( .A1(n45669), .A2(n46885), .ZN(n21803) );
  NAND2_X1 U16084 ( .A1(n47853), .A2(n61909), .ZN(n18265) );
  NOR2_X1 U16085 ( .A1(n12648), .A2(n47880), .ZN(n2250) );
  NAND3_X1 U16089 ( .A1(n4315), .A2(n63734), .A3(n46078), .ZN(n46079) );
  INV_X2 U16095 ( .I(n48567), .ZN(n47123) );
  INV_X1 U16096 ( .I(n46790), .ZN(n21198) );
  OAI22_X1 U16098 ( .A1(n25480), .A2(n48624), .B1(n571), .B2(n22635), .ZN(
        n21567) );
  NAND2_X1 U16100 ( .A1(n48629), .A2(n48615), .ZN(n15145) );
  INV_X1 U16101 ( .I(n47420), .ZN(n12025) );
  INV_X1 U16102 ( .I(n47682), .ZN(n20005) );
  INV_X1 U16103 ( .I(n11492), .ZN(n6194) );
  NOR2_X1 U16104 ( .A1(n46875), .A2(n45491), .ZN(n13729) );
  NAND2_X1 U16107 ( .A1(n1385), .A2(n47806), .ZN(n47807) );
  INV_X1 U16108 ( .I(n46737), .ZN(n46740) );
  INV_X1 U16109 ( .I(n48209), .ZN(n48210) );
  NAND3_X1 U16111 ( .A1(n24820), .A2(n5771), .A3(n47530), .ZN(n12227) );
  INV_X1 U16114 ( .I(n45674), .ZN(n44872) );
  AND2_X1 U16115 ( .A1(n8758), .A2(n9851), .Z(n11025) );
  AND2_X1 U16116 ( .A1(n57852), .A2(n263), .Z(n16296) );
  NOR2_X1 U16117 ( .A1(n47299), .A2(n47298), .ZN(n7235) );
  OR2_X1 U16118 ( .A1(n47119), .A2(n48559), .Z(n47120) );
  AND2_X1 U16119 ( .A1(n45696), .A2(n18196), .Z(n14911) );
  NOR2_X1 U16120 ( .A1(n48562), .A2(n60848), .ZN(n9794) );
  OAI22_X1 U16121 ( .A1(n47243), .A2(n45576), .B1(n60979), .B2(n45988), .ZN(
        n45008) );
  OAI22_X1 U16122 ( .A1(n48640), .A2(n48162), .B1(n64791), .B2(n48642), .ZN(
        n46562) );
  INV_X1 U16125 ( .I(n12993), .ZN(n48164) );
  INV_X1 U16126 ( .I(n17805), .ZN(n12709) );
  OR2_X1 U16127 ( .A1(n17318), .A2(n48659), .Z(n12708) );
  NAND2_X1 U16130 ( .A1(n8200), .A2(n48481), .ZN(n8199) );
  AND2_X1 U16131 ( .A1(n47434), .A2(n62788), .Z(n47443) );
  AOI22_X1 U16132 ( .A1(n20111), .A2(n47380), .B1(n23718), .B2(n10172), .ZN(
        n10675) );
  OR2_X1 U16134 ( .A1(n47251), .A2(n47259), .Z(n45668) );
  INV_X1 U16135 ( .I(n46893), .ZN(n15566) );
  NAND2_X1 U16141 ( .A1(n48239), .A2(n48234), .ZN(n19557) );
  AOI21_X1 U16142 ( .A1(n5532), .A2(n47565), .B(n5465), .ZN(n5464) );
  INV_X1 U16143 ( .I(n25480), .ZN(n6903) );
  AND2_X1 U16145 ( .A1(n21719), .A2(n21718), .Z(n47095) );
  NAND2_X1 U16146 ( .A1(n21689), .A2(n48166), .ZN(n12990) );
  NAND2_X1 U16148 ( .A1(n45794), .A2(n47411), .ZN(n45796) );
  NAND2_X1 U16149 ( .A1(n16493), .A2(n1480), .ZN(n46263) );
  NOR2_X1 U16152 ( .A1(n47874), .A2(n64548), .ZN(n11906) );
  NAND2_X1 U16154 ( .A1(n3105), .A2(n1479), .ZN(n3287) );
  NOR2_X1 U16155 ( .A1(n59821), .A2(n46913), .ZN(n24313) );
  NOR2_X1 U16156 ( .A1(n47110), .A2(n12698), .ZN(n47113) );
  NAND2_X1 U16158 ( .A1(n45966), .A2(n47605), .ZN(n18911) );
  NAND2_X1 U16159 ( .A1(n21689), .A2(n16286), .ZN(n12997) );
  NOR2_X1 U16160 ( .A1(n23185), .A2(n20340), .ZN(n48548) );
  NAND2_X1 U16161 ( .A1(n47209), .A2(n5090), .ZN(n47092) );
  OR2_X1 U16163 ( .A1(n10397), .A2(n57740), .Z(n11628) );
  NOR2_X1 U16165 ( .A1(n4090), .A2(n47367), .ZN(n46826) );
  INV_X1 U16166 ( .I(n63853), .ZN(n21712) );
  AND2_X1 U16168 ( .A1(n45957), .A2(n47329), .Z(n45951) );
  AND2_X1 U16169 ( .A1(n47729), .A2(n47728), .Z(n15919) );
  OR2_X1 U16170 ( .A1(n48518), .A2(n48514), .Z(n16286) );
  NAND2_X1 U16171 ( .A1(n48511), .A2(n23263), .ZN(n48496) );
  NAND2_X1 U16172 ( .A1(n22635), .A2(n25482), .ZN(n46358) );
  NAND2_X1 U16175 ( .A1(n48624), .A2(n47542), .ZN(n47165) );
  AND2_X1 U16176 ( .A1(n46951), .A2(n64960), .Z(n16225) );
  INV_X1 U16177 ( .I(n47261), .ZN(n15567) );
  AND2_X1 U16178 ( .A1(n47529), .A2(n62115), .Z(n15835) );
  NAND2_X1 U16179 ( .A1(n3203), .A2(n46919), .ZN(n46060) );
  NOR2_X1 U16180 ( .A1(n47316), .A2(n47307), .ZN(n8270) );
  NAND2_X1 U16181 ( .A1(n47174), .A2(n571), .ZN(n46365) );
  INV_X1 U16188 ( .I(n47247), .ZN(n45669) );
  NOR2_X1 U16189 ( .A1(n48624), .A2(n14419), .ZN(n46463) );
  AND2_X1 U16190 ( .A1(n838), .A2(n15157), .Z(n14454) );
  AND2_X1 U16192 ( .A1(n64042), .A2(n47838), .Z(n47560) );
  INV_X1 U16195 ( .I(n5090), .ZN(n47083) );
  OAI21_X1 U16197 ( .A1(n48620), .A2(n14419), .B(n3341), .ZN(n48225) );
  CLKBUF_X2 U16198 ( .I(n47156), .Z(n9851) );
  NAND2_X1 U16199 ( .A1(n1085), .A2(n1483), .ZN(n44864) );
  NOR2_X1 U16200 ( .A1(n4214), .A2(n25477), .ZN(n2150) );
  NOR2_X1 U16202 ( .A1(n3367), .A2(n3366), .ZN(n46102) );
  NAND2_X1 U16206 ( .A1(n3368), .A2(n8152), .ZN(n8155) );
  NAND2_X1 U16208 ( .A1(n47180), .A2(n571), .ZN(n48613) );
  AND2_X1 U16209 ( .A1(n48614), .A2(n48620), .Z(n15324) );
  NAND2_X1 U16210 ( .A1(n8639), .A2(n3341), .ZN(n48610) );
  NAND2_X1 U16212 ( .A1(n8639), .A2(n14418), .ZN(n47169) );
  NAND2_X1 U16213 ( .A1(n47593), .A2(n23186), .ZN(n3637) );
  NOR2_X1 U16215 ( .A1(n47736), .A2(n59008), .ZN(n5132) );
  OAI21_X1 U16216 ( .A1(n47735), .A2(n62788), .B(n63647), .ZN(n47436) );
  NAND3_X1 U16217 ( .A1(n15360), .A2(n47244), .A3(n47623), .ZN(n45577) );
  AOI21_X1 U16218 ( .A1(n47381), .A2(n23934), .B(n20112), .ZN(n20111) );
  AND2_X2 U16219 ( .A1(n5803), .A2(n5265), .Z(n3686) );
  NOR2_X1 U16220 ( .A1(n47502), .A2(n9331), .ZN(n17808) );
  NOR2_X1 U16221 ( .A1(n47437), .A2(n63647), .ZN(n15418) );
  AND2_X1 U16222 ( .A1(n47487), .A2(n62853), .Z(n16077) );
  OR2_X1 U16225 ( .A1(n48085), .A2(n11708), .Z(n10979) );
  AND2_X1 U16226 ( .A1(n23894), .A2(n61025), .Z(n16068) );
  AND2_X1 U16227 ( .A1(n64548), .A2(n47876), .Z(n14120) );
  OR2_X1 U16228 ( .A1(n48543), .A2(n57973), .Z(n16012) );
  AOI21_X1 U16229 ( .A1(n47240), .A2(n60979), .B(n47239), .ZN(n47241) );
  AOI22_X1 U16230 ( .A1(n47565), .A2(n5554), .B1(n47834), .B2(n47830), .ZN(
        n16375) );
  INV_X1 U16232 ( .I(n46027), .ZN(n6247) );
  AND2_X1 U16234 ( .A1(n19040), .A2(n48654), .Z(n47001) );
  NAND2_X1 U16235 ( .A1(n6957), .A2(n44770), .ZN(n2170) );
  INV_X2 U16236 ( .I(n46944), .ZN(n47233) );
  CLKBUF_X2 U16238 ( .I(n45075), .Z(n47309) );
  NAND3_X1 U16240 ( .A1(n47274), .A2(n45551), .A3(n47270), .ZN(n3638) );
  CLKBUF_X2 U16243 ( .I(n15824), .Z(n10627) );
  INV_X2 U16244 ( .I(n21452), .ZN(n47252) );
  INV_X1 U16246 ( .I(n47251), .ZN(n4315) );
  AND2_X2 U16248 ( .A1(n46244), .A2(n10364), .Z(n18570) );
  INV_X2 U16254 ( .I(n14929), .ZN(n47156) );
  NAND2_X1 U16256 ( .A1(n6497), .A2(n47985), .ZN(n6645) );
  AND2_X1 U16261 ( .A1(n1267), .A2(n46913), .Z(n6290) );
  INV_X1 U16262 ( .I(n48560), .ZN(n24113) );
  INV_X1 U16263 ( .I(n10475), .ZN(n16486) );
  INV_X1 U16265 ( .I(n65275), .ZN(n47499) );
  NOR2_X1 U16266 ( .A1(n64888), .A2(n45718), .ZN(n13728) );
  BUF_X2 U16268 ( .I(n46244), .Z(n48667) );
  CLKBUF_X2 U16272 ( .I(n47832), .Z(n10420) );
  INV_X1 U16276 ( .I(n9860), .ZN(n22536) );
  CLKBUF_X2 U16277 ( .I(n45191), .Z(n23167) );
  CLKBUF_X2 U16279 ( .I(n43748), .Z(n47730) );
  CLKBUF_X2 U16280 ( .I(n46262), .Z(n23035) );
  CLKBUF_X2 U16282 ( .I(n45520), .Z(n20917) );
  INV_X2 U16288 ( .I(n15823), .ZN(n46770) );
  BUF_X2 U16295 ( .I(n46513), .Z(n48642) );
  INV_X1 U16297 ( .I(n44670), .ZN(n3271) );
  CLKBUF_X2 U16300 ( .I(n14888), .Z(n22908) );
  INV_X1 U16303 ( .I(n44294), .ZN(n5663) );
  CLKBUF_X2 U16304 ( .I(n25166), .Z(n47838) );
  INV_X2 U16306 ( .I(n24161), .ZN(n47472) );
  INV_X2 U16307 ( .I(n21241), .ZN(n5299) );
  INV_X1 U16311 ( .I(n44387), .ZN(n5573) );
  INV_X1 U16312 ( .I(n46149), .ZN(n44857) );
  INV_X1 U16313 ( .I(n25208), .ZN(n18124) );
  INV_X1 U16317 ( .I(n44923), .ZN(n2778) );
  INV_X1 U16318 ( .I(n25957), .ZN(n9874) );
  CLKBUF_X2 U16319 ( .I(n25982), .Z(n4761) );
  INV_X1 U16320 ( .I(n25602), .ZN(n46706) );
  INV_X1 U16321 ( .I(n46580), .ZN(n10812) );
  INV_X1 U16322 ( .I(n3913), .ZN(n44539) );
  INV_X1 U16324 ( .I(n4900), .ZN(n24979) );
  INV_X1 U16325 ( .I(n45815), .ZN(n9736) );
  INV_X1 U16326 ( .I(n45358), .ZN(n10700) );
  INV_X1 U16327 ( .I(n44626), .ZN(n7164) );
  INV_X1 U16328 ( .I(n21989), .ZN(n14873) );
  INV_X1 U16331 ( .I(n20324), .ZN(n12342) );
  INV_X1 U16332 ( .I(n7999), .ZN(n18986) );
  NAND2_X1 U16335 ( .A1(n6587), .A2(n5359), .ZN(n44976) );
  INV_X1 U16338 ( .I(n6204), .ZN(n44881) );
  CLKBUF_X2 U16339 ( .I(n4546), .Z(n10139) );
  INV_X1 U16343 ( .I(n20044), .ZN(n4218) );
  INV_X1 U16346 ( .I(n45859), .ZN(n12452) );
  INV_X1 U16347 ( .I(n23534), .ZN(n3474) );
  CLKBUF_X2 U16349 ( .I(n44129), .Z(n6967) );
  INV_X1 U16351 ( .I(n46163), .ZN(n44246) );
  INV_X1 U16353 ( .I(n1198), .ZN(n11185) );
  NAND2_X1 U16356 ( .A1(n2599), .A2(n2598), .ZN(n2597) );
  INV_X1 U16358 ( .I(n23131), .ZN(n46188) );
  CLKBUF_X2 U16361 ( .I(n46620), .Z(n10620) );
  INV_X1 U16362 ( .I(n44254), .ZN(n4800) );
  INV_X1 U16365 ( .I(n23696), .ZN(n12501) );
  INV_X1 U16368 ( .I(n46229), .ZN(n5809) );
  INV_X1 U16369 ( .I(n46312), .ZN(n13513) );
  INV_X1 U16371 ( .I(n19071), .ZN(n6755) );
  INV_X4 U16374 ( .I(n2722), .ZN(n46197) );
  INV_X1 U16379 ( .I(n46558), .ZN(n11877) );
  INV_X2 U16380 ( .I(n20824), .ZN(n1676) );
  INV_X2 U16381 ( .I(n19433), .ZN(n1677) );
  INV_X2 U16383 ( .I(n24068), .ZN(n1678) );
  CLKBUF_X2 U16393 ( .I(n19155), .Z(n4529) );
  NAND2_X1 U16403 ( .A1(n46342), .A2(n46341), .ZN(n46656) );
  INV_X1 U16404 ( .I(n244), .ZN(n8869) );
  NAND2_X1 U16405 ( .A1(n12666), .A2(n42746), .ZN(n4317) );
  NOR2_X1 U16406 ( .A1(n20329), .A2(n20330), .ZN(n6785) );
  OAI21_X1 U16409 ( .A1(n16942), .A2(n19961), .B(n1503), .ZN(n16549) );
  NOR2_X1 U16412 ( .A1(n19486), .A2(n19487), .ZN(n5853) );
  INV_X1 U16413 ( .I(n6423), .ZN(n6420) );
  NOR2_X1 U16418 ( .A1(n6969), .A2(n16201), .ZN(n6968) );
  CLKBUF_X2 U16421 ( .I(n46166), .Z(n23059) );
  NOR2_X1 U16429 ( .A1(n11406), .A2(n43950), .ZN(n10159) );
  INV_X1 U16431 ( .I(n46187), .ZN(n15015) );
  INV_X1 U16432 ( .I(n45070), .ZN(n2453) );
  CLKBUF_X2 U16434 ( .I(n46529), .Z(n23872) );
  NAND2_X1 U16443 ( .A1(n41531), .A2(n8425), .ZN(n41534) );
  OAI22_X1 U16444 ( .A1(n43949), .A2(n43304), .B1(n42798), .B2(n59709), .ZN(
        n42799) );
  INV_X1 U16446 ( .I(n13912), .ZN(n13911) );
  NAND2_X1 U16455 ( .A1(n43296), .A2(n43951), .ZN(n16942) );
  NAND2_X1 U16456 ( .A1(n9668), .A2(n42672), .ZN(n7827) );
  NAND2_X1 U16458 ( .A1(n24591), .A2(n43322), .ZN(n14657) );
  AOI21_X1 U16461 ( .A1(n42745), .A2(n42744), .B(n42743), .ZN(n42746) );
  NAND2_X1 U16463 ( .A1(n6639), .A2(n11986), .ZN(n3004) );
  INV_X1 U16468 ( .I(n42743), .ZN(n13450) );
  NAND2_X1 U16470 ( .A1(n6427), .A2(n6426), .ZN(n6422) );
  OAI21_X1 U16471 ( .A1(n43855), .A2(n43854), .B(n43853), .ZN(n11156) );
  NOR2_X1 U16475 ( .A1(n21935), .A2(n43119), .ZN(n9748) );
  NAND2_X1 U16477 ( .A1(n43424), .A2(n22087), .ZN(n6022) );
  NAND2_X1 U16479 ( .A1(n21916), .A2(n21917), .ZN(n20722) );
  NAND2_X1 U16480 ( .A1(n6070), .A2(n6067), .ZN(n5327) );
  NAND2_X1 U16485 ( .A1(n42932), .A2(n42928), .ZN(n15492) );
  NOR2_X1 U16487 ( .A1(n15813), .A2(n21376), .ZN(n9438) );
  INV_X1 U16488 ( .I(n41563), .ZN(n21347) );
  OAI21_X1 U16489 ( .A1(n43699), .A2(n14214), .B(n12447), .ZN(n12446) );
  INV_X1 U16490 ( .I(n14262), .ZN(n43228) );
  AOI21_X1 U16498 ( .A1(n12971), .A2(n43612), .B(n12969), .ZN(n13108) );
  NAND2_X1 U16509 ( .A1(n8430), .A2(n8429), .ZN(n12137) );
  NAND2_X1 U16511 ( .A1(n12389), .A2(n42376), .ZN(n41533) );
  INV_X1 U16513 ( .I(n41330), .ZN(n7215) );
  NAND2_X1 U16515 ( .A1(n43477), .A2(n18650), .ZN(n43479) );
  OAI22_X1 U16516 ( .A1(n42538), .A2(n42539), .B1(n20380), .B2(n43956), .ZN(
        n6639) );
  NAND2_X1 U16520 ( .A1(n43895), .A2(n43894), .ZN(n43896) );
  OAI22_X1 U16521 ( .A1(n40085), .A2(n40084), .B1(n13750), .B2(n40082), .ZN(
        n12143) );
  NAND2_X1 U16522 ( .A1(n43997), .A2(n43996), .ZN(n3209) );
  NOR2_X1 U16525 ( .A1(n21798), .A2(n43982), .ZN(n3210) );
  NAND2_X1 U16526 ( .A1(n7177), .A2(n42823), .ZN(n9668) );
  AOI22_X1 U16534 ( .A1(n20632), .A2(n42837), .B1(n21426), .B2(n42827), .ZN(
        n7829) );
  NOR2_X1 U16536 ( .A1(n43955), .A2(n9248), .ZN(n9247) );
  NAND2_X1 U16537 ( .A1(n43070), .A2(n22673), .ZN(n21917) );
  OAI21_X1 U16539 ( .A1(n10991), .A2(n10989), .B(n4689), .ZN(n21916) );
  OAI21_X1 U16549 ( .A1(n10299), .A2(n43028), .B(n10298), .ZN(n25757) );
  AOI21_X1 U16551 ( .A1(n1333), .A2(n43891), .B(n43232), .ZN(n43240) );
  NAND2_X1 U16552 ( .A1(n9503), .A2(n39428), .ZN(n39433) );
  NOR2_X1 U16553 ( .A1(n12903), .A2(n12902), .ZN(n12901) );
  INV_X1 U16557 ( .I(n22109), .ZN(n5851) );
  NAND2_X1 U16559 ( .A1(n11365), .A2(n11364), .ZN(n11363) );
  NOR2_X1 U16560 ( .A1(n15502), .A2(n43850), .ZN(n5849) );
  OAI21_X1 U16561 ( .A1(n43652), .A2(n3484), .B(n43889), .ZN(n10199) );
  NAND2_X1 U16562 ( .A1(n13452), .A2(n13454), .ZN(n6421) );
  AOI21_X1 U16569 ( .A1(n43143), .A2(n13037), .B(n3452), .ZN(n3451) );
  NAND2_X1 U16574 ( .A1(n23196), .A2(n3696), .ZN(n3450) );
  INV_X1 U16575 ( .I(n43850), .ZN(n43855) );
  INV_X1 U16577 ( .I(n13832), .ZN(n42752) );
  NAND2_X1 U16583 ( .A1(n42856), .A2(n2587), .ZN(n42857) );
  OAI21_X1 U16585 ( .A1(n15219), .A2(n15218), .B(n15217), .ZN(n16340) );
  INV_X1 U16586 ( .I(n41579), .ZN(n42548) );
  INV_X1 U16587 ( .I(n16148), .ZN(n9032) );
  NAND2_X1 U16588 ( .A1(n41522), .A2(n42703), .ZN(n13978) );
  NAND2_X1 U16590 ( .A1(n43580), .A2(n6866), .ZN(n2690) );
  NAND2_X1 U16591 ( .A1(n43653), .A2(n3485), .ZN(n3484) );
  INV_X1 U16593 ( .I(n42881), .ZN(n4573) );
  AND2_X1 U16595 ( .A1(n43689), .A2(n4229), .Z(n4228) );
  NOR2_X1 U16596 ( .A1(n40279), .A2(n64663), .ZN(n5543) );
  INV_X1 U16598 ( .I(n24216), .ZN(n6067) );
  OAI22_X1 U16599 ( .A1(n4609), .A2(n41729), .B1(n6706), .B2(n42146), .ZN(
        n41371) );
  INV_X1 U16602 ( .I(n42184), .ZN(n10299) );
  INV_X1 U16603 ( .I(n42112), .ZN(n10466) );
  NAND2_X1 U16605 ( .A1(n40600), .A2(n40599), .ZN(n8612) );
  INV_X1 U16610 ( .I(n9511), .ZN(n11059) );
  AOI21_X1 U16613 ( .A1(n43256), .A2(n21800), .B(n20294), .ZN(n20293) );
  NOR2_X1 U16614 ( .A1(n43305), .A2(n44229), .ZN(n20322) );
  AND2_X1 U16615 ( .A1(n16298), .A2(n17755), .Z(n42798) );
  INV_X1 U16616 ( .I(n43107), .ZN(n40881) );
  NAND2_X1 U16622 ( .A1(n9697), .A2(n41044), .ZN(n6973) );
  AOI21_X1 U16624 ( .A1(n2448), .A2(n23838), .B(n4322), .ZN(n2446) );
  OAI21_X1 U16626 ( .A1(n43312), .A2(n43714), .B(n44230), .ZN(n43314) );
  NOR2_X1 U16627 ( .A1(n41320), .A2(n1332), .ZN(n25795) );
  NOR2_X1 U16628 ( .A1(n43213), .A2(n13882), .ZN(n43215) );
  NAND2_X1 U16630 ( .A1(n14404), .A2(n12694), .ZN(n11536) );
  INV_X1 U16632 ( .I(n39938), .ZN(n3227) );
  NAND2_X1 U16633 ( .A1(n46326), .A2(n13680), .ZN(n13679) );
  INV_X1 U16634 ( .I(n42557), .ZN(n9600) );
  NAND2_X1 U16637 ( .A1(n5949), .A2(n41584), .ZN(n5948) );
  INV_X1 U16638 ( .I(n3965), .ZN(n3964) );
  OAI21_X1 U16639 ( .A1(n41555), .A2(n4588), .B(n4587), .ZN(n41563) );
  NOR2_X1 U16644 ( .A1(n16997), .A2(n43696), .ZN(n8191) );
  INV_X1 U16649 ( .I(n41484), .ZN(n43324) );
  INV_X1 U16655 ( .I(n41481), .ZN(n12576) );
  NOR2_X1 U16658 ( .A1(n42033), .A2(n42034), .ZN(n2707) );
  NOR2_X1 U16659 ( .A1(n20451), .A2(n43157), .ZN(n43158) );
  NAND2_X1 U16660 ( .A1(n24191), .A2(n43959), .ZN(n9248) );
  OAI22_X1 U16661 ( .A1(n43976), .A2(n6007), .B1(n43977), .B2(n9163), .ZN(
        n43983) );
  INV_X1 U16662 ( .I(n24191), .ZN(n7144) );
  NOR2_X1 U16664 ( .A1(n15337), .A2(n42839), .ZN(n42829) );
  OAI22_X1 U16665 ( .A1(n42780), .A2(n16262), .B1(n24762), .B2(n43022), .ZN(
        n24764) );
  NOR2_X1 U16668 ( .A1(n43868), .A2(n1492), .ZN(n11067) );
  NAND2_X1 U16670 ( .A1(n43430), .A2(n43437), .ZN(n15376) );
  OR2_X1 U16671 ( .A1(n8343), .A2(n43094), .Z(n4657) );
  AND2_X1 U16674 ( .A1(n43426), .A2(n42366), .Z(n18405) );
  AOI21_X1 U16675 ( .A1(n25711), .A2(n25710), .B(n25709), .ZN(n25708) );
  NOR2_X1 U16677 ( .A1(n42761), .A2(n19271), .ZN(n23013) );
  NAND2_X1 U16678 ( .A1(n16148), .A2(n42076), .ZN(n8430) );
  NAND2_X1 U16679 ( .A1(n8171), .A2(n43342), .ZN(n8876) );
  INV_X1 U16680 ( .I(n57410), .ZN(n42801) );
  NAND2_X1 U16681 ( .A1(n42622), .A2(n13201), .ZN(n13200) );
  NOR2_X1 U16682 ( .A1(n43190), .A2(n24492), .ZN(n24491) );
  AOI21_X1 U16683 ( .A1(n42312), .A2(n43986), .B(n42311), .ZN(n21138) );
  NAND2_X1 U16685 ( .A1(n43146), .A2(n43144), .ZN(n3452) );
  INV_X1 U16687 ( .I(n8981), .ZN(n43106) );
  OAI21_X1 U16689 ( .A1(n41711), .A2(n21408), .B(n21950), .ZN(n11364) );
  NAND2_X1 U16691 ( .A1(n43994), .A2(n15639), .ZN(n43996) );
  INV_X1 U16692 ( .I(n43091), .ZN(n14261) );
  INV_X1 U16694 ( .I(n43297), .ZN(n42533) );
  OAI22_X1 U16695 ( .A1(n39015), .A2(n1297), .B1(n42927), .B2(n13074), .ZN(
        n12902) );
  INV_X1 U16698 ( .I(n14408), .ZN(n42539) );
  NAND2_X1 U16699 ( .A1(n43625), .A2(n43552), .ZN(n43556) );
  NAND2_X1 U16700 ( .A1(n42097), .A2(n21527), .ZN(n41956) );
  INV_X1 U16701 ( .I(n7877), .ZN(n41701) );
  OAI21_X1 U16703 ( .A1(n41790), .A2(n8028), .B(n43268), .ZN(n39798) );
  INV_X1 U16704 ( .I(n20685), .ZN(n43245) );
  AND3_X1 U16707 ( .A1(n42753), .A2(n42759), .A3(n22182), .Z(n16459) );
  AND2_X1 U16709 ( .A1(n43651), .A2(n61951), .Z(n43652) );
  AND2_X1 U16710 ( .A1(n60583), .A2(n22673), .Z(n43840) );
  NAND2_X1 U16711 ( .A1(n39802), .A2(n63529), .ZN(n15217) );
  AND2_X1 U16712 ( .A1(n43457), .A2(n43478), .Z(n16156) );
  INV_X1 U16717 ( .I(n12154), .ZN(n5340) );
  NAND2_X1 U16719 ( .A1(n42553), .A2(n23702), .ZN(n42101) );
  NOR2_X1 U16721 ( .A1(n16998), .A2(n42019), .ZN(n8192) );
  NAND2_X1 U16723 ( .A1(n43317), .A2(n1298), .ZN(n20688) );
  AND2_X1 U16724 ( .A1(n43948), .A2(n43957), .Z(n15334) );
  AND2_X1 U16726 ( .A1(n42050), .A2(n18143), .Z(n18406) );
  NAND2_X1 U16729 ( .A1(n6563), .A2(n1493), .ZN(n42424) );
  INV_X1 U16730 ( .I(n13621), .ZN(n40868) );
  OR2_X1 U16732 ( .A1(n43289), .A2(n2735), .Z(n20067) );
  OR2_X1 U16733 ( .A1(n43303), .A2(n43957), .Z(n20380) );
  INV_X1 U16734 ( .I(n42942), .ZN(n9850) );
  INV_X1 U16735 ( .I(n43986), .ZN(n44232) );
  NAND2_X1 U16740 ( .A1(n24685), .A2(n24684), .ZN(n40894) );
  NOR2_X1 U16741 ( .A1(n8962), .A2(n15219), .ZN(n41320) );
  OAI21_X1 U16742 ( .A1(n41734), .A2(n20784), .B(n21469), .ZN(n41735) );
  NAND3_X1 U16743 ( .A1(n62043), .A2(n61745), .A3(n43042), .ZN(n43045) );
  NOR2_X1 U16744 ( .A1(n43286), .A2(n15020), .ZN(n43275) );
  NAND2_X1 U16746 ( .A1(n41341), .A2(n14896), .ZN(n41342) );
  NAND2_X1 U16748 ( .A1(n64291), .A2(n42607), .ZN(n9212) );
  NAND2_X1 U16750 ( .A1(n42642), .A2(n13678), .ZN(n13677) );
  INV_X1 U16751 ( .I(n46331), .ZN(n13680) );
  NAND2_X1 U16753 ( .A1(n3630), .A2(n42670), .ZN(n3628) );
  INV_X1 U16754 ( .I(n41651), .ZN(n41652) );
  NAND2_X1 U16755 ( .A1(n41556), .A2(n9914), .ZN(n4587) );
  INV_X1 U16756 ( .I(n43892), .ZN(n42860) );
  NAND2_X1 U16759 ( .A1(n43085), .A2(n11476), .ZN(n39878) );
  NAND3_X1 U16760 ( .A1(n39171), .A2(n41990), .A3(n39170), .ZN(n39172) );
  NAND2_X1 U16761 ( .A1(n42926), .A2(n1297), .ZN(n8907) );
  NAND3_X1 U16762 ( .A1(n42926), .A2(n13074), .A3(n13073), .ZN(n12904) );
  NOR2_X1 U16763 ( .A1(n42968), .A2(n13476), .ZN(n40081) );
  AOI21_X1 U16764 ( .A1(n61186), .A2(n2496), .B(n19428), .ZN(n42802) );
  NOR2_X1 U16765 ( .A1(n42836), .A2(n42827), .ZN(n11866) );
  OR2_X1 U16767 ( .A1(n1299), .A2(n1503), .Z(n16298) );
  OR2_X1 U16768 ( .A1(n62546), .A2(n42543), .Z(n7032) );
  NAND2_X1 U16771 ( .A1(n42403), .A2(n64492), .ZN(n9034) );
  INV_X1 U16772 ( .I(n23195), .ZN(n7490) );
  INV_X1 U16775 ( .I(n43121), .ZN(n43127) );
  NOR2_X1 U16777 ( .A1(n25439), .A2(n25440), .ZN(n7049) );
  NOR2_X1 U16780 ( .A1(n13595), .A2(n41322), .ZN(n9886) );
  INV_X1 U16781 ( .I(n43869), .ZN(n38353) );
  NAND2_X1 U16782 ( .A1(n43018), .A2(n43020), .ZN(n9643) );
  NOR2_X1 U16783 ( .A1(n1493), .A2(n15020), .ZN(n43280) );
  INV_X1 U16785 ( .I(n1908), .ZN(n41519) );
  INV_X1 U16786 ( .I(n42108), .ZN(n42103) );
  INV_X1 U16788 ( .I(n42842), .ZN(n18022) );
  OAI22_X1 U16791 ( .A1(n37537), .A2(n9295), .B1(n12378), .B2(n42593), .ZN(
        n37538) );
  INV_X1 U16794 ( .I(n2121), .ZN(n41797) );
  AND2_X1 U16800 ( .A1(n19761), .A2(n43980), .Z(n16144) );
  OR2_X1 U16801 ( .A1(n13385), .A2(n42655), .Z(n2448) );
  NAND2_X1 U16802 ( .A1(n23279), .A2(n7516), .ZN(n13167) );
  AND2_X1 U16805 ( .A1(n43178), .A2(n20888), .Z(n16076) );
  OR2_X1 U16806 ( .A1(n13100), .A2(n8350), .Z(n8349) );
  NAND2_X1 U16808 ( .A1(n41981), .A2(n1500), .ZN(n12927) );
  NOR2_X1 U16813 ( .A1(n42940), .A2(n43438), .ZN(n16260) );
  INV_X1 U16814 ( .I(n43875), .ZN(n5801) );
  INV_X1 U16817 ( .I(n42540), .ZN(n13073) );
  NAND2_X1 U16818 ( .A1(n3674), .A2(n61107), .ZN(n3675) );
  AND2_X1 U16820 ( .A1(n42415), .A2(n13750), .Z(n15122) );
  NAND3_X1 U16821 ( .A1(n1393), .A2(n4805), .A3(n42386), .ZN(n42388) );
  INV_X1 U16825 ( .I(n42747), .ZN(n7996) );
  NAND2_X1 U16826 ( .A1(n42910), .A2(n42911), .ZN(n42913) );
  AND2_X1 U16830 ( .A1(n42064), .A2(n43916), .Z(n1934) );
  NAND2_X1 U16831 ( .A1(n1336), .A2(n13749), .ZN(n43469) );
  INV_X1 U16832 ( .I(n43093), .ZN(n25537) );
  NAND2_X1 U16833 ( .A1(n42998), .A2(n4659), .ZN(n42999) );
  INV_X1 U16835 ( .I(n25440), .ZN(n2580) );
  NAND2_X1 U16836 ( .A1(n20276), .A2(n12089), .ZN(n43539) );
  NOR2_X1 U16838 ( .A1(n16864), .A2(n12089), .ZN(n43536) );
  NOR2_X1 U16840 ( .A1(n42553), .A2(n42555), .ZN(n15233) );
  INV_X1 U16842 ( .I(n17176), .ZN(n42794) );
  NOR2_X1 U16843 ( .A1(n42553), .A2(n42554), .ZN(n5280) );
  NAND2_X1 U16845 ( .A1(n11727), .A2(n7620), .ZN(n39797) );
  NOR2_X1 U16847 ( .A1(n40284), .A2(n22999), .ZN(n4648) );
  AND2_X1 U16848 ( .A1(n22087), .A2(n57810), .Z(n43554) );
  NOR2_X1 U16850 ( .A1(n59746), .A2(n2994), .ZN(n41139) );
  NAND2_X1 U16851 ( .A1(n1497), .A2(n42837), .ZN(n11625) );
  NAND2_X1 U16852 ( .A1(n6706), .A2(n42672), .ZN(n22225) );
  INV_X1 U16854 ( .I(n41340), .ZN(n14896) );
  INV_X1 U16856 ( .I(n41325), .ZN(n41791) );
  NOR2_X1 U16858 ( .A1(n42067), .A2(n43474), .ZN(n7366) );
  INV_X1 U16859 ( .I(n42371), .ZN(n42935) );
  AND2_X1 U16860 ( .A1(n43582), .A2(n2995), .Z(n6866) );
  INV_X1 U16861 ( .I(n43605), .ZN(n12970) );
  INV_X1 U16862 ( .I(n43026), .ZN(n9822) );
  AOI21_X1 U16864 ( .A1(n10970), .A2(n20244), .B(n42694), .ZN(n40175) );
  OR2_X1 U16866 ( .A1(n11747), .A2(n10990), .Z(n10989) );
  OR2_X1 U16867 ( .A1(n41715), .A2(n42551), .Z(n6338) );
  INV_X1 U16871 ( .I(n60583), .ZN(n43058) );
  INV_X1 U16872 ( .I(n42014), .ZN(n43097) );
  INV_X1 U16876 ( .I(n42976), .ZN(n10882) );
  CLKBUF_X2 U16877 ( .I(n43561), .Z(n5001) );
  INV_X1 U16879 ( .I(n41584), .ZN(n42544) );
  INV_X2 U16880 ( .I(n43989), .ZN(n43309) );
  NAND2_X1 U16881 ( .A1(n42655), .A2(n60846), .ZN(n40366) );
  INV_X1 U16884 ( .I(n43734), .ZN(n42119) );
  INV_X1 U16885 ( .I(n42167), .ZN(n42166) );
  NAND2_X1 U16886 ( .A1(n42875), .A2(n1502), .ZN(n42869) );
  INV_X1 U16890 ( .I(n42551), .ZN(n9566) );
  INV_X2 U16891 ( .I(n43657), .ZN(n2588) );
  OR2_X1 U16892 ( .A1(n42397), .A2(n41689), .Z(n6268) );
  INV_X1 U16893 ( .I(n41532), .ZN(n12389) );
  NOR2_X1 U16894 ( .A1(n8352), .A2(n42016), .ZN(n13100) );
  AND2_X1 U16897 ( .A1(n2557), .A2(n63529), .Z(n3328) );
  BUF_X4 U16898 ( .I(n23984), .Z(n15540) );
  OR2_X1 U16899 ( .A1(n42120), .A2(n19358), .Z(n43212) );
  INV_X1 U16905 ( .I(n43098), .ZN(n7577) );
  NOR2_X1 U16906 ( .A1(n42151), .A2(n8912), .ZN(n21426) );
  INV_X1 U16913 ( .I(n43102), .ZN(n43086) );
  OR2_X1 U16921 ( .A1(n22446), .A2(n42155), .Z(n13105) );
  NAND2_X1 U16922 ( .A1(n22716), .A2(n6007), .ZN(n43708) );
  NOR2_X1 U16926 ( .A1(n61107), .A2(n6297), .ZN(n8215) );
  INV_X1 U16927 ( .I(n19517), .ZN(n41692) );
  INV_X1 U16928 ( .I(n43957), .ZN(n18723) );
  INV_X4 U16930 ( .I(n5125), .ZN(n37536) );
  AND2_X1 U16931 ( .A1(n42827), .A2(n42672), .Z(n16134) );
  INV_X1 U16933 ( .I(n43490), .ZN(n12644) );
  INV_X2 U16935 ( .I(n9427), .ZN(n8911) );
  NAND2_X1 U16936 ( .A1(n10203), .A2(n7285), .ZN(n43226) );
  OR2_X1 U16937 ( .A1(n41353), .A2(n43225), .Z(n16231) );
  NAND2_X1 U16939 ( .A1(n1502), .A2(n42868), .ZN(n41503) );
  NOR3_X1 U16941 ( .A1(n22446), .A2(n43601), .A3(n42155), .ZN(n13107) );
  INV_X4 U16942 ( .I(n43124), .ZN(n1701) );
  INV_X1 U16946 ( .I(n7749), .ZN(n5796) );
  NOR2_X1 U16954 ( .A1(n19642), .A2(n18755), .ZN(n18754) );
  NAND2_X1 U16956 ( .A1(n19386), .A2(n19384), .ZN(n39956) );
  CLKBUF_X2 U16962 ( .I(n42993), .Z(n10203) );
  INV_X2 U16965 ( .I(n42104), .ZN(n4077) );
  INV_X2 U16966 ( .I(n40839), .ZN(n24360) );
  INV_X1 U16969 ( .I(n14620), .ZN(n4107) );
  INV_X1 U16971 ( .I(n577), .ZN(n8937) );
  NAND2_X1 U16975 ( .A1(n18593), .A2(n41463), .ZN(n5211) );
  NAND2_X1 U16976 ( .A1(n4455), .A2(n734), .ZN(n20392) );
  OAI21_X1 U16979 ( .A1(n4967), .A2(n40034), .B(n40355), .ZN(n18755) );
  NOR2_X1 U16985 ( .A1(n39610), .A2(n40382), .ZN(n12244) );
  NAND2_X1 U16986 ( .A1(n17751), .A2(n5847), .ZN(n14497) );
  NOR2_X1 U16987 ( .A1(n40163), .A2(n11129), .ZN(n11128) );
  NAND2_X1 U16989 ( .A1(n41450), .A2(n41449), .ZN(n12187) );
  NAND2_X1 U16990 ( .A1(n19387), .A2(n39954), .ZN(n19386) );
  INV_X1 U16991 ( .I(n41313), .ZN(n17043) );
  BUF_X4 U16994 ( .I(n42583), .Z(n1716) );
  OAI21_X1 U16995 ( .A1(n4952), .A2(n4951), .B(n25358), .ZN(n2561) );
  AOI22_X1 U16997 ( .A1(n40037), .A2(n40039), .B1(n9798), .B2(n19331), .ZN(
        n40044) );
  NAND3_X1 U17005 ( .A1(n40168), .A2(n64948), .A3(n6576), .ZN(n40169) );
  NAND2_X1 U17006 ( .A1(n40168), .A2(n40242), .ZN(n7392) );
  NAND2_X1 U17007 ( .A1(n40233), .A2(n40159), .ZN(n2166) );
  OR2_X1 U17008 ( .A1(n41647), .A2(n6855), .Z(n24792) );
  INV_X4 U17011 ( .I(n6797), .ZN(n43572) );
  NOR2_X1 U17012 ( .A1(n42475), .A2(n40038), .ZN(n18041) );
  INV_X1 U17014 ( .I(n23380), .ZN(n15159) );
  NOR2_X1 U17016 ( .A1(n12736), .A2(n12731), .ZN(n12730) );
  INV_X1 U17017 ( .I(n39849), .ZN(n13863) );
  AOI21_X1 U17019 ( .A1(n6838), .A2(n10074), .B(n17019), .ZN(n17536) );
  AOI21_X1 U17027 ( .A1(n41094), .A2(n5516), .B(n40580), .ZN(n5515) );
  NAND2_X1 U17028 ( .A1(n42228), .A2(n63435), .ZN(n8404) );
  AOI21_X1 U17029 ( .A1(n41061), .A2(n39796), .B(n39794), .ZN(n9350) );
  NOR2_X1 U17030 ( .A1(n41181), .A2(n41180), .ZN(n6707) );
  AOI21_X1 U17031 ( .A1(n18304), .A2(n11244), .B(n25305), .ZN(n4967) );
  NAND2_X1 U17032 ( .A1(n7502), .A2(n7501), .ZN(n7500) );
  INV_X1 U17034 ( .I(n4132), .ZN(n4131) );
  NOR2_X1 U17035 ( .A1(n24400), .A2(n42266), .ZN(n5509) );
  NAND2_X1 U17039 ( .A1(n40714), .A2(n60810), .ZN(n40718) );
  NAND2_X1 U17041 ( .A1(n39923), .A2(n39922), .ZN(n22259) );
  NOR2_X1 U17043 ( .A1(n39054), .A2(n17130), .ZN(n39055) );
  INV_X1 U17044 ( .I(n16643), .ZN(n17355) );
  NOR2_X1 U17045 ( .A1(n42258), .A2(n42260), .ZN(n5514) );
  OAI21_X1 U17046 ( .A1(n42290), .A2(n3457), .B(n3455), .ZN(n41249) );
  OAI22_X1 U17048 ( .A1(n40379), .A2(n11646), .B1(n41445), .B2(n41428), .ZN(
        n11645) );
  INV_X1 U17051 ( .I(n41441), .ZN(n12194) );
  NAND3_X1 U17054 ( .A1(n25219), .A2(n42205), .A3(n15814), .ZN(n25218) );
  NOR2_X1 U17055 ( .A1(n5797), .A2(n13756), .ZN(n5795) );
  NOR2_X1 U17056 ( .A1(n7951), .A2(n22290), .ZN(n38275) );
  AOI21_X1 U17058 ( .A1(n40675), .A2(n41460), .B(n25777), .ZN(n25776) );
  OAI21_X1 U17059 ( .A1(n25596), .A2(n42447), .B(n1401), .ZN(n10106) );
  NOR2_X1 U17061 ( .A1(n41837), .A2(n1273), .ZN(n16297) );
  NAND3_X1 U17067 ( .A1(n40380), .A2(n23406), .A3(n19385), .ZN(n19384) );
  INV_X1 U17070 ( .I(n42205), .ZN(n20669) );
  OAI21_X1 U17071 ( .A1(n40590), .A2(n40589), .B(n64592), .ZN(n14621) );
  NAND2_X1 U17073 ( .A1(n25286), .A2(n25285), .ZN(n14906) );
  AOI21_X1 U17079 ( .A1(n41836), .A2(n16079), .B(n24751), .ZN(n24750) );
  AOI21_X1 U17080 ( .A1(n38934), .A2(n40405), .B(n38933), .ZN(n12948) );
  NAND3_X1 U17081 ( .A1(n2586), .A2(n42209), .A3(n23501), .ZN(n41291) );
  AOI22_X1 U17082 ( .A1(n40216), .A2(n5394), .B1(n40211), .B2(n40212), .ZN(
        n3135) );
  AOI22_X1 U17084 ( .A1(n41839), .A2(n42474), .B1(n9627), .B2(n14524), .ZN(
        n41840) );
  INV_X1 U17089 ( .I(n41260), .ZN(n3060) );
  AOI22_X1 U17091 ( .A1(n40307), .A2(n40306), .B1(n40302), .B2(n40301), .ZN(
        n26205) );
  OAI21_X1 U17092 ( .A1(n42210), .A2(n65199), .B(n1506), .ZN(n42220) );
  OAI21_X1 U17093 ( .A1(n42474), .A2(n11101), .B(n18045), .ZN(n12851) );
  AOI21_X1 U17094 ( .A1(n42492), .A2(n42491), .B(n12464), .ZN(n12680) );
  AOI22_X1 U17097 ( .A1(n42429), .A2(n14863), .B1(n4248), .B2(n4150), .ZN(
        n4763) );
  INV_X1 U17098 ( .I(n12101), .ZN(n41827) );
  OAI22_X1 U17099 ( .A1(n39844), .A2(n39843), .B1(n41433), .B2(n15441), .ZN(
        n10878) );
  AOI22_X1 U17102 ( .A1(n42234), .A2(n41945), .B1(n41800), .B2(n8841), .ZN(
        n8840) );
  OAI21_X1 U17105 ( .A1(n22154), .A2(n40650), .B(n22004), .ZN(n22003) );
  NAND2_X1 U17106 ( .A1(n20638), .A2(n13511), .ZN(n7869) );
  AOI22_X1 U17110 ( .A1(n40608), .A2(n16467), .B1(n40612), .B2(n20054), .ZN(
        n16466) );
  OAI21_X1 U17111 ( .A1(n61986), .A2(n38039), .B(n38038), .ZN(n38044) );
  AOI22_X1 U17112 ( .A1(n4358), .A2(n9790), .B1(n40853), .B2(n4357), .ZN(
        n20585) );
  AOI21_X1 U17113 ( .A1(n8070), .A2(n40362), .B(n8069), .ZN(n8068) );
  AOI22_X1 U17116 ( .A1(n64948), .A2(n40238), .B1(n40075), .B2(n40239), .ZN(
        n40077) );
  OAI21_X1 U17117 ( .A1(n37933), .A2(n65206), .B(n40472), .ZN(n37937) );
  OR2_X1 U17119 ( .A1(n6839), .A2(n39999), .Z(n6838) );
  NAND2_X1 U17120 ( .A1(n41037), .A2(n40519), .ZN(n13133) );
  INV_X1 U17123 ( .I(n10133), .ZN(n41176) );
  NAND2_X1 U17124 ( .A1(n40126), .A2(n16396), .ZN(n16394) );
  NOR2_X1 U17125 ( .A1(n2895), .A2(n6843), .ZN(n13551) );
  OR2_X1 U17127 ( .A1(n1932), .A2(n11995), .Z(n20094) );
  NAND2_X1 U17130 ( .A1(n40655), .A2(n11193), .ZN(n40674) );
  NAND2_X1 U17133 ( .A1(n40561), .A2(n40790), .ZN(n15633) );
  AOI21_X1 U17134 ( .A1(n41813), .A2(n11994), .B(n41820), .ZN(n1979) );
  AOI21_X1 U17136 ( .A1(n38676), .A2(n9589), .B(n22330), .ZN(n9588) );
  OAI22_X1 U17137 ( .A1(n40709), .A2(n40708), .B1(n40713), .B2(n25839), .ZN(
        n40711) );
  NAND2_X1 U17141 ( .A1(n6305), .A2(n22289), .ZN(n41300) );
  NAND2_X1 U17142 ( .A1(n40835), .A2(n9909), .ZN(n7502) );
  NAND2_X1 U17144 ( .A1(n41175), .A2(n24881), .ZN(n41181) );
  NAND3_X1 U17145 ( .A1(n5241), .A2(n41110), .A3(n41111), .ZN(n41115) );
  NAND2_X1 U17148 ( .A1(n41003), .A2(n37528), .ZN(n25286) );
  AOI22_X1 U17153 ( .A1(n39097), .A2(n36107), .B1(n21162), .B2(n1400), .ZN(
        n21161) );
  NAND2_X1 U17154 ( .A1(n7848), .A2(n41433), .ZN(n18085) );
  NOR2_X1 U17162 ( .A1(n41080), .A2(n18365), .ZN(n41089) );
  NOR2_X1 U17164 ( .A1(n38689), .A2(n40726), .ZN(n24486) );
  NAND2_X1 U17170 ( .A1(n14654), .A2(n4359), .ZN(n4358) );
  NAND2_X1 U17174 ( .A1(n22224), .A2(n59252), .ZN(n20638) );
  OAI21_X1 U17176 ( .A1(n40239), .A2(n25661), .B(n40238), .ZN(n40240) );
  NAND2_X1 U17177 ( .A1(n1001), .A2(n14815), .ZN(n14814) );
  NOR2_X1 U17178 ( .A1(n15344), .A2(n8919), .ZN(n8918) );
  INV_X1 U17181 ( .I(n41442), .ZN(n10879) );
  INV_X1 U17183 ( .I(n12805), .ZN(n38934) );
  NOR2_X1 U17184 ( .A1(n22758), .A2(n41414), .ZN(n6879) );
  NAND2_X1 U17185 ( .A1(n42497), .A2(n42496), .ZN(n16015) );
  AOI21_X1 U17187 ( .A1(n39098), .A2(n1400), .B(n9188), .ZN(n21383) );
  OAI21_X1 U17188 ( .A1(n6200), .A2(n61746), .B(n6199), .ZN(n6198) );
  AND2_X1 U17190 ( .A1(n40238), .A2(n40070), .Z(n39420) );
  INV_X1 U17191 ( .I(n42279), .ZN(n42283) );
  NOR2_X1 U17192 ( .A1(n40404), .A2(n41414), .ZN(n6874) );
  NAND2_X1 U17193 ( .A1(n40143), .A2(n6623), .ZN(n39330) );
  NAND2_X1 U17194 ( .A1(n40538), .A2(n3870), .ZN(n3869) );
  NOR2_X1 U17196 ( .A1(n40204), .A2(n40203), .ZN(n40209) );
  NAND2_X1 U17197 ( .A1(n41134), .A2(n11016), .ZN(n9870) );
  NAND2_X1 U17199 ( .A1(n39919), .A2(n40292), .ZN(n10972) );
  OAI21_X1 U17200 ( .A1(n57245), .A2(n41412), .B(n21001), .ZN(n13266) );
  NAND2_X1 U17203 ( .A1(n39012), .A2(n57925), .ZN(n5061) );
  INV_X1 U17204 ( .I(n39009), .ZN(n5063) );
  NAND2_X1 U17205 ( .A1(n41426), .A2(n41425), .ZN(n25417) );
  INV_X1 U17206 ( .I(n2338), .ZN(n2337) );
  AOI21_X1 U17207 ( .A1(n41440), .A2(n6993), .B(n41439), .ZN(n41441) );
  NAND3_X1 U17208 ( .A1(n11718), .A2(n41435), .A3(n41436), .ZN(n12192) );
  INV_X1 U17209 ( .I(n14987), .ZN(n14986) );
  AOI22_X1 U17210 ( .A1(n41471), .A2(n58047), .B1(n18661), .B2(n41476), .ZN(
        n14982) );
  NAND2_X1 U17211 ( .A1(n42527), .A2(n14279), .ZN(n42207) );
  NAND3_X1 U17212 ( .A1(n40335), .A2(n40336), .A3(n7694), .ZN(n40342) );
  OAI21_X1 U17213 ( .A1(n8246), .A2(n8245), .B(n22638), .ZN(n8244) );
  NOR2_X1 U17214 ( .A1(n23551), .A2(n39101), .ZN(n25272) );
  INV_X1 U17217 ( .I(n41467), .ZN(n8944) );
  NAND2_X1 U17218 ( .A1(n5393), .A2(n5392), .ZN(n3134) );
  NAND2_X1 U17219 ( .A1(n1001), .A2(n8116), .ZN(n37596) );
  NAND2_X1 U17220 ( .A1(n22346), .A2(n22345), .ZN(n40307) );
  AOI21_X1 U17222 ( .A1(n41193), .A2(n8536), .B(n15496), .ZN(n15495) );
  OAI22_X1 U17223 ( .A1(n10452), .A2(n65021), .B1(n41166), .B2(n41161), .ZN(
        n22224) );
  NAND2_X1 U17224 ( .A1(n2713), .A2(n40211), .ZN(n39326) );
  INV_X1 U17227 ( .I(n5508), .ZN(n5505) );
  OAI21_X1 U17228 ( .A1(n40309), .A2(n40310), .B(n42427), .ZN(n15670) );
  OAI21_X1 U17230 ( .A1(n41171), .A2(n24883), .B(n24882), .ZN(n24881) );
  OAI21_X1 U17232 ( .A1(n976), .A2(n22290), .B(n60143), .ZN(n41801) );
  NOR2_X1 U17234 ( .A1(n41230), .A2(n1303), .ZN(n15344) );
  NAND2_X1 U17236 ( .A1(n25651), .A2(n64566), .ZN(n22996) );
  INV_X1 U17240 ( .I(n42516), .ZN(n41832) );
  NAND2_X1 U17241 ( .A1(n18417), .A2(n59637), .ZN(n18414) );
  INV_X1 U17243 ( .I(n41394), .ZN(n11587) );
  NOR2_X1 U17244 ( .A1(n40415), .A2(n8942), .ZN(n7188) );
  NAND3_X1 U17245 ( .A1(n41807), .A2(n41806), .A3(n1510), .ZN(n41808) );
  OAI22_X1 U17246 ( .A1(n60229), .A2(n40258), .B1(n60172), .B2(n40257), .ZN(
        n39163) );
  OAI21_X1 U17247 ( .A1(n40516), .A2(n13136), .B(n20726), .ZN(n13135) );
  NAND2_X1 U17249 ( .A1(n60229), .A2(n40924), .ZN(n39165) );
  AOI21_X1 U17250 ( .A1(n41121), .A2(n17020), .B(n10074), .ZN(n17019) );
  NAND2_X1 U17251 ( .A1(n40287), .A2(n58970), .ZN(n14555) );
  NAND2_X1 U17252 ( .A1(n1504), .A2(n41035), .ZN(n8486) );
  NAND2_X1 U17253 ( .A1(n11718), .A2(n41445), .ZN(n39608) );
  OAI21_X1 U17254 ( .A1(n41272), .A2(n42299), .B(n2800), .ZN(n41273) );
  AND3_X1 U17255 ( .A1(n42289), .A2(n42287), .A3(n6412), .Z(n16055) );
  AOI21_X1 U17257 ( .A1(n24743), .A2(n41001), .B(n16468), .ZN(n16467) );
  NAND2_X1 U17259 ( .A1(n41261), .A2(n59531), .ZN(n3061) );
  INV_X1 U17260 ( .I(n3109), .ZN(n40120) );
  AOI22_X1 U17261 ( .A1(n40210), .A2(n18706), .B1(n61986), .B2(n10542), .ZN(
        n5391) );
  INV_X1 U17262 ( .I(n40948), .ZN(n18611) );
  INV_X1 U17264 ( .I(n42249), .ZN(n42255) );
  OAI21_X1 U17266 ( .A1(n40310), .A2(n24505), .B(n62018), .ZN(n13888) );
  NAND2_X1 U17268 ( .A1(n40124), .A2(n40125), .ZN(n20246) );
  NAND3_X1 U17269 ( .A1(n40065), .A2(n41817), .A3(n42446), .ZN(n1982) );
  NAND2_X1 U17271 ( .A1(n13725), .A2(n57207), .ZN(n13724) );
  INV_X1 U17273 ( .I(n6702), .ZN(n40317) );
  NAND2_X1 U17274 ( .A1(n63233), .A2(n65199), .ZN(n41295) );
  OAI21_X1 U17275 ( .A1(n42436), .A2(n42433), .B(n41825), .ZN(n4248) );
  OAI21_X1 U17279 ( .A1(n17930), .A2(n15655), .B(n38340), .ZN(n11436) );
  NOR2_X1 U17281 ( .A1(n42446), .A2(n10999), .ZN(n38339) );
  NOR2_X1 U17284 ( .A1(n39505), .A2(n18338), .ZN(n6800) );
  NAND2_X1 U17285 ( .A1(n41125), .A2(n21230), .ZN(n39698) );
  AND2_X1 U17288 ( .A1(n11016), .A2(n39505), .Z(n11015) );
  NAND2_X1 U17290 ( .A1(n37828), .A2(n41889), .ZN(n18892) );
  AND3_X1 U17292 ( .A1(n42288), .A2(n42287), .A3(n62134), .Z(n15894) );
  INV_X1 U17294 ( .I(n37196), .ZN(n11044) );
  INV_X1 U17297 ( .I(n15439), .ZN(n41443) );
  INV_X1 U17299 ( .I(n40698), .ZN(n18086) );
  NAND2_X1 U17301 ( .A1(n15369), .A2(n15367), .ZN(n19230) );
  NOR2_X1 U17302 ( .A1(n10956), .A2(n61986), .ZN(n10955) );
  OAI21_X1 U17303 ( .A1(n41232), .A2(n58046), .B(n39050), .ZN(n39012) );
  AOI21_X1 U17304 ( .A1(n42303), .A2(n13168), .B(n38270), .ZN(n38271) );
  INV_X1 U17305 ( .I(n39485), .ZN(n40572) );
  NAND2_X1 U17307 ( .A1(n61746), .A2(n7094), .ZN(n7681) );
  NAND2_X1 U17309 ( .A1(n39785), .A2(n2693), .ZN(n18744) );
  NAND2_X1 U17312 ( .A1(n1981), .A2(n40314), .ZN(n39929) );
  NOR2_X1 U17316 ( .A1(n41195), .A2(n41194), .ZN(n17471) );
  NAND2_X1 U17317 ( .A1(n3282), .A2(n983), .ZN(n18365) );
  NAND2_X1 U17321 ( .A1(n41868), .A2(n42211), .ZN(n9998) );
  NAND2_X1 U17322 ( .A1(n6626), .A2(n6624), .ZN(n6623) );
  AOI21_X1 U17323 ( .A1(n18741), .A2(n14965), .B(n40849), .ZN(n40851) );
  NAND2_X1 U17324 ( .A1(n40636), .A2(n38675), .ZN(n40639) );
  OAI21_X1 U17325 ( .A1(n41100), .A2(n40573), .B(n41113), .ZN(n4141) );
  OAI21_X1 U17327 ( .A1(n40390), .A2(n41083), .B(n14131), .ZN(n40391) );
  INV_X1 U17330 ( .I(n40346), .ZN(n18045) );
  NOR2_X1 U17331 ( .A1(n14616), .A2(n41384), .ZN(n13848) );
  INV_X1 U17337 ( .I(n2233), .ZN(n40241) );
  INV_X1 U17338 ( .I(n17077), .ZN(n37719) );
  NAND2_X1 U17340 ( .A1(n23890), .A2(n40557), .ZN(n14099) );
  NAND2_X1 U17342 ( .A1(n12466), .A2(n25246), .ZN(n10801) );
  NOR2_X1 U17344 ( .A1(n13050), .A2(n13049), .ZN(n13048) );
  AND2_X1 U17346 ( .A1(n21736), .A2(n25570), .Z(n16284) );
  NAND2_X1 U17347 ( .A1(n22617), .A2(n22913), .ZN(n13310) );
  NOR2_X1 U17349 ( .A1(n17212), .A2(n41376), .ZN(n13002) );
  OAI21_X1 U17351 ( .A1(n10936), .A2(n37061), .B(n61986), .ZN(n6754) );
  NAND2_X1 U17352 ( .A1(n40311), .A2(n17930), .ZN(n11045) );
  NAND2_X1 U17353 ( .A1(n12409), .A2(n40213), .ZN(n6626) );
  AOI21_X1 U17357 ( .A1(n41854), .A2(n12264), .B(n42507), .ZN(n39931) );
  AND2_X1 U17360 ( .A1(n40029), .A2(n40291), .Z(n39919) );
  AND2_X1 U17361 ( .A1(n59252), .A2(n7011), .Z(n3870) );
  AND2_X1 U17363 ( .A1(n57258), .A2(n64592), .Z(n12345) );
  NAND2_X1 U17364 ( .A1(n41425), .A2(n65184), .ZN(n5938) );
  OAI21_X1 U17365 ( .A1(n1748), .A2(n8688), .B(n18396), .ZN(n39834) );
  INV_X1 U17369 ( .I(n40727), .ZN(n41204) );
  INV_X1 U17370 ( .I(n42286), .ZN(n15051) );
  INV_X1 U17371 ( .I(n38049), .ZN(n40110) );
  NOR2_X1 U17372 ( .A1(n1272), .A2(n984), .ZN(n14655) );
  CLKBUF_X2 U17373 ( .I(n15258), .Z(n23967) );
  INV_X1 U17374 ( .I(n41928), .ZN(n7995) );
  NAND2_X1 U17375 ( .A1(n2867), .A2(n222), .ZN(n40584) );
  AND2_X1 U17376 ( .A1(n41400), .A2(n24523), .Z(n15345) );
  OR2_X1 U17379 ( .A1(n22502), .A2(n41906), .Z(n10670) );
  INV_X1 U17380 ( .I(n42215), .ZN(n21992) );
  NOR2_X1 U17381 ( .A1(n6260), .A2(n42453), .ZN(n6259) );
  NAND3_X1 U17382 ( .A1(n13169), .A2(n6058), .A3(n57207), .ZN(n41849) );
  AND2_X1 U17383 ( .A1(n40517), .A2(n21736), .Z(n15799) );
  NOR2_X1 U17384 ( .A1(n60139), .A2(n20984), .ZN(n41148) );
  NAND2_X1 U17385 ( .A1(n63849), .A2(n40582), .ZN(n40576) );
  OR2_X1 U17386 ( .A1(n40747), .A2(n40748), .Z(n40752) );
  NAND2_X1 U17387 ( .A1(n16306), .A2(n4359), .ZN(n4357) );
  NOR2_X1 U17388 ( .A1(n40061), .A2(n10479), .ZN(n38337) );
  INV_X1 U17390 ( .I(n41884), .ZN(n41063) );
  NAND2_X1 U17391 ( .A1(n40147), .A2(n59062), .ZN(n40148) );
  INV_X1 U17392 ( .I(n37934), .ZN(n40463) );
  AND2_X1 U17394 ( .A1(n41149), .A2(n1516), .Z(n16285) );
  INV_X1 U17396 ( .I(n11525), .ZN(n37593) );
  AND2_X1 U17401 ( .A1(n41163), .A2(n23884), .Z(n20637) );
  AND2_X1 U17402 ( .A1(n41122), .A2(n61638), .Z(n39993) );
  OR2_X1 U17403 ( .A1(n9790), .A2(n40595), .Z(n16306) );
  INV_X1 U17404 ( .I(n25777), .ZN(n41461) );
  OR2_X1 U17407 ( .A1(n42446), .A2(n11994), .Z(n11995) );
  NOR2_X1 U17408 ( .A1(n40641), .A2(n10587), .ZN(n7963) );
  AND2_X1 U17409 ( .A1(n59601), .A2(n41109), .Z(n16292) );
  NAND2_X1 U17410 ( .A1(n61950), .A2(n41411), .ZN(n15585) );
  INV_X1 U17412 ( .I(n40519), .ZN(n6348) );
  NAND2_X1 U17414 ( .A1(n64592), .A2(n41889), .ZN(n39791) );
  NAND2_X1 U17415 ( .A1(n6625), .A2(n10542), .ZN(n6624) );
  OR2_X1 U17416 ( .A1(n22776), .A2(n16680), .Z(n16171) );
  NOR2_X1 U17418 ( .A1(n23855), .A2(n4364), .ZN(n4489) );
  INV_X1 U17421 ( .I(n17349), .ZN(n38346) );
  AND3_X1 U17422 ( .A1(n22713), .A2(n16680), .A3(n22776), .Z(n16189) );
  NAND3_X1 U17423 ( .A1(n1512), .A2(n60928), .A3(n12523), .ZN(n22565) );
  INV_X1 U17424 ( .I(n40108), .ZN(n37463) );
  OR2_X1 U17427 ( .A1(n41255), .A2(n286), .Z(n40792) );
  AND2_X1 U17428 ( .A1(n971), .A2(n59601), .Z(n11819) );
  OR3_X1 U17430 ( .A1(n40944), .A2(n40949), .A3(n15558), .Z(n15915) );
  INV_X1 U17431 ( .I(n38604), .ZN(n40528) );
  NAND2_X1 U17432 ( .A1(n23616), .A2(n11787), .ZN(n38479) );
  CLKBUF_X2 U17433 ( .I(n38495), .Z(n22913) );
  INV_X1 U17434 ( .I(n38498), .ZN(n39092) );
  INV_X1 U17435 ( .I(n18338), .ZN(n39506) );
  NAND3_X1 U17441 ( .A1(n14863), .A2(n22285), .A3(n42427), .ZN(n15655) );
  AND2_X1 U17444 ( .A1(n40308), .A2(n1307), .Z(n1963) );
  INV_X1 U17445 ( .I(n1518), .ZN(n40075) );
  AND2_X1 U17446 ( .A1(n57208), .A2(n1517), .Z(n39920) );
  CLKBUF_X2 U17450 ( .I(n25920), .Z(n23298) );
  NOR2_X1 U17452 ( .A1(n61005), .A2(n10954), .ZN(n40142) );
  CLKBUF_X2 U17453 ( .I(n40294), .Z(n4364) );
  INV_X1 U17456 ( .I(n40087), .ZN(n1738) );
  CLKBUF_X2 U17459 ( .I(n3178), .Z(n9969) );
  BUF_X4 U17461 ( .I(n41165), .Z(n14462) );
  NAND2_X1 U17479 ( .A1(n64592), .A2(n64732), .ZN(n7511) );
  CLKBUF_X2 U17482 ( .I(n38480), .Z(n39146) );
  INV_X2 U17493 ( .I(n19065), .ZN(n38134) );
  INV_X1 U17495 ( .I(n39565), .ZN(n7106) );
  INV_X1 U17503 ( .I(n37842), .ZN(n13220) );
  INV_X1 U17505 ( .I(n39627), .ZN(n20533) );
  INV_X1 U17506 ( .I(n6749), .ZN(n1994) );
  INV_X1 U17507 ( .I(n38245), .ZN(n25248) );
  INV_X1 U17508 ( .I(n37496), .ZN(n4147) );
  INV_X1 U17509 ( .I(n38859), .ZN(n38484) );
  INV_X1 U17510 ( .I(n39647), .ZN(n10356) );
  INV_X1 U17512 ( .I(n9805), .ZN(n6997) );
  INV_X1 U17516 ( .I(n38319), .ZN(n2870) );
  INV_X1 U17518 ( .I(n3753), .ZN(n39239) );
  INV_X1 U17519 ( .I(n39290), .ZN(n6160) );
  BUF_X2 U17520 ( .I(n19441), .Z(n3479) );
  INV_X1 U17521 ( .I(n37727), .ZN(n14696) );
  INV_X2 U17523 ( .I(n12980), .ZN(n1749) );
  INV_X1 U17525 ( .I(n38621), .ZN(n2107) );
  INV_X1 U17528 ( .I(n39372), .ZN(n8234) );
  INV_X1 U17529 ( .I(n24435), .ZN(n9121) );
  INV_X1 U17534 ( .I(n25995), .ZN(n5973) );
  INV_X1 U17536 ( .I(n25161), .ZN(n24468) );
  INV_X1 U17537 ( .I(n38175), .ZN(n5822) );
  INV_X1 U17541 ( .I(n37888), .ZN(n9412) );
  INV_X1 U17542 ( .I(n38361), .ZN(n3277) );
  INV_X1 U17543 ( .I(n19381), .ZN(n8205) );
  BUF_X2 U17544 ( .I(n37697), .Z(n17594) );
  BUF_X2 U17545 ( .I(n37802), .Z(n16449) );
  INV_X1 U17547 ( .I(n38987), .ZN(n38986) );
  INV_X1 U17548 ( .I(n14553), .ZN(n22344) );
  INV_X1 U17549 ( .I(n37553), .ZN(n1753) );
  INV_X1 U17550 ( .I(n18132), .ZN(n38105) );
  INV_X1 U17551 ( .I(n38364), .ZN(n9362) );
  INV_X1 U17552 ( .I(n39564), .ZN(n4395) );
  CLKBUF_X2 U17553 ( .I(n16632), .Z(n22535) );
  AND2_X1 U17554 ( .A1(n12171), .A2(n1523), .Z(n5479) );
  INV_X1 U17555 ( .I(n38807), .ZN(n13905) );
  INV_X1 U17557 ( .I(n18268), .ZN(n38220) );
  BUF_X2 U17565 ( .I(n39586), .Z(n5779) );
  INV_X1 U17566 ( .I(n39562), .ZN(n39563) );
  INV_X1 U17567 ( .I(n38968), .ZN(n1909) );
  INV_X1 U17569 ( .I(n38253), .ZN(n1755) );
  INV_X1 U17571 ( .I(n62852), .ZN(n10780) );
  NAND2_X1 U17572 ( .A1(n2319), .A2(n2318), .ZN(n37820) );
  CLKBUF_X2 U17573 ( .I(n38286), .Z(n9269) );
  CLKBUF_X2 U17574 ( .I(n38123), .Z(n23332) );
  CLKBUF_X2 U17575 ( .I(n39386), .Z(n22697) );
  INV_X1 U17576 ( .I(n3480), .ZN(n15664) );
  INV_X1 U17578 ( .I(n15704), .ZN(n8601) );
  INV_X1 U17580 ( .I(n10351), .ZN(n2682) );
  INV_X1 U17583 ( .I(n37726), .ZN(n13618) );
  INV_X1 U17586 ( .I(n22988), .ZN(n3752) );
  NOR2_X1 U17587 ( .A1(n10804), .A2(n18991), .ZN(n6731) );
  CLKBUF_X2 U17589 ( .I(n36298), .Z(n22480) );
  INV_X1 U17591 ( .I(n2320), .ZN(n2319) );
  CLKBUF_X2 U17592 ( .I(n38304), .Z(n20087) );
  INV_X1 U17593 ( .I(n9931), .ZN(n12128) );
  AOI21_X1 U17594 ( .A1(n14891), .A2(n14894), .B(n38993), .ZN(n8233) );
  INV_X1 U17595 ( .I(n57836), .ZN(n8684) );
  INV_X1 U17600 ( .I(n13321), .ZN(n11792) );
  INV_X1 U17601 ( .I(n15579), .ZN(n39206) );
  INV_X1 U17602 ( .I(n39276), .ZN(n38867) );
  INV_X2 U17603 ( .I(n21688), .ZN(n1760) );
  NAND2_X1 U17604 ( .A1(n14909), .A2(n14908), .ZN(n3399) );
  INV_X1 U17605 ( .I(n38325), .ZN(n8149) );
  CLKBUF_X2 U17607 ( .I(n38188), .Z(n22916) );
  INV_X1 U17609 ( .I(n39527), .ZN(n9922) );
  NAND2_X1 U17616 ( .A1(n10671), .A2(n36263), .ZN(n2685) );
  OAI21_X1 U17619 ( .A1(n36164), .A2(n24366), .B(n37364), .ZN(n6836) );
  NAND2_X1 U17620 ( .A1(n37494), .A2(n34850), .ZN(n18991) );
  INV_X1 U17621 ( .I(n18671), .ZN(n18670) );
  INV_X2 U17623 ( .I(n19261), .ZN(n1762) );
  NAND2_X1 U17627 ( .A1(n4510), .A2(n4509), .ZN(n10803) );
  NAND2_X1 U17629 ( .A1(n15581), .A2(n15580), .ZN(n15579) );
  INV_X1 U17630 ( .I(n24018), .ZN(n14590) );
  NOR2_X1 U17631 ( .A1(n23750), .A2(n23748), .ZN(n32156) );
  NOR2_X1 U17633 ( .A1(n24627), .A2(n17960), .ZN(n24626) );
  NOR2_X1 U17640 ( .A1(n6770), .A2(n35460), .ZN(n5383) );
  NAND2_X1 U17641 ( .A1(n37961), .A2(n62010), .ZN(n15580) );
  AOI21_X1 U17642 ( .A1(n15583), .A2(n15582), .B(n39524), .ZN(n15581) );
  AND2_X1 U17644 ( .A1(n36065), .A2(n17197), .Z(n17196) );
  NAND2_X1 U17650 ( .A1(n35728), .A2(n57542), .ZN(n5558) );
  INV_X1 U17651 ( .I(n39230), .ZN(n10813) );
  NAND2_X1 U17652 ( .A1(n8763), .A2(n8762), .ZN(n8761) );
  NOR3_X1 U17656 ( .A1(n37332), .A2(n37331), .A3(n37330), .ZN(n37346) );
  AOI21_X1 U17657 ( .A1(n8861), .A2(n8859), .B(n8858), .ZN(n36880) );
  NAND2_X1 U17660 ( .A1(n9086), .A2(n26243), .ZN(n15970) );
  AND3_X1 U17664 ( .A1(n32449), .A2(n32448), .A3(n32450), .Z(n7714) );
  INV_X1 U17665 ( .I(n12879), .ZN(n12860) );
  NOR2_X1 U17668 ( .A1(n21773), .A2(n34856), .ZN(n18990) );
  OAI21_X1 U17669 ( .A1(n36411), .A2(n14688), .B(n55), .ZN(n14687) );
  NAND2_X1 U17673 ( .A1(n36333), .A2(n36820), .ZN(n13996) );
  NAND2_X1 U17675 ( .A1(n35362), .A2(n18312), .ZN(n35365) );
  NAND3_X1 U17684 ( .A1(n4499), .A2(n34487), .A3(n19064), .ZN(n21674) );
  AOI21_X1 U17685 ( .A1(n4834), .A2(n37192), .B(n37191), .ZN(n37193) );
  OAI21_X1 U17689 ( .A1(n4009), .A2(n20373), .B(n36552), .ZN(n3999) );
  OAI21_X1 U17693 ( .A1(n11730), .A2(n57275), .B(n10394), .ZN(n11728) );
  NOR2_X1 U17695 ( .A1(n37005), .A2(n37004), .ZN(n22954) );
  INV_X1 U17698 ( .I(n8976), .ZN(n35268) );
  INV_X1 U17700 ( .I(n37129), .ZN(n6630) );
  NAND2_X1 U17701 ( .A1(n36259), .A2(n35183), .ZN(n34107) );
  NAND2_X1 U17702 ( .A1(n11040), .A2(n21675), .ZN(n4499) );
  NOR2_X1 U17703 ( .A1(n18616), .A2(n18614), .ZN(n18613) );
  NOR2_X1 U17704 ( .A1(n21742), .A2(n21741), .ZN(n21544) );
  NOR2_X1 U17705 ( .A1(n12834), .A2(n35604), .ZN(n14029) );
  OAI22_X1 U17706 ( .A1(n36177), .A2(n21615), .B1(n36430), .B2(n36173), .ZN(
        n8546) );
  NOR2_X1 U17707 ( .A1(n37098), .A2(n37097), .ZN(n11753) );
  AOI22_X1 U17708 ( .A1(n34111), .A2(n34108), .B1(n34110), .B2(n34109), .ZN(
        n34112) );
  NAND2_X1 U17713 ( .A1(n36117), .A2(n4263), .ZN(n8763) );
  NOR2_X1 U17717 ( .A1(n34287), .A2(n34286), .ZN(n8637) );
  INV_X1 U17718 ( .I(n35878), .ZN(n5462) );
  NOR2_X1 U17728 ( .A1(n32149), .A2(n8010), .ZN(n23749) );
  OAI21_X1 U17729 ( .A1(n34202), .A2(n35986), .B(n36706), .ZN(n34207) );
  INV_X1 U17731 ( .I(n36409), .ZN(n14688) );
  OAI21_X1 U17734 ( .A1(n37286), .A2(n25187), .B(n16153), .ZN(n34459) );
  NAND2_X1 U17736 ( .A1(n7759), .A2(n37222), .ZN(n37223) );
  AOI21_X1 U17739 ( .A1(n34492), .A2(n685), .B(n34493), .ZN(n34494) );
  AOI21_X1 U17740 ( .A1(n63900), .A2(n36761), .B(n36760), .ZN(n6834) );
  AOI22_X1 U17741 ( .A1(n36642), .A2(n36641), .B1(n36640), .B2(n20251), .ZN(
        n36643) );
  NAND2_X1 U17743 ( .A1(n37495), .A2(n37489), .ZN(n10804) );
  NAND2_X1 U17745 ( .A1(n37189), .A2(n24658), .ZN(n37191) );
  INV_X1 U17748 ( .I(n36260), .ZN(n2683) );
  NOR2_X1 U17749 ( .A1(n17193), .A2(n32858), .ZN(n5385) );
  NOR2_X1 U17750 ( .A1(n37244), .A2(n13647), .ZN(n14485) );
  OAI21_X1 U17753 ( .A1(n17144), .A2(n3764), .B(n3763), .ZN(n3762) );
  NAND2_X1 U17754 ( .A1(n20793), .A2(n9869), .ZN(n5556) );
  NOR3_X1 U17755 ( .A1(n2628), .A2(n37410), .A3(n36834), .ZN(n8099) );
  NAND2_X1 U17758 ( .A1(n18061), .A2(n36600), .ZN(n25294) );
  NAND2_X1 U17759 ( .A1(n37312), .A2(n2242), .ZN(n10556) );
  AOI21_X1 U17762 ( .A1(n6050), .A2(n21148), .B(n6049), .ZN(n21146) );
  NAND2_X1 U17763 ( .A1(n35485), .A2(n14914), .ZN(n31547) );
  NAND2_X1 U17764 ( .A1(n36184), .A2(n14264), .ZN(n36187) );
  INV_X1 U17767 ( .I(n19677), .ZN(n37287) );
  AOI22_X1 U17770 ( .A1(n19347), .A2(n37336), .B1(n37337), .B2(n37338), .ZN(
        n37345) );
  OAI22_X1 U17771 ( .A1(n6985), .A2(n37400), .B1(n6984), .B2(n36332), .ZN(
        n36333) );
  NOR2_X1 U17772 ( .A1(n1308), .A2(n10708), .ZN(n10707) );
  INV_X1 U17774 ( .I(n36156), .ZN(n15161) );
  OAI22_X1 U17775 ( .A1(n37391), .A2(n8808), .B1(n36865), .B2(n16885), .ZN(
        n35339) );
  NAND2_X1 U17776 ( .A1(n36899), .A2(n36057), .ZN(n35386) );
  OAI21_X1 U17777 ( .A1(n34928), .A2(n35954), .B(n62041), .ZN(n3156) );
  NAND2_X1 U17779 ( .A1(n8039), .A2(n8520), .ZN(n9836) );
  AOI21_X1 U17781 ( .A1(n35927), .A2(n36866), .B(n37387), .ZN(n35928) );
  NOR2_X1 U17783 ( .A1(n36913), .A2(n37423), .ZN(n8636) );
  NOR2_X1 U17786 ( .A1(n36364), .A2(n25775), .ZN(n7725) );
  NAND2_X1 U17788 ( .A1(n37027), .A2(n37026), .ZN(n25343) );
  INV_X1 U17789 ( .I(n36672), .ZN(n5287) );
  NAND2_X1 U17793 ( .A1(n3234), .A2(n11272), .ZN(n3316) );
  NAND2_X1 U17795 ( .A1(n9842), .A2(n12899), .ZN(n20309) );
  OAI21_X1 U17800 ( .A1(n36329), .A2(n6540), .B(n37410), .ZN(n35263) );
  AOI21_X1 U17801 ( .A1(n36004), .A2(n36003), .B(n36002), .ZN(n36005) );
  NAND2_X1 U17803 ( .A1(n21881), .A2(n37389), .ZN(n5871) );
  NAND2_X1 U17805 ( .A1(n25489), .A2(n64405), .ZN(n25488) );
  OAI21_X1 U17806 ( .A1(n35566), .A2(n35565), .B(n16690), .ZN(n13302) );
  NOR2_X1 U17807 ( .A1(n14753), .A2(n11564), .ZN(n11563) );
  INV_X1 U17808 ( .I(n36093), .ZN(n36091) );
  NAND2_X1 U17812 ( .A1(n8102), .A2(n36835), .ZN(n2628) );
  INV_X1 U17813 ( .I(n16027), .ZN(n23471) );
  NOR2_X1 U17814 ( .A1(n35488), .A2(n14298), .ZN(n12494) );
  INV_X1 U17815 ( .I(n11302), .ZN(n11301) );
  OAI22_X1 U17818 ( .A1(n37243), .A2(n37249), .B1(n37240), .B2(n13647), .ZN(
        n14445) );
  AOI22_X1 U17819 ( .A1(n36438), .A2(n36439), .B1(n61940), .B2(n36440), .ZN(
        n10394) );
  INV_X1 U17820 ( .I(n18811), .ZN(n36957) );
  NOR2_X1 U17825 ( .A1(n15191), .A2(n15192), .ZN(n15178) );
  AND2_X1 U17826 ( .A1(n20530), .A2(n20531), .Z(n20373) );
  NOR2_X1 U17829 ( .A1(n35162), .A2(n15036), .ZN(n32440) );
  NOR2_X1 U17831 ( .A1(n12882), .A2(n10484), .ZN(n12861) );
  NAND2_X1 U17833 ( .A1(n35556), .A2(n10413), .ZN(n11040) );
  AOI21_X1 U17835 ( .A1(n11722), .A2(n35534), .B(n11720), .ZN(n36095) );
  NOR2_X1 U17836 ( .A1(n33669), .A2(n35142), .ZN(n6050) );
  INV_X1 U17840 ( .I(n36828), .ZN(n36826) );
  NOR2_X1 U17842 ( .A1(n31542), .A2(n20433), .ZN(n20432) );
  OR2_X1 U17843 ( .A1(n36329), .A2(n8195), .Z(n20790) );
  INV_X1 U17852 ( .I(n36109), .ZN(n35360) );
  NAND3_X1 U17853 ( .A1(n34474), .A2(n35147), .A3(n35962), .ZN(n4308) );
  INV_X1 U17855 ( .I(n35503), .ZN(n4980) );
  NAND2_X1 U17856 ( .A1(n32910), .A2(n32911), .ZN(n4981) );
  OR2_X1 U17857 ( .A1(n18313), .A2(n36193), .Z(n18312) );
  NAND2_X1 U17861 ( .A1(n4571), .A2(n20530), .ZN(n4006) );
  NAND2_X1 U17862 ( .A1(n20783), .A2(n36961), .ZN(n12489) );
  NAND2_X1 U17864 ( .A1(n4853), .A2(n4852), .ZN(n36015) );
  NAND2_X1 U17865 ( .A1(n17660), .A2(n36821), .ZN(n6985) );
  NAND2_X1 U17867 ( .A1(n7805), .A2(n7803), .ZN(n31788) );
  NAND2_X1 U17868 ( .A1(n35446), .A2(n12572), .ZN(n12571) );
  NAND2_X1 U17869 ( .A1(n3471), .A2(n17596), .ZN(n36876) );
  INV_X1 U17870 ( .I(n35608), .ZN(n35348) );
  INV_X1 U17873 ( .I(n36213), .ZN(n14243) );
  NAND2_X1 U17877 ( .A1(n36114), .A2(n22474), .ZN(n8760) );
  NOR2_X1 U17878 ( .A1(n37958), .A2(n15582), .ZN(n35484) );
  AND2_X1 U17879 ( .A1(n36412), .A2(n36193), .Z(n36113) );
  AOI21_X1 U17880 ( .A1(n576), .A2(n36027), .B(n35583), .ZN(n17193) );
  INV_X1 U17881 ( .I(n21912), .ZN(n21911) );
  AOI21_X1 U17883 ( .A1(n33457), .A2(n36893), .B(n24310), .ZN(n24309) );
  NAND2_X1 U17885 ( .A1(n21880), .A2(n10765), .ZN(n35335) );
  NOR2_X1 U17888 ( .A1(n34929), .A2(n59229), .ZN(n15191) );
  INV_X1 U17890 ( .I(n11780), .ZN(n11778) );
  AND3_X1 U17892 ( .A1(n3907), .A2(n11273), .A3(n11271), .Z(n36155) );
  NAND2_X1 U17893 ( .A1(n11835), .A2(n24356), .ZN(n11833) );
  AND2_X1 U17894 ( .A1(n34925), .A2(n63406), .Z(n23601) );
  NAND2_X1 U17895 ( .A1(n32816), .A2(n23626), .ZN(n32855) );
  INV_X1 U17897 ( .I(n11271), .ZN(n3234) );
  NAND2_X1 U17900 ( .A1(n34920), .A2(n7682), .ZN(n11836) );
  NOR2_X1 U17903 ( .A1(n2094), .A2(n2093), .ZN(n2092) );
  NOR2_X1 U17905 ( .A1(n36172), .A2(n60949), .ZN(n8547) );
  NAND2_X1 U17906 ( .A1(n36424), .A2(n2761), .ZN(n8549) );
  INV_X1 U17909 ( .I(n4680), .ZN(n4679) );
  INV_X1 U17910 ( .I(n37187), .ZN(n17537) );
  NAND3_X1 U17912 ( .A1(n59809), .A2(n59147), .A3(n2418), .ZN(n34806) );
  NOR2_X1 U17915 ( .A1(n34934), .A2(n36725), .ZN(n9769) );
  AND3_X1 U17917 ( .A1(n35548), .A2(n35966), .A3(n23577), .Z(n16114) );
  NOR2_X1 U17922 ( .A1(n60196), .A2(n18144), .ZN(n36391) );
  OAI21_X1 U17924 ( .A1(n36140), .A2(n34577), .B(n36801), .ZN(n34578) );
  NOR2_X1 U17927 ( .A1(n35445), .A2(n13983), .ZN(n12572) );
  INV_X1 U17929 ( .I(n16054), .ZN(n11337) );
  NAND2_X1 U17931 ( .A1(n21771), .A2(n10165), .ZN(n4509) );
  NOR2_X1 U17932 ( .A1(n16268), .A2(n18130), .ZN(n21672) );
  NAND2_X1 U17933 ( .A1(n57656), .A2(n2057), .ZN(n23241) );
  NOR2_X1 U17934 ( .A1(n5976), .A2(n18969), .ZN(n5975) );
  NOR2_X1 U17936 ( .A1(n34097), .A2(n3217), .ZN(n34098) );
  NAND2_X1 U17938 ( .A1(n36495), .A2(n12408), .ZN(n12407) );
  AND2_X1 U17939 ( .A1(n37354), .A2(n37293), .Z(n11221) );
  NAND2_X1 U17941 ( .A1(n36461), .A2(n64087), .ZN(n3315) );
  NAND2_X1 U17944 ( .A1(n39523), .A2(n37957), .ZN(n15583) );
  INV_X1 U17945 ( .I(n37044), .ZN(n35100) );
  AND2_X1 U17948 ( .A1(n14915), .A2(n58026), .Z(n14914) );
  INV_X1 U17949 ( .I(n36431), .ZN(n14685) );
  NOR2_X1 U17951 ( .A1(n9494), .A2(n36926), .ZN(n7429) );
  NOR2_X1 U17952 ( .A1(n33783), .A2(n18615), .ZN(n18614) );
  AOI21_X1 U17959 ( .A1(n36892), .A2(n36891), .B(n5524), .ZN(n5523) );
  AOI21_X1 U17961 ( .A1(n34862), .A2(n20431), .B(n7861), .ZN(n24010) );
  NAND2_X1 U17962 ( .A1(n36942), .A2(n6167), .ZN(n11756) );
  INV_X1 U17964 ( .I(n36049), .ZN(n10708) );
  NAND2_X1 U17965 ( .A1(n24660), .A2(n11811), .ZN(n37337) );
  NAND2_X1 U17967 ( .A1(n8363), .A2(n36239), .ZN(n4495) );
  NAND2_X1 U17968 ( .A1(n1415), .A2(n36257), .ZN(n36258) );
  INV_X1 U17970 ( .I(n9947), .ZN(n14298) );
  OAI22_X1 U17971 ( .A1(n64181), .A2(n32977), .B1(n32978), .B2(n22785), .ZN(
        n25489) );
  INV_X1 U17972 ( .I(n36967), .ZN(n36970) );
  NOR2_X1 U17973 ( .A1(n37333), .A2(n12301), .ZN(n37338) );
  NAND2_X1 U17976 ( .A1(n60980), .A2(n9783), .ZN(n37373) );
  NAND3_X1 U17977 ( .A1(n3588), .A2(n60659), .A3(n22524), .ZN(n1911) );
  AND2_X1 U17979 ( .A1(n35900), .A2(n24118), .Z(n34492) );
  NAND2_X1 U17982 ( .A1(n10067), .A2(n1415), .ZN(n34109) );
  NAND3_X1 U17986 ( .A1(n34094), .A2(n34093), .A3(n34092), .ZN(n34095) );
  OR2_X1 U17987 ( .A1(n1525), .A2(n10413), .Z(n35557) );
  OAI21_X1 U17988 ( .A1(n12863), .A2(n14189), .B(n36748), .ZN(n20281) );
  OR2_X1 U17990 ( .A1(n22461), .A2(n34815), .Z(n3764) );
  AND2_X1 U17993 ( .A1(n35447), .A2(n36959), .Z(n20783) );
  INV_X1 U17997 ( .I(n13647), .ZN(n37442) );
  AND2_X1 U17999 ( .A1(n23842), .A2(n18969), .Z(n18983) );
  OAI21_X1 U18000 ( .A1(n24041), .A2(n6984), .B(n10550), .ZN(n37412) );
  NOR2_X1 U18003 ( .A1(n36921), .A2(n36926), .ZN(n32906) );
  NOR2_X1 U18005 ( .A1(n10226), .A2(n64620), .ZN(n16192) );
  INV_X1 U18008 ( .I(n35607), .ZN(n36730) );
  INV_X1 U18009 ( .I(n37132), .ZN(n5978) );
  INV_X1 U18010 ( .I(n7656), .ZN(n35598) );
  NOR2_X1 U18011 ( .A1(n18048), .A2(n10829), .ZN(n32772) );
  INV_X1 U18012 ( .I(n36626), .ZN(n35056) );
  AOI21_X1 U18013 ( .A1(n36460), .A2(n36152), .B(n60462), .ZN(n2301) );
  NAND2_X1 U18016 ( .A1(n57209), .A2(n8438), .ZN(n7446) );
  INV_X1 U18017 ( .I(n5483), .ZN(n6713) );
  OAI21_X1 U18018 ( .A1(n36956), .A2(n1781), .B(n60694), .ZN(n36958) );
  NOR2_X1 U18019 ( .A1(n36966), .A2(n63643), .ZN(n11592) );
  CLKBUF_X2 U18020 ( .I(n36394), .Z(n22454) );
  NOR2_X1 U18021 ( .A1(n35910), .A2(n37035), .ZN(n3588) );
  INV_X1 U18022 ( .I(n34821), .ZN(n32816) );
  INV_X1 U18023 ( .I(n8132), .ZN(n35927) );
  NAND2_X1 U18024 ( .A1(n61066), .A2(n36040), .ZN(n32859) );
  INV_X1 U18026 ( .I(n3460), .ZN(n4036) );
  NAND2_X1 U18027 ( .A1(n34908), .A2(n1421), .ZN(n33449) );
  INV_X1 U18029 ( .I(n35507), .ZN(n35504) );
  INV_X1 U18030 ( .I(n2792), .ZN(n34925) );
  NOR2_X1 U18031 ( .A1(n34930), .A2(n35506), .ZN(n15192) );
  INV_X1 U18034 ( .I(n37289), .ZN(n37104) );
  NOR2_X1 U18035 ( .A1(n36890), .A2(n1421), .ZN(n5524) );
  NAND2_X1 U18036 ( .A1(n35066), .A2(n35067), .ZN(n4654) );
  NOR2_X1 U18038 ( .A1(n12004), .A2(n1417), .ZN(n35070) );
  INV_X1 U18040 ( .I(n21802), .ZN(n36428) );
  INV_X1 U18041 ( .I(n20951), .ZN(n12458) );
  INV_X1 U18044 ( .I(n25163), .ZN(n36172) );
  AND2_X1 U18045 ( .A1(n8356), .A2(n4035), .Z(n11722) );
  NAND2_X1 U18046 ( .A1(n37334), .A2(n8010), .ZN(n6123) );
  AND2_X1 U18050 ( .A1(n61180), .A2(n20147), .Z(n35982) );
  OAI21_X1 U18051 ( .A1(n61940), .A2(n7656), .B(n36434), .ZN(n34704) );
  INV_X1 U18052 ( .I(n36597), .ZN(n36507) );
  NAND2_X1 U18054 ( .A1(n36310), .A2(n57211), .ZN(n36141) );
  OAI21_X1 U18055 ( .A1(n36374), .A2(n23677), .B(n36096), .ZN(n36101) );
  INV_X1 U18058 ( .I(n35387), .ZN(n35389) );
  NOR2_X1 U18060 ( .A1(n62041), .A2(n1777), .ZN(n35953) );
  NAND2_X1 U18064 ( .A1(n12393), .A2(n2885), .ZN(n36134) );
  NOR2_X1 U18067 ( .A1(n34927), .A2(n24198), .ZN(n4305) );
  INV_X1 U18070 ( .I(n36924), .ZN(n11564) );
  AND2_X1 U18073 ( .A1(n36262), .A2(n63897), .Z(n34108) );
  AND2_X1 U18074 ( .A1(n3218), .A2(n7933), .Z(n3217) );
  INV_X1 U18075 ( .I(n36340), .ZN(n35068) );
  NAND2_X1 U18079 ( .A1(n3218), .A2(n22113), .ZN(n2093) );
  INV_X1 U18081 ( .I(n35404), .ZN(n35493) );
  AND2_X1 U18084 ( .A1(n5936), .A2(n1421), .Z(n11393) );
  NAND2_X1 U18090 ( .A1(n37359), .A2(n19573), .ZN(n37360) );
  AND2_X1 U18093 ( .A1(n64609), .A2(n22524), .Z(n15831) );
  INV_X1 U18096 ( .I(n34077), .ZN(n36745) );
  NAND2_X1 U18098 ( .A1(n1777), .A2(n34927), .ZN(n32895) );
  AND2_X1 U18100 ( .A1(n36151), .A2(n60462), .Z(n10789) );
  OR2_X1 U18102 ( .A1(n2958), .A2(n37335), .Z(n11811) );
  NOR2_X1 U18103 ( .A1(n35860), .A2(n14189), .ZN(n35864) );
  OR2_X1 U18104 ( .A1(n36344), .A2(n17364), .Z(n12881) );
  OR2_X1 U18105 ( .A1(n36483), .A2(n10829), .Z(n12408) );
  OR2_X1 U18106 ( .A1(n3218), .A2(n59379), .Z(n3789) );
  INV_X1 U18107 ( .I(n36171), .ZN(n36419) );
  NOR2_X1 U18108 ( .A1(n35532), .A2(n36555), .ZN(n36564) );
  INV_X1 U18109 ( .I(n36252), .ZN(n1775) );
  NAND2_X1 U18110 ( .A1(n10498), .A2(n36470), .ZN(n36474) );
  INV_X1 U18112 ( .I(n36441), .ZN(n36450) );
  INV_X2 U18114 ( .I(n17132), .ZN(n2958) );
  AND2_X1 U18123 ( .A1(n22113), .A2(n10498), .Z(n36154) );
  NAND2_X1 U18136 ( .A1(n10498), .A2(n1217), .ZN(n2719) );
  INV_X4 U18144 ( .I(n24249), .ZN(n37363) );
  INV_X1 U18150 ( .I(n37184), .ZN(n6779) );
  INV_X2 U18153 ( .I(n24365), .ZN(n22317) );
  NOR2_X1 U18162 ( .A1(n16234), .A2(n15821), .ZN(n21781) );
  NAND2_X1 U18165 ( .A1(n33535), .A2(n59121), .ZN(n12748) );
  NAND3_X1 U18166 ( .A1(n31953), .A2(n31952), .A3(n35315), .ZN(n10495) );
  AND2_X1 U18168 ( .A1(n35361), .A2(n36193), .Z(n33608) );
  NAND2_X1 U18172 ( .A1(n10640), .A2(n10639), .ZN(n31525) );
  NOR2_X1 U18174 ( .A1(n18933), .A2(n18932), .ZN(n22073) );
  INV_X1 U18175 ( .I(n4249), .ZN(n33813) );
  NOR2_X1 U18177 ( .A1(n3994), .A2(n63624), .ZN(n32815) );
  NAND2_X1 U18187 ( .A1(n35257), .A2(n35261), .ZN(n6541) );
  NOR2_X1 U18188 ( .A1(n19449), .A2(n19448), .ZN(n21278) );
  AOI22_X1 U18192 ( .A1(n12514), .A2(n19457), .B1(n12511), .B2(n33775), .ZN(
        n12817) );
  INV_X1 U18195 ( .I(n34472), .ZN(n11319) );
  OAI21_X1 U18200 ( .A1(n16990), .A2(n16145), .B(n16989), .ZN(n10698) );
  AOI22_X1 U18210 ( .A1(n35808), .A2(n35809), .B1(n35810), .B2(n11186), .ZN(
        n20596) );
  AOI21_X1 U18212 ( .A1(n10632), .A2(n33703), .B(n33351), .ZN(n33352) );
  NOR2_X1 U18213 ( .A1(n35312), .A2(n35259), .ZN(n12011) );
  NAND2_X1 U18214 ( .A1(n26229), .A2(n16243), .ZN(n24497) );
  NOR2_X1 U18215 ( .A1(n34441), .A2(n35764), .ZN(n12012) );
  NAND2_X1 U18223 ( .A1(n4891), .A2(n7317), .ZN(n32786) );
  INV_X1 U18224 ( .I(n19240), .ZN(n10640) );
  NOR2_X1 U18226 ( .A1(n35029), .A2(n14246), .ZN(n14245) );
  NOR2_X1 U18228 ( .A1(n57294), .A2(n11181), .ZN(n13405) );
  OR2_X1 U18230 ( .A1(n31778), .A2(n10277), .Z(n16198) );
  OAI21_X1 U18231 ( .A1(n33927), .A2(n35777), .B(n5583), .ZN(n5582) );
  INV_X1 U18236 ( .I(n20062), .ZN(n20061) );
  NAND2_X1 U18238 ( .A1(n2308), .A2(n20660), .ZN(n2307) );
  AOI21_X1 U18239 ( .A1(n18243), .A2(n18244), .B(n57172), .ZN(n16096) );
  NOR2_X1 U18242 ( .A1(n35281), .A2(n63163), .ZN(n21765) );
  NOR2_X1 U18243 ( .A1(n34768), .A2(n34769), .ZN(n25910) );
  NAND2_X1 U18244 ( .A1(n35631), .A2(n7342), .ZN(n32681) );
  OAI21_X1 U18245 ( .A1(n33533), .A2(n33532), .B(n6398), .ZN(n6397) );
  OAI21_X1 U18246 ( .A1(n25900), .A2(n15574), .B(n15573), .ZN(n15572) );
  OAI22_X1 U18247 ( .A1(n1541), .A2(n2908), .B1(n19265), .B2(n904), .ZN(n34412) );
  NOR2_X1 U18249 ( .A1(n33403), .A2(n3549), .ZN(n3548) );
  OAI21_X1 U18253 ( .A1(n35334), .A2(n22835), .B(n25946), .ZN(n11668) );
  NOR2_X1 U18257 ( .A1(n34293), .A2(n34227), .ZN(n2386) );
  NOR2_X1 U18258 ( .A1(n17071), .A2(n17070), .ZN(n17069) );
  NOR2_X1 U18260 ( .A1(n32460), .A2(n33611), .ZN(n11349) );
  OAI21_X1 U18261 ( .A1(n5083), .A2(n5084), .B(n58998), .ZN(n4430) );
  NAND2_X1 U18264 ( .A1(n19444), .A2(n19443), .ZN(n22297) );
  AOI22_X1 U18265 ( .A1(n13851), .A2(n34334), .B1(n13850), .B2(n33925), .ZN(
        n16727) );
  NOR2_X1 U18266 ( .A1(n18647), .A2(n15143), .ZN(n15142) );
  NAND2_X1 U18267 ( .A1(n8115), .A2(n8114), .ZN(n17427) );
  BUF_X4 U18268 ( .I(n29875), .Z(n1793) );
  OR2_X1 U18273 ( .A1(n445), .A2(n18180), .Z(n18179) );
  NAND3_X1 U18274 ( .A1(n34710), .A2(n35818), .A3(n21485), .ZN(n21484) );
  OAI21_X1 U18278 ( .A1(n9797), .A2(n9796), .B(n7359), .ZN(n33706) );
  NAND2_X1 U18283 ( .A1(n35788), .A2(n5874), .ZN(n35789) );
  NAND2_X1 U18286 ( .A1(n4639), .A2(n33339), .ZN(n15287) );
  NAND2_X1 U18289 ( .A1(n34180), .A2(n14913), .ZN(n34181) );
  NAND2_X1 U18291 ( .A1(n12776), .A2(n34273), .ZN(n13127) );
  AOI22_X1 U18299 ( .A1(n11401), .A2(n11402), .B1(n57165), .B2(n11403), .ZN(
        n11400) );
  INV_X1 U18302 ( .I(n34300), .ZN(n35278) );
  INV_X1 U18303 ( .I(n25196), .ZN(n10118) );
  NOR2_X1 U18304 ( .A1(n32428), .A2(n21455), .ZN(n11542) );
  NAND2_X1 U18308 ( .A1(n34960), .A2(n32918), .ZN(n9278) );
  OAI21_X1 U18313 ( .A1(n4911), .A2(n34445), .B(n34444), .ZN(n16729) );
  OAI21_X1 U18314 ( .A1(n9127), .A2(n5477), .B(n9125), .ZN(n9129) );
  NAND2_X1 U18315 ( .A1(n34638), .A2(n61449), .ZN(n34650) );
  NAND2_X1 U18317 ( .A1(n14669), .A2(n32887), .ZN(n3130) );
  OAI21_X1 U18322 ( .A1(n35615), .A2(n58533), .B(n22976), .ZN(n35641) );
  AOI21_X1 U18323 ( .A1(n17548), .A2(n17547), .B(n4892), .ZN(n4891) );
  NAND3_X1 U18327 ( .A1(n33967), .A2(n9542), .A3(n118), .ZN(n9539) );
  INV_X1 U18331 ( .I(n16919), .ZN(n18801) );
  NAND2_X1 U18332 ( .A1(n34318), .A2(n35826), .ZN(n22642) );
  NAND2_X1 U18333 ( .A1(n5159), .A2(n1312), .ZN(n5162) );
  NAND2_X1 U18335 ( .A1(n7415), .A2(n7414), .ZN(n14246) );
  AOI22_X1 U18337 ( .A1(n33438), .A2(n8005), .B1(n64283), .B2(n4075), .ZN(
        n16422) );
  OAI22_X1 U18339 ( .A1(n33944), .A2(n33945), .B1(n2695), .B2(n34116), .ZN(
        n33952) );
  OAI21_X1 U18340 ( .A1(n20064), .A2(n20063), .B(n33951), .ZN(n20062) );
  AOI22_X1 U18341 ( .A1(n20923), .A2(n32847), .B1(n34146), .B2(n64100), .ZN(
        n32852) );
  INV_X1 U18342 ( .I(n20955), .ZN(n9720) );
  NOR2_X1 U18343 ( .A1(n34330), .A2(n16721), .ZN(n16720) );
  NAND2_X1 U18345 ( .A1(n21040), .A2(n20895), .ZN(n10108) );
  NAND2_X1 U18348 ( .A1(n33644), .A2(n59121), .ZN(n33368) );
  NAND2_X1 U18352 ( .A1(n34086), .A2(n23119), .ZN(n34087) );
  NAND2_X1 U18356 ( .A1(n33483), .A2(n33482), .ZN(n2308) );
  NAND2_X1 U18357 ( .A1(n14811), .A2(n16579), .ZN(n16578) );
  NAND2_X1 U18358 ( .A1(n31237), .A2(n35045), .ZN(n15821) );
  INV_X1 U18359 ( .I(n18681), .ZN(n10932) );
  NAND2_X1 U18360 ( .A1(n33498), .A2(n33728), .ZN(n7150) );
  AOI22_X1 U18362 ( .A1(n4700), .A2(n33517), .B1(n20439), .B2(n11083), .ZN(
        n3223) );
  INV_X1 U18363 ( .I(n12081), .ZN(n3222) );
  NOR2_X1 U18367 ( .A1(n12403), .A2(n12406), .ZN(n14231) );
  INV_X1 U18368 ( .I(n21611), .ZN(n14083) );
  AND2_X1 U18369 ( .A1(n34152), .A2(n19986), .Z(n16254) );
  NOR2_X1 U18370 ( .A1(n31540), .A2(n3582), .ZN(n10639) );
  OAI21_X1 U18373 ( .A1(n35776), .A2(n5874), .B(n64984), .ZN(n35780) );
  INV_X1 U18374 ( .I(n15466), .ZN(n35041) );
  NAND2_X1 U18376 ( .A1(n9910), .A2(n32893), .ZN(n31514) );
  OAI21_X1 U18378 ( .A1(n34065), .A2(n34066), .B(n34076), .ZN(n8344) );
  NAND2_X1 U18381 ( .A1(n10322), .A2(n21432), .ZN(n2395) );
  NAND2_X1 U18382 ( .A1(n34514), .A2(n34515), .ZN(n12914) );
  NOR2_X1 U18383 ( .A1(n2401), .A2(n1539), .ZN(n2399) );
  INV_X1 U18384 ( .I(n33589), .ZN(n11089) );
  OAI21_X1 U18385 ( .A1(n9814), .A2(n9813), .B(n34550), .ZN(n14190) );
  NOR2_X1 U18386 ( .A1(n34543), .A2(n34542), .ZN(n3722) );
  NOR2_X1 U18389 ( .A1(n33379), .A2(n33219), .ZN(n16083) );
  OAI21_X1 U18390 ( .A1(n15286), .A2(n20887), .B(n15285), .ZN(n15284) );
  NAND3_X1 U18392 ( .A1(n10658), .A2(n63888), .A3(n11061), .ZN(n4639) );
  NAND2_X1 U18393 ( .A1(n34016), .A2(n22495), .ZN(n18647) );
  INV_X1 U18394 ( .I(n34770), .ZN(n8115) );
  NAND2_X1 U18396 ( .A1(n5518), .A2(n35042), .ZN(n9134) );
  NAND2_X1 U18398 ( .A1(n33644), .A2(n33643), .ZN(n7465) );
  NAND2_X1 U18399 ( .A1(n9132), .A2(n33446), .ZN(n9128) );
  NOR2_X1 U18404 ( .A1(n33700), .A2(n33701), .ZN(n9797) );
  NAND3_X1 U18410 ( .A1(n34778), .A2(n10016), .A3(n18506), .ZN(n18505) );
  NAND2_X1 U18412 ( .A1(n21813), .A2(n14535), .ZN(n21812) );
  NOR2_X1 U18414 ( .A1(n16991), .A2(n11874), .ZN(n16990) );
  AOI21_X1 U18415 ( .A1(n7207), .A2(n7206), .B(n63305), .ZN(n34630) );
  NOR2_X1 U18416 ( .A1(n3442), .A2(n3441), .ZN(n18945) );
  NAND2_X1 U18417 ( .A1(n4170), .A2(n35213), .ZN(n4164) );
  NAND2_X1 U18418 ( .A1(n32947), .A2(n32946), .ZN(n16133) );
  NAND2_X1 U18421 ( .A1(n34214), .A2(n34215), .ZN(n18896) );
  NOR2_X1 U18423 ( .A1(n33623), .A2(n14329), .ZN(n10103) );
  NAND2_X1 U18426 ( .A1(n34568), .A2(n33757), .ZN(n21807) );
  NAND2_X1 U18428 ( .A1(n57268), .A2(n14702), .ZN(n34663) );
  OAI21_X1 U18429 ( .A1(n32453), .A2(n32452), .B(n33010), .ZN(n32456) );
  INV_X1 U18433 ( .I(n34775), .ZN(n25909) );
  NAND2_X1 U18434 ( .A1(n33538), .A2(n33644), .ZN(n7042) );
  NAND2_X1 U18436 ( .A1(n33530), .A2(n63103), .ZN(n7043) );
  AND3_X1 U18438 ( .A1(n34572), .A2(n32964), .A3(n32300), .Z(n7593) );
  NAND3_X1 U18440 ( .A1(n33980), .A2(n2635), .A3(n33981), .ZN(n33982) );
  NAND2_X1 U18442 ( .A1(n33977), .A2(n33978), .ZN(n19450) );
  AOI22_X1 U18443 ( .A1(n10608), .A2(n35283), .B1(n61496), .B2(n10566), .ZN(
        n35284) );
  AOI21_X1 U18444 ( .A1(n15656), .A2(n1535), .B(n1534), .ZN(n13254) );
  INV_X1 U18445 ( .I(n25216), .ZN(n33779) );
  NAND2_X1 U18449 ( .A1(n34743), .A2(n21464), .ZN(n19443) );
  OAI22_X1 U18451 ( .A1(n33683), .A2(n17759), .B1(n6033), .B2(n22601), .ZN(
        n33682) );
  NOR2_X1 U18456 ( .A1(n33627), .A2(n33623), .ZN(n33625) );
  NAND2_X1 U18459 ( .A1(n10337), .A2(n34385), .ZN(n8631) );
  NOR2_X1 U18461 ( .A1(n33437), .A2(n20835), .ZN(n5158) );
  NAND2_X1 U18463 ( .A1(n9028), .A2(n33801), .ZN(n9843) );
  CLKBUF_X2 U18464 ( .I(n33690), .Z(n10267) );
  NAND2_X1 U18466 ( .A1(n24488), .A2(n26242), .ZN(n18368) );
  NAND2_X1 U18468 ( .A1(n35737), .A2(n16215), .ZN(n13652) );
  OAI22_X1 U18473 ( .A1(n35044), .A2(n9130), .B1(n13068), .B2(n5927), .ZN(
        n35049) );
  NAND2_X1 U18474 ( .A1(n33295), .A2(n9029), .ZN(n33296) );
  NAND2_X1 U18475 ( .A1(n32887), .A2(n34161), .ZN(n31473) );
  AND2_X1 U18476 ( .A1(n21259), .A2(n33947), .Z(n21258) );
  INV_X1 U18477 ( .I(n33956), .ZN(n10641) );
  OAI21_X1 U18478 ( .A1(n32973), .A2(n10016), .B(n7116), .ZN(n2508) );
  NOR2_X1 U18479 ( .A1(n34033), .A2(n19621), .ZN(n34046) );
  OR2_X1 U18482 ( .A1(n3560), .A2(n34080), .Z(n3559) );
  OAI22_X1 U18483 ( .A1(n35777), .A2(n35778), .B1(n11659), .B2(n35786), .ZN(
        n35779) );
  OR2_X1 U18484 ( .A1(n24942), .A2(n16347), .Z(n16264) );
  NAND2_X1 U18485 ( .A1(n32921), .A2(n58076), .ZN(n4747) );
  AOI22_X1 U18486 ( .A1(n35813), .A2(n35306), .B1(n35307), .B2(n8405), .ZN(
        n35311) );
  OAI21_X1 U18487 ( .A1(n32875), .A2(n7453), .B(n33432), .ZN(n11433) );
  INV_X1 U18488 ( .I(n14308), .ZN(n32798) );
  NAND2_X1 U18489 ( .A1(n7174), .A2(n7172), .ZN(n7171) );
  AND2_X1 U18491 ( .A1(n33455), .A2(n34518), .Z(n9460) );
  NAND2_X1 U18493 ( .A1(n1537), .A2(n12169), .ZN(n12168) );
  NOR2_X1 U18496 ( .A1(n7727), .A2(n34959), .ZN(n11582) );
  INV_X1 U18501 ( .I(n9169), .ZN(n34152) );
  OAI21_X1 U18502 ( .A1(n23148), .A2(n22176), .B(n19024), .ZN(n13131) );
  NOR2_X1 U18503 ( .A1(n9169), .A2(n65052), .ZN(n33673) );
  NOR2_X1 U18505 ( .A1(n22419), .A2(n13818), .ZN(n34974) );
  AOI21_X1 U18507 ( .A1(n8689), .A2(n34239), .B(n23556), .ZN(n21483) );
  OAI21_X1 U18508 ( .A1(n12170), .A2(n34949), .B(n34948), .ZN(n9889) );
  NAND2_X1 U18509 ( .A1(n61699), .A2(n33542), .ZN(n32677) );
  NAND2_X1 U18510 ( .A1(n32460), .A2(n15989), .ZN(n32464) );
  INV_X1 U18512 ( .I(n6842), .ZN(n35664) );
  INV_X1 U18514 ( .I(n10866), .ZN(n35331) );
  NOR2_X1 U18517 ( .A1(n33307), .A2(n33596), .ZN(n9717) );
  AND2_X1 U18518 ( .A1(n15927), .A2(n33780), .Z(n12776) );
  OR2_X1 U18519 ( .A1(n33493), .A2(n57710), .Z(n26232) );
  NAND2_X1 U18520 ( .A1(n5902), .A2(n35047), .ZN(n34636) );
  NAND3_X1 U18521 ( .A1(n21538), .A2(n32218), .A3(n34752), .ZN(n32219) );
  INV_X1 U18525 ( .I(n34758), .ZN(n32947) );
  NAND2_X1 U18527 ( .A1(n6579), .A2(n60604), .ZN(n9391) );
  OR2_X1 U18528 ( .A1(n19435), .A2(n61197), .Z(n12587) );
  NAND2_X1 U18530 ( .A1(n9131), .A2(n9130), .ZN(n9126) );
  INV_X1 U18531 ( .I(n12406), .ZN(n34568) );
  OR2_X1 U18532 ( .A1(n22909), .A2(n7531), .Z(n9027) );
  AOI21_X1 U18533 ( .A1(n64958), .A2(n33754), .B(n33753), .ZN(n21809) );
  NAND2_X1 U18535 ( .A1(n34531), .A2(n34971), .ZN(n34532) );
  NOR2_X1 U18536 ( .A1(n30469), .A2(n2273), .ZN(n30470) );
  NAND2_X1 U18537 ( .A1(n33681), .A2(n34157), .ZN(n9039) );
  AOI21_X1 U18538 ( .A1(n15547), .A2(n1538), .B(n34029), .ZN(n12081) );
  OAI22_X1 U18539 ( .A1(n34559), .A2(n35020), .B1(n2208), .B2(n18136), .ZN(
        n29871) );
  OR2_X1 U18540 ( .A1(n19053), .A2(n61449), .Z(n23777) );
  NAND2_X1 U18542 ( .A1(n29558), .A2(n64708), .ZN(n11825) );
  INV_X1 U18544 ( .I(n35708), .ZN(n3903) );
  OR2_X1 U18545 ( .A1(n34997), .A2(n34790), .Z(n15574) );
  NOR2_X1 U18547 ( .A1(n34517), .A2(n3467), .ZN(n8402) );
  AND2_X1 U18550 ( .A1(n8009), .A2(n10769), .Z(n20466) );
  NOR2_X1 U18551 ( .A1(n34523), .A2(n24543), .ZN(n8400) );
  NAND2_X1 U18553 ( .A1(n11423), .A2(n63344), .ZN(n33483) );
  INV_X1 U18554 ( .I(n34017), .ZN(n15141) );
  NAND2_X1 U18556 ( .A1(n12405), .A2(n12404), .ZN(n12403) );
  NAND2_X1 U18557 ( .A1(n34989), .A2(n903), .ZN(n13576) );
  NAND2_X1 U18559 ( .A1(n57268), .A2(n5411), .ZN(n34182) );
  NOR2_X1 U18561 ( .A1(n15547), .A2(n34557), .ZN(n12237) );
  NOR2_X1 U18562 ( .A1(n33476), .A2(n34956), .ZN(n2305) );
  NOR2_X1 U18564 ( .A1(n33484), .A2(n58472), .ZN(n5612) );
  AND2_X1 U18565 ( .A1(n2476), .A2(n12350), .Z(n2825) );
  OAI22_X1 U18567 ( .A1(n33436), .A2(n57165), .B1(n24153), .B2(n33432), .ZN(
        n11434) );
  NAND2_X1 U18568 ( .A1(n33485), .A2(n34510), .ZN(n5609) );
  INV_X1 U18569 ( .I(n57166), .ZN(n9899) );
  NOR2_X1 U18570 ( .A1(n34504), .A2(n35047), .ZN(n15143) );
  OR2_X1 U18572 ( .A1(n14247), .A2(n18136), .Z(n7414) );
  NAND2_X1 U18574 ( .A1(n64100), .A2(n34156), .ZN(n19925) );
  NAND2_X1 U18576 ( .A1(n23125), .A2(n2207), .ZN(n7415) );
  INV_X1 U18580 ( .I(n35663), .ZN(n35219) );
  NAND2_X1 U18581 ( .A1(n33450), .A2(n34056), .ZN(n7174) );
  NAND2_X1 U18583 ( .A1(n24083), .A2(n3467), .ZN(n7172) );
  AND2_X1 U18585 ( .A1(n63375), .A2(n33573), .Z(n6983) );
  NOR2_X1 U18587 ( .A1(n63671), .A2(n63072), .ZN(n33895) );
  NOR2_X1 U18590 ( .A1(n34646), .A2(n35032), .ZN(n9127) );
  NOR2_X1 U18592 ( .A1(n35647), .A2(n22909), .ZN(n3441) );
  NOR2_X1 U18593 ( .A1(n15330), .A2(n15329), .ZN(n15328) );
  NAND2_X1 U18594 ( .A1(n5477), .A2(n34632), .ZN(n5519) );
  INV_X1 U18595 ( .I(n8800), .ZN(n34269) );
  INV_X1 U18596 ( .I(n2968), .ZN(n34685) );
  OR2_X1 U18601 ( .A1(n34324), .A2(n35303), .Z(n16179) );
  AOI21_X1 U18604 ( .A1(n60456), .A2(n4356), .B(n4355), .ZN(n15285) );
  OR2_X1 U18605 ( .A1(n33489), .A2(n7661), .Z(n7660) );
  NAND2_X1 U18606 ( .A1(n24799), .A2(n61748), .ZN(n13895) );
  OAI22_X1 U18607 ( .A1(n33479), .A2(n5529), .B1(n59432), .B2(n1545), .ZN(
        n2304) );
  NAND2_X1 U18609 ( .A1(n35770), .A2(n35775), .ZN(n33918) );
  NOR2_X1 U18610 ( .A1(n32884), .A2(n33), .ZN(n32886) );
  NOR2_X1 U18612 ( .A1(n34413), .A2(n18835), .ZN(n2286) );
  NOR2_X1 U18616 ( .A1(n7849), .A2(n2635), .ZN(n21969) );
  AOI21_X1 U18617 ( .A1(n33), .A2(n60628), .B(n15028), .ZN(n31468) );
  NAND2_X1 U18618 ( .A1(n10822), .A2(n13043), .ZN(n18773) );
  NOR2_X1 U18620 ( .A1(n35795), .A2(n13043), .ZN(n34383) );
  INV_X1 U18621 ( .I(n21041), .ZN(n19563) );
  INV_X2 U18623 ( .I(n7849), .ZN(n34040) );
  NOR2_X1 U18624 ( .A1(n64838), .A2(n6304), .ZN(n3551) );
  INV_X1 U18625 ( .I(n33408), .ZN(n8142) );
  CLKBUF_X2 U18627 ( .I(n35756), .Z(n10504) );
  NAND2_X1 U18628 ( .A1(n61702), .A2(n35745), .ZN(n5996) );
  NOR2_X1 U18629 ( .A1(n20835), .A2(n1312), .ZN(n5161) );
  NAND2_X1 U18630 ( .A1(n33534), .A2(n25428), .ZN(n33371) );
  AOI22_X1 U18631 ( .A1(n34115), .A2(n34116), .B1(n34114), .B2(n60808), .ZN(
        n9852) );
  NAND2_X1 U18632 ( .A1(n34604), .A2(n19512), .ZN(n20444) );
  INV_X1 U18633 ( .I(n34405), .ZN(n34402) );
  NAND4_X1 U18635 ( .A1(n34021), .A2(n34020), .A3(n8694), .A4(n2208), .ZN(
        n34022) );
  NOR2_X1 U18636 ( .A1(n35645), .A2(n35654), .ZN(n7562) );
  INV_X1 U18638 ( .I(n32678), .ZN(n35197) );
  AOI22_X1 U18639 ( .A1(n32944), .A2(n34305), .B1(n57619), .B2(n32946), .ZN(
        n7818) );
  INV_X1 U18640 ( .I(n34994), .ZN(n34510) );
  NAND3_X1 U18641 ( .A1(n33974), .A2(n33975), .A3(n33984), .ZN(n23506) );
  OAI21_X1 U18642 ( .A1(n64708), .A2(n64499), .B(n18136), .ZN(n34028) );
  NAND2_X1 U18643 ( .A1(n9389), .A2(n34726), .ZN(n9302) );
  NAND2_X1 U18644 ( .A1(n14703), .A2(n5410), .ZN(n14614) );
  INV_X1 U18647 ( .I(n4938), .ZN(n9814) );
  AND2_X1 U18649 ( .A1(n16614), .A2(n33561), .Z(n18281) );
  AND2_X1 U18650 ( .A1(n34019), .A2(n57774), .Z(n14192) );
  INV_X1 U18652 ( .I(n35625), .ZN(n33547) );
  AND2_X1 U18653 ( .A1(n33599), .A2(n24688), .Z(n5356) );
  NOR2_X1 U18657 ( .A1(n10656), .A2(n23313), .ZN(n33337) );
  INV_X1 U18662 ( .I(n31358), .ZN(n34664) );
  AND2_X1 U18664 ( .A1(n33752), .A2(n22185), .Z(n7155) );
  NAND2_X1 U18666 ( .A1(n34164), .A2(n5410), .ZN(n3013) );
  AOI21_X1 U18668 ( .A1(n34798), .A2(n61748), .B(n35003), .ZN(n22026) );
  INV_X1 U18670 ( .I(n34997), .ZN(n15575) );
  OR2_X1 U18673 ( .A1(n33406), .A2(n58998), .Z(n3524) );
  CLKBUF_X2 U18674 ( .I(n32454), .Z(n7311) );
  CLKBUF_X2 U18675 ( .I(n24054), .Z(n21096) );
  INV_X1 U18677 ( .I(n35037), .ZN(n5478) );
  INV_X1 U18679 ( .I(n10091), .ZN(n3790) );
  OR2_X1 U18680 ( .A1(n35764), .A2(n35762), .Z(n16243) );
  INV_X1 U18682 ( .I(n22226), .ZN(n9517) );
  INV_X2 U18688 ( .I(n25389), .ZN(n8405) );
  NOR2_X1 U18689 ( .A1(n7321), .A2(n24286), .ZN(n6980) );
  NOR2_X1 U18691 ( .A1(n12506), .A2(n57986), .ZN(n33574) );
  INV_X1 U18694 ( .I(n61496), .ZN(n15408) );
  INV_X1 U18699 ( .I(n33534), .ZN(n12849) );
  INV_X1 U18701 ( .I(n8997), .ZN(n32459) );
  INV_X1 U18703 ( .I(n32965), .ZN(n34959) );
  INV_X1 U18705 ( .I(n35745), .ZN(n35699) );
  INV_X1 U18707 ( .I(n33614), .ZN(n33001) );
  CLKBUF_X2 U18711 ( .I(n61196), .Z(n23351) );
  NAND2_X1 U18713 ( .A1(n3790), .A2(n7534), .ZN(n34072) );
  OR2_X1 U18715 ( .A1(n22723), .A2(n33338), .Z(n16301) );
  NAND2_X1 U18717 ( .A1(n34613), .A2(n33420), .ZN(n14320) );
  INV_X1 U18722 ( .I(n63617), .ZN(n34565) );
  INV_X1 U18723 ( .I(n34529), .ZN(n3669) );
  CLKBUF_X2 U18725 ( .I(n33464), .Z(n9766) );
  AND3_X1 U18734 ( .A1(n10769), .A2(n23717), .A3(n35775), .Z(n16724) );
  INV_X1 U18735 ( .I(n33277), .ZN(n34447) );
  NAND2_X1 U18739 ( .A1(n14110), .A2(n35002), .ZN(n33464) );
  BUF_X2 U18745 ( .I(n2271), .Z(n2033) );
  INV_X2 U18756 ( .I(n24872), .ZN(n1815) );
  INV_X1 U18757 ( .I(n33971), .ZN(n34585) );
  INV_X1 U18759 ( .I(n32571), .ZN(n4933) );
  INV_X2 U18761 ( .I(n33810), .ZN(n35762) );
  CLKBUF_X2 U18766 ( .I(n33336), .Z(n22723) );
  INV_X1 U18767 ( .I(n35001), .ZN(n14110) );
  INV_X1 U18771 ( .I(n33161), .ZN(n24780) );
  INV_X1 U18773 ( .I(n33154), .ZN(n2616) );
  INV_X2 U18774 ( .I(n21939), .ZN(n1817) );
  INV_X1 U18775 ( .I(n17510), .ZN(n9429) );
  INV_X1 U18776 ( .I(n58841), .ZN(n9529) );
  INV_X1 U18777 ( .I(n15629), .ZN(n15288) );
  INV_X1 U18778 ( .I(n32720), .ZN(n11341) );
  INV_X1 U18780 ( .I(n32422), .ZN(n4669) );
  INV_X1 U18782 ( .I(n33192), .ZN(n13428) );
  INV_X1 U18783 ( .I(n2937), .ZN(n33254) );
  INV_X1 U18786 ( .I(n31744), .ZN(n2412) );
  INV_X1 U18787 ( .I(n33132), .ZN(n2173) );
  INV_X2 U18789 ( .I(n16935), .ZN(n1818) );
  INV_X1 U18790 ( .I(n31697), .ZN(n2780) );
  INV_X1 U18793 ( .I(n13475), .ZN(n18720) );
  INV_X1 U18794 ( .I(n24790), .ZN(n11220) );
  INV_X1 U18795 ( .I(n24145), .ZN(n33231) );
  INV_X1 U18796 ( .I(n9179), .ZN(n9462) );
  CLKBUF_X2 U18797 ( .I(n28983), .Z(n10430) );
  INV_X1 U18798 ( .I(n31456), .ZN(n22145) );
  INV_X1 U18800 ( .I(n11265), .ZN(n1952) );
  INV_X1 U18801 ( .I(n8590), .ZN(n14129) );
  INV_X1 U18802 ( .I(n31013), .ZN(n15662) );
  INV_X1 U18805 ( .I(n32572), .ZN(n12665) );
  INV_X1 U18808 ( .I(n25822), .ZN(n32565) );
  INV_X1 U18809 ( .I(n31675), .ZN(n3798) );
  CLKBUF_X2 U18810 ( .I(n16581), .Z(n7225) );
  INV_X1 U18813 ( .I(n61610), .ZN(n12762) );
  INV_X1 U18814 ( .I(n32035), .ZN(n6482) );
  INV_X1 U18815 ( .I(n31288), .ZN(n31289) );
  INV_X1 U18820 ( .I(n33030), .ZN(n17232) );
  CLKBUF_X2 U18821 ( .I(n16458), .Z(n7578) );
  INV_X1 U18822 ( .I(n1347), .ZN(n13277) );
  INV_X1 U18824 ( .I(n33164), .ZN(n9683) );
  CLKBUF_X2 U18825 ( .I(n32244), .Z(n22257) );
  INV_X1 U18828 ( .I(n6322), .ZN(n12123) );
  INV_X2 U18832 ( .I(n32514), .ZN(n19093) );
  INV_X1 U18833 ( .I(n16439), .ZN(n6040) );
  CLKBUF_X4 U18834 ( .I(n32467), .Z(n23389) );
  INV_X1 U18835 ( .I(n15102), .ZN(n31550) );
  NOR2_X1 U18836 ( .A1(n3301), .A2(n3300), .ZN(n3299) );
  CLKBUF_X2 U18837 ( .I(n21986), .Z(n23260) );
  NOR2_X1 U18842 ( .A1(n14544), .A2(n14545), .ZN(n3311) );
  INV_X1 U18843 ( .I(n31630), .ZN(n12520) );
  CLKBUF_X2 U18846 ( .I(n16037), .Z(n9636) );
  INV_X2 U18849 ( .I(n32653), .ZN(n1823) );
  INV_X2 U18850 ( .I(n9283), .ZN(n32475) );
  INV_X1 U18852 ( .I(n15510), .ZN(n11485) );
  NAND2_X1 U18853 ( .A1(n6445), .A2(n24064), .ZN(n6444) );
  INV_X2 U18854 ( .I(n24517), .ZN(n9108) );
  NOR2_X1 U18858 ( .A1(n7909), .A2(n30956), .ZN(n7908) );
  INV_X1 U18859 ( .I(n31629), .ZN(n31855) );
  INV_X1 U18861 ( .I(n31440), .ZN(n12780) );
  INV_X1 U18863 ( .I(n33904), .ZN(n22566) );
  NAND2_X1 U18864 ( .A1(n25083), .A2(n30792), .ZN(n25082) );
  CLKBUF_X2 U18866 ( .I(n33904), .Z(n20838) );
  INV_X2 U18868 ( .I(n16037), .ZN(n1825) );
  INV_X1 U18869 ( .I(n22583), .ZN(n7361) );
  INV_X2 U18871 ( .I(n5402), .ZN(n1826) );
  INV_X1 U18873 ( .I(n24017), .ZN(n9666) );
  INV_X1 U18875 ( .I(n11360), .ZN(n8564) );
  NAND2_X1 U18876 ( .A1(n4778), .A2(n30534), .ZN(n5296) );
  NAND2_X1 U18877 ( .A1(n15527), .A2(n15530), .ZN(n7615) );
  INV_X2 U18880 ( .I(n21944), .ZN(n32494) );
  CLKBUF_X2 U18881 ( .I(n24839), .Z(n10378) );
  INV_X1 U18886 ( .I(n18765), .ZN(n7909) );
  AOI21_X1 U18889 ( .A1(n13813), .A2(n30236), .B(n30235), .ZN(n13812) );
  INV_X1 U18890 ( .I(n1990), .ZN(n1987) );
  CLKBUF_X2 U18892 ( .I(n33239), .Z(n20673) );
  NAND2_X1 U18893 ( .A1(n884), .A2(n2282), .ZN(n2281) );
  NOR2_X1 U18894 ( .A1(n16831), .A2(n16830), .ZN(n23154) );
  NAND2_X1 U18896 ( .A1(n16683), .A2(n16684), .ZN(n15586) );
  NOR2_X1 U18897 ( .A1(n23136), .A2(n30814), .ZN(n23135) );
  NOR2_X1 U18899 ( .A1(n16146), .A2(n16646), .ZN(n25083) );
  CLKBUF_X2 U18900 ( .I(n31873), .Z(n23791) );
  INV_X1 U18905 ( .I(n32543), .ZN(n1831) );
  INV_X2 U18906 ( .I(n20058), .ZN(n1832) );
  NAND2_X2 U18907 ( .A1(n24560), .A2(n24559), .ZN(n32412) );
  NAND4_X1 U18913 ( .A1(n14273), .A2(n14272), .A3(n14275), .A4(n14271), .ZN(
        n24282) );
  INV_X1 U18914 ( .I(n30399), .ZN(n3298) );
  NOR2_X1 U18915 ( .A1(n30399), .A2(n55150), .ZN(n3300) );
  INV_X1 U18920 ( .I(n24008), .ZN(n9698) );
  NAND2_X1 U18921 ( .A1(n12878), .A2(n28908), .ZN(n7569) );
  CLKBUF_X2 U18922 ( .I(n32318), .Z(n22820) );
  NOR2_X1 U18924 ( .A1(n5689), .A2(n5799), .ZN(n5031) );
  CLKBUF_X2 U18929 ( .I(n32057), .Z(n23042) );
  INV_X1 U18933 ( .I(n14271), .ZN(n14270) );
  NOR2_X1 U18936 ( .A1(n13086), .A2(n13085), .ZN(n13084) );
  INV_X1 U18937 ( .I(n27738), .ZN(n5633) );
  INV_X1 U18938 ( .I(n16759), .ZN(n15685) );
  NOR2_X1 U18942 ( .A1(n28743), .A2(n28744), .ZN(n6475) );
  NOR2_X1 U18944 ( .A1(n21061), .A2(n2730), .ZN(n2726) );
  OAI21_X1 U18945 ( .A1(n30731), .A2(n14396), .B(n28775), .ZN(n14395) );
  AOI21_X1 U18946 ( .A1(n28992), .A2(n28993), .B(n5491), .ZN(n5490) );
  NAND3_X1 U18947 ( .A1(n22762), .A2(n30230), .A3(n6539), .ZN(n6538) );
  NAND2_X1 U18950 ( .A1(n28787), .A2(n1554), .ZN(n9340) );
  NOR2_X1 U18951 ( .A1(n27775), .A2(n27774), .ZN(n27778) );
  INV_X1 U18952 ( .I(n29498), .ZN(n17790) );
  OAI21_X1 U18954 ( .A1(n30774), .A2(n30775), .B(n16832), .ZN(n16831) );
  INV_X1 U18956 ( .I(n14274), .ZN(n14273) );
  NAND3_X1 U18960 ( .A1(n8947), .A2(n8945), .A3(n30680), .ZN(n13813) );
  AND2_X1 U18961 ( .A1(n26845), .A2(n26846), .Z(n25635) );
  NOR2_X1 U18965 ( .A1(n7605), .A2(n7603), .ZN(n15623) );
  INV_X1 U18967 ( .I(n30053), .ZN(n2253) );
  AOI22_X1 U18968 ( .A1(n7878), .A2(n8020), .B1(n29864), .B2(n29863), .ZN(
        n8019) );
  NAND2_X1 U18972 ( .A1(n23137), .A2(n30825), .ZN(n23136) );
  NOR2_X1 U18974 ( .A1(n9892), .A2(n9890), .ZN(n29852) );
  NAND2_X1 U18979 ( .A1(n24563), .A2(n20538), .ZN(n24562) );
  OAI21_X1 U18980 ( .A1(n30682), .A2(n30681), .B(n6536), .ZN(n6535) );
  OAI21_X1 U18981 ( .A1(n29774), .A2(n11464), .B(n1552), .ZN(n29775) );
  NAND2_X1 U18982 ( .A1(n18476), .A2(n7594), .ZN(n7605) );
  AOI21_X1 U18983 ( .A1(n29012), .A2(n5859), .B(n29011), .ZN(n4868) );
  OAI21_X1 U18987 ( .A1(n8335), .A2(n9281), .B(n30074), .ZN(n30080) );
  INV_X1 U18999 ( .I(n5654), .ZN(n5653) );
  NAND3_X1 U19001 ( .A1(n30952), .A2(n27780), .A3(n61825), .ZN(n27779) );
  NAND2_X1 U19003 ( .A1(n29883), .A2(n25978), .ZN(n21704) );
  NAND2_X1 U19004 ( .A1(n7037), .A2(n14217), .ZN(n24559) );
  NAND2_X1 U19006 ( .A1(n3988), .A2(n19597), .ZN(n3987) );
  OAI21_X1 U19009 ( .A1(n29965), .A2(n30769), .B(n29964), .ZN(n29966) );
  NOR2_X1 U19011 ( .A1(n16291), .A2(n29815), .ZN(n25631) );
  OAI22_X1 U19012 ( .A1(n29812), .A2(n29811), .B1(n1555), .B2(n30222), .ZN(
        n25317) );
  NOR2_X1 U19016 ( .A1(n17482), .A2(n17481), .ZN(n11672) );
  AOI21_X1 U19017 ( .A1(n28902), .A2(n11988), .B(n28903), .ZN(n5862) );
  NAND2_X1 U19018 ( .A1(n30773), .A2(n11465), .ZN(n16832) );
  INV_X1 U19026 ( .I(n30075), .ZN(n30073) );
  NOR2_X1 U19028 ( .A1(n2734), .A2(n2733), .ZN(n2730) );
  NAND2_X1 U19029 ( .A1(n21063), .A2(n21062), .ZN(n21061) );
  AOI21_X1 U19030 ( .A1(n8753), .A2(n30326), .B(n29273), .ZN(n8752) );
  NAND2_X1 U19033 ( .A1(n3265), .A2(n3264), .ZN(n3263) );
  NAND2_X1 U19035 ( .A1(n9280), .A2(n30075), .ZN(n2729) );
  NAND2_X1 U19036 ( .A1(n29495), .A2(n29497), .ZN(n17784) );
  INV_X1 U19038 ( .I(n25236), .ZN(n17791) );
  NOR2_X1 U19040 ( .A1(n15908), .A2(n15774), .ZN(n17786) );
  OAI21_X1 U19041 ( .A1(n29722), .A2(n29721), .B(n30885), .ZN(n10777) );
  AOI21_X1 U19042 ( .A1(n30589), .A2(n8584), .B(n24913), .ZN(n30592) );
  NOR2_X1 U19045 ( .A1(n28877), .A2(n62892), .ZN(n4483) );
  OAI21_X1 U19047 ( .A1(n12442), .A2(n30502), .B(n30886), .ZN(n30506) );
  INV_X1 U19049 ( .I(n31169), .ZN(n1986) );
  NOR2_X1 U19051 ( .A1(n30241), .A2(n30240), .ZN(n13814) );
  NAND2_X1 U19055 ( .A1(n10492), .A2(n25882), .ZN(n13085) );
  INV_X1 U19057 ( .I(n8424), .ZN(n30318) );
  OAI21_X1 U19058 ( .A1(n28116), .A2(n29453), .B(n29460), .ZN(n8706) );
  NAND2_X1 U19059 ( .A1(n28208), .A2(n31119), .ZN(n9819) );
  INV_X1 U19060 ( .I(n14216), .ZN(n13109) );
  NAND2_X1 U19062 ( .A1(n29519), .A2(n29520), .ZN(n14163) );
  AOI21_X1 U19064 ( .A1(n30350), .A2(n30349), .B(n15979), .ZN(n20387) );
  INV_X1 U19066 ( .I(n25237), .ZN(n1836) );
  NAND2_X1 U19068 ( .A1(n20079), .A2(n30886), .ZN(n20078) );
  NOR2_X1 U19069 ( .A1(n4101), .A2(n4100), .ZN(n4099) );
  INV_X1 U19071 ( .I(n29255), .ZN(n7944) );
  INV_X1 U19072 ( .I(n15136), .ZN(n29211) );
  NOR2_X1 U19073 ( .A1(n31043), .A2(n3989), .ZN(n3988) );
  NAND2_X1 U19075 ( .A1(n19697), .A2(n31116), .ZN(n11662) );
  AOI21_X1 U19077 ( .A1(n30448), .A2(n30449), .B(n19028), .ZN(n15256) );
  NAND2_X1 U19078 ( .A1(n495), .A2(n7965), .ZN(n7964) );
  INV_X1 U19081 ( .I(n7423), .ZN(n2734) );
  OAI21_X1 U19083 ( .A1(n31184), .A2(n31185), .B(n31183), .ZN(n31572) );
  OAI22_X1 U19084 ( .A1(n30190), .A2(n5631), .B1(n29043), .B2(n2177), .ZN(
        n29047) );
  NAND2_X1 U19085 ( .A1(n31033), .A2(n31032), .ZN(n3991) );
  NAND2_X1 U19086 ( .A1(n21777), .A2(n21528), .ZN(n21776) );
  NAND3_X1 U19087 ( .A1(n6256), .A2(n21176), .A3(n31038), .ZN(n29024) );
  NAND3_X1 U19089 ( .A1(n30721), .A2(n14386), .A3(n14384), .ZN(n14388) );
  OAI21_X1 U19091 ( .A1(n9351), .A2(n25241), .B(n29798), .ZN(n20960) );
  OAI21_X1 U19094 ( .A1(n30779), .A2(n4076), .B(n30782), .ZN(n10123) );
  NAND2_X1 U19095 ( .A1(n26783), .A2(n29205), .ZN(n7466) );
  OR2_X1 U19096 ( .A1(n3098), .A2(n30455), .Z(n3097) );
  OAI21_X1 U19097 ( .A1(n28901), .A2(n62647), .B(n28900), .ZN(n5863) );
  NOR2_X1 U19100 ( .A1(n30414), .A2(n30646), .ZN(n30418) );
  NAND2_X1 U19103 ( .A1(n29846), .A2(n29451), .ZN(n28096) );
  NOR3_X1 U19104 ( .A1(n30305), .A2(n4633), .A3(n28428), .ZN(n21401) );
  NAND3_X1 U19105 ( .A1(n30865), .A2(n30864), .A3(n30863), .ZN(n30866) );
  OAI21_X1 U19106 ( .A1(n25513), .A2(n30001), .B(n12656), .ZN(n12657) );
  NOR2_X1 U19109 ( .A1(n28793), .A2(n28794), .ZN(n18102) );
  NAND3_X1 U19110 ( .A1(n18462), .A2(n20315), .A3(n30524), .ZN(n18461) );
  OAI21_X1 U19112 ( .A1(n30324), .A2(n30000), .B(n29999), .ZN(n3108) );
  INV_X1 U19115 ( .I(n28091), .ZN(n8700) );
  NAND3_X1 U19119 ( .A1(n29890), .A2(n11909), .A3(n30885), .ZN(n29891) );
  NAND4_X1 U19120 ( .A1(n11909), .A2(n12893), .A3(n31245), .A4(n5933), .ZN(
        n20282) );
  NOR2_X1 U19121 ( .A1(n30891), .A2(n5933), .ZN(n12808) );
  INV_X1 U19124 ( .I(n30094), .ZN(n11174) );
  INV_X1 U19125 ( .I(n5866), .ZN(n29008) );
  NAND2_X1 U19128 ( .A1(n30233), .A2(n30244), .ZN(n15138) );
  NAND2_X1 U19130 ( .A1(n6769), .A2(n29935), .ZN(n20762) );
  INV_X1 U19131 ( .I(n28748), .ZN(n27781) );
  NAND3_X1 U19133 ( .A1(n6720), .A2(n28751), .A3(n61187), .ZN(n28752) );
  INV_X1 U19134 ( .I(n14921), .ZN(n12376) );
  NOR2_X1 U19136 ( .A1(n12893), .A2(n30888), .ZN(n20079) );
  NAND3_X1 U19137 ( .A1(n29522), .A2(n16228), .A3(n29523), .ZN(n14164) );
  NAND3_X1 U19138 ( .A1(n29234), .A2(n61187), .A3(n11830), .ZN(n29930) );
  INV_X1 U19139 ( .I(n30887), .ZN(n20080) );
  INV_X1 U19140 ( .I(n31093), .ZN(n28208) );
  NAND2_X1 U19141 ( .A1(n30783), .A2(n10122), .ZN(n10121) );
  INV_X1 U19142 ( .I(n30025), .ZN(n3934) );
  INV_X1 U19144 ( .I(n30519), .ZN(n11464) );
  NOR2_X1 U19147 ( .A1(n19216), .A2(n29571), .ZN(n21313) );
  OR3_X1 U19148 ( .A1(n14921), .A2(n65), .A3(n59841), .Z(n9834) );
  OR2_X1 U19150 ( .A1(n30684), .A2(n30685), .Z(n6539) );
  NAND2_X1 U19152 ( .A1(n13361), .A2(n29080), .ZN(n8268) );
  INV_X1 U19153 ( .I(n31035), .ZN(n30134) );
  OR2_X1 U19154 ( .A1(n30313), .A2(n1278), .Z(n28876) );
  NOR2_X1 U19155 ( .A1(n29026), .A2(n17627), .ZN(n17626) );
  NAND2_X1 U19156 ( .A1(n11387), .A2(n30476), .ZN(n9702) );
  OAI22_X1 U19158 ( .A1(n9786), .A2(n9785), .B1(n30158), .B2(n58999), .ZN(
        n20990) );
  INV_X1 U19159 ( .I(n30489), .ZN(n11388) );
  NAND2_X1 U19160 ( .A1(n12470), .A2(n4477), .ZN(n4476) );
  NAND2_X1 U19161 ( .A1(n29843), .A2(n29844), .ZN(n9891) );
  INV_X1 U19162 ( .I(n8961), .ZN(n8960) );
  OR2_X1 U19164 ( .A1(n29033), .A2(n7683), .Z(n26235) );
  NAND2_X1 U19165 ( .A1(n26781), .A2(n8946), .ZN(n8945) );
  OR2_X1 U19166 ( .A1(n30246), .A2(n19461), .Z(n15802) );
  NAND2_X1 U19167 ( .A1(n11206), .A2(n11204), .ZN(n28922) );
  AND2_X1 U19170 ( .A1(n28973), .A2(n13448), .Z(n28974) );
  AOI21_X1 U19173 ( .A1(n29499), .A2(n24852), .B(n3180), .ZN(n5654) );
  NAND2_X1 U19177 ( .A1(n30259), .A2(n30258), .ZN(n6552) );
  INV_X1 U19179 ( .I(n12858), .ZN(n30590) );
  NAND2_X1 U19180 ( .A1(n14602), .A2(n29256), .ZN(n13119) );
  NOR2_X1 U19181 ( .A1(n30684), .A2(n30679), .ZN(n25182) );
  INV_X1 U19182 ( .I(n30475), .ZN(n11387) );
  NAND2_X1 U19183 ( .A1(n30780), .A2(n21886), .ZN(n4076) );
  NAND2_X1 U19184 ( .A1(n23988), .A2(n9865), .ZN(n2429) );
  INV_X1 U19185 ( .I(n30684), .ZN(n25184) );
  INV_X1 U19186 ( .I(n29487), .ZN(n12247) );
  OAI21_X1 U19188 ( .A1(n29749), .A2(n2965), .B(n30786), .ZN(n29750) );
  AND3_X1 U19189 ( .A1(n13810), .A2(n19218), .A3(n30681), .Z(n15964) );
  NAND2_X1 U19190 ( .A1(n30763), .A2(n57806), .ZN(n30014) );
  NOR2_X1 U19191 ( .A1(n16613), .A2(n30303), .ZN(n16612) );
  NAND3_X1 U19193 ( .A1(n2042), .A2(n30885), .A3(n58621), .ZN(n29396) );
  OAI21_X1 U19194 ( .A1(n29985), .A2(n29984), .B(n29992), .ZN(n2103) );
  INV_X1 U19196 ( .I(n5179), .ZN(n27765) );
  NAND2_X1 U19197 ( .A1(n30631), .A2(n1432), .ZN(n12656) );
  INV_X1 U19199 ( .I(n28681), .ZN(n31203) );
  INV_X1 U19200 ( .I(n29538), .ZN(n28907) );
  NOR2_X1 U19201 ( .A1(n28115), .A2(n14399), .ZN(n28097) );
  INV_X1 U19204 ( .I(n29007), .ZN(n4442) );
  NAND3_X1 U19206 ( .A1(n19535), .A2(n30002), .A3(n13280), .ZN(n19534) );
  OR2_X1 U19207 ( .A1(n31119), .A2(n60327), .Z(n11954) );
  OR3_X1 U19209 ( .A1(n30303), .A2(n11206), .A3(n29268), .Z(n28982) );
  NAND3_X1 U19210 ( .A1(n30707), .A2(n15626), .A3(n21176), .ZN(n30146) );
  AOI21_X1 U19211 ( .A1(n30488), .A2(n29814), .B(n29813), .ZN(n29815) );
  NOR2_X1 U19212 ( .A1(n29453), .A2(n7980), .ZN(n27245) );
  AND3_X1 U19213 ( .A1(n30747), .A2(n9979), .A3(n58644), .Z(n30635) );
  INV_X1 U19214 ( .I(n28207), .ZN(n30578) );
  NAND2_X1 U19216 ( .A1(n28771), .A2(n29036), .ZN(n14386) );
  NAND2_X1 U19219 ( .A1(n23072), .A2(n30135), .ZN(n30137) );
  NOR2_X1 U19220 ( .A1(n29842), .A2(n29841), .ZN(n9892) );
  INV_X1 U19221 ( .I(n31045), .ZN(n9786) );
  OR2_X1 U19226 ( .A1(n30375), .A2(n30374), .Z(n10151) );
  AND3_X1 U19227 ( .A1(n6537), .A2(n30678), .A3(n30677), .Z(n6536) );
  INV_X1 U19230 ( .I(n26781), .ZN(n30233) );
  NAND2_X1 U19233 ( .A1(n8892), .A2(n57790), .ZN(n16363) );
  INV_X1 U19234 ( .I(n30299), .ZN(n19216) );
  INV_X1 U19235 ( .I(n8770), .ZN(n8773) );
  NOR2_X1 U19236 ( .A1(n30076), .A2(n9335), .ZN(n14548) );
  NAND2_X1 U19237 ( .A1(n21359), .A2(n21358), .ZN(n21357) );
  AOI21_X1 U19238 ( .A1(n19451), .A2(n62647), .B(n29530), .ZN(n29531) );
  NAND2_X1 U19240 ( .A1(n64894), .A2(n20859), .ZN(n3813) );
  INV_X1 U19241 ( .I(n29060), .ZN(n3820) );
  NAND2_X1 U19242 ( .A1(n25722), .A2(n61928), .ZN(n2440) );
  INV_X1 U19246 ( .I(n29256), .ZN(n13339) );
  AND3_X1 U19247 ( .A1(n7943), .A2(n27610), .A3(n13336), .Z(n13335) );
  NAND2_X1 U19248 ( .A1(n29487), .A2(n23004), .ZN(n30586) );
  INV_X1 U19250 ( .I(n30701), .ZN(n31036) );
  INV_X1 U19251 ( .I(n9581), .ZN(n1839) );
  NOR2_X1 U19252 ( .A1(n31034), .A2(n31040), .ZN(n3985) );
  AOI21_X1 U19253 ( .A1(n11105), .A2(n22742), .B(n11104), .ZN(n6084) );
  NAND2_X1 U19256 ( .A1(n30438), .A2(n29411), .ZN(n17550) );
  NOR2_X1 U19257 ( .A1(n31042), .A2(n31040), .ZN(n20121) );
  AOI21_X1 U19258 ( .A1(n30392), .A2(n4037), .B(n30391), .ZN(n27631) );
  INV_X1 U19259 ( .I(n30737), .ZN(n13033) );
  NAND2_X1 U19260 ( .A1(n17495), .A2(n1551), .ZN(n7087) );
  AND2_X1 U19261 ( .A1(n21640), .A2(n9618), .Z(n16164) );
  INV_X1 U19264 ( .I(n6509), .ZN(n30104) );
  NAND2_X1 U19265 ( .A1(n28077), .A2(n1553), .ZN(n6793) );
  NOR2_X1 U19266 ( .A1(n2119), .A2(n29824), .ZN(n16949) );
  INV_X1 U19267 ( .I(n30857), .ZN(n30856) );
  INV_X1 U19268 ( .I(n31275), .ZN(n8181) );
  NOR2_X1 U19269 ( .A1(n28078), .A2(n7776), .ZN(n28081) );
  AND2_X1 U19271 ( .A1(n30108), .A2(n22322), .Z(n30109) );
  INV_X1 U19272 ( .I(n3706), .ZN(n29829) );
  AND3_X1 U19275 ( .A1(n31073), .A2(n28584), .A3(n61629), .Z(n26231) );
  AOI21_X1 U19276 ( .A1(n1315), .A2(n12907), .B(n30702), .ZN(n29022) );
  OAI21_X1 U19277 ( .A1(n1315), .A2(n12907), .B(n6349), .ZN(n29021) );
  NOR3_X1 U19284 ( .A1(n8584), .A2(n1316), .A3(n31141), .ZN(n8583) );
  NAND2_X1 U19285 ( .A1(n30480), .A2(n1352), .ZN(n27766) );
  NOR2_X1 U19287 ( .A1(n24164), .A2(n24163), .ZN(n30778) );
  INV_X1 U19288 ( .I(n16920), .ZN(n16800) );
  NOR2_X1 U19289 ( .A1(n30618), .A2(n30348), .ZN(n6270) );
  INV_X1 U19291 ( .I(n30226), .ZN(n10371) );
  NOR2_X1 U19292 ( .A1(n28427), .A2(n30296), .ZN(n30305) );
  NAND2_X1 U19294 ( .A1(n20172), .A2(n31201), .ZN(n13243) );
  INV_X1 U19295 ( .I(n30181), .ZN(n22091) );
  INV_X1 U19297 ( .I(n30302), .ZN(n21359) );
  NAND2_X1 U19299 ( .A1(n30077), .A2(n64589), .ZN(n28785) );
  NOR2_X1 U19300 ( .A1(n1554), .A2(n30085), .ZN(n9328) );
  INV_X1 U19301 ( .I(n31082), .ZN(n31081) );
  INV_X1 U19302 ( .I(n30321), .ZN(n21421) );
  INV_X1 U19305 ( .I(n31271), .ZN(n30876) );
  INV_X1 U19306 ( .I(n31166), .ZN(n12471) );
  NAND2_X1 U19307 ( .A1(n21559), .A2(n62231), .ZN(n20343) );
  NAND2_X1 U19309 ( .A1(n13444), .A2(n1353), .ZN(n24251) );
  OAI21_X1 U19311 ( .A1(n14064), .A2(n24097), .B(n29251), .ZN(n28950) );
  INV_X1 U19312 ( .I(n29561), .ZN(n11262) );
  OR2_X1 U19316 ( .A1(n30214), .A2(n30211), .Z(n16219) );
  INV_X1 U19318 ( .I(n7683), .ZN(n18841) );
  INV_X1 U19319 ( .I(n62892), .ZN(n30668) );
  INV_X1 U19321 ( .I(n21134), .ZN(n29513) );
  AND2_X1 U19322 ( .A1(n30296), .A2(n11205), .Z(n16182) );
  INV_X1 U19325 ( .I(n28781), .ZN(n30232) );
  INV_X1 U19326 ( .I(n29821), .ZN(n29985) );
  INV_X1 U19328 ( .I(n30369), .ZN(n26112) );
  OAI21_X1 U19329 ( .A1(n7943), .A2(n29254), .B(n12894), .ZN(n29257) );
  AOI21_X1 U19330 ( .A1(n29996), .A2(n29995), .B(n24896), .ZN(n2100) );
  AND2_X1 U19331 ( .A1(n9197), .A2(n22903), .Z(n9351) );
  INV_X2 U19334 ( .I(n846), .ZN(n29268) );
  INV_X1 U19336 ( .I(n30320), .ZN(n2101) );
  INV_X1 U19337 ( .I(n23397), .ZN(n7776) );
  AND2_X1 U19338 ( .A1(n22014), .A2(n9047), .Z(n11719) );
  INV_X1 U19339 ( .I(n18867), .ZN(n8811) );
  INV_X1 U19341 ( .I(n29246), .ZN(n29784) );
  AND2_X1 U19343 ( .A1(n29846), .A2(n20809), .Z(n14868) );
  AND2_X1 U19345 ( .A1(n18075), .A2(n8891), .Z(n8892) );
  INV_X4 U19351 ( .I(n31098), .ZN(n1856) );
  CLKBUF_X2 U19352 ( .I(n30395), .Z(n22742) );
  CLKBUF_X2 U19353 ( .I(n29988), .Z(n10345) );
  AND2_X1 U19354 ( .A1(n23055), .A2(n22416), .Z(n9000) );
  INV_X1 U19358 ( .I(n29245), .ZN(n9476) );
  INV_X4 U19359 ( .I(n30695), .ZN(n1858) );
  CLKBUF_X2 U19360 ( .I(n30145), .Z(n21019) );
  NAND2_X1 U19363 ( .A1(n23269), .A2(n6316), .ZN(n31165) );
  CLKBUF_X4 U19364 ( .I(n15808), .Z(n23053) );
  BUF_X4 U19370 ( .I(n30486), .Z(n24402) );
  AND2_X1 U19371 ( .A1(n30084), .A2(n131), .Z(n29802) );
  BUF_X4 U19375 ( .I(n30761), .Z(n7426) );
  BUF_X4 U19379 ( .I(n27905), .Z(n29905) );
  BUF_X4 U19383 ( .I(n23705), .Z(n16808) );
  CLKBUF_X2 U19384 ( .I(n30347), .Z(n10240) );
  BUF_X4 U19390 ( .I(n29391), .Z(n31247) );
  NOR2_X1 U19392 ( .A1(n7917), .A2(n7914), .ZN(n7913) );
  NAND2_X1 U19394 ( .A1(n26542), .A2(n26541), .ZN(n23083) );
  NAND2_X1 U19396 ( .A1(n23085), .A2(n26543), .ZN(n23084) );
  NOR2_X1 U19401 ( .A1(n26885), .A2(n26884), .ZN(n26891) );
  NAND3_X1 U19403 ( .A1(n25574), .A2(n25575), .A3(n26725), .ZN(n6555) );
  INV_X1 U19407 ( .I(n9472), .ZN(n9471) );
  AOI21_X1 U19412 ( .A1(n26465), .A2(n26464), .B(n26463), .ZN(n26475) );
  NOR2_X1 U19413 ( .A1(n26496), .A2(n4840), .ZN(n4568) );
  OAI22_X1 U19414 ( .A1(n28377), .A2(n16184), .B1(n23251), .B2(n28378), .ZN(
        n28393) );
  INV_X1 U19416 ( .I(n11638), .ZN(n8169) );
  NOR2_X1 U19417 ( .A1(n7125), .A2(n27950), .ZN(n11095) );
  INV_X1 U19423 ( .I(n27535), .ZN(n15422) );
  OAI21_X1 U19424 ( .A1(n16792), .A2(n26477), .B(n9946), .ZN(n16791) );
  NOR2_X1 U19426 ( .A1(n10305), .A2(n29669), .ZN(n10643) );
  NOR2_X1 U19431 ( .A1(n13006), .A2(n13004), .ZN(n13003) );
  NOR2_X1 U19434 ( .A1(n27418), .A2(n11658), .ZN(n11657) );
  NOR2_X1 U19436 ( .A1(n26538), .A2(n26537), .ZN(n26542) );
  NAND2_X1 U19438 ( .A1(n29359), .A2(n29334), .ZN(n26699) );
  OAI21_X1 U19441 ( .A1(n28145), .A2(n6374), .B(n6372), .ZN(n6371) );
  INV_X1 U19445 ( .I(n14135), .ZN(n26611) );
  INV_X1 U19450 ( .I(n7585), .ZN(n7584) );
  NOR2_X1 U19452 ( .A1(n13762), .A2(n27290), .ZN(n9582) );
  OAI21_X1 U19453 ( .A1(n19548), .A2(n19547), .B(n555), .ZN(n19546) );
  NAND2_X1 U19457 ( .A1(n13516), .A2(n13514), .ZN(n15769) );
  NOR3_X1 U19462 ( .A1(n3197), .A2(n25633), .A3(n26798), .ZN(n3196) );
  NOR2_X1 U19467 ( .A1(n26300), .A2(n16283), .ZN(n20649) );
  NAND2_X1 U19470 ( .A1(n20051), .A2(n20050), .ZN(n20049) );
  NOR2_X1 U19471 ( .A1(n18471), .A2(n18470), .ZN(n21888) );
  NAND2_X1 U19475 ( .A1(n4393), .A2(n4392), .ZN(n26463) );
  AOI21_X1 U19478 ( .A1(n13805), .A2(n13804), .B(n29129), .ZN(n13803) );
  NOR2_X1 U19480 ( .A1(n26006), .A2(n26003), .ZN(n15208) );
  NOR2_X1 U19482 ( .A1(n21629), .A2(n21628), .ZN(n21627) );
  NOR2_X1 U19483 ( .A1(n26806), .A2(n3202), .ZN(n3201) );
  OAI21_X1 U19484 ( .A1(n27663), .A2(n27662), .B(n28499), .ZN(n27673) );
  NOR2_X1 U19486 ( .A1(n14534), .A2(n22992), .ZN(n14531) );
  OAI22_X1 U19488 ( .A1(n29604), .A2(n14938), .B1(n29620), .B2(n14937), .ZN(
        n14936) );
  NOR2_X1 U19491 ( .A1(n19369), .A2(n28486), .ZN(n28487) );
  OAI22_X1 U19492 ( .A1(n8372), .A2(n8371), .B1(n17931), .B2(n28001), .ZN(
        n2113) );
  NAND2_X1 U19494 ( .A1(n28605), .A2(n28451), .ZN(n20051) );
  NAND2_X1 U19496 ( .A1(n16570), .A2(n16794), .ZN(n16792) );
  AOI21_X1 U19498 ( .A1(n9364), .A2(n9363), .B(n23840), .ZN(n14677) );
  AOI21_X1 U19499 ( .A1(n28024), .A2(n28023), .B(n21946), .ZN(n28028) );
  NAND2_X1 U19500 ( .A1(n26378), .A2(n3434), .ZN(n2006) );
  NAND2_X1 U19501 ( .A1(n13188), .A2(n12071), .ZN(n13187) );
  NAND2_X1 U19502 ( .A1(n15770), .A2(n26907), .ZN(n20052) );
  NAND2_X1 U19503 ( .A1(n15985), .A2(n21300), .ZN(n6823) );
  NAND2_X1 U19504 ( .A1(n13378), .A2(n13379), .ZN(n13377) );
  AOI21_X1 U19507 ( .A1(n27943), .A2(n11605), .B(n3793), .ZN(n13761) );
  NAND2_X1 U19509 ( .A1(n26462), .A2(n8518), .ZN(n4392) );
  INV_X1 U19510 ( .I(n44345), .ZN(n23253) );
  NAND2_X1 U19512 ( .A1(n26461), .A2(n26460), .ZN(n4393) );
  NOR2_X1 U19513 ( .A1(n14149), .A2(n14150), .ZN(n5414) );
  NAND2_X1 U19515 ( .A1(n26423), .A2(n8973), .ZN(n8824) );
  NOR2_X1 U19516 ( .A1(n8823), .A2(n22505), .ZN(n8822) );
  NOR2_X1 U19517 ( .A1(n29681), .A2(n29682), .ZN(n29688) );
  OAI22_X1 U19518 ( .A1(n28798), .A2(n6778), .B1(n6777), .B2(n17522), .ZN(
        n6776) );
  NOR2_X1 U19519 ( .A1(n14028), .A2(n27592), .ZN(n12281) );
  AOI21_X1 U19520 ( .A1(n29369), .A2(n6775), .B(n28812), .ZN(n6774) );
  AOI21_X1 U19522 ( .A1(n27963), .A2(n28278), .B(n8778), .ZN(n8779) );
  NAND2_X1 U19523 ( .A1(n4447), .A2(n27657), .ZN(n27663) );
  AND2_X1 U19524 ( .A1(n27864), .A2(n5268), .Z(n27865) );
  NAND2_X1 U19525 ( .A1(n60542), .A2(n23916), .ZN(n27662) );
  AOI21_X1 U19526 ( .A1(n27134), .A2(n27133), .B(n27132), .ZN(n27146) );
  OAI21_X1 U19527 ( .A1(n27956), .A2(n27957), .B(n63850), .ZN(n11093) );
  AOI21_X1 U19528 ( .A1(n27312), .A2(n27311), .B(n12741), .ZN(n9784) );
  INV_X1 U19531 ( .I(n28361), .ZN(n26538) );
  NAND3_X1 U19532 ( .A1(n57270), .A2(n29669), .A3(n29649), .ZN(n29656) );
  AOI22_X1 U19534 ( .A1(n28304), .A2(n16088), .B1(n28308), .B2(n28309), .ZN(
        n24898) );
  NOR3_X1 U19535 ( .A1(n26365), .A2(n26502), .A3(n26364), .ZN(n26369) );
  NOR2_X1 U19537 ( .A1(n27598), .A2(n27597), .ZN(n12276) );
  OAI21_X1 U19538 ( .A1(n26968), .A2(n7437), .B(n19857), .ZN(n26972) );
  NOR2_X1 U19540 ( .A1(n7363), .A2(n18035), .ZN(n18034) );
  OAI21_X1 U19541 ( .A1(n2920), .A2(n2919), .B(n63533), .ZN(n15516) );
  AOI21_X1 U19542 ( .A1(n12280), .A2(n12279), .B(n27609), .ZN(n12278) );
  OAI21_X1 U19543 ( .A1(n26384), .A2(n26385), .B(n27295), .ZN(n16656) );
  AND3_X1 U19544 ( .A1(n27342), .A2(n57270), .A3(n27341), .Z(n27343) );
  OAI21_X1 U19545 ( .A1(n27571), .A2(n27570), .B(n27569), .ZN(n27590) );
  OAI21_X1 U19546 ( .A1(n27715), .A2(n27714), .B(n27713), .ZN(n27721) );
  INV_X1 U19548 ( .I(n26867), .ZN(n11066) );
  OAI21_X1 U19551 ( .A1(n28618), .A2(n13005), .B(n28434), .ZN(n13004) );
  INV_X1 U19554 ( .I(n28185), .ZN(n13414) );
  NOR2_X1 U19555 ( .A1(n27432), .A2(n27618), .ZN(n14177) );
  AOI22_X1 U19556 ( .A1(n29602), .A2(n1567), .B1(n12659), .B2(n29612), .ZN(
        n14941) );
  AND3_X1 U19557 ( .A1(n555), .A2(n19581), .A3(n59935), .Z(n15958) );
  NOR2_X1 U19558 ( .A1(n29183), .A2(n29184), .ZN(n24968) );
  AOI21_X1 U19559 ( .A1(n28286), .A2(n28285), .B(n28284), .ZN(n18501) );
  NAND3_X1 U19560 ( .A1(n19625), .A2(n28845), .A3(n19626), .ZN(n6376) );
  OAI21_X1 U19561 ( .A1(n7920), .A2(n7919), .B(n5153), .ZN(n7918) );
  AOI21_X1 U19562 ( .A1(n28146), .A2(n21203), .B(n6373), .ZN(n6372) );
  AOI21_X1 U19563 ( .A1(n10483), .A2(n10482), .B(n28805), .ZN(n17462) );
  NAND2_X1 U19565 ( .A1(n6603), .A2(n6602), .ZN(n29646) );
  INV_X1 U19566 ( .I(n17634), .ZN(n28809) );
  NAND2_X1 U19567 ( .A1(n7258), .A2(n830), .ZN(n26351) );
  NOR2_X1 U19568 ( .A1(n27417), .A2(n12181), .ZN(n12180) );
  NAND2_X1 U19569 ( .A1(n24818), .A2(n24817), .ZN(n24816) );
  NOR2_X1 U19571 ( .A1(n27477), .A2(n27547), .ZN(n27489) );
  INV_X1 U19572 ( .I(n29117), .ZN(n11513) );
  NAND2_X1 U19574 ( .A1(n27981), .A2(n7499), .ZN(n26750) );
  OAI21_X1 U19575 ( .A1(n26323), .A2(n26324), .B(n21042), .ZN(n26325) );
  OAI21_X1 U19576 ( .A1(n264), .A2(n28168), .B(n64145), .ZN(n28170) );
  NAND2_X1 U19577 ( .A1(n20215), .A2(n15995), .ZN(n28875) );
  OAI21_X1 U19579 ( .A1(n27162), .A2(n10458), .B(n22481), .ZN(n9088) );
  INV_X1 U19580 ( .I(n28667), .ZN(n28173) );
  INV_X1 U19581 ( .I(n29653), .ZN(n29651) );
  INV_X1 U19582 ( .I(n27376), .ZN(n2142) );
  NAND2_X1 U19584 ( .A1(n20511), .A2(n20510), .ZN(n26940) );
  OAI22_X1 U19587 ( .A1(n27444), .A2(n27443), .B1(n27442), .B2(n6759), .ZN(
        n27445) );
  NAND2_X1 U19588 ( .A1(n28508), .A2(n27853), .ZN(n7808) );
  INV_X1 U19589 ( .I(n19857), .ZN(n11875) );
  INV_X1 U19590 ( .I(n14580), .ZN(n6017) );
  NAND2_X1 U19591 ( .A1(n26675), .A2(n26676), .ZN(n9261) );
  NAND2_X1 U19593 ( .A1(n13097), .A2(n12072), .ZN(n12071) );
  NAND2_X1 U19594 ( .A1(n26614), .A2(n26613), .ZN(n13516) );
  NAND2_X1 U19597 ( .A1(n27606), .A2(n27605), .ZN(n9363) );
  INV_X1 U19598 ( .I(n28672), .ZN(n12637) );
  AOI21_X1 U19599 ( .A1(n28233), .A2(n28232), .B(n18224), .ZN(n14580) );
  AOI21_X1 U19600 ( .A1(n28447), .A2(n27854), .B(n13398), .ZN(n13400) );
  INV_X1 U19601 ( .I(n27413), .ZN(n4907) );
  OAI21_X1 U19604 ( .A1(n28664), .A2(n27314), .B(n29603), .ZN(n27316) );
  OAI21_X1 U19605 ( .A1(n6369), .A2(n28151), .B(n19643), .ZN(n27346) );
  INV_X1 U19606 ( .I(n26253), .ZN(n2091) );
  INV_X1 U19607 ( .I(n44290), .ZN(n46276) );
  INV_X1 U19608 ( .I(n27581), .ZN(n27585) );
  NOR2_X1 U19609 ( .A1(n29164), .A2(n13097), .ZN(n12181) );
  AOI21_X1 U19610 ( .A1(n27416), .A2(n5371), .B(n28260), .ZN(n27417) );
  NAND2_X1 U19611 ( .A1(n16492), .A2(n26024), .ZN(n7807) );
  OAI21_X1 U19612 ( .A1(n27268), .A2(n28216), .B(n27970), .ZN(n27269) );
  INV_X1 U19613 ( .I(n2639), .ZN(n16199) );
  NOR2_X1 U19614 ( .A1(n12740), .A2(n6303), .ZN(n27315) );
  NAND2_X1 U19617 ( .A1(n6616), .A2(n27217), .ZN(n6718) );
  NAND2_X1 U19620 ( .A1(n28013), .A2(n7558), .ZN(n10223) );
  INV_X1 U19621 ( .I(n23767), .ZN(n13773) );
  NAND2_X1 U19622 ( .A1(n26499), .A2(n26657), .ZN(n13380) );
  INV_X1 U19624 ( .I(n46437), .ZN(n10810) );
  NOR2_X1 U19625 ( .A1(n7976), .A2(n18780), .ZN(n27984) );
  INV_X1 U19627 ( .I(n20148), .ZN(n8973) );
  INV_X1 U19628 ( .I(n28506), .ZN(n8823) );
  INV_X1 U19629 ( .I(n27715), .ZN(n26837) );
  INV_X1 U19630 ( .I(n33899), .ZN(n38177) );
  NAND2_X1 U19632 ( .A1(n27931), .A2(n6913), .ZN(n2655) );
  INV_X1 U19634 ( .I(n27370), .ZN(n27955) );
  AND2_X1 U19635 ( .A1(n10309), .A2(n13194), .Z(n13193) );
  NAND2_X1 U19636 ( .A1(n28258), .A2(n5306), .ZN(n14258) );
  AND2_X1 U19637 ( .A1(n29647), .A2(n10756), .Z(n10755) );
  AOI22_X1 U19638 ( .A1(n10919), .A2(n8072), .B1(n19279), .B2(n28873), .ZN(
        n10918) );
  NAND2_X1 U19642 ( .A1(n10625), .A2(n14968), .ZN(n10483) );
  NAND2_X1 U19643 ( .A1(n10747), .A2(n7760), .ZN(n15896) );
  NOR2_X1 U19645 ( .A1(n12660), .A2(n12741), .ZN(n12659) );
  NAND2_X1 U19646 ( .A1(n29135), .A2(n29134), .ZN(n3405) );
  NAND2_X1 U19647 ( .A1(n29136), .A2(n6519), .ZN(n3406) );
  NAND2_X1 U19648 ( .A1(n24233), .A2(n29306), .ZN(n24784) );
  NOR2_X1 U19650 ( .A1(n28050), .A2(n11637), .ZN(n28056) );
  NOR2_X1 U19652 ( .A1(n26661), .A2(n21132), .ZN(n27184) );
  NOR2_X1 U19653 ( .A1(n27180), .A2(n1354), .ZN(n8015) );
  NOR2_X1 U19654 ( .A1(n6369), .A2(n4812), .ZN(n6373) );
  NOR2_X1 U19655 ( .A1(n28149), .A2(n28846), .ZN(n19626) );
  NAND2_X1 U19656 ( .A1(n1354), .A2(n1572), .ZN(n18113) );
  INV_X1 U19657 ( .I(n6293), .ZN(n19548) );
  INV_X1 U19658 ( .I(n27169), .ZN(n9468) );
  OAI21_X1 U19659 ( .A1(n20148), .A2(n1569), .B(n28504), .ZN(n28505) );
  OAI22_X1 U19660 ( .A1(n28515), .A2(n8302), .B1(n26043), .B2(n28514), .ZN(
        n28522) );
  INV_X1 U19661 ( .I(n27036), .ZN(n11137) );
  INV_X1 U19662 ( .I(n26529), .ZN(n11136) );
  AND2_X1 U19664 ( .A1(n28618), .A2(n23487), .Z(n15770) );
  NAND2_X1 U19665 ( .A1(n15953), .A2(n21184), .ZN(n26298) );
  NOR2_X1 U19666 ( .A1(n27492), .A2(n12030), .ZN(n7919) );
  NOR3_X1 U19667 ( .A1(n13097), .A2(n28264), .A3(n17909), .ZN(n13098) );
  NAND3_X1 U19669 ( .A1(n19170), .A2(n10404), .A3(n3626), .ZN(n5091) );
  INV_X1 U19671 ( .I(n45286), .ZN(n3242) );
  INV_X1 U19672 ( .I(n26682), .ZN(n7258) );
  AOI22_X1 U19673 ( .A1(n29607), .A2(n27698), .B1(n26878), .B2(n11975), .ZN(
        n26879) );
  AOI21_X1 U19674 ( .A1(n11772), .A2(n57412), .B(n27163), .ZN(n11770) );
  NOR2_X1 U19675 ( .A1(n15651), .A2(n27121), .ZN(n27118) );
  NOR2_X1 U19676 ( .A1(n27131), .A2(n27130), .ZN(n27134) );
  NOR2_X1 U19677 ( .A1(n6863), .A2(n28034), .ZN(n6862) );
  NAND2_X1 U19678 ( .A1(n26799), .A2(n27869), .ZN(n3198) );
  NAND2_X1 U19679 ( .A1(n64614), .A2(n23037), .ZN(n14780) );
  INV_X1 U19680 ( .I(n26992), .ZN(n6777) );
  NAND3_X1 U19681 ( .A1(n28453), .A2(n28607), .A3(n63330), .ZN(n28454) );
  NOR2_X1 U19682 ( .A1(n27851), .A2(n27846), .ZN(n26416) );
  CLKBUF_X2 U19684 ( .I(n52592), .Z(n23249) );
  NOR2_X1 U19686 ( .A1(n29286), .A2(n60894), .ZN(n23430) );
  AOI21_X1 U19688 ( .A1(n28622), .A2(n28621), .B(n28632), .ZN(n28629) );
  OAI21_X1 U19689 ( .A1(n22312), .A2(n28609), .B(n4869), .ZN(n27651) );
  INV_X1 U19690 ( .I(n52470), .ZN(n8279) );
  INV_X1 U19691 ( .I(n28219), .ZN(n29116) );
  NAND2_X1 U19692 ( .A1(n29670), .A2(n25221), .ZN(n11948) );
  OAI21_X1 U19693 ( .A1(n7477), .A2(n27573), .B(n27577), .ZN(n8014) );
  INV_X1 U19694 ( .I(n28460), .ZN(n28614) );
  NAND2_X1 U19695 ( .A1(n29107), .A2(n3904), .ZN(n5407) );
  INV_X1 U19696 ( .I(n28617), .ZN(n13005) );
  CLKBUF_X2 U19698 ( .I(n845), .Z(n9826) );
  INV_X1 U19699 ( .I(n21203), .ZN(n29638) );
  NOR2_X1 U19701 ( .A1(n5218), .A2(n26966), .ZN(n26967) );
  AND2_X1 U19703 ( .A1(n18231), .A2(n29144), .Z(n9098) );
  NOR2_X1 U19704 ( .A1(n28257), .A2(n28256), .ZN(n4822) );
  INV_X1 U19705 ( .I(n29105), .ZN(n14150) );
  INV_X1 U19706 ( .I(n19709), .ZN(n6374) );
  CLKBUF_X2 U19707 ( .I(n46219), .Z(n23767) );
  CLKBUF_X2 U19708 ( .I(n37584), .Z(n22458) );
  AOI21_X1 U19710 ( .A1(n27360), .A2(n23797), .B(n28161), .ZN(n27361) );
  INV_X1 U19711 ( .I(n27850), .ZN(n26734) );
  INV_X1 U19713 ( .I(n11225), .ZN(n26597) );
  OR2_X1 U19714 ( .A1(n5153), .A2(n1360), .Z(n5908) );
  AND2_X1 U19715 ( .A1(n856), .A2(n7538), .Z(n15684) );
  AOI22_X1 U19716 ( .A1(n28460), .A2(n22312), .B1(n28617), .B2(n12263), .ZN(
        n6257) );
  INV_X1 U19717 ( .I(n32583), .ZN(n32112) );
  INV_X1 U19718 ( .I(n4869), .ZN(n27863) );
  INV_X1 U19719 ( .I(n1971), .ZN(n29703) );
  OAI22_X1 U19721 ( .A1(n28380), .A2(n28379), .B1(n28381), .B2(n7886), .ZN(
        n28382) );
  INV_X1 U19722 ( .I(n29134), .ZN(n26381) );
  INV_X1 U19723 ( .I(n27927), .ZN(n12705) );
  INV_X1 U19724 ( .I(n27136), .ZN(n27141) );
  NOR2_X1 U19727 ( .A1(n16845), .A2(n22351), .ZN(n29176) );
  NAND2_X1 U19728 ( .A1(n1569), .A2(n23753), .ZN(n27710) );
  AND2_X1 U19729 ( .A1(n25090), .A2(n27485), .Z(n15779) );
  NOR3_X1 U19732 ( .A1(n23170), .A2(n24060), .A3(n5430), .ZN(n27015) );
  INV_X1 U19733 ( .I(n29107), .ZN(n2112) );
  OAI21_X1 U19734 ( .A1(n28000), .A2(n23166), .B(n19170), .ZN(n8371) );
  INV_X1 U19736 ( .I(n41498), .ZN(n17703) );
  NOR2_X1 U19737 ( .A1(n9908), .A2(n18497), .ZN(n17813) );
  NAND2_X1 U19739 ( .A1(n27262), .A2(n26376), .ZN(n4687) );
  AND2_X1 U19740 ( .A1(n18515), .A2(n23824), .Z(n23930) );
  NAND2_X1 U19742 ( .A1(n14968), .A2(n17460), .ZN(n17457) );
  OR2_X1 U19744 ( .A1(n29668), .A2(n1363), .Z(n15995) );
  NOR2_X1 U19745 ( .A1(n10324), .A2(n27491), .ZN(n25311) );
  NAND2_X1 U19746 ( .A1(n27213), .A2(n59552), .ZN(n24945) );
  OR2_X1 U19748 ( .A1(n26327), .A2(n26536), .Z(n15953) );
  NAND2_X1 U19749 ( .A1(n28665), .A2(n61307), .ZN(n12660) );
  INV_X2 U19750 ( .I(n29173), .ZN(n1878) );
  INV_X1 U19751 ( .I(n11374), .ZN(n29378) );
  NOR2_X1 U19752 ( .A1(n27583), .A2(n10049), .ZN(n12978) );
  NAND2_X1 U19753 ( .A1(n26605), .A2(n26606), .ZN(n12422) );
  NAND2_X1 U19755 ( .A1(n29665), .A2(n29662), .ZN(n10756) );
  AND2_X1 U19756 ( .A1(n22234), .A2(n10321), .Z(n26311) );
  NAND2_X1 U19757 ( .A1(n29643), .A2(n20907), .ZN(n6602) );
  AND2_X1 U19759 ( .A1(n26301), .A2(n26612), .Z(n16283) );
  INV_X1 U19760 ( .I(n24001), .ZN(n12346) );
  AOI21_X1 U19761 ( .A1(n27099), .A2(n6215), .B(n27098), .ZN(n27100) );
  NAND2_X1 U19762 ( .A1(n8420), .A2(n19170), .ZN(n28220) );
  NAND2_X1 U19765 ( .A1(n28842), .A2(n19581), .ZN(n19709) );
  NOR2_X1 U19769 ( .A1(n26958), .A2(n59552), .ZN(n26960) );
  NAND2_X1 U19770 ( .A1(n9661), .A2(n22203), .ZN(n6856) );
  NAND2_X1 U19771 ( .A1(n13194), .A2(n28259), .ZN(n13192) );
  CLKBUF_X2 U19772 ( .I(n38981), .Z(n23020) );
  CLKBUF_X2 U19773 ( .I(n27574), .Z(n23225) );
  INV_X1 U19775 ( .I(n30932), .ZN(n1881) );
  INV_X1 U19776 ( .I(n19593), .ZN(n6381) );
  NOR3_X1 U19777 ( .A1(n28381), .A2(n23007), .A3(n23917), .ZN(n26624) );
  INV_X1 U19779 ( .I(n19581), .ZN(n6515) );
  OR2_X1 U19782 ( .A1(n13399), .A2(n28606), .Z(n13398) );
  NOR2_X1 U19784 ( .A1(n28381), .A2(n23007), .ZN(n2705) );
  INV_X1 U19786 ( .I(n49787), .ZN(n4064) );
  NOR2_X1 U19787 ( .A1(n11873), .A2(n29609), .ZN(n13483) );
  AND2_X1 U19788 ( .A1(n1363), .A2(n29661), .Z(n15893) );
  CLKBUF_X2 U19789 ( .I(n16308), .Z(n22252) );
  AND2_X1 U19790 ( .A1(n28854), .A2(n23797), .Z(n16218) );
  NAND2_X1 U19791 ( .A1(n23797), .A2(n9987), .ZN(n19966) );
  NOR2_X1 U19792 ( .A1(n28673), .A2(n28674), .ZN(n4717) );
  NOR2_X1 U19796 ( .A1(n29295), .A2(n29304), .ZN(n7921) );
  INV_X1 U19797 ( .I(n55139), .ZN(n6815) );
  AND2_X1 U19800 ( .A1(n61035), .A2(n9908), .Z(n16290) );
  INV_X1 U19803 ( .I(n27228), .ZN(n25793) );
  NOR2_X1 U19804 ( .A1(n2066), .A2(n28872), .ZN(n28868) );
  OR2_X1 U19805 ( .A1(n23825), .A2(n28630), .Z(n16241) );
  OR2_X1 U19808 ( .A1(n29372), .A2(n29371), .Z(n16278) );
  INV_X1 U19809 ( .I(n9940), .ZN(n16532) );
  INV_X1 U19813 ( .I(n28328), .ZN(n28054) );
  CLKBUF_X2 U19815 ( .I(n64903), .Z(n21065) );
  CLKBUF_X2 U19817 ( .I(n27189), .Z(n24124) );
  CLKBUF_X2 U19819 ( .I(n29370), .Z(n22158) );
  OR2_X1 U19826 ( .A1(n20240), .A2(n29663), .Z(n28871) );
  INV_X1 U19827 ( .I(n51881), .ZN(n17430) );
  INV_X1 U19828 ( .I(n60797), .ZN(n51610) );
  INV_X1 U19829 ( .I(n16709), .ZN(n12206) );
  CLKBUF_X2 U19830 ( .I(n9548), .Z(n23362) );
  INV_X1 U19831 ( .I(n44613), .ZN(n25934) );
  INV_X1 U19833 ( .I(n15710), .ZN(n1887) );
  CLKBUF_X2 U19834 ( .I(n23800), .Z(n19423) );
  INV_X1 U19836 ( .I(n27859), .ZN(n23814) );
  CLKBUF_X2 U19837 ( .I(n27661), .Z(n22721) );
  INV_X1 U19838 ( .I(n9434), .ZN(n9435) );
  CLKBUF_X2 U19839 ( .I(n26730), .Z(n29120) );
  INV_X2 U19840 ( .I(n59604), .ZN(n29684) );
  CLKBUF_X2 U19842 ( .I(n28632), .Z(n7112) );
  INV_X1 U19843 ( .I(n52511), .ZN(n13114) );
  CLKBUF_X2 U19844 ( .I(n23943), .Z(n9661) );
  INV_X1 U19845 ( .I(n29174), .ZN(n14504) );
  INV_X2 U19847 ( .I(n64155), .ZN(n1890) );
  CLKBUF_X2 U19848 ( .I(n28273), .Z(n23876) );
  CLKBUF_X2 U19850 ( .I(n22352), .Z(n4847) );
  INV_X1 U19854 ( .I(n44467), .ZN(n21779) );
  INV_X2 U19855 ( .I(n29338), .ZN(n1892) );
  INV_X1 U19859 ( .I(n56879), .ZN(n11856) );
  CLKBUF_X4 U19864 ( .I(n27501), .Z(n23496) );
  INV_X1 U19865 ( .I(n56180), .ZN(n11336) );
  BUF_X2 U19867 ( .I(n28303), .Z(n23636) );
  INV_X1 U19868 ( .I(n55580), .ZN(n4525) );
  CLKBUF_X2 U19869 ( .I(n28806), .Z(n23824) );
  INV_X2 U19870 ( .I(n17311), .ZN(n22352) );
  INV_X1 U19871 ( .I(n26275), .ZN(n2941) );
  CLKBUF_X2 U19880 ( .I(n27709), .Z(n23753) );
  INV_X1 U19881 ( .I(n54376), .ZN(n54377) );
  INV_X1 U19882 ( .I(n23158), .ZN(n10747) );
  INV_X1 U19883 ( .I(n56124), .ZN(n56125) );
  INV_X1 U19884 ( .I(n52734), .ZN(n52735) );
  INV_X1 U19885 ( .I(n51569), .ZN(n5890) );
  INV_X1 U19886 ( .I(n54896), .ZN(n2202) );
  CLKBUF_X2 U19887 ( .I(n58420), .Z(n22604) );
  INV_X1 U19888 ( .I(n53154), .ZN(n53155) );
  INV_X1 U19889 ( .I(n53713), .ZN(n53714) );
  INV_X1 U19891 ( .I(n53318), .ZN(n53319) );
  INV_X1 U19893 ( .I(n55777), .ZN(n55778) );
  INV_X1 U19894 ( .I(n56683), .ZN(n56684) );
  INV_X1 U19895 ( .I(n53641), .ZN(n53642) );
  CLKBUF_X2 U19896 ( .I(n27336), .Z(n29663) );
  INV_X1 U19898 ( .I(n54143), .ZN(n52511) );
  INV_X2 U19899 ( .I(n25054), .ZN(n29641) );
  INV_X1 U19900 ( .I(n53748), .ZN(n53749) );
  INV_X1 U19902 ( .I(n53530), .ZN(n53531) );
  CLKBUF_X2 U19903 ( .I(Key[98]), .Z(n55126) );
  CLKBUF_X4 U19905 ( .I(Key[68]), .Z(n54386) );
  CLKBUF_X4 U19906 ( .I(Key[125]), .Z(n55655) );
  CLKBUF_X4 U19909 ( .I(Key[189]), .Z(n57131) );
  CLKBUF_X4 U19910 ( .I(Key[57]), .Z(n54168) );
  INV_X2 U19912 ( .I(n56849), .ZN(n1900) );
  CLKBUF_X4 U19914 ( .I(Key[135]), .Z(n22773) );
  CLKBUF_X2 U19917 ( .I(Key[126]), .Z(n23851) );
  CLKBUF_X4 U19918 ( .I(Key[27]), .Z(n53499) );
  CLKBUF_X2 U19919 ( .I(Key[78]), .Z(n54676) );
  CLKBUF_X4 U19920 ( .I(Key[12]), .Z(n53246) );
  INV_X1 U19921 ( .I(Ciphertext[56]), .ZN(n7123) );
  CLKBUF_X2 U19923 ( .I(Key[82]), .Z(n54748) );
  CLKBUF_X2 U19926 ( .I(Key[167]), .Z(n56745) );
  CLKBUF_X4 U19927 ( .I(Key[14]), .Z(n53262) );
  INV_X1 U19930 ( .I(n57131), .ZN(n21266) );
  CLKBUF_X2 U19932 ( .I(Key[64]), .Z(n4921) );
  CLKBUF_X2 U19934 ( .I(Key[155]), .Z(n24098) );
  CLKBUF_X2 U19935 ( .I(Key[13]), .Z(n22691) );
  CLKBUF_X2 U19936 ( .I(Key[112]), .Z(n19171) );
  CLKBUF_X2 U19937 ( .I(Key[187]), .Z(n20818) );
  CLKBUF_X2 U19939 ( .I(Key[60]), .Z(n20814) );
  XOR2_X1 U19947 ( .A1(n16028), .A2(n1033), .Z(n1905) );
  XOR2_X1 U19949 ( .A1(n11339), .A2(n4215), .Z(n1906) );
  XOR2_X1 U19951 ( .A1(n57187), .A2(n52317), .Z(n1907) );
  AOI21_X1 U19953 ( .A1(n42874), .A2(n1908), .B(n42873), .ZN(n42884) );
  XOR2_X1 U19955 ( .A1(n1910), .A2(n1909), .Z(n12015) );
  NOR2_X2 U19960 ( .A1(n21579), .A2(n2294), .ZN(n19314) );
  NAND2_X2 U19964 ( .A1(n1913), .A2(n1912), .ZN(n45281) );
  XOR2_X1 U19974 ( .A1(n5728), .A2(n39312), .Z(n24241) );
  NOR2_X2 U19975 ( .A1(n7641), .A2(n41020), .ZN(n40500) );
  NAND3_X1 U19977 ( .A1(n20752), .A2(n19300), .A3(n63022), .ZN(n16016) );
  NAND2_X2 U19978 ( .A1(n4336), .A2(n1919), .ZN(n19300) );
  INV_X2 U19979 ( .I(n7955), .ZN(n4336) );
  NOR2_X2 U19984 ( .A1(n28090), .A2(n1923), .ZN(n1922) );
  AND2_X1 U19985 ( .A1(n27306), .A2(n23053), .Z(n1923) );
  OAI22_X1 U19989 ( .A1(n14947), .A2(n57954), .B1(n29123), .B2(n3473), .ZN(
        n13654) );
  NOR2_X1 U19990 ( .A1(n1565), .A2(n57954), .ZN(n15110) );
  INV_X4 U19991 ( .I(n3580), .ZN(n1926) );
  NAND2_X2 U19992 ( .A1(n8287), .A2(n22533), .ZN(n50420) );
  NAND2_X2 U19995 ( .A1(n1252), .A2(n23425), .ZN(n41684) );
  NAND2_X1 U19996 ( .A1(n19946), .A2(n15556), .ZN(n41996) );
  XOR2_X1 U19999 ( .A1(n1928), .A2(n37151), .Z(n37199) );
  XOR2_X1 U20000 ( .A1(n12068), .A2(n9693), .Z(n1928) );
  XOR2_X1 U20002 ( .A1(n1929), .A2(n43773), .Z(n11676) );
  XOR2_X1 U20010 ( .A1(n43912), .A2(n1933), .Z(n1938) );
  XOR2_X1 U20016 ( .A1(n25629), .A2(n1672), .Z(n2881) );
  XOR2_X1 U20017 ( .A1(n12084), .A2(n52570), .Z(n1943) );
  XOR2_X1 U20020 ( .A1(n1946), .A2(n4589), .Z(n6717) );
  XOR2_X1 U20021 ( .A1(n12449), .A2(n50643), .Z(n52570) );
  XOR2_X1 U20023 ( .A1(n24368), .A2(n5626), .Z(n1946) );
  XOR2_X1 U20024 ( .A1(n1948), .A2(n866), .Z(n1947) );
  XOR2_X1 U20025 ( .A1(n25754), .A2(n14742), .Z(n1948) );
  XOR2_X1 U20026 ( .A1(n25828), .A2(n827), .Z(n52322) );
  XOR2_X1 U20030 ( .A1(n1953), .A2(n31683), .Z(n31685) );
  XOR2_X1 U20031 ( .A1(n1951), .A2(n22145), .Z(n31683) );
  XOR2_X1 U20032 ( .A1(n13638), .A2(n1952), .Z(n1951) );
  XOR2_X1 U20035 ( .A1(n31681), .A2(n33177), .Z(n1955) );
  NAND2_X1 U20036 ( .A1(n13614), .A2(n1956), .ZN(n45923) );
  NAND2_X1 U20037 ( .A1(n49948), .A2(n1956), .ZN(n15549) );
  NAND2_X2 U20038 ( .A1(n1379), .A2(n1956), .ZN(n50268) );
  NOR2_X1 U20039 ( .A1(n11623), .A2(n1956), .ZN(n5806) );
  INV_X2 U20040 ( .I(n50271), .ZN(n1956) );
  NAND2_X2 U20041 ( .A1(n1958), .A2(n1957), .ZN(n4898) );
  INV_X2 U20045 ( .I(n2894), .ZN(n47748) );
  NAND2_X1 U20048 ( .A1(n30538), .A2(n1962), .ZN(n29415) );
  AOI21_X1 U20049 ( .A1(n1277), .A2(n1253), .B(n23478), .ZN(n1962) );
  INV_X2 U20052 ( .I(n23126), .ZN(n2153) );
  XOR2_X1 U20053 ( .A1(n8983), .A2(n21767), .Z(n39342) );
  INV_X2 U20065 ( .I(n24165), .ZN(n55443) );
  XOR2_X1 U20066 ( .A1(n1973), .A2(n1972), .Z(n24165) );
  XOR2_X1 U20067 ( .A1(n1620), .A2(n1974), .Z(n1972) );
  XOR2_X1 U20069 ( .A1(n52058), .A2(n1975), .Z(n1974) );
  XOR2_X1 U20070 ( .A1(n6512), .A2(n1119), .Z(n1976) );
  NOR2_X1 U20074 ( .A1(n35731), .A2(n2287), .ZN(n35729) );
  OAI21_X1 U20075 ( .A1(n35747), .A2(n35743), .B(n2287), .ZN(n35744) );
  OAI21_X1 U20076 ( .A1(n35749), .A2(n2287), .B(n904), .ZN(n12935) );
  INV_X4 U20077 ( .I(n34415), .ZN(n2287) );
  INV_X2 U20078 ( .I(n1981), .ZN(n11994) );
  NOR2_X2 U20079 ( .A1(n1307), .A2(n57173), .ZN(n1981) );
  NAND2_X2 U20081 ( .A1(n35266), .A2(n35265), .ZN(n4512) );
  NOR2_X2 U20084 ( .A1(n1989), .A2(n1988), .ZN(n33185) );
  XOR2_X1 U20088 ( .A1(n3755), .A2(n14442), .Z(n1995) );
  INV_X1 U20090 ( .I(n12084), .ZN(n1996) );
  INV_X2 U20096 ( .I(n53196), .ZN(n2001) );
  AND2_X2 U20099 ( .A1(n24334), .A2(n16894), .Z(n29959) );
  INV_X2 U20102 ( .I(n2013), .ZN(n6789) );
  OAI21_X1 U20103 ( .A1(n1178), .A2(n2013), .B(n2012), .ZN(n53266) );
  NAND2_X1 U20104 ( .A1(n2013), .A2(n53303), .ZN(n2012) );
  NOR2_X2 U20105 ( .A1(n53294), .A2(n19735), .ZN(n2013) );
  NOR2_X1 U20106 ( .A1(n6789), .A2(n2014), .ZN(n19578) );
  XOR2_X1 U20110 ( .A1(n7205), .A2(n33162), .Z(n2017) );
  INV_X1 U20111 ( .I(n2018), .ZN(n12439) );
  NOR2_X1 U20113 ( .A1(n25067), .A2(n2018), .ZN(n52839) );
  AOI21_X1 U20114 ( .A1(n53605), .A2(n2018), .B(n25067), .ZN(n52752) );
  NAND2_X2 U20116 ( .A1(n23401), .A2(n15713), .ZN(n2018) );
  XOR2_X1 U20126 ( .A1(n2029), .A2(n17473), .Z(n2028) );
  XOR2_X1 U20127 ( .A1(n37824), .A2(n39582), .Z(n2029) );
  XOR2_X1 U20130 ( .A1(n39300), .A2(n17772), .Z(n2032) );
  XOR2_X1 U20131 ( .A1(n2035), .A2(n2034), .Z(n2271) );
  XOR2_X1 U20132 ( .A1(n23760), .A2(n17727), .Z(n2034) );
  XOR2_X1 U20133 ( .A1(n32281), .A2(n17201), .Z(n2035) );
  XOR2_X1 U20134 ( .A1(n2070), .A2(n52525), .Z(n7292) );
  XOR2_X1 U20135 ( .A1(n9230), .A2(n50606), .Z(n52525) );
  NAND3_X2 U20141 ( .A1(n2709), .A2(n2708), .A3(n2707), .ZN(n6564) );
  XOR2_X1 U20142 ( .A1(n43863), .A2(n43862), .Z(n3501) );
  XOR2_X1 U20143 ( .A1(n20230), .A2(n11111), .Z(n43863) );
  INV_X2 U20150 ( .I(n8464), .ZN(n11231) );
  INV_X2 U20153 ( .I(n7627), .ZN(n32393) );
  OAI22_X1 U20165 ( .A1(n16024), .A2(n19294), .B1(n2047), .B2(n6323), .ZN(
        n3921) );
  NAND2_X1 U20166 ( .A1(n47922), .A2(n49057), .ZN(n2046) );
  NAND2_X2 U20168 ( .A1(n54904), .A2(n2329), .ZN(n54892) );
  NOR2_X1 U20173 ( .A1(n33785), .A2(n15045), .ZN(n2056) );
  NOR2_X1 U20177 ( .A1(n22295), .A2(n2059), .ZN(n36180) );
  NOR2_X1 U20179 ( .A1(n36170), .A2(n2059), .ZN(n2057) );
  OAI22_X1 U20180 ( .A1(n36129), .A2(n2059), .B1(n12804), .B2(n21802), .ZN(
        n13345) );
  OAI22_X1 U20187 ( .A1(n6312), .A2(n54815), .B1(n15023), .B2(n14358), .ZN(
        n54097) );
  INV_X1 U20188 ( .I(n58806), .ZN(n2062) );
  INV_X1 U20190 ( .I(n2064), .ZN(n2063) );
  NOR2_X1 U20191 ( .A1(n34251), .A2(n2064), .ZN(n32930) );
  OAI22_X1 U20192 ( .A1(n34252), .A2(n64965), .B1(n34254), .B2(n2064), .ZN(
        n34255) );
  OAI21_X1 U20193 ( .A1(n33745), .A2(n33744), .B(n2064), .ZN(n33749) );
  INV_X2 U20196 ( .I(n10908), .ZN(n23805) );
  NOR2_X1 U20198 ( .A1(n2068), .A2(n22446), .ZN(n42584) );
  NAND2_X1 U20209 ( .A1(n2081), .A2(n18418), .ZN(n4139) );
  XOR2_X1 U20211 ( .A1(n2083), .A2(n2082), .Z(n2769) );
  XOR2_X1 U20212 ( .A1(n44733), .A2(n8862), .Z(n2082) );
  INV_X2 U20214 ( .I(n46178), .ZN(n8862) );
  XOR2_X1 U20219 ( .A1(n2747), .A2(n44028), .Z(n2086) );
  XOR2_X1 U20220 ( .A1(n25348), .A2(n12835), .Z(n2747) );
  XOR2_X1 U20221 ( .A1(n25364), .A2(n3389), .Z(n33132) );
  NOR2_X2 U20223 ( .A1(n2408), .A2(n52704), .ZN(n56545) );
  XOR2_X1 U20224 ( .A1(Ciphertext[63]), .A2(Key[142]), .Z(n21656) );
  NOR2_X2 U20225 ( .A1(n2087), .A2(n9588), .ZN(n42916) );
  OAI21_X1 U20229 ( .A1(n2091), .A2(n28270), .B(n62663), .ZN(n28272) );
  NAND2_X2 U20232 ( .A1(n11414), .A2(n22113), .ZN(n36583) );
  NOR2_X2 U20239 ( .A1(n5708), .A2(n5706), .ZN(n38612) );
  XOR2_X1 U20241 ( .A1(n6889), .A2(n39246), .Z(n2108) );
  XOR2_X1 U20242 ( .A1(n23949), .A2(n23093), .Z(n39246) );
  XOR2_X1 U20249 ( .A1(n12563), .A2(n2109), .Z(n11852) );
  XNOR2_X1 U20250 ( .A1(n6342), .A2(n26245), .ZN(n11446) );
  NAND3_X2 U20251 ( .A1(n5679), .A2(n5680), .A3(n5681), .ZN(n26245) );
  INV_X2 U20253 ( .I(n37118), .ZN(n38757) );
  XOR2_X1 U20254 ( .A1(n37118), .A2(n62273), .Z(n2114) );
  NAND2_X2 U20256 ( .A1(n2303), .A2(n2307), .ZN(n4893) );
  NOR2_X1 U20258 ( .A1(n29275), .A2(n2120), .ZN(n4104) );
  NAND2_X2 U20260 ( .A1(n18423), .A2(n2295), .ZN(n28281) );
  NOR2_X1 U20265 ( .A1(n2122), .A2(n61256), .ZN(n32208) );
  NOR2_X2 U20266 ( .A1(n3308), .A2(n2122), .ZN(n33493) );
  NOR2_X1 U20267 ( .A1(n2617), .A2(n2122), .ZN(n12513) );
  NAND2_X2 U20268 ( .A1(n34784), .A2(n64387), .ZN(n2122) );
  NAND2_X2 U20269 ( .A1(n29200), .A2(n29203), .ZN(n30845) );
  NAND2_X1 U20270 ( .A1(n60171), .A2(n14102), .ZN(n29112) );
  XOR2_X1 U20277 ( .A1(n39248), .A2(n22757), .Z(n2125) );
  XOR2_X1 U20278 ( .A1(n38220), .A2(n23518), .Z(n39248) );
  XOR2_X1 U20280 ( .A1(n11508), .A2(n11545), .Z(n2127) );
  INV_X2 U20281 ( .I(n15873), .ZN(n17801) );
  XOR2_X1 U20286 ( .A1(n32163), .A2(n2133), .Z(n2132) );
  XOR2_X1 U20287 ( .A1(n2130), .A2(n32568), .Z(n32163) );
  INV_X2 U20291 ( .I(n14740), .ZN(n15153) );
  XOR2_X1 U20292 ( .A1(n20719), .A2(n16706), .Z(n2133) );
  NAND2_X2 U20295 ( .A1(n2137), .A2(n2134), .ZN(n29053) );
  AND2_X1 U20303 ( .A1(n44943), .A2(n46024), .Z(n2151) );
  INV_X2 U20304 ( .I(n2152), .ZN(n24757) );
  XOR2_X1 U20305 ( .A1(n2154), .A2(n24757), .Z(n52628) );
  XOR2_X1 U20309 ( .A1(n2153), .A2(n2155), .Z(n2154) );
  XOR2_X1 U20310 ( .A1(n52627), .A2(n52626), .Z(n2155) );
  INV_X2 U20311 ( .I(n19300), .ZN(n3188) );
  NOR2_X2 U20312 ( .A1(n19982), .A2(n17349), .ZN(n38344) );
  INV_X2 U20315 ( .I(n57330), .ZN(n37118) );
  XOR2_X1 U20317 ( .A1(n2928), .A2(n59895), .Z(n38470) );
  XOR2_X1 U20318 ( .A1(n1411), .A2(n57330), .Z(n37553) );
  NAND2_X2 U20319 ( .A1(n2157), .A2(n49700), .ZN(n48354) );
  NOR2_X1 U20322 ( .A1(n2158), .A2(n19573), .ZN(n34456) );
  XOR2_X1 U20323 ( .A1(n2158), .A2(n19573), .Z(n17998) );
  NAND2_X2 U20324 ( .A1(n20124), .A2(n37359), .ZN(n2158) );
  NAND3_X1 U20326 ( .A1(n12174), .A2(n17410), .A3(n2267), .ZN(n12160) );
  OAI21_X1 U20329 ( .A1(n29759), .A2(n30051), .B(n2267), .ZN(n29761) );
  NAND2_X2 U20332 ( .A1(n2161), .A2(n40170), .ZN(n42695) );
  XOR2_X1 U20337 ( .A1(n1189), .A2(n7246), .Z(n25395) );
  XOR2_X1 U20339 ( .A1(n5798), .A2(n2173), .Z(n2172) );
  XOR2_X1 U20341 ( .A1(n2175), .A2(n8236), .Z(n2174) );
  XOR2_X1 U20342 ( .A1(n33885), .A2(n17847), .Z(n2175) );
  NAND2_X1 U20346 ( .A1(n30099), .A2(n2177), .ZN(n7604) );
  NOR2_X2 U20348 ( .A1(n25841), .A2(n24615), .ZN(n2179) );
  NAND2_X1 U20350 ( .A1(n18766), .A2(n2178), .ZN(n8574) );
  AOI21_X1 U20351 ( .A1(n47798), .A2(n2178), .B(n23180), .ZN(n47804) );
  OAI21_X1 U20352 ( .A1(n47706), .A2(n61756), .B(n2178), .ZN(n45306) );
  XOR2_X1 U20356 ( .A1(n51302), .A2(n2184), .Z(n2183) );
  INV_X2 U20361 ( .I(n2192), .ZN(n3625) );
  NAND2_X1 U20362 ( .A1(n41127), .A2(n2193), .ZN(n41128) );
  XOR2_X1 U20366 ( .A1(n2391), .A2(n31750), .Z(n7008) );
  AOI21_X1 U20368 ( .A1(n19652), .A2(n45808), .B(n47368), .ZN(n10673) );
  NOR2_X1 U20370 ( .A1(n17155), .A2(n7200), .ZN(n55182) );
  INV_X2 U20371 ( .I(n5214), .ZN(n5989) );
  INV_X1 U20375 ( .I(n18862), .ZN(n20278) );
  NAND2_X2 U20380 ( .A1(n42006), .A2(n24250), .ZN(n2197) );
  AND2_X1 U20383 ( .A1(n8444), .A2(n30252), .Z(n2370) );
  NAND2_X1 U20384 ( .A1(n8443), .A2(n30255), .ZN(n8444) );
  XOR2_X1 U20386 ( .A1(n2203), .A2(n2202), .Z(Plaintext[86]) );
  XOR2_X1 U20390 ( .A1(n52147), .A2(n12419), .Z(n11307) );
  XOR2_X1 U20391 ( .A1(n18512), .A2(n2212), .Z(n52147) );
  XOR2_X1 U20392 ( .A1(n12299), .A2(n23283), .Z(n2212) );
  XOR2_X1 U20394 ( .A1(n52323), .A2(n14730), .Z(n2215) );
  INV_X2 U20396 ( .I(n17317), .ZN(n47568) );
  OAI22_X2 U20397 ( .A1(n47905), .A2(n47902), .B1(n47576), .B2(n2571), .ZN(
        n17317) );
  INV_X2 U20398 ( .I(n2217), .ZN(n22142) );
  XOR2_X1 U20402 ( .A1(n39480), .A2(n14646), .Z(n2219) );
  XOR2_X1 U20417 ( .A1(n51749), .A2(n23022), .Z(n50992) );
  XOR2_X1 U20424 ( .A1(n879), .A2(n4279), .Z(n11981) );
  NOR2_X1 U20428 ( .A1(n2240), .A2(n53281), .ZN(n53276) );
  INV_X2 U20429 ( .I(n17904), .ZN(n28223) );
  NAND2_X1 U20431 ( .A1(n28224), .A2(n17904), .ZN(n29104) );
  XOR2_X1 U20432 ( .A1(n32098), .A2(n4278), .Z(n4280) );
  INV_X2 U20433 ( .I(n18490), .ZN(n4278) );
  NAND2_X2 U20436 ( .A1(n16380), .A2(n20251), .ZN(n37942) );
  NAND2_X2 U20444 ( .A1(n49542), .A2(n49529), .ZN(n49379) );
  OAI22_X1 U20448 ( .A1(n40805), .A2(n41906), .B1(n40579), .B2(n2247), .ZN(
        n40580) );
  OAI21_X1 U20452 ( .A1(n47883), .A2(n47882), .B(n2250), .ZN(n47889) );
  NAND2_X2 U20454 ( .A1(n2269), .A2(n9047), .ZN(n30050) );
  INV_X1 U20463 ( .I(n63263), .ZN(n52549) );
  XOR2_X1 U20465 ( .A1(n15487), .A2(n63263), .Z(n2257) );
  XOR2_X1 U20468 ( .A1(n2258), .A2(n22795), .Z(n52550) );
  XOR2_X1 U20469 ( .A1(n52443), .A2(n52444), .Z(n2258) );
  INV_X2 U20473 ( .I(n24301), .ZN(n22807) );
  NOR2_X1 U20475 ( .A1(n50212), .A2(n2262), .ZN(n50013) );
  OAI21_X1 U20476 ( .A1(n50216), .A2(n2262), .B(n1383), .ZN(n50016) );
  NAND2_X1 U20477 ( .A1(n8120), .A2(n2262), .ZN(n50214) );
  XOR2_X1 U20479 ( .A1(n2266), .A2(n2263), .Z(n3039) );
  XOR2_X1 U20480 ( .A1(n2264), .A2(n2265), .Z(n2263) );
  INV_X2 U20486 ( .I(n14721), .ZN(n41007) );
  NAND2_X2 U20488 ( .A1(n41007), .A2(n41019), .ZN(n40603) );
  XOR2_X1 U20489 ( .A1(n2842), .A2(n9108), .Z(n11506) );
  INV_X2 U20490 ( .I(n24522), .ZN(n9012) );
  XOR2_X1 U20492 ( .A1(n6306), .A2(n23583), .Z(n21299) );
  NAND3_X2 U20493 ( .A1(n36007), .A2(n36006), .A3(n36005), .ZN(n38145) );
  NOR3_X1 U20500 ( .A1(n2286), .A2(n35729), .A3(n60527), .ZN(n2288) );
  XOR2_X1 U20501 ( .A1(n2289), .A2(n5899), .Z(n3894) );
  XOR2_X1 U20504 ( .A1(n26062), .A2(n33175), .Z(n33877) );
  NAND2_X2 U20508 ( .A1(n2291), .A2(n2688), .ZN(n2686) );
  NOR3_X2 U20509 ( .A1(n2293), .A2(n1025), .A3(n2292), .ZN(n2291) );
  XOR2_X1 U20511 ( .A1(n14), .A2(n804), .Z(n15839) );
  NAND2_X2 U20516 ( .A1(n2297), .A2(n2296), .ZN(n23491) );
  NOR4_X2 U20523 ( .A1(n33480), .A2(n2306), .A3(n2305), .A4(n2304), .ZN(n2303)
         );
  INV_X2 U20524 ( .I(n2309), .ZN(n45551) );
  NOR2_X2 U20529 ( .A1(n2312), .A2(n13969), .ZN(n15692) );
  XOR2_X1 U20532 ( .A1(n24859), .A2(n37820), .Z(n2317) );
  NAND3_X1 U20534 ( .A1(n3650), .A2(n3647), .A3(n50606), .ZN(n2318) );
  AOI21_X1 U20535 ( .A1(n3650), .A2(n3647), .B(n50606), .ZN(n2320) );
  INV_X2 U20541 ( .I(n17018), .ZN(n24522) );
  INV_X2 U20543 ( .I(n2324), .ZN(n2867) );
  XOR2_X1 U20547 ( .A1(n44144), .A2(n43138), .Z(n2327) );
  XOR2_X1 U20548 ( .A1(n10893), .A2(n2540), .Z(n2328) );
  NAND2_X2 U20550 ( .A1(n54813), .A2(n58843), .ZN(n5140) );
  INV_X2 U20551 ( .I(n6873), .ZN(n54813) );
  NOR2_X2 U20553 ( .A1(n1225), .A2(n1701), .ZN(n43131) );
  INV_X2 U20558 ( .I(n2342), .ZN(n16707) );
  XOR2_X1 U20561 ( .A1(n6056), .A2(n6684), .Z(n2345) );
  NAND3_X1 U20563 ( .A1(n61900), .A2(n2350), .A3(n30224), .ZN(n24973) );
  INV_X1 U20568 ( .I(n22698), .ZN(n2356) );
  NAND3_X2 U20576 ( .A1(n25360), .A2(n26174), .A3(n44946), .ZN(n22962) );
  INV_X2 U20577 ( .I(n3118), .ZN(n21984) );
  XOR2_X1 U20585 ( .A1(n1828), .A2(n31371), .Z(n2364) );
  XOR2_X1 U20589 ( .A1(n17618), .A2(n45357), .Z(n2365) );
  INV_X2 U20597 ( .I(n25300), .ZN(n27966) );
  NAND2_X2 U20599 ( .A1(n29054), .A2(n30048), .ZN(n12174) );
  NAND2_X2 U20600 ( .A1(n22014), .A2(n2269), .ZN(n29054) );
  NOR2_X1 U20602 ( .A1(n2372), .A2(n56885), .ZN(n17362) );
  INV_X1 U20605 ( .I(n29876), .ZN(n2374) );
  NAND2_X2 U20612 ( .A1(n2385), .A2(n2384), .ZN(n9806) );
  OR2_X1 U20614 ( .A1(n34226), .A2(n34225), .Z(n2385) );
  NAND2_X2 U20619 ( .A1(n2400), .A2(n2397), .ZN(n19765) );
  INV_X2 U20626 ( .I(n2409), .ZN(n52704) );
  XOR2_X1 U20627 ( .A1(n51317), .A2(n51315), .Z(n2410) );
  XOR2_X1 U20629 ( .A1(n2413), .A2(n2412), .Z(n4592) );
  XOR2_X1 U20630 ( .A1(n6309), .A2(n17701), .Z(n2413) );
  AOI21_X1 U20635 ( .A1(n63589), .A2(n30197), .B(n59798), .ZN(n2416) );
  NAND2_X2 U20637 ( .A1(n5099), .A2(n5604), .ZN(n34221) );
  OR2_X1 U20639 ( .A1(n34780), .A2(n19025), .Z(n2420) );
  NOR2_X1 U20640 ( .A1(n2422), .A2(n56734), .ZN(n56727) );
  NAND2_X1 U20643 ( .A1(n9559), .A2(n2422), .ZN(n8827) );
  NAND3_X2 U20644 ( .A1(n56725), .A2(n20696), .A3(n56697), .ZN(n2422) );
  XOR2_X1 U20650 ( .A1(n46522), .A2(n45127), .Z(n2425) );
  NOR2_X2 U20654 ( .A1(n29271), .A2(n23216), .ZN(n16959) );
  XOR2_X1 U20655 ( .A1(n25037), .A2(n31863), .Z(n33178) );
  INV_X2 U20657 ( .I(n2428), .ZN(n24951) );
  XNOR2_X1 U20658 ( .A1(Ciphertext[33]), .A2(Key[124]), .ZN(n2428) );
  NAND2_X2 U20659 ( .A1(n8218), .A2(n1317), .ZN(n29266) );
  INV_X1 U20660 ( .I(n13817), .ZN(n21814) );
  NAND2_X1 U20662 ( .A1(n45555), .A2(n2432), .ZN(n2431) );
  NOR2_X2 U20663 ( .A1(n45558), .A2(n2434), .ZN(n23514) );
  AND2_X1 U20664 ( .A1(n45978), .A2(n47275), .Z(n2432) );
  NOR2_X1 U20670 ( .A1(n15936), .A2(n2435), .ZN(n9405) );
  NOR2_X2 U20672 ( .A1(n48135), .A2(n24545), .ZN(n46455) );
  NAND2_X2 U20674 ( .A1(n23114), .A2(n4897), .ZN(n47087) );
  AOI21_X1 U20677 ( .A1(n42655), .A2(n14920), .B(n6426), .ZN(n2451) );
  XOR2_X1 U20679 ( .A1(n2452), .A2(n2453), .Z(n8554) );
  XOR2_X1 U20681 ( .A1(n63027), .A2(n23579), .Z(n15766) );
  XOR2_X1 U20682 ( .A1(n63027), .A2(n44805), .Z(n2481) );
  XOR2_X1 U20685 ( .A1(n2457), .A2(n6166), .Z(n4220) );
  XOR2_X1 U20687 ( .A1(n3530), .A2(n2457), .Z(n3529) );
  XOR2_X1 U20689 ( .A1(n2457), .A2(n5184), .Z(n5183) );
  XOR2_X1 U20690 ( .A1(n2458), .A2(n17800), .Z(n11242) );
  NAND2_X1 U20693 ( .A1(n2459), .A2(n42452), .ZN(n40360) );
  NAND2_X1 U20694 ( .A1(n2459), .A2(n22759), .ZN(n42449) );
  NAND2_X2 U20695 ( .A1(n1733), .A2(n19291), .ZN(n2459) );
  INV_X1 U20696 ( .I(n2460), .ZN(n18216) );
  NOR2_X1 U20697 ( .A1(n12885), .A2(n2460), .ZN(n12884) );
  NOR2_X2 U20699 ( .A1(n36742), .A2(n20812), .ZN(n2460) );
  INV_X2 U20700 ( .I(n3639), .ZN(n34035) );
  XOR2_X1 U20701 ( .A1(n880), .A2(n2461), .Z(n3639) );
  XOR2_X1 U20702 ( .A1(n31020), .A2(n33266), .Z(n2461) );
  XOR2_X1 U20703 ( .A1(n2465), .A2(n25530), .Z(n4703) );
  XOR2_X1 U20706 ( .A1(n44892), .A2(n44804), .Z(n2465) );
  NOR2_X2 U20709 ( .A1(n54605), .A2(n54778), .ZN(n54955) );
  INV_X2 U20711 ( .I(n2469), .ZN(n39011) );
  NAND2_X2 U20718 ( .A1(n2329), .A2(n13671), .ZN(n54898) );
  NAND3_X1 U20719 ( .A1(n2476), .A2(n34512), .A3(n34068), .ZN(n8346) );
  NAND2_X2 U20720 ( .A1(n2322), .A2(n1424), .ZN(n2476) );
  NAND2_X1 U20724 ( .A1(n696), .A2(n48983), .ZN(n14069) );
  INV_X2 U20726 ( .I(n24887), .ZN(n47901) );
  XOR2_X1 U20727 ( .A1(n2480), .A2(n2478), .Z(n24887) );
  XOR2_X1 U20728 ( .A1(n1023), .A2(n2479), .Z(n2478) );
  XOR2_X1 U20730 ( .A1(n2482), .A2(n2481), .Z(n2480) );
  XOR2_X1 U20734 ( .A1(n2487), .A2(n2484), .Z(n2485) );
  XOR2_X1 U20736 ( .A1(n52370), .A2(n17143), .Z(n2484) );
  XOR2_X1 U20737 ( .A1(n51583), .A2(n8007), .Z(n17143) );
  INV_X2 U20739 ( .I(n2487), .ZN(n3214) );
  XOR2_X1 U20740 ( .A1(n2485), .A2(n2486), .Z(n8517) );
  INV_X1 U20745 ( .I(n51606), .ZN(n2489) );
  AOI21_X1 U20746 ( .A1(n2493), .A2(n54926), .B(n2490), .ZN(n54882) );
  NAND3_X1 U20747 ( .A1(n2491), .A2(n63022), .A3(n7680), .ZN(n2490) );
  XOR2_X1 U20748 ( .A1(n2494), .A2(n16452), .Z(n10019) );
  XOR2_X1 U20750 ( .A1(n11766), .A2(n15865), .Z(n2494) );
  NAND2_X1 U20753 ( .A1(n2499), .A2(n22574), .ZN(n48131) );
  NAND2_X1 U20754 ( .A1(n48472), .A2(n2499), .ZN(n14611) );
  NOR2_X1 U20757 ( .A1(n14521), .A2(n2499), .ZN(n8870) );
  XOR2_X1 U20759 ( .A1(n2500), .A2(n22795), .Z(n51605) );
  XOR2_X1 U20760 ( .A1(n26028), .A2(n23218), .Z(n2500) );
  NOR2_X2 U20761 ( .A1(n2502), .A2(n2501), .ZN(n26028) );
  INV_X2 U20762 ( .I(n38648), .ZN(n25277) );
  XOR2_X1 U20766 ( .A1(n2505), .A2(n1679), .Z(n2504) );
  XOR2_X1 U20767 ( .A1(n1684), .A2(n46426), .Z(n2505) );
  XOR2_X1 U20768 ( .A1(n60350), .A2(n46429), .Z(n2506) );
  INV_X1 U20769 ( .I(n9274), .ZN(n36555) );
  OR2_X1 U20771 ( .A1(n34780), .A2(n19457), .Z(n2510) );
  NAND2_X1 U20775 ( .A1(n36639), .A2(n2512), .ZN(n36644) );
  NAND2_X1 U20776 ( .A1(n2513), .A2(n60171), .ZN(n27376) );
  NAND3_X1 U20777 ( .A1(n2514), .A2(n49117), .A3(n49790), .ZN(n20979) );
  AOI21_X1 U20779 ( .A1(n45997), .A2(n2514), .B(n48443), .ZN(n45998) );
  NAND2_X1 U20783 ( .A1(n4336), .A2(n63020), .ZN(n8307) );
  INV_X1 U20788 ( .I(n30846), .ZN(n2519) );
  NOR2_X1 U20789 ( .A1(n23589), .A2(n21512), .ZN(n30846) );
  XOR2_X1 U20792 ( .A1(n2191), .A2(n15615), .Z(n2522) );
  INV_X1 U20793 ( .I(n2524), .ZN(n55298) );
  NAND2_X1 U20795 ( .A1(n2524), .A2(n55685), .ZN(n19902) );
  NAND3_X1 U20797 ( .A1(n55696), .A2(n2524), .A3(n55684), .ZN(n19903) );
  XOR2_X1 U20807 ( .A1(n57630), .A2(n43723), .Z(n43724) );
  XOR2_X1 U20809 ( .A1(n13359), .A2(n2540), .Z(n9007) );
  NAND2_X1 U20812 ( .A1(n58645), .A2(n4780), .ZN(n2543) );
  INV_X4 U20814 ( .I(n58645), .ZN(n20971) );
  NAND2_X2 U20817 ( .A1(n27406), .A2(n27970), .ZN(n2907) );
  XOR2_X1 U20819 ( .A1(n31519), .A2(n2551), .Z(n2550) );
  XOR2_X1 U20820 ( .A1(n8625), .A2(n57435), .Z(n2551) );
  XOR2_X1 U20822 ( .A1(n14866), .A2(n21779), .Z(n2553) );
  NAND2_X2 U20828 ( .A1(n21945), .A2(n34127), .ZN(n2695) );
  XOR2_X1 U20829 ( .A1(n8979), .A2(n44828), .Z(n2565) );
  XOR2_X1 U20830 ( .A1(n44821), .A2(n6715), .Z(n2567) );
  OAI21_X1 U20831 ( .A1(n5645), .A2(n2568), .B(n1901), .ZN(n5644) );
  NAND2_X1 U20832 ( .A1(n3117), .A2(n2569), .ZN(n3331) );
  NAND2_X1 U20835 ( .A1(n28418), .A2(n58792), .ZN(n28419) );
  NAND2_X1 U20836 ( .A1(n27088), .A2(n2569), .ZN(n22965) );
  NOR2_X1 U20837 ( .A1(n2571), .A2(n47894), .ZN(n17367) );
  NOR2_X1 U20838 ( .A1(n2571), .A2(n47900), .ZN(n17970) );
  INV_X1 U20840 ( .I(n2571), .ZN(n2570) );
  INV_X4 U20842 ( .I(n2572), .ZN(n24948) );
  INV_X2 U20845 ( .I(n2574), .ZN(n2960) );
  NAND3_X2 U20847 ( .A1(n42612), .A2(n42610), .A3(n42611), .ZN(n10339) );
  INV_X2 U20849 ( .I(n7602), .ZN(n13664) );
  INV_X2 U20864 ( .I(n20770), .ZN(n25522) );
  NAND2_X2 U20866 ( .A1(n23701), .A2(n53226), .ZN(n53009) );
  NOR2_X2 U20868 ( .A1(n3696), .A2(n2588), .ZN(n2797) );
  OAI21_X1 U20869 ( .A1(n7516), .A2(n3696), .B(n2588), .ZN(n43246) );
  NOR2_X1 U20870 ( .A1(n43144), .A2(n2588), .ZN(n26190) );
  NOR2_X1 U20876 ( .A1(n63532), .A2(n29153), .ZN(n3823) );
  OAI22_X1 U20877 ( .A1(n27976), .A2(n6522), .B1(n65111), .B2(n29152), .ZN(
        n27979) );
  AOI22_X1 U20880 ( .A1(n29151), .A2(n27392), .B1(n29150), .B2(n63532), .ZN(
        n27258) );
  XOR2_X1 U20882 ( .A1(n2596), .A2(n44355), .Z(n25363) );
  XOR2_X1 U20883 ( .A1(n2597), .A2(n15355), .Z(n2596) );
  NAND3_X1 U20884 ( .A1(n43249), .A2(n43248), .A3(n44097), .ZN(n2598) );
  INV_X1 U20885 ( .I(n2600), .ZN(n2599) );
  AOI21_X1 U20886 ( .A1(n43249), .A2(n43248), .B(n44097), .ZN(n2600) );
  NAND2_X2 U20887 ( .A1(n25148), .A2(n20090), .ZN(n7318) );
  XOR2_X1 U20888 ( .A1(n38819), .A2(n2601), .Z(n38081) );
  XOR2_X1 U20889 ( .A1(n60489), .A2(n2602), .Z(n2601) );
  XOR2_X1 U20890 ( .A1(n18452), .A2(n38577), .Z(n2602) );
  NAND2_X1 U20897 ( .A1(n2607), .A2(n22461), .ZN(n37430) );
  NOR2_X1 U20898 ( .A1(n35935), .A2(n2607), .ZN(n34810) );
  NOR2_X2 U20900 ( .A1(n8177), .A2(n63549), .ZN(n2607) );
  NAND3_X1 U20902 ( .A1(n49476), .A2(n260), .A3(n2608), .ZN(n49478) );
  XOR2_X1 U20905 ( .A1(n24178), .A2(n32282), .Z(n2612) );
  NAND2_X2 U20910 ( .A1(n20381), .A2(n53695), .ZN(n2619) );
  XOR2_X1 U20911 ( .A1(n2620), .A2(n1048), .Z(n6844) );
  XOR2_X1 U20912 ( .A1(n2621), .A2(n7778), .Z(n2620) );
  XOR2_X1 U20913 ( .A1(n2622), .A2(n11185), .Z(n2621) );
  NOR2_X2 U20922 ( .A1(n17922), .A2(n34035), .ZN(n34045) );
  NAND2_X1 U20923 ( .A1(n61622), .A2(n2636), .ZN(n2846) );
  XOR2_X1 U20924 ( .A1(n2638), .A2(n44800), .Z(n2637) );
  XOR2_X1 U20925 ( .A1(n62136), .A2(n44798), .Z(n2638) );
  NOR3_X1 U20926 ( .A1(n27968), .A2(n27405), .A3(n60298), .ZN(n2639) );
  XOR2_X1 U20936 ( .A1(n11620), .A2(n15087), .Z(n2650) );
  XOR2_X1 U20937 ( .A1(n20469), .A2(n32186), .Z(n32715) );
  XOR2_X1 U20938 ( .A1(n32292), .A2(n32186), .Z(n3878) );
  NOR3_X2 U20940 ( .A1(n2651), .A2(n5983), .A3(n24851), .ZN(n24868) );
  NOR3_X2 U20943 ( .A1(n2660), .A2(n2659), .A3(n2654), .ZN(n7022) );
  NOR2_X1 U20944 ( .A1(n24940), .A2(n23591), .ZN(n2658) );
  NAND2_X2 U20945 ( .A1(n18231), .A2(n6913), .ZN(n6519) );
  INV_X2 U20946 ( .I(n7006), .ZN(n17047) );
  NOR2_X1 U20949 ( .A1(n46946), .A2(n2664), .ZN(n46053) );
  INV_X2 U20951 ( .I(n2665), .ZN(n40193) );
  NAND2_X2 U20953 ( .A1(n40193), .A2(n1238), .ZN(n40200) );
  NAND3_X2 U20955 ( .A1(n10751), .A2(n10752), .A3(n15918), .ZN(n24243) );
  XOR2_X1 U20960 ( .A1(n44611), .A2(n2669), .Z(n6571) );
  XOR2_X1 U20961 ( .A1(n63667), .A2(n44618), .Z(n2669) );
  XOR2_X1 U20962 ( .A1(n59694), .A2(n2036), .Z(n44611) );
  NAND3_X1 U20975 ( .A1(n2675), .A2(n54960), .A3(n55089), .ZN(n55090) );
  AOI22_X1 U20976 ( .A1(n55098), .A2(n2675), .B1(n4087), .B2(n5051), .ZN(n4416) );
  OAI21_X1 U20979 ( .A1(n2676), .A2(n54395), .B(n54408), .ZN(n54399) );
  XOR2_X1 U20982 ( .A1(n2677), .A2(n8539), .Z(n25144) );
  XOR2_X1 U20984 ( .A1(n63008), .A2(n6307), .Z(n2677) );
  XOR2_X1 U20986 ( .A1(n61137), .A2(n3741), .Z(n50575) );
  NOR2_X1 U20988 ( .A1(n54798), .A2(n25215), .ZN(n54296) );
  XOR2_X1 U20989 ( .A1(n2680), .A2(n11357), .Z(n25580) );
  XOR2_X1 U20990 ( .A1(n32505), .A2(n2681), .Z(n31346) );
  XOR2_X1 U20991 ( .A1(n32292), .A2(n2681), .Z(n13255) );
  XOR2_X1 U20992 ( .A1(n23768), .A2(n33150), .Z(n2681) );
  XOR2_X1 U20993 ( .A1(n37967), .A2(n2682), .Z(n6308) );
  NAND2_X1 U20999 ( .A1(n49751), .A2(n2692), .ZN(n5345) );
  NAND2_X1 U21000 ( .A1(n3237), .A2(n2692), .ZN(n3236) );
  AOI22_X1 U21001 ( .A1(n49159), .A2(n49160), .B1(n2692), .B2(n49229), .ZN(
        n49163) );
  NOR2_X1 U21008 ( .A1(n3971), .A2(n2810), .ZN(n49046) );
  NAND2_X2 U21011 ( .A1(n22409), .A2(n45728), .ZN(n10636) );
  NOR2_X1 U21012 ( .A1(n1504), .A2(n22617), .ZN(n9188) );
  NOR3_X1 U21013 ( .A1(n18241), .A2(n22786), .A3(n38497), .ZN(n36107) );
  NAND2_X1 U21014 ( .A1(n12575), .A2(n2698), .ZN(n53248) );
  AOI21_X1 U21015 ( .A1(n22889), .A2(n2698), .B(n61361), .ZN(n19637) );
  NOR2_X2 U21016 ( .A1(n4283), .A2(n1232), .ZN(n2698) );
  XOR2_X1 U21017 ( .A1(n2701), .A2(n2700), .Z(n35152) );
  XOR2_X1 U21018 ( .A1(n2703), .A2(n37496), .Z(n2700) );
  XOR2_X1 U21019 ( .A1(n57458), .A2(n61061), .Z(n37496) );
  NAND3_X1 U21021 ( .A1(n2706), .A2(n23039), .A3(n7886), .ZN(n28388) );
  OAI21_X1 U21022 ( .A1(n27562), .A2(n2706), .B(n27561), .ZN(n27563) );
  XOR2_X1 U21024 ( .A1(n2710), .A2(n6750), .Z(n25292) );
  XOR2_X1 U21025 ( .A1(n36903), .A2(n6749), .Z(n2710) );
  XOR2_X1 U21026 ( .A1(n920), .A2(n3754), .Z(n6749) );
  AOI21_X1 U21030 ( .A1(n2712), .A2(n50810), .B(n15415), .ZN(n50811) );
  XOR2_X1 U21034 ( .A1(n2714), .A2(n32342), .Z(n32343) );
  XOR2_X1 U21035 ( .A1(n2714), .A2(n32749), .Z(n32760) );
  XOR2_X1 U21036 ( .A1(n1823), .A2(n33204), .Z(n2714) );
  NAND2_X2 U21038 ( .A1(n2717), .A2(n2716), .ZN(n24151) );
  NAND2_X2 U21041 ( .A1(n36462), .A2(n36463), .ZN(n11081) );
  OAI21_X1 U21044 ( .A1(n34796), .A2(n2721), .B(n33759), .ZN(n33761) );
  NAND2_X2 U21045 ( .A1(n14111), .A2(n15588), .ZN(n2721) );
  XOR2_X1 U21050 ( .A1(n13801), .A2(n42984), .Z(n11858) );
  XOR2_X1 U21053 ( .A1(n22566), .A2(n32267), .Z(n32653) );
  NAND2_X2 U21054 ( .A1(n2727), .A2(n2726), .ZN(n32267) );
  INV_X1 U21055 ( .I(n9280), .ZN(n30089) );
  NAND2_X1 U21057 ( .A1(n21950), .A2(n2735), .ZN(n3003) );
  NOR2_X1 U21060 ( .A1(n24576), .A2(n2735), .ZN(n39431) );
  INV_X2 U21062 ( .I(n2737), .ZN(n47851) );
  XNOR2_X1 U21064 ( .A1(n43826), .A2(n43825), .ZN(n2737) );
  XOR2_X1 U21065 ( .A1(n2740), .A2(n2738), .Z(n25007) );
  XOR2_X1 U21066 ( .A1(n2739), .A2(n44116), .Z(n2738) );
  XOR2_X1 U21067 ( .A1(n43967), .A2(n43806), .Z(n2739) );
  NAND2_X1 U21071 ( .A1(n19834), .A2(n2742), .ZN(n19833) );
  NAND2_X1 U21075 ( .A1(n9328), .A2(n3150), .ZN(n9326) );
  OAI22_X1 U21080 ( .A1(n53679), .A2(n53687), .B1(n53678), .B2(n2746), .ZN(
        n53680) );
  AOI22_X1 U21081 ( .A1(n53675), .A2(n2746), .B1(n53688), .B2(n53673), .ZN(
        n53656) );
  NOR2_X1 U21082 ( .A1(n53646), .A2(n2746), .ZN(n11936) );
  NAND2_X2 U21083 ( .A1(n53700), .A2(n53688), .ZN(n2746) );
  NOR2_X2 U21089 ( .A1(n2757), .A2(n2756), .ZN(n22805) );
  NOR2_X1 U21092 ( .A1(n2760), .A2(n64475), .ZN(n41074) );
  NOR2_X1 U21093 ( .A1(n2760), .A2(n41083), .ZN(n2759) );
  INV_X2 U21095 ( .I(n25772), .ZN(n21008) );
  XOR2_X1 U21096 ( .A1(n2762), .A2(n738), .Z(n25772) );
  XOR2_X1 U21098 ( .A1(n1823), .A2(n30407), .Z(n2763) );
  OR2_X1 U21099 ( .A1(n34992), .A2(n2765), .Z(n2764) );
  INV_X2 U21100 ( .I(n2767), .ZN(n47467) );
  XOR2_X1 U21104 ( .A1(n1051), .A2(n3373), .Z(n44931) );
  XOR2_X1 U21106 ( .A1(n37002), .A2(n2771), .Z(n2770) );
  XOR2_X1 U21107 ( .A1(n2772), .A2(n37001), .Z(n2771) );
  XOR2_X1 U21108 ( .A1(n39735), .A2(n37382), .Z(n2772) );
  XOR2_X1 U21111 ( .A1(n38796), .A2(n20042), .Z(n6604) );
  XOR2_X1 U21112 ( .A1(n14967), .A2(n7614), .Z(n51302) );
  XOR2_X1 U21116 ( .A1(n1253), .A2(n1434), .Z(n13594) );
  XOR2_X1 U21120 ( .A1(n2781), .A2(n2780), .Z(n2779) );
  XOR2_X1 U21121 ( .A1(n31334), .A2(n23726), .Z(n31697) );
  XOR2_X1 U21122 ( .A1(n33866), .A2(n31332), .Z(n2781) );
  XOR2_X1 U21123 ( .A1(n2783), .A2(n33233), .Z(n2782) );
  XOR2_X1 U21124 ( .A1(n32479), .A2(n16273), .Z(n2783) );
  XOR2_X1 U21125 ( .A1(n31333), .A2(n32572), .Z(n32479) );
  AOI21_X1 U21126 ( .A1(n2784), .A2(n55147), .B(n55168), .ZN(n52647) );
  OAI22_X1 U21128 ( .A1(n1167), .A2(n55140), .B1(n7986), .B2(n2784), .ZN(n7985) );
  NAND2_X1 U21134 ( .A1(n24357), .A2(n24609), .ZN(n2792) );
  INV_X2 U21138 ( .I(n3256), .ZN(n2790) );
  NAND2_X2 U21139 ( .A1(n3117), .A2(n24951), .ZN(n3256) );
  NOR2_X2 U21142 ( .A1(n24852), .A2(n1557), .ZN(n30391) );
  INV_X2 U21145 ( .I(n2798), .ZN(n6417) );
  AND2_X2 U21146 ( .A1(n4413), .A2(n6417), .Z(n9758) );
  XOR2_X1 U21148 ( .A1(n19622), .A2(n31943), .Z(n21128) );
  NAND3_X2 U21149 ( .A1(n30379), .A2(n30381), .A3(n30380), .ZN(n31943) );
  NAND2_X2 U21152 ( .A1(n25553), .A2(n30399), .ZN(n31686) );
  XOR2_X1 U21156 ( .A1(n11426), .A2(n2804), .Z(n2803) );
  XOR2_X1 U21157 ( .A1(n51163), .A2(n22521), .Z(n11426) );
  XOR2_X1 U21159 ( .A1(n2805), .A2(n13574), .Z(n2804) );
  XOR2_X1 U21160 ( .A1(n50580), .A2(n19785), .Z(n2805) );
  INV_X2 U21161 ( .I(n2806), .ZN(n30294) );
  NAND2_X1 U21162 ( .A1(n12612), .A2(n2806), .ZN(n28926) );
  OAI22_X1 U21163 ( .A1(n28977), .A2(n2806), .B1(n10129), .B2(n11205), .ZN(
        n28978) );
  XOR2_X1 U21171 ( .A1(n2817), .A2(n38212), .Z(n2816) );
  NAND2_X1 U21175 ( .A1(n2820), .A2(n23856), .ZN(n52228) );
  INV_X2 U21177 ( .I(n2821), .ZN(n45400) );
  NAND3_X2 U21183 ( .A1(n60808), .A2(n32794), .A3(n32795), .ZN(n14308) );
  NAND2_X2 U21184 ( .A1(n6867), .A2(n34993), .ZN(n12350) );
  NAND2_X1 U21188 ( .A1(n53645), .A2(n53644), .ZN(n2831) );
  NOR2_X1 U21189 ( .A1(n53688), .A2(n53695), .ZN(n53666) );
  NAND2_X2 U21192 ( .A1(n53643), .A2(n53655), .ZN(n53644) );
  NOR2_X1 U21194 ( .A1(n29051), .A2(n30197), .ZN(n2841) );
  XOR2_X1 U21199 ( .A1(n2850), .A2(n12307), .Z(n25998) );
  XOR2_X1 U21213 ( .A1(n2863), .A2(n6040), .Z(n2858) );
  NOR2_X2 U21220 ( .A1(n54939), .A2(n21877), .ZN(n54945) );
  XOR2_X1 U21222 ( .A1(n52419), .A2(n52418), .Z(n52510) );
  XOR2_X1 U21223 ( .A1(n51418), .A2(n52202), .Z(n52419) );
  XOR2_X1 U21226 ( .A1(n19519), .A2(n50796), .Z(n24074) );
  NAND2_X1 U21227 ( .A1(n40845), .A2(n2325), .ZN(n40846) );
  NAND3_X1 U21228 ( .A1(n62357), .A2(n64592), .A3(n2325), .ZN(n41879) );
  OAI21_X1 U21229 ( .A1(n15890), .A2(n2867), .B(n41055), .ZN(n41056) );
  XOR2_X1 U21232 ( .A1(n31629), .A2(n16709), .Z(n18965) );
  XOR2_X1 U21237 ( .A1(n25794), .A2(n2950), .Z(n51924) );
  NAND2_X1 U21239 ( .A1(n2789), .A2(n28405), .ZN(n27092) );
  NAND2_X1 U21242 ( .A1(n2877), .A2(n16285), .ZN(n8312) );
  NAND2_X1 U21245 ( .A1(n541), .A2(n42681), .ZN(n42821) );
  NAND2_X2 U21248 ( .A1(n8911), .A2(n2879), .ZN(n42825) );
  NAND2_X2 U21251 ( .A1(n5212), .A2(n5211), .ZN(n2879) );
  XOR2_X1 U21252 ( .A1(n2880), .A2(n2882), .Z(n2894) );
  XOR2_X1 U21253 ( .A1(n2881), .A2(n44038), .Z(n2880) );
  XOR2_X1 U21254 ( .A1(n15216), .A2(n43674), .Z(n2882) );
  XOR2_X1 U21262 ( .A1(n11853), .A2(n26009), .Z(n2886) );
  NOR2_X1 U21265 ( .A1(n62663), .A2(n61035), .ZN(n17418) );
  NOR2_X1 U21267 ( .A1(n7719), .A2(n62663), .ZN(n23779) );
  NAND3_X1 U21268 ( .A1(n26251), .A2(n27959), .A3(n62663), .ZN(n26252) );
  NOR2_X1 U21269 ( .A1(n11892), .A2(n2889), .ZN(n11891) );
  NAND2_X1 U21271 ( .A1(n2890), .A2(n10938), .ZN(n17376) );
  NAND2_X1 U21272 ( .A1(n2890), .A2(n1453), .ZN(n51710) );
  NOR2_X1 U21273 ( .A1(n2890), .A2(n23704), .ZN(n54104) );
  NAND2_X1 U21276 ( .A1(n53870), .A2(n2890), .ZN(n49819) );
  NAND2_X1 U21280 ( .A1(n47749), .A2(n2894), .ZN(n47432) );
  XOR2_X1 U21282 ( .A1(n2896), .A2(n3475), .Z(n43867) );
  XOR2_X1 U21283 ( .A1(n3477), .A2(n4956), .Z(n2896) );
  OAI21_X1 U21286 ( .A1(n42719), .A2(n2898), .B(n42718), .ZN(n42720) );
  INV_X2 U21293 ( .I(n47799), .ZN(n47809) );
  NAND2_X2 U21294 ( .A1(n45199), .A2(n11417), .ZN(n47799) );
  NAND2_X1 U21297 ( .A1(n19151), .A2(n61405), .ZN(n2903) );
  NAND2_X2 U21300 ( .A1(n12197), .A2(n12199), .ZN(n49529) );
  XOR2_X1 U21303 ( .A1(n31063), .A2(n2906), .Z(n9319) );
  INV_X2 U21310 ( .I(n6832), .ZN(n6703) );
  XOR2_X1 U21311 ( .A1(n4947), .A2(n61450), .Z(n39628) );
  NAND2_X1 U21316 ( .A1(n14741), .A2(n61543), .ZN(n2914) );
  NAND3_X1 U21317 ( .A1(n24114), .A2(n47828), .A3(n15157), .ZN(n2916) );
  XOR2_X1 U21319 ( .A1(n2917), .A2(n5000), .Z(n4440) );
  XOR2_X1 U21320 ( .A1(n2917), .A2(n44279), .Z(n18065) );
  NAND2_X1 U21322 ( .A1(n35933), .A2(n2918), .ZN(n23546) );
  AND2_X1 U21327 ( .A1(n19359), .A2(n3211), .Z(n2920) );
  XOR2_X1 U21328 ( .A1(n22377), .A2(n26430), .Z(n19359) );
  NAND2_X1 U21329 ( .A1(n20179), .A2(n62999), .ZN(n17483) );
  NOR2_X2 U21333 ( .A1(n43569), .A2(n2994), .ZN(n43581) );
  INV_X2 U21336 ( .I(n2922), .ZN(n2989) );
  NAND2_X2 U21337 ( .A1(n2924), .A2(n2989), .ZN(n10526) );
  XNOR2_X1 U21338 ( .A1(n2992), .A2(n2990), .ZN(n2922) );
  XOR2_X1 U21340 ( .A1(n22940), .A2(n51588), .Z(n11507) );
  XOR2_X1 U21341 ( .A1(n22940), .A2(n11480), .Z(n11479) );
  NOR2_X1 U21342 ( .A1(n53041), .A2(n2925), .ZN(n20369) );
  AOI22_X2 U21346 ( .A1(n1521), .A2(n6781), .B1(n2928), .B2(n6782), .ZN(n14588) );
  XOR2_X1 U21349 ( .A1(n2930), .A2(n868), .Z(n2929) );
  XOR2_X1 U21350 ( .A1(n2934), .A2(n748), .Z(n2930) );
  XOR2_X1 U21353 ( .A1(n50833), .A2(n26072), .Z(n2934) );
  XOR2_X1 U21354 ( .A1(n52440), .A2(n62084), .Z(n2935) );
  XOR2_X1 U21356 ( .A1(n1819), .A2(n33191), .Z(n2937) );
  INV_X2 U21357 ( .I(n35329), .ZN(n3939) );
  XOR2_X1 U21360 ( .A1(n32120), .A2(n32117), .Z(n2939) );
  XOR2_X1 U21361 ( .A1(n32116), .A2(n32270), .Z(n2940) );
  INV_X2 U21363 ( .I(n27056), .ZN(n6215) );
  XOR2_X1 U21369 ( .A1(n2947), .A2(n44895), .Z(n8230) );
  XOR2_X1 U21370 ( .A1(n2998), .A2(n31757), .Z(n2947) );
  XOR2_X1 U21377 ( .A1(n64095), .A2(n52607), .Z(n14862) );
  XOR2_X1 U21378 ( .A1(n2876), .A2(n45475), .Z(n45476) );
  XOR2_X1 U21379 ( .A1(n23758), .A2(n64095), .Z(n23939) );
  XOR2_X1 U21380 ( .A1(n2876), .A2(n52321), .Z(n50839) );
  XOR2_X1 U21382 ( .A1(n22584), .A2(n2876), .Z(n24031) );
  NOR2_X2 U21383 ( .A1(n2754), .A2(n22533), .ZN(n50428) );
  NAND2_X2 U21384 ( .A1(n54102), .A2(n2951), .ZN(n54108) );
  INV_X2 U21391 ( .I(n39841), .ZN(n43225) );
  NAND2_X2 U21396 ( .A1(n37181), .A2(n2958), .ZN(n5442) );
  NAND2_X1 U21397 ( .A1(n61574), .A2(n64620), .ZN(n32144) );
  XOR2_X1 U21398 ( .A1(n63343), .A2(n51335), .Z(n51744) );
  XOR2_X1 U21399 ( .A1(n63343), .A2(n9154), .Z(n50907) );
  XOR2_X1 U21400 ( .A1(n63343), .A2(n10344), .Z(n11861) );
  INV_X2 U21401 ( .I(n41889), .ZN(n41065) );
  NOR2_X2 U21402 ( .A1(n40842), .A2(n2867), .ZN(n41889) );
  XOR2_X1 U21403 ( .A1(n2952), .A2(n32082), .Z(n32083) );
  INV_X2 U21405 ( .I(n2961), .ZN(n17919) );
  NAND2_X1 U21411 ( .A1(n2962), .A2(n35410), .ZN(n35411) );
  NAND2_X2 U21415 ( .A1(n2965), .A2(n29747), .ZN(n30782) );
  NOR2_X2 U21418 ( .A1(n3023), .A2(n9687), .ZN(n2968) );
  INV_X2 U21419 ( .I(n57173), .ZN(n10554) );
  NOR2_X1 U21424 ( .A1(n22726), .A2(n2971), .ZN(n3822) );
  NOR2_X2 U21425 ( .A1(n29154), .A2(n27397), .ZN(n2971) );
  NAND3_X1 U21430 ( .A1(n3637), .A2(n3638), .A3(n2973), .ZN(n45552) );
  XOR2_X1 U21434 ( .A1(n28983), .A2(n24756), .Z(n26178) );
  XOR2_X1 U21440 ( .A1(n2991), .A2(n21642), .Z(n2990) );
  XOR2_X1 U21442 ( .A1(n5981), .A2(n17182), .Z(n2993) );
  NOR2_X1 U21444 ( .A1(n2996), .A2(n11263), .ZN(n28956) );
  OAI22_X1 U21445 ( .A1(n28958), .A2(n15593), .B1(n2996), .B2(n29442), .ZN(
        n15592) );
  NOR2_X2 U21446 ( .A1(n14202), .A2(n31129), .ZN(n2996) );
  NAND2_X2 U21456 ( .A1(n34203), .A2(n61517), .ZN(n8041) );
  INV_X4 U21457 ( .I(n23766), .ZN(n6918) );
  NOR2_X2 U21458 ( .A1(n34161), .A2(n23947), .ZN(n15028) );
  XOR2_X1 U21460 ( .A1(n3244), .A2(n37123), .Z(n3015) );
  XOR2_X1 U21464 ( .A1(n3018), .A2(n44294), .Z(n18214) );
  XOR2_X1 U21465 ( .A1(n3019), .A2(n18139), .Z(n44294) );
  XOR2_X1 U21466 ( .A1(n15773), .A2(n44731), .Z(n3019) );
  NAND2_X1 U21469 ( .A1(n56936), .A2(n3021), .ZN(n56939) );
  AOI22_X1 U21470 ( .A1(n56918), .A2(n56957), .B1(n56917), .B2(n3021), .ZN(
        n56922) );
  NAND2_X1 U21471 ( .A1(n3022), .A2(n27022), .ZN(n27023) );
  NOR2_X1 U21472 ( .A1(n3022), .A2(n57872), .ZN(n28042) );
  NOR2_X1 U21474 ( .A1(n34520), .A2(n3023), .ZN(n24544) );
  XNOR2_X1 U21479 ( .A1(Ciphertext[38]), .A2(Key[63]), .ZN(n3027) );
  XOR2_X1 U21485 ( .A1(n25660), .A2(n44504), .Z(n3033) );
  XOR2_X1 U21488 ( .A1(n44973), .A2(n56949), .Z(n3037) );
  INV_X2 U21490 ( .I(n3039), .ZN(n24749) );
  INV_X2 U21491 ( .I(n24748), .ZN(n55486) );
  INV_X2 U21494 ( .I(n41147), .ZN(n4819) );
  NAND2_X2 U21496 ( .A1(n3055), .A2(n50056), .ZN(n50058) );
  NOR2_X2 U21499 ( .A1(n7952), .A2(n1643), .ZN(n3123) );
  OR3_X1 U21501 ( .A1(n15436), .A2(n50308), .A3(n50304), .Z(n3046) );
  NOR2_X2 U21514 ( .A1(n3050), .A2(n3049), .ZN(n15045) );
  XOR2_X1 U21518 ( .A1(n25854), .A2(n24886), .Z(n11737) );
  NAND2_X1 U21519 ( .A1(n3052), .A2(n16694), .ZN(n29418) );
  NAND2_X1 U21520 ( .A1(n1839), .A2(n28092), .ZN(n13573) );
  AOI21_X1 U21521 ( .A1(n30440), .A2(n30439), .B(n3052), .ZN(n30446) );
  XOR2_X1 U21522 ( .A1(n37699), .A2(n37701), .Z(n5786) );
  NOR2_X2 U21532 ( .A1(n34563), .A2(n34562), .ZN(n8697) );
  NAND2_X2 U21533 ( .A1(n24195), .A2(n43242), .ZN(n13037) );
  XOR2_X1 U21538 ( .A1(n37801), .A2(n3069), .Z(n37886) );
  XOR2_X1 U21542 ( .A1(n3071), .A2(n853), .Z(n12505) );
  XOR2_X1 U21545 ( .A1(n3073), .A2(n767), .Z(n18562) );
  XOR2_X1 U21546 ( .A1(n8228), .A2(n3334), .Z(n3073) );
  OAI21_X1 U21550 ( .A1(n22474), .A2(n3076), .B(n18313), .ZN(n8762) );
  NOR2_X1 U21552 ( .A1(n54590), .A2(n3077), .ZN(n6464) );
  NOR2_X2 U21553 ( .A1(n3769), .A2(n54087), .ZN(n3077) );
  NOR2_X2 U21555 ( .A1(n22776), .A2(n3078), .ZN(n41248) );
  AOI21_X1 U21557 ( .A1(n42275), .A2(n42286), .B(n3078), .ZN(n42278) );
  INV_X2 U21559 ( .I(n3080), .ZN(n46049) );
  OR2_X2 U21573 ( .A1(n1203), .A2(n24850), .Z(n48614) );
  XOR2_X1 U21575 ( .A1(n2952), .A2(n45359), .Z(n24095) );
  OAI22_X1 U21578 ( .A1(n3098), .A2(n60162), .B1(n60170), .B2(n21159), .ZN(
        n21604) );
  INV_X2 U21579 ( .I(n5265), .ZN(n48103) );
  XOR2_X1 U21583 ( .A1(n3101), .A2(n19854), .Z(n25595) );
  NOR3_X2 U21584 ( .A1(n3103), .A2(n35489), .A3(n3102), .ZN(n12491) );
  XOR2_X1 U21589 ( .A1(n3104), .A2(n12507), .Z(n45284) );
  XOR2_X1 U21590 ( .A1(n3104), .A2(n16518), .Z(n46322) );
  XOR2_X1 U21591 ( .A1(n3104), .A2(n23534), .Z(n42179) );
  XOR2_X1 U21592 ( .A1(n42715), .A2(n3104), .Z(n18900) );
  NOR2_X1 U21595 ( .A1(n8218), .A2(n1317), .ZN(n21358) );
  NAND2_X2 U21596 ( .A1(n39106), .A2(n40951), .ZN(n3109) );
  NAND2_X1 U21598 ( .A1(n3111), .A2(n48471), .ZN(n48477) );
  AOI21_X1 U21600 ( .A1(n48466), .A2(n3111), .B(n48465), .ZN(n48470) );
  XOR2_X1 U21604 ( .A1(n10442), .A2(n19013), .Z(n3113) );
  XOR2_X1 U21607 ( .A1(n19411), .A2(n46421), .Z(n3116) );
  NOR3_X1 U21608 ( .A1(n36938), .A2(n35426), .A3(n1421), .ZN(n24963) );
  XOR2_X1 U21610 ( .A1(Ciphertext[30]), .A2(Key[7]), .Z(n3385) );
  XNOR2_X1 U21612 ( .A1(n25794), .A2(n52107), .ZN(n3118) );
  NAND2_X2 U21613 ( .A1(n4013), .A2(n4010), .ZN(n52107) );
  NAND2_X1 U21618 ( .A1(n9523), .A2(n20922), .ZN(n9522) );
  AND2_X1 U21619 ( .A1(n3122), .A2(n33437), .Z(n16229) );
  NOR2_X2 U21620 ( .A1(n1342), .A2(n10064), .ZN(n10358) );
  NAND2_X2 U21621 ( .A1(n61749), .A2(n34586), .ZN(n17420) );
  NAND3_X1 U21623 ( .A1(n50140), .A2(n3123), .A3(n50141), .ZN(n50146) );
  XOR2_X1 U21627 ( .A1(n63024), .A2(n22922), .Z(n11167) );
  INV_X2 U21632 ( .I(n9967), .ZN(n12129) );
  NAND2_X2 U21635 ( .A1(n52786), .A2(n7095), .ZN(n3127) );
  XOR2_X1 U21639 ( .A1(n3136), .A2(n13244), .Z(n12772) );
  XOR2_X1 U21642 ( .A1(n9615), .A2(n51003), .Z(n3139) );
  INV_X2 U21646 ( .I(n3142), .ZN(n39324) );
  XOR2_X1 U21650 ( .A1(n3354), .A2(n10795), .Z(n3145) );
  XOR2_X1 U21651 ( .A1(n5440), .A2(n5438), .Z(n3142) );
  NOR2_X1 U21659 ( .A1(n35980), .A2(n58853), .ZN(n36709) );
  NAND2_X1 U21661 ( .A1(n34205), .A2(n58853), .ZN(n34206) );
  NAND2_X2 U21666 ( .A1(n50427), .A2(n50426), .ZN(n49256) );
  AOI22_X1 U21667 ( .A1(n34904), .A2(n36947), .B1(n34902), .B2(n34903), .ZN(
        n3154) );
  NAND4_X2 U21671 ( .A1(n3155), .A2(n34919), .A3(n34918), .A4(n3154), .ZN(
        n38770) );
  XOR2_X1 U21676 ( .A1(n3162), .A2(n3159), .Z(n12151) );
  XOR2_X1 U21677 ( .A1(n46611), .A2(n3161), .Z(n3159) );
  XOR2_X1 U21680 ( .A1(n25244), .A2(n43974), .Z(n3161) );
  XOR2_X1 U21681 ( .A1(n45271), .A2(n46680), .Z(n3162) );
  XOR2_X1 U21682 ( .A1(Ciphertext[32]), .A2(Key[21]), .Z(n3177) );
  INV_X2 U21683 ( .I(n6241), .ZN(n6747) );
  INV_X2 U21684 ( .I(n5833), .ZN(n12249) );
  XOR2_X1 U21687 ( .A1(n10024), .A2(n3163), .Z(n15489) );
  XOR2_X1 U21689 ( .A1(n23690), .A2(n33034), .Z(n3164) );
  XOR2_X1 U21690 ( .A1(n31385), .A2(n24283), .Z(n3165) );
  AOI22_X1 U21694 ( .A1(n4036), .A2(n37230), .B1(n3171), .B2(n36350), .ZN(
        n36354) );
  NAND2_X1 U21701 ( .A1(n33017), .A2(n33597), .ZN(n3173) );
  INV_X2 U21704 ( .I(n24701), .ZN(n28410) );
  XOR2_X1 U21705 ( .A1(n24702), .A2(Key[138]), .Z(n24701) );
  INV_X2 U21706 ( .I(n3177), .ZN(n24039) );
  AOI21_X1 U21710 ( .A1(n30394), .A2(n3180), .B(n30393), .ZN(n30397) );
  NAND4_X1 U21711 ( .A1(n1500), .A2(n1499), .A3(n42355), .A4(n41980), .ZN(
        n41617) );
  XOR2_X1 U21714 ( .A1(n3183), .A2(n3518), .Z(n3182) );
  XOR2_X1 U21717 ( .A1(n50620), .A2(n25969), .Z(n3185) );
  XOR2_X1 U21720 ( .A1(n7388), .A2(n63009), .Z(n3187) );
  OAI21_X1 U21721 ( .A1(n3188), .A2(n7956), .B(n54904), .ZN(n54903) );
  AOI21_X1 U21722 ( .A1(n12690), .A2(n54930), .B(n3188), .ZN(n12689) );
  OAI21_X1 U21723 ( .A1(n54927), .A2(n3188), .B(n54926), .ZN(n54933) );
  XOR2_X1 U21726 ( .A1(n3191), .A2(n7528), .Z(n3190) );
  XOR2_X1 U21727 ( .A1(n61178), .A2(n6336), .Z(n3191) );
  XOR2_X1 U21728 ( .A1(n52631), .A2(n21700), .Z(n52413) );
  XOR2_X1 U21729 ( .A1(n7847), .A2(n8076), .Z(n52631) );
  XNOR2_X1 U21732 ( .A1(n50036), .A2(n8674), .ZN(n12119) );
  NAND3_X2 U21735 ( .A1(n3201), .A2(n3199), .A3(n3196), .ZN(n28792) );
  NAND2_X1 U21736 ( .A1(n59670), .A2(n6933), .ZN(n47322) );
  NAND2_X1 U21737 ( .A1(n3203), .A2(n47307), .ZN(n45620) );
  NAND2_X1 U21739 ( .A1(n43984), .A2(n3204), .ZN(n43987) );
  NAND2_X1 U21740 ( .A1(n3204), .A2(n16880), .ZN(n43993) );
  OAI21_X1 U21741 ( .A1(n43985), .A2(n3204), .B(n43306), .ZN(n43307) );
  AOI21_X2 U21745 ( .A1(n54838), .A2(n6235), .B(n52477), .ZN(n54871) );
  NOR2_X2 U21746 ( .A1(n3207), .A2(n3206), .ZN(n8348) );
  AOI21_X1 U21747 ( .A1(n54845), .A2(n54844), .B(n54843), .ZN(n3206) );
  NAND3_X2 U21748 ( .A1(n20173), .A2(n3210), .A3(n3209), .ZN(n6136) );
  INV_X2 U21749 ( .I(n26802), .ZN(n28533) );
  XOR2_X1 U21751 ( .A1(n3212), .A2(Ciphertext[98]), .Z(n26802) );
  INV_X1 U21752 ( .I(Key[99]), .ZN(n3212) );
  INV_X2 U21753 ( .I(n3213), .ZN(n7728) );
  XOR2_X1 U21755 ( .A1(n12015), .A2(n9415), .Z(n38491) );
  NAND2_X2 U21756 ( .A1(n34278), .A2(n15927), .ZN(n3325) );
  NAND2_X2 U21757 ( .A1(n1815), .A2(n32972), .ZN(n34278) );
  NAND2_X2 U21762 ( .A1(n20004), .A2(n7086), .ZN(n8679) );
  NAND2_X2 U21763 ( .A1(n10498), .A2(n36471), .ZN(n3218) );
  NAND2_X2 U21764 ( .A1(n23542), .A2(n48481), .ZN(n48177) );
  NAND2_X2 U21766 ( .A1(n23813), .A2(n24185), .ZN(n48176) );
  NAND3_X2 U21768 ( .A1(n3224), .A2(n3223), .A3(n3222), .ZN(n36579) );
  XOR2_X1 U21771 ( .A1(n3231), .A2(n3230), .Z(n3229) );
  XOR2_X1 U21772 ( .A1(n3244), .A2(n38257), .Z(n3230) );
  NOR3_X2 U21778 ( .A1(n3240), .A2(n5567), .A3(n3235), .ZN(n25535) );
  NAND2_X2 U21781 ( .A1(n34783), .A2(n1430), .ZN(n19894) );
  XOR2_X1 U21782 ( .A1(n32267), .A2(n3242), .Z(n7397) );
  XOR2_X1 U21786 ( .A1(n3248), .A2(n934), .Z(n3247) );
  NAND2_X2 U21791 ( .A1(n3251), .A2(n55387), .ZN(n16503) );
  NAND2_X2 U21793 ( .A1(n3250), .A2(n55389), .ZN(n55372) );
  NOR2_X2 U21795 ( .A1(n9421), .A2(n3251), .ZN(n55382) );
  INV_X2 U21796 ( .I(n24529), .ZN(n3251) );
  XOR2_X1 U21799 ( .A1(n61947), .A2(n38366), .Z(n4073) );
  INV_X2 U21800 ( .I(n3257), .ZN(n13029) );
  XOR2_X1 U21802 ( .A1(n7811), .A2(n16883), .Z(n46528) );
  XOR2_X1 U21803 ( .A1(n16898), .A2(n16899), .Z(n3259) );
  NAND2_X1 U21807 ( .A1(n3266), .A2(n14202), .ZN(n3264) );
  NOR2_X2 U21808 ( .A1(n27797), .A2(n29916), .ZN(n29434) );
  NOR2_X1 U21810 ( .A1(n6041), .A2(n3267), .ZN(n3266) );
  INV_X1 U21811 ( .I(n29916), .ZN(n3267) );
  NAND2_X2 U21812 ( .A1(n29915), .A2(n4706), .ZN(n31127) );
  INV_X1 U21813 ( .I(n58765), .ZN(n29559) );
  NOR2_X2 U21814 ( .A1(n25269), .A2(n29432), .ZN(n6041) );
  XOR2_X1 U21815 ( .A1(n3268), .A2(n1268), .Z(n44768) );
  INV_X1 U21818 ( .I(n22143), .ZN(n3269) );
  INV_X2 U21822 ( .I(n3272), .ZN(n34149) );
  XOR2_X1 U21830 ( .A1(n3279), .A2(n3277), .Z(n19713) );
  XOR2_X1 U21831 ( .A1(n10802), .A2(n3480), .Z(n38361) );
  XOR2_X1 U21833 ( .A1(n11005), .A2(n24169), .Z(n3279) );
  NAND2_X1 U21836 ( .A1(n2820), .A2(n3285), .ZN(n53157) );
  AOI21_X1 U21837 ( .A1(n53136), .A2(n3285), .B(n53135), .ZN(n3507) );
  OAI21_X2 U21842 ( .A1(n48460), .A2(n47208), .B(n48463), .ZN(n3289) );
  XOR2_X1 U21846 ( .A1(n17919), .A2(n8158), .Z(n3291) );
  INV_X1 U21848 ( .I(n12015), .ZN(n12068) );
  NAND2_X2 U21849 ( .A1(n3299), .A2(n3296), .ZN(n32515) );
  XOR2_X1 U21850 ( .A1(n23259), .A2(n32515), .Z(n32165) );
  INV_X1 U21852 ( .I(n3303), .ZN(n50012) );
  NAND2_X1 U21853 ( .A1(n50011), .A2(n3303), .ZN(n25504) );
  AOI21_X1 U21854 ( .A1(n3303), .A2(n49348), .B(n49345), .ZN(n49346) );
  OAI21_X1 U21857 ( .A1(n11044), .A2(n3306), .B(n3305), .ZN(n9202) );
  OAI21_X1 U21858 ( .A1(n11043), .A2(n11042), .B(n3306), .ZN(n3305) );
  NAND2_X2 U21860 ( .A1(n21411), .A2(n21410), .ZN(n23646) );
  NAND2_X1 U21863 ( .A1(n34776), .A2(n3308), .ZN(n34778) );
  XOR2_X1 U21871 ( .A1(n10994), .A2(n3318), .Z(n10993) );
  XOR2_X1 U21873 ( .A1(n3323), .A2(n3324), .Z(n3322) );
  XOR2_X1 U21874 ( .A1(n11736), .A2(n11735), .Z(n3323) );
  NAND2_X2 U21875 ( .A1(n1203), .A2(n24850), .ZN(n9140) );
  XOR2_X1 U21876 ( .A1(n18890), .A2(n46322), .Z(n3324) );
  XOR2_X1 U21878 ( .A1(n32045), .A2(n3329), .Z(n12504) );
  XOR2_X1 U21879 ( .A1(n31998), .A2(n12520), .Z(n3329) );
  XOR2_X1 U21880 ( .A1(n32044), .A2(n32412), .Z(n31998) );
  NAND2_X2 U21881 ( .A1(n30328), .A2(n24671), .ZN(n32044) );
  NAND2_X2 U21885 ( .A1(n1893), .A2(n58927), .ZN(n8202) );
  XOR2_X1 U21887 ( .A1(n3333), .A2(n15649), .Z(n11165) );
  XOR2_X1 U21891 ( .A1(n23173), .A2(n3333), .Z(n50202) );
  XOR2_X1 U21892 ( .A1(n4265), .A2(n3334), .Z(n50704) );
  XOR2_X1 U21895 ( .A1(n10678), .A2(n3339), .Z(n11734) );
  NAND2_X2 U21898 ( .A1(n3345), .A2(n40595), .ZN(n7907) );
  INV_X2 U21903 ( .I(n3346), .ZN(n6889) );
  CLKBUF_X4 U21907 ( .I(n48676), .Z(n3348) );
  NOR2_X2 U21912 ( .A1(n42709), .A2(n22554), .ZN(n20754) );
  XOR2_X1 U21913 ( .A1(n43866), .A2(n3474), .Z(n3353) );
  NAND3_X1 U21917 ( .A1(n40150), .A2(n59062), .A3(n61005), .ZN(n25865) );
  XOR2_X1 U21923 ( .A1(n21100), .A2(n3334), .Z(n12791) );
  XOR2_X1 U21924 ( .A1(n18854), .A2(n3334), .Z(n52371) );
  NAND2_X1 U21928 ( .A1(n14308), .A2(n3363), .ZN(n20063) );
  AOI21_X1 U21929 ( .A1(n34121), .A2(n34122), .B(n3363), .ZN(n34123) );
  NAND2_X1 U21934 ( .A1(n16846), .A2(n5570), .ZN(n8062) );
  INV_X2 U21935 ( .I(n4898), .ZN(n9067) );
  NAND2_X1 U21936 ( .A1(n674), .A2(n9067), .ZN(n9066) );
  INV_X2 U21940 ( .I(n55088), .ZN(n55101) );
  XOR2_X1 U21941 ( .A1(n44539), .A2(n3374), .Z(n3373) );
  XOR2_X1 U21942 ( .A1(n44254), .A2(n3449), .Z(n3374) );
  XOR2_X1 U21943 ( .A1(n45015), .A2(n44735), .Z(n3517) );
  XOR2_X1 U21944 ( .A1(n14299), .A2(n3375), .Z(n3690) );
  XOR2_X1 U21946 ( .A1(n61538), .A2(n32095), .Z(n20670) );
  XOR2_X1 U21947 ( .A1(n31599), .A2(n54587), .Z(n9977) );
  XOR2_X1 U21953 ( .A1(n3717), .A2(n22344), .Z(n3380) );
  INV_X2 U21955 ( .I(n6116), .ZN(n25213) );
  XOR2_X1 U21969 ( .A1(n11310), .A2(n3396), .Z(n3395) );
  XOR2_X1 U21970 ( .A1(n38711), .A2(n10499), .Z(n11310) );
  NAND2_X2 U21975 ( .A1(n3398), .A2(n11210), .ZN(n38072) );
  NAND3_X1 U21981 ( .A1(n41263), .A2(n64768), .A3(n4635), .ZN(n40798) );
  NOR2_X2 U21984 ( .A1(n3410), .A2(n3404), .ZN(n8470) );
  INV_X2 U21986 ( .I(n13173), .ZN(n24068) );
  XOR2_X1 U21989 ( .A1(n13173), .A2(n22923), .Z(n3416) );
  XOR2_X1 U21990 ( .A1(n3418), .A2(n44498), .Z(n3417) );
  XOR2_X1 U21992 ( .A1(n17112), .A2(n3419), .Z(n11842) );
  XOR2_X1 U21994 ( .A1(n24258), .A2(n13181), .Z(n3420) );
  XOR2_X1 U21995 ( .A1(n18490), .A2(n3422), .Z(n3421) );
  XOR2_X1 U21996 ( .A1(n23343), .A2(n840), .Z(n3422) );
  XOR2_X1 U21999 ( .A1(n19220), .A2(n11529), .Z(n3424) );
  INV_X2 U22002 ( .I(n3427), .ZN(n14424) );
  NAND2_X1 U22003 ( .A1(n3428), .A2(n28652), .ZN(n28645) );
  XOR2_X1 U22004 ( .A1(n3429), .A2(n39490), .Z(n22299) );
  XOR2_X1 U22005 ( .A1(n3429), .A2(n36321), .Z(n36322) );
  XOR2_X1 U22006 ( .A1(n3429), .A2(n38833), .Z(n38834) );
  XOR2_X1 U22008 ( .A1(n24908), .A2(n3430), .Z(n33054) );
  INV_X1 U22009 ( .I(n3431), .ZN(n3430) );
  AOI22_X1 U22012 ( .A1(n12108), .A2(n16862), .B1(n16908), .B2(n4436), .ZN(
        n12215) );
  INV_X2 U22017 ( .I(n3436), .ZN(n25247) );
  XOR2_X1 U22020 ( .A1(n3438), .A2(n38870), .Z(n39750) );
  XOR2_X1 U22023 ( .A1(n1760), .A2(n953), .Z(n3440) );
  NAND2_X2 U22026 ( .A1(n35656), .A2(n63773), .ZN(n35645) );
  INV_X4 U22027 ( .I(n35651), .ZN(n35656) );
  NAND2_X2 U22028 ( .A1(n19701), .A2(n13280), .ZN(n28681) );
  NAND3_X2 U22031 ( .A1(n3453), .A2(n3451), .A3(n3450), .ZN(n46269) );
  NOR2_X1 U22032 ( .A1(n60949), .A2(n3459), .ZN(n12358) );
  NAND2_X2 U22033 ( .A1(n58250), .A2(n37224), .ZN(n3460) );
  NAND2_X2 U22036 ( .A1(n13798), .A2(n25924), .ZN(n42387) );
  NOR2_X2 U22037 ( .A1(n27292), .A2(n25202), .ZN(n7371) );
  XOR2_X1 U22038 ( .A1(n26807), .A2(n26808), .Z(n3470) );
  OAI22_X1 U22039 ( .A1(n29121), .A2(n29128), .B1(n29118), .B2(n3473), .ZN(
        n27409) );
  INV_X1 U22042 ( .I(n10776), .ZN(n44421) );
  XOR2_X1 U22043 ( .A1(n45128), .A2(n46653), .Z(n3475) );
  XOR2_X1 U22044 ( .A1(n3476), .A2(n60458), .Z(n46653) );
  XOR2_X1 U22048 ( .A1(n32060), .A2(n32164), .Z(n32757) );
  XOR2_X1 U22049 ( .A1(n31322), .A2(n32335), .Z(n32164) );
  NOR2_X2 U22050 ( .A1(n31213), .A2(n31212), .ZN(n32335) );
  XOR2_X1 U22052 ( .A1(n33248), .A2(n22978), .Z(n32010) );
  INV_X1 U22054 ( .I(n7564), .ZN(n3482) );
  NAND2_X2 U22055 ( .A1(n10908), .A2(n10739), .ZN(n8113) );
  XOR2_X1 U22057 ( .A1(Ciphertext[144]), .A2(Key[37]), .Z(n12049) );
  NAND2_X2 U22061 ( .A1(n42452), .A2(n21920), .ZN(n41805) );
  XOR2_X1 U22066 ( .A1(n3715), .A2(n22698), .Z(n15371) );
  XOR2_X1 U22067 ( .A1(n4563), .A2(n3499), .Z(n39395) );
  XOR2_X1 U22071 ( .A1(n16519), .A2(n1881), .Z(n3500) );
  NAND2_X1 U22072 ( .A1(n9801), .A2(n62435), .ZN(n24685) );
  NOR2_X1 U22073 ( .A1(n40278), .A2(n9801), .ZN(n5541) );
  XOR2_X1 U22074 ( .A1(n8599), .A2(n46271), .Z(n3777) );
  NAND2_X1 U22076 ( .A1(n3505), .A2(n64566), .ZN(n40331) );
  NAND2_X1 U22077 ( .A1(n40267), .A2(n3505), .ZN(n40268) );
  NAND2_X1 U22078 ( .A1(n40328), .A2(n3505), .ZN(n40330) );
  NAND2_X1 U22079 ( .A1(n40329), .A2(n3505), .ZN(n18015) );
  XOR2_X1 U22086 ( .A1(n3776), .A2(n3775), .Z(n8525) );
  NAND2_X1 U22088 ( .A1(n36422), .A2(n1227), .ZN(n36176) );
  NAND2_X2 U22089 ( .A1(n21808), .A2(n21806), .ZN(n36178) );
  NAND3_X2 U22090 ( .A1(n3512), .A2(n3515), .A3(n3511), .ZN(n33721) );
  INV_X2 U22092 ( .I(n3516), .ZN(n3580) );
  XNOR2_X1 U22093 ( .A1(Ciphertext[76]), .A2(Key[137]), .ZN(n3516) );
  XOR2_X1 U22094 ( .A1(n3517), .A2(n44389), .Z(n6715) );
  XOR2_X1 U22096 ( .A1(n16376), .A2(n51522), .Z(n3518) );
  XOR2_X1 U22100 ( .A1(n3522), .A2(n3521), .Z(n3520) );
  XOR2_X1 U22101 ( .A1(n8526), .A2(n13475), .Z(n3521) );
  XOR2_X1 U22109 ( .A1(Ciphertext[75]), .A2(Key[34]), .Z(n15092) );
  XOR2_X1 U22114 ( .A1(n6889), .A2(n37865), .Z(n3527) );
  XOR2_X1 U22116 ( .A1(n38214), .A2(n38218), .Z(n3530) );
  XOR2_X1 U22118 ( .A1(n18268), .A2(n38219), .Z(n3532) );
  XOR2_X1 U22120 ( .A1(n25856), .A2(n3533), .Z(n24517) );
  AOI22_X2 U22122 ( .A1(n29066), .A2(n29065), .B1(n22325), .B2(n29067), .ZN(
        n18356) );
  XOR2_X1 U22129 ( .A1(n32615), .A2(n5489), .Z(n31637) );
  NAND2_X2 U22130 ( .A1(n52230), .A2(n5614), .ZN(n53126) );
  NAND2_X2 U22133 ( .A1(n3547), .A2(n3550), .ZN(n36256) );
  NOR2_X1 U22137 ( .A1(n3555), .A2(n29129), .ZN(n3553) );
  INV_X2 U22138 ( .I(n3556), .ZN(n25721) );
  NAND2_X1 U22142 ( .A1(n23478), .A2(n1253), .ZN(n29412) );
  NAND2_X1 U22143 ( .A1(n3560), .A2(n64534), .ZN(n7207) );
  NAND2_X1 U22148 ( .A1(n35509), .A2(n3561), .ZN(n32907) );
  NAND3_X1 U22149 ( .A1(n11780), .A2(n35507), .A3(n3561), .ZN(n11779) );
  AOI21_X1 U22151 ( .A1(n14753), .A2(n32895), .B(n3561), .ZN(n32905) );
  AOI21_X1 U22152 ( .A1(n35504), .A2(n3561), .B(n36921), .ZN(n34928) );
  NOR2_X1 U22153 ( .A1(n47615), .A2(n3562), .ZN(n7286) );
  AOI21_X1 U22154 ( .A1(n45985), .A2(n3562), .B(n47615), .ZN(n45573) );
  NAND2_X1 U22155 ( .A1(n47241), .A2(n3562), .ZN(n8650) );
  OAI22_X1 U22156 ( .A1(n45578), .A2(n47618), .B1(n45579), .B2(n3562), .ZN(
        n45580) );
  NAND2_X2 U22157 ( .A1(n45988), .A2(n15806), .ZN(n3562) );
  INV_X2 U22158 ( .I(n42262), .ZN(n5581) );
  XOR2_X1 U22166 ( .A1(n25856), .A2(n13771), .Z(n18391) );
  XOR2_X1 U22167 ( .A1(n59163), .A2(n844), .Z(n13291) );
  XOR2_X1 U22171 ( .A1(n3574), .A2(n3571), .Z(n3570) );
  XOR2_X1 U22172 ( .A1(n3573), .A2(n3572), .Z(n3571) );
  XOR2_X1 U22173 ( .A1(n13883), .A2(n44963), .Z(n3572) );
  XOR2_X1 U22175 ( .A1(n21253), .A2(n26011), .Z(n3574) );
  INV_X2 U22180 ( .I(n3579), .ZN(n25849) );
  NAND2_X2 U22181 ( .A1(n30376), .A2(n847), .ZN(n31144) );
  INV_X2 U22182 ( .I(n14767), .ZN(n30376) );
  NAND2_X2 U22183 ( .A1(n5769), .A2(n27647), .ZN(n14767) );
  XOR2_X1 U22186 ( .A1(n5897), .A2(n59811), .Z(n45110) );
  XNOR2_X1 U22187 ( .A1(n16909), .A2(n25432), .ZN(n5897) );
  NAND2_X1 U22194 ( .A1(n3591), .A2(n28616), .ZN(n27642) );
  NAND2_X1 U22195 ( .A1(n10085), .A2(n3591), .ZN(n27650) );
  NOR2_X1 U22196 ( .A1(n23487), .A2(n3591), .ZN(n28437) );
  NOR2_X1 U22197 ( .A1(n65039), .A2(n3591), .ZN(n26793) );
  AOI21_X1 U22198 ( .A1(n28612), .A2(n23033), .B(n3591), .ZN(n13014) );
  NAND2_X2 U22199 ( .A1(n23649), .A2(n23814), .ZN(n3591) );
  XOR2_X1 U22202 ( .A1(n62987), .A2(n58945), .Z(n50976) );
  NAND2_X2 U22204 ( .A1(n3596), .A2(n5481), .ZN(n49842) );
  NAND3_X1 U22205 ( .A1(n10405), .A2(n47852), .A3(n3597), .ZN(n43833) );
  XOR2_X1 U22207 ( .A1(n3605), .A2(n928), .Z(n3600) );
  INV_X2 U22209 ( .I(n3602), .ZN(n25204) );
  XOR2_X1 U22211 ( .A1(n3604), .A2(n21826), .Z(n3603) );
  XOR2_X1 U22212 ( .A1(n3499), .A2(n38837), .Z(n3605) );
  NAND2_X2 U22216 ( .A1(n62314), .A2(n42807), .ZN(n3606) );
  NOR2_X2 U22217 ( .A1(n24003), .A2(n52131), .ZN(n17708) );
  NAND2_X2 U22218 ( .A1(n1840), .A2(n23502), .ZN(n6178) );
  XOR2_X1 U22223 ( .A1(n32036), .A2(n18211), .Z(n25307) );
  NOR2_X1 U22228 ( .A1(n3613), .A2(n56350), .ZN(n56339) );
  OAI21_X1 U22229 ( .A1(n3613), .A2(n1591), .B(n56296), .ZN(n56283) );
  AOI22_X1 U22230 ( .A1(n56320), .A2(n3613), .B1(n11427), .B2(n22430), .ZN(
        n11918) );
  NAND2_X2 U22231 ( .A1(n3616), .A2(n24944), .ZN(n11521) );
  NAND2_X1 U22234 ( .A1(n5672), .A2(n3616), .ZN(n5670) );
  INV_X4 U22235 ( .I(n8122), .ZN(n3616) );
  XOR2_X1 U22236 ( .A1(Ciphertext[79]), .A2(Key[62]), .Z(n7322) );
  XOR2_X1 U22237 ( .A1(n37488), .A2(n23518), .Z(n24752) );
  XOR2_X1 U22238 ( .A1(n11234), .A2(n23518), .Z(n18784) );
  NAND3_X2 U22239 ( .A1(n41000), .A2(n40999), .A3(n19351), .ZN(n42175) );
  NOR2_X2 U22240 ( .A1(n3619), .A2(n3618), .ZN(n6764) );
  INV_X1 U22242 ( .I(n3620), .ZN(n21771) );
  AOI21_X1 U22245 ( .A1(n36767), .A2(n3620), .B(n36766), .ZN(n9597) );
  OAI21_X1 U22246 ( .A1(n3620), .A2(n36771), .B(n36770), .ZN(n9596) );
  XOR2_X1 U22248 ( .A1(n12005), .A2(n51924), .Z(n3621) );
  AOI21_X1 U22251 ( .A1(n48374), .A2(n3596), .B(n3772), .ZN(n45613) );
  NAND3_X1 U22252 ( .A1(n49851), .A2(n22756), .A3(n62927), .ZN(n49852) );
  XOR2_X1 U22253 ( .A1(n3625), .A2(n51881), .Z(n38901) );
  XOR2_X1 U22254 ( .A1(n3625), .A2(n38091), .Z(n38092) );
  OR2_X1 U22257 ( .A1(n3626), .A2(n24060), .Z(n17931) );
  NOR2_X2 U22259 ( .A1(n41158), .A2(n41160), .ZN(n39066) );
  NAND2_X2 U22260 ( .A1(n41164), .A2(n23634), .ZN(n41166) );
  OAI22_X1 U22267 ( .A1(n47299), .A2(n47301), .B1(n46025), .B2(n3641), .ZN(
        n45937) );
  NOR2_X1 U22268 ( .A1(n3641), .A2(n47302), .ZN(n7234) );
  NOR2_X1 U22281 ( .A1(n9566), .A2(n3653), .ZN(n9565) );
  NAND2_X1 U22285 ( .A1(n2433), .A2(n3654), .ZN(n25473) );
  XOR2_X1 U22290 ( .A1(n21724), .A2(n44022), .Z(n44084) );
  NOR2_X2 U22292 ( .A1(n22131), .A2(n22130), .ZN(n44022) );
  NOR2_X2 U22296 ( .A1(n7077), .A2(n3662), .ZN(n49637) );
  OAI21_X1 U22298 ( .A1(n47604), .A2(n47827), .B(n3663), .ZN(n47606) );
  NAND2_X2 U22301 ( .A1(n47604), .A2(n14199), .ZN(n3663) );
  INV_X1 U22304 ( .I(n3665), .ZN(n8354) );
  XOR2_X1 U22305 ( .A1(n3665), .A2(n18809), .Z(n9930) );
  NAND3_X1 U22307 ( .A1(n20984), .A2(n41453), .A3(n3667), .ZN(n38841) );
  XOR2_X1 U22311 ( .A1(n24258), .A2(n31063), .Z(n31019) );
  OAI21_X1 U22316 ( .A1(n3966), .A2(n3962), .B(n1574), .ZN(n3671) );
  OR2_X1 U22317 ( .A1(n3962), .A2(n1574), .Z(n3672) );
  NAND2_X2 U22318 ( .A1(n61745), .A2(n15784), .ZN(n42543) );
  NOR2_X1 U22319 ( .A1(n3675), .A2(n15784), .ZN(n41577) );
  XOR2_X1 U22325 ( .A1(n51917), .A2(n51385), .Z(n51589) );
  XOR2_X1 U22331 ( .A1(n3690), .A2(n3866), .Z(n4915) );
  XOR2_X1 U22332 ( .A1(n6816), .A2(n3690), .Z(n6106) );
  NOR2_X1 U22336 ( .A1(n13819), .A2(n49195), .ZN(n3695) );
  CLKBUF_X4 U22337 ( .I(n41287), .Z(n3696) );
  NOR2_X2 U22338 ( .A1(n43657), .A2(n41287), .ZN(n11635) );
  AOI21_X1 U22341 ( .A1(n1586), .A2(n271), .B(n5476), .ZN(n4989) );
  OAI21_X1 U22343 ( .A1(n29276), .A2(n29277), .B(n3706), .ZN(n29279) );
  NOR2_X1 U22344 ( .A1(n3708), .A2(n62768), .ZN(n54095) );
  OAI21_X1 U22346 ( .A1(n62648), .A2(n3708), .B(n54658), .ZN(n5057) );
  NAND2_X2 U22355 ( .A1(n3716), .A2(n47309), .ZN(n47313) );
  NAND2_X2 U22361 ( .A1(n14230), .A2(n1208), .ZN(n29992) );
  NAND2_X1 U22362 ( .A1(n30319), .A2(n1208), .ZN(n29995) );
  NAND2_X2 U22364 ( .A1(n29820), .A2(n29993), .ZN(n16026) );
  XOR2_X1 U22367 ( .A1(n14230), .A2(n1208), .Z(n4103) );
  XOR2_X1 U22371 ( .A1(n3724), .A2(n44036), .Z(n9257) );
  INV_X2 U22373 ( .I(n57061), .ZN(n57063) );
  NAND2_X2 U22375 ( .A1(n39509), .A2(n1745), .ZN(n8394) );
  INV_X1 U22377 ( .I(n3725), .ZN(n39508) );
  NOR2_X2 U22378 ( .A1(n3302), .A2(n18742), .ZN(n8373) );
  INV_X1 U22381 ( .I(n3733), .ZN(n8953) );
  NAND3_X1 U22382 ( .A1(n47886), .A2(n3732), .A3(n47362), .ZN(n47363) );
  OAI22_X1 U22388 ( .A1(n49102), .A2(n60428), .B1(n49101), .B2(n61362), .ZN(
        n49103) );
  NAND2_X2 U22389 ( .A1(n7587), .A2(n10045), .ZN(n3734) );
  NOR2_X2 U22390 ( .A1(n24455), .A2(n55668), .ZN(n4830) );
  INV_X2 U22391 ( .I(n32919), .ZN(n34962) );
  INV_X2 U22392 ( .I(n3735), .ZN(n34972) );
  INV_X2 U22395 ( .I(n63015), .ZN(n4897) );
  NAND2_X2 U22397 ( .A1(n3739), .A2(n47333), .ZN(n49923) );
  INV_X1 U22400 ( .I(n5897), .ZN(n15266) );
  NAND3_X1 U22402 ( .A1(n22745), .A2(n58644), .A3(n9979), .ZN(n30633) );
  INV_X1 U22403 ( .I(n30748), .ZN(n9979) );
  XOR2_X1 U22405 ( .A1(n51804), .A2(n65016), .Z(n50530) );
  XOR2_X1 U22406 ( .A1(n51804), .A2(n51803), .Z(n17370) );
  XOR2_X1 U22407 ( .A1(n3741), .A2(n51123), .Z(n51124) );
  XOR2_X1 U22408 ( .A1(n3741), .A2(n24758), .Z(n51368) );
  XOR2_X1 U22409 ( .A1(n59787), .A2(n51374), .Z(n8426) );
  XOR2_X1 U22410 ( .A1(n59787), .A2(n50317), .Z(n50318) );
  XOR2_X1 U22411 ( .A1(n22650), .A2(n64013), .Z(n44584) );
  XOR2_X1 U22412 ( .A1(n64013), .A2(n23267), .Z(n44464) );
  XOR2_X1 U22413 ( .A1(n8673), .A2(n64013), .Z(n13228) );
  NOR3_X2 U22415 ( .A1(n25571), .A2(n21010), .A3(n60659), .ZN(n7861) );
  XOR2_X1 U22416 ( .A1(n3751), .A2(n39342), .Z(n3755) );
  XOR2_X1 U22418 ( .A1(n5522), .A2(n1758), .Z(n3754) );
  XOR2_X1 U22419 ( .A1(Ciphertext[131]), .A2(Key[42]), .Z(n3773) );
  XOR2_X1 U22422 ( .A1(n3757), .A2(n8422), .Z(n21899) );
  INV_X2 U22424 ( .I(n21899), .ZN(n24083) );
  XOR2_X1 U22425 ( .A1(n19527), .A2(n16324), .Z(n13046) );
  NAND2_X2 U22428 ( .A1(n14217), .A2(n3761), .ZN(n19721) );
  NAND2_X2 U22429 ( .A1(n30746), .A2(n3761), .ZN(n14641) );
  NAND2_X1 U22435 ( .A1(n54089), .A2(n3769), .ZN(n54090) );
  NAND3_X1 U22436 ( .A1(n51702), .A2(n54595), .A3(n3769), .ZN(n51704) );
  NOR2_X2 U22438 ( .A1(n25519), .A2(n54323), .ZN(n54325) );
  AOI22_X1 U22439 ( .A1(n12198), .A2(n3770), .B1(n59629), .B2(n47611), .ZN(
        n12197) );
  NAND2_X1 U22440 ( .A1(n49843), .A2(n3772), .ZN(n49454) );
  INV_X2 U22443 ( .I(n3773), .ZN(n29690) );
  NAND2_X2 U22444 ( .A1(n29695), .A2(n25341), .ZN(n28651) );
  XOR2_X1 U22446 ( .A1(n20448), .A2(n8596), .Z(n3775) );
  XOR2_X1 U22448 ( .A1(n21316), .A2(n23006), .Z(n20448) );
  NAND2_X1 U22452 ( .A1(n14776), .A2(n3780), .ZN(n21443) );
  NOR2_X1 U22453 ( .A1(n57156), .A2(n58277), .ZN(n3780) );
  INV_X1 U22455 ( .I(n14776), .ZN(n3781) );
  NAND3_X1 U22456 ( .A1(n22182), .A2(n11198), .A3(n41568), .ZN(n3782) );
  NAND2_X2 U22463 ( .A1(n43381), .A2(n43373), .ZN(n42756) );
  INV_X1 U22467 ( .I(n3793), .ZN(n27945) );
  XOR2_X1 U22469 ( .A1(n31632), .A2(n3799), .Z(n14215) );
  XOR2_X1 U22470 ( .A1(n17182), .A2(n3800), .Z(n3799) );
  XOR2_X1 U22471 ( .A1(n31675), .A2(n841), .Z(n3800) );
  NAND2_X2 U22472 ( .A1(n6444), .A2(n19070), .ZN(n31675) );
  NAND2_X2 U22475 ( .A1(n10013), .A2(n16738), .ZN(n24258) );
  NAND2_X2 U22476 ( .A1(n42407), .A2(n19241), .ZN(n42082) );
  INV_X1 U22482 ( .I(n3809), .ZN(n36373) );
  NAND3_X1 U22483 ( .A1(n36379), .A2(n3809), .A3(n64181), .ZN(n32979) );
  NAND2_X1 U22484 ( .A1(n36090), .A2(n3809), .ZN(n35535) );
  NAND2_X1 U22491 ( .A1(n18397), .A2(n29980), .ZN(n3817) );
  NAND2_X2 U22495 ( .A1(n26742), .A2(n29154), .ZN(n6522) );
  XOR2_X1 U22497 ( .A1(n3830), .A2(n3829), .Z(n16756) );
  XOR2_X1 U22498 ( .A1(n24580), .A2(n19769), .Z(n3829) );
  XOR2_X1 U22500 ( .A1(n46580), .A2(n19767), .Z(n3831) );
  XOR2_X1 U22503 ( .A1(n44362), .A2(n5989), .Z(n24580) );
  XOR2_X1 U22505 ( .A1(n46551), .A2(n46550), .Z(n46580) );
  NAND2_X2 U22512 ( .A1(n7854), .A2(n26226), .ZN(n12968) );
  XOR2_X1 U22517 ( .A1(n60654), .A2(n32356), .Z(n3840) );
  XOR2_X1 U22520 ( .A1(n3842), .A2(n52497), .Z(n21412) );
  XOR2_X1 U22523 ( .A1(n3843), .A2(n13739), .Z(n17765) );
  OAI21_X1 U22529 ( .A1(n46098), .A2(n62220), .B(n48600), .ZN(n46099) );
  XOR2_X1 U22531 ( .A1(n25149), .A2(n3863), .Z(n9878) );
  XNOR2_X1 U22532 ( .A1(n50648), .A2(n51621), .ZN(n25149) );
  NAND2_X2 U22536 ( .A1(n3862), .A2(n3861), .ZN(n51621) );
  NOR2_X2 U22538 ( .A1(n23716), .A2(n28221), .ZN(n10404) );
  XOR2_X1 U22541 ( .A1(Ciphertext[61]), .A2(Key[128]), .Z(n4506) );
  XOR2_X1 U22542 ( .A1(n58750), .A2(n45086), .Z(n3875) );
  XOR2_X1 U22550 ( .A1(n33053), .A2(n30912), .Z(n3881) );
  INV_X2 U22554 ( .I(n8989), .ZN(n9255) );
  INV_X2 U22562 ( .I(n3887), .ZN(n53845) );
  INV_X2 U22568 ( .I(n3890), .ZN(n11443) );
  NAND2_X1 U22575 ( .A1(n3895), .A2(n53824), .ZN(n53045) );
  NOR2_X2 U22577 ( .A1(n11092), .A2(n23140), .ZN(n30331) );
  AOI21_X1 U22580 ( .A1(n63850), .A2(n27996), .B(n3904), .ZN(n5415) );
  XNOR2_X1 U22581 ( .A1(n19155), .A2(n44991), .ZN(n46354) );
  NAND3_X2 U22583 ( .A1(n40371), .A2(n40372), .A3(n40370), .ZN(n3905) );
  XOR2_X1 U22585 ( .A1(n44386), .A2(n7365), .Z(n3913) );
  NAND2_X2 U22587 ( .A1(n11037), .A2(n21320), .ZN(n17379) );
  INV_X1 U22590 ( .I(n10363), .ZN(n33171) );
  AOI21_X1 U22591 ( .A1(n3908), .A2(n24949), .B(n29007), .ZN(n27632) );
  INV_X2 U22592 ( .I(n3911), .ZN(n29106) );
  NOR2_X1 U22593 ( .A1(n23716), .A2(n3911), .ZN(n3910) );
  NOR2_X2 U22594 ( .A1(n27374), .A2(n435), .ZN(n3911) );
  INV_X2 U22595 ( .I(n32283), .ZN(n32710) );
  XOR2_X1 U22599 ( .A1(n23668), .A2(n9079), .Z(n3914) );
  OR2_X1 U22602 ( .A1(n4908), .A2(n48067), .Z(n3923) );
  XOR2_X1 U22606 ( .A1(n29204), .A2(n3928), .Z(n3927) );
  INV_X1 U22607 ( .I(n33880), .ZN(n3928) );
  XOR2_X1 U22608 ( .A1(n26178), .A2(n3930), .Z(n3929) );
  XOR2_X1 U22609 ( .A1(n11484), .A2(n11483), .Z(n3930) );
  NOR2_X2 U22611 ( .A1(n27097), .A2(n3932), .ZN(n28034) );
  XOR2_X1 U22612 ( .A1(Ciphertext[42]), .A2(Key[91]), .Z(n6589) );
  NAND2_X1 U22614 ( .A1(n28984), .A2(n25898), .ZN(n3933) );
  OR2_X2 U22616 ( .A1(n3935), .A2(n24589), .Z(n35003) );
  NAND2_X1 U22618 ( .A1(n3939), .A2(n35774), .ZN(n35776) );
  NOR2_X2 U22619 ( .A1(n35775), .A2(n3939), .ZN(n34423) );
  OAI21_X1 U22622 ( .A1(n33924), .A2(n3939), .B(n3938), .ZN(n32139) );
  NAND2_X1 U22623 ( .A1(n35770), .A2(n3939), .ZN(n3938) );
  NAND2_X1 U22624 ( .A1(n5874), .A2(n3940), .ZN(n34428) );
  NAND2_X1 U22625 ( .A1(n1806), .A2(n10769), .ZN(n3940) );
  XOR2_X1 U22626 ( .A1(n3941), .A2(n45284), .Z(n18695) );
  XOR2_X1 U22628 ( .A1(n23783), .A2(n3941), .Z(n19656) );
  NAND2_X1 U22630 ( .A1(n45781), .A2(n3942), .ZN(n44698) );
  NAND2_X1 U22631 ( .A1(n13655), .A2(n61166), .ZN(n45537) );
  NAND2_X1 U22633 ( .A1(n44699), .A2(n61166), .ZN(n44403) );
  NAND2_X2 U22638 ( .A1(n1402), .A2(n15731), .ZN(n3946) );
  NAND2_X2 U22639 ( .A1(n3946), .A2(n22776), .ZN(n41936) );
  NAND2_X1 U22640 ( .A1(n40818), .A2(n3946), .ZN(n40819) );
  XOR2_X1 U22641 ( .A1(n51509), .A2(n20723), .Z(n19711) );
  XOR2_X1 U22647 ( .A1(n15938), .A2(n24248), .Z(n3950) );
  XOR2_X1 U22648 ( .A1(n4667), .A2(n1899), .Z(n15938) );
  NAND3_X2 U22649 ( .A1(n3954), .A2(n3952), .A3(n3951), .ZN(n44156) );
  NOR3_X2 U22650 ( .A1(n13832), .A2(n42749), .A3(n42748), .ZN(n3951) );
  NAND2_X1 U22652 ( .A1(n65147), .A2(n60843), .ZN(n3953) );
  NAND2_X1 U22654 ( .A1(n43052), .A2(n43874), .ZN(n3958) );
  NOR2_X1 U22655 ( .A1(n48419), .A2(n201), .ZN(n48420) );
  OAI22_X1 U22656 ( .A1(n48415), .A2(n12595), .B1(n201), .B2(n48416), .ZN(
        n12838) );
  XOR2_X1 U22657 ( .A1(n32332), .A2(n3959), .Z(n11633) );
  XOR2_X1 U22658 ( .A1(n32268), .A2(n1824), .Z(n3959) );
  XOR2_X1 U22659 ( .A1(n3960), .A2(n32655), .Z(n32332) );
  XOR2_X1 U22660 ( .A1(n31686), .A2(n32754), .Z(n3960) );
  NOR2_X2 U22668 ( .A1(n48069), .A2(n48070), .ZN(n49053) );
  NAND2_X1 U22678 ( .A1(n21550), .A2(n3979), .ZN(n26099) );
  NAND2_X1 U22679 ( .A1(n47978), .A2(n3979), .ZN(n4300) );
  AOI22_X1 U22681 ( .A1(n3980), .A2(n15784), .B1(n41577), .B2(n42545), .ZN(
        n13102) );
  OR2_X1 U22683 ( .A1(n31042), .A2(n31041), .Z(n3986) );
  AOI21_X1 U22686 ( .A1(n36532), .A2(n36548), .B(n20530), .ZN(n4009) );
  NAND3_X2 U22688 ( .A1(n46090), .A2(n47068), .A3(n4015), .ZN(n4014) );
  INV_X1 U22694 ( .I(n6943), .ZN(n20484) );
  OAI22_X1 U22695 ( .A1(n53242), .A2(n53238), .B1(n61730), .B2(n61572), .ZN(
        n4023) );
  INV_X1 U22698 ( .I(n61730), .ZN(n4025) );
  INV_X1 U22703 ( .I(n21572), .ZN(n4029) );
  NOR2_X1 U22709 ( .A1(n12855), .A2(n4033), .ZN(n53053) );
  INV_X1 U22712 ( .I(n32527), .ZN(n4034) );
  NAND2_X1 U22713 ( .A1(n36565), .A2(n4035), .ZN(n19559) );
  NOR2_X2 U22716 ( .A1(n25755), .A2(n22742), .ZN(n4037) );
  INV_X2 U22717 ( .I(n4038), .ZN(n5536) );
  XOR2_X1 U22718 ( .A1(n12379), .A2(n20998), .Z(n50633) );
  NOR2_X2 U22721 ( .A1(n37452), .A2(n37453), .ZN(n37600) );
  AOI22_X1 U22723 ( .A1(n29683), .A2(n28182), .B1(n17274), .B2(n28639), .ZN(
        n4043) );
  NOR2_X1 U22724 ( .A1(n42916), .A2(n4077), .ZN(n42921) );
  NAND2_X1 U22725 ( .A1(n9191), .A2(n57808), .ZN(n41714) );
  NOR2_X1 U22726 ( .A1(n9191), .A2(n57808), .ZN(n42111) );
  INV_X1 U22727 ( .I(n4046), .ZN(n34804) );
  NAND3_X1 U22728 ( .A1(n4046), .A2(n1418), .A3(n59147), .ZN(n21742) );
  NAND2_X2 U22731 ( .A1(n4048), .A2(n4047), .ZN(n7971) );
  OAI21_X1 U22740 ( .A1(n29509), .A2(n4270), .B(n29508), .ZN(n4051) );
  XOR2_X1 U22742 ( .A1(n37821), .A2(n38106), .Z(n4052) );
  NAND2_X2 U22743 ( .A1(n25918), .A2(n25915), .ZN(n38106) );
  INV_X2 U22744 ( .I(n4054), .ZN(n55950) );
  XOR2_X1 U22747 ( .A1(n25106), .A2(n17781), .Z(n18156) );
  INV_X1 U22757 ( .I(n24329), .ZN(n52403) );
  XOR2_X1 U22758 ( .A1(n51028), .A2(n50107), .Z(n21970) );
  XOR2_X1 U22759 ( .A1(n24329), .A2(n4064), .Z(n50107) );
  XOR2_X1 U22764 ( .A1(n21650), .A2(n18648), .Z(n4068) );
  XOR2_X1 U22767 ( .A1(n38360), .A2(n1759), .Z(n4072) );
  XOR2_X1 U22769 ( .A1(n52403), .A2(n52402), .Z(n52405) );
  XOR2_X1 U22770 ( .A1(n52403), .A2(n50919), .Z(n50920) );
  XOR2_X1 U22771 ( .A1(n52403), .A2(n51725), .Z(n51726) );
  XOR2_X1 U22772 ( .A1(n52403), .A2(n50321), .Z(n50322) );
  NAND3_X2 U22774 ( .A1(n3128), .A2(n35508), .A3(n24198), .ZN(n18509) );
  NAND2_X2 U22775 ( .A1(n5473), .A2(n5475), .ZN(n42104) );
  XOR2_X1 U22778 ( .A1(n4079), .A2(n9419), .Z(n22594) );
  XOR2_X1 U22779 ( .A1(n8862), .A2(n1673), .Z(n4080) );
  NAND2_X1 U22780 ( .A1(n1566), .A2(n28648), .ZN(n16185) );
  NAND2_X1 U22781 ( .A1(n28188), .A2(n4081), .ZN(n18823) );
  AOI22_X1 U22782 ( .A1(n11352), .A2(n4081), .B1(n28188), .B2(n29697), .ZN(
        n14924) );
  NAND2_X2 U22783 ( .A1(n28187), .A2(n11655), .ZN(n4081) );
  NOR2_X2 U22784 ( .A1(n23918), .A2(n31147), .ZN(n22627) );
  XOR2_X1 U22786 ( .A1(n14027), .A2(n5626), .Z(n4085) );
  NAND2_X2 U22787 ( .A1(n4086), .A2(n46033), .ZN(n46872) );
  INV_X4 U22790 ( .I(n25092), .ZN(n4086) );
  NAND2_X1 U22794 ( .A1(n1072), .A2(n4090), .ZN(n14569) );
  NAND2_X1 U22799 ( .A1(n39926), .A2(n21207), .ZN(n4096) );
  NAND2_X2 U22801 ( .A1(n34119), .A2(n15783), .ZN(n4097) );
  XOR2_X1 U22806 ( .A1(n4105), .A2(n16475), .Z(n19821) );
  XOR2_X1 U22807 ( .A1(n4105), .A2(n51407), .Z(n23174) );
  XOR2_X1 U22808 ( .A1(n4105), .A2(n54917), .Z(n37552) );
  AOI22_X2 U22811 ( .A1(n43338), .A2(n42587), .B1(n4106), .B2(n42155), .ZN(
        n42589) );
  NAND2_X2 U22812 ( .A1(n18882), .A2(n60163), .ZN(n4109) );
  OAI21_X1 U22813 ( .A1(n4109), .A2(n50240), .B(n14353), .ZN(n19618) );
  XOR2_X1 U22814 ( .A1(n46691), .A2(n4111), .Z(n45044) );
  XOR2_X1 U22815 ( .A1(n4111), .A2(n45114), .Z(n45116) );
  INV_X1 U22820 ( .I(n29295), .ZN(n5259) );
  NAND2_X2 U22821 ( .A1(n1445), .A2(n22410), .ZN(n22144) );
  NAND2_X2 U22824 ( .A1(n4117), .A2(n4116), .ZN(n52808) );
  OAI22_X1 U22831 ( .A1(n27962), .A2(n60993), .B1(n22043), .B2(n64374), .ZN(
        n27403) );
  OAI21_X1 U22832 ( .A1(n28275), .A2(n28274), .B(n64374), .ZN(n28276) );
  XOR2_X1 U22836 ( .A1(n4130), .A2(n5434), .Z(n4129) );
  XOR2_X1 U22837 ( .A1(n5437), .A2(n25887), .Z(n4130) );
  NOR2_X2 U22838 ( .A1(n4135), .A2(n4131), .ZN(n11818) );
  OAI21_X1 U22839 ( .A1(n19343), .A2(n20856), .B(n18418), .ZN(n4133) );
  NAND3_X2 U22840 ( .A1(n4141), .A2(n4138), .A3(n4136), .ZN(n4135) );
  XOR2_X1 U22842 ( .A1(n8214), .A2(n18584), .Z(n4142) );
  MUX2_X1 U22843 ( .I0(n10456), .I1(n49388), .S(n49382), .Z(n44011) );
  XOR2_X1 U22848 ( .A1(n7102), .A2(n4145), .Z(n4144) );
  XOR2_X1 U22849 ( .A1(n4148), .A2(n4147), .Z(n4146) );
  NAND3_X1 U22851 ( .A1(n42129), .A2(n21376), .A3(n42667), .ZN(n4149) );
  XOR2_X1 U22854 ( .A1(n23878), .A2(n61178), .Z(n50600) );
  INV_X2 U22856 ( .I(n19765), .ZN(n34926) );
  NAND2_X1 U22857 ( .A1(n20752), .A2(n4336), .ZN(n54921) );
  INV_X1 U22858 ( .I(n4154), .ZN(n54384) );
  INV_X1 U22859 ( .I(n4153), .ZN(n24193) );
  OAI21_X1 U22860 ( .A1(n4154), .A2(n1586), .B(n54410), .ZN(n4153) );
  XOR2_X1 U22864 ( .A1(n8473), .A2(n51144), .Z(n5272) );
  XOR2_X1 U22865 ( .A1(n4157), .A2(n14640), .Z(n7634) );
  XOR2_X1 U22866 ( .A1(n4158), .A2(n23267), .Z(n4157) );
  XOR2_X1 U22867 ( .A1(n16318), .A2(n4343), .Z(n4158) );
  OR2_X1 U22869 ( .A1(n35666), .A2(n17401), .Z(n4170) );
  NAND2_X1 U22873 ( .A1(n24984), .A2(n64077), .ZN(n24985) );
  NOR2_X1 U22875 ( .A1(n4173), .A2(n49732), .ZN(n4172) );
  OAI21_X1 U22881 ( .A1(n49024), .A2(n62405), .B(n49030), .ZN(n49028) );
  OAI22_X1 U22882 ( .A1(n21017), .A2(n49425), .B1(n63238), .B2(n62405), .ZN(
        n21892) );
  INV_X2 U22885 ( .I(n4175), .ZN(n25339) );
  OAI21_X1 U22891 ( .A1(n46641), .A2(n4176), .B(n47096), .ZN(n46643) );
  XOR2_X1 U22893 ( .A1(n21424), .A2(n15476), .Z(n4178) );
  NAND2_X2 U22897 ( .A1(n41160), .A2(n41161), .ZN(n40645) );
  INV_X2 U22898 ( .I(n53214), .ZN(n57030) );
  MUX2_X1 U22899 ( .I0(n52236), .I1(n4183), .S(n4181), .Z(n4182) );
  NAND2_X2 U22904 ( .A1(n11617), .A2(n13079), .ZN(n21086) );
  NOR2_X2 U22905 ( .A1(n1321), .A2(n26034), .ZN(n12072) );
  OAI21_X1 U22908 ( .A1(n21263), .A2(n4188), .B(n30192), .ZN(n21262) );
  OAI21_X1 U22911 ( .A1(n4191), .A2(n1473), .B(n50373), .ZN(n4190) );
  NOR2_X1 U22912 ( .A1(n4193), .A2(n4192), .ZN(n4191) );
  INV_X1 U22914 ( .I(n8599), .ZN(n46270) );
  NAND2_X2 U22917 ( .A1(n23053), .A2(n1277), .ZN(n4196) );
  OAI22_X1 U22918 ( .A1(n4196), .A2(n1253), .B1(n13572), .B2(n28094), .ZN(
        n13571) );
  OAI21_X1 U22919 ( .A1(n30443), .A2(n30444), .B(n4196), .ZN(n30445) );
  INV_X1 U22923 ( .I(n48148), .ZN(n48549) );
  AOI22_X1 U22927 ( .A1(n21737), .A2(n48953), .B1(n48952), .B2(n49777), .ZN(
        n4202) );
  NAND2_X1 U22928 ( .A1(n21550), .A2(n49777), .ZN(n4207) );
  NAND2_X1 U22929 ( .A1(n21550), .A2(n48949), .ZN(n4208) );
  NOR2_X2 U22930 ( .A1(n49783), .A2(n57735), .ZN(n48949) );
  XOR2_X1 U22931 ( .A1(n4209), .A2(n10283), .Z(n13244) );
  NOR2_X2 U22935 ( .A1(n25470), .A2(n20025), .ZN(n4210) );
  NAND3_X1 U22939 ( .A1(n20666), .A2(n46016), .A3(n25477), .ZN(n19533) );
  XOR2_X1 U22940 ( .A1(n4217), .A2(n13369), .Z(n4215) );
  INV_X2 U22941 ( .I(n4216), .ZN(n11380) );
  XOR2_X1 U22942 ( .A1(n15621), .A2(n4218), .Z(n4217) );
  XOR2_X1 U22943 ( .A1(n4220), .A2(n4219), .Z(n4221) );
  XOR2_X1 U22944 ( .A1(n8629), .A2(n38292), .Z(n4219) );
  XOR2_X1 U22945 ( .A1(n4221), .A2(n18122), .Z(n10519) );
  XOR2_X1 U22946 ( .A1(n11755), .A2(n11751), .Z(n6166) );
  OR3_X1 U22948 ( .A1(n52781), .A2(n53856), .A3(n53025), .Z(n4224) );
  XOR2_X1 U22955 ( .A1(Ciphertext[185]), .A2(Key[36]), .Z(n19340) );
  NOR3_X2 U22958 ( .A1(n24323), .A2(n24322), .A3(n24324), .ZN(n24365) );
  NAND2_X1 U22960 ( .A1(n4231), .A2(n33600), .ZN(n10660) );
  OAI21_X1 U22961 ( .A1(n4231), .A2(n22723), .B(n35691), .ZN(n33306) );
  NOR2_X1 U22962 ( .A1(n35688), .A2(n4231), .ZN(n12121) );
  OAI21_X1 U22963 ( .A1(n35688), .A2(n33338), .B(n4231), .ZN(n4356) );
  XOR2_X1 U22965 ( .A1(n52107), .A2(n1887), .Z(n16119) );
  INV_X2 U22968 ( .I(n54570), .ZN(n22217) );
  INV_X4 U22970 ( .I(n4233), .ZN(n13566) );
  NOR2_X1 U22971 ( .A1(n4233), .A2(n62571), .ZN(n46031) );
  NAND2_X1 U22972 ( .A1(n4233), .A2(n62571), .ZN(n46034) );
  NAND2_X1 U22973 ( .A1(n14300), .A2(n4233), .ZN(n19375) );
  NAND2_X1 U22974 ( .A1(n46858), .A2(n4233), .ZN(n6248) );
  XOR2_X1 U22976 ( .A1(n4234), .A2(n29407), .Z(n52423) );
  XOR2_X1 U22977 ( .A1(n4234), .A2(n10461), .Z(n51554) );
  XOR2_X1 U22980 ( .A1(n32564), .A2(n32562), .Z(n4237) );
  XOR2_X1 U22981 ( .A1(n18837), .A2(n19886), .Z(n32562) );
  OAI21_X1 U22984 ( .A1(n2198), .A2(n22544), .B(n4239), .ZN(n4238) );
  XOR2_X1 U22987 ( .A1(n26028), .A2(n803), .Z(n52332) );
  XOR2_X1 U22988 ( .A1(n26028), .A2(n1290), .Z(n50583) );
  XOR2_X1 U22989 ( .A1(n23697), .A2(n4245), .Z(n21342) );
  XOR2_X1 U22990 ( .A1(n13285), .A2(n4245), .Z(n50729) );
  XOR2_X1 U22991 ( .A1(n5390), .A2(n4245), .Z(n25316) );
  INV_X2 U22992 ( .I(n38338), .ZN(n21207) );
  NAND2_X2 U22993 ( .A1(n52235), .A2(n57030), .ZN(n21582) );
  NOR2_X2 U22994 ( .A1(n12777), .A2(n25936), .ZN(n52235) );
  INV_X2 U22995 ( .I(n14636), .ZN(n25936) );
  NAND2_X2 U22996 ( .A1(n1794), .A2(n35320), .ZN(n4249) );
  AOI21_X2 U22998 ( .A1(n4249), .A2(n35317), .B(n61547), .ZN(n11671) );
  XOR2_X1 U23000 ( .A1(n4252), .A2(n51160), .Z(n13720) );
  XOR2_X1 U23001 ( .A1(n11354), .A2(n19888), .Z(n4252) );
  NAND2_X1 U23002 ( .A1(n11041), .A2(n23974), .ZN(n4255) );
  XOR2_X1 U23004 ( .A1(n4256), .A2(n44316), .Z(n44317) );
  XOR2_X1 U23006 ( .A1(n15095), .A2(n4256), .Z(n9496) );
  NAND2_X1 U23008 ( .A1(n10052), .A2(n31270), .ZN(n31166) );
  NAND2_X1 U23010 ( .A1(n23269), .A2(n4257), .ZN(n31263) );
  NAND2_X2 U23011 ( .A1(n23909), .A2(n29701), .ZN(n10052) );
  INV_X2 U23012 ( .I(n49779), .ZN(n21737) );
  NAND2_X1 U23018 ( .A1(n21839), .A2(n1413), .ZN(n17596) );
  INV_X2 U23019 ( .I(n18053), .ZN(n18313) );
  XOR2_X1 U23026 ( .A1(n4294), .A2(n51526), .Z(n51527) );
  XOR2_X1 U23027 ( .A1(n52172), .A2(n4294), .Z(n13897) );
  XOR2_X1 U23028 ( .A1(n7166), .A2(n4265), .Z(n51198) );
  NAND2_X2 U23031 ( .A1(n13459), .A2(n37415), .ZN(n38989) );
  NAND3_X2 U23032 ( .A1(n13206), .A2(n6138), .A3(n6139), .ZN(n38453) );
  AOI21_X2 U23033 ( .A1(n8150), .A2(n38989), .B(n4269), .ZN(n7418) );
  INV_X2 U23034 ( .I(n25755), .ZN(n24852) );
  NAND2_X2 U23035 ( .A1(n10631), .A2(n26530), .ZN(n25755) );
  XOR2_X1 U23039 ( .A1(n44504), .A2(n44506), .Z(n4273) );
  XOR2_X1 U23040 ( .A1(n44747), .A2(n44318), .Z(n44506) );
  XOR2_X1 U23043 ( .A1(n4280), .A2(n16142), .Z(n4279) );
  XOR2_X1 U23046 ( .A1(n9883), .A2(n31675), .Z(n4281) );
  NAND2_X1 U23048 ( .A1(n4282), .A2(n43714), .ZN(n10302) );
  NAND2_X2 U23049 ( .A1(n4284), .A2(n53229), .ZN(n23862) );
  OAI21_X2 U23050 ( .A1(n44077), .A2(n12835), .B(n4287), .ZN(n16700) );
  NOR2_X2 U23054 ( .A1(n34253), .A2(n493), .ZN(n33737) );
  XOR2_X1 U23056 ( .A1(n4290), .A2(n4292), .Z(n4289) );
  XOR2_X1 U23057 ( .A1(n324), .A2(n4291), .Z(n4290) );
  XOR2_X1 U23058 ( .A1(n38084), .A2(n800), .Z(n4291) );
  XOR2_X1 U23059 ( .A1(n4293), .A2(n38083), .Z(n4292) );
  XOR2_X1 U23060 ( .A1(n23070), .A2(n38999), .Z(n4293) );
  AND2_X1 U23061 ( .A1(n21943), .A2(n61959), .Z(n4302) );
  NAND3_X1 U23063 ( .A1(n13258), .A2(n58233), .A3(n4678), .ZN(n46069) );
  NOR2_X2 U23064 ( .A1(n58313), .A2(n24782), .ZN(n4678) );
  INV_X2 U23065 ( .I(n5662), .ZN(n24782) );
  NOR2_X2 U23066 ( .A1(n35508), .A2(n4304), .ZN(n36924) );
  NAND2_X2 U23067 ( .A1(n53214), .A2(n57017), .ZN(n12573) );
  AOI21_X2 U23077 ( .A1(n4312), .A2(n53362), .B(n53345), .ZN(n12667) );
  OAI21_X1 U23078 ( .A1(n53363), .A2(n53364), .B(n4312), .ZN(n53358) );
  XOR2_X1 U23081 ( .A1(n62873), .A2(n5068), .Z(n45004) );
  NAND2_X2 U23082 ( .A1(n40994), .A2(n10954), .ZN(n5362) );
  INV_X2 U23086 ( .I(n15871), .ZN(n47259) );
  NOR2_X1 U23087 ( .A1(n15871), .A2(n63793), .ZN(n16212) );
  NAND2_X2 U23088 ( .A1(n46897), .A2(n25403), .ZN(n6148) );
  NAND4_X1 U23089 ( .A1(n54753), .A2(n54751), .A3(n54752), .A4(n4316), .ZN(
        n54775) );
  OR2_X1 U23091 ( .A1(n42741), .A2(n4774), .Z(n4318) );
  NAND2_X1 U23092 ( .A1(n14467), .A2(n4319), .ZN(n13334) );
  XOR2_X1 U23095 ( .A1(n13934), .A2(n32563), .Z(n4321) );
  NOR2_X2 U23100 ( .A1(n40344), .A2(n40345), .ZN(n24024) );
  NOR2_X1 U23102 ( .A1(n13645), .A2(n4323), .ZN(n8435) );
  NOR2_X2 U23106 ( .A1(n27188), .A2(n28106), .ZN(n4324) );
  AOI21_X1 U23107 ( .A1(n23383), .A2(n4324), .B(n1572), .ZN(n8022) );
  AOI21_X1 U23108 ( .A1(n62784), .A2(n4324), .B(n12978), .ZN(n23747) );
  NOR2_X1 U23111 ( .A1(n4326), .A2(n1542), .ZN(n31657) );
  NOR3_X1 U23112 ( .A1(n5086), .A2(n5085), .A3(n4326), .ZN(n5084) );
  NAND2_X1 U23116 ( .A1(n54883), .A2(n4152), .ZN(n54884) );
  INV_X4 U23118 ( .I(n4897), .ZN(n20996) );
  XOR2_X1 U23126 ( .A1(n9179), .A2(n17035), .Z(n4340) );
  XOR2_X1 U23127 ( .A1(n16303), .A2(n21094), .Z(n4341) );
  NAND3_X2 U23128 ( .A1(n4342), .A2(n52479), .A3(n5569), .ZN(n55271) );
  NOR2_X1 U23130 ( .A1(n21169), .A2(n55261), .ZN(n4342) );
  XOR2_X1 U23133 ( .A1(n26148), .A2(n4350), .Z(n4349) );
  XOR2_X1 U23134 ( .A1(n17336), .A2(n51293), .Z(n51786) );
  INV_X2 U23135 ( .I(n4351), .ZN(n11355) );
  XOR2_X1 U23136 ( .A1(n4351), .A2(n39436), .Z(n39438) );
  XOR2_X1 U23137 ( .A1(n4351), .A2(n37684), .Z(n37685) );
  NAND2_X2 U23144 ( .A1(n64738), .A2(n24509), .ZN(n21030) );
  NAND2_X1 U23152 ( .A1(n11569), .A2(n21159), .ZN(n11568) );
  NAND2_X2 U23153 ( .A1(n5371), .A2(n1321), .ZN(n28256) );
  XOR2_X1 U23156 ( .A1(n4365), .A2(n773), .Z(n4565) );
  XOR2_X1 U23157 ( .A1(n20535), .A2(n20534), .Z(n4365) );
  OR2_X2 U23158 ( .A1(n9289), .A2(n33005), .Z(n5082) );
  NAND2_X1 U23159 ( .A1(n40806), .A2(n63849), .ZN(n4366) );
  NAND2_X1 U23160 ( .A1(n40807), .A2(n42266), .ZN(n4367) );
  NOR2_X1 U23166 ( .A1(n14656), .A2(n14655), .ZN(n14654) );
  XOR2_X1 U23168 ( .A1(n14249), .A2(n4369), .Z(n16951) );
  AND3_X1 U23170 ( .A1(n19367), .A2(n19832), .A3(n49254), .Z(n7554) );
  XOR2_X1 U23173 ( .A1(n44905), .A2(n16247), .Z(n6252) );
  BUF_X2 U23180 ( .I(n32734), .Z(n24103) );
  AND3_X1 U23182 ( .A1(n29087), .A2(n29088), .A3(n29086), .Z(n19584) );
  INV_X2 U23183 ( .I(n4378), .ZN(n9256) );
  NAND3_X1 U23188 ( .A1(n35022), .A2(n35021), .A3(n35020), .ZN(n16576) );
  OR2_X1 U23189 ( .A1(n18375), .A2(n27936), .Z(n18388) );
  BUF_X4 U23192 ( .I(n23294), .Z(n6606) );
  OR2_X1 U23194 ( .A1(n29862), .A2(n11395), .Z(n28746) );
  AOI22_X1 U23201 ( .A1(n30509), .A2(n25989), .B1(n31269), .B2(n31279), .ZN(
        n4387) );
  XOR2_X1 U23214 ( .A1(Key[111]), .A2(Ciphertext[182]), .Z(n4394) );
  XOR2_X1 U23217 ( .A1(n11501), .A2(n15322), .Z(n51201) );
  OAI21_X1 U23218 ( .A1(n61282), .A2(n2104), .B(n52935), .ZN(n52937) );
  NAND2_X2 U23221 ( .A1(n8029), .A2(n14703), .ZN(n10699) );
  XOR2_X1 U23224 ( .A1(n4398), .A2(n44245), .Z(n7266) );
  INV_X2 U23232 ( .I(n4403), .ZN(n8023) );
  XOR2_X1 U23234 ( .A1(n4404), .A2(n46300), .Z(n46309) );
  XOR2_X1 U23235 ( .A1(n46299), .A2(n46298), .Z(n4404) );
  NAND2_X1 U23237 ( .A1(n48607), .A2(n47546), .ZN(n47543) );
  OAI21_X1 U23238 ( .A1(n27408), .A2(n27409), .B(n27407), .ZN(n9761) );
  NAND3_X1 U23239 ( .A1(n9761), .A2(n22120), .A3(n16199), .ZN(n17215) );
  XOR2_X1 U23241 ( .A1(n32187), .A2(n32188), .Z(n32196) );
  NOR2_X1 U23246 ( .A1(n18460), .A2(n6005), .ZN(n44234) );
  NOR2_X1 U23247 ( .A1(n42090), .A2(n42089), .ZN(n6452) );
  XOR2_X1 U23248 ( .A1(n30980), .A2(n792), .Z(n44100) );
  XOR2_X1 U23249 ( .A1(n37635), .A2(n61034), .Z(n30980) );
  OAI22_X1 U23252 ( .A1(n56339), .A2(n56340), .B1(n56338), .B2(n60353), .ZN(
        n56358) );
  NAND2_X1 U23258 ( .A1(n64990), .A2(n49910), .ZN(n4418) );
  NAND2_X2 U23263 ( .A1(n52479), .A2(n8023), .ZN(n5277) );
  AOI22_X1 U23269 ( .A1(n54524), .A2(n22572), .B1(n54511), .B2(n54512), .ZN(
        n54515) );
  NAND2_X2 U23276 ( .A1(n10165), .A2(n3622), .ZN(n36769) );
  NAND2_X2 U23277 ( .A1(n20872), .A2(n12263), .ZN(n28609) );
  INV_X4 U23282 ( .I(n19609), .ZN(n34614) );
  XOR2_X1 U23283 ( .A1(n31989), .A2(n21885), .Z(n12634) );
  NAND2_X1 U23288 ( .A1(n33982), .A2(n19450), .ZN(n19449) );
  INV_X4 U23291 ( .I(n17016), .ZN(n16766) );
  BUF_X2 U23292 ( .I(n15775), .Z(n20788) );
  XOR2_X1 U23296 ( .A1(n32077), .A2(n4433), .Z(n17239) );
  XOR2_X1 U23297 ( .A1(n13044), .A2(n31795), .Z(n4433) );
  NAND3_X2 U23298 ( .A1(n30130), .A2(n22353), .A3(n30131), .ZN(n32470) );
  AND2_X1 U23299 ( .A1(n36275), .A2(n7446), .Z(n5528) );
  NOR2_X2 U23303 ( .A1(n28278), .A2(n22043), .ZN(n28284) );
  NAND2_X2 U23304 ( .A1(n14470), .A2(n14471), .ZN(n15742) );
  NAND2_X1 U23306 ( .A1(n10247), .A2(n10248), .ZN(n23435) );
  NOR2_X2 U23307 ( .A1(n14890), .A2(n24958), .ZN(n10248) );
  OAI21_X1 U23309 ( .A1(n36160), .A2(n35922), .B(n35921), .ZN(n35923) );
  OAI21_X1 U23311 ( .A1(n53192), .A2(n25467), .B(n9963), .ZN(n52759) );
  AND2_X1 U23312 ( .A1(n42806), .A2(n43326), .Z(n8657) );
  XOR2_X1 U23313 ( .A1(n24274), .A2(n51128), .Z(n12294) );
  AOI22_X1 U23314 ( .A1(n47724), .A2(n47723), .B1(n47717), .B2(n47716), .ZN(
        n9227) );
  XOR2_X1 U23315 ( .A1(n12374), .A2(n4441), .Z(n16280) );
  NOR2_X2 U23316 ( .A1(n58999), .A2(n31051), .ZN(n20918) );
  NAND2_X1 U23325 ( .A1(n43493), .A2(n43914), .ZN(n20100) );
  NAND3_X1 U23328 ( .A1(n62270), .A2(n60545), .A3(n27656), .ZN(n4447) );
  INV_X4 U23332 ( .I(n1592), .ZN(n55550) );
  XOR2_X1 U23334 ( .A1(n8570), .A2(n51404), .Z(n4451) );
  NOR2_X2 U23336 ( .A1(n13487), .A2(n892), .ZN(n34395) );
  XOR2_X1 U23340 ( .A1(n233), .A2(n51543), .Z(n39237) );
  NOR3_X1 U23341 ( .A1(n55525), .A2(n4454), .A3(n55526), .ZN(n55532) );
  NOR2_X1 U23342 ( .A1(n55530), .A2(n55565), .ZN(n4454) );
  NAND2_X2 U23343 ( .A1(n64042), .A2(n64944), .ZN(n47831) );
  NAND2_X1 U23345 ( .A1(n39125), .A2(n64571), .ZN(n4455) );
  NAND4_X1 U23348 ( .A1(n4457), .A2(n27980), .A3(n29156), .A4(n1320), .ZN(
        n27265) );
  INV_X1 U23350 ( .I(n4459), .ZN(n36674) );
  AOI21_X1 U23351 ( .A1(n36670), .A2(n36671), .B(n4460), .ZN(n4459) );
  NAND2_X1 U23352 ( .A1(n36672), .A2(n36673), .ZN(n4460) );
  XOR2_X1 U23355 ( .A1(n38596), .A2(n19360), .Z(n18849) );
  XOR2_X1 U23356 ( .A1(n37149), .A2(n37150), .Z(n38596) );
  INV_X1 U23362 ( .I(n29543), .ZN(n4824) );
  NAND2_X1 U23371 ( .A1(n4465), .A2(n4463), .ZN(n13077) );
  NAND2_X1 U23372 ( .A1(n56489), .A2(n4464), .ZN(n4463) );
  INV_X1 U23373 ( .I(n4466), .ZN(n4465) );
  OAI21_X1 U23374 ( .A1(n56489), .A2(n56502), .B(n56510), .ZN(n4466) );
  NAND3_X1 U23383 ( .A1(n12150), .A2(n34333), .A3(n12149), .ZN(n12148) );
  OAI21_X1 U23394 ( .A1(n20659), .A2(n20658), .B(n53109), .ZN(n53087) );
  OR2_X1 U23401 ( .A1(n30509), .A2(n25989), .Z(n4477) );
  XOR2_X1 U23404 ( .A1(n51808), .A2(n51730), .Z(n51120) );
  XOR2_X1 U23406 ( .A1(n16521), .A2(n7394), .Z(n4479) );
  NOR2_X2 U23407 ( .A1(n1426), .A2(n35774), .ZN(n34427) );
  AOI22_X1 U23408 ( .A1(n56756), .A2(n56755), .B1(n61971), .B2(n56813), .ZN(
        n56760) );
  NOR4_X1 U23412 ( .A1(n17526), .A2(n17118), .A3(n17117), .A4(n27920), .ZN(
        n17116) );
  XOR2_X1 U23413 ( .A1(n10098), .A2(n44977), .Z(n11149) );
  NAND3_X2 U23416 ( .A1(n11321), .A2(n14877), .A3(n35355), .ZN(n39345) );
  NAND2_X1 U23417 ( .A1(n24670), .A2(n4485), .ZN(n55392) );
  INV_X2 U23418 ( .I(n10022), .ZN(n40494) );
  NAND2_X2 U23420 ( .A1(n14199), .A2(n22386), .ZN(n10088) );
  INV_X2 U23422 ( .I(n4487), .ZN(n40218) );
  XNOR2_X1 U23423 ( .A1(n39453), .A2(n39271), .ZN(n4487) );
  INV_X4 U23424 ( .I(n25427), .ZN(n23086) );
  AND3_X1 U23425 ( .A1(n53986), .A2(n53987), .A3(n53994), .Z(n23685) );
  NAND3_X1 U23426 ( .A1(n33376), .A2(n33377), .A3(n33629), .ZN(n33380) );
  XOR2_X1 U23427 ( .A1(n39391), .A2(n55610), .Z(n20684) );
  AND2_X1 U23429 ( .A1(n41556), .A2(n42140), .Z(n41344) );
  OR2_X1 U23431 ( .A1(n35184), .A2(n36259), .Z(n20945) );
  XOR2_X1 U23433 ( .A1(n39260), .A2(n39259), .Z(n25624) );
  XOR2_X1 U23434 ( .A1(n25623), .A2(n25622), .Z(n39260) );
  AND2_X1 U23441 ( .A1(n23881), .A2(n4495), .Z(n36240) );
  NAND2_X2 U23443 ( .A1(n3785), .A2(n24884), .ZN(n41699) );
  AOI21_X2 U23445 ( .A1(n26539), .A2(n26531), .B(n64174), .ZN(n27122) );
  XNOR2_X1 U23446 ( .A1(n38943), .A2(n38942), .ZN(n13390) );
  XOR2_X1 U23450 ( .A1(n51807), .A2(n17060), .Z(n17061) );
  INV_X2 U23456 ( .I(n4506), .ZN(n27366) );
  NOR3_X1 U23460 ( .A1(n61699), .A2(n35625), .A3(n445), .ZN(n32680) );
  INV_X1 U23463 ( .I(n24512), .ZN(n53844) );
  XOR2_X1 U23464 ( .A1(n4514), .A2(n5127), .Z(n12974) );
  INV_X1 U23465 ( .I(n30032), .ZN(n7180) );
  INV_X1 U23467 ( .I(n20310), .ZN(n9842) );
  AOI21_X1 U23468 ( .A1(n5092), .A2(n5091), .B(n23166), .ZN(n22591) );
  NAND3_X2 U23478 ( .A1(n46787), .A2(n46785), .A3(n46786), .ZN(n50088) );
  OAI21_X1 U23480 ( .A1(n20649), .A2(n26302), .B(n26330), .ZN(n26303) );
  XOR2_X1 U23485 ( .A1(n18641), .A2(n18638), .Z(n51606) );
  NOR3_X1 U23486 ( .A1(n30198), .A2(n30197), .A3(n59798), .ZN(n30194) );
  XOR2_X1 U23493 ( .A1(n10620), .A2(n44304), .Z(n44754) );
  NOR3_X2 U23494 ( .A1(n55013), .A2(n55014), .A3(n55012), .ZN(n55015) );
  AOI22_X1 U23496 ( .A1(n41349), .A2(n43078), .B1(n43072), .B2(n63792), .ZN(
        n4522) );
  INV_X2 U23499 ( .I(n13298), .ZN(n48564) );
  INV_X1 U23500 ( .I(n60930), .ZN(n13824) );
  NAND2_X2 U23503 ( .A1(n13864), .A2(n13865), .ZN(n14373) );
  OR3_X1 U23504 ( .A1(n5318), .A2(n54825), .A3(n54657), .Z(n54335) );
  XOR2_X1 U23507 ( .A1(n10847), .A2(n31688), .Z(n10408) );
  OR2_X1 U23520 ( .A1(n48558), .A2(n64036), .Z(n46787) );
  NAND2_X1 U23523 ( .A1(n26012), .A2(n8312), .ZN(n8311) );
  NAND2_X2 U23528 ( .A1(n34208), .A2(n34771), .ZN(n34759) );
  XOR2_X1 U23529 ( .A1(n4532), .A2(n9024), .Z(n19904) );
  INV_X2 U23533 ( .I(n4533), .ZN(n25867) );
  NAND3_X1 U23543 ( .A1(n56358), .A2(n4810), .A3(n56357), .ZN(n4809) );
  OR2_X1 U23544 ( .A1(n64155), .A2(n28410), .Z(n26514) );
  XOR2_X1 U23547 ( .A1(n15511), .A2(n20058), .Z(n32129) );
  NAND2_X2 U23548 ( .A1(n5858), .A2(n5855), .ZN(n20058) );
  INV_X2 U23552 ( .I(n28518), .ZN(n10239) );
  AND2_X1 U23553 ( .A1(n27717), .A2(n28518), .Z(n27718) );
  OAI21_X1 U23554 ( .A1(n4539), .A2(n4538), .B(n53809), .ZN(n53771) );
  NOR2_X1 U23555 ( .A1(n53776), .A2(n53790), .ZN(n4539) );
  OAI21_X1 U23556 ( .A1(n34450), .A2(n35644), .B(n22909), .ZN(n34451) );
  XNOR2_X1 U23560 ( .A1(n43621), .A2(n61662), .ZN(n4751) );
  XOR2_X1 U23561 ( .A1(n4543), .A2(n17217), .Z(n7019) );
  NAND2_X2 U23562 ( .A1(n4428), .A2(n12100), .ZN(n8632) );
  XOR2_X1 U23564 ( .A1(n44143), .A2(n6715), .Z(n5224) );
  NOR2_X1 U23565 ( .A1(n15883), .A2(n19526), .ZN(n17507) );
  NOR2_X2 U23568 ( .A1(n55569), .A2(n21272), .ZN(n55567) );
  NAND2_X2 U23570 ( .A1(n30752), .A2(n19929), .ZN(n18581) );
  XOR2_X1 U23575 ( .A1(n38707), .A2(n955), .Z(n4549) );
  INV_X2 U23579 ( .I(n12462), .ZN(n21100) );
  NAND2_X2 U23581 ( .A1(n28048), .A2(n64903), .ZN(n15156) );
  XOR2_X1 U23587 ( .A1(n51972), .A2(n61571), .Z(n51158) );
  NAND3_X2 U23588 ( .A1(n48090), .A2(n48091), .A3(n48092), .ZN(n48141) );
  INV_X4 U23592 ( .I(n27305), .ZN(n30538) );
  XOR2_X1 U23596 ( .A1(n44723), .A2(n4556), .Z(n25695) );
  XOR2_X1 U23600 ( .A1(n44817), .A2(n43009), .Z(n4558) );
  INV_X2 U23601 ( .I(n25405), .ZN(n40394) );
  INV_X2 U23603 ( .I(n55261), .ZN(n54996) );
  INV_X2 U23608 ( .I(n4560), .ZN(n6001) );
  NOR2_X1 U23610 ( .A1(n48801), .A2(n59004), .ZN(n48806) );
  NAND2_X2 U23613 ( .A1(n4685), .A2(n19373), .ZN(n9329) );
  OAI22_X1 U23619 ( .A1(n8015), .A2(n8014), .B1(n26655), .B2(n27577), .ZN(
        n10412) );
  NAND2_X1 U23620 ( .A1(n26451), .A2(n5292), .ZN(n5291) );
  NOR2_X1 U23621 ( .A1(n15941), .A2(n16685), .ZN(n20368) );
  INV_X4 U23626 ( .I(n4567), .ZN(n30799) );
  NAND2_X2 U23627 ( .A1(n4568), .A2(n26498), .ZN(n4567) );
  XOR2_X1 U23630 ( .A1(n33914), .A2(n15678), .Z(n15677) );
  INV_X2 U23631 ( .I(n4570), .ZN(n11084) );
  NAND2_X2 U23634 ( .A1(n976), .A2(n42230), .ZN(n17077) );
  XOR2_X1 U23636 ( .A1(n15733), .A2(n4572), .Z(n32522) );
  XOR2_X1 U23637 ( .A1(n32590), .A2(n32521), .Z(n4572) );
  NAND2_X1 U23638 ( .A1(n56101), .A2(n24092), .ZN(n20876) );
  NOR2_X2 U23639 ( .A1(n33718), .A2(n12350), .ZN(n34509) );
  XOR2_X1 U23644 ( .A1(n4576), .A2(n44847), .Z(n5898) );
  XOR2_X1 U23645 ( .A1(n44383), .A2(n7424), .Z(n4576) );
  AND3_X1 U23650 ( .A1(n24121), .A2(n32774), .A3(n23881), .Z(n32778) );
  NOR2_X1 U23651 ( .A1(n12285), .A2(n40337), .ZN(n40339) );
  NAND2_X2 U23653 ( .A1(n18335), .A2(n56393), .ZN(n56574) );
  NAND3_X1 U23655 ( .A1(n12285), .A2(n19611), .A3(n9802), .ZN(n40336) );
  XNOR2_X1 U23657 ( .A1(n45852), .A2(n7034), .ZN(n4859) );
  XNOR2_X1 U23658 ( .A1(n45096), .A2(n1021), .ZN(n7145) );
  NOR2_X2 U23665 ( .A1(n5258), .A2(n23839), .ZN(n50238) );
  OR2_X1 U23668 ( .A1(n41554), .A2(n9914), .Z(n4588) );
  XOR2_X1 U23669 ( .A1(n59854), .A2(n62985), .Z(n4589) );
  INV_X2 U23676 ( .I(n47843), .ZN(n47828) );
  INV_X4 U23679 ( .I(n49548), .ZN(n15319) );
  XOR2_X1 U23681 ( .A1(n9826), .A2(n4595), .Z(n44932) );
  XOR2_X1 U23682 ( .A1(n32396), .A2(n22950), .Z(n4595) );
  NAND2_X2 U23683 ( .A1(n13926), .A2(n24136), .ZN(n24138) );
  OAI21_X1 U23692 ( .A1(n5619), .A2(n53066), .B(n53109), .ZN(n4601) );
  INV_X2 U23699 ( .I(n4604), .ZN(n26691) );
  NAND3_X2 U23701 ( .A1(n16611), .A2(n16608), .A3(n16236), .ZN(n23216) );
  XOR2_X1 U23705 ( .A1(n19204), .A2(n14665), .Z(n24827) );
  INV_X1 U23706 ( .I(n34136), .ZN(n19538) );
  AND2_X1 U23709 ( .A1(n1417), .A2(n36742), .Z(n35072) );
  XOR2_X1 U23711 ( .A1(n37518), .A2(n4691), .Z(n37527) );
  XOR2_X1 U23712 ( .A1(n24787), .A2(n26087), .Z(n12603) );
  OAI21_X1 U23718 ( .A1(n10218), .A2(n14560), .B(n59599), .ZN(n52291) );
  BUF_X4 U23719 ( .I(n14409), .Z(n12677) );
  NAND3_X2 U23722 ( .A1(n23094), .A2(n20988), .A3(n28079), .ZN(n29994) );
  NOR2_X1 U23730 ( .A1(n12304), .A2(n11717), .ZN(n11714) );
  XOR2_X1 U23731 ( .A1(n19204), .A2(n50494), .Z(n32667) );
  XOR2_X1 U23736 ( .A1(n39371), .A2(n5183), .Z(n4616) );
  XOR2_X1 U23746 ( .A1(n4621), .A2(n20302), .Z(n52005) );
  XOR2_X1 U23747 ( .A1(n22338), .A2(n52004), .Z(n4621) );
  NAND2_X2 U23748 ( .A1(n5794), .A2(n5791), .ZN(n5787) );
  XOR2_X1 U23749 ( .A1(n4622), .A2(n54386), .Z(Plaintext[68]) );
  NAND2_X2 U23753 ( .A1(n34914), .A2(n9456), .ZN(n36940) );
  NOR2_X2 U23754 ( .A1(n4629), .A2(n47872), .ZN(n47873) );
  XOR2_X1 U23756 ( .A1(n4630), .A2(n4631), .Z(n20739) );
  NAND2_X1 U23758 ( .A1(n28323), .A2(n28325), .ZN(n14534) );
  NOR3_X1 U23759 ( .A1(n30302), .A2(n30296), .A3(n28921), .ZN(n4633) );
  OAI22_X1 U23761 ( .A1(n61909), .A2(n10653), .B1(n47858), .B2(n23311), .ZN(
        n47856) );
  INV_X1 U23767 ( .I(n34440), .ZN(n12065) );
  NAND2_X1 U23769 ( .A1(n20439), .A2(n14192), .ZN(n14191) );
  NOR2_X1 U23781 ( .A1(n35339), .A2(n35338), .ZN(n6131) );
  XNOR2_X1 U23782 ( .A1(n38647), .A2(n38646), .ZN(n9781) );
  NAND2_X1 U23784 ( .A1(n19068), .A2(n52845), .ZN(n12289) );
  NAND2_X2 U23789 ( .A1(n4642), .A2(n22746), .ZN(n40891) );
  INV_X1 U23790 ( .I(n33509), .ZN(n34539) );
  OR2_X1 U23797 ( .A1(n23095), .A2(n56541), .Z(n56382) );
  XOR2_X1 U23802 ( .A1(n43782), .A2(n21142), .Z(n18012) );
  XOR2_X1 U23803 ( .A1(n64714), .A2(n15354), .Z(n43782) );
  NOR2_X1 U23804 ( .A1(n18574), .A2(n17392), .ZN(n17391) );
  OR2_X2 U23809 ( .A1(n19609), .A2(n31026), .Z(n7849) );
  NOR2_X2 U23812 ( .A1(n8248), .A2(n52952), .ZN(n20177) );
  AND2_X1 U23813 ( .A1(n19845), .A2(n8256), .Z(n8254) );
  NAND3_X2 U23823 ( .A1(n4664), .A2(n49907), .A3(n49906), .ZN(n49917) );
  NAND3_X1 U23827 ( .A1(n53569), .A2(n53568), .A3(n53567), .ZN(n4666) );
  OAI21_X1 U23829 ( .A1(n45177), .A2(n61510), .B(n5940), .ZN(n45178) );
  NOR2_X1 U23830 ( .A1(n43115), .A2(n16385), .ZN(n9749) );
  AND3_X2 U23832 ( .A1(n29678), .A2(n29680), .A3(n29679), .Z(n10585) );
  NOR2_X1 U23836 ( .A1(n42227), .A2(n42228), .ZN(n12736) );
  XOR2_X1 U23837 ( .A1(n38287), .A2(n38144), .Z(n6332) );
  NAND2_X2 U23843 ( .A1(n47502), .A2(n21044), .ZN(n45479) );
  XOR2_X1 U23846 ( .A1(n4671), .A2(n20742), .Z(n13721) );
  XOR2_X1 U23847 ( .A1(n58738), .A2(n11269), .Z(n4671) );
  OR2_X1 U23853 ( .A1(n5705), .A2(n48540), .Z(n5704) );
  XOR2_X1 U23855 ( .A1(n7678), .A2(n44834), .Z(n4674) );
  XOR2_X1 U23858 ( .A1(n4675), .A2(n39657), .Z(n24932) );
  XOR2_X1 U23859 ( .A1(n39658), .A2(n6113), .Z(n4675) );
  NAND2_X2 U23864 ( .A1(n29154), .A2(n27397), .ZN(n8528) );
  NAND2_X1 U23870 ( .A1(n4683), .A2(n1510), .ZN(n4682) );
  INV_X4 U23873 ( .I(n6100), .ZN(n22657) );
  INV_X1 U23875 ( .I(n18883), .ZN(n9818) );
  XOR2_X1 U23880 ( .A1(n22561), .A2(n16122), .Z(n39497) );
  INV_X2 U23881 ( .I(n17097), .ZN(n21090) );
  NOR2_X2 U23883 ( .A1(n1608), .A2(n54324), .ZN(n8375) );
  INV_X1 U23890 ( .I(n38419), .ZN(n5305) );
  NOR3_X1 U23897 ( .A1(n11715), .A2(n11714), .A3(n51015), .ZN(n11713) );
  AND2_X1 U23901 ( .A1(n26638), .A2(n26632), .Z(n20195) );
  NAND2_X2 U23902 ( .A1(n23734), .A2(n24316), .ZN(n30293) );
  AND2_X1 U23904 ( .A1(n49361), .A2(n49362), .Z(n4695) );
  XOR2_X1 U23905 ( .A1(n4696), .A2(n15241), .Z(n6592) );
  INV_X2 U23907 ( .I(n50045), .ZN(n20199) );
  XOR2_X1 U23908 ( .A1(n39371), .A2(n4697), .Z(n8004) );
  INV_X1 U23909 ( .I(n39369), .ZN(n4697) );
  INV_X4 U23913 ( .I(n21187), .ZN(n34841) );
  NOR2_X2 U23916 ( .A1(n23636), .A2(n26641), .ZN(n27178) );
  OAI21_X1 U23921 ( .A1(n41434), .A2(n11645), .B(n41433), .ZN(n12188) );
  NAND3_X2 U23922 ( .A1(n7933), .A2(n36472), .A3(n36477), .ZN(n36151) );
  XOR2_X1 U23924 ( .A1(Ciphertext[46]), .A2(Key[119]), .Z(n6012) );
  NOR2_X1 U23930 ( .A1(n54326), .A2(n64681), .ZN(n6465) );
  NOR2_X1 U23938 ( .A1(n64135), .A2(n62139), .ZN(n17087) );
  NOR2_X1 U23943 ( .A1(n21421), .A2(n2119), .ZN(n30323) );
  NOR2_X2 U23947 ( .A1(n25532), .A2(n29295), .ZN(n7437) );
  NAND2_X1 U23949 ( .A1(n57912), .A2(n11887), .ZN(n11888) );
  NAND2_X1 U23950 ( .A1(n11888), .A2(n11886), .ZN(n11885) );
  INV_X2 U23955 ( .I(n20508), .ZN(n20509) );
  NOR2_X1 U23960 ( .A1(n45947), .A2(n13356), .ZN(n4713) );
  NAND2_X2 U23965 ( .A1(n42324), .A2(n41675), .ZN(n43012) );
  XOR2_X1 U23972 ( .A1(n41440), .A2(n23967), .Z(n40701) );
  XOR2_X1 U23974 ( .A1(n31884), .A2(n33884), .Z(n31886) );
  INV_X2 U23978 ( .I(n53014), .ZN(n53795) );
  XOR2_X1 U23985 ( .A1(n4726), .A2(n9674), .Z(n44420) );
  XOR2_X1 U23986 ( .A1(n5360), .A2(n44611), .Z(n4726) );
  XOR2_X1 U23988 ( .A1(n60717), .A2(n13365), .Z(n4727) );
  XOR2_X1 U23990 ( .A1(n4728), .A2(n7687), .Z(n7686) );
  XOR2_X1 U23991 ( .A1(n38179), .A2(n5822), .Z(n4728) );
  NOR2_X1 U23992 ( .A1(n15968), .A2(n17367), .ZN(n21705) );
  AND2_X1 U24000 ( .A1(n44194), .A2(n6081), .Z(n44776) );
  AND2_X1 U24004 ( .A1(n4729), .A2(n40326), .Z(n23250) );
  NAND2_X1 U24005 ( .A1(n40318), .A2(n20751), .ZN(n4729) );
  AND4_X1 U24007 ( .A1(n38423), .A2(n38424), .A3(n38422), .A4(n21295), .Z(
        n5474) );
  XOR2_X1 U24010 ( .A1(n2452), .A2(n44337), .Z(n4732) );
  INV_X2 U24014 ( .I(n4737), .ZN(n15809) );
  XNOR2_X1 U24015 ( .A1(n9180), .A2(n14715), .ZN(n4737) );
  OAI21_X1 U24017 ( .A1(n44773), .A2(n44661), .B(n4738), .ZN(n11526) );
  NAND2_X2 U24019 ( .A1(n27948), .A2(n23770), .ZN(n19059) );
  NOR2_X1 U24020 ( .A1(n14418), .A2(n47541), .ZN(n46460) );
  NOR2_X2 U24021 ( .A1(n56191), .A2(n56182), .ZN(n56169) );
  NAND3_X2 U24023 ( .A1(n25370), .A2(n25371), .A3(n29953), .ZN(n31345) );
  INV_X1 U24024 ( .I(n28256), .ZN(n27943) );
  OR2_X1 U24025 ( .A1(n28256), .A2(n12070), .Z(n27944) );
  NAND2_X2 U24031 ( .A1(n1575), .A2(n27494), .ZN(n29304) );
  NOR2_X2 U24032 ( .A1(n47123), .A2(n48557), .ZN(n48089) );
  NAND3_X1 U24034 ( .A1(n18841), .A2(n60187), .A3(n30167), .ZN(n18840) );
  AND2_X1 U24036 ( .A1(n30068), .A2(n30067), .Z(n4744) );
  OR2_X1 U24037 ( .A1(n48239), .A2(n60560), .Z(n18633) );
  NAND2_X1 U24038 ( .A1(n6718), .A2(n24945), .ZN(n5164) );
  INV_X1 U24042 ( .I(n29608), .ZN(n28665) );
  XOR2_X1 U24047 ( .A1(n24548), .A2(n33272), .Z(n7141) );
  NAND2_X1 U24050 ( .A1(n12007), .A2(n12764), .ZN(n12006) );
  OR2_X1 U24051 ( .A1(n61177), .A2(n27098), .Z(n6857) );
  NOR2_X2 U24052 ( .A1(n13858), .A2(n55885), .ZN(n55895) );
  NAND2_X1 U24056 ( .A1(n33968), .A2(n33969), .ZN(n9541) );
  INV_X4 U24060 ( .I(n9536), .ZN(n9593) );
  NOR2_X1 U24061 ( .A1(n19604), .A2(n6348), .ZN(n6347) );
  NAND3_X1 U24065 ( .A1(n26991), .A2(n28810), .A3(n26990), .ZN(n27000) );
  OAI21_X2 U24067 ( .A1(n52772), .A2(n52771), .B(n6792), .ZN(n52776) );
  OAI21_X1 U24070 ( .A1(n34861), .A2(n4756), .B(n37029), .ZN(n19158) );
  NAND2_X1 U24071 ( .A1(n35907), .A2(n7598), .ZN(n4756) );
  XOR2_X1 U24072 ( .A1(n51507), .A2(n4757), .Z(n49416) );
  XOR2_X1 U24074 ( .A1(n12669), .A2(n2823), .Z(n4759) );
  INV_X1 U24075 ( .I(n45267), .ZN(n4760) );
  XOR2_X1 U24078 ( .A1(n4762), .A2(n38741), .Z(n36370) );
  NAND2_X2 U24081 ( .A1(n30699), .A2(n30698), .ZN(n32663) );
  XOR2_X1 U24083 ( .A1(n8385), .A2(n9009), .Z(n11801) );
  NAND2_X1 U24084 ( .A1(n4765), .A2(n60593), .ZN(n16992) );
  NOR3_X1 U24087 ( .A1(n23063), .A2(n22042), .A3(n50426), .ZN(n45443) );
  XOR2_X1 U24091 ( .A1(n9729), .A2(n4771), .Z(n47011) );
  XOR2_X1 U24092 ( .A1(n16932), .A2(n19947), .Z(n4771) );
  OAI22_X1 U24094 ( .A1(n42733), .A2(n43359), .B1(n1491), .B2(n42734), .ZN(
        n4774) );
  INV_X1 U24096 ( .I(n30785), .ZN(n16648) );
  OAI21_X1 U24098 ( .A1(n26789), .A2(n26788), .B(n26787), .ZN(n17529) );
  OR2_X1 U24100 ( .A1(n36052), .A2(n17775), .Z(n34855) );
  XOR2_X1 U24101 ( .A1(n4775), .A2(n31236), .Z(n23027) );
  XOR2_X1 U24102 ( .A1(n5521), .A2(n1823), .Z(n31236) );
  XOR2_X1 U24105 ( .A1(n33189), .A2(n33188), .Z(n4776) );
  NAND2_X2 U24109 ( .A1(n30802), .A2(n29934), .ZN(n18120) );
  OAI22_X1 U24111 ( .A1(n61697), .A2(n56173), .B1(n56191), .B2(n56162), .ZN(
        n18173) );
  NOR3_X1 U24115 ( .A1(n5429), .A2(n5428), .A3(n16922), .ZN(n5427) );
  NAND2_X1 U24116 ( .A1(n49681), .A2(n5427), .ZN(n5426) );
  XOR2_X1 U24123 ( .A1(n37385), .A2(n37384), .Z(n4782) );
  INV_X2 U24125 ( .I(n4784), .ZN(n17747) );
  NAND2_X2 U24128 ( .A1(n57471), .A2(n4785), .ZN(n16389) );
  NAND3_X1 U24130 ( .A1(n34393), .A2(n19312), .A3(n16240), .ZN(n34400) );
  XOR2_X1 U24135 ( .A1(n4790), .A2(n9149), .Z(n9531) );
  XOR2_X1 U24136 ( .A1(n26025), .A2(n13658), .Z(n4790) );
  NAND2_X1 U24137 ( .A1(n47267), .A2(n65145), .ZN(n47268) );
  OR2_X2 U24140 ( .A1(n50461), .A2(n24390), .Z(n53858) );
  XOR2_X1 U24141 ( .A1(n11860), .A2(n16760), .Z(n50461) );
  INV_X2 U24142 ( .I(n34777), .ZN(n34273) );
  NAND2_X2 U24143 ( .A1(n19457), .A2(n34783), .ZN(n34777) );
  XOR2_X1 U24151 ( .A1(n52602), .A2(n14861), .Z(n14096) );
  NAND2_X1 U24153 ( .A1(n46908), .A2(n44196), .ZN(n17032) );
  NOR2_X2 U24154 ( .A1(n28256), .A2(n29161), .ZN(n28266) );
  XOR2_X1 U24156 ( .A1(n10477), .A2(n23124), .Z(n4797) );
  NAND4_X2 U24158 ( .A1(n18389), .A2(n28268), .A3(n28262), .A4(n18388), .ZN(
        n4799) );
  OAI21_X1 U24171 ( .A1(n45545), .A2(n47971), .B(n13645), .ZN(n5697) );
  XOR2_X1 U24174 ( .A1(n24348), .A2(n24349), .Z(n24347) );
  XOR2_X1 U24178 ( .A1(n4809), .A2(n24098), .Z(Plaintext[155]) );
  AND2_X1 U24179 ( .A1(n56356), .A2(n56355), .Z(n4810) );
  XOR2_X1 U24180 ( .A1(n4811), .A2(n50592), .Z(n50593) );
  XOR2_X1 U24183 ( .A1(n8527), .A2(n4953), .Z(n8526) );
  INV_X2 U24189 ( .I(n4813), .ZN(n9601) );
  XOR2_X1 U24191 ( .A1(n25337), .A2(n4814), .Z(n25897) );
  XOR2_X1 U24194 ( .A1(n4816), .A2(n37689), .Z(n38636) );
  NOR2_X2 U24199 ( .A1(n60202), .A2(n23140), .ZN(n30410) );
  XOR2_X1 U24207 ( .A1(n51250), .A2(n23939), .Z(n14078) );
  XOR2_X1 U24208 ( .A1(n24368), .A2(n49985), .Z(n51250) );
  NOR2_X2 U24212 ( .A1(n41152), .A2(n4819), .ZN(n40716) );
  XOR2_X1 U24215 ( .A1(n46442), .A2(n45145), .Z(n20905) );
  NAND2_X2 U24216 ( .A1(n14444), .A2(n40917), .ZN(n46442) );
  AND3_X1 U24218 ( .A1(n28707), .A2(n58448), .A3(n15269), .Z(n12060) );
  NOR2_X1 U24229 ( .A1(n25650), .A2(n23298), .ZN(n22995) );
  AND2_X1 U24236 ( .A1(n40316), .A2(n23654), .Z(n16017) );
  NOR2_X1 U24238 ( .A1(n40095), .A2(n42413), .ZN(n13408) );
  NAND2_X2 U24239 ( .A1(n4832), .A2(n19546), .ZN(n25051) );
  XOR2_X1 U24241 ( .A1(n4833), .A2(n21869), .Z(n21868) );
  XOR2_X1 U24242 ( .A1(n33898), .A2(n32009), .Z(n4833) );
  XNOR2_X1 U24243 ( .A1(n52030), .A2(n52029), .ZN(n14458) );
  XOR2_X1 U24244 ( .A1(n24689), .A2(n46511), .Z(n13719) );
  NAND2_X2 U24245 ( .A1(n20985), .A2(n22782), .ZN(n5476) );
  XOR2_X1 U24250 ( .A1(n52445), .A2(n51929), .Z(n10994) );
  NAND2_X2 U24251 ( .A1(n14858), .A2(n14859), .ZN(n52445) );
  INV_X4 U24256 ( .I(n31470), .ZN(n5410) );
  OAI21_X1 U24257 ( .A1(n55374), .A2(n9065), .B(n55373), .ZN(n55375) );
  NAND3_X1 U24259 ( .A1(n42544), .A2(n42545), .A3(n42543), .ZN(n10073) );
  NAND2_X1 U24260 ( .A1(n26494), .A2(n26495), .ZN(n4840) );
  OR2_X1 U24266 ( .A1(n53561), .A2(n1599), .Z(n53560) );
  XOR2_X1 U24268 ( .A1(n4842), .A2(n23858), .Z(Plaintext[33]) );
  XOR2_X1 U24274 ( .A1(n38960), .A2(n4845), .Z(n13062) );
  XOR2_X1 U24275 ( .A1(n23181), .A2(n790), .Z(n4845) );
  INV_X4 U24277 ( .I(n14165), .ZN(n41400) );
  INV_X4 U24278 ( .I(n17977), .ZN(n43155) );
  INV_X2 U24280 ( .I(n4850), .ZN(n8228) );
  AND2_X1 U24282 ( .A1(n39419), .A2(n11126), .Z(n11130) );
  XOR2_X1 U24283 ( .A1(n9217), .A2(n9219), .Z(n4854) );
  NAND2_X1 U24284 ( .A1(n56266), .A2(n5670), .ZN(n5669) );
  NAND2_X1 U24286 ( .A1(n61696), .A2(n4855), .ZN(n53804) );
  NAND2_X1 U24287 ( .A1(n53789), .A2(n53793), .ZN(n4855) );
  XOR2_X1 U24291 ( .A1(n63031), .A2(n19330), .Z(n46092) );
  XOR2_X1 U24293 ( .A1(n4871), .A2(n4859), .Z(n4858) );
  NOR3_X2 U24297 ( .A1(n19907), .A2(n4863), .A3(n19446), .ZN(n51891) );
  NAND2_X2 U24298 ( .A1(n22694), .A2(n49940), .ZN(n48318) );
  XOR2_X1 U24303 ( .A1(n10292), .A2(n53375), .Z(n8229) );
  NOR2_X2 U24304 ( .A1(n61452), .A2(n4851), .ZN(n5902) );
  XNOR2_X1 U24306 ( .A1(n6516), .A2(n39547), .ZN(n5854) );
  NAND4_X2 U24308 ( .A1(n4873), .A2(n10374), .A3(n10373), .A4(n40955), .ZN(
        n9525) );
  NAND4_X1 U24310 ( .A1(n4874), .A2(n55585), .A3(n55584), .A4(n55583), .ZN(
        n22851) );
  XOR2_X1 U24312 ( .A1(n15074), .A2(n45356), .Z(n4876) );
  OAI21_X1 U24313 ( .A1(n56777), .A2(n56790), .B(n23030), .ZN(n56782) );
  AND2_X2 U24317 ( .A1(n13752), .A2(n26067), .Z(n23399) );
  NOR2_X2 U24318 ( .A1(n7760), .A2(n13955), .ZN(n7110) );
  NAND2_X2 U24319 ( .A1(n33643), .A2(n33370), .ZN(n33219) );
  INV_X2 U24320 ( .I(n39886), .ZN(n42489) );
  NAND2_X2 U24321 ( .A1(n21050), .A2(n39886), .ZN(n6467) );
  XNOR2_X1 U24322 ( .A1(n10781), .A2(n10778), .ZN(n39886) );
  OAI21_X2 U24334 ( .A1(n4884), .A2(n60860), .B(n20248), .ZN(n19537) );
  NAND4_X2 U24336 ( .A1(n10970), .A2(n41972), .A3(n42694), .A4(n20244), .ZN(
        n42707) );
  XOR2_X1 U24337 ( .A1(n6688), .A2(n4886), .Z(n6686) );
  XOR2_X1 U24338 ( .A1(n17201), .A2(n24346), .Z(n4886) );
  NAND2_X2 U24340 ( .A1(n23350), .A2(n20244), .ZN(n42699) );
  XOR2_X1 U24341 ( .A1(n4887), .A2(n15841), .Z(n34359) );
  INV_X2 U24344 ( .I(n55316), .ZN(n54999) );
  XOR2_X1 U24346 ( .A1(n39006), .A2(n39005), .Z(n11462) );
  NAND2_X1 U24347 ( .A1(n36484), .A2(n19038), .ZN(n23881) );
  XOR2_X1 U24351 ( .A1(n5234), .A2(n20633), .Z(n24858) );
  NAND2_X2 U24353 ( .A1(n7517), .A2(n18339), .ZN(n33613) );
  NOR2_X1 U24354 ( .A1(n47931), .A2(n47930), .ZN(n15605) );
  NOR2_X2 U24356 ( .A1(n37198), .A2(n40934), .ZN(n4968) );
  INV_X1 U24358 ( .I(n41141), .ZN(n6969) );
  NAND2_X1 U24360 ( .A1(n22313), .A2(n22314), .ZN(n49121) );
  NAND2_X2 U24369 ( .A1(n12598), .A2(n25838), .ZN(n51264) );
  NOR2_X1 U24370 ( .A1(n34683), .A2(n34684), .ZN(n7300) );
  NAND2_X1 U24371 ( .A1(n28423), .A2(n63890), .ZN(n8089) );
  XNOR2_X1 U24376 ( .A1(n8417), .A2(n20478), .ZN(n4899) );
  INV_X1 U24377 ( .I(n45757), .ZN(n6661) );
  NAND2_X2 U24378 ( .A1(n37292), .A2(n15449), .ZN(n37858) );
  AND2_X1 U24391 ( .A1(n7692), .A2(n48826), .Z(n7653) );
  XOR2_X1 U24392 ( .A1(n4904), .A2(n1122), .Z(n12810) );
  NOR2_X1 U24403 ( .A1(n22886), .A2(n43214), .ZN(n11537) );
  OAI21_X1 U24404 ( .A1(n19563), .A2(n34979), .B(n33508), .ZN(n10046) );
  NOR2_X2 U24405 ( .A1(n40063), .A2(n40308), .ZN(n17930) );
  AND3_X2 U24410 ( .A1(n15395), .A2(n26241), .A3(n26027), .Z(n15394) );
  NAND3_X2 U24415 ( .A1(n12492), .A2(n12491), .A3(n7434), .ZN(n25326) );
  NAND2_X2 U24423 ( .A1(n52862), .A2(n52861), .ZN(n52665) );
  AND2_X1 U24426 ( .A1(n19287), .A2(n17689), .Z(n15986) );
  OR2_X1 U24428 ( .A1(n5872), .A2(n62720), .Z(n21816) );
  XOR2_X1 U24430 ( .A1(n23852), .A2(n52623), .Z(n9236) );
  XOR2_X1 U24432 ( .A1(n21098), .A2(n57420), .Z(n4922) );
  OAI21_X1 U24438 ( .A1(n55685), .A2(n55487), .B(n11164), .ZN(n19133) );
  AND2_X1 U24444 ( .A1(n8222), .A2(n5553), .Z(n52312) );
  XOR2_X1 U24446 ( .A1(n13359), .A2(n13228), .Z(n18190) );
  NAND2_X2 U24452 ( .A1(n5944), .A2(n61502), .ZN(n6333) );
  INV_X2 U24455 ( .I(n42619), .ZN(n43548) );
  XOR2_X1 U24460 ( .A1(n4928), .A2(n16206), .Z(n9872) );
  NAND2_X1 U24461 ( .A1(n18183), .A2(n44789), .ZN(n18182) );
  NOR2_X1 U24462 ( .A1(n18182), .A2(n18181), .ZN(n9825) );
  OAI22_X1 U24466 ( .A1(n21020), .A2(n6033), .B1(n33683), .B2(n12413), .ZN(
        n33686) );
  NAND3_X1 U24468 ( .A1(n1490), .A2(n12196), .A3(n11223), .ZN(n11222) );
  XOR2_X1 U24470 ( .A1(n56988), .A2(n13920), .Z(n4929) );
  INV_X2 U24472 ( .I(n4930), .ZN(n8121) );
  OR2_X1 U24477 ( .A1(n26502), .A2(n18112), .Z(n16174) );
  XOR2_X1 U24478 ( .A1(n51011), .A2(n52549), .Z(n12040) );
  XOR2_X1 U24479 ( .A1(n50114), .A2(n50113), .Z(n51011) );
  INV_X1 U24480 ( .I(n7915), .ZN(n7914) );
  NOR2_X2 U24481 ( .A1(n4934), .A2(n27006), .ZN(n31122) );
  XOR2_X1 U24488 ( .A1(n36863), .A2(n16052), .Z(n4936) );
  XOR2_X1 U24489 ( .A1(n4937), .A2(n21316), .Z(n8384) );
  XOR2_X1 U24490 ( .A1(n45254), .A2(n64837), .Z(n4937) );
  AOI22_X1 U24492 ( .A1(n14837), .A2(n56018), .B1(n56020), .B2(n60672), .ZN(
        n4940) );
  NAND2_X2 U24495 ( .A1(n19852), .A2(n27071), .ZN(n11621) );
  NOR2_X2 U24503 ( .A1(n28039), .A2(n9685), .ZN(n28228) );
  XOR2_X1 U24504 ( .A1(n11700), .A2(n1449), .Z(n17939) );
  NOR3_X2 U24510 ( .A1(n3691), .A2(n37210), .A3(n37225), .ZN(n36613) );
  INV_X2 U24511 ( .I(n5263), .ZN(n14919) );
  INV_X4 U24512 ( .I(n14919), .ZN(n55401) );
  NOR2_X2 U24525 ( .A1(n17496), .A2(n19830), .ZN(n8982) );
  XOR2_X1 U24526 ( .A1(n4950), .A2(n12022), .Z(n8668) );
  XOR2_X1 U24527 ( .A1(n7079), .A2(n23491), .Z(n4950) );
  NOR2_X2 U24528 ( .A1(n24940), .A2(n26720), .ZN(n29134) );
  INV_X2 U24530 ( .I(n33144), .ZN(n4953) );
  INV_X1 U24531 ( .I(n25982), .ZN(n20385) );
  OAI22_X1 U24534 ( .A1(n4955), .A2(n55372), .B1(n55362), .B2(n15703), .ZN(
        n55337) );
  XOR2_X1 U24536 ( .A1(n4958), .A2(n21993), .Z(n48060) );
  XOR2_X1 U24538 ( .A1(n50038), .A2(n51813), .Z(n6299) );
  XOR2_X1 U24539 ( .A1(n50964), .A2(n6004), .Z(n50038) );
  XOR2_X1 U24540 ( .A1(n31687), .A2(n32596), .Z(n10847) );
  XOR2_X1 U24541 ( .A1(n31317), .A2(n32591), .Z(n31687) );
  XOR2_X1 U24544 ( .A1(n4960), .A2(n11191), .Z(n10243) );
  OAI22_X1 U24549 ( .A1(n16334), .A2(n63202), .B1(n16543), .B2(n16333), .ZN(
        n49996) );
  NAND3_X2 U24550 ( .A1(n4961), .A2(n10777), .A3(n29723), .ZN(n22978) );
  AND2_X1 U24551 ( .A1(n29724), .A2(n29886), .Z(n4961) );
  NAND2_X2 U24555 ( .A1(n21228), .A2(n21227), .ZN(n5435) );
  NOR2_X2 U24556 ( .A1(n4962), .A2(n53432), .ZN(n53462) );
  NAND2_X1 U24557 ( .A1(n23437), .A2(n22689), .ZN(n4962) );
  XOR2_X1 U24559 ( .A1(n32412), .A2(n32318), .Z(n21986) );
  OAI21_X1 U24561 ( .A1(n53472), .A2(n53473), .B(n53514), .ZN(n4963) );
  BUF_X4 U24562 ( .I(n16420), .Z(n16337) );
  XOR2_X1 U24572 ( .A1(n32582), .A2(n24666), .Z(n5252) );
  INV_X4 U24574 ( .I(n23874), .ZN(n53355) );
  NAND3_X1 U24579 ( .A1(n8582), .A2(n45966), .A3(n45960), .ZN(n45227) );
  OAI21_X1 U24580 ( .A1(n4978), .A2(n55820), .B(n4977), .ZN(n55783) );
  XOR2_X1 U24581 ( .A1(n22933), .A2(n21403), .Z(n4978) );
  NOR2_X2 U24583 ( .A1(n9200), .A2(n65230), .ZN(n41540) );
  AND2_X1 U24587 ( .A1(n31095), .A2(n31094), .Z(n4982) );
  XOR2_X1 U24588 ( .A1(n21088), .A2(n8821), .Z(n10285) );
  INV_X4 U24593 ( .I(n15215), .ZN(n39028) );
  AND2_X1 U24602 ( .A1(n6519), .A2(n27292), .Z(n18177) );
  NOR2_X1 U24603 ( .A1(n5669), .A2(n5667), .ZN(n22302) );
  NAND2_X1 U24604 ( .A1(n28150), .A2(n28847), .ZN(n4988) );
  XOR2_X1 U24606 ( .A1(n7862), .A2(n4991), .Z(n5293) );
  NOR2_X1 U24612 ( .A1(n16381), .A2(n6184), .ZN(n49159) );
  INV_X2 U24617 ( .I(n17494), .ZN(n46307) );
  BUF_X2 U24630 ( .I(n16971), .Z(n4999) );
  XOR2_X1 U24634 ( .A1(n50863), .A2(n1465), .Z(n16376) );
  INV_X2 U24637 ( .I(n27105), .ZN(n27565) );
  AND2_X1 U24639 ( .A1(n42749), .A2(n65147), .Z(n7373) );
  AND2_X1 U24641 ( .A1(n37407), .A2(n16426), .Z(n5003) );
  XOR2_X1 U24652 ( .A1(n5867), .A2(n21990), .Z(n5868) );
  INV_X1 U24655 ( .I(n8475), .ZN(n47364) );
  OR2_X1 U24656 ( .A1(n8475), .A2(n1387), .Z(n9451) );
  NOR2_X1 U24657 ( .A1(n26713), .A2(n26718), .ZN(n26716) );
  NOR2_X1 U24663 ( .A1(n56245), .A2(n14601), .ZN(n14600) );
  XOR2_X1 U24671 ( .A1(n5023), .A2(n46127), .Z(n15457) );
  INV_X1 U24672 ( .I(n12697), .ZN(n51937) );
  XOR2_X1 U24675 ( .A1(n5028), .A2(n19798), .Z(n41147) );
  OAI22_X2 U24680 ( .A1(n10998), .A2(n39938), .B1(n59650), .B2(n43836), .ZN(
        n5030) );
  NAND2_X2 U24683 ( .A1(n5690), .A2(n5031), .ZN(n22674) );
  XOR2_X1 U24687 ( .A1(n5155), .A2(n6745), .Z(n5037) );
  XOR2_X1 U24689 ( .A1(n38323), .A2(n39384), .Z(n5039) );
  NAND4_X2 U24691 ( .A1(n12066), .A2(n12010), .A3(n12065), .A4(n8050), .ZN(
        n37288) );
  AOI21_X2 U24692 ( .A1(n16966), .A2(n16965), .B(n44487), .ZN(n49901) );
  NOR2_X2 U24693 ( .A1(n5042), .A2(n13445), .ZN(n16966) );
  INV_X1 U24701 ( .I(n47039), .ZN(n10572) );
  XOR2_X1 U24703 ( .A1(n12315), .A2(n735), .Z(n5048) );
  INV_X4 U24707 ( .I(n36951), .ZN(n34914) );
  NAND2_X2 U24708 ( .A1(n57426), .A2(n5050), .ZN(n47812) );
  INV_X2 U24715 ( .I(n25171), .ZN(n5054) );
  INV_X2 U24720 ( .I(n5318), .ZN(n5711) );
  INV_X2 U24721 ( .I(n8553), .ZN(n6512) );
  INV_X2 U24729 ( .I(n12755), .ZN(n18726) );
  NOR2_X1 U24730 ( .A1(n24946), .A2(n26964), .ZN(n5069) );
  NAND2_X1 U24741 ( .A1(n5368), .A2(n1501), .ZN(n24684) );
  NAND2_X1 U24742 ( .A1(n41721), .A2(n5368), .ZN(n11497) );
  XOR2_X1 U24743 ( .A1(n17624), .A2(n33258), .Z(n31977) );
  XOR2_X1 U24744 ( .A1(n20621), .A2(n52226), .Z(n5080) );
  NAND2_X2 U24747 ( .A1(n31659), .A2(n1542), .ZN(n25509) );
  INV_X2 U24748 ( .I(n30421), .ZN(n31076) );
  NAND2_X2 U24750 ( .A1(n25644), .A2(n26973), .ZN(n9153) );
  XOR2_X1 U24754 ( .A1(n31851), .A2(n5089), .Z(n18782) );
  INV_X1 U24755 ( .I(n27011), .ZN(n5092) );
  INV_X1 U24757 ( .I(n8342), .ZN(n23957) );
  XOR2_X1 U24759 ( .A1(n46577), .A2(n46380), .Z(n13938) );
  NOR2_X1 U24770 ( .A1(n30492), .A2(n9411), .ZN(n27759) );
  AND2_X1 U24773 ( .A1(n5124), .A2(n24735), .Z(n5117) );
  NAND2_X2 U24774 ( .A1(n9017), .A2(n1894), .ZN(n24735) );
  XOR2_X1 U24776 ( .A1(n23587), .A2(n46430), .Z(n8158) );
  XOR2_X1 U24777 ( .A1(n5118), .A2(n46634), .Z(n46635) );
  XOR2_X1 U24778 ( .A1(n4990), .A2(n5118), .Z(n43673) );
  XOR2_X1 U24779 ( .A1(n5360), .A2(n5118), .Z(n10664) );
  INV_X2 U24780 ( .I(n5120), .ZN(n11912) );
  AOI22_X1 U24785 ( .A1(n5122), .A2(n55878), .B1(n55837), .B2(n60092), .ZN(
        n55838) );
  NOR2_X2 U24786 ( .A1(n17774), .A2(n55893), .ZN(n5122) );
  AOI22_X1 U24787 ( .A1(n28352), .A2(n28351), .B1(n28350), .B2(n5124), .ZN(
        n28353) );
  NOR2_X2 U24789 ( .A1(n21166), .A2(n21168), .ZN(n5125) );
  XOR2_X1 U24790 ( .A1(n25005), .A2(n22241), .Z(n5127) );
  XOR2_X1 U24791 ( .A1(n17801), .A2(n63003), .Z(n22241) );
  XOR2_X1 U24792 ( .A1(n5665), .A2(n24368), .Z(n25005) );
  INV_X2 U24796 ( .I(n22739), .ZN(n41020) );
  NAND2_X2 U24797 ( .A1(n9543), .A2(n26686), .ZN(n23569) );
  OR2_X1 U24798 ( .A1(n34628), .A2(n22226), .Z(n5134) );
  NOR2_X1 U24800 ( .A1(n61735), .A2(n22128), .ZN(n6721) );
  XOR2_X1 U24801 ( .A1(n31734), .A2(n15489), .Z(n5139) );
  XOR2_X1 U24802 ( .A1(n11470), .A2(n5142), .Z(n11469) );
  XOR2_X1 U24803 ( .A1(n5144), .A2(n5143), .Z(n5142) );
  XOR2_X1 U24804 ( .A1(n22332), .A2(n51580), .Z(n5144) );
  NOR2_X1 U24805 ( .A1(n47838), .A2(n5145), .ZN(n42618) );
  NOR2_X1 U24806 ( .A1(n22537), .A2(n5145), .ZN(n45215) );
  AOI21_X1 U24808 ( .A1(n59695), .A2(n15157), .B(n5145), .ZN(n17135) );
  OAI21_X2 U24815 ( .A1(n5150), .A2(n25326), .B(n5149), .ZN(n14755) );
  NOR2_X1 U24820 ( .A1(n27224), .A2(n5153), .ZN(n26971) );
  NAND2_X2 U24822 ( .A1(n26446), .A2(n1445), .ZN(n5218) );
  XNOR2_X1 U24823 ( .A1(n46547), .A2(n25926), .ZN(n9150) );
  NAND3_X1 U24827 ( .A1(n22674), .A2(n12878), .A3(n28908), .ZN(n5156) );
  NAND2_X1 U24829 ( .A1(n47798), .A2(n47800), .ZN(n6192) );
  NAND2_X1 U24830 ( .A1(n1312), .A2(n58702), .ZN(n34597) );
  INV_X2 U24831 ( .I(n11192), .ZN(n5349) );
  XOR2_X1 U24833 ( .A1(n5166), .A2(n15096), .Z(n5165) );
  XOR2_X1 U24834 ( .A1(n23552), .A2(n15505), .Z(n5166) );
  NAND2_X2 U24835 ( .A1(n46011), .A2(n20622), .ZN(n15505) );
  INV_X4 U24836 ( .I(n732), .ZN(n17148) );
  NAND2_X1 U24837 ( .A1(n22797), .A2(n732), .ZN(n34240) );
  INV_X2 U24841 ( .I(n9437), .ZN(n48612) );
  XOR2_X1 U24842 ( .A1(n46272), .A2(n46281), .Z(n5170) );
  NOR2_X1 U24843 ( .A1(n43219), .A2(n5171), .ZN(n8678) );
  NAND2_X2 U24845 ( .A1(n52124), .A2(n50931), .ZN(n52120) );
  XOR2_X1 U24848 ( .A1(n31748), .A2(n6744), .Z(n6275) );
  XOR2_X1 U24849 ( .A1(n64035), .A2(n6744), .Z(n12814) );
  XOR2_X1 U24851 ( .A1(n5180), .A2(n46673), .Z(n46676) );
  XOR2_X1 U24853 ( .A1(n8539), .A2(n5182), .Z(n5181) );
  XOR2_X1 U24854 ( .A1(n38977), .A2(n38975), .Z(n5182) );
  XOR2_X1 U24855 ( .A1(n306), .A2(n38976), .Z(n5184) );
  INV_X2 U24856 ( .I(n12974), .ZN(n7055) );
  XOR2_X1 U24857 ( .A1(n5458), .A2(n17129), .Z(n37633) );
  NOR2_X2 U24859 ( .A1(n35031), .A2(n15756), .ZN(n34646) );
  INV_X4 U24868 ( .I(n54901), .ZN(n54904) );
  NAND2_X2 U24869 ( .A1(n15798), .A2(n16149), .ZN(n54901) );
  AOI21_X1 U24873 ( .A1(n29303), .A2(n26965), .B(n5206), .ZN(n26963) );
  NAND2_X1 U24878 ( .A1(n5218), .A2(n29297), .ZN(n26688) );
  NAND2_X1 U24879 ( .A1(n5218), .A2(n29296), .ZN(n26445) );
  NOR2_X2 U24881 ( .A1(n44408), .A2(n5219), .ZN(n48036) );
  NAND2_X2 U24882 ( .A1(n48323), .A2(n49014), .ZN(n5219) );
  XOR2_X1 U24888 ( .A1(n7699), .A2(n5223), .Z(n5222) );
  XOR2_X1 U24890 ( .A1(n9079), .A2(n44142), .Z(n5223) );
  OAI22_X1 U24892 ( .A1(n44782), .A2(n46905), .B1(n5225), .B2(n44783), .ZN(
        n44785) );
  NAND2_X1 U24893 ( .A1(n5225), .A2(n1070), .ZN(n17033) );
  NAND2_X1 U24894 ( .A1(n5225), .A2(n23480), .ZN(n45511) );
  INV_X2 U24896 ( .I(n5228), .ZN(n31470) );
  XNOR2_X1 U24900 ( .A1(n5231), .A2(n25034), .ZN(n5228) );
  XOR2_X1 U24901 ( .A1(n59274), .A2(n5232), .Z(n25034) );
  XOR2_X1 U24902 ( .A1(n21369), .A2(n5744), .Z(n5232) );
  XOR2_X1 U24905 ( .A1(n10599), .A2(n46348), .Z(n5234) );
  NOR2_X1 U24908 ( .A1(n64121), .A2(n5235), .ZN(n14366) );
  NAND2_X2 U24910 ( .A1(n25148), .A2(n20091), .ZN(n5235) );
  NOR2_X1 U24912 ( .A1(n22977), .A2(n5236), .ZN(n5672) );
  NAND3_X1 U24914 ( .A1(n52218), .A2(n9111), .A3(n58373), .ZN(n12304) );
  NAND2_X2 U24917 ( .A1(n20738), .A2(n55656), .ZN(n5236) );
  NAND2_X1 U24918 ( .A1(n64155), .A2(n28400), .ZN(n28402) );
  OR2_X1 U24919 ( .A1(n42341), .A2(n43582), .Z(n5238) );
  XOR2_X1 U24922 ( .A1(n5266), .A2(n17042), .Z(n6331) );
  XOR2_X1 U24924 ( .A1(n9530), .A2(n44826), .Z(n5245) );
  NAND2_X1 U24926 ( .A1(n20110), .A2(n5246), .ZN(n20109) );
  NAND2_X1 U24927 ( .A1(n46827), .A2(n5246), .ZN(n46828) );
  XOR2_X1 U24928 ( .A1(n32574), .A2(n33848), .Z(n12663) );
  XOR2_X1 U24929 ( .A1(n33848), .A2(n829), .Z(n31698) );
  XOR2_X1 U24931 ( .A1(n31329), .A2(n33848), .Z(n16273) );
  INV_X2 U24934 ( .I(n5251), .ZN(n22477) );
  XNOR2_X1 U24937 ( .A1(n24108), .A2(n5252), .ZN(n5251) );
  XOR2_X1 U24940 ( .A1(n2801), .A2(n51505), .Z(n17803) );
  XOR2_X1 U24941 ( .A1(n19323), .A2(n2801), .Z(n19357) );
  OR2_X2 U24943 ( .A1(n24301), .A2(n5263), .Z(n55415) );
  NOR2_X1 U24946 ( .A1(n22598), .A2(n12768), .ZN(n31713) );
  NAND2_X1 U24947 ( .A1(n34143), .A2(n12768), .ZN(n6923) );
  XOR2_X1 U24951 ( .A1(n39207), .A2(n22), .Z(n7212) );
  NAND4_X2 U24952 ( .A1(n16606), .A2(n13303), .A3(n16605), .A4(n16604), .ZN(
        n21130) );
  NOR2_X2 U24959 ( .A1(n37529), .A2(n1409), .ZN(n22738) );
  XOR2_X1 U24961 ( .A1(n64454), .A2(n4156), .Z(n52468) );
  XOR2_X1 U24962 ( .A1(n8273), .A2(n4156), .Z(n51851) );
  XOR2_X1 U24963 ( .A1(n51943), .A2(n4156), .Z(n52497) );
  XOR2_X1 U24964 ( .A1(n50452), .A2(n4156), .Z(n50884) );
  XOR2_X1 U24965 ( .A1(n12603), .A2(n4156), .Z(n51274) );
  NOR2_X1 U24969 ( .A1(n28608), .A2(n4869), .ZN(n13013) );
  NAND2_X1 U24971 ( .A1(n19634), .A2(n1632), .ZN(n50443) );
  NAND2_X2 U24974 ( .A1(n5283), .A2(n62334), .ZN(n17818) );
  NAND2_X1 U24978 ( .A1(n5285), .A2(n30374), .ZN(n27724) );
  NAND2_X1 U24979 ( .A1(n5285), .A2(n30375), .ZN(n30368) );
  NOR2_X1 U24980 ( .A1(n5285), .A2(n1316), .ZN(n20187) );
  AOI22_X1 U24981 ( .A1(n20606), .A2(n29482), .B1(n8583), .B2(n5285), .ZN(
        n29484) );
  INV_X2 U24987 ( .I(n5293), .ZN(n23634) );
  NAND2_X2 U24990 ( .A1(n45075), .A2(n21241), .ZN(n46919) );
  XOR2_X1 U24991 ( .A1(n6342), .A2(n45014), .Z(n45016) );
  AOI21_X1 U24993 ( .A1(n32835), .A2(n33992), .B(n1539), .ZN(n32838) );
  INV_X1 U24996 ( .I(n47808), .ZN(n5307) );
  NOR2_X2 U24997 ( .A1(n5310), .A2(n5309), .ZN(n5308) );
  NAND2_X2 U24998 ( .A1(n47816), .A2(n5311), .ZN(n5310) );
  INV_X1 U24999 ( .I(n44385), .ZN(n41553) );
  XNOR2_X1 U25000 ( .A1(n6342), .A2(n44385), .ZN(n43408) );
  INV_X1 U25001 ( .I(n41602), .ZN(n5316) );
  XOR2_X1 U25004 ( .A1(n37735), .A2(n37299), .Z(n37302) );
  NAND2_X1 U25006 ( .A1(n5319), .A2(n41898), .ZN(n41901) );
  NAND2_X1 U25007 ( .A1(n41894), .A2(n5319), .ZN(n41897) );
  NOR2_X1 U25008 ( .A1(n24644), .A2(n5319), .ZN(n5508) );
  NOR2_X2 U25013 ( .A1(n23170), .A2(n27996), .ZN(n29107) );
  XOR2_X1 U25015 ( .A1(n3389), .A2(n21884), .Z(n22787) );
  INV_X2 U25018 ( .I(n36220), .ZN(n36442) );
  NAND2_X2 U25019 ( .A1(n24539), .A2(n24538), .ZN(n36220) );
  NAND2_X2 U25020 ( .A1(n10983), .A2(n15804), .ZN(n52222) );
  NAND2_X2 U25022 ( .A1(n12282), .A2(n56234), .ZN(n56557) );
  XOR2_X1 U25025 ( .A1(n12084), .A2(n5333), .Z(n5332) );
  NAND2_X2 U25027 ( .A1(n23354), .A2(n32222), .ZN(n34736) );
  NOR2_X2 U25028 ( .A1(n34752), .A2(n31976), .ZN(n32222) );
  INV_X1 U25034 ( .I(n43571), .ZN(n5341) );
  XOR2_X1 U25035 ( .A1(n32278), .A2(n5342), .Z(n15416) );
  XOR2_X1 U25036 ( .A1(n742), .A2(n5342), .Z(n32356) );
  XOR2_X1 U25037 ( .A1(n21332), .A2(n5342), .Z(n31893) );
  XOR2_X1 U25038 ( .A1(n30573), .A2(n5342), .Z(n30598) );
  NAND2_X1 U25040 ( .A1(n30393), .A2(n2795), .ZN(n5343) );
  NAND2_X2 U25041 ( .A1(n45189), .A2(n45190), .ZN(n5945) );
  MUX2_X1 U25042 ( .I0(n30364), .I1(n29060), .S(n1558), .Z(n28296) );
  XOR2_X1 U25045 ( .A1(n5349), .A2(n6224), .Z(n51528) );
  XOR2_X1 U25048 ( .A1(n5353), .A2(n12283), .Z(n5352) );
  NAND2_X2 U25050 ( .A1(n1442), .A2(n11617), .ZN(n12070) );
  AOI21_X1 U25054 ( .A1(n40982), .A2(n6768), .B(n5362), .ZN(n40984) );
  XOR2_X1 U25057 ( .A1(n16404), .A2(n5363), .Z(n38116) );
  XOR2_X1 U25060 ( .A1(n5371), .A2(n28259), .Z(n27028) );
  NOR2_X2 U25061 ( .A1(n28254), .A2(n5371), .ZN(n29173) );
  XOR2_X1 U25065 ( .A1(n38232), .A2(n38322), .Z(n5374) );
  XOR2_X1 U25066 ( .A1(n17512), .A2(n16404), .Z(n38322) );
  XOR2_X1 U25076 ( .A1(n14847), .A2(n13153), .Z(n32370) );
  INV_X2 U25077 ( .I(n36031), .ZN(n35388) );
  NAND2_X2 U25078 ( .A1(n8474), .A2(n4802), .ZN(n36031) );
  NAND2_X1 U25087 ( .A1(n7016), .A2(n5389), .ZN(n31775) );
  XOR2_X1 U25089 ( .A1(n52453), .A2(n51394), .Z(n5390) );
  NAND2_X2 U25090 ( .A1(n24683), .A2(n11594), .ZN(n52453) );
  NOR2_X2 U25091 ( .A1(n12410), .A2(n40996), .ZN(n40217) );
  XOR2_X1 U25093 ( .A1(n8599), .A2(n24401), .Z(n8419) );
  NAND2_X1 U25094 ( .A1(n5396), .A2(n24613), .ZN(n10025) );
  NAND2_X2 U25095 ( .A1(n4888), .A2(n49465), .ZN(n24613) );
  AND2_X1 U25100 ( .A1(n41117), .A2(n41115), .Z(n5400) );
  OAI21_X2 U25101 ( .A1(n5402), .A2(n30229), .B(n5401), .ZN(n32230) );
  XOR2_X1 U25105 ( .A1(n51590), .A2(n11507), .Z(n5404) );
  XOR2_X1 U25107 ( .A1(n62455), .A2(n52436), .Z(n5405) );
  NOR2_X2 U25109 ( .A1(n45199), .A2(n11417), .ZN(n8047) );
  XOR2_X1 U25110 ( .A1(n5824), .A2(n17517), .Z(n8170) );
  XOR2_X1 U25111 ( .A1(n15075), .A2(n5408), .Z(n5824) );
  INV_X4 U25117 ( .I(n11424), .ZN(n16971) );
  INV_X2 U25118 ( .I(n13204), .ZN(n15727) );
  INV_X2 U25120 ( .I(n5417), .ZN(n9883) );
  OAI21_X1 U25122 ( .A1(n22473), .A2(n56256), .B(n51888), .ZN(n5418) );
  NOR2_X2 U25125 ( .A1(n49367), .A2(n49671), .ZN(n48007) );
  XOR2_X1 U25126 ( .A1(n5432), .A2(n44501), .Z(n46201) );
  XOR2_X1 U25127 ( .A1(n10678), .A2(n57586), .Z(n5432) );
  XOR2_X1 U25130 ( .A1(n24292), .A2(n31314), .Z(n5433) );
  XOR2_X1 U25131 ( .A1(n5435), .A2(n11930), .Z(n5434) );
  XOR2_X1 U25132 ( .A1(n38587), .A2(n5439), .Z(n5438) );
  XOR2_X1 U25133 ( .A1(n36993), .A2(n36992), .Z(n5439) );
  NOR2_X1 U25136 ( .A1(n37329), .A2(n5442), .ZN(n32153) );
  NOR2_X1 U25137 ( .A1(n37333), .A2(n5442), .ZN(n32150) );
  NOR2_X1 U25138 ( .A1(n17537), .A2(n5442), .ZN(n12176) );
  OAI22_X1 U25139 ( .A1(n37325), .A2(n5442), .B1(n37326), .B2(n17444), .ZN(
        n37332) );
  NOR2_X2 U25142 ( .A1(n56817), .A2(n56757), .ZN(n56788) );
  NOR2_X1 U25143 ( .A1(n56815), .A2(n5447), .ZN(n5446) );
  NAND2_X1 U25144 ( .A1(n56816), .A2(n56817), .ZN(n5447) );
  XOR2_X1 U25146 ( .A1(n10619), .A2(n8480), .Z(n5449) );
  XOR2_X1 U25147 ( .A1(n5450), .A2(n22199), .Z(n11372) );
  XOR2_X1 U25148 ( .A1(n5451), .A2(n5452), .Z(n5450) );
  XOR2_X1 U25149 ( .A1(n41741), .A2(n41742), .Z(n5452) );
  INV_X2 U25150 ( .I(n5457), .ZN(n20446) );
  NAND2_X2 U25152 ( .A1(n5459), .A2(n25688), .ZN(n23637) );
  NOR2_X1 U25158 ( .A1(n49674), .A2(n5463), .ZN(n48709) );
  NAND2_X2 U25161 ( .A1(n5469), .A2(n5467), .ZN(n30649) );
  NOR2_X1 U25163 ( .A1(n10769), .A2(n58020), .ZN(n35330) );
  NAND2_X1 U25164 ( .A1(n35769), .A2(n58020), .ZN(n33926) );
  OAI21_X1 U25165 ( .A1(n60152), .A2(n58020), .B(n34422), .ZN(n34330) );
  OAI22_X1 U25166 ( .A1(n22835), .A2(n58020), .B1(n58231), .B2(n35777), .ZN(
        n34420) );
  AND2_X1 U25167 ( .A1(n38425), .A2(n38426), .Z(n5475) );
  NAND2_X1 U25168 ( .A1(n5773), .A2(n1718), .ZN(n42918) );
  OAI21_X1 U25169 ( .A1(n5324), .A2(n5476), .B(n54410), .ZN(n54412) );
  NOR2_X2 U25172 ( .A1(n13068), .A2(n25999), .ZN(n5477) );
  NAND2_X2 U25173 ( .A1(n24300), .A2(n12171), .ZN(n18700) );
  OAI22_X1 U25178 ( .A1(n28987), .A2(n20025), .B1(n30021), .B2(n30020), .ZN(
        n5491) );
  AND3_X1 U25184 ( .A1(n40583), .A2(n40802), .A3(n40582), .Z(n5512) );
  INV_X2 U25186 ( .I(n10353), .ZN(n5517) );
  INV_X2 U25187 ( .I(n34632), .ZN(n35047) );
  XOR2_X1 U25188 ( .A1(n5520), .A2(n14292), .Z(n14294) );
  OAI21_X1 U25194 ( .A1(n12653), .A2(n36628), .B(n36627), .ZN(n5527) );
  NAND2_X2 U25203 ( .A1(n1419), .A2(n7705), .ZN(n35591) );
  XOR2_X1 U25205 ( .A1(n23440), .A2(n63941), .Z(n44954) );
  INV_X2 U25207 ( .I(n5533), .ZN(n6082) );
  NOR2_X2 U25208 ( .A1(n45768), .A2(n6082), .ZN(n6081) );
  NAND2_X1 U25212 ( .A1(n4496), .A2(n35691), .ZN(n32764) );
  OAI21_X1 U25213 ( .A1(n4496), .A2(n22723), .B(n35691), .ZN(n33014) );
  OAI22_X1 U25224 ( .A1(n27106), .A2(n22234), .B1(n23917), .B2(n5548), .ZN(
        n27107) );
  NAND2_X1 U25227 ( .A1(n55659), .A2(n5550), .ZN(n55661) );
  NAND2_X1 U25233 ( .A1(n5553), .A2(n55639), .ZN(n5552) );
  NAND3_X2 U25236 ( .A1(n35854), .A2(n5557), .A3(n5556), .ZN(n14798) );
  AND2_X1 U25239 ( .A1(n37221), .A2(n36264), .Z(n5561) );
  OAI22_X1 U25241 ( .A1(n5565), .A2(n62600), .B1(n43573), .B2(n43577), .ZN(
        n5564) );
  XOR2_X1 U25242 ( .A1(n1391), .A2(n5398), .Z(n5565) );
  XOR2_X1 U25243 ( .A1(n2748), .A2(n45253), .Z(n45254) );
  XOR2_X1 U25244 ( .A1(n44252), .A2(n2748), .Z(n41659) );
  INV_X1 U25245 ( .I(n35747), .ZN(n10900) );
  INV_X4 U25247 ( .I(n5571), .ZN(n43995) );
  XOR2_X1 U25250 ( .A1(n5574), .A2(n5573), .Z(n5572) );
  XOR2_X1 U25251 ( .A1(n16700), .A2(n1390), .Z(n44387) );
  XOR2_X1 U25256 ( .A1(n14798), .A2(n38648), .Z(n16450) );
  XOR2_X1 U25257 ( .A1(n16706), .A2(n54249), .Z(n31850) );
  NAND2_X1 U25258 ( .A1(n49750), .A2(n49749), .ZN(n5578) );
  NOR2_X1 U25259 ( .A1(n5581), .A2(n40804), .ZN(n40807) );
  NAND4_X1 U25260 ( .A1(n41895), .A2(n41897), .A3(n5581), .A4(n41896), .ZN(
        n41903) );
  INV_X2 U25268 ( .I(n5586), .ZN(n22508) );
  NAND2_X2 U25269 ( .A1(n22508), .A2(n17464), .ZN(n47700) );
  AOI21_X1 U25273 ( .A1(n19042), .A2(n15724), .B(n4724), .ZN(n49303) );
  INV_X1 U25275 ( .I(Key[83]), .ZN(n5593) );
  XOR2_X1 U25276 ( .A1(n5593), .A2(Ciphertext[178]), .Z(n5935) );
  INV_X2 U25278 ( .I(n14324), .ZN(n11524) );
  NAND2_X2 U25279 ( .A1(n15804), .A2(n56268), .ZN(n56264) );
  INV_X2 U25281 ( .I(n11310), .ZN(n37874) );
  XOR2_X1 U25283 ( .A1(n25721), .A2(n5596), .Z(n5595) );
  XOR2_X1 U25284 ( .A1(n5597), .A2(n38578), .Z(n5596) );
  XOR2_X1 U25285 ( .A1(n23931), .A2(n37872), .Z(n5597) );
  XOR2_X1 U25290 ( .A1(n52335), .A2(n5603), .Z(n9619) );
  XOR2_X1 U25292 ( .A1(n16984), .A2(n5603), .Z(n50847) );
  XOR2_X1 U25293 ( .A1(n22783), .A2(n5603), .Z(n51177) );
  XOR2_X1 U25294 ( .A1(n51483), .A2(n5603), .Z(n51484) );
  XOR2_X1 U25295 ( .A1(n5603), .A2(n20332), .Z(n50730) );
  INV_X2 U25300 ( .I(n5622), .ZN(n32295) );
  XOR2_X1 U25306 ( .A1(n5626), .A2(n50497), .Z(n5694) );
  XOR2_X1 U25307 ( .A1(n5626), .A2(n50721), .Z(n50722) );
  XOR2_X1 U25308 ( .A1(n58834), .A2(n51494), .Z(n51293) );
  XOR2_X1 U25309 ( .A1(n1197), .A2(n62084), .Z(n14441) );
  NAND2_X1 U25310 ( .A1(n28221), .A2(n27366), .ZN(n5627) );
  NOR2_X2 U25316 ( .A1(n5631), .A2(n64950), .ZN(n14944) );
  NOR2_X2 U25318 ( .A1(n21791), .A2(n1739), .ZN(n41220) );
  NAND4_X2 U25320 ( .A1(n5633), .A2(n11621), .A3(n24826), .A4(n5632), .ZN(
        n33856) );
  XOR2_X1 U25321 ( .A1(Ciphertext[64]), .A2(Key[53]), .Z(n5716) );
  XOR2_X1 U25323 ( .A1(n38466), .A2(n21462), .Z(n5638) );
  XOR2_X1 U25324 ( .A1(n13620), .A2(n5640), .Z(n5639) );
  XOR2_X1 U25326 ( .A1(n13619), .A2(n13618), .Z(n13620) );
  AOI21_X1 U25327 ( .A1(n5641), .A2(n33788), .B(n59261), .ZN(n13342) );
  NAND3_X1 U25328 ( .A1(n5646), .A2(n5644), .A3(n5643), .ZN(Plaintext[53]) );
  NAND2_X1 U25329 ( .A1(n5650), .A2(n1901), .ZN(n5643) );
  NAND2_X1 U25330 ( .A1(n54014), .A2(n61695), .ZN(n5645) );
  NAND4_X1 U25331 ( .A1(n5647), .A2(n61695), .A3(n54014), .A4(n24061), .ZN(
        n5646) );
  AND2_X1 U25332 ( .A1(n53903), .A2(n53902), .Z(n5649) );
  NAND2_X1 U25334 ( .A1(n12915), .A2(n54001), .ZN(n5651) );
  XOR2_X1 U25335 ( .A1(n23525), .A2(n32406), .Z(n13213) );
  XOR2_X1 U25336 ( .A1(n63892), .A2(n5652), .Z(n32406) );
  NAND2_X2 U25337 ( .A1(n6151), .A2(n6150), .ZN(n25106) );
  XOR2_X1 U25338 ( .A1(n22161), .A2(n22162), .Z(n5652) );
  NAND2_X1 U25341 ( .A1(n24111), .A2(n5656), .ZN(n53868) );
  NAND2_X1 U25342 ( .A1(n53868), .A2(n54108), .ZN(n53869) );
  NAND2_X1 U25345 ( .A1(n56867), .A2(n5658), .ZN(n56862) );
  NAND3_X1 U25347 ( .A1(n56837), .A2(n56885), .A3(n5658), .ZN(n52726) );
  OAI22_X1 U25348 ( .A1(n56841), .A2(n56853), .B1(n56845), .B2(n5658), .ZN(
        n17650) );
  AOI21_X1 U25349 ( .A1(n5659), .A2(n28195), .B(n57781), .ZN(n27339) );
  NOR2_X1 U25350 ( .A1(n20126), .A2(n5659), .ZN(n28662) );
  XOR2_X1 U25351 ( .A1(n5660), .A2(n38524), .Z(n23907) );
  OAI21_X1 U25353 ( .A1(n5661), .A2(n48825), .B(n59808), .ZN(n48826) );
  XOR2_X1 U25356 ( .A1(n7136), .A2(n1077), .Z(n5664) );
  XOR2_X1 U25357 ( .A1(n14648), .A2(n5666), .Z(n5665) );
  NAND2_X2 U25359 ( .A1(n25558), .A2(n25561), .ZN(n51504) );
  NOR2_X2 U25360 ( .A1(n60077), .A2(n17382), .ZN(n23610) );
  XOR2_X1 U25363 ( .A1(n5682), .A2(n7302), .Z(n5969) );
  XOR2_X1 U25364 ( .A1(n11884), .A2(n53705), .Z(n5682) );
  NAND4_X2 U25365 ( .A1(n6020), .A2(n6021), .A3(n6022), .A4(n20592), .ZN(
        n11884) );
  XNOR2_X1 U25367 ( .A1(n15066), .A2(n16389), .ZN(n26035) );
  NAND2_X2 U25368 ( .A1(n15065), .A2(n15067), .ZN(n15066) );
  XOR2_X1 U25371 ( .A1(n6744), .A2(n29885), .Z(n5685) );
  INV_X1 U25377 ( .I(n5705), .ZN(n21953) );
  NOR2_X1 U25378 ( .A1(n48529), .A2(n5705), .ZN(n25954) );
  XOR2_X1 U25382 ( .A1(n31675), .A2(n5155), .Z(n30597) );
  OR2_X1 U25385 ( .A1(n8026), .A2(n40661), .Z(n5707) );
  INV_X1 U25387 ( .I(n43226), .ZN(n42995) );
  XOR2_X1 U25390 ( .A1(n5710), .A2(n23497), .Z(n9072) );
  XOR2_X1 U25391 ( .A1(n1331), .A2(n44147), .Z(n5710) );
  XOR2_X1 U25393 ( .A1(n5712), .A2(n44431), .Z(n44432) );
  XOR2_X1 U25394 ( .A1(n21142), .A2(n62569), .Z(n9855) );
  XOR2_X1 U25395 ( .A1(n5712), .A2(n25530), .Z(n15056) );
  XOR2_X1 U25396 ( .A1(n13959), .A2(n5712), .Z(n13958) );
  NAND3_X1 U25399 ( .A1(n5713), .A2(n48957), .A3(n49177), .ZN(n10873) );
  NOR2_X1 U25400 ( .A1(n5714), .A2(n6896), .ZN(n49185) );
  NOR3_X1 U25401 ( .A1(n23151), .A2(n60843), .A3(n15044), .ZN(n5715) );
  NOR2_X2 U25402 ( .A1(n21240), .A2(n43874), .ZN(n6144) );
  XOR2_X1 U25406 ( .A1(n8625), .A2(n31429), .Z(n31430) );
  INV_X2 U25408 ( .I(n5716), .ZN(n28221) );
  AND2_X1 U25409 ( .A1(n42411), .A2(n42072), .Z(n5720) );
  NOR2_X1 U25411 ( .A1(n46944), .A2(n60038), .ZN(n47986) );
  NAND2_X1 U25412 ( .A1(n5722), .A2(n59922), .ZN(n5721) );
  INV_X1 U25413 ( .I(n9512), .ZN(n5722) );
  XOR2_X1 U25415 ( .A1(n5725), .A2(n50967), .Z(n5724) );
  XOR2_X1 U25417 ( .A1(n1831), .A2(n5727), .Z(n24348) );
  XOR2_X1 U25418 ( .A1(n24677), .A2(n1573), .Z(n5730) );
  NAND2_X2 U25419 ( .A1(n16638), .A2(n16637), .ZN(n24677) );
  NAND2_X1 U25422 ( .A1(n5734), .A2(n1416), .ZN(n8664) );
  NOR2_X2 U25424 ( .A1(n61443), .A2(n54074), .ZN(n54471) );
  NAND2_X2 U25428 ( .A1(n19342), .A2(n43101), .ZN(n44455) );
  INV_X2 U25433 ( .I(n5743), .ZN(n49266) );
  NAND2_X1 U25434 ( .A1(n48957), .A2(n4647), .ZN(n10070) );
  XOR2_X1 U25435 ( .A1(n5745), .A2(n25034), .Z(n13950) );
  XOR2_X1 U25436 ( .A1(n33178), .A2(n4795), .Z(n5744) );
  XOR2_X1 U25439 ( .A1(n16936), .A2(n11930), .Z(n33190) );
  XOR2_X1 U25441 ( .A1(n5748), .A2(n43594), .Z(n43595) );
  XOR2_X1 U25443 ( .A1(n19348), .A2(n9179), .Z(n5749) );
  XOR2_X1 U25446 ( .A1(n5752), .A2(n9759), .Z(n14337) );
  XOR2_X1 U25447 ( .A1(n32495), .A2(n21094), .Z(n5752) );
  XOR2_X1 U25449 ( .A1(n32570), .A2(n25822), .Z(n5754) );
  INV_X1 U25451 ( .I(n35457), .ZN(n5758) );
  NAND2_X2 U25453 ( .A1(n5757), .A2(n35461), .ZN(n6441) );
  INV_X2 U25460 ( .I(n5766), .ZN(n45333) );
  INV_X2 U25462 ( .I(n14427), .ZN(n5767) );
  NOR2_X1 U25463 ( .A1(n27648), .A2(n27649), .ZN(n5770) );
  INV_X2 U25466 ( .I(n11980), .ZN(n13770) );
  OR2_X2 U25469 ( .A1(n9711), .A2(n5774), .Z(n40663) );
  NAND2_X2 U25471 ( .A1(n25427), .A2(n25428), .ZN(n33623) );
  AOI22_X1 U25473 ( .A1(n54611), .A2(n5777), .B1(n54431), .B2(n54436), .ZN(
        n52382) );
  INV_X2 U25475 ( .I(n7991), .ZN(n5778) );
  XOR2_X1 U25476 ( .A1(n5781), .A2(n5782), .Z(n5780) );
  XOR2_X1 U25477 ( .A1(n4563), .A2(n2905), .Z(n5781) );
  XOR2_X1 U25478 ( .A1(n16476), .A2(n61651), .Z(n5782) );
  XOR2_X1 U25481 ( .A1(n37697), .A2(n24189), .Z(n39768) );
  XOR2_X1 U25483 ( .A1(n5786), .A2(n37702), .Z(n38619) );
  NAND4_X1 U25484 ( .A1(n38274), .A2(n42237), .A3(n22290), .A4(n41942), .ZN(
        n5790) );
  NAND2_X1 U25486 ( .A1(n37336), .A2(n37182), .ZN(n22552) );
  XOR2_X1 U25490 ( .A1(n45399), .A2(n5811), .Z(n5810) );
  XOR2_X1 U25491 ( .A1(n45325), .A2(n45324), .Z(n5811) );
  XOR2_X1 U25492 ( .A1(n11074), .A2(n54143), .Z(n45399) );
  XOR2_X1 U25493 ( .A1(n11529), .A2(n33891), .Z(n5818) );
  XOR2_X1 U25494 ( .A1(n31911), .A2(n32181), .Z(n5819) );
  XOR2_X1 U25498 ( .A1(n3480), .A2(n52575), .Z(n38175) );
  NAND3_X2 U25500 ( .A1(n5826), .A2(n5825), .A3(n43055), .ZN(n44592) );
  XOR2_X1 U25501 ( .A1(n5830), .A2(n5828), .Z(n13857) );
  XOR2_X1 U25502 ( .A1(n5829), .A2(n33059), .Z(n5828) );
  XOR2_X1 U25503 ( .A1(n32129), .A2(n19388), .Z(n33059) );
  XOR2_X1 U25504 ( .A1(n60902), .A2(n32130), .Z(n5829) );
  XOR2_X1 U25505 ( .A1(n61152), .A2(n32393), .Z(n32130) );
  XOR2_X1 U25509 ( .A1(n6324), .A2(n44606), .Z(n5834) );
  INV_X2 U25511 ( .I(n5836), .ZN(n39241) );
  INV_X2 U25514 ( .I(n18473), .ZN(n5837) );
  NOR2_X1 U25515 ( .A1(n16244), .A2(n21517), .ZN(n17301) );
  XOR2_X1 U25517 ( .A1(n23089), .A2(n10043), .Z(n46395) );
  NAND3_X2 U25519 ( .A1(n41976), .A2(n41977), .A3(n22951), .ZN(n46224) );
  XOR2_X1 U25522 ( .A1(n39222), .A2(n39223), .Z(n5841) );
  XOR2_X1 U25523 ( .A1(n5842), .A2(n37998), .Z(n39224) );
  XOR2_X1 U25524 ( .A1(n38856), .A2(n51019), .Z(n5842) );
  NAND2_X2 U25530 ( .A1(n12878), .A2(n28908), .ZN(n25176) );
  XOR2_X1 U25531 ( .A1(n38131), .A2(n38130), .Z(n5867) );
  XOR2_X1 U25532 ( .A1(n38160), .A2(n38877), .Z(n38131) );
  NAND2_X2 U25534 ( .A1(n5870), .A2(n5869), .ZN(n20351) );
  NAND2_X2 U25535 ( .A1(n43486), .A2(n43487), .ZN(n43778) );
  NAND2_X2 U25536 ( .A1(n24750), .A2(n20006), .ZN(n21073) );
  INV_X1 U25538 ( .I(n49744), .ZN(n5883) );
  XOR2_X1 U25545 ( .A1(n44377), .A2(n46354), .Z(n5899) );
  INV_X1 U25547 ( .I(n5900), .ZN(n36363) );
  OAI22_X1 U25549 ( .A1(n36963), .A2(n36964), .B1(n5900), .B2(n19052), .ZN(
        n19051) );
  NOR2_X1 U25553 ( .A1(n9130), .A2(n5903), .ZN(n33447) );
  NOR2_X1 U25556 ( .A1(n34500), .A2(n5903), .ZN(n34499) );
  NAND2_X1 U25559 ( .A1(n14226), .A2(n5907), .ZN(n19819) );
  INV_X1 U25560 ( .I(n50094), .ZN(n47928) );
  NAND2_X2 U25563 ( .A1(n46753), .A2(n20344), .ZN(n20340) );
  XOR2_X1 U25565 ( .A1(n5913), .A2(n5914), .Z(n7036) );
  XOR2_X1 U25566 ( .A1(n52065), .A2(n5878), .Z(n5914) );
  NOR2_X2 U25567 ( .A1(n41132), .A2(n11243), .ZN(n10041) );
  XOR2_X1 U25577 ( .A1(n33837), .A2(n33231), .Z(n16809) );
  XOR2_X1 U25578 ( .A1(n20623), .A2(n22652), .Z(n24145) );
  NOR2_X2 U25579 ( .A1(n22715), .A2(n25082), .ZN(n22652) );
  XOR2_X1 U25584 ( .A1(n11234), .A2(n5920), .Z(n5919) );
  XOR2_X1 U25585 ( .A1(n5922), .A2(n19101), .Z(n5920) );
  XOR2_X1 U25586 ( .A1(n13548), .A2(n39544), .Z(n5922) );
  XOR2_X1 U25587 ( .A1(n5923), .A2(n44434), .Z(n44435) );
  XOR2_X1 U25589 ( .A1(n25872), .A2(n10443), .Z(n5924) );
  XOR2_X1 U25590 ( .A1(n44608), .A2(n61498), .Z(n10443) );
  NOR2_X2 U25594 ( .A1(n5933), .A2(n5931), .ZN(n30885) );
  NAND2_X2 U25595 ( .A1(n11161), .A2(n11163), .ZN(n21838) );
  MUX2_X1 U25598 ( .I0(n22993), .I1(n36952), .S(n5936), .Z(n36954) );
  NAND2_X2 U25600 ( .A1(n47209), .A2(n9045), .ZN(n48463) );
  NOR2_X2 U25601 ( .A1(n19928), .A2(n23350), .ZN(n42386) );
  OAI22_X1 U25603 ( .A1(n47635), .A2(n14473), .B1(n7579), .B2(n5940), .ZN(
        n47638) );
  NAND3_X2 U25604 ( .A1(n47876), .A2(n47882), .A3(n12647), .ZN(n5940) );
  XOR2_X1 U25605 ( .A1(n51731), .A2(n5941), .Z(n6117) );
  XOR2_X1 U25606 ( .A1(n51806), .A2(n5943), .Z(n5941) );
  XOR2_X1 U25607 ( .A1(n6364), .A2(n6217), .Z(n51806) );
  INV_X1 U25609 ( .I(n51730), .ZN(n5943) );
  NAND3_X1 U25613 ( .A1(n58491), .A2(n61502), .A3(n5944), .ZN(n54482) );
  INV_X2 U25616 ( .I(n5950), .ZN(n23875) );
  XOR2_X1 U25620 ( .A1(n38828), .A2(n25021), .Z(n5952) );
  INV_X2 U25621 ( .I(n5953), .ZN(n6938) );
  XOR2_X1 U25623 ( .A1(n17907), .A2(n5955), .Z(n5954) );
  XOR2_X1 U25624 ( .A1(n43664), .A2(n44273), .Z(n5955) );
  XOR2_X1 U25626 ( .A1(n6174), .A2(n12038), .Z(n5957) );
  NOR2_X2 U25627 ( .A1(n34914), .A2(n22737), .ZN(n35430) );
  AND2_X1 U25628 ( .A1(n35425), .A2(n22993), .Z(n5960) );
  NAND2_X1 U25630 ( .A1(n1581), .A2(n53489), .ZN(n5963) );
  XOR2_X1 U25634 ( .A1(n5969), .A2(n43724), .Z(n18955) );
  XOR2_X1 U25638 ( .A1(n18545), .A2(n24753), .Z(n17078) );
  OAI21_X2 U25639 ( .A1(n39689), .A2(n39275), .B(n16731), .ZN(n24753) );
  NAND3_X2 U25641 ( .A1(n16734), .A2(n16735), .A3(n5974), .ZN(n39689) );
  NOR2_X1 U25642 ( .A1(n5977), .A2(n5975), .ZN(n5974) );
  NAND2_X1 U25643 ( .A1(n26052), .A2(n63430), .ZN(n5976) );
  INV_X2 U25644 ( .I(n24007), .ZN(n46950) );
  INV_X2 U25645 ( .I(n12735), .ZN(n42235) );
  XOR2_X1 U25646 ( .A1(n19069), .A2(n31810), .Z(n5981) );
  NAND2_X1 U25648 ( .A1(n47229), .A2(n9758), .ZN(n44653) );
  NOR2_X2 U25650 ( .A1(n3932), .A2(n20753), .ZN(n5982) );
  XOR2_X1 U25651 ( .A1(n5710), .A2(n5990), .Z(n5986) );
  XOR2_X1 U25652 ( .A1(n5988), .A2(n44819), .Z(n5987) );
  XOR2_X1 U25653 ( .A1(n5992), .A2(n22212), .Z(n44819) );
  XOR2_X1 U25654 ( .A1(n5991), .A2(n44593), .Z(n5988) );
  XOR2_X1 U25655 ( .A1(n46550), .A2(n22247), .Z(n5991) );
  XOR2_X1 U25656 ( .A1(n45246), .A2(n21940), .Z(n5992) );
  OAI21_X1 U25657 ( .A1(n43030), .A2(n43029), .B(n57256), .ZN(n43031) );
  INV_X2 U25662 ( .I(n6012), .ZN(n14834) );
  XOR2_X1 U25665 ( .A1(n51910), .A2(n51909), .Z(n51996) );
  AOI21_X1 U25667 ( .A1(n42293), .A2(n42299), .B(n6016), .ZN(n38270) );
  NAND3_X1 U25668 ( .A1(n42506), .A2(n13725), .A3(n6016), .ZN(n42513) );
  NAND2_X2 U25669 ( .A1(n22882), .A2(n41856), .ZN(n6016) );
  NAND3_X2 U25670 ( .A1(n15609), .A2(n6018), .A3(n6017), .ZN(n11424) );
  OAI21_X2 U25671 ( .A1(n1200), .A2(n38994), .B(n6019), .ZN(n6092) );
  NAND2_X2 U25672 ( .A1(n14891), .A2(n14894), .ZN(n38994) );
  AOI21_X1 U25674 ( .A1(n54825), .A2(n5711), .B(n15761), .ZN(n54826) );
  AOI21_X1 U25675 ( .A1(n54096), .A2(n5711), .B(n54443), .ZN(n51636) );
  NAND3_X1 U25678 ( .A1(n7818), .A2(n32948), .A3(n6025), .ZN(n7817) );
  INV_X2 U25681 ( .I(n26568), .ZN(n28231) );
  NAND2_X2 U25682 ( .A1(n28035), .A2(n14834), .ZN(n26568) );
  XOR2_X1 U25683 ( .A1(n58433), .A2(n1549), .Z(n11845) );
  INV_X2 U25685 ( .I(n6027), .ZN(n49905) );
  NOR2_X1 U25686 ( .A1(n48732), .A2(n6027), .ZN(n48733) );
  NAND2_X2 U25688 ( .A1(n21406), .A2(n49901), .ZN(n6027) );
  XOR2_X1 U25691 ( .A1(n6756), .A2(n6755), .Z(n6031) );
  NOR2_X2 U25692 ( .A1(n53525), .A2(n6032), .ZN(n53503) );
  NOR2_X1 U25693 ( .A1(n53500), .A2(n6032), .ZN(n6078) );
  OAI21_X1 U25694 ( .A1(n53521), .A2(n6032), .B(n53497), .ZN(n6077) );
  NAND2_X2 U25695 ( .A1(n25789), .A2(n53492), .ZN(n6032) );
  NAND2_X1 U25696 ( .A1(n6033), .A2(n33670), .ZN(n31598) );
  NAND2_X1 U25697 ( .A1(n61746), .A2(n6170), .ZN(n38196) );
  NAND3_X1 U25698 ( .A1(n42447), .A2(n59674), .A3(n61746), .ZN(n6197) );
  XOR2_X1 U25704 ( .A1(n6036), .A2(n44321), .Z(n6035) );
  XOR2_X1 U25705 ( .A1(n24262), .A2(n46650), .Z(n44321) );
  XOR2_X1 U25706 ( .A1(n18624), .A2(n44506), .Z(n6036) );
  XOR2_X1 U25707 ( .A1(n16439), .A2(n7522), .Z(n10645) );
  NAND2_X1 U25710 ( .A1(n6041), .A2(n29566), .ZN(n28951) );
  XOR2_X1 U25718 ( .A1(n13975), .A2(n6133), .Z(n6045) );
  INV_X1 U25721 ( .I(n6048), .ZN(n6047) );
  NOR3_X2 U25726 ( .A1(n19950), .A2(n19949), .A3(n24410), .ZN(n24180) );
  NAND2_X2 U25727 ( .A1(n11347), .A2(n6054), .ZN(n35353) );
  XOR2_X1 U25728 ( .A1(n10893), .A2(n14514), .Z(n45375) );
  NOR4_X2 U25731 ( .A1(n61910), .A2(n6060), .A3(n1084), .A4(n47010), .ZN(n6059) );
  NAND2_X2 U25736 ( .A1(n5731), .A2(n24181), .ZN(n11064) );
  XOR2_X1 U25738 ( .A1(n14878), .A2(n38255), .Z(n6062) );
  XOR2_X1 U25739 ( .A1(n38791), .A2(n38252), .Z(n6065) );
  NAND2_X2 U25740 ( .A1(n63435), .A2(n6305), .ZN(n41947) );
  NAND2_X2 U25744 ( .A1(n26034), .A2(n814), .ZN(n10187) );
  NAND3_X2 U25746 ( .A1(n271), .A2(n4688), .A3(n11275), .ZN(n54408) );
  INV_X1 U25748 ( .I(n54408), .ZN(n54413) );
  XOR2_X1 U25749 ( .A1(n6092), .A2(n55840), .Z(n6846) );
  CLKBUF_X4 U25751 ( .I(n12127), .Z(n6095) );
  NAND2_X2 U25752 ( .A1(n2232), .A2(n1533), .ZN(n35765) );
  XOR2_X1 U25753 ( .A1(n6097), .A2(n43673), .Z(n6096) );
  NOR2_X2 U25754 ( .A1(n6101), .A2(n39824), .ZN(n6100) );
  OR2_X1 U25755 ( .A1(n39826), .A2(n40000), .Z(n6103) );
  XOR2_X1 U25760 ( .A1(n15938), .A2(n6780), .Z(n6113) );
  XOR2_X1 U25761 ( .A1(n6114), .A2(n952), .Z(n10811) );
  NAND2_X2 U25763 ( .A1(n29432), .A2(n28959), .ZN(n29442) );
  NAND2_X2 U25764 ( .A1(n27104), .A2(n6120), .ZN(n29432) );
  NAND2_X1 U25765 ( .A1(n31846), .A2(n10337), .ZN(n6125) );
  XOR2_X1 U25766 ( .A1(n8288), .A2(n6126), .Z(n31840) );
  XOR2_X1 U25767 ( .A1(n6127), .A2(n23143), .Z(n6126) );
  INV_X2 U25769 ( .I(n6129), .ZN(n53615) );
  NAND2_X2 U25773 ( .A1(n8690), .A2(n43989), .ZN(n19761) );
  NOR2_X2 U25774 ( .A1(n42222), .A2(n42223), .ZN(n43989) );
  NAND3_X1 U25776 ( .A1(n6135), .A2(n54012), .A3(n53992), .ZN(n53971) );
  OAI21_X1 U25778 ( .A1(n53931), .A2(n6135), .B(n58817), .ZN(n53930) );
  XOR2_X1 U25779 ( .A1(n45040), .A2(n6136), .Z(n20328) );
  XOR2_X1 U25780 ( .A1(n3208), .A2(n44217), .Z(n44218) );
  XOR2_X1 U25781 ( .A1(n20950), .A2(n6136), .Z(n44384) );
  INV_X2 U25783 ( .I(n23469), .ZN(n28035) );
  XOR2_X1 U25785 ( .A1(n9876), .A2(n54587), .Z(n50616) );
  XOR2_X1 U25787 ( .A1(n8228), .A2(n1465), .Z(n52175) );
  XOR2_X1 U25788 ( .A1(n6143), .A2(n6142), .Z(n6141) );
  XOR2_X1 U25789 ( .A1(n6336), .A2(n52537), .Z(n6142) );
  XOR2_X1 U25790 ( .A1(n52173), .A2(n23173), .Z(n6143) );
  NAND2_X1 U25792 ( .A1(n38348), .A2(n6144), .ZN(n7348) );
  AOI22_X1 U25793 ( .A1(n38352), .A2(n43350), .B1(n6144), .B2(n38353), .ZN(
        n7139) );
  XOR2_X1 U25796 ( .A1(n36370), .A2(n22953), .Z(n38861) );
  NAND3_X2 U25799 ( .A1(n6146), .A2(n15402), .A3(n10557), .ZN(n11074) );
  INV_X2 U25801 ( .I(n25106), .ZN(n22160) );
  INV_X2 U25811 ( .I(n31840), .ZN(n35802) );
  XOR2_X1 U25816 ( .A1(n6161), .A2(n6160), .Z(n39293) );
  INV_X1 U25820 ( .I(n42363), .ZN(n6164) );
  XOR2_X1 U25821 ( .A1(n31773), .A2(n13833), .Z(n7205) );
  XOR2_X1 U25822 ( .A1(n6166), .A2(n37971), .Z(n37972) );
  NAND2_X2 U25825 ( .A1(n6170), .A2(n1733), .ZN(n7094) );
  XOR2_X1 U25826 ( .A1(n46178), .A2(n1214), .Z(n6171) );
  XOR2_X1 U25827 ( .A1(n62574), .A2(n47940), .Z(n21994) );
  XOR2_X1 U25828 ( .A1(n62574), .A2(n51361), .Z(n50708) );
  NAND2_X2 U25831 ( .A1(n44651), .A2(n46049), .ZN(n46048) );
  NAND2_X2 U25832 ( .A1(n6173), .A2(n15697), .ZN(n44651) );
  XOR2_X1 U25834 ( .A1(n43265), .A2(n45316), .Z(n6174) );
  XOR2_X1 U25835 ( .A1(n59694), .A2(n54563), .Z(n45316) );
  NAND2_X2 U25838 ( .A1(n1664), .A2(n7579), .ZN(n14289) );
  OR2_X1 U25839 ( .A1(n14289), .A2(n45183), .Z(n45177) );
  INV_X1 U25847 ( .I(n53294), .ZN(n19594) );
  XOR2_X1 U25851 ( .A1(n22551), .A2(n6204), .Z(n44419) );
  XOR2_X1 U25852 ( .A1(n6204), .A2(n22994), .Z(n46629) );
  XOR2_X1 U25853 ( .A1(n10713), .A2(n6204), .Z(n44612) );
  XOR2_X1 U25855 ( .A1(n24918), .A2(n22697), .Z(n6207) );
  XOR2_X1 U25856 ( .A1(n6208), .A2(n19889), .Z(n51676) );
  XOR2_X1 U25857 ( .A1(n60448), .A2(n6209), .Z(n6208) );
  XOR2_X1 U25858 ( .A1(n6210), .A2(n19888), .Z(n19890) );
  XOR2_X1 U25859 ( .A1(n51972), .A2(n51664), .Z(n6209) );
  XOR2_X1 U25861 ( .A1(n51762), .A2(n51087), .Z(n51972) );
  NAND4_X2 U25863 ( .A1(n737), .A2(n6214), .A3(n19520), .A4(n6213), .ZN(n19519) );
  OAI21_X1 U25866 ( .A1(n6857), .A2(n6215), .B(n6856), .ZN(n6859) );
  NAND2_X1 U25868 ( .A1(n54501), .A2(n1610), .ZN(n24512) );
  XOR2_X1 U25870 ( .A1(n6216), .A2(n51729), .Z(n6217) );
  NOR2_X2 U25872 ( .A1(n6366), .A2(n6365), .ZN(n18191) );
  AOI22_X1 U25874 ( .A1(n27057), .A2(n6222), .B1(n27056), .B2(n9685), .ZN(
        n27058) );
  NAND2_X1 U25876 ( .A1(n56560), .A2(n1596), .ZN(n56663) );
  XOR2_X1 U25877 ( .A1(n58819), .A2(n50794), .Z(n6224) );
  NAND2_X2 U25879 ( .A1(n43917), .A2(n6225), .ZN(n18919) );
  NOR2_X2 U25880 ( .A1(n48688), .A2(n10636), .ZN(n49057) );
  NAND3_X2 U25882 ( .A1(n6233), .A2(n43780), .A3(n6232), .ZN(n44329) );
  NAND3_X2 U25884 ( .A1(n55267), .A2(n55265), .A3(n64255), .ZN(n6235) );
  INV_X2 U25887 ( .I(n4512), .ZN(n35915) );
  INV_X2 U25891 ( .I(n6747), .ZN(n22852) );
  NOR2_X2 U25892 ( .A1(n18651), .A2(n35735), .ZN(n20865) );
  INV_X2 U25898 ( .I(n6245), .ZN(n35756) );
  XOR2_X1 U25902 ( .A1(n6251), .A2(n32509), .Z(n32510) );
  XOR2_X1 U25904 ( .A1(n6252), .A2(n44532), .Z(n46874) );
  XOR2_X1 U25905 ( .A1(n45044), .A2(n7202), .Z(n6253) );
  INV_X4 U25909 ( .I(n12908), .ZN(n16279) );
  OAI21_X1 U25914 ( .A1(n29592), .A2(n6270), .B(n6269), .ZN(n28914) );
  NAND2_X2 U25916 ( .A1(n23723), .A2(n16235), .ZN(n30347) );
  OAI21_X1 U25918 ( .A1(n35980), .A2(n10849), .B(n57210), .ZN(n22895) );
  NAND2_X2 U25923 ( .A1(n23033), .A2(n6273), .ZN(n21854) );
  XOR2_X1 U25925 ( .A1(n20715), .A2(n433), .Z(n31744) );
  XOR2_X1 U25926 ( .A1(n24911), .A2(n6275), .Z(n6274) );
  NOR2_X1 U25927 ( .A1(n60172), .A2(n6276), .ZN(n37935) );
  INV_X1 U25931 ( .I(n18229), .ZN(n54559) );
  NAND2_X2 U25934 ( .A1(n44779), .A2(n25444), .ZN(n45766) );
  NOR2_X2 U25936 ( .A1(n24198), .A2(n57939), .ZN(n35507) );
  XOR2_X1 U25944 ( .A1(n5913), .A2(n411), .Z(n6294) );
  XOR2_X1 U25946 ( .A1(n18537), .A2(n10252), .Z(n6296) );
  XOR2_X1 U25947 ( .A1(n25721), .A2(n23062), .Z(n11439) );
  XOR2_X1 U25948 ( .A1(n25721), .A2(n38298), .Z(n9492) );
  XOR2_X1 U25949 ( .A1(n6301), .A2(n13949), .Z(n6300) );
  INV_X1 U25950 ( .I(n45513), .ZN(n44197) );
  NAND2_X2 U25952 ( .A1(n5346), .A2(n44779), .ZN(n18361) );
  INV_X1 U25954 ( .I(n6302), .ZN(n38210) );
  AOI21_X1 U25957 ( .A1(n29611), .A2(n11975), .B(n6303), .ZN(n14940) );
  OAI21_X1 U25958 ( .A1(n26888), .A2(n6303), .B(n28172), .ZN(n26889) );
  NAND3_X2 U25959 ( .A1(n6304), .A2(n33004), .A3(n65256), .ZN(n33616) );
  NAND2_X2 U25960 ( .A1(n33408), .A2(n6304), .ZN(n33405) );
  XOR2_X1 U25963 ( .A1(n6308), .A2(n26063), .Z(n6307) );
  XOR2_X1 U25964 ( .A1(n6309), .A2(n20554), .Z(n14597) );
  NOR2_X1 U25966 ( .A1(n6313), .A2(n49739), .ZN(n16239) );
  XOR2_X1 U25969 ( .A1(n16595), .A2(n6314), .Z(n49155) );
  AOI21_X1 U25971 ( .A1(n48398), .A2(n6314), .B(n48397), .ZN(n8579) );
  OAI21_X1 U25973 ( .A1(n61601), .A2(n47623), .B(n47244), .ZN(n45993) );
  AOI22_X2 U25974 ( .A1(n40367), .A2(n1490), .B1(n43366), .B2(n42735), .ZN(
        n40372) );
  INV_X2 U25976 ( .I(n31276), .ZN(n6317) );
  NOR2_X1 U25987 ( .A1(n6329), .A2(n36492), .ZN(n36499) );
  NAND2_X1 U25998 ( .A1(n7912), .A2(n6341), .ZN(n20663) );
  AND2_X1 U25999 ( .A1(n6341), .A2(n58205), .Z(n6340) );
  CLKBUF_X4 U26000 ( .I(n19619), .Z(n6345) );
  INV_X2 U26001 ( .I(n19426), .ZN(n19619) );
  CLKBUF_X4 U26006 ( .I(n19598), .Z(n6349) );
  NAND3_X2 U26010 ( .A1(n18487), .A2(n20319), .A3(n6351), .ZN(n53181) );
  NOR2_X1 U26012 ( .A1(n53177), .A2(n63126), .ZN(n20353) );
  XOR2_X1 U26015 ( .A1(n1347), .A2(n32722), .Z(n21522) );
  XOR2_X1 U26018 ( .A1(n6353), .A2(n54536), .Z(Plaintext[74]) );
  OR2_X1 U26019 ( .A1(n54540), .A2(n6356), .Z(n6355) );
  XOR2_X1 U26020 ( .A1(n18012), .A2(n18011), .Z(n6358) );
  INV_X2 U26022 ( .I(n6721), .ZN(n34080) );
  NAND2_X2 U26026 ( .A1(n6375), .A2(n6371), .ZN(n19624) );
  AOI22_X1 U26029 ( .A1(n61787), .A2(n56573), .B1(n6379), .B2(n51251), .ZN(
        n6391) );
  NAND2_X1 U26031 ( .A1(n6345), .A2(n6380), .ZN(n26848) );
  NAND2_X1 U26032 ( .A1(n6381), .A2(n26856), .ZN(n6380) );
  XOR2_X1 U26035 ( .A1(n22979), .A2(n6383), .Z(n6385) );
  INV_X2 U26037 ( .I(n6386), .ZN(n9011) );
  NAND2_X1 U26041 ( .A1(n42918), .A2(n6388), .ZN(n14183) );
  NAND2_X2 U26042 ( .A1(n42554), .A2(n42916), .ZN(n6388) );
  INV_X2 U26043 ( .I(n15697), .ZN(n47985) );
  AND2_X1 U26044 ( .A1(n46048), .A2(n46940), .Z(n44643) );
  XOR2_X1 U26045 ( .A1(n8563), .A2(n1835), .Z(n10270) );
  NOR2_X2 U26047 ( .A1(n6392), .A2(n6390), .ZN(n56144) );
  MUX2_X1 U26048 ( .I0(n6394), .I1(n18386), .S(n8367), .Z(n6393) );
  NAND2_X1 U26049 ( .A1(n18255), .A2(n56564), .ZN(n6394) );
  XOR2_X1 U26054 ( .A1(n7761), .A2(n22373), .Z(n6403) );
  INV_X2 U26055 ( .I(n6404), .ZN(n18335) );
  XOR2_X1 U26056 ( .A1(n31556), .A2(n31804), .Z(n32574) );
  NOR2_X2 U26057 ( .A1(n6406), .A2(n30316), .ZN(n31804) );
  XOR2_X1 U26062 ( .A1(n6415), .A2(n6414), .Z(n6617) );
  XOR2_X1 U26063 ( .A1(n45100), .A2(n21989), .Z(n6414) );
  XOR2_X1 U26064 ( .A1(n46385), .A2(n19766), .Z(n45100) );
  XOR2_X1 U26065 ( .A1(n5710), .A2(n44153), .Z(n6416) );
  NAND2_X1 U26066 ( .A1(n41547), .A2(n42736), .ZN(n6427) );
  XOR2_X1 U26075 ( .A1(n59926), .A2(n36733), .Z(n6437) );
  NAND2_X1 U26077 ( .A1(n6439), .A2(n6611), .ZN(n32454) );
  XOR2_X1 U26078 ( .A1(n14215), .A2(n849), .Z(n6611) );
  INV_X2 U26079 ( .I(n60014), .ZN(n36385) );
  XOR2_X1 U26083 ( .A1(n4947), .A2(n50832), .Z(n38142) );
  XOR2_X1 U26084 ( .A1(n6441), .A2(n51290), .Z(n15320) );
  XOR2_X1 U26085 ( .A1(n4947), .A2(n39253), .Z(n39004) );
  NAND2_X1 U26088 ( .A1(n40857), .A2(n63119), .ZN(n40398) );
  INV_X1 U26099 ( .I(n42088), .ZN(n6453) );
  XOR2_X1 U26100 ( .A1(n31647), .A2(n6455), .Z(n6454) );
  XOR2_X1 U26101 ( .A1(n65197), .A2(n31646), .Z(n6455) );
  XOR2_X1 U26102 ( .A1(n32271), .A2(n6457), .Z(n6456) );
  NOR2_X1 U26106 ( .A1(n6467), .A2(n19102), .ZN(n40089) );
  NOR2_X1 U26107 ( .A1(n25246), .A2(n6467), .ZN(n12679) );
  NOR2_X1 U26111 ( .A1(n21134), .A2(n1838), .ZN(n6473) );
  XOR2_X1 U26119 ( .A1(n23667), .A2(n6482), .Z(n6481) );
  XOR2_X1 U26120 ( .A1(n17608), .A2(n31995), .Z(n6483) );
  OR2_X1 U26123 ( .A1(n23127), .A2(n25509), .Z(n15989) );
  INV_X2 U26125 ( .I(n19883), .ZN(n29643) );
  AOI21_X1 U26126 ( .A1(n19581), .A2(n28847), .B(n28846), .ZN(n19549) );
  NAND2_X2 U26127 ( .A1(n28842), .A2(n26856), .ZN(n28595) );
  NAND2_X2 U26128 ( .A1(n26061), .A2(n19883), .ZN(n28588) );
  NOR2_X1 U26129 ( .A1(n34740), .A2(n23354), .ZN(n34743) );
  NOR2_X2 U26132 ( .A1(n51863), .A2(n54025), .ZN(n53031) );
  NAND2_X2 U26134 ( .A1(n43305), .A2(n20526), .ZN(n43710) );
  NAND2_X2 U26138 ( .A1(n24359), .A2(n21090), .ZN(n46943) );
  NAND3_X2 U26140 ( .A1(n19620), .A2(n23386), .A3(n28598), .ZN(n28845) );
  NAND2_X1 U26141 ( .A1(n22443), .A2(n28598), .ZN(n22442) );
  XOR2_X1 U26145 ( .A1(n6501), .A2(n24699), .Z(n6500) );
  INV_X2 U26147 ( .I(n7835), .ZN(n56983) );
  NAND2_X2 U26148 ( .A1(n8597), .A2(n7835), .ZN(n56606) );
  XOR2_X1 U26151 ( .A1(n18191), .A2(n19488), .Z(n6502) );
  INV_X2 U26152 ( .I(n15545), .ZN(n15815) );
  INV_X2 U26153 ( .I(n11766), .ZN(n7663) );
  XOR2_X1 U26155 ( .A1(n6504), .A2(n9040), .Z(n33230) );
  XOR2_X1 U26156 ( .A1(n32495), .A2(n129), .Z(n6504) );
  XOR2_X1 U26157 ( .A1(n16502), .A2(n11766), .Z(n6505) );
  XOR2_X1 U26158 ( .A1(n9179), .A2(n7887), .Z(n11766) );
  INV_X1 U26159 ( .I(n64667), .ZN(n34437) );
  AOI21_X1 U26162 ( .A1(n33815), .A2(n64667), .B(n65205), .ZN(n33816) );
  NOR3_X1 U26165 ( .A1(n18827), .A2(n6508), .A3(n39057), .ZN(n18853) );
  XOR2_X1 U26166 ( .A1(n25137), .A2(n40613), .Z(n6508) );
  XOR2_X1 U26170 ( .A1(n8553), .A2(n1288), .Z(n6959) );
  NAND2_X2 U26176 ( .A1(n19593), .A2(n29641), .ZN(n6513) );
  XOR2_X1 U26177 ( .A1(n703), .A2(n38888), .Z(n19101) );
  XOR2_X1 U26178 ( .A1(n6517), .A2(n17406), .Z(n6516) );
  XOR2_X1 U26179 ( .A1(n39188), .A2(n39187), .Z(n6517) );
  XOR2_X1 U26180 ( .A1(n11700), .A2(n9376), .Z(n39547) );
  XOR2_X1 U26183 ( .A1(n18276), .A2(n23518), .Z(n39189) );
  NOR2_X1 U26186 ( .A1(n65205), .A2(n35762), .ZN(n35763) );
  NAND2_X1 U26187 ( .A1(n65205), .A2(n35318), .ZN(n34433) );
  NAND2_X1 U26188 ( .A1(n35259), .A2(n65205), .ZN(n35260) );
  AOI22_X1 U26190 ( .A1(n21720), .A2(n6522), .B1(n29152), .B2(n27397), .ZN(
        n21633) );
  NAND3_X1 U26192 ( .A1(n6523), .A2(n47281), .A3(n47590), .ZN(n16510) );
  AOI22_X1 U26193 ( .A1(n47594), .A2(n45681), .B1(n548), .B2(n6523), .ZN(
        n45686) );
  XOR2_X1 U26196 ( .A1(n63004), .A2(n776), .Z(n15957) );
  XOR2_X1 U26197 ( .A1(n63004), .A2(n733), .Z(n22015) );
  XOR2_X1 U26198 ( .A1(n6524), .A2(n36994), .Z(n38292) );
  XOR2_X1 U26199 ( .A1(n6524), .A2(n13733), .Z(n13732) );
  NOR2_X2 U26202 ( .A1(n6527), .A2(n32678), .ZN(n6526) );
  NAND2_X2 U26203 ( .A1(n32684), .A2(n61647), .ZN(n6527) );
  NAND3_X2 U26206 ( .A1(n39433), .A2(n39432), .A3(n6532), .ZN(n44851) );
  NAND3_X2 U26207 ( .A1(n24179), .A2(n15020), .A3(n43286), .ZN(n43107) );
  NAND2_X2 U26208 ( .A1(n1493), .A2(n20844), .ZN(n43282) );
  NOR2_X1 U26210 ( .A1(n61892), .A2(n8602), .ZN(n6546) );
  NOR2_X2 U26212 ( .A1(n30242), .A2(n1862), .ZN(n30230) );
  NOR2_X2 U26213 ( .A1(n6555), .A2(n6554), .ZN(n22374) );
  XOR2_X1 U26214 ( .A1(n32657), .A2(n32654), .Z(n15676) );
  XOR2_X1 U26215 ( .A1(n32522), .A2(n32654), .Z(n32523) );
  NAND3_X1 U26217 ( .A1(n54400), .A2(n7138), .A3(n54390), .ZN(n6561) );
  NAND3_X1 U26218 ( .A1(n54394), .A2(n54403), .A3(n54414), .ZN(n6562) );
  NOR2_X2 U26219 ( .A1(n24275), .A2(n6565), .ZN(n18468) );
  XOR2_X1 U26220 ( .A1(n1464), .A2(n30908), .Z(n6566) );
  XOR2_X1 U26221 ( .A1(n21896), .A2(n44612), .Z(n6567) );
  XOR2_X1 U26222 ( .A1(n21895), .A2(n58964), .Z(n6568) );
  INV_X2 U26224 ( .I(n6570), .ZN(n17869) );
  XOR2_X1 U26226 ( .A1(n6578), .A2(n21608), .Z(n21607) );
  NOR2_X1 U26227 ( .A1(n59821), .A2(n18361), .ZN(n16245) );
  NAND2_X2 U26228 ( .A1(n36926), .A2(n35508), .ZN(n34924) );
  NAND2_X1 U26229 ( .A1(n6580), .A2(n14457), .ZN(n54463) );
  NAND2_X2 U26230 ( .A1(n46969), .A2(n48425), .ZN(n6583) );
  NAND2_X1 U26232 ( .A1(n23502), .A2(n6586), .ZN(n6585) );
  NAND3_X1 U26233 ( .A1(n6588), .A2(n1330), .A3(n24262), .ZN(n6587) );
  XOR2_X1 U26237 ( .A1(n25935), .A2(n25934), .Z(n31766) );
  XOR2_X1 U26239 ( .A1(n31316), .A2(n32592), .Z(n6593) );
  NAND2_X2 U26240 ( .A1(n40996), .A2(n40994), .ZN(n7257) );
  NOR2_X2 U26241 ( .A1(n34119), .A2(n15783), .ZN(n33953) );
  XOR2_X1 U26242 ( .A1(n2823), .A2(n23695), .Z(n23175) );
  XOR2_X1 U26243 ( .A1(n2823), .A2(n38507), .Z(n38509) );
  NOR2_X2 U26247 ( .A1(n20047), .A2(n16962), .ZN(n6598) );
  INV_X2 U26249 ( .I(n6605), .ZN(n32495) );
  XOR2_X1 U26251 ( .A1(n58839), .A2(n5729), .Z(n12593) );
  INV_X2 U26255 ( .I(n7814), .ZN(n18339) );
  NOR2_X2 U26256 ( .A1(n11207), .A2(n51866), .ZN(n54344) );
  NOR2_X2 U26257 ( .A1(n54026), .A2(n54017), .ZN(n54348) );
  NAND2_X2 U26261 ( .A1(n42407), .A2(n42404), .ZN(n42398) );
  INV_X2 U26263 ( .I(n6617), .ZN(n45768) );
  XOR2_X1 U26265 ( .A1(n64117), .A2(n45296), .Z(n45297) );
  XOR2_X1 U26266 ( .A1(n64117), .A2(n44329), .Z(n43781) );
  NOR2_X1 U26267 ( .A1(n54912), .A2(n22486), .ZN(n6621) );
  NAND2_X2 U26271 ( .A1(n11264), .A2(n39324), .ZN(n40213) );
  NAND2_X2 U26272 ( .A1(n6627), .A2(n36788), .ZN(n38548) );
  NAND2_X2 U26273 ( .A1(n37475), .A2(n6632), .ZN(n6627) );
  NAND2_X2 U26276 ( .A1(n37491), .A2(n37276), .ZN(n38544) );
  NAND2_X2 U26277 ( .A1(n37476), .A2(n61890), .ZN(n38546) );
  NAND2_X2 U26278 ( .A1(n36783), .A2(n36782), .ZN(n37476) );
  NOR2_X2 U26280 ( .A1(n47983), .A2(n18465), .ZN(n48790) );
  NAND2_X1 U26281 ( .A1(n55022), .A2(n6635), .ZN(n54854) );
  NAND3_X1 U26282 ( .A1(n55023), .A2(n55022), .A3(n6635), .ZN(n55026) );
  NAND2_X1 U26283 ( .A1(n18484), .A2(n6635), .ZN(n54643) );
  AOI22_X1 U26284 ( .A1(n7800), .A2(n3916), .B1(n7148), .B2(n6635), .ZN(n54330) );
  INV_X2 U26286 ( .I(n6636), .ZN(n7999) );
  INV_X1 U26287 ( .I(n42535), .ZN(n6638) );
  OAI21_X1 U26289 ( .A1(n40881), .A2(n40880), .B(n6640), .ZN(n40884) );
  NAND2_X2 U26290 ( .A1(n43290), .A2(n19591), .ZN(n6640) );
  INV_X2 U26291 ( .I(n6641), .ZN(n54292) );
  XOR2_X1 U26294 ( .A1(n6643), .A2(n51763), .Z(n52523) );
  XOR2_X1 U26296 ( .A1(n51762), .A2(n52423), .Z(n6644) );
  NAND2_X1 U26298 ( .A1(n54397), .A2(n61829), .ZN(n6647) );
  NOR2_X2 U26299 ( .A1(n7138), .A2(n5324), .ZN(n54383) );
  NAND2_X1 U26300 ( .A1(n6647), .A2(n54391), .ZN(n24194) );
  XOR2_X1 U26304 ( .A1(n6663), .A2(n55610), .Z(Plaintext[122]) );
  NAND2_X2 U26305 ( .A1(n6667), .A2(n6666), .ZN(n52223) );
  NOR2_X2 U26312 ( .A1(n23799), .A2(n31224), .ZN(n6680) );
  NAND2_X2 U26316 ( .A1(n4969), .A2(n36517), .ZN(n36515) );
  XOR2_X1 U26318 ( .A1(n46186), .A2(n9723), .Z(n6684) );
  NOR2_X1 U26319 ( .A1(n1702), .A2(n6685), .ZN(n41636) );
  NAND2_X2 U26320 ( .A1(n15091), .A2(n8986), .ZN(n6685) );
  XOR2_X1 U26326 ( .A1(n6691), .A2(n6690), .Z(n11209) );
  XOR2_X1 U26327 ( .A1(n51845), .A2(n20370), .Z(n6690) );
  XOR2_X1 U26328 ( .A1(n22305), .A2(n4846), .Z(n51845) );
  XOR2_X1 U26329 ( .A1(n6692), .A2(n6694), .Z(n6691) );
  XOR2_X1 U26330 ( .A1(n6693), .A2(n62818), .Z(n6692) );
  XOR2_X1 U26331 ( .A1(n21097), .A2(n15447), .Z(n6693) );
  MUX2_X1 U26335 ( .I0(n23485), .I1(n43057), .S(n59650), .Z(n43064) );
  XOR2_X1 U26346 ( .A1(n6701), .A2(n32539), .Z(n10539) );
  XOR2_X1 U26347 ( .A1(n6701), .A2(n25176), .Z(n28930) );
  XOR2_X1 U26348 ( .A1(n33141), .A2(n6701), .Z(n31603) );
  XOR2_X1 U26349 ( .A1(n24008), .A2(n6701), .Z(n31987) );
  XOR2_X1 U26350 ( .A1(n33269), .A2(n6701), .Z(n33140) );
  NAND3_X1 U26351 ( .A1(n6702), .A2(n13985), .A3(n59851), .ZN(n39893) );
  NOR2_X2 U26352 ( .A1(n25742), .A2(n24389), .ZN(n13985) );
  XOR2_X1 U26354 ( .A1(n6849), .A2(n6703), .Z(n38289) );
  NOR2_X1 U26355 ( .A1(n49488), .A2(n6704), .ZN(n9353) );
  NOR2_X2 U26356 ( .A1(n10571), .A2(n47040), .ZN(n49500) );
  XOR2_X1 U26357 ( .A1(n7699), .A2(n1673), .Z(n17692) );
  XOR2_X1 U26368 ( .A1(n6711), .A2(n23120), .Z(n11190) );
  AOI21_X1 U26370 ( .A1(n1338), .A2(n6713), .B(n35053), .ZN(n35054) );
  NOR2_X1 U26371 ( .A1(n48030), .A2(n9853), .ZN(n15469) );
  NOR2_X1 U26372 ( .A1(n1472), .A2(n9853), .ZN(n49009) );
  AOI21_X1 U26375 ( .A1(n45512), .A2(n1070), .B(n46911), .ZN(n44784) );
  NOR2_X2 U26376 ( .A1(n22144), .A2(n27494), .ZN(n29302) );
  NAND2_X2 U26377 ( .A1(n29295), .A2(n6727), .ZN(n24233) );
  NAND2_X2 U26379 ( .A1(n24123), .A2(n11830), .ZN(n6720) );
  NOR2_X1 U26380 ( .A1(n6720), .A2(n30812), .ZN(n29237) );
  NAND2_X2 U26385 ( .A1(n64603), .A2(n25849), .ZN(n11992) );
  AOI21_X2 U26387 ( .A1(n33141), .A2(n32541), .B(n6723), .ZN(n10823) );
  XOR2_X1 U26392 ( .A1(n52360), .A2(n55889), .Z(n6725) );
  INV_X2 U26395 ( .I(n6728), .ZN(n12725) );
  INV_X2 U26396 ( .I(n8170), .ZN(n8337) );
  XOR2_X1 U26398 ( .A1(n4846), .A2(n50888), .Z(n50889) );
  XOR2_X1 U26399 ( .A1(n4311), .A2(n8569), .Z(n52361) );
  NOR2_X1 U26400 ( .A1(n6730), .A2(n47857), .ZN(n47862) );
  INV_X2 U26405 ( .I(n22509), .ZN(n49383) );
  NAND2_X2 U26406 ( .A1(n11609), .A2(n43053), .ZN(n43868) );
  OAI21_X1 U26407 ( .A1(n33224), .A2(n33531), .B(n20092), .ZN(n6736) );
  INV_X1 U26408 ( .I(n4835), .ZN(n54029) );
  MUX2_X1 U26409 ( .I0(n53881), .I1(n6737), .S(n54340), .Z(n53033) );
  XOR2_X1 U26414 ( .A1(n23571), .A2(n50611), .Z(n51808) );
  NOR2_X2 U26415 ( .A1(n19976), .A2(n15879), .ZN(n50611) );
  XOR2_X1 U26418 ( .A1(n51581), .A2(n53328), .Z(n6740) );
  NOR2_X2 U26420 ( .A1(n6743), .A2(n6742), .ZN(n19085) );
  NAND2_X1 U26421 ( .A1(n24482), .A2(n53034), .ZN(n53041) );
  NAND3_X1 U26422 ( .A1(n53040), .A2(n10527), .A3(n53039), .ZN(n16685) );
  XOR2_X1 U26424 ( .A1(n43135), .A2(n31602), .Z(n6745) );
  XOR2_X1 U26425 ( .A1(n51817), .A2(n38448), .Z(n43135) );
  BUF_X2 U26427 ( .I(n25292), .Z(n6748) );
  XOR2_X1 U26428 ( .A1(n14878), .A2(n36936), .Z(n6750) );
  XOR2_X1 U26430 ( .A1(n64373), .A2(n44092), .Z(n19071) );
  NOR2_X2 U26431 ( .A1(n42577), .A2(n42576), .ZN(n44092) );
  NOR2_X1 U26435 ( .A1(n6760), .A2(n24737), .ZN(n8005) );
  NAND2_X1 U26436 ( .A1(n20800), .A2(n6760), .ZN(n7206) );
  OAI22_X1 U26437 ( .A1(n34621), .A2(n6760), .B1(n34623), .B2(n34622), .ZN(
        n20206) );
  AOI21_X1 U26438 ( .A1(n32893), .A2(n6760), .B(n34623), .ZN(n25197) );
  AOI22_X1 U26439 ( .A1(n12539), .A2(n34085), .B1(n34084), .B2(n6760), .ZN(
        n10758) );
  NOR2_X1 U26440 ( .A1(n31524), .A2(n6760), .ZN(n31540) );
  INV_X2 U26444 ( .I(n6765), .ZN(n24908) );
  INV_X2 U26446 ( .I(n3356), .ZN(n40997) );
  NAND2_X2 U26447 ( .A1(n6776), .A2(n6772), .ZN(n29834) );
  AOI21_X1 U26448 ( .A1(n28802), .A2(n26994), .B(n10625), .ZN(n6778) );
  INV_X2 U26449 ( .I(n32076), .ZN(n37328) );
  INV_X1 U26454 ( .I(n37697), .ZN(n17512) );
  XNOR2_X1 U26458 ( .A1(n19155), .A2(n44182), .ZN(n15095) );
  NAND2_X2 U26460 ( .A1(n6785), .A2(n6784), .ZN(n20950) );
  INV_X2 U26461 ( .I(n15095), .ZN(n18133) );
  XOR2_X1 U26465 ( .A1(n2748), .A2(n54208), .Z(n44736) );
  NAND2_X2 U26466 ( .A1(n4283), .A2(n1232), .ZN(n6790) );
  NOR2_X1 U26467 ( .A1(n6790), .A2(n2014), .ZN(n53257) );
  NOR2_X1 U26468 ( .A1(n6789), .A2(n53279), .ZN(n13240) );
  NAND2_X1 U26472 ( .A1(n6792), .A2(n21082), .ZN(n7428) );
  NAND2_X1 U26473 ( .A1(n6792), .A2(n52768), .ZN(n22542) );
  INV_X2 U26476 ( .I(n8368), .ZN(n25685) );
  XOR2_X1 U26479 ( .A1(n22975), .A2(n45318), .Z(n6803) );
  INV_X2 U26480 ( .I(n6805), .ZN(n46814) );
  INV_X2 U26481 ( .I(n6808), .ZN(n25340) );
  NAND2_X2 U26482 ( .A1(n15748), .A2(n45436), .ZN(n11202) );
  INV_X2 U26484 ( .I(n6809), .ZN(n15748) );
  INV_X2 U26485 ( .I(n6810), .ZN(n23347) );
  XOR2_X1 U26490 ( .A1(n6812), .A2(n31707), .Z(n17821) );
  XOR2_X1 U26491 ( .A1(n6813), .A2(n61497), .Z(n6812) );
  XOR2_X1 U26492 ( .A1(n23152), .A2(n32494), .Z(n6813) );
  NOR2_X1 U26493 ( .A1(n18677), .A2(n6918), .ZN(n36707) );
  OAI21_X1 U26494 ( .A1(n11020), .A2(n6918), .B(n18205), .ZN(n35476) );
  XOR2_X1 U26496 ( .A1(n1522), .A2(n8665), .Z(n8497) );
  XOR2_X1 U26497 ( .A1(n23931), .A2(n6815), .Z(n8665) );
  NAND2_X2 U26498 ( .A1(n34606), .A2(n34035), .ZN(n34604) );
  NAND2_X1 U26505 ( .A1(n28038), .A2(n10537), .ZN(n6827) );
  NOR2_X2 U26510 ( .A1(n24373), .A2(n29148), .ZN(n29155) );
  NAND2_X1 U26511 ( .A1(n6829), .A2(n35247), .ZN(n35248) );
  OAI22_X1 U26513 ( .A1(n33278), .A2(n6829), .B1(n63773), .B2(n33802), .ZN(
        n33294) );
  NAND3_X1 U26514 ( .A1(n11089), .A2(n8879), .A3(n6829), .ZN(n8880) );
  NAND2_X1 U26517 ( .A1(n23226), .A2(n6831), .ZN(n37290) );
  NAND3_X1 U26519 ( .A1(n21536), .A2(n37360), .A3(n6831), .ZN(n18775) );
  INV_X4 U26521 ( .I(n4541), .ZN(n6831) );
  NAND3_X2 U26523 ( .A1(n6835), .A2(n6834), .A3(n6833), .ZN(n39709) );
  INV_X2 U26525 ( .I(n6839), .ZN(n41119) );
  NOR3_X2 U26529 ( .A1(n48587), .A2(n19200), .A3(n48487), .ZN(n48491) );
  INV_X2 U26530 ( .I(n48189), .ZN(n19200) );
  NAND2_X1 U26531 ( .A1(n41051), .A2(n41887), .ZN(n6843) );
  INV_X2 U26532 ( .I(n6844), .ZN(n46148) );
  INV_X2 U26533 ( .I(n6845), .ZN(n15934) );
  XOR2_X1 U26534 ( .A1(n6846), .A2(n16449), .Z(n38707) );
  XOR2_X1 U26535 ( .A1(n37807), .A2(n37806), .Z(n6847) );
  XOR2_X1 U26536 ( .A1(n38289), .A2(n39480), .Z(n6848) );
  XOR2_X1 U26537 ( .A1(n10767), .A2(n24058), .Z(n6849) );
  XOR2_X1 U26538 ( .A1(n37801), .A2(n6850), .Z(n39480) );
  XOR2_X1 U26539 ( .A1(n16450), .A2(n39626), .Z(n6850) );
  NAND2_X2 U26541 ( .A1(n6853), .A2(n22525), .ZN(n12806) );
  OAI22_X1 U26542 ( .A1(n39867), .A2(n4383), .B1(n9935), .B2(n61850), .ZN(
        n39868) );
  NAND2_X2 U26544 ( .A1(n1739), .A2(n40408), .ZN(n6853) );
  NAND2_X1 U26545 ( .A1(n6855), .A2(n41051), .ZN(n40844) );
  NAND2_X1 U26546 ( .A1(n41877), .A2(n6855), .ZN(n24791) );
  NAND2_X1 U26550 ( .A1(n6861), .A2(n61643), .ZN(n6860) );
  OAI21_X1 U26551 ( .A1(n16981), .A2(n15650), .B(n28035), .ZN(n6861) );
  NOR2_X1 U26555 ( .A1(n34994), .A2(n6867), .ZN(n13536) );
  XOR2_X1 U26557 ( .A1(n7203), .A2(n1671), .Z(n6871) );
  NAND2_X1 U26562 ( .A1(n6881), .A2(n9677), .ZN(n18383) );
  INV_X2 U26566 ( .I(n44466), .ZN(n44465) );
  XOR2_X1 U26567 ( .A1(n1268), .A2(n19864), .Z(n44466) );
  XOR2_X1 U26568 ( .A1(n44190), .A2(n44465), .Z(n44191) );
  INV_X2 U26570 ( .I(n6886), .ZN(n29148) );
  NOR2_X1 U26573 ( .A1(n1648), .A2(n46905), .ZN(n16238) );
  NAND2_X2 U26578 ( .A1(n20477), .A2(n1583), .ZN(n6902) );
  INV_X1 U26581 ( .I(n12177), .ZN(n19798) );
  NAND2_X1 U26587 ( .A1(n35086), .A2(n24370), .ZN(n35081) );
  NAND2_X1 U26589 ( .A1(n42479), .A2(n19638), .ZN(n6911) );
  NOR2_X1 U26594 ( .A1(n26383), .A2(n6913), .ZN(n26384) );
  OAI21_X1 U26595 ( .A1(n35677), .A2(n6914), .B(n24614), .ZN(n6956) );
  NAND2_X1 U26596 ( .A1(n35674), .A2(n17400), .ZN(n18382) );
  NOR2_X1 U26597 ( .A1(n35674), .A2(n17400), .ZN(n6915) );
  INV_X2 U26599 ( .I(n6917), .ZN(n51986) );
  NOR3_X2 U26601 ( .A1(n6920), .A2(n941), .A3(n19664), .ZN(n6919) );
  NAND2_X1 U26602 ( .A1(n42614), .A2(n6926), .ZN(n8788) );
  NAND2_X1 U26606 ( .A1(n40296), .A2(n58970), .ZN(n9092) );
  NAND2_X1 U26607 ( .A1(n14016), .A2(n6932), .ZN(n14015) );
  NAND2_X2 U26611 ( .A1(n23588), .A2(n6934), .ZN(n6933) );
  XOR2_X1 U26613 ( .A1(n1038), .A2(n6936), .Z(n26158) );
  XOR2_X1 U26614 ( .A1(n46499), .A2(n14251), .Z(n6936) );
  INV_X2 U26615 ( .I(n20817), .ZN(n41982) );
  INV_X2 U26618 ( .I(n6940), .ZN(n11213) );
  XOR2_X1 U26620 ( .A1(n11213), .A2(n30897), .Z(n6941) );
  OR2_X1 U26626 ( .A1(n17555), .A2(n57017), .Z(n53219) );
  NAND2_X1 U26629 ( .A1(n35667), .A2(n33573), .ZN(n6955) );
  NOR2_X1 U26630 ( .A1(n46106), .A2(n25231), .ZN(n48661) );
  XOR2_X1 U26635 ( .A1(n8426), .A2(n51186), .Z(n6963) );
  XOR2_X1 U26636 ( .A1(n24953), .A2(n51128), .Z(n51186) );
  NOR2_X2 U26643 ( .A1(n6974), .A2(n6973), .ZN(n43820) );
  NOR2_X1 U26644 ( .A1(n41045), .A2(n42344), .ZN(n6974) );
  INV_X4 U26650 ( .I(n18599), .ZN(n50360) );
  OAI22_X1 U26660 ( .A1(n37398), .A2(n36835), .B1(n58285), .B2(n37408), .ZN(
        n35271) );
  INV_X2 U26663 ( .I(n6988), .ZN(n51388) );
  NAND3_X1 U26664 ( .A1(n24595), .A2(n11227), .A3(n9967), .ZN(n6990) );
  NOR2_X1 U26670 ( .A1(n23625), .A2(n6991), .ZN(n56610) );
  NAND2_X2 U26672 ( .A1(n15258), .A2(n24302), .ZN(n41447) );
  INV_X2 U26673 ( .I(n14638), .ZN(n15258) );
  XOR2_X1 U26674 ( .A1(n6994), .A2(n20115), .Z(n20114) );
  XOR2_X1 U26679 ( .A1(n17486), .A2(n6999), .Z(n6998) );
  XOR2_X1 U26680 ( .A1(n37688), .A2(n20193), .Z(n6999) );
  NAND2_X1 U26682 ( .A1(n58683), .A2(n17503), .ZN(n30830) );
  NAND3_X1 U26683 ( .A1(n60054), .A2(n34668), .A3(n25465), .ZN(n33456) );
  INV_X2 U26687 ( .I(n9084), .ZN(n24537) );
  NOR2_X2 U26690 ( .A1(n24941), .A2(n62623), .ZN(n7006) );
  INV_X1 U26694 ( .I(n48031), .ZN(n11641) );
  NAND2_X1 U26696 ( .A1(n48323), .A2(n49006), .ZN(n48325) );
  NAND2_X1 U26700 ( .A1(n53492), .A2(n7021), .ZN(n53494) );
  NAND2_X1 U26702 ( .A1(n25675), .A2(n7021), .ZN(n53471) );
  NOR2_X2 U26705 ( .A1(n53459), .A2(n19353), .ZN(n7020) );
  INV_X4 U26706 ( .I(n7022), .ZN(n19830) );
  INV_X1 U26707 ( .I(n30517), .ZN(n7025) );
  NOR2_X2 U26708 ( .A1(n1872), .A2(n18075), .ZN(n30517) );
  NOR2_X1 U26715 ( .A1(n10705), .A2(n34853), .ZN(n16988) );
  XOR2_X1 U26716 ( .A1(n19103), .A2(n7036), .Z(n24166) );
  OR3_X1 U26717 ( .A1(n15333), .A2(n18839), .A3(n30167), .Z(n18842) );
  NOR3_X1 U26718 ( .A1(n20881), .A2(n52649), .A3(n55112), .ZN(n52657) );
  INV_X1 U26720 ( .I(n1593), .ZN(n7986) );
  BUF_X2 U26729 ( .I(n23055), .Z(n7040) );
  OR2_X1 U26730 ( .A1(n36412), .A2(n18313), .Z(n16181) );
  INV_X4 U26731 ( .I(n7595), .ZN(n20922) );
  INV_X2 U26732 ( .I(n20462), .ZN(n45929) );
  NAND3_X1 U26735 ( .A1(n49330), .A2(n49329), .A3(n61513), .ZN(n11844) );
  XNOR2_X1 U26736 ( .A1(n37554), .A2(n35367), .ZN(n23356) );
  NAND3_X2 U26739 ( .A1(n11657), .A2(n12180), .A3(n12182), .ZN(n30255) );
  NOR2_X1 U26740 ( .A1(n13014), .A2(n13013), .ZN(n13012) );
  NOR2_X1 U26741 ( .A1(n43325), .A2(n14605), .ZN(n7048) );
  NOR2_X1 U26749 ( .A1(n46095), .A2(n12227), .ZN(n12226) );
  AND2_X2 U26750 ( .A1(n19638), .A2(n26067), .Z(n40039) );
  NOR2_X1 U26751 ( .A1(n56776), .A2(n56793), .ZN(n56777) );
  AOI21_X1 U26756 ( .A1(n43912), .A2(n43922), .B(n43911), .ZN(n43921) );
  INV_X2 U26764 ( .I(n7063), .ZN(n12100) );
  AND2_X1 U26765 ( .A1(n11073), .A2(n8518), .Z(n11052) );
  XOR2_X1 U26766 ( .A1(n7064), .A2(n31983), .Z(n7935) );
  XOR2_X1 U26767 ( .A1(n25876), .A2(n5489), .Z(n7064) );
  AOI22_X1 U26770 ( .A1(n43912), .A2(n43528), .B1(n43530), .B2(n61743), .ZN(
        n43535) );
  NOR2_X1 U26772 ( .A1(n23006), .A2(n25495), .ZN(n25493) );
  XOR2_X1 U26773 ( .A1(n7509), .A2(n39477), .Z(n7065) );
  INV_X4 U26774 ( .I(n7067), .ZN(n21701) );
  NAND2_X2 U26778 ( .A1(n25412), .A2(n42634), .ZN(n41702) );
  NAND2_X1 U26781 ( .A1(n42200), .A2(n57545), .ZN(n15814) );
  NOR3_X2 U26784 ( .A1(n7068), .A2(n15572), .A3(n15571), .ZN(n36469) );
  NOR2_X1 U26787 ( .A1(n23595), .A2(n20525), .ZN(n15922) );
  XOR2_X1 U26791 ( .A1(n18155), .A2(n31683), .Z(n7071) );
  INV_X4 U26792 ( .I(n8470), .ZN(n21512) );
  INV_X1 U26794 ( .I(n10200), .ZN(n14302) );
  INV_X2 U26797 ( .I(n7080), .ZN(n15536) );
  XOR2_X1 U26798 ( .A1(n15537), .A2(n1128), .Z(n7080) );
  NOR2_X2 U26800 ( .A1(n18531), .A2(n7081), .ZN(n28711) );
  XOR2_X1 U26801 ( .A1(n32107), .A2(n32106), .Z(n33291) );
  XOR2_X1 U26804 ( .A1(n39621), .A2(n980), .Z(n7082) );
  XOR2_X1 U26805 ( .A1(n32114), .A2(n32170), .Z(n32115) );
  XOR2_X1 U26806 ( .A1(n7084), .A2(n20041), .Z(n37383) );
  XOR2_X1 U26807 ( .A1(n38988), .A2(n37381), .Z(n7084) );
  XOR2_X1 U26808 ( .A1(n37637), .A2(n30402), .Z(n37257) );
  XOR2_X1 U26809 ( .A1(n51261), .A2(n55638), .Z(n30402) );
  INV_X2 U26813 ( .I(n12606), .ZN(n25168) );
  NOR2_X2 U26815 ( .A1(n18839), .A2(n17627), .ZN(n29029) );
  NAND2_X1 U26827 ( .A1(n30054), .A2(n9047), .ZN(n29056) );
  NAND2_X1 U26829 ( .A1(n53118), .A2(n53056), .ZN(n20525) );
  NAND2_X2 U26831 ( .A1(n18700), .A2(n22081), .ZN(n14259) );
  NAND2_X2 U26832 ( .A1(n8676), .A2(n42008), .ZN(n43092) );
  NAND2_X2 U26833 ( .A1(n13862), .A2(n13863), .ZN(n42008) );
  INV_X2 U26837 ( .I(n7096), .ZN(n12779) );
  INV_X2 U26841 ( .I(n7099), .ZN(n19291) );
  XOR2_X1 U26843 ( .A1(n44045), .A2(n16518), .Z(n9025) );
  NAND2_X2 U26844 ( .A1(n47934), .A2(n15603), .ZN(n15177) );
  NAND2_X2 U26845 ( .A1(n9924), .A2(n50090), .ZN(n47934) );
  NAND2_X1 U26847 ( .A1(n59052), .A2(n14357), .ZN(n7100) );
  AOI21_X1 U26853 ( .A1(n11625), .A2(n1395), .B(n20784), .ZN(n41364) );
  XOR2_X1 U26855 ( .A1(n7105), .A2(n2259), .Z(n33049) );
  XOR2_X1 U26856 ( .A1(n33048), .A2(n33047), .Z(n7105) );
  NAND2_X2 U26858 ( .A1(n20090), .A2(n12779), .ZN(n24820) );
  OR2_X2 U26862 ( .A1(n13694), .A2(n9940), .Z(n28381) );
  XOR2_X1 U26863 ( .A1(n31872), .A2(n23412), .Z(n31883) );
  INV_X4 U26869 ( .I(n37405), .ZN(n8195) );
  NAND3_X1 U26872 ( .A1(n21401), .A2(n28432), .A3(n8091), .ZN(n8090) );
  NOR2_X2 U26873 ( .A1(n21957), .A2(n56245), .ZN(n56407) );
  NAND2_X2 U26875 ( .A1(n23480), .A2(n46914), .ZN(n46905) );
  NAND2_X1 U26876 ( .A1(n7151), .A2(n7152), .ZN(n7117) );
  OR2_X1 U26878 ( .A1(n11035), .A2(n50218), .Z(n47996) );
  AOI21_X1 U26880 ( .A1(n11945), .A2(n28197), .B(n5659), .ZN(n11943) );
  XOR2_X1 U26884 ( .A1(n19703), .A2(n25415), .Z(n12088) );
  NAND2_X2 U26885 ( .A1(n25747), .A2(n53226), .ZN(n25746) );
  BUF_X4 U26886 ( .I(n29991), .Z(n16961) );
  XOR2_X1 U26888 ( .A1(Key[189]), .A2(n7123), .Z(n28273) );
  NAND2_X1 U26891 ( .A1(n7886), .A2(n28381), .ZN(n28374) );
  XOR2_X1 U26893 ( .A1(Ciphertext[20]), .A2(Key[129]), .Z(n20716) );
  OR2_X2 U26896 ( .A1(n30159), .A2(n58999), .Z(n30165) );
  INV_X1 U26899 ( .I(n33096), .ZN(n32814) );
  XOR2_X1 U26903 ( .A1(n20623), .A2(n32226), .Z(n32227) );
  XOR2_X1 U26905 ( .A1(n23618), .A2(n7137), .Z(n44990) );
  XOR2_X1 U26910 ( .A1(n7141), .A2(n33273), .Z(n9665) );
  XOR2_X1 U26912 ( .A1(n7143), .A2(n11577), .Z(n51366) );
  XOR2_X1 U26913 ( .A1(n51933), .A2(n15735), .Z(n7143) );
  NOR3_X1 U26916 ( .A1(n49793), .A2(n10015), .A3(n49789), .ZN(n46008) );
  NAND2_X1 U26918 ( .A1(n54404), .A2(n54403), .ZN(n7151) );
  NAND2_X1 U26919 ( .A1(n54405), .A2(n7153), .ZN(n7152) );
  INV_X1 U26920 ( .I(n54403), .ZN(n7153) );
  INV_X4 U26923 ( .I(n15759), .ZN(n23331) );
  OAI21_X1 U26932 ( .A1(n9065), .A2(n55359), .B(n9238), .ZN(n55360) );
  INV_X1 U26935 ( .I(n5299), .ZN(n47308) );
  XOR2_X1 U26938 ( .A1(n46123), .A2(n10099), .Z(n7162) );
  XOR2_X1 U26939 ( .A1(n7163), .A2(n25975), .Z(n17097) );
  XOR2_X1 U26940 ( .A1(n25847), .A2(n7164), .Z(n7163) );
  NAND2_X2 U26942 ( .A1(n24075), .A2(n55401), .ZN(n55246) );
  XOR2_X1 U26943 ( .A1(n22350), .A2(n51197), .Z(n7166) );
  NOR3_X2 U26945 ( .A1(n21416), .A2(n21415), .A3(n7167), .ZN(n22959) );
  NAND4_X2 U26946 ( .A1(n16510), .A2(n16509), .A3(n45983), .A4(n45982), .ZN(
        n7167) );
  OAI21_X1 U26947 ( .A1(n7168), .A2(n36423), .B(n36121), .ZN(n35134) );
  NOR2_X2 U26949 ( .A1(n19646), .A2(n15220), .ZN(n49797) );
  XOR2_X1 U26950 ( .A1(n32369), .A2(n13570), .Z(n13569) );
  INV_X1 U26952 ( .I(n39902), .ZN(n18046) );
  NOR2_X2 U26959 ( .A1(n49195), .A2(n48845), .ZN(n11781) );
  XOR2_X1 U26960 ( .A1(n7178), .A2(n14161), .Z(n11538) );
  XOR2_X1 U26967 ( .A1(n7184), .A2(n56475), .Z(Plaintext[158]) );
  AND2_X1 U26968 ( .A1(n56474), .A2(n56512), .Z(n7185) );
  NAND2_X2 U26969 ( .A1(n53493), .A2(n23611), .ZN(n53525) );
  NAND2_X1 U26970 ( .A1(n23002), .A2(n30273), .ZN(n14396) );
  NAND3_X1 U26972 ( .A1(n16253), .A2(n23747), .A3(n22948), .ZN(n22378) );
  NAND2_X2 U26975 ( .A1(n22668), .A2(n24581), .ZN(n20337) );
  NAND3_X1 U26976 ( .A1(n34806), .A2(n36721), .A3(n34805), .ZN(n34808) );
  XOR2_X1 U26977 ( .A1(n7190), .A2(n51261), .Z(Plaintext[148]) );
  INV_X1 U26982 ( .I(n44182), .ZN(n21463) );
  INV_X2 U26983 ( .I(n14335), .ZN(n7587) );
  NAND2_X2 U26985 ( .A1(n24715), .A2(n24884), .ZN(n42759) );
  XOR2_X1 U26986 ( .A1(n7192), .A2(n51056), .Z(n56210) );
  NOR3_X1 U26991 ( .A1(n60510), .A2(n26223), .A3(n47356), .ZN(n20941) );
  NOR2_X1 U26994 ( .A1(n49255), .A2(n63876), .ZN(n45468) );
  XOR2_X1 U26997 ( .A1(n37145), .A2(n7195), .Z(n37146) );
  XOR2_X1 U26998 ( .A1(n21494), .A2(n17154), .Z(n7195) );
  NAND2_X1 U27005 ( .A1(n25712), .A2(n25708), .ZN(n42840) );
  INV_X4 U27013 ( .I(n18606), .ZN(n50123) );
  NAND2_X1 U27015 ( .A1(n21788), .A2(n21787), .ZN(n21786) );
  NOR2_X2 U27016 ( .A1(n47435), .A2(n9046), .ZN(n47737) );
  NAND2_X2 U27017 ( .A1(n8784), .A2(n51351), .ZN(n57014) );
  NOR4_X2 U27018 ( .A1(n27682), .A2(n27896), .A3(n27681), .A4(n27680), .ZN(
        n27686) );
  NAND2_X1 U27019 ( .A1(n22040), .A2(n22041), .ZN(n22039) );
  INV_X4 U27020 ( .I(n12539), .ZN(n12859) );
  BUF_X4 U27022 ( .I(n19507), .Z(n7598) );
  NAND2_X2 U27023 ( .A1(n16655), .A2(n16656), .ZN(n18129) );
  XOR2_X1 U27027 ( .A1(n8625), .A2(n32158), .Z(n31965) );
  AOI22_X1 U27033 ( .A1(n9561), .A2(n27392), .B1(n27391), .B2(n29150), .ZN(
        n27393) );
  XOR2_X1 U27034 ( .A1(n7216), .A2(n15001), .Z(n15078) );
  NOR2_X2 U27039 ( .A1(n52388), .A2(n7801), .ZN(n55151) );
  INV_X4 U27041 ( .I(n15227), .ZN(n26213) );
  OR2_X1 U27043 ( .A1(n52948), .A2(n55264), .Z(n8058) );
  INV_X1 U27052 ( .I(n62128), .ZN(n27958) );
  XOR2_X1 U27056 ( .A1(n7231), .A2(n50689), .Z(n13681) );
  XOR2_X1 U27057 ( .A1(n50694), .A2(n7232), .Z(n7231) );
  INV_X1 U27060 ( .I(n9066), .ZN(n55098) );
  OAI21_X1 U27061 ( .A1(n7235), .A2(n7234), .B(n24047), .ZN(n15383) );
  XOR2_X1 U27065 ( .A1(n18578), .A2(n37662), .Z(n7238) );
  AOI21_X1 U27066 ( .A1(n53782), .A2(n53783), .B(n7239), .ZN(n53784) );
  AND2_X1 U27067 ( .A1(n25879), .A2(n27534), .Z(n15423) );
  OAI22_X1 U27068 ( .A1(n28346), .A2(n18931), .B1(n24735), .B2(n23362), .ZN(
        n10010) );
  NOR2_X2 U27071 ( .A1(n17619), .A2(n17824), .ZN(n17343) );
  OAI22_X1 U27082 ( .A1(n7247), .A2(n10522), .B1(n54587), .B2(n44455), .ZN(
        n44459) );
  NAND2_X1 U27084 ( .A1(n35298), .A2(n20103), .ZN(n20102) );
  NOR3_X2 U27085 ( .A1(n18733), .A2(n1136), .A3(n7249), .ZN(n18478) );
  NOR2_X1 U27087 ( .A1(n13673), .A2(n40575), .ZN(n14622) );
  OAI21_X1 U27089 ( .A1(n10127), .A2(n1775), .B(n35604), .ZN(n33412) );
  INV_X4 U27090 ( .I(n22508), .ZN(n47803) );
  INV_X4 U27092 ( .I(n29566), .ZN(n11263) );
  NOR2_X1 U27093 ( .A1(n1425), .A2(n14464), .ZN(n14463) );
  OR4_X1 U27094 ( .A1(n36450), .A2(n36452), .A3(n23257), .A4(n9633), .Z(n11730) );
  NOR2_X1 U27095 ( .A1(n17362), .A2(n17361), .ZN(n17360) );
  XOR2_X1 U27096 ( .A1(n38777), .A2(n7263), .Z(n16052) );
  XOR2_X1 U27097 ( .A1(n6782), .A2(n36862), .Z(n7263) );
  NAND3_X1 U27098 ( .A1(n11688), .A2(n11686), .A3(n11687), .ZN(n11685) );
  BUF_X2 U27102 ( .I(n30968), .Z(n7264) );
  XOR2_X1 U27105 ( .A1(n7266), .A2(n44248), .Z(n44249) );
  XOR2_X1 U27106 ( .A1(n7267), .A2(n32202), .Z(n16366) );
  XOR2_X1 U27107 ( .A1(n32105), .A2(n32101), .Z(n7267) );
  OAI21_X1 U27112 ( .A1(n1971), .A2(n29706), .B(n29705), .ZN(n29707) );
  NAND2_X1 U27114 ( .A1(n12499), .A2(n10508), .ZN(n25345) );
  NAND3_X2 U27116 ( .A1(n15304), .A2(n57026), .A3(n15435), .ZN(n57018) );
  AND2_X1 U27120 ( .A1(n56594), .A2(n56595), .Z(n7277) );
  OR3_X1 U27122 ( .A1(n60397), .A2(n50307), .A3(n3055), .Z(n50310) );
  NOR2_X1 U27123 ( .A1(n47632), .A2(n13054), .ZN(n47641) );
  AND2_X2 U27124 ( .A1(n26228), .A2(n21276), .Z(n14056) );
  AND2_X2 U27129 ( .A1(n35756), .A2(n11981), .Z(n10503) );
  INV_X4 U27132 ( .I(n7283), .ZN(n20391) );
  OR2_X1 U27135 ( .A1(n12797), .A2(n12798), .Z(n7284) );
  OAI21_X1 U27136 ( .A1(n7287), .A2(n7286), .B(n45006), .ZN(n14411) );
  NOR2_X1 U27137 ( .A1(n22468), .A2(n1069), .ZN(n7287) );
  XOR2_X1 U27144 ( .A1(n7292), .A2(n50610), .Z(n50613) );
  XOR2_X1 U27148 ( .A1(n16814), .A2(n7295), .Z(n16813) );
  XOR2_X1 U27149 ( .A1(n50768), .A2(n8856), .Z(n7295) );
  NAND2_X2 U27151 ( .A1(n35816), .A2(n34316), .ZN(n25389) );
  NOR2_X2 U27152 ( .A1(n1741), .A2(n20552), .ZN(n42252) );
  BUF_X2 U27160 ( .I(n53415), .Z(n7303) );
  INV_X4 U27161 ( .I(n25204), .ZN(n40713) );
  XOR2_X1 U27165 ( .A1(n1411), .A2(n38523), .Z(n16561) );
  XOR2_X1 U27166 ( .A1(n14550), .A2(n24533), .Z(n38523) );
  NOR2_X2 U27169 ( .A1(n42257), .A2(n7304), .ZN(n44227) );
  NAND3_X2 U27170 ( .A1(n42254), .A2(n42256), .A3(n7305), .ZN(n7304) );
  AND2_X1 U27171 ( .A1(n42253), .A2(n42255), .Z(n7305) );
  AND2_X1 U27174 ( .A1(n48422), .A2(n18469), .Z(n16047) );
  OAI22_X1 U27176 ( .A1(n54724), .A2(n7307), .B1(n54709), .B2(n54752), .ZN(
        n54679) );
  NAND2_X1 U27189 ( .A1(n23993), .A2(n20566), .ZN(n20565) );
  NAND2_X1 U27190 ( .A1(n20498), .A2(n20497), .ZN(n20496) );
  XOR2_X1 U27191 ( .A1(n7313), .A2(n33163), .Z(n33215) );
  NAND2_X1 U27192 ( .A1(n18343), .A2(n1042), .ZN(n18020) );
  XOR2_X1 U27194 ( .A1(n7315), .A2(n9609), .Z(n33160) );
  XOR2_X1 U27195 ( .A1(n9254), .A2(n46684), .Z(n7315) );
  NAND3_X1 U27196 ( .A1(n10010), .A2(n4998), .A3(n27533), .ZN(n25879) );
  XOR2_X1 U27202 ( .A1(n19189), .A2(n24040), .Z(n7320) );
  NOR2_X1 U27203 ( .A1(n43870), .A2(n43869), .ZN(n11068) );
  NOR2_X1 U27204 ( .A1(n11068), .A2(n11067), .ZN(n10557) );
  NAND3_X1 U27207 ( .A1(n25646), .A2(n7324), .A3(n25645), .ZN(n22630) );
  OAI21_X1 U27208 ( .A1(n7437), .A2(n26964), .B(n26963), .ZN(n7324) );
  NAND2_X1 U27213 ( .A1(n12581), .A2(n50381), .ZN(n9487) );
  NAND2_X2 U27217 ( .A1(n25214), .A2(n54292), .ZN(n54798) );
  NAND2_X1 U27218 ( .A1(n14746), .A2(n28118), .ZN(n8710) );
  OAI21_X1 U27219 ( .A1(n9407), .A2(n22379), .B(n56627), .ZN(n7333) );
  NOR2_X2 U27224 ( .A1(n25858), .A2(n26834), .ZN(n28507) );
  OR2_X1 U27226 ( .A1(n29158), .A2(n820), .Z(n26379) );
  NOR2_X2 U27227 ( .A1(n43626), .A2(n57810), .ZN(n43633) );
  AND2_X1 U27230 ( .A1(n63220), .A2(n34433), .Z(n26229) );
  OR2_X1 U27234 ( .A1(n45984), .A2(n64470), .Z(n45986) );
  XOR2_X1 U27235 ( .A1(n7340), .A2(n7341), .Z(n7842) );
  NOR2_X1 U27238 ( .A1(n55020), .A2(n61472), .ZN(n7346) );
  XOR2_X1 U27243 ( .A1(n44990), .A2(n44989), .Z(n11358) );
  XOR2_X1 U27245 ( .A1(n24798), .A2(n1674), .Z(n22725) );
  AND2_X1 U27247 ( .A1(n38273), .A2(n60587), .Z(n41800) );
  INV_X1 U27251 ( .I(n48823), .ZN(n11290) );
  XOR2_X1 U27252 ( .A1(n16909), .A2(n10076), .Z(n44119) );
  NOR2_X2 U27255 ( .A1(n1541), .A2(n34414), .ZN(n18834) );
  NAND3_X1 U27256 ( .A1(n55498), .A2(n55300), .A3(n55303), .ZN(n52049) );
  INV_X2 U27258 ( .I(n7352), .ZN(n16936) );
  NOR2_X1 U27261 ( .A1(n18070), .A2(n11024), .ZN(n32804) );
  INV_X1 U27264 ( .I(n24376), .ZN(n15497) );
  XOR2_X1 U27266 ( .A1(n7360), .A2(n32514), .Z(n21866) );
  XOR2_X1 U27267 ( .A1(n30715), .A2(n7361), .Z(n7360) );
  XOR2_X1 U27268 ( .A1(n32587), .A2(n31585), .Z(n7362) );
  NOR2_X1 U27272 ( .A1(n29703), .A2(n22648), .ZN(n7363) );
  INV_X4 U27280 ( .I(n14199), .ZN(n19329) );
  OR2_X1 U27284 ( .A1(n28300), .A2(n27179), .Z(n12280) );
  AND2_X1 U27289 ( .A1(n7710), .A2(n34395), .Z(n35234) );
  XOR2_X1 U27290 ( .A1(n7375), .A2(n57162), .Z(Plaintext[191]) );
  NOR3_X2 U27291 ( .A1(n57055), .A2(n57054), .A3(n57056), .ZN(n57109) );
  XOR2_X1 U27292 ( .A1(n7377), .A2(n33170), .Z(n23590) );
  XOR2_X1 U27298 ( .A1(n25421), .A2(n39661), .Z(n25420) );
  XOR2_X1 U27305 ( .A1(n7685), .A2(n1674), .Z(n7385) );
  AND2_X1 U27309 ( .A1(n12188), .A2(n12187), .Z(n11854) );
  NAND2_X1 U27311 ( .A1(n31782), .A2(n10494), .ZN(n31783) );
  INV_X4 U27312 ( .I(n53532), .ZN(n13370) );
  NOR2_X2 U27317 ( .A1(n18637), .A2(n18634), .ZN(n17913) );
  XOR2_X1 U27320 ( .A1(n16884), .A2(n1550), .Z(n7390) );
  NOR2_X2 U27321 ( .A1(n14518), .A2(n48460), .ZN(n47079) );
  NOR2_X1 U27324 ( .A1(n26179), .A2(n20023), .ZN(n19919) );
  NAND2_X2 U27326 ( .A1(n9201), .A2(n9202), .ZN(n42598) );
  XOR2_X1 U27328 ( .A1(n32077), .A2(n17026), .Z(n7394) );
  XOR2_X1 U27329 ( .A1(n1213), .A2(n17934), .Z(n17933) );
  NAND2_X1 U27331 ( .A1(n56078), .A2(n56079), .ZN(Plaintext[141]) );
  NAND2_X1 U27332 ( .A1(n56060), .A2(n1184), .ZN(n56077) );
  XOR2_X1 U27333 ( .A1(n20057), .A2(n20056), .Z(n9755) );
  XOR2_X1 U27336 ( .A1(n25165), .A2(n7396), .Z(n25164) );
  XOR2_X1 U27337 ( .A1(n17875), .A2(n7397), .Z(n7396) );
  XOR2_X1 U27338 ( .A1(n7398), .A2(n16983), .Z(n17133) );
  NOR2_X1 U27345 ( .A1(n9481), .A2(n9480), .ZN(n19674) );
  NOR2_X2 U27348 ( .A1(n20372), .A2(n62530), .ZN(n42620) );
  AND2_X1 U27351 ( .A1(n58907), .A2(n25128), .Z(n16157) );
  XOR2_X1 U27354 ( .A1(n52026), .A2(n7743), .Z(n9062) );
  AOI21_X1 U27361 ( .A1(n55827), .A2(n20710), .B(n12434), .ZN(n12433) );
  NAND2_X2 U27365 ( .A1(n34585), .A2(n15809), .ZN(n34185) );
  XOR2_X1 U27367 ( .A1(n13458), .A2(n25376), .Z(n38877) );
  NAND2_X2 U27368 ( .A1(n16533), .A2(n47490), .ZN(n48209) );
  XOR2_X1 U27369 ( .A1(n21985), .A2(n30354), .Z(n27008) );
  XOR2_X1 U27372 ( .A1(n7417), .A2(n27630), .Z(n33519) );
  NAND2_X1 U27378 ( .A1(n7463), .A2(n7462), .ZN(n8825) );
  XOR2_X1 U27380 ( .A1(n50693), .A2(n51548), .Z(n50694) );
  NAND3_X2 U27386 ( .A1(n18979), .A2(n47741), .A3(n47740), .ZN(n18978) );
  NOR2_X1 U27394 ( .A1(n55472), .A2(n55478), .ZN(n7894) );
  NAND2_X2 U27398 ( .A1(n12131), .A2(n29201), .ZN(n30844) );
  NAND2_X2 U27403 ( .A1(n43679), .A2(n65203), .ZN(n43564) );
  INV_X2 U27406 ( .I(n31710), .ZN(n33663) );
  NAND3_X2 U27410 ( .A1(n40029), .A2(n4364), .A3(n40304), .ZN(n40226) );
  NAND2_X1 U27417 ( .A1(n22825), .A2(n22824), .ZN(n52496) );
  INV_X2 U27419 ( .I(n7439), .ZN(n14624) );
  INV_X2 U27421 ( .I(n25085), .ZN(n52861) );
  NOR2_X2 U27422 ( .A1(n34132), .A2(n157), .ZN(n34142) );
  NAND2_X1 U27424 ( .A1(n13126), .A2(n34288), .ZN(n34815) );
  NAND2_X1 U27427 ( .A1(n7441), .A2(n18179), .ZN(n33556) );
  OAI22_X1 U27428 ( .A1(n33546), .A2(n33547), .B1(n33549), .B2(n33548), .ZN(
        n7441) );
  XOR2_X1 U27429 ( .A1(n39348), .A2(n39643), .Z(n10781) );
  XOR2_X1 U27431 ( .A1(n7442), .A2(n58740), .Z(n44970) );
  XOR2_X1 U27433 ( .A1(n1436), .A2(n1435), .Z(n7444) );
  AOI21_X1 U27436 ( .A1(n7445), .A2(n56438), .B(n61368), .ZN(n56439) );
  NAND2_X1 U27437 ( .A1(n56437), .A2(n9022), .ZN(n7445) );
  NOR3_X2 U27443 ( .A1(n20474), .A2(n20863), .A3(n15159), .ZN(n15029) );
  NOR2_X1 U27444 ( .A1(n17564), .A2(n17563), .ZN(n17562) );
  XOR2_X1 U27446 ( .A1(n38817), .A2(n927), .Z(n12545) );
  XOR2_X1 U27448 ( .A1(n31293), .A2(n7456), .Z(n31294) );
  XOR2_X1 U27449 ( .A1(n22734), .A2(n8625), .Z(n7456) );
  XOR2_X1 U27451 ( .A1(n60528), .A2(n33144), .Z(n8884) );
  NAND2_X2 U27454 ( .A1(n56255), .A2(n7274), .ZN(n56582) );
  INV_X4 U27455 ( .I(n7767), .ZN(n8361) );
  INV_X1 U27458 ( .I(n28202), .ZN(n11949) );
  INV_X1 U27460 ( .I(n54952), .ZN(n7654) );
  NAND2_X2 U27462 ( .A1(n45940), .A2(n45939), .ZN(n47347) );
  XOR2_X1 U27470 ( .A1(n8805), .A2(n51343), .Z(n51689) );
  OR2_X2 U27472 ( .A1(n8794), .A2(n46148), .Z(n48189) );
  NAND2_X1 U27473 ( .A1(n55244), .A2(n54978), .ZN(n7469) );
  AND3_X1 U27475 ( .A1(n56957), .A2(n56967), .A3(n56959), .Z(n9653) );
  NAND3_X1 U27480 ( .A1(n1394), .A2(n42692), .A3(n42697), .ZN(n42708) );
  NAND3_X2 U27485 ( .A1(n54728), .A2(n22122), .A3(n22385), .ZN(n54724) );
  AND2_X1 U27489 ( .A1(n13909), .A2(n41173), .Z(n24882) );
  OAI21_X1 U27490 ( .A1(n24985), .A2(n40092), .B(n10801), .ZN(n40130) );
  OR2_X1 U27491 ( .A1(n1777), .A2(n35508), .Z(n7483) );
  NAND3_X1 U27493 ( .A1(n40086), .A2(n39887), .A3(n25246), .ZN(n39412) );
  INV_X1 U27494 ( .I(n47996), .ZN(n10889) );
  NOR3_X1 U27495 ( .A1(n53768), .A2(n53766), .A3(n53767), .ZN(n7486) );
  INV_X2 U27498 ( .I(n7487), .ZN(n46262) );
  XOR2_X1 U27499 ( .A1(n18065), .A2(n18066), .Z(n7487) );
  INV_X2 U27500 ( .I(n7489), .ZN(n15093) );
  XOR2_X1 U27501 ( .A1(Ciphertext[72]), .A2(Key[109]), .Z(n7489) );
  XOR2_X1 U27502 ( .A1(n32163), .A2(n31550), .Z(n31612) );
  INV_X2 U27503 ( .I(n19491), .ZN(n54728) );
  AND3_X1 U27506 ( .A1(n18918), .A2(n49547), .A3(n49170), .Z(n48278) );
  INV_X4 U27508 ( .I(n12725), .ZN(n20912) );
  NOR3_X2 U27512 ( .A1(n29365), .A2(n29363), .A3(n29364), .ZN(n29392) );
  INV_X1 U27517 ( .I(n17708), .ZN(n8489) );
  XOR2_X1 U27518 ( .A1(n7496), .A2(n63487), .Z(n8294) );
  XOR2_X1 U27519 ( .A1(n39626), .A2(n53641), .Z(n7496) );
  NOR2_X1 U27521 ( .A1(n7692), .A2(n20941), .ZN(n13259) );
  NAND2_X2 U27522 ( .A1(n53823), .A2(n15928), .ZN(n53793) );
  XOR2_X1 U27529 ( .A1(n7508), .A2(n53642), .Z(Plaintext[30]) );
  NOR4_X1 U27530 ( .A1(n53638), .A2(n53640), .A3(n53639), .A4(n53648), .ZN(
        n7508) );
  XOR2_X1 U27532 ( .A1(n5244), .A2(n18999), .Z(n7509) );
  XOR2_X1 U27533 ( .A1(n7510), .A2(n15672), .Z(n26105) );
  NAND2_X2 U27537 ( .A1(n10747), .A2(n8889), .ZN(n8948) );
  NAND2_X1 U27538 ( .A1(n41170), .A2(n13510), .ZN(n7870) );
  INV_X1 U27541 ( .I(n18348), .ZN(n36484) );
  XOR2_X1 U27543 ( .A1(n32665), .A2(n7512), .Z(n20081) );
  XOR2_X1 U27544 ( .A1(n31926), .A2(n59546), .Z(n7512) );
  AND2_X1 U27545 ( .A1(n7775), .A2(n28036), .Z(n15985) );
  NOR2_X1 U27547 ( .A1(n7515), .A2(n7514), .ZN(n7513) );
  NOR2_X1 U27548 ( .A1(n43899), .A2(n7516), .ZN(n7515) );
  OAI21_X1 U27549 ( .A1(n61394), .A2(n41951), .B(n59280), .ZN(n7928) );
  AND2_X1 U27552 ( .A1(n16373), .A2(n838), .Z(n15983) );
  INV_X2 U27554 ( .I(n18478), .ZN(n22940) );
  NOR2_X1 U27555 ( .A1(n14677), .A2(n747), .ZN(n10288) );
  NOR2_X1 U27556 ( .A1(n15897), .A2(n19562), .ZN(n19460) );
  AND2_X1 U27557 ( .A1(n7735), .A2(n20960), .Z(n21404) );
  OAI21_X2 U27559 ( .A1(n1113), .A2(n18813), .B(n49540), .ZN(n18815) );
  AND2_X1 U27561 ( .A1(n27179), .A2(n23840), .Z(n24877) );
  XOR2_X1 U27563 ( .A1(n7525), .A2(n54587), .Z(Plaintext[77]) );
  XOR2_X1 U27564 ( .A1(n45293), .A2(n9259), .Z(n9258) );
  NAND2_X1 U27573 ( .A1(n51443), .A2(n51444), .ZN(n51445) );
  INV_X1 U27575 ( .I(n48540), .ZN(n48118) );
  BUF_X2 U27576 ( .I(n11501), .Z(n7528) );
  BUF_X2 U27578 ( .I(n15815), .Z(n7531) );
  NAND4_X1 U27583 ( .A1(n35654), .A2(n33275), .A3(n33274), .A4(n35656), .ZN(
        n21046) );
  INV_X4 U27586 ( .I(n40443), .ZN(n25358) );
  XOR2_X1 U27591 ( .A1(n33070), .A2(n32035), .Z(n7535) );
  NAND2_X2 U27592 ( .A1(n54938), .A2(n21877), .ZN(n22544) );
  AOI21_X2 U27593 ( .A1(n14619), .A2(n57233), .B(n57124), .ZN(n57104) );
  NOR2_X2 U27594 ( .A1(n23940), .A2(n13672), .ZN(n11073) );
  XOR2_X1 U27597 ( .A1(n7540), .A2(n7539), .Z(n8249) );
  XOR2_X1 U27608 ( .A1(n7551), .A2(n8498), .Z(n19518) );
  XOR2_X1 U27609 ( .A1(n8497), .A2(n35957), .Z(n7551) );
  XOR2_X1 U27610 ( .A1(n44188), .A2(n7552), .Z(n7685) );
  NOR3_X2 U27613 ( .A1(n55180), .A2(n55179), .A3(n55178), .ZN(n55189) );
  OAI21_X1 U27615 ( .A1(n30411), .A2(n30412), .B(n30410), .ZN(n7556) );
  BUF_X2 U27616 ( .I(n10229), .Z(n7557) );
  NOR2_X1 U27617 ( .A1(n32679), .A2(n33323), .ZN(n32690) );
  AND3_X2 U27620 ( .A1(n46933), .A2(n46935), .A3(n46934), .Z(n18364) );
  NAND3_X1 U27621 ( .A1(n17971), .A2(n40619), .A3(n40618), .ZN(n15427) );
  NOR2_X2 U27624 ( .A1(n48612), .A2(n8639), .ZN(n48623) );
  XOR2_X1 U27626 ( .A1(n14671), .A2(n22434), .Z(n24519) );
  NOR2_X2 U27629 ( .A1(n28633), .A2(n27823), .ZN(n7561) );
  XOR2_X1 U27631 ( .A1(Ciphertext[147]), .A2(Key[154]), .Z(n7564) );
  NAND2_X2 U27633 ( .A1(n13234), .A2(n7567), .ZN(n16528) );
  XNOR2_X1 U27635 ( .A1(n51761), .A2(n51760), .ZN(n9704) );
  XNOR2_X1 U27636 ( .A1(n45429), .A2(n43946), .ZN(n14889) );
  INV_X2 U27641 ( .I(n7574), .ZN(n45682) );
  OR2_X2 U27642 ( .A1(n990), .A2(n11090), .Z(n10044) );
  XOR2_X1 U27645 ( .A1(n7575), .A2(n23464), .Z(n18971) );
  NAND3_X2 U27648 ( .A1(n47641), .A2(n47639), .A3(n47640), .ZN(n10472) );
  XOR2_X1 U27649 ( .A1(n7581), .A2(n55150), .Z(Plaintext[100]) );
  XOR2_X1 U27652 ( .A1(n2960), .A2(n8900), .Z(n8899) );
  NAND2_X1 U27654 ( .A1(n1383), .A2(n61362), .ZN(n7586) );
  NOR2_X1 U27655 ( .A1(n50211), .A2(n7588), .ZN(n47222) );
  NOR2_X1 U27656 ( .A1(n49100), .A2(n64751), .ZN(n18081) );
  OAI22_X1 U27658 ( .A1(n1890), .A2(n28400), .B1(n28414), .B2(n3117), .ZN(
        n26256) );
  XOR2_X1 U27660 ( .A1(n7589), .A2(n39732), .Z(n14144) );
  XOR2_X1 U27661 ( .A1(n7589), .A2(n38666), .Z(n38667) );
  NAND3_X2 U27662 ( .A1(n34705), .A2(n34706), .A3(n34704), .ZN(n7589) );
  NAND2_X2 U27665 ( .A1(n22798), .A2(n26159), .ZN(n7595) );
  NOR2_X1 U27666 ( .A1(n7596), .A2(n31277), .ZN(n30510) );
  INV_X2 U27670 ( .I(n61714), .ZN(n24359) );
  NOR2_X1 U27672 ( .A1(n43990), .A2(n1706), .ZN(n43718) );
  NAND2_X2 U27675 ( .A1(n9137), .A2(n10938), .ZN(n51716) );
  OAI21_X1 U27676 ( .A1(n22796), .A2(n1846), .B(n7604), .ZN(n7603) );
  INV_X2 U27678 ( .I(n7607), .ZN(n10969) );
  NAND2_X2 U27682 ( .A1(n15815), .A2(n24571), .ZN(n35646) );
  NAND3_X1 U27687 ( .A1(n7616), .A2(n15527), .A3(n15530), .ZN(n7888) );
  XOR2_X1 U27688 ( .A1(n19993), .A2(n1897), .Z(n32632) );
  XOR2_X1 U27689 ( .A1(n7616), .A2(n2952), .Z(n30797) );
  INV_X4 U27694 ( .I(n30730), .ZN(n23317) );
  NAND3_X2 U27696 ( .A1(n24823), .A2(n27458), .A3(n27459), .ZN(n30730) );
  NOR2_X2 U27698 ( .A1(n58598), .A2(n15815), .ZN(n33589) );
  INV_X1 U27699 ( .I(n39482), .ZN(n14645) );
  XOR2_X1 U27700 ( .A1(n7626), .A2(n1830), .Z(n8263) );
  XOR2_X1 U27701 ( .A1(n7627), .A2(n32026), .Z(n7626) );
  XOR2_X1 U27705 ( .A1(n62065), .A2(n46163), .Z(n7628) );
  INV_X2 U27706 ( .I(n41462), .ZN(n40712) );
  NOR2_X2 U27707 ( .A1(n4819), .A2(n17382), .ZN(n41462) );
  XOR2_X1 U27711 ( .A1(n7635), .A2(n7633), .Z(n16666) );
  XOR2_X1 U27712 ( .A1(n20448), .A2(n7634), .Z(n7633) );
  NAND2_X2 U27716 ( .A1(n10315), .A2(n22539), .ZN(n52424) );
  XOR2_X1 U27718 ( .A1(n10899), .A2(n24912), .Z(n7639) );
  XOR2_X1 U27720 ( .A1(n38718), .A2(n21299), .Z(n38630) );
  OAI22_X1 U27723 ( .A1(n40609), .A2(n40605), .B1(n40603), .B2(n60957), .ZN(
        n39119) );
  INV_X2 U27725 ( .I(n7642), .ZN(n8225) );
  XOR2_X1 U27728 ( .A1(n59854), .A2(n52439), .Z(n8066) );
  INV_X2 U27732 ( .I(n7650), .ZN(n22498) );
  INV_X2 U27733 ( .I(n22709), .ZN(n7651) );
  INV_X2 U27734 ( .I(n28526), .ZN(n28543) );
  XNOR2_X1 U27736 ( .A1(Ciphertext[99]), .A2(Key[10]), .ZN(n7650) );
  NOR3_X2 U27737 ( .A1(n7653), .A2(n48824), .A3(n10469), .ZN(n12604) );
  NAND2_X1 U27738 ( .A1(n7654), .A2(n54951), .ZN(n52385) );
  NAND2_X1 U27739 ( .A1(n7654), .A2(n54436), .ZN(n52957) );
  NAND2_X1 U27740 ( .A1(n7654), .A2(n60439), .ZN(n54782) );
  XOR2_X1 U27743 ( .A1(n2952), .A2(n32494), .Z(n7658) );
  INV_X2 U27744 ( .I(n29991), .ZN(n29820) );
  NAND2_X2 U27745 ( .A1(n28080), .A2(n28079), .ZN(n29991) );
  XOR2_X1 U27746 ( .A1(n62502), .A2(n1761), .Z(n38818) );
  OAI22_X1 U27747 ( .A1(n7662), .A2(n37090), .B1(n37940), .B2(n59825), .ZN(
        n37094) );
  AOI21_X1 U27748 ( .A1(n37316), .A2(n7662), .B(n37315), .ZN(n37317) );
  XOR2_X1 U27749 ( .A1(n7663), .A2(n9429), .Z(n9428) );
  NAND3_X2 U27754 ( .A1(n17835), .A2(n17834), .A3(n23271), .ZN(n52041) );
  INV_X2 U27755 ( .I(n52041), .ZN(n11789) );
  NAND2_X1 U27757 ( .A1(n15759), .A2(n4428), .ZN(n47132) );
  NAND4_X2 U27759 ( .A1(n7677), .A2(n41327), .A3(n41321), .A4(n25795), .ZN(
        n44834) );
  XOR2_X1 U27762 ( .A1(n45041), .A2(n7679), .Z(n44219) );
  XOR2_X1 U27763 ( .A1(n7679), .A2(n21463), .Z(n8108) );
  NAND2_X2 U27764 ( .A1(n8081), .A2(n8080), .ZN(n7679) );
  INV_X2 U27768 ( .I(n46912), .ZN(n45765) );
  INV_X2 U27770 ( .I(n17776), .ZN(n34627) );
  XOR2_X1 U27772 ( .A1(n38367), .A2(n1411), .Z(n7687) );
  XOR2_X1 U27774 ( .A1(n21891), .A2(n38263), .Z(n7688) );
  XOR2_X1 U27775 ( .A1(n38180), .A2(n7689), .Z(n38263) );
  INV_X1 U27776 ( .I(n22321), .ZN(n7689) );
  XOR2_X1 U27778 ( .A1(n14589), .A2(n18428), .Z(n24184) );
  XOR2_X1 U27779 ( .A1(n59370), .A2(n7691), .Z(n7997) );
  NOR2_X2 U27782 ( .A1(n8195), .A2(n1235), .ZN(n36329) );
  OAI21_X1 U27784 ( .A1(n36828), .A2(n1235), .B(n36827), .ZN(n36833) );
  INV_X1 U27785 ( .I(n20047), .ZN(n7694) );
  AOI21_X1 U27786 ( .A1(n7697), .A2(n54460), .B(n54858), .ZN(n52642) );
  OAI22_X1 U27788 ( .A1(n54637), .A2(n7697), .B1(n62760), .B2(n59713), .ZN(
        n54639) );
  OAI21_X1 U27790 ( .A1(n32965), .A2(n5529), .B(n1537), .ZN(n11652) );
  NAND2_X1 U27791 ( .A1(n8552), .A2(n5529), .ZN(n21811) );
  XOR2_X1 U27793 ( .A1(n63016), .A2(n8865), .Z(n7702) );
  XOR2_X1 U27795 ( .A1(n1051), .A2(n8862), .Z(n7703) );
  NAND2_X1 U27800 ( .A1(n34406), .A2(n7710), .ZN(n34407) );
  AOI22_X1 U27801 ( .A1(n34394), .A2(n35224), .B1(n7710), .B2(n35713), .ZN(
        n34398) );
  XOR2_X1 U27804 ( .A1(n7711), .A2(n18492), .Z(n18491) );
  XOR2_X1 U27806 ( .A1(n18340), .A2(n22277), .Z(n37888) );
  NOR2_X1 U27808 ( .A1(n21949), .A2(n7719), .ZN(n7718) );
  NAND2_X1 U27810 ( .A1(n43351), .A2(n7720), .ZN(n43354) );
  OAI21_X2 U27812 ( .A1(n7725), .A2(n7724), .B(n7722), .ZN(n16120) );
  NAND2_X2 U27815 ( .A1(n3348), .A2(n20428), .ZN(n20311) );
  XOR2_X1 U27816 ( .A1(n38457), .A2(n20032), .Z(n19991) );
  NOR2_X2 U27821 ( .A1(n61729), .A2(n22903), .ZN(n12420) );
  XOR2_X1 U27823 ( .A1(n7743), .A2(n50915), .Z(n8955) );
  NOR2_X2 U27831 ( .A1(n7757), .A2(n7756), .ZN(n8110) );
  NAND2_X2 U27832 ( .A1(n8963), .A2(n7758), .ZN(n7757) );
  NOR2_X2 U27833 ( .A1(n49389), .A2(n49395), .ZN(n49213) );
  NAND2_X1 U27834 ( .A1(n65224), .A2(n9256), .ZN(n19989) );
  NAND2_X1 U27835 ( .A1(n47468), .A2(n65224), .ZN(n9175) );
  XOR2_X1 U27837 ( .A1(n51591), .A2(n51249), .Z(n7761) );
  NAND2_X2 U27839 ( .A1(n4819), .A2(n17382), .ZN(n25777) );
  XOR2_X1 U27840 ( .A1(n45237), .A2(n7768), .Z(n44021) );
  XOR2_X1 U27841 ( .A1(n7769), .A2(n46288), .Z(n7768) );
  XOR2_X1 U27842 ( .A1(n43764), .A2(n785), .Z(n7769) );
  NAND4_X2 U27843 ( .A1(n15636), .A2(n15638), .A3(n43315), .A4(n43314), .ZN(
        n45019) );
  XOR2_X1 U27845 ( .A1(n59701), .A2(n33153), .Z(n7773) );
  OAI21_X2 U27847 ( .A1(n16961), .A2(n29993), .B(n29994), .ZN(n7774) );
  NAND2_X1 U27848 ( .A1(n28032), .A2(n7775), .ZN(n26578) );
  NAND2_X1 U27849 ( .A1(n27052), .A2(n7775), .ZN(n27053) );
  OAI22_X1 U27850 ( .A1(n23498), .A2(n26581), .B1(n28233), .B2(n7775), .ZN(
        n23938) );
  NAND2_X2 U27851 ( .A1(n3932), .A2(n20753), .ZN(n7775) );
  INV_X2 U27853 ( .I(n7452), .ZN(n22043) );
  XOR2_X1 U27855 ( .A1(n46591), .A2(n11014), .Z(n7778) );
  NOR2_X2 U27860 ( .A1(n34566), .A2(n32295), .ZN(n34958) );
  OAI21_X1 U27862 ( .A1(n48487), .A2(n48488), .B(n60232), .ZN(n48489) );
  NAND3_X1 U27863 ( .A1(n48590), .A2(n48591), .A3(n64634), .ZN(n48592) );
  NAND2_X1 U27866 ( .A1(n20832), .A2(n7799), .ZN(n20831) );
  AOI22_X1 U27867 ( .A1(n24217), .A2(n41947), .B1(n41803), .B2(n59280), .ZN(
        n17296) );
  NAND2_X2 U27871 ( .A1(n26119), .A2(n26117), .ZN(n55133) );
  INV_X2 U27872 ( .I(n35882), .ZN(n35887) );
  INV_X2 U27873 ( .I(n7810), .ZN(n7811) );
  XOR2_X1 U27875 ( .A1(n46626), .A2(n46436), .Z(n23345) );
  XOR2_X1 U27876 ( .A1(n46440), .A2(n46441), .Z(n46626) );
  AOI21_X2 U27877 ( .A1(n2722), .A2(n14536), .B(n61670), .ZN(n46440) );
  OR2_X1 U27878 ( .A1(n48467), .A2(n48134), .Z(n8137) );
  XOR2_X1 U27880 ( .A1(n15102), .A2(n7823), .Z(n15017) );
  XOR2_X1 U27881 ( .A1(n13449), .A2(n31848), .Z(n7823) );
  XOR2_X1 U27882 ( .A1(Ciphertext[106]), .A2(Key[155]), .Z(n9556) );
  NAND3_X2 U27885 ( .A1(n7827), .A2(n42153), .A3(n7830), .ZN(n7826) );
  NAND2_X1 U27891 ( .A1(n48514), .A2(n7834), .ZN(n21689) );
  NAND2_X1 U27893 ( .A1(n48494), .A2(n7834), .ZN(n46566) );
  NAND2_X2 U27894 ( .A1(n1212), .A2(n11380), .ZN(n7834) );
  INV_X2 U27895 ( .I(n15536), .ZN(n7836) );
  INV_X2 U27896 ( .I(n15536), .ZN(n56990) );
  OAI22_X1 U27897 ( .A1(n33000), .A2(n33613), .B1(n9085), .B2(n5082), .ZN(
        n7841) );
  INV_X2 U27898 ( .I(n7842), .ZN(n51191) );
  OR2_X1 U27900 ( .A1(n25777), .A2(n1507), .Z(n7845) );
  NOR2_X2 U27903 ( .A1(n16766), .A2(n7846), .ZN(n50215) );
  NAND2_X1 U27904 ( .A1(n50209), .A2(n7336), .ZN(n49100) );
  NOR2_X1 U27905 ( .A1(n10889), .A2(n7336), .ZN(n47992) );
  NAND2_X2 U27906 ( .A1(n11390), .A2(n47221), .ZN(n7846) );
  XOR2_X1 U27907 ( .A1(n58989), .A2(n23878), .Z(n52374) );
  NOR2_X1 U27910 ( .A1(n7849), .A2(n33984), .ZN(n33979) );
  NAND2_X1 U27911 ( .A1(n7849), .A2(n34042), .ZN(n34044) );
  OAI22_X1 U27912 ( .A1(n34036), .A2(n7849), .B1(n34603), .B2(n60763), .ZN(
        n34037) );
  XOR2_X1 U27913 ( .A1(n7850), .A2(n45016), .Z(n45018) );
  XOR2_X1 U27916 ( .A1(n7853), .A2(n36647), .Z(n39565) );
  XOR2_X1 U27917 ( .A1(n61279), .A2(n7578), .Z(n30992) );
  XOR2_X1 U27918 ( .A1(n31431), .A2(n7578), .Z(n8506) );
  OAI21_X2 U27920 ( .A1(n31305), .A2(n36605), .B(n35100), .ZN(n36609) );
  XOR2_X1 U27924 ( .A1(n15500), .A2(n7863), .Z(n14085) );
  XOR2_X1 U27925 ( .A1(n7864), .A2(n38645), .Z(n7863) );
  XOR2_X1 U27926 ( .A1(n37285), .A2(n52206), .Z(n7864) );
  NAND2_X1 U27929 ( .A1(n7868), .A2(n60622), .ZN(n50237) );
  NOR2_X1 U27932 ( .A1(n5258), .A2(n7866), .ZN(n7867) );
  NOR3_X2 U27933 ( .A1(n50444), .A2(n50019), .A3(n7868), .ZN(n50448) );
  OAI22_X1 U27934 ( .A1(n50231), .A2(n7868), .B1(n50232), .B2(n25966), .ZN(
        n23372) );
  NAND2_X2 U27937 ( .A1(n6705), .A2(n42681), .ZN(n42149) );
  NOR2_X2 U27938 ( .A1(n7870), .A2(n7869), .ZN(n42681) );
  XOR2_X1 U27939 ( .A1(n7871), .A2(n31383), .Z(n9587) );
  XOR2_X1 U27940 ( .A1(n7872), .A2(n31384), .Z(n7871) );
  XOR2_X1 U27941 ( .A1(n9179), .A2(n9483), .Z(n31384) );
  AND2_X1 U27945 ( .A1(n55149), .A2(n55154), .Z(n7875) );
  INV_X1 U27946 ( .I(n21390), .ZN(n7876) );
  XOR2_X1 U27950 ( .A1(n7880), .A2(n7881), .Z(n7879) );
  XOR2_X1 U27951 ( .A1(n10555), .A2(n43795), .Z(n7881) );
  INV_X2 U27954 ( .I(n7885), .ZN(n24368) );
  INV_X2 U27956 ( .I(n26035), .ZN(n8179) );
  AOI21_X1 U27957 ( .A1(n1230), .A2(n7886), .B(n28379), .ZN(n26312) );
  XOR2_X1 U27958 ( .A1(n6544), .A2(n22751), .Z(n7887) );
  NAND2_X2 U27959 ( .A1(n7889), .A2(n13812), .ZN(n22751) );
  NAND2_X2 U27960 ( .A1(n7617), .A2(n7888), .ZN(n9179) );
  NAND2_X2 U27964 ( .A1(n15550), .A2(n1956), .ZN(n48315) );
  XOR2_X1 U27968 ( .A1(n15458), .A2(n7902), .Z(n39554) );
  XOR2_X1 U27969 ( .A1(n7903), .A2(n16972), .Z(n7902) );
  NAND2_X1 U27974 ( .A1(n7907), .A2(n40854), .ZN(n39782) );
  OAI21_X2 U27975 ( .A1(n40593), .A2(n7907), .B(n41073), .ZN(n41069) );
  NOR2_X1 U27976 ( .A1(n40393), .A2(n7907), .ZN(n40397) );
  XOR2_X1 U27977 ( .A1(n23719), .A2(n32572), .Z(n30958) );
  NAND2_X2 U27978 ( .A1(n7908), .A2(n30957), .ZN(n32572) );
  AOI21_X2 U27979 ( .A1(n1066), .A2(n8025), .B(n7910), .ZN(n8024) );
  NAND3_X2 U27980 ( .A1(n7911), .A2(n48493), .A3(n48492), .ZN(n7910) );
  OAI21_X1 U27981 ( .A1(n49452), .A2(n7912), .B(n22756), .ZN(n48973) );
  OR2_X1 U27982 ( .A1(n27493), .A2(n7921), .Z(n7920) );
  NOR2_X2 U27985 ( .A1(n25412), .A2(n62353), .ZN(n41567) );
  NOR2_X1 U27986 ( .A1(n41300), .A2(n42236), .ZN(n7927) );
  OAI21_X1 U27987 ( .A1(n26196), .A2(n41951), .B(n7951), .ZN(n7929) );
  NOR2_X1 U27991 ( .A1(n7931), .A2(n47797), .ZN(n10005) );
  XOR2_X1 U28000 ( .A1(n62998), .A2(n39729), .Z(n39731) );
  INV_X2 U28002 ( .I(n39781), .ZN(n40595) );
  INV_X4 U28003 ( .I(n24230), .ZN(n54197) );
  NOR2_X1 U28005 ( .A1(n23603), .A2(n24230), .ZN(n54175) );
  XOR2_X1 U28009 ( .A1(n9773), .A2(n7942), .Z(n7941) );
  XOR2_X1 U28010 ( .A1(n24053), .A2(n52405), .Z(n7942) );
  NAND2_X2 U28011 ( .A1(n29244), .A2(n27626), .ZN(n28938) );
  XOR2_X1 U28013 ( .A1(n16625), .A2(n7949), .Z(n7948) );
  NAND2_X1 U28014 ( .A1(n8139), .A2(n7950), .ZN(n43872) );
  INV_X4 U28017 ( .I(n5787), .ZN(n7950) );
  INV_X1 U28018 ( .I(n7951), .ZN(n41303) );
  CLKBUF_X4 U28019 ( .I(n26169), .Z(n7952) );
  XOR2_X1 U28022 ( .A1(n7960), .A2(n31368), .Z(n7959) );
  XOR2_X1 U28023 ( .A1(n31367), .A2(n9055), .Z(n7960) );
  NAND2_X1 U28024 ( .A1(n1437), .A2(n61007), .ZN(n7965) );
  NOR2_X2 U28027 ( .A1(n36012), .A2(n61747), .ZN(n36663) );
  OAI21_X1 U28036 ( .A1(n55006), .A2(n7973), .B(n55001), .ZN(n55002) );
  INV_X1 U28038 ( .I(n7975), .ZN(n13047) );
  OAI21_X1 U28039 ( .A1(n26592), .A2(n7975), .B(n27525), .ZN(n26593) );
  NAND2_X2 U28040 ( .A1(n9465), .A2(n23835), .ZN(n7975) );
  XOR2_X1 U28041 ( .A1(n46147), .A2(n9888), .Z(n24653) );
  INV_X1 U28042 ( .I(n7977), .ZN(n56735) );
  NAND3_X1 U28043 ( .A1(n7977), .A2(n56674), .A3(n56731), .ZN(n56651) );
  AOI22_X1 U28044 ( .A1(n56706), .A2(n17532), .B1(n7977), .B2(n56705), .ZN(
        n56713) );
  OAI22_X1 U28050 ( .A1(n29451), .A2(n29453), .B1(n22230), .B2(n7979), .ZN(
        n28727) );
  OAI21_X1 U28053 ( .A1(n55131), .A2(n7984), .B(n55136), .ZN(n7982) );
  INV_X1 U28054 ( .I(n55148), .ZN(n7989) );
  INV_X2 U28056 ( .I(n24477), .ZN(n42275) );
  XOR2_X1 U28057 ( .A1(n7997), .A2(n17777), .Z(n17776) );
  INV_X2 U28058 ( .I(n9373), .ZN(n16935) );
  XOR2_X1 U28060 ( .A1(n7999), .A2(n45400), .Z(n8000) );
  XOR2_X1 U28061 ( .A1(n4651), .A2(n1828), .Z(n8002) );
  XOR2_X1 U28066 ( .A1(n8004), .A2(n9050), .Z(n9049) );
  XOR2_X1 U28067 ( .A1(n25136), .A2(n16125), .Z(n39371) );
  XOR2_X1 U28068 ( .A1(n13548), .A2(n25721), .Z(n25136) );
  XOR2_X1 U28071 ( .A1(n24005), .A2(n18715), .Z(n51583) );
  XOR2_X1 U28072 ( .A1(n23852), .A2(n18191), .Z(n8007) );
  XOR2_X1 U28073 ( .A1(n8006), .A2(n26010), .Z(n8008) );
  NAND2_X2 U28074 ( .A1(n8010), .A2(n15743), .ZN(n37326) );
  OR2_X1 U28075 ( .A1(n37013), .A2(n8010), .Z(n23051) );
  NAND2_X2 U28077 ( .A1(n16527), .A2(n42019), .ZN(n19975) );
  NAND2_X1 U28079 ( .A1(n41928), .A2(n109), .ZN(n16072) );
  NAND2_X1 U28080 ( .A1(n43897), .A2(n43242), .ZN(n43658) );
  AND2_X1 U28082 ( .A1(n29865), .A2(n8019), .Z(n12984) );
  NOR2_X1 U28083 ( .A1(n17413), .A2(n12979), .ZN(n8020) );
  NAND3_X1 U28085 ( .A1(n48798), .A2(n22570), .A3(n1469), .ZN(n48808) );
  NOR2_X2 U28088 ( .A1(n24124), .A2(n27188), .ZN(n26660) );
  XOR2_X1 U28091 ( .A1(n8329), .A2(n32470), .Z(n32736) );
  NOR2_X1 U28093 ( .A1(n8026), .A2(n41177), .ZN(n24883) );
  NOR3_X1 U28094 ( .A1(n8026), .A2(n41173), .A3(n9393), .ZN(n14704) );
  NOR2_X1 U28096 ( .A1(n41183), .A2(n8026), .ZN(n23134) );
  OAI21_X1 U28097 ( .A1(n39145), .A2(n8026), .B(n709), .ZN(n39152) );
  NAND2_X2 U28100 ( .A1(n11245), .A2(n26332), .ZN(n14547) );
  NAND2_X1 U28103 ( .A1(n8029), .A2(n34003), .ZN(n15656) );
  NOR3_X1 U28104 ( .A1(n34165), .A2(n34658), .A3(n8029), .ZN(n34166) );
  XOR2_X1 U28106 ( .A1(n8031), .A2(n9474), .Z(n8030) );
  XOR2_X1 U28107 ( .A1(n8032), .A2(n38465), .Z(n8031) );
  XOR2_X1 U28108 ( .A1(n23853), .A2(n38464), .Z(n8032) );
  XOR2_X1 U28110 ( .A1(n38903), .A2(n39715), .Z(n8033) );
  XOR2_X1 U28111 ( .A1(n38084), .A2(n52226), .Z(n39715) );
  XOR2_X1 U28112 ( .A1(n7998), .A2(n8036), .Z(n8035) );
  XOR2_X1 U28113 ( .A1(n37807), .A2(n37661), .Z(n8036) );
  OAI22_X1 U28116 ( .A1(n35930), .A2(n8039), .B1(n21839), .B2(n1416), .ZN(
        n35931) );
  INV_X1 U28117 ( .I(n8040), .ZN(n47515) );
  INV_X1 U28121 ( .I(n8041), .ZN(n35981) );
  XNOR2_X1 U28125 ( .A1(n44098), .A2(n16519), .ZN(n8042) );
  NAND2_X2 U28131 ( .A1(n11291), .A2(n25077), .ZN(n48414) );
  XOR2_X1 U28132 ( .A1(n52115), .A2(n8179), .Z(n52116) );
  XOR2_X1 U28133 ( .A1(n2452), .A2(n17228), .Z(n17227) );
  NOR2_X1 U28137 ( .A1(n18918), .A2(n15319), .ZN(n48020) );
  AOI21_X1 U28138 ( .A1(n24393), .A2(n61089), .B(n13633), .ZN(n13632) );
  OAI21_X1 U28140 ( .A1(n10809), .A2(n77), .B(n8049), .ZN(n10808) );
  OAI21_X1 U28141 ( .A1(n12011), .A2(n12012), .B(n8049), .ZN(n12010) );
  NAND3_X2 U28144 ( .A1(n8059), .A2(n8056), .A3(n8054), .ZN(n55223) );
  XOR2_X1 U28145 ( .A1(n12299), .A2(n55516), .Z(n8065) );
  XOR2_X1 U28147 ( .A1(n15873), .A2(n8065), .Z(n8064) );
  NAND2_X1 U28151 ( .A1(n42455), .A2(n1746), .ZN(n8070) );
  AOI22_X1 U28152 ( .A1(n11374), .A2(n10805), .B1(n8072), .B2(n8296), .ZN(
        n27342) );
  INV_X2 U28154 ( .I(n8306), .ZN(n19551) );
  XOR2_X1 U28156 ( .A1(n8076), .A2(n834), .Z(n51819) );
  XOR2_X1 U28157 ( .A1(n52172), .A2(n8077), .Z(n51721) );
  XOR2_X1 U28160 ( .A1(n45045), .A2(n3208), .Z(n14061) );
  XOR2_X1 U28167 ( .A1(n51804), .A2(n50878), .Z(n8086) );
  NAND2_X2 U28168 ( .A1(n8738), .A2(n50316), .ZN(n51804) );
  NOR2_X1 U28176 ( .A1(n65233), .A2(n8097), .ZN(n30621) );
  NOR2_X2 U28177 ( .A1(n26226), .A2(n7854), .ZN(n23263) );
  INV_X2 U28178 ( .I(n16756), .ZN(n26226) );
  NAND2_X1 U28179 ( .A1(n36822), .A2(n8100), .ZN(n8101) );
  NAND4_X1 U28180 ( .A1(n36829), .A2(n17660), .A3(n24041), .A4(n37400), .ZN(
        n8100) );
  INV_X2 U28181 ( .I(n8103), .ZN(n14199) );
  NAND2_X2 U28186 ( .A1(n15693), .A2(n49384), .ZN(n49325) );
  NOR2_X2 U28187 ( .A1(n25282), .A2(n25284), .ZN(n49384) );
  XOR2_X1 U28189 ( .A1(n3523), .A2(n15735), .Z(n31983) );
  XOR2_X1 U28192 ( .A1(n14296), .A2(n33153), .Z(n8111) );
  NAND2_X1 U28194 ( .A1(n8113), .A2(n29663), .ZN(n29664) );
  NAND2_X1 U28195 ( .A1(n29375), .A2(n8113), .ZN(n29377) );
  OAI22_X1 U28196 ( .A1(n29667), .A2(n8113), .B1(n29668), .B2(n29669), .ZN(
        n29677) );
  NAND2_X1 U28198 ( .A1(n8017), .A2(n8117), .ZN(n42280) );
  XOR2_X1 U28204 ( .A1(n51012), .A2(n52028), .Z(n8125) );
  INV_X1 U28207 ( .I(n47409), .ZN(n8126) );
  NOR2_X1 U28209 ( .A1(n21881), .A2(n8132), .ZN(n36688) );
  NAND3_X2 U28212 ( .A1(n25824), .A2(n25825), .A3(n38341), .ZN(n9135) );
  AOI21_X1 U28213 ( .A1(n59476), .A2(n61134), .B(n8139), .ZN(n42747) );
  XOR2_X1 U28217 ( .A1(n26060), .A2(n8143), .Z(n8144) );
  XOR2_X1 U28218 ( .A1(n25224), .A2(n11270), .Z(n26060) );
  NAND4_X2 U28219 ( .A1(n13316), .A2(n49199), .A3(n24144), .A4(n49200), .ZN(
        n25224) );
  INV_X2 U28220 ( .I(n15041), .ZN(n19868) );
  XOR2_X1 U28224 ( .A1(n24203), .A2(n3318), .Z(n10770) );
  XOR2_X1 U28227 ( .A1(n39274), .A2(n8149), .Z(n8148) );
  NAND2_X2 U28229 ( .A1(n37917), .A2(n4275), .ZN(n43703) );
  INV_X4 U28230 ( .I(n9256), .ZN(n46982) );
  XOR2_X1 U28236 ( .A1(n11265), .A2(n31653), .Z(n8161) );
  XOR2_X1 U28237 ( .A1(n33283), .A2(n32068), .Z(n8162) );
  XOR2_X1 U28240 ( .A1(n46702), .A2(n44592), .Z(n44145) );
  XOR2_X1 U28242 ( .A1(n3523), .A2(n32192), .Z(n32194) );
  INV_X2 U28243 ( .I(n55486), .ZN(n51961) );
  NOR2_X1 U28244 ( .A1(n29586), .A2(n8167), .ZN(n8166) );
  INV_X1 U28245 ( .I(n29084), .ZN(n8167) );
  NOR2_X1 U28246 ( .A1(n29586), .A2(n8169), .ZN(n8168) );
  XOR2_X1 U28249 ( .A1(n23801), .A2(n8177), .Z(n35516) );
  INV_X2 U28250 ( .I(n8178), .ZN(n23914) );
  NOR2_X2 U28252 ( .A1(n31264), .A2(n31277), .ZN(n31268) );
  NAND2_X2 U28254 ( .A1(n20585), .A2(n20584), .ZN(n20586) );
  NAND2_X2 U28255 ( .A1(n1716), .A2(n8185), .ZN(n43335) );
  NOR2_X1 U28256 ( .A1(n1716), .A2(n8185), .ZN(n43337) );
  NAND2_X1 U28257 ( .A1(n14620), .A2(n20586), .ZN(n41627) );
  XOR2_X1 U28260 ( .A1(n26920), .A2(n8186), .Z(n31561) );
  XOR2_X1 U28261 ( .A1(n30949), .A2(n8186), .Z(n30950) );
  XOR2_X1 U28262 ( .A1(n8186), .A2(n17463), .Z(n32673) );
  XOR2_X1 U28265 ( .A1(n8196), .A2(n39553), .Z(n11091) );
  NOR2_X1 U28267 ( .A1(n1742), .A2(n1407), .ZN(n25180) );
  NAND2_X1 U28268 ( .A1(n40832), .A2(n64450), .ZN(n15084) );
  XOR2_X1 U28272 ( .A1(n32634), .A2(n8197), .Z(n32635) );
  XOR2_X1 U28273 ( .A1(n33031), .A2(n32633), .Z(n8197) );
  NAND3_X2 U28276 ( .A1(n18327), .A2(n37665), .A3(n1004), .ZN(n18482) );
  OAI21_X1 U28280 ( .A1(n55699), .A2(n55698), .B(n8203), .ZN(n55700) );
  XOR2_X1 U28283 ( .A1(n23464), .A2(n37650), .Z(n39270) );
  XOR2_X1 U28285 ( .A1(n37554), .A2(n39646), .Z(n37657) );
  XOR2_X1 U28288 ( .A1(n8209), .A2(n38861), .Z(n8208) );
  NOR3_X1 U28290 ( .A1(n20378), .A2(n8211), .A3(n31208), .ZN(n11968) );
  XOR2_X1 U28293 ( .A1(n11252), .A2(n44223), .Z(n14783) );
  AOI21_X1 U28295 ( .A1(n8619), .A2(n43341), .B(n25368), .ZN(n42163) );
  INV_X2 U28299 ( .I(n8219), .ZN(n9628) );
  XOR2_X1 U28300 ( .A1(n12377), .A2(n9628), .Z(n19947) );
  INV_X2 U28302 ( .I(n11090), .ZN(n20552) );
  OAI21_X1 U28303 ( .A1(n41924), .A2(n287), .B(n59531), .ZN(n40560) );
  XOR2_X1 U28305 ( .A1(n31759), .A2(n32640), .Z(n8221) );
  OAI21_X1 U28309 ( .A1(n17660), .A2(n8223), .B(n37404), .ZN(n37406) );
  NAND3_X1 U28310 ( .A1(n36828), .A2(n8195), .A3(n8223), .ZN(n36832) );
  XOR2_X1 U28312 ( .A1(n11167), .A2(n8226), .Z(n50968) );
  XOR2_X1 U28314 ( .A1(n8229), .A2(n23422), .Z(n21133) );
  NAND3_X1 U28316 ( .A1(n14891), .A2(n38993), .A3(n14894), .ZN(n8231) );
  INV_X1 U28317 ( .I(n8233), .ZN(n8232) );
  XOR2_X1 U28319 ( .A1(n3798), .A2(n33140), .Z(n8236) );
  NAND2_X1 U28323 ( .A1(n36513), .A2(n36524), .ZN(n8241) );
  XOR2_X1 U28326 ( .A1(n10291), .A2(n1902), .Z(n24248) );
  NAND2_X2 U28327 ( .A1(n41445), .A2(n39847), .ZN(n41442) );
  NAND2_X2 U28328 ( .A1(n42939), .A2(n43444), .ZN(n42947) );
  NOR2_X2 U28329 ( .A1(n8247), .A2(n43437), .ZN(n42939) );
  INV_X2 U28331 ( .I(n8249), .ZN(n13639) );
  OAI21_X2 U28332 ( .A1(n52176), .A2(n7331), .B(n8250), .ZN(n13622) );
  NOR2_X2 U28335 ( .A1(n1926), .A2(n8478), .ZN(n8437) );
  NAND2_X1 U28337 ( .A1(n14549), .A2(n55651), .ZN(n8256) );
  NOR2_X1 U28338 ( .A1(n26183), .A2(n8258), .ZN(n8257) );
  INV_X1 U28343 ( .I(n8261), .ZN(n9238) );
  XOR2_X1 U28344 ( .A1(n32029), .A2(n8263), .Z(n8262) );
  XOR2_X1 U28345 ( .A1(n1313), .A2(n32710), .Z(n32029) );
  NAND2_X2 U28349 ( .A1(n8275), .A2(n8274), .ZN(n19540) );
  XOR2_X1 U28351 ( .A1(n8277), .A2(n19540), .Z(n13687) );
  XOR2_X1 U28352 ( .A1(n52472), .A2(n8278), .Z(n8277) );
  XOR2_X1 U28353 ( .A1(n63001), .A2(n8279), .Z(n8278) );
  INV_X1 U28357 ( .I(n14752), .ZN(n25612) );
  XOR2_X1 U28358 ( .A1(n17869), .A2(n8281), .Z(n8280) );
  XOR2_X1 U28359 ( .A1(n14760), .A2(n8282), .Z(n8281) );
  XOR2_X1 U28360 ( .A1(n23548), .A2(n45062), .Z(n8282) );
  XOR2_X1 U28364 ( .A1(n14857), .A2(n55087), .Z(n45058) );
  XOR2_X1 U28365 ( .A1(n12879), .A2(n870), .Z(n39560) );
  XOR2_X1 U28366 ( .A1(n12879), .A2(n1900), .Z(n39640) );
  NOR2_X2 U28367 ( .A1(n23743), .A2(n34708), .ZN(n35307) );
  XOR2_X1 U28370 ( .A1(n1329), .A2(n43484), .Z(n45249) );
  XOR2_X1 U28371 ( .A1(n31836), .A2(n18541), .Z(n8288) );
  XOR2_X1 U28372 ( .A1(n9373), .A2(n18543), .Z(n31836) );
  INV_X2 U28373 ( .I(n8289), .ZN(n15091) );
  NAND2_X2 U28374 ( .A1(n40823), .A2(n40824), .ZN(n8289) );
  INV_X2 U28376 ( .I(n19806), .ZN(n22332) );
  XOR2_X1 U28377 ( .A1(n12697), .A2(n52531), .Z(n9773) );
  XOR2_X1 U28378 ( .A1(n19806), .A2(n25158), .Z(n52531) );
  NAND2_X2 U28379 ( .A1(n8292), .A2(n11217), .ZN(n25158) );
  NOR3_X1 U28381 ( .A1(n37236), .A2(n36883), .A3(n37444), .ZN(n8295) );
  NOR2_X1 U28382 ( .A1(n8298), .A2(n63954), .ZN(n49831) );
  NOR2_X1 U28383 ( .A1(n20458), .A2(n8298), .ZN(n49836) );
  OAI21_X1 U28385 ( .A1(n65135), .A2(n8298), .B(n11705), .ZN(n45701) );
  AOI21_X1 U28386 ( .A1(n65135), .A2(n8298), .B(n11950), .ZN(n45702) );
  NAND2_X1 U28387 ( .A1(n20458), .A2(n8298), .ZN(n49827) );
  OAI22_X1 U28389 ( .A1(n49079), .A2(n62861), .B1(n49078), .B2(n49077), .ZN(
        n49080) );
  XOR2_X1 U28392 ( .A1(n7573), .A2(n37577), .Z(n8301) );
  NAND3_X1 U28394 ( .A1(n12975), .A2(n8303), .A3(n22776), .ZN(n41930) );
  NAND2_X1 U28395 ( .A1(n16870), .A2(n8303), .ZN(n40817) );
  NAND2_X1 U28396 ( .A1(n34666), .A2(n8304), .ZN(n12339) );
  NOR2_X1 U28397 ( .A1(n21906), .A2(n8304), .ZN(n33450) );
  NAND2_X2 U28400 ( .A1(n5787), .A2(n11609), .ZN(n43350) );
  XOR2_X1 U28402 ( .A1(n19551), .A2(n16706), .Z(n31432) );
  NOR2_X2 U28404 ( .A1(n47314), .A2(n15824), .ZN(n47328) );
  NAND2_X2 U28405 ( .A1(n8902), .A2(n25502), .ZN(n8905) );
  NAND2_X2 U28407 ( .A1(n15311), .A2(n15313), .ZN(n55387) );
  NAND3_X2 U28416 ( .A1(n8328), .A2(n8327), .A3(n8326), .ZN(n55135) );
  XOR2_X1 U28418 ( .A1(n8333), .A2(n8330), .Z(n8594) );
  XOR2_X1 U28419 ( .A1(n8331), .A2(n8332), .Z(n8330) );
  XOR2_X1 U28420 ( .A1(n9283), .A2(n32560), .Z(n8331) );
  XOR2_X1 U28421 ( .A1(n1825), .A2(n8329), .Z(n8332) );
  NOR2_X2 U28424 ( .A1(n23216), .A2(n29271), .ZN(n19654) );
  INV_X2 U28427 ( .I(n8341), .ZN(n41386) );
  INV_X4 U28428 ( .I(n41386), .ZN(n41122) );
  XOR2_X1 U28429 ( .A1(n39677), .A2(n39676), .Z(n8341) );
  NOR2_X1 U28431 ( .A1(n22657), .A2(n59381), .ZN(n42994) );
  INV_X2 U28436 ( .I(n49564), .ZN(n48832) );
  NAND2_X2 U28437 ( .A1(n58907), .A2(n8347), .ZN(n49564) );
  NAND2_X1 U28440 ( .A1(n61107), .A2(n15784), .ZN(n8352) );
  AOI21_X2 U28444 ( .A1(n34565), .A2(n32971), .B(n32970), .ZN(n36377) );
  INV_X2 U28446 ( .I(n8359), .ZN(n27622) );
  NOR2_X2 U28447 ( .A1(n15758), .A2(n19522), .ZN(n8359) );
  NAND2_X1 U28451 ( .A1(n8367), .A2(n51268), .ZN(n18270) );
  NAND3_X1 U28454 ( .A1(n56398), .A2(n8367), .A3(n62769), .ZN(n56399) );
  NOR2_X2 U28455 ( .A1(n55936), .A2(n12605), .ZN(n8367) );
  AOI21_X1 U28457 ( .A1(n23568), .A2(n27998), .B(n27997), .ZN(n8372) );
  OAI21_X1 U28458 ( .A1(n8373), .A2(n43270), .B(n43268), .ZN(n8785) );
  NOR2_X1 U28459 ( .A1(n23541), .A2(n8373), .ZN(n41792) );
  NAND2_X1 U28460 ( .A1(n43131), .A2(n8373), .ZN(n25439) );
  INV_X1 U28462 ( .I(n54471), .ZN(n54322) );
  NAND2_X2 U28468 ( .A1(n13614), .A2(n1209), .ZN(n50267) );
  NOR2_X1 U28469 ( .A1(n8378), .A2(n30455), .ZN(n29061) );
  NAND3_X1 U28470 ( .A1(n18402), .A2(n8378), .A3(n30455), .ZN(n29060) );
  NAND2_X1 U28471 ( .A1(n60170), .A2(n8378), .ZN(n29431) );
  NAND2_X1 U28477 ( .A1(n48943), .A2(n8380), .ZN(n13923) );
  XOR2_X1 U28483 ( .A1(n17657), .A2(n8387), .Z(n8386) );
  XOR2_X1 U28485 ( .A1(n37579), .A2(n11751), .Z(n37634) );
  NAND2_X2 U28488 ( .A1(n23822), .A2(n10403), .ZN(n8389) );
  INV_X1 U28491 ( .I(n30832), .ZN(n23400) );
  NAND2_X1 U28493 ( .A1(n8405), .A2(n64458), .ZN(n8689) );
  NAND2_X1 U28494 ( .A1(n8405), .A2(n26242), .ZN(n34241) );
  XOR2_X1 U28498 ( .A1(n10531), .A2(n2952), .Z(n31964) );
  XOR2_X1 U28500 ( .A1(n12034), .A2(n42019), .Z(n8415) );
  NOR2_X1 U28508 ( .A1(n23170), .A2(n27996), .ZN(n8420) );
  XOR2_X1 U28510 ( .A1(n31762), .A2(n8423), .Z(n8422) );
  NAND2_X2 U28511 ( .A1(n14151), .A2(n14148), .ZN(n18306) );
  NOR2_X1 U28512 ( .A1(n8424), .A2(n30319), .ZN(n28697) );
  INV_X2 U28515 ( .I(n8427), .ZN(n38021) );
  NOR2_X2 U28517 ( .A1(n42080), .A2(n25071), .ZN(n42395) );
  NAND2_X1 U28519 ( .A1(n8431), .A2(n34530), .ZN(n33722) );
  INV_X1 U28523 ( .I(n28216), .ZN(n27968) );
  XOR2_X1 U28524 ( .A1(Ciphertext[73]), .A2(Key[20]), .Z(n15043) );
  NAND3_X2 U28526 ( .A1(n12633), .A2(n13023), .A3(n19474), .ZN(n19473) );
  NOR2_X2 U28527 ( .A1(n16852), .A2(n57536), .ZN(n40106) );
  NAND2_X2 U28528 ( .A1(n20046), .A2(n40100), .ZN(n20047) );
  INV_X2 U28529 ( .I(n8443), .ZN(n10205) );
  XOR2_X1 U28533 ( .A1(n8449), .A2(n16315), .Z(n8450) );
  NOR2_X1 U28534 ( .A1(n63311), .A2(n19040), .ZN(n48657) );
  NOR2_X2 U28537 ( .A1(n34149), .A2(n32846), .ZN(n34156) );
  NAND2_X2 U28539 ( .A1(n19773), .A2(n20199), .ZN(n50046) );
  NAND2_X2 U28543 ( .A1(n15546), .A2(n28947), .ZN(n12898) );
  XOR2_X1 U28551 ( .A1(n8472), .A2(n10101), .Z(n51653) );
  XOR2_X1 U28552 ( .A1(n8472), .A2(n51756), .Z(n51759) );
  NOR2_X2 U28553 ( .A1(n49917), .A2(n49916), .ZN(n8473) );
  NAND2_X2 U28554 ( .A1(n57701), .A2(n61646), .ZN(n18884) );
  NAND2_X1 U28555 ( .A1(n10254), .A2(n8474), .ZN(n36039) );
  NOR2_X1 U28556 ( .A1(n8474), .A2(n10254), .ZN(n35580) );
  NAND2_X1 U28559 ( .A1(n32857), .A2(n8474), .ZN(n17191) );
  NOR2_X1 U28560 ( .A1(n8475), .A2(n10225), .ZN(n45179) );
  NAND3_X1 U28561 ( .A1(n8924), .A2(n47882), .A3(n8475), .ZN(n8923) );
  XOR2_X1 U28562 ( .A1(n20270), .A2(n14737), .Z(n12381) );
  XOR2_X1 U28563 ( .A1(n19540), .A2(n8477), .Z(n8848) );
  INV_X2 U28566 ( .I(n15043), .ZN(n8478) );
  INV_X4 U28567 ( .I(n15101), .ZN(n40943) );
  XOR2_X1 U28571 ( .A1(n8480), .A2(n43334), .Z(n23566) );
  XOR2_X1 U28572 ( .A1(n13883), .A2(n8480), .Z(n45108) );
  OR2_X1 U28573 ( .A1(n38498), .A2(n9189), .Z(n8483) );
  NAND2_X2 U28574 ( .A1(n18240), .A2(n38023), .ZN(n38498) );
  NAND2_X2 U28576 ( .A1(n38495), .A2(n41034), .ZN(n9189) );
  NAND2_X2 U28577 ( .A1(n24455), .A2(n55668), .ZN(n55293) );
  XOR2_X1 U28579 ( .A1(n30935), .A2(n8492), .Z(n30936) );
  NAND2_X1 U28584 ( .A1(n19629), .A2(n19632), .ZN(n8496) );
  NOR2_X2 U28586 ( .A1(n15152), .A2(n24664), .ZN(n34661) );
  XOR2_X1 U28587 ( .A1(n8499), .A2(n929), .Z(n8498) );
  XOR2_X1 U28588 ( .A1(n8500), .A2(n35912), .Z(n8499) );
  XOR2_X1 U28592 ( .A1(n31708), .A2(n8505), .Z(n10197) );
  XOR2_X1 U28593 ( .A1(n32493), .A2(n32084), .Z(n8505) );
  NAND3_X2 U28594 ( .A1(n48499), .A2(n3091), .A3(n48514), .ZN(n48639) );
  INV_X2 U28596 ( .I(n28059), .ZN(n24896) );
  NAND2_X1 U28597 ( .A1(n28059), .A2(n22556), .ZN(n29821) );
  NAND2_X2 U28598 ( .A1(n8511), .A2(n9775), .ZN(n28059) );
  NAND2_X2 U28599 ( .A1(n55287), .A2(n55470), .ZN(n8513) );
  INV_X2 U28600 ( .I(n8514), .ZN(n35738) );
  OAI21_X1 U28605 ( .A1(n26597), .A2(n26598), .B(n8518), .ZN(n26601) );
  NAND2_X2 U28606 ( .A1(n11767), .A2(n14439), .ZN(n8518) );
  OAI21_X1 U28610 ( .A1(n61187), .A2(n10830), .B(n30812), .ZN(n10573) );
  AOI21_X1 U28616 ( .A1(n30333), .A2(n11092), .B(n8522), .ZN(n27991) );
  NAND2_X1 U28617 ( .A1(n30409), .A2(n8522), .ZN(n30411) );
  NAND3_X1 U28619 ( .A1(n29945), .A2(n29944), .A3(n8522), .ZN(n29946) );
  NOR2_X1 U28621 ( .A1(n5980), .A2(n8523), .ZN(n8841) );
  XOR2_X1 U28622 ( .A1(n9787), .A2(n45878), .Z(n8527) );
  NOR2_X1 U28624 ( .A1(n27262), .A2(n8528), .ZN(n27973) );
  NOR2_X1 U28626 ( .A1(n1886), .A2(n4457), .ZN(n18536) );
  XOR2_X1 U28627 ( .A1(n22361), .A2(n16401), .Z(n8529) );
  NAND2_X2 U28628 ( .A1(n24273), .A2(n19512), .ZN(n34610) );
  NAND2_X1 U28629 ( .A1(n856), .A2(n29297), .ZN(n29298) );
  NAND2_X1 U28630 ( .A1(n57830), .A2(n36259), .ZN(n8535) );
  NAND2_X2 U28631 ( .A1(n39035), .A2(n8538), .ZN(n8537) );
  XOR2_X1 U28636 ( .A1(n8543), .A2(n8542), .Z(n8541) );
  INV_X2 U28641 ( .I(n8551), .ZN(n8805) );
  XNOR2_X1 U28642 ( .A1(n52443), .A2(n50582), .ZN(n8550) );
  NAND4_X2 U28643 ( .A1(n47350), .A2(n19848), .A3(n47349), .A4(n47348), .ZN(
        n52443) );
  NOR2_X2 U28644 ( .A1(n19850), .A2(n49444), .ZN(n50582) );
  XOR2_X1 U28653 ( .A1(n8561), .A2(n8560), .Z(n8559) );
  XOR2_X1 U28654 ( .A1(n15729), .A2(n16404), .Z(n8560) );
  XOR2_X1 U28655 ( .A1(n39221), .A2(n17583), .Z(n8561) );
  XOR2_X1 U28656 ( .A1(n4470), .A2(n1576), .Z(n8562) );
  XOR2_X1 U28659 ( .A1(n7253), .A2(n8564), .Z(n8563) );
  NAND2_X1 U28660 ( .A1(n892), .A2(n13487), .ZN(n34405) );
  INV_X4 U28661 ( .I(n25068), .ZN(n42080) );
  INV_X2 U28664 ( .I(n8567), .ZN(n8590) );
  XOR2_X1 U28665 ( .A1(n8590), .A2(n29557), .Z(n14808) );
  XOR2_X1 U28667 ( .A1(n17497), .A2(n65280), .Z(n8843) );
  XOR2_X1 U28668 ( .A1(n52177), .A2(n8569), .Z(n25542) );
  XOR2_X1 U28669 ( .A1(n48946), .A2(n23371), .Z(n8570) );
  XOR2_X1 U28670 ( .A1(n44991), .A2(n7424), .Z(n44528) );
  XOR2_X1 U28671 ( .A1(n23067), .A2(n7424), .Z(n43967) );
  XOR2_X1 U28672 ( .A1(n44223), .A2(n7424), .Z(n44190) );
  XOR2_X1 U28673 ( .A1(n4953), .A2(n16307), .Z(n8575) );
  INV_X1 U28674 ( .I(n42160), .ZN(n42161) );
  INV_X4 U28676 ( .I(n31141), .ZN(n30585) );
  NAND2_X2 U28677 ( .A1(n8586), .A2(n1836), .ZN(n24746) );
  XOR2_X1 U28678 ( .A1(n8587), .A2(n1135), .Z(n26070) );
  XOR2_X1 U28679 ( .A1(n8588), .A2(n810), .Z(n8587) );
  NOR2_X1 U28683 ( .A1(n43845), .A2(n8589), .ZN(n43072) );
  NAND2_X1 U28684 ( .A1(n24002), .A2(n22112), .ZN(n43841) );
  NAND2_X2 U28685 ( .A1(n39918), .A2(n10972), .ZN(n8589) );
  XOR2_X1 U28686 ( .A1(n8593), .A2(n8591), .Z(n9118) );
  XOR2_X1 U28688 ( .A1(n8590), .A2(n31654), .Z(n33051) );
  NAND2_X2 U28692 ( .A1(n13757), .A2(n15536), .ZN(n8597) );
  INV_X2 U28694 ( .I(n8600), .ZN(n23464) );
  XOR2_X1 U28696 ( .A1(n23464), .A2(n8601), .Z(n37727) );
  NOR2_X2 U28698 ( .A1(n40578), .A2(n42259), .ZN(n42266) );
  NAND2_X1 U28701 ( .A1(n30252), .A2(n10205), .ZN(n30262) );
  XOR2_X1 U28703 ( .A1(n9011), .A2(n17233), .Z(n18308) );
  NOR2_X2 U28704 ( .A1(n1292), .A2(n24332), .ZN(n17523) );
  XOR2_X1 U28712 ( .A1(n43941), .A2(n1576), .Z(n44130) );
  NOR2_X2 U28713 ( .A1(n20851), .A2(n8612), .ZN(n43941) );
  XOR2_X1 U28720 ( .A1(n46189), .A2(n8620), .Z(n46190) );
  XOR2_X1 U28723 ( .A1(n31816), .A2(n8624), .Z(n8623) );
  XOR2_X1 U28724 ( .A1(n23768), .A2(n31821), .Z(n8624) );
  CLKBUF_X4 U28725 ( .I(n6544), .Z(n8625) );
  XOR2_X1 U28726 ( .A1(n20719), .A2(n8625), .Z(n31768) );
  INV_X2 U28727 ( .I(n5604), .ZN(n34385) );
  XOR2_X1 U28732 ( .A1(n37158), .A2(n38004), .Z(n25211) );
  NOR2_X1 U28737 ( .A1(n17747), .A2(n27298), .ZN(n27299) );
  NOR2_X1 U28738 ( .A1(n27301), .A2(n17747), .ZN(n22679) );
  NAND2_X2 U28740 ( .A1(n8772), .A2(n23140), .ZN(n8770) );
  XOR2_X1 U28742 ( .A1(n19993), .A2(n15726), .Z(n31795) );
  XOR2_X1 U28743 ( .A1(n15413), .A2(n8652), .Z(n15412) );
  NOR2_X2 U28749 ( .A1(n8659), .A2(n8658), .ZN(n14955) );
  NOR2_X2 U28751 ( .A1(n40683), .A2(n8662), .ZN(n12567) );
  NAND2_X2 U28752 ( .A1(n10968), .A2(n54112), .ZN(n10938) );
  INV_X1 U28756 ( .I(n20923), .ZN(n33357) );
  NOR2_X2 U28758 ( .A1(n34155), .A2(n61196), .ZN(n20923) );
  MUX2_X1 U28759 ( .I0(n47018), .I1(n1651), .S(n8666), .Z(n12231) );
  AND2_X1 U28765 ( .A1(n8672), .A2(n27512), .Z(n8671) );
  AND2_X1 U28766 ( .A1(n27511), .A2(n29358), .Z(n8672) );
  XOR2_X1 U28767 ( .A1(n18311), .A2(n25836), .Z(n18310) );
  XOR2_X1 U28768 ( .A1(n44120), .A2(n62065), .Z(n25836) );
  XOR2_X1 U28770 ( .A1(n45094), .A2(n8673), .Z(n45095) );
  XOR2_X1 U28771 ( .A1(n31982), .A2(n32028), .Z(n21105) );
  XOR2_X1 U28774 ( .A1(n52373), .A2(n56202), .Z(n8674) );
  XOR2_X1 U28776 ( .A1(n4659), .A2(n11476), .Z(n39876) );
  NAND3_X1 U28779 ( .A1(n48956), .A2(n10873), .A3(n8679), .ZN(n12674) );
  XOR2_X1 U28780 ( .A1(n13579), .A2(n3665), .Z(n11911) );
  XOR2_X1 U28781 ( .A1(n37677), .A2(n8684), .Z(n13579) );
  NAND2_X2 U28783 ( .A1(n43130), .A2(n1701), .ZN(n8687) );
  XOR2_X1 U28784 ( .A1(n46133), .A2(n46137), .Z(n8795) );
  INV_X2 U28786 ( .I(n41112), .ZN(n23046) );
  INV_X2 U28787 ( .I(n19761), .ZN(n24071) );
  INV_X1 U28788 ( .I(n47659), .ZN(n47561) );
  INV_X2 U28799 ( .I(n8716), .ZN(n10502) );
  AOI22_X2 U28800 ( .A1(n42646), .A2(n4467), .B1(n43534), .B2(n43538), .ZN(
        n43780) );
  XOR2_X1 U28801 ( .A1(n3717), .A2(n65046), .Z(n8720) );
  NOR2_X2 U28802 ( .A1(n8722), .A2(n25987), .ZN(n56955) );
  OAI22_X1 U28803 ( .A1(n56926), .A2(n8722), .B1(n56925), .B2(n56924), .ZN(
        n56931) );
  NOR2_X1 U28807 ( .A1(n8734), .A2(n56008), .ZN(n21711) );
  NAND3_X1 U28808 ( .A1(n8734), .A2(n21293), .A3(n56008), .ZN(n21708) );
  INV_X2 U28811 ( .I(n33005), .ZN(n32461) );
  XOR2_X1 U28812 ( .A1(n46625), .A2(n62065), .Z(n46714) );
  XOR2_X1 U28813 ( .A1(n8735), .A2(n9874), .Z(n25956) );
  XOR2_X1 U28814 ( .A1(n8736), .A2(n25958), .Z(n8735) );
  XOR2_X1 U28818 ( .A1(n11261), .A2(n22265), .Z(n23669) );
  NAND3_X2 U28822 ( .A1(n48541), .A2(n8750), .A3(n8748), .ZN(n23194) );
  NAND2_X2 U28825 ( .A1(n8754), .A2(n18366), .ZN(n37067) );
  XOR2_X1 U28826 ( .A1(n15406), .A2(n39192), .Z(n8766) );
  XOR2_X1 U28827 ( .A1(n63133), .A2(n15615), .Z(n39192) );
  INV_X2 U28828 ( .I(n8767), .ZN(n43218) );
  XOR2_X1 U28829 ( .A1(n43218), .A2(n797), .Z(n44334) );
  XOR2_X1 U28830 ( .A1(n21142), .A2(n8769), .Z(n21143) );
  INV_X1 U28831 ( .I(n43218), .ZN(n8769) );
  INV_X4 U28832 ( .I(n30649), .ZN(n23140) );
  INV_X1 U28833 ( .I(n27988), .ZN(n8772) );
  INV_X2 U28834 ( .I(n27988), .ZN(n30333) );
  OAI22_X1 U28842 ( .A1(n36054), .A2(n18144), .B1(n36385), .B2(n8781), .ZN(
        n33125) );
  OAI21_X1 U28843 ( .A1(n24078), .A2(n65075), .B(n8781), .ZN(n33111) );
  AOI21_X1 U28844 ( .A1(n24078), .A2(n8781), .B(n33124), .ZN(n33126) );
  XOR2_X1 U28850 ( .A1(n16901), .A2(n8796), .Z(n16900) );
  NAND2_X1 U28858 ( .A1(n65276), .A2(n48779), .ZN(n47913) );
  INV_X4 U28860 ( .I(n8803), .ZN(n29452) );
  NOR2_X1 U28862 ( .A1(n29453), .A2(n22230), .ZN(n29848) );
  INV_X4 U28863 ( .I(n29452), .ZN(n22230) );
  NAND2_X2 U28864 ( .A1(n9469), .A2(n9466), .ZN(n8803) );
  NOR2_X1 U28865 ( .A1(n22591), .A2(n8806), .ZN(n20828) );
  NAND2_X2 U28866 ( .A1(n23636), .A2(n26641), .ZN(n27179) );
  INV_X1 U28870 ( .I(n37677), .ZN(n19060) );
  XOR2_X1 U28871 ( .A1(n37677), .A2(n35956), .Z(n35957) );
  NAND2_X1 U28876 ( .A1(n41945), .A2(n8812), .ZN(n16775) );
  AOI21_X1 U28877 ( .A1(n12735), .A2(n8812), .B(n61435), .ZN(n12734) );
  XOR2_X1 U28878 ( .A1(n9570), .A2(n31981), .Z(n21740) );
  XOR2_X1 U28881 ( .A1(n8825), .A2(n56702), .Z(Plaintext[165]) );
  NOR2_X2 U28882 ( .A1(n21893), .A2(n56624), .ZN(n56619) );
  NAND2_X1 U28883 ( .A1(n56621), .A2(n56622), .ZN(n8829) );
  MUX2_X1 U28884 ( .I0(n28505), .I1(n28506), .S(n27853), .Z(n28513) );
  NAND3_X2 U28885 ( .A1(n21056), .A2(n34752), .A3(n34753), .ZN(n21863) );
  NOR2_X2 U28886 ( .A1(n17958), .A2(n8832), .ZN(n34753) );
  INV_X1 U28887 ( .I(n34342), .ZN(n8832) );
  XOR2_X1 U28888 ( .A1(n13294), .A2(n50623), .Z(n51056) );
  XOR2_X1 U28889 ( .A1(n24929), .A2(n185), .Z(n50623) );
  XOR2_X1 U28890 ( .A1(n8837), .A2(n8835), .Z(n34336) );
  XOR2_X1 U28891 ( .A1(n63029), .A2(n32038), .Z(n8835) );
  XOR2_X1 U28892 ( .A1(n8836), .A2(n9712), .Z(n32038) );
  XOR2_X1 U28893 ( .A1(n31336), .A2(n1314), .Z(n8836) );
  XOR2_X1 U28896 ( .A1(n31998), .A2(n31999), .Z(n8839) );
  NAND2_X1 U28897 ( .A1(n48665), .A2(n8842), .ZN(n20404) );
  NAND2_X1 U28898 ( .A1(n48667), .A2(n8842), .ZN(n20679) );
  AOI21_X1 U28899 ( .A1(n15757), .A2(n16628), .B(n8842), .ZN(n48672) );
  XOR2_X1 U28901 ( .A1(n8844), .A2(n8843), .Z(n22092) );
  XOR2_X1 U28903 ( .A1(n51986), .A2(n51069), .Z(n8847) );
  XOR2_X1 U28904 ( .A1(n8848), .A2(n12599), .Z(n51226) );
  NOR2_X1 U28906 ( .A1(n52786), .A2(n57046), .ZN(n8850) );
  INV_X2 U28908 ( .I(n57046), .ZN(n8851) );
  NAND2_X1 U28909 ( .A1(n8852), .A2(n15283), .ZN(n40276) );
  NOR2_X1 U28910 ( .A1(n8852), .A2(n12402), .ZN(n24569) );
  INV_X2 U28914 ( .I(n8854), .ZN(n13232) );
  AOI22_X1 U28916 ( .A1(n8860), .A2(n59924), .B1(n10765), .B2(n36871), .ZN(
        n8859) );
  OR2_X1 U28917 ( .A1(n36870), .A2(n25396), .Z(n8860) );
  XOR2_X1 U28918 ( .A1(n46668), .A2(n46186), .Z(n8864) );
  XOR2_X1 U28920 ( .A1(n46185), .A2(n3449), .Z(n8865) );
  XOR2_X1 U28922 ( .A1(n44354), .A2(n19071), .Z(n44338) );
  XOR2_X1 U28923 ( .A1(n44549), .A2(n8869), .Z(n8868) );
  NOR2_X1 U28927 ( .A1(n8877), .A2(n8876), .ZN(n8875) );
  NAND2_X1 U28928 ( .A1(n42588), .A2(n42589), .ZN(n8877) );
  XOR2_X1 U28932 ( .A1(n25111), .A2(n51019), .Z(n33261) );
  XOR2_X1 U28933 ( .A1(n18391), .A2(n10409), .Z(n8885) );
  NOR2_X1 U28934 ( .A1(n8887), .A2(n10030), .ZN(n45236) );
  OR2_X1 U28935 ( .A1(n8887), .A2(n49150), .Z(n49151) );
  INV_X2 U28936 ( .I(n17496), .ZN(n13943) );
  NAND2_X2 U28937 ( .A1(n8893), .A2(n19829), .ZN(n17496) );
  NOR2_X2 U28938 ( .A1(n18882), .A2(n60163), .ZN(n49811) );
  NAND2_X2 U28939 ( .A1(n60360), .A2(n5258), .ZN(n50437) );
  XOR2_X1 U28940 ( .A1(n43218), .A2(n46233), .Z(n8900) );
  NAND2_X1 U28944 ( .A1(n55910), .A2(n15454), .ZN(n17601) );
  NAND2_X2 U28945 ( .A1(n1326), .A2(n55909), .ZN(n55910) );
  NAND2_X2 U28949 ( .A1(n9229), .A2(n59633), .ZN(n16543) );
  XOR2_X1 U28956 ( .A1(n46243), .A2(n46235), .Z(n8929) );
  XOR2_X1 U28957 ( .A1(n44965), .A2(n45402), .Z(n46235) );
  XOR2_X1 U28958 ( .A1(n25872), .A2(n46137), .Z(n46243) );
  XOR2_X1 U28961 ( .A1(n25531), .A2(n57892), .Z(n44965) );
  XOR2_X1 U28962 ( .A1(n46237), .A2(n46236), .Z(n8932) );
  OAI21_X1 U28965 ( .A1(n1837), .A2(n19461), .B(n30230), .ZN(n8947) );
  XOR2_X1 U28966 ( .A1(n8951), .A2(n33838), .Z(n8950) );
  XOR2_X1 U28967 ( .A1(n25203), .A2(n33158), .Z(n8951) );
  XOR2_X1 U28968 ( .A1(n13365), .A2(n13449), .Z(n8952) );
  INV_X2 U28969 ( .I(n13026), .ZN(n55722) );
  XOR2_X1 U28971 ( .A1(n51737), .A2(n8955), .Z(n8954) );
  OAI21_X1 U28974 ( .A1(n35834), .A2(n35709), .B(n8956), .ZN(n35711) );
  NAND3_X1 U28975 ( .A1(n35834), .A2(n33807), .A3(n34404), .ZN(n8956) );
  OAI22_X1 U28976 ( .A1(n2168), .A2(n34395), .B1(n21252), .B2(n8957), .ZN(
        n33210) );
  NAND2_X2 U28977 ( .A1(n27921), .A2(n62231), .ZN(n16504) );
  XOR2_X1 U28983 ( .A1(n16691), .A2(n24758), .Z(n51125) );
  XOR2_X1 U28984 ( .A1(n49809), .A2(n8975), .Z(n8974) );
  INV_X2 U28990 ( .I(n8982), .ZN(n27921) );
  XOR2_X1 U28991 ( .A1(n8984), .A2(n65210), .Z(n36647) );
  AOI21_X1 U28993 ( .A1(n56130), .A2(n56174), .B(n8985), .ZN(n56131) );
  NAND3_X1 U28994 ( .A1(n19853), .A2(n56169), .A3(n8985), .ZN(n56140) );
  NAND2_X2 U28997 ( .A1(n43741), .A2(n8986), .ZN(n13630) );
  XOR2_X1 U29003 ( .A1(n46270), .A2(n1019), .Z(n9005) );
  NAND2_X1 U29004 ( .A1(n21008), .A2(n9012), .ZN(n33719) );
  NAND2_X2 U29006 ( .A1(n21237), .A2(n26354), .ZN(n29801) );
  NAND2_X1 U29008 ( .A1(n825), .A2(n40949), .ZN(n9015) );
  INV_X1 U29010 ( .I(Key[162]), .ZN(n9018) );
  INV_X2 U29012 ( .I(n27524), .ZN(n27526) );
  INV_X2 U29014 ( .I(n9019), .ZN(n12880) );
  NAND3_X2 U29015 ( .A1(n37284), .A2(n37282), .A3(n37283), .ZN(n38063) );
  XNOR2_X1 U29016 ( .A1(n23464), .A2(n12880), .ZN(n17710) );
  XOR2_X1 U29017 ( .A1(n718), .A2(n26010), .Z(n11486) );
  OAI21_X1 U29018 ( .A1(n18597), .A2(n9022), .B(n56434), .ZN(n9056) );
  NAND2_X2 U29021 ( .A1(n64712), .A2(n23836), .ZN(n56997) );
  AOI21_X1 U29023 ( .A1(n53234), .A2(n64712), .B(n62515), .ZN(n53235) );
  XOR2_X1 U29024 ( .A1(n20228), .A2(n11665), .Z(n9024) );
  NAND2_X2 U29025 ( .A1(n18919), .A2(n16864), .ZN(n42646) );
  NOR2_X2 U29026 ( .A1(n35920), .A2(n9026), .ZN(n37411) );
  INV_X1 U29027 ( .I(n9035), .ZN(n56928) );
  NAND2_X1 U29028 ( .A1(n9035), .A2(n1583), .ZN(n56937) );
  NAND2_X1 U29029 ( .A1(n17850), .A2(n9035), .ZN(n56945) );
  NAND2_X1 U29031 ( .A1(n10038), .A2(n9035), .ZN(n10383) );
  OAI22_X1 U29032 ( .A1(n56929), .A2(n9035), .B1(n63420), .B2(n56952), .ZN(
        n56930) );
  XOR2_X1 U29039 ( .A1(n9044), .A2(n51291), .Z(n14946) );
  OAI21_X1 U29041 ( .A1(n24081), .A2(n62788), .B(n59008), .ZN(n47750) );
  NOR2_X1 U29042 ( .A1(n47434), .A2(n62788), .ZN(n45907) );
  NOR2_X1 U29043 ( .A1(n47431), .A2(n62788), .ZN(n15419) );
  INV_X2 U29044 ( .I(n43748), .ZN(n9046) );
  INV_X1 U29045 ( .I(n14773), .ZN(n25661) );
  INV_X2 U29048 ( .I(n9049), .ZN(n19102) );
  XOR2_X1 U29049 ( .A1(n13272), .A2(n57174), .Z(n9050) );
  XOR2_X1 U29055 ( .A1(n9055), .A2(n32508), .Z(n32509) );
  XOR2_X1 U29056 ( .A1(n13740), .A2(n9055), .Z(n12415) );
  XOR2_X1 U29057 ( .A1(n9060), .A2(n9057), .Z(n24226) );
  XOR2_X1 U29058 ( .A1(n9058), .A2(n50849), .Z(n9057) );
  XOR2_X1 U29059 ( .A1(n354), .A2(n64316), .Z(n9058) );
  XOR2_X1 U29060 ( .A1(n9059), .A2(n47652), .Z(n50849) );
  XOR2_X1 U29061 ( .A1(n52325), .A2(n24076), .Z(n9059) );
  NOR2_X1 U29065 ( .A1(n10562), .A2(n10277), .ZN(n19417) );
  NAND2_X1 U29067 ( .A1(n9068), .A2(n5051), .ZN(n55061) );
  NAND2_X1 U29070 ( .A1(n55075), .A2(n9068), .ZN(n9096) );
  XOR2_X1 U29074 ( .A1(n9072), .A2(n25012), .Z(n9071) );
  NOR2_X1 U29075 ( .A1(n65283), .A2(n1609), .ZN(n9075) );
  XOR2_X1 U29077 ( .A1(n3449), .A2(n46271), .Z(n14910) );
  XOR2_X1 U29078 ( .A1(n9079), .A2(n8813), .Z(n46677) );
  OAI21_X1 U29080 ( .A1(n22900), .A2(n24009), .B(n9082), .ZN(n55019) );
  NAND2_X1 U29081 ( .A1(n9082), .A2(n7148), .ZN(n52639) );
  NAND3_X1 U29082 ( .A1(n9082), .A2(n59713), .A3(n17935), .ZN(n54638) );
  NOR2_X1 U29083 ( .A1(n47449), .A2(n11950), .ZN(n21335) );
  INV_X1 U29086 ( .I(n10677), .ZN(n15476) );
  XOR2_X1 U29087 ( .A1(n44886), .A2(n19543), .Z(n21624) );
  INV_X4 U29088 ( .I(n17978), .ZN(n19118) );
  NOR2_X2 U29090 ( .A1(n7118), .A2(n20867), .ZN(n36201) );
  INV_X4 U29092 ( .I(n38273), .ZN(n42230) );
  INV_X1 U29093 ( .I(n43350), .ZN(n43355) );
  NAND2_X2 U29098 ( .A1(n40026), .A2(n23477), .ZN(n40303) );
  INV_X1 U29101 ( .I(n18231), .ZN(n18200) );
  XOR2_X1 U29102 ( .A1(n4651), .A2(n9110), .Z(n9109) );
  XOR2_X1 U29103 ( .A1(n33258), .A2(n15735), .Z(n9110) );
  AOI22_X1 U29105 ( .A1(n55925), .A2(n10040), .B1(n9111), .B2(n55926), .ZN(
        n55928) );
  OAI21_X1 U29106 ( .A1(n61627), .A2(n56313), .B(n20957), .ZN(n9117) );
  INV_X2 U29107 ( .I(n9118), .ZN(n9524) );
  NOR2_X2 U29108 ( .A1(n24138), .A2(n13912), .ZN(n45386) );
  INV_X2 U29110 ( .I(n12129), .ZN(n18829) );
  XOR2_X1 U29111 ( .A1(n14553), .A2(n19410), .Z(n39368) );
  XOR2_X1 U29112 ( .A1(n39246), .A2(n39245), .Z(n9120) );
  NAND2_X2 U29117 ( .A1(n13982), .A2(n34632), .ZN(n35032) );
  NAND3_X1 U29121 ( .A1(n29335), .A2(n29351), .A3(n58977), .ZN(n9138) );
  NAND2_X2 U29123 ( .A1(n19452), .A2(n27501), .ZN(n29338) );
  INV_X2 U29127 ( .I(n35146), .ZN(n35144) );
  NOR2_X2 U29128 ( .A1(n34478), .A2(n35970), .ZN(n35146) );
  NAND2_X2 U29129 ( .A1(n21018), .A2(n15754), .ZN(n35970) );
  XOR2_X1 U29131 ( .A1(n9148), .A2(n9145), .Z(n38336) );
  XOR2_X1 U29132 ( .A1(n9147), .A2(n9146), .Z(n9145) );
  XOR2_X1 U29133 ( .A1(n60489), .A2(n17938), .Z(n9146) );
  XOR2_X1 U29134 ( .A1(n19145), .A2(n38299), .Z(n9147) );
  XOR2_X1 U29135 ( .A1(n44268), .A2(n44267), .Z(n9149) );
  XOR2_X1 U29137 ( .A1(n11614), .A2(n21521), .Z(n13658) );
  NOR2_X2 U29140 ( .A1(n9152), .A2(n48594), .ZN(n47017) );
  AOI22_X1 U29143 ( .A1(n47529), .A2(n9152), .B1(n47535), .B2(n62115), .ZN(
        n44694) );
  XOR2_X1 U29145 ( .A1(n11448), .A2(n9154), .Z(n11447) );
  XOR2_X1 U29146 ( .A1(n55624), .A2(n9154), .Z(n51475) );
  XOR2_X1 U29147 ( .A1(n23213), .A2(n9154), .Z(n50590) );
  NOR2_X2 U29149 ( .A1(n21759), .A2(n21758), .ZN(n44077) );
  XOR2_X1 U29150 ( .A1(n9158), .A2(n25787), .Z(n9159) );
  NAND2_X1 U29151 ( .A1(n25267), .A2(n53795), .ZN(n53780) );
  NAND3_X2 U29153 ( .A1(n1706), .A2(n43980), .A3(n23314), .ZN(n9163) );
  NOR2_X2 U29154 ( .A1(n1547), .A2(n5410), .ZN(n34003) );
  NAND2_X2 U29159 ( .A1(n25619), .A2(n10403), .ZN(n26977) );
  NOR2_X2 U29167 ( .A1(n35898), .A2(n9721), .ZN(n35561) );
  XOR2_X1 U29170 ( .A1(n7573), .A2(n37485), .Z(n37487) );
  XOR2_X1 U29171 ( .A1(n7573), .A2(n22170), .Z(n38580) );
  XOR2_X1 U29172 ( .A1(n32648), .A2(n750), .Z(n14715) );
  INV_X2 U29175 ( .I(n9216), .ZN(n36648) );
  NOR2_X1 U29178 ( .A1(n1859), .A2(n9186), .ZN(n29413) );
  NOR2_X1 U29181 ( .A1(n22786), .A2(n9189), .ZN(n39091) );
  AOI21_X1 U29182 ( .A1(n41030), .A2(n22617), .B(n9189), .ZN(n41032) );
  NAND2_X1 U29183 ( .A1(n40517), .A2(n9189), .ZN(n40518) );
  XOR2_X1 U29189 ( .A1(n9193), .A2(n9192), .Z(n9519) );
  XOR2_X1 U29190 ( .A1(n50937), .A2(n51960), .Z(n9194) );
  NAND2_X2 U29196 ( .A1(n9197), .A2(n61729), .ZN(n23111) );
  NAND2_X1 U29197 ( .A1(n30084), .A2(n9197), .ZN(n9335) );
  OAI21_X1 U29199 ( .A1(n27916), .A2(n9197), .B(n9287), .ZN(n27917) );
  INV_X4 U29200 ( .I(n29794), .ZN(n9197) );
  NAND2_X2 U29201 ( .A1(n12863), .A2(n20812), .ZN(n35422) );
  XOR2_X1 U29202 ( .A1(n20573), .A2(n15662), .Z(n17921) );
  NAND3_X2 U29204 ( .A1(n42607), .A2(n42608), .A3(n429), .ZN(n9211) );
  XOR2_X1 U29211 ( .A1(n46701), .A2(n21940), .Z(n15561) );
  XOR2_X1 U29212 ( .A1(n9222), .A2(n1045), .Z(n9221) );
  XOR2_X1 U29213 ( .A1(n8381), .A2(n25594), .Z(n9222) );
  NAND2_X1 U29214 ( .A1(n47719), .A2(n47718), .ZN(n9226) );
  XOR2_X1 U29220 ( .A1(n46228), .A2(n14674), .Z(n9244) );
  XOR2_X1 U29221 ( .A1(n45237), .A2(n15562), .Z(n46228) );
  XOR2_X1 U29223 ( .A1(n46227), .A2(n46226), .Z(n9246) );
  OAI22_X1 U29226 ( .A1(n29786), .A2(n9250), .B1(n29254), .B2(n29251), .ZN(
        n29252) );
  OAI22_X1 U29227 ( .A1(n29781), .A2(n9250), .B1(n29787), .B2(n29782), .ZN(
        n29791) );
  INV_X2 U29230 ( .I(n9254), .ZN(n33828) );
  XOR2_X1 U29231 ( .A1(n44035), .A2(n44037), .Z(n9259) );
  NAND2_X1 U29232 ( .A1(n26673), .A2(n26674), .ZN(n9260) );
  XOR2_X1 U29233 ( .A1(n61498), .A2(n44033), .Z(n44034) );
  XOR2_X1 U29234 ( .A1(n61498), .A2(n44742), .Z(n44743) );
  XOR2_X1 U29235 ( .A1(n61498), .A2(n46596), .Z(n46597) );
  AND2_X1 U29243 ( .A1(n32920), .A2(n32921), .Z(n9277) );
  NAND2_X2 U29245 ( .A1(n15622), .A2(n30092), .ZN(n32324) );
  INV_X2 U29247 ( .I(n9285), .ZN(n55671) );
  NAND2_X2 U29248 ( .A1(n24091), .A2(n55671), .ZN(n23900) );
  NAND3_X1 U29252 ( .A1(n9291), .A2(n64341), .A3(n17334), .ZN(n9290) );
  NAND2_X1 U29253 ( .A1(n49498), .A2(n49501), .ZN(n9291) );
  NAND2_X1 U29254 ( .A1(n42600), .A2(n60657), .ZN(n9295) );
  NAND2_X1 U29255 ( .A1(n53591), .A2(n9296), .ZN(n53592) );
  XOR2_X1 U29257 ( .A1(n51387), .A2(n9298), .Z(n9297) );
  XOR2_X1 U29258 ( .A1(n50576), .A2(n12006), .Z(n51003) );
  XOR2_X1 U29259 ( .A1(n19785), .A2(n50167), .Z(n51387) );
  XOR2_X1 U29260 ( .A1(n51033), .A2(n1576), .Z(n19785) );
  NAND2_X1 U29261 ( .A1(n45740), .A2(n9299), .ZN(n10184) );
  NOR3_X2 U29263 ( .A1(n9390), .A2(n19017), .A3(n9301), .ZN(n19018) );
  NAND3_X2 U29264 ( .A1(n57164), .A2(n34731), .A3(n9302), .ZN(n9301) );
  NOR3_X2 U29266 ( .A1(n18554), .A2(n18553), .A3(n37923), .ZN(n46497) );
  NOR2_X1 U29269 ( .A1(n21467), .A2(n9304), .ZN(n36199) );
  NAND2_X1 U29270 ( .A1(n36724), .A2(n9304), .ZN(n36727) );
  OAI22_X1 U29271 ( .A1(n36204), .A2(n9304), .B1(n26243), .B2(n36203), .ZN(
        n36205) );
  XOR2_X1 U29274 ( .A1(n18434), .A2(n32324), .Z(n22162) );
  INV_X2 U29275 ( .I(n9307), .ZN(n19556) );
  NAND2_X1 U29282 ( .A1(n17620), .A2(n23163), .ZN(n56477) );
  XOR2_X1 U29285 ( .A1(n24012), .A2(n9315), .Z(n9345) );
  XOR2_X1 U29286 ( .A1(n9317), .A2(n9316), .Z(n9315) );
  XOR2_X1 U29287 ( .A1(n62740), .A2(n32629), .Z(n9316) );
  XOR2_X1 U29288 ( .A1(n9318), .A2(n20554), .Z(n9317) );
  XOR2_X1 U29289 ( .A1(n23706), .A2(n32627), .Z(n9318) );
  INV_X1 U29291 ( .I(n48280), .ZN(n48829) );
  INV_X1 U29294 ( .I(n48828), .ZN(n9321) );
  INV_X1 U29295 ( .I(n48022), .ZN(n9322) );
  INV_X1 U29296 ( .I(n9339), .ZN(n9327) );
  OAI21_X1 U29298 ( .A1(n39801), .A2(n39800), .B(n14846), .ZN(n9365) );
  AOI21_X1 U29300 ( .A1(n28786), .A2(n28785), .B(n17794), .ZN(n9339) );
  XOR2_X1 U29303 ( .A1(n10352), .A2(n12791), .Z(n9342) );
  XOR2_X1 U29304 ( .A1(n12524), .A2(n811), .Z(n16898) );
  XOR2_X1 U29305 ( .A1(n24247), .A2(n9343), .Z(n24162) );
  INV_X1 U29306 ( .I(n12524), .ZN(n9343) );
  INV_X1 U29307 ( .I(n9344), .ZN(n27593) );
  NAND2_X1 U29308 ( .A1(n28302), .A2(n9344), .ZN(n27598) );
  OAI21_X1 U29309 ( .A1(n27081), .A2(n27080), .B(n9344), .ZN(n27082) );
  NAND2_X2 U29310 ( .A1(n20437), .A2(n26641), .ZN(n9344) );
  INV_X2 U29311 ( .I(n9345), .ZN(n19373) );
  NAND2_X2 U29312 ( .A1(n17255), .A2(n19373), .ZN(n33542) );
  INV_X1 U29313 ( .I(n40864), .ZN(n41638) );
  INV_X2 U29315 ( .I(n9355), .ZN(n24318) );
  INV_X2 U29316 ( .I(n25997), .ZN(n57048) );
  XOR2_X1 U29318 ( .A1(n9357), .A2(n32395), .Z(n9356) );
  XOR2_X1 U29319 ( .A1(n31749), .A2(n32399), .Z(n9357) );
  NAND3_X2 U29322 ( .A1(n23659), .A2(n49306), .A3(n49305), .ZN(n52174) );
  AND2_X1 U29323 ( .A1(n41751), .A2(n9366), .Z(n22753) );
  NAND2_X2 U29324 ( .A1(n25232), .A2(n23900), .ZN(n15244) );
  NAND2_X1 U29325 ( .A1(n14142), .A2(n23900), .ZN(n14141) );
  OAI21_X1 U29326 ( .A1(n16018), .A2(n60553), .B(n23900), .ZN(n24903) );
  OAI22_X2 U29329 ( .A1(n15183), .A2(n1536), .B1(n15184), .B2(n63250), .ZN(
        n15182) );
  XOR2_X1 U29331 ( .A1(n21494), .A2(n9370), .Z(n12774) );
  XOR2_X1 U29332 ( .A1(n38106), .A2(n9371), .Z(n9370) );
  NAND2_X2 U29335 ( .A1(n19018), .A2(n34732), .ZN(n9372) );
  XNOR2_X1 U29336 ( .A1(n16936), .A2(n24292), .ZN(n9373) );
  NAND2_X2 U29338 ( .A1(n9375), .A2(n23333), .ZN(n37866) );
  NAND3_X2 U29341 ( .A1(n10153), .A2(n10152), .A3(n13123), .ZN(n9378) );
  XOR2_X1 U29342 ( .A1(n1684), .A2(n59382), .Z(n10776) );
  OR2_X1 U29343 ( .A1(n9386), .A2(n52053), .Z(n9381) );
  NAND2_X2 U29348 ( .A1(n63249), .A2(n32934), .ZN(n34730) );
  NAND2_X1 U29351 ( .A1(n11987), .A2(n9392), .ZN(n27764) );
  OAI21_X1 U29352 ( .A1(n5070), .A2(n9392), .B(n28898), .ZN(n28901) );
  NOR2_X1 U29353 ( .A1(n29816), .A2(n9392), .ZN(n29817) );
  INV_X2 U29355 ( .I(n12426), .ZN(n17967) );
  NAND2_X2 U29360 ( .A1(n20000), .A2(n56423), .ZN(n23163) );
  INV_X2 U29361 ( .I(n37556), .ZN(n39259) );
  XOR2_X1 U29362 ( .A1(n9399), .A2(n9397), .Z(n38466) );
  XOR2_X1 U29363 ( .A1(n9400), .A2(n9398), .Z(n9399) );
  NAND2_X2 U29364 ( .A1(n37194), .A2(n37193), .ZN(n22988) );
  XOR2_X1 U29366 ( .A1(n9401), .A2(n55349), .Z(Plaintext[110]) );
  NOR2_X1 U29368 ( .A1(n55346), .A2(n55345), .ZN(n9404) );
  NAND2_X2 U29369 ( .A1(n9410), .A2(n22891), .ZN(n56347) );
  OAI22_X1 U29370 ( .A1(n56300), .A2(n11654), .B1(n20957), .B2(n9410), .ZN(
        n56301) );
  NAND2_X2 U29372 ( .A1(n11987), .A2(n463), .ZN(n30475) );
  XOR2_X1 U29373 ( .A1(n21508), .A2(n9412), .Z(n9415) );
  XOR2_X1 U29374 ( .A1(n9413), .A2(n21494), .Z(n21508) );
  XOR2_X1 U29375 ( .A1(n57452), .A2(n38106), .Z(n9413) );
  INV_X4 U29376 ( .I(n7728), .ZN(n42251) );
  XOR2_X1 U29377 ( .A1(n9417), .A2(n23069), .Z(n52086) );
  XOR2_X1 U29378 ( .A1(n19349), .A2(n11070), .Z(n9417) );
  OAI21_X1 U29379 ( .A1(n9418), .A2(n18258), .B(n55438), .ZN(n18257) );
  INV_X2 U29381 ( .I(n18145), .ZN(n9418) );
  XOR2_X1 U29382 ( .A1(n9420), .A2(n23902), .Z(n9419) );
  XOR2_X1 U29383 ( .A1(n45341), .A2(n44538), .Z(n9420) );
  NAND2_X2 U29389 ( .A1(n8912), .A2(n42827), .ZN(n41369) );
  XOR2_X1 U29392 ( .A1(n9428), .A2(n31611), .Z(n9430) );
  XOR2_X1 U29394 ( .A1(n9433), .A2(n30993), .Z(n9432) );
  XOR2_X1 U29395 ( .A1(n30992), .A2(n25401), .Z(n9433) );
  XOR2_X1 U29396 ( .A1(n53764), .A2(n4921), .Z(n51407) );
  XOR2_X1 U29397 ( .A1(n54563), .A2(n9434), .Z(n39349) );
  XOR2_X1 U29398 ( .A1(n55638), .A2(n9435), .Z(n44270) );
  XOR2_X1 U29399 ( .A1(n56508), .A2(n9435), .Z(n37254) );
  XOR2_X1 U29400 ( .A1(n44796), .A2(n9434), .Z(n33195) );
  XOR2_X1 U29401 ( .A1(n37499), .A2(n9434), .Z(n48954) );
  XOR2_X1 U29402 ( .A1(n33203), .A2(n9434), .Z(n19479) );
  XOR2_X1 U29404 ( .A1(n22640), .A2(n9434), .Z(Plaintext[64]) );
  INV_X1 U29409 ( .I(n47718), .ZN(n9453) );
  INV_X1 U29410 ( .I(n9455), .ZN(n48963) );
  NOR2_X1 U29411 ( .A1(n9455), .A2(n49410), .ZN(n49268) );
  NAND2_X2 U29414 ( .A1(n9461), .A2(n9457), .ZN(n24228) );
  XOR2_X1 U29415 ( .A1(n31518), .A2(n9462), .Z(n13833) );
  AOI21_X1 U29418 ( .A1(n26592), .A2(n16021), .B(n9465), .ZN(n26588) );
  NAND2_X2 U29420 ( .A1(n25785), .A2(n27478), .ZN(n9473) );
  OAI21_X1 U29421 ( .A1(n9473), .A2(n27543), .B(n27479), .ZN(n26477) );
  OAI21_X1 U29422 ( .A1(n9473), .A2(n26935), .B(n14869), .ZN(n26476) );
  NOR2_X1 U29423 ( .A1(n23474), .A2(n9473), .ZN(n27472) );
  NAND2_X2 U29424 ( .A1(n20509), .A2(n9473), .ZN(n16788) );
  NOR2_X1 U29425 ( .A1(n26936), .A2(n9473), .ZN(n26482) );
  AOI22_X1 U29426 ( .A1(n26705), .A2(n9473), .B1(n27538), .B2(n4617), .ZN(
        n16794) );
  XOR2_X1 U29429 ( .A1(n14878), .A2(n38467), .Z(n24891) );
  AOI21_X1 U29433 ( .A1(n61186), .A2(n59139), .B(n43327), .ZN(n41464) );
  NOR2_X2 U29435 ( .A1(n9475), .A2(n58710), .ZN(n29778) );
  NOR2_X1 U29437 ( .A1(n48642), .A2(n3091), .ZN(n48647) );
  NAND2_X1 U29438 ( .A1(n23416), .A2(n3091), .ZN(n48166) );
  INV_X2 U29440 ( .I(n23862), .ZN(n53265) );
  INV_X4 U29441 ( .I(n9482), .ZN(n15171) );
  NAND2_X2 U29443 ( .A1(n9482), .A2(n3129), .ZN(n36921) );
  INV_X1 U29444 ( .I(n10884), .ZN(n9483) );
  XOR2_X1 U29445 ( .A1(n31382), .A2(n843), .Z(n9484) );
  XOR2_X1 U29446 ( .A1(n23069), .A2(n9485), .Z(n50941) );
  XOR2_X1 U29447 ( .A1(n19349), .A2(n1900), .Z(n9485) );
  INV_X2 U29449 ( .I(n9488), .ZN(n41019) );
  NOR2_X2 U29451 ( .A1(n1512), .A2(n12523), .ZN(n41006) );
  XNOR2_X1 U29452 ( .A1(n14681), .A2(n14682), .ZN(n9488) );
  XOR2_X1 U29454 ( .A1(n9492), .A2(n9491), .Z(n12596) );
  XOR2_X1 U29455 ( .A1(n37866), .A2(n51604), .Z(n36992) );
  XOR2_X1 U29458 ( .A1(n9497), .A2(n9496), .Z(n25847) );
  NAND2_X1 U29466 ( .A1(n9504), .A2(n42572), .ZN(n42574) );
  NAND2_X2 U29469 ( .A1(n22549), .A2(n47270), .ZN(n9505) );
  XOR2_X1 U29471 ( .A1(n9506), .A2(n50988), .Z(n50989) );
  XOR2_X1 U29472 ( .A1(n51626), .A2(n9506), .Z(n51627) );
  INV_X2 U29474 ( .I(n9508), .ZN(n51860) );
  NOR2_X2 U29475 ( .A1(n51860), .A2(n51870), .ZN(n54028) );
  XNOR2_X1 U29476 ( .A1(n9510), .A2(n9509), .ZN(n9508) );
  XOR2_X1 U29478 ( .A1(n60448), .A2(n50862), .Z(n9510) );
  XOR2_X1 U29479 ( .A1(n11209), .A2(n11208), .Z(n54021) );
  OAI21_X1 U29481 ( .A1(n9511), .A2(n22989), .B(n4274), .ZN(n20283) );
  NOR2_X1 U29486 ( .A1(n18522), .A2(n9514), .ZN(n18521) );
  AOI21_X1 U29488 ( .A1(n52782), .A2(n53622), .B(n9514), .ZN(n52783) );
  INV_X2 U29490 ( .I(n32975), .ZN(n34786) );
  NOR3_X1 U29491 ( .A1(n33776), .A2(n7116), .A3(n18503), .ZN(n9515) );
  INV_X2 U29492 ( .I(n26039), .ZN(n32560) );
  NAND2_X1 U29493 ( .A1(n53322), .A2(n63931), .ZN(n53323) );
  OAI22_X1 U29495 ( .A1(n15405), .A2(n63931), .B1(n17012), .B2(n53348), .ZN(
        n15404) );
  INV_X2 U29497 ( .I(n9519), .ZN(n52126) );
  NAND2_X1 U29500 ( .A1(n42358), .A2(n9522), .ZN(n23340) );
  XOR2_X1 U29501 ( .A1(n42355), .A2(n1301), .Z(n9523) );
  INV_X4 U29504 ( .I(n9525), .ZN(n16850) );
  INV_X1 U29507 ( .I(n4422), .ZN(n19502) );
  XOR2_X1 U29508 ( .A1(n4422), .A2(n37300), .Z(n37980) );
  NAND2_X1 U29510 ( .A1(n14306), .A2(n57199), .ZN(n40507) );
  XOR2_X1 U29511 ( .A1(n46493), .A2(n55833), .Z(n9530) );
  NAND2_X2 U29512 ( .A1(n41574), .A2(n41575), .ZN(n46493) );
  INV_X2 U29513 ( .I(n9531), .ZN(n47501) );
  INV_X2 U29516 ( .I(n26185), .ZN(n52559) );
  XOR2_X1 U29517 ( .A1(n52612), .A2(n52620), .Z(n21963) );
  XOR2_X1 U29518 ( .A1(n9546), .A2(n9545), .Z(n52612) );
  XOR2_X1 U29519 ( .A1(n26185), .A2(n9547), .Z(n9546) );
  XOR2_X1 U29520 ( .A1(n52325), .A2(n53090), .Z(n9547) );
  XOR2_X1 U29521 ( .A1(Ciphertext[6]), .A2(Key[31]), .Z(n13826) );
  INV_X1 U29528 ( .I(n185), .ZN(n51593) );
  NAND2_X2 U29529 ( .A1(n9553), .A2(n9552), .ZN(n25192) );
  XOR2_X1 U29531 ( .A1(n59063), .A2(n44955), .Z(n14295) );
  XOR2_X1 U29532 ( .A1(n9554), .A2(n24449), .Z(n44955) );
  XOR2_X1 U29533 ( .A1(n23162), .A2(n24098), .Z(n9554) );
  INV_X1 U29534 ( .I(n9555), .ZN(n56379) );
  OAI22_X1 U29535 ( .A1(n52241), .A2(n13489), .B1(n23095), .B2(n9555), .ZN(
        n52246) );
  NAND2_X1 U29537 ( .A1(n56529), .A2(n9555), .ZN(n22370) );
  AOI21_X1 U29538 ( .A1(n21732), .A2(n9555), .B(n56545), .ZN(n16689) );
  XOR2_X1 U29540 ( .A1(n52031), .A2(n51172), .Z(n9557) );
  OR2_X1 U29542 ( .A1(n56738), .A2(n56718), .Z(n9559) );
  NAND3_X1 U29543 ( .A1(n20269), .A2(n56733), .A3(n23785), .ZN(n56699) );
  OAI21_X1 U29544 ( .A1(n20128), .A2(n56733), .B(n56698), .ZN(n9560) );
  NOR2_X2 U29545 ( .A1(n56719), .A2(n56733), .ZN(n56738) );
  XOR2_X1 U29550 ( .A1(n9575), .A2(n9571), .Z(n9610) );
  XOR2_X1 U29551 ( .A1(n19411), .A2(n9572), .Z(n9571) );
  XOR2_X1 U29552 ( .A1(n9574), .A2(n9573), .Z(n9572) );
  XOR2_X1 U29553 ( .A1(n44738), .A2(n21141), .Z(n9573) );
  XOR2_X1 U29554 ( .A1(n45401), .A2(n44743), .Z(n9574) );
  NAND2_X1 U29556 ( .A1(n30441), .A2(n23053), .ZN(n9581) );
  NAND2_X2 U29557 ( .A1(n9583), .A2(n9582), .ZN(n15808) );
  XOR2_X1 U29560 ( .A1(n26142), .A2(n15865), .Z(n9586) );
  INV_X2 U29561 ( .I(n10583), .ZN(n15865) );
  NOR2_X2 U29564 ( .A1(n13029), .A2(n22283), .ZN(n16882) );
  INV_X1 U29566 ( .I(n9590), .ZN(n9589) );
  NOR2_X1 U29567 ( .A1(n17280), .A2(n60839), .ZN(n46105) );
  NAND2_X1 U29568 ( .A1(n48247), .A2(n60839), .ZN(n16418) );
  NAND2_X1 U29569 ( .A1(n9593), .A2(n20060), .ZN(n34853) );
  NOR2_X1 U29570 ( .A1(n9593), .A2(n36777), .ZN(n34857) );
  OAI21_X1 U29572 ( .A1(n9593), .A2(n36775), .B(n36777), .ZN(n20310) );
  NOR2_X2 U29575 ( .A1(n25791), .A2(n25790), .ZN(n49493) );
  NOR2_X2 U29576 ( .A1(n53492), .A2(n9595), .ZN(n53526) );
  XOR2_X1 U29579 ( .A1(n11665), .A2(n38658), .Z(n9603) );
  INV_X2 U29582 ( .I(n9607), .ZN(n10064) );
  XOR2_X1 U29583 ( .A1(n20719), .A2(n16625), .Z(n31518) );
  INV_X2 U29584 ( .I(n9610), .ZN(n22283) );
  NAND2_X1 U29587 ( .A1(n50337), .A2(n49973), .ZN(n20857) );
  XOR2_X1 U29590 ( .A1(n52154), .A2(n50765), .Z(n9615) );
  NOR2_X2 U29593 ( .A1(n11959), .A2(n38672), .ZN(n24977) );
  XNOR2_X1 U29595 ( .A1(n17803), .A2(n17802), .ZN(n9659) );
  NAND3_X1 U29596 ( .A1(n41189), .A2(n41190), .A3(n64858), .ZN(n22330) );
  INV_X2 U29597 ( .I(n18376), .ZN(n19953) );
  NAND2_X2 U29598 ( .A1(n15717), .A2(n11789), .ZN(n18376) );
  OAI21_X1 U29601 ( .A1(n39946), .A2(n10041), .B(n23420), .ZN(n39953) );
  AND2_X1 U29604 ( .A1(n16525), .A2(n27841), .Z(n16524) );
  XOR2_X1 U29605 ( .A1(n3715), .A2(n37564), .Z(n17346) );
  INV_X1 U29606 ( .I(n30121), .ZN(n29772) );
  INV_X1 U29608 ( .I(n28795), .ZN(n13945) );
  INV_X4 U29610 ( .I(n47034), .ZN(n20299) );
  XOR2_X1 U29616 ( .A1(Ciphertext[112]), .A2(Key[5]), .Z(n10347) );
  XOR2_X1 U29617 ( .A1(n9621), .A2(n45858), .Z(n11725) );
  XOR2_X1 U29618 ( .A1(n45859), .A2(n14373), .Z(n9621) );
  XOR2_X1 U29619 ( .A1(n17983), .A2(n9622), .Z(n44368) );
  XOR2_X1 U29620 ( .A1(n24021), .A2(n44366), .Z(n9622) );
  NAND2_X1 U29621 ( .A1(n19266), .A2(n28935), .ZN(n25181) );
  OR3_X2 U29627 ( .A1(n42123), .A2(n42122), .A3(n42124), .Z(n13912) );
  NAND2_X1 U29629 ( .A1(n29517), .A2(n29858), .ZN(n9821) );
  OAI22_X1 U29630 ( .A1(n17458), .A2(n28802), .B1(n17459), .B2(n10625), .ZN(
        n9629) );
  XOR2_X1 U29632 ( .A1(n22160), .A2(n31835), .Z(n18542) );
  XOR2_X1 U29636 ( .A1(n44155), .A2(n43672), .Z(n9637) );
  NAND3_X2 U29637 ( .A1(n9638), .A2(n11333), .A3(n26891), .ZN(n30148) );
  AND3_X1 U29638 ( .A1(n26889), .A2(n26892), .A3(n26890), .Z(n9638) );
  OR2_X1 U29639 ( .A1(n55310), .A2(n55442), .Z(n55318) );
  NAND3_X2 U29642 ( .A1(n9641), .A2(n30711), .A3(n30713), .ZN(n33906) );
  AND2_X1 U29643 ( .A1(n30714), .A2(n30712), .Z(n9641) );
  BUF_X2 U29647 ( .I(n4734), .Z(n9646) );
  XOR2_X1 U29649 ( .A1(n15261), .A2(n51701), .Z(n15260) );
  INV_X4 U29650 ( .I(n15060), .ZN(n21364) );
  NOR2_X2 U29651 ( .A1(n40654), .A2(n41183), .ZN(n39141) );
  INV_X2 U29652 ( .I(n25956), .ZN(n48536) );
  OAI21_X1 U29653 ( .A1(n9653), .A2(n25987), .B(n9652), .ZN(n52292) );
  NAND2_X1 U29654 ( .A1(n56924), .A2(n25987), .ZN(n9652) );
  BUF_X2 U29655 ( .I(n52278), .Z(n9655) );
  AND2_X1 U29659 ( .A1(n41254), .A2(n24195), .Z(n43892) );
  INV_X1 U29660 ( .I(n38343), .ZN(n9894) );
  NOR2_X1 U29661 ( .A1(n36136), .A2(n36137), .ZN(n36144) );
  XOR2_X1 U29662 ( .A1(n11242), .A2(n9659), .Z(n11241) );
  INV_X2 U29665 ( .I(n19040), .ZN(n47482) );
  NAND2_X2 U29666 ( .A1(n26145), .A2(n16616), .ZN(n19040) );
  XOR2_X1 U29667 ( .A1(n9662), .A2(n12762), .Z(n12186) );
  XOR2_X1 U29668 ( .A1(n20670), .A2(n32098), .Z(n9662) );
  OR3_X1 U29670 ( .A1(n42978), .A2(n43326), .A3(n59139), .Z(n42982) );
  XOR2_X1 U29673 ( .A1(n63033), .A2(n24379), .Z(n9664) );
  XOR2_X1 U29674 ( .A1(n9665), .A2(n15332), .Z(n33277) );
  NAND2_X1 U29676 ( .A1(n27254), .A2(n26761), .ZN(n26762) );
  XOR2_X1 U29677 ( .A1(n9666), .A2(n20617), .Z(n11382) );
  XOR2_X1 U29678 ( .A1(n11231), .A2(n11230), .Z(n11233) );
  XOR2_X1 U29679 ( .A1(n37777), .A2(n9667), .Z(n37783) );
  NOR2_X2 U29682 ( .A1(n24337), .A2(n24336), .ZN(n25952) );
  NAND2_X2 U29683 ( .A1(n25953), .A2(n22761), .ZN(n24337) );
  XOR2_X1 U29684 ( .A1(n51941), .A2(n9673), .Z(n51942) );
  XOR2_X1 U29685 ( .A1(n52472), .A2(n22614), .Z(n9673) );
  XOR2_X1 U29687 ( .A1(n44417), .A2(n14760), .Z(n9674) );
  NOR2_X2 U29688 ( .A1(n17452), .A2(n23331), .ZN(n21177) );
  NOR2_X1 U29691 ( .A1(n7588), .A2(n12474), .ZN(n12473) );
  NAND2_X1 U29694 ( .A1(n27436), .A2(n10625), .ZN(n26998) );
  NAND2_X2 U29695 ( .A1(n23773), .A2(n27435), .ZN(n18515) );
  BUF_X2 U29696 ( .I(n22597), .Z(n9679) );
  OAI22_X1 U29698 ( .A1(n29672), .A2(n29673), .B1(n29675), .B2(n29674), .ZN(
        n29676) );
  BUF_X4 U29700 ( .I(n49565), .Z(n18975) );
  MUX2_X1 U29701 ( .I0(n31951), .I1(n35251), .S(n7345), .Z(n31953) );
  XOR2_X1 U29704 ( .A1(n10229), .A2(n19282), .Z(n13947) );
  NOR2_X2 U29706 ( .A1(n27441), .A2(n27435), .ZN(n17824) );
  XOR2_X1 U29707 ( .A1(n33042), .A2(n9682), .Z(n22921) );
  XOR2_X1 U29708 ( .A1(n30998), .A2(n9683), .Z(n9682) );
  INV_X4 U29709 ( .I(n22556), .ZN(n29824) );
  AND3_X1 U29712 ( .A1(n20767), .A2(n43710), .A3(n43711), .Z(n12742) );
  XOR2_X1 U29714 ( .A1(n51084), .A2(n9690), .Z(n51085) );
  XOR2_X1 U29715 ( .A1(n51761), .A2(n51083), .Z(n9690) );
  XOR2_X1 U29717 ( .A1(n9691), .A2(n14251), .Z(n23740) );
  XOR2_X1 U29718 ( .A1(n44898), .A2(n12607), .Z(n9691) );
  NAND2_X1 U29720 ( .A1(n10563), .A2(n64823), .ZN(n9692) );
  BUF_X2 U29721 ( .I(n25332), .Z(n25331) );
  XOR2_X1 U29723 ( .A1(n37146), .A2(n37147), .Z(n9693) );
  OR2_X2 U29725 ( .A1(n47552), .A2(n47553), .Z(n25857) );
  NAND3_X2 U29726 ( .A1(n24384), .A2(n13994), .A3(n13996), .ZN(n39579) );
  INV_X1 U29728 ( .I(n35910), .ZN(n35905) );
  XNOR2_X1 U29729 ( .A1(n31454), .A2(n31453), .ZN(n24831) );
  XOR2_X1 U29731 ( .A1(n26202), .A2(n32724), .Z(n12107) );
  INV_X2 U29736 ( .I(n9703), .ZN(n11655) );
  XOR2_X1 U29737 ( .A1(Ciphertext[129]), .A2(Key[28]), .Z(n9703) );
  XOR2_X1 U29741 ( .A1(n32714), .A2(n10430), .Z(n9707) );
  XOR2_X1 U29742 ( .A1(n14037), .A2(n9708), .Z(n14292) );
  XOR2_X1 U29743 ( .A1(n43409), .A2(n41501), .Z(n9708) );
  XOR2_X1 U29745 ( .A1(n9710), .A2(n45285), .Z(n9709) );
  XOR2_X1 U29748 ( .A1(n17463), .A2(n23726), .Z(n9712) );
  XOR2_X1 U29752 ( .A1(n32615), .A2(n9714), .Z(n32712) );
  AND2_X1 U29756 ( .A1(n29209), .A2(n26740), .Z(n28781) );
  NOR2_X1 U29757 ( .A1(n41035), .A2(n36106), .ZN(n21162) );
  NAND2_X2 U29759 ( .A1(n45628), .A2(n10078), .ZN(n49076) );
  XOR2_X1 U29760 ( .A1(n38501), .A2(n37743), .Z(n23147) );
  AOI21_X1 U29763 ( .A1(n17619), .A2(n28801), .B(n9719), .ZN(n26991) );
  INV_X4 U29764 ( .I(n26041), .ZN(n52977) );
  XOR2_X1 U29765 ( .A1(n39705), .A2(n37878), .Z(n44634) );
  XOR2_X1 U29766 ( .A1(n38277), .A2(n38651), .Z(n39705) );
  NAND2_X1 U29769 ( .A1(n11662), .A2(n31117), .ZN(n14271) );
  NOR2_X2 U29770 ( .A1(n12051), .A2(n13392), .ZN(n14276) );
  OAI21_X1 U29771 ( .A1(n39416), .A2(n39417), .B(n2234), .ZN(n21283) );
  OAI21_X1 U29772 ( .A1(n21285), .A2(n21284), .B(n21283), .ZN(n21282) );
  OR2_X1 U29774 ( .A1(n63014), .A2(n1717), .Z(n43188) );
  XOR2_X1 U29775 ( .A1(n44083), .A2(n3504), .Z(n9723) );
  INV_X4 U29777 ( .I(n15258), .ZN(n41430) );
  OR2_X1 U29779 ( .A1(n12687), .A2(n65275), .Z(n44286) );
  XOR2_X1 U29790 ( .A1(n57630), .A2(n45872), .Z(n45873) );
  INV_X1 U29799 ( .I(n6170), .ZN(n39905) );
  XOR2_X1 U29808 ( .A1(n17272), .A2(n20303), .Z(n9745) );
  XOR2_X1 U29809 ( .A1(n17237), .A2(n17273), .Z(n9746) );
  NAND3_X2 U29812 ( .A1(n24395), .A2(n24396), .A3(n20019), .ZN(n49549) );
  BUF_X2 U29816 ( .I(n15736), .Z(n9752) );
  XOR2_X1 U29820 ( .A1(n9755), .A2(n37997), .Z(n17149) );
  NAND2_X2 U29823 ( .A1(n13840), .A2(n47779), .ZN(n44558) );
  NAND3_X2 U29825 ( .A1(n13406), .A2(n13404), .A3(n13405), .ZN(n37130) );
  XOR2_X1 U29826 ( .A1(n21083), .A2(n32494), .Z(n9759) );
  OR2_X1 U29830 ( .A1(n5008), .A2(n53451), .Z(n49627) );
  NOR2_X2 U29831 ( .A1(n9616), .A2(n53726), .ZN(n53716) );
  NOR2_X1 U29832 ( .A1(n47928), .A2(n47927), .ZN(n15601) );
  INV_X2 U29833 ( .I(n9762), .ZN(n19005) );
  XOR2_X1 U29835 ( .A1(n9763), .A2(n56335), .Z(Plaintext[154]) );
  INV_X1 U29836 ( .I(n30944), .ZN(n34529) );
  NAND2_X2 U29837 ( .A1(n10486), .A2(n25549), .ZN(n20593) );
  NAND3_X1 U29838 ( .A1(n54923), .A2(n54922), .A3(n17959), .ZN(n54935) );
  XOR2_X1 U29840 ( .A1(n18091), .A2(n8065), .Z(n23841) );
  INV_X2 U29842 ( .I(n9767), .ZN(n25377) );
  NAND2_X2 U29844 ( .A1(n8758), .A2(n48584), .ZN(n48482) );
  INV_X2 U29845 ( .I(n9770), .ZN(n15759) );
  INV_X2 U29846 ( .I(n9771), .ZN(n27930) );
  XNOR2_X1 U29847 ( .A1(Ciphertext[89]), .A2(Key[132]), .ZN(n9771) );
  INV_X4 U29849 ( .I(n14930), .ZN(n23816) );
  AOI21_X1 U29852 ( .A1(n10275), .A2(n16911), .B(n17176), .ZN(n42991) );
  NAND4_X2 U29853 ( .A1(n15495), .A2(n15497), .A3(n9776), .A4(n65272), .ZN(
        n24375) );
  XOR2_X1 U29856 ( .A1(n38635), .A2(n9781), .Z(n9780) );
  NAND2_X1 U29857 ( .A1(n45896), .A2(n59216), .ZN(n45899) );
  NOR2_X2 U29862 ( .A1(n38480), .A2(n24890), .ZN(n41186) );
  NOR2_X2 U29863 ( .A1(n25866), .A2(n25867), .ZN(n10397) );
  NOR2_X2 U29864 ( .A1(n27318), .A2(n9784), .ZN(n31051) );
  XOR2_X1 U29870 ( .A1(n9791), .A2(n12206), .Z(Plaintext[6]) );
  NAND4_X2 U29872 ( .A1(n36816), .A2(n36815), .A3(n36814), .A4(n36817), .ZN(
        n37681) );
  NAND2_X2 U29879 ( .A1(n22711), .A2(n48140), .ZN(n50331) );
  XOR2_X1 U29880 ( .A1(n46386), .A2(n63745), .Z(n14349) );
  XOR2_X1 U29882 ( .A1(n43764), .A2(n46549), .Z(n26212) );
  BUF_X4 U29886 ( .I(n26667), .Z(n11987) );
  BUF_X2 U29887 ( .I(n1301), .Z(n9801) );
  AND2_X2 U29889 ( .A1(n28870), .A2(n28201), .Z(n19279) );
  AND3_X2 U29890 ( .A1(n27720), .A2(n27722), .A3(n27721), .Z(n13976) );
  XOR2_X1 U29893 ( .A1(n38869), .A2(n38868), .Z(n9803) );
  XOR2_X1 U29894 ( .A1(n9804), .A2(n14480), .Z(n20963) );
  XOR2_X1 U29895 ( .A1(n20355), .A2(n39209), .Z(n9804) );
  NAND2_X1 U29898 ( .A1(n24059), .A2(n35848), .ZN(n20257) );
  XOR2_X1 U29902 ( .A1(n11676), .A2(n11675), .Z(n9809) );
  XOR2_X1 U29904 ( .A1(n39629), .A2(n9810), .Z(n10295) );
  XOR2_X1 U29905 ( .A1(n39688), .A2(n22855), .Z(n9811) );
  AOI22_X1 U29906 ( .A1(n34966), .A2(n59293), .B1(n34976), .B2(n34977), .ZN(
        n13023) );
  OR2_X1 U29912 ( .A1(n65161), .A2(n47380), .Z(n47146) );
  NAND3_X1 U29913 ( .A1(n56287), .A2(n56288), .A3(n24120), .ZN(n56289) );
  NAND4_X2 U29914 ( .A1(n9821), .A2(n14163), .A3(n29524), .A4(n14164), .ZN(
        n15587) );
  INV_X2 U29915 ( .I(n33098), .ZN(n16856) );
  XOR2_X1 U29917 ( .A1(n9823), .A2(n20703), .Z(n11384) );
  XOR2_X1 U29918 ( .A1(n21006), .A2(n33144), .Z(n9823) );
  NAND2_X2 U29922 ( .A1(n15971), .A2(n20544), .ZN(n49803) );
  NOR2_X2 U29923 ( .A1(n9828), .A2(n39331), .ZN(n39427) );
  AND2_X1 U29925 ( .A1(n48301), .A2(n48300), .Z(n9829) );
  INV_X2 U29926 ( .I(n23297), .ZN(n27478) );
  OR2_X1 U29927 ( .A1(n17930), .A2(n11994), .Z(n15679) );
  XOR2_X1 U29928 ( .A1(n21661), .A2(n21662), .Z(n21660) );
  XOR2_X1 U29931 ( .A1(n9831), .A2(n55060), .Z(Plaintext[92]) );
  XOR2_X1 U29932 ( .A1(n9832), .A2(n45100), .Z(n21420) );
  XOR2_X1 U29933 ( .A1(n22483), .A2(n45098), .Z(n9832) );
  NOR2_X2 U29934 ( .A1(n52857), .A2(n57079), .ZN(n52668) );
  NAND2_X1 U29935 ( .A1(n35926), .A2(n9836), .ZN(n35929) );
  NOR2_X2 U29940 ( .A1(n45805), .A2(n57400), .ZN(n46816) );
  INV_X4 U29941 ( .I(n1381), .ZN(n50081) );
  AND2_X1 U29942 ( .A1(n16504), .A2(n60214), .Z(n16152) );
  INV_X2 U29948 ( .I(n26641), .ZN(n28299) );
  OAI22_X1 U29949 ( .A1(n26037), .A2(n12184), .B1(n11659), .B2(n35785), .ZN(
        n34424) );
  XOR2_X1 U29958 ( .A1(n58834), .A2(n14648), .Z(n24739) );
  NAND2_X1 U29962 ( .A1(n18842), .A2(n18840), .ZN(n30056) );
  XOR2_X1 U29966 ( .A1(n12377), .A2(n23005), .Z(n9861) );
  XOR2_X1 U29968 ( .A1(n14508), .A2(n38756), .Z(n38759) );
  NAND2_X1 U29971 ( .A1(n30766), .A2(n19525), .ZN(n14526) );
  XOR2_X1 U29973 ( .A1(n9864), .A2(n51430), .Z(n50032) );
  XOR2_X1 U29974 ( .A1(n51764), .A2(n50031), .Z(n9864) );
  NOR2_X2 U29975 ( .A1(n25866), .A2(n47682), .ZN(n47687) );
  XOR2_X1 U29976 ( .A1(n39642), .A2(n39643), .Z(n13437) );
  XOR2_X1 U29977 ( .A1(n10782), .A2(n39347), .Z(n39643) );
  XOR2_X1 U29982 ( .A1(n18114), .A2(n45399), .Z(n11201) );
  OR2_X2 U29986 ( .A1(n20716), .A2(n14876), .Z(n28375) );
  XOR2_X1 U29987 ( .A1(n31592), .A2(n1827), .Z(n26078) );
  XOR2_X1 U29988 ( .A1(n13520), .A2(n54563), .Z(n31592) );
  OR2_X1 U29989 ( .A1(n26610), .A2(n12423), .Z(n13514) );
  AOI22_X1 U29990 ( .A1(n47382), .A2(n11202), .B1(n47380), .B2(n47381), .ZN(
        n12499) );
  NOR2_X2 U29991 ( .A1(n22736), .A2(n23347), .ZN(n47380) );
  XOR2_X1 U29994 ( .A1(n8983), .A2(n16432), .Z(n9873) );
  AND2_X1 U29995 ( .A1(n35465), .A2(n58267), .Z(n15892) );
  OR2_X1 U29998 ( .A1(n55820), .A2(n21403), .Z(n55793) );
  AOI22_X1 U29999 ( .A1(n56464), .A2(n19827), .B1(n56465), .B2(n56481), .ZN(
        n56468) );
  INV_X2 U30003 ( .I(n9880), .ZN(n14039) );
  XOR2_X1 U30004 ( .A1(n17765), .A2(n17763), .Z(n9880) );
  NAND3_X1 U30007 ( .A1(n37220), .A2(n37221), .A3(n60431), .ZN(n20646) );
  OAI21_X1 U30008 ( .A1(n21852), .A2(n56368), .B(n12720), .ZN(n52283) );
  XOR2_X1 U30009 ( .A1(n14961), .A2(n9882), .Z(n14828) );
  OR2_X1 U30010 ( .A1(n49861), .A2(n8732), .Z(n14436) );
  INV_X1 U30011 ( .I(n52665), .ZN(n57058) );
  XOR2_X1 U30013 ( .A1(n16308), .A2(n30564), .Z(n44290) );
  NAND2_X1 U30015 ( .A1(n48278), .A2(n48277), .ZN(n13388) );
  NOR2_X1 U30017 ( .A1(n16811), .A2(n28549), .ZN(n16810) );
  XOR2_X1 U30021 ( .A1(n21895), .A2(n46146), .Z(n9888) );
  NAND2_X1 U30022 ( .A1(n53671), .A2(n53670), .ZN(n53684) );
  NOR2_X1 U30023 ( .A1(n9907), .A2(n23035), .ZN(n44281) );
  INV_X1 U30025 ( .I(n55285), .ZN(n15317) );
  NOR2_X2 U30031 ( .A1(n522), .A2(n26217), .ZN(n29191) );
  NAND3_X1 U30041 ( .A1(n56988), .A2(n56987), .A3(n56989), .ZN(n56995) );
  NAND2_X1 U30042 ( .A1(n49262), .A2(n49261), .ZN(n13783) );
  BUF_X4 U30043 ( .I(n41043), .Z(n41779) );
  NAND2_X1 U30045 ( .A1(n12693), .A2(n15084), .ZN(n9909) );
  NOR3_X2 U30049 ( .A1(n52047), .A2(n9913), .A3(n9912), .ZN(n21410) );
  NAND2_X1 U30052 ( .A1(n20563), .A2(n20562), .ZN(n50435) );
  XOR2_X1 U30056 ( .A1(n45845), .A2(n10253), .Z(n13299) );
  XOR2_X1 U30058 ( .A1(n14707), .A2(n38458), .Z(n9917) );
  XOR2_X1 U30059 ( .A1(n9918), .A2(n55546), .Z(Plaintext[116]) );
  NAND3_X1 U30060 ( .A1(n55544), .A2(n55543), .A3(n55545), .ZN(n9918) );
  NOR2_X1 U30062 ( .A1(n43987), .A2(n19346), .ZN(n21798) );
  AOI22_X1 U30063 ( .A1(n55812), .A2(n9920), .B1(n55760), .B2(n55820), .ZN(
        n55747) );
  INV_X1 U30064 ( .I(n55780), .ZN(n9920) );
  NOR2_X2 U30065 ( .A1(n21403), .A2(n55821), .ZN(n55780) );
  NAND4_X2 U30067 ( .A1(n32137), .A2(n32136), .A3(n32134), .A4(n32135), .ZN(
        n32141) );
  AND2_X1 U30068 ( .A1(n13187), .A2(n28265), .Z(n13203) );
  NOR4_X2 U30072 ( .A1(n55125), .A2(n55124), .A3(n55123), .A4(n55122), .ZN(
        n55128) );
  XOR2_X1 U30077 ( .A1(n21963), .A2(n21962), .Z(n52622) );
  NOR2_X1 U30078 ( .A1(n1597), .A2(n19497), .ZN(n19496) );
  XOR2_X1 U30079 ( .A1(n13581), .A2(n38977), .Z(n13580) );
  XOR2_X1 U30080 ( .A1(n62502), .A2(n37633), .Z(n38977) );
  XOR2_X1 U30081 ( .A1(n9928), .A2(n64316), .Z(n23221) );
  INV_X2 U30090 ( .I(n9936), .ZN(n26100) );
  NAND3_X2 U30092 ( .A1(n13264), .A2(n13266), .A3(n13265), .ZN(n23230) );
  OAI21_X1 U30093 ( .A1(n29675), .A2(n11948), .B(n10738), .ZN(n11947) );
  NOR2_X1 U30094 ( .A1(n11947), .A2(n11943), .ZN(n11942) );
  XOR2_X1 U30098 ( .A1(n26310), .A2(Key[143]), .Z(n9940) );
  XOR2_X1 U30100 ( .A1(n21170), .A2(n42731), .Z(n46318) );
  XOR2_X1 U30104 ( .A1(n18901), .A2(n1041), .Z(n9945) );
  AOI21_X1 U30105 ( .A1(n16787), .A2(n27460), .B(n16786), .ZN(n9946) );
  XOR2_X1 U30108 ( .A1(n9948), .A2(n10417), .Z(n25059) );
  AOI21_X1 U30110 ( .A1(n17037), .A2(n17036), .B(n54023), .ZN(n18621) );
  OR2_X1 U30116 ( .A1(n53066), .A2(n53110), .Z(n53068) );
  XOR2_X1 U30129 ( .A1(n44583), .A2(n44584), .Z(n44585) );
  NAND2_X1 U30134 ( .A1(n21930), .A2(n64608), .ZN(n21929) );
  NAND3_X1 U30138 ( .A1(n48394), .A2(n48393), .A3(n6704), .ZN(n17773) );
  OR2_X2 U30139 ( .A1(n34203), .A2(n18205), .Z(n35983) );
  NAND2_X2 U30141 ( .A1(n11558), .A2(n34921), .ZN(n35503) );
  NAND3_X1 U30142 ( .A1(n42248), .A2(n61785), .A3(n42247), .ZN(n42256) );
  XOR2_X1 U30144 ( .A1(n24064), .A2(n14565), .Z(n13748) );
  NAND3_X2 U30145 ( .A1(n30596), .A2(n20186), .A3(n30595), .ZN(n14565) );
  NOR2_X2 U30146 ( .A1(n58852), .A2(n1437), .ZN(n18810) );
  NOR2_X2 U30147 ( .A1(n18033), .A2(n18036), .ZN(n23004) );
  NOR3_X2 U30151 ( .A1(n9976), .A2(n9975), .A3(n9974), .ZN(n15886) );
  OAI21_X1 U30153 ( .A1(n40089), .A2(n9978), .B(n16118), .ZN(n39895) );
  NOR2_X1 U30154 ( .A1(n40090), .A2(n60971), .ZN(n9978) );
  OAI21_X1 U30162 ( .A1(n19789), .A2(n35663), .B(n33128), .ZN(n33129) );
  NOR2_X1 U30163 ( .A1(n33129), .A2(n9677), .ZN(n24324) );
  NOR3_X2 U30168 ( .A1(n10410), .A2(n10411), .A3(n26239), .ZN(n26667) );
  NAND2_X1 U30169 ( .A1(n54617), .A2(n20701), .ZN(n19500) );
  BUF_X2 U30172 ( .I(n36404), .Z(n9984) );
  INV_X4 U30174 ( .I(n37067), .ZN(n36691) );
  BUF_X2 U30175 ( .I(n25092), .Z(n9988) );
  XOR2_X1 U30177 ( .A1(n9989), .A2(n15865), .Z(n32052) );
  XNOR2_X1 U30180 ( .A1(n37526), .A2(n38458), .ZN(n14681) );
  XOR2_X1 U30184 ( .A1(n9991), .A2(n16128), .Z(n33628) );
  NAND3_X1 U30188 ( .A1(n26879), .A2(n26880), .A3(n28672), .ZN(n26893) );
  INV_X2 U30193 ( .I(n9995), .ZN(n26912) );
  XOR2_X1 U30200 ( .A1(n39225), .A2(n9997), .Z(n16248) );
  XOR2_X1 U30201 ( .A1(n37770), .A2(n960), .Z(n9997) );
  INV_X1 U30202 ( .I(n17994), .ZN(n13471) );
  AND2_X1 U30203 ( .A1(n53491), .A2(n17110), .Z(n53504) );
  NAND2_X1 U30204 ( .A1(n47483), .A2(n47488), .ZN(n13040) );
  NAND2_X1 U30205 ( .A1(n53398), .A2(n53397), .ZN(n13423) );
  NAND2_X2 U30210 ( .A1(n4283), .A2(n61361), .ZN(n53296) );
  INV_X2 U30212 ( .I(n23113), .ZN(n45751) );
  AND2_X1 U30213 ( .A1(n16436), .A2(n16435), .Z(n10000) );
  AND2_X1 U30218 ( .A1(n43566), .A2(n43548), .Z(n10003) );
  NOR2_X2 U30219 ( .A1(n63635), .A2(n56229), .ZN(n56424) );
  INV_X2 U30220 ( .I(n30803), .ZN(n29932) );
  XOR2_X1 U30224 ( .A1(n15677), .A2(n57321), .Z(n15675) );
  AOI22_X1 U30227 ( .A1(n9139), .A2(n26492), .B1(n20930), .B2(n1892), .ZN(
        n26495) );
  NOR2_X2 U30230 ( .A1(n28243), .A2(n27380), .ZN(n27389) );
  NOR2_X2 U30231 ( .A1(n11110), .A2(n28067), .ZN(n28243) );
  INV_X2 U30237 ( .I(n10019), .ZN(n16451) );
  XOR2_X1 U30245 ( .A1(n25741), .A2(n1314), .Z(n10024) );
  NOR2_X2 U30252 ( .A1(n10027), .A2(n53447), .ZN(n53448) );
  NOR2_X2 U30255 ( .A1(n38264), .A2(n65271), .ZN(n42508) );
  NOR2_X1 U30257 ( .A1(n56682), .A2(n56681), .ZN(n56685) );
  XOR2_X1 U30259 ( .A1(n10035), .A2(n12342), .Z(n17868) );
  XOR2_X1 U30260 ( .A1(n44104), .A2(n17869), .Z(n10035) );
  XOR2_X1 U30261 ( .A1(n52372), .A2(n15353), .Z(n10791) );
  XOR2_X1 U30263 ( .A1(n10036), .A2(n22953), .Z(n39272) );
  XOR2_X1 U30264 ( .A1(n21688), .A2(n38741), .Z(n10036) );
  NAND2_X1 U30266 ( .A1(n37182), .A2(n37183), .ZN(n34884) );
  XOR2_X1 U30275 ( .A1(n11661), .A2(n32085), .Z(n32315) );
  INV_X4 U30276 ( .I(n14705), .ZN(n23191) );
  NAND2_X1 U30278 ( .A1(n43738), .A2(n43734), .ZN(n13524) );
  INV_X4 U30281 ( .I(n10174), .ZN(n56554) );
  OR2_X1 U30282 ( .A1(n29692), .A2(n491), .Z(n17849) );
  INV_X2 U30284 ( .I(n10053), .ZN(n43750) );
  XOR2_X1 U30286 ( .A1(n39449), .A2(n10056), .Z(n16513) );
  XOR2_X1 U30287 ( .A1(n16514), .A2(n39452), .Z(n10056) );
  INV_X2 U30288 ( .I(n52044), .ZN(n55300) );
  NAND3_X1 U30289 ( .A1(n12471), .A2(n1853), .A3(n31279), .ZN(n12470) );
  XOR2_X1 U30290 ( .A1(n44038), .A2(n10058), .Z(n22433) );
  XOR2_X1 U30291 ( .A1(n44154), .A2(n60458), .Z(n10058) );
  XOR2_X1 U30293 ( .A1(n10060), .A2(n53175), .Z(Plaintext[10]) );
  XOR2_X1 U30295 ( .A1(n10618), .A2(n50568), .Z(n10062) );
  XOR2_X1 U30299 ( .A1(n10065), .A2(n51056), .Z(n13288) );
  AND2_X1 U30302 ( .A1(n19223), .A2(n27698), .Z(n12740) );
  INV_X2 U30305 ( .I(n12423), .ZN(n10946) );
  OR2_X1 U30306 ( .A1(n12423), .A2(n23191), .Z(n28361) );
  XOR2_X1 U30308 ( .A1(n39468), .A2(n39467), .Z(n10069) );
  AOI21_X1 U30312 ( .A1(n10072), .A2(n34338), .B(n34752), .ZN(n20955) );
  AND2_X1 U30315 ( .A1(n14189), .A2(n17364), .Z(n36336) );
  NOR2_X2 U30316 ( .A1(n10075), .A2(n34091), .ZN(n20280) );
  XOR2_X1 U30317 ( .A1(n46251), .A2(n56065), .Z(n10076) );
  XNOR2_X1 U30318 ( .A1(n14755), .A2(n18862), .ZN(n38828) );
  AND4_X1 U30319 ( .A1(n55208), .A2(n16978), .A3(n55222), .A4(n16943), .Z(
        n55178) );
  BUF_X2 U30325 ( .I(n22317), .Z(n10087) );
  XOR2_X1 U30328 ( .A1(n10090), .A2(n1618), .Z(n52075) );
  OAI21_X1 U30330 ( .A1(n1413), .A2(n21839), .B(n37393), .ZN(n16910) );
  NOR2_X2 U30335 ( .A1(n23773), .A2(n23800), .ZN(n15414) );
  AND2_X1 U30337 ( .A1(n43675), .A2(n5001), .Z(n22089) );
  XOR2_X1 U30339 ( .A1(n10579), .A2(n50172), .Z(n10095) );
  NAND2_X1 U30341 ( .A1(n53698), .A2(n12323), .ZN(n12322) );
  NOR3_X2 U30347 ( .A1(n48432), .A2(n23802), .A3(n24209), .ZN(n49795) );
  NOR2_X2 U30349 ( .A1(n21135), .A2(n53848), .ZN(n54312) );
  INV_X1 U30352 ( .I(n19549), .ZN(n19529) );
  NAND2_X1 U30357 ( .A1(n11701), .A2(n31100), .ZN(n10732) );
  XOR2_X1 U30359 ( .A1(n44947), .A2(n23957), .Z(n10597) );
  NAND2_X1 U30362 ( .A1(n14548), .A2(n60262), .ZN(n28790) );
  XOR2_X1 U30365 ( .A1(n10105), .A2(n52508), .Z(n52509) );
  OR2_X1 U30366 ( .A1(n29576), .A2(n29269), .Z(n28921) );
  NAND2_X1 U30369 ( .A1(n32966), .A2(n15088), .ZN(n32967) );
  INV_X1 U30370 ( .I(n42490), .ZN(n12467) );
  INV_X2 U30372 ( .I(n60009), .ZN(n30523) );
  INV_X1 U30374 ( .I(n13248), .ZN(n12783) );
  XOR2_X1 U30375 ( .A1(n13757), .A2(n56990), .Z(n22211) );
  NOR2_X2 U30376 ( .A1(n23904), .A2(n40132), .ZN(n40136) );
  INV_X1 U30382 ( .I(n36823), .ZN(n15200) );
  INV_X2 U30383 ( .I(n22594), .ZN(n25092) );
  INV_X1 U30384 ( .I(n20546), .ZN(n15648) );
  NAND2_X2 U30385 ( .A1(n14278), .A2(n23558), .ZN(n42521) );
  OAI21_X1 U30386 ( .A1(n4635), .A2(n42240), .B(n40786), .ZN(n40787) );
  OAI21_X1 U30387 ( .A1(n40787), .A2(n40788), .B(n286), .ZN(n13915) );
  XOR2_X1 U30388 ( .A1(n23719), .A2(n14666), .Z(n13353) );
  NAND4_X2 U30389 ( .A1(n10112), .A2(n47959), .A3(n47958), .A4(n47957), .ZN(
        n47963) );
  NAND2_X1 U30394 ( .A1(n48554), .A2(n48553), .ZN(n10117) );
  NAND2_X1 U30395 ( .A1(n10123), .A2(n10121), .ZN(n30792) );
  INV_X1 U30396 ( .I(n30782), .ZN(n10122) );
  BUF_X2 U30399 ( .I(n22564), .Z(n10126) );
  INV_X1 U30400 ( .I(n45590), .ZN(n25557) );
  NAND4_X2 U30406 ( .A1(n43639), .A2(n43638), .A3(n43636), .A4(n43637), .ZN(
        n46446) );
  AND2_X1 U30408 ( .A1(n21397), .A2(n48149), .Z(n10132) );
  AND2_X1 U30410 ( .A1(n20860), .A2(n29663), .Z(n10919) );
  NAND2_X2 U30416 ( .A1(n1866), .A2(n1353), .ZN(n13411) );
  XOR2_X1 U30418 ( .A1(n44432), .A2(n44433), .Z(n10141) );
  NOR2_X2 U30420 ( .A1(n31549), .A2(n31548), .ZN(n39223) );
  NAND2_X2 U30422 ( .A1(n22765), .A2(n23337), .ZN(n27717) );
  OR2_X1 U30423 ( .A1(n16788), .A2(n23474), .Z(n16071) );
  INV_X4 U30424 ( .I(n15394), .ZN(n22717) );
  XOR2_X1 U30427 ( .A1(n9397), .A2(n10145), .Z(n14432) );
  NOR2_X2 U30434 ( .A1(n20527), .A2(n42308), .ZN(n22881) );
  INV_X1 U30436 ( .I(n20375), .ZN(n14841) );
  AOI21_X1 U30437 ( .A1(n20635), .A2(n20636), .B(n14841), .ZN(n14840) );
  OAI22_X1 U30440 ( .A1(n41166), .A2(n40645), .B1(n39066), .B2(n20925), .ZN(
        n10150) );
  INV_X1 U30441 ( .I(n28870), .ZN(n20241) );
  NAND2_X1 U30443 ( .A1(n24465), .A2(n24464), .ZN(n24463) );
  NAND2_X2 U30444 ( .A1(n61747), .A2(n26213), .ZN(n36842) );
  XOR2_X1 U30445 ( .A1(n38781), .A2(n39448), .Z(n38372) );
  XOR2_X1 U30446 ( .A1(n37555), .A2(n22988), .Z(n38781) );
  AND2_X1 U30448 ( .A1(n26719), .A2(n27292), .Z(n29136) );
  INV_X1 U30453 ( .I(Key[180]), .ZN(n11268) );
  NAND2_X1 U30454 ( .A1(n28282), .A2(n28283), .ZN(n28285) );
  AOI21_X1 U30456 ( .A1(n48539), .A2(n48540), .B(n21178), .ZN(n10155) );
  NAND2_X2 U30457 ( .A1(n1422), .A2(n58748), .ZN(n36808) );
  INV_X2 U30460 ( .I(n10156), .ZN(n14705) );
  XOR2_X1 U30461 ( .A1(Key[157]), .A2(Ciphertext[24]), .Z(n10156) );
  XOR2_X1 U30463 ( .A1(n22191), .A2(n20699), .Z(n24577) );
  NOR2_X2 U30464 ( .A1(n50296), .A2(n3054), .ZN(n50056) );
  INV_X1 U30465 ( .I(n42472), .ZN(n14499) );
  NOR4_X2 U30467 ( .A1(n13124), .A2(n13125), .A3(n998), .A4(n997), .ZN(n10167)
         );
  NAND3_X1 U30470 ( .A1(n56581), .A2(n10169), .A3(n10168), .ZN(n56251) );
  NAND2_X1 U30472 ( .A1(n56248), .A2(n56587), .ZN(n10169) );
  OAI21_X1 U30473 ( .A1(n1546), .A2(n21096), .B(n10327), .ZN(n35258) );
  XOR2_X1 U30475 ( .A1(n10171), .A2(n38918), .Z(n12890) );
  XOR2_X1 U30476 ( .A1(n38919), .A2(n12891), .Z(n10171) );
  XOR2_X1 U30479 ( .A1(n17598), .A2(n51124), .Z(n51127) );
  OAI22_X1 U30484 ( .A1(n10178), .A2(n61426), .B1(n31126), .B2(n10176), .ZN(
        n31132) );
  INV_X1 U30485 ( .I(n10177), .ZN(n10176) );
  AOI21_X1 U30486 ( .A1(n31128), .A2(n31127), .B(n31129), .ZN(n10177) );
  INV_X1 U30487 ( .I(n20556), .ZN(n20389) );
  NOR2_X2 U30489 ( .A1(n35318), .A2(n35762), .ZN(n35252) );
  NAND2_X1 U30491 ( .A1(n17723), .A2(n17722), .ZN(n17721) );
  OAI21_X1 U30493 ( .A1(n43993), .A2(n21799), .B(n43992), .ZN(n43997) );
  NAND2_X1 U30495 ( .A1(n20875), .A2(n26666), .ZN(n10410) );
  OAI21_X1 U30499 ( .A1(n12321), .A2(n53689), .B(n53688), .ZN(n12320) );
  NAND2_X1 U30501 ( .A1(n12155), .A2(n12156), .ZN(n12157) );
  NAND2_X1 U30502 ( .A1(n22302), .A2(n55923), .ZN(n10185) );
  OAI21_X1 U30504 ( .A1(n53296), .A2(n53303), .B(n53301), .ZN(n53300) );
  NAND3_X1 U30506 ( .A1(n53186), .A2(n53184), .A3(n53185), .ZN(n53188) );
  XOR2_X1 U30507 ( .A1(n24053), .A2(n53958), .Z(n22911) );
  INV_X2 U30509 ( .I(n10192), .ZN(n14930) );
  XOR2_X1 U30510 ( .A1(Ciphertext[132]), .A2(Key[145]), .Z(n10192) );
  XNOR2_X1 U30511 ( .A1(n46268), .A2(n46118), .ZN(n12260) );
  CLKBUF_X2 U30520 ( .I(Key[19]), .Z(n24067) );
  AND2_X1 U30521 ( .A1(n52809), .A2(n52810), .Z(n52811) );
  INV_X2 U30523 ( .I(n10198), .ZN(n28119) );
  XNOR2_X1 U30524 ( .A1(Key[93]), .A2(Ciphertext[152]), .ZN(n10198) );
  XOR2_X1 U30527 ( .A1(n46318), .A2(n12375), .Z(n11735) );
  AND2_X1 U30535 ( .A1(n56374), .A2(n17860), .Z(n15902) );
  XOR2_X1 U30541 ( .A1(n51917), .A2(n23222), .Z(n51502) );
  XOR2_X1 U30543 ( .A1(n32317), .A2(n32483), .Z(n30848) );
  XOR2_X1 U30551 ( .A1(n20758), .A2(n43255), .Z(n23579) );
  AOI21_X2 U30552 ( .A1(n44541), .A2(n44540), .B(n44542), .ZN(n43255) );
  NOR4_X2 U30555 ( .A1(n27587), .A2(n27586), .A3(n27585), .A4(n27584), .ZN(
        n27588) );
  NOR2_X2 U30556 ( .A1(n44226), .A2(n23314), .ZN(n43709) );
  NAND2_X2 U30557 ( .A1(n13467), .A2(n13468), .ZN(n22898) );
  XOR2_X1 U30558 ( .A1(n50967), .A2(n50966), .Z(n10217) );
  OR2_X1 U30561 ( .A1(n30832), .A2(n34679), .Z(n34675) );
  NAND4_X1 U30562 ( .A1(n53715), .A2(n53717), .A3(n53716), .A4(n17286), .ZN(
        n53723) );
  OAI21_X1 U30567 ( .A1(n10224), .A2(n7558), .B(n10223), .ZN(n28017) );
  NAND2_X2 U30568 ( .A1(n2674), .A2(n21592), .ZN(n33534) );
  INV_X1 U30569 ( .I(n29258), .ZN(n13086) );
  XOR2_X1 U30570 ( .A1(n37562), .A2(n39221), .Z(n23390) );
  NAND2_X1 U30571 ( .A1(n24488), .A2(n32071), .ZN(n10227) );
  NOR2_X2 U30572 ( .A1(n24259), .A2(n56659), .ZN(n56359) );
  XOR2_X1 U30579 ( .A1(n13663), .A2(n21970), .Z(n10543) );
  AOI22_X1 U30582 ( .A1(n23025), .A2(n21082), .B1(n53456), .B2(n53590), .ZN(
        n53457) );
  NOR2_X2 U30583 ( .A1(n14603), .A2(n14604), .ZN(n27470) );
  BUF_X2 U30584 ( .I(n35152), .Z(n22617) );
  NAND2_X1 U30586 ( .A1(n10383), .A2(n56911), .ZN(n10233) );
  NOR2_X1 U30589 ( .A1(n28519), .A2(n28520), .ZN(n28521) );
  NAND2_X1 U30597 ( .A1(n45706), .A2(n48046), .ZN(n10244) );
  INV_X2 U30604 ( .I(n34524), .ZN(n25251) );
  AND2_X1 U30608 ( .A1(n13347), .A2(n13346), .Z(n12803) );
  XOR2_X1 U30611 ( .A1(n1035), .A2(n10552), .Z(n10253) );
  XOR2_X1 U30612 ( .A1(n39363), .A2(n55368), .Z(n17339) );
  XOR2_X1 U30613 ( .A1(n55624), .A2(n55139), .Z(n39363) );
  OR2_X1 U30620 ( .A1(n20734), .A2(n20975), .Z(n28395) );
  NAND2_X2 U30625 ( .A1(n28669), .A2(n28171), .ZN(n28667) );
  INV_X2 U30626 ( .I(n10265), .ZN(n19926) );
  AND3_X1 U30628 ( .A1(n51871), .A2(n21696), .A3(n51873), .Z(n24013) );
  NOR3_X1 U30630 ( .A1(n10269), .A2(n10268), .A3(n58889), .ZN(n11452) );
  NOR2_X1 U30631 ( .A1(n4760), .A2(n63686), .ZN(n10268) );
  INV_X1 U30632 ( .I(n46754), .ZN(n10269) );
  XOR2_X1 U30633 ( .A1(n33145), .A2(n10270), .Z(n15512) );
  OAI21_X2 U30634 ( .A1(n34461), .A2(n10271), .B(n576), .ZN(n37620) );
  INV_X2 U30636 ( .I(n43923), .ZN(n43538) );
  XOR2_X1 U30637 ( .A1(n10273), .A2(n52090), .Z(n19639) );
  XOR2_X1 U30639 ( .A1(n10274), .A2(n20954), .Z(n16947) );
  XOR2_X1 U30640 ( .A1(n1619), .A2(n52531), .Z(n10274) );
  XOR2_X1 U30648 ( .A1(n10278), .A2(n61071), .Z(n23131) );
  NOR2_X1 U30652 ( .A1(n20850), .A2(n1324), .ZN(n20570) );
  XOR2_X1 U30653 ( .A1(n13904), .A2(n14706), .Z(n13903) );
  XOR2_X1 U30655 ( .A1(n8179), .A2(n16969), .Z(n10283) );
  NAND2_X2 U30656 ( .A1(n10284), .A2(n21674), .ZN(n39732) );
  NAND2_X1 U30658 ( .A1(n12956), .A2(n23248), .ZN(n12789) );
  NOR2_X1 U30661 ( .A1(n21857), .A2(n24534), .ZN(n56383) );
  AND4_X1 U30664 ( .A1(n29019), .A2(n23111), .A3(n8336), .A4(n23370), .Z(
        n16110) );
  BUF_X4 U30665 ( .I(n52700), .Z(n56547) );
  XOR2_X1 U30668 ( .A1(n10293), .A2(n31502), .Z(n22250) );
  XOR2_X1 U30669 ( .A1(n30973), .A2(n11265), .Z(n10293) );
  XOR2_X1 U30672 ( .A1(n32279), .A2(n15416), .Z(n14081) );
  NOR2_X1 U30677 ( .A1(n30376), .A2(n23918), .ZN(n14764) );
  INV_X4 U30678 ( .I(n25811), .ZN(n14315) );
  AND2_X1 U30682 ( .A1(n52641), .A2(n55024), .Z(n22518) );
  XOR2_X1 U30686 ( .A1(n25314), .A2(n4278), .Z(n33266) );
  XOR2_X1 U30688 ( .A1(n10314), .A2(n4311), .Z(n17442) );
  XOR2_X1 U30694 ( .A1(n10319), .A2(n14663), .Z(n14662) );
  NAND2_X2 U30695 ( .A1(n23486), .A2(n54031), .ZN(n54032) );
  AND2_X1 U30697 ( .A1(n54349), .A2(n9613), .Z(n15945) );
  INV_X1 U30699 ( .I(n41716), .ZN(n38683) );
  XOR2_X1 U30700 ( .A1(n23481), .A2(n951), .Z(n10320) );
  OAI21_X1 U30701 ( .A1(n38494), .A2(n13138), .B(n1400), .ZN(n13137) );
  NOR2_X1 U30702 ( .A1(n31532), .A2(n31526), .ZN(n22078) );
  OR2_X1 U30703 ( .A1(n19417), .A2(n18390), .Z(n10322) );
  NAND3_X1 U30708 ( .A1(n56744), .A2(n56742), .A3(n56743), .ZN(n56746) );
  OR2_X1 U30711 ( .A1(n48089), .A2(n60651), .Z(n10329) );
  OR2_X1 U30713 ( .A1(n50237), .A2(n1632), .Z(n10334) );
  NAND2_X2 U30717 ( .A1(n47127), .A2(n48560), .ZN(n10624) );
  OR2_X1 U30720 ( .A1(n34057), .A2(n17503), .Z(n15998) );
  NAND3_X2 U30721 ( .A1(n17005), .A2(n17009), .A3(n17008), .ZN(n16838) );
  NOR2_X2 U30725 ( .A1(n25636), .A2(n55460), .ZN(n55503) );
  NAND2_X2 U30726 ( .A1(n28051), .A2(n26281), .ZN(n28044) );
  INV_X1 U30729 ( .I(n21254), .ZN(n46696) );
  XOR2_X1 U30730 ( .A1(n21254), .A2(n45355), .Z(n14747) );
  INV_X2 U30732 ( .I(n10347), .ZN(n28488) );
  XOR2_X1 U30736 ( .A1(n10348), .A2(n53531), .Z(Plaintext[29]) );
  NOR4_X2 U30737 ( .A1(n17098), .A2(n14022), .A3(n14020), .A4(n17100), .ZN(
        n10348) );
  INV_X2 U30739 ( .I(n10349), .ZN(n24885) );
  XOR2_X1 U30740 ( .A1(Ciphertext[13]), .A2(Key[176]), .Z(n10349) );
  INV_X4 U30741 ( .I(n43155), .ZN(n43161) );
  NAND2_X2 U30744 ( .A1(n21106), .A2(n60763), .ZN(n31528) );
  XOR2_X1 U30745 ( .A1(n51387), .A2(n18846), .Z(n12258) );
  INV_X4 U30746 ( .I(n48546), .ZN(n24364) );
  NAND2_X1 U30748 ( .A1(n33361), .A2(n33360), .ZN(n22724) );
  NAND2_X2 U30749 ( .A1(n49910), .A2(n14315), .ZN(n10353) );
  NOR2_X2 U30750 ( .A1(n26114), .A2(n28655), .ZN(n30748) );
  XOR2_X1 U30754 ( .A1(n17284), .A2(n10356), .Z(n22288) );
  INV_X2 U30755 ( .I(n10357), .ZN(n15824) );
  NAND2_X1 U30758 ( .A1(n24901), .A2(n24900), .ZN(n14532) );
  XOR2_X1 U30760 ( .A1(n17594), .A2(n38618), .Z(n10360) );
  INV_X2 U30761 ( .I(n10361), .ZN(n16102) );
  XOR2_X1 U30762 ( .A1(n17592), .A2(n17591), .Z(n10361) );
  INV_X2 U30764 ( .I(n21625), .ZN(n41213) );
  NAND2_X1 U30765 ( .A1(n12310), .A2(n10842), .ZN(n10841) );
  NOR2_X1 U30766 ( .A1(n10843), .A2(n10841), .ZN(n10840) );
  XOR2_X1 U30769 ( .A1(n16622), .A2(n46257), .Z(n10364) );
  INV_X2 U30770 ( .I(n25640), .ZN(n40934) );
  NAND2_X1 U30772 ( .A1(n43705), .A2(n37921), .ZN(n18553) );
  XOR2_X1 U30774 ( .A1(n33176), .A2(n10366), .Z(n30973) );
  XOR2_X1 U30775 ( .A1(n30972), .A2(n30971), .Z(n10366) );
  XOR2_X1 U30776 ( .A1(n10367), .A2(n16349), .Z(n52117) );
  NOR2_X2 U30778 ( .A1(n25922), .A2(n13797), .ZN(n13798) );
  XOR2_X1 U30780 ( .A1(n44303), .A2(n44302), .Z(n10370) );
  NOR2_X1 U30781 ( .A1(n10880), .A2(n37187), .ZN(n26221) );
  INV_X2 U30783 ( .I(n10372), .ZN(n15101) );
  XOR2_X1 U30784 ( .A1(n37266), .A2(n37265), .Z(n10372) );
  NAND2_X2 U30785 ( .A1(n10377), .A2(n10376), .ZN(n16985) );
  INV_X4 U30786 ( .I(n57015), .ZN(n57156) );
  XOR2_X1 U30788 ( .A1(n23883), .A2(n50010), .Z(n11354) );
  INV_X1 U30789 ( .I(n33782), .ZN(n35371) );
  OR2_X1 U30790 ( .A1(n36123), .A2(n33782), .Z(n15082) );
  INV_X4 U30792 ( .I(n14934), .ZN(n57015) );
  XOR2_X1 U30799 ( .A1(n10390), .A2(n24055), .Z(n43933) );
  NOR2_X2 U30800 ( .A1(n41339), .A2(n64532), .ZN(n41556) );
  XOR2_X1 U30801 ( .A1(n13748), .A2(n31365), .Z(n13747) );
  OR2_X1 U30803 ( .A1(n31105), .A2(n31097), .Z(n14334) );
  NOR2_X2 U30804 ( .A1(n56045), .A2(n56104), .ZN(n56035) );
  NAND4_X2 U30805 ( .A1(n30582), .A2(n19396), .A3(n31113), .A4(n30581), .ZN(
        n30583) );
  NOR2_X1 U30809 ( .A1(n24562), .A2(n24561), .ZN(n24560) );
  NAND2_X2 U30817 ( .A1(n31246), .A2(n58621), .ZN(n29397) );
  CLKBUF_X8 U30818 ( .I(n35030), .Z(n36959) );
  XOR2_X1 U30824 ( .A1(n10408), .A2(n31693), .Z(n33661) );
  OAI22_X2 U30826 ( .A1(n19270), .A2(n48093), .B1(n11699), .B2(n46814), .ZN(
        n48122) );
  XOR2_X1 U30828 ( .A1(n10416), .A2(n9854), .Z(n10927) );
  XOR2_X1 U30830 ( .A1(n39257), .A2(n18939), .Z(n10417) );
  NOR2_X2 U30831 ( .A1(n16750), .A2(n21029), .ZN(n30344) );
  NAND2_X1 U30832 ( .A1(n12340), .A2(n12339), .ZN(n34665) );
  XOR2_X1 U30833 ( .A1(n37970), .A2(n37969), .Z(n37971) );
  XOR2_X1 U30837 ( .A1(n16747), .A2(n49754), .Z(n15385) );
  NOR2_X2 U30842 ( .A1(n16654), .A2(n23591), .ZN(n26719) );
  NAND2_X1 U30846 ( .A1(n41093), .A2(n41894), .ZN(n10434) );
  AND2_X1 U30848 ( .A1(n42259), .A2(n25837), .Z(n16158) );
  AND2_X1 U30849 ( .A1(n57161), .A2(n57150), .Z(n10436) );
  OR2_X1 U30852 ( .A1(n43139), .A2(n43247), .Z(n23196) );
  INV_X2 U30853 ( .I(n21830), .ZN(n57124) );
  NAND2_X1 U30854 ( .A1(n20071), .A2(n17849), .ZN(n29700) );
  NAND2_X2 U30857 ( .A1(n14517), .A2(n48134), .ZN(n48468) );
  XOR2_X1 U30859 ( .A1(n10443), .A2(n46418), .Z(n10442) );
  NAND2_X1 U30860 ( .A1(n24194), .A2(n54414), .ZN(n10445) );
  OAI21_X2 U30862 ( .A1(n17343), .A2(n23829), .B(n17522), .ZN(n27324) );
  NOR2_X2 U30863 ( .A1(n20204), .A2(n48757), .ZN(n47456) );
  NAND2_X2 U30865 ( .A1(n16411), .A2(n1633), .ZN(n48923) );
  NAND2_X1 U30867 ( .A1(n40560), .A2(n12057), .ZN(n40561) );
  NAND2_X2 U30868 ( .A1(n10446), .A2(n14531), .ZN(n28920) );
  INV_X1 U30869 ( .I(n56542), .ZN(n57011) );
  OR2_X1 U30870 ( .A1(n56542), .A2(n22029), .Z(n22041) );
  XOR2_X1 U30871 ( .A1(n60931), .A2(n32158), .Z(n19800) );
  NAND2_X2 U30872 ( .A1(n15152), .A2(n60765), .ZN(n34165) );
  INV_X2 U30873 ( .I(n10453), .ZN(n16020) );
  XOR2_X1 U30874 ( .A1(n19233), .A2(n21363), .Z(n10453) );
  NAND2_X1 U30879 ( .A1(n49332), .A2(n49333), .ZN(n10454) );
  OAI21_X1 U30880 ( .A1(n56160), .A2(n56191), .B(n15663), .ZN(n24806) );
  NOR3_X1 U30881 ( .A1(n11522), .A2(n52222), .A3(n11521), .ZN(n11715) );
  AOI21_X1 U30885 ( .A1(n54970), .A2(n54292), .B(n24192), .ZN(n54295) );
  NOR2_X1 U30886 ( .A1(n26190), .A2(n43655), .ZN(n42864) );
  NAND2_X2 U30888 ( .A1(n27661), .A2(n28488), .ZN(n27664) );
  XOR2_X1 U30889 ( .A1(n23618), .A2(n46403), .Z(n45822) );
  NOR2_X2 U30898 ( .A1(n54197), .A2(n54032), .ZN(n10464) );
  NAND2_X1 U30903 ( .A1(n49218), .A2(n49217), .ZN(n13973) );
  OAI22_X1 U30908 ( .A1(n17380), .A2(n48819), .B1(n48412), .B2(n201), .ZN(
        n10469) );
  XOR2_X1 U30909 ( .A1(n10470), .A2(n52429), .Z(n20693) );
  XOR2_X1 U30910 ( .A1(n52201), .A2(n52200), .Z(n10470) );
  INV_X2 U30917 ( .I(n11202), .ZN(n21102) );
  INV_X2 U30919 ( .I(n43053), .ZN(n17950) );
  NAND2_X2 U30920 ( .A1(n11069), .A2(n11082), .ZN(n43053) );
  NOR3_X2 U30921 ( .A1(n31027), .A2(n31028), .A3(n10478), .ZN(n35092) );
  INV_X2 U30923 ( .I(n38145), .ZN(n36994) );
  NAND2_X1 U30924 ( .A1(n28816), .A2(n17824), .ZN(n10482) );
  AND2_X1 U30927 ( .A1(n34319), .A2(n23556), .Z(n15984) );
  XOR2_X1 U30930 ( .A1(n13695), .A2(n39599), .Z(n10488) );
  NOR2_X1 U30931 ( .A1(n13590), .A2(n13589), .ZN(n56783) );
  NAND2_X1 U30934 ( .A1(n29250), .A2(n58237), .ZN(n10492) );
  NOR2_X2 U30935 ( .A1(n27574), .A2(n26618), .ZN(n26665) );
  XOR2_X1 U30936 ( .A1(n26355), .A2(Key[181]), .Z(n26359) );
  OR2_X1 U30939 ( .A1(n7802), .A2(n23584), .Z(n10494) );
  NAND3_X1 U30940 ( .A1(n47852), .A2(n637), .A3(n7395), .ZN(n47675) );
  NAND2_X1 U30942 ( .A1(n10957), .A2(n10955), .ZN(n15514) );
  NAND4_X2 U30943 ( .A1(n47522), .A2(n47523), .A3(n47520), .A4(n47521), .ZN(
        n47524) );
  NAND2_X2 U30949 ( .A1(n34209), .A2(n25372), .ZN(n13081) );
  NAND2_X1 U30951 ( .A1(n13915), .A2(n24855), .ZN(n13650) );
  INV_X4 U30952 ( .I(n21400), .ZN(n24361) );
  XOR2_X1 U30953 ( .A1(n10501), .A2(n22209), .Z(n50460) );
  INV_X4 U30959 ( .I(n23816), .ZN(n12741) );
  NAND2_X1 U30960 ( .A1(n26893), .A2(n28675), .ZN(n11333) );
  NAND2_X1 U30961 ( .A1(n10505), .A2(n26427), .ZN(n26428) );
  OAI21_X1 U30962 ( .A1(n26426), .A2(n26425), .B(n27846), .ZN(n10505) );
  NAND2_X1 U30969 ( .A1(n31091), .A2(n31090), .ZN(n14420) );
  NAND2_X2 U30973 ( .A1(n16726), .A2(n33927), .ZN(n34329) );
  XOR2_X1 U30974 ( .A1(n13622), .A2(n10510), .Z(n23032) );
  NAND2_X2 U30977 ( .A1(n38550), .A2(n18496), .ZN(n37126) );
  INV_X1 U30978 ( .I(n56042), .ZN(n56064) );
  NAND2_X1 U30979 ( .A1(n56050), .A2(n56106), .ZN(n56042) );
  XOR2_X1 U30980 ( .A1(n23192), .A2(n10513), .Z(n24140) );
  XOR2_X1 U30981 ( .A1(n25415), .A2(n51995), .Z(n10513) );
  XOR2_X1 U30982 ( .A1(n11190), .A2(n11774), .Z(n11188) );
  XOR2_X1 U30993 ( .A1(n10519), .A2(n963), .Z(n11764) );
  XOR2_X1 U30996 ( .A1(n10521), .A2(n39274), .Z(n39403) );
  XOR2_X1 U30997 ( .A1(n23573), .A2(n55242), .Z(n10521) );
  NAND2_X2 U30998 ( .A1(n19329), .A2(n14630), .ZN(n47826) );
  NAND2_X1 U30999 ( .A1(n44452), .A2(n44456), .ZN(n10522) );
  INV_X2 U31002 ( .I(n47302), .ZN(n46024) );
  NOR2_X1 U31007 ( .A1(n20024), .A2(n17479), .ZN(n17478) );
  NAND3_X2 U31008 ( .A1(n24959), .A2(n24960), .A3(n55683), .ZN(n55818) );
  INV_X2 U31010 ( .I(n23475), .ZN(n54112) );
  INV_X2 U31012 ( .I(n10533), .ZN(n16616) );
  XOR2_X1 U31013 ( .A1(n16618), .A2(n44726), .Z(n10533) );
  XOR2_X1 U31015 ( .A1(n10538), .A2(n44253), .Z(n10540) );
  XOR2_X1 U31017 ( .A1(n10539), .A2(n19069), .Z(n24346) );
  XOR2_X1 U31018 ( .A1(n10540), .A2(n44260), .Z(n11649) );
  NOR2_X2 U31022 ( .A1(n55372), .A2(n15703), .ZN(n55355) );
  XOR2_X1 U31023 ( .A1(n10543), .A2(n18435), .Z(n13662) );
  XOR2_X1 U31024 ( .A1(n10545), .A2(n20916), .Z(n23124) );
  XOR2_X1 U31025 ( .A1(n14356), .A2(n23758), .Z(n10545) );
  NAND2_X2 U31027 ( .A1(n1379), .A2(n22694), .ZN(n13988) );
  XOR2_X1 U31031 ( .A1(n43796), .A2(n43794), .Z(n10555) );
  NOR2_X2 U31033 ( .A1(n13352), .A2(n34278), .ZN(n22176) );
  INV_X2 U31036 ( .I(n19910), .ZN(n55864) );
  NAND2_X2 U31037 ( .A1(n55896), .A2(n20892), .ZN(n19910) );
  NAND2_X2 U31040 ( .A1(n12158), .A2(n473), .ZN(n41126) );
  NOR2_X1 U31041 ( .A1(n27410), .A2(n1565), .ZN(n10567) );
  NOR2_X2 U31043 ( .A1(n53700), .A2(n53688), .ZN(n20381) );
  XOR2_X1 U31045 ( .A1(n14349), .A2(n46394), .Z(n14348) );
  INV_X1 U31048 ( .I(n47087), .ZN(n47091) );
  XOR2_X1 U31056 ( .A1(n18186), .A2(n51210), .Z(n10575) );
  XOR2_X1 U31059 ( .A1(n24739), .A2(n14836), .Z(n25845) );
  AND2_X1 U31062 ( .A1(n34504), .A2(n34505), .Z(n10578) );
  OAI21_X2 U31063 ( .A1(n40076), .A2(n1721), .B(n6576), .ZN(n36654) );
  INV_X4 U31067 ( .I(n36139), .ZN(n36803) );
  XOR2_X1 U31075 ( .A1(n10597), .A2(n12728), .Z(n12727) );
  XOR2_X1 U31077 ( .A1(n26022), .A2(n49879), .Z(n10595) );
  INV_X2 U31082 ( .I(n10600), .ZN(n45075) );
  OR2_X1 U31084 ( .A1(n61736), .A2(n54300), .Z(n54294) );
  AND2_X1 U31085 ( .A1(n24240), .A2(n24239), .Z(n10602) );
  XOR2_X1 U31087 ( .A1(n45365), .A2(n12714), .Z(n10606) );
  NAND2_X2 U31088 ( .A1(n56600), .A2(n24647), .ZN(n51444) );
  NAND3_X2 U31097 ( .A1(n30112), .A2(n26918), .A3(n30142), .ZN(n26919) );
  XOR2_X1 U31101 ( .A1(n12296), .A2(n25098), .Z(n10613) );
  NOR2_X2 U31103 ( .A1(n20720), .A2(n17364), .ZN(n35863) );
  NOR2_X2 U31105 ( .A1(n15498), .A2(n57075), .ZN(n57067) );
  NAND2_X1 U31106 ( .A1(n10615), .A2(n61930), .ZN(n24611) );
  NAND2_X1 U31107 ( .A1(n39932), .A2(n1403), .ZN(n10615) );
  NAND2_X1 U31111 ( .A1(n12573), .A2(n15434), .ZN(n53216) );
  NAND2_X2 U31112 ( .A1(n14667), .A2(n27246), .ZN(n14665) );
  OAI21_X1 U31115 ( .A1(n59827), .A2(n25359), .B(n56239), .ZN(n56241) );
  NAND2_X2 U31116 ( .A1(n28496), .A2(n27661), .ZN(n27668) );
  NAND2_X1 U31117 ( .A1(n31712), .A2(n31711), .ZN(n25821) );
  OAI21_X2 U31118 ( .A1(n30143), .A2(n1315), .B(n30142), .ZN(n22311) );
  NAND3_X1 U31119 ( .A1(n54903), .A2(n16016), .A3(n14635), .ZN(n54908) );
  OAI22_X1 U31121 ( .A1(n23795), .A2(n46788), .B1(n61863), .B2(n21820), .ZN(
        n46640) );
  NOR2_X2 U31123 ( .A1(n48555), .A2(n48546), .ZN(n47101) );
  OAI21_X1 U31124 ( .A1(n61704), .A2(n36510), .B(n36509), .ZN(n36513) );
  BUF_X4 U31127 ( .I(n53115), .Z(n19080) );
  AND2_X2 U31129 ( .A1(n16532), .A2(n13694), .Z(n18751) );
  NOR2_X2 U31131 ( .A1(n56962), .A2(n56953), .ZN(n56957) );
  NOR2_X2 U31135 ( .A1(n51268), .A2(n56568), .ZN(n17211) );
  INV_X2 U31136 ( .I(n25838), .ZN(n56568) );
  XOR2_X1 U31137 ( .A1(n20962), .A2(n23417), .Z(n25838) );
  AND2_X1 U31140 ( .A1(n56311), .A2(n11144), .Z(n56338) );
  NOR2_X1 U31141 ( .A1(n25717), .A2(n25720), .ZN(n25716) );
  AND2_X2 U31142 ( .A1(n24165), .A2(n24166), .Z(n52952) );
  XOR2_X1 U31145 ( .A1(n51912), .A2(n10630), .Z(n12096) );
  XOR2_X1 U31146 ( .A1(n19970), .A2(n12097), .Z(n10630) );
  OAI22_X1 U31147 ( .A1(n33347), .A2(n61523), .B1(n63624), .B2(n33559), .ZN(
        n10632) );
  OR2_X1 U31148 ( .A1(n53366), .A2(n53365), .Z(n53371) );
  INV_X4 U31151 ( .I(n11795), .ZN(n49177) );
  XOR2_X1 U31153 ( .A1(n10634), .A2(n32504), .Z(n21085) );
  AOI21_X1 U31157 ( .A1(n54415), .A2(n61829), .B(n54414), .ZN(n54422) );
  INV_X4 U31159 ( .I(n25804), .ZN(n51959) );
  OAI21_X2 U31168 ( .A1(n10643), .A2(n10642), .B(n27344), .ZN(n23015) );
  OAI21_X1 U31172 ( .A1(n28953), .A2(n14202), .B(n29561), .ZN(n27799) );
  INV_X2 U31176 ( .I(n14774), .ZN(n23469) );
  NOR2_X1 U31177 ( .A1(n14834), .A2(n14774), .ZN(n28230) );
  INV_X1 U31178 ( .I(n24858), .ZN(n32716) );
  XOR2_X1 U31180 ( .A1(n10649), .A2(n10648), .Z(n10647) );
  XOR2_X1 U31181 ( .A1(n25925), .A2(n63791), .Z(n10648) );
  XOR2_X1 U31184 ( .A1(n62923), .A2(n1755), .Z(n10654) );
  XOR2_X1 U31187 ( .A1(n10531), .A2(n32718), .Z(n25925) );
  INV_X2 U31188 ( .I(n22662), .ZN(n19511) );
  XOR2_X1 U31189 ( .A1(n10662), .A2(n45387), .Z(n10663) );
  XOR2_X1 U31190 ( .A1(n10665), .A2(n10664), .Z(n45387) );
  XOR2_X1 U31191 ( .A1(n17919), .A2(n23534), .Z(n10665) );
  INV_X2 U31193 ( .I(n24284), .ZN(n51268) );
  NAND2_X2 U31194 ( .A1(n18119), .A2(n59180), .ZN(n56290) );
  XOR2_X1 U31199 ( .A1(n10325), .A2(n33840), .Z(n10684) );
  XOR2_X1 U31200 ( .A1(n31432), .A2(n10686), .Z(n10685) );
  XOR2_X1 U31201 ( .A1(n10687), .A2(n7225), .Z(n10686) );
  XOR2_X1 U31202 ( .A1(n31430), .A2(n19800), .Z(n10687) );
  XOR2_X1 U31203 ( .A1(n10691), .A2(n10689), .Z(n10688) );
  XOR2_X1 U31204 ( .A1(n7365), .A2(n10690), .Z(n10689) );
  XOR2_X1 U31205 ( .A1(n44735), .A2(n801), .Z(n10690) );
  XOR2_X1 U31206 ( .A1(n20073), .A2(n44826), .Z(n10691) );
  OR2_X1 U31208 ( .A1(n14809), .A2(n64406), .Z(n10694) );
  XOR2_X1 U31218 ( .A1(n11501), .A2(n22979), .Z(n22256) );
  XOR2_X1 U31219 ( .A1(n1622), .A2(n7528), .Z(n51652) );
  XOR2_X1 U31221 ( .A1(n23415), .A2(n22883), .Z(n43260) );
  AND2_X1 U31222 ( .A1(n45798), .A2(n47413), .Z(n25864) );
  OR2_X1 U31224 ( .A1(n10716), .A2(n48745), .Z(n10715) );
  INV_X2 U31228 ( .I(n10719), .ZN(n25866) );
  XOR2_X1 U31232 ( .A1(n10727), .A2(n17757), .Z(n10722) );
  XOR2_X1 U31236 ( .A1(n10726), .A2(n17756), .Z(n10725) );
  XOR2_X1 U31237 ( .A1(n51959), .A2(n51958), .Z(n10726) );
  AOI22_X1 U31241 ( .A1(n28199), .A2(n29660), .B1(n28198), .B2(n29383), .ZN(
        n10738) );
  XOR2_X1 U31244 ( .A1(n45293), .A2(n10744), .Z(n10743) );
  XOR2_X1 U31245 ( .A1(n45299), .A2(n45298), .Z(n10744) );
  XOR2_X1 U31246 ( .A1(Ciphertext[102]), .A2(Key[127]), .Z(n23158) );
  NAND2_X1 U31249 ( .A1(n20978), .A2(n34627), .ZN(n10750) );
  XOR2_X1 U31251 ( .A1(n3129), .A2(n35508), .Z(n10753) );
  INV_X1 U31255 ( .I(n10754), .ZN(n29647) );
  NAND2_X1 U31256 ( .A1(n10754), .A2(n28196), .ZN(n11946) );
  NAND2_X2 U31257 ( .A1(n20241), .A2(n25222), .ZN(n10754) );
  INV_X2 U31258 ( .I(n10761), .ZN(n49606) );
  NAND2_X1 U31259 ( .A1(n47445), .A2(n10761), .ZN(n26030) );
  INV_X1 U31261 ( .I(n11088), .ZN(n10766) );
  XOR2_X1 U31265 ( .A1(n10771), .A2(n10770), .Z(n51746) );
  XOR2_X1 U31266 ( .A1(n52611), .A2(n51742), .Z(n10771) );
  NAND2_X2 U31268 ( .A1(n25866), .A2(n25867), .ZN(n47429) );
  XOR2_X1 U31269 ( .A1(n60133), .A2(n44421), .Z(n45285) );
  XOR2_X1 U31270 ( .A1(n23771), .A2(n22978), .Z(n32118) );
  XOR2_X1 U31273 ( .A1(n7619), .A2(n39344), .Z(n10782) );
  XOR2_X1 U31274 ( .A1(n10784), .A2(n10783), .Z(n51303) );
  XOR2_X1 U31275 ( .A1(n51786), .A2(n21545), .Z(n10783) );
  XOR2_X1 U31277 ( .A1(n51388), .A2(n14946), .Z(n10786) );
  XOR2_X1 U31278 ( .A1(n10792), .A2(n10791), .Z(n52380) );
  XOR2_X1 U31279 ( .A1(n52371), .A2(n15321), .Z(n10793) );
  INV_X1 U31280 ( .I(n10794), .ZN(n37356) );
  OAI21_X1 U31281 ( .A1(n36759), .A2(n10794), .B(n37117), .ZN(n36760) );
  XOR2_X1 U31282 ( .A1(n64268), .A2(n10796), .Z(n10795) );
  XOR2_X1 U31283 ( .A1(n9956), .A2(n36739), .Z(n10796) );
  NAND2_X1 U31286 ( .A1(n37920), .A2(n10806), .ZN(n43705) );
  XOR2_X1 U31287 ( .A1(n25741), .A2(n10810), .Z(n32037) );
  XOR2_X1 U31289 ( .A1(n46581), .A2(n10812), .Z(n20345) );
  XOR2_X1 U31290 ( .A1(n10536), .A2(n23687), .Z(n45377) );
  XOR2_X1 U31291 ( .A1(n19261), .A2(n10813), .Z(n39231) );
  INV_X2 U31295 ( .I(n30804), .ZN(n25448) );
  NAND2_X2 U31296 ( .A1(n31842), .A2(n22236), .ZN(n13043) );
  OAI22_X2 U31298 ( .A1(n13962), .A2(n13961), .B1(n17617), .B2(n24746), .ZN(
        n17781) );
  NOR2_X2 U31300 ( .A1(n10970), .A2(n2160), .ZN(n41969) );
  XOR2_X1 U31303 ( .A1(n10398), .A2(n51955), .Z(n51957) );
  XOR2_X1 U31304 ( .A1(n10398), .A2(n50973), .Z(n50974) );
  XOR2_X1 U31305 ( .A1(n10461), .A2(n10398), .Z(n51833) );
  XOR2_X1 U31306 ( .A1(n49231), .A2(n10398), .Z(n49241) );
  XOR2_X1 U31307 ( .A1(n50851), .A2(n10398), .Z(n51973) );
  XOR2_X1 U31309 ( .A1(n15189), .A2(n39314), .Z(n39553) );
  OAI21_X1 U31310 ( .A1(n41503), .A2(n19174), .B(n10827), .ZN(n41504) );
  AOI22_X1 U31311 ( .A1(n10828), .A2(n23954), .B1(n25619), .B2(n28887), .ZN(
        n28888) );
  AOI21_X1 U31314 ( .A1(n22527), .A2(n10829), .B(n36483), .ZN(n34487) );
  NOR2_X1 U31316 ( .A1(n30817), .A2(n10830), .ZN(n30819) );
  NAND2_X1 U31317 ( .A1(n61187), .A2(n10830), .ZN(n26508) );
  OAI21_X1 U31319 ( .A1(n29832), .A2(n30820), .B(n10830), .ZN(n28756) );
  OAI21_X1 U31320 ( .A1(n30531), .A2(n30532), .B(n10830), .ZN(n30533) );
  INV_X4 U31321 ( .I(n30799), .ZN(n10830) );
  NOR2_X1 U31322 ( .A1(n52300), .A2(n55643), .ZN(n10834) );
  NOR2_X2 U31323 ( .A1(n52298), .A2(n63520), .ZN(n55630) );
  NAND2_X2 U31324 ( .A1(n10840), .A2(n10836), .ZN(n25259) );
  INV_X2 U31330 ( .I(n10859), .ZN(n10863) );
  XOR2_X1 U31333 ( .A1(n63791), .A2(n33840), .Z(n31772) );
  NAND2_X2 U31334 ( .A1(n6606), .A2(n13768), .ZN(n35147) );
  NOR2_X1 U31335 ( .A1(n35548), .A2(n13768), .ZN(n35550) );
  NAND2_X1 U31336 ( .A1(n35966), .A2(n13768), .ZN(n21148) );
  NAND2_X1 U31337 ( .A1(n33669), .A2(n23577), .ZN(n35544) );
  AOI21_X1 U31338 ( .A1(n64024), .A2(n35357), .B(n13768), .ZN(n21695) );
  XOR2_X1 U31339 ( .A1(n2823), .A2(n37745), .Z(n37159) );
  XOR2_X1 U31340 ( .A1(n37517), .A2(n2823), .Z(n37518) );
  INV_X1 U31341 ( .I(n10865), .ZN(n42130) );
  NOR2_X2 U31342 ( .A1(n42127), .A2(n11883), .ZN(n10865) );
  INV_X4 U31344 ( .I(n40550), .ZN(n42662) );
  NOR2_X2 U31345 ( .A1(n40499), .A2(n40498), .ZN(n40550) );
  NAND2_X1 U31346 ( .A1(n10769), .A2(n10866), .ZN(n12149) );
  INV_X2 U31350 ( .I(n10868), .ZN(n15931) );
  INV_X2 U31351 ( .I(n10870), .ZN(n20547) );
  NAND2_X2 U31352 ( .A1(n20547), .A2(n19434), .ZN(n53533) );
  NAND2_X1 U31354 ( .A1(n37003), .A2(n37326), .ZN(n10880) );
  NAND2_X1 U31358 ( .A1(n10885), .A2(n34598), .ZN(n32880) );
  INV_X4 U31363 ( .I(n11035), .ZN(n50220) );
  INV_X1 U31364 ( .I(n13801), .ZN(n23445) );
  INV_X1 U31366 ( .I(n14880), .ZN(n10891) );
  NAND2_X2 U31369 ( .A1(n48770), .A2(n64764), .ZN(n49274) );
  NOR2_X2 U31371 ( .A1(n22457), .A2(n49276), .ZN(n48770) );
  NAND2_X1 U31374 ( .A1(n57032), .A2(n15435), .ZN(n16801) );
  NOR2_X2 U31375 ( .A1(n14332), .A2(n23796), .ZN(n57032) );
  XOR2_X1 U31378 ( .A1(n46630), .A2(n7811), .Z(n10902) );
  NAND4_X2 U31381 ( .A1(n13887), .A2(n18239), .A3(n59004), .A4(n10906), .ZN(
        n22846) );
  INV_X2 U31390 ( .I(n11767), .ZN(n23352) );
  INV_X2 U31394 ( .I(n23138), .ZN(n29241) );
  NAND2_X2 U31395 ( .A1(n25448), .A2(n29242), .ZN(n29238) );
  NAND2_X2 U31396 ( .A1(n1433), .A2(n30799), .ZN(n29242) );
  INV_X2 U31398 ( .I(n18295), .ZN(n18296) );
  XOR2_X1 U31399 ( .A1(n32121), .A2(n10622), .Z(n15241) );
  NAND2_X1 U31400 ( .A1(n45694), .A2(n10193), .ZN(n45695) );
  NOR2_X2 U31401 ( .A1(n23730), .A2(n60583), .ZN(n22695) );
  INV_X1 U31403 ( .I(n10938), .ZN(n53870) );
  OAI21_X1 U31404 ( .A1(n13815), .A2(n10938), .B(n54107), .ZN(n54109) );
  NAND3_X1 U31405 ( .A1(n53869), .A2(n23704), .A3(n10938), .ZN(n53873) );
  INV_X2 U31407 ( .I(n10941), .ZN(n23656) );
  NOR2_X1 U31408 ( .A1(n10941), .A2(n49307), .ZN(n49614) );
  NAND2_X1 U31409 ( .A1(n49609), .A2(n10941), .ZN(n48705) );
  NAND4_X1 U31413 ( .A1(n42563), .A2(n42562), .A3(n42564), .A4(n60079), .ZN(
        n42569) );
  OAI22_X1 U31414 ( .A1(n22269), .A2(n42889), .B1(n43170), .B2(n60079), .ZN(
        n42908) );
  AOI21_X1 U31416 ( .A1(n28370), .A2(n10946), .B(n28369), .ZN(n28371) );
  NAND3_X2 U31418 ( .A1(n18227), .A2(n11627), .A3(n47407), .ZN(n47406) );
  OR2_X1 U31419 ( .A1(n52121), .A2(n10949), .Z(n20017) );
  NOR2_X2 U31421 ( .A1(n53795), .A2(n53823), .ZN(n53800) );
  XOR2_X1 U31422 ( .A1(n10950), .A2(n32494), .Z(n31288) );
  XOR2_X1 U31423 ( .A1(n7522), .A2(n756), .Z(n10950) );
  XOR2_X1 U31425 ( .A1(n10953), .A2(n50908), .Z(n10952) );
  NAND2_X1 U31427 ( .A1(n40997), .A2(n10954), .ZN(n10957) );
  NAND2_X2 U31431 ( .A1(n41350), .A2(n60583), .ZN(n43068) );
  NAND2_X1 U31434 ( .A1(n64036), .A2(n46771), .ZN(n10977) );
  MUX2_X1 U31438 ( .I0(n45631), .I1(n45632), .S(n47295), .Z(n45650) );
  XOR2_X1 U31439 ( .A1(n10985), .A2(n10984), .Z(n11673) );
  XOR2_X1 U31440 ( .A1(n25208), .A2(n45843), .Z(n10984) );
  XOR2_X1 U31441 ( .A1(n45047), .A2(n19727), .Z(n25208) );
  NAND2_X1 U31444 ( .A1(n10986), .A2(n64100), .ZN(n31607) );
  OAI21_X1 U31445 ( .A1(n10986), .A2(n23351), .B(n34155), .ZN(n33680) );
  XOR2_X1 U31447 ( .A1(n10620), .A2(n46619), .Z(n46622) );
  XOR2_X1 U31448 ( .A1(n10620), .A2(n44516), .Z(n44517) );
  XOR2_X1 U31452 ( .A1(n23495), .A2(n58084), .Z(n11755) );
  XOR2_X1 U31453 ( .A1(n10993), .A2(n52609), .Z(n10997) );
  INV_X2 U31454 ( .I(n26029), .ZN(n52609) );
  XOR2_X1 U31455 ( .A1(n26028), .A2(n52453), .Z(n26029) );
  INV_X2 U31456 ( .I(n41806), .ZN(n42448) );
  INV_X1 U31457 ( .I(n8805), .ZN(n52031) );
  XOR2_X1 U31459 ( .A1(n8805), .A2(n1116), .Z(n52146) );
  XOR2_X1 U31461 ( .A1(n51930), .A2(n10997), .Z(n10996) );
  INV_X2 U31463 ( .I(n43205), .ZN(n10998) );
  NAND2_X1 U31465 ( .A1(n1517), .A2(n21207), .ZN(n42434) );
  NOR2_X1 U31466 ( .A1(n10554), .A2(n65128), .ZN(n10999) );
  NOR2_X2 U31467 ( .A1(n18817), .A2(n48906), .ZN(n16571) );
  INV_X1 U31468 ( .I(n11006), .ZN(n36824) );
  NOR2_X1 U31469 ( .A1(n11009), .A2(n11008), .ZN(n11007) );
  INV_X1 U31470 ( .I(n36829), .ZN(n11009) );
  XOR2_X1 U31472 ( .A1(n37842), .A2(n15446), .Z(n11013) );
  XOR2_X1 U31473 ( .A1(n23552), .A2(n50637), .Z(n50638) );
  XOR2_X1 U31474 ( .A1(n46343), .A2(n25518), .Z(n46135) );
  XOR2_X1 U31475 ( .A1(n20044), .A2(n46136), .Z(n11014) );
  NAND2_X1 U31476 ( .A1(n18441), .A2(n7501), .ZN(n11017) );
  INV_X4 U31483 ( .I(n35605), .ZN(n36262) );
  NAND2_X1 U31487 ( .A1(n11036), .A2(n14931), .ZN(n12472) );
  AOI21_X1 U31495 ( .A1(n53197), .A2(n53605), .B(n11041), .ZN(n53200) );
  AOI21_X1 U31496 ( .A1(n53388), .A2(n11041), .B(n53387), .ZN(n53389) );
  NOR2_X1 U31498 ( .A1(n61159), .A2(n63303), .ZN(n11043) );
  NAND3_X1 U31500 ( .A1(n21207), .A2(n42432), .A3(n10554), .ZN(n11046) );
  OR2_X1 U31501 ( .A1(n34886), .A2(n36247), .Z(n11049) );
  NAND2_X2 U31502 ( .A1(n33353), .A2(n33352), .ZN(n35605) );
  XOR2_X1 U31503 ( .A1(n32486), .A2(n32485), .Z(n32487) );
  XOR2_X1 U31505 ( .A1(n57313), .A2(n39732), .Z(n21688) );
  XOR2_X1 U31509 ( .A1(Ciphertext[190]), .A2(Key[167]), .Z(n27160) );
  XOR2_X1 U31512 ( .A1(n50717), .A2(n15066), .Z(n50833) );
  NAND2_X2 U31513 ( .A1(n10820), .A2(n61187), .ZN(n29239) );
  NAND2_X1 U31518 ( .A1(n11073), .A2(n19122), .ZN(n18916) );
  NAND2_X1 U31519 ( .A1(n11073), .A2(n57412), .ZN(n26604) );
  XOR2_X1 U31520 ( .A1(n46598), .A2(n62569), .Z(n46599) );
  NAND3_X1 U31521 ( .A1(n36587), .A2(n11077), .A3(n36588), .ZN(n36592) );
  NAND3_X2 U31526 ( .A1(n11095), .A2(n11094), .A3(n11093), .ZN(n30413) );
  INV_X2 U31528 ( .I(n12546), .ZN(n13413) );
  INV_X2 U31529 ( .I(n11098), .ZN(n18452) );
  NOR2_X1 U31534 ( .A1(n28240), .A2(n4443), .ZN(n28242) );
  AOI22_X1 U31536 ( .A1(n26267), .A2(n22094), .B1(n28241), .B2(n4443), .ZN(
        n26269) );
  INV_X2 U31539 ( .I(n11119), .ZN(n11121) );
  NOR2_X2 U31540 ( .A1(n55934), .A2(n25168), .ZN(n11989) );
  NOR4_X2 U31542 ( .A1(n11139), .A2(n14797), .A3(n11135), .A4(n11133), .ZN(
        n14796) );
  NAND2_X1 U31543 ( .A1(n28238), .A2(n28241), .ZN(n11138) );
  XOR2_X1 U31546 ( .A1(n19687), .A2(n37650), .Z(n11147) );
  OR2_X1 U31552 ( .A1(n5463), .A2(n49671), .Z(n11154) );
  NOR3_X2 U31555 ( .A1(n29301), .A2(n29300), .A3(n11162), .ZN(n11161) );
  NAND2_X1 U31556 ( .A1(n1285), .A2(n55690), .ZN(n55487) );
  INV_X2 U31557 ( .I(n5531), .ZN(n37532) );
  XOR2_X1 U31558 ( .A1(n11165), .A2(n50066), .Z(n50967) );
  NOR3_X2 U31562 ( .A1(n23580), .A2(n11175), .A3(n11174), .ZN(n32317) );
  OAI22_X1 U31564 ( .A1(n37281), .A2(n37272), .B1(n37134), .B2(n11178), .ZN(
        n37140) );
  XOR2_X1 U31570 ( .A1(n12097), .A2(n52630), .Z(n20577) );
  XOR2_X1 U31571 ( .A1(n51136), .A2(n12097), .Z(n22981) );
  XOR2_X1 U31572 ( .A1(n50352), .A2(n12097), .Z(n25434) );
  XOR2_X1 U31576 ( .A1(n11201), .A2(n23559), .Z(n11200) );
  INV_X4 U31577 ( .I(n18098), .ZN(n18114) );
  NOR2_X1 U31578 ( .A1(n46747), .A2(n11202), .ZN(n46748) );
  AOI21_X2 U31579 ( .A1(n26031), .A2(n26030), .B(n11820), .ZN(n11594) );
  NAND2_X2 U31582 ( .A1(n40541), .A2(n40641), .ZN(n39069) );
  XOR2_X1 U31584 ( .A1(n38071), .A2(n38973), .Z(n11211) );
  INV_X2 U31586 ( .I(n11213), .ZN(n22363) );
  NAND2_X1 U31588 ( .A1(n11225), .A2(n64445), .ZN(n11772) );
  AOI21_X1 U31590 ( .A1(n11225), .A2(n27623), .B(n27622), .ZN(n27624) );
  OAI22_X1 U31591 ( .A1(n28402), .A2(n28416), .B1(n28401), .B2(n11226), .ZN(
        n28403) );
  XNOR2_X1 U31592 ( .A1(n11382), .A2(n11232), .ZN(n11230) );
  XOR2_X1 U31594 ( .A1(n21522), .A2(n23260), .Z(n33032) );
  XOR2_X1 U31596 ( .A1(n11240), .A2(n18797), .Z(n15446) );
  XOR2_X1 U31597 ( .A1(n11239), .A2(n37645), .Z(n11240) );
  INV_X2 U31598 ( .I(n11241), .ZN(n24259) );
  AOI22_X1 U31599 ( .A1(n61547), .A2(n7345), .B1(n10503), .B2(n35252), .ZN(
        n34439) );
  NOR2_X1 U31602 ( .A1(n11246), .A2(n48688), .ZN(n48689) );
  NOR2_X1 U31603 ( .A1(n48685), .A2(n11246), .ZN(n46974) );
  OAI21_X1 U31604 ( .A1(n34539), .A2(n34534), .B(n11247), .ZN(n32918) );
  NAND2_X1 U31605 ( .A1(n34526), .A2(n11247), .ZN(n32915) );
  XOR2_X1 U31608 ( .A1(n11255), .A2(n22530), .Z(n11254) );
  NAND2_X1 U31611 ( .A1(n12423), .A2(n64174), .ZN(n26320) );
  NOR3_X2 U31612 ( .A1(n21958), .A2(n15633), .A3(n11260), .ZN(n42583) );
  XOR2_X1 U31613 ( .A1(n11261), .A2(n32248), .Z(n32261) );
  NOR3_X1 U31614 ( .A1(n11263), .A2(n9904), .A3(n31129), .ZN(n29433) );
  NOR2_X1 U31615 ( .A1(n11262), .A2(n29566), .ZN(n16140) );
  NAND3_X1 U31616 ( .A1(n27151), .A2(n24000), .A3(n11263), .ZN(n27152) );
  MUX2_X1 U31617 ( .I0(n29909), .I1(n29916), .S(n11263), .Z(n29437) );
  XOR2_X1 U31618 ( .A1(n11265), .A2(n33177), .Z(n32408) );
  NOR2_X1 U31621 ( .A1(n22110), .A2(n26606), .ZN(n11267) );
  XOR2_X1 U31623 ( .A1(n11268), .A2(Ciphertext[41]), .Z(n28328) );
  XOR2_X1 U31624 ( .A1(n11269), .A2(n51769), .Z(n51770) );
  XOR2_X1 U31626 ( .A1(n23069), .A2(n11269), .Z(n48725) );
  XOR2_X1 U31627 ( .A1(n22790), .A2(n11269), .Z(n52085) );
  NAND2_X2 U31628 ( .A1(n18174), .A2(n5172), .ZN(n56176) );
  AND2_X1 U31629 ( .A1(n11275), .A2(n7138), .Z(n11276) );
  MUX2_X1 U31630 ( .I0(n54355), .I1(n54379), .S(n54391), .Z(n54358) );
  AOI21_X2 U31632 ( .A1(n47383), .A2(n25346), .B(n25345), .ZN(n25320) );
  NOR2_X1 U31634 ( .A1(n18228), .A2(n24179), .ZN(n11280) );
  NOR2_X2 U31635 ( .A1(n16378), .A2(n19454), .ZN(n43277) );
  XOR2_X1 U31638 ( .A1(n11285), .A2(n11283), .Z(n11287) );
  XOR2_X1 U31639 ( .A1(n11284), .A2(n11788), .Z(n11283) );
  XOR2_X1 U31640 ( .A1(n17216), .A2(n11286), .Z(n11285) );
  XOR2_X1 U31641 ( .A1(n44273), .A2(n19215), .Z(n11286) );
  INV_X2 U31642 ( .I(n11287), .ZN(n45484) );
  INV_X2 U31643 ( .I(n45484), .ZN(n16493) );
  XOR2_X1 U31646 ( .A1(n49623), .A2(n19029), .Z(n49624) );
  NAND2_X1 U31647 ( .A1(n47510), .A2(n10333), .ZN(n11297) );
  XOR2_X1 U31648 ( .A1(n11305), .A2(n16205), .Z(n22307) );
  XOR2_X1 U31651 ( .A1(Key[103]), .A2(Ciphertext[126]), .Z(n24197) );
  INV_X2 U31652 ( .I(n24197), .ZN(n28187) );
  XOR2_X1 U31654 ( .A1(n7999), .A2(n46136), .Z(n11309) );
  INV_X1 U31655 ( .I(n17238), .ZN(n14161) );
  XOR2_X1 U31656 ( .A1(n17238), .A2(n11309), .Z(n18067) );
  NAND2_X1 U31657 ( .A1(n7086), .A2(n11314), .ZN(n12673) );
  XOR2_X1 U31659 ( .A1(n11318), .A2(n12716), .Z(n14089) );
  INV_X1 U31660 ( .I(n33051), .ZN(n26165) );
  XOR2_X1 U31661 ( .A1(n23371), .A2(n15460), .Z(n51846) );
  XOR2_X1 U31664 ( .A1(n51502), .A2(n25814), .Z(n11323) );
  INV_X2 U31666 ( .I(n11557), .ZN(n54424) );
  NAND3_X1 U31668 ( .A1(n56806), .A2(n60851), .A3(n56808), .ZN(n11328) );
  XOR2_X1 U31670 ( .A1(Ciphertext[127]), .A2(Key[14]), .Z(n20786) );
  NOR2_X2 U31672 ( .A1(n31040), .A2(n31038), .ZN(n30705) );
  INV_X2 U31675 ( .I(n30148), .ZN(n31040) );
  NAND2_X2 U31678 ( .A1(n7213), .A2(n12469), .ZN(n56360) );
  INV_X2 U31683 ( .I(n23581), .ZN(n49005) );
  INV_X2 U31684 ( .I(n57031), .ZN(n57019) );
  NOR2_X2 U31686 ( .A1(n17274), .A2(n20473), .ZN(n28188) );
  NAND2_X2 U31687 ( .A1(n47970), .A2(n8044), .ZN(n12595) );
  NAND3_X1 U31690 ( .A1(n11356), .A2(n47621), .A3(n1069), .ZN(n11553) );
  OAI21_X1 U31691 ( .A1(n22468), .A2(n45576), .B(n22239), .ZN(n11356) );
  XOR2_X1 U31693 ( .A1(n11358), .A2(n46159), .Z(n11357) );
  XOR2_X1 U31694 ( .A1(n718), .A2(n32614), .Z(n32616) );
  XOR2_X1 U31697 ( .A1(n10619), .A2(n43904), .Z(n43905) );
  XOR2_X1 U31698 ( .A1(n23905), .A2(n10619), .Z(n44722) );
  XOR2_X1 U31699 ( .A1(n23906), .A2(n10619), .Z(n46296) );
  NOR2_X1 U31702 ( .A1(n31247), .A2(n23008), .ZN(n11378) );
  XOR2_X1 U31706 ( .A1(n11384), .A2(n33059), .Z(n11383) );
  OAI21_X1 U31707 ( .A1(n54380), .A2(n54424), .B(n5324), .ZN(n54394) );
  NOR2_X2 U31717 ( .A1(n52828), .A2(n25936), .ZN(n15435) );
  NAND2_X2 U31718 ( .A1(n23796), .A2(n14332), .ZN(n57026) );
  INV_X2 U31719 ( .I(n47036), .ZN(n45538) );
  INV_X2 U31721 ( .I(n25897), .ZN(n11417) );
  XOR2_X1 U31722 ( .A1(n11419), .A2(n11418), .Z(n25298) );
  XOR2_X1 U31723 ( .A1(n25062), .A2(n14806), .Z(n11418) );
  XOR2_X1 U31724 ( .A1(n61410), .A2(n18986), .Z(n25062) );
  XOR2_X1 U31726 ( .A1(n1198), .A2(n1009), .Z(n11420) );
  OAI22_X1 U31730 ( .A1(n19027), .A2(n30455), .B1(n30457), .B2(n30456), .ZN(
        n15387) );
  AOI21_X1 U31731 ( .A1(n56285), .A2(n11427), .B(n14383), .ZN(n56287) );
  NOR2_X1 U31732 ( .A1(n11654), .A2(n23318), .ZN(n11427) );
  AND2_X1 U31734 ( .A1(n15099), .A2(n34583), .Z(n11435) );
  NOR2_X2 U31738 ( .A1(n25066), .A2(n45781), .ZN(n45529) );
  NAND2_X2 U31739 ( .A1(n11443), .A2(n47034), .ZN(n45781) );
  NOR2_X2 U31740 ( .A1(n45532), .A2(n1294), .ZN(n45785) );
  OR2_X1 U31741 ( .A1(n33493), .A2(n11445), .Z(n12239) );
  NAND3_X1 U31742 ( .A1(n1781), .A2(n1786), .A3(n12652), .ZN(n36281) );
  XOR2_X1 U31743 ( .A1(n51013), .A2(n11447), .Z(n24849) );
  INV_X2 U31748 ( .I(n25984), .ZN(n38870) );
  XOR2_X1 U31749 ( .A1(n38979), .A2(n38671), .Z(n24409) );
  XOR2_X1 U31750 ( .A1(n25984), .A2(n916), .Z(n38979) );
  XOR2_X1 U31751 ( .A1(n38168), .A2(n16120), .Z(n25984) );
  NOR2_X1 U31753 ( .A1(n41583), .A2(n59309), .ZN(n12932) );
  XOR2_X1 U31757 ( .A1(n32284), .A2(n32291), .Z(n11457) );
  INV_X2 U31758 ( .I(n47181), .ZN(n48622) );
  NAND2_X2 U31762 ( .A1(n8891), .A2(n1351), .ZN(n30519) );
  OR2_X1 U31763 ( .A1(n47983), .A2(n22085), .Z(n11467) );
  NAND2_X2 U31764 ( .A1(n47982), .A2(n11468), .ZN(n47983) );
  XOR2_X1 U31766 ( .A1(n11471), .A2(n51582), .Z(n11470) );
  NOR2_X1 U31772 ( .A1(n43087), .A2(n11476), .ZN(n43088) );
  NAND2_X1 U31773 ( .A1(n11477), .A2(n24077), .ZN(n33427) );
  INV_X4 U31774 ( .I(n22940), .ZN(n52154) );
  XOR2_X1 U31776 ( .A1(n11479), .A2(n15149), .Z(n11478) );
  XOR2_X1 U31778 ( .A1(n11486), .A2(n31485), .Z(n11483) );
  XOR2_X1 U31780 ( .A1(n11486), .A2(n15510), .Z(n32293) );
  XOR2_X1 U31782 ( .A1(n11488), .A2(n15736), .Z(n20972) );
  OAI21_X1 U31783 ( .A1(n11492), .A2(n45201), .B(n47803), .ZN(n44001) );
  NAND2_X1 U31784 ( .A1(n47800), .A2(n11492), .ZN(n47695) );
  NOR2_X2 U31785 ( .A1(n47797), .A2(n25895), .ZN(n11492) );
  AOI21_X2 U31787 ( .A1(n42684), .A2(n42683), .B(n42682), .ZN(n44540) );
  NAND2_X2 U31789 ( .A1(n23986), .A2(n40943), .ZN(n39104) );
  AND2_X1 U31791 ( .A1(n30471), .A2(n30472), .Z(n11495) );
  XOR2_X1 U31793 ( .A1(n11500), .A2(n25273), .Z(n11499) );
  INV_X2 U31794 ( .I(n38759), .ZN(n41469) );
  AND2_X1 U31796 ( .A1(n40756), .A2(n18623), .Z(n11505) );
  OR2_X2 U31797 ( .A1(n38759), .A2(n14994), .Z(n18623) );
  XOR2_X1 U31799 ( .A1(n13079), .A2(n11617), .Z(n17103) );
  INV_X2 U31800 ( .I(n26161), .ZN(n11617) );
  XOR2_X1 U31801 ( .A1(Ciphertext[66]), .A2(Key[67]), .Z(n26161) );
  NOR4_X2 U31802 ( .A1(n11517), .A2(n42375), .A3(n42374), .A4(n43450), .ZN(
        n11516) );
  XOR2_X1 U31804 ( .A1(n11519), .A2(n46311), .Z(n45218) );
  NAND2_X2 U31807 ( .A1(n22422), .A2(n15535), .ZN(n15533) );
  NAND2_X1 U31810 ( .A1(n11524), .A2(n11523), .ZN(n11522) );
  OAI22_X1 U31811 ( .A1(n27889), .A2(n27890), .B1(n27888), .B2(n1889), .ZN(
        n27895) );
  XOR2_X1 U31812 ( .A1(n11527), .A2(n17320), .Z(n14819) );
  XOR2_X1 U31813 ( .A1(n11528), .A2(n5727), .Z(n19757) );
  XOR2_X1 U31818 ( .A1(n11534), .A2(n60141), .Z(n39267) );
  INV_X2 U31823 ( .I(n36453), .ZN(n36444) );
  XOR2_X1 U31825 ( .A1(n63011), .A2(n11546), .Z(n11545) );
  XOR2_X1 U31826 ( .A1(n10992), .A2(n817), .Z(n11546) );
  XOR2_X1 U31827 ( .A1(n39543), .A2(n18354), .Z(n18355) );
  XOR2_X1 U31828 ( .A1(n51284), .A2(n1618), .Z(n51761) );
  XOR2_X1 U31830 ( .A1(n61462), .A2(n11529), .Z(n11551) );
  NAND3_X1 U31831 ( .A1(n42404), .A2(n25534), .A3(n19241), .ZN(n42406) );
  NAND4_X2 U31832 ( .A1(n11553), .A2(n47628), .A3(n47626), .A4(n47627), .ZN(
        n11552) );
  XOR2_X1 U31836 ( .A1(n1558), .A2(n30455), .Z(n11569) );
  OAI21_X1 U31838 ( .A1(n11571), .A2(n1457), .B(n53184), .ZN(n50476) );
  NOR2_X2 U31840 ( .A1(n20349), .A2(n19567), .ZN(n11571) );
  AOI21_X2 U31841 ( .A1(n28266), .A2(n28265), .B(n11572), .ZN(n18389) );
  XOR2_X1 U31844 ( .A1(n61960), .A2(n24449), .Z(n11575) );
  INV_X2 U31846 ( .I(n11589), .ZN(n26791) );
  XNOR2_X1 U31847 ( .A1(Ciphertext[116]), .A2(Key[33]), .ZN(n11589) );
  XOR2_X1 U31850 ( .A1(n10536), .A2(n44016), .Z(n44017) );
  NAND2_X2 U31852 ( .A1(n34566), .A2(n32295), .ZN(n34956) );
  INV_X2 U31853 ( .I(n21725), .ZN(n34566) );
  NAND2_X1 U31855 ( .A1(n11599), .A2(n18227), .ZN(n43829) );
  NAND3_X1 U31856 ( .A1(n18265), .A2(n47671), .A3(n11599), .ZN(n18264) );
  NOR2_X1 U31857 ( .A1(n47870), .A2(n11599), .ZN(n12738) );
  NOR2_X1 U31861 ( .A1(n29172), .A2(n62005), .ZN(n15196) );
  NAND2_X2 U31862 ( .A1(n13079), .A2(n11514), .ZN(n13763) );
  XOR2_X1 U31864 ( .A1(n18490), .A2(n11610), .Z(n32278) );
  XOR2_X1 U31865 ( .A1(n57167), .A2(n11529), .Z(n11610) );
  XOR2_X1 U31866 ( .A1(Ciphertext[69]), .A2(Key[184]), .Z(n11616) );
  INV_X2 U31868 ( .I(n11616), .ZN(n13079) );
  INV_X1 U31873 ( .I(n11557), .ZN(n11622) );
  NAND2_X1 U31874 ( .A1(n11623), .A2(n61624), .ZN(n49946) );
  INV_X2 U31877 ( .I(n14038), .ZN(n14037) );
  XOR2_X1 U31878 ( .A1(n33838), .A2(n13365), .Z(n31796) );
  INV_X2 U31879 ( .I(n15413), .ZN(n13365) );
  XOR2_X1 U31880 ( .A1(n11634), .A2(n11633), .Z(n11632) );
  NAND2_X1 U31882 ( .A1(n43654), .A2(n11635), .ZN(n43661) );
  XOR2_X1 U31884 ( .A1(n11142), .A2(n60141), .Z(n39765) );
  XOR2_X1 U31885 ( .A1(n11636), .A2(n37812), .Z(n39450) );
  XOR2_X1 U31886 ( .A1(n36933), .A2(n60141), .Z(n36935) );
  XOR2_X1 U31890 ( .A1(n62477), .A2(n796), .Z(n45821) );
  NAND2_X1 U31894 ( .A1(n34001), .A2(n11643), .ZN(n16991) );
  INV_X2 U31896 ( .I(n11644), .ZN(n41856) );
  XOR2_X1 U31901 ( .A1(n30985), .A2(n23253), .Z(n32336) );
  XOR2_X1 U31902 ( .A1(n30985), .A2(n30933), .Z(n32517) );
  XOR2_X1 U31905 ( .A1(n63010), .A2(n51755), .Z(n51756) );
  NAND2_X2 U31908 ( .A1(n31121), .A2(n10235), .ZN(n32001) );
  NAND2_X1 U31910 ( .A1(n42339), .A2(n1391), .ZN(n41655) );
  OAI21_X1 U31911 ( .A1(n11654), .A2(n56350), .B(n56349), .ZN(n56356) );
  NAND2_X2 U31914 ( .A1(n1816), .A2(n24331), .ZN(n35770) );
  XOR2_X1 U31916 ( .A1(n14666), .A2(n25331), .Z(n11661) );
  XOR2_X1 U31918 ( .A1(n10292), .A2(n13830), .Z(n13949) );
  XOR2_X1 U31920 ( .A1(n59163), .A2(n32128), .Z(n11663) );
  INV_X2 U31923 ( .I(n11673), .ZN(n15823) );
  INV_X4 U31924 ( .I(n55820), .ZN(n55829) );
  MUX2_X1 U31925 ( .I0(n58018), .I1(n3686), .S(n2955), .Z(n11693) );
  XOR2_X1 U31927 ( .A1(n20408), .A2(n788), .Z(n39472) );
  NOR2_X2 U31928 ( .A1(n1868), .A2(n31105), .ZN(n31119) );
  NAND2_X2 U31929 ( .A1(n11702), .A2(n28180), .ZN(n31105) );
  NAND2_X1 U31931 ( .A1(n11704), .A2(n64450), .ZN(n39948) );
  NAND2_X1 U31932 ( .A1(n11704), .A2(n60693), .ZN(n12693) );
  NAND2_X1 U31934 ( .A1(n1468), .A2(n11705), .ZN(n49078) );
  NOR2_X2 U31935 ( .A1(n48082), .A2(n48076), .ZN(n48561) );
  NAND2_X2 U31942 ( .A1(n11726), .A2(n23554), .ZN(n55351) );
  NOR2_X2 U31943 ( .A1(n55362), .A2(n24063), .ZN(n11726) );
  XOR2_X1 U31946 ( .A1(n32228), .A2(n11732), .Z(n18732) );
  XOR2_X1 U31947 ( .A1(n32227), .A2(n1833), .Z(n11732) );
  XOR2_X1 U31949 ( .A1(n11515), .A2(n45856), .Z(n45857) );
  XOR2_X1 U31950 ( .A1(n11515), .A2(n799), .Z(n15054) );
  XOR2_X1 U31952 ( .A1(n46209), .A2(n17902), .Z(n18890) );
  INV_X1 U31954 ( .I(n11741), .ZN(n50734) );
  XOR2_X1 U31955 ( .A1(n11741), .A2(n50741), .Z(n50742) );
  XOR2_X1 U31956 ( .A1(n16984), .A2(n11741), .Z(n51231) );
  XOR2_X1 U31957 ( .A1(n11741), .A2(n21425), .Z(n50626) );
  MUX2_X1 U31959 ( .I0(n11743), .I1(n48225), .S(n62308), .Z(n48226) );
  INV_X2 U31961 ( .I(n47541), .ZN(n25481) );
  AND2_X1 U31962 ( .A1(n37087), .A2(n37940), .Z(n11754) );
  NAND2_X1 U31963 ( .A1(n27433), .A2(n18747), .ZN(n11761) );
  INV_X2 U31964 ( .I(n34614), .ZN(n34039) );
  NAND2_X2 U31965 ( .A1(n19291), .A2(n39904), .ZN(n11765) );
  INV_X2 U31966 ( .I(n11764), .ZN(n39904) );
  XOR2_X1 U31968 ( .A1(n11768), .A2(n19688), .Z(n51068) );
  XOR2_X1 U31969 ( .A1(n11768), .A2(n21994), .Z(n21993) );
  INV_X1 U31970 ( .I(n27429), .ZN(n11773) );
  XOR2_X1 U31971 ( .A1(n12056), .A2(n11775), .Z(n11774) );
  XOR2_X1 U31972 ( .A1(n25911), .A2(n11776), .Z(n11775) );
  INV_X1 U31973 ( .I(n38447), .ZN(n11776) );
  INV_X1 U31974 ( .I(n11781), .ZN(n13319) );
  NAND2_X1 U31975 ( .A1(n11781), .A2(n58975), .ZN(n14207) );
  NOR2_X1 U31976 ( .A1(n49196), .A2(n11781), .ZN(n49200) );
  AND2_X1 U31978 ( .A1(n55888), .A2(n11784), .Z(n11783) );
  OR2_X1 U31979 ( .A1(n55867), .A2(n60092), .Z(n11784) );
  OR2_X1 U31980 ( .A1(n19075), .A2(n55834), .Z(n11785) );
  XOR2_X1 U31984 ( .A1(n9628), .A2(n44321), .Z(n11788) );
  NAND2_X2 U31985 ( .A1(n13860), .A2(n13859), .ZN(n55892) );
  XOR2_X1 U31990 ( .A1(n33158), .A2(n44112), .Z(n11797) );
  NAND2_X2 U31994 ( .A1(n11229), .A2(n43601), .ZN(n43339) );
  NOR2_X1 U31996 ( .A1(n17860), .A2(n61202), .ZN(n56233) );
  OR2_X1 U31998 ( .A1(n55670), .A2(n55972), .Z(n11805) );
  NAND2_X2 U31999 ( .A1(n52036), .A2(n20891), .ZN(n55967) );
  NOR2_X2 U32002 ( .A1(n47516), .A2(n47494), .ZN(n47493) );
  NAND2_X1 U32005 ( .A1(n11825), .A2(n11822), .ZN(n29874) );
  NAND2_X1 U32006 ( .A1(n11824), .A2(n11823), .ZN(n11822) );
  NOR2_X1 U32007 ( .A1(n64708), .A2(n14247), .ZN(n11823) );
  NAND2_X1 U32008 ( .A1(n34553), .A2(n64499), .ZN(n11824) );
  INV_X4 U32009 ( .I(n11831), .ZN(n50576) );
  INV_X2 U32011 ( .I(n52719), .ZN(n56624) );
  XOR2_X1 U32013 ( .A1(n9885), .A2(n37120), .Z(n37121) );
  NAND2_X2 U32014 ( .A1(n16736), .A2(n24331), .ZN(n16403) );
  XOR2_X1 U32015 ( .A1(n10282), .A2(n46376), .Z(n46379) );
  XOR2_X1 U32016 ( .A1(n14513), .A2(n46377), .Z(n14514) );
  XOR2_X1 U32022 ( .A1(n11842), .A2(n12186), .Z(n12185) );
  XOR2_X1 U32024 ( .A1(n61927), .A2(n31901), .Z(n11847) );
  NOR2_X2 U32027 ( .A1(n11849), .A2(n19522), .ZN(n26670) );
  XOR2_X1 U32030 ( .A1(n23069), .A2(n10335), .Z(n52588) );
  XOR2_X1 U32032 ( .A1(n51677), .A2(n52610), .Z(n11853) );
  INV_X2 U32033 ( .I(n11855), .ZN(n41437) );
  NOR3_X1 U32034 ( .A1(n41428), .A2(n23967), .A3(n11855), .ZN(n39601) );
  AOI21_X1 U32035 ( .A1(n40698), .A2(n23967), .B(n11855), .ZN(n40376) );
  INV_X2 U32037 ( .I(n24154), .ZN(n32585) );
  XOR2_X1 U32038 ( .A1(n23613), .A2(n32749), .Z(n13429) );
  XOR2_X1 U32039 ( .A1(n30401), .A2(n62548), .Z(n32749) );
  XOR2_X1 U32040 ( .A1(n24154), .A2(n11856), .Z(n30401) );
  XNOR2_X1 U32041 ( .A1(n38966), .A2(n18132), .ZN(n39578) );
  XOR2_X1 U32042 ( .A1(n38848), .A2(n39769), .Z(n38966) );
  NAND2_X2 U32043 ( .A1(n36284), .A2(n36285), .ZN(n38848) );
  NAND2_X2 U32044 ( .A1(n24309), .A2(n24306), .ZN(n39769) );
  XOR2_X1 U32045 ( .A1(n39391), .A2(n22277), .Z(n18132) );
  INV_X1 U32047 ( .I(n27895), .ZN(n11859) );
  XOR2_X1 U32048 ( .A1(n11861), .A2(n26009), .Z(n52442) );
  NAND2_X1 U32050 ( .A1(n30135), .A2(n12907), .ZN(n11863) );
  NAND2_X2 U32053 ( .A1(n23056), .A2(n31039), .ZN(n31032) );
  NOR2_X2 U32057 ( .A1(n53421), .A2(n4481), .ZN(n53857) );
  NAND2_X1 U32060 ( .A1(n41169), .A2(n40645), .ZN(n13510) );
  NAND3_X1 U32063 ( .A1(n18608), .A2(n1471), .A3(n1384), .ZN(n46777) );
  XOR2_X1 U32066 ( .A1(n7410), .A2(n11877), .Z(n11879) );
  XOR2_X1 U32070 ( .A1(n5676), .A2(n44027), .Z(n44028) );
  XOR2_X1 U32072 ( .A1(n5676), .A2(n44394), .Z(n44395) );
  NOR2_X2 U32073 ( .A1(n57949), .A2(n49395), .ZN(n49330) );
  OAI21_X1 U32074 ( .A1(n20598), .A2(n64732), .B(n11895), .ZN(n40585) );
  NOR2_X2 U32078 ( .A1(n1436), .A2(n1561), .ZN(n11909) );
  XOR2_X1 U32080 ( .A1(n12596), .A2(n11911), .Z(n13553) );
  OR2_X1 U32081 ( .A1(n56318), .A2(n58755), .Z(n11916) );
  OR2_X1 U32082 ( .A1(n61727), .A2(n24032), .Z(n11917) );
  XOR2_X1 U32083 ( .A1(n11922), .A2(n11924), .Z(n42421) );
  XOR2_X1 U32084 ( .A1(n64714), .A2(n11925), .Z(n11924) );
  XOR2_X1 U32085 ( .A1(n11931), .A2(n18596), .Z(n18595) );
  XOR2_X1 U32086 ( .A1(n25443), .A2(n11930), .Z(n11931) );
  XOR2_X1 U32088 ( .A1(n19090), .A2(n11933), .Z(n31465) );
  XOR2_X1 U32089 ( .A1(n11934), .A2(n31692), .Z(n11933) );
  XOR2_X1 U32090 ( .A1(n31592), .A2(n11935), .Z(n11934) );
  XOR2_X1 U32091 ( .A1(n32387), .A2(n31426), .Z(n11935) );
  NOR2_X1 U32093 ( .A1(n29375), .A2(n11946), .ZN(n11945) );
  XOR2_X1 U32097 ( .A1(n14058), .A2(n11955), .Z(n51316) );
  XOR2_X1 U32098 ( .A1(n16280), .A2(n61883), .Z(n11956) );
  XOR2_X1 U32099 ( .A1(n12586), .A2(n20656), .Z(n11957) );
  XOR2_X1 U32101 ( .A1(n63487), .A2(n813), .Z(n11961) );
  NAND2_X1 U32103 ( .A1(n58983), .A2(n10422), .ZN(n49380) );
  AOI21_X1 U32104 ( .A1(n49377), .A2(n10422), .B(n49543), .ZN(n48781) );
  NAND2_X2 U32105 ( .A1(n47850), .A2(n15596), .ZN(n15595) );
  XOR2_X1 U32109 ( .A1(n24739), .A2(n11971), .Z(n11970) );
  XOR2_X1 U32110 ( .A1(n15096), .A2(n23678), .Z(n11971) );
  XOR2_X1 U32114 ( .A1(n11978), .A2(n16210), .Z(n28674) );
  XOR2_X1 U32115 ( .A1(n56155), .A2(n61380), .Z(n11978) );
  XOR2_X1 U32116 ( .A1(n62518), .A2(n56879), .Z(n42115) );
  XOR2_X1 U32117 ( .A1(n57448), .A2(n38305), .Z(n38306) );
  INV_X1 U32118 ( .I(n11984), .ZN(n53701) );
  NOR2_X1 U32119 ( .A1(n11984), .A2(n19475), .ZN(n53669) );
  OAI21_X1 U32120 ( .A1(n53696), .A2(n53697), .B(n11984), .ZN(n12323) );
  AOI21_X1 U32121 ( .A1(n53634), .A2(n11984), .B(n53633), .ZN(n53639) );
  INV_X2 U32122 ( .I(n11985), .ZN(n47680) );
  NOR2_X1 U32125 ( .A1(n59647), .A2(n51268), .ZN(n11990) );
  NOR2_X1 U32126 ( .A1(n11989), .A2(n10389), .ZN(n51251) );
  XOR2_X1 U32129 ( .A1(n11993), .A2(n12565), .Z(n12564) );
  NAND2_X1 U32130 ( .A1(n11994), .A2(n9725), .ZN(n15680) );
  NOR2_X1 U32131 ( .A1(n11994), .A2(n65128), .ZN(n40309) );
  NOR2_X1 U32132 ( .A1(n53600), .A2(n19062), .ZN(n11997) );
  NAND3_X2 U32133 ( .A1(n11999), .A2(n53609), .A3(n53608), .ZN(n11998) );
  XOR2_X1 U32136 ( .A1(n22940), .A2(n781), .Z(n12005) );
  XOR2_X1 U32140 ( .A1(n33192), .A2(n33191), .Z(n33202) );
  XOR2_X1 U32141 ( .A1(n12014), .A2(n12013), .Z(n33192) );
  XNOR2_X1 U32142 ( .A1(n33242), .A2(n22978), .ZN(n12014) );
  NAND3_X2 U32143 ( .A1(n29719), .A2(n29720), .A3(n19524), .ZN(n33242) );
  XOR2_X1 U32144 ( .A1(Key[70]), .A2(Ciphertext[135]), .Z(n12758) );
  INV_X1 U32147 ( .I(n59274), .ZN(n20810) );
  XOR2_X1 U32148 ( .A1(n12016), .A2(n32738), .Z(n32739) );
  XOR2_X1 U32149 ( .A1(n12019), .A2(n12017), .Z(n12016) );
  XOR2_X1 U32150 ( .A1(n12018), .A2(n32735), .Z(n12017) );
  INV_X1 U32151 ( .I(n57984), .ZN(n12018) );
  XOR2_X1 U32153 ( .A1(n20385), .A2(n14284), .Z(n12020) );
  NAND2_X2 U32154 ( .A1(n1863), .A2(n61383), .ZN(n30676) );
  NOR2_X2 U32155 ( .A1(n13935), .A2(n26780), .ZN(n28932) );
  XOR2_X1 U32156 ( .A1(n22350), .A2(n1623), .Z(n18644) );
  XOR2_X1 U32160 ( .A1(n32732), .A2(n12022), .Z(n25991) );
  INV_X1 U32161 ( .I(n32733), .ZN(n32468) );
  XOR2_X1 U32162 ( .A1(n32733), .A2(n33174), .Z(n33044) );
  XOR2_X1 U32163 ( .A1(n12022), .A2(n30918), .Z(n30920) );
  NAND2_X2 U32164 ( .A1(n41257), .A2(n7728), .ZN(n40797) );
  NAND2_X1 U32169 ( .A1(n26689), .A2(n12030), .ZN(n21840) );
  NAND2_X1 U32170 ( .A1(n26967), .A2(n12030), .ZN(n25645) );
  XOR2_X1 U32172 ( .A1(n6092), .A2(n39203), .Z(n39204) );
  NAND2_X2 U32174 ( .A1(n6654), .A2(n65222), .ZN(n49019) );
  XOR2_X1 U32176 ( .A1(n22551), .A2(n45057), .Z(n12038) );
  XOR2_X1 U32178 ( .A1(n44850), .A2(n51394), .Z(n12044) );
  NAND3_X1 U32183 ( .A1(n23651), .A2(n37940), .A3(n12050), .ZN(n33938) );
  AOI21_X1 U32185 ( .A1(n49314), .A2(n49608), .B(n49607), .ZN(n25040) );
  XOR2_X1 U32187 ( .A1(n52521), .A2(n50974), .Z(n23627) );
  XOR2_X1 U32188 ( .A1(n12052), .A2(n23069), .Z(n52521) );
  XOR2_X1 U32189 ( .A1(n52424), .A2(n51832), .Z(n12052) );
  XOR2_X1 U32193 ( .A1(n20931), .A2(n20554), .Z(n12055) );
  XOR2_X1 U32194 ( .A1(n324), .A2(n38445), .Z(n12056) );
  INV_X2 U32196 ( .I(n12062), .ZN(n23666) );
  XOR2_X1 U32198 ( .A1(n11448), .A2(n51239), .Z(n51240) );
  XOR2_X1 U32199 ( .A1(n11448), .A2(n50125), .Z(n14610) );
  XOR2_X1 U32200 ( .A1(n52334), .A2(n11448), .Z(n51490) );
  XOR2_X1 U32201 ( .A1(n11448), .A2(n52615), .Z(n52618) );
  XOR2_X1 U32202 ( .A1(n11448), .A2(n51395), .Z(n51396) );
  NOR2_X1 U32204 ( .A1(n10309), .A2(n29170), .ZN(n15195) );
  NAND2_X2 U32206 ( .A1(n12076), .A2(n12900), .ZN(n50283) );
  XOR2_X1 U32207 ( .A1(n12080), .A2(n12077), .Z(n33431) );
  XOR2_X1 U32208 ( .A1(n12078), .A2(n28931), .Z(n12077) );
  INV_X1 U32214 ( .I(n12085), .ZN(n27408) );
  INV_X2 U32215 ( .I(n12086), .ZN(n50601) );
  XOR2_X1 U32217 ( .A1(n52066), .A2(n50600), .Z(n12087) );
  NAND2_X2 U32218 ( .A1(n35027), .A2(n10340), .ZN(n18136) );
  NAND2_X2 U32219 ( .A1(n12112), .A2(n14523), .ZN(n29207) );
  XOR2_X1 U32223 ( .A1(n52544), .A2(n19969), .Z(n12092) );
  XOR2_X1 U32225 ( .A1(n51996), .A2(n12096), .Z(n12095) );
  INV_X2 U32226 ( .I(n11501), .ZN(n12097) );
  NAND2_X1 U32229 ( .A1(n12101), .A2(n38342), .ZN(n25824) );
  INV_X2 U32230 ( .I(n12102), .ZN(n17299) );
  XOR2_X1 U32232 ( .A1(n12105), .A2(n12104), .Z(n12103) );
  XOR2_X1 U32233 ( .A1(n32722), .A2(n43937), .Z(n12104) );
  XOR2_X1 U32234 ( .A1(n33033), .A2(n32721), .Z(n12105) );
  XOR2_X1 U32235 ( .A1(n20673), .A2(n14665), .Z(n33033) );
  XOR2_X1 U32236 ( .A1(n32725), .A2(n12107), .Z(n12106) );
  XOR2_X1 U32237 ( .A1(n17299), .A2(n12665), .Z(n32725) );
  NOR2_X1 U32242 ( .A1(n35602), .A2(n12116), .ZN(n25225) );
  NAND3_X1 U32243 ( .A1(n35602), .A2(n36262), .A3(n12116), .ZN(n34885) );
  NAND3_X1 U32244 ( .A1(n1311), .A2(n3856), .A3(n12116), .ZN(n35180) );
  NAND2_X1 U32246 ( .A1(n33413), .A2(n12116), .ZN(n24625) );
  NAND2_X1 U32248 ( .A1(n12125), .A2(n4257), .ZN(n31280) );
  AND2_X1 U32252 ( .A1(n29203), .A2(n12131), .Z(n12130) );
  INV_X1 U32254 ( .I(n12141), .ZN(n17686) );
  OAI22_X1 U32255 ( .A1(n35417), .A2(n35418), .B1(n35416), .B2(n12141), .ZN(
        n35419) );
  OAI21_X1 U32256 ( .A1(n13591), .A2(n56773), .B(n12142), .ZN(n13590) );
  NAND2_X2 U32257 ( .A1(n51563), .A2(n7209), .ZN(n12142) );
  OAI21_X1 U32260 ( .A1(n35327), .A2(n23717), .B(n12148), .ZN(n32142) );
  NAND2_X2 U32266 ( .A1(n41384), .A2(n41386), .ZN(n17212) );
  XOR2_X1 U32271 ( .A1(n32281), .A2(n12172), .Z(n13552) );
  XOR2_X1 U32272 ( .A1(n32280), .A2(n12781), .Z(n12172) );
  INV_X2 U32274 ( .I(n29170), .ZN(n28267) );
  NAND2_X2 U32275 ( .A1(n29171), .A2(n23769), .ZN(n29170) );
  INV_X2 U32276 ( .I(n12179), .ZN(n18098) );
  INV_X2 U32278 ( .I(n12185), .ZN(n16736) );
  INV_X2 U32279 ( .I(n13857), .ZN(n24331) );
  NAND2_X2 U32283 ( .A1(n1715), .A2(n22282), .ZN(n43359) );
  OAI22_X1 U32284 ( .A1(n7050), .A2(n47825), .B1(n1652), .B2(n10088), .ZN(
        n12198) );
  NOR2_X1 U32288 ( .A1(n22861), .A2(n13826), .ZN(n12221) );
  XOR2_X1 U32289 ( .A1(n25695), .A2(n13179), .Z(n44817) );
  XOR2_X1 U32291 ( .A1(n25982), .A2(n43067), .Z(n46127) );
  NAND2_X1 U32292 ( .A1(n12231), .A2(n7104), .ZN(n12230) );
  XOR2_X1 U32294 ( .A1(n44388), .A2(n44082), .Z(n12232) );
  NAND2_X2 U32296 ( .A1(n25438), .A2(n43132), .ZN(n43133) );
  OR2_X1 U32302 ( .A1(n57001), .A2(n10237), .Z(n12251) );
  NAND2_X2 U32303 ( .A1(n19735), .A2(n9338), .ZN(n53301) );
  INV_X2 U32304 ( .I(n12254), .ZN(n25804) );
  XOR2_X1 U32306 ( .A1(n26060), .A2(n13674), .Z(n12257) );
  XOR2_X1 U32310 ( .A1(n244), .A2(n44352), .Z(n44353) );
  XOR2_X1 U32311 ( .A1(n244), .A2(n59984), .Z(n44433) );
  XOR2_X1 U32312 ( .A1(n244), .A2(n45069), .Z(n45071) );
  INV_X2 U32314 ( .I(n23649), .ZN(n28452) );
  XOR2_X1 U32315 ( .A1(n26785), .A2(Key[47]), .Z(n27859) );
  INV_X1 U32316 ( .I(n28604), .ZN(n12263) );
  NOR2_X2 U32318 ( .A1(n17951), .A2(n45437), .ZN(n47372) );
  NAND2_X1 U32321 ( .A1(n27605), .A2(n28299), .ZN(n12279) );
  INV_X1 U32322 ( .I(n20883), .ZN(n25969) );
  XOR2_X1 U32323 ( .A1(n40100), .A2(n12285), .Z(n12284) );
  OAI21_X1 U32325 ( .A1(n36170), .A2(n12288), .B(n36121), .ZN(n36122) );
  AOI21_X1 U32328 ( .A1(n35131), .A2(n12288), .B(n36170), .ZN(n35133) );
  NAND2_X1 U32329 ( .A1(n36175), .A2(n12288), .ZN(n36183) );
  MUX2_X1 U32330 ( .I0(n22295), .I1(n21801), .S(n12288), .Z(n35136) );
  INV_X4 U32331 ( .I(n22169), .ZN(n12288) );
  NOR2_X2 U32333 ( .A1(n13810), .A2(n30677), .ZN(n30685) );
  NAND4_X2 U32334 ( .A1(n1099), .A2(n22690), .A3(n12292), .A4(n12291), .ZN(
        n51828) );
  NAND2_X1 U32335 ( .A1(n48731), .A2(n48737), .ZN(n12291) );
  XOR2_X1 U32337 ( .A1(n50670), .A2(n51548), .Z(n12297) );
  XOR2_X1 U32338 ( .A1(n23883), .A2(n50669), .Z(n12298) );
  NOR3_X2 U32343 ( .A1(n12302), .A2(n32141), .A3(n34329), .ZN(n17132) );
  INV_X2 U32345 ( .I(n25701), .ZN(n22236) );
  INV_X2 U32351 ( .I(n14876), .ZN(n23917) );
  NOR2_X1 U32357 ( .A1(n42415), .A2(n42065), .ZN(n12313) );
  INV_X4 U32358 ( .I(n12314), .ZN(n19611) );
  XOR2_X1 U32360 ( .A1(n25804), .A2(n49825), .Z(n12315) );
  XOR2_X1 U32361 ( .A1(n19125), .A2(n20742), .Z(n12317) );
  XOR2_X1 U32362 ( .A1(n14970), .A2(n14971), .Z(n39720) );
  XOR2_X1 U32363 ( .A1(n12318), .A2(n17221), .Z(Plaintext[35]) );
  XOR2_X1 U32364 ( .A1(n53687), .A2(n53692), .Z(n12321) );
  INV_X1 U32365 ( .I(n17869), .ZN(n24744) );
  NOR3_X2 U32368 ( .A1(n12336), .A2(n12334), .A3(n12332), .ZN(n12331) );
  NAND3_X1 U32369 ( .A1(n48004), .A2(n49195), .A3(n65005), .ZN(n12333) );
  NAND2_X1 U32370 ( .A1(n1261), .A2(n49525), .ZN(n12335) );
  XOR2_X1 U32373 ( .A1(n33828), .A2(n793), .Z(n27794) );
  XOR2_X1 U32374 ( .A1(n9254), .A2(n30795), .Z(n30796) );
  NAND2_X1 U32375 ( .A1(n46096), .A2(n61422), .ZN(n44134) );
  NAND2_X1 U32376 ( .A1(n47014), .A2(n61422), .ZN(n23676) );
  NOR3_X1 U32379 ( .A1(n62784), .A2(n12346), .A3(n26665), .ZN(n27571) );
  INV_X2 U32382 ( .I(n12349), .ZN(n25427) );
  NAND2_X1 U32383 ( .A1(n12350), .A2(n34994), .ZN(n30458) );
  AOI21_X1 U32384 ( .A1(n21008), .A2(n12350), .B(n12983), .ZN(n12982) );
  NAND4_X2 U32386 ( .A1(n35959), .A2(n11272), .A3(n36472), .A4(n12352), .ZN(
        n35960) );
  AOI21_X1 U32389 ( .A1(n21811), .A2(n22189), .B(n12354), .ZN(n21810) );
  NOR2_X2 U32392 ( .A1(n47304), .A2(n26180), .ZN(n47292) );
  INV_X2 U32394 ( .I(n25471), .ZN(n47304) );
  NOR2_X2 U32395 ( .A1(n45929), .A2(n61932), .ZN(n12360) );
  NAND2_X2 U32396 ( .A1(n57377), .A2(n12361), .ZN(n25349) );
  AOI21_X1 U32400 ( .A1(n20034), .A2(n19290), .B(n29621), .ZN(n12365) );
  NOR2_X1 U32401 ( .A1(n29280), .A2(n28125), .ZN(n12366) );
  NOR2_X1 U32402 ( .A1(n12369), .A2(n12368), .ZN(n12367) );
  OAI22_X1 U32403 ( .A1(n25967), .A2(n47921), .B1(n49049), .B2(n47920), .ZN(
        n12369) );
  XOR2_X1 U32404 ( .A1(n12371), .A2(n44931), .Z(n20462) );
  XOR2_X1 U32405 ( .A1(n13359), .A2(n44930), .Z(n12372) );
  XOR2_X1 U32407 ( .A1(n46650), .A2(n46317), .Z(n12375) );
  NAND3_X2 U32412 ( .A1(n21862), .A2(n21861), .A3(n42165), .ZN(n46321) );
  NAND2_X2 U32414 ( .A1(n37536), .A2(n42598), .ZN(n12378) );
  AOI21_X1 U32418 ( .A1(n41029), .A2(n12384), .B(n13139), .ZN(n13138) );
  INV_X1 U32419 ( .I(n62593), .ZN(n48916) );
  NOR2_X2 U32420 ( .A1(n62200), .A2(n16411), .ZN(n47073) );
  NAND2_X1 U32421 ( .A1(n43286), .A2(n10111), .ZN(n18172) );
  INV_X1 U32422 ( .I(n43282), .ZN(n41710) );
  INV_X1 U32424 ( .I(n35460), .ZN(n12387) );
  NAND2_X1 U32425 ( .A1(n42387), .A2(n40174), .ZN(n41532) );
  NAND2_X2 U32427 ( .A1(n48227), .A2(n48226), .ZN(n50359) );
  XOR2_X1 U32429 ( .A1(n1622), .A2(n1901), .Z(n51320) );
  INV_X1 U32436 ( .I(n42354), .ZN(n41988) );
  INV_X2 U32437 ( .I(n33116), .ZN(n21592) );
  NAND2_X2 U32440 ( .A1(n12413), .A2(n14039), .ZN(n17759) );
  XOR2_X1 U32441 ( .A1(n31637), .A2(n12415), .Z(n13739) );
  NAND2_X1 U32443 ( .A1(n12420), .A2(n29803), .ZN(n21063) );
  NOR2_X1 U32444 ( .A1(n16082), .A2(n12420), .ZN(n21023) );
  NOR2_X1 U32445 ( .A1(n12423), .A2(n26606), .ZN(n26331) );
  XOR2_X1 U32451 ( .A1(n2905), .A2(n12436), .Z(n17473) );
  XOR2_X1 U32452 ( .A1(n25422), .A2(n21826), .Z(n25421) );
  NOR2_X2 U32458 ( .A1(n31247), .A2(n1435), .ZN(n12443) );
  OR2_X1 U32459 ( .A1(n43697), .A2(n43698), .Z(n12444) );
  OR2_X1 U32460 ( .A1(n43696), .A2(n43695), .Z(n12445) );
  XOR2_X1 U32461 ( .A1(n1197), .A2(n50639), .Z(n12448) );
  XOR2_X1 U32462 ( .A1(n52154), .A2(n22747), .Z(n12449) );
  AOI21_X1 U32463 ( .A1(n57389), .A2(n12453), .B(n41054), .ZN(n41641) );
  NAND4_X2 U32468 ( .A1(n12461), .A2(n12460), .A3(n36974), .A4(n37252), .ZN(
        n12459) );
  NAND2_X1 U32471 ( .A1(n48287), .A2(n1380), .ZN(n22931) );
  AOI21_X1 U32472 ( .A1(n50424), .A2(n50417), .B(n1380), .ZN(n50418) );
  OAI21_X1 U32473 ( .A1(n48755), .A2(n1380), .B(n2878), .ZN(n45462) );
  NAND2_X1 U32481 ( .A1(n18757), .A2(n16533), .ZN(n12482) );
  XOR2_X1 U32482 ( .A1(n3523), .A2(n43902), .Z(n33882) );
  XOR2_X1 U32483 ( .A1(n3523), .A2(n32551), .Z(n32553) );
  INV_X2 U32484 ( .I(n24953), .ZN(n52165) );
  NAND2_X2 U32487 ( .A1(n1429), .A2(n24083), .ZN(n31358) );
  NOR2_X2 U32488 ( .A1(n12493), .A2(n12494), .ZN(n12492) );
  INV_X2 U32495 ( .I(n33780), .ZN(n13352) );
  NOR2_X2 U32496 ( .A1(n16451), .A2(n64387), .ZN(n33780) );
  NOR2_X2 U32497 ( .A1(n22169), .A2(n36121), .ZN(n36420) );
  XOR2_X1 U32501 ( .A1(n32176), .A2(n12505), .Z(n12519) );
  XOR2_X1 U32503 ( .A1(n17299), .A2(n18748), .Z(n32666) );
  INV_X1 U32505 ( .I(n13620), .ZN(n37849) );
  AOI21_X1 U32507 ( .A1(n12506), .A2(n24286), .B(n18879), .ZN(n33128) );
  XOR2_X1 U32508 ( .A1(n12507), .A2(n46143), .Z(n46144) );
  XOR2_X1 U32509 ( .A1(n12507), .A2(n44101), .Z(n44102) );
  XOR2_X1 U32510 ( .A1(n46651), .A2(n12507), .Z(n46652) );
  NAND2_X1 U32511 ( .A1(n20491), .A2(n59755), .ZN(n30869) );
  OAI21_X1 U32512 ( .A1(n33774), .A2(n61108), .B(n12512), .ZN(n12511) );
  NOR2_X1 U32513 ( .A1(n12513), .A2(n22176), .ZN(n12512) );
  AND2_X2 U32521 ( .A1(n20716), .A2(n14876), .Z(n27111) );
  NAND2_X1 U32523 ( .A1(n23339), .A2(n42357), .ZN(n22208) );
  INV_X4 U32525 ( .I(n33319), .ZN(n32684) );
  AND2_X1 U32526 ( .A1(n209), .A2(n48653), .Z(n15828) );
  NAND2_X1 U32527 ( .A1(n17686), .A2(n36777), .ZN(n17685) );
  INV_X2 U32532 ( .I(n20739), .ZN(n24485) );
  NAND2_X2 U32537 ( .A1(n1353), .A2(n31189), .ZN(n31177) );
  INV_X4 U32538 ( .I(n19329), .ZN(n47827) );
  INV_X4 U32540 ( .I(n42259), .ZN(n41906) );
  INV_X1 U32541 ( .I(n25156), .ZN(n23880) );
  NOR2_X2 U32542 ( .A1(n28854), .A2(n29310), .ZN(n29325) );
  INV_X4 U32548 ( .I(n18852), .ZN(n55820) );
  NOR2_X1 U32551 ( .A1(n29197), .A2(n29198), .ZN(n14301) );
  INV_X1 U32556 ( .I(Ciphertext[150]), .ZN(n14104) );
  OAI21_X1 U32557 ( .A1(n49874), .A2(n12917), .B(n63679), .ZN(n17288) );
  INV_X4 U32560 ( .I(n27533), .ZN(n27523) );
  OAI22_X1 U32561 ( .A1(n53269), .A2(n14267), .B1(n53268), .B2(n22889), .ZN(
        n53270) );
  INV_X1 U32562 ( .I(n27206), .ZN(n26594) );
  NOR3_X1 U32567 ( .A1(n26299), .A2(n23041), .A3(n26298), .ZN(n26304) );
  NOR2_X1 U32569 ( .A1(n28356), .A2(n28357), .ZN(n13055) );
  NOR2_X1 U32570 ( .A1(n42071), .A2(n1193), .ZN(n20039) );
  INV_X4 U32577 ( .I(n51911), .ZN(n52630) );
  INV_X4 U32583 ( .I(n48555), .ZN(n48544) );
  INV_X2 U32584 ( .I(n19926), .ZN(n19994) );
  BUF_X4 U32585 ( .I(n39427), .Z(n43290) );
  AOI22_X1 U32586 ( .A1(n41409), .A2(n41408), .B1(n41404), .B2(n17063), .ZN(
        n13264) );
  NOR3_X2 U32587 ( .A1(n24167), .A2(n48719), .A3(n50291), .ZN(n48724) );
  NAND2_X2 U32589 ( .A1(n1814), .A2(n15756), .ZN(n35038) );
  NAND2_X2 U32591 ( .A1(n43626), .A2(n43415), .ZN(n43553) );
  NAND2_X2 U32593 ( .A1(n14708), .A2(n56942), .ZN(n56916) );
  NAND3_X1 U32594 ( .A1(n12531), .A2(n12528), .A3(n56164), .ZN(n12527) );
  INV_X1 U32595 ( .I(n12582), .ZN(n32949) );
  INV_X4 U32610 ( .I(n15378), .ZN(n40295) );
  INV_X4 U32611 ( .I(n36070), .ZN(n36304) );
  NOR2_X1 U32613 ( .A1(n11108), .A2(n50267), .ZN(n21834) );
  INV_X2 U32615 ( .I(n21510), .ZN(n25202) );
  NOR2_X2 U32619 ( .A1(n56084), .A2(n56106), .ZN(n56048) );
  NAND2_X1 U32622 ( .A1(n56163), .A2(n12525), .ZN(n12526) );
  XOR2_X1 U32623 ( .A1(n12527), .A2(n56165), .Z(Plaintext[146]) );
  XOR2_X1 U32624 ( .A1(n51590), .A2(n19029), .Z(n12533) );
  NOR2_X2 U32626 ( .A1(n23130), .A2(n27786), .ZN(n20623) );
  XOR2_X1 U32627 ( .A1(n12542), .A2(n12541), .Z(n12540) );
  XOR2_X1 U32628 ( .A1(n18276), .A2(n13705), .Z(n12541) );
  XOR2_X1 U32629 ( .A1(n12545), .A2(n929), .Z(n12542) );
  INV_X1 U32632 ( .I(n18276), .ZN(n38819) );
  XOR2_X1 U32633 ( .A1(n1412), .A2(n38574), .Z(n39257) );
  INV_X1 U32635 ( .I(n12548), .ZN(n17502) );
  NOR4_X2 U32636 ( .A1(n17796), .A2(n12554), .A3(n12550), .A4(n12549), .ZN(
        n17671) );
  NAND2_X2 U32641 ( .A1(n12562), .A2(n12561), .ZN(n33034) );
  INV_X2 U32642 ( .I(n12564), .ZN(n12605) );
  XOR2_X1 U32643 ( .A1(n51200), .A2(n12566), .Z(n12565) );
  XOR2_X1 U32646 ( .A1(n32315), .A2(n10535), .Z(n12568) );
  XOR2_X1 U32647 ( .A1(n32246), .A2(n59546), .Z(n32420) );
  XOR2_X1 U32648 ( .A1(n32726), .A2(n32316), .Z(n12569) );
  NAND2_X1 U32652 ( .A1(n36965), .A2(n1527), .ZN(n35445) );
  INV_X2 U32653 ( .I(n20902), .ZN(n17951) );
  NOR3_X1 U32654 ( .A1(n21706), .A2(n1372), .A3(n12573), .ZN(n52829) );
  NOR2_X1 U32656 ( .A1(n12574), .A2(n57039), .ZN(n53207) );
  NAND2_X1 U32658 ( .A1(n12574), .A2(n57051), .ZN(n50806) );
  OAI21_X1 U32659 ( .A1(n12575), .A2(n53255), .B(n53275), .ZN(n53261) );
  XOR2_X1 U32661 ( .A1(n39001), .A2(n39534), .Z(n12578) );
  XOR2_X1 U32664 ( .A1(n12585), .A2(n12583), .Z(n25803) );
  XOR2_X1 U32665 ( .A1(n12584), .A2(n51973), .Z(n12583) );
  XOR2_X1 U32666 ( .A1(n50795), .A2(n11071), .Z(n12584) );
  NAND2_X1 U32668 ( .A1(n12588), .A2(n12587), .ZN(n31604) );
  OAI22_X1 U32669 ( .A1(n26881), .A2(n12589), .B1(n28168), .B2(n29608), .ZN(
        n26882) );
  INV_X2 U32671 ( .I(n12590), .ZN(n19282) );
  XOR2_X1 U32672 ( .A1(n12591), .A2(n17703), .Z(n17702) );
  XOR2_X1 U32673 ( .A1(n12591), .A2(n58077), .Z(n33138) );
  XOR2_X1 U32674 ( .A1(n32503), .A2(n17700), .Z(n19250) );
  NOR2_X1 U32675 ( .A1(n12592), .A2(n61986), .ZN(n40210) );
  AOI21_X1 U32676 ( .A1(n22459), .A2(n40215), .B(n12592), .ZN(n40216) );
  MUX2_X1 U32677 ( .I0(n38040), .I1(n38035), .S(n6581), .Z(n38039) );
  OAI21_X1 U32678 ( .A1(n26104), .A2(n48420), .B(n12595), .ZN(n26103) );
  NAND2_X1 U32680 ( .A1(n37455), .A2(n10907), .ZN(n36882) );
  AOI22_X1 U32681 ( .A1(n35832), .A2(n37444), .B1(n62992), .B2(n10907), .ZN(
        n35851) );
  XOR2_X1 U32684 ( .A1(n58341), .A2(n23288), .Z(n12599) );
  OAI21_X2 U32687 ( .A1(n50948), .A2(n50949), .B(n12602), .ZN(n24787) );
  NOR2_X2 U32688 ( .A1(n25168), .A2(n12605), .ZN(n25167) );
  XOR2_X1 U32689 ( .A1(n12608), .A2(n1888), .Z(n45812) );
  XOR2_X1 U32691 ( .A1(n12607), .A2(n61010), .Z(n46254) );
  INV_X2 U32693 ( .I(n12609), .ZN(n39007) );
  XNOR2_X1 U32695 ( .A1(n39407), .A2(n12610), .ZN(n12609) );
  XOR2_X1 U32696 ( .A1(n12611), .A2(n937), .Z(n12610) );
  XOR2_X1 U32698 ( .A1(Ciphertext[9]), .A2(Key[148]), .Z(n22861) );
  OR2_X1 U32699 ( .A1(n21315), .A2(n12612), .Z(n16236) );
  XOR2_X1 U32700 ( .A1(n20429), .A2(n1106), .Z(n12614) );
  NAND2_X1 U32702 ( .A1(n12615), .A2(n24861), .ZN(n15073) );
  NAND2_X2 U32704 ( .A1(n35794), .A2(n61458), .ZN(n34388) );
  NAND2_X2 U32707 ( .A1(n20349), .A2(n19567), .ZN(n53535) );
  OAI21_X1 U32708 ( .A1(n12580), .A2(n49722), .B(n12626), .ZN(n12625) );
  XOR2_X1 U32712 ( .A1(n9602), .A2(n30898), .Z(n32497) );
  NOR3_X2 U32714 ( .A1(n12638), .A2(n12637), .A3(n12636), .ZN(n12635) );
  NOR4_X1 U32718 ( .A1(n12645), .A2(n43925), .A3(n61743), .A4(n12644), .ZN(
        n12643) );
  NOR2_X2 U32719 ( .A1(n23565), .A2(n43600), .ZN(n12646) );
  NAND2_X1 U32722 ( .A1(n14289), .A2(n12647), .ZN(n18003) );
  NAND3_X1 U32723 ( .A1(n64548), .A2(n59967), .A3(n12647), .ZN(n47720) );
  NAND3_X1 U32724 ( .A1(n11901), .A2(n47882), .A3(n12648), .ZN(n43598) );
  NAND2_X1 U32725 ( .A1(n51717), .A2(n53877), .ZN(n12651) );
  OR2_X1 U32726 ( .A1(n54243), .A2(n54209), .Z(n15991) );
  INV_X2 U32728 ( .I(n35019), .ZN(n25124) );
  NAND3_X2 U32729 ( .A1(n35018), .A2(n35017), .A3(n35016), .ZN(n35019) );
  XOR2_X1 U32731 ( .A1(n63016), .A2(n12655), .Z(n12654) );
  XOR2_X1 U32732 ( .A1(n46279), .A2(n43499), .Z(n12655) );
  XNOR2_X1 U32733 ( .A1(n43496), .A2(n14514), .ZN(n44587) );
  NOR2_X1 U32734 ( .A1(n12741), .A2(n29609), .ZN(n29607) );
  XOR2_X1 U32735 ( .A1(n32513), .A2(n60372), .Z(n33076) );
  XOR2_X1 U32736 ( .A1(n33242), .A2(n23771), .Z(n32513) );
  NAND3_X2 U32737 ( .A1(n12661), .A2(n24842), .A3(n19628), .ZN(n23771) );
  XOR2_X1 U32739 ( .A1(n12663), .A2(n32581), .Z(n12662) );
  INV_X2 U32741 ( .I(n12668), .ZN(n39406) );
  XOR2_X1 U32742 ( .A1(n39406), .A2(n39405), .Z(n39590) );
  INV_X2 U32745 ( .I(n12676), .ZN(n15758) );
  XNOR2_X1 U32746 ( .A1(Ciphertext[187]), .A2(Key[50]), .ZN(n12676) );
  NAND2_X2 U32748 ( .A1(n35570), .A2(n36026), .ZN(n34822) );
  XOR2_X1 U32752 ( .A1(n12681), .A2(n25060), .Z(n13290) );
  XOR2_X1 U32753 ( .A1(n60642), .A2(n50148), .Z(n50149) );
  XOR2_X1 U32757 ( .A1(n19282), .A2(n31672), .Z(n12686) );
  NOR2_X2 U32761 ( .A1(n6095), .A2(n54461), .ZN(n12692) );
  NOR2_X2 U32762 ( .A1(n12694), .A2(n8290), .ZN(n43742) );
  XOR2_X1 U32764 ( .A1(n6927), .A2(n62487), .Z(n39191) );
  NOR2_X2 U32765 ( .A1(n7086), .A2(n49177), .ZN(n21367) );
  NOR2_X1 U32766 ( .A1(n11060), .A2(n33600), .ZN(n33305) );
  NOR2_X1 U32768 ( .A1(n33012), .A2(n11060), .ZN(n33013) );
  NAND2_X1 U32769 ( .A1(n59534), .A2(n63888), .ZN(n33298) );
  NOR2_X2 U32771 ( .A1(n12696), .A2(n55445), .ZN(n21395) );
  NAND2_X1 U32772 ( .A1(n12696), .A2(n55306), .ZN(n55307) );
  NAND3_X1 U32773 ( .A1(n12696), .A2(n55440), .A3(n55442), .ZN(n52490) );
  NAND2_X1 U32774 ( .A1(n55322), .A2(n12696), .ZN(n55008) );
  NAND3_X1 U32776 ( .A1(n19819), .A2(n19818), .A3(n12696), .ZN(n19817) );
  NAND2_X1 U32777 ( .A1(n55309), .A2(n12696), .ZN(n12695) );
  NAND2_X2 U32778 ( .A1(n55443), .A2(n55444), .ZN(n12696) );
  NAND2_X1 U32781 ( .A1(n25680), .A2(n2754), .ZN(n50417) );
  NOR3_X1 U32782 ( .A1(n45464), .A2(n23063), .A3(n2754), .ZN(n45444) );
  INV_X4 U32783 ( .I(n15743), .ZN(n37181) );
  NAND2_X2 U32785 ( .A1(n21499), .A2(n25202), .ZN(n29145) );
  XOR2_X1 U32787 ( .A1(n12710), .A2(n763), .Z(n32046) );
  XOR2_X1 U32788 ( .A1(n32045), .A2(n12711), .Z(n12710) );
  XOR2_X1 U32789 ( .A1(n17299), .A2(n32043), .Z(n12711) );
  XOR2_X1 U32793 ( .A1(n46251), .A2(n12715), .Z(n12714) );
  XOR2_X1 U32794 ( .A1(n46150), .A2(n45364), .Z(n12715) );
  XOR2_X1 U32795 ( .A1(n12716), .A2(n50642), .Z(n50643) );
  NAND2_X1 U32797 ( .A1(n42601), .A2(n429), .ZN(n12717) );
  NAND2_X2 U32798 ( .A1(n12739), .A2(n4613), .ZN(n28174) );
  XOR2_X1 U32800 ( .A1(n13989), .A2(n64837), .Z(n12728) );
  NAND2_X1 U32802 ( .A1(n33409), .A2(n57830), .ZN(n33410) );
  NAND2_X2 U32804 ( .A1(n23816), .A2(n15790), .ZN(n19223) );
  NAND2_X1 U32808 ( .A1(n49195), .A2(n48845), .ZN(n12753) );
  XOR2_X1 U32809 ( .A1(n12754), .A2(n1062), .Z(n13438) );
  INV_X2 U32811 ( .I(n12758), .ZN(n15790) );
  NAND2_X2 U32812 ( .A1(n15790), .A2(n14930), .ZN(n29603) );
  OAI21_X1 U32813 ( .A1(n47045), .A2(n13072), .B(n1480), .ZN(n17810) );
  NAND2_X2 U32814 ( .A1(n23301), .A2(n48586), .ZN(n47154) );
  XOR2_X1 U32816 ( .A1(n786), .A2(n14882), .Z(n12771) );
  INV_X2 U32817 ( .I(n12772), .ZN(n24353) );
  XOR2_X1 U32818 ( .A1(n39661), .A2(n57403), .Z(n39677) );
  XOR2_X1 U32819 ( .A1(n39494), .A2(n3604), .Z(n39661) );
  XOR2_X1 U32821 ( .A1(n23600), .A2(n15735), .Z(n12773) );
  NAND2_X2 U32823 ( .A1(n17029), .A2(n16081), .ZN(n17623) );
  INV_X1 U32824 ( .I(n52235), .ZN(n52827) );
  INV_X2 U32826 ( .I(n37755), .ZN(n42267) );
  XOR2_X1 U32827 ( .A1(n19282), .A2(n12780), .Z(n13368) );
  XOR2_X1 U32828 ( .A1(n22363), .A2(n12781), .Z(n18211) );
  INV_X1 U32830 ( .I(n17233), .ZN(n18307) );
  INV_X2 U32835 ( .I(n7074), .ZN(n12797) );
  XOR2_X1 U32837 ( .A1(n12799), .A2(n50516), .Z(n50517) );
  XOR2_X1 U32838 ( .A1(n12799), .A2(n51946), .Z(n50560) );
  XOR2_X1 U32839 ( .A1(n12799), .A2(n51983), .Z(n51984) );
  INV_X1 U32840 ( .I(n61702), .ZN(n35737) );
  XOR2_X1 U32852 ( .A1(n12813), .A2(n20836), .Z(n12812) );
  XOR2_X1 U32854 ( .A1(n33138), .A2(n32182), .Z(n12815) );
  NOR2_X1 U32856 ( .A1(n1232), .A2(n9338), .ZN(n12827) );
  OR2_X1 U32861 ( .A1(n36194), .A2(n36412), .Z(n12831) );
  NAND3_X2 U32862 ( .A1(n19081), .A2(n19083), .A3(n12832), .ZN(n53115) );
  XOR2_X1 U32867 ( .A1(n12854), .A2(n46311), .Z(n46314) );
  XOR2_X1 U32868 ( .A1(n12853), .A2(n12852), .Z(n46311) );
  XOR2_X1 U32869 ( .A1(n41333), .A2(n20900), .Z(n12852) );
  XOR2_X1 U32870 ( .A1(n15734), .A2(n44993), .Z(n12853) );
  XOR2_X1 U32871 ( .A1(n46310), .A2(n19335), .Z(n12854) );
  NAND2_X2 U32872 ( .A1(n28504), .A2(n27846), .ZN(n28517) );
  XOR2_X1 U32873 ( .A1(n12857), .A2(n774), .Z(n12856) );
  XOR2_X1 U32874 ( .A1(n55765), .A2(n53989), .Z(n12857) );
  XOR2_X1 U32879 ( .A1(n37979), .A2(n12860), .Z(n39337) );
  XOR2_X1 U32883 ( .A1(n50939), .A2(n50940), .Z(n12869) );
  XOR2_X1 U32884 ( .A1(n21513), .A2(n24211), .Z(n19759) );
  XOR2_X1 U32885 ( .A1(n15755), .A2(n12880), .Z(n21513) );
  INV_X1 U32888 ( .I(n12871), .ZN(n30710) );
  NAND2_X2 U32890 ( .A1(n31038), .A2(n31040), .ZN(n12871) );
  NAND2_X1 U32897 ( .A1(n1787), .A2(n18385), .ZN(n35575) );
  XOR2_X1 U32898 ( .A1(n36338), .A2(n36742), .Z(n12883) );
  NAND2_X1 U32899 ( .A1(n46944), .A2(n10193), .ZN(n45731) );
  NOR2_X2 U32900 ( .A1(n25604), .A2(n23874), .ZN(n12923) );
  INV_X1 U32902 ( .I(n37509), .ZN(n12889) );
  XOR2_X1 U32903 ( .A1(n38921), .A2(n38920), .Z(n12891) );
  NAND3_X2 U32907 ( .A1(n38940), .A2(n12947), .A3(n12948), .ZN(n12960) );
  NAND2_X1 U32908 ( .A1(n12895), .A2(n64364), .ZN(n40406) );
  NAND2_X1 U32909 ( .A1(n12895), .A2(n22525), .ZN(n41420) );
  AOI21_X1 U32910 ( .A1(n12895), .A2(n10173), .B(n65184), .ZN(n41214) );
  NAND2_X1 U32911 ( .A1(n20652), .A2(n62272), .ZN(n39870) );
  NAND2_X2 U32913 ( .A1(n20053), .A2(n20052), .ZN(n12908) );
  XOR2_X1 U32918 ( .A1(n45282), .A2(n12911), .Z(n45300) );
  XOR2_X1 U32919 ( .A1(n61662), .A2(n1013), .Z(n12911) );
  NAND2_X2 U32923 ( .A1(n53871), .A2(n12917), .ZN(n53549) );
  XOR2_X1 U32925 ( .A1(n12921), .A2(n46590), .Z(n15377) );
  XOR2_X1 U32926 ( .A1(n12920), .A2(n19766), .Z(n46590) );
  XOR2_X1 U32927 ( .A1(n23652), .A2(n46216), .Z(n12920) );
  NAND2_X1 U32930 ( .A1(n53321), .A2(n12923), .ZN(n16776) );
  INV_X2 U32936 ( .I(n14672), .ZN(n23343) );
  XOR2_X1 U32938 ( .A1(n12940), .A2(n20234), .Z(n38574) );
  NOR3_X2 U32941 ( .A1(n15302), .A2(n15300), .A3(n15299), .ZN(n51081) );
  XOR2_X1 U32943 ( .A1(n15885), .A2(n21107), .Z(n12945) );
  XOR2_X1 U32945 ( .A1(n3717), .A2(n20411), .Z(n20410) );
  INV_X2 U32946 ( .I(n12954), .ZN(n23834) );
  NAND2_X2 U32947 ( .A1(n12953), .A2(n551), .ZN(n33720) );
  NAND2_X2 U32948 ( .A1(n34980), .A2(n12953), .ZN(n33486) );
  INV_X2 U32949 ( .I(n18214), .ZN(n48082) );
  XOR2_X1 U32952 ( .A1(n12963), .A2(n39465), .Z(n38924) );
  XOR2_X1 U32953 ( .A1(n38877), .A2(n25375), .Z(n39465) );
  OAI22_X1 U32956 ( .A1(n61676), .A2(n20199), .B1(n49575), .B2(n12966), .ZN(
        n49578) );
  INV_X1 U32958 ( .I(n12968), .ZN(n48637) );
  NOR2_X1 U32959 ( .A1(n48636), .A2(n12968), .ZN(n19774) );
  NOR2_X1 U32960 ( .A1(n48632), .A2(n12968), .ZN(n48633) );
  AOI21_X1 U32962 ( .A1(n48631), .A2(n12968), .B(n48511), .ZN(n47215) );
  NOR2_X1 U32966 ( .A1(n12975), .A2(n41934), .ZN(n41250) );
  NAND2_X1 U32967 ( .A1(n15051), .A2(n12975), .ZN(n17094) );
  INV_X2 U32968 ( .I(n889), .ZN(n34970) );
  XOR2_X1 U32969 ( .A1(n30934), .A2(n19478), .Z(n12976) );
  OR2_X2 U32971 ( .A1(n22378), .A2(n26621), .Z(n29860) );
  OAI21_X1 U32972 ( .A1(n10091), .A2(n2323), .B(n63421), .ZN(n12983) );
  NOR2_X2 U32973 ( .A1(n60693), .A2(n41132), .ZN(n17915) );
  XOR2_X1 U32976 ( .A1(n19530), .A2(n12987), .Z(n12986) );
  XOR2_X1 U32977 ( .A1(n11070), .A2(n50183), .Z(n12987) );
  XOR2_X1 U32978 ( .A1(n10335), .A2(n50936), .Z(n13974) );
  XOR2_X1 U32979 ( .A1(n61423), .A2(n52587), .Z(n51154) );
  NOR3_X2 U32980 ( .A1(n12995), .A2(n48635), .A3(n12992), .ZN(n12991) );
  NAND2_X1 U32983 ( .A1(n28615), .A2(n63330), .ZN(n13007) );
  NAND3_X1 U32984 ( .A1(n28605), .A2(n21854), .A3(n23649), .ZN(n13011) );
  INV_X1 U32986 ( .I(n25886), .ZN(n31502) );
  INV_X1 U32987 ( .I(n13022), .ZN(n56263) );
  NOR2_X1 U32990 ( .A1(n21427), .A2(n13024), .ZN(n21428) );
  NAND2_X2 U32993 ( .A1(n13042), .A2(n13039), .ZN(n17994) );
  INV_X2 U32994 ( .I(n19527), .ZN(n32568) );
  XOR2_X1 U32995 ( .A1(n13045), .A2(n13046), .Z(n13044) );
  NOR2_X1 U32998 ( .A1(n22856), .A2(n13047), .ZN(n26057) );
  NAND2_X1 U32999 ( .A1(n26594), .A2(n13047), .ZN(n26348) );
  INV_X1 U33000 ( .I(n61094), .ZN(n41223) );
  NAND3_X1 U33001 ( .A1(n20652), .A2(n13048), .A3(n58794), .ZN(n13052) );
  NAND2_X2 U33004 ( .A1(n1714), .A2(n61107), .ZN(n14051) );
  OR2_X1 U33006 ( .A1(n60962), .A2(n24696), .Z(n13057) );
  AND2_X1 U33007 ( .A1(n56553), .A2(n56554), .Z(n13059) );
  XOR2_X1 U33008 ( .A1(n39383), .A2(n13061), .Z(n13270) );
  XOR2_X1 U33011 ( .A1(n24859), .A2(n13062), .Z(n13061) );
  XOR2_X1 U33014 ( .A1(n32027), .A2(n882), .Z(n13064) );
  XOR2_X1 U33015 ( .A1(n32186), .A2(n20617), .Z(n32027) );
  INV_X1 U33016 ( .I(n12468), .ZN(n13067) );
  INV_X1 U33018 ( .I(n61107), .ZN(n13074) );
  NAND2_X2 U33019 ( .A1(n1763), .A2(n13078), .ZN(n19410) );
  NAND2_X2 U33020 ( .A1(n31147), .A2(n31141), .ZN(n22579) );
  XOR2_X1 U33021 ( .A1(n52087), .A2(n52086), .Z(n52088) );
  INV_X2 U33022 ( .I(n43553), .ZN(n17245) );
  INV_X2 U33023 ( .I(n13082), .ZN(n21878) );
  INV_X2 U33024 ( .I(n19876), .ZN(n34783) );
  NAND3_X1 U33028 ( .A1(n61940), .A2(n60562), .A3(n36224), .ZN(n34700) );
  AOI22_X1 U33031 ( .A1(n32444), .A2(n35591), .B1(n61940), .B2(n32445), .ZN(
        n32450) );
  NAND2_X1 U33034 ( .A1(n29171), .A2(n28260), .ZN(n28264) );
  INV_X1 U33035 ( .I(n13100), .ZN(n42546) );
  XOR2_X1 U33036 ( .A1(n42115), .A2(n25426), .Z(n44273) );
  INV_X1 U33037 ( .I(n13103), .ZN(n13600) );
  OAI21_X1 U33038 ( .A1(n53875), .A2(n13815), .B(n53545), .ZN(n13103) );
  OAI22_X2 U33043 ( .A1(n61723), .A2(n13112), .B1(n54435), .B2(n52957), .ZN(
        n52963) );
  XOR2_X1 U33045 ( .A1(n13809), .A2(n13114), .Z(n38780) );
  XOR2_X1 U33046 ( .A1(n61506), .A2(n13115), .Z(n36934) );
  NAND2_X1 U33047 ( .A1(n24788), .A2(n47970), .ZN(n48822) );
  OR2_X1 U33048 ( .A1(n47025), .A2(n18321), .Z(n47033) );
  NAND2_X2 U33049 ( .A1(n13655), .A2(n47034), .ZN(n18321) );
  NAND2_X2 U33050 ( .A1(n13122), .A2(n22526), .ZN(n49467) );
  NAND3_X2 U33051 ( .A1(n41423), .A2(n66), .A3(n38935), .ZN(n13125) );
  INV_X1 U33058 ( .I(n49882), .ZN(n13148) );
  XOR2_X1 U33061 ( .A1(n1057), .A2(n44906), .Z(n13151) );
  XOR2_X1 U33062 ( .A1(n45147), .A2(n44829), .Z(n13152) );
  XOR2_X1 U33063 ( .A1(n64971), .A2(n23872), .Z(n45147) );
  XOR2_X1 U33065 ( .A1(n16582), .A2(n850), .Z(n13153) );
  XOR2_X1 U33066 ( .A1(n43807), .A2(n64050), .Z(n43623) );
  XOR2_X1 U33068 ( .A1(n51082), .A2(n13155), .Z(n51083) );
  NAND2_X1 U33069 ( .A1(n1359), .A2(n17909), .ZN(n27416) );
  NAND2_X1 U33070 ( .A1(n1359), .A2(n29162), .ZN(n13188) );
  NOR2_X2 U33075 ( .A1(n43750), .A2(n26166), .ZN(n47729) );
  NAND2_X2 U33077 ( .A1(n31777), .A2(n16198), .ZN(n35886) );
  XOR2_X1 U33079 ( .A1(n5244), .A2(n38892), .Z(n22166) );
  INV_X1 U33081 ( .I(n42509), .ZN(n13168) );
  NAND2_X1 U33087 ( .A1(n13174), .A2(n29726), .ZN(n30021) );
  INV_X1 U33089 ( .I(n35886), .ZN(n35881) );
  NAND2_X1 U33091 ( .A1(n15828), .A2(n22233), .ZN(n13178) );
  XOR2_X1 U33092 ( .A1(n44488), .A2(n13179), .Z(n44938) );
  XOR2_X1 U33093 ( .A1(n21724), .A2(n13179), .Z(n41742) );
  INV_X1 U33094 ( .I(n38526), .ZN(n13183) );
  INV_X2 U33095 ( .I(n13184), .ZN(n25214) );
  XOR2_X1 U33098 ( .A1(n10635), .A2(n22152), .Z(n48703) );
  INV_X1 U33104 ( .I(n13196), .ZN(n13197) );
  INV_X2 U33109 ( .I(n13205), .ZN(n44779) );
  XOR2_X1 U33110 ( .A1(n38453), .A2(n23695), .Z(n37708) );
  NAND2_X2 U33113 ( .A1(n43309), .A2(n23314), .ZN(n43992) );
  NAND2_X1 U33114 ( .A1(n13210), .A2(n63247), .ZN(n13209) );
  XOR2_X1 U33116 ( .A1(n13213), .A2(n13214), .Z(n32409) );
  XOR2_X1 U33119 ( .A1(n51930), .A2(n51599), .Z(n51600) );
  INV_X2 U33120 ( .I(n13218), .ZN(n54657) );
  XOR2_X1 U33121 ( .A1(n13221), .A2(n13220), .Z(n13219) );
  XOR2_X1 U33124 ( .A1(n20304), .A2(n16041), .Z(n19146) );
  INV_X2 U33129 ( .I(n33486), .ZN(n34995) );
  OAI21_X1 U33130 ( .A1(n41495), .A2(n14214), .B(n13229), .ZN(n14044) );
  NAND2_X2 U33131 ( .A1(n13232), .A2(n25803), .ZN(n57046) );
  XOR2_X1 U33132 ( .A1(n51406), .A2(n50768), .Z(n13233) );
  NOR2_X2 U33133 ( .A1(n14214), .A2(n4274), .ZN(n13242) );
  INV_X2 U33134 ( .I(n17994), .ZN(n49525) );
  XOR2_X1 U33136 ( .A1(n1189), .A2(n16119), .Z(n13246) );
  XOR2_X1 U33143 ( .A1(n46680), .A2(n44315), .Z(n13257) );
  OAI21_X1 U33146 ( .A1(n54210), .A2(n54209), .B(n13263), .ZN(n23236) );
  NAND4_X1 U33147 ( .A1(n15991), .A2(n17433), .A3(n13263), .A4(n51880), .ZN(
        n17432) );
  XOR2_X1 U33148 ( .A1(n39368), .A2(n39367), .Z(n13272) );
  XOR2_X1 U33150 ( .A1(n13274), .A2(n26167), .Z(n19335) );
  XOR2_X1 U33151 ( .A1(n13513), .A2(n24992), .Z(n13274) );
  XOR2_X1 U33153 ( .A1(n31924), .A2(n13277), .Z(n13276) );
  NOR2_X2 U33156 ( .A1(n25047), .A2(n25467), .ZN(n53381) );
  INV_X2 U33157 ( .I(n13288), .ZN(n25047) );
  XOR2_X1 U33158 ( .A1(n22111), .A2(n1898), .Z(n44355) );
  XOR2_X1 U33159 ( .A1(n13801), .A2(n13281), .Z(n46312) );
  XOR2_X1 U33160 ( .A1(n13283), .A2(n46127), .Z(n48483) );
  NAND2_X1 U33162 ( .A1(n42638), .A2(n13284), .ZN(n43200) );
  OAI21_X1 U33163 ( .A1(n13284), .A2(n43189), .B(n61744), .ZN(n40782) );
  NOR2_X2 U33164 ( .A1(n43188), .A2(n43513), .ZN(n13284) );
  XOR2_X1 U33166 ( .A1(n13286), .A2(n54168), .Z(n50500) );
  XOR2_X1 U33167 ( .A1(n13286), .A2(n23754), .Z(n51232) );
  XOR2_X1 U33170 ( .A1(n63021), .A2(n13285), .Z(n51052) );
  XOR2_X1 U33176 ( .A1(n31917), .A2(n13291), .Z(n20457) );
  NAND2_X2 U33180 ( .A1(n22352), .A2(n28552), .ZN(n26217) );
  MUX2_X1 U33182 ( .I0(n13292), .I1(n53598), .S(n23169), .Z(n53193) );
  XOR2_X1 U33184 ( .A1(n24076), .A2(n13295), .Z(n13294) );
  XOR2_X1 U33185 ( .A1(n11448), .A2(n50622), .Z(n13295) );
  NAND2_X2 U33190 ( .A1(n13305), .A2(n13304), .ZN(n13306) );
  NAND2_X1 U33191 ( .A1(n21057), .A2(n38023), .ZN(n13308) );
  INV_X1 U33194 ( .I(n38061), .ZN(n13315) );
  NAND2_X2 U33195 ( .A1(n15533), .A2(n13320), .ZN(n27789) );
  XOR2_X1 U33197 ( .A1(n324), .A2(n16300), .Z(n13324) );
  NAND2_X2 U33199 ( .A1(n13326), .A2(n27523), .ZN(n27525) );
  AND3_X1 U33200 ( .A1(n9548), .A2(n20929), .A3(n28349), .Z(n13326) );
  AND2_X1 U33201 ( .A1(n19159), .A2(n27525), .Z(n16101) );
  NAND2_X2 U33203 ( .A1(n1604), .A2(n54945), .ZN(n13328) );
  NOR2_X2 U33204 ( .A1(n13331), .A2(n13330), .ZN(n54570) );
  NAND3_X2 U33206 ( .A1(n27588), .A2(n27589), .A3(n27590), .ZN(n27591) );
  OR2_X1 U33209 ( .A1(n13345), .A2(n36431), .Z(n13343) );
  AOI21_X1 U33212 ( .A1(n46764), .A2(n10624), .B(n46763), .ZN(n13347) );
  INV_X2 U33213 ( .I(n48561), .ZN(n13348) );
  NOR2_X2 U33217 ( .A1(n40416), .A2(n7165), .ZN(n41466) );
  INV_X2 U33218 ( .I(n25132), .ZN(n40416) );
  NOR2_X1 U33222 ( .A1(n13356), .A2(n59959), .ZN(n17315) );
  NOR2_X1 U33223 ( .A1(n47903), .A2(n13356), .ZN(n22412) );
  NAND2_X2 U33224 ( .A1(n23969), .A2(n1483), .ZN(n13356) );
  NOR2_X2 U33225 ( .A1(n27661), .A2(n28488), .ZN(n26824) );
  NOR2_X1 U33228 ( .A1(n1530), .A2(n13358), .ZN(n36624) );
  XOR2_X1 U33229 ( .A1(n13365), .A2(n10531), .Z(n20789) );
  XOR2_X1 U33230 ( .A1(n33271), .A2(n13368), .Z(n13367) );
  XOR2_X1 U33231 ( .A1(n31366), .A2(n31365), .Z(n33271) );
  XOR2_X1 U33232 ( .A1(n64610), .A2(n25530), .Z(n13369) );
  INV_X1 U33233 ( .I(n21238), .ZN(n23181) );
  XOR2_X1 U33234 ( .A1(n21238), .A2(n789), .Z(n36659) );
  NAND2_X1 U33238 ( .A1(n23071), .A2(n23737), .ZN(n13375) );
  INV_X2 U33239 ( .I(n13383), .ZN(n14317) );
  XOR2_X1 U33242 ( .A1(n19859), .A2(n51018), .Z(n52055) );
  AND2_X1 U33243 ( .A1(n1868), .A2(n31098), .Z(n28205) );
  NAND2_X1 U33245 ( .A1(n13781), .A2(n25362), .ZN(n32955) );
  NAND2_X2 U33246 ( .A1(n61703), .A2(n36220), .ZN(n36436) );
  INV_X1 U33250 ( .I(n25912), .ZN(n13397) );
  NOR2_X2 U33252 ( .A1(n28448), .A2(n28446), .ZN(n13399) );
  INV_X2 U33254 ( .I(n37130), .ZN(n38551) );
  OR2_X1 U33256 ( .A1(n16628), .A2(n15757), .Z(n18498) );
  XOR2_X1 U33257 ( .A1(n13409), .A2(n15379), .Z(n13479) );
  XOR2_X1 U33259 ( .A1(Ciphertext[114]), .A2(Key[19]), .Z(n13439) );
  NAND2_X1 U33262 ( .A1(n13413), .A2(n21304), .ZN(n21639) );
  INV_X4 U33265 ( .I(n13418), .ZN(n20138) );
  XOR2_X1 U33266 ( .A1(n44754), .A2(n62065), .Z(n24133) );
  XOR2_X1 U33270 ( .A1(n13429), .A2(n13427), .Z(n24965) );
  XOR2_X1 U33271 ( .A1(n31692), .A2(n13428), .Z(n13427) );
  XOR2_X1 U33274 ( .A1(n13435), .A2(n39647), .Z(n13436) );
  XOR2_X1 U33275 ( .A1(n39646), .A2(n39645), .Z(n13435) );
  XNOR2_X1 U33276 ( .A1(n13437), .A2(n13436), .ZN(n13434) );
  INV_X2 U33277 ( .I(n23458), .ZN(n45401) );
  INV_X2 U33278 ( .I(n13439), .ZN(n28448) );
  NAND3_X2 U33280 ( .A1(n17080), .A2(n48638), .A3(n17079), .ZN(n49582) );
  NAND2_X2 U33281 ( .A1(n3335), .A2(n13440), .ZN(n49355) );
  INV_X2 U33286 ( .I(n13456), .ZN(n23904) );
  XOR2_X1 U33289 ( .A1(n39273), .A2(n39272), .Z(n13457) );
  XOR2_X1 U33291 ( .A1(n10449), .A2(n794), .Z(n46125) );
  XOR2_X1 U33292 ( .A1(n10255), .A2(n13463), .Z(n44018) );
  XOR2_X1 U33293 ( .A1(n44341), .A2(n13463), .Z(n44342) );
  XOR2_X1 U33298 ( .A1(n33034), .A2(n50634), .Z(n13464) );
  NAND2_X2 U33299 ( .A1(n48847), .A2(n13471), .ZN(n49512) );
  NOR2_X1 U33302 ( .A1(n29514), .A2(n1838), .ZN(n18762) );
  OAI22_X1 U33304 ( .A1(n21134), .A2(n17413), .B1(n17414), .B2(n1838), .ZN(
        n29854) );
  MUX2_X1 U33305 ( .I0(n30955), .I1(n30954), .S(n1838), .Z(n30957) );
  NAND2_X2 U33306 ( .A1(n7311), .A2(n33614), .ZN(n32460) );
  XOR2_X1 U33308 ( .A1(Ciphertext[19]), .A2(Key[26]), .Z(n13694) );
  INV_X2 U33310 ( .I(n13479), .ZN(n15378) );
  XOR2_X1 U33311 ( .A1(n13480), .A2(n38942), .Z(n39312) );
  XOR2_X1 U33312 ( .A1(n19803), .A2(n50943), .Z(n13480) );
  XOR2_X1 U33313 ( .A1(n11577), .A2(n49405), .Z(n22675) );
  XOR2_X1 U33314 ( .A1(n9231), .A2(n11577), .Z(n50323) );
  XOR2_X1 U33315 ( .A1(n11577), .A2(n51024), .Z(n51025) );
  AOI22_X1 U33316 ( .A1(n31048), .A2(n31049), .B1(n31047), .B2(n13481), .ZN(
        n14724) );
  INV_X2 U33317 ( .I(n47704), .ZN(n24615) );
  NOR2_X1 U33318 ( .A1(n22229), .A2(n13489), .ZN(n22875) );
  NAND2_X1 U33319 ( .A1(n57011), .A2(n13489), .ZN(n17455) );
  AOI21_X1 U33320 ( .A1(n56386), .A2(n13489), .B(n56542), .ZN(n56387) );
  XOR2_X1 U33323 ( .A1(n13508), .A2(n13507), .Z(n13781) );
  AOI21_X1 U33324 ( .A1(n13509), .A2(n18836), .B(n20637), .ZN(n13511) );
  NOR2_X1 U33325 ( .A1(n41168), .A2(n41167), .ZN(n13509) );
  XOR2_X1 U33327 ( .A1(n13515), .A2(n23989), .Z(n26610) );
  XOR2_X1 U33328 ( .A1(n26292), .A2(n54748), .Z(n13515) );
  XOR2_X1 U33331 ( .A1(n13518), .A2(n13519), .Z(n25868) );
  XOR2_X1 U33332 ( .A1(n50737), .A2(n52031), .Z(n13518) );
  XOR2_X1 U33333 ( .A1(n52145), .A2(n50732), .Z(n13519) );
  XOR2_X1 U33334 ( .A1(n13520), .A2(n32753), .Z(n32755) );
  XOR2_X1 U33335 ( .A1(n13520), .A2(n32660), .Z(n32662) );
  XOR2_X1 U33336 ( .A1(n63099), .A2(n13520), .Z(n33075) );
  NOR2_X2 U33340 ( .A1(n13525), .A2(n287), .ZN(n42249) );
  OAI21_X1 U33344 ( .A1(n914), .A2(n13536), .B(n34995), .ZN(n34996) );
  XOR2_X1 U33346 ( .A1(n51721), .A2(n13541), .Z(n13539) );
  XOR2_X1 U33347 ( .A1(n23422), .A2(n51720), .Z(n13541) );
  INV_X1 U33356 ( .I(n14005), .ZN(n49280) );
  NAND2_X2 U33360 ( .A1(n48688), .A2(n2810), .ZN(n48690) );
  NOR2_X1 U33361 ( .A1(n13558), .A2(n61900), .ZN(n29812) );
  INV_X2 U33365 ( .I(n25362), .ZN(n13559) );
  AND2_X1 U33368 ( .A1(n21805), .A2(n29120), .Z(n13565) );
  NAND2_X1 U33369 ( .A1(n13566), .A2(n45715), .ZN(n45720) );
  OAI21_X1 U33372 ( .A1(n47772), .A2(n64878), .B(n13566), .ZN(n47778) );
  OAI22_X1 U33375 ( .A1(n52249), .A2(n57068), .B1(n21079), .B2(n13567), .ZN(
        n52250) );
  INV_X4 U33377 ( .I(n57079), .ZN(n13567) );
  XOR2_X1 U33379 ( .A1(n32370), .A2(n18855), .Z(n13568) );
  XOR2_X1 U33380 ( .A1(n32368), .A2(n15187), .Z(n13570) );
  XOR2_X1 U33381 ( .A1(n15186), .A2(n9609), .Z(n32368) );
  NOR3_X2 U33385 ( .A1(n27910), .A2(n27908), .A3(n27909), .ZN(n13578) );
  XOR2_X1 U33390 ( .A1(n13579), .A2(n13580), .Z(n19648) );
  XOR2_X1 U33393 ( .A1(n15444), .A2(n58234), .Z(n13584) );
  NAND4_X2 U33394 ( .A1(n13586), .A2(n48592), .A3(n48593), .A4(n13585), .ZN(
        n48944) );
  OR2_X1 U33396 ( .A1(n48583), .A2(n13587), .Z(n13586) );
  NOR2_X2 U33399 ( .A1(n56775), .A2(n23030), .ZN(n51563) );
  INV_X2 U33400 ( .I(n13592), .ZN(n48586) );
  NAND2_X2 U33404 ( .A1(n13608), .A2(n13607), .ZN(n35265) );
  NAND2_X1 U33405 ( .A1(n15408), .A2(n904), .ZN(n13607) );
  INV_X1 U33406 ( .I(n13609), .ZN(n13608) );
  AOI21_X1 U33407 ( .A1(n35195), .A2(n35286), .B(n15408), .ZN(n13609) );
  XOR2_X1 U33409 ( .A1(n20886), .A2(n23267), .Z(n13613) );
  XOR2_X1 U33410 ( .A1(n37742), .A2(n13616), .Z(n13615) );
  XOR2_X1 U33411 ( .A1(n59788), .A2(n783), .Z(n13616) );
  XOR2_X1 U33412 ( .A1(n39451), .A2(n24147), .Z(n13619) );
  XOR2_X1 U33413 ( .A1(n6749), .A2(n63019), .Z(n21368) );
  XOR2_X1 U33415 ( .A1(n44242), .A2(n43944), .Z(n24992) );
  XOR2_X1 U33420 ( .A1(n14299), .A2(n1621), .Z(n18537) );
  NAND2_X2 U33423 ( .A1(n18918), .A2(n49548), .ZN(n23612) );
  XOR2_X1 U33424 ( .A1(n37848), .A2(n38062), .Z(n13634) );
  XOR2_X1 U33425 ( .A1(n38323), .A2(n39292), .Z(n13635) );
  XOR2_X1 U33427 ( .A1(n51284), .A2(n50518), .Z(n13642) );
  XOR2_X1 U33430 ( .A1(n51748), .A2(n52465), .Z(n51943) );
  INV_X1 U33434 ( .I(n8478), .ZN(n29123) );
  NAND2_X2 U33437 ( .A1(n13666), .A2(n1783), .ZN(n37943) );
  NAND2_X1 U33439 ( .A1(n13667), .A2(n53355), .ZN(n53329) );
  OAI21_X1 U33440 ( .A1(n16778), .A2(n13667), .B(n53373), .ZN(n16777) );
  AOI22_X1 U33441 ( .A1(n29247), .A2(n29778), .B1(n29246), .B2(n61175), .ZN(
        n25882) );
  NAND2_X1 U33442 ( .A1(n29779), .A2(n13336), .ZN(n29782) );
  NAND2_X1 U33443 ( .A1(n29783), .A2(n13336), .ZN(n29785) );
  OR2_X2 U33445 ( .A1(n13675), .A2(n48435), .Z(n52421) );
  OAI21_X1 U33446 ( .A1(n25528), .A2(n25529), .B(n48444), .ZN(n13675) );
  XNOR2_X1 U33447 ( .A1(n52421), .A2(n52587), .ZN(n13674) );
  NAND2_X2 U33448 ( .A1(n48458), .A2(n48457), .ZN(n52587) );
  XOR2_X1 U33449 ( .A1(n13720), .A2(n13681), .Z(n53213) );
  OR2_X1 U33450 ( .A1(n50261), .A2(n50336), .Z(n13682) );
  XOR2_X1 U33452 ( .A1(n24248), .A2(n38945), .Z(n13685) );
  XOR2_X1 U33453 ( .A1(n38941), .A2(n39358), .Z(n13686) );
  XOR2_X1 U33454 ( .A1(n24018), .A2(n30402), .Z(n38941) );
  XOR2_X1 U33455 ( .A1(n51987), .A2(n51986), .Z(n52473) );
  OAI21_X1 U33457 ( .A1(n48365), .A2(n13692), .B(n48364), .ZN(n48371) );
  XOR2_X1 U33458 ( .A1(n21152), .A2(n13696), .Z(n15950) );
  OR2_X1 U33459 ( .A1(n24737), .A2(n33961), .Z(n13698) );
  NAND2_X1 U33461 ( .A1(n34952), .A2(n57166), .ZN(n33753) );
  MUX2_X1 U33462 ( .I0(n26622), .I1(n26623), .S(n28383), .Z(n26632) );
  XOR2_X1 U33465 ( .A1(n3208), .A2(n46352), .Z(n21568) );
  NOR2_X1 U33466 ( .A1(n54193), .A2(n54194), .ZN(n13714) );
  XOR2_X1 U33470 ( .A1(n15719), .A2(n13721), .Z(n51160) );
  OR2_X1 U33471 ( .A1(n45492), .A2(n13728), .Z(n13727) );
  NAND2_X2 U33472 ( .A1(n13730), .A2(n43778), .ZN(n43913) );
  NAND2_X2 U33474 ( .A1(n18693), .A2(n41863), .ZN(n43924) );
  NOR2_X1 U33476 ( .A1(n8808), .A2(n13734), .ZN(n21880) );
  AOI21_X1 U33477 ( .A1(n13767), .A2(n13734), .B(n4798), .ZN(n37070) );
  NOR2_X2 U33478 ( .A1(n28349), .A2(n27533), .ZN(n28350) );
  XOR2_X1 U33479 ( .A1(n14730), .A2(n49670), .Z(n26072) );
  XOR2_X1 U33482 ( .A1(n21084), .A2(n61874), .Z(n13740) );
  INV_X2 U33483 ( .I(n54110), .ZN(n13743) );
  INV_X2 U33485 ( .I(n13747), .ZN(n20554) );
  INV_X2 U33486 ( .I(n48711), .ZN(n49671) );
  NAND2_X1 U33490 ( .A1(n42968), .A2(n13750), .ZN(n13749) );
  NAND2_X1 U33491 ( .A1(n12312), .A2(n13751), .ZN(n43459) );
  NAND2_X1 U33492 ( .A1(n43467), .A2(n13751), .ZN(n41758) );
  AOI21_X1 U33493 ( .A1(n42966), .A2(n13751), .B(n43471), .ZN(n42967) );
  INV_X2 U33494 ( .I(n13752), .ZN(n19638) );
  NOR2_X1 U33499 ( .A1(n61435), .A2(n1727), .ZN(n16289) );
  OAI21_X1 U33501 ( .A1(n36688), .A2(n13767), .B(n37393), .ZN(n36689) );
  NAND2_X1 U33504 ( .A1(n35316), .A2(n13770), .ZN(n31951) );
  AOI22_X1 U33505 ( .A1(n7345), .A2(n77), .B1(n35763), .B2(n13770), .ZN(n35766) );
  XOR2_X1 U33506 ( .A1(n43332), .A2(n13772), .Z(n13771) );
  XOR2_X1 U33507 ( .A1(n44085), .A2(n13773), .Z(n13772) );
  XOR2_X1 U33508 ( .A1(n845), .A2(n32286), .Z(n43332) );
  AND2_X1 U33509 ( .A1(n36182), .A2(n36183), .Z(n13780) );
  XOR2_X1 U33511 ( .A1(n18730), .A2(n18729), .Z(n32308) );
  INV_X1 U33512 ( .I(n13782), .ZN(n47668) );
  NOR2_X2 U33516 ( .A1(n48028), .A2(n48024), .ZN(n13787) );
  NAND2_X2 U33518 ( .A1(n13891), .A2(n13893), .ZN(n13799) );
  NAND2_X1 U33521 ( .A1(n22929), .A2(n26732), .ZN(n13804) );
  NOR2_X2 U33524 ( .A1(n15674), .A2(n43100), .ZN(n42007) );
  NAND2_X2 U33526 ( .A1(n1894), .A2(n27524), .ZN(n27204) );
  XOR2_X1 U33527 ( .A1(n11142), .A2(n39636), .Z(n39637) );
  XOR2_X1 U33528 ( .A1(n24151), .A2(n54888), .Z(n39448) );
  XOR2_X1 U33529 ( .A1(n19418), .A2(n11142), .Z(n37267) );
  NAND3_X2 U33530 ( .A1(n11627), .A2(n24893), .A3(n47674), .ZN(n47401) );
  NOR2_X2 U33532 ( .A1(n13824), .A2(n13823), .ZN(n42027) );
  XOR2_X1 U33535 ( .A1(n18204), .A2(n17985), .Z(n33154) );
  XOR2_X1 U33536 ( .A1(n10292), .A2(n782), .Z(n50071) );
  XOR2_X1 U33537 ( .A1(n13831), .A2(n4265), .Z(n51064) );
  NAND2_X1 U33541 ( .A1(n55659), .A2(n61321), .ZN(n55660) );
  XOR2_X1 U33545 ( .A1(n45393), .A2(n45316), .Z(n13841) );
  OAI21_X1 U33546 ( .A1(n13848), .A2(n13847), .B(n10294), .ZN(n13846) );
  NOR2_X1 U33547 ( .A1(n41126), .A2(n17212), .ZN(n13847) );
  INV_X1 U33548 ( .I(n19570), .ZN(n13850) );
  NAND3_X2 U33551 ( .A1(n37495), .A2(n13856), .A3(n13855), .ZN(n19008) );
  AND2_X1 U33552 ( .A1(n37489), .A2(n17038), .Z(n13855) );
  NOR2_X2 U33555 ( .A1(n16782), .A2(n33929), .ZN(n33933) );
  OAI22_X1 U33556 ( .A1(n7132), .A2(n10160), .B1(n57300), .B2(n13866), .ZN(
        n13870) );
  NAND3_X1 U33557 ( .A1(n15118), .A2(n13874), .A3(n15117), .ZN(n13873) );
  INV_X1 U33558 ( .I(n16569), .ZN(n13874) );
  NOR2_X2 U33560 ( .A1(n18886), .A2(n1326), .ZN(n52122) );
  NAND2_X1 U33566 ( .A1(n1475), .A2(n14630), .ZN(n13881) );
  NOR3_X1 U33567 ( .A1(n13882), .A2(n20700), .A3(n42119), .ZN(n42123) );
  XOR2_X1 U33569 ( .A1(n44359), .A2(n13883), .Z(n20226) );
  XOR2_X1 U33571 ( .A1(n23687), .A2(n13883), .Z(n44494) );
  OAI22_X1 U33574 ( .A1(n49865), .A2(n50262), .B1(n49867), .B2(n49866), .ZN(
        n13886) );
  NAND2_X1 U33575 ( .A1(n48430), .A2(n48431), .ZN(n13887) );
  XOR2_X1 U33577 ( .A1(n52415), .A2(n51576), .Z(n13896) );
  XOR2_X1 U33578 ( .A1(n21700), .A2(n13897), .Z(n52637) );
  NOR2_X2 U33579 ( .A1(n1154), .A2(n13901), .ZN(n13900) );
  XOR2_X1 U33581 ( .A1(n13906), .A2(n13903), .Z(n15723) );
  XOR2_X1 U33582 ( .A1(n38990), .A2(n13905), .Z(n13904) );
  XOR2_X1 U33586 ( .A1(n17463), .A2(n31446), .Z(n30354) );
  INV_X1 U33591 ( .I(n1133), .ZN(n13921) );
  NAND2_X1 U33592 ( .A1(n48663), .A2(n26139), .ZN(n13932) );
  INV_X2 U33594 ( .I(n41920), .ZN(n24990) );
  NAND2_X2 U33595 ( .A1(n28780), .A2(n28779), .ZN(n28933) );
  XOR2_X1 U33597 ( .A1(n58839), .A2(n946), .Z(n13936) );
  NOR2_X1 U33600 ( .A1(n19438), .A2(n23654), .ZN(n39397) );
  NAND2_X2 U33601 ( .A1(n21050), .A2(n42489), .ZN(n19438) );
  XNOR2_X1 U33604 ( .A1(n49817), .A2(n51030), .ZN(n13944) );
  XOR2_X1 U33607 ( .A1(n23389), .A2(n13956), .Z(n18544) );
  XOR2_X1 U33608 ( .A1(n19886), .A2(n13956), .Z(n31760) );
  XOR2_X1 U33609 ( .A1(n2259), .A2(n13956), .Z(n31930) );
  XOR2_X1 U33610 ( .A1(n33285), .A2(n13956), .Z(n33288) );
  XOR2_X1 U33611 ( .A1(n31861), .A2(n13956), .Z(n31862) );
  XOR2_X1 U33612 ( .A1(n13958), .A2(n44894), .Z(n13957) );
  NOR2_X1 U33615 ( .A1(n13960), .A2(n56108), .ZN(n56032) );
  XOR2_X1 U33622 ( .A1(n13974), .A2(n52429), .Z(n50937) );
  NOR2_X1 U33626 ( .A1(n13978), .A2(n42385), .ZN(n41529) );
  INV_X2 U33627 ( .I(n14714), .ZN(n25657) );
  XOR2_X1 U33629 ( .A1(n13986), .A2(n52106), .Z(n54998) );
  XOR2_X1 U33630 ( .A1(n13987), .A2(n20674), .Z(n13986) );
  XOR2_X1 U33631 ( .A1(n52094), .A2(n52093), .Z(n13987) );
  XOR2_X1 U33635 ( .A1(n33044), .A2(n19058), .Z(n13992) );
  MUX2_X1 U33638 ( .I0(n36326), .I1(n36819), .S(n36831), .Z(n13994) );
  XOR2_X1 U33641 ( .A1(n46677), .A2(n46676), .Z(n13998) );
  XOR2_X1 U33645 ( .A1(n14003), .A2(n39383), .Z(n14002) );
  XOR2_X1 U33646 ( .A1(n39396), .A2(n39394), .Z(n14003) );
  NAND2_X1 U33650 ( .A1(n1472), .A2(n14007), .ZN(n48033) );
  OR2_X1 U33654 ( .A1(n40029), .A2(n14018), .Z(n14017) );
  XOR2_X1 U33655 ( .A1(Ciphertext[117]), .A2(Key[136]), .Z(n28446) );
  XOR2_X1 U33658 ( .A1(n2666), .A2(n51814), .Z(n30898) );
  XOR2_X1 U33660 ( .A1(n14023), .A2(n37078), .Z(n37173) );
  XOR2_X1 U33663 ( .A1(n32129), .A2(n20357), .Z(n33145) );
  XOR2_X1 U33664 ( .A1(n20573), .A2(n32130), .Z(n14025) );
  XOR2_X1 U33665 ( .A1(n23283), .A2(n53641), .Z(n14027) );
  NAND2_X1 U33667 ( .A1(n22764), .A2(n59200), .ZN(n49733) );
  NAND2_X1 U33668 ( .A1(n49730), .A2(n59200), .ZN(n24680) );
  NOR2_X1 U33672 ( .A1(n50296), .A2(n50309), .ZN(n14047) );
  INV_X2 U33674 ( .I(n14049), .ZN(n25876) );
  XOR2_X1 U33675 ( .A1(n63041), .A2(n51652), .Z(n14052) );
  NAND2_X1 U33678 ( .A1(n1158), .A2(n7159), .ZN(n49820) );
  OAI21_X1 U33679 ( .A1(n14375), .A2(n17372), .B(n7159), .ZN(n14374) );
  XOR2_X1 U33680 ( .A1(n672), .A2(n45315), .Z(n45393) );
  INV_X1 U33681 ( .I(n14056), .ZN(n20850) );
  NAND2_X1 U33682 ( .A1(n14056), .A2(n101), .ZN(n52123) );
  NOR2_X1 U33683 ( .A1(n55425), .A2(n14056), .ZN(n15485) );
  NOR2_X2 U33684 ( .A1(n39090), .A2(n14060), .ZN(n44627) );
  MUX2_X1 U33687 ( .I0(n47666), .I1(n47665), .S(n2640), .Z(n24396) );
  XOR2_X1 U33690 ( .A1(n14075), .A2(n14076), .Z(n14074) );
  XOR2_X1 U33691 ( .A1(n14441), .A2(n64142), .Z(n14075) );
  XOR2_X1 U33692 ( .A1(n14079), .A2(n16969), .Z(n14076) );
  INV_X2 U33693 ( .I(n14077), .ZN(n26041) );
  XOR2_X1 U33694 ( .A1(n14967), .A2(n14440), .Z(n14079) );
  NAND2_X2 U33695 ( .A1(n14084), .A2(n14083), .ZN(n24864) );
  XOR2_X1 U33697 ( .A1(n8179), .A2(n14089), .Z(n14088) );
  NAND3_X1 U33698 ( .A1(n53701), .A2(n53699), .A3(n53700), .ZN(n14090) );
  XOR2_X1 U33702 ( .A1(n52603), .A2(n17504), .Z(n14095) );
  INV_X2 U33704 ( .I(n25171), .ZN(n22362) );
  NOR2_X2 U33705 ( .A1(n14101), .A2(n14100), .ZN(n25171) );
  AOI22_X1 U33707 ( .A1(n32297), .A2(n18077), .B1(n34569), .B2(n7797), .ZN(
        n32300) );
  XOR2_X1 U33709 ( .A1(n14106), .A2(n25005), .Z(n22429) );
  NAND2_X1 U33710 ( .A1(n34652), .A2(n14107), .ZN(n34655) );
  XOR2_X1 U33713 ( .A1(n24656), .A2(n32343), .Z(n35001) );
  AOI21_X1 U33714 ( .A1(n14115), .A2(n9792), .B(n17848), .ZN(n14114) );
  NOR2_X2 U33716 ( .A1(n63666), .A2(n42785), .ZN(n17371) );
  NAND2_X2 U33717 ( .A1(n17848), .A2(n41660), .ZN(n43027) );
  NOR2_X1 U33718 ( .A1(n43318), .A2(n19428), .ZN(n14118) );
  NAND2_X2 U33720 ( .A1(n14136), .A2(n21010), .ZN(n15488) );
  XOR2_X1 U33721 ( .A1(n14144), .A2(n14143), .Z(n14145) );
  INV_X2 U33723 ( .I(n14145), .ZN(n38990) );
  XOR2_X1 U33724 ( .A1(n39213), .A2(n38990), .Z(n38991) );
  XOR2_X1 U33726 ( .A1(Ciphertext[65]), .A2(Key[156]), .Z(n17904) );
  XOR2_X1 U33728 ( .A1(n14154), .A2(n61662), .Z(n14153) );
  XOR2_X1 U33730 ( .A1(n18133), .A2(n1018), .Z(n14155) );
  XOR2_X1 U33733 ( .A1(n14158), .A2(n39765), .Z(n14157) );
  XOR2_X1 U33736 ( .A1(n14160), .A2(n38253), .Z(n25407) );
  XOR2_X1 U33737 ( .A1(Ciphertext[52]), .A2(Key[161]), .Z(n24989) );
  XOR2_X1 U33738 ( .A1(n14162), .A2(n22188), .Z(n23254) );
  NAND2_X1 U33740 ( .A1(n49357), .A2(n14167), .ZN(n14166) );
  NOR2_X1 U33741 ( .A1(n14169), .A2(n14168), .ZN(n14167) );
  AOI21_X1 U33742 ( .A1(n50043), .A2(n3348), .B(n1637), .ZN(n14169) );
  XOR2_X1 U33746 ( .A1(n20972), .A2(n50324), .Z(n14181) );
  XOR2_X1 U33748 ( .A1(n14187), .A2(n14186), .Z(n22918) );
  XOR2_X1 U33749 ( .A1(n16559), .A2(n15458), .Z(n14186) );
  OR2_X1 U33751 ( .A1(n14627), .A2(n14628), .Z(n14881) );
  XOR2_X1 U33752 ( .A1(n14188), .A2(n15579), .Z(n17712) );
  INV_X1 U33753 ( .I(n22435), .ZN(n14188) );
  NOR2_X1 U33755 ( .A1(n49465), .A2(n57608), .ZN(n49751) );
  NOR2_X1 U33757 ( .A1(n36743), .A2(n14189), .ZN(n36744) );
  NOR2_X2 U33764 ( .A1(n14630), .A2(n14199), .ZN(n45964) );
  NAND3_X1 U33765 ( .A1(n27799), .A2(n27798), .A3(n14200), .ZN(n25095) );
  NAND2_X1 U33766 ( .A1(n28952), .A2(n14202), .ZN(n14201) );
  NAND3_X2 U33770 ( .A1(n49523), .A2(n14208), .A3(n14207), .ZN(n14206) );
  NAND2_X2 U33771 ( .A1(n27690), .A2(n20627), .ZN(n14212) );
  NAND2_X1 U33774 ( .A1(n29918), .A2(n14213), .ZN(n17714) );
  NAND2_X2 U33775 ( .A1(n29916), .A2(n31129), .ZN(n14213) );
  NAND3_X2 U33776 ( .A1(n32466), .A2(n14219), .A3(n32465), .ZN(n18348) );
  XOR2_X1 U33780 ( .A1(n10896), .A2(n57226), .Z(n51619) );
  NOR2_X1 U33782 ( .A1(n14225), .A2(n14226), .ZN(n55435) );
  NOR2_X1 U33784 ( .A1(n55317), .A2(n14226), .ZN(n21393) );
  OAI21_X1 U33785 ( .A1(n52492), .A2(n14225), .B(n14226), .ZN(n52494) );
  XOR2_X1 U33786 ( .A1(n14228), .A2(n50984), .Z(n37682) );
  XOR2_X1 U33787 ( .A1(n14228), .A2(n778), .Z(n15955) );
  AOI21_X1 U33791 ( .A1(n3971), .A2(n2810), .B(n13554), .ZN(n49061) );
  NAND2_X2 U33794 ( .A1(n36139), .A2(n1422), .ZN(n35396) );
  INV_X2 U33795 ( .I(n60930), .ZN(n42605) );
  NAND2_X1 U33800 ( .A1(n20787), .A2(n21803), .ZN(n14236) );
  XOR2_X1 U33802 ( .A1(n38300), .A2(n14238), .Z(n20022) );
  XOR2_X1 U33803 ( .A1(n61944), .A2(n16313), .Z(n14238) );
  XOR2_X1 U33807 ( .A1(n14252), .A2(n43593), .Z(n43594) );
  XOR2_X1 U33808 ( .A1(n14251), .A2(n20772), .Z(n14252) );
  XOR2_X1 U33809 ( .A1(n14253), .A2(n46207), .Z(n46209) );
  XOR2_X1 U33810 ( .A1(n14253), .A2(n43671), .Z(n43672) );
  XOR2_X1 U33811 ( .A1(n14760), .A2(n58740), .Z(n18711) );
  NAND2_X1 U33813 ( .A1(n49947), .A2(n14254), .ZN(n48741) );
  OAI22_X1 U33814 ( .A1(n27938), .A2(n27937), .B1(n1359), .B2(n14258), .ZN(
        n14257) );
  XOR2_X1 U33815 ( .A1(n21369), .A2(n31864), .Z(n32405) );
  XOR2_X1 U33817 ( .A1(n14259), .A2(n784), .Z(n16106) );
  INV_X1 U33818 ( .I(n43087), .ZN(n43096) );
  NAND3_X2 U33821 ( .A1(n31101), .A2(n30579), .A3(n60327), .ZN(n31113) );
  INV_X2 U33822 ( .I(n42217), .ZN(n14278) );
  NOR2_X2 U33823 ( .A1(n14280), .A2(n14279), .ZN(n42217) );
  XOR2_X1 U33828 ( .A1(n19433), .A2(n45245), .Z(n14284) );
  AOI21_X1 U33830 ( .A1(n47882), .A2(n14289), .B(n11899), .ZN(n47724) );
  XOR2_X1 U33833 ( .A1(n6904), .A2(n14295), .Z(n14293) );
  XOR2_X1 U33834 ( .A1(n17986), .A2(n33152), .Z(n14296) );
  NOR2_X1 U33836 ( .A1(n14300), .A2(n20426), .ZN(n45487) );
  XOR2_X1 U33838 ( .A1(n51828), .A2(n19519), .Z(n51762) );
  NOR2_X1 U33839 ( .A1(n42893), .A2(n14305), .ZN(n42888) );
  XOR2_X1 U33842 ( .A1(n24314), .A2(n51161), .Z(n14977) );
  XOR2_X1 U33845 ( .A1(n5767), .A2(n1489), .Z(n44371) );
  INV_X2 U33847 ( .I(n5767), .ZN(n17102) );
  XOR2_X1 U33850 ( .A1(n60466), .A2(n53375), .Z(n31438) );
  INV_X2 U33852 ( .I(n53518), .ZN(n17225) );
  NOR2_X1 U33853 ( .A1(n14324), .A2(n22977), .ZN(n55921) );
  NAND2_X1 U33854 ( .A1(n11524), .A2(n1370), .ZN(n14325) );
  NAND3_X1 U33855 ( .A1(n1338), .A2(n36956), .A3(n60694), .ZN(n36273) );
  NOR2_X1 U33859 ( .A1(n14334), .A2(n31098), .ZN(n30577) );
  INV_X1 U33861 ( .I(n44759), .ZN(n14339) );
  NOR2_X1 U33862 ( .A1(n29785), .A2(n29784), .ZN(n29789) );
  NOR2_X2 U33863 ( .A1(n1871), .A2(n58710), .ZN(n29246) );
  INV_X2 U33864 ( .I(n15242), .ZN(n15783) );
  INV_X2 U33866 ( .I(n13719), .ZN(n47576) );
  AOI21_X2 U33867 ( .A1(n14857), .A2(n59694), .B(n14856), .ZN(n18624) );
  XOR2_X1 U33870 ( .A1(n30985), .A2(n32266), .Z(n14345) );
  INV_X1 U33875 ( .I(n14352), .ZN(n55735) );
  NAND2_X1 U33877 ( .A1(n6531), .A2(n61247), .ZN(n14351) );
  OAI22_X1 U33878 ( .A1(n52926), .A2(n52927), .B1(n52925), .B2(n14352), .ZN(
        n52928) );
  NAND2_X2 U33879 ( .A1(n2180), .A2(n52211), .ZN(n14352) );
  NAND2_X1 U33887 ( .A1(n14358), .A2(n62768), .ZN(n25446) );
  NOR2_X1 U33888 ( .A1(n14358), .A2(n23849), .ZN(n54817) );
  NAND2_X1 U33889 ( .A1(n19137), .A2(n14358), .ZN(n54691) );
  NOR2_X1 U33890 ( .A1(n14358), .A2(n62768), .ZN(n14357) );
  NOR2_X2 U33892 ( .A1(n23554), .A2(n58828), .ZN(n14360) );
  NAND2_X2 U33893 ( .A1(n14361), .A2(n21487), .ZN(n35827) );
  XOR2_X1 U33899 ( .A1(n14373), .A2(n45138), .Z(n45139) );
  XOR2_X1 U33900 ( .A1(n14379), .A2(n19959), .Z(n14378) );
  XOR2_X1 U33901 ( .A1(n32184), .A2(n25314), .Z(n14379) );
  XOR2_X1 U33902 ( .A1(n30936), .A2(n31768), .Z(n14380) );
  XOR2_X1 U33904 ( .A1(n21688), .A2(n12669), .Z(n14382) );
  NAND3_X2 U33905 ( .A1(n14395), .A2(n14388), .A3(n14387), .ZN(n32543) );
  INV_X1 U33909 ( .I(n63389), .ZN(n48455) );
  AOI21_X2 U33910 ( .A1(n15475), .A2(n25459), .B(n14403), .ZN(n14402) );
  OAI21_X2 U33911 ( .A1(n49010), .A2(n25459), .B(n15474), .ZN(n14403) );
  NOR2_X2 U33912 ( .A1(n48323), .A2(n23738), .ZN(n49010) );
  NAND2_X1 U33915 ( .A1(n25481), .A2(n14419), .ZN(n46357) );
  AOI21_X1 U33916 ( .A1(n31084), .A2(n31083), .B(n31082), .ZN(n14421) );
  XOR2_X1 U33918 ( .A1(n50625), .A2(n50624), .Z(n14425) );
  INV_X2 U33920 ( .I(n44639), .ZN(n46299) );
  XOR2_X1 U33921 ( .A1(n20413), .A2(n14426), .Z(n25602) );
  XOR2_X1 U33922 ( .A1(n14427), .A2(n44639), .Z(n14426) );
  NAND3_X2 U33923 ( .A1(n42960), .A2(n44237), .A3(n42959), .ZN(n44639) );
  INV_X2 U33925 ( .I(n55356), .ZN(n55389) );
  NAND2_X2 U33926 ( .A1(n14429), .A2(n24673), .ZN(n55356) );
  INV_X2 U33928 ( .I(n29282), .ZN(n18062) );
  INV_X1 U33930 ( .I(n14433), .ZN(n29624) );
  INV_X1 U33931 ( .I(n26948), .ZN(n28837) );
  NOR2_X1 U33933 ( .A1(n28127), .A2(n23549), .ZN(n14434) );
  INV_X2 U33934 ( .I(n24350), .ZN(n14439) );
  XOR2_X1 U33935 ( .A1(n24025), .A2(n848), .Z(n14440) );
  XOR2_X1 U33936 ( .A1(n38310), .A2(n38309), .Z(n14442) );
  XOR2_X1 U33937 ( .A1(n38531), .A2(n38313), .Z(n14443) );
  XOR2_X1 U33938 ( .A1(n46712), .A2(n46713), .Z(n14447) );
  XOR2_X1 U33940 ( .A1(n14449), .A2(n38823), .Z(n19956) );
  XOR2_X1 U33941 ( .A1(n1750), .A2(n922), .Z(n14449) );
  NOR2_X1 U33942 ( .A1(n1564), .A2(n16707), .ZN(n14450) );
  NAND2_X1 U33943 ( .A1(n26771), .A2(n522), .ZN(n26776) );
  NOR2_X2 U33944 ( .A1(n47843), .A2(n9860), .ZN(n47839) );
  NOR2_X2 U33946 ( .A1(n15520), .A2(n5051), .ZN(n55074) );
  XOR2_X1 U33947 ( .A1(n14459), .A2(n52326), .Z(n54615) );
  XOR2_X1 U33948 ( .A1(n8805), .A2(n14458), .Z(n52326) );
  NAND2_X2 U33952 ( .A1(n28717), .A2(n21887), .ZN(n30781) );
  INV_X1 U33953 ( .I(n32295), .ZN(n34564) );
  NAND2_X1 U33954 ( .A1(n32295), .A2(n21725), .ZN(n14464) );
  XOR2_X1 U33956 ( .A1(n14465), .A2(n17383), .Z(n14958) );
  XOR2_X1 U33957 ( .A1(n14466), .A2(n936), .Z(n14465) );
  INV_X1 U33959 ( .I(n20909), .ZN(n14471) );
  NOR2_X1 U33963 ( .A1(n58983), .A2(n49538), .ZN(n49539) );
  OR2_X1 U33968 ( .A1(n42476), .A2(n42479), .Z(n14478) );
  XOR2_X1 U33969 ( .A1(n14482), .A2(n14481), .Z(n14480) );
  XOR2_X1 U33970 ( .A1(n39216), .A2(n39215), .Z(n14481) );
  XOR2_X1 U33971 ( .A1(n22953), .A2(n39405), .Z(n14482) );
  AOI21_X1 U33972 ( .A1(n14484), .A2(n56919), .B(n64845), .ZN(n56911) );
  NOR2_X1 U33973 ( .A1(n17850), .A2(n14484), .ZN(n14560) );
  NAND2_X2 U33975 ( .A1(n7055), .A2(n55722), .ZN(n55908) );
  XOR2_X1 U33979 ( .A1(n14489), .A2(n54563), .Z(Plaintext[76]) );
  NAND3_X1 U33980 ( .A1(n14493), .A2(n14492), .A3(n14490), .ZN(n14489) );
  INV_X1 U33981 ( .I(n54562), .ZN(n14492) );
  AOI22_X1 U33982 ( .A1(n54559), .A2(n1174), .B1(n14551), .B2(n54579), .ZN(
        n14493) );
  INV_X2 U33983 ( .I(n26184), .ZN(n29317) );
  NAND2_X2 U33984 ( .A1(n14496), .A2(n14498), .ZN(n43302) );
  AND2_X1 U33987 ( .A1(n28554), .A2(n14502), .Z(n16751) );
  NAND3_X1 U33988 ( .A1(n28553), .A2(n19328), .A3(n29178), .ZN(n14502) );
  NOR2_X1 U33989 ( .A1(n14504), .A2(n24419), .ZN(n14503) );
  NAND2_X2 U33990 ( .A1(n23608), .A2(n22352), .ZN(n28548) );
  INV_X2 U33992 ( .I(n27125), .ZN(n27142) );
  NOR2_X2 U33993 ( .A1(n64903), .A2(n28048), .ZN(n27125) );
  XOR2_X1 U33994 ( .A1(Ciphertext[36]), .A2(Key[49]), .Z(n26278) );
  AND2_X1 U33996 ( .A1(n28780), .A2(n28779), .Z(n14523) );
  OAI21_X1 U33997 ( .A1(n25304), .A2(n25305), .B(n14524), .ZN(n18137) );
  XOR2_X1 U34000 ( .A1(n14528), .A2(n14527), .Z(n14530) );
  XOR2_X1 U34001 ( .A1(n25582), .A2(n14824), .Z(n14527) );
  INV_X2 U34003 ( .I(n14530), .ZN(n15871) );
  INV_X2 U34004 ( .I(n30292), .ZN(n29575) );
  NAND3_X2 U34005 ( .A1(n14532), .A2(n24898), .A3(n24897), .ZN(n30292) );
  NAND2_X2 U34008 ( .A1(n15540), .A2(n18724), .ZN(n17755) );
  OR2_X1 U34010 ( .A1(n14881), .A2(n42983), .Z(n14536) );
  OAI21_X2 U34012 ( .A1(n48881), .A2(n22320), .B(n48880), .ZN(n52360) );
  XOR2_X1 U34014 ( .A1(n32744), .A2(n1834), .Z(n23667) );
  XOR2_X1 U34016 ( .A1(n17204), .A2(n23611), .Z(n53433) );
  XOR2_X1 U34018 ( .A1(n38794), .A2(n38793), .Z(n39209) );
  XOR2_X1 U34022 ( .A1(n15102), .A2(n32367), .Z(n15188) );
  AOI21_X1 U34023 ( .A1(n52217), .A2(n55927), .B(n55920), .ZN(n14539) );
  NAND2_X1 U34024 ( .A1(n55926), .A2(n14541), .ZN(n52219) );
  INV_X1 U34025 ( .I(n28694), .ZN(n14544) );
  INV_X1 U34026 ( .I(n14546), .ZN(n14545) );
  NAND2_X1 U34029 ( .A1(n14552), .A2(n54575), .ZN(n14551) );
  XOR2_X1 U34031 ( .A1(n63011), .A2(n828), .Z(n36993) );
  INV_X1 U34033 ( .I(n40136), .ZN(n14556) );
  NOR2_X2 U34038 ( .A1(n1583), .A2(n1257), .ZN(n56936) );
  NAND2_X1 U34039 ( .A1(n19435), .A2(n34155), .ZN(n31608) );
  AOI22_X1 U34041 ( .A1(n17759), .A2(n34151), .B1(n34150), .B2(n19435), .ZN(
        n19986) );
  INV_X2 U34042 ( .I(n16590), .ZN(n48421) );
  NAND2_X1 U34045 ( .A1(n14565), .A2(n14564), .ZN(n19070) );
  OR2_X1 U34046 ( .A1(n30584), .A2(n30583), .Z(n14564) );
  XOR2_X1 U34047 ( .A1(n32352), .A2(n14563), .Z(n32353) );
  XOR2_X1 U34048 ( .A1(n22781), .A2(n14563), .Z(n32280) );
  NOR2_X2 U34049 ( .A1(n14570), .A2(n14566), .ZN(n15741) );
  NOR2_X2 U34050 ( .A1(n14578), .A2(n14576), .ZN(n14709) );
  NOR2_X1 U34051 ( .A1(n14583), .A2(n28031), .ZN(n14582) );
  XOR2_X1 U34053 ( .A1(Ciphertext[43]), .A2(Key[2]), .Z(n14774) );
  XOR2_X1 U34055 ( .A1(n24184), .A2(n14587), .Z(n14586) );
  XOR2_X1 U34056 ( .A1(n60062), .A2(n17533), .Z(n14587) );
  XOR2_X1 U34057 ( .A1(n23174), .A2(n14590), .Z(n14589) );
  XOR2_X1 U34060 ( .A1(n52621), .A2(n354), .Z(n14593) );
  XOR2_X1 U34061 ( .A1(n51490), .A2(n51489), .Z(n14594) );
  XOR2_X1 U34062 ( .A1(n14596), .A2(n14595), .Z(n14733) );
  XOR2_X1 U34064 ( .A1(n5200), .A2(n24169), .Z(n35075) );
  XOR2_X1 U34065 ( .A1(n5200), .A2(n39755), .Z(n39655) );
  NAND2_X2 U34066 ( .A1(n47167), .A2(n47166), .ZN(n48616) );
  XOR2_X1 U34070 ( .A1(n51792), .A2(n51179), .Z(n14607) );
  XOR2_X1 U34071 ( .A1(n51181), .A2(n51178), .Z(n14608) );
  XOR2_X1 U34072 ( .A1(n14610), .A2(n24076), .Z(n51181) );
  XOR2_X1 U34073 ( .A1(n23375), .A2(n16984), .Z(n14609) );
  XOR2_X1 U34074 ( .A1(n46288), .A2(n46287), .Z(n46289) );
  XOR2_X1 U34075 ( .A1(n65170), .A2(n46288), .Z(n25697) );
  INV_X2 U34076 ( .I(n14612), .ZN(n20897) );
  OAI22_X1 U34077 ( .A1(n17212), .A2(n39994), .B1(n14616), .B2(n41122), .ZN(
        n39997) );
  NOR2_X1 U34078 ( .A1(n39819), .A2(n14616), .ZN(n39820) );
  XOR2_X1 U34079 ( .A1(n46549), .A2(n45106), .Z(n45107) );
  NOR2_X1 U34081 ( .A1(n14619), .A2(n63784), .ZN(n57091) );
  AOI21_X1 U34082 ( .A1(n25146), .A2(n14619), .B(n19054), .ZN(n25145) );
  NAND2_X2 U34083 ( .A1(n21570), .A2(n21569), .ZN(n14619) );
  INV_X2 U34085 ( .I(n14620), .ZN(n23561) );
  INV_X2 U34093 ( .I(n23474), .ZN(n16523) );
  NOR2_X2 U34094 ( .A1(n27233), .A2(n20519), .ZN(n14633) );
  NOR3_X1 U34097 ( .A1(n57278), .A2(n36794), .A3(n36808), .ZN(n15946) );
  INV_X2 U34098 ( .I(n14639), .ZN(n15074) );
  XOR2_X1 U34100 ( .A1(n12356), .A2(n1573), .Z(n16038) );
  XOR2_X1 U34103 ( .A1(n23668), .A2(n23440), .Z(n14640) );
  NAND3_X2 U34104 ( .A1(n14644), .A2(n18655), .A3(n22915), .ZN(n18652) );
  XOR2_X1 U34106 ( .A1(n39481), .A2(n25911), .Z(n14646) );
  INV_X2 U34107 ( .I(n21495), .ZN(n45437) );
  INV_X2 U34108 ( .I(n16666), .ZN(n20902) );
  NAND2_X1 U34110 ( .A1(n57026), .A2(n53212), .ZN(n16767) );
  NAND2_X1 U34117 ( .A1(n2489), .A2(n5140), .ZN(n14661) );
  INV_X2 U34118 ( .I(n14662), .ZN(n41078) );
  XOR2_X1 U34119 ( .A1(n1239), .A2(n39731), .Z(n14663) );
  CLKBUF_X4 U34120 ( .I(n15714), .Z(n14666) );
  XOR2_X1 U34121 ( .A1(n24827), .A2(n31335), .Z(n21988) );
  XOR2_X1 U34122 ( .A1(n31556), .A2(n15714), .Z(n31335) );
  NAND3_X2 U34123 ( .A1(n30306), .A2(n21312), .A3(n30307), .ZN(n15714) );
  AOI22_X2 U34126 ( .A1(n15277), .A2(n14991), .B1(n45041), .B2(n60486), .ZN(
        n25432) );
  XOR2_X1 U34128 ( .A1(n2666), .A2(n17728), .Z(n17727) );
  XOR2_X1 U34130 ( .A1(n46212), .A2(n46214), .Z(n14674) );
  XOR2_X1 U34131 ( .A1(n23807), .A2(n46215), .Z(n14675) );
  XOR2_X1 U34133 ( .A1(n37527), .A2(n37793), .Z(n14682) );
  XOR2_X1 U34134 ( .A1(n37625), .A2(n39687), .Z(n15932) );
  NAND3_X1 U34135 ( .A1(n36424), .A2(n36422), .A3(n36423), .ZN(n14686) );
  NAND2_X2 U34137 ( .A1(n14692), .A2(n14689), .ZN(n15708) );
  NOR2_X2 U34138 ( .A1(n48213), .A2(n48204), .ZN(n47492) );
  XOR2_X1 U34139 ( .A1(n16511), .A2(n14696), .Z(n17320) );
  NOR2_X1 U34145 ( .A1(n34658), .A2(n5411), .ZN(n14702) );
  NOR3_X1 U34146 ( .A1(n14954), .A2(n34165), .A3(n14703), .ZN(n14953) );
  NOR2_X1 U34148 ( .A1(n39146), .A2(n11787), .ZN(n39040) );
  NOR2_X2 U34150 ( .A1(n23942), .A2(n14705), .ZN(n26531) );
  XOR2_X1 U34151 ( .A1(n38455), .A2(n38500), .Z(n14706) );
  XOR2_X1 U34152 ( .A1(n24753), .A2(n37525), .Z(n38458) );
  XOR2_X1 U34153 ( .A1(n38456), .A2(n38452), .Z(n14707) );
  NAND3_X2 U34154 ( .A1(n15624), .A2(n15623), .A3(n30101), .ZN(n18434) );
  INV_X2 U34155 ( .I(n52287), .ZN(n56961) );
  NAND2_X2 U34158 ( .A1(n14710), .A2(n52240), .ZN(n56965) );
  XNOR2_X1 U34159 ( .A1(n14716), .A2(n14715), .ZN(n14714) );
  INV_X2 U34160 ( .I(n14717), .ZN(n22953) );
  XNOR2_X1 U34161 ( .A1(n38325), .A2(n38510), .ZN(n14717) );
  NAND2_X2 U34162 ( .A1(n23681), .A2(n34112), .ZN(n38325) );
  NAND2_X1 U34163 ( .A1(n25050), .A2(n34204), .ZN(n14719) );
  XOR2_X1 U34166 ( .A1(n61410), .A2(n45394), .Z(n14807) );
  XOR2_X1 U34168 ( .A1(n50638), .A2(n14730), .Z(n50639) );
  NOR2_X1 U34171 ( .A1(n58651), .A2(n30441), .ZN(n30438) );
  NOR3_X1 U34173 ( .A1(n30439), .A2(n30537), .A3(n58651), .ZN(n30436) );
  XOR2_X1 U34175 ( .A1(n14736), .A2(n44273), .Z(n14735) );
  XOR2_X1 U34176 ( .A1(n18624), .A2(n24173), .Z(n14736) );
  XOR2_X1 U34177 ( .A1(n14737), .A2(n37723), .Z(n20291) );
  XOR2_X1 U34179 ( .A1(n37682), .A2(n58725), .Z(n20191) );
  NAND2_X1 U34181 ( .A1(n14739), .A2(n30537), .ZN(n29979) );
  OAI22_X1 U34182 ( .A1(n28092), .A2(n30439), .B1(n16694), .B2(n14739), .ZN(
        n16695) );
  AOI21_X1 U34184 ( .A1(n35953), .A2(n14743), .B(n26125), .ZN(n26124) );
  NAND2_X1 U34186 ( .A1(n28098), .A2(n29000), .ZN(n14744) );
  NAND2_X1 U34187 ( .A1(n28097), .A2(n28096), .ZN(n14746) );
  XOR2_X1 U34188 ( .A1(n14748), .A2(n14747), .Z(n48097) );
  XOR2_X1 U34190 ( .A1(n45246), .A2(n802), .Z(n45353) );
  XOR2_X1 U34191 ( .A1(n324), .A2(n14751), .Z(n21762) );
  XOR2_X1 U34192 ( .A1(n12377), .A2(n22994), .Z(n17898) );
  NAND2_X2 U34193 ( .A1(n13672), .A2(n19522), .ZN(n27615) );
  NAND2_X2 U34196 ( .A1(n27241), .A2(n27240), .ZN(n20809) );
  XOR2_X1 U34197 ( .A1(n18468), .A2(n46522), .Z(n46527) );
  XOR2_X1 U34198 ( .A1(n14760), .A2(n46650), .Z(n21896) );
  NAND2_X2 U34199 ( .A1(n18144), .A2(n36057), .ZN(n14763) );
  NAND2_X2 U34203 ( .A1(n1518), .A2(n14773), .ZN(n40238) );
  XOR2_X1 U34205 ( .A1(n24621), .A2(n51388), .Z(n19810) );
  XOR2_X1 U34206 ( .A1(Ciphertext[134]), .A2(Key[159]), .Z(n29619) );
  INV_X1 U34207 ( .I(n49811), .ZN(n17549) );
  NOR2_X1 U34208 ( .A1(n14778), .A2(n63784), .ZN(n21437) );
  NOR2_X1 U34209 ( .A1(n14778), .A2(n21829), .ZN(n57099) );
  OAI21_X1 U34210 ( .A1(n14778), .A2(n57156), .B(n57433), .ZN(n57086) );
  NAND2_X1 U34213 ( .A1(n57136), .A2(n14778), .ZN(n57137) );
  AOI21_X1 U34214 ( .A1(n57154), .A2(n14778), .B(n57153), .ZN(n57155) );
  INV_X4 U34215 ( .I(n21570), .ZN(n14778) );
  NAND2_X2 U34216 ( .A1(n28400), .A2(n3117), .ZN(n28406) );
  XOR2_X1 U34217 ( .A1(n14783), .A2(n14251), .Z(n45815) );
  NAND3_X1 U34218 ( .A1(n33518), .A2(n35024), .A3(n20785), .ZN(n14792) );
  XOR2_X1 U34219 ( .A1(n246), .A2(n50954), .Z(n14793) );
  XOR2_X1 U34220 ( .A1(n63026), .A2(n50715), .Z(n14794) );
  XOR2_X1 U34222 ( .A1(n5555), .A2(n63000), .Z(n38083) );
  AOI21_X1 U34225 ( .A1(n38762), .A2(n41478), .B(n38761), .ZN(n14801) );
  AND2_X1 U34226 ( .A1(n15132), .A2(n62261), .Z(n14804) );
  XOR2_X1 U34228 ( .A1(n61490), .A2(n45402), .Z(n46666) );
  XOR2_X1 U34229 ( .A1(n44966), .A2(n10745), .Z(n45394) );
  XOR2_X1 U34230 ( .A1(n18156), .A2(n14808), .Z(n32738) );
  NOR2_X1 U34231 ( .A1(n61835), .A2(n14809), .ZN(n48382) );
  OR2_X1 U34235 ( .A1(n1001), .A2(n22713), .Z(n14816) );
  XOR2_X1 U34236 ( .A1(n14818), .A2(n32034), .Z(n19960) );
  XOR2_X1 U34237 ( .A1(n14818), .A2(n13181), .Z(n20715) );
  NOR2_X2 U34239 ( .A1(n15892), .A2(n57459), .ZN(n18208) );
  XOR2_X1 U34241 ( .A1(n14826), .A2(n14824), .Z(n14825) );
  INV_X1 U34245 ( .I(n56099), .ZN(n14837) );
  XOR2_X1 U34247 ( .A1(n58310), .A2(n20224), .Z(n20223) );
  XOR2_X1 U34248 ( .A1(n14839), .A2(n50831), .Z(Plaintext[38]) );
  INV_X2 U34250 ( .I(n53727), .ZN(n25117) );
  NAND2_X2 U34251 ( .A1(n21999), .A2(n21996), .ZN(n53727) );
  NOR2_X1 U34253 ( .A1(n22385), .A2(n63473), .ZN(n54766) );
  XOR2_X1 U34256 ( .A1(n14855), .A2(n46525), .Z(n46526) );
  XOR2_X1 U34258 ( .A1(n14855), .A2(n16518), .Z(n46140) );
  XOR2_X1 U34259 ( .A1(n21984), .A2(n14862), .Z(n14861) );
  XOR2_X1 U34265 ( .A1(n33840), .A2(n14866), .Z(n21563) );
  OAI22_X1 U34268 ( .A1(n27229), .A2(n27483), .B1(n27485), .B2(n14869), .ZN(
        n27226) );
  XOR2_X1 U34271 ( .A1(n52092), .A2(n25192), .Z(n52093) );
  XOR2_X1 U34273 ( .A1(n25623), .A2(n37649), .Z(n24148) );
  NOR2_X2 U34274 ( .A1(n20944), .A2(n22896), .ZN(n25623) );
  INV_X1 U34275 ( .I(n14875), .ZN(n47474) );
  NOR2_X1 U34276 ( .A1(n14875), .A2(n46979), .ZN(n46981) );
  MUX2_X1 U34277 ( .I0(n3368), .I1(n45517), .S(n14875), .Z(n44070) );
  MUX2_X1 U34278 ( .I0(n65224), .I1(n47473), .S(n14875), .Z(n45745) );
  NAND3_X1 U34279 ( .A1(n45523), .A2(n45522), .A3(n14875), .ZN(n45525) );
  AOI21_X1 U34280 ( .A1(n44685), .A2(n44686), .B(n14875), .ZN(n44687) );
  XNOR2_X1 U34282 ( .A1(Ciphertext[23]), .A2(Key[54]), .ZN(n14876) );
  OAI21_X1 U34289 ( .A1(n27219), .A2(n63883), .B(n14887), .ZN(n27220) );
  XNOR2_X1 U34291 ( .A1(n45152), .A2(n14889), .ZN(n14888) );
  INV_X1 U34292 ( .I(n55826), .ZN(n20710) );
  NAND2_X1 U34293 ( .A1(n37399), .A2(n36160), .ZN(n14895) );
  NAND2_X2 U34296 ( .A1(n45835), .A2(n45836), .ZN(n43909) );
  XNOR2_X1 U34298 ( .A1(Ciphertext[10]), .A2(Key[59]), .ZN(n14903) );
  NAND2_X2 U34303 ( .A1(n1856), .A2(n1868), .ZN(n14921) );
  NOR2_X1 U34304 ( .A1(n14927), .A2(n55316), .ZN(n55320) );
  NAND3_X1 U34305 ( .A1(n55321), .A2(n14927), .A3(n55440), .ZN(n52955) );
  NOR2_X2 U34308 ( .A1(n55433), .A2(n55306), .ZN(n14927) );
  NAND2_X2 U34314 ( .A1(n14943), .A2(n56539), .ZN(n16329) );
  NAND3_X1 U34315 ( .A1(n56534), .A2(n22870), .A3(n14943), .ZN(n56384) );
  NAND2_X1 U34317 ( .A1(n63589), .A2(n14944), .ZN(n26305) );
  INV_X2 U34322 ( .I(n16021), .ZN(n28346) );
  NOR2_X2 U34323 ( .A1(n27524), .A2(n1894), .ZN(n16021) );
  INV_X2 U34324 ( .I(n14958), .ZN(n17382) );
  NOR2_X1 U34330 ( .A1(n14965), .A2(n41072), .ZN(n41075) );
  OR2_X1 U34331 ( .A1(n40849), .A2(n14965), .Z(n39967) );
  XOR2_X1 U34334 ( .A1(n60964), .A2(n824), .Z(n18446) );
  XOR2_X1 U34336 ( .A1(n12985), .A2(n14974), .Z(n50541) );
  XOR2_X1 U34337 ( .A1(n51552), .A2(n14974), .Z(n52195) );
  XOR2_X1 U34338 ( .A1(n51672), .A2(n14974), .Z(n51673) );
  XOR2_X1 U34339 ( .A1(n52597), .A2(n14974), .Z(n52598) );
  XOR2_X1 U34340 ( .A1(n51327), .A2(n14974), .Z(n51328) );
  XOR2_X1 U34344 ( .A1(n14981), .A2(n31590), .Z(n30987) );
  XOR2_X1 U34345 ( .A1(n14981), .A2(n45123), .Z(n33193) );
  XOR2_X1 U34346 ( .A1(n14981), .A2(n22472), .Z(n30733) );
  XOR2_X1 U34350 ( .A1(n61571), .A2(n14993), .Z(n50980) );
  NAND2_X1 U34356 ( .A1(n53368), .A2(n23874), .ZN(n53348) );
  NOR2_X2 U34357 ( .A1(n40850), .A2(n64459), .ZN(n40857) );
  NAND2_X2 U34359 ( .A1(n15000), .A2(n56238), .ZN(n18096) );
  INV_X2 U34360 ( .I(n52285), .ZN(n15000) );
  XOR2_X1 U34365 ( .A1(n1411), .A2(n49088), .Z(n15003) );
  AND2_X1 U34366 ( .A1(n50294), .A2(n3054), .Z(n15006) );
  OR2_X1 U34369 ( .A1(n36227), .A2(n36228), .Z(n15010) );
  NOR2_X2 U34370 ( .A1(n33297), .A2(n15012), .ZN(n36517) );
  XOR2_X1 U34371 ( .A1(n59218), .A2(n43390), .Z(n23239) );
  XOR2_X1 U34372 ( .A1(n15015), .A2(n23828), .Z(n43390) );
  XOR2_X1 U34374 ( .A1(n31849), .A2(n15017), .Z(n15016) );
  XOR2_X1 U34377 ( .A1(n15022), .A2(n52413), .Z(n51362) );
  XOR2_X1 U34378 ( .A1(n51361), .A2(n23628), .Z(n15022) );
  NAND3_X1 U34379 ( .A1(n2699), .A2(n25671), .A3(n14138), .ZN(n35488) );
  NOR2_X1 U34380 ( .A1(n20431), .A2(n14138), .ZN(n20433) );
  NAND2_X1 U34389 ( .A1(n1227), .A2(n15045), .ZN(n18538) );
  NOR2_X2 U34391 ( .A1(n29128), .A2(n10399), .ZN(n27406) );
  INV_X2 U34392 ( .I(n15046), .ZN(n32425) );
  XOR2_X1 U34397 ( .A1(n46344), .A2(n15054), .Z(n15053) );
  NOR2_X1 U34400 ( .A1(n53180), .A2(n15059), .ZN(n52750) );
  XNOR2_X1 U34403 ( .A1(n15262), .A2(n15260), .ZN(n15060) );
  NAND2_X1 U34409 ( .A1(n34067), .A2(n15085), .ZN(n34076) );
  AOI21_X1 U34410 ( .A1(n34511), .A2(n15085), .B(n34510), .ZN(n34515) );
  NOR2_X1 U34411 ( .A1(n24875), .A2(n15086), .ZN(n24874) );
  AND2_X1 U34412 ( .A1(n33486), .A2(n15085), .Z(n15086) );
  INV_X4 U34415 ( .I(n17661), .ZN(n20942) );
  NAND2_X1 U34418 ( .A1(n54543), .A2(n18063), .ZN(n54541) );
  OAI21_X2 U34419 ( .A1(n40952), .A2(n40949), .B(n58351), .ZN(n38045) );
  OAI21_X1 U34421 ( .A1(n22929), .A2(n24080), .B(n22928), .ZN(n15116) );
  NAND2_X2 U34422 ( .A1(n23895), .A2(n44013), .ZN(n23283) );
  OR2_X1 U34423 ( .A1(n20427), .A2(n15124), .Z(n49573) );
  AOI22_X1 U34424 ( .A1(n49360), .A2(n49441), .B1(n15124), .B2(n19773), .ZN(
        n49361) );
  XOR2_X1 U34427 ( .A1(n44092), .A2(n1682), .Z(n15125) );
  NAND2_X1 U34428 ( .A1(n15126), .A2(n15727), .ZN(n28287) );
  NAND2_X1 U34429 ( .A1(n15126), .A2(n11425), .ZN(n29423) );
  NOR2_X1 U34431 ( .A1(n30361), .A2(n3478), .ZN(n15433) );
  NAND2_X1 U34432 ( .A1(n15132), .A2(n51905), .ZN(n55706) );
  NAND2_X1 U34435 ( .A1(n55988), .A2(n15132), .ZN(n16621) );
  NAND2_X1 U34436 ( .A1(n55714), .A2(n15132), .ZN(n16331) );
  OAI22_X1 U34437 ( .A1(n55703), .A2(n15132), .B1(n56227), .B2(n55986), .ZN(
        n51906) );
  AOI22_X1 U34438 ( .A1(n55989), .A2(n15132), .B1(n64850), .B2(n55990), .ZN(
        n55991) );
  NOR2_X2 U34439 ( .A1(n1616), .A2(n56435), .ZN(n15132) );
  NAND2_X2 U34443 ( .A1(n15139), .A2(n20856), .ZN(n41109) );
  XOR2_X1 U34447 ( .A1(n22540), .A2(n50832), .Z(n31123) );
  XOR2_X1 U34448 ( .A1(n17463), .A2(n32578), .Z(n32580) );
  XOR2_X1 U34449 ( .A1(n17463), .A2(n33237), .Z(n33238) );
  XOR2_X1 U34450 ( .A1(n33168), .A2(n17463), .Z(n33169) );
  XOR2_X1 U34451 ( .A1(n22558), .A2(n17463), .Z(n32418) );
  NAND2_X2 U34454 ( .A1(n18651), .A2(n35283), .ZN(n15148) );
  XOR2_X1 U34456 ( .A1(n23152), .A2(n15153), .Z(n32049) );
  INV_X1 U34457 ( .I(n15156), .ZN(n28322) );
  NOR2_X1 U34458 ( .A1(n57872), .A2(n15156), .ZN(n27130) );
  NAND3_X1 U34459 ( .A1(n28320), .A2(n28321), .A3(n15156), .ZN(n26561) );
  NAND2_X1 U34460 ( .A1(n15157), .A2(n64944), .ZN(n47562) );
  NAND2_X1 U34461 ( .A1(n47664), .A2(n15157), .ZN(n47660) );
  MUX2_X1 U34462 ( .I0(n36741), .I1(n36742), .S(n17595), .Z(n36752) );
  NAND2_X2 U34466 ( .A1(n48533), .A2(n23331), .ZN(n21894) );
  INV_X2 U34468 ( .I(n24679), .ZN(n51911) );
  INV_X1 U34469 ( .I(n24508), .ZN(n19985) );
  XOR2_X1 U34470 ( .A1(n44480), .A2(n22731), .Z(n15173) );
  AOI21_X2 U34477 ( .A1(n15185), .A2(n34249), .B(n15182), .ZN(n34259) );
  XOR2_X1 U34479 ( .A1(n15188), .A2(n32494), .Z(n15187) );
  INV_X4 U34480 ( .I(n22963), .ZN(n29915) );
  NAND2_X2 U34481 ( .A1(n22964), .A2(n22965), .ZN(n22963) );
  INV_X2 U34482 ( .I(n15201), .ZN(n18524) );
  NAND2_X2 U34485 ( .A1(n15209), .A2(n15208), .ZN(n30547) );
  INV_X1 U34486 ( .I(n27269), .ZN(n15206) );
  INV_X1 U34488 ( .I(n19866), .ZN(n15213) );
  NAND2_X2 U34489 ( .A1(n15214), .A2(n23709), .ZN(n42572) );
  XOR2_X1 U34490 ( .A1(n15220), .A2(n49109), .Z(n48438) );
  NAND2_X1 U34491 ( .A1(n1642), .A2(n15220), .ZN(n20529) );
  NOR2_X1 U34492 ( .A1(n48440), .A2(n15220), .ZN(n46002) );
  NAND2_X1 U34493 ( .A1(n49789), .A2(n15220), .ZN(n49117) );
  XOR2_X1 U34494 ( .A1(n48436), .A2(n15220), .Z(n48439) );
  NOR2_X1 U34496 ( .A1(n49110), .A2(n15220), .ZN(n47942) );
  INV_X4 U34497 ( .I(n22959), .ZN(n15220) );
  XOR2_X1 U34500 ( .A1(n25911), .A2(n39534), .Z(n15222) );
  INV_X1 U34501 ( .I(n20278), .ZN(n25911) );
  XOR2_X1 U34504 ( .A1(n15615), .A2(n39535), .Z(n15225) );
  INV_X2 U34507 ( .I(n18854), .ZN(n52066) );
  NAND3_X1 U34508 ( .A1(n64147), .A2(n13307), .A3(n22786), .ZN(n39096) );
  NAND3_X1 U34509 ( .A1(n64147), .A2(n13307), .A3(n25570), .ZN(n41038) );
  NAND3_X1 U34510 ( .A1(n64147), .A2(n59255), .A3(n38024), .ZN(n21167) );
  NOR2_X1 U34511 ( .A1(n31315), .A2(n15242), .ZN(n33950) );
  NAND3_X1 U34512 ( .A1(n15244), .A2(n55976), .A3(n15730), .ZN(n52133) );
  NAND3_X1 U34514 ( .A1(n15244), .A2(n55976), .A3(n55668), .ZN(n55448) );
  XOR2_X1 U34517 ( .A1(n64268), .A2(n62380), .Z(n39255) );
  XOR2_X1 U34519 ( .A1(n44969), .A2(n16270), .Z(n15351) );
  XOR2_X1 U34520 ( .A1(n20044), .A2(n44895), .Z(n44969) );
  XOR2_X1 U34523 ( .A1(n2603), .A2(n721), .Z(n18456) );
  NOR3_X1 U34526 ( .A1(n15249), .A2(n54601), .A3(n64307), .ZN(n54327) );
  OAI21_X1 U34527 ( .A1(n54475), .A2(n15249), .B(n54474), .ZN(n54476) );
  OAI22_X1 U34528 ( .A1(n54593), .A2(n15249), .B1(n54603), .B2(n54604), .ZN(
        n15690) );
  NAND2_X1 U34529 ( .A1(n24779), .A2(n15252), .ZN(n41485) );
  NAND2_X1 U34530 ( .A1(n20690), .A2(n60432), .ZN(n20689) );
  NAND3_X2 U34533 ( .A1(n15256), .A2(n15387), .A3(n19026), .ZN(n18295) );
  INV_X2 U34534 ( .I(n15257), .ZN(n24302) );
  OAI21_X1 U34535 ( .A1(n36627), .A2(n35445), .B(n63616), .ZN(n35441) );
  XOR2_X1 U34536 ( .A1(n51693), .A2(n64142), .Z(n15261) );
  XOR2_X1 U34538 ( .A1(n25798), .A2(n8179), .Z(n51700) );
  NOR2_X1 U34540 ( .A1(n13182), .A2(n28705), .ZN(n15267) );
  NOR2_X1 U34542 ( .A1(n24688), .A2(n15318), .ZN(n20896) );
  NOR2_X1 U34543 ( .A1(n10682), .A2(n15318), .ZN(n32765) );
  NOR2_X1 U34546 ( .A1(n15282), .A2(n49376), .ZN(n18225) );
  XOR2_X1 U34551 ( .A1(n15291), .A2(n32747), .Z(n15290) );
  XOR2_X1 U34552 ( .A1(Key[46]), .A2(Ciphertext[159]), .Z(n15338) );
  INV_X2 U34553 ( .I(n38021), .ZN(n16852) );
  XOR2_X1 U34555 ( .A1(n62477), .A2(n46250), .Z(n15297) );
  INV_X2 U34556 ( .I(n20600), .ZN(n22842) );
  NOR2_X2 U34558 ( .A1(n33697), .A2(n32807), .ZN(n15298) );
  NAND3_X1 U34559 ( .A1(n32764), .A2(n32763), .A3(n15303), .ZN(n32768) );
  NAND2_X1 U34560 ( .A1(n15304), .A2(n15435), .ZN(n19834) );
  NOR2_X2 U34561 ( .A1(n18826), .A2(n15305), .ZN(n28646) );
  INV_X1 U34562 ( .I(n15306), .ZN(n22102) );
  XOR2_X1 U34563 ( .A1(n14316), .A2(n52525), .Z(n20954) );
  NAND2_X1 U34564 ( .A1(n42027), .A2(n37536), .ZN(n42592) );
  NOR2_X2 U34565 ( .A1(n62606), .A2(n48847), .ZN(n49511) );
  CLKBUF_X4 U34567 ( .I(n15309), .Z(n15308) );
  XOR2_X1 U34568 ( .A1(n15309), .A2(n10402), .Z(n36637) );
  XOR2_X1 U34570 ( .A1(n15309), .A2(n23927), .Z(n37300) );
  XOR2_X1 U34572 ( .A1(n38062), .A2(n15308), .Z(n38069) );
  NAND2_X2 U34582 ( .A1(n15319), .A2(n49166), .ZN(n49561) );
  NOR2_X1 U34583 ( .A1(n55295), .A2(n55299), .ZN(n19455) );
  XOR2_X1 U34584 ( .A1(n15320), .A2(n9660), .Z(n39481) );
  XOR2_X1 U34585 ( .A1(n15323), .A2(n15322), .Z(n15321) );
  XOR2_X1 U34586 ( .A1(n51911), .A2(n52379), .Z(n15323) );
  NAND3_X1 U34587 ( .A1(n15325), .A2(n48613), .A3(n15324), .ZN(n48617) );
  XOR2_X1 U34589 ( .A1(n33266), .A2(n33265), .Z(n15332) );
  NOR2_X1 U34590 ( .A1(n15333), .A2(n31059), .ZN(n31060) );
  OAI21_X1 U34592 ( .A1(n30064), .A2(n15333), .B(n30176), .ZN(n29035) );
  NOR2_X2 U34593 ( .A1(n42514), .A2(n42515), .ZN(n42985) );
  XOR2_X1 U34597 ( .A1(n8144), .A2(n52209), .Z(n52349) );
  XOR2_X1 U34598 ( .A1(n52205), .A2(n8144), .Z(n51331) );
  INV_X2 U34601 ( .I(n15338), .ZN(n26192) );
  AND2_X1 U34602 ( .A1(n28162), .A2(n22514), .Z(n27452) );
  NOR2_X2 U34603 ( .A1(n29310), .A2(n28858), .ZN(n28162) );
  XOR2_X1 U34605 ( .A1(n45151), .A2(n43648), .Z(n43649) );
  INV_X2 U34607 ( .I(n10291), .ZN(n39307) );
  OAI21_X1 U34608 ( .A1(n49547), .A2(n15349), .B(n49167), .ZN(n15348) );
  XOR2_X1 U34612 ( .A1(n14299), .A2(n52374), .Z(n15353) );
  XOR2_X1 U34613 ( .A1(n21141), .A2(n15355), .Z(n46237) );
  XOR2_X1 U34614 ( .A1(n25531), .A2(n15355), .Z(n46344) );
  OAI22_X1 U34615 ( .A1(n58108), .A2(n29311), .B1(n29316), .B2(n15358), .ZN(
        n29313) );
  OAI21_X1 U34616 ( .A1(n28163), .A2(n15358), .B(n28162), .ZN(n28166) );
  AOI22_X1 U34617 ( .A1(n28863), .A2(n28864), .B1(n29325), .B2(n15358), .ZN(
        n28865) );
  NAND2_X1 U34618 ( .A1(n65208), .A2(n9395), .ZN(n46368) );
  NAND2_X1 U34619 ( .A1(n49411), .A2(n9395), .ZN(n49181) );
  NAND2_X2 U34621 ( .A1(n42503), .A2(n41270), .ZN(n41852) );
  XOR2_X1 U34624 ( .A1(n31603), .A2(n4278), .Z(n15372) );
  INV_X2 U34626 ( .I(n23278), .ZN(n24759) );
  INV_X4 U34627 ( .I(n53368), .ZN(n53345) );
  INV_X1 U34630 ( .I(n19865), .ZN(n15379) );
  XOR2_X1 U34632 ( .A1(n15381), .A2(n901), .Z(n18317) );
  NAND2_X2 U34636 ( .A1(n19758), .A2(n41712), .ZN(n21940) );
  XOR2_X1 U34638 ( .A1(n18295), .A2(n33905), .Z(n22187) );
  NAND2_X2 U34643 ( .A1(n25760), .A2(n41385), .ZN(n39821) );
  NAND2_X2 U34644 ( .A1(n22384), .A2(n41120), .ZN(n25760) );
  INV_X2 U34645 ( .I(n26100), .ZN(n23883) );
  XOR2_X1 U34646 ( .A1(n19299), .A2(n15399), .Z(n15398) );
  XOR2_X1 U34647 ( .A1(n61490), .A2(n24112), .Z(n15399) );
  AOI22_X1 U34655 ( .A1(n31052), .A2(n18839), .B1(n31050), .B2(n15407), .ZN(
        n31058) );
  OAI21_X1 U34656 ( .A1(n30066), .A2(n30065), .B(n60112), .ZN(n30067) );
  INV_X2 U34657 ( .I(n30159), .ZN(n15407) );
  NAND2_X1 U34658 ( .A1(n48330), .A2(n14315), .ZN(n48334) );
  XOR2_X1 U34660 ( .A1(n33827), .A2(n15412), .Z(n16688) );
  NAND2_X2 U34663 ( .A1(n49816), .A2(n18876), .ZN(n49817) );
  NAND2_X2 U34664 ( .A1(n24252), .A2(n46731), .ZN(n20031) );
  NOR2_X2 U34665 ( .A1(n40619), .A2(n39058), .ZN(n40526) );
  INV_X2 U34666 ( .I(n15429), .ZN(n23796) );
  XOR2_X1 U34667 ( .A1(n411), .A2(n50708), .Z(n15430) );
  NAND2_X1 U34669 ( .A1(n35140), .A2(n6052), .ZN(n15432) );
  XOR2_X1 U34670 ( .A1(n32158), .A2(n2952), .Z(n31555) );
  XOR2_X1 U34674 ( .A1(n50436), .A2(n50943), .Z(n51069) );
  XOR2_X1 U34676 ( .A1(n15447), .A2(n52503), .Z(n52504) );
  XOR2_X1 U34677 ( .A1(n15447), .A2(n52580), .Z(n52582) );
  XOR2_X1 U34678 ( .A1(n57908), .A2(n15447), .Z(n50993) );
  XOR2_X1 U34679 ( .A1(n65143), .A2(n15447), .Z(n49960) );
  NAND2_X2 U34684 ( .A1(n55915), .A2(n15454), .ZN(n55718) );
  OAI21_X1 U34685 ( .A1(n23919), .A2(n15454), .B(n55914), .ZN(n55916) );
  NAND2_X1 U34686 ( .A1(n10113), .A2(n15454), .ZN(n55912) );
  OAI21_X1 U34687 ( .A1(n55915), .A2(n15454), .B(n55716), .ZN(n55717) );
  INV_X1 U34689 ( .I(n50682), .ZN(n15460) );
  XOR2_X1 U34690 ( .A1(n51081), .A2(n50685), .Z(n15461) );
  XOR2_X1 U34691 ( .A1(n50948), .A2(n22658), .Z(n15462) );
  XOR2_X1 U34692 ( .A1(n25887), .A2(n15464), .Z(n29259) );
  NOR2_X2 U34696 ( .A1(n8343), .A2(n41354), .ZN(n43219) );
  NAND2_X1 U34699 ( .A1(n27591), .A2(n13320), .ZN(n29783) );
  NAND2_X1 U34700 ( .A1(n15477), .A2(n10419), .ZN(n27558) );
  NAND2_X1 U34703 ( .A1(n28382), .A2(n15477), .ZN(n28391) );
  NAND2_X1 U34707 ( .A1(n25104), .A2(n37463), .ZN(n15483) );
  XOR2_X1 U34708 ( .A1(n15487), .A2(n50583), .Z(n51400) );
  XOR2_X1 U34709 ( .A1(n15489), .A2(n31386), .Z(n25740) );
  OAI21_X1 U34711 ( .A1(n1858), .A2(n60111), .B(n30167), .ZN(n30057) );
  NAND2_X1 U34712 ( .A1(n30174), .A2(n1858), .ZN(n30064) );
  AOI21_X1 U34713 ( .A1(n30696), .A2(n579), .B(n1858), .ZN(n22839) );
  NOR2_X1 U34719 ( .A1(n15501), .A2(n29316), .ZN(n26179) );
  NAND2_X1 U34720 ( .A1(n28853), .A2(n19972), .ZN(n15501) );
  NOR2_X1 U34723 ( .A1(n42428), .A2(n9725), .ZN(n41818) );
  NAND2_X2 U34724 ( .A1(n40063), .A2(n42441), .ZN(n15503) );
  XOR2_X1 U34726 ( .A1(n15505), .A2(n16326), .Z(n22455) );
  AOI21_X1 U34728 ( .A1(n16583), .A2(n16585), .B(n101), .ZN(n15509) );
  XOR2_X1 U34729 ( .A1(n32709), .A2(n15510), .Z(n32711) );
  XOR2_X1 U34730 ( .A1(n15510), .A2(n24698), .Z(n32552) );
  XOR2_X1 U34731 ( .A1(n25653), .A2(n15510), .Z(n25652) );
  INV_X1 U34732 ( .I(n15512), .ZN(n33256) );
  AND2_X1 U34735 ( .A1(n26437), .A2(n26436), .Z(n15515) );
  AND3_X1 U34737 ( .A1(n55088), .A2(n22362), .A3(n4898), .Z(n15519) );
  INV_X2 U34739 ( .I(n15524), .ZN(n15806) );
  XOR2_X1 U34740 ( .A1(n45342), .A2(n17692), .Z(n15525) );
  NAND2_X2 U34741 ( .A1(n1373), .A2(n54860), .ZN(n17499) );
  AOI22_X1 U34743 ( .A1(n27617), .A2(n27618), .B1(n27616), .B2(n10458), .ZN(
        n15535) );
  XOR2_X1 U34744 ( .A1(n51367), .A2(n51366), .Z(n15538) );
  XOR2_X1 U34746 ( .A1(Ciphertext[18]), .A2(Key[115]), .Z(n27559) );
  INV_X2 U34748 ( .I(n15544), .ZN(n15545) );
  NAND2_X2 U34749 ( .A1(n15545), .A2(n35240), .ZN(n35653) );
  OAI21_X1 U34756 ( .A1(n15554), .A2(n15553), .B(n47683), .ZN(n25861) );
  NOR2_X1 U34757 ( .A1(n15555), .A2(n45794), .ZN(n15554) );
  NOR2_X2 U34760 ( .A1(n25860), .A2(n25862), .ZN(n48742) );
  INV_X2 U34761 ( .I(n15560), .ZN(n21253) );
  XOR2_X1 U34762 ( .A1(n46550), .A2(n15563), .Z(n15562) );
  XOR2_X1 U34763 ( .A1(n46549), .A2(n15564), .Z(n15563) );
  INV_X1 U34766 ( .I(n15576), .ZN(n31125) );
  NOR2_X1 U34767 ( .A1(n29442), .A2(n29566), .ZN(n15576) );
  INV_X4 U34768 ( .I(n4706), .ZN(n29916) );
  OR2_X1 U34769 ( .A1(n5194), .A2(n56129), .Z(n19161) );
  XOR2_X1 U34770 ( .A1(n24258), .A2(n24008), .Z(n17728) );
  OAI21_X1 U34771 ( .A1(n15585), .A2(n23108), .B(n40744), .ZN(n39009) );
  XOR2_X1 U34772 ( .A1(n15589), .A2(n32330), .Z(n35002) );
  NOR2_X1 U34775 ( .A1(n28962), .A2(n15592), .ZN(n23187) );
  OAI21_X1 U34776 ( .A1(n29909), .A2(n29566), .B(n9904), .ZN(n15593) );
  XOR2_X1 U34777 ( .A1(n38946), .A2(n9397), .Z(n19249) );
  XOR2_X1 U34778 ( .A1(n19418), .A2(n38307), .Z(n38946) );
  INV_X2 U34780 ( .I(n15597), .ZN(n17128) );
  NOR2_X2 U34781 ( .A1(n47830), .A2(n17128), .ZN(n47664) );
  NOR2_X2 U34782 ( .A1(n26579), .A2(n26580), .ZN(n28229) );
  XOR2_X1 U34783 ( .A1(n15611), .A2(n32499), .Z(n15610) );
  INV_X1 U34788 ( .I(n19564), .ZN(n15621) );
  OR2_X2 U34790 ( .A1(n21067), .A2(n21279), .Z(n25702) );
  XOR2_X1 U34791 ( .A1(n32247), .A2(n57218), .Z(n32563) );
  XOR2_X1 U34795 ( .A1(n15630), .A2(n39479), .Z(n18999) );
  XOR2_X1 U34796 ( .A1(n15631), .A2(n55516), .Z(n38088) );
  XOR2_X1 U34797 ( .A1(n15630), .A2(n37954), .Z(n37955) );
  XOR2_X1 U34798 ( .A1(n15630), .A2(n37307), .Z(n37308) );
  XOR2_X1 U34799 ( .A1(n16594), .A2(n15630), .Z(n38704) );
  XOR2_X1 U34800 ( .A1(n15074), .A2(n15889), .Z(n25957) );
  AND2_X1 U34801 ( .A1(n43313), .A2(n15637), .Z(n15636) );
  NAND2_X1 U34802 ( .A1(n43307), .A2(n43308), .ZN(n15638) );
  NAND2_X1 U34803 ( .A1(n16880), .A2(n1334), .ZN(n15639) );
  XOR2_X1 U34805 ( .A1(n15644), .A2(n56202), .Z(n39455) );
  XOR2_X1 U34806 ( .A1(n15644), .A2(n38866), .Z(n38006) );
  XOR2_X1 U34807 ( .A1(n15644), .A2(n39736), .Z(n39745) );
  INV_X2 U34808 ( .I(n15645), .ZN(n42285) );
  XNOR2_X1 U34810 ( .A1(n15646), .A2(n15950), .ZN(n15645) );
  XOR2_X1 U34811 ( .A1(n19531), .A2(n63081), .Z(n15646) );
  XOR2_X1 U34814 ( .A1(n18452), .A2(n17939), .Z(n39247) );
  NAND2_X1 U34815 ( .A1(n1569), .A2(n16470), .ZN(n20546) );
  NAND2_X2 U34816 ( .A1(n10747), .A2(n23337), .ZN(n16470) );
  INV_X2 U34818 ( .I(n15650), .ZN(n28032) );
  XOR2_X1 U34819 ( .A1(n15654), .A2(n15653), .Z(n15652) );
  XOR2_X1 U34820 ( .A1(n721), .A2(n50959), .Z(n15654) );
  NAND2_X1 U34821 ( .A1(n41636), .A2(n43217), .ZN(n15658) );
  INV_X2 U34823 ( .I(n44145), .ZN(n46385) );
  XOR2_X1 U34826 ( .A1(n22338), .A2(n62989), .Z(n51380) );
  XOR2_X1 U34827 ( .A1(n62989), .A2(n50163), .Z(n50164) );
  XOR2_X1 U34828 ( .A1(n62989), .A2(n24757), .Z(n50954) );
  INV_X1 U34830 ( .I(n24367), .ZN(n45805) );
  INV_X2 U34831 ( .I(n36116), .ZN(n21591) );
  INV_X2 U34832 ( .I(n15675), .ZN(n15807) );
  XOR2_X1 U34834 ( .A1(n32664), .A2(n33194), .Z(n15678) );
  NAND2_X1 U34835 ( .A1(n15683), .A2(n55416), .ZN(n15682) );
  OAI21_X1 U34836 ( .A1(n65010), .A2(n55412), .B(n55256), .ZN(n15683) );
  XOR2_X1 U34838 ( .A1(n30985), .A2(n15685), .Z(n16953) );
  NOR2_X2 U34839 ( .A1(n29584), .A2(n15686), .ZN(n30985) );
  INV_X2 U34840 ( .I(n15687), .ZN(n32748) );
  INV_X1 U34841 ( .I(n24448), .ZN(n29570) );
  NAND2_X2 U34842 ( .A1(n28920), .A2(n30292), .ZN(n21832) );
  INV_X2 U34844 ( .I(n54670), .ZN(n54768) );
  NAND3_X1 U34845 ( .A1(n21992), .A2(n41870), .A3(n42527), .ZN(n23558) );
  INV_X1 U34846 ( .I(n16025), .ZN(n25161) );
  BUF_X4 U34847 ( .I(n16900), .Z(n16402) );
  NAND2_X2 U34848 ( .A1(n18051), .A2(n19248), .ZN(n42397) );
  INV_X4 U34852 ( .I(n38758), .ZN(n40749) );
  CLKBUF_X2 U34853 ( .I(Key[49]), .Z(n53945) );
  INV_X2 U34856 ( .I(n44435), .ZN(n46897) );
  INV_X1 U34861 ( .I(n34586), .ZN(n22333) );
  BUF_X4 U34863 ( .I(n30953), .Z(n17414) );
  NAND2_X1 U34864 ( .A1(n40319), .A2(n40087), .ZN(n39411) );
  AOI21_X2 U34865 ( .A1(n1121), .A2(n48315), .B(n48745), .ZN(n48028) );
  INV_X4 U34866 ( .I(n21492), .ZN(n42287) );
  BUF_X4 U34868 ( .I(n30620), .Z(n16750) );
  NAND3_X1 U34870 ( .A1(n54921), .A2(n13671), .A3(n2049), .ZN(n54922) );
  INV_X1 U34871 ( .I(n26334), .ZN(n26640) );
  NAND2_X2 U34872 ( .A1(n27171), .A2(n28312), .ZN(n27602) );
  INV_X2 U34873 ( .I(n35201), .ZN(n35611) );
  INV_X4 U34875 ( .I(n17632), .ZN(n28127) );
  INV_X4 U34876 ( .I(n30558), .ZN(n31083) );
  BUF_X4 U34879 ( .I(n25595), .Z(n21945) );
  NAND2_X1 U34880 ( .A1(n18945), .A2(n18944), .ZN(n18943) );
  AOI21_X1 U34882 ( .A1(n34871), .A2(n16690), .B(n19814), .ZN(n19629) );
  NOR2_X2 U34883 ( .A1(n37269), .A2(n17243), .ZN(n34849) );
  OR2_X2 U34887 ( .A1(n39317), .A2(n22069), .Z(n40224) );
  OAI21_X1 U34888 ( .A1(n50604), .A2(n52670), .B(n50603), .ZN(n17170) );
  NAND2_X2 U34892 ( .A1(n29628), .A2(n28119), .ZN(n28125) );
  NOR2_X1 U34893 ( .A1(n22208), .A2(n23340), .ZN(n42364) );
  OAI21_X1 U34895 ( .A1(n16410), .A2(n43690), .B(n16409), .ZN(n37833) );
  INV_X1 U34897 ( .I(n33372), .ZN(n33115) );
  NOR2_X1 U34898 ( .A1(n34041), .A2(n33984), .ZN(n21242) );
  NAND2_X1 U34899 ( .A1(n34197), .A2(n5386), .ZN(n24160) );
  NAND2_X1 U34900 ( .A1(n27015), .A2(n28222), .ZN(n27016) );
  INV_X1 U34901 ( .I(n23695), .ZN(n19983) );
  INV_X1 U34902 ( .I(n28280), .ZN(n27404) );
  INV_X1 U34903 ( .I(n50850), .ZN(n17941) );
  INV_X1 U34904 ( .I(n21488), .ZN(n18302) );
  INV_X1 U34905 ( .I(n32065), .ZN(n18543) );
  INV_X1 U34907 ( .I(n33231), .ZN(n24043) );
  NOR2_X1 U34908 ( .A1(n24549), .A2(n35648), .ZN(n33592) );
  NOR2_X1 U34909 ( .A1(n24550), .A2(n33802), .ZN(n24549) );
  NAND2_X1 U34910 ( .A1(n35660), .A2(n33801), .ZN(n24550) );
  NOR2_X1 U34913 ( .A1(n24664), .A2(n5410), .ZN(n32884) );
  NAND2_X1 U34915 ( .A1(n21292), .A2(n61896), .ZN(n21291) );
  NOR2_X1 U34916 ( .A1(n33702), .A2(n16856), .ZN(n32531) );
  NAND2_X1 U34917 ( .A1(n32526), .A2(n32525), .ZN(n19467) );
  NAND2_X1 U34919 ( .A1(n20706), .A2(n35276), .ZN(n17297) );
  NOR3_X1 U34920 ( .A1(n504), .A2(n5936), .A3(n36946), .ZN(n34904) );
  INV_X1 U34924 ( .I(n36105), .ZN(n38496) );
  INV_X2 U34927 ( .I(n24989), .ZN(n26270) );
  NAND2_X1 U34928 ( .A1(n29491), .A2(n28209), .ZN(n31094) );
  INV_X1 U34930 ( .I(n39681), .ZN(n18555) );
  INV_X1 U34932 ( .I(n28395), .ZN(n26343) );
  AOI21_X1 U34933 ( .A1(n59015), .A2(n64277), .B(n41167), .ZN(n40539) );
  NAND2_X1 U34934 ( .A1(n42286), .A2(n16680), .ZN(n42289) );
  NAND2_X1 U34935 ( .A1(n16171), .A2(n42273), .ZN(n16806) );
  NOR2_X1 U34936 ( .A1(n58307), .A2(n17752), .ZN(n17751) );
  NAND2_X1 U34939 ( .A1(n19742), .A2(n22228), .ZN(n18725) );
  NOR2_X1 U34942 ( .A1(n20911), .A2(n49682), .ZN(n18007) );
  INV_X1 U34944 ( .I(n48652), .ZN(n22233) );
  INV_X1 U34945 ( .I(n48648), .ZN(n17082) );
  OAI21_X1 U34946 ( .A1(n48647), .A2(n48646), .B(n18282), .ZN(n17083) );
  OAI21_X1 U34947 ( .A1(n48631), .A2(n12993), .B(n48630), .ZN(n48634) );
  NAND2_X1 U34952 ( .A1(n45750), .A2(n15076), .ZN(n45501) );
  NAND2_X1 U34953 ( .A1(n45480), .A2(n45481), .ZN(n25077) );
  NAND3_X1 U34954 ( .A1(n45783), .A2(n45782), .A3(n45784), .ZN(n20184) );
  NOR2_X1 U34955 ( .A1(n47531), .A2(n24801), .ZN(n47533) );
  NAND2_X1 U34956 ( .A1(n47536), .A2(n47532), .ZN(n25387) );
  INV_X1 U34959 ( .I(n45809), .ZN(n45810) );
  NOR2_X1 U34960 ( .A1(n46821), .A2(n21451), .ZN(n20110) );
  NOR2_X1 U34961 ( .A1(n47288), .A2(n22908), .ZN(n22011) );
  AOI21_X1 U34964 ( .A1(n23661), .A2(n18570), .B(n48668), .ZN(n18569) );
  NAND2_X1 U34965 ( .A1(n64969), .A2(n45517), .ZN(n19987) );
  OAI21_X1 U34968 ( .A1(n1291), .A2(n21870), .B(n50348), .ZN(n17899) );
  INV_X1 U34972 ( .I(n46092), .ZN(n23208) );
  INV_X1 U34973 ( .I(n7229), .ZN(n24132) );
  NOR2_X1 U34975 ( .A1(n55434), .A2(n55436), .ZN(n52491) );
  NOR2_X1 U34976 ( .A1(n20177), .A2(n20176), .ZN(n20175) );
  INV_X1 U34977 ( .I(n55323), .ZN(n20176) );
  OAI21_X1 U34978 ( .A1(n55318), .A2(n52487), .B(n55006), .ZN(n22825) );
  NAND2_X1 U34979 ( .A1(n52489), .A2(n24454), .ZN(n22824) );
  INV_X1 U34981 ( .I(n33155), .ZN(n17120) );
  NOR2_X1 U34983 ( .A1(n34752), .A2(n21731), .ZN(n21730) );
  INV_X1 U34986 ( .I(n20989), .ZN(n21849) );
  OAI21_X1 U34988 ( .A1(n7342), .A2(n445), .B(n35612), .ZN(n33551) );
  NAND3_X1 U34990 ( .A1(n59432), .A2(n34564), .A3(n33752), .ZN(n33754) );
  NAND2_X1 U34991 ( .A1(n34571), .A2(n34564), .ZN(n22189) );
  INV_X1 U34992 ( .I(n31537), .ZN(n18933) );
  NAND3_X1 U34993 ( .A1(n35302), .A2(n17614), .A3(n35301), .ZN(n20107) );
  INV_X1 U34994 ( .I(n35299), .ZN(n20105) );
  INV_X1 U34995 ( .I(n34957), .ZN(n21613) );
  NAND2_X1 U34996 ( .A1(n18300), .A2(n58472), .ZN(n34067) );
  NAND2_X1 U34997 ( .A1(n34056), .A2(n34679), .ZN(n16661) );
  NAND2_X1 U35000 ( .A1(n34624), .A2(n20279), .ZN(n20207) );
  NAND2_X1 U35001 ( .A1(n20206), .A2(n22226), .ZN(n20205) );
  INV_X1 U35002 ( .I(n16347), .ZN(n34232) );
  NAND2_X1 U35004 ( .A1(n17538), .A2(n34268), .ZN(n32218) );
  NOR2_X1 U35005 ( .A1(n34741), .A2(n22278), .ZN(n24540) );
  NAND2_X1 U35008 ( .A1(n33645), .A2(n33541), .ZN(n20799) );
  NAND3_X1 U35010 ( .A1(n34029), .A2(n34028), .A3(n34027), .ZN(n34030) );
  INV_X1 U35011 ( .I(n33324), .ZN(n33323) );
  NAND2_X1 U35013 ( .A1(n32022), .A2(n32021), .ZN(n24457) );
  INV_X1 U35014 ( .I(n35280), .ZN(n34391) );
  OAI22_X1 U35016 ( .A1(n33985), .A2(n21106), .B1(n31023), .B2(n21242), .ZN(
        n33986) );
  NAND2_X1 U35019 ( .A1(n33946), .A2(n33947), .ZN(n20064) );
  NAND2_X1 U35020 ( .A1(n20524), .A2(n62931), .ZN(n33954) );
  NAND2_X1 U35024 ( .A1(n33593), .A2(n33590), .ZN(n24925) );
  OAI21_X1 U35025 ( .A1(n34360), .A2(n21461), .B(n21460), .ZN(n21193) );
  OAI22_X1 U35028 ( .A1(n33499), .A2(n34964), .B1(n57423), .B2(n19563), .ZN(
        n30964) );
  NAND3_X1 U35029 ( .A1(n63578), .A2(n60628), .A3(n60554), .ZN(n20550) );
  AOI21_X1 U35031 ( .A1(n21484), .A2(n23556), .B(n21483), .ZN(n21482) );
  AOI21_X1 U35034 ( .A1(n34196), .A2(n60684), .B(n21291), .ZN(n24410) );
  NAND2_X1 U35035 ( .A1(n33808), .A2(n35220), .ZN(n20256) );
  NAND2_X1 U35037 ( .A1(n33317), .A2(n33316), .ZN(n24635) );
  AOI21_X1 U35039 ( .A1(n33559), .A2(n32511), .B(n19467), .ZN(n32535) );
  AOI22_X1 U35040 ( .A1(n32532), .A2(n33559), .B1(n32531), .B2(n33695), .ZN(
        n32533) );
  INV_X1 U35042 ( .I(n39368), .ZN(n21609) );
  NAND2_X1 U35043 ( .A1(n36722), .A2(n36723), .ZN(n25919) );
  INV_X1 U35045 ( .I(n38780), .ZN(n24662) );
  NAND3_X1 U35047 ( .A1(n60990), .A2(n60894), .A3(n27320), .ZN(n17991) );
  NOR2_X1 U35048 ( .A1(n1970), .A2(n7112), .ZN(n20609) );
  NAND3_X1 U35049 ( .A1(n19287), .A2(n28620), .A3(n27689), .ZN(n18038) );
  NAND2_X1 U35055 ( .A1(n40765), .A2(n18661), .ZN(n18660) );
  NAND2_X1 U35057 ( .A1(n23823), .A2(n64994), .ZN(n26938) );
  NAND2_X1 U35058 ( .A1(n9098), .A2(n17451), .ZN(n29140) );
  NAND2_X1 U35059 ( .A1(n23430), .A2(n22945), .ZN(n23973) );
  INV_X1 U35060 ( .I(n28161), .ZN(n29323) );
  AOI21_X1 U35062 ( .A1(n26574), .A2(n26573), .B(n28039), .ZN(n26576) );
  NAND2_X1 U35063 ( .A1(n27982), .A2(n27981), .ZN(n18528) );
  AND3_X1 U35065 ( .A1(n27384), .A2(n27045), .A3(n16042), .Z(n16150) );
  NAND3_X1 U35067 ( .A1(n28044), .A2(n22671), .A3(n22670), .ZN(n26284) );
  NAND2_X1 U35068 ( .A1(n27025), .A2(n24836), .ZN(n22670) );
  NAND2_X1 U35071 ( .A1(n27470), .A2(n27464), .ZN(n27227) );
  NOR3_X1 U35073 ( .A1(n23053), .A2(n30538), .A3(n15205), .ZN(n16696) );
  NAND2_X1 U35076 ( .A1(n39899), .A2(n17945), .ZN(n17357) );
  NOR2_X1 U35077 ( .A1(n19592), .A2(n17752), .ZN(n17354) );
  INV_X1 U35078 ( .I(n39242), .ZN(n18304) );
  NAND2_X1 U35079 ( .A1(n20190), .A2(n38273), .ZN(n38274) );
  NAND2_X1 U35082 ( .A1(n39097), .A2(n39096), .ZN(n21386) );
  NAND2_X1 U35083 ( .A1(n40514), .A2(n15799), .ZN(n21384) );
  NOR2_X1 U35084 ( .A1(n39318), .A2(n23515), .ZN(n23550) );
  NOR2_X1 U35086 ( .A1(n18704), .A2(n60820), .ZN(n40972) );
  NOR2_X1 U35088 ( .A1(n64940), .A2(n63891), .ZN(n18764) );
  NOR2_X1 U35089 ( .A1(n30817), .A2(n29835), .ZN(n29234) );
  OAI21_X1 U35090 ( .A1(n27933), .A2(n27932), .B(n27931), .ZN(n17250) );
  NOR2_X1 U35091 ( .A1(n62083), .A2(n26610), .ZN(n27117) );
  NAND2_X1 U35092 ( .A1(n25774), .A2(n28076), .ZN(n17174) );
  NAND2_X1 U35094 ( .A1(n27614), .A2(n22958), .ZN(n22957) );
  AOI21_X1 U35096 ( .A1(n28026), .A2(n60885), .B(n15836), .ZN(n25301) );
  NAND2_X1 U35097 ( .A1(n27066), .A2(n28024), .ZN(n27068) );
  NOR2_X1 U35098 ( .A1(n26563), .A2(n26562), .ZN(n25756) );
  OAI21_X1 U35099 ( .A1(n26566), .A2(n26567), .B(n26092), .ZN(n22560) );
  NAND2_X1 U35100 ( .A1(n27150), .A2(n25096), .ZN(n27800) );
  NAND2_X1 U35102 ( .A1(n26132), .A2(n26131), .ZN(n26130) );
  NOR2_X1 U35103 ( .A1(n40066), .A2(n25661), .ZN(n25469) );
  NAND3_X1 U35104 ( .A1(n6576), .A2(n40070), .A3(n40069), .ZN(n40072) );
  NOR3_X1 U35107 ( .A1(n43956), .A2(n43957), .A3(n1299), .ZN(n25670) );
  INV_X1 U35108 ( .I(n43418), .ZN(n43625) );
  NAND2_X1 U35110 ( .A1(n42278), .A2(n22713), .ZN(n16881) );
  OAI21_X1 U35111 ( .A1(n14280), .A2(n1273), .B(n42517), .ZN(n42203) );
  INV_X1 U35112 ( .I(n38413), .ZN(n25423) );
  OAI21_X1 U35113 ( .A1(n43695), .A2(n4274), .B(n22989), .ZN(n20285) );
  OAI21_X1 U35117 ( .A1(n41834), .A2(n41835), .B(n41833), .ZN(n20006) );
  NOR2_X1 U35118 ( .A1(n41798), .A2(n42228), .ZN(n17294) );
  NAND2_X1 U35119 ( .A1(n42671), .A2(n42670), .ZN(n17963) );
  INV_X1 U35120 ( .I(n30454), .ZN(n19027) );
  NOR2_X1 U35121 ( .A1(n21095), .A2(n58448), .ZN(n30452) );
  NAND2_X1 U35125 ( .A1(n40131), .A2(n60860), .ZN(n16400) );
  OAI21_X1 U35126 ( .A1(n40324), .A2(n16397), .B(n40087), .ZN(n16396) );
  NOR2_X1 U35127 ( .A1(n60929), .A2(n61264), .ZN(n16397) );
  NAND2_X1 U35129 ( .A1(n43037), .A2(n4276), .ZN(n22130) );
  AOI22_X1 U35131 ( .A1(n43379), .A2(n43378), .B1(n43376), .B2(n43377), .ZN(
        n24129) );
  NAND2_X1 U35132 ( .A1(n43568), .A2(n20331), .ZN(n20330) );
  NAND2_X1 U35133 ( .A1(n43554), .A2(n17245), .ZN(n20331) );
  NOR2_X1 U35134 ( .A1(n43555), .A2(n17245), .ZN(n20329) );
  NAND4_X1 U35135 ( .A1(n47703), .A2(n47811), .A3(n8048), .A4(n47384), .ZN(
        n47395) );
  NOR2_X1 U35136 ( .A1(n16538), .A2(n16628), .ZN(n48215) );
  NAND3_X1 U35137 ( .A1(n16533), .A2(n47490), .A3(n48668), .ZN(n25930) );
  INV_X1 U35139 ( .I(n21803), .ZN(n21977) );
  NAND2_X1 U35140 ( .A1(n45672), .A2(n21976), .ZN(n21975) );
  OAI21_X1 U35141 ( .A1(n4315), .A2(n47261), .B(n9730), .ZN(n21980) );
  NAND2_X1 U35143 ( .A1(n45984), .A2(n47615), .ZN(n19739) );
  NAND2_X1 U35144 ( .A1(n47240), .A2(n62739), .ZN(n19740) );
  NOR2_X1 U35146 ( .A1(n1295), .A2(n10088), .ZN(n18351) );
  NAND2_X1 U35147 ( .A1(n47612), .A2(n47613), .ZN(n18349) );
  OAI21_X1 U35149 ( .A1(n23850), .A2(n46810), .B(n16950), .ZN(n17771) );
  NOR2_X1 U35151 ( .A1(n22599), .A2(n18099), .ZN(n20687) );
  OAI21_X1 U35152 ( .A1(n48146), .A2(n22599), .B(n23185), .ZN(n21398) );
  OAI21_X1 U35155 ( .A1(n47862), .A2(n47861), .B(n10405), .ZN(n47865) );
  NOR2_X1 U35156 ( .A1(n15825), .A2(n15748), .ZN(n47145) );
  AND3_X1 U35157 ( .A1(n46830), .A2(n46829), .A3(n46828), .Z(n46831) );
  NAND2_X1 U35158 ( .A1(n19558), .A2(n4428), .ZN(n48231) );
  INV_X1 U35159 ( .I(n63098), .ZN(n45749) );
  INV_X1 U35161 ( .I(n47492), .ZN(n17006) );
  OAI22_X1 U35163 ( .A1(n47202), .A2(n20679), .B1(n47197), .B2(n48194), .ZN(
        n46258) );
  INV_X1 U35164 ( .I(n46260), .ZN(n17009) );
  NOR2_X1 U35165 ( .A1(n14473), .A2(n14121), .ZN(n47716) );
  NAND2_X1 U35166 ( .A1(n44573), .A2(n44711), .ZN(n18320) );
  OAI22_X1 U35167 ( .A1(n45301), .A2(n62321), .B1(n63686), .B2(n59528), .ZN(
        n20568) );
  AOI21_X1 U35168 ( .A1(n63700), .A2(n46064), .B(n46926), .ZN(n21558) );
  NAND2_X1 U35169 ( .A1(n33434), .A2(n23223), .ZN(n17419) );
  OAI21_X1 U35171 ( .A1(n48530), .A2(n21177), .B(n18118), .ZN(n47192) );
  NOR2_X1 U35173 ( .A1(n50398), .A2(n50395), .ZN(n49029) );
  NAND3_X1 U35174 ( .A1(n48552), .A2(n47096), .A3(n21820), .ZN(n46802) );
  OAI21_X1 U35175 ( .A1(n57670), .A2(n45786), .B(n45785), .ZN(n20185) );
  AOI21_X1 U35176 ( .A1(n47895), .A2(n47900), .B(n17970), .ZN(n45949) );
  AND3_X1 U35178 ( .A1(n45995), .A2(n45994), .A3(n45993), .Z(n15971) );
  NAND2_X1 U35180 ( .A1(n64548), .A2(n14473), .ZN(n47892) );
  NOR2_X1 U35182 ( .A1(n19867), .A2(n18918), .ZN(n48275) );
  NAND2_X1 U35183 ( .A1(n34978), .A2(n34979), .ZN(n19474) );
  NAND3_X1 U35185 ( .A1(n53219), .A2(n57030), .A3(n50739), .ZN(n25110) );
  NAND2_X1 U35190 ( .A1(n56441), .A2(n56435), .ZN(n55986) );
  NAND2_X1 U35191 ( .A1(n20757), .A2(n55695), .ZN(n20756) );
  NAND2_X1 U35192 ( .A1(n55696), .A2(n55299), .ZN(n20757) );
  NOR3_X1 U35193 ( .A1(n55496), .A2(n17979), .A3(n64019), .ZN(n23272) );
  NAND3_X1 U35195 ( .A1(n23047), .A2(n1457), .A3(n23857), .ZN(n50480) );
  AOI21_X1 U35196 ( .A1(n53548), .A2(n16487), .B(n21971), .ZN(n21972) );
  OAI21_X1 U35199 ( .A1(n54949), .A2(n54783), .B(n54610), .ZN(n19494) );
  NOR3_X1 U35201 ( .A1(n18192), .A2(n53396), .A3(n20630), .ZN(n18193) );
  NAND2_X1 U35202 ( .A1(n58763), .A2(n1457), .ZN(n18192) );
  INV_X1 U35203 ( .I(n53177), .ZN(n17260) );
  OAI21_X1 U35204 ( .A1(n3916), .A2(n54457), .B(n54331), .ZN(n26118) );
  NAND2_X1 U35206 ( .A1(n9613), .A2(n19401), .ZN(n53886) );
  AOI22_X1 U35207 ( .A1(n54018), .A2(n53881), .B1(n23482), .B2(n54346), .ZN(
        n17036) );
  NAND2_X1 U35212 ( .A1(n54495), .A2(n21297), .ZN(n51839) );
  NOR2_X1 U35214 ( .A1(n55854), .A2(n55885), .ZN(n55846) );
  INV_X1 U35215 ( .I(n55264), .ZN(n54995) );
  INV_X1 U35216 ( .I(n33070), .ZN(n20931) );
  INV_X1 U35217 ( .I(n13181), .ZN(n18675) );
  INV_X1 U35219 ( .I(n23950), .ZN(n17104) );
  OAI22_X1 U35223 ( .A1(n33724), .A2(n22419), .B1(n33725), .B2(n127), .ZN(
        n33726) );
  NAND2_X1 U35227 ( .A1(n34752), .A2(n17538), .ZN(n32019) );
  NAND2_X1 U35228 ( .A1(n33500), .A2(n32919), .ZN(n32920) );
  NAND2_X1 U35229 ( .A1(n34741), .A2(n34742), .ZN(n19444) );
  NAND2_X1 U35231 ( .A1(n33406), .A2(n3549), .ZN(n17548) );
  AOI21_X1 U35232 ( .A1(n5082), .A2(n1542), .B(n1796), .ZN(n17547) );
  NAND2_X1 U35233 ( .A1(n23556), .A2(n25389), .ZN(n35308) );
  NOR2_X1 U35235 ( .A1(n34320), .A2(n23556), .ZN(n18799) );
  INV_X1 U35237 ( .I(n33981), .ZN(n18935) );
  NAND3_X1 U35238 ( .A1(n18390), .A2(n32890), .A3(n18277), .ZN(n17039) );
  AOI21_X1 U35239 ( .A1(n34200), .A2(n18680), .B(n31775), .ZN(n19826) );
  NAND2_X1 U35240 ( .A1(n4834), .A2(n10226), .ZN(n19347) );
  INV_X1 U35241 ( .I(n33798), .ZN(n33794) );
  NOR2_X1 U35244 ( .A1(n34348), .A2(n34347), .ZN(n19007) );
  AOI21_X1 U35245 ( .A1(n34746), .A2(n34752), .B(n34346), .ZN(n34347) );
  NOR2_X1 U35246 ( .A1(n1811), .A2(n61090), .ZN(n33321) );
  INV_X1 U35247 ( .I(n35624), .ZN(n33316) );
  INV_X1 U35249 ( .I(n36627), .ZN(n36365) );
  NOR2_X1 U35250 ( .A1(n36423), .A2(n36169), .ZN(n22184) );
  NOR2_X1 U35252 ( .A1(n57200), .A2(n35670), .ZN(n22402) );
  INV_X1 U35253 ( .I(n8438), .ZN(n25775) );
  NOR2_X1 U35255 ( .A1(n35379), .A2(n24078), .ZN(n35460) );
  NOR2_X1 U35256 ( .A1(n2383), .A2(n37425), .ZN(n35510) );
  NOR2_X1 U35257 ( .A1(n37435), .A2(n22461), .ZN(n16442) );
  OAI21_X1 U35259 ( .A1(n22595), .A2(n2383), .B(n58220), .ZN(n35512) );
  NOR2_X1 U35260 ( .A1(n18092), .A2(n18130), .ZN(n36500) );
  NAND2_X1 U35261 ( .A1(n16268), .A2(n36483), .ZN(n18092) );
  NAND2_X1 U35262 ( .A1(n21186), .A2(n22733), .ZN(n21185) );
  INV_X1 U35266 ( .I(n21880), .ZN(n37392) );
  INV_X1 U35267 ( .I(n36764), .ZN(n34851) );
  NAND3_X1 U35268 ( .A1(n32220), .A2(n32219), .A3(n31976), .ZN(n24538) );
  NAND2_X1 U35270 ( .A1(n7092), .A2(n36847), .ZN(n35408) );
  NAND3_X1 U35273 ( .A1(n8808), .A2(n4798), .A3(n21881), .ZN(n36869) );
  NAND2_X1 U35275 ( .A1(n59910), .A2(n36777), .ZN(n34007) );
  AOI21_X1 U35276 ( .A1(n23584), .A2(n35567), .B(n24118), .ZN(n35564) );
  NAND2_X1 U35279 ( .A1(n34869), .A2(n35901), .ZN(n16690) );
  NAND3_X1 U35280 ( .A1(n21150), .A2(n35148), .A3(n62026), .ZN(n20131) );
  NAND2_X1 U35281 ( .A1(n35975), .A2(n35543), .ZN(n21147) );
  NAND2_X1 U35282 ( .A1(n33717), .A2(n23577), .ZN(n20136) );
  INV_X1 U35283 ( .I(n33412), .ZN(n24627) );
  NAND3_X1 U35285 ( .A1(n36493), .A2(n18348), .A3(n24028), .ZN(n36235) );
  NAND3_X1 U35287 ( .A1(n36162), .A2(n36597), .A3(n36590), .ZN(n36164) );
  OAI21_X1 U35289 ( .A1(n35424), .A2(n25154), .B(n17720), .ZN(n25152) );
  NOR2_X1 U35291 ( .A1(n18602), .A2(n36408), .ZN(n18574) );
  NAND2_X1 U35292 ( .A1(n33606), .A2(n21591), .ZN(n17394) );
  OAI22_X1 U35295 ( .A1(n17851), .A2(n36473), .B1(n36475), .B2(n36474), .ZN(
        n36476) );
  NOR2_X1 U35297 ( .A1(n34903), .A2(n35431), .ZN(n36950) );
  NAND2_X1 U35298 ( .A1(n23449), .A2(n37225), .ZN(n36615) );
  NOR2_X1 U35299 ( .A1(n28632), .A2(n28630), .ZN(n20629) );
  AOI21_X1 U35301 ( .A1(n32856), .A2(n34462), .B(n32857), .ZN(n17192) );
  NOR2_X1 U35303 ( .A1(n24775), .A2(n35994), .ZN(n36604) );
  NAND2_X1 U35304 ( .A1(n17633), .A2(n25151), .ZN(n27322) );
  NOR2_X1 U35305 ( .A1(n28802), .A2(n22158), .ZN(n25151) );
  NAND3_X1 U35306 ( .A1(n20097), .A2(n26912), .A3(n29694), .ZN(n19163) );
  NOR2_X1 U35307 ( .A1(n64128), .A2(n31115), .ZN(n16388) );
  NAND2_X1 U35308 ( .A1(n28227), .A2(n28226), .ZN(n18263) );
  NAND3_X1 U35309 ( .A1(n26544), .A2(n26606), .A3(n28367), .ZN(n23085) );
  INV_X1 U35310 ( .I(n27696), .ZN(n26885) );
  INV_X1 U35311 ( .I(n29179), .ZN(n17278) );
  NAND2_X1 U35312 ( .A1(n28258), .A2(n17909), .ZN(n27937) );
  INV_X1 U35313 ( .I(n17103), .ZN(n27938) );
  AOI22_X1 U35314 ( .A1(n28163), .A2(n29316), .B1(n29322), .B2(n28860), .ZN(
        n26925) );
  NAND2_X1 U35316 ( .A1(n28239), .A2(n97), .ZN(n24818) );
  OAI21_X1 U35317 ( .A1(n29711), .A2(n29710), .B(n17688), .ZN(n20088) );
  NAND2_X1 U35318 ( .A1(n28858), .A2(n29310), .ZN(n27449) );
  NOR2_X1 U35319 ( .A1(n29714), .A2(n7112), .ZN(n28634) );
  NOR3_X1 U35321 ( .A1(n29176), .A2(n29175), .A3(n29174), .ZN(n29185) );
  NOR2_X1 U35322 ( .A1(n29182), .A2(n29181), .ZN(n23892) );
  AOI21_X1 U35323 ( .A1(n29291), .A2(n17988), .B(n23732), .ZN(n17987) );
  NOR2_X1 U35324 ( .A1(n40092), .A2(n40090), .ZN(n39398) );
  NOR2_X1 U35325 ( .A1(n41031), .A2(n59255), .ZN(n38025) );
  OAI21_X1 U35326 ( .A1(n39948), .A2(n40825), .B(n39947), .ZN(n39952) );
  INV_X1 U35327 ( .I(n41077), .ZN(n40393) );
  NOR2_X1 U35329 ( .A1(n28375), .A2(n23039), .ZN(n16619) );
  NAND2_X1 U35331 ( .A1(n20561), .A2(n23540), .ZN(n20608) );
  NOR2_X1 U35333 ( .A1(n21158), .A2(n23586), .ZN(n28235) );
  NAND2_X1 U35334 ( .A1(n28245), .A2(n21158), .ZN(n28246) );
  NAND2_X1 U35335 ( .A1(n28869), .A2(n29668), .ZN(n20215) );
  NAND3_X1 U35336 ( .A1(n27970), .A2(n28212), .A3(n63714), .ZN(n27971) );
  NOR2_X1 U35337 ( .A1(n31092), .A2(n24199), .ZN(n30383) );
  NAND2_X1 U35338 ( .A1(n27389), .A2(n28239), .ZN(n28064) );
  NAND2_X1 U35341 ( .A1(n26871), .A2(n17688), .ZN(n26872) );
  NAND2_X1 U35344 ( .A1(n28805), .A2(n28804), .ZN(n17459) );
  AOI22_X1 U35345 ( .A1(n28801), .A2(n18515), .B1(n23773), .B2(n28813), .ZN(
        n17458) );
  NAND2_X1 U35346 ( .A1(n17634), .A2(n28812), .ZN(n28819) );
  NOR2_X1 U35347 ( .A1(n26970), .A2(n26969), .ZN(n27493) );
  NAND3_X1 U35348 ( .A1(n27853), .A2(n27849), .A3(n28510), .ZN(n26418) );
  OAI21_X1 U35349 ( .A1(n23386), .A2(n29634), .B(n19462), .ZN(n29640) );
  NAND3_X1 U35351 ( .A1(n1566), .A2(n27897), .A3(n29689), .ZN(n20071) );
  AOI21_X1 U35353 ( .A1(n28661), .A2(n28660), .B(n28659), .ZN(n20171) );
  NOR2_X1 U35355 ( .A1(n26819), .A2(n26820), .ZN(n17604) );
  NAND2_X1 U35356 ( .A1(n27843), .A2(n28490), .ZN(n26402) );
  NAND2_X1 U35357 ( .A1(n27261), .A2(n29153), .ZN(n23000) );
  NAND2_X1 U35358 ( .A1(n16419), .A2(n28510), .ZN(n28511) );
  OR2_X1 U35359 ( .A1(n28531), .A2(n64809), .Z(n16235) );
  NAND2_X1 U35360 ( .A1(n22115), .A2(n62083), .ZN(n17723) );
  NAND2_X1 U35362 ( .A1(n15953), .A2(n27122), .ZN(n17724) );
  NAND2_X1 U35363 ( .A1(n39007), .A2(n18856), .ZN(n39850) );
  INV_X1 U35364 ( .I(n41234), .ZN(n39852) );
  INV_X1 U35366 ( .I(n40126), .ZN(n20245) );
  NOR3_X1 U35369 ( .A1(n40052), .A2(n18649), .A3(n40337), .ZN(n40053) );
  NOR2_X1 U35370 ( .A1(n39110), .A2(n23932), .ZN(n39115) );
  INV_X1 U35372 ( .I(n61712), .ZN(n39109) );
  NAND2_X1 U35373 ( .A1(n41189), .A2(n64858), .ZN(n22728) );
  NOR2_X1 U35374 ( .A1(n21355), .A2(n21354), .ZN(n21374) );
  NAND2_X1 U35375 ( .A1(n40518), .A2(n40519), .ZN(n21355) );
  NAND2_X1 U35376 ( .A1(n41163), .A2(n10452), .ZN(n39068) );
  NAND2_X1 U35378 ( .A1(n40528), .A2(n40617), .ZN(n25140) );
  NAND2_X1 U35380 ( .A1(n61435), .A2(n41944), .ZN(n41302) );
  INV_X1 U35381 ( .I(n40647), .ZN(n22007) );
  NAND3_X1 U35382 ( .A1(n40723), .A2(n62175), .A3(n22304), .ZN(n17576) );
  NOR3_X1 U35383 ( .A1(n57462), .A2(n40728), .A3(n41197), .ZN(n40629) );
  OAI21_X1 U35384 ( .A1(n41022), .A2(n60166), .B(n17450), .ZN(n16462) );
  AND3_X1 U35385 ( .A1(n38768), .A2(n38767), .A3(n38766), .Z(n15899) );
  NAND2_X1 U35386 ( .A1(n9802), .A2(n16962), .ZN(n40335) );
  AOI22_X1 U35387 ( .A1(n1736), .A2(n40338), .B1(n40339), .B2(n25511), .ZN(
        n40340) );
  NAND2_X1 U35388 ( .A1(n40503), .A2(n1275), .ZN(n19295) );
  NAND3_X1 U35390 ( .A1(n40004), .A2(n41375), .A3(n41382), .ZN(n39822) );
  OAI21_X1 U35391 ( .A1(n61638), .A2(n39821), .B(n39820), .ZN(n23971) );
  NAND2_X1 U35392 ( .A1(n10294), .A2(n39994), .ZN(n39826) );
  AOI21_X1 U35393 ( .A1(n41845), .A2(n41844), .B(n58307), .ZN(n41846) );
  NAND2_X1 U35394 ( .A1(n42526), .A2(n1273), .ZN(n19675) );
  AOI21_X1 U35395 ( .A1(n1273), .A2(n21520), .B(n41838), .ZN(n24751) );
  NAND2_X1 U35396 ( .A1(n64986), .A2(n23501), .ZN(n21520) );
  NAND2_X1 U35397 ( .A1(n39959), .A2(n16292), .ZN(n18411) );
  NAND2_X1 U35399 ( .A1(n16071), .A2(n26941), .ZN(n19339) );
  INV_X1 U35400 ( .I(n26985), .ZN(n25620) );
  NAND2_X1 U35402 ( .A1(n27108), .A2(n64481), .ZN(n25801) );
  AOI21_X1 U35403 ( .A1(n30654), .A2(n30659), .B(n17903), .ZN(n30414) );
  AND2_X1 U35405 ( .A1(n25017), .A2(n20714), .Z(n16138) );
  NAND2_X1 U35406 ( .A1(n31244), .A2(n603), .ZN(n24240) );
  INV_X1 U35407 ( .I(n30888), .ZN(n31240) );
  NAND2_X1 U35408 ( .A1(n29144), .A2(n18231), .ZN(n17247) );
  NAND2_X1 U35409 ( .A1(n19967), .A2(n19966), .ZN(n19965) );
  INV_X1 U35410 ( .I(n29496), .ZN(n17788) );
  NAND2_X1 U35411 ( .A1(n19571), .A2(n29494), .ZN(n29495) );
  NOR3_X1 U35412 ( .A1(n30651), .A2(n30333), .A3(n62285), .ZN(n28710) );
  NAND2_X1 U35413 ( .A1(n26619), .A2(n26653), .ZN(n22948) );
  OR2_X1 U35414 ( .A1(n26620), .A2(n21132), .Z(n16253) );
  NAND2_X1 U35415 ( .A1(n23071), .A2(n21132), .ZN(n26615) );
  NAND2_X1 U35418 ( .A1(n29222), .A2(n30285), .ZN(n30720) );
  NOR2_X1 U35419 ( .A1(n10629), .A2(n59798), .ZN(n21876) );
  NAND2_X1 U35420 ( .A1(n29461), .A2(n61421), .ZN(n28731) );
  NAND2_X1 U35421 ( .A1(n21601), .A2(n27404), .ZN(n21631) );
  NOR2_X1 U35422 ( .A1(n27093), .A2(n16222), .ZN(n22964) );
  INV_X1 U35424 ( .I(n23837), .ZN(n16425) );
  OAI21_X1 U35426 ( .A1(n28462), .A2(n26793), .B(n28617), .ZN(n17527) );
  INV_X1 U35429 ( .I(n28717), .ZN(n24164) );
  NAND2_X1 U35433 ( .A1(n41350), .A2(n60706), .ZN(n41348) );
  OAI21_X1 U35438 ( .A1(n19112), .A2(n16154), .B(n25666), .ZN(n21645) );
  OAI21_X1 U35441 ( .A1(n38498), .A2(n22523), .B(n17965), .ZN(n36108) );
  NAND2_X1 U35443 ( .A1(n41888), .A2(n2325), .ZN(n19439) );
  NAND2_X1 U35446 ( .A1(n39901), .A2(n18278), .ZN(n18043) );
  NAND2_X1 U35447 ( .A1(n41463), .A2(n41462), .ZN(n21349) );
  AOI21_X1 U35450 ( .A1(n13357), .A2(n41145), .B(n40713), .ZN(n23381) );
  NAND2_X1 U35451 ( .A1(n20601), .A2(n20602), .ZN(n41766) );
  NAND2_X1 U35453 ( .A1(n43513), .A2(n43504), .ZN(n43507) );
  NAND2_X1 U35455 ( .A1(n42281), .A2(n17981), .ZN(n41937) );
  INV_X1 U35456 ( .I(n60525), .ZN(n32282) );
  NOR2_X1 U35457 ( .A1(n29952), .A2(n29951), .ZN(n25370) );
  NAND2_X1 U35459 ( .A1(n29063), .A2(n21095), .ZN(n17000) );
  AOI21_X1 U35460 ( .A1(n27102), .A2(n27101), .B(n27100), .ZN(n27104) );
  NOR2_X1 U35462 ( .A1(n30658), .A2(n30638), .ZN(n30646) );
  OAI21_X1 U35464 ( .A1(n27117), .A2(n12421), .B(n26609), .ZN(n17780) );
  NOR2_X1 U35466 ( .A1(n26601), .A2(n26600), .ZN(n18760) );
  NAND2_X1 U35467 ( .A1(n30816), .A2(n30815), .ZN(n23137) );
  NAND2_X1 U35468 ( .A1(n25533), .A2(n29835), .ZN(n18906) );
  NOR2_X1 U35469 ( .A1(n30808), .A2(n30807), .ZN(n25533) );
  NOR2_X1 U35471 ( .A1(n30809), .A2(n30812), .ZN(n18905) );
  NAND2_X1 U35472 ( .A1(n30813), .A2(n30812), .ZN(n26138) );
  OAI21_X1 U35477 ( .A1(n1719), .A2(n43979), .B(n21800), .ZN(n43981) );
  OAI22_X1 U35478 ( .A1(n21566), .A2(n43988), .B1(n43985), .B2(n43986), .ZN(
        n20987) );
  INV_X1 U35483 ( .I(n43508), .ZN(n24494) );
  NOR2_X1 U35484 ( .A1(n43506), .A2(n43518), .ZN(n24492) );
  NAND2_X1 U35485 ( .A1(n30452), .A2(n17268), .ZN(n19026) );
  OAI22_X1 U35486 ( .A1(n18234), .A2(n13810), .B1(n30679), .B2(n30684), .ZN(
        n18233) );
  INV_X1 U35487 ( .I(n16398), .ZN(n16395) );
  NAND3_X1 U35489 ( .A1(n41702), .A2(n65228), .A3(n22367), .ZN(n25373) );
  NOR2_X1 U35490 ( .A1(n41328), .A2(n42694), .ZN(n19720) );
  OAI22_X1 U35491 ( .A1(n41329), .A2(n42381), .B1(n41972), .B2(n42703), .ZN(
        n19719) );
  INV_X1 U35496 ( .I(n17736), .ZN(n44372) );
  NOR2_X1 U35497 ( .A1(n47288), .A2(n47593), .ZN(n21418) );
  NAND2_X1 U35498 ( .A1(n62247), .A2(n59406), .ZN(n25046) );
  INV_X1 U35501 ( .I(n48102), .ZN(n45368) );
  AOI22_X1 U35502 ( .A1(n19533), .A2(n47302), .B1(n46023), .B2(n24047), .ZN(
        n19532) );
  NAND2_X1 U35503 ( .A1(n33440), .A2(n22226), .ZN(n16421) );
  AOI21_X1 U35508 ( .A1(n44858), .A2(n24290), .B(n25557), .ZN(n44859) );
  INV_X1 U35509 ( .I(n47901), .ZN(n44840) );
  INV_X1 U35510 ( .I(n21705), .ZN(n17366) );
  NAND2_X1 U35511 ( .A1(n63294), .A2(n20832), .ZN(n45080) );
  NAND2_X1 U35513 ( .A1(n47634), .A2(n14473), .ZN(n47359) );
  NAND2_X1 U35515 ( .A1(n48490), .A2(n48585), .ZN(n48492) );
  NAND2_X1 U35516 ( .A1(n48484), .A2(n48481), .ZN(n21548) );
  NAND2_X1 U35521 ( .A1(n46100), .A2(n46099), .ZN(n16840) );
  NAND2_X1 U35522 ( .A1(n48649), .A2(n46103), .ZN(n46109) );
  AOI21_X1 U35528 ( .A1(n47282), .A2(n47283), .B(n19176), .ZN(n45159) );
  NAND2_X1 U35529 ( .A1(n11172), .A2(n1638), .ZN(n48307) );
  NAND2_X1 U35531 ( .A1(n46992), .A2(n48667), .ZN(n26085) );
  AOI21_X1 U35532 ( .A1(n21977), .A2(n21975), .B(n47249), .ZN(n21974) );
  NOR2_X1 U35534 ( .A1(n406), .A2(n49525), .ZN(n24802) );
  NOR2_X1 U35535 ( .A1(n33418), .A2(n34615), .ZN(n21109) );
  OAI22_X1 U35536 ( .A1(n33419), .A2(n19610), .B1(n33975), .B2(n34039), .ZN(
        n33425) );
  OAI21_X1 U35537 ( .A1(n47616), .A2(n45210), .B(n45209), .ZN(n45211) );
  NOR2_X1 U35539 ( .A1(n48223), .A2(n21567), .ZN(n48227) );
  NAND2_X1 U35540 ( .A1(n48578), .A2(n59269), .ZN(n18221) );
  NOR2_X1 U35544 ( .A1(n48071), .A2(n45791), .ZN(n17682) );
  NOR2_X1 U35545 ( .A1(n19294), .A2(n64167), .ZN(n17684) );
  NOR2_X1 U35547 ( .A1(n22457), .A2(n16411), .ZN(n44790) );
  INV_X1 U35548 ( .I(n18625), .ZN(n47969) );
  OAI21_X1 U35549 ( .A1(n47271), .A2(n47579), .B(n22009), .ZN(n22008) );
  INV_X1 U35550 ( .I(n1643), .ZN(n50303) );
  INV_X1 U35552 ( .I(n25773), .ZN(n49427) );
  NAND2_X1 U35555 ( .A1(n48825), .A2(n48064), .ZN(n19899) );
  NAND2_X1 U35556 ( .A1(n24582), .A2(n1627), .ZN(n19445) );
  NAND2_X1 U35559 ( .A1(n11314), .A2(n10874), .ZN(n49409) );
  NAND3_X1 U35560 ( .A1(n18756), .A2(n48665), .A3(n48194), .ZN(n17008) );
  OAI21_X1 U35562 ( .A1(n46431), .A2(n48136), .B(n23663), .ZN(n46458) );
  AOI21_X1 U35563 ( .A1(n23021), .A2(n48136), .B(n48475), .ZN(n23663) );
  INV_X1 U35564 ( .I(n48471), .ZN(n23021) );
  NAND2_X1 U35569 ( .A1(n23612), .A2(n19867), .ZN(n20901) );
  INV_X1 U35571 ( .I(n47306), .ZN(n18843) );
  NAND2_X1 U35573 ( .A1(n20199), .A2(n1637), .ZN(n49575) );
  AND2_X1 U35574 ( .A1(n18142), .A2(n50077), .Z(n15990) );
  NOR2_X1 U35576 ( .A1(n19107), .A2(n16411), .ZN(n16908) );
  NOR3_X1 U35577 ( .A1(n48004), .A2(n49512), .A3(n58975), .ZN(n18430) );
  INV_X1 U35579 ( .I(n51553), .ZN(n22219) );
  NAND2_X1 U35581 ( .A1(n1612), .A2(n57022), .ZN(n16772) );
  NOR2_X1 U35582 ( .A1(n53212), .A2(n23796), .ZN(n16770) );
  NOR2_X1 U35584 ( .A1(n54589), .A2(n51705), .ZN(n51706) );
  NAND2_X1 U35585 ( .A1(n54596), .A2(n23736), .ZN(n51702) );
  OAI22_X1 U35587 ( .A1(n55914), .A2(n55911), .B1(n55912), .B2(n13025), .ZN(
        n24142) );
  INV_X1 U35588 ( .I(n54016), .ZN(n16866) );
  NAND2_X1 U35589 ( .A1(n51864), .A2(n53881), .ZN(n16865) );
  NAND2_X1 U35591 ( .A1(n56374), .A2(n56660), .ZN(n21852) );
  INV_X1 U35592 ( .I(n55271), .ZN(n55259) );
  OAI21_X1 U35594 ( .A1(n16117), .A2(n55693), .B(n19971), .ZN(n55701) );
  NOR2_X1 U35595 ( .A1(n53451), .A2(n53223), .ZN(n16436) );
  NAND3_X1 U35598 ( .A1(n26095), .A2(n2198), .A3(n54433), .ZN(n26096) );
  NAND2_X1 U35600 ( .A1(n55658), .A2(n19958), .ZN(n24403) );
  OAI21_X1 U35601 ( .A1(n51903), .A2(n1369), .B(n16621), .ZN(n16620) );
  NAND3_X1 U35603 ( .A1(n53835), .A2(n64978), .A3(n60794), .ZN(n54496) );
  OAI21_X1 U35608 ( .A1(n13815), .A2(n53878), .B(n53880), .ZN(n51714) );
  NAND2_X1 U35609 ( .A1(n15929), .A2(n9137), .ZN(n51713) );
  NAND2_X1 U35611 ( .A1(n64978), .A2(n17057), .ZN(n54309) );
  NAND2_X1 U35613 ( .A1(n54318), .A2(n21135), .ZN(n54319) );
  INV_X1 U35614 ( .I(n64978), .ZN(n54311) );
  AOI22_X1 U35616 ( .A1(n51864), .A2(n16175), .B1(n54026), .B2(n54346), .ZN(
        n21696) );
  INV_X1 U35617 ( .I(n21225), .ZN(n52251) );
  NOR3_X1 U35619 ( .A1(n55436), .A2(n55434), .A3(n14225), .ZN(n25719) );
  NAND2_X1 U35620 ( .A1(n54818), .A2(n15761), .ZN(n21051) );
  NOR2_X1 U35621 ( .A1(n53424), .A2(n53423), .ZN(n22689) );
  OAI21_X1 U35623 ( .A1(n21747), .A2(n53042), .B(n23206), .ZN(n21746) );
  NAND2_X1 U35624 ( .A1(n53807), .A2(n53809), .ZN(n21747) );
  NOR2_X1 U35627 ( .A1(n51258), .A2(n56229), .ZN(n16332) );
  NAND2_X1 U35628 ( .A1(n54784), .A2(n54949), .ZN(n25502) );
  INV_X1 U35629 ( .I(n54794), .ZN(n54979) );
  NAND2_X1 U35630 ( .A1(n24032), .A2(n61627), .ZN(n56319) );
  NOR2_X1 U35631 ( .A1(n53237), .A2(n52872), .ZN(n52876) );
  NOR2_X1 U35632 ( .A1(n23272), .A2(n51965), .ZN(n23271) );
  NOR2_X1 U35633 ( .A1(n56583), .A2(n56584), .ZN(n56597) );
  NOR2_X1 U35636 ( .A1(n49873), .A2(n54102), .ZN(n17289) );
  AOI21_X1 U35637 ( .A1(n54611), .A2(n54612), .B(n19494), .ZN(n19493) );
  NOR2_X1 U35638 ( .A1(n21998), .A2(n21997), .ZN(n21996) );
  NOR2_X1 U35640 ( .A1(n26118), .A2(n22518), .ZN(n26117) );
  NAND3_X1 U35641 ( .A1(n55264), .A2(n55270), .A3(n65101), .ZN(n54841) );
  NAND2_X1 U35643 ( .A1(n53887), .A2(n53886), .ZN(n18620) );
  NAND2_X1 U35644 ( .A1(n54345), .A2(n54344), .ZN(n17037) );
  NAND2_X1 U35645 ( .A1(n56476), .A2(n23920), .ZN(n56483) );
  NAND2_X1 U35648 ( .A1(n55439), .A2(n18256), .ZN(n21274) );
  NAND2_X1 U35652 ( .A1(n64788), .A2(n63873), .ZN(n54242) );
  NAND2_X1 U35653 ( .A1(n20570), .A2(n55906), .ZN(n52127) );
  OAI21_X1 U35654 ( .A1(n19133), .A2(n19132), .B(n52049), .ZN(n21411) );
  INV_X2 U35655 ( .I(n56689), .ZN(n56708) );
  NOR2_X1 U35657 ( .A1(n20319), .A2(n53533), .ZN(n19485) );
  NOR2_X1 U35658 ( .A1(n53738), .A2(n24326), .ZN(n53712) );
  NOR2_X1 U35659 ( .A1(n53726), .A2(n25011), .ZN(n24326) );
  NAND3_X1 U35660 ( .A1(n1260), .A2(n22381), .A3(n55966), .ZN(n19030) );
  NAND2_X1 U35661 ( .A1(n53755), .A2(n53728), .ZN(n50830) );
  INV_X1 U35662 ( .I(n33172), .ZN(n22215) );
  INV_X1 U35663 ( .I(n31858), .ZN(n18962) );
  INV_X1 U35664 ( .I(n34438), .ZN(n16906) );
  NAND2_X1 U35666 ( .A1(n18390), .A2(n33995), .ZN(n17048) );
  INV_X1 U35667 ( .I(n64234), .ZN(n33969) );
  NOR2_X1 U35668 ( .A1(n34190), .A2(n118), .ZN(n23177) );
  NAND2_X1 U35670 ( .A1(n34433), .A2(n35322), .ZN(n34435) );
  NAND3_X1 U35672 ( .A1(n34148), .A2(n19435), .A3(n34147), .ZN(n34154) );
  AOI22_X1 U35673 ( .A1(n24287), .A2(n22601), .B1(n20923), .B2(n23757), .ZN(
        n34153) );
  OAI22_X1 U35675 ( .A1(n26242), .A2(n34713), .B1(n35303), .B2(n35309), .ZN(
        n34716) );
  NAND3_X1 U35676 ( .A1(n12338), .A2(n34670), .A3(n34669), .ZN(n34672) );
  NOR2_X1 U35678 ( .A1(n30960), .A2(n21041), .ZN(n21040) );
  NOR2_X1 U35680 ( .A1(n18440), .A2(n34306), .ZN(n17070) );
  NAND3_X1 U35681 ( .A1(n34559), .A2(n34020), .A3(n20785), .ZN(n17552) );
  NAND2_X1 U35682 ( .A1(n33518), .A2(n23125), .ZN(n34029) );
  INV_X1 U35684 ( .I(n34307), .ZN(n34312) );
  NAND2_X1 U35686 ( .A1(n897), .A2(n34385), .ZN(n18273) );
  INV_X1 U35688 ( .I(n34965), .ZN(n34960) );
  NAND2_X1 U35690 ( .A1(n32949), .A2(n21317), .ZN(n32950) );
  NOR2_X1 U35691 ( .A1(n21317), .A2(n20157), .ZN(n22023) );
  NAND2_X1 U35692 ( .A1(n34353), .A2(n34358), .ZN(n32932) );
  NAND3_X1 U35696 ( .A1(n21407), .A2(n33945), .A3(n33949), .ZN(n32792) );
  NOR3_X1 U35697 ( .A1(n139), .A2(n1812), .A3(n32795), .ZN(n21407) );
  NAND3_X1 U35699 ( .A1(n16087), .A2(n34753), .A3(n21538), .ZN(n34754) );
  OAI21_X1 U35702 ( .A1(n35711), .A2(n35842), .B(n21252), .ZN(n35719) );
  NAND3_X1 U35704 ( .A1(n34358), .A2(n32927), .A3(n34246), .ZN(n32426) );
  NOR2_X1 U35705 ( .A1(n31609), .A2(n19925), .ZN(n19464) );
  OAI21_X1 U35706 ( .A1(n34602), .A2(n24273), .B(n34603), .ZN(n19602) );
  INV_X1 U35707 ( .I(n18877), .ZN(n36827) );
  NOR2_X1 U35708 ( .A1(n34724), .A2(n1536), .ZN(n19017) );
  INV_X1 U35710 ( .I(n32792), .ZN(n20676) );
  NAND2_X1 U35711 ( .A1(n33715), .A2(n15754), .ZN(n35961) );
  NAND2_X1 U35712 ( .A1(n34952), .A2(n34564), .ZN(n33479) );
  INV_X1 U35713 ( .I(n35450), .ZN(n36271) );
  NAND2_X1 U35715 ( .A1(n36026), .A2(n36020), .ZN(n36037) );
  NAND2_X1 U35716 ( .A1(n33821), .A2(n19789), .ZN(n24371) );
  OAI21_X1 U35717 ( .A1(n19772), .A2(n57337), .B(n23556), .ZN(n18366) );
  NAND2_X1 U35718 ( .A1(n61090), .A2(n17254), .ZN(n35633) );
  INV_X1 U35719 ( .I(n20182), .ZN(n35635) );
  INV_X1 U35720 ( .I(n37051), .ZN(n35095) );
  AOI21_X1 U35722 ( .A1(n35327), .A2(n35326), .B(n35774), .ZN(n21883) );
  INV_X1 U35723 ( .I(n20616), .ZN(n34912) );
  INV_X1 U35724 ( .I(n34907), .ZN(n34906) );
  NOR2_X1 U35730 ( .A1(n34817), .A2(n34815), .ZN(n34287) );
  NOR2_X1 U35731 ( .A1(n35961), .A2(n35548), .ZN(n35975) );
  INV_X1 U35734 ( .I(n34937), .ZN(n36720) );
  INV_X1 U35735 ( .I(n36766), .ZN(n21768) );
  INV_X1 U35736 ( .I(n36048), .ZN(n21769) );
  INV_X1 U35737 ( .I(n18705), .ZN(n21773) );
  INV_X1 U35738 ( .I(n32943), .ZN(n21380) );
  OAI22_X1 U35742 ( .A1(n33449), .A2(n64101), .B1(n33458), .B2(n36945), .ZN(
        n24310) );
  OAI21_X1 U35744 ( .A1(n37343), .A2(n37342), .B(n37341), .ZN(n37344) );
  NOR2_X1 U35746 ( .A1(n60297), .A2(n22317), .ZN(n34374) );
  NAND2_X1 U35748 ( .A1(n16566), .A2(n37116), .ZN(n16565) );
  NOR2_X1 U35749 ( .A1(n19677), .A2(n16563), .ZN(n16562) );
  NAND2_X1 U35751 ( .A1(n37268), .A2(n17243), .ZN(n34847) );
  NAND2_X1 U35754 ( .A1(n63817), .A2(n4541), .ZN(n34455) );
  INV_X1 U35755 ( .I(n34432), .ZN(n25187) );
  NAND2_X1 U35756 ( .A1(n20571), .A2(n25366), .ZN(n34819) );
  AOI21_X1 U35757 ( .A1(n1772), .A2(n21913), .B(n37051), .ZN(n21912) );
  NAND3_X1 U35758 ( .A1(n37050), .A2(n1793), .A3(n35096), .ZN(n21913) );
  NAND2_X1 U35759 ( .A1(n31307), .A2(n37055), .ZN(n25334) );
  NAND2_X1 U35760 ( .A1(n1793), .A2(n35096), .ZN(n31303) );
  NOR2_X1 U35763 ( .A1(n37044), .A2(n31306), .ZN(n22578) );
  NAND2_X1 U35764 ( .A1(n36046), .A2(n36774), .ZN(n34008) );
  NAND2_X1 U35765 ( .A1(n37333), .A2(n37181), .ZN(n24659) );
  AOI21_X1 U35767 ( .A1(n36728), .A2(n59147), .B(n36729), .ZN(n36206) );
  NAND2_X1 U35769 ( .A1(n35496), .A2(n35495), .ZN(n19608) );
  NAND2_X1 U35772 ( .A1(n36904), .A2(n58220), .ZN(n36905) );
  NAND2_X1 U35773 ( .A1(n37419), .A2(n2383), .ZN(n36907) );
  NOR2_X1 U35775 ( .A1(n35277), .A2(n35278), .ZN(n17298) );
  NAND2_X1 U35776 ( .A1(n33547), .A2(n35620), .ZN(n32992) );
  AOI21_X1 U35779 ( .A1(n12863), .A2(n35860), .B(n1417), .ZN(n16664) );
  INV_X1 U35780 ( .I(n23648), .ZN(n35865) );
  NAND2_X1 U35781 ( .A1(n24028), .A2(n36485), .ZN(n21675) );
  NOR2_X1 U35782 ( .A1(n1525), .A2(n1782), .ZN(n21671) );
  INV_X1 U35783 ( .I(n38708), .ZN(n38207) );
  OAI21_X1 U35784 ( .A1(n34842), .A2(n23842), .B(n17243), .ZN(n34843) );
  NAND2_X1 U35785 ( .A1(n35609), .A2(n36721), .ZN(n21542) );
  NOR3_X1 U35790 ( .A1(n36927), .A2(n36924), .A3(n35506), .ZN(n25850) );
  OAI21_X1 U35791 ( .A1(n13403), .A2(n17243), .B(n37268), .ZN(n36083) );
  NAND2_X1 U35793 ( .A1(n37136), .A2(n23842), .ZN(n36087) );
  INV_X1 U35795 ( .I(n38333), .ZN(n21687) );
  NOR2_X1 U35797 ( .A1(n20255), .A2(n20254), .ZN(n20253) );
  NOR2_X1 U35800 ( .A1(n35151), .A2(n16639), .ZN(n16638) );
  INV_X1 U35801 ( .I(n34818), .ZN(n19690) );
  INV_X1 U35802 ( .I(n19813), .ZN(n19633) );
  OAI21_X1 U35803 ( .A1(n23648), .A2(n23647), .B(n36334), .ZN(n35866) );
  OAI22_X1 U35804 ( .A1(n29311), .A2(n20093), .B1(n28854), .B2(n27360), .ZN(
        n25156) );
  NAND2_X1 U35805 ( .A1(n30165), .A2(n30691), .ZN(n29030) );
  NAND2_X1 U35806 ( .A1(n20918), .A2(n31054), .ZN(n29026) );
  NAND2_X1 U35807 ( .A1(n10125), .A2(n63094), .ZN(n27657) );
  NAND2_X1 U35808 ( .A1(n29178), .A2(n24419), .ZN(n16845) );
  NAND3_X1 U35809 ( .A1(n28516), .A2(n27850), .A3(n27717), .ZN(n16492) );
  NAND2_X1 U35810 ( .A1(n1569), .A2(n27852), .ZN(n26024) );
  NOR2_X1 U35812 ( .A1(n19138), .A2(n19139), .ZN(n18059) );
  INV_X1 U35813 ( .I(n18049), .ZN(n19044) );
  INV_X1 U35814 ( .I(n38321), .ZN(n37702) );
  NOR2_X1 U35815 ( .A1(n36231), .A2(n18352), .ZN(n36242) );
  INV_X1 U35820 ( .I(n39303), .ZN(n17975) );
  INV_X1 U35821 ( .I(n19303), .ZN(n38857) );
  NOR2_X1 U35823 ( .A1(n36615), .A2(n37222), .ZN(n20680) );
  INV_X1 U35824 ( .I(n39759), .ZN(n25409) );
  OAI21_X1 U35825 ( .A1(n9098), .A2(n266), .B(n22177), .ZN(n27293) );
  NOR2_X1 U35826 ( .A1(n29138), .A2(n29142), .ZN(n22177) );
  NAND2_X1 U35827 ( .A1(n27272), .A2(n24967), .ZN(n19678) );
  NAND2_X1 U35828 ( .A1(n13672), .A2(n20721), .ZN(n27162) );
  NOR2_X1 U35829 ( .A1(n22205), .A2(n97), .ZN(n25733) );
  NAND2_X1 U35830 ( .A1(n27387), .A2(n28239), .ZN(n22205) );
  OAI21_X1 U35831 ( .A1(n27382), .A2(n28071), .B(n27381), .ZN(n27383) );
  INV_X1 U35832 ( .I(n28241), .ZN(n27382) );
  NAND2_X1 U35834 ( .A1(n26431), .A2(n28534), .ZN(n26801) );
  INV_X1 U35835 ( .I(n28516), .ZN(n28520) );
  NOR2_X1 U35836 ( .A1(n27247), .A2(n28527), .ZN(n26003) );
  NAND2_X1 U35837 ( .A1(n40970), .A2(n40962), .ZN(n38604) );
  NOR2_X1 U35839 ( .A1(n39099), .A2(n59255), .ZN(n21354) );
  NOR2_X1 U35840 ( .A1(n42207), .A2(n23501), .ZN(n22248) );
  NAND3_X1 U35841 ( .A1(n41871), .A2(n38136), .A3(n42519), .ZN(n20074) );
  NAND2_X1 U35844 ( .A1(n18076), .A2(n36958), .ZN(n18812) );
  NAND2_X1 U35845 ( .A1(n41375), .A2(n10074), .ZN(n40425) );
  INV_X1 U35846 ( .I(n39779), .ZN(n17888) );
  NAND2_X1 U35847 ( .A1(n40712), .A2(n41149), .ZN(n40710) );
  NOR2_X1 U35850 ( .A1(n22832), .A2(n22638), .ZN(n41449) );
  NOR2_X1 U35851 ( .A1(n59961), .A2(n18622), .ZN(n39983) );
  NOR2_X1 U35852 ( .A1(n31279), .A2(n6317), .ZN(n31167) );
  INV_X1 U35854 ( .I(n31118), .ZN(n30386) );
  OAI21_X1 U35855 ( .A1(n1857), .A2(n1853), .B(n30871), .ZN(n19524) );
  OAI22_X1 U35856 ( .A1(n30586), .A2(n30585), .B1(n495), .B2(n22579), .ZN(
        n25236) );
  NAND3_X1 U35858 ( .A1(n28261), .A2(n62005), .A3(n29173), .ZN(n17918) );
  NOR2_X1 U35859 ( .A1(n23716), .A2(n23166), .ZN(n27949) );
  NOR2_X1 U35862 ( .A1(n28549), .A2(n29187), .ZN(n17279) );
  NAND2_X1 U35863 ( .A1(n60885), .A2(n17813), .ZN(n27963) );
  NOR2_X1 U35864 ( .A1(n28517), .A2(n25858), .ZN(n27708) );
  INV_X1 U35865 ( .I(n61729), .ZN(n29016) );
  NOR2_X1 U35866 ( .A1(n21614), .A2(n17418), .ZN(n21628) );
  INV_X1 U35867 ( .I(n27403), .ZN(n21632) );
  NOR2_X1 U35869 ( .A1(n19872), .A2(n30585), .ZN(n30378) );
  OAI21_X1 U35870 ( .A1(n23940), .A2(n22643), .B(n22952), .ZN(n26672) );
  NOR3_X1 U35872 ( .A1(n57424), .A2(n28855), .A3(n27449), .ZN(n28164) );
  NOR4_X1 U35873 ( .A1(n27448), .A2(n57424), .A3(n9987), .A4(n27447), .ZN(
        n27453) );
  NOR2_X1 U35874 ( .A1(n28678), .A2(n30743), .ZN(n18871) );
  NAND2_X1 U35876 ( .A1(n30702), .A2(n21019), .ZN(n30149) );
  INV_X1 U35877 ( .I(n39828), .ZN(n26132) );
  INV_X1 U35878 ( .I(n42266), .ZN(n40581) );
  NAND2_X1 U35879 ( .A1(n12806), .A2(n41425), .ZN(n22758) );
  NAND2_X1 U35880 ( .A1(n40818), .A2(n38345), .ZN(n17093) );
  AOI21_X1 U35881 ( .A1(n40403), .A2(n41422), .B(n22168), .ZN(n38928) );
  AOI22_X1 U35882 ( .A1(n41422), .A2(n38935), .B1(n41425), .B2(n1739), .ZN(
        n20820) );
  INV_X1 U35883 ( .I(n41511), .ZN(n40941) );
  NAND3_X1 U35884 ( .A1(n62107), .A2(n61417), .A3(n12158), .ZN(n40007) );
  NAND2_X1 U35886 ( .A1(n21036), .A2(n40355), .ZN(n19112) );
  NAND2_X1 U35888 ( .A1(n39911), .A2(n39910), .ZN(n39917) );
  NAND3_X1 U35889 ( .A1(n40228), .A2(n40291), .A3(n64613), .ZN(n39910) );
  NAND2_X1 U35891 ( .A1(n41646), .A2(n24792), .ZN(n41649) );
  INV_X1 U35893 ( .I(n18407), .ZN(n43435) );
  INV_X1 U35894 ( .I(n40841), .ZN(n24606) );
  NAND2_X1 U35896 ( .A1(n41412), .A2(n41402), .ZN(n21001) );
  NOR2_X1 U35897 ( .A1(n41031), .A2(n40517), .ZN(n38494) );
  OR2_X1 U35898 ( .A1(n41168), .A2(n14462), .Z(n25227) );
  NAND2_X1 U35899 ( .A1(n17450), .A2(n37532), .ZN(n38425) );
  NAND2_X1 U35902 ( .A1(n15584), .A2(n41400), .ZN(n20889) );
  NOR2_X1 U35903 ( .A1(n61417), .A2(n41382), .ZN(n17020) );
  NOR2_X1 U35904 ( .A1(n41802), .A2(n41801), .ZN(n17295) );
  NAND2_X1 U35905 ( .A1(n40379), .A2(n22638), .ZN(n19385) );
  AOI21_X1 U35908 ( .A1(n27390), .A2(n7499), .B(n29153), .ZN(n26749) );
  NAND2_X1 U35909 ( .A1(n30224), .A2(n22416), .ZN(n30839) );
  NOR2_X1 U35911 ( .A1(n30214), .A2(n1869), .ZN(n21775) );
  NOR2_X1 U35912 ( .A1(n30223), .A2(n30840), .ZN(n21528) );
  INV_X1 U35913 ( .I(n30217), .ZN(n21777) );
  NAND3_X1 U35914 ( .A1(n3426), .A2(n770), .A3(n7040), .ZN(n21778) );
  NOR2_X1 U35915 ( .A1(n16800), .A2(n63691), .ZN(n30219) );
  NAND2_X1 U35916 ( .A1(n30517), .A2(n1351), .ZN(n18462) );
  OAI22_X1 U35917 ( .A1(n28252), .A2(n60020), .B1(n24498), .B2(n22095), .ZN(
        n28253) );
  NOR2_X1 U35918 ( .A1(n23269), .A2(n4257), .ZN(n31282) );
  NAND2_X1 U35919 ( .A1(n31238), .A2(n31239), .ZN(n24239) );
  NOR2_X1 U35922 ( .A1(n19255), .A2(n1435), .ZN(n29887) );
  NAND2_X1 U35924 ( .A1(n27614), .A2(n18747), .ZN(n26598) );
  NOR2_X1 U35925 ( .A1(n26599), .A2(n22273), .ZN(n26600) );
  OAI21_X1 U35927 ( .A1(n24172), .A2(n25240), .B(n25238), .ZN(n25237) );
  NAND2_X1 U35928 ( .A1(n5768), .A2(n30585), .ZN(n25240) );
  NOR2_X1 U35929 ( .A1(n59810), .A2(n1316), .ZN(n25239) );
  NAND2_X1 U35930 ( .A1(n23829), .A2(n9719), .ZN(n27438) );
  INV_X1 U35933 ( .I(n26485), .ZN(n25454) );
  NAND2_X1 U35935 ( .A1(n28844), .A2(n28845), .ZN(n19547) );
  NAND2_X1 U35936 ( .A1(n27493), .A2(n24947), .ZN(n24785) );
  NOR2_X1 U35938 ( .A1(n30558), .A2(n31086), .ZN(n31080) );
  NAND2_X1 U35940 ( .A1(n59841), .A2(n28209), .ZN(n30581) );
  NAND2_X1 U35942 ( .A1(n24975), .A2(n29805), .ZN(n24974) );
  NAND3_X1 U35943 ( .A1(n20123), .A2(n29024), .A3(n21019), .ZN(n20122) );
  INV_X1 U35944 ( .I(n31033), .ZN(n20123) );
  AOI21_X1 U35945 ( .A1(n27484), .A2(n27543), .B(n15999), .ZN(n27488) );
  OAI21_X1 U35949 ( .A1(n16648), .A2(n30787), .B(n30786), .ZN(n16647) );
  NAND2_X1 U35951 ( .A1(n29878), .A2(n20028), .ZN(n29730) );
  NAND2_X1 U35952 ( .A1(n30164), .A2(n31054), .ZN(n30166) );
  INV_X1 U35954 ( .I(n42438), .ZN(n40065) );
  NAND2_X1 U35957 ( .A1(n16527), .A2(n4274), .ZN(n41491) );
  NOR2_X1 U35958 ( .A1(n40956), .A2(n40528), .ZN(n40530) );
  NAND2_X1 U35959 ( .A1(n12089), .A2(n61743), .ZN(n19844) );
  NOR2_X1 U35960 ( .A1(n43155), .A2(n43156), .ZN(n20452) );
  NAND2_X1 U35963 ( .A1(n43130), .A2(n43270), .ZN(n43122) );
  NOR2_X1 U35964 ( .A1(n43042), .A2(n43043), .ZN(n19955) );
  NOR2_X1 U35965 ( .A1(n43041), .A2(n41583), .ZN(n19954) );
  NOR2_X1 U35966 ( .A1(n22087), .A2(n22553), .ZN(n43635) );
  INV_X1 U35968 ( .I(n39789), .ZN(n18746) );
  NOR2_X1 U35969 ( .A1(n43273), .A2(n16671), .ZN(n16670) );
  NAND2_X1 U35970 ( .A1(n43120), .A2(n2330), .ZN(n16671) );
  INV_X1 U35971 ( .I(n57178), .ZN(n43217) );
  AOI22_X1 U35973 ( .A1(n18796), .A2(n58850), .B1(n18793), .B2(n43445), .ZN(
        n18792) );
  NOR2_X1 U35975 ( .A1(n43444), .A2(n18794), .ZN(n18793) );
  NOR2_X1 U35977 ( .A1(n20220), .A2(n12089), .ZN(n20219) );
  NOR2_X1 U35978 ( .A1(n20351), .A2(n21073), .ZN(n20220) );
  NOR2_X1 U35979 ( .A1(n43490), .A2(n43912), .ZN(n20222) );
  NAND2_X1 U35981 ( .A1(n42040), .A2(n42041), .ZN(n22777) );
  INV_X1 U35982 ( .I(n43181), .ZN(n42041) );
  NAND2_X1 U35983 ( .A1(n42914), .A2(n42554), .ZN(n41604) );
  INV_X1 U35985 ( .I(n41547), .ZN(n42742) );
  NAND2_X1 U35986 ( .A1(n42371), .A2(n43444), .ZN(n42942) );
  AOI21_X1 U35987 ( .A1(n39053), .A2(n41412), .B(n41230), .ZN(n39054) );
  NAND2_X1 U35991 ( .A1(n25816), .A2(n62241), .ZN(n41062) );
  OAI21_X1 U35993 ( .A1(n23184), .A2(n60792), .B(n62389), .ZN(n41995) );
  NOR2_X1 U35995 ( .A1(n30022), .A2(n30021), .ZN(n21657) );
  NAND2_X1 U35996 ( .A1(n29268), .A2(n1317), .ZN(n16610) );
  NAND2_X1 U35997 ( .A1(n30296), .A2(n29579), .ZN(n16613) );
  NAND2_X1 U35998 ( .A1(n23988), .A2(n1317), .ZN(n21315) );
  INV_X1 U36002 ( .I(n29331), .ZN(n24263) );
  OAI21_X1 U36003 ( .A1(n29912), .A2(n1844), .B(n17714), .ZN(n17713) );
  NAND2_X1 U36004 ( .A1(n30078), .A2(n29794), .ZN(n28787) );
  AOI21_X1 U36005 ( .A1(n30317), .A2(n16897), .B(n2118), .ZN(n16896) );
  NOR2_X1 U36006 ( .A1(n2119), .A2(n10345), .ZN(n16897) );
  INV_X1 U36007 ( .I(n30326), .ZN(n29272) );
  AOI21_X1 U36008 ( .A1(n30521), .A2(n22877), .B(n62231), .ZN(n17118) );
  NOR3_X1 U36009 ( .A1(n30124), .A2(n22877), .A3(n1872), .ZN(n17117) );
  NAND2_X1 U36010 ( .A1(n60214), .A2(n57790), .ZN(n22873) );
  NAND3_X1 U36014 ( .A1(n30681), .A2(n30244), .A3(n19218), .ZN(n30247) );
  NAND2_X1 U36017 ( .A1(n29736), .A2(n30197), .ZN(n19089) );
  INV_X1 U36018 ( .I(n21876), .ZN(n19087) );
  NAND2_X1 U36020 ( .A1(n21864), .A2(n22799), .ZN(n29738) );
  INV_X1 U36021 ( .I(n30099), .ZN(n21864) );
  NOR2_X1 U36022 ( .A1(n27243), .A2(n27242), .ZN(n25466) );
  AND4_X1 U36024 ( .A1(n25095), .A2(n27803), .A3(n27802), .A4(n29910), .Z(
        n16040) );
  INV_X1 U36025 ( .I(n32611), .ZN(n24756) );
  OAI21_X1 U36027 ( .A1(n42487), .A2(n40319), .B(n40091), .ZN(n16398) );
  INV_X1 U36028 ( .I(n42491), .ZN(n42487) );
  INV_X1 U36029 ( .I(n42138), .ZN(n25235) );
  AOI22_X1 U36032 ( .A1(n17744), .A2(n41348), .B1(n22673), .B2(n43854), .ZN(
        n41352) );
  OAI21_X1 U36033 ( .A1(n43207), .A2(n59650), .B(n23730), .ZN(n41351) );
  INV_X1 U36034 ( .I(n42825), .ZN(n42152) );
  NOR2_X1 U36035 ( .A1(n20602), .A2(n43155), .ZN(n40685) );
  NAND2_X1 U36036 ( .A1(n16473), .A2(n43154), .ZN(n16472) );
  NAND2_X1 U36038 ( .A1(n41988), .A2(n1500), .ZN(n40895) );
  OAI22_X1 U36039 ( .A1(n40887), .A2(n1499), .B1(n1500), .B2(n62435), .ZN(
        n40888) );
  INV_X1 U36041 ( .I(n43446), .ZN(n42051) );
  NOR3_X1 U36042 ( .A1(n42935), .A2(n43449), .A3(n43447), .ZN(n40024) );
  OAI21_X1 U36044 ( .A1(n21644), .A2(n42735), .B(n22417), .ZN(n40371) );
  NOR2_X1 U36045 ( .A1(n42655), .A2(n22418), .ZN(n22417) );
  NAND2_X1 U36046 ( .A1(n1335), .A2(n22282), .ZN(n22418) );
  INV_X1 U36047 ( .I(n17501), .ZN(n41360) );
  NAND2_X1 U36048 ( .A1(n42151), .A2(n60131), .ZN(n41367) );
  AOI22_X1 U36051 ( .A1(n1700), .A2(n42687), .B1(n42688), .B2(n42689), .ZN(
        n42690) );
  INV_X1 U36055 ( .I(n43392), .ZN(n16410) );
  INV_X1 U36056 ( .I(n20243), .ZN(n37832) );
  AND2_X1 U36057 ( .A1(n42018), .A2(n4274), .Z(n16261) );
  NAND2_X1 U36058 ( .A1(n41490), .A2(n16527), .ZN(n22693) );
  INV_X1 U36059 ( .I(n19975), .ZN(n37915) );
  OAI21_X1 U36060 ( .A1(n43317), .A2(n20689), .B(n20688), .ZN(n43329) );
  NAND2_X1 U36061 ( .A1(n41781), .A2(n42169), .ZN(n24623) );
  AOI21_X1 U36062 ( .A1(n57178), .A2(n23811), .B(n16713), .ZN(n25000) );
  OAI21_X1 U36063 ( .A1(n40878), .A2(n64629), .B(n40877), .ZN(n19336) );
  NAND2_X1 U36064 ( .A1(n59394), .A2(n41689), .ZN(n38058) );
  AND2_X1 U36065 ( .A1(n24954), .A2(n29533), .Z(n16291) );
  INV_X1 U36066 ( .I(n25526), .ZN(n24954) );
  AND2_X1 U36067 ( .A1(n29521), .A2(n29860), .Z(n16228) );
  AOI21_X1 U36068 ( .A1(n29514), .A2(n64565), .B(n1838), .ZN(n21209) );
  INV_X1 U36069 ( .I(n63050), .ZN(n18314) );
  INV_X1 U36071 ( .I(n43256), .ZN(n43259) );
  NOR2_X1 U36073 ( .A1(n62264), .A2(n42383), .ZN(n19718) );
  NAND2_X1 U36074 ( .A1(n42699), .A2(n62264), .ZN(n41329) );
  INV_X1 U36075 ( .I(n4546), .ZN(n19268) );
  OAI21_X1 U36076 ( .A1(n42965), .A2(n42964), .B(n42963), .ZN(n17150) );
  NAND2_X1 U36078 ( .A1(n19808), .A2(n19807), .ZN(n41690) );
  AOI21_X1 U36081 ( .A1(n42988), .A2(n43957), .B(n43295), .ZN(n25550) );
  NAND2_X1 U36085 ( .A1(n42587), .A2(n8185), .ZN(n16705) );
  NAND2_X1 U36086 ( .A1(n20380), .A2(n43302), .ZN(n19100) );
  NAND2_X1 U36087 ( .A1(n41764), .A2(n24494), .ZN(n24493) );
  NOR2_X1 U36088 ( .A1(n16554), .A2(n16552), .ZN(n16551) );
  AOI21_X1 U36089 ( .A1(n16553), .A2(n16237), .B(n42865), .ZN(n16552) );
  AOI21_X1 U36090 ( .A1(n41528), .A2(n2160), .B(n41330), .ZN(n40186) );
  INV_X1 U36091 ( .I(n46697), .ZN(n23807) );
  INV_X1 U36092 ( .I(n46520), .ZN(n18648) );
  NAND2_X1 U36094 ( .A1(n46925), .A2(n45954), .ZN(n46059) );
  INV_X1 U36095 ( .I(n31763), .ZN(n22104) );
  INV_X1 U36096 ( .I(n33174), .ZN(n25442) );
  INV_X1 U36097 ( .I(n34634), .ZN(n35039) );
  NAND2_X1 U36099 ( .A1(n3510), .A2(n45568), .ZN(n45569) );
  NAND2_X1 U36100 ( .A1(n17568), .A2(n45561), .ZN(n17567) );
  OAI21_X1 U36101 ( .A1(n47821), .A2(n3510), .B(n8603), .ZN(n17568) );
  NOR2_X1 U36102 ( .A1(n45225), .A2(n18911), .ZN(n18910) );
  NAND3_X1 U36106 ( .A1(n45630), .A2(n45633), .A3(n44921), .ZN(n44942) );
  NAND2_X1 U36107 ( .A1(n47297), .A2(n25477), .ZN(n44921) );
  NOR2_X1 U36108 ( .A1(n46059), .A2(n47324), .ZN(n20264) );
  NAND2_X1 U36109 ( .A1(n45452), .A2(n46745), .ZN(n45913) );
  NAND2_X1 U36111 ( .A1(n47853), .A2(n47851), .ZN(n23311) );
  INV_X1 U36112 ( .I(n48528), .ZN(n25955) );
  INV_X1 U36113 ( .I(n21894), .ZN(n48534) );
  NAND3_X1 U36115 ( .A1(n47417), .A2(n47416), .A3(n47415), .ZN(n47419) );
  NAND2_X1 U36116 ( .A1(n47687), .A2(n45267), .ZN(n47416) );
  INV_X1 U36117 ( .I(n47545), .ZN(n47174) );
  INV_X1 U36120 ( .I(n48139), .ZN(n22712) );
  OAI22_X1 U36124 ( .A1(n45153), .A2(n47581), .B1(n47593), .B2(n22549), .ZN(
        n19176) );
  NAND2_X1 U36126 ( .A1(n47378), .A2(n15825), .ZN(n45435) );
  INV_X1 U36127 ( .I(n47376), .ZN(n45439) );
  NOR2_X1 U36130 ( .A1(n46892), .A2(n17208), .ZN(n17207) );
  NAND2_X1 U36131 ( .A1(n63294), .A2(n10627), .ZN(n46929) );
  NOR2_X1 U36132 ( .A1(n23903), .A2(n47034), .ZN(n20297) );
  NAND2_X1 U36136 ( .A1(n33520), .A2(n34553), .ZN(n21474) );
  OAI22_X1 U36137 ( .A1(n64158), .A2(n560), .B1(n61262), .B2(n21317), .ZN(
        n35011) );
  NAND2_X1 U36140 ( .A1(n47211), .A2(n47079), .ZN(n24428) );
  INV_X1 U36141 ( .I(n48081), .ZN(n48562) );
  NAND2_X1 U36142 ( .A1(n48087), .A2(n48086), .ZN(n48088) );
  NAND3_X1 U36143 ( .A1(n47885), .A2(n47886), .A3(n59967), .ZN(n47887) );
  INV_X1 U36149 ( .I(n45231), .ZN(n49153) );
  NOR2_X1 U36150 ( .A1(n47019), .A2(n47018), .ZN(n19786) );
  NAND2_X1 U36151 ( .A1(n49458), .A2(n1205), .ZN(n49225) );
  INV_X1 U36152 ( .I(n19998), .ZN(n48992) );
  AOI22_X1 U36155 ( .A1(n44704), .A2(n16974), .B1(n44705), .B2(n23903), .ZN(
        n44708) );
  NAND2_X1 U36156 ( .A1(n17573), .A2(n47186), .ZN(n47188) );
  NAND2_X1 U36157 ( .A1(n18117), .A2(n48118), .ZN(n18116) );
  INV_X1 U36158 ( .I(n47185), .ZN(n18117) );
  AOI21_X1 U36159 ( .A1(n61025), .A2(n16933), .B(n18349), .ZN(n18106) );
  OAI22_X1 U36160 ( .A1(n47602), .A2(n7050), .B1(n47824), .B2(n47820), .ZN(
        n16933) );
  NOR2_X1 U36162 ( .A1(n48948), .A2(n26102), .ZN(n26098) );
  NAND3_X1 U36163 ( .A1(n50349), .A2(n60467), .A3(n50348), .ZN(n49866) );
  AOI21_X1 U36165 ( .A1(n49366), .A2(n49367), .B(n49365), .ZN(n24622) );
  NOR2_X1 U36166 ( .A1(n49550), .A2(n49551), .ZN(n18374) );
  OAI22_X1 U36167 ( .A1(n49558), .A2(n49557), .B1(n49556), .B2(n49555), .ZN(
        n49563) );
  NAND2_X1 U36168 ( .A1(n21127), .A2(n8347), .ZN(n49558) );
  INV_X1 U36169 ( .I(n20575), .ZN(n19378) );
  NOR2_X1 U36171 ( .A1(n23533), .A2(n50283), .ZN(n50117) );
  NAND2_X1 U36172 ( .A1(n17886), .A2(n18882), .ZN(n47149) );
  NAND2_X1 U36173 ( .A1(n49905), .A2(n25812), .ZN(n24304) );
  INV_X1 U36174 ( .I(n49441), .ZN(n17072) );
  NAND2_X1 U36175 ( .A1(n50091), .A2(n50090), .ZN(n22268) );
  NAND2_X1 U36178 ( .A1(n49348), .A2(n61362), .ZN(n49350) );
  NAND2_X1 U36180 ( .A1(n45302), .A2(n16296), .ZN(n45303) );
  NAND2_X1 U36181 ( .A1(n60510), .A2(n17379), .ZN(n17380) );
  INV_X1 U36183 ( .I(n50210), .ZN(n50207) );
  AOI21_X1 U36186 ( .A1(n49946), .A2(n61083), .B(n15550), .ZN(n48744) );
  INV_X1 U36187 ( .I(n49426), .ZN(n25869) );
  INV_X1 U36188 ( .I(n50048), .ZN(n16917) );
  NAND2_X1 U36190 ( .A1(n48675), .A2(n16256), .ZN(n48677) );
  NOR2_X1 U36192 ( .A1(n50142), .A2(n3055), .ZN(n49145) );
  NOR2_X1 U36193 ( .A1(n50348), .A2(n13684), .ZN(n24770) );
  NAND2_X1 U36194 ( .A1(n49110), .A2(n63605), .ZN(n22314) );
  INV_X1 U36195 ( .I(n48870), .ZN(n48871) );
  OAI21_X1 U36196 ( .A1(n50019), .A2(n50444), .B(n19653), .ZN(n50021) );
  NAND2_X1 U36197 ( .A1(n50019), .A2(n59621), .ZN(n19653) );
  NAND3_X1 U36198 ( .A1(n617), .A2(n49323), .A3(n18950), .ZN(n47063) );
  NAND2_X1 U36200 ( .A1(n49784), .A2(n49783), .ZN(n20011) );
  NAND2_X1 U36201 ( .A1(n49782), .A2(n25048), .ZN(n20010) );
  NAND2_X1 U36203 ( .A1(n48065), .A2(n48066), .ZN(n19896) );
  NAND2_X1 U36204 ( .A1(n49229), .A2(n19756), .ZN(n45233) );
  NOR2_X1 U36205 ( .A1(n48839), .A2(n48847), .ZN(n20741) );
  INV_X1 U36206 ( .I(n50543), .ZN(n19149) );
  INV_X1 U36207 ( .I(n65142), .ZN(n21600) );
  NAND3_X1 U36208 ( .A1(n18598), .A2(n49476), .A3(n25932), .ZN(n48270) );
  NAND2_X1 U36210 ( .A1(n23299), .A2(n19634), .ZN(n50447) );
  OAI22_X1 U36211 ( .A1(n20901), .A2(n49174), .B1(n23612), .B2(n49167), .ZN(
        n48837) );
  INV_X1 U36212 ( .I(n48836), .ZN(n18480) );
  AOI22_X1 U36213 ( .A1(n49026), .A2(n63084), .B1(n49028), .B2(n49027), .ZN(
        n25938) );
  OAI21_X1 U36214 ( .A1(n50400), .A2(n50076), .B(n19262), .ZN(n50087) );
  NAND2_X1 U36217 ( .A1(n48056), .A2(n48300), .ZN(n20417) );
  INV_X1 U36218 ( .I(n51684), .ZN(n18642) );
  OAI21_X1 U36223 ( .A1(n21835), .A2(n21834), .B(n49953), .ZN(n21833) );
  NAND2_X1 U36224 ( .A1(n35450), .A2(n36626), .ZN(n25784) );
  NAND3_X1 U36226 ( .A1(n17373), .A2(n54108), .A3(n13815), .ZN(n17372) );
  NAND2_X1 U36227 ( .A1(n23704), .A2(n53547), .ZN(n17373) );
  NAND2_X1 U36228 ( .A1(n10362), .A2(n55690), .ZN(n18293) );
  INV_X1 U36229 ( .I(n57008), .ZN(n23544) );
  NAND2_X1 U36232 ( .A1(n61282), .A2(n22499), .ZN(n52935) );
  OAI21_X1 U36234 ( .A1(n22039), .A2(n57010), .B(n56530), .ZN(n22510) );
  NOR3_X1 U36235 ( .A1(n55452), .A2(n3567), .A3(n55290), .ZN(n55291) );
  NAND3_X1 U36239 ( .A1(n1602), .A2(n52265), .A3(n52870), .ZN(n52267) );
  NAND2_X1 U36240 ( .A1(n61730), .A2(n1325), .ZN(n52266) );
  NOR2_X1 U36242 ( .A1(n53858), .A2(n53622), .ZN(n19412) );
  NAND2_X1 U36243 ( .A1(n187), .A2(n62769), .ZN(n18386) );
  INV_X1 U36244 ( .I(n55684), .ZN(n18108) );
  INV_X1 U36245 ( .I(n17753), .ZN(n17754) );
  NAND2_X1 U36247 ( .A1(n54688), .A2(n15040), .ZN(n25447) );
  NAND2_X1 U36248 ( .A1(n18219), .A2(n25437), .ZN(n17181) );
  OR2_X1 U36251 ( .A1(n24003), .A2(n20891), .Z(n52130) );
  NOR2_X1 U36252 ( .A1(n56638), .A2(n58846), .ZN(n22379) );
  INV_X1 U36254 ( .I(n56258), .ZN(n22294) );
  OAI22_X1 U36255 ( .A1(n25792), .A2(n54950), .B1(n54952), .B2(n54951), .ZN(
        n54953) );
  NAND2_X1 U36261 ( .A1(n54500), .A2(n21011), .ZN(n54064) );
  NAND2_X1 U36262 ( .A1(n55737), .A2(n55278), .ZN(n55285) );
  NAND2_X1 U36264 ( .A1(n19403), .A2(n59970), .ZN(n19402) );
  INV_X1 U36266 ( .I(n56172), .ZN(n19945) );
  OAI21_X1 U36268 ( .A1(n53280), .A2(n53303), .B(n53295), .ZN(n19577) );
  NOR2_X1 U36269 ( .A1(n16046), .A2(n56411), .ZN(n24312) );
  NOR2_X1 U36270 ( .A1(n54409), .A2(n1367), .ZN(n54417) );
  NOR2_X1 U36271 ( .A1(n22401), .A2(n5324), .ZN(n54425) );
  NAND2_X1 U36272 ( .A1(n52952), .A2(n55440), .ZN(n55309) );
  NOR2_X1 U36273 ( .A1(n56342), .A2(n1591), .ZN(n56293) );
  NAND2_X1 U36277 ( .A1(n54251), .A2(n14354), .ZN(n54267) );
  NAND3_X1 U36278 ( .A1(n55266), .A2(n55267), .A3(n55265), .ZN(n24524) );
  NAND2_X1 U36279 ( .A1(n53793), .A2(n53817), .ZN(n53776) );
  NAND3_X1 U36282 ( .A1(n55247), .A2(n55404), .A3(n55246), .ZN(n55253) );
  NAND2_X1 U36284 ( .A1(n53096), .A2(n53119), .ZN(n52895) );
  NAND2_X1 U36285 ( .A1(n55007), .A2(n55006), .ZN(n20541) );
  NAND2_X1 U36288 ( .A1(n52762), .A2(n25604), .ZN(n53335) );
  NAND2_X1 U36292 ( .A1(n62421), .A2(n9311), .ZN(n56481) );
  NOR2_X1 U36293 ( .A1(n57014), .A2(n24669), .ZN(n51352) );
  NAND2_X1 U36298 ( .A1(n56845), .A2(n56867), .ZN(n56851) );
  NAND2_X1 U36299 ( .A1(n55497), .A2(n55299), .ZN(n24980) );
  NOR2_X1 U36300 ( .A1(n53517), .A2(n53514), .ZN(n17101) );
  NAND2_X1 U36302 ( .A1(n5227), .A2(n54095), .ZN(n18861) );
  BUF_X4 U36303 ( .I(n54032), .Z(n54189) );
  NOR2_X1 U36305 ( .A1(n53793), .A2(n58811), .ZN(n53017) );
  INV_X1 U36306 ( .I(n19693), .ZN(n19692) );
  OAI21_X1 U36307 ( .A1(n21), .A2(n53797), .B(n53042), .ZN(n19694) );
  AOI21_X1 U36308 ( .A1(n53047), .A2(n53798), .B(n53046), .ZN(n17055) );
  NAND3_X1 U36309 ( .A1(n53043), .A2(n53800), .A3(n53045), .ZN(n17056) );
  INV_X1 U36310 ( .I(n53812), .ZN(n19154) );
  NAND2_X1 U36311 ( .A1(n53813), .A2(n53807), .ZN(n53810) );
  NOR2_X1 U36314 ( .A1(n61687), .A2(n25147), .ZN(n25146) );
  AND2_X1 U36315 ( .A1(n21828), .A2(n19203), .Z(n57133) );
  INV_X1 U36316 ( .I(n57108), .ZN(n19203) );
  NAND2_X1 U36317 ( .A1(n1591), .A2(n60353), .ZN(n18254) );
  NOR2_X1 U36318 ( .A1(n53107), .A2(n63767), .ZN(n53091) );
  NAND2_X1 U36319 ( .A1(n18376), .A2(n55895), .ZN(n18557) );
  NAND4_X1 U36320 ( .A1(n23856), .A2(n2820), .A3(n53147), .A4(n2037), .ZN(
        n53141) );
  NAND3_X1 U36321 ( .A1(n54755), .A2(n54764), .A3(n65124), .ZN(n54730) );
  NAND2_X1 U36325 ( .A1(n55790), .A2(n10248), .ZN(n22858) );
  INV_X1 U36327 ( .I(n55883), .ZN(n19076) );
  NAND2_X1 U36328 ( .A1(n10381), .A2(n55650), .ZN(n19023) );
  NAND2_X1 U36329 ( .A1(n55639), .A2(n59610), .ZN(n55645) );
  NAND2_X1 U36332 ( .A1(n55111), .A2(n55121), .ZN(n25682) );
  INV_X1 U36334 ( .I(n17287), .ZN(n16471) );
  AOI21_X1 U36335 ( .A1(n53737), .A2(n61933), .B(n53726), .ZN(n20635) );
  NAND2_X1 U36336 ( .A1(n50828), .A2(n53712), .ZN(n16592) );
  NAND4_X1 U36337 ( .A1(n54266), .A2(n54268), .A3(n54280), .A4(n54271), .ZN(
        n17433) );
  NOR2_X1 U36338 ( .A1(n51874), .A2(n51875), .ZN(n17437) );
  NOR2_X1 U36339 ( .A1(n54256), .A2(n64788), .ZN(n51875) );
  INV_X1 U36341 ( .I(n53889), .ZN(n18618) );
  INV_X1 U36342 ( .I(n53888), .ZN(n18619) );
  INV_X1 U36343 ( .I(n17861), .ZN(n18808) );
  NAND2_X1 U36344 ( .A1(n1590), .A2(n61228), .ZN(n18176) );
  NOR2_X1 U36345 ( .A1(n55598), .A2(n55597), .ZN(n24297) );
  NAND2_X1 U36346 ( .A1(n55595), .A2(n1592), .ZN(n55571) );
  NOR2_X1 U36347 ( .A1(n53480), .A2(n17111), .ZN(n17110) );
  NAND2_X1 U36348 ( .A1(n53492), .A2(n53514), .ZN(n17111) );
  NOR2_X1 U36349 ( .A1(n53490), .A2(n53493), .ZN(n17109) );
  NAND2_X1 U36350 ( .A1(n53525), .A2(n53526), .ZN(n17242) );
  INV_X1 U36353 ( .I(n56730), .ZN(n22024) );
  INV_X1 U36355 ( .I(n32164), .ZN(n23259) );
  NOR2_X1 U36356 ( .A1(n3082), .A2(n65189), .ZN(n17368) );
  NAND2_X1 U36358 ( .A1(n21751), .A2(n17538), .ZN(n34338) );
  NAND2_X1 U36361 ( .A1(n34196), .A2(n18390), .ZN(n17341) );
  INV_X1 U36362 ( .I(n33469), .ZN(n33760) );
  AND2_X1 U36363 ( .A1(n31976), .A2(n34752), .Z(n16087) );
  NOR2_X1 U36364 ( .A1(n31976), .A2(n20326), .ZN(n17614) );
  NAND3_X1 U36365 ( .A1(n18395), .A2(n35755), .A3(n35314), .ZN(n18394) );
  OAI21_X1 U36366 ( .A1(n59432), .A2(n34565), .B(n34564), .ZN(n34567) );
  NAND2_X1 U36367 ( .A1(n31299), .A2(n33442), .ZN(n22580) );
  AOI21_X1 U36371 ( .A1(n34118), .A2(n139), .B(n20524), .ZN(n34122) );
  INV_X1 U36372 ( .I(n34718), .ZN(n17163) );
  AND2_X1 U36373 ( .A1(n34669), .A2(n9687), .Z(n16155) );
  NOR2_X1 U36374 ( .A1(n9687), .A2(n242), .ZN(n21910) );
  NOR2_X1 U36375 ( .A1(n31356), .A2(n1429), .ZN(n24084) );
  NAND2_X1 U36377 ( .A1(n34604), .A2(n1798), .ZN(n24072) );
  NOR3_X1 U36378 ( .A1(n34952), .A2(n34564), .A3(n34947), .ZN(n32297) );
  NAND2_X1 U36379 ( .A1(n31767), .A2(n17199), .ZN(n19825) );
  NOR2_X1 U36381 ( .A1(n35229), .A2(n33807), .ZN(n35835) );
  INV_X1 U36383 ( .I(n34395), .ZN(n20356) );
  INV_X1 U36384 ( .I(n17614), .ZN(n34346) );
  NOR2_X1 U36387 ( .A1(n21388), .A2(n34307), .ZN(n34315) );
  INV_X1 U36392 ( .I(n25509), .ZN(n33003) );
  INV_X1 U36395 ( .I(n34172), .ZN(n34653) );
  NOR2_X1 U36397 ( .A1(n35670), .A2(n18382), .ZN(n18381) );
  NAND2_X1 U36399 ( .A1(n21252), .A2(n35224), .ZN(n16507) );
  INV_X1 U36400 ( .I(n17304), .ZN(n33212) );
  OAI21_X1 U36402 ( .A1(n35296), .A2(n35297), .B(n22278), .ZN(n20103) );
  NAND2_X1 U36403 ( .A1(n35680), .A2(n9679), .ZN(n23231) );
  NAND2_X1 U36405 ( .A1(n34525), .A2(n34668), .ZN(n23363) );
  OAI21_X1 U36406 ( .A1(n32934), .A2(n34247), .B(n34725), .ZN(n32424) );
  NOR3_X1 U36407 ( .A1(n34082), .A2(n18450), .A3(n34621), .ZN(n17697) );
  NOR2_X1 U36408 ( .A1(n34618), .A2(n33960), .ZN(n18450) );
  INV_X1 U36411 ( .I(n34423), .ZN(n26037) );
  AOI21_X1 U36412 ( .A1(n23281), .A2(n34358), .B(n34357), .ZN(n21460) );
  NAND2_X1 U36413 ( .A1(n34194), .A2(n17199), .ZN(n18679) );
  NOR4_X1 U36414 ( .A1(n16066), .A2(n61896), .A3(n10401), .A4(n20181), .ZN(
        n18682) );
  NAND2_X1 U36416 ( .A1(n61896), .A2(n34198), .ZN(n25731) );
  NAND2_X1 U36418 ( .A1(n35802), .A2(n35805), .ZN(n35795) );
  NAND2_X1 U36419 ( .A1(n35086), .A2(n37090), .ZN(n37310) );
  NOR2_X1 U36420 ( .A1(n23859), .A2(n35712), .ZN(n20259) );
  OAI21_X1 U36421 ( .A1(n23859), .A2(n33807), .B(n35712), .ZN(n33808) );
  OAI21_X1 U36422 ( .A1(n33801), .A2(n35247), .B(n35651), .ZN(n33800) );
  NOR2_X1 U36424 ( .A1(n33549), .A2(n35620), .ZN(n33315) );
  OAI21_X1 U36425 ( .A1(n33561), .A2(n33568), .B(n7273), .ZN(n33562) );
  INV_X1 U36426 ( .I(n21058), .ZN(n36495) );
  INV_X1 U36427 ( .I(n35003), .ZN(n33460) );
  NAND2_X1 U36429 ( .A1(n37361), .A2(n37359), .ZN(n22822) );
  NAND2_X1 U36430 ( .A1(n59011), .A2(n19573), .ZN(n34432) );
  NOR2_X1 U36432 ( .A1(n7092), .A2(n36847), .ZN(n36677) );
  NAND2_X1 U36433 ( .A1(n36676), .A2(n36847), .ZN(n36680) );
  INV_X1 U36434 ( .I(n34213), .ZN(n34214) );
  NAND2_X1 U36435 ( .A1(n35909), .A2(n35490), .ZN(n20915) );
  NOR2_X1 U36437 ( .A1(n24028), .A2(n19616), .ZN(n35558) );
  NAND2_X1 U36439 ( .A1(n33950), .A2(n19119), .ZN(n31354) );
  NOR2_X1 U36440 ( .A1(n60892), .A2(n15783), .ZN(n21311) );
  AOI21_X1 U36441 ( .A1(n18151), .A2(n35404), .B(n23146), .ZN(n36858) );
  AOI21_X1 U36442 ( .A1(n37044), .A2(n37055), .B(n37043), .ZN(n37045) );
  NOR2_X1 U36444 ( .A1(n36979), .A2(n61935), .ZN(n36990) );
  INV_X1 U36446 ( .I(n36980), .ZN(n37205) );
  NAND3_X1 U36447 ( .A1(n36212), .A2(n26243), .A3(n35348), .ZN(n34935) );
  NOR2_X1 U36448 ( .A1(n36211), .A2(n20867), .ZN(n21741) );
  NAND2_X1 U36453 ( .A1(n36857), .A2(n36856), .ZN(n18147) );
  NAND3_X1 U36455 ( .A1(n18149), .A2(n18151), .A3(n63697), .ZN(n18148) );
  NOR2_X1 U36456 ( .A1(n35404), .A2(n23146), .ZN(n18149) );
  NOR3_X1 U36460 ( .A1(n4834), .A2(n58561), .A3(n24661), .ZN(n37006) );
  NOR2_X1 U36461 ( .A1(n37007), .A2(n58561), .ZN(n24840) );
  NAND2_X1 U36462 ( .A1(n20951), .A2(n37161), .ZN(n37162) );
  INV_X1 U36463 ( .I(n17139), .ZN(n35809) );
  NOR3_X1 U36464 ( .A1(n35995), .A2(n21039), .A3(n62010), .ZN(n36000) );
  NOR2_X1 U36465 ( .A1(n1793), .A2(n37050), .ZN(n21039) );
  AOI21_X1 U36476 ( .A1(n10317), .A2(n35560), .B(n18885), .ZN(n26194) );
  NAND2_X1 U36477 ( .A1(n36484), .A2(n1525), .ZN(n18885) );
  NAND2_X1 U36478 ( .A1(n36472), .A2(n36471), .ZN(n36473) );
  NOR2_X1 U36479 ( .A1(n37110), .A2(n37111), .ZN(n22968) );
  NAND2_X1 U36480 ( .A1(n37106), .A2(n37359), .ZN(n37109) );
  NOR2_X1 U36481 ( .A1(n1524), .A2(n20124), .ZN(n17911) );
  OAI21_X1 U36483 ( .A1(n32442), .A2(n35163), .B(n32441), .ZN(n32451) );
  INV_X1 U36484 ( .I(n36420), .ZN(n18615) );
  NOR2_X1 U36485 ( .A1(n33784), .A2(n36420), .ZN(n18616) );
  NAND2_X1 U36488 ( .A1(n35146), .A2(n35965), .ZN(n16634) );
  NAND2_X1 U36489 ( .A1(n16114), .A2(n62026), .ZN(n35145) );
  NAND2_X1 U36491 ( .A1(n35905), .A2(n35911), .ZN(n25663) );
  OAI21_X1 U36492 ( .A1(n24118), .A2(n34878), .B(n35568), .ZN(n19813) );
  NOR3_X1 U36493 ( .A1(n35561), .A2(n35883), .A3(n10596), .ZN(n34871) );
  OAI22_X1 U36494 ( .A1(n34879), .A2(n7802), .B1(n34877), .B2(n34876), .ZN(
        n19814) );
  NAND2_X1 U36496 ( .A1(n34870), .A2(n15870), .ZN(n19632) );
  INV_X1 U36501 ( .I(n28469), .ZN(n17689) );
  NOR2_X1 U36502 ( .A1(n34477), .A2(n35352), .ZN(n25385) );
  NAND2_X1 U36503 ( .A1(n36416), .A2(n36408), .ZN(n19138) );
  INV_X1 U36504 ( .I(n39626), .ZN(n24204) );
  INV_X1 U36506 ( .I(n21348), .ZN(n38140) );
  NAND2_X1 U36507 ( .A1(n36403), .A2(n25592), .ZN(n25591) );
  OAI21_X1 U36508 ( .A1(n35456), .A2(n36061), .B(n58888), .ZN(n35457) );
  NOR2_X1 U36512 ( .A1(n37219), .A2(n37224), .ZN(n24824) );
  NAND2_X1 U36515 ( .A1(n36011), .A2(n4754), .ZN(n19554) );
  NAND2_X1 U36516 ( .A1(n17667), .A2(n36012), .ZN(n17666) );
  NAND2_X1 U36517 ( .A1(n36924), .A2(n36923), .ZN(n25386) );
  OAI21_X1 U36518 ( .A1(n34852), .A2(n36775), .B(n36776), .ZN(n22520) );
  NAND2_X1 U36521 ( .A1(n35896), .A2(n35897), .ZN(n19245) );
  INV_X1 U36522 ( .I(n51512), .ZN(n21578) );
  INV_X1 U36525 ( .I(n35065), .ZN(n36342) );
  NAND2_X1 U36527 ( .A1(n23648), .A2(n36343), .ZN(n24726) );
  NAND2_X1 U36528 ( .A1(n7933), .A2(n64087), .ZN(n33523) );
  NAND3_X1 U36529 ( .A1(n18130), .A2(n32692), .A3(n1525), .ZN(n32770) );
  OAI21_X1 U36530 ( .A1(n16733), .A2(n16732), .B(n39689), .ZN(n16731) );
  INV_X1 U36531 ( .I(n17924), .ZN(n16733) );
  INV_X1 U36532 ( .I(n17923), .ZN(n16732) );
  NAND3_X1 U36533 ( .A1(n23471), .A2(n23842), .A3(n18969), .ZN(n17038) );
  INV_X1 U36534 ( .I(n36565), .ZN(n36568) );
  INV_X1 U36535 ( .I(n34819), .ZN(n34463) );
  BUF_X2 U36536 ( .I(n24257), .Z(n17164) );
  INV_X1 U36541 ( .I(n27094), .ZN(n26569) );
  NAND2_X1 U36542 ( .A1(n27361), .A2(n19916), .ZN(n19915) );
  NAND2_X1 U36543 ( .A1(n27448), .A2(n20665), .ZN(n19916) );
  NOR2_X1 U36544 ( .A1(n28843), .A2(n6513), .ZN(n28150) );
  NOR2_X1 U36545 ( .A1(n28066), .A2(n21158), .ZN(n27044) );
  INV_X1 U36548 ( .I(n57113), .ZN(n25622) );
  INV_X1 U36549 ( .I(n38307), .ZN(n21767) );
  NAND3_X1 U36550 ( .A1(n36742), .A2(n23648), .A3(n17364), .ZN(n34092) );
  INV_X1 U36551 ( .I(n39357), .ZN(n19217) );
  INV_X1 U36552 ( .I(n1519), .ZN(n20523) );
  INV_X1 U36554 ( .I(n25479), .ZN(n21967) );
  INV_X1 U36555 ( .I(n38382), .ZN(n25374) );
  BUF_X2 U36557 ( .I(n38836), .Z(n17347) );
  INV_X1 U36558 ( .I(n39208), .ZN(n18868) );
  INV_X1 U36559 ( .I(n17164), .ZN(n26121) );
  NOR2_X1 U36561 ( .A1(n18333), .A2(n1745), .ZN(n39512) );
  NAND2_X1 U36562 ( .A1(n35120), .A2(n35119), .ZN(n16956) );
  NAND2_X1 U36563 ( .A1(n35118), .A2(n18313), .ZN(n16955) );
  NOR2_X1 U36564 ( .A1(n18617), .A2(n20130), .ZN(n16849) );
  INV_X1 U36565 ( .I(n37979), .ZN(n39639) );
  INV_X1 U36568 ( .I(n18305), .ZN(n18071) );
  NAND3_X1 U36569 ( .A1(n36895), .A2(n35384), .A3(n7103), .ZN(n23765) );
  INV_X1 U36570 ( .I(n39735), .ZN(n18056) );
  INV_X1 U36571 ( .I(n48954), .ZN(n16475) );
  NAND2_X1 U36573 ( .A1(n40258), .A2(n40464), .ZN(n37924) );
  NOR2_X1 U36574 ( .A1(n23932), .A2(n40199), .ZN(n38046) );
  NOR2_X1 U36575 ( .A1(n42448), .A2(n22759), .ZN(n41811) );
  NAND2_X1 U36576 ( .A1(n28414), .A2(n64614), .ZN(n28415) );
  NAND3_X1 U36578 ( .A1(n26935), .A2(n27471), .A3(n20509), .ZN(n20511) );
  NAND2_X1 U36579 ( .A1(n29303), .A2(n26968), .ZN(n26961) );
  NAND2_X1 U36581 ( .A1(n27406), .A2(n8436), .ZN(n22119) );
  INV_X1 U36582 ( .I(n28217), .ZN(n29121) );
  NOR2_X1 U36583 ( .A1(n1858), .A2(n58999), .ZN(n29027) );
  NAND2_X1 U36584 ( .A1(n29163), .A2(n28260), .ZN(n28261) );
  NOR2_X1 U36586 ( .A1(n24080), .A2(n21955), .ZN(n27268) );
  NAND2_X1 U36587 ( .A1(n28212), .A2(n8478), .ZN(n27405) );
  NAND2_X1 U36589 ( .A1(n18751), .A2(n64481), .ZN(n26622) );
  INV_X1 U36590 ( .I(n29379), .ZN(n29380) );
  NOR2_X1 U36591 ( .A1(n23383), .A2(n21132), .ZN(n26503) );
  INV_X1 U36592 ( .I(n28587), .ZN(n28148) );
  INV_X1 U36593 ( .I(n29286), .ZN(n28138) );
  NAND2_X1 U36594 ( .A1(n7772), .A2(n28510), .ZN(n26424) );
  NAND3_X1 U36595 ( .A1(n27025), .A2(n28054), .A3(n22408), .ZN(n25391) );
  INV_X1 U36596 ( .I(n27380), .ZN(n22094) );
  AOI21_X1 U36597 ( .A1(n26254), .A2(n22043), .B(n61049), .ZN(n21948) );
  NAND2_X1 U36599 ( .A1(n60993), .A2(n23876), .ZN(n21614) );
  INV_X1 U36600 ( .I(n25532), .ZN(n26958) );
  NAND2_X1 U36601 ( .A1(n29322), .A2(n19972), .ZN(n19995) );
  NOR2_X1 U36603 ( .A1(n27485), .A2(n27483), .ZN(n27471) );
  INV_X1 U36605 ( .I(n27657), .ZN(n28491) );
  NAND2_X1 U36606 ( .A1(n26903), .A2(n26074), .ZN(n28489) );
  AOI22_X1 U36608 ( .A1(n24967), .A2(n26411), .B1(n29176), .B2(n26410), .ZN(
        n21890) );
  INV_X1 U36609 ( .I(n28554), .ZN(n18471) );
  NOR2_X1 U36610 ( .A1(n27875), .A2(n1443), .ZN(n28529) );
  NOR2_X1 U36611 ( .A1(n24909), .A2(n28532), .ZN(n23724) );
  INV_X1 U36613 ( .I(n29712), .ZN(n27814) );
  NAND2_X1 U36615 ( .A1(n17741), .A2(n29713), .ZN(n17740) );
  NOR2_X1 U36616 ( .A1(n20743), .A2(n28620), .ZN(n17741) );
  NAND2_X1 U36617 ( .A1(n1895), .A2(n26606), .ZN(n27113) );
  NAND3_X1 U36618 ( .A1(n40578), .A2(n23145), .A3(n42259), .ZN(n40579) );
  INV_X1 U36619 ( .I(n40047), .ZN(n25651) );
  INV_X1 U36621 ( .I(n38838), .ZN(n17591) );
  NAND2_X1 U36622 ( .A1(n42287), .A2(n22776), .ZN(n17095) );
  NAND2_X1 U36623 ( .A1(n41386), .A2(n41382), .ZN(n39998) );
  NOR2_X1 U36624 ( .A1(n42449), .A2(n41306), .ZN(n38199) );
  AOI21_X1 U36625 ( .A1(n59583), .A2(n59409), .B(n20598), .ZN(n39792) );
  NOR2_X1 U36626 ( .A1(n42449), .A2(n42448), .ZN(n25596) );
  INV_X1 U36629 ( .I(n23481), .ZN(n37580) );
  INV_X1 U36630 ( .I(n38636), .ZN(n22287) );
  INV_X1 U36631 ( .I(n39769), .ZN(n17220) );
  INV_X1 U36638 ( .I(n38661), .ZN(n24407) );
  NAND2_X1 U36640 ( .A1(n25246), .A2(n13984), .ZN(n40322) );
  OAI22_X1 U36641 ( .A1(n40840), .A2(n41063), .B1(n40588), .B2(n62241), .ZN(
        n40590) );
  OAI21_X1 U36642 ( .A1(n23112), .A2(n41382), .B(n41122), .ZN(n39819) );
  NAND2_X1 U36643 ( .A1(n18664), .A2(n40763), .ZN(n18669) );
  NOR2_X1 U36644 ( .A1(n39998), .A2(n16461), .ZN(n41127) );
  NOR2_X1 U36645 ( .A1(n1737), .A2(n61994), .ZN(n39323) );
  NAND2_X1 U36646 ( .A1(n40293), .A2(n23516), .ZN(n23515) );
  INV_X1 U36647 ( .I(n40223), .ZN(n23516) );
  INV_X1 U36648 ( .I(n22916), .ZN(n16432) );
  INV_X1 U36650 ( .I(n41111), .ZN(n25943) );
  INV_X1 U36654 ( .I(n27544), .ZN(n20797) );
  NOR2_X1 U36655 ( .A1(n19755), .A2(n61251), .ZN(n19754) );
  AND2_X1 U36656 ( .A1(n29027), .A2(n60187), .Z(n16060) );
  NAND4_X1 U36658 ( .A1(n28204), .A2(n28206), .A3(n28205), .A4(n28207), .ZN(
        n28210) );
  NAND2_X1 U36659 ( .A1(n22857), .A2(n27526), .ZN(n22856) );
  NOR2_X1 U36663 ( .A1(n15779), .A2(n26482), .ZN(n26483) );
  NAND2_X1 U36664 ( .A1(n24080), .A2(n21956), .ZN(n21562) );
  INV_X1 U36665 ( .I(n17285), .ZN(n26772) );
  NAND2_X1 U36666 ( .A1(n61169), .A2(n58971), .ZN(n26770) );
  NOR2_X1 U36667 ( .A1(n27087), .A2(n21379), .ZN(n26518) );
  NAND2_X1 U36669 ( .A1(n27618), .A2(n26669), .ZN(n18915) );
  NOR2_X1 U36670 ( .A1(n27431), .A2(n22810), .ZN(n22958) );
  NAND2_X1 U36672 ( .A1(n27162), .A2(n27622), .ZN(n17996) );
  AOI21_X1 U36673 ( .A1(n27433), .A2(n27161), .B(n61992), .ZN(n22481) );
  NOR2_X1 U36674 ( .A1(n23940), .A2(n27611), .ZN(n27161) );
  NAND3_X1 U36675 ( .A1(n29887), .A2(n9654), .A3(n31241), .ZN(n29888) );
  NOR2_X1 U36677 ( .A1(n25786), .A2(n27469), .ZN(n27540) );
  INV_X1 U36678 ( .I(n27554), .ZN(n21000) );
  OAI21_X1 U36680 ( .A1(n27603), .A2(n16094), .B(n27604), .ZN(n23837) );
  AOI22_X1 U36681 ( .A1(n30352), .A2(n30351), .B1(n30343), .B2(n30344), .ZN(
        n20556) );
  INV_X1 U36682 ( .I(n16788), .ZN(n16793) );
  AOI21_X1 U36683 ( .A1(n27506), .A2(n29333), .B(n29340), .ZN(n27513) );
  NOR2_X1 U36685 ( .A1(n27249), .A2(n27868), .ZN(n25633) );
  OAI22_X1 U36686 ( .A1(n57792), .A2(n16136), .B1(n26801), .B2(n23528), .ZN(
        n26806) );
  NAND2_X1 U36687 ( .A1(n57792), .A2(n23529), .ZN(n23528) );
  NAND2_X1 U36688 ( .A1(n64337), .A2(n23303), .ZN(n23529) );
  NAND2_X1 U36689 ( .A1(n30585), .A2(n23918), .ZN(n24171) );
  NOR2_X1 U36691 ( .A1(n20539), .A2(n27109), .ZN(n26637) );
  NAND2_X1 U36692 ( .A1(n24734), .A2(n27526), .ZN(n19159) );
  NAND2_X1 U36693 ( .A1(n29930), .A2(n29929), .ZN(n30532) );
  OAI21_X1 U36695 ( .A1(n9618), .A2(n30523), .B(n29767), .ZN(n26839) );
  NAND2_X1 U36696 ( .A1(n57451), .A2(n40645), .ZN(n17213) );
  OAI22_X1 U36697 ( .A1(n1732), .A2(n40571), .B1(n39957), .B2(n16980), .ZN(
        n39830) );
  OAI22_X1 U36699 ( .A1(n40791), .A2(n64895), .B1(n61785), .B2(n61047), .ZN(
        n40564) );
  NAND4_X1 U36700 ( .A1(n42479), .A2(n61708), .A3(n25666), .A4(n5837), .ZN(
        n16669) );
  NOR2_X1 U36702 ( .A1(n40691), .A2(n23967), .ZN(n19574) );
  NOR2_X1 U36703 ( .A1(n42519), .A2(n64986), .ZN(n19962) );
  AOI22_X1 U36704 ( .A1(n16284), .A2(n21057), .B1(n22523), .B2(n23319), .ZN(
        n19604) );
  NAND2_X1 U36707 ( .A1(n25976), .A2(n41435), .ZN(n40698) );
  INV_X1 U36712 ( .I(n22045), .ZN(n41912) );
  NAND2_X1 U36713 ( .A1(n42444), .A2(n42443), .ZN(n24344) );
  INV_X1 U36714 ( .I(n42434), .ZN(n42435) );
  NAND4_X1 U36715 ( .A1(n42474), .A2(n42473), .A3(n18242), .A4(n25666), .ZN(
        n42476) );
  NAND4_X1 U36719 ( .A1(n41857), .A2(n3534), .A3(n41859), .A4(n41858), .ZN(
        n19276) );
  NAND2_X1 U36720 ( .A1(n60820), .A2(n40617), .ZN(n40618) );
  NOR2_X1 U36721 ( .A1(n57451), .A2(n40650), .ZN(n22005) );
  NAND3_X1 U36722 ( .A1(n38603), .A2(n38602), .A3(n40616), .ZN(n38610) );
  INV_X1 U36723 ( .I(n40526), .ZN(n40616) );
  OAI21_X1 U36724 ( .A1(n40974), .A2(n38607), .B(n40968), .ZN(n38608) );
  OAI22_X1 U36725 ( .A1(n59961), .A2(n41472), .B1(n19019), .B2(n64308), .ZN(
        n38762) );
  INV_X1 U36726 ( .I(n40754), .ZN(n19019) );
  NOR2_X1 U36728 ( .A1(n42403), .A2(n19793), .ZN(n42409) );
  NAND2_X1 U36729 ( .A1(n41276), .A2(n22608), .ZN(n22607) );
  NAND2_X1 U36730 ( .A1(n22609), .A2(n3534), .ZN(n22608) );
  NAND2_X1 U36732 ( .A1(n64277), .A2(n10587), .ZN(n39073) );
  NAND2_X1 U36733 ( .A1(n39067), .A2(n40650), .ZN(n24767) );
  INV_X1 U36735 ( .I(n17845), .ZN(n37610) );
  NAND2_X1 U36737 ( .A1(n38017), .A2(n19611), .ZN(n25072) );
  NOR3_X1 U36740 ( .A1(n39960), .A2(n18741), .A3(n40592), .ZN(n39962) );
  NOR2_X1 U36741 ( .A1(n984), .A2(n18741), .ZN(n39972) );
  INV_X1 U36742 ( .I(n18112), .ZN(n18937) );
  INV_X1 U36743 ( .I(n31268), .ZN(n31161) );
  NAND2_X1 U36744 ( .A1(n31268), .A2(n25989), .ZN(n18573) );
  OAI21_X1 U36745 ( .A1(n31163), .A2(n61251), .B(n20821), .ZN(n31170) );
  NAND2_X1 U36746 ( .A1(n31164), .A2(n61251), .ZN(n20821) );
  NAND2_X1 U36748 ( .A1(n28518), .A2(n26834), .ZN(n24440) );
  INV_X1 U36749 ( .I(n28899), .ZN(n28900) );
  NAND2_X1 U36750 ( .A1(n29877), .A2(n23315), .ZN(n21702) );
  INV_X1 U36751 ( .I(n29100), .ZN(n29092) );
  INV_X1 U36752 ( .I(n31110), .ZN(n31111) );
  INV_X1 U36754 ( .I(n31046), .ZN(n31047) );
  NAND2_X1 U36755 ( .A1(n21019), .A2(n12907), .ZN(n19597) );
  NAND2_X1 U36756 ( .A1(n19665), .A2(n30276), .ZN(n28775) );
  AOI21_X1 U36757 ( .A1(n25053), .A2(n25052), .B(n30004), .ZN(n28877) );
  NAND2_X1 U36759 ( .A1(n28039), .A2(n61643), .ZN(n27101) );
  NOR2_X1 U36760 ( .A1(n25052), .A2(n31224), .ZN(n30667) );
  NOR2_X1 U36761 ( .A1(n22322), .A2(n16279), .ZN(n31037) );
  NAND2_X1 U36764 ( .A1(n15727), .A2(n11425), .ZN(n29062) );
  NAND2_X1 U36765 ( .A1(n21262), .A2(n21261), .ZN(n30182) );
  NAND2_X1 U36766 ( .A1(n5631), .A2(n30181), .ZN(n21261) );
  NAND3_X1 U36767 ( .A1(n16116), .A2(n30243), .A3(n30242), .ZN(n30248) );
  INV_X1 U36768 ( .I(n30681), .ZN(n30243) );
  NAND2_X1 U36769 ( .A1(n30006), .A2(n23799), .ZN(n19525) );
  AOI21_X1 U36770 ( .A1(n30749), .A2(n57806), .B(n23799), .ZN(n19526) );
  INV_X1 U36771 ( .I(n30685), .ZN(n30683) );
  NAND2_X1 U36776 ( .A1(n30760), .A2(n7426), .ZN(n30308) );
  NAND2_X1 U36777 ( .A1(n30322), .A2(n23397), .ZN(n23396) );
  NOR2_X1 U36778 ( .A1(n28728), .A2(n12632), .ZN(n17293) );
  NAND2_X1 U36783 ( .A1(n31129), .A2(n60575), .ZN(n28953) );
  NOR3_X1 U36786 ( .A1(n61048), .A2(n29422), .A3(n21095), .ZN(n19207) );
  OAI21_X1 U36787 ( .A1(n19721), .A2(n19536), .B(n19534), .ZN(n30003) );
  NAND2_X1 U36788 ( .A1(n1432), .A2(n59096), .ZN(n19536) );
  OAI21_X1 U36789 ( .A1(n29594), .A2(n30616), .B(n62495), .ZN(n29596) );
  NOR2_X1 U36792 ( .A1(n21559), .A2(n9618), .ZN(n17605) );
  NAND2_X1 U36793 ( .A1(n26843), .A2(n27922), .ZN(n26844) );
  NOR2_X1 U36794 ( .A1(n22322), .A2(n1315), .ZN(n30150) );
  NOR2_X1 U36795 ( .A1(n25246), .A2(n20751), .ZN(n40324) );
  NAND2_X1 U36796 ( .A1(n25511), .A2(n16852), .ZN(n40101) );
  OAI21_X1 U36797 ( .A1(n4789), .A2(n43161), .B(n20602), .ZN(n43149) );
  NAND2_X1 U36799 ( .A1(n43375), .A2(n42630), .ZN(n25933) );
  NAND2_X1 U36800 ( .A1(n39036), .A2(n39037), .ZN(n23133) );
  NOR2_X1 U36801 ( .A1(n10415), .A2(n64363), .ZN(n42558) );
  NAND2_X1 U36802 ( .A1(n41755), .A2(n42971), .ZN(n40097) );
  OAI21_X1 U36803 ( .A1(n42968), .A2(n43460), .B(n65129), .ZN(n24027) );
  INV_X1 U36804 ( .I(n40897), .ZN(n25169) );
  NOR2_X1 U36806 ( .A1(n43336), .A2(n11229), .ZN(n22030) );
  INV_X1 U36807 ( .I(n43437), .ZN(n24087) );
  INV_X2 U36808 ( .I(n38345), .ZN(n41934) );
  OAI21_X1 U36809 ( .A1(n11229), .A2(n23561), .B(n1708), .ZN(n41630) );
  NAND2_X1 U36813 ( .A1(n42634), .A2(n11198), .ZN(n42757) );
  NAND3_X1 U36815 ( .A1(n42834), .A2(n41363), .A3(n65185), .ZN(n25712) );
  NAND3_X1 U36820 ( .A1(n42687), .A2(n42694), .A3(n42377), .ZN(n41524) );
  INV_X1 U36821 ( .I(n25929), .ZN(n41635) );
  NOR2_X1 U36826 ( .A1(n40956), .A2(n40613), .ZN(n19015) );
  NAND2_X1 U36827 ( .A1(n1500), .A2(n42354), .ZN(n42358) );
  INV_X1 U36828 ( .I(n43712), .ZN(n43312) );
  AOI22_X1 U36829 ( .A1(n43583), .A2(n1397), .B1(n41961), .B2(n2995), .ZN(
        n41962) );
  INV_X1 U36830 ( .I(n31073), .ZN(n31075) );
  NAND3_X1 U36831 ( .A1(n28114), .A2(n29457), .A3(n28113), .ZN(n28730) );
  NAND2_X1 U36836 ( .A1(n2310), .A2(n18785), .ZN(n23080) );
  NOR2_X1 U36837 ( .A1(n30250), .A2(n30252), .ZN(n18785) );
  AND3_X1 U36838 ( .A1(n25121), .A2(n25120), .A3(n31218), .Z(n16065) );
  NAND3_X1 U36839 ( .A1(n31273), .A2(n327), .A3(n31282), .ZN(n20365) );
  INV_X1 U36842 ( .I(n31079), .ZN(n29467) );
  AOI21_X1 U36843 ( .A1(n29887), .A2(n23008), .B(n9654), .ZN(n29393) );
  NAND2_X1 U36844 ( .A1(n30891), .A2(n31256), .ZN(n29394) );
  NAND2_X1 U36845 ( .A1(n31238), .A2(n9654), .ZN(n29402) );
  NAND2_X1 U36846 ( .A1(n30051), .A2(n61622), .ZN(n30052) );
  AOI22_X1 U36847 ( .A1(n30416), .A2(n30331), .B1(n62285), .B2(n30651), .ZN(
        n28715) );
  NOR2_X1 U36848 ( .A1(n19665), .A2(n30276), .ZN(n27518) );
  NAND2_X1 U36851 ( .A1(n60170), .A2(n21159), .ZN(n28289) );
  NOR3_X1 U36854 ( .A1(n29062), .A2(n29059), .A3(n18402), .ZN(n28294) );
  OAI21_X1 U36855 ( .A1(n27990), .A2(n17903), .B(n23901), .ZN(n27992) );
  NAND2_X1 U36858 ( .A1(n63237), .A2(n30724), .ZN(n30726) );
  NAND2_X1 U36860 ( .A1(n30718), .A2(n30719), .ZN(n19471) );
  NAND2_X1 U36861 ( .A1(n30683), .A2(n23349), .ZN(n22762) );
  INV_X1 U36863 ( .I(n29878), .ZN(n28990) );
  NAND2_X1 U36864 ( .A1(n29731), .A2(n20026), .ZN(n28992) );
  OAI21_X1 U36866 ( .A1(n1841), .A2(n1349), .B(n1842), .ZN(n29760) );
  INV_X1 U36867 ( .I(n23693), .ZN(n22070) );
  AOI21_X1 U36869 ( .A1(n29451), .A2(n60030), .B(n20808), .ZN(n29450) );
  OAI21_X1 U36870 ( .A1(n30772), .A2(n30771), .B(n30770), .ZN(n16830) );
  OAI21_X1 U36871 ( .A1(n21886), .A2(n20179), .B(n20178), .ZN(n30775) );
  AND2_X1 U36872 ( .A1(n30790), .A2(n30789), .Z(n16146) );
  AOI21_X1 U36873 ( .A1(n29730), .A2(n30018), .B(n29877), .ZN(n24651) );
  NAND2_X1 U36874 ( .A1(n31131), .A2(n29566), .ZN(n24158) );
  NAND2_X1 U36875 ( .A1(n1393), .A2(n42383), .ZN(n19292) );
  NAND2_X1 U36878 ( .A1(n41683), .A2(n62389), .ZN(n22469) );
  AOI21_X1 U36880 ( .A1(n43703), .A2(n43393), .B(n20243), .ZN(n19442) );
  NAND2_X1 U36881 ( .A1(n23488), .A2(n19844), .ZN(n19843) );
  INV_X1 U36883 ( .I(n42564), .ZN(n43164) );
  INV_X1 U36884 ( .I(n42972), .ZN(n17152) );
  NAND2_X1 U36885 ( .A1(n10111), .A2(n20844), .ZN(n21932) );
  NOR2_X1 U36887 ( .A1(n64363), .A2(n42917), .ZN(n41605) );
  AOI21_X1 U36888 ( .A1(n42607), .A2(n429), .B(n42593), .ZN(n41542) );
  NOR2_X1 U36890 ( .A1(n41562), .A2(n42849), .ZN(n41783) );
  INV_X1 U36892 ( .I(n23151), .ZN(n41591) );
  AOI21_X1 U36893 ( .A1(n17755), .A2(n11986), .B(n12864), .ZN(n19961) );
  NAND2_X1 U36895 ( .A1(n19241), .A2(n42404), .ZN(n19809) );
  NAND2_X1 U36897 ( .A1(n43506), .A2(n43502), .ZN(n40781) );
  INV_X1 U36899 ( .I(n42042), .ZN(n42038) );
  NAND2_X1 U36901 ( .A1(n21376), .A2(n65141), .ZN(n41334) );
  NAND3_X1 U36902 ( .A1(n43286), .A2(n10111), .A3(n24179), .ZN(n39429) );
  INV_X1 U36903 ( .I(n41705), .ZN(n22367) );
  NOR2_X1 U36905 ( .A1(n41906), .A2(n41904), .ZN(n25365) );
  NAND2_X1 U36907 ( .A1(n19742), .A2(n43948), .ZN(n42538) );
  NOR3_X1 U36908 ( .A1(n5261), .A2(n23184), .A3(n42324), .ZN(n42326) );
  NOR2_X1 U36911 ( .A1(n20526), .A2(n16144), .ZN(n42309) );
  OAI21_X1 U36912 ( .A1(n17245), .A2(n43625), .B(n43624), .ZN(n43639) );
  INV_X1 U36916 ( .I(n11362), .ZN(n16385) );
  NOR2_X1 U36917 ( .A1(n43108), .A2(n43107), .ZN(n43109) );
  NOR2_X1 U36918 ( .A1(n43114), .A2(n11362), .ZN(n16386) );
  NAND2_X1 U36920 ( .A1(n43184), .A2(n43513), .ZN(n20497) );
  NOR2_X1 U36923 ( .A1(n279), .A2(n43538), .ZN(n21518) );
  NAND2_X1 U36924 ( .A1(n41865), .A2(n20222), .ZN(n20221) );
  INV_X1 U36928 ( .I(n43303), .ZN(n17267) );
  AOI21_X1 U36929 ( .A1(n43301), .A2(n16890), .B(n43949), .ZN(n19098) );
  NAND3_X1 U36933 ( .A1(n42070), .A2(n1193), .A3(n1336), .ZN(n20038) );
  NAND2_X1 U36935 ( .A1(n42168), .A2(n19174), .ZN(n16553) );
  AOI21_X1 U36937 ( .A1(n42176), .A2(n64346), .B(n42876), .ZN(n16554) );
  OR2_X1 U36938 ( .A1(n43000), .A2(n16649), .Z(n16090) );
  INV_X2 U36939 ( .I(n58874), .ZN(n43089) );
  NAND2_X1 U36940 ( .A1(n23730), .A2(n60706), .ZN(n22677) );
  NAND2_X1 U36941 ( .A1(n1500), .A2(n22999), .ZN(n40278) );
  INV_X1 U36943 ( .I(n43515), .ZN(n42045) );
  OAI21_X1 U36944 ( .A1(n40882), .A2(n42423), .B(n22645), .ZN(n18299) );
  NAND3_X1 U36945 ( .A1(n43105), .A2(n10111), .A3(n43104), .ZN(n40883) );
  INV_X2 U36947 ( .I(n17300), .ZN(n44596) );
  INV_X1 U36948 ( .I(n42872), .ZN(n42873) );
  NAND2_X1 U36949 ( .A1(n43925), .A2(n20276), .ZN(n43927) );
  INV_X1 U36950 ( .I(n29414), .ZN(n18159) );
  OAI21_X1 U36953 ( .A1(n30093), .A2(n62585), .B(n19260), .ZN(n30101) );
  NAND2_X1 U36954 ( .A1(n30094), .A2(n62585), .ZN(n19260) );
  AOI22_X1 U36955 ( .A1(n17856), .A2(n30212), .B1(n23589), .B2(n61900), .ZN(
        n17855) );
  AOI22_X1 U36956 ( .A1(n30846), .A2(n17853), .B1(n30842), .B2(n30841), .ZN(
        n17852) );
  NOR2_X1 U36958 ( .A1(n30320), .A2(n30319), .ZN(n30325) );
  NAND2_X1 U36959 ( .A1(n31148), .A2(n59810), .ZN(n31149) );
  OAI22_X1 U36960 ( .A1(n18763), .A2(n18762), .B1(n18736), .B2(n740), .ZN(
        n18761) );
  INV_X1 U36961 ( .I(n31327), .ZN(n30990) );
  INV_X1 U36962 ( .I(n31850), .ZN(n25401) );
  INV_X1 U36963 ( .I(n30284), .ZN(n20009) );
  AOI22_X1 U36964 ( .A1(n29769), .A2(n29768), .B1(n29770), .B2(n16363), .ZN(
        n29777) );
  NAND2_X1 U36965 ( .A1(n29738), .A2(n62588), .ZN(n19179) );
  NOR2_X1 U36967 ( .A1(n30701), .A2(n30700), .ZN(n30714) );
  AOI21_X1 U36968 ( .A1(n29057), .A2(n29056), .B(n29055), .ZN(n29058) );
  NOR2_X1 U36969 ( .A1(n20343), .A2(n30524), .ZN(n20152) );
  NAND3_X1 U36970 ( .A1(n29533), .A2(n18917), .A3(n19451), .ZN(n29535) );
  NAND3_X1 U36974 ( .A1(n43252), .A2(n42665), .A3(n42660), .ZN(n40545) );
  NOR3_X1 U36976 ( .A1(n41670), .A2(n42788), .A3(n41665), .ZN(n43026) );
  NOR2_X1 U36977 ( .A1(n43024), .A2(n62620), .ZN(n43025) );
  INV_X1 U36978 ( .I(n45054), .ZN(n18727) );
  OAI21_X1 U36980 ( .A1(n42674), .A2(n6706), .B(n22225), .ZN(n41245) );
  NAND2_X1 U36981 ( .A1(n40685), .A2(n43150), .ZN(n22844) );
  AND2_X1 U36982 ( .A1(n42946), .A2(n42947), .Z(n16002) );
  INV_X1 U36983 ( .I(n44122), .ZN(n18311) );
  NAND2_X1 U36985 ( .A1(n42794), .A2(n43295), .ZN(n20847) );
  INV_X1 U36987 ( .I(n45844), .ZN(n44225) );
  NAND2_X1 U36988 ( .A1(n43701), .A2(n37917), .ZN(n43689) );
  OAI21_X1 U36991 ( .A1(n42691), .A2(n42697), .B(n42690), .ZN(n42709) );
  NAND2_X1 U36993 ( .A1(n64324), .A2(n43626), .ZN(n42096) );
  INV_X1 U36995 ( .I(n44143), .ZN(n46496) );
  OAI21_X1 U36998 ( .A1(n24071), .A2(n42958), .B(n42957), .ZN(n42959) );
  NAND2_X1 U36999 ( .A1(n43814), .A2(n19174), .ZN(n43815) );
  OAI21_X1 U37000 ( .A1(n29213), .A2(n18238), .B(n30679), .ZN(n18237) );
  INV_X1 U37001 ( .I(n31200), .ZN(n31403) );
  INV_X1 U37002 ( .I(n31518), .ZN(n31517) );
  OAI21_X1 U37003 ( .A1(n29513), .A2(n29512), .B(n21209), .ZN(n16684) );
  OAI21_X1 U37004 ( .A1(n29513), .A2(n29857), .B(n64940), .ZN(n16683) );
  INV_X1 U37006 ( .I(n51261), .ZN(n17403) );
  BUF_X2 U37007 ( .I(n23771), .Z(n19627) );
  NAND3_X1 U37008 ( .A1(n30122), .A2(n30519), .A3(n30525), .ZN(n30130) );
  INV_X1 U37009 ( .I(n61071), .ZN(n17735) );
  INV_X1 U37010 ( .I(n44360), .ZN(n20225) );
  INV_X1 U37013 ( .I(n46519), .ZN(n17228) );
  INV_X1 U37015 ( .I(n46592), .ZN(n21447) );
  OAI21_X1 U37017 ( .A1(n42779), .A2(n42778), .B(n61344), .ZN(n42789) );
  NAND2_X1 U37018 ( .A1(n24114), .A2(n10420), .ZN(n47833) );
  INV_X1 U37019 ( .I(n44754), .ZN(n19727) );
  INV_X1 U37020 ( .I(n42955), .ZN(n45843) );
  NAND2_X1 U37022 ( .A1(n48242), .A2(n48653), .ZN(n48243) );
  INV_X1 U37024 ( .I(n48645), .ZN(n18282) );
  INV_X1 U37027 ( .I(n46702), .ZN(n23073) );
  INV_X1 U37029 ( .I(n177), .ZN(n47577) );
  NAND2_X1 U37030 ( .A1(n47035), .A2(n20299), .ZN(n45530) );
  NAND2_X1 U37033 ( .A1(n47324), .A2(n6934), .ZN(n20830) );
  NAND2_X1 U37034 ( .A1(n6957), .A2(n209), .ZN(n19041) );
  INV_X1 U37036 ( .I(n46890), .ZN(n17208) );
  INV_X1 U37037 ( .I(n44181), .ZN(n46914) );
  NOR2_X1 U37041 ( .A1(n47316), .A2(n47315), .ZN(n47319) );
  INV_X1 U37043 ( .I(n32331), .ZN(n22471) );
  NOR2_X1 U37044 ( .A1(n47494), .A2(n12825), .ZN(n19568) );
  NAND2_X1 U37049 ( .A1(n25026), .A2(n47882), .ZN(n47631) );
  NAND2_X1 U37050 ( .A1(n637), .A2(n1266), .ZN(n43828) );
  NAND2_X1 U37052 ( .A1(n47818), .A2(n45972), .ZN(n23326) );
  NOR2_X1 U37053 ( .A1(n48594), .A2(n59056), .ZN(n47532) );
  AOI21_X1 U37054 ( .A1(n47691), .A2(n47682), .B(n47681), .ZN(n23077) );
  NAND2_X1 U37057 ( .A1(n47013), .A2(n24820), .ZN(n47526) );
  NAND3_X1 U37058 ( .A1(n687), .A2(n2357), .A3(n49698), .ZN(n45167) );
  NAND2_X1 U37061 ( .A1(n209), .A2(n48654), .ZN(n17280) );
  OAI21_X1 U37063 ( .A1(n48658), .A2(n47482), .B(n63311), .ZN(n47483) );
  NAND2_X1 U37065 ( .A1(n8692), .A2(n59695), .ZN(n47663) );
  NAND2_X1 U37069 ( .A1(n47707), .A2(n47706), .ZN(n19422) );
  NAND3_X1 U37071 ( .A1(n18787), .A2(n48209), .A3(n18570), .ZN(n47203) );
  NAND2_X1 U37073 ( .A1(n48118), .A2(n47137), .ZN(n25265) );
  NAND2_X1 U37074 ( .A1(n21894), .A2(n48239), .ZN(n17840) );
  OAI21_X1 U37075 ( .A1(n60753), .A2(n24558), .B(n59418), .ZN(n46077) );
  AOI21_X1 U37077 ( .A1(n48543), .A2(n48544), .B(n24364), .ZN(n24363) );
  INV_X1 U37078 ( .I(n47098), .ZN(n47097) );
  NOR2_X1 U37079 ( .A1(n34953), .A2(n34952), .ZN(n20846) );
  NOR2_X1 U37080 ( .A1(n22342), .A2(n63617), .ZN(n20845) );
  NAND2_X1 U37082 ( .A1(n47699), .A2(n1657), .ZN(n17610) );
  NOR2_X1 U37083 ( .A1(n45196), .A2(n45197), .ZN(n17611) );
  NOR2_X1 U37084 ( .A1(n13655), .A2(n47034), .ZN(n44706) );
  NOR2_X1 U37085 ( .A1(n47132), .A2(n48530), .ZN(n47187) );
  NAND2_X1 U37086 ( .A1(n25004), .A2(n47252), .ZN(n47256) );
  NAND2_X1 U37088 ( .A1(n42618), .A2(n47565), .ZN(n47564) );
  INV_X1 U37093 ( .I(n46771), .ZN(n48077) );
  NAND2_X1 U37097 ( .A1(n6313), .A2(n49739), .ZN(n48396) );
  NAND3_X1 U37098 ( .A1(n46082), .A2(n12845), .A3(n48953), .ZN(n46084) );
  INV_X1 U37100 ( .I(n46730), .ZN(n46735) );
  AOI21_X1 U37101 ( .A1(n47431), .A2(n47736), .B(n21786), .ZN(n21785) );
  NAND2_X1 U37102 ( .A1(n64096), .A2(n59008), .ZN(n21787) );
  INV_X1 U37103 ( .I(n46745), .ZN(n21788) );
  NOR2_X1 U37105 ( .A1(n22549), .A2(n47580), .ZN(n22009) );
  INV_X1 U37106 ( .I(n50306), .ZN(n50301) );
  AOI21_X1 U37107 ( .A1(n18821), .A2(n49377), .B(n23576), .ZN(n23575) );
  INV_X1 U37110 ( .I(n49216), .ZN(n44005) );
  OAI21_X1 U37111 ( .A1(n23661), .A2(n47197), .B(n48212), .ZN(n18756) );
  INV_X1 U37112 ( .I(n46591), .ZN(n19013) );
  INV_X1 U37113 ( .I(n47870), .ZN(n21951) );
  NOR2_X1 U37114 ( .A1(n59698), .A2(n47654), .ZN(n47657) );
  OAI22_X1 U37115 ( .A1(n47660), .A2(n47659), .B1(n23361), .B2(n47831), .ZN(
        n47661) );
  AOI21_X1 U37116 ( .A1(n48379), .A2(n48979), .B(n16379), .ZN(n20662) );
  NAND2_X1 U37119 ( .A1(n49851), .A2(n16379), .ZN(n17422) );
  OAI21_X1 U37121 ( .A1(n63294), .A2(n45623), .B(n47310), .ZN(n45624) );
  NAND2_X1 U37122 ( .A1(n48679), .A2(n9863), .ZN(n24916) );
  NAND3_X1 U37123 ( .A1(n49702), .A2(n49757), .A3(n48678), .ZN(n20730) );
  NOR2_X1 U37124 ( .A1(n47418), .A2(n23995), .ZN(n23994) );
  OAI21_X1 U37125 ( .A1(n46755), .A2(n45267), .B(n47690), .ZN(n20566) );
  AOI21_X1 U37126 ( .A1(n49556), .A2(n19867), .B(n24394), .ZN(n48274) );
  NAND2_X1 U37127 ( .A1(n18609), .A2(n1471), .ZN(n49884) );
  NOR2_X1 U37129 ( .A1(n48577), .A2(n64267), .ZN(n45892) );
  NAND2_X1 U37130 ( .A1(n49512), .A2(n1261), .ZN(n49513) );
  OAI22_X1 U37131 ( .A1(n21189), .A2(n21188), .B1(n1377), .B2(n46777), .ZN(
        n21190) );
  AOI22_X1 U37134 ( .A1(n49797), .A2(n1642), .B1(n47343), .B2(n49114), .ZN(
        n19849) );
  OAI21_X1 U37135 ( .A1(n49797), .A2(n1642), .B(n62724), .ZN(n47344) );
  INV_X1 U37138 ( .I(n16589), .ZN(n16588) );
  OAI21_X1 U37139 ( .A1(n16591), .A2(n46963), .B(n46947), .ZN(n16589) );
  NOR2_X1 U37140 ( .A1(n48421), .A2(n22570), .ZN(n16586) );
  INV_X1 U37141 ( .I(n47058), .ZN(n20594) );
  NAND2_X1 U37142 ( .A1(n49986), .A2(n60209), .ZN(n16333) );
  NOR2_X1 U37147 ( .A1(n59293), .A2(n34974), .ZN(n34976) );
  NOR2_X1 U37148 ( .A1(n44669), .A2(n19751), .ZN(n19750) );
  OAI21_X1 U37150 ( .A1(n49908), .A2(n14314), .B(n63357), .ZN(n19747) );
  NAND2_X1 U37151 ( .A1(n49792), .A2(n47347), .ZN(n48436) );
  OAI21_X1 U37153 ( .A1(n45920), .A2(n45921), .B(n61083), .ZN(n45922) );
  NOR2_X1 U37154 ( .A1(n48024), .A2(n21835), .ZN(n45927) );
  NOR2_X1 U37155 ( .A1(n7866), .A2(n49810), .ZN(n47760) );
  OAI21_X1 U37156 ( .A1(n47818), .A2(n45969), .B(n45568), .ZN(n25779) );
  NOR2_X1 U37157 ( .A1(n47605), .A2(n47827), .ZN(n47608) );
  NOR3_X1 U37161 ( .A1(n24692), .A2(n19379), .A3(n49918), .ZN(n19510) );
  INV_X1 U37163 ( .I(n63009), .ZN(n51138) );
  AOI21_X1 U37164 ( .A1(n63663), .A2(n48811), .B(n48431), .ZN(n17091) );
  NOR2_X1 U37165 ( .A1(n48923), .A2(n48924), .ZN(n48928) );
  NOR3_X1 U37166 ( .A1(n48925), .A2(n57194), .A3(n49278), .ZN(n48926) );
  NOR2_X1 U37167 ( .A1(n48984), .A2(n21526), .ZN(n21525) );
  OAI21_X1 U37169 ( .A1(n17126), .A2(n49843), .B(n48970), .ZN(n48057) );
  INV_X1 U37170 ( .I(n24583), .ZN(n47931) );
  AOI21_X1 U37175 ( .A1(n48363), .A2(n16986), .B(n16411), .ZN(n48364) );
  NAND3_X1 U37176 ( .A1(n59493), .A2(n49789), .A3(n46004), .ZN(n49791) );
  NOR2_X1 U37177 ( .A1(n49287), .A2(n49276), .ZN(n48931) );
  NOR2_X1 U37182 ( .A1(n17874), .A2(n49317), .ZN(n19998) );
  NAND2_X1 U37183 ( .A1(n49355), .A2(n50042), .ZN(n22235) );
  NAND2_X1 U37185 ( .A1(n17514), .A2(n49842), .ZN(n17513) );
  NAND3_X1 U37188 ( .A1(n48704), .A2(n8129), .A3(n49607), .ZN(n17948) );
  NAND2_X1 U37189 ( .A1(n49494), .A2(n6704), .ZN(n20671) );
  NAND2_X1 U37190 ( .A1(n7866), .A2(n18882), .ZN(n19219) );
  NAND2_X1 U37191 ( .A1(n17885), .A2(n22264), .ZN(n50231) );
  NOR2_X1 U37192 ( .A1(n23299), .A2(n18882), .ZN(n50234) );
  AOI21_X1 U37193 ( .A1(n50296), .A2(n3054), .B(n1643), .ZN(n50055) );
  INV_X1 U37194 ( .I(n49473), .ZN(n25932) );
  INV_X1 U37195 ( .I(n49201), .ZN(n49131) );
  NOR2_X1 U37196 ( .A1(n9229), .A2(n50360), .ZN(n17200) );
  NAND2_X1 U37198 ( .A1(n25813), .A2(n25810), .ZN(n49907) );
  NOR2_X1 U37199 ( .A1(n50348), .A2(n21052), .ZN(n50258) );
  OAI21_X1 U37203 ( .A1(n25812), .A2(n48341), .B(n63357), .ZN(n47074) );
  OAI21_X1 U37205 ( .A1(n23992), .A2(n50420), .B(n2878), .ZN(n20562) );
  NOR2_X1 U37206 ( .A1(n50418), .A2(n50419), .ZN(n50434) );
  NAND2_X1 U37207 ( .A1(n50215), .A2(n50221), .ZN(n49102) );
  NOR2_X1 U37208 ( .A1(n49101), .A2(n1383), .ZN(n18079) );
  INV_X1 U37210 ( .I(n19530), .ZN(n51327) );
  NAND2_X1 U37211 ( .A1(n64135), .A2(n6411), .ZN(n49712) );
  NAND2_X1 U37212 ( .A1(n47987), .A2(n47988), .ZN(n22085) );
  NAND2_X1 U37213 ( .A1(n23500), .A2(n17334), .ZN(n24235) );
  NOR2_X1 U37214 ( .A1(n9594), .A2(n17335), .ZN(n49299) );
  NOR2_X1 U37216 ( .A1(n62724), .A2(n48441), .ZN(n25528) );
  NAND2_X1 U37221 ( .A1(n15693), .A2(n4815), .ZN(n49216) );
  NAND2_X1 U37222 ( .A1(n26099), .A2(n49781), .ZN(n26101) );
  NAND2_X1 U37223 ( .A1(n48705), .A2(n49612), .ZN(n25041) );
  NAND2_X1 U37224 ( .A1(n25967), .A2(n49055), .ZN(n48684) );
  NOR2_X1 U37225 ( .A1(n50305), .A2(n50304), .ZN(n48579) );
  NAND2_X1 U37227 ( .A1(n44790), .A2(n1633), .ZN(n18181) );
  NOR3_X1 U37229 ( .A1(n49554), .A2(n49553), .A3(n49570), .ZN(n18373) );
  INV_X1 U37231 ( .I(n47358), .ZN(n24928) );
  INV_X1 U37232 ( .I(n30402), .ZN(n52350) );
  NAND2_X1 U37233 ( .A1(n49649), .A2(n1643), .ZN(n21373) );
  NOR2_X1 U37234 ( .A1(n4734), .A2(n1643), .ZN(n21372) );
  AOI21_X1 U37236 ( .A1(n24691), .A2(n15826), .B(n1641), .ZN(n24690) );
  AOI21_X1 U37237 ( .A1(n49618), .A2(n50373), .B(n49617), .ZN(n49622) );
  NAND2_X1 U37238 ( .A1(n1374), .A2(n48851), .ZN(n24804) );
  INV_X1 U37239 ( .I(n51604), .ZN(n23218) );
  BUF_X2 U37240 ( .I(n52444), .Z(n20332) );
  INV_X1 U37241 ( .I(n61518), .ZN(n24203) );
  INV_X1 U37244 ( .I(n49434), .ZN(n24880) );
  INV_X1 U37245 ( .I(n50916), .ZN(n21668) );
  INV_X1 U37246 ( .I(n17446), .ZN(n50440) );
  NAND2_X1 U37248 ( .A1(n48741), .A2(n49950), .ZN(n22424) );
  NAND3_X1 U37249 ( .A1(n49834), .A2(n49833), .A3(n49832), .ZN(n49840) );
  INV_X1 U37250 ( .I(n51199), .ZN(n51200) );
  INV_X1 U37251 ( .I(n50952), .ZN(n18222) );
  NAND3_X1 U37252 ( .A1(n49937), .A2(n23414), .A3(n60467), .ZN(n24768) );
  INV_X1 U37254 ( .I(n50929), .ZN(n21480) );
  BUF_X2 U37255 ( .I(n51140), .Z(n25415) );
  INV_X2 U37256 ( .I(n25099), .ZN(n51548) );
  OAI22_X1 U37257 ( .A1(n50232), .A2(n60360), .B1(n25966), .B2(n50447), .ZN(
        n50020) );
  AOI22_X1 U37262 ( .A1(n49173), .A2(n49174), .B1(n49566), .B2(n49175), .ZN(
        n22539) );
  INV_X1 U37263 ( .I(n51748), .ZN(n24713) );
  INV_X1 U37264 ( .I(n51274), .ZN(n51540) );
  NOR2_X1 U37265 ( .A1(n56547), .A2(n56544), .ZN(n56534) );
  INV_X1 U37266 ( .I(n50166), .ZN(n20303) );
  OAI21_X1 U37267 ( .A1(n54027), .A2(n54026), .B(n23482), .ZN(n21930) );
  INV_X1 U37269 ( .I(n51539), .ZN(n21107) );
  NAND2_X1 U37270 ( .A1(n57042), .A2(n52825), .ZN(n52821) );
  BUF_X2 U37271 ( .I(n52373), .Z(n23878) );
  NOR2_X1 U37273 ( .A1(n21296), .A2(n4473), .ZN(n52988) );
  NAND2_X1 U37274 ( .A1(n54436), .A2(n52958), .ZN(n54618) );
  AOI21_X1 U37277 ( .A1(n53624), .A2(n18521), .B(n18520), .ZN(n18519) );
  INV_X1 U37279 ( .I(n4226), .ZN(n18522) );
  NAND2_X1 U37280 ( .A1(n53616), .A2(n61560), .ZN(n18523) );
  NAND2_X1 U37281 ( .A1(n18247), .A2(n55017), .ZN(n55018) );
  NAND2_X1 U37282 ( .A1(n55264), .A2(n16848), .ZN(n16847) );
  NAND2_X1 U37283 ( .A1(n54034), .A2(n54058), .ZN(n53914) );
  NAND2_X1 U37284 ( .A1(n53616), .A2(n62664), .ZN(n18499) );
  INV_X1 U37285 ( .I(n59970), .ZN(n19401) );
  NOR2_X1 U37290 ( .A1(n61736), .A2(n61502), .ZN(n54619) );
  NAND2_X1 U37292 ( .A1(n23095), .A2(n52706), .ZN(n52699) );
  OAI21_X1 U37293 ( .A1(n53196), .A2(n50676), .B(n23891), .ZN(n25461) );
  NAND2_X1 U37298 ( .A1(n54860), .A2(n24009), .ZN(n54848) );
  NAND3_X1 U37301 ( .A1(n52767), .A2(n52768), .A3(n16708), .ZN(n52770) );
  NAND2_X1 U37303 ( .A1(n55501), .A2(n55500), .ZN(n20926) );
  NAND2_X1 U37304 ( .A1(n55684), .A2(n18109), .ZN(n55495) );
  NAND2_X1 U37305 ( .A1(n65283), .A2(n55695), .ZN(n20958) );
  NOR2_X1 U37306 ( .A1(n55690), .A2(n52044), .ZN(n51964) );
  INV_X1 U37309 ( .I(n50782), .ZN(n22310) );
  INV_X1 U37314 ( .I(n50616), .ZN(n17234) );
  INV_X1 U37315 ( .I(n24923), .ZN(n19403) );
  NOR2_X1 U37316 ( .A1(n57018), .A2(n25160), .ZN(n21575) );
  NAND2_X1 U37317 ( .A1(n52706), .A2(n14943), .ZN(n52247) );
  NAND2_X1 U37318 ( .A1(n18270), .A2(n11121), .ZN(n18269) );
  NAND2_X1 U37319 ( .A1(n53176), .A2(n53541), .ZN(n19562) );
  INV_X1 U37320 ( .I(n20630), .ZN(n53182) );
  NOR2_X1 U37321 ( .A1(n61554), .A2(n56404), .ZN(n22388) );
  NAND2_X1 U37322 ( .A1(n54039), .A2(n53907), .ZN(n26198) );
  INV_X1 U37323 ( .I(n16708), .ZN(n53005) );
  OAI21_X1 U37324 ( .A1(n51961), .A2(n18109), .B(n20849), .ZN(n52918) );
  NAND2_X1 U37326 ( .A1(n56588), .A2(n56587), .ZN(n20129) );
  NAND2_X1 U37327 ( .A1(n56582), .A2(n56581), .ZN(n56583) );
  NAND2_X1 U37328 ( .A1(n16767), .A2(n21728), .ZN(n52234) );
  AOI21_X1 U37329 ( .A1(n10425), .A2(n59831), .B(n53545), .ZN(n53546) );
  OAI22_X1 U37330 ( .A1(n53016), .A2(n53015), .B1(n64076), .B2(n13940), .ZN(
        n25268) );
  INV_X1 U37334 ( .I(n54346), .ZN(n24636) );
  AOI21_X1 U37335 ( .A1(n49087), .A2(n54023), .B(n49086), .ZN(n21997) );
  INV_X1 U37336 ( .I(n52497), .ZN(n52498) );
  NOR2_X1 U37337 ( .A1(n65175), .A2(n56404), .ZN(n19356) );
  AOI21_X1 U37338 ( .A1(n55005), .A2(n18145), .B(n55310), .ZN(n55007) );
  AOI21_X1 U37340 ( .A1(n55435), .A2(n55436), .B(n18257), .ZN(n18256) );
  NOR2_X1 U37341 ( .A1(n55437), .A2(n55440), .ZN(n18258) );
  NAND2_X1 U37342 ( .A1(n55442), .A2(n55443), .ZN(n19818) );
  OAI21_X1 U37345 ( .A1(n17935), .A2(n54459), .B(n18247), .ZN(n54455) );
  AOI22_X1 U37346 ( .A1(n54590), .A2(n54589), .B1(n54588), .B2(n818), .ZN(
        n54591) );
  NOR2_X1 U37348 ( .A1(n55681), .A2(n55451), .ZN(n24466) );
  NOR2_X1 U37349 ( .A1(n64978), .A2(n60794), .ZN(n19197) );
  NOR2_X1 U37351 ( .A1(n55425), .A2(n55721), .ZN(n52121) );
  NAND2_X1 U37353 ( .A1(n21081), .A2(n55986), .ZN(n55990) );
  NAND2_X1 U37354 ( .A1(n55938), .A2(n18194), .ZN(n55939) );
  NOR2_X1 U37355 ( .A1(n57047), .A2(n57050), .ZN(n19614) );
  NAND2_X1 U37356 ( .A1(n53242), .A2(n21453), .ZN(n20362) );
  NAND2_X1 U37359 ( .A1(n20163), .A2(n53860), .ZN(n53429) );
  NAND2_X1 U37360 ( .A1(n65282), .A2(n22201), .ZN(n20163) );
  OAI22_X1 U37361 ( .A1(n21732), .A2(n56541), .B1(n56545), .B2(n56542), .ZN(
        n56543) );
  NAND2_X1 U37367 ( .A1(n518), .A2(n53284), .ZN(n53285) );
  NAND2_X1 U37368 ( .A1(n56328), .A2(n56342), .ZN(n24585) );
  INV_X1 U37369 ( .I(n53200), .ZN(n20691) );
  INV_X1 U37371 ( .I(n51884), .ZN(n51886) );
  NAND2_X1 U37374 ( .A1(n15820), .A2(n52125), .ZN(n16585) );
  AOI21_X1 U37375 ( .A1(n16584), .A2(n52122), .B(n52121), .ZN(n16583) );
  NOR2_X1 U37376 ( .A1(n55908), .A2(n52126), .ZN(n16584) );
  NAND2_X1 U37377 ( .A1(n21287), .A2(n54268), .ZN(n19884) );
  NOR2_X1 U37379 ( .A1(n17799), .A2(n62711), .ZN(n55232) );
  NAND2_X1 U37380 ( .A1(n17799), .A2(n18786), .ZN(n55177) );
  NOR2_X1 U37382 ( .A1(n56839), .A2(n56838), .ZN(n17651) );
  NOR2_X1 U37385 ( .A1(n55136), .A2(n8027), .ZN(n20881) );
  NOR3_X1 U37386 ( .A1(n55131), .A2(n11353), .A3(n55166), .ZN(n52649) );
  NOR2_X1 U37387 ( .A1(n55639), .A2(n52309), .ZN(n52310) );
  NAND4_X1 U37389 ( .A1(n19943), .A2(n19942), .A3(n56173), .A4(n19941), .ZN(
        n56178) );
  OAI21_X1 U37390 ( .A1(n19945), .A2(n19944), .B(n19853), .ZN(n19943) );
  AOI21_X1 U37391 ( .A1(n56496), .A2(n16217), .B(n25705), .ZN(n25704) );
  NOR2_X1 U37392 ( .A1(n56497), .A2(n19827), .ZN(n25705) );
  NAND2_X1 U37393 ( .A1(n54417), .A2(n15202), .ZN(n54418) );
  INV_X1 U37394 ( .I(n54425), .ZN(n54423) );
  NAND2_X1 U37395 ( .A1(n54565), .A2(n22572), .ZN(n25763) );
  NOR2_X1 U37398 ( .A1(n53085), .A2(n53084), .ZN(n20659) );
  NAND2_X1 U37399 ( .A1(n53129), .A2(n5614), .ZN(n52227) );
  INV_X1 U37400 ( .I(n55338), .ZN(n18288) );
  NOR2_X1 U37401 ( .A1(n55626), .A2(n52309), .ZN(n26183) );
  AOI21_X1 U37402 ( .A1(n56133), .A2(n17408), .B(n56191), .ZN(n56136) );
  NAND2_X1 U37404 ( .A1(n60203), .A2(n55882), .ZN(n55847) );
  OAI21_X1 U37405 ( .A1(n56351), .A2(n22891), .B(n56343), .ZN(n56346) );
  NAND2_X1 U37407 ( .A1(n60092), .A2(n63830), .ZN(n19032) );
  INV_X1 U37408 ( .I(n19037), .ZN(n19036) );
  NAND2_X1 U37409 ( .A1(n16168), .A2(n138), .ZN(n19708) );
  NOR2_X1 U37411 ( .A1(n21210), .A2(n15703), .ZN(n17270) );
  NAND2_X1 U37412 ( .A1(n55886), .A2(n55879), .ZN(n19073) );
  INV_X1 U37413 ( .I(n55880), .ZN(n19075) );
  INV_X1 U37414 ( .I(n25344), .ZN(n53985) );
  OR3_X1 U37416 ( .A1(n53741), .A2(n53715), .A3(n50470), .Z(n50471) );
  NAND2_X1 U37417 ( .A1(n54710), .A2(n23448), .ZN(n22491) );
  NAND3_X1 U37418 ( .A1(n54723), .A2(n54741), .A3(n54709), .ZN(n54710) );
  OAI21_X1 U37419 ( .A1(n52895), .A2(n53109), .B(n53048), .ZN(n23594) );
  NAND2_X1 U37422 ( .A1(n53332), .A2(n53331), .ZN(n53333) );
  NAND2_X1 U37423 ( .A1(n61872), .A2(n56963), .ZN(n21477) );
  NOR2_X1 U37425 ( .A1(n1583), .A2(n64845), .ZN(n56909) );
  INV_X1 U37426 ( .I(n55835), .ZN(n20416) );
  OAI21_X1 U37427 ( .A1(n15800), .A2(n55881), .B(n52042), .ZN(n17844) );
  INV_X1 U37428 ( .I(n53995), .ZN(n53979) );
  OAI21_X1 U37429 ( .A1(n21438), .A2(n21437), .B(n57134), .ZN(n21436) );
  NOR2_X1 U37430 ( .A1(n15877), .A2(n4030), .ZN(n21438) );
  NOR2_X1 U37431 ( .A1(n54569), .A2(n54530), .ZN(n19376) );
  NAND4_X1 U37433 ( .A1(n56480), .A2(n56483), .A3(n56482), .A4(n56481), .ZN(
        n56488) );
  NAND2_X1 U37437 ( .A1(n20438), .A2(n56775), .ZN(n56774) );
  AOI21_X1 U37439 ( .A1(n55570), .A2(n55569), .B(n15933), .ZN(n55572) );
  INV_X1 U37440 ( .I(n55867), .ZN(n55887) );
  NAND3_X1 U37443 ( .A1(n56851), .A2(n64833), .A3(n56850), .ZN(n56852) );
  INV_X1 U37444 ( .I(n19797), .ZN(n55332) );
  NAND2_X1 U37445 ( .A1(n54256), .A2(n64788), .ZN(n54261) );
  NOR2_X1 U37446 ( .A1(n20438), .A2(n56808), .ZN(n56797) );
  NAND2_X1 U37447 ( .A1(n20631), .A2(n53702), .ZN(n53703) );
  INV_X1 U37449 ( .I(n53819), .ZN(n21750) );
  AOI22_X1 U37450 ( .A1(n56147), .A2(n56173), .B1(n56148), .B2(n1590), .ZN(
        n24809) );
  OAI21_X1 U37451 ( .A1(n22221), .A2(n22222), .B(n53101), .ZN(n19254) );
  INV_X1 U37454 ( .I(n55106), .ZN(n55107) );
  INV_X1 U37456 ( .I(n55789), .ZN(n22859) );
  AOI21_X1 U37457 ( .A1(n64075), .A2(n54265), .B(n54264), .ZN(n21037) );
  NAND2_X1 U37458 ( .A1(n55652), .A2(n55651), .ZN(n16573) );
  AOI21_X1 U37459 ( .A1(n55153), .A2(n55113), .B(n55112), .ZN(n25684) );
  NAND2_X1 U37460 ( .A1(n16471), .A2(n50829), .ZN(n20376) );
  NAND2_X1 U37461 ( .A1(n9953), .A2(n57158), .ZN(n18802) );
  INV_X1 U37462 ( .I(n18804), .ZN(n18803) );
  NAND3_X1 U37463 ( .A1(n54264), .A2(n64075), .A3(n22545), .ZN(n54246) );
  AOI21_X1 U37464 ( .A1(n17110), .A2(n53493), .B(n17109), .ZN(n17108) );
  NOR2_X1 U37465 ( .A1(n17242), .A2(n53524), .ZN(n17100) );
  INV_X1 U37466 ( .I(n23882), .ZN(n53662) );
  AND2_X2 U37468 ( .A1(n32075), .A2(n21482), .Z(n15743) );
  AND2_X1 U37469 ( .A1(n61816), .A2(n43072), .Z(n15745) );
  INV_X1 U37471 ( .I(n16755), .ZN(n42486) );
  XNOR2_X1 U37473 ( .A1(n37979), .A2(n22452), .ZN(n15755) );
  AND2_X1 U37475 ( .A1(n24633), .A2(n5837), .Z(n15762) );
  NOR2_X2 U37476 ( .A1(n19999), .A2(n65216), .ZN(n15765) );
  OR2_X1 U37477 ( .A1(n21817), .A2(n21445), .Z(n15768) );
  AND2_X1 U37478 ( .A1(n53286), .A2(n16057), .Z(n15771) );
  OAI21_X1 U37479 ( .A1(n64493), .A2(n41460), .B(n23381), .ZN(n23380) );
  NOR2_X2 U37482 ( .A1(n17415), .A2(n26649), .ZN(n15791) );
  XOR2_X1 U37483 ( .A1(n25367), .A2(n37746), .Z(n15795) );
  AND2_X1 U37484 ( .A1(n54805), .A2(n54804), .Z(n15798) );
  INV_X1 U37488 ( .I(n24735), .ZN(n18930) );
  INV_X1 U37489 ( .I(n29451), .ZN(n29449) );
  INV_X1 U37490 ( .I(n54317), .ZN(n54073) );
  NAND2_X1 U37491 ( .A1(n1561), .A2(n31254), .ZN(n29889) );
  OR2_X1 U37495 ( .A1(n21614), .A2(n16290), .Z(n15836) );
  INV_X1 U37497 ( .I(n41831), .ZN(n42526) );
  NAND2_X1 U37498 ( .A1(n26208), .A2(n16539), .ZN(n49132) );
  XNOR2_X1 U37499 ( .A1(n32380), .A2(n32379), .ZN(n15841) );
  AND2_X1 U37502 ( .A1(n16981), .A2(n28034), .Z(n15845) );
  NOR2_X1 U37503 ( .A1(n24117), .A2(n58808), .ZN(n15846) );
  AND4_X1 U37504 ( .A1(n50040), .A2(n1637), .A3(n50039), .A4(n16915), .Z(
        n15850) );
  XNOR2_X1 U37507 ( .A1(n64360), .A2(n32106), .ZN(n15854) );
  AND2_X1 U37509 ( .A1(n29856), .A2(n29855), .Z(n15860) );
  BUF_X2 U37510 ( .I(n31508), .Z(n34083) );
  AND2_X1 U37511 ( .A1(n40049), .A2(n40103), .Z(n15861) );
  XOR2_X1 U37512 ( .A1(n24580), .A2(n21989), .Z(n15862) );
  AND2_X1 U37513 ( .A1(n54539), .A2(n4232), .Z(n15863) );
  XNOR2_X1 U37518 ( .A1(n61464), .A2(n51363), .ZN(n15881) );
  XOR2_X1 U37520 ( .A1(n51147), .A2(n51146), .Z(n15885) );
  XNOR2_X1 U37521 ( .A1(n38820), .A2(n14645), .ZN(n15888) );
  XNOR2_X1 U37522 ( .A1(n44959), .A2(n22340), .ZN(n15889) );
  INV_X2 U37523 ( .I(n52211), .ZN(n55727) );
  OR2_X1 U37527 ( .A1(n33439), .A2(n20978), .Z(n15907) );
  AND2_X1 U37528 ( .A1(n4993), .A2(n59841), .Z(n15908) );
  OR2_X1 U37529 ( .A1(n5569), .A2(n54996), .Z(n15909) );
  OR2_X1 U37533 ( .A1(n24767), .A2(n61707), .Z(n15913) );
  INV_X1 U37534 ( .I(n30006), .ZN(n30751) );
  OAI21_X1 U37535 ( .A1(n58307), .A2(n61708), .B(n16669), .ZN(n19642) );
  XOR2_X1 U37536 ( .A1(n52632), .A2(n52638), .Z(n15916) );
  NAND3_X1 U37537 ( .A1(n35428), .A2(n5936), .A3(n504), .ZN(n15917) );
  AOI21_X1 U37538 ( .A1(n41408), .A2(n41230), .B(n17063), .ZN(n40738) );
  AND2_X1 U37539 ( .A1(n56734), .A2(n56670), .Z(n15920) );
  AND2_X1 U37540 ( .A1(n56997), .A2(n57004), .Z(n15924) );
  INV_X1 U37542 ( .I(n18244), .ZN(n33645) );
  XNOR2_X1 U37545 ( .A1(n21680), .A2(n15950), .ZN(n15930) );
  OR2_X2 U37546 ( .A1(n20319), .A2(n53537), .Z(n15935) );
  INV_X2 U37548 ( .I(n29003), .ZN(n29506) );
  INV_X1 U37550 ( .I(n65228), .ZN(n42635) );
  XNOR2_X1 U37556 ( .A1(n45003), .A2(n45002), .ZN(n15960) );
  XNOR2_X1 U37558 ( .A1(n21365), .A2(n31974), .ZN(n15962) );
  XOR2_X1 U37559 ( .A1(n16681), .A2(n39465), .Z(n15963) );
  AND2_X1 U37561 ( .A1(n63874), .A2(n177), .Z(n15968) );
  AND2_X1 U37562 ( .A1(n23248), .A2(n7095), .Z(n15975) );
  AND2_X1 U37566 ( .A1(n56590), .A2(n64187), .Z(n15981) );
  OR2_X1 U37570 ( .A1(n56979), .A2(n56983), .Z(n15996) );
  AND2_X1 U37574 ( .A1(n32904), .A2(n20923), .Z(n16001) );
  AND2_X1 U37576 ( .A1(n46821), .A2(n47367), .Z(n16004) );
  XOR2_X1 U37577 ( .A1(n51520), .A2(n51519), .Z(n16006) );
  AND2_X1 U37578 ( .A1(n20122), .A2(n20118), .Z(n16007) );
  AND2_X1 U37579 ( .A1(n18861), .A2(n5056), .Z(n16008) );
  AND2_X1 U37581 ( .A1(n52130), .A2(n52129), .Z(n16010) );
  NAND2_X1 U37582 ( .A1(n25785), .A2(n27228), .ZN(n27486) );
  XOR2_X1 U37583 ( .A1(n39256), .A2(n39255), .Z(n16011) );
  OR2_X1 U37584 ( .A1(n30000), .A2(n23396), .Z(n16014) );
  OR2_X1 U37585 ( .A1(n55680), .A2(n20891), .Z(n16018) );
  INV_X1 U37586 ( .I(n28589), .ZN(n29636) );
  XNOR2_X1 U37589 ( .A1(n46614), .A2(n46613), .ZN(n16032) );
  XNOR2_X1 U37591 ( .A1(n50613), .A2(n50612), .ZN(n16034) );
  XNOR2_X1 U37592 ( .A1(n37610), .A2(n37569), .ZN(n16035) );
  INV_X1 U37593 ( .I(n18355), .ZN(n39475) );
  INV_X1 U37596 ( .I(n20431), .ZN(n37026) );
  XNOR2_X1 U37597 ( .A1(n58972), .A2(n16972), .ZN(n16039) );
  XNOR2_X1 U37598 ( .A1(n23126), .A2(n23571), .ZN(n16041) );
  XNOR2_X1 U37599 ( .A1(n17908), .A2(n25667), .ZN(n16045) );
  XNOR2_X1 U37600 ( .A1(n44918), .A2(n44917), .ZN(n16048) );
  XNOR2_X1 U37601 ( .A1(n18054), .A2(n37718), .ZN(n16049) );
  XNOR2_X1 U37602 ( .A1(n57586), .A2(n23987), .ZN(n16050) );
  AND2_X1 U37605 ( .A1(n30071), .A2(n30077), .Z(n16062) );
  AND2_X1 U37606 ( .A1(n49951), .A2(n48740), .Z(n16063) );
  AND2_X1 U37608 ( .A1(n28070), .A2(n22094), .Z(n16069) );
  INV_X1 U37609 ( .I(n21511), .ZN(n27295) );
  OR2_X1 U37612 ( .A1(n41396), .A2(n41395), .Z(n16081) );
  OR2_X1 U37613 ( .A1(n52267), .A2(n64424), .Z(n16086) );
  NOR2_X1 U37614 ( .A1(n24586), .A2(n65155), .ZN(n16091) );
  OR2_X1 U37615 ( .A1(n27602), .A2(n28314), .Z(n16094) );
  NOR2_X1 U37616 ( .A1(n33944), .A2(n139), .ZN(n16098) );
  INV_X1 U37618 ( .I(n25760), .ZN(n39995) );
  INV_X1 U37619 ( .I(n24472), .ZN(n55704) );
  NAND3_X1 U37623 ( .A1(n55855), .A2(n55885), .A3(n19307), .ZN(n55834) );
  INV_X1 U37624 ( .I(n55834), .ZN(n55881) );
  AND2_X1 U37626 ( .A1(n45913), .A2(n45912), .Z(n16109) );
  INV_X2 U37627 ( .I(n23829), .ZN(n28802) );
  INV_X1 U37629 ( .I(n65194), .ZN(n17425) );
  AND2_X1 U37631 ( .A1(n26561), .A2(n26560), .Z(n16113) );
  AND2_X1 U37632 ( .A1(n55695), .A2(n18292), .Z(n16117) );
  INV_X1 U37634 ( .I(n38924), .ZN(n41419) );
  INV_X1 U37637 ( .I(n11459), .ZN(n24523) );
  XNOR2_X1 U37638 ( .A1(n38411), .A2(n23680), .ZN(n16122) );
  XNOR2_X1 U37639 ( .A1(n21294), .A2(n31761), .ZN(n16123) );
  XNOR2_X1 U37641 ( .A1(n63004), .A2(n38978), .ZN(n16125) );
  XNOR2_X1 U37642 ( .A1(n14038), .A2(n46576), .ZN(n16126) );
  XNOR2_X1 U37643 ( .A1(n32589), .A2(n32588), .ZN(n16128) );
  OR2_X1 U37648 ( .A1(n26800), .A2(n63533), .Z(n16136) );
  XNOR2_X1 U37650 ( .A1(n61610), .A2(n31916), .ZN(n16142) );
  AND2_X1 U37652 ( .A1(n34454), .A2(n36756), .Z(n16153) );
  AND2_X1 U37653 ( .A1(n40354), .A2(n40353), .Z(n16154) );
  INV_X4 U37654 ( .I(n18087), .ZN(n43516) );
  AND2_X1 U37656 ( .A1(n27023), .A2(n27024), .Z(n16172) );
  AND2_X1 U37657 ( .A1(n40134), .A2(n40135), .Z(n16173) );
  NOR2_X1 U37660 ( .A1(n47455), .A2(n47454), .ZN(n16177) );
  OR2_X1 U37661 ( .A1(n23252), .A2(n16619), .Z(n16184) );
  OR2_X1 U37663 ( .A1(n16588), .A2(n16587), .Z(n16187) );
  INV_X1 U37664 ( .I(n17902), .ZN(n46208) );
  NAND2_X1 U37665 ( .A1(n49299), .A2(n9177), .ZN(n16188) );
  INV_X1 U37666 ( .I(n7225), .ZN(n26026) );
  AND2_X1 U37667 ( .A1(n49687), .A2(n62248), .Z(n16193) );
  INV_X1 U37668 ( .I(n47456), .ZN(n48755) );
  XNOR2_X1 U37671 ( .A1(n45139), .A2(n46592), .ZN(n16195) );
  INV_X1 U37675 ( .I(n35071), .ZN(n36749) );
  BUF_X4 U37676 ( .I(n35071), .Z(n36742) );
  XNOR2_X1 U37679 ( .A1(n39766), .A2(n37990), .ZN(n16205) );
  XNOR2_X1 U37680 ( .A1(n38174), .A2(n38173), .ZN(n16206) );
  XNOR2_X1 U37682 ( .A1(n36369), .A2(n38170), .ZN(n16207) );
  XNOR2_X1 U37683 ( .A1(n18516), .A2(n51631), .ZN(n16208) );
  XNOR2_X1 U37686 ( .A1(n37462), .A2(n37461), .ZN(n16209) );
  XNOR2_X1 U37687 ( .A1(Ciphertext[135]), .A2(Ciphertext[132]), .ZN(n16210) );
  XNOR2_X1 U37688 ( .A1(n25161), .A2(n38942), .ZN(n16213) );
  INV_X1 U37692 ( .I(n36493), .ZN(n36238) );
  AND2_X1 U37693 ( .A1(n57852), .A2(n4760), .Z(n16230) );
  AND2_X1 U37694 ( .A1(n43742), .A2(n43741), .Z(n16232) );
  NAND2_X1 U37696 ( .A1(n42167), .A2(n295), .ZN(n16237) );
  OAI21_X1 U37697 ( .A1(n37361), .A2(n37359), .B(n4541), .ZN(n37116) );
  XNOR2_X1 U37700 ( .A1(n32048), .A2(n45403), .ZN(n16246) );
  XNOR2_X1 U37701 ( .A1(n44530), .A2(n44529), .ZN(n16247) );
  XNOR2_X1 U37704 ( .A1(n39438), .A2(n39437), .ZN(n16250) );
  XNOR2_X1 U37705 ( .A1(n38118), .A2(n968), .ZN(n16251) );
  XNOR2_X1 U37706 ( .A1(n32492), .A2(n33839), .ZN(n16252) );
  INV_X1 U37708 ( .I(n35803), .ZN(n34224) );
  INV_X1 U37711 ( .I(n31841), .ZN(n35810) );
  INV_X1 U37712 ( .I(n27329), .ZN(n29367) );
  NAND2_X1 U37713 ( .A1(n27435), .A2(n28806), .ZN(n27329) );
  NAND2_X1 U37715 ( .A1(n40776), .A2(n64462), .ZN(n43502) );
  NAND2_X1 U37716 ( .A1(n35294), .A2(n32222), .ZN(n16267) );
  INV_X1 U37718 ( .I(n23583), .ZN(n22170) );
  BUF_X2 U37719 ( .I(n45115), .Z(n24030) );
  XNOR2_X1 U37720 ( .A1(n46229), .A2(n44968), .ZN(n16270) );
  XNOR2_X1 U37721 ( .A1(n23181), .A2(n16404), .ZN(n16271) );
  INV_X1 U37722 ( .I(n61717), .ZN(n47895) );
  XNOR2_X1 U37725 ( .A1(n51746), .A2(n51745), .ZN(n16274) );
  INV_X1 U37726 ( .I(n48770), .ZN(n18185) );
  INV_X1 U37729 ( .I(n4591), .ZN(n33743) );
  INV_X1 U37731 ( .I(n18969), .ZN(n18984) );
  INV_X1 U37735 ( .I(n52986), .ZN(n54490) );
  INV_X2 U37736 ( .I(n53809), .ZN(n53794) );
  INV_X1 U37737 ( .I(n59125), .ZN(n33538) );
  XNOR2_X1 U37743 ( .A1(n33261), .A2(n33262), .ZN(n16287) );
  XOR2_X1 U37744 ( .A1(n38576), .A2(n39625), .Z(n16288) );
  INV_X1 U37746 ( .I(n48818), .ZN(n24788) );
  INV_X2 U37747 ( .I(n27479), .ZN(n27483) );
  XNOR2_X1 U37749 ( .A1(n46550), .A2(n44964), .ZN(n16293) );
  OR2_X1 U37750 ( .A1(n37623), .A2(n37622), .Z(n16295) );
  XOR2_X1 U37753 ( .A1(n44414), .A2(n32167), .Z(n16299) );
  INV_X1 U37754 ( .I(n47902), .ZN(n24290) );
  XNOR2_X1 U37755 ( .A1(n35541), .A2(n25277), .ZN(n16300) );
  INV_X1 U37762 ( .I(n53860), .ZN(n53624) );
  INV_X1 U37763 ( .I(n38493), .ZN(n40661) );
  XNOR2_X1 U37764 ( .A1(n51680), .A2(n32161), .ZN(n16302) );
  XNOR2_X1 U37765 ( .A1(n31618), .A2(n38430), .ZN(n16303) );
  BUF_X2 U37766 ( .I(n37492), .Z(n23842) );
  XOR2_X1 U37767 ( .A1(n16404), .A2(n39220), .Z(n16304) );
  XNOR2_X1 U37768 ( .A1(n45278), .A2(n31771), .ZN(n16305) );
  XNOR2_X1 U37771 ( .A1(n50102), .A2(n43759), .ZN(n16307) );
  XOR2_X1 U37772 ( .A1(n32274), .A2(n24920), .Z(n16308) );
  INV_X2 U37773 ( .I(n25569), .ZN(n34127) );
  XNOR2_X1 U37776 ( .A1(n31948), .A2(n46603), .ZN(n16309) );
  XNOR2_X1 U37777 ( .A1(n32303), .A2(n43588), .ZN(n16310) );
  BUF_X2 U37778 ( .I(Key[32]), .Z(n23882) );
  BUF_X2 U37779 ( .I(Key[44]), .Z(n53805) );
  XNOR2_X1 U37781 ( .A1(n49877), .A2(n34835), .ZN(n16311) );
  XNOR2_X1 U37782 ( .A1(n37760), .A2(n52150), .ZN(n16312) );
  XNOR2_X1 U37783 ( .A1(n51142), .A2(n48967), .ZN(n16313) );
  XNOR2_X1 U37784 ( .A1(n52003), .A2(n49403), .ZN(n16314) );
  XNOR2_X1 U37785 ( .A1(n52182), .A2(n37995), .ZN(n16315) );
  XNOR2_X1 U37786 ( .A1(n51642), .A2(n38854), .ZN(n16316) );
  XNOR2_X1 U37788 ( .A1(n45340), .A2(n45339), .ZN(n16317) );
  XNOR2_X1 U37789 ( .A1(n45372), .A2(n45371), .ZN(n16318) );
  XNOR2_X1 U37790 ( .A1(n50987), .A2(n42021), .ZN(n16319) );
  XNOR2_X1 U37791 ( .A1(n46417), .A2(n46416), .ZN(n16320) );
  XNOR2_X1 U37792 ( .A1(n45317), .A2(n56335), .ZN(n16321) );
  XNOR2_X1 U37793 ( .A1(n44271), .A2(n51278), .ZN(n16322) );
  XNOR2_X1 U37794 ( .A1(n43195), .A2(n43194), .ZN(n16323) );
  XNOR2_X1 U37795 ( .A1(n39536), .A2(n31794), .ZN(n16324) );
  INV_X1 U37796 ( .I(n45404), .ZN(n17129) );
  BUF_X2 U37797 ( .I(Key[40]), .Z(n53764) );
  XNOR2_X1 U37798 ( .A1(n51188), .A2(n51187), .ZN(n16325) );
  XNOR2_X1 U37799 ( .A1(n50228), .A2(n50227), .ZN(n16326) );
  XNOR2_X1 U37800 ( .A1(n50573), .A2(n50572), .ZN(n16327) );
  XNOR2_X1 U37801 ( .A1(n51935), .A2(n51934), .ZN(n16328) );
  BUF_X2 U37802 ( .I(Key[6]), .Z(n51493) );
  INV_X1 U37803 ( .I(n51493), .ZN(n16709) );
  BUF_X2 U37805 ( .I(Key[120]), .Z(n52226) );
  INV_X1 U37806 ( .I(n53705), .ZN(n17221) );
  NOR3_X2 U37807 ( .A1(n16329), .A2(n57013), .A3(n56545), .ZN(n57009) );
  NAND2_X1 U37808 ( .A1(n16329), .A2(n56530), .ZN(n17198) );
  OAI21_X1 U37809 ( .A1(n16329), .A2(n22870), .B(n56530), .ZN(n52245) );
  OAI21_X2 U37811 ( .A1(n16332), .A2(n15951), .B(n16330), .ZN(n18174) );
  NAND2_X2 U37813 ( .A1(n24553), .A2(n51902), .ZN(n56432) );
  NAND2_X2 U37814 ( .A1(n26208), .A2(n16336), .ZN(n49986) );
  NAND2_X1 U37819 ( .A1(n55715), .A2(n56424), .ZN(n16344) );
  XOR2_X1 U37824 ( .A1(n2167), .A2(n52116), .Z(n16349) );
  NAND2_X2 U37826 ( .A1(n37436), .A2(n37426), .ZN(n35946) );
  XOR2_X1 U37828 ( .A1(n32514), .A2(n16361), .Z(n16360) );
  XOR2_X1 U37833 ( .A1(n33190), .A2(n16366), .Z(n16365) );
  XOR2_X1 U37834 ( .A1(n16368), .A2(n32100), .Z(n16367) );
  XOR2_X1 U37835 ( .A1(n22227), .A2(n29407), .Z(n32202) );
  XOR2_X1 U37836 ( .A1(n17668), .A2(n5436), .Z(n16368) );
  XOR2_X1 U37838 ( .A1(n16476), .A2(n16304), .Z(n16370) );
  NOR3_X1 U37844 ( .A1(n24613), .A2(n16595), .A3(n57608), .ZN(n48399) );
  INV_X2 U37847 ( .I(n17798), .ZN(n16383) );
  NAND3_X1 U37849 ( .A1(n16017), .A2(n1738), .A3(n40086), .ZN(n16391) );
  XOR2_X1 U37851 ( .A1(n21094), .A2(n16302), .Z(n32162) );
  XOR2_X1 U37852 ( .A1(n24943), .A2(n21094), .Z(n33023) );
  NOR2_X2 U37854 ( .A1(n1426), .A2(n23717), .ZN(n35769) );
  XOR2_X1 U37855 ( .A1(n9896), .A2(n16404), .Z(n18540) );
  XOR2_X1 U37856 ( .A1(n39671), .A2(n16404), .Z(n39672) );
  NAND2_X2 U37857 ( .A1(n6095), .A2(n55017), .ZN(n26200) );
  NAND4_X2 U37862 ( .A1(n33441), .A2(n15907), .A3(n16422), .A4(n16421), .ZN(
        n16420) );
  XOR2_X1 U37865 ( .A1(n46121), .A2(n46122), .Z(n46546) );
  NAND2_X2 U37868 ( .A1(n53726), .A2(n53729), .ZN(n53752) );
  NOR2_X2 U37869 ( .A1(n17261), .A2(n17256), .ZN(n53729) );
  OAI21_X1 U37871 ( .A1(n24286), .A2(n33573), .B(n35662), .ZN(n33575) );
  INV_X2 U37873 ( .I(n24378), .ZN(n24286) );
  XOR2_X1 U37875 ( .A1(n16430), .A2(n46200), .Z(n16428) );
  XOR2_X1 U37876 ( .A1(n62065), .A2(n57918), .Z(n46200) );
  XOR2_X1 U37877 ( .A1(n673), .A2(n46199), .Z(n16430) );
  XOR2_X1 U37878 ( .A1(n46706), .A2(n46190), .Z(n16431) );
  XOR2_X1 U37879 ( .A1(n920), .A2(n38786), .Z(n39647) );
  NAND2_X2 U37881 ( .A1(n20747), .A2(n26084), .ZN(n31092) );
  NAND2_X1 U37887 ( .A1(n16461), .A2(n21229), .ZN(n41121) );
  NOR2_X1 U37888 ( .A1(n16461), .A2(n41379), .ZN(n41124) );
  INV_X2 U37892 ( .I(n16470), .ZN(n28509) );
  NAND2_X1 U37893 ( .A1(n16470), .A2(n1568), .ZN(n28515) );
  OAI21_X1 U37897 ( .A1(n42412), .A2(n16480), .B(n1193), .ZN(n42418) );
  NAND2_X1 U37898 ( .A1(n16481), .A2(n61458), .ZN(n17140) );
  NAND2_X1 U37899 ( .A1(n35802), .A2(n16481), .ZN(n34389) );
  AOI21_X1 U37900 ( .A1(n18848), .A2(n28517), .B(n25858), .ZN(n16485) );
  NAND2_X2 U37901 ( .A1(n28510), .A2(n23753), .ZN(n18848) );
  NAND2_X1 U37904 ( .A1(n42968), .A2(n57198), .ZN(n41755) );
  NAND2_X2 U37905 ( .A1(n13478), .A2(n43464), .ZN(n41757) );
  OAI21_X1 U37906 ( .A1(n39920), .A2(n16497), .B(n16496), .ZN(n39924) );
  NAND2_X1 U37907 ( .A1(n42428), .A2(n16497), .ZN(n16496) );
  NAND2_X2 U37909 ( .A1(n40308), .A2(n40063), .ZN(n16497) );
  INV_X1 U37911 ( .I(n38292), .ZN(n17938) );
  NOR2_X1 U37912 ( .A1(n55381), .A2(n16503), .ZN(n23129) );
  NOR2_X1 U37913 ( .A1(n29774), .A2(n16504), .ZN(n18101) );
  XOR2_X1 U37918 ( .A1(n39453), .A2(n16513), .Z(n16657) );
  XOR2_X1 U37921 ( .A1(n39448), .A2(n39447), .Z(n16514) );
  OAI21_X1 U37926 ( .A1(n27550), .A2(n16523), .B(n27549), .ZN(n27551) );
  NOR2_X1 U37928 ( .A1(n16525), .A2(n10125), .ZN(n27832) );
  OAI22_X1 U37929 ( .A1(n26393), .A2(n28483), .B1(n16525), .B2(n18006), .ZN(
        n26394) );
  NAND2_X2 U37932 ( .A1(n17589), .A2(n28485), .ZN(n16525) );
  NAND2_X1 U37933 ( .A1(n16526), .A2(n14820), .ZN(n41251) );
  NAND3_X1 U37935 ( .A1(n16806), .A2(n42287), .A3(n16526), .ZN(n16803) );
  NOR2_X1 U37936 ( .A1(n50004), .A2(n6977), .ZN(n49138) );
  NAND2_X1 U37937 ( .A1(n23394), .A2(n6977), .ZN(n49473) );
  XOR2_X1 U37938 ( .A1(n62323), .A2(n31008), .Z(n31009) );
  XOR2_X1 U37941 ( .A1(n16536), .A2(n39240), .Z(n16535) );
  XOR2_X1 U37944 ( .A1(n38782), .A2(n24147), .Z(n39233) );
  NAND2_X1 U37945 ( .A1(n18273), .A2(n34386), .ZN(n16556) );
  XOR2_X1 U37946 ( .A1(n15698), .A2(n15766), .Z(n44434) );
  XOR2_X1 U37948 ( .A1(n16346), .A2(n38470), .Z(n16559) );
  AND3_X1 U37950 ( .A1(n16565), .A2(n16564), .A3(n16562), .Z(n16626) );
  NOR2_X1 U37951 ( .A1(n16567), .A2(n37291), .ZN(n16566) );
  NAND2_X1 U37952 ( .A1(n22823), .A2(n22822), .ZN(n16567) );
  INV_X1 U37954 ( .I(n16571), .ZN(n48911) );
  NAND3_X2 U37957 ( .A1(n27552), .A2(n27553), .A3(n27551), .ZN(n27626) );
  NOR2_X1 U37958 ( .A1(n49712), .A2(n16586), .ZN(n16587) );
  OR2_X1 U37959 ( .A1(n18469), .A2(n6633), .Z(n16591) );
  INV_X2 U37960 ( .I(n17913), .ZN(n31385) );
  NOR3_X2 U37961 ( .A1(n25852), .A2(n25853), .A3(n15861), .ZN(n20893) );
  NAND2_X2 U37962 ( .A1(n36979), .A2(n23742), .ZN(n37227) );
  NAND2_X1 U37964 ( .A1(n11243), .A2(n60693), .ZN(n39511) );
  AOI21_X1 U37965 ( .A1(n29460), .A2(n29455), .B(n60028), .ZN(n28100) );
  NAND2_X1 U37973 ( .A1(n34770), .A2(n59724), .ZN(n34774) );
  NOR2_X1 U37978 ( .A1(n32512), .A2(n16856), .ZN(n16614) );
  XOR2_X1 U37980 ( .A1(n26025), .A2(n16196), .Z(n16618) );
  INV_X1 U37981 ( .I(n21728), .ZN(n57036) );
  NAND2_X1 U37982 ( .A1(n17555), .A2(n25160), .ZN(n21728) );
  OAI21_X1 U37985 ( .A1(n27984), .A2(n27985), .B(n1320), .ZN(n18530) );
  OAI22_X1 U37987 ( .A1(n46991), .A2(n16628), .B1(n48212), .B2(n63913), .ZN(
        n46992) );
  NAND2_X1 U37988 ( .A1(n18569), .A2(n16628), .ZN(n48670) );
  MUX2_X1 U37990 ( .I0(n43395), .I1(n43034), .S(n62326), .Z(n43035) );
  XOR2_X1 U37993 ( .A1(n49817), .A2(n15735), .Z(n16641) );
  NOR2_X2 U37995 ( .A1(n37454), .A2(n37233), .ZN(n37446) );
  NAND2_X2 U37997 ( .A1(n35850), .A2(n23160), .ZN(n37441) );
  NAND2_X1 U37999 ( .A1(n18129), .A2(n21887), .ZN(n24163) );
  INV_X2 U38000 ( .I(n16657), .ZN(n23933) );
  NOR2_X2 U38004 ( .A1(n34095), .A2(n16662), .ZN(n38988) );
  NOR2_X1 U38008 ( .A1(n28375), .A2(n10419), .ZN(n26625) );
  XOR2_X1 U38010 ( .A1(n16668), .A2(n33838), .Z(n17510) );
  XOR2_X1 U38011 ( .A1(n20623), .A2(n52327), .Z(n16668) );
  OR2_X2 U38013 ( .A1(n24834), .A2(n15963), .Z(n40441) );
  XOR2_X1 U38014 ( .A1(n25377), .A2(n25374), .Z(n38878) );
  NAND2_X2 U38019 ( .A1(n56547), .A2(n56544), .ZN(n57013) );
  NAND2_X2 U38021 ( .A1(n53820), .A2(n58811), .ZN(n53826) );
  NOR2_X2 U38022 ( .A1(n13504), .A2(n58811), .ZN(n53811) );
  OAI21_X1 U38025 ( .A1(n28558), .A2(n16707), .B(n16812), .ZN(n28559) );
  NOR2_X2 U38029 ( .A1(n17302), .A2(n17303), .ZN(n20371) );
  NOR2_X1 U38032 ( .A1(n50004), .A2(n16712), .ZN(n16711) );
  NAND2_X2 U38039 ( .A1(n53483), .A2(n53516), .ZN(n53501) );
  INV_X2 U38040 ( .I(n25676), .ZN(n53516) );
  NAND2_X1 U38041 ( .A1(n16718), .A2(n48665), .ZN(n46259) );
  NOR2_X1 U38042 ( .A1(n20788), .A2(n16717), .ZN(n46993) );
  NAND2_X1 U38043 ( .A1(n48199), .A2(n48668), .ZN(n16717) );
  OAI21_X1 U38044 ( .A1(n20788), .A2(n16718), .B(n48668), .ZN(n48669) );
  NAND3_X2 U38046 ( .A1(n16727), .A2(n16725), .A3(n16719), .ZN(n34846) );
  NOR2_X1 U38047 ( .A1(n12184), .A2(n35786), .ZN(n16721) );
  NAND2_X1 U38048 ( .A1(n12184), .A2(n16724), .ZN(n16723) );
  NAND3_X1 U38049 ( .A1(n25313), .A2(n49490), .A3(n16730), .ZN(n25312) );
  NAND2_X2 U38050 ( .A1(n17924), .A2(n17923), .ZN(n39275) );
  NAND3_X1 U38054 ( .A1(n34362), .A2(n37273), .A3(n37136), .ZN(n16734) );
  XOR2_X1 U38056 ( .A1(n64945), .A2(n46592), .Z(n17520) );
  XOR2_X1 U38057 ( .A1(n16741), .A2(n25530), .Z(n46592) );
  XOR2_X1 U38058 ( .A1(n57892), .A2(n25531), .Z(n16741) );
  OAI21_X1 U38059 ( .A1(n59859), .A2(n16742), .B(n25477), .ZN(n45635) );
  NAND2_X2 U38060 ( .A1(n25429), .A2(n24047), .ZN(n16742) );
  NAND2_X2 U38061 ( .A1(n49177), .A2(n20600), .ZN(n16745) );
  NAND2_X1 U38063 ( .A1(n20844), .A2(n1493), .ZN(n21666) );
  NAND2_X1 U38064 ( .A1(n43117), .A2(n1493), .ZN(n43119) );
  XOR2_X1 U38069 ( .A1(n16758), .A2(n30932), .Z(n30933) );
  XOR2_X1 U38070 ( .A1(n16758), .A2(n33073), .Z(n33074) );
  XOR2_X1 U38071 ( .A1(n32121), .A2(n16758), .Z(n32122) );
  XOR2_X1 U38072 ( .A1(n32011), .A2(n16758), .Z(n31880) );
  XOR2_X1 U38073 ( .A1(n16761), .A2(n16762), .Z(n16760) );
  XOR2_X1 U38074 ( .A1(n51790), .A2(n50265), .Z(n16761) );
  XOR2_X1 U38075 ( .A1(n50266), .A2(n354), .Z(n16762) );
  NAND2_X1 U38076 ( .A1(n4428), .A2(n46716), .ZN(n48109) );
  NAND2_X1 U38077 ( .A1(n48533), .A2(n4428), .ZN(n48233) );
  NAND2_X2 U38079 ( .A1(n29188), .A2(n14451), .ZN(n17285) );
  OR2_X1 U38082 ( .A1(n57029), .A2(n16770), .Z(n16769) );
  XOR2_X1 U38084 ( .A1(n39259), .A2(n37694), .Z(n37695) );
  NOR2_X1 U38085 ( .A1(n16882), .A2(n16783), .ZN(n24128) );
  INV_X1 U38086 ( .I(n27231), .ZN(n16786) );
  NOR3_X1 U38087 ( .A1(n27229), .A2(n26705), .A3(n23823), .ZN(n16787) );
  NAND2_X1 U38089 ( .A1(n16788), .A2(n20519), .ZN(n27477) );
  INV_X2 U38091 ( .I(n26091), .ZN(n27661) );
  NAND4_X2 U38097 ( .A1(n16802), .A2(n16803), .A3(n16804), .A4(n16881), .ZN(
        n42313) );
  XOR2_X1 U38098 ( .A1(n16809), .A2(n15865), .Z(n32634) );
  INV_X2 U38100 ( .I(n16813), .ZN(n57075) );
  NAND2_X1 U38103 ( .A1(n10874), .A2(n23912), .ZN(n48960) );
  NAND2_X1 U38104 ( .A1(n39992), .A2(n12158), .ZN(n41394) );
  NAND2_X1 U38106 ( .A1(n10074), .A2(n12158), .ZN(n40427) );
  XOR2_X1 U38109 ( .A1(n59355), .A2(n31850), .Z(n32305) );
  NOR2_X2 U38113 ( .A1(n16838), .A2(n16837), .ZN(n20600) );
  NAND2_X2 U38114 ( .A1(n16836), .A2(n61668), .ZN(n48199) );
  NAND2_X2 U38115 ( .A1(n55261), .A2(n24870), .ZN(n55275) );
  INV_X4 U38122 ( .I(n25071), .ZN(n42404) );
  NAND2_X2 U38123 ( .A1(n16853), .A2(n25069), .ZN(n25071) );
  INV_X1 U38124 ( .I(n16939), .ZN(n33703) );
  XOR2_X1 U38130 ( .A1(n16207), .A2(n13695), .Z(n36371) );
  XOR2_X1 U38131 ( .A1(n16873), .A2(n16872), .Z(n17018) );
  XOR2_X1 U38132 ( .A1(n1549), .A2(n16275), .Z(n16872) );
  XOR2_X1 U38134 ( .A1(n9628), .A2(n44748), .Z(n16883) );
  NAND2_X1 U38135 ( .A1(n16885), .A2(n36870), .ZN(n37395) );
  XOR2_X1 U38137 ( .A1(n16893), .A2(n17999), .Z(n16892) );
  XOR2_X1 U38138 ( .A1(n61732), .A2(n32164), .Z(n31641) );
  XOR2_X1 U38140 ( .A1(n16895), .A2(n7225), .Z(n21823) );
  XOR2_X1 U38141 ( .A1(n59355), .A2(n129), .Z(n16895) );
  NAND2_X2 U38142 ( .A1(n29830), .A2(n16896), .ZN(n31590) );
  XOR2_X1 U38143 ( .A1(n19511), .A2(n1679), .Z(n16899) );
  INV_X2 U38145 ( .I(n25209), .ZN(n46621) );
  XOR2_X1 U38146 ( .A1(n31950), .A2(n16951), .Z(n16901) );
  XOR2_X1 U38147 ( .A1(n46196), .A2(n50494), .Z(n43940) );
  XOR2_X1 U38148 ( .A1(n46196), .A2(n55335), .Z(n44121) );
  AND2_X1 U38149 ( .A1(n28065), .A2(n26529), .Z(n25546) );
  NAND2_X1 U38150 ( .A1(n35313), .A2(n35320), .ZN(n16904) );
  NAND2_X1 U38153 ( .A1(n16911), .A2(n15540), .ZN(n43294) );
  NOR3_X1 U38154 ( .A1(n17755), .A2(n59709), .A3(n16911), .ZN(n16941) );
  NAND2_X1 U38156 ( .A1(n63438), .A2(n30334), .ZN(n30639) );
  NOR2_X1 U38157 ( .A1(n13144), .A2(n63438), .ZN(n30335) );
  NAND2_X1 U38159 ( .A1(n20199), .A2(n50042), .ZN(n16915) );
  INV_X2 U38167 ( .I(n26067), .ZN(n18473) );
  NAND2_X2 U38169 ( .A1(n45538), .A2(n21755), .ZN(n47028) );
  AOI21_X1 U38172 ( .A1(n33701), .A2(n59681), .B(n16939), .ZN(n33571) );
  XOR2_X1 U38176 ( .A1(n16944), .A2(n52532), .Z(n55248) );
  XOR2_X1 U38177 ( .A1(n16947), .A2(n16945), .Z(n16944) );
  NAND3_X1 U38179 ( .A1(n55406), .A2(n55407), .A3(n10551), .ZN(n55408) );
  NAND3_X1 U38180 ( .A1(n55417), .A2(n55416), .A3(n10551), .ZN(n55420) );
  NAND2_X2 U38181 ( .A1(n55397), .A2(n55250), .ZN(n16948) );
  NAND2_X1 U38182 ( .A1(n48102), .A2(n16950), .ZN(n47116) );
  OAI21_X1 U38183 ( .A1(n23099), .A2(n21304), .B(n16950), .ZN(n46759) );
  NAND2_X2 U38184 ( .A1(n38021), .A2(n19990), .ZN(n23711) );
  AOI21_X2 U38186 ( .A1(n16966), .A2(n16965), .B(n44487), .ZN(n16963) );
  OAI22_X1 U38189 ( .A1(n61048), .A2(n30451), .B1(n60162), .B2(n4999), .ZN(
        n19028) );
  OAI22_X1 U38190 ( .A1(n28287), .A2(n16971), .B1(n21159), .B2(n21095), .ZN(
        n28288) );
  NOR2_X2 U38191 ( .A1(n36193), .A2(n16968), .ZN(n36413) );
  INV_X2 U38193 ( .I(n18004), .ZN(n20753) );
  NOR2_X1 U38197 ( .A1(n16980), .A2(n41103), .ZN(n41108) );
  NAND2_X1 U38198 ( .A1(n19765), .A2(n24609), .ZN(n35949) );
  XOR2_X1 U38202 ( .A1(n52333), .A2(n23128), .Z(n52339) );
  XOR2_X1 U38203 ( .A1(n51688), .A2(n16984), .Z(n52333) );
  XOR2_X1 U38209 ( .A1(n21233), .A2(n21232), .Z(n17002) );
  NAND2_X1 U38210 ( .A1(n49438), .A2(n1637), .ZN(n49439) );
  NOR2_X2 U38212 ( .A1(n5873), .A2(n25396), .ZN(n37064) );
  XOR2_X1 U38213 ( .A1(n1200), .A2(n39624), .Z(n21234) );
  NAND2_X1 U38214 ( .A1(n17003), .A2(n52786), .ZN(n52816) );
  OAI21_X1 U38216 ( .A1(n833), .A2(n17003), .B(n57037), .ZN(n57038) );
  NOR2_X1 U38219 ( .A1(n6530), .A2(n15807), .ZN(n35620) );
  NOR2_X2 U38221 ( .A1(n53368), .A2(n17012), .ZN(n53334) );
  XOR2_X1 U38225 ( .A1(n21581), .A2(n33230), .Z(n17024) );
  XOR2_X1 U38226 ( .A1(n6322), .A2(n62658), .Z(n17025) );
  XOR2_X1 U38227 ( .A1(n17119), .A2(n33840), .Z(n32077) );
  XOR2_X1 U38228 ( .A1(n17120), .A2(n32083), .Z(n17026) );
  NAND2_X2 U38230 ( .A1(n37269), .A2(n58580), .ZN(n17030) );
  OAI21_X1 U38232 ( .A1(n23990), .A2(n46914), .B(n1070), .ZN(n17034) );
  INV_X2 U38233 ( .I(n18277), .ZN(n34196) );
  INV_X1 U38234 ( .I(n25326), .ZN(n17042) );
  XOR2_X1 U38236 ( .A1(n11070), .A2(n50667), .Z(n50668) );
  INV_X2 U38240 ( .I(n17058), .ZN(n57074) );
  INV_X4 U38243 ( .I(n63014), .ZN(n20888) );
  NAND2_X1 U38245 ( .A1(n17072), .A2(n50041), .ZN(n50040) );
  NAND2_X2 U38246 ( .A1(n50044), .A2(n9799), .ZN(n50039) );
  NAND2_X2 U38247 ( .A1(n37268), .A2(n37269), .ZN(n18969) );
  XOR2_X1 U38250 ( .A1(n17102), .A2(n44126), .Z(n44127) );
  XOR2_X1 U38251 ( .A1(n17102), .A2(n44173), .Z(n44174) );
  XOR2_X1 U38252 ( .A1(n17102), .A2(n18726), .Z(n17160) );
  NAND3_X1 U38253 ( .A1(n17103), .A2(n28267), .A3(n17909), .ZN(n28268) );
  XOR2_X1 U38254 ( .A1(n17105), .A2(n17104), .Z(n32098) );
  XOR2_X1 U38255 ( .A1(n19348), .A2(n24943), .Z(n17119) );
  INV_X2 U38256 ( .I(n5458), .ZN(n38577) );
  NOR2_X1 U38260 ( .A1(n45549), .A2(n24114), .ZN(n17137) );
  NAND2_X1 U38262 ( .A1(n10526), .A2(n17140), .ZN(n17139) );
  NOR2_X1 U38263 ( .A1(n10526), .A2(n35799), .ZN(n34227) );
  AOI21_X1 U38266 ( .A1(n34295), .A2(n17141), .B(n31844), .ZN(n31845) );
  INV_X4 U38269 ( .I(n54717), .ZN(n54767) );
  AOI21_X1 U38270 ( .A1(n62106), .A2(n40443), .B(n41106), .ZN(n18416) );
  NAND2_X2 U38271 ( .A1(n17148), .A2(n34233), .ZN(n35822) );
  NAND2_X1 U38272 ( .A1(n17148), .A2(n22633), .ZN(n34318) );
  NAND2_X1 U38273 ( .A1(n17148), .A2(n35820), .ZN(n34707) );
  NAND3_X1 U38274 ( .A1(n35308), .A2(n35309), .A3(n17148), .ZN(n35310) );
  NAND2_X1 U38281 ( .A1(n43462), .A2(n62686), .ZN(n42417) );
  NOR2_X1 U38282 ( .A1(n20038), .A2(n62686), .ZN(n20037) );
  NAND2_X2 U38283 ( .A1(n18501), .A2(n18500), .ZN(n18401) );
  NAND2_X2 U38284 ( .A1(n25576), .A2(n40875), .ZN(n46187) );
  NAND2_X2 U38285 ( .A1(n17151), .A2(n17150), .ZN(n44909) );
  XOR2_X1 U38287 ( .A1(n17154), .A2(n38106), .Z(n38158) );
  XOR2_X1 U38288 ( .A1(n17347), .A2(n17154), .Z(n38486) );
  XOR2_X1 U38289 ( .A1(n17220), .A2(n17154), .Z(n17218) );
  NAND4_X2 U38290 ( .A1(n15970), .A2(n21543), .A3(n21542), .A4(n21541), .ZN(
        n37583) );
  NAND3_X2 U38292 ( .A1(n29069), .A2(n29068), .A3(n18356), .ZN(n22244) );
  XOR2_X1 U38295 ( .A1(n17160), .A2(n17161), .Z(n17157) );
  XOR2_X1 U38297 ( .A1(n20271), .A2(n45052), .Z(n17159) );
  XOR2_X1 U38298 ( .A1(n45051), .A2(n45047), .Z(n17161) );
  XOR2_X1 U38303 ( .A1(n24257), .A2(n39343), .Z(n39344) );
  XOR2_X1 U38304 ( .A1(n17164), .A2(n38784), .Z(n38785) );
  XOR2_X1 U38305 ( .A1(n17164), .A2(n37506), .Z(n37507) );
  XOR2_X1 U38306 ( .A1(n38373), .A2(n17164), .Z(n38540) );
  NOR2_X1 U38308 ( .A1(n22934), .A2(n8182), .ZN(n29717) );
  XOR2_X1 U38310 ( .A1(n31858), .A2(n31738), .Z(n31740) );
  XOR2_X1 U38311 ( .A1(n31858), .A2(n31331), .Z(n31332) );
  AND2_X1 U38314 ( .A1(n60885), .A2(n60993), .Z(n28021) );
  XOR2_X1 U38318 ( .A1(n17171), .A2(n50858), .Z(n50859) );
  XOR2_X1 U38319 ( .A1(n52340), .A2(n17171), .Z(n19430) );
  XOR2_X1 U38321 ( .A1(n17171), .A2(n9635), .Z(n50940) );
  NOR2_X2 U38325 ( .A1(n42464), .A2(n17184), .ZN(n42986) );
  XOR2_X1 U38326 ( .A1(n1548), .A2(n31741), .Z(n31742) );
  NAND3_X1 U38328 ( .A1(n33111), .A2(n22454), .A3(n58924), .ZN(n17197) );
  NAND2_X1 U38329 ( .A1(n17720), .A2(n63593), .ZN(n24725) );
  NOR3_X1 U38331 ( .A1(n18216), .A2(n24721), .A3(n63593), .ZN(n24723) );
  NOR2_X1 U38334 ( .A1(n14561), .A2(n6633), .ZN(n48794) );
  XOR2_X1 U38335 ( .A1(n17218), .A2(n38412), .Z(n17217) );
  XOR2_X1 U38336 ( .A1(n17845), .A2(n38414), .Z(n17219) );
  NOR2_X2 U38337 ( .A1(n40026), .A2(n23477), .ZN(n40025) );
  NAND2_X1 U38339 ( .A1(n17225), .A2(n53516), .ZN(n53467) );
  OAI21_X1 U38340 ( .A1(n53460), .A2(n17225), .B(n53507), .ZN(n53461) );
  XOR2_X1 U38341 ( .A1(n59585), .A2(n17227), .Z(n17226) );
  XOR2_X1 U38343 ( .A1(n17233), .A2(n51820), .Z(n51821) );
  XOR2_X1 U38346 ( .A1(n21348), .A2(n942), .Z(n17241) );
  NAND2_X2 U38349 ( .A1(n50360), .A2(n60975), .ZN(n49201) );
  NAND2_X2 U38350 ( .A1(n13370), .A2(n19555), .ZN(n20630) );
  NOR2_X1 U38355 ( .A1(n17255), .A2(n19373), .ZN(n35624) );
  NAND2_X1 U38356 ( .A1(n33319), .A2(n33550), .ZN(n17254) );
  NAND2_X2 U38361 ( .A1(n54102), .A2(n54110), .ZN(n54107) );
  NOR2_X1 U38363 ( .A1(n18178), .A2(n15703), .ZN(n55386) );
  XOR2_X1 U38364 ( .A1(n32616), .A2(n32611), .Z(n17271) );
  NAND2_X1 U38366 ( .A1(n6977), .A2(n9229), .ZN(n49133) );
  XOR2_X1 U38367 ( .A1(n19647), .A2(n18435), .Z(n50921) );
  XOR2_X1 U38368 ( .A1(n50325), .A2(n20306), .Z(n17273) );
  NAND2_X1 U38369 ( .A1(n17274), .A2(n29695), .ZN(n29696) );
  AOI22_X1 U38370 ( .A1(n27891), .A2(n17274), .B1(n29694), .B2(n20473), .ZN(
        n27893) );
  XNOR2_X1 U38371 ( .A1(n52510), .A2(n52435), .ZN(n17275) );
  XOR2_X1 U38372 ( .A1(n61462), .A2(n12591), .Z(n32095) );
  MUX2_X1 U38373 ( .I0(n32992), .I1(n32991), .S(n61090), .Z(n32998) );
  NOR2_X2 U38376 ( .A1(n27283), .A2(n14504), .ZN(n29179) );
  NAND2_X1 U38379 ( .A1(n17285), .A2(n29179), .ZN(n29182) );
  NOR2_X1 U38380 ( .A1(n1564), .A2(n17285), .ZN(n26816) );
  OAI21_X1 U38381 ( .A1(n26405), .A2(n1355), .B(n17285), .ZN(n26406) );
  INV_X2 U38382 ( .I(n17292), .ZN(n26034) );
  XNOR2_X1 U38383 ( .A1(Ciphertext[67]), .A2(Key[170]), .ZN(n17292) );
  XNOR2_X1 U38387 ( .A1(Ciphertext[94]), .A2(Key[71]), .ZN(n17311) );
  NOR2_X1 U38390 ( .A1(n59427), .A2(n40199), .ZN(n40205) );
  XOR2_X1 U38391 ( .A1(n17402), .A2(n33198), .Z(n33199) );
  XOR2_X1 U38392 ( .A1(n63050), .A2(n17403), .Z(n17402) );
  INV_X2 U38394 ( .I(n25654), .ZN(n20519) );
  XOR2_X1 U38395 ( .A1(n38781), .A2(n38957), .Z(n17321) );
  NAND2_X1 U38400 ( .A1(n52894), .A2(n52893), .ZN(n17329) );
  NAND2_X1 U38402 ( .A1(n20678), .A2(n17824), .ZN(n17333) );
  INV_X1 U38405 ( .I(n32513), .ZN(n24225) );
  AOI21_X1 U38408 ( .A1(n34126), .A2(n34125), .B(n62931), .ZN(n20909) );
  XOR2_X1 U38411 ( .A1(n17339), .A2(n39469), .Z(n38074) );
  XOR2_X1 U38412 ( .A1(n61045), .A2(n44759), .Z(n44470) );
  XOR2_X1 U38413 ( .A1(n61045), .A2(n56495), .Z(n52328) );
  XOR2_X1 U38414 ( .A1(n39539), .A2(n61045), .Z(n39540) );
  XOR2_X1 U38415 ( .A1(n37795), .A2(n61045), .Z(n31551) );
  XOR2_X1 U38417 ( .A1(n17344), .A2(n16035), .Z(n42284) );
  XOR2_X1 U38418 ( .A1(n17345), .A2(n38413), .Z(n17344) );
  XOR2_X1 U38419 ( .A1(n37568), .A2(n17346), .Z(n17345) );
  XOR2_X1 U38420 ( .A1(n37563), .A2(n38836), .Z(n38117) );
  NAND4_X2 U38421 ( .A1(n56831), .A2(n56832), .A3(n17348), .A4(n24177), .ZN(
        n25347) );
  NAND4_X1 U38423 ( .A1(n56833), .A2(n56832), .A3(n17348), .A4(n56831), .ZN(
        n56834) );
  INV_X1 U38426 ( .I(n40817), .ZN(n17351) );
  NAND2_X1 U38430 ( .A1(n17371), .A2(n62620), .ZN(n42189) );
  XOR2_X1 U38432 ( .A1(n39382), .A2(n39192), .Z(n17378) );
  XOR2_X1 U38434 ( .A1(n60889), .A2(n24234), .Z(n17383) );
  INV_X2 U38435 ( .I(n17384), .ZN(n54110) );
  AND2_X1 U38437 ( .A1(n41505), .A2(n41504), .Z(n17398) );
  XOR2_X1 U38439 ( .A1(n33074), .A2(n17402), .Z(n23451) );
  XOR2_X1 U38440 ( .A1(n39207), .A2(n17712), .Z(n17405) );
  XOR2_X1 U38442 ( .A1(n19410), .A2(n11751), .Z(n17406) );
  NOR2_X2 U38443 ( .A1(n26935), .A2(n27233), .ZN(n27538) );
  OAI22_X1 U38444 ( .A1(n23474), .A2(n27232), .B1(n27537), .B2(n64994), .ZN(
        n27234) );
  NAND2_X2 U38445 ( .A1(n1793), .A2(n17407), .ZN(n35482) );
  NOR3_X2 U38450 ( .A1(n18760), .A2(n18758), .A3(n18759), .ZN(n30953) );
  NAND2_X2 U38451 ( .A1(n17416), .A2(n26056), .ZN(n29862) );
  NAND2_X1 U38455 ( .A1(n34589), .A2(n59522), .ZN(n33968) );
  AOI22_X1 U38458 ( .A1(n61917), .A2(n17420), .B1(n64234), .B2(n34583), .ZN(
        n34593) );
  NAND2_X2 U38460 ( .A1(n27621), .A2(n20721), .ZN(n18747) );
  NAND2_X1 U38463 ( .A1(n22239), .A2(n17423), .ZN(n45579) );
  INV_X1 U38464 ( .I(n15360), .ZN(n17423) );
  INV_X1 U38465 ( .I(n17429), .ZN(n17428) );
  NOR4_X1 U38466 ( .A1(n21800), .A2(n22716), .A3(n17429), .A4(n43309), .ZN(
        n20323) );
  NAND2_X2 U38467 ( .A1(n44226), .A2(n43995), .ZN(n17429) );
  XOR2_X1 U38468 ( .A1(n17431), .A2(n17430), .Z(Plaintext[60]) );
  XOR2_X1 U38470 ( .A1(n17439), .A2(n16208), .Z(n51632) );
  NAND3_X1 U38475 ( .A1(n37188), .A2(n37187), .A3(n17444), .ZN(n37192) );
  NOR2_X1 U38476 ( .A1(n37003), .A2(n17444), .ZN(n37004) );
  NAND2_X2 U38479 ( .A1(n25022), .A2(n56942), .ZN(n56964) );
  XOR2_X1 U38482 ( .A1(n38942), .A2(n38634), .Z(n17447) );
  XOR2_X1 U38485 ( .A1(n11239), .A2(n65079), .Z(n39653) );
  INV_X1 U38486 ( .I(n37563), .ZN(n37511) );
  XOR2_X1 U38487 ( .A1(n17463), .A2(n32723), .Z(n32724) );
  XOR2_X1 U38489 ( .A1(n43942), .A2(n44247), .Z(n17466) );
  NAND2_X1 U38490 ( .A1(n23349), .A2(n30679), .ZN(n30245) );
  XOR2_X1 U38494 ( .A1(n25816), .A2(n62241), .Z(n17476) );
  AOI21_X1 U38498 ( .A1(n18200), .A2(n27292), .B(n17489), .ZN(n26713) );
  AOI21_X1 U38501 ( .A1(n18075), .A2(n13943), .B(n17495), .ZN(n19940) );
  XOR2_X1 U38502 ( .A1(n26022), .A2(n50947), .Z(n17497) );
  NOR2_X2 U38504 ( .A1(n29371), .A2(n29370), .ZN(n17522) );
  NAND2_X2 U38505 ( .A1(n55639), .A2(n55627), .ZN(n17500) );
  NAND3_X2 U38506 ( .A1(n41732), .A2(n41733), .A3(n17501), .ZN(n42834) );
  NAND2_X1 U38508 ( .A1(n12338), .A2(n34669), .ZN(n34055) );
  XOR2_X1 U38509 ( .A1(n62985), .A2(n24040), .Z(n17504) );
  NAND3_X1 U38510 ( .A1(n47407), .A2(n18227), .A3(n47669), .ZN(n45906) );
  NAND3_X1 U38511 ( .A1(n30758), .A2(n30757), .A3(n30760), .ZN(n17508) );
  XOR2_X1 U38512 ( .A1(n31432), .A2(n17509), .Z(n17511) );
  XOR2_X1 U38513 ( .A1(n17510), .A2(n30798), .Z(n17509) );
  INV_X2 U38514 ( .I(n25668), .ZN(n30895) );
  XOR2_X1 U38515 ( .A1(n17511), .A2(n16045), .Z(n25668) );
  XOR2_X1 U38516 ( .A1(n19828), .A2(n31668), .Z(n31750) );
  NAND2_X2 U38517 ( .A1(n18886), .A2(n1326), .ZN(n18750) );
  XOR2_X1 U38520 ( .A1(n18891), .A2(n51490), .Z(n51737) );
  XOR2_X1 U38521 ( .A1(n17521), .A2(n17520), .Z(n21653) );
  INV_X2 U38522 ( .I(n25129), .ZN(n29371) );
  INV_X1 U38523 ( .I(n19940), .ZN(n17526) );
  INV_X2 U38524 ( .I(n30125), .ZN(n24987) );
  NAND3_X2 U38525 ( .A1(n17529), .A2(n17528), .A3(n17527), .ZN(n30125) );
  NOR2_X1 U38526 ( .A1(n48122), .A2(n17530), .ZN(n17900) );
  NAND2_X1 U38531 ( .A1(n10353), .A2(n48341), .ZN(n25810) );
  NAND2_X1 U38532 ( .A1(n49902), .A2(n63186), .ZN(n25813) );
  OR2_X1 U38539 ( .A1(n40758), .A2(n40759), .Z(n17557) );
  AND2_X1 U38540 ( .A1(n49364), .A2(n3348), .Z(n17558) );
  NOR3_X1 U38541 ( .A1(n15834), .A2(n43502), .A3(n17560), .ZN(n17559) );
  NAND2_X2 U38542 ( .A1(n19000), .A2(n61442), .ZN(n43506) );
  NAND2_X1 U38543 ( .A1(n17573), .A2(n57728), .ZN(n46715) );
  NAND2_X1 U38544 ( .A1(n17573), .A2(n64605), .ZN(n47193) );
  XOR2_X1 U38548 ( .A1(n17584), .A2(n44434), .Z(n18357) );
  OR2_X2 U38553 ( .A1(n27844), .A2(n27845), .Z(n22444) );
  XOR2_X1 U38557 ( .A1(n24479), .A2(n23197), .Z(n24848) );
  XOR2_X1 U38558 ( .A1(n17598), .A2(n50920), .Z(n17599) );
  INV_X2 U38560 ( .I(n20326), .ZN(n21056) );
  AOI21_X2 U38563 ( .A1(n17602), .A2(n26833), .B(n26832), .ZN(n24993) );
  AOI21_X1 U38564 ( .A1(n56194), .A2(n17606), .B(n23258), .ZN(n56195) );
  XOR2_X1 U38565 ( .A1(n58440), .A2(n10378), .Z(n17608) );
  NOR2_X2 U38566 ( .A1(n41052), .A2(n41874), .ZN(n41885) );
  NAND2_X1 U38568 ( .A1(n45200), .A2(n17610), .ZN(n17613) );
  OAI21_X1 U38569 ( .A1(n10734), .A2(n12051), .B(n10427), .ZN(n28206) );
  NOR2_X1 U38570 ( .A1(n20747), .A2(n12051), .ZN(n29491) );
  NOR2_X1 U38571 ( .A1(n31118), .A2(n65), .ZN(n31120) );
  XOR2_X1 U38572 ( .A1(n32638), .A2(n32064), .Z(n21661) );
  XOR2_X1 U38573 ( .A1(n17617), .A2(n17616), .Z(n32064) );
  NAND2_X2 U38574 ( .A1(n41052), .A2(n41874), .ZN(n19466) );
  AOI22_X1 U38576 ( .A1(n29366), .A2(n27435), .B1(n17619), .B2(n27436), .ZN(
        n27440) );
  NOR2_X1 U38579 ( .A1(n30168), .A2(n60111), .ZN(n17628) );
  NAND2_X2 U38580 ( .A1(n39994), .A2(n41383), .ZN(n41376) );
  XOR2_X1 U38585 ( .A1(n26942), .A2(Key[107]), .Z(n29282) );
  NAND2_X2 U38587 ( .A1(n23578), .A2(n18062), .ZN(n29284) );
  NAND2_X1 U38589 ( .A1(n53044), .A2(n53809), .ZN(n17637) );
  NOR2_X1 U38590 ( .A1(n17642), .A2(n17639), .ZN(n17638) );
  OAI21_X1 U38591 ( .A1(n24535), .A2(n17644), .B(n17643), .ZN(n17642) );
  NAND3_X1 U38592 ( .A1(n53044), .A2(n53809), .A3(n53046), .ZN(n17643) );
  NAND2_X1 U38593 ( .A1(n19692), .A2(n19694), .ZN(n17644) );
  NAND2_X1 U38594 ( .A1(n56887), .A2(n56848), .ZN(n17645) );
  MUX2_X1 U38595 ( .I0(n17648), .I1(n17647), .S(n56885), .Z(n17646) );
  OAI22_X2 U38598 ( .A1(n56840), .A2(n56872), .B1(n56846), .B2(n23074), .ZN(
        n17655) );
  XOR2_X1 U38601 ( .A1(n45402), .A2(n43775), .Z(n17656) );
  XOR2_X1 U38602 ( .A1(n16691), .A2(n16325), .Z(n51189) );
  NAND2_X1 U38605 ( .A1(n36010), .A2(n61747), .ZN(n17667) );
  NOR2_X1 U38607 ( .A1(n17364), .A2(n1417), .ZN(n35067) );
  NAND2_X2 U38609 ( .A1(n34083), .A2(n34627), .ZN(n24737) );
  XOR2_X1 U38611 ( .A1(n11448), .A2(n52446), .Z(n21340) );
  NAND2_X1 U38612 ( .A1(n17672), .A2(n17683), .ZN(n17679) );
  NAND4_X2 U38613 ( .A1(n17681), .A2(n45793), .A3(n17680), .A4(n17679), .ZN(
        n17678) );
  INV_X2 U38615 ( .I(n43778), .ZN(n43925) );
  XOR2_X1 U38616 ( .A1(n43924), .A2(n43778), .Z(n42064) );
  AOI21_X1 U38617 ( .A1(n17945), .A2(n42480), .B(n42479), .ZN(n41839) );
  XOR2_X1 U38618 ( .A1(n44728), .A2(n17702), .Z(n17701) );
  OAI21_X1 U38619 ( .A1(n49594), .A2(n17874), .B(n49593), .ZN(n49595) );
  XOR2_X1 U38620 ( .A1(n17704), .A2(n51976), .Z(n55672) );
  XOR2_X1 U38621 ( .A1(n51763), .A2(n50941), .Z(n17705) );
  NAND2_X1 U38622 ( .A1(n17708), .A2(n1260), .ZN(n52008) );
  NAND2_X1 U38623 ( .A1(n17708), .A2(n55668), .ZN(n25336) );
  OAI21_X1 U38624 ( .A1(n55447), .A2(n55670), .B(n17708), .ZN(n55450) );
  XOR2_X1 U38626 ( .A1(n39234), .A2(n37267), .Z(n17711) );
  NAND2_X1 U38627 ( .A1(n1263), .A2(n47414), .ZN(n47417) );
  NAND2_X2 U38628 ( .A1(n11084), .A2(n11279), .ZN(n24633) );
  XOR2_X1 U38633 ( .A1(n44050), .A2(n44051), .Z(n17733) );
  XOR2_X1 U38634 ( .A1(n15810), .A2(n17735), .Z(n17736) );
  XOR2_X1 U38635 ( .A1(n17736), .A2(n44059), .Z(n44060) );
  NAND2_X2 U38640 ( .A1(n28630), .A2(n27691), .ZN(n19287) );
  NAND2_X2 U38641 ( .A1(n28633), .A2(n27823), .ZN(n20627) );
  NOR2_X1 U38642 ( .A1(n17745), .A2(n30767), .ZN(n29546) );
  XOR2_X1 U38643 ( .A1(n30767), .A2(n17745), .Z(n29956) );
  INV_X4 U38645 ( .I(n24335), .ZN(n17745) );
  INV_X2 U38646 ( .I(n19196), .ZN(n26720) );
  OAI21_X1 U38649 ( .A1(n35383), .A2(n36063), .B(n60196), .ZN(n36895) );
  XOR2_X1 U38654 ( .A1(n52589), .A2(n51960), .Z(n17756) );
  XOR2_X1 U38655 ( .A1(n52086), .A2(n15719), .Z(n17757) );
  NAND2_X1 U38657 ( .A1(n17759), .A2(n34155), .ZN(n33358) );
  NAND3_X1 U38658 ( .A1(n34156), .A2(n23351), .A3(n17759), .ZN(n32850) );
  NAND2_X1 U38661 ( .A1(n58424), .A2(n29521), .ZN(n29100) );
  NAND2_X2 U38662 ( .A1(n17778), .A2(n17780), .ZN(n26650) );
  NAND2_X2 U38664 ( .A1(n14705), .A2(n23942), .ZN(n27121) );
  XOR2_X1 U38665 ( .A1(n17764), .A2(n31750), .Z(n17763) );
  XOR2_X1 U38667 ( .A1(n23181), .A2(n37515), .Z(n17772) );
  XOR2_X1 U38668 ( .A1(n64241), .A2(n17583), .Z(n39300) );
  INV_X2 U38669 ( .I(n20892), .ZN(n19307) );
  XOR2_X1 U38670 ( .A1(n25843), .A2(n18696), .Z(n17777) );
  INV_X1 U38672 ( .I(n17794), .ZN(n26371) );
  XOR2_X1 U38675 ( .A1(n51503), .A2(n51501), .Z(n17802) );
  NAND2_X1 U38676 ( .A1(n49493), .A2(n49486), .ZN(n48854) );
  XOR2_X1 U38680 ( .A1(n18832), .A2(n17817), .Z(n37578) );
  OAI21_X1 U38683 ( .A1(n3031), .A2(n50373), .B(n17818), .ZN(n50381) );
  XOR2_X1 U38685 ( .A1(n37082), .A2(n38578), .Z(n37099) );
  NOR2_X2 U38687 ( .A1(n56565), .A2(n51268), .ZN(n18323) );
  INV_X1 U38689 ( .I(n31702), .ZN(n33162) );
  NOR2_X1 U38690 ( .A1(n17824), .A2(n28811), .ZN(n27437) );
  NOR2_X1 U38691 ( .A1(n27328), .A2(n17824), .ZN(n26457) );
  AOI22_X1 U38692 ( .A1(n27330), .A2(n29367), .B1(n17824), .B2(n28801), .ZN(
        n27331) );
  NAND3_X1 U38696 ( .A1(n19968), .A2(n55295), .A3(n51964), .ZN(n17837) );
  AOI21_X1 U38698 ( .A1(n48529), .A2(n22255), .B(n17840), .ZN(n25266) );
  XOR2_X1 U38699 ( .A1(n17841), .A2(n22773), .Z(Plaintext[135]) );
  XOR2_X1 U38700 ( .A1(n17347), .A2(n22698), .Z(n38414) );
  XOR2_X1 U38701 ( .A1(n38411), .A2(n38410), .Z(n17846) );
  XOR2_X1 U38702 ( .A1(n33138), .A2(n33137), .Z(n17847) );
  NAND4_X2 U38705 ( .A1(n39078), .A2(n15913), .A3(n24765), .A4(n39079), .ZN(
        n23364) );
  INV_X1 U38708 ( .I(n491), .ZN(n20097) );
  XOR2_X1 U38711 ( .A1(Ciphertext[164]), .A2(Key[177]), .Z(n28806) );
  NAND2_X1 U38712 ( .A1(n21828), .A2(n58277), .ZN(n17861) );
  NOR2_X1 U38713 ( .A1(n17862), .A2(n57116), .ZN(n18804) );
  NOR2_X1 U38714 ( .A1(n17862), .A2(n57233), .ZN(n21440) );
  XOR2_X1 U38717 ( .A1(n17863), .A2(n47769), .Z(n51813) );
  AOI22_X1 U38721 ( .A1(n30697), .A2(n30696), .B1(n60187), .B2(n60142), .ZN(
        n30698) );
  XOR2_X1 U38722 ( .A1(n16299), .A2(n32170), .Z(n17875) );
  NAND2_X2 U38724 ( .A1(n17880), .A2(n17876), .ZN(n31242) );
  NAND3_X1 U38726 ( .A1(n49935), .A2(n21870), .A3(n49936), .ZN(n17883) );
  NAND3_X1 U38728 ( .A1(n50333), .A2(n50336), .A3(n7098), .ZN(n17884) );
  NAND3_X2 U38732 ( .A1(n47130), .A2(n47129), .A3(n47131), .ZN(n50236) );
  INV_X2 U38733 ( .I(n51407), .ZN(n52470) );
  XOR2_X1 U38734 ( .A1(n30402), .A2(n8279), .Z(n39650) );
  XOR2_X1 U38736 ( .A1(n17890), .A2(n37892), .Z(n17889) );
  XOR2_X1 U38737 ( .A1(n38117), .A2(n37893), .Z(n17890) );
  NOR2_X1 U38740 ( .A1(n21932), .A2(n15020), .ZN(n21933) );
  NOR4_X2 U38741 ( .A1(n28295), .A2(n28294), .A3(n28293), .A4(n28705), .ZN(
        n28297) );
  NAND4_X1 U38748 ( .A1(n54601), .A2(n23897), .A3(n64129), .A4(n54597), .ZN(
        n54326) );
  NOR2_X1 U38751 ( .A1(n42836), .A2(n65185), .ZN(n25709) );
  NOR2_X2 U38752 ( .A1(n16103), .A2(n42836), .ZN(n42148) );
  INV_X1 U38754 ( .I(n35950), .ZN(n34920) );
  NAND4_X1 U38756 ( .A1(n22945), .A2(n28831), .A3(n28136), .A4(n22720), .ZN(
        n28140) );
  NOR3_X1 U38759 ( .A1(n4436), .A2(n49274), .A3(n64488), .ZN(n25559) );
  OAI21_X1 U38760 ( .A1(n56167), .A2(n56191), .B(n56196), .ZN(n19944) );
  OAI21_X1 U38762 ( .A1(n32457), .A2(n33406), .B(n32782), .ZN(n32453) );
  NAND2_X1 U38764 ( .A1(n20508), .A2(n27483), .ZN(n27231) );
  NAND2_X1 U38765 ( .A1(n56170), .A2(n56169), .ZN(n19942) );
  NAND2_X1 U38767 ( .A1(n36342), .A2(n35863), .ZN(n24722) );
  NOR2_X1 U38768 ( .A1(n36338), .A2(n36340), .ZN(n36345) );
  OAI21_X1 U38771 ( .A1(n33625), .A2(n33626), .B(n33624), .ZN(n20769) );
  NAND2_X1 U38772 ( .A1(n33624), .A2(n33627), .ZN(n18243) );
  NAND2_X1 U38773 ( .A1(n24093), .A2(n33540), .ZN(n33220) );
  NAND2_X2 U38774 ( .A1(n43839), .A2(n57591), .ZN(n43851) );
  OAI21_X1 U38776 ( .A1(n18249), .A2(n1383), .B(n50220), .ZN(n18250) );
  INV_X1 U38777 ( .I(n38070), .ZN(n22451) );
  NAND3_X1 U38779 ( .A1(n56175), .A2(n56176), .A3(n15872), .ZN(n18601) );
  NOR3_X1 U38780 ( .A1(n56185), .A2(n56191), .A3(n56146), .ZN(n56147) );
  OAI22_X1 U38782 ( .A1(n19045), .A2(n64732), .B1(n41064), .B2(n40588), .ZN(
        n40589) );
  NOR2_X1 U38784 ( .A1(n39795), .A2(n64732), .ZN(n37825) );
  BUF_X2 U38785 ( .I(n38992), .Z(n18054) );
  AOI22_X1 U38786 ( .A1(n25184), .A2(n30230), .B1(n30681), .B2(n30237), .ZN(
        n25183) );
  NOR2_X1 U38787 ( .A1(n30239), .A2(n30230), .ZN(n19266) );
  INV_X1 U38788 ( .I(n44820), .ZN(n18139) );
  NAND2_X1 U38790 ( .A1(n8640), .A2(n11092), .ZN(n30638) );
  NAND2_X1 U38793 ( .A1(n19023), .A2(n19022), .ZN(n55652) );
  NAND2_X1 U38794 ( .A1(n19021), .A2(n21099), .ZN(n55626) );
  BUF_X4 U38795 ( .I(n21099), .Z(n19020) );
  NAND2_X1 U38796 ( .A1(n28383), .A2(n27111), .ZN(n26549) );
  NAND3_X1 U38797 ( .A1(n1790), .A2(n1217), .A3(n2362), .ZN(n34096) );
  AOI21_X1 U38799 ( .A1(n56511), .A2(n56512), .B(n17893), .ZN(n56513) );
  NOR2_X2 U38802 ( .A1(n1543), .A2(n35026), .ZN(n34026) );
  NOR2_X1 U38803 ( .A1(n34558), .A2(n64954), .ZN(n17897) );
  NAND2_X1 U38804 ( .A1(n17906), .A2(n49685), .ZN(n47642) );
  NAND3_X1 U38805 ( .A1(n17906), .A2(n58645), .A3(n16922), .ZN(n49368) );
  NOR3_X2 U38808 ( .A1(n34062), .A2(n34063), .A3(n34064), .ZN(n36746) );
  XOR2_X1 U38809 ( .A1(n19204), .A2(n17914), .Z(n31805) );
  XOR2_X1 U38810 ( .A1(n17463), .A2(n17914), .Z(n32313) );
  NAND2_X1 U38811 ( .A1(n17915), .A2(n61233), .ZN(n17916) );
  NAND2_X1 U38812 ( .A1(n1730), .A2(n39509), .ZN(n17917) );
  XOR2_X1 U38814 ( .A1(n20441), .A2(n17921), .Z(n17920) );
  XOR2_X1 U38815 ( .A1(n17922), .A2(n34613), .Z(n33421) );
  NAND2_X1 U38816 ( .A1(n34616), .A2(n60763), .ZN(n31025) );
  NAND3_X2 U38818 ( .A1(n21278), .A2(n33983), .A3(n33986), .ZN(n26147) );
  INV_X1 U38819 ( .I(n17928), .ZN(n22886) );
  XOR2_X1 U38822 ( .A1(n33883), .A2(n1830), .Z(n17932) );
  XOR2_X1 U38823 ( .A1(n31753), .A2(n22390), .Z(n17934) );
  XOR2_X1 U38824 ( .A1(n20308), .A2(n56692), .Z(n33883) );
  INV_X2 U38825 ( .I(n18230), .ZN(n24009) );
  XOR2_X1 U38827 ( .A1(n17942), .A2(n50921), .Z(n26228) );
  XOR2_X1 U38828 ( .A1(n15722), .A2(n51368), .Z(n17943) );
  NAND2_X1 U38830 ( .A1(n60843), .A2(n8305), .ZN(n17949) );
  AND3_X1 U38831 ( .A1(n50285), .A2(n1384), .A3(n57182), .Z(n17954) );
  OR2_X2 U38832 ( .A1(n34342), .A2(n34336), .Z(n22278) );
  OAI21_X1 U38833 ( .A1(n15937), .A2(n17959), .B(n54915), .ZN(n54894) );
  AOI22_X1 U38834 ( .A1(n54879), .A2(n15937), .B1(n17959), .B2(n54912), .ZN(
        n54886) );
  NAND2_X1 U38836 ( .A1(n41556), .A2(n17963), .ZN(n17962) );
  NAND2_X1 U38839 ( .A1(n17971), .A2(n38601), .ZN(n38603) );
  NAND2_X2 U38841 ( .A1(n29625), .A2(n20714), .ZN(n17972) );
  XOR2_X1 U38846 ( .A1(n17980), .A2(n38374), .Z(n38376) );
  XOR2_X1 U38847 ( .A1(n39455), .A2(n17980), .Z(n37576) );
  NAND2_X1 U38849 ( .A1(n62358), .A2(n22526), .ZN(n49160) );
  AOI21_X1 U38850 ( .A1(n62358), .A2(n16595), .B(n57610), .ZN(n49749) );
  NAND3_X1 U38851 ( .A1(n42280), .A2(n42281), .A3(n21493), .ZN(n40812) );
  NAND3_X1 U38853 ( .A1(n7571), .A2(n41248), .A3(n59019), .ZN(n37598) );
  XOR2_X1 U38854 ( .A1(n17983), .A2(n44300), .Z(n44301) );
  XOR2_X1 U38855 ( .A1(n17983), .A2(n44447), .Z(n44448) );
  XOR2_X1 U38856 ( .A1(n17983), .A2(n43938), .Z(n43939) );
  XOR2_X1 U38857 ( .A1(n17983), .A2(n43401), .Z(n43402) );
  XOR2_X1 U38858 ( .A1(n22207), .A2(n17983), .Z(n43640) );
  XOR2_X1 U38859 ( .A1(n24017), .A2(n785), .Z(n17985) );
  XOR2_X1 U38860 ( .A1(n5009), .A2(n60528), .Z(n17986) );
  OAI21_X1 U38861 ( .A1(n31716), .A2(n31715), .B(n61646), .ZN(n25819) );
  AOI21_X1 U38863 ( .A1(n29621), .A2(n22945), .B(n29627), .ZN(n17988) );
  NOR2_X2 U38865 ( .A1(n19290), .A2(n28119), .ZN(n17989) );
  XOR2_X1 U38866 ( .A1(n26951), .A2(n26952), .Z(n29629) );
  NAND3_X1 U38868 ( .A1(n49195), .A2(n48847), .A3(n13038), .ZN(n48841) );
  INV_X2 U38869 ( .I(n25713), .ZN(n23853) );
  XOR2_X1 U38870 ( .A1(n39232), .A2(n39261), .Z(n17999) );
  XOR2_X1 U38871 ( .A1(n39337), .A2(n19381), .Z(n39232) );
  AND2_X1 U38872 ( .A1(n45192), .A2(n47905), .Z(n18000) );
  XNOR2_X1 U38874 ( .A1(Ciphertext[45]), .A2(Key[16]), .ZN(n18004) );
  AOI21_X1 U38877 ( .A1(n28484), .A2(n28485), .B(n18006), .ZN(n19369) );
  AND2_X1 U38879 ( .A1(n20599), .A2(n56361), .Z(n18010) );
  XOR2_X1 U38880 ( .A1(n46520), .A2(n16323), .Z(n18011) );
  XOR2_X1 U38881 ( .A1(n27796), .A2(n18014), .Z(n18013) );
  XOR2_X1 U38882 ( .A1(n24858), .A2(n30992), .Z(n18014) );
  AOI21_X1 U38885 ( .A1(n36185), .A2(n36403), .B(n4263), .ZN(n36186) );
  NAND3_X1 U38886 ( .A1(n18029), .A2(n18027), .A3(n25929), .ZN(n18603) );
  INV_X2 U38891 ( .I(n18039), .ZN(n44802) );
  XOR2_X1 U38893 ( .A1(n18050), .A2(n7713), .Z(n37763) );
  XOR2_X1 U38894 ( .A1(n18049), .A2(n21098), .Z(n18050) );
  XOR2_X1 U38896 ( .A1(n15932), .A2(n37785), .Z(n39468) );
  XOR2_X1 U38899 ( .A1(n2036), .A2(n18058), .Z(n24173) );
  XOR2_X1 U38900 ( .A1(n18887), .A2(n16319), .Z(n18058) );
  NOR2_X2 U38901 ( .A1(n30799), .A2(n29835), .ZN(n30815) );
  NAND2_X2 U38905 ( .A1(n17632), .A2(n18062), .ZN(n20034) );
  NOR2_X2 U38906 ( .A1(n17632), .A2(n18062), .ZN(n20714) );
  NOR2_X1 U38907 ( .A1(n28125), .A2(n18062), .ZN(n28833) );
  NOR2_X1 U38908 ( .A1(n29291), .A2(n18062), .ZN(n28142) );
  XOR2_X1 U38913 ( .A1(n44744), .A2(n18067), .Z(n18066) );
  XOR2_X1 U38918 ( .A1(n18073), .A2(n37608), .Z(n37609) );
  NAND3_X2 U38920 ( .A1(n26817), .A2(n23598), .A3(n26818), .ZN(n23024) );
  AOI21_X1 U38921 ( .A1(n20660), .A2(n18077), .B(n34950), .ZN(n34951) );
  NOR2_X2 U38923 ( .A1(n40706), .A2(n40705), .ZN(n18087) );
  AND3_X1 U38925 ( .A1(n51559), .A2(n56360), .A3(n51558), .Z(n18097) );
  NAND3_X1 U38929 ( .A1(n18104), .A2(n41640), .A3(n41646), .ZN(n41644) );
  OAI21_X1 U38930 ( .A1(n41648), .A2(n41649), .B(n18104), .ZN(n41650) );
  NOR2_X2 U38932 ( .A1(n55494), .A2(n20849), .ZN(n55685) );
  XOR2_X1 U38936 ( .A1(n3665), .A2(n23518), .Z(n18122) );
  XOR2_X1 U38938 ( .A1(n6967), .A2(n44130), .Z(n20668) );
  OR2_X2 U38939 ( .A1(n52719), .A2(n56210), .Z(n56417) );
  XOR2_X1 U38940 ( .A1(n51478), .A2(n51054), .Z(n18125) );
  INV_X1 U38941 ( .I(n10088), .ZN(n47609) );
  NAND2_X1 U38942 ( .A1(n43309), .A2(n19346), .ZN(n42956) );
  NAND2_X2 U38943 ( .A1(n43995), .A2(n22716), .ZN(n19346) );
  NAND2_X2 U38944 ( .A1(n1782), .A2(n22527), .ZN(n18130) );
  NAND2_X2 U38946 ( .A1(n30418), .A2(n22971), .ZN(n19048) );
  NAND2_X1 U38947 ( .A1(n18134), .A2(n55378), .ZN(n55380) );
  NAND3_X2 U38955 ( .A1(n20485), .A2(n20486), .A3(n16086), .ZN(n18582) );
  NAND3_X1 U38959 ( .A1(n36848), .A2(n36850), .A3(n61747), .ZN(n18150) );
  NOR2_X2 U38960 ( .A1(n41384), .A2(n39994), .ZN(n41118) );
  XOR2_X1 U38961 ( .A1(n39238), .A2(n39239), .Z(n39240) );
  XOR2_X1 U38962 ( .A1(n39232), .A2(n39238), .Z(n18656) );
  INV_X2 U38967 ( .I(n18167), .ZN(n34606) );
  XOR2_X1 U38969 ( .A1(n39227), .A2(n57448), .Z(n18169) );
  XOR2_X1 U38970 ( .A1(n63032), .A2(n15955), .Z(n18170) );
  NAND2_X1 U38971 ( .A1(n55377), .A2(n18178), .ZN(n18283) );
  XOR2_X1 U38972 ( .A1(n57194), .A2(n19107), .Z(n18183) );
  INV_X2 U38973 ( .I(n26047), .ZN(n51763) );
  XOR2_X1 U38975 ( .A1(n18189), .A2(n51203), .Z(n18187) );
  XOR2_X1 U38976 ( .A1(n18188), .A2(n49188), .Z(n51203) );
  XOR2_X1 U38977 ( .A1(n52201), .A2(n9635), .Z(n18188) );
  NOR2_X1 U38978 ( .A1(n53391), .A2(n18193), .ZN(n50206) );
  NOR2_X1 U38979 ( .A1(n11119), .A2(n18195), .ZN(n56570) );
  AOI21_X1 U38980 ( .A1(n64295), .A2(n55934), .B(n18195), .ZN(n55935) );
  AOI21_X1 U38981 ( .A1(n51265), .A2(n10183), .B(n18195), .ZN(n51252) );
  NOR2_X1 U38982 ( .A1(n56389), .A2(n51268), .ZN(n18194) );
  NOR2_X1 U38984 ( .A1(n18199), .A2(n35817), .ZN(n19772) );
  INV_X1 U38985 ( .I(n18202), .ZN(n48810) );
  NAND2_X1 U38987 ( .A1(n18203), .A2(n28539), .ZN(n27251) );
  OAI21_X1 U38988 ( .A1(n27868), .A2(n18203), .B(n26753), .ZN(n26754) );
  NOR2_X1 U38989 ( .A1(n28527), .A2(n18203), .ZN(n28528) );
  AOI21_X1 U38990 ( .A1(n26757), .A2(n18203), .B(n26798), .ZN(n26758) );
  INV_X2 U38991 ( .I(n34203), .ZN(n21584) );
  INV_X1 U38993 ( .I(n18213), .ZN(n28434) );
  NOR2_X1 U38994 ( .A1(n28460), .A2(n65039), .ZN(n28461) );
  OR2_X1 U38997 ( .A1(n34395), .A2(n24089), .Z(n18218) );
  NOR2_X2 U38998 ( .A1(n52044), .A2(n55299), .ZN(n55684) );
  XOR2_X1 U38999 ( .A1(n18222), .A2(n51937), .Z(n50953) );
  INV_X2 U39000 ( .I(n24577), .ZN(n55017) );
  OAI21_X1 U39001 ( .A1(n28033), .A2(n21301), .B(n18223), .ZN(n28029) );
  NAND2_X1 U39002 ( .A1(n61643), .A2(n28033), .ZN(n18223) );
  NOR2_X2 U39006 ( .A1(n18247), .A2(n24009), .ZN(n55016) );
  NAND2_X1 U39008 ( .A1(n30230), .A2(n10431), .ZN(n18234) );
  NOR2_X1 U39013 ( .A1(n18242), .A2(n24633), .ZN(n40035) );
  NAND2_X1 U39014 ( .A1(n54330), .A2(n54331), .ZN(n18246) );
  NAND2_X1 U39016 ( .A1(n17935), .A2(n18247), .ZN(n54452) );
  XOR2_X1 U39017 ( .A1(n18248), .A2(n30911), .Z(n30912) );
  XOR2_X1 U39018 ( .A1(n65112), .A2(n32617), .Z(n32193) );
  XOR2_X1 U39019 ( .A1(n65112), .A2(n22476), .Z(n32399) );
  XOR2_X1 U39020 ( .A1(n65112), .A2(n31980), .Z(n31981) );
  NOR2_X1 U39021 ( .A1(n20971), .A2(n62248), .ZN(n48009) );
  AOI22_X1 U39022 ( .A1(n48712), .A2(n62248), .B1(n49677), .B2(n49675), .ZN(
        n48713) );
  XOR2_X1 U39024 ( .A1(n18259), .A2(n18262), .Z(n20962) );
  XOR2_X1 U39025 ( .A1(n18261), .A2(n18260), .Z(n18259) );
  XOR2_X1 U39026 ( .A1(n51229), .A2(n51227), .Z(n18261) );
  XOR2_X1 U39027 ( .A1(n52360), .A2(n51628), .Z(n51227) );
  XOR2_X1 U39028 ( .A1(n51224), .A2(n51228), .Z(n18262) );
  XOR2_X1 U39029 ( .A1(n13325), .A2(n7459), .Z(n51228) );
  INV_X1 U39031 ( .I(n19331), .ZN(n40350) );
  XNOR2_X1 U39032 ( .A1(n466), .A2(n11829), .ZN(n18268) );
  NAND2_X1 U39033 ( .A1(n61697), .A2(n11716), .ZN(n56159) );
  NAND4_X1 U39035 ( .A1(n9424), .A2(n24063), .A3(n55362), .A4(n58828), .ZN(
        n18287) );
  NAND2_X1 U39036 ( .A1(n55384), .A2(n9424), .ZN(n55338) );
  NOR2_X1 U39037 ( .A1(n18109), .A2(n55690), .ZN(n18291) );
  NOR2_X1 U39038 ( .A1(n65283), .A2(n18294), .ZN(n55689) );
  NOR2_X1 U39039 ( .A1(n18109), .A2(n18293), .ZN(n18292) );
  NOR2_X1 U39040 ( .A1(n55694), .A2(n18294), .ZN(n55699) );
  XOR2_X1 U39041 ( .A1(n18296), .A2(n22806), .Z(n31935) );
  XOR2_X1 U39042 ( .A1(n10622), .A2(n15733), .Z(n31234) );
  NAND2_X2 U39043 ( .A1(n15871), .A2(n21792), .ZN(n47262) );
  NAND2_X1 U39045 ( .A1(n7501), .A2(n64390), .ZN(n41135) );
  XOR2_X1 U39046 ( .A1(n18303), .A2(n18302), .Z(n23781) );
  XOR2_X1 U39047 ( .A1(n25164), .A2(n32171), .Z(n18303) );
  OAI22_X1 U39048 ( .A1(n33330), .A2(n36589), .B1(n36163), .B2(n34378), .ZN(
        n18305) );
  NOR2_X1 U39050 ( .A1(n9346), .A2(n7086), .ZN(n48958) );
  NOR2_X1 U39052 ( .A1(n18313), .A2(n35361), .ZN(n36119) );
  NOR3_X1 U39053 ( .A1(n18313), .A2(n36193), .A3(n10601), .ZN(n35124) );
  NOR2_X1 U39055 ( .A1(n18602), .A2(n18313), .ZN(n19139) );
  XOR2_X1 U39058 ( .A1(n18316), .A2(n18334), .Z(n18315) );
  INV_X2 U39060 ( .I(n18317), .ZN(n23410) );
  INV_X2 U39063 ( .I(n26081), .ZN(n32654) );
  NAND2_X1 U39064 ( .A1(n18323), .A2(n56573), .ZN(n56279) );
  XOR2_X1 U39068 ( .A1(n39582), .A2(n37823), .Z(n18334) );
  XOR2_X1 U39072 ( .A1(n5779), .A2(n37888), .Z(n37611) );
  XOR2_X1 U39073 ( .A1(n39391), .A2(n56692), .Z(n18340) );
  NAND3_X1 U39075 ( .A1(n46907), .A2(n59892), .A3(n18361), .ZN(n45769) );
  XOR2_X1 U39077 ( .A1(n24112), .A2(n44168), .Z(n18362) );
  OAI21_X1 U39079 ( .A1(n55878), .A2(n60203), .B(n18376), .ZN(n19951) );
  OAI22_X1 U39080 ( .A1(n18561), .A2(n18560), .B1(n55894), .B2(n18376), .ZN(
        n18559) );
  INV_X1 U39081 ( .I(n47694), .ZN(n47693) );
  NAND2_X1 U39082 ( .A1(n47810), .A2(n47798), .ZN(n47694) );
  NOR2_X2 U39083 ( .A1(n8048), .A2(n45199), .ZN(n47798) );
  AOI21_X1 U39084 ( .A1(n17235), .A2(n18377), .B(n29139), .ZN(n26726) );
  NAND3_X1 U39085 ( .A1(n1350), .A2(n61928), .A3(n30226), .ZN(n30227) );
  AOI21_X1 U39088 ( .A1(n61066), .A2(n4802), .B(n36040), .ZN(n36024) );
  OAI21_X1 U39089 ( .A1(n34465), .A2(n36040), .B(n61066), .ZN(n37617) );
  NOR2_X1 U39090 ( .A1(n18390), .A2(n31767), .ZN(n20181) );
  NAND2_X1 U39091 ( .A1(n33994), .A2(n18390), .ZN(n20314) );
  NOR3_X2 U39093 ( .A1(n18481), .A2(n18480), .A3(n48837), .ZN(n52176) );
  NAND2_X2 U39096 ( .A1(n43438), .A2(n43433), .ZN(n43434) );
  AND2_X1 U39099 ( .A1(n18418), .A2(n25358), .Z(n18417) );
  NAND2_X1 U39101 ( .A1(n23046), .A2(n40443), .ZN(n18420) );
  MUX2_X1 U39103 ( .I0(n41032), .I1(n41033), .S(n36106), .Z(n41042) );
  XOR2_X1 U39105 ( .A1(n60502), .A2(n16311), .Z(n18426) );
  INV_X1 U39107 ( .I(n49192), .ZN(n48283) );
  XOR2_X1 U39108 ( .A1(n4795), .A2(n25887), .Z(n31568) );
  XOR2_X1 U39109 ( .A1(n1288), .A2(n1102), .Z(n50612) );
  NAND3_X1 U39110 ( .A1(n1304), .A2(n41133), .A3(n18441), .ZN(n41136) );
  XOR2_X1 U39112 ( .A1(n18443), .A2(n18442), .Z(n25275) );
  XOR2_X1 U39113 ( .A1(n32405), .A2(n31865), .Z(n18442) );
  XOR2_X1 U39114 ( .A1(n18444), .A2(n52345), .Z(n21616) );
  NAND2_X1 U39117 ( .A1(n43394), .A2(n43692), .ZN(n18448) );
  INV_X1 U39118 ( .I(n19442), .ZN(n18447) );
  XOR2_X1 U39120 ( .A1(n38578), .A2(n24700), .Z(n18453) );
  XOR2_X1 U39121 ( .A1(n18456), .A2(n18455), .Z(n51936) );
  XOR2_X1 U39122 ( .A1(n9231), .A2(n16328), .Z(n18455) );
  XOR2_X1 U39123 ( .A1(n18458), .A2(n18457), .Z(n25715) );
  XOR2_X1 U39124 ( .A1(n46714), .A2(n46626), .Z(n18457) );
  OR2_X1 U39127 ( .A1(n47108), .A2(n47107), .Z(n18459) );
  NOR3_X1 U39131 ( .A1(n29138), .A2(n24940), .A3(n26719), .ZN(n26717) );
  NOR2_X1 U39132 ( .A1(n29137), .A2(n24940), .ZN(n26723) );
  XOR2_X1 U39134 ( .A1(n43332), .A2(n37889), .Z(n50712) );
  XOR2_X1 U39135 ( .A1(n51638), .A2(n43332), .Z(n46585) );
  XOR2_X1 U39136 ( .A1(n43332), .A2(n43333), .Z(n43334) );
  INV_X1 U39137 ( .I(n19766), .ZN(n25599) );
  XOR2_X1 U39140 ( .A1(n18467), .A2(n53805), .Z(n49787) );
  XOR2_X1 U39141 ( .A1(n44014), .A2(n18467), .Z(n46387) );
  XOR2_X1 U39142 ( .A1(n46219), .A2(n18467), .Z(n38850) );
  XOR2_X1 U39143 ( .A1(n31369), .A2(n18467), .Z(n32988) );
  XOR2_X1 U39144 ( .A1(n46284), .A2(n18467), .Z(n46285) );
  XOR2_X1 U39145 ( .A1(n54153), .A2(n23882), .Z(n18467) );
  NOR2_X1 U39147 ( .A1(n28553), .A2(n1564), .ZN(n18470) );
  NAND2_X1 U39150 ( .A1(n19089), .A2(n18476), .ZN(n19088) );
  NAND3_X1 U39151 ( .A1(n45511), .A2(n45510), .A3(n18477), .ZN(n45516) );
  NOR2_X1 U39153 ( .A1(n4275), .A2(n12034), .ZN(n20284) );
  NOR2_X1 U39155 ( .A1(n16527), .A2(n4275), .ZN(n37919) );
  OAI21_X1 U39157 ( .A1(n54640), .A2(n18247), .B(n54848), .ZN(n18484) );
  XOR2_X1 U39158 ( .A1(n50892), .A2(n18485), .Z(n50893) );
  NAND2_X1 U39160 ( .A1(n11571), .A2(n18487), .ZN(n53543) );
  XOR2_X1 U39161 ( .A1(n18490), .A2(n33269), .Z(n31884) );
  XOR2_X1 U39162 ( .A1(n1094), .A2(n62818), .Z(n18492) );
  XOR2_X1 U39163 ( .A1(n19540), .A2(n19541), .Z(n18493) );
  XOR2_X1 U39164 ( .A1(n18495), .A2(n50188), .Z(n18494) );
  XOR2_X1 U39165 ( .A1(n50194), .A2(n19374), .Z(n18495) );
  NAND2_X1 U39166 ( .A1(n23589), .A2(n22416), .ZN(n30840) );
  NOR2_X2 U39167 ( .A1(n18497), .A2(n21154), .ZN(n28270) );
  OAI21_X1 U39168 ( .A1(n28271), .A2(n61035), .B(n18497), .ZN(n27061) );
  XOR2_X1 U39169 ( .A1(n25377), .A2(n16295), .Z(n37624) );
  INV_X1 U39170 ( .I(n18508), .ZN(n18503) );
  NAND2_X1 U39172 ( .A1(n34777), .A2(n34786), .ZN(n18506) );
  XOR2_X1 U39174 ( .A1(n25363), .A2(n25872), .Z(n18513) );
  XOR2_X1 U39175 ( .A1(n39193), .A2(n38572), .Z(n18514) );
  XOR2_X1 U39178 ( .A1(n43161), .A2(n20601), .Z(n42563) );
  INV_X2 U39180 ( .I(n2998), .ZN(n19389) );
  XOR2_X1 U39183 ( .A1(n38159), .A2(n19044), .Z(n18539) );
  XOR2_X1 U39184 ( .A1(n18542), .A2(n18544), .Z(n18541) );
  OAI22_X1 U39185 ( .A1(n34376), .A2(n37371), .B1(n36512), .B2(n2592), .ZN(
        n18546) );
  MUX2_X1 U39186 ( .I0(n55850), .I1(n55851), .S(n19953), .Z(n55860) );
  NOR3_X1 U39187 ( .A1(n55900), .A2(n55899), .A3(n55898), .ZN(n18558) );
  NAND2_X1 U39188 ( .A1(n55898), .A2(n55893), .ZN(n18560) );
  NAND2_X2 U39191 ( .A1(n54767), .A2(n54768), .ZN(n54759) );
  XOR2_X1 U39195 ( .A1(n18580), .A2(n16106), .Z(n21608) );
  XOR2_X1 U39196 ( .A1(n18584), .A2(n46612), .Z(n46613) );
  NAND2_X1 U39197 ( .A1(n63261), .A2(n18585), .ZN(n49993) );
  NOR2_X1 U39201 ( .A1(n47434), .A2(n18590), .ZN(n47442) );
  NOR2_X1 U39202 ( .A1(n45450), .A2(n18590), .ZN(n43752) );
  NAND2_X1 U39208 ( .A1(n18597), .A2(n56229), .ZN(n56231) );
  OAI21_X1 U39209 ( .A1(n18597), .A2(n24473), .B(n56436), .ZN(n51901) );
  NAND2_X2 U39210 ( .A1(n18600), .A2(n9229), .ZN(n18598) );
  NOR2_X1 U39211 ( .A1(n41634), .A2(n18603), .ZN(n25928) );
  XOR2_X1 U39213 ( .A1(n64258), .A2(n18605), .Z(n46693) );
  XOR2_X1 U39214 ( .A1(n4529), .A2(n46689), .Z(n18605) );
  NAND2_X2 U39216 ( .A1(n18609), .A2(n1224), .ZN(n50288) );
  NAND2_X2 U39219 ( .A1(n21784), .A2(n23106), .ZN(n18606) );
  INV_X2 U39220 ( .I(n53998), .ZN(n53992) );
  NAND3_X2 U39221 ( .A1(n53998), .A2(n18619), .A3(n18618), .ZN(n53995) );
  NOR2_X2 U39222 ( .A1(n18621), .A2(n18620), .ZN(n53998) );
  NOR2_X2 U39223 ( .A1(n40754), .A2(n18623), .ZN(n40759) );
  NOR2_X1 U39224 ( .A1(n18623), .A2(n40749), .ZN(n41467) );
  OR2_X1 U39225 ( .A1(n40417), .A2(n18623), .Z(n18622) );
  XOR2_X1 U39226 ( .A1(n18624), .A2(n46629), .Z(n20806) );
  XOR2_X1 U39229 ( .A1(n32540), .A2(n17104), .Z(n32499) );
  INV_X1 U39232 ( .I(n12004), .ZN(n35063) );
  XOR2_X1 U39234 ( .A1(n18639), .A2(n18640), .Z(n18638) );
  XOR2_X1 U39235 ( .A1(n51593), .A2(n18642), .Z(n18640) );
  NAND3_X1 U39242 ( .A1(n40103), .A2(n18649), .A3(n40104), .ZN(n25923) );
  NAND2_X1 U39244 ( .A1(n40048), .A2(n18649), .ZN(n40050) );
  CLKBUF_X4 U39245 ( .I(n33847), .Z(n18651) );
  NAND2_X1 U39247 ( .A1(n54197), .A2(n54198), .ZN(n54205) );
  XOR2_X1 U39250 ( .A1(n33892), .A2(n18674), .Z(n21937) );
  XOR2_X1 U39251 ( .A1(n18676), .A2(n18675), .Z(n18674) );
  XOR2_X1 U39252 ( .A1(n21531), .A2(n33890), .Z(n18676) );
  AOI21_X1 U39254 ( .A1(n15720), .A2(n18205), .B(n18677), .ZN(n34891) );
  NAND3_X1 U39255 ( .A1(n60684), .A2(n34196), .A3(n21409), .ZN(n18681) );
  XOR2_X1 U39257 ( .A1(n18686), .A2(n51334), .Z(n18685) );
  XOR2_X1 U39258 ( .A1(n51684), .A2(n51340), .Z(n18686) );
  XOR2_X1 U39259 ( .A1(n7070), .A2(n51341), .Z(n18687) );
  NOR2_X2 U39262 ( .A1(n8474), .A2(n4802), .ZN(n35583) );
  AOI22_X1 U39263 ( .A1(n18690), .A2(n48832), .B1(n48279), .B2(n24393), .ZN(
        n47753) );
  NOR2_X1 U39266 ( .A1(n18691), .A2(n30408), .ZN(n30412) );
  XOR2_X1 U39268 ( .A1(n18708), .A2(n31503), .Z(n18696) );
  NAND3_X1 U39269 ( .A1(n18700), .A2(n22081), .A3(n55034), .ZN(n22080) );
  INV_X2 U39270 ( .I(n18701), .ZN(n23217) );
  XOR2_X1 U39273 ( .A1(n18707), .A2(n25886), .Z(n18708) );
  XOR2_X1 U39274 ( .A1(n59622), .A2(n31507), .Z(n18707) );
  INV_X1 U39275 ( .I(n19285), .ZN(n22227) );
  AOI21_X1 U39278 ( .A1(n18716), .A2(n29516), .B(n29521), .ZN(n29517) );
  AOI21_X2 U39283 ( .A1(n40080), .A2(n40079), .B(n25468), .ZN(n43468) );
  INV_X2 U39284 ( .I(n42986), .ZN(n43947) );
  INV_X1 U39285 ( .I(n15810), .ZN(n44993) );
  INV_X1 U39286 ( .I(n30936), .ZN(n18729) );
  XOR2_X1 U39287 ( .A1(n23246), .A2(n9040), .Z(n18730) );
  NAND2_X2 U39290 ( .A1(n18737), .A2(n55264), .ZN(n54842) );
  NOR2_X1 U39293 ( .A1(n18747), .A2(n27615), .ZN(n27616) );
  INV_X1 U39296 ( .I(n29514), .ZN(n30952) );
  NAND2_X1 U39297 ( .A1(n42942), .A2(n18770), .ZN(n41753) );
  INV_X2 U39298 ( .I(n18774), .ZN(n55494) );
  NAND4_X1 U39299 ( .A1(n1524), .A2(n21536), .A3(n20124), .A4(n37359), .ZN(
        n18777) );
  NOR2_X1 U39300 ( .A1(n7499), .A2(n18780), .ZN(n27978) );
  NAND2_X2 U39304 ( .A1(n55203), .A2(n18786), .ZN(n55219) );
  OAI21_X1 U39305 ( .A1(n18786), .A2(n55222), .B(n55225), .ZN(n22466) );
  NOR2_X1 U39306 ( .A1(n57628), .A2(n18789), .ZN(n18788) );
  INV_X1 U39307 ( .I(n35821), .ZN(n18789) );
  XOR2_X1 U39308 ( .A1(n19008), .A2(n38944), .Z(n38945) );
  XOR2_X1 U39309 ( .A1(n18797), .A2(n49897), .Z(n37720) );
  XOR2_X1 U39310 ( .A1(n38300), .A2(n18797), .Z(n38104) );
  INV_X1 U39315 ( .I(n18810), .ZN(n31140) );
  NAND2_X1 U39316 ( .A1(n29487), .A2(n18810), .ZN(n29483) );
  NOR2_X1 U39320 ( .A1(n49546), .A2(n49545), .ZN(n18819) );
  INV_X2 U39321 ( .I(n11329), .ZN(n20473) );
  XOR2_X1 U39322 ( .A1(n65046), .A2(n38586), .Z(n18830) );
  NAND2_X1 U39323 ( .A1(n35744), .A2(n18835), .ZN(n25309) );
  NOR2_X1 U39324 ( .A1(n18836), .A2(n7012), .ZN(n40642) );
  AOI21_X1 U39325 ( .A1(n40540), .A2(n39073), .B(n18836), .ZN(n39077) );
  XOR2_X1 U39326 ( .A1(n32470), .A2(n46336), .Z(n18837) );
  XOR2_X1 U39327 ( .A1(n51386), .A2(n51589), .Z(n18846) );
  XOR2_X1 U39328 ( .A1(n46216), .A2(n46558), .Z(n46217) );
  XOR2_X1 U39329 ( .A1(n17300), .A2(n46216), .Z(n44498) );
  MUX2_X1 U39331 ( .I0(n28522), .I1(n28521), .S(n18848), .Z(n28523) );
  INV_X2 U39332 ( .I(n38600), .ZN(n40523) );
  INV_X1 U39333 ( .I(n18850), .ZN(n36378) );
  NAND2_X1 U39334 ( .A1(n35533), .A2(n18850), .ZN(n35536) );
  OAI21_X1 U39335 ( .A1(n36380), .A2(n36572), .B(n18850), .ZN(n35188) );
  OAI21_X1 U39336 ( .A1(n19364), .A2(n36572), .B(n18850), .ZN(n32985) );
  XOR2_X1 U39338 ( .A1(n32493), .A2(n21563), .Z(n18855) );
  INV_X2 U39339 ( .I(n54191), .ZN(n54207) );
  XNOR2_X1 U39340 ( .A1(n21986), .A2(n31797), .ZN(n18964) );
  XOR2_X1 U39341 ( .A1(n30833), .A2(n32044), .Z(n31797) );
  NOR2_X1 U39342 ( .A1(n29610), .A2(n12741), .ZN(n29601) );
  OAI21_X1 U39343 ( .A1(n11873), .A2(n28665), .B(n12741), .ZN(n27700) );
  NAND2_X1 U39344 ( .A1(n28664), .A2(n12741), .ZN(n28668) );
  NAND2_X1 U39349 ( .A1(n24041), .A2(n18877), .ZN(n36160) );
  AND2_X1 U39352 ( .A1(n28671), .A2(n28668), .Z(n18881) );
  XOR2_X1 U39360 ( .A1(n18899), .A2(n18897), .Z(n24617) );
  XOR2_X1 U39361 ( .A1(n60532), .A2(n18898), .Z(n18897) );
  XOR2_X1 U39362 ( .A1(n38580), .A2(n38579), .Z(n18898) );
  XOR2_X1 U39364 ( .A1(n46145), .A2(n43863), .Z(n18902) );
  NOR2_X1 U39366 ( .A1(n5082), .A2(n1542), .ZN(n20137) );
  OAI21_X1 U39367 ( .A1(n23127), .A2(n5082), .B(n33405), .ZN(n31656) );
  NAND2_X1 U39368 ( .A1(n49556), .A2(n18918), .ZN(n49557) );
  XOR2_X1 U39370 ( .A1(n19121), .A2(n23927), .Z(n38309) );
  XOR2_X1 U39371 ( .A1(n19926), .A2(n18920), .Z(n45119) );
  XOR2_X1 U39372 ( .A1(n45281), .A2(n42790), .Z(n18920) );
  XOR2_X1 U39374 ( .A1(n18924), .A2(n37508), .Z(n18923) );
  XOR2_X1 U39375 ( .A1(n38310), .A2(n35194), .Z(n37509) );
  XOR2_X1 U39376 ( .A1(n37507), .A2(n39238), .Z(n18924) );
  NOR2_X1 U39378 ( .A1(n5227), .A2(n15782), .ZN(n18926) );
  NAND2_X1 U39380 ( .A1(n18930), .A2(n28342), .ZN(n28354) );
  NOR2_X1 U39383 ( .A1(n27579), .A2(n27567), .ZN(n18938) );
  XOR2_X1 U39387 ( .A1(n23907), .A2(n38527), .Z(n18941) );
  NAND3_X1 U39388 ( .A1(n35657), .A2(n35655), .A3(n35656), .ZN(n18947) );
  NAND2_X1 U39393 ( .A1(n22647), .A2(n18951), .ZN(n45077) );
  XOR2_X1 U39397 ( .A1(n14037), .A2(n43725), .Z(n18954) );
  XOR2_X1 U39398 ( .A1(n45017), .A2(n45018), .Z(n18956) );
  XOR2_X1 U39399 ( .A1(n44386), .A2(n41553), .Z(n18957) );
  XOR2_X1 U39400 ( .A1(n18964), .A2(n18959), .Z(n18963) );
  XOR2_X1 U39401 ( .A1(n32000), .A2(n19306), .Z(n18959) );
  XOR2_X1 U39402 ( .A1(n18965), .A2(n25331), .Z(n32000) );
  XOR2_X1 U39404 ( .A1(n31859), .A2(n18961), .Z(n18960) );
  XOR2_X1 U39405 ( .A1(n18962), .A2(n59546), .Z(n18961) );
  XOR2_X1 U39407 ( .A1(n18967), .A2(n38538), .Z(n18966) );
  XOR2_X1 U39408 ( .A1(n38531), .A2(n18968), .Z(n18967) );
  XOR2_X1 U39409 ( .A1(n23330), .A2(n38530), .Z(n18968) );
  XOR2_X1 U39411 ( .A1(n39561), .A2(n39563), .Z(n18972) );
  NAND2_X1 U39412 ( .A1(n22700), .A2(n24081), .ZN(n18973) );
  NOR2_X2 U39413 ( .A1(n47435), .A2(n47730), .ZN(n22700) );
  INV_X2 U39414 ( .I(n49565), .ZN(n19867) );
  NOR2_X2 U39415 ( .A1(n18982), .A2(n18978), .ZN(n49565) );
  XOR2_X1 U39418 ( .A1(n787), .A2(n43688), .Z(n18987) );
  NAND2_X2 U39419 ( .A1(n43980), .A2(n16880), .ZN(n43306) );
  NOR3_X1 U39420 ( .A1(n25131), .A2(n41469), .A3(n40749), .ZN(n40751) );
  NOR2_X2 U39421 ( .A1(n11229), .A2(n42160), .ZN(n43338) );
  XOR2_X1 U39422 ( .A1(n18998), .A2(n18996), .Z(n25884) );
  XOR2_X1 U39423 ( .A1(n18997), .A2(n746), .Z(n18996) );
  XOR2_X1 U39424 ( .A1(n38750), .A2(n38749), .Z(n18997) );
  XOR2_X1 U39427 ( .A1(n19002), .A2(n21094), .Z(n33229) );
  XOR2_X1 U39428 ( .A1(n10531), .A2(n26237), .Z(n19002) );
  NOR2_X2 U39430 ( .A1(n41779), .A2(n42878), .ZN(n19004) );
  AOI22_X1 U39433 ( .A1(n19004), .A2(n42869), .B1(n43817), .B2(n42870), .ZN(
        n42885) );
  INV_X2 U39434 ( .I(n19006), .ZN(n34308) );
  NOR2_X2 U39435 ( .A1(n34308), .A2(n34761), .ZN(n34307) );
  XOR2_X1 U39436 ( .A1(n19009), .A2(n19008), .Z(n23044) );
  NAND2_X1 U39441 ( .A1(n15700), .A2(n19020), .ZN(n19022) );
  INV_X1 U39443 ( .I(n19894), .ZN(n19024) );
  NOR2_X1 U39444 ( .A1(n19894), .A2(n34779), .ZN(n19025) );
  XOR2_X1 U39446 ( .A1(n19034), .A2(n55898), .Z(n19033) );
  NAND3_X1 U39447 ( .A1(n15716), .A2(n55842), .A3(n60203), .ZN(n19037) );
  NAND2_X1 U39448 ( .A1(n49499), .A2(n19043), .ZN(n25313) );
  INV_X1 U39449 ( .I(n19048), .ZN(n22806) );
  XOR2_X1 U39450 ( .A1(n63099), .A2(n19048), .Z(n33205) );
  XOR2_X1 U39451 ( .A1(n23786), .A2(n19048), .Z(n32119) );
  NAND3_X1 U39452 ( .A1(n33442), .A2(n33446), .A3(n19053), .ZN(n33443) );
  INV_X1 U39453 ( .I(n19054), .ZN(n57105) );
  NOR2_X2 U39455 ( .A1(n21570), .A2(n21569), .ZN(n19054) );
  XOR2_X1 U39456 ( .A1(n32620), .A2(n19056), .Z(n19055) );
  XOR2_X1 U39457 ( .A1(n60902), .A2(n19057), .Z(n19056) );
  XOR2_X1 U39458 ( .A1(n16959), .A2(n31198), .Z(n19058) );
  XOR2_X1 U39459 ( .A1(n64285), .A2(n13705), .Z(n25642) );
  MUX2_X1 U39460 ( .I0(n48778), .I1(n49545), .S(n18769), .Z(n48788) );
  XOR2_X1 U39462 ( .A1(n39359), .A2(n20317), .Z(n19067) );
  NOR3_X1 U39463 ( .A1(n53601), .A2(n19068), .A3(n53196), .ZN(n53201) );
  INV_X1 U39465 ( .I(n19078), .ZN(n41004) );
  NAND2_X1 U39466 ( .A1(n19078), .A2(n23355), .ZN(n40608) );
  NOR2_X2 U39469 ( .A1(n23666), .A2(n47680), .ZN(n47425) );
  XOR2_X1 U39470 ( .A1(n31421), .A2(n19091), .Z(n19090) );
  XOR2_X1 U39471 ( .A1(n31316), .A2(n19092), .Z(n19091) );
  XOR2_X1 U39472 ( .A1(n32661), .A2(n32118), .Z(n19092) );
  XOR2_X1 U39474 ( .A1(n25063), .A2(n18296), .Z(n19094) );
  XOR2_X1 U39479 ( .A1(n22212), .A2(n46391), .Z(n46393) );
  XOR2_X1 U39480 ( .A1(n22212), .A2(n44088), .Z(n44089) );
  NAND3_X2 U39482 ( .A1(n40050), .A2(n40333), .A3(n19105), .ZN(n25853) );
  NAND4_X1 U39483 ( .A1(n54573), .A2(n58810), .A3(n18425), .A4(n18422), .ZN(
        n54520) );
  XOR2_X1 U39484 ( .A1(n19106), .A2(n16032), .Z(n25714) );
  XOR2_X1 U39485 ( .A1(n46610), .A2(n22876), .Z(n19106) );
  NAND3_X2 U39486 ( .A1(n24555), .A2(n15949), .A3(n56432), .ZN(n24552) );
  NAND2_X1 U39487 ( .A1(n25141), .A2(n13811), .ZN(n40047) );
  NOR2_X1 U39488 ( .A1(n34436), .A2(n34435), .ZN(n19108) );
  AND2_X1 U39489 ( .A1(n54546), .A2(n58896), .Z(n54566) );
  NOR2_X1 U39490 ( .A1(n28753), .A2(n58816), .ZN(n19191) );
  NOR3_X1 U39493 ( .A1(n40034), .A2(n41844), .A3(n25665), .ZN(n25664) );
  AOI22_X1 U39494 ( .A1(n19109), .A2(n36226), .B1(n35161), .B2(n35162), .ZN(
        n35167) );
  NOR2_X1 U39495 ( .A1(n35160), .A2(n23257), .ZN(n19109) );
  NAND2_X1 U39496 ( .A1(n40383), .A2(n40385), .ZN(n19212) );
  BUF_X4 U39497 ( .I(n51461), .Z(n56775) );
  NAND2_X1 U39498 ( .A1(n40693), .A2(n40694), .ZN(n40706) );
  XOR2_X1 U39502 ( .A1(n31577), .A2(n32408), .Z(n20834) );
  OAI22_X1 U39503 ( .A1(n19114), .A2(n49245), .B1(n2878), .B2(n47456), .ZN(
        n48763) );
  OR2_X1 U39504 ( .A1(n48754), .A2(n25680), .Z(n19114) );
  XOR2_X1 U39505 ( .A1(n38193), .A2(n38637), .Z(n19352) );
  AND2_X1 U39506 ( .A1(n39093), .A2(n39092), .Z(n25567) );
  NOR2_X2 U39511 ( .A1(n57281), .A2(n43190), .ZN(n20492) );
  NAND2_X1 U39514 ( .A1(n52212), .A2(n52213), .ZN(n19409) );
  XOR2_X1 U39516 ( .A1(n35358), .A2(n39345), .Z(n19121) );
  MUX2_X1 U39517 ( .I0(n1811), .I1(n32684), .S(n35200), .Z(n33554) );
  AOI22_X1 U39518 ( .A1(n19123), .A2(n34142), .B1(n34138), .B2(n19416), .ZN(
        n32820) );
  NAND2_X1 U39519 ( .A1(n34133), .A2(n65232), .ZN(n19123) );
  NOR2_X2 U39520 ( .A1(n35709), .A2(n34404), .ZN(n35235) );
  BUF_X4 U39521 ( .I(n40651), .Z(n20602) );
  XOR2_X1 U39525 ( .A1(n23929), .A2(n55191), .Z(n19126) );
  XOR2_X1 U39526 ( .A1(n32279), .A2(n31744), .Z(n25973) );
  XOR2_X1 U39527 ( .A1(n44355), .A2(n44353), .Z(n20335) );
  NAND3_X1 U39529 ( .A1(n36488), .A2(n1525), .A3(n22527), .ZN(n19127) );
  INV_X2 U39530 ( .I(n32699), .ZN(n34138) );
  NAND2_X1 U39533 ( .A1(n47344), .A2(n19849), .ZN(n19848) );
  XOR2_X1 U39535 ( .A1(n19129), .A2(n47448), .Z(n47462) );
  XOR2_X1 U39536 ( .A1(n47351), .A2(n47352), .Z(n19129) );
  NOR3_X1 U39538 ( .A1(n20740), .A2(n54452), .A3(n55020), .ZN(n19131) );
  XOR2_X1 U39539 ( .A1(n19372), .A2(n19134), .Z(n23592) );
  XOR2_X1 U39540 ( .A1(n21985), .A2(n33860), .Z(n19134) );
  NAND2_X2 U39541 ( .A1(n47036), .A2(n16938), .ZN(n19595) );
  NAND2_X1 U39544 ( .A1(n19137), .A2(n54657), .ZN(n21617) );
  NOR2_X2 U39545 ( .A1(n43757), .A2(n49323), .ZN(n49388) );
  NAND2_X1 U39548 ( .A1(n42380), .A2(n19292), .ZN(n42382) );
  XOR2_X1 U39550 ( .A1(n19140), .A2(n23306), .Z(Plaintext[73]) );
  NAND2_X2 U39558 ( .A1(n23479), .A2(n29371), .ZN(n27328) );
  XOR2_X1 U39559 ( .A1(n22697), .A2(n23019), .Z(n39393) );
  NAND3_X1 U39560 ( .A1(n26989), .A2(n29372), .A3(n26988), .ZN(n24476) );
  XOR2_X1 U39561 ( .A1(n51320), .A2(n1621), .Z(n21757) );
  OR2_X1 U39562 ( .A1(n61008), .A2(n41058), .Z(n20024) );
  NOR2_X1 U39563 ( .A1(n47385), .A2(n47798), .ZN(n47389) );
  AOI21_X1 U39565 ( .A1(n54368), .A2(n22782), .B(n5323), .ZN(n26109) );
  OAI22_X1 U39568 ( .A1(n53757), .A2(n53758), .B1(n53756), .B2(n16489), .ZN(
        n19147) );
  AND2_X1 U39569 ( .A1(n22093), .A2(n63953), .Z(n19685) );
  OAI21_X1 U39571 ( .A1(n47411), .A2(n47690), .B(n21199), .ZN(n19150) );
  NAND2_X2 U39574 ( .A1(n20277), .A2(n38264), .ZN(n41854) );
  XOR2_X1 U39575 ( .A1(n19152), .A2(n23754), .Z(Plaintext[45]) );
  INV_X1 U39578 ( .I(n50755), .ZN(n50756) );
  OR2_X1 U39584 ( .A1(n20925), .A2(n14462), .Z(n38417) );
  INV_X1 U39585 ( .I(n20994), .ZN(n25839) );
  NAND4_X1 U39589 ( .A1(n36833), .A2(n36832), .A3(n36831), .A4(n36830), .ZN(
        n19165) );
  NAND2_X2 U39590 ( .A1(n58559), .A2(n28495), .ZN(n28494) );
  XOR2_X1 U39591 ( .A1(n20717), .A2(n21024), .Z(n23388) );
  NOR2_X1 U39592 ( .A1(n21576), .A2(n21575), .ZN(n19301) );
  OAI21_X2 U39593 ( .A1(n27735), .A2(n27734), .B(n30018), .ZN(n27737) );
  XOR2_X1 U39596 ( .A1(n19177), .A2(n56495), .Z(Plaintext[159]) );
  INV_X1 U39598 ( .I(n55499), .ZN(n20927) );
  XOR2_X1 U39599 ( .A1(n18191), .A2(n16327), .Z(n21686) );
  OR3_X1 U39602 ( .A1(n22947), .A2(n54997), .A3(n52477), .Z(n19187) );
  NAND2_X2 U39603 ( .A1(n3055), .A2(n4734), .ZN(n20763) );
  INV_X4 U39606 ( .I(n48082), .ZN(n48559) );
  NOR2_X1 U39608 ( .A1(n28752), .A2(n29241), .ZN(n19192) );
  BUF_X4 U39611 ( .I(n35651), .Z(n22909) );
  NAND3_X1 U39617 ( .A1(n54314), .A2(n21296), .A3(n1610), .ZN(n19208) );
  NOR2_X1 U39619 ( .A1(n41006), .A2(n1275), .ZN(n19209) );
  XOR2_X1 U39624 ( .A1(n13639), .A2(n52067), .Z(n20545) );
  NOR2_X1 U39625 ( .A1(n43159), .A2(n43158), .ZN(n19214) );
  XOR2_X1 U39626 ( .A1(n46206), .A2(n44272), .Z(n19215) );
  NAND2_X1 U39627 ( .A1(n36234), .A2(n19617), .ZN(n32769) );
  NAND2_X1 U39631 ( .A1(n25010), .A2(n5936), .ZN(n19221) );
  BUF_X2 U39632 ( .I(n26086), .Z(n19224) );
  NAND2_X2 U39635 ( .A1(n40239), .A2(n40070), .ZN(n40163) );
  NOR2_X1 U39637 ( .A1(n28394), .A2(n28395), .ZN(n19227) );
  NAND3_X1 U39638 ( .A1(n22534), .A2(n47197), .A3(n48196), .ZN(n47200) );
  NAND4_X2 U39640 ( .A1(n19230), .A2(n42307), .A3(n42305), .A4(n42306), .ZN(
        n20527) );
  OR2_X2 U39641 ( .A1(n58825), .A2(n25267), .Z(n53797) );
  OAI21_X2 U39642 ( .A1(n47812), .A2(n47811), .B(n47810), .ZN(n47816) );
  XOR2_X1 U39644 ( .A1(n45874), .A2(n21316), .Z(n19237) );
  XOR2_X1 U39645 ( .A1(n24593), .A2(n46590), .Z(n24592) );
  XOR2_X1 U39646 ( .A1(n19238), .A2(n46588), .Z(n46589) );
  XOR2_X1 U39647 ( .A1(n21516), .A2(n10449), .Z(n19238) );
  AND3_X1 U39651 ( .A1(n48694), .A2(n48693), .A3(n48692), .Z(n19242) );
  NAND2_X2 U39653 ( .A1(n59020), .A2(n15434), .ZN(n53220) );
  NAND3_X1 U39654 ( .A1(n40304), .A2(n40296), .A3(n40029), .ZN(n40030) );
  INV_X1 U39655 ( .I(n61895), .ZN(n55402) );
  INV_X1 U39657 ( .I(n38304), .ZN(n22266) );
  NAND2_X2 U39660 ( .A1(n1458), .A2(n55300), .ZN(n55296) );
  NAND2_X1 U39663 ( .A1(n32598), .A2(n33639), .ZN(n32599) );
  XOR2_X1 U39665 ( .A1(n19254), .A2(n53103), .Z(Plaintext[4]) );
  NAND2_X2 U39666 ( .A1(n58267), .A2(n21584), .ZN(n34896) );
  NAND2_X2 U39668 ( .A1(n27885), .A2(n27884), .ZN(n27905) );
  AND2_X2 U39669 ( .A1(n28542), .A2(n28537), .Z(n27871) );
  NAND2_X1 U39671 ( .A1(n19263), .A2(n19042), .ZN(n25783) );
  INV_X4 U39673 ( .I(n16102), .ZN(n38675) );
  INV_X2 U39674 ( .I(n19269), .ZN(n21720) );
  XOR2_X1 U39675 ( .A1(n21721), .A2(Ciphertext[82]), .Z(n19269) );
  NAND3_X1 U39679 ( .A1(n30525), .A2(n1351), .A3(n20364), .ZN(n20155) );
  NAND2_X2 U39680 ( .A1(n24987), .A2(n18075), .ZN(n20364) );
  OAI21_X1 U39682 ( .A1(n27457), .A2(n27358), .B(n57424), .ZN(n19917) );
  NAND2_X1 U39683 ( .A1(n19917), .A2(n19915), .ZN(n19914) );
  AOI22_X1 U39684 ( .A1(n41362), .A2(n60131), .B1(n42151), .B2(n41369), .ZN(
        n41365) );
  NOR3_X2 U39685 ( .A1(n24461), .A2(n19275), .A3(n24460), .ZN(n24459) );
  INV_X1 U39686 ( .I(n35547), .ZN(n21694) );
  NAND2_X1 U39690 ( .A1(n35397), .A2(n35398), .ZN(n19281) );
  XOR2_X1 U39692 ( .A1(n19285), .A2(n31193), .Z(n25886) );
  NOR2_X1 U39695 ( .A1(n24717), .A2(n24723), .ZN(n24716) );
  NOR2_X1 U39698 ( .A1(n19588), .A2(n31104), .ZN(n19289) );
  OR2_X1 U39700 ( .A1(n23108), .A2(n11459), .Z(n39851) );
  OAI21_X1 U39701 ( .A1(n23411), .A2(n53253), .B(n53250), .ZN(n19676) );
  XNOR2_X1 U39702 ( .A1(n11922), .A2(n42627), .ZN(n25250) );
  NAND2_X2 U39704 ( .A1(n64391), .A2(n42080), .ZN(n42405) );
  XOR2_X1 U39705 ( .A1(n20145), .A2(n31700), .Z(n20144) );
  OR2_X1 U39709 ( .A1(n54920), .A2(n19300), .Z(n54923) );
  NAND4_X2 U39710 ( .A1(n33311), .A2(n33310), .A3(n33309), .A4(n33308), .ZN(
        n33312) );
  NAND3_X1 U39713 ( .A1(n55974), .A2(n55976), .A3(n55973), .ZN(n55978) );
  NAND3_X1 U39714 ( .A1(n55974), .A2(n55976), .A3(n1600), .ZN(n55458) );
  NAND3_X1 U39716 ( .A1(n27474), .A2(n27473), .A3(n27475), .ZN(n23200) );
  NOR2_X2 U39717 ( .A1(n29316), .A2(n23596), .ZN(n27448) );
  XOR2_X1 U39718 ( .A1(n33075), .A2(n30987), .Z(n29868) );
  INV_X1 U39719 ( .I(n48145), .ZN(n46751) );
  INV_X4 U39720 ( .I(n21409), .ZN(n31767) );
  XOR2_X1 U39721 ( .A1(n24090), .A2(n29407), .Z(n25518) );
  XOR2_X1 U39724 ( .A1(n26920), .A2(n31857), .Z(n19306) );
  AOI22_X1 U39727 ( .A1(n42675), .A2(n60131), .B1(n6706), .B2(n42674), .ZN(
        n42680) );
  NAND4_X2 U39729 ( .A1(n22954), .A2(n37015), .A3(n37014), .A4(n23050), .ZN(
        n38742) );
  XOR2_X1 U39733 ( .A1(n50184), .A2(n50185), .Z(n50186) );
  NAND3_X1 U39737 ( .A1(n19319), .A2(n42348), .A3(n42349), .ZN(n42350) );
  XOR2_X1 U39738 ( .A1(n10553), .A2(n31802), .Z(n31803) );
  INV_X1 U39739 ( .I(n57018), .ZN(n19321) );
  XOR2_X1 U39743 ( .A1(n17801), .A2(n51171), .Z(n19323) );
  AOI21_X1 U39744 ( .A1(n34908), .A2(n35425), .B(n11393), .ZN(n24399) );
  XOR2_X1 U39745 ( .A1(n39257), .A2(n16011), .Z(n22067) );
  NAND2_X1 U39746 ( .A1(n53421), .A2(n53616), .ZN(n52782) );
  NOR3_X2 U39747 ( .A1(n48050), .A2(n48051), .A3(n48049), .ZN(n19324) );
  NAND4_X2 U39749 ( .A1(n19378), .A2(n19377), .A3(n15768), .A4(n21821), .ZN(
        n23533) );
  NAND2_X2 U39750 ( .A1(n23112), .A2(n26182), .ZN(n39992) );
  XOR2_X1 U39755 ( .A1(n21361), .A2(n52321), .Z(n19330) );
  NAND2_X2 U39756 ( .A1(n19646), .A2(n47347), .ZN(n47343) );
  NAND2_X2 U39757 ( .A1(n45493), .A2(n2024), .ZN(n23113) );
  XNOR2_X1 U39758 ( .A1(n51675), .A2(n51674), .ZN(n19889) );
  AND2_X1 U39759 ( .A1(n20423), .A2(n64878), .Z(n19392) );
  NAND3_X2 U39762 ( .A1(n28866), .A2(n28865), .A3(n28867), .ZN(n30664) );
  OAI21_X1 U39763 ( .A1(n19337), .A2(n24072), .B(n33424), .ZN(n31027) );
  NAND2_X1 U39765 ( .A1(n20797), .A2(n27475), .ZN(n19338) );
  INV_X2 U39766 ( .I(n19340), .ZN(n27479) );
  XOR2_X1 U39768 ( .A1(n63955), .A2(n23690), .Z(n19341) );
  NOR3_X2 U39769 ( .A1(n33817), .A2(n33816), .A3(n19344), .ZN(n33818) );
  NOR3_X1 U39770 ( .A1(n35754), .A2(n1546), .A3(n59930), .ZN(n19344) );
  NAND2_X2 U39776 ( .A1(n42175), .A2(n42871), .ZN(n43816) );
  OR3_X1 U39777 ( .A1(n47505), .A2(n45479), .A3(n1480), .Z(n44671) );
  AND2_X1 U39778 ( .A1(n43851), .A2(n10990), .Z(n43853) );
  NOR2_X2 U39779 ( .A1(n26765), .A2(n23303), .ZN(n26764) );
  XOR2_X1 U39782 ( .A1(n3604), .A2(n38595), .Z(n19360) );
  INV_X1 U39783 ( .I(n52645), .ZN(n55161) );
  NAND3_X1 U39784 ( .A1(n55095), .A2(n55096), .A3(n55097), .ZN(n55104) );
  NAND2_X1 U39786 ( .A1(n21775), .A2(n16920), .ZN(n19432) );
  NOR2_X1 U39787 ( .A1(n53157), .A2(n53158), .ZN(n53173) );
  NAND2_X2 U39788 ( .A1(n7979), .A2(n29458), .ZN(n29448) );
  XOR2_X1 U39793 ( .A1(n33866), .A2(n33865), .Z(n19372) );
  XOR2_X1 U39795 ( .A1(n50193), .A2(n7459), .Z(n19374) );
  OAI22_X1 U39798 ( .A1(n53114), .A2(n53113), .B1(n53116), .B2(n19080), .ZN(
        n53121) );
  INV_X1 U39802 ( .I(n19838), .ZN(n19835) );
  INV_X2 U39804 ( .I(n28670), .ZN(n28168) );
  NAND2_X2 U39809 ( .A1(n49538), .A2(n6015), .ZN(n49376) );
  XOR2_X1 U39810 ( .A1(n51053), .A2(n51475), .Z(n49456) );
  XOR2_X1 U39811 ( .A1(n20774), .A2(n1290), .Z(n51053) );
  XOR2_X1 U39812 ( .A1(n50683), .A2(n10101), .Z(n51284) );
  XOR2_X1 U39815 ( .A1(n19390), .A2(n9660), .Z(n36157) );
  XOR2_X1 U39816 ( .A1(n24058), .A2(n36148), .Z(n19390) );
  OR2_X2 U39817 ( .A1(n43460), .A2(n10457), .Z(n42067) );
  INV_X2 U39820 ( .I(n19393), .ZN(n19567) );
  NOR2_X2 U39822 ( .A1(n20426), .A2(n46033), .ZN(n46028) );
  NAND2_X1 U39823 ( .A1(n26716), .A2(n26715), .ZN(n25574) );
  XOR2_X1 U39824 ( .A1(n21084), .A2(n32393), .Z(n19395) );
  AOI21_X1 U39827 ( .A1(n19397), .A2(n19000), .B(n43517), .ZN(n40779) );
  XOR2_X1 U39829 ( .A1(n46620), .A2(n46432), .Z(n44910) );
  NAND2_X2 U39836 ( .A1(n7092), .A2(n36853), .ZN(n35404) );
  AND3_X1 U39847 ( .A1(n56619), .A2(n58846), .A3(n60129), .Z(n20002) );
  NOR3_X1 U39848 ( .A1(n64751), .A2(n50211), .A3(n50213), .ZN(n47995) );
  NOR2_X1 U39849 ( .A1(n35468), .A2(n15720), .ZN(n35467) );
  INV_X4 U39852 ( .I(n23086), .ZN(n33375) );
  BUF_X2 U39855 ( .I(n52416), .Z(n20512) );
  XOR2_X1 U39858 ( .A1(n51159), .A2(n50980), .Z(n50981) );
  XOR2_X1 U39859 ( .A1(Ciphertext[139]), .A2(Key[98]), .Z(n19426) );
  OR3_X1 U39862 ( .A1(n20895), .A2(n19246), .A3(n34534), .Z(n34536) );
  NAND2_X1 U39864 ( .A1(n20207), .A2(n20205), .ZN(n20455) );
  XOR2_X1 U39867 ( .A1(n19530), .A2(n19430), .Z(n50544) );
  BUF_X2 U39868 ( .I(n46547), .Z(n19433) );
  NAND2_X1 U39870 ( .A1(n53098), .A2(n53104), .ZN(n22222) );
  NAND2_X1 U39874 ( .A1(n35340), .A2(n59809), .ZN(n34936) );
  NAND2_X1 U39875 ( .A1(n19440), .A2(n19439), .ZN(n37831) );
  NAND2_X1 U39876 ( .A1(n37830), .A2(n41054), .ZN(n19440) );
  AND2_X1 U39882 ( .A1(n33979), .A2(n34604), .Z(n19448) );
  XOR2_X1 U39883 ( .A1(n19453), .A2(n53273), .Z(Plaintext[15]) );
  NOR2_X1 U39884 ( .A1(n53201), .A2(n53199), .ZN(n20692) );
  INV_X2 U39888 ( .I(n34341), .ZN(n31976) );
  XOR2_X1 U39889 ( .A1(n31975), .A2(n15962), .Z(n34341) );
  INV_X2 U39901 ( .I(n24850), .ZN(n47181) );
  NAND2_X2 U39906 ( .A1(n19476), .A2(n19484), .ZN(n53677) );
  NOR2_X2 U39907 ( .A1(n53691), .A2(n19475), .ZN(n20631) );
  XOR2_X1 U39908 ( .A1(n32517), .A2(n33897), .Z(n19478) );
  XOR2_X1 U39909 ( .A1(n19479), .A2(n19627), .Z(n33897) );
  INV_X1 U39911 ( .I(n51379), .ZN(n19488) );
  XOR2_X1 U39912 ( .A1(n38541), .A2(n19502), .Z(n19501) );
  XOR2_X1 U39913 ( .A1(n19504), .A2(n9397), .Z(n19503) );
  XOR2_X1 U39914 ( .A1(n38727), .A2(n37175), .Z(n19504) );
  XOR2_X1 U39917 ( .A1(n19622), .A2(n779), .Z(n31765) );
  XOR2_X1 U39918 ( .A1(n19622), .A2(n1574), .Z(n32387) );
  XOR2_X1 U39919 ( .A1(n32007), .A2(n19514), .Z(n32008) );
  NOR2_X2 U39920 ( .A1(n19516), .A2(n19515), .ZN(n19622) );
  XOR2_X1 U39921 ( .A1(n36104), .A2(n19518), .Z(n36105) );
  XOR2_X1 U39924 ( .A1(n52340), .A2(n52201), .Z(n50851) );
  NAND2_X2 U39926 ( .A1(n49187), .A2(n49186), .ZN(n52201) );
  AND2_X1 U39929 ( .A1(n5939), .A2(n2160), .Z(n42692) );
  NOR2_X1 U39930 ( .A1(n34128), .A2(n19538), .ZN(n33655) );
  NAND4_X1 U39932 ( .A1(n32773), .A2(n36484), .A3(n64093), .A4(n10413), .ZN(
        n32774) );
  INV_X1 U39933 ( .I(n21097), .ZN(n19541) );
  NAND2_X2 U39935 ( .A1(n49770), .A2(n49780), .ZN(n47068) );
  NOR2_X2 U39936 ( .A1(n19544), .A2(n62700), .ZN(n49780) );
  NOR2_X2 U39938 ( .A1(n19555), .A2(n53532), .ZN(n53539) );
  INV_X1 U39941 ( .I(n24090), .ZN(n19564) );
  NAND3_X1 U39943 ( .A1(n34424), .A2(n35769), .A3(n19570), .ZN(n34425) );
  NOR2_X1 U39944 ( .A1(n31092), .A2(n24199), .ZN(n19571) );
  AND2_X1 U39945 ( .A1(n36756), .A2(n19573), .Z(n25296) );
  OAI21_X1 U39946 ( .A1(n19575), .A2(n19574), .B(n60653), .ZN(n40384) );
  AOI21_X1 U39951 ( .A1(n29635), .A2(n19581), .B(n20907), .ZN(n28146) );
  NAND3_X1 U39952 ( .A1(n10102), .A2(n26084), .A3(n19590), .ZN(n28204) );
  OAI21_X1 U39953 ( .A1(n5837), .A2(n39900), .B(n19592), .ZN(n39901) );
  XOR2_X1 U39954 ( .A1(Ciphertext[140]), .A2(Key[9]), .Z(n28589) );
  NAND2_X1 U39955 ( .A1(n19595), .A2(n64063), .ZN(n45531) );
  XOR2_X1 U39957 ( .A1(n51390), .A2(n19599), .Z(n25497) );
  XOR2_X1 U39958 ( .A1(n50750), .A2(n19600), .Z(n19599) );
  XOR2_X1 U39959 ( .A1(n19601), .A2(n22795), .Z(n19600) );
  XOR2_X1 U39960 ( .A1(n52103), .A2(n50749), .Z(n19601) );
  XOR2_X1 U39961 ( .A1(n46196), .A2(n46195), .Z(n46198) );
  XOR2_X1 U39962 ( .A1(n46196), .A2(n44752), .Z(n44753) );
  XOR2_X1 U39963 ( .A1(n19606), .A2(n50498), .Z(n38821) );
  NOR2_X2 U39964 ( .A1(n41034), .A2(n23720), .ZN(n22523) );
  INV_X1 U39968 ( .I(n39720), .ZN(n19612) );
  XOR2_X1 U39969 ( .A1(n37966), .A2(n25514), .Z(n19613) );
  NAND2_X1 U39973 ( .A1(n1782), .A2(n36483), .ZN(n19617) );
  INV_X2 U39975 ( .I(n23410), .ZN(n23746) );
  XOR2_X1 U39976 ( .A1(n19530), .A2(n54888), .Z(n51430) );
  XOR2_X1 U39977 ( .A1(n19530), .A2(n50692), .Z(n50693) );
  XOR2_X1 U39978 ( .A1(n19530), .A2(n10335), .Z(n50372) );
  INV_X1 U39979 ( .I(n34003), .ZN(n32882) );
  AND2_X1 U39980 ( .A1(n34873), .A2(n35897), .Z(n19631) );
  INV_X2 U39983 ( .I(n50230), .ZN(n19634) );
  AND2_X1 U39984 ( .A1(n29238), .A2(n29237), .Z(n19636) );
  XOR2_X1 U39985 ( .A1(n19640), .A2(n50545), .Z(n52090) );
  XOR2_X1 U39986 ( .A1(n50544), .A2(n19888), .Z(n19640) );
  XOR2_X1 U39987 ( .A1(n19389), .A2(n42626), .Z(n42627) );
  XOR2_X1 U39988 ( .A1(n44897), .A2(n19389), .Z(n43208) );
  AOI21_X1 U39989 ( .A1(n27029), .A2(n11605), .B(n28256), .ZN(n27031) );
  OAI21_X1 U39991 ( .A1(n1615), .A2(n55721), .B(n10113), .ZN(n55427) );
  NAND2_X1 U39993 ( .A1(n15817), .A2(n15748), .ZN(n45809) );
  OAI21_X1 U39994 ( .A1(n47371), .A2(n23718), .B(n15748), .ZN(n46827) );
  XOR2_X1 U39998 ( .A1(n31597), .A2(n32394), .Z(n21923) );
  NOR2_X2 U39999 ( .A1(n32695), .A2(n33654), .ZN(n33390) );
  INV_X1 U40000 ( .I(n30266), .ZN(n19665) );
  NAND2_X1 U40003 ( .A1(n41830), .A2(n19675), .ZN(n41835) );
  INV_X2 U40004 ( .I(n29322), .ZN(n28862) );
  NOR2_X2 U40005 ( .A1(n28858), .A2(n29317), .ZN(n29322) );
  XNOR2_X1 U40007 ( .A1(n38535), .A2(n35395), .ZN(n19687) );
  INV_X1 U40009 ( .I(n58822), .ZN(n19865) );
  INV_X2 U40010 ( .I(n21276), .ZN(n55909) );
  NAND2_X1 U40011 ( .A1(n25512), .A2(n58644), .ZN(n24563) );
  NOR2_X1 U40015 ( .A1(n47964), .A2(n19681), .ZN(n19706) );
  AOI21_X1 U40016 ( .A1(n28603), .A2(n19709), .B(n28602), .ZN(n24411) );
  OAI21_X2 U40017 ( .A1(n19720), .A2(n19719), .B(n19717), .ZN(n24278) );
  XOR2_X1 U40018 ( .A1(n33833), .A2(n19722), .Z(n33834) );
  INV_X1 U40019 ( .I(n32568), .ZN(n19722) );
  XOR2_X1 U40020 ( .A1(n5727), .A2(n12591), .Z(n19723) );
  XOR2_X1 U40022 ( .A1(n45047), .A2(n44906), .Z(n44908) );
  XOR2_X1 U40023 ( .A1(n23118), .A2(n21580), .Z(n21596) );
  NAND2_X1 U40026 ( .A1(n56444), .A2(n19827), .ZN(n19729) );
  AOI21_X1 U40027 ( .A1(n56509), .A2(n15238), .B(n20587), .ZN(n19730) );
  NOR2_X2 U40028 ( .A1(n19731), .A2(n61964), .ZN(n56509) );
  AOI21_X1 U40030 ( .A1(n53183), .A2(n53182), .B(n20353), .ZN(n19736) );
  NAND2_X1 U40032 ( .A1(n45576), .A2(n45992), .ZN(n47240) );
  OAI21_X1 U40034 ( .A1(n49910), .A2(n49908), .B(n13839), .ZN(n19751) );
  XOR2_X1 U40035 ( .A1(n31270), .A2(n31277), .Z(n19755) );
  NAND2_X2 U40036 ( .A1(n31155), .A2(n31156), .ZN(n31270) );
  XOR2_X1 U40037 ( .A1(n24663), .A2(n38069), .Z(n19760) );
  NAND2_X1 U40038 ( .A1(n19761), .A2(n43995), .ZN(n21799) );
  OR3_X1 U40039 ( .A1(n36920), .A2(n19764), .A3(n36924), .Z(n19763) );
  NAND2_X2 U40041 ( .A1(n29636), .A2(n6345), .ZN(n28596) );
  NAND2_X2 U40042 ( .A1(n23955), .A2(n20747), .ZN(n28207) );
  XOR2_X1 U40043 ( .A1(n19768), .A2(n46552), .Z(n19767) );
  XOR2_X1 U40044 ( .A1(n1678), .A2(n46560), .Z(n19769) );
  XOR2_X1 U40046 ( .A1(n38636), .A2(n20506), .Z(n19771) );
  AND2_X1 U40047 ( .A1(n6345), .A2(n19593), .Z(n29645) );
  XOR2_X1 U40049 ( .A1(n61506), .A2(n38370), .Z(n38371) );
  INV_X2 U40052 ( .I(n13306), .ZN(n25534) );
  NAND2_X2 U40053 ( .A1(n35882), .A2(n35173), .ZN(n35901) );
  NOR2_X1 U40057 ( .A1(n15754), .A2(n23577), .ZN(n21150) );
  OAI22_X1 U40058 ( .A1(n35970), .A2(n23577), .B1(n6606), .B2(n35971), .ZN(
        n35973) );
  OAI21_X1 U40059 ( .A1(n15754), .A2(n35964), .B(n23577), .ZN(n35968) );
  NAND3_X1 U40060 ( .A1(n17945), .A2(n17752), .A3(n9627), .ZN(n40348) );
  XOR2_X1 U40062 ( .A1(n1835), .A2(n32617), .Z(n19828) );
  NOR2_X1 U40063 ( .A1(n22042), .A2(n50426), .ZN(n48287) );
  OAI21_X1 U40064 ( .A1(n60853), .A2(n48757), .B(n50427), .ZN(n48288) );
  OAI22_X1 U40065 ( .A1(n45466), .A2(n2878), .B1(n49253), .B2(n60853), .ZN(
        n45467) );
  INV_X1 U40066 ( .I(n15435), .ZN(n53218) );
  NAND2_X1 U40068 ( .A1(n22745), .A2(n19701), .ZN(n19841) );
  NOR2_X2 U40071 ( .A1(n56128), .A2(n56127), .ZN(n56189) );
  OR2_X2 U40073 ( .A1(n25595), .A2(n25569), .Z(n34113) );
  XOR2_X1 U40074 ( .A1(n26141), .A2(n31324), .Z(n19854) );
  NOR2_X1 U40075 ( .A1(n2786), .A2(n6934), .ZN(n19856) );
  NAND2_X2 U40076 ( .A1(n20263), .A2(n20266), .ZN(n49792) );
  XOR2_X1 U40078 ( .A1(n33229), .A2(n26026), .Z(n19860) );
  AOI21_X1 U40081 ( .A1(n1285), .A2(n18109), .B(n55299), .ZN(n52919) );
  NAND2_X1 U40082 ( .A1(n49170), .A2(n19867), .ZN(n48018) );
  AOI21_X1 U40084 ( .A1(n49559), .A2(n19867), .B(n23612), .ZN(n49169) );
  OAI22_X1 U40085 ( .A1(n42), .A2(n49560), .B1(n49559), .B2(n19867), .ZN(
        n49562) );
  XOR2_X1 U40086 ( .A1(n64039), .A2(n14251), .Z(n46510) );
  AOI21_X2 U40088 ( .A1(n24088), .A2(n24264), .B(n29331), .ZN(n31254) );
  NOR2_X2 U40090 ( .A1(n41532), .A2(n42699), .ZN(n41528) );
  OR3_X1 U40092 ( .A1(n30593), .A2(n31141), .A3(n1437), .Z(n19871) );
  NAND2_X1 U40093 ( .A1(n1843), .A2(n8584), .ZN(n19872) );
  OAI22_X1 U40094 ( .A1(n31143), .A2(n847), .B1(n23918), .B2(n1437), .ZN(
        n29011) );
  NOR3_X1 U40095 ( .A1(n30374), .A2(n30588), .A3(n1437), .ZN(n30377) );
  XOR2_X1 U40096 ( .A1(n39566), .A2(n38616), .Z(n38617) );
  AND2_X1 U40097 ( .A1(n37433), .A2(n37434), .Z(n19874) );
  INV_X1 U40100 ( .I(n32564), .ZN(n19878) );
  MUX2_X1 U40102 ( .I0(n35943), .I1(n58220), .S(n22461), .Z(n35945) );
  INV_X2 U40103 ( .I(n62546), .ZN(n19882) );
  XOR2_X1 U40104 ( .A1(Key[23]), .A2(Ciphertext[142]), .Z(n19883) );
  NOR2_X1 U40105 ( .A1(n19884), .A2(n54252), .ZN(n54253) );
  XOR2_X1 U40107 ( .A1(n31461), .A2(n1822), .Z(n31973) );
  XOR2_X1 U40108 ( .A1(n61304), .A2(n19886), .Z(n32200) );
  XOR2_X1 U40109 ( .A1(n2259), .A2(n19886), .Z(n32407) );
  XOR2_X1 U40110 ( .A1(n31866), .A2(n19886), .Z(n31867) );
  NAND2_X1 U40113 ( .A1(n19893), .A2(n37424), .ZN(n37427) );
  NAND2_X1 U40116 ( .A1(n15793), .A2(n50334), .ZN(n49970) );
  NAND3_X1 U40117 ( .A1(n49980), .A2(n49979), .A3(n15793), .ZN(n49981) );
  NAND3_X2 U40118 ( .A1(n19909), .A2(n20239), .A3(n19908), .ZN(n19907) );
  AOI21_X1 U40120 ( .A1(n19953), .A2(n19910), .B(n22681), .ZN(n19952) );
  NAND2_X1 U40122 ( .A1(n19995), .A2(n19913), .ZN(n19912) );
  AOI21_X1 U40123 ( .A1(n28862), .A2(n57424), .B(n28855), .ZN(n19913) );
  XOR2_X1 U40127 ( .A1(n19927), .A2(n20288), .Z(n20289) );
  CLKBUF_X4 U40129 ( .I(n42693), .Z(n19928) );
  INV_X2 U40132 ( .I(n55497), .ZN(n55696) );
  XOR2_X1 U40136 ( .A1(n46346), .A2(n44116), .Z(n19936) );
  INV_X1 U40137 ( .I(n46161), .ZN(n44116) );
  XOR2_X1 U40138 ( .A1(n22725), .A2(n44117), .Z(n19937) );
  OAI22_X1 U40139 ( .A1(n56572), .A2(n10183), .B1(n56567), .B2(n18255), .ZN(
        n56569) );
  NAND3_X1 U40140 ( .A1(n56167), .A2(n56185), .A3(n56191), .ZN(n19941) );
  NOR2_X2 U40141 ( .A1(n39169), .A2(n39162), .ZN(n19946) );
  NOR2_X2 U40142 ( .A1(n13858), .A2(n15717), .ZN(n55878) );
  XOR2_X1 U40143 ( .A1(n15615), .A2(n38092), .Z(n38820) );
  OAI21_X1 U40144 ( .A1(n39023), .A2(n39022), .B(n63464), .ZN(n26012) );
  AND2_X1 U40145 ( .A1(n58050), .A2(n60370), .Z(n19958) );
  XOR2_X1 U40146 ( .A1(n19960), .A2(n32035), .Z(n19959) );
  INV_X1 U40147 ( .I(n28852), .ZN(n29319) );
  NOR2_X1 U40148 ( .A1(n28852), .A2(n19965), .ZN(n19964) );
  XOR2_X1 U40149 ( .A1(n20512), .A2(n26201), .Z(n19969) );
  XOR2_X1 U40150 ( .A1(n51911), .A2(n51916), .Z(n19970) );
  INV_X1 U40151 ( .I(n19995), .ZN(n27455) );
  NAND2_X1 U40154 ( .A1(n61016), .A2(n1640), .ZN(n26223) );
  NAND2_X1 U40155 ( .A1(n11058), .A2(n1640), .ZN(n48415) );
  OAI21_X1 U40156 ( .A1(n19705), .A2(n24788), .B(n1640), .ZN(n47965) );
  XOR2_X1 U40157 ( .A1(n22953), .A2(n19983), .Z(n21153) );
  XOR2_X1 U40158 ( .A1(n1760), .A2(n22953), .Z(n37385) );
  XOR2_X1 U40159 ( .A1(n2686), .A2(n44046), .Z(n19984) );
  XOR2_X1 U40161 ( .A1(n19994), .A2(n46607), .Z(n46608) );
  NOR2_X2 U40163 ( .A1(n10769), .A2(n35775), .ZN(n35325) );
  NOR2_X1 U40164 ( .A1(n11172), .A2(n25032), .ZN(n49599) );
  NOR2_X1 U40165 ( .A1(n1638), .A2(n11172), .ZN(n48998) );
  XOR2_X1 U40166 ( .A1(n61949), .A2(n38295), .Z(n38297) );
  XOR2_X1 U40168 ( .A1(n38577), .A2(n61949), .Z(n37100) );
  XOR2_X1 U40169 ( .A1(n10992), .A2(n61949), .Z(n38214) );
  NAND2_X1 U40172 ( .A1(n48960), .A2(n58856), .ZN(n48961) );
  NAND3_X1 U40173 ( .A1(n6896), .A2(n65208), .A3(n58856), .ZN(n48966) );
  XOR2_X1 U40175 ( .A1(n50611), .A2(n51508), .Z(n23970) );
  NAND3_X2 U40176 ( .A1(n20012), .A2(n20011), .A3(n20010), .ZN(n51508) );
  OAI21_X1 U40178 ( .A1(n22514), .A2(n28858), .B(n23797), .ZN(n20023) );
  OAI21_X1 U40180 ( .A1(n27749), .A2(n30021), .B(n20025), .ZN(n27751) );
  NAND3_X2 U40181 ( .A1(n20828), .A2(n21715), .A3(n21714), .ZN(n21713) );
  XOR2_X1 U40182 ( .A1(n4663), .A2(n25176), .Z(n31070) );
  XOR2_X1 U40183 ( .A1(n4663), .A2(n23096), .Z(n31986) );
  NOR2_X1 U40184 ( .A1(n21702), .A2(n20028), .ZN(n20029) );
  INV_X1 U40186 ( .I(n20031), .ZN(n47433) );
  OAI21_X1 U40187 ( .A1(n64096), .A2(n20031), .B(n43750), .ZN(n47739) );
  AOI22_X1 U40188 ( .A1(n47743), .A2(n47744), .B1(n47745), .B2(n20031), .ZN(
        n20970) );
  XOR2_X1 U40189 ( .A1(n39680), .A2(n38015), .Z(n20032) );
  NAND2_X2 U40190 ( .A1(n15237), .A2(n62421), .ZN(n26162) );
  NAND2_X1 U40191 ( .A1(n9311), .A2(n15237), .ZN(n56486) );
  NOR2_X1 U40193 ( .A1(n20034), .A2(n23578), .ZN(n28126) );
  XOR2_X1 U40196 ( .A1(n20041), .A2(n37790), .Z(n37791) );
  XOR2_X1 U40197 ( .A1(n20041), .A2(n39211), .Z(n39212) );
  XOR2_X1 U40198 ( .A1(n20041), .A2(n38239), .Z(n38240) );
  XOR2_X1 U40199 ( .A1(n39743), .A2(n20041), .Z(n37742) );
  NAND2_X1 U40200 ( .A1(n20047), .A2(n25511), .ZN(n40269) );
  XOR2_X1 U40202 ( .A1(n1520), .A2(n39291), .Z(n20056) );
  XOR2_X1 U40203 ( .A1(n39224), .A2(n38003), .Z(n20057) );
  NAND2_X2 U40205 ( .A1(n20065), .A2(n20061), .ZN(n36768) );
  INV_X2 U40207 ( .I(n47622), .ZN(n47236) );
  AOI21_X1 U40208 ( .A1(n33001), .A2(n20068), .B(n33000), .ZN(n33002) );
  NOR2_X2 U40209 ( .A1(n20473), .A2(n10598), .ZN(n29689) );
  XOR2_X1 U40210 ( .A1(n62740), .A2(n31675), .Z(n31676) );
  XOR2_X1 U40211 ( .A1(n20073), .A2(n44729), .Z(n44730) );
  XOR2_X1 U40212 ( .A1(n46494), .A2(n20073), .Z(n20481) );
  XOR2_X1 U40215 ( .A1(n30951), .A2(n30958), .Z(n20084) );
  NAND2_X1 U40217 ( .A1(n36955), .A2(n1530), .ZN(n20085) );
  AOI22_X1 U40219 ( .A1(n29714), .A2(n29713), .B1(n29712), .B2(n20627), .ZN(
        n20089) );
  XOR2_X1 U40220 ( .A1(n21083), .A2(n16310), .Z(n32304) );
  NAND4_X2 U40224 ( .A1(n921), .A2(n20108), .A3(n20107), .A4(n21863), .ZN(
        n20106) );
  XOR2_X1 U40225 ( .A1(n20116), .A2(n20114), .Z(n20127) );
  XOR2_X1 U40226 ( .A1(n22981), .A2(n861), .Z(n20115) );
  INV_X1 U40229 ( .I(n46816), .ZN(n48093) );
  XOR2_X1 U40231 ( .A1(n19381), .A2(n39336), .Z(n39339) );
  XOR2_X1 U40232 ( .A1(n39259), .A2(n19381), .Z(n38313) );
  XOR2_X1 U40233 ( .A1(n38725), .A2(n19381), .Z(n38726) );
  XOR2_X1 U40234 ( .A1(n38956), .A2(n19381), .Z(n38958) );
  NAND2_X2 U40236 ( .A1(n20125), .A2(n25252), .ZN(n56408) );
  INV_X2 U40237 ( .I(n20126), .ZN(n29381) );
  NAND2_X2 U40238 ( .A1(n20240), .A2(n25222), .ZN(n20126) );
  AOI21_X1 U40240 ( .A1(n42929), .A2(n19882), .B(n41579), .ZN(n41582) );
  INV_X2 U40241 ( .I(n20127), .ZN(n25252) );
  NOR2_X2 U40242 ( .A1(n25252), .A2(n55950), .ZN(n56593) );
  NAND3_X1 U40243 ( .A1(n20128), .A2(n56703), .A3(n20696), .ZN(n56653) );
  NOR2_X2 U40244 ( .A1(n20269), .A2(n56719), .ZN(n20128) );
  NAND2_X1 U40245 ( .A1(n48320), .A2(n24330), .ZN(n51581) );
  NAND2_X2 U40246 ( .A1(n8889), .A2(n22765), .ZN(n26834) );
  NOR2_X1 U40250 ( .A1(n11608), .A2(n11606), .ZN(n38352) );
  XOR2_X1 U40252 ( .A1(n20142), .A2(n20144), .Z(n31701) );
  XOR2_X1 U40253 ( .A1(n31699), .A2(n22986), .Z(n20142) );
  XOR2_X1 U40254 ( .A1(n20143), .A2(n22257), .Z(n31699) );
  XOR2_X1 U40256 ( .A1(n32418), .A2(n23826), .Z(n20145) );
  NAND2_X1 U40262 ( .A1(n22989), .A2(n43695), .ZN(n41495) );
  NOR2_X1 U40263 ( .A1(n36578), .A2(n36577), .ZN(n20166) );
  INV_X2 U40264 ( .I(n24222), .ZN(n42224) );
  XOR2_X1 U40265 ( .A1(n50036), .A2(n22887), .Z(n50371) );
  XOR2_X1 U40266 ( .A1(Ciphertext[105]), .A2(Key[52]), .Z(n20553) );
  NAND2_X1 U40271 ( .A1(n26835), .A2(n1570), .ZN(n26836) );
  NOR2_X1 U40272 ( .A1(n27712), .A2(n1570), .ZN(n27714) );
  OAI22_X1 U40274 ( .A1(n43142), .A2(n20685), .B1(n43141), .B2(n43892), .ZN(
        n43143) );
  XOR2_X1 U40275 ( .A1(n38175), .A2(n37685), .Z(n20193) );
  OR2_X1 U40276 ( .A1(n57390), .A2(n20982), .Z(n20201) );
  XOR2_X1 U40277 ( .A1(n22061), .A2(n39582), .Z(n20202) );
  NOR2_X1 U40278 ( .A1(n20203), .A2(n63697), .ZN(n36682) );
  NOR2_X1 U40283 ( .A1(n49256), .A2(n20204), .ZN(n48756) );
  XOR2_X1 U40285 ( .A1(n20213), .A2(n31513), .Z(n20212) );
  XOR2_X1 U40286 ( .A1(n31512), .A2(n31630), .Z(n20213) );
  NOR2_X1 U40287 ( .A1(n23805), .A2(n20240), .ZN(n29648) );
  NOR2_X1 U40288 ( .A1(n28657), .A2(n20214), .ZN(n28658) );
  NAND2_X1 U40290 ( .A1(n20736), .A2(n897), .ZN(n35798) );
  NAND3_X2 U40291 ( .A1(n20221), .A2(n20218), .A3(n20217), .ZN(n21517) );
  XOR2_X1 U40292 ( .A1(n20226), .A2(n20225), .Z(n20224) );
  XOR2_X1 U40293 ( .A1(n20230), .A2(n16322), .Z(n44272) );
  XOR2_X1 U40294 ( .A1(n20230), .A2(n16321), .Z(n45318) );
  XOR2_X1 U40297 ( .A1(n20234), .A2(n37669), .Z(n37671) );
  NAND2_X2 U40299 ( .A1(n20286), .A2(n20241), .ZN(n29659) );
  XOR2_X1 U40300 ( .A1(Ciphertext[145]), .A2(Key[140]), .Z(n28870) );
  NAND2_X2 U40301 ( .A1(n20250), .A2(n33809), .ZN(n37090) );
  NAND3_X2 U40302 ( .A1(n20253), .A2(n20252), .A3(n33809), .ZN(n20251) );
  XOR2_X1 U40303 ( .A1(n58814), .A2(n50832), .Z(n51036) );
  XOR2_X1 U40304 ( .A1(n46621), .A2(n46307), .Z(n20271) );
  XOR2_X1 U40306 ( .A1(n1519), .A2(n16213), .Z(n20272) );
  NAND2_X1 U40307 ( .A1(n44666), .A2(n44665), .ZN(n20275) );
  INV_X2 U40308 ( .I(n24390), .ZN(n53023) );
  NOR2_X2 U40310 ( .A1(n31246), .A2(n58621), .ZN(n30891) );
  INV_X1 U40312 ( .I(n20292), .ZN(n20286) );
  XOR2_X1 U40313 ( .A1(n20289), .A2(n20290), .Z(n22097) );
  XOR2_X1 U40314 ( .A1(n7370), .A2(n20291), .Z(n20290) );
  INV_X1 U40315 ( .I(n28201), .ZN(n20292) );
  NOR2_X1 U40316 ( .A1(n1363), .A2(n28872), .ZN(n28193) );
  NAND3_X1 U40317 ( .A1(n25221), .A2(n23805), .A3(n1363), .ZN(n29379) );
  XOR2_X1 U40318 ( .A1(n31344), .A2(n23950), .Z(n31810) );
  NAND2_X1 U40322 ( .A1(n20300), .A2(n53716), .ZN(n20375) );
  AOI21_X1 U40323 ( .A1(n20300), .A2(n25117), .B(n53709), .ZN(n22020) );
  XOR2_X1 U40324 ( .A1(n32470), .A2(n31461), .Z(n31654) );
  XOR2_X1 U40325 ( .A1(n20304), .A2(n20305), .Z(n50166) );
  INV_X2 U40326 ( .I(n23970), .ZN(n20304) );
  XOR2_X1 U40327 ( .A1(n20302), .A2(n2604), .Z(n20305) );
  XOR2_X1 U40328 ( .A1(n15736), .A2(n50164), .Z(n20306) );
  XOR2_X1 U40329 ( .A1(n51932), .A2(n50165), .Z(n50325) );
  XOR2_X1 U40330 ( .A1(n33879), .A2(n19388), .Z(n20357) );
  XOR2_X1 U40331 ( .A1(n24698), .A2(n19388), .Z(n31011) );
  XOR2_X1 U40332 ( .A1(n38102), .A2(n38104), .Z(n20317) );
  XOR2_X1 U40333 ( .A1(n38103), .A2(n38361), .Z(n20318) );
  NOR2_X1 U40334 ( .A1(n20319), .A2(n1457), .ZN(n53187) );
  NOR4_X2 U40336 ( .A1(n20323), .A2(n20322), .A3(n20321), .A4(n20320), .ZN(
        n21754) );
  NAND2_X1 U40338 ( .A1(n32222), .A2(n20326), .ZN(n34262) );
  XOR2_X1 U40339 ( .A1(n20328), .A2(n20950), .Z(n44479) );
  XOR2_X1 U40340 ( .A1(n1290), .A2(n20332), .Z(n50266) );
  XOR2_X1 U40341 ( .A1(n52444), .A2(n52335), .Z(n52336) );
  XOR2_X1 U40344 ( .A1(n44354), .A2(n45400), .Z(n20334) );
  INV_X4 U40346 ( .I(n20337), .ZN(n21467) );
  NAND3_X1 U40349 ( .A1(n18099), .A2(n47096), .A3(n20340), .ZN(n46799) );
  AOI21_X1 U40350 ( .A1(n48150), .A2(n64231), .B(n48147), .ZN(n20575) );
  NOR2_X1 U40353 ( .A1(n53188), .A2(n53187), .ZN(n20354) );
  OAI21_X1 U40355 ( .A1(n36292), .A2(n34457), .B(n37357), .ZN(n20360) );
  NOR2_X1 U40356 ( .A1(n20124), .A2(n37359), .ZN(n34457) );
  NOR2_X1 U40357 ( .A1(n60214), .A2(n57790), .ZN(n27920) );
  NAND2_X2 U40359 ( .A1(n20369), .A2(n20368), .ZN(n53807) );
  XOR2_X1 U40360 ( .A1(n23016), .A2(n48969), .Z(n20370) );
  INV_X2 U40362 ( .I(n47017), .ZN(n48597) );
  NAND2_X1 U40367 ( .A1(n38543), .A2(n20374), .ZN(n38597) );
  NAND2_X2 U40369 ( .A1(n25341), .A2(n491), .ZN(n29698) );
  INV_X4 U40370 ( .I(n28639), .ZN(n25341) );
  OAI21_X1 U40373 ( .A1(n53658), .A2(n23935), .B(n20381), .ZN(n53659) );
  AOI22_X1 U40374 ( .A1(n53668), .A2(n53672), .B1(n20381), .B2(n53655), .ZN(
        n53657) );
  NAND3_X1 U40379 ( .A1(n43017), .A2(n20400), .A3(n43016), .ZN(n43018) );
  NAND3_X2 U40381 ( .A1(n31149), .A2(n31151), .A3(n31150), .ZN(n20403) );
  XOR2_X1 U40383 ( .A1(n39730), .A2(n20407), .Z(n20406) );
  XOR2_X1 U40384 ( .A1(n20408), .A2(n38710), .Z(n20407) );
  XOR2_X1 U40386 ( .A1(n20412), .A2(n20410), .Z(n20409) );
  XOR2_X1 U40387 ( .A1(n23655), .A2(n38715), .Z(n20411) );
  NAND2_X2 U40390 ( .A1(n54814), .A2(n54659), .ZN(n54825) );
  NAND2_X1 U40391 ( .A1(n55837), .A2(n55878), .ZN(n20415) );
  NOR2_X1 U40392 ( .A1(n40963), .A2(n60820), .ZN(n40964) );
  XNOR2_X1 U40393 ( .A1(n39276), .A2(n38742), .ZN(n38123) );
  XOR2_X1 U40395 ( .A1(n26100), .A2(n20421), .Z(n52345) );
  XOR2_X1 U40396 ( .A1(n25888), .A2(n51607), .Z(n20421) );
  NOR3_X1 U40398 ( .A1(n45450), .A2(n15421), .A3(n47732), .ZN(n43747) );
  OAI21_X1 U40399 ( .A1(n45725), .A2(n4569), .B(n20426), .ZN(n20423) );
  XOR2_X1 U40401 ( .A1(n51320), .A2(n50492), .Z(n20430) );
  INV_X2 U40402 ( .I(n21679), .ZN(n39095) );
  NAND2_X1 U40404 ( .A1(n22684), .A2(n63926), .ZN(n48595) );
  NAND2_X2 U40406 ( .A1(n20436), .A2(n31541), .ZN(n20908) );
  NAND2_X1 U40408 ( .A1(n28310), .A2(n20437), .ZN(n27600) );
  XOR2_X1 U40410 ( .A1(n20442), .A2(n31012), .Z(n20441) );
  XOR2_X1 U40411 ( .A1(n31010), .A2(n31011), .Z(n20442) );
  OAI21_X1 U40413 ( .A1(n34041), .A2(n19512), .B(n20444), .ZN(n31530) );
  XOR2_X1 U40414 ( .A1(n1522), .A2(n39475), .Z(n36243) );
  NAND2_X1 U40415 ( .A1(n55812), .A2(n20447), .ZN(n55784) );
  NOR2_X1 U40416 ( .A1(n16342), .A2(n20447), .ZN(n55802) );
  NOR2_X1 U40417 ( .A1(n55811), .A2(n20447), .ZN(n55773) );
  INV_X2 U40419 ( .I(n20449), .ZN(n52044) );
  XOR2_X1 U40421 ( .A1(n20457), .A2(n20573), .Z(n20456) );
  NOR2_X1 U40422 ( .A1(n20466), .A2(n33918), .ZN(n33919) );
  XOR2_X1 U40425 ( .A1(n38901), .A2(n20472), .Z(n20471) );
  XOR2_X1 U40426 ( .A1(n60499), .A2(n9956), .Z(n20472) );
  INV_X1 U40427 ( .I(n20477), .ZN(n56926) );
  XOR2_X1 U40429 ( .A1(n20479), .A2(n46496), .Z(n20478) );
  XOR2_X1 U40430 ( .A1(n20481), .A2(n20480), .Z(n20479) );
  INV_X1 U40431 ( .I(n45085), .ZN(n20480) );
  XOR2_X1 U40434 ( .A1(n19303), .A2(n15729), .Z(n37893) );
  NAND2_X1 U40435 ( .A1(n22737), .A2(n35427), .ZN(n34907) );
  NAND2_X2 U40436 ( .A1(n35431), .A2(n22737), .ZN(n35426) );
  NAND2_X2 U40437 ( .A1(n21108), .A2(n21112), .ZN(n22737) );
  NAND2_X1 U40438 ( .A1(n36939), .A2(n5936), .ZN(n20504) );
  INV_X1 U40439 ( .I(n36947), .ZN(n20505) );
  INV_X1 U40440 ( .I(n38637), .ZN(n20506) );
  INV_X2 U40443 ( .I(n20513), .ZN(n47884) );
  NAND2_X2 U40446 ( .A1(n20519), .A2(n27233), .ZN(n27543) );
  OAI21_X1 U40449 ( .A1(n34519), .A2(n34518), .B(n23363), .ZN(n20520) );
  NOR2_X1 U40451 ( .A1(n53086), .A2(n20525), .ZN(n20658) );
  INV_X2 U40453 ( .I(n20528), .ZN(n38264) );
  XOR2_X1 U40454 ( .A1(Ciphertext[184]), .A2(Key[125]), .Z(n25654) );
  XOR2_X1 U40459 ( .A1(n33076), .A2(n32517), .Z(n20534) );
  INV_X2 U40462 ( .I(n49794), .ZN(n48440) );
  NAND2_X2 U40463 ( .A1(n49792), .A2(n48440), .ZN(n48434) );
  NAND3_X1 U40465 ( .A1(n24441), .A2(n24440), .A3(n20546), .ZN(n24439) );
  INV_X2 U40466 ( .I(n20553), .ZN(n23337) );
  OAI21_X1 U40467 ( .A1(n40626), .A2(n20555), .B(n40625), .ZN(n40627) );
  NAND2_X1 U40468 ( .A1(n30345), .A2(n30339), .ZN(n20557) );
  INV_X2 U40474 ( .I(n24830), .ZN(n23689) );
  XOR2_X1 U40477 ( .A1(n7034), .A2(n43673), .Z(n43674) );
  XOR2_X1 U40481 ( .A1(n20579), .A2(n50930), .Z(n20578) );
  NOR2_X1 U40482 ( .A1(n20581), .A2(n29682), .ZN(n27890) );
  NAND2_X1 U40483 ( .A1(n20581), .A2(n10473), .ZN(n26913) );
  NAND2_X1 U40484 ( .A1(n10598), .A2(n20581), .ZN(n29685) );
  NAND2_X1 U40485 ( .A1(n60603), .A2(n20581), .ZN(n28189) );
  INV_X1 U40486 ( .I(n21189), .ZN(n49890) );
  INV_X2 U40487 ( .I(n56516), .ZN(n56510) );
  NAND2_X1 U40492 ( .A1(n39037), .A2(n63174), .ZN(n39039) );
  NOR2_X1 U40493 ( .A1(n20610), .A2(n54024), .ZN(n21998) );
  NOR2_X1 U40495 ( .A1(n20613), .A2(n53549), .ZN(n49931) );
  XOR2_X1 U40496 ( .A1(n19994), .A2(n20772), .Z(n20614) );
  NAND2_X1 U40497 ( .A1(n53674), .A2(n20615), .ZN(n53682) );
  NAND2_X1 U40499 ( .A1(n34457), .A2(n59011), .ZN(n37286) );
  NAND2_X2 U40500 ( .A1(n24174), .A2(n24176), .ZN(n40776) );
  XOR2_X1 U40501 ( .A1(n38468), .A2(n11239), .Z(n38099) );
  XOR2_X1 U40504 ( .A1(n46520), .A2(n46518), .Z(n20626) );
  NOR2_X1 U40506 ( .A1(n20627), .A2(n29709), .ZN(n29711) );
  NAND2_X1 U40507 ( .A1(n16241), .A2(n20627), .ZN(n28635) );
  NOR2_X1 U40508 ( .A1(n20630), .A2(n1457), .ZN(n50477) );
  NOR2_X1 U40509 ( .A1(n20630), .A2(n58763), .ZN(n52745) );
  OAI22_X1 U40510 ( .A1(n53533), .A2(n23784), .B1(n20630), .B2(n53396), .ZN(
        n53398) );
  NOR4_X2 U40511 ( .A1(n23935), .A2(n53666), .A3(n53700), .A4(n20631), .ZN(
        n53648) );
  INV_X1 U40512 ( .I(n20882), .ZN(n20633) );
  NOR2_X1 U40515 ( .A1(n46812), .A2(n23099), .ZN(n21318) );
  BUF_X4 U40518 ( .I(n56210), .Z(n21893) );
  OR2_X1 U40519 ( .A1(n37069), .A2(n62720), .Z(n36868) );
  INV_X2 U40520 ( .I(n22945), .ZN(n29625) );
  NAND2_X2 U40521 ( .A1(n23549), .A2(n23578), .ZN(n22945) );
  BUF_X4 U40523 ( .I(n37817), .Z(n41874) );
  NOR2_X2 U40524 ( .A1(n21881), .A2(n25396), .ZN(n36864) );
  OAI21_X1 U40525 ( .A1(n20643), .A2(n41054), .B(n41877), .ZN(n41057) );
  OR2_X1 U40527 ( .A1(n40788), .A2(n20645), .Z(n37912) );
  AND2_X1 U40529 ( .A1(n36268), .A2(n36269), .Z(n20648) );
  NAND3_X1 U40530 ( .A1(n42258), .A2(n40801), .A3(n40800), .ZN(n40810) );
  NOR2_X2 U40534 ( .A1(n49498), .A2(n19175), .ZN(n48859) );
  XOR2_X1 U40537 ( .A1(n33150), .A2(n10409), .Z(n20656) );
  AND2_X1 U40538 ( .A1(n52697), .A2(n62517), .Z(n20657) );
  INV_X1 U40540 ( .I(n28176), .ZN(n27692) );
  OR3_X1 U40541 ( .A1(n19223), .A2(n28176), .A3(n29609), .Z(n28672) );
  NAND4_X1 U40542 ( .A1(n23688), .A2(n55040), .A3(n55041), .A4(n55084), .ZN(
        n55051) );
  AND3_X1 U40543 ( .A1(n1695), .A2(n12073), .A3(n40874), .Z(n25579) );
  XOR2_X1 U40546 ( .A1(n21214), .A2(n52104), .Z(n20674) );
  NOR2_X2 U40547 ( .A1(n18348), .A2(n36493), .ZN(n21058) );
  NAND2_X1 U40550 ( .A1(n1599), .A2(n53557), .ZN(n20993) );
  NAND2_X1 U40554 ( .A1(n11244), .A2(n15921), .ZN(n25304) );
  XOR2_X1 U40555 ( .A1(n20675), .A2(n50683), .Z(n22331) );
  AND2_X1 U40558 ( .A1(n29395), .A2(n29397), .Z(n20683) );
  XOR2_X1 U40561 ( .A1(n25149), .A2(n8273), .Z(n52188) );
  XOR2_X1 U40562 ( .A1(n14665), .A2(n14666), .Z(n31153) );
  INV_X2 U40564 ( .I(n32199), .ZN(n32326) );
  INV_X2 U40566 ( .I(n25298), .ZN(n47036) );
  NAND2_X1 U40568 ( .A1(n30626), .A2(n30625), .ZN(n25036) );
  NAND4_X2 U40572 ( .A1(n53202), .A2(n53203), .A3(n20692), .A4(n20691), .ZN(
        n53204) );
  NAND4_X2 U40573 ( .A1(n31475), .A2(n31474), .A3(n31473), .A4(n31472), .ZN(
        n31476) );
  XOR2_X1 U40574 ( .A1(n20693), .A2(n52202), .Z(n52203) );
  XOR2_X1 U40575 ( .A1(n46212), .A2(n46384), .Z(n20694) );
  XOR2_X1 U40576 ( .A1(n15876), .A2(n52628), .Z(n20699) );
  NOR2_X1 U40577 ( .A1(n22281), .A2(n50811), .ZN(n22280) );
  NAND3_X1 U40579 ( .A1(n59879), .A2(n54616), .A3(n54945), .ZN(n20701) );
  XOR2_X1 U40582 ( .A1(n50712), .A2(n33057), .Z(n20703) );
  INV_X1 U40583 ( .I(n21417), .ZN(n21416) );
  OAI21_X1 U40585 ( .A1(n26515), .A2(n16266), .B(n20711), .ZN(n21223) );
  AOI22_X1 U40586 ( .A1(n28399), .A2(n180), .B1(n26345), .B2(n26346), .ZN(
        n20711) );
  NAND2_X2 U40587 ( .A1(n14307), .A2(n56403), .ZN(n56404) );
  XOR2_X1 U40588 ( .A1(n22845), .A2(n62985), .Z(n51693) );
  OR2_X1 U40590 ( .A1(n35692), .A2(n20896), .Z(n35695) );
  NAND3_X1 U40592 ( .A1(n55321), .A2(n55322), .A3(n55437), .ZN(n55324) );
  XOR2_X1 U40593 ( .A1(n23078), .A2(n10043), .Z(n46123) );
  NAND2_X1 U40594 ( .A1(n54302), .A2(n54303), .ZN(n20968) );
  INV_X1 U40596 ( .I(n39924), .ZN(n22260) );
  MUX2_X1 U40597 ( .I0(n35771), .I1(n35772), .S(n1423), .Z(n35792) );
  NOR2_X1 U40598 ( .A1(n26351), .A2(n26350), .ZN(n21237) );
  BUF_X4 U40599 ( .I(n35793), .Z(n37233) );
  AOI21_X1 U40603 ( .A1(n57005), .A2(n57004), .B(n23544), .ZN(n25023) );
  NAND3_X1 U40604 ( .A1(n41546), .A2(n40876), .A3(n40879), .ZN(n21682) );
  AND2_X1 U40605 ( .A1(n36448), .A2(n36449), .Z(n20728) );
  OAI21_X1 U40607 ( .A1(n38610), .A2(n38609), .B(n38608), .ZN(n21738) );
  XOR2_X1 U40609 ( .A1(n37002), .A2(n38861), .Z(n21280) );
  NAND2_X1 U40611 ( .A1(n54305), .A2(n54304), .ZN(n20969) );
  XOR2_X1 U40612 ( .A1(n20733), .A2(n24407), .Z(n25020) );
  XOR2_X1 U40613 ( .A1(n24409), .A2(n24408), .Z(n20733) );
  NOR2_X1 U40619 ( .A1(n43294), .A2(n11986), .ZN(n20841) );
  BUF_X2 U40620 ( .I(n25224), .Z(n20742) );
  XOR2_X1 U40622 ( .A1(n32585), .A2(n32336), .Z(n32269) );
  OR2_X1 U40623 ( .A1(n20807), .A2(n23904), .Z(n22345) );
  XOR2_X1 U40624 ( .A1(n20745), .A2(n50458), .Z(n50459) );
  XOR2_X1 U40625 ( .A1(n51662), .A2(n23022), .Z(n20745) );
  NAND3_X1 U40627 ( .A1(n31173), .A2(n30858), .A3(n31177), .ZN(n24156) );
  NAND2_X1 U40633 ( .A1(n52923), .A2(n55730), .ZN(n20749) );
  INV_X1 U40634 ( .I(n52924), .ZN(n20750) );
  NOR2_X2 U40636 ( .A1(n55470), .A2(n2180), .ZN(n55740) );
  AOI21_X1 U40637 ( .A1(n22274), .A2(n56840), .B(n22415), .ZN(n22414) );
  NOR2_X1 U40643 ( .A1(n20761), .A2(n33341), .ZN(n33344) );
  XOR2_X1 U40646 ( .A1(n45270), .A2(n20919), .Z(n45813) );
  XOR2_X1 U40647 ( .A1(n20764), .A2(n44826), .Z(n43496) );
  XOR2_X1 U40648 ( .A1(n44082), .A2(n43485), .Z(n20764) );
  INV_X4 U40649 ( .I(n22002), .ZN(n43156) );
  XOR2_X1 U40651 ( .A1(n20766), .A2(n24065), .Z(Plaintext[97]) );
  XOR2_X1 U40652 ( .A1(n43977), .A2(n21800), .Z(n20767) );
  XOR2_X1 U40654 ( .A1(n46630), .A2(n20806), .Z(n21424) );
  AND2_X1 U40655 ( .A1(n54459), .A2(n24009), .Z(n54852) );
  NAND2_X1 U40656 ( .A1(n35187), .A2(n20945), .ZN(n20944) );
  NAND3_X1 U40658 ( .A1(n46640), .A2(n46639), .A3(n20773), .ZN(n46645) );
  AOI22_X1 U40659 ( .A1(n64779), .A2(n46638), .B1(n63423), .B2(n48146), .ZN(
        n20773) );
  OR2_X1 U40660 ( .A1(n20946), .A2(n19512), .Z(n22086) );
  INV_X1 U40661 ( .I(n25759), .ZN(n25758) );
  NOR2_X2 U40664 ( .A1(n17155), .A2(n55231), .ZN(n55208) );
  XOR2_X1 U40666 ( .A1(n23042), .A2(n65171), .Z(n31870) );
  AOI22_X1 U40667 ( .A1(n27827), .A2(n28497), .B1(n27828), .B2(n27829), .ZN(
        n27836) );
  XOR2_X1 U40669 ( .A1(n32391), .A2(n32390), .Z(n20776) );
  NAND3_X1 U40670 ( .A1(n55140), .A2(n55153), .A3(n8027), .ZN(n20778) );
  NOR2_X1 U40671 ( .A1(n18525), .A2(n9783), .ZN(n20779) );
  INV_X2 U40672 ( .I(n34288), .ZN(n36909) );
  AND2_X2 U40673 ( .A1(n26303), .A2(n26304), .Z(n22106) );
  NOR2_X1 U40676 ( .A1(n61335), .A2(n30778), .ZN(n28722) );
  BUF_X2 U40677 ( .I(n27283), .Z(n20782) );
  INV_X1 U40683 ( .I(n35851), .ZN(n20793) );
  NOR2_X1 U40685 ( .A1(n24345), .A2(n24344), .ZN(n24325) );
  NAND2_X1 U40689 ( .A1(n34830), .A2(n34829), .ZN(n24341) );
  NAND4_X2 U40690 ( .A1(n33923), .A2(n35773), .A3(n33922), .A4(n33921), .ZN(
        n33929) );
  XOR2_X1 U40693 ( .A1(n37570), .A2(n20803), .Z(n43720) );
  XOR2_X1 U40694 ( .A1(n39738), .A2(n22252), .Z(n20803) );
  OR2_X1 U40697 ( .A1(n43460), .A2(n26020), .Z(n42415) );
  NOR2_X1 U40698 ( .A1(n27235), .A2(n27234), .ZN(n27236) );
  XOR2_X1 U40699 ( .A1(n44909), .A2(n44910), .Z(n46713) );
  XOR2_X1 U40700 ( .A1(n30837), .A2(n30836), .Z(n31386) );
  XOR2_X1 U40701 ( .A1(Ciphertext[183]), .A2(Key[22]), .Z(n23297) );
  OR3_X1 U40702 ( .A1(n40220), .A2(n23855), .A3(n40025), .Z(n40032) );
  NAND3_X1 U40703 ( .A1(n35258), .A2(n35320), .A3(n31956), .ZN(n20815) );
  OR2_X2 U40704 ( .A1(n52383), .A2(n52381), .Z(n54952) );
  INV_X4 U40705 ( .I(n47803), .ZN(n47811) );
  NAND2_X1 U40706 ( .A1(n20816), .A2(n31278), .ZN(n31287) );
  XOR2_X1 U40707 ( .A1(n31277), .A2(n6316), .Z(n20816) );
  NAND2_X1 U40710 ( .A1(n32018), .A2(n35302), .ZN(n20819) );
  OAI22_X1 U40711 ( .A1(n41424), .A2(n64826), .B1(n38925), .B2(n20820), .ZN(
        n38930) );
  NAND2_X1 U40712 ( .A1(n34567), .A2(n21613), .ZN(n21612) );
  INV_X2 U40715 ( .I(n20826), .ZN(n25841) );
  XOR2_X1 U40716 ( .A1(n26129), .A2(n26128), .Z(n20826) );
  AND2_X1 U40717 ( .A1(n45727), .A2(n45729), .Z(n22409) );
  AOI21_X1 U40720 ( .A1(n30557), .A2(n30556), .B(n31073), .ZN(n25031) );
  XOR2_X1 U40721 ( .A1(n58841), .A2(n20834), .Z(n31584) );
  XOR2_X1 U40724 ( .A1(n32378), .A2(n32280), .Z(n20836) );
  XOR2_X1 U40725 ( .A1(n20837), .A2(n32376), .Z(n32380) );
  XOR2_X1 U40726 ( .A1(n32377), .A2(n14818), .Z(n20837) );
  XOR2_X1 U40727 ( .A1(n45120), .A2(n45119), .Z(n21101) );
  NAND2_X2 U40729 ( .A1(n28032), .A2(n22203), .ZN(n27047) );
  INV_X1 U40732 ( .I(n26181), .ZN(n46628) );
  OR2_X1 U40738 ( .A1(n40408), .A2(n41213), .Z(n38926) );
  NOR2_X1 U40739 ( .A1(n23871), .A2(n53312), .ZN(n23870) );
  INV_X2 U40744 ( .I(n41675), .ZN(n42328) );
  NAND3_X1 U40745 ( .A1(n30266), .A2(n22139), .A3(n14389), .ZN(n23002) );
  OR2_X1 U40750 ( .A1(n52770), .A2(n53588), .Z(n20869) );
  OR2_X1 U40751 ( .A1(n53552), .A2(n52973), .Z(n20870) );
  XNOR2_X1 U40752 ( .A1(n44939), .A2(n45032), .ZN(n24598) );
  NAND3_X1 U40754 ( .A1(n33624), .A2(n33534), .A3(n33375), .ZN(n32598) );
  XOR2_X1 U40755 ( .A1(n52442), .A2(n52457), .Z(n21244) );
  AND2_X1 U40756 ( .A1(n27538), .A2(n27482), .Z(n22456) );
  INV_X4 U40757 ( .I(n21169), .ZN(n52477) );
  OR2_X2 U40758 ( .A1(n15258), .A2(n24302), .Z(n41445) );
  INV_X2 U40759 ( .I(n27189), .ZN(n28106) );
  BUF_X4 U40760 ( .I(n49549), .Z(n24394) );
  INV_X2 U40761 ( .I(n25649), .ZN(n52866) );
  NAND2_X2 U40762 ( .A1(n48559), .A2(n48076), .ZN(n48557) );
  XOR2_X1 U40763 ( .A1(n21340), .A2(n21341), .Z(n21339) );
  NAND2_X1 U40766 ( .A1(n36046), .A2(n24427), .ZN(n36045) );
  INV_X2 U40772 ( .I(n28488), .ZN(n28496) );
  OAI21_X1 U40773 ( .A1(n34172), .A2(n34661), .B(n34171), .ZN(n34173) );
  NOR2_X2 U40774 ( .A1(n55209), .A2(n22683), .ZN(n55203) );
  XOR2_X1 U40775 ( .A1(Ciphertext[53]), .A2(Key[72]), .Z(n22190) );
  XOR2_X1 U40777 ( .A1(n39343), .A2(n39346), .Z(n37650) );
  AOI21_X1 U40779 ( .A1(n49490), .A2(n48857), .B(n48856), .ZN(n22654) );
  NOR2_X1 U40780 ( .A1(n28062), .A2(n28250), .ZN(n21961) );
  XOR2_X1 U40782 ( .A1(n38659), .A2(n39592), .Z(n38745) );
  AND3_X2 U40783 ( .A1(n45220), .A2(n45221), .A3(n45219), .Z(n25162) );
  BUF_X2 U40788 ( .I(n46433), .Z(n20900) );
  OAI21_X1 U40790 ( .A1(n54341), .A2(n54350), .B(n24483), .ZN(n24482) );
  NOR2_X2 U40792 ( .A1(n24047), .A2(n44944), .ZN(n47297) );
  AOI21_X1 U40795 ( .A1(n45665), .A2(n45664), .B(n45668), .ZN(n25002) );
  NAND2_X1 U40797 ( .A1(n20913), .A2(n33375), .ZN(n32601) );
  NAND2_X2 U40800 ( .A1(n54581), .A2(n18422), .ZN(n54549) );
  XOR2_X1 U40802 ( .A1(n535), .A2(n51736), .Z(n20916) );
  NAND2_X2 U40804 ( .A1(n17538), .A2(n17958), .ZN(n35297) );
  INV_X1 U40808 ( .I(n24630), .ZN(n24629) );
  XOR2_X1 U40814 ( .A1(n39237), .A2(n37811), .Z(n20932) );
  OAI22_X1 U40815 ( .A1(n25966), .A2(n50022), .B1(n50023), .B2(n50441), .ZN(
        n20935) );
  NAND2_X1 U40816 ( .A1(n20936), .A2(n48630), .ZN(n47213) );
  NAND3_X1 U40817 ( .A1(n48495), .A2(n48642), .A3(n48164), .ZN(n20936) );
  BUF_X2 U40818 ( .I(n46513), .Z(n20937) );
  XOR2_X1 U40819 ( .A1(n64794), .A2(n23042), .Z(n20940) );
  BUF_X2 U40823 ( .I(n20818), .Z(n57113) );
  AND3_X1 U40824 ( .A1(n55252), .A2(n65011), .A3(n55412), .Z(n24675) );
  NOR2_X2 U40825 ( .A1(n40664), .A2(n41182), .ZN(n41177) );
  XOR2_X1 U40826 ( .A1(n52473), .A2(n51988), .Z(n51989) );
  NOR2_X1 U40828 ( .A1(n27039), .A2(n27038), .ZN(n20947) );
  INV_X2 U40835 ( .I(n63037), .ZN(n25999) );
  XOR2_X1 U40836 ( .A1(n25628), .A2(n39584), .Z(n39604) );
  NOR2_X1 U40840 ( .A1(n57020), .A2(n57019), .ZN(n21576) );
  INV_X1 U40841 ( .I(n21331), .ZN(n39528) );
  OAI21_X1 U40843 ( .A1(n55695), .A2(n51961), .B(n20958), .ZN(n55489) );
  AOI21_X2 U40845 ( .A1(n55493), .A2(n55492), .B(n25089), .ZN(n55594) );
  INV_X2 U40847 ( .I(n20963), .ZN(n25258) );
  XOR2_X1 U40848 ( .A1(n7264), .A2(n20964), .Z(n44094) );
  XOR2_X1 U40849 ( .A1(n31311), .A2(n31310), .Z(n20964) );
  INV_X1 U40850 ( .I(n38878), .ZN(n25375) );
  OAI21_X1 U40852 ( .A1(n54268), .A2(n54280), .B(n54282), .ZN(n24515) );
  OAI21_X1 U40853 ( .A1(n1845), .A2(n64589), .B(n28788), .ZN(n28791) );
  NAND3_X2 U40856 ( .A1(n42949), .A2(n16002), .A3(n42948), .ZN(n43944) );
  INV_X2 U40857 ( .I(n20975), .ZN(n25992) );
  XOR2_X1 U40858 ( .A1(Ciphertext[34]), .A2(Key[35]), .Z(n20975) );
  XOR2_X1 U40862 ( .A1(n33898), .A2(n31935), .Z(n31937) );
  NOR2_X1 U40863 ( .A1(n21729), .A2(n49302), .ZN(n24236) );
  NOR2_X1 U40869 ( .A1(n53266), .A2(n62199), .ZN(n20980) );
  NAND2_X1 U40870 ( .A1(n36152), .A2(n7933), .ZN(n35959) );
  OAI21_X1 U40874 ( .A1(n39076), .A2(n39077), .B(n59252), .ZN(n39078) );
  INV_X1 U40875 ( .I(n34103), .ZN(n25753) );
  INV_X4 U40880 ( .I(n25874), .ZN(n40804) );
  XOR2_X1 U40881 ( .A1(n46590), .A2(n16293), .Z(n21363) );
  OR2_X1 U40883 ( .A1(n22380), .A2(n23884), .Z(n20991) );
  AND2_X1 U40884 ( .A1(n35235), .A2(n33807), .Z(n24059) );
  NAND2_X2 U40885 ( .A1(n7285), .A2(n42008), .ZN(n43087) );
  NAND4_X1 U40886 ( .A1(n53560), .A2(n20993), .A3(n53559), .A4(n54053), .ZN(
        n53569) );
  NAND3_X2 U40887 ( .A1(n39859), .A2(n39858), .A3(n39860), .ZN(n43099) );
  XOR2_X1 U40892 ( .A1(n50499), .A2(n6597), .Z(n20998) );
  NOR2_X2 U40894 ( .A1(n21005), .A2(n54094), .ZN(n24229) );
  NAND2_X2 U40896 ( .A1(n40257), .A2(n37198), .ZN(n39158) );
  INV_X1 U40898 ( .I(n28272), .ZN(n23418) );
  AOI22_X1 U40899 ( .A1(n28457), .A2(n28615), .B1(n28458), .B2(n28459), .ZN(
        n28464) );
  AND2_X1 U40901 ( .A1(n46771), .A2(n48076), .Z(n47124) );
  OR2_X1 U40903 ( .A1(n54063), .A2(n22372), .Z(n21011) );
  NOR3_X1 U40906 ( .A1(n56122), .A2(n56121), .A3(n56123), .ZN(n56126) );
  NAND2_X1 U40907 ( .A1(n26256), .A2(n28401), .ZN(n26257) );
  INV_X2 U40910 ( .I(n21021), .ZN(n24418) );
  XOR2_X1 U40911 ( .A1(Ciphertext[138]), .A2(Key[187]), .Z(n21021) );
  INV_X4 U40912 ( .I(n21362), .ZN(n49783) );
  XOR2_X1 U40915 ( .A1(n44907), .A2(n23385), .Z(n21024) );
  XOR2_X1 U40918 ( .A1(n9628), .A2(n46140), .Z(n46210) );
  OAI21_X1 U40919 ( .A1(n26744), .A2(n26747), .B(n22482), .ZN(n26746) );
  OAI21_X1 U40921 ( .A1(n16010), .A2(n61182), .B(n52134), .ZN(n21271) );
  NAND2_X1 U40924 ( .A1(n21032), .A2(n55628), .ZN(n55623) );
  NAND2_X1 U40926 ( .A1(n40803), .A2(n25365), .ZN(n40808) );
  NAND2_X1 U40929 ( .A1(n27400), .A2(n28281), .ZN(n21629) );
  INV_X1 U40931 ( .I(Key[179]), .ZN(n21721) );
  INV_X1 U40932 ( .I(Ciphertext[35]), .ZN(n24702) );
  NOR2_X1 U40933 ( .A1(n47112), .A2(n47113), .ZN(n23597) );
  NAND2_X2 U40935 ( .A1(n49109), .A2(n47347), .ZN(n49790) );
  INV_X1 U40936 ( .I(n22866), .ZN(n22276) );
  BUF_X4 U40938 ( .I(n50096), .Z(n23650) );
  NOR2_X2 U40941 ( .A1(n21346), .A2(n5250), .ZN(n33224) );
  NAND2_X2 U40943 ( .A1(n1237), .A2(n16629), .ZN(n56433) );
  OAI21_X1 U40945 ( .A1(n21419), .A2(n21418), .B(n23186), .ZN(n21417) );
  NOR2_X1 U40946 ( .A1(n47279), .A2(n45978), .ZN(n45980) );
  OAI21_X1 U40948 ( .A1(n27411), .A2(n27412), .B(n29128), .ZN(n22120) );
  NAND2_X2 U40950 ( .A1(n42666), .A2(n43254), .ZN(n42849) );
  XOR2_X1 U40951 ( .A1(n21060), .A2(n57269), .Z(n52189) );
  XNOR2_X1 U40953 ( .A1(n31236), .A2(n22470), .ZN(n21900) );
  NAND3_X1 U40954 ( .A1(n27169), .A2(n22706), .A3(n26337), .ZN(n24879) );
  OAI21_X1 U40955 ( .A1(n56478), .A2(n56479), .B(n56502), .ZN(n56480) );
  XOR2_X1 U40958 ( .A1(Ciphertext[55]), .A2(Key[86]), .Z(n21064) );
  NOR4_X2 U40959 ( .A1(n26521), .A2(n26520), .A3(n26519), .A4(n26518), .ZN(
        n26522) );
  NOR2_X2 U40960 ( .A1(n56719), .A2(n56708), .ZN(n56730) );
  INV_X1 U40962 ( .I(n56825), .ZN(n21847) );
  NOR2_X2 U40966 ( .A1(n2180), .A2(n55727), .ZN(n55463) );
  INV_X4 U40967 ( .I(n45199), .ZN(n47797) );
  AND2_X1 U40968 ( .A1(n30075), .A2(n26370), .Z(n22127) );
  NOR2_X2 U40970 ( .A1(n45596), .A2(n45595), .ZN(n47899) );
  NAND2_X2 U40972 ( .A1(n61741), .A2(n49538), .ZN(n49430) );
  NAND2_X2 U40973 ( .A1(n54860), .A2(n54640), .ZN(n55020) );
  MUX2_X1 U40974 ( .I0(n54332), .I1(n61829), .S(n54414), .Z(n54359) );
  XOR2_X1 U40975 ( .A1(n21085), .A2(n32497), .Z(n32527) );
  BUF_X4 U40976 ( .I(n53233), .Z(n22114) );
  BUF_X2 U40981 ( .I(n30450), .Z(n21095) );
  NAND2_X1 U40982 ( .A1(n1260), .A2(n60553), .ZN(n52033) );
  INV_X4 U40984 ( .I(n21099), .ZN(n55639) );
  NOR2_X2 U40985 ( .A1(n23934), .A2(n21451), .ZN(n45807) );
  NOR2_X1 U40986 ( .A1(n11789), .A2(n19307), .ZN(n55883) );
  NOR2_X1 U40989 ( .A1(n53903), .A2(n23292), .ZN(n21115) );
  AND2_X1 U40990 ( .A1(n53962), .A2(n59662), .Z(n21118) );
  NAND2_X1 U40991 ( .A1(n53953), .A2(n53995), .ZN(n21122) );
  NOR2_X2 U40993 ( .A1(n28067), .A2(n24853), .ZN(n28250) );
  NAND2_X2 U40995 ( .A1(n18975), .A2(n49548), .ZN(n21127) );
  NOR2_X1 U40996 ( .A1(n55864), .A2(n60092), .ZN(n21129) );
  NAND2_X2 U40997 ( .A1(n27185), .A2(n26360), .ZN(n27583) );
  XOR2_X1 U41000 ( .A1(n21143), .A2(n46136), .Z(n43686) );
  XOR2_X1 U41002 ( .A1(n21153), .A2(n39598), .Z(n21152) );
  XOR2_X1 U41004 ( .A1(n31836), .A2(n21157), .Z(n21156) );
  INV_X1 U41005 ( .I(n31762), .ZN(n21157) );
  OAI21_X1 U41007 ( .A1(n21160), .A2(n36108), .B(n21381), .ZN(n21163) );
  INV_X1 U41008 ( .I(n39097), .ZN(n21160) );
  NAND2_X1 U41009 ( .A1(n21163), .A2(n21161), .ZN(n21168) );
  XOR2_X1 U41012 ( .A1(n21170), .A2(n46430), .Z(n44103) );
  XOR2_X1 U41013 ( .A1(n21170), .A2(n51261), .Z(n42178) );
  XOR2_X1 U41014 ( .A1(n46428), .A2(n21170), .Z(n46429) );
  NAND2_X2 U41018 ( .A1(n13403), .A2(n37492), .ZN(n37271) );
  AOI21_X1 U41019 ( .A1(n26052), .A2(n13403), .B(n21185), .ZN(n34844) );
  NAND2_X1 U41020 ( .A1(n18496), .A2(n37268), .ZN(n21186) );
  XOR2_X1 U41021 ( .A1(n26052), .A2(n13403), .Z(n36082) );
  NAND3_X1 U41022 ( .A1(n34847), .A2(n38550), .A3(n13403), .ZN(n37490) );
  NOR3_X1 U41025 ( .A1(n33216), .A2(n33213), .A3(n2168), .ZN(n33214) );
  OAI22_X1 U41026 ( .A1(n35844), .A2(n35845), .B1(n64884), .B2(n2168), .ZN(
        n35846) );
  XOR2_X1 U41027 ( .A1(n14), .A2(n21578), .Z(n39585) );
  XOR2_X1 U41028 ( .A1(n14), .A2(n16314), .Z(n37567) );
  XOR2_X1 U41029 ( .A1(n14), .A2(n16316), .Z(n38855) );
  NAND3_X1 U41033 ( .A1(n21204), .A2(n26539), .A3(n26540), .ZN(n26541) );
  OAI22_X1 U41034 ( .A1(n28360), .A2(n21204), .B1(n22735), .B2(n28361), .ZN(
        n28363) );
  AOI21_X1 U41035 ( .A1(n1335), .A2(n14920), .B(n4322), .ZN(n40368) );
  NOR2_X1 U41036 ( .A1(n22282), .A2(n14920), .ZN(n43362) );
  NOR2_X1 U41038 ( .A1(n43358), .A2(n14920), .ZN(n42744) );
  XOR2_X1 U41041 ( .A1(n52558), .A2(n24076), .Z(n21214) );
  XOR2_X1 U41042 ( .A1(n52103), .A2(n24051), .Z(n52558) );
  INV_X2 U41043 ( .I(n21219), .ZN(n21220) );
  XOR2_X1 U41044 ( .A1(n21220), .A2(n1463), .Z(n26211) );
  XOR2_X1 U41045 ( .A1(n21220), .A2(n21668), .Z(n50762) );
  XOR2_X1 U41048 ( .A1(n1318), .A2(n25241), .Z(n27914) );
  OR2_X1 U41052 ( .A1(n41120), .A2(n473), .Z(n21229) );
  OR2_X1 U41053 ( .A1(n41384), .A2(n41120), .Z(n21230) );
  XOR2_X1 U41054 ( .A1(n51941), .A2(n7459), .Z(n50990) );
  XOR2_X1 U41055 ( .A1(n39626), .A2(n38999), .Z(n21232) );
  XOR2_X1 U41056 ( .A1(n21234), .A2(n39625), .Z(n21233) );
  NAND3_X1 U41057 ( .A1(n62886), .A2(n58815), .A3(n21235), .ZN(n57081) );
  NAND2_X1 U41058 ( .A1(n52256), .A2(n21235), .ZN(n51463) );
  NAND2_X2 U41059 ( .A1(n52861), .A2(n50601), .ZN(n21235) );
  XOR2_X1 U41060 ( .A1(n57755), .A2(n39566), .Z(n37698) );
  XOR2_X1 U41061 ( .A1(n57755), .A2(n38114), .Z(n38115) );
  XOR2_X1 U41062 ( .A1(n17597), .A2(n5778), .Z(n50614) );
  XOR2_X1 U41063 ( .A1(n51389), .A2(n52611), .Z(n52457) );
  AND3_X1 U41065 ( .A1(n46998), .A2(n46994), .A3(n47199), .Z(n21257) );
  XNOR2_X1 U41066 ( .A1(Ciphertext[59]), .A2(Key[114]), .ZN(n21264) );
  XOR2_X1 U41069 ( .A1(n46353), .A2(n51596), .Z(n23860) );
  NOR2_X2 U41071 ( .A1(n21099), .A2(n55648), .ZN(n55625) );
  NOR2_X2 U41072 ( .A1(n21271), .A2(n21270), .ZN(n55648) );
  NAND2_X2 U41074 ( .A1(n21275), .A2(n21274), .ZN(n55582) );
  XOR2_X1 U41076 ( .A1(n21280), .A2(n36371), .Z(n36649) );
  NAND2_X1 U41077 ( .A1(n21281), .A2(n28308), .ZN(n26644) );
  NAND3_X1 U41078 ( .A1(n21281), .A2(n27179), .A3(n28313), .ZN(n27604) );
  INV_X1 U41079 ( .I(n1280), .ZN(n54271) );
  INV_X1 U41080 ( .I(n54235), .ZN(n54252) );
  AOI21_X1 U41081 ( .A1(n54233), .A2(n54235), .B(n21286), .ZN(n54216) );
  NOR3_X1 U41082 ( .A1(n54259), .A2(n1280), .A3(n21288), .ZN(n21287) );
  NAND2_X1 U41085 ( .A1(n34198), .A2(n10401), .ZN(n21292) );
  NOR2_X1 U41086 ( .A1(n21293), .A2(n56008), .ZN(n21710) );
  NAND2_X1 U41087 ( .A1(n22565), .A2(n21295), .ZN(n37531) );
  NAND2_X1 U41089 ( .A1(n21298), .A2(n7532), .ZN(n21297) );
  INV_X1 U41090 ( .I(n54065), .ZN(n21298) );
  XOR2_X1 U41096 ( .A1(n21309), .A2(n21310), .Z(n21308) );
  XOR2_X1 U41098 ( .A1(n23687), .A2(n23905), .Z(n21310) );
  AOI22_X1 U41102 ( .A1(n21317), .A2(n60960), .B1(n9766), .B2(n35003), .ZN(
        n32358) );
  NAND2_X2 U41103 ( .A1(n32951), .A2(n14111), .ZN(n21317) );
  INV_X4 U41104 ( .I(n36567), .ZN(n22785) );
  XOR2_X1 U41105 ( .A1(n24223), .A2(n37696), .Z(n24224) );
  XOR2_X1 U41106 ( .A1(n21319), .A2(n21733), .Z(n21585) );
  NOR2_X2 U41107 ( .A1(n38495), .A2(n41034), .ZN(n39094) );
  INV_X2 U41108 ( .I(n23720), .ZN(n38495) );
  AOI21_X1 U41113 ( .A1(n35575), .A2(n23626), .B(n21329), .ZN(n35578) );
  AOI21_X1 U41114 ( .A1(n36039), .A2(n36040), .B(n21329), .ZN(n36042) );
  INV_X1 U41115 ( .I(n21330), .ZN(n51351) );
  NOR2_X1 U41116 ( .A1(n22229), .A2(n21330), .ZN(n56538) );
  NAND2_X1 U41118 ( .A1(n24534), .A2(n21330), .ZN(n22072) );
  XOR2_X1 U41120 ( .A1(n43409), .A2(n43408), .Z(n22702) );
  XOR2_X1 U41121 ( .A1(n7365), .A2(n1448), .Z(n43409) );
  XOR2_X1 U41123 ( .A1(n52444), .A2(n51788), .Z(n21341) );
  XOR2_X1 U41124 ( .A1(n33334), .A2(n33335), .Z(n21344) );
  XOR2_X1 U41125 ( .A1(n22561), .A2(n16271), .Z(n38847) );
  INV_X1 U41127 ( .I(n21345), .ZN(n35111) );
  NAND2_X1 U41128 ( .A1(n55650), .A2(n15700), .ZN(n55607) );
  OAI21_X1 U41130 ( .A1(n43259), .A2(n42956), .B(n21360), .ZN(n44237) );
  NOR2_X2 U41131 ( .A1(n21978), .A2(n21974), .ZN(n21362) );
  XOR2_X1 U41132 ( .A1(n21253), .A2(n24068), .Z(n21989) );
  XOR2_X1 U41133 ( .A1(n37578), .A2(n37634), .Z(n21366) );
  XOR2_X1 U41134 ( .A1(n21368), .A2(n37816), .Z(n37817) );
  NAND2_X1 U41135 ( .A1(n138), .A2(n14708), .ZN(n56925) );
  NAND3_X1 U41137 ( .A1(n50306), .A2(n62035), .A3(n21372), .ZN(n21371) );
  NOR2_X2 U41138 ( .A1(n21375), .A2(n21374), .ZN(n21377) );
  NAND2_X1 U41141 ( .A1(n28409), .A2(n28401), .ZN(n21379) );
  INV_X1 U41142 ( .I(n25566), .ZN(n21387) );
  NAND2_X2 U41144 ( .A1(n21385), .A2(n21382), .ZN(n23425) );
  MUX2_X1 U41145 ( .I0(n21384), .I1(n21383), .S(n21381), .Z(n21382) );
  INV_X2 U41147 ( .I(n25275), .ZN(n23470) );
  NAND2_X1 U41148 ( .A1(n21389), .A2(n52645), .ZN(n52646) );
  NAND2_X1 U41149 ( .A1(n21389), .A2(n7890), .ZN(n55115) );
  XOR2_X1 U41152 ( .A1(n7370), .A2(n11355), .Z(n37834) );
  INV_X2 U41153 ( .I(n21402), .ZN(n33662) );
  CLKBUF_X4 U41155 ( .I(n22925), .Z(n21403) );
  NAND3_X2 U41156 ( .A1(n55701), .A2(n55702), .A3(n55700), .ZN(n22925) );
  NAND2_X1 U41157 ( .A1(n43116), .A2(n21408), .ZN(n22645) );
  NOR2_X1 U41158 ( .A1(n29507), .A2(n11106), .ZN(n21413) );
  AOI21_X1 U41159 ( .A1(n45977), .A2(n47597), .B(n23186), .ZN(n21415) );
  NOR2_X1 U41160 ( .A1(n45980), .A2(n45979), .ZN(n21419) );
  XOR2_X1 U41161 ( .A1(n21420), .A2(n1063), .Z(n21530) );
  XOR2_X1 U41162 ( .A1(n21599), .A2(n52105), .Z(n21422) );
  NOR2_X2 U41164 ( .A1(n1416), .A2(n17615), .ZN(n36875) );
  XOR2_X1 U41166 ( .A1(n21430), .A2(n39736), .Z(n21429) );
  XOR2_X1 U41167 ( .A1(n38377), .A2(n49273), .Z(n21430) );
  NAND2_X1 U41168 ( .A1(n57136), .A2(n58277), .ZN(n21434) );
  NOR2_X1 U41170 ( .A1(n57159), .A2(n57121), .ZN(n21441) );
  NAND2_X1 U41171 ( .A1(n57130), .A2(n21443), .ZN(n21442) );
  XOR2_X1 U41172 ( .A1(n21448), .A2(n21447), .Z(n21446) );
  XOR2_X1 U41173 ( .A1(n46591), .A2(n46599), .Z(n21448) );
  NAND4_X1 U41175 ( .A1(n36444), .A2(n7705), .A3(n36442), .A4(n15038), .ZN(
        n36446) );
  NAND2_X2 U41176 ( .A1(n18496), .A2(n34841), .ZN(n37133) );
  NAND2_X1 U41179 ( .A1(n60170), .A2(n11425), .ZN(n30447) );
  OAI22_X1 U41181 ( .A1(n34736), .A2(n21464), .B1(n31976), .B2(n35297), .ZN(
        n34737) );
  XOR2_X1 U41182 ( .A1(n25351), .A2(n26144), .Z(n26143) );
  OR2_X1 U41184 ( .A1(n42677), .A2(n18858), .Z(n21469) );
  NAND3_X1 U41188 ( .A1(n30029), .A2(n22748), .A3(n21478), .ZN(n28987) );
  NAND2_X1 U41189 ( .A1(n30025), .A2(n21478), .ZN(n21659) );
  NAND3_X1 U41190 ( .A1(n29879), .A2(n29878), .A3(n21478), .ZN(n24826) );
  NAND2_X2 U41192 ( .A1(n49937), .A2(n21479), .ZN(n49980) );
  NOR2_X1 U41193 ( .A1(n61064), .A2(n22043), .ZN(n26255) );
  XOR2_X1 U41194 ( .A1(n24537), .A2(n21480), .Z(n50326) );
  XOR2_X1 U41195 ( .A1(n23173), .A2(n21481), .Z(n51991) );
  AND2_X1 U41200 ( .A1(n57470), .A2(n23836), .Z(n53236) );
  XOR2_X1 U41201 ( .A1(n45376), .A2(n21496), .Z(n21498) );
  XOR2_X1 U41202 ( .A1(n46558), .A2(n45383), .Z(n21496) );
  XOR2_X1 U41203 ( .A1(n45377), .A2(n22340), .Z(n21497) );
  NAND2_X1 U41205 ( .A1(n18661), .A2(n21506), .ZN(n38766) );
  XOR2_X1 U41206 ( .A1(Ciphertext[85]), .A2(Key[104]), .Z(n21510) );
  NAND2_X1 U41207 ( .A1(n43412), .A2(n62997), .ZN(n43413) );
  XOR2_X1 U41209 ( .A1(n17300), .A2(n44360), .Z(n21521) );
  XOR2_X1 U41210 ( .A1(n21509), .A2(n31799), .Z(n32422) );
  INV_X2 U41212 ( .I(n21530), .ZN(n47274) );
  CLKBUF_X4 U41213 ( .I(n24023), .Z(n21531) );
  NOR2_X1 U41215 ( .A1(n22544), .A2(n25792), .ZN(n54608) );
  XOR2_X1 U41218 ( .A1(n1683), .A2(n17301), .Z(n21535) );
  NAND2_X2 U41219 ( .A1(n27930), .A2(n29133), .ZN(n29141) );
  INV_X1 U41220 ( .I(n21537), .ZN(n49657) );
  NOR2_X1 U41221 ( .A1(n50302), .A2(n21537), .ZN(n50315) );
  OR2_X1 U41222 ( .A1(n26243), .A2(n36207), .Z(n21541) );
  XOR2_X1 U41223 ( .A1(n21984), .A2(n51292), .Z(n21546) );
  OAI22_X1 U41225 ( .A1(n42587), .A2(n41624), .B1(n23561), .B2(n25368), .ZN(
        n40597) );
  NAND2_X2 U41226 ( .A1(n21551), .A2(n21558), .ZN(n49779) );
  INV_X1 U41229 ( .I(n21561), .ZN(n56998) );
  OAI21_X1 U41230 ( .A1(n56999), .A2(n21561), .B(n57000), .ZN(n21572) );
  AND2_X1 U41235 ( .A1(n43990), .A2(n1495), .Z(n21566) );
  XOR2_X1 U41236 ( .A1(n46353), .A2(n21568), .Z(n46355) );
  NOR3_X1 U41237 ( .A1(n6491), .A2(n1524), .A3(n21536), .ZN(n36289) );
  INV_X2 U41241 ( .I(n21585), .ZN(n23720) );
  INV_X1 U41244 ( .I(n21588), .ZN(n30650) );
  XOR2_X1 U41248 ( .A1(n26009), .A2(n21600), .Z(n21599) );
  OR2_X1 U41249 ( .A1(n21601), .A2(n61021), .Z(n23419) );
  NOR2_X2 U41256 ( .A1(n21630), .A2(n21627), .ZN(n22181) );
  XOR2_X1 U41257 ( .A1(n19410), .A2(n52095), .Z(n38716) );
  XOR2_X1 U41259 ( .A1(n25639), .A2(n13943), .Z(n21640) );
  XOR2_X1 U41260 ( .A1(n59773), .A2(n3260), .Z(n21642) );
  NOR2_X2 U41261 ( .A1(n56541), .A2(n56539), .ZN(n21643) );
  NAND2_X1 U41262 ( .A1(n17635), .A2(n21643), .ZN(n22040) );
  NAND2_X2 U41264 ( .A1(n37287), .A2(n37286), .ZN(n37856) );
  INV_X2 U41267 ( .I(n21653), .ZN(n44944) );
  NAND2_X2 U41268 ( .A1(n44944), .A2(n24047), .ZN(n46016) );
  INV_X2 U41269 ( .I(n25979), .ZN(n32636) );
  XOR2_X1 U41271 ( .A1(n25979), .A2(n21663), .Z(n21662) );
  XOR2_X1 U41272 ( .A1(n33283), .A2(n31972), .Z(n21663) );
  NAND2_X1 U41273 ( .A1(n48199), .A2(n15757), .ZN(n48200) );
  NAND2_X1 U41275 ( .A1(n21669), .A2(n57079), .ZN(n52671) );
  NAND2_X1 U41276 ( .A1(n52849), .A2(n21669), .ZN(n52851) );
  NAND2_X2 U41277 ( .A1(n39095), .A2(n15930), .ZN(n41035) );
  XOR2_X1 U41278 ( .A1(n34809), .A2(n746), .Z(n21680) );
  INV_X1 U41279 ( .I(n47265), .ZN(n21683) );
  XOR2_X1 U41282 ( .A1(n1760), .A2(n21687), .Z(n34495) );
  INV_X1 U41283 ( .I(n21690), .ZN(n54222) );
  NAND2_X1 U41284 ( .A1(n64788), .A2(n21690), .ZN(n54223) );
  NOR2_X1 U41285 ( .A1(n54251), .A2(n21690), .ZN(n54286) );
  NAND2_X2 U41286 ( .A1(n54277), .A2(n1280), .ZN(n21690) );
  NAND2_X1 U41287 ( .A1(n35972), .A2(n35551), .ZN(n21693) );
  NOR2_X1 U41289 ( .A1(n51863), .A2(n62102), .ZN(n21697) );
  INV_X2 U41290 ( .I(n41153), .ZN(n41455) );
  NAND2_X2 U41294 ( .A1(n21795), .A2(n21796), .ZN(n30229) );
  NAND2_X2 U41295 ( .A1(n21709), .A2(n21708), .ZN(n37807) );
  NAND2_X1 U41297 ( .A1(n22874), .A2(n48549), .ZN(n21718) );
  XOR2_X1 U41298 ( .A1(n21723), .A2(n39238), .Z(n21722) );
  XOR2_X1 U41299 ( .A1(n35377), .A2(n38780), .Z(n21723) );
  OR2_X1 U41300 ( .A1(n41713), .A2(n42923), .Z(n25962) );
  XOR2_X1 U41301 ( .A1(n42923), .A2(n1269), .Z(n41606) );
  NOR2_X1 U41302 ( .A1(n23500), .A2(n9594), .ZN(n21729) );
  XOR2_X1 U41303 ( .A1(n21734), .A2(n21735), .Z(n21733) );
  XOR2_X1 U41304 ( .A1(n16449), .A2(n38892), .Z(n21735) );
  NAND2_X2 U41305 ( .A1(n21737), .A2(n49767), .ZN(n48947) );
  NAND2_X2 U41308 ( .A1(n21743), .A2(n60049), .ZN(n53410) );
  MUX2_X1 U41309 ( .I0(n52976), .I1(n53911), .S(n21743), .Z(n52982) );
  NAND2_X2 U41310 ( .A1(n53915), .A2(n23217), .ZN(n21743) );
  NAND2_X1 U41311 ( .A1(n21749), .A2(n53815), .ZN(n21748) );
  OAI21_X1 U41312 ( .A1(n53811), .A2(n9161), .B(n53828), .ZN(n21749) );
  NOR2_X1 U41314 ( .A1(n34748), .A2(n21751), .ZN(n32018) );
  NAND3_X1 U41316 ( .A1(n32020), .A2(n32019), .A3(n59676), .ZN(n32021) );
  NAND2_X1 U41319 ( .A1(n3619), .A2(n42347), .ZN(n25126) );
  NOR2_X1 U41320 ( .A1(n42868), .A2(n3619), .ZN(n42870) );
  OAI21_X1 U41321 ( .A1(n41047), .A2(n43814), .B(n19174), .ZN(n41048) );
  XOR2_X1 U41325 ( .A1(n21761), .A2(n23329), .Z(n21760) );
  XOR2_X1 U41326 ( .A1(n21762), .A2(n16449), .Z(n21761) );
  INV_X1 U41327 ( .I(n32011), .ZN(n32012) );
  NAND2_X1 U41328 ( .A1(n63691), .A2(n22596), .ZN(n30217) );
  XOR2_X1 U41331 ( .A1(n22305), .A2(n21097), .Z(n51630) );
  XOR2_X1 U41332 ( .A1(n51621), .A2(n21097), .Z(n50649) );
  INV_X1 U41334 ( .I(n21799), .ZN(n43991) );
  NAND2_X1 U41336 ( .A1(n59545), .A2(n18607), .ZN(n50290) );
  NAND2_X1 U41341 ( .A1(n22516), .A2(n21829), .ZN(n57138) );
  XNOR2_X1 U41343 ( .A1(Ciphertext[40]), .A2(Key[77]), .ZN(n21831) );
  XOR2_X1 U41344 ( .A1(n50683), .A2(n49897), .Z(n49898) );
  NAND3_X1 U41347 ( .A1(n23008), .A2(n31247), .A3(n19255), .ZN(n31248) );
  INV_X2 U41348 ( .I(n51779), .ZN(n54625) );
  NOR2_X2 U41349 ( .A1(n46366), .A2(n21841), .ZN(n49263) );
  NAND4_X2 U41350 ( .A1(n46364), .A2(n46362), .A3(n46363), .A4(n46365), .ZN(
        n21841) );
  NAND2_X2 U41351 ( .A1(n52691), .A2(n21844), .ZN(n21843) );
  NAND2_X1 U41353 ( .A1(n34337), .A2(n21849), .ZN(n21848) );
  NAND2_X2 U41354 ( .A1(n21942), .A2(n21941), .ZN(n23232) );
  INV_X1 U41356 ( .I(n56368), .ZN(n56661) );
  INV_X2 U41360 ( .I(n21866), .ZN(n33079) );
  XOR2_X1 U41361 ( .A1(n21867), .A2(n32016), .Z(n32017) );
  XOR2_X1 U41362 ( .A1(n21868), .A2(n33079), .Z(n21867) );
  XOR2_X1 U41363 ( .A1(n32059), .A2(n32008), .Z(n21869) );
  XOR2_X1 U41364 ( .A1(n21098), .A2(n39297), .Z(n39298) );
  AND3_X1 U41366 ( .A1(n49928), .A2(n49927), .A3(n21875), .Z(n22761) );
  XOR2_X1 U41369 ( .A1(n21884), .A2(n31017), .Z(n31018) );
  XOR2_X1 U41370 ( .A1(n24034), .A2(n21884), .Z(n24919) );
  XOR2_X1 U41371 ( .A1(n23706), .A2(n21884), .Z(n30536) );
  INV_X2 U41372 ( .I(n50395), .ZN(n50400) );
  NAND2_X2 U41373 ( .A1(n21066), .A2(n21893), .ZN(n56630) );
  NAND2_X1 U41374 ( .A1(n48234), .A2(n21894), .ZN(n21954) );
  OR2_X1 U41375 ( .A1(n55339), .A2(n60974), .Z(n21897) );
  OR2_X1 U41377 ( .A1(n35103), .A2(n21915), .Z(n21904) );
  OAI21_X2 U41382 ( .A1(n21931), .A2(n51865), .B(n21929), .ZN(n22626) );
  XOR2_X1 U41384 ( .A1(n23232), .A2(n38113), .Z(n38114) );
  XOR2_X1 U41385 ( .A1(n9875), .A2(n1273), .Z(n41288) );
  NOR3_X1 U41388 ( .A1(n50000), .A2(n260), .A3(n50005), .ZN(n50001) );
  MUX2_X1 U41389 ( .I0(n49128), .I1(n49129), .S(n63202), .Z(n49141) );
  XOR2_X1 U41390 ( .A1(n21531), .A2(n19220), .Z(n21952) );
  NAND2_X1 U41393 ( .A1(n24958), .A2(n14890), .ZN(n55769) );
  NOR2_X2 U41396 ( .A1(n14307), .A2(n21957), .ZN(n56248) );
  INV_X2 U41397 ( .I(n29576), .ZN(n29580) );
  NAND2_X2 U41398 ( .A1(n28372), .A2(n28371), .ZN(n29576) );
  XOR2_X1 U41399 ( .A1(Ciphertext[27]), .A2(Key[82]), .Z(n21959) );
  NOR2_X1 U41401 ( .A1(n21961), .A2(n27040), .ZN(n25548) );
  NOR2_X1 U41402 ( .A1(n27381), .A2(n24498), .ZN(n28062) );
  NOR2_X1 U41403 ( .A1(n54582), .A2(n18425), .ZN(n54564) );
  NAND2_X1 U41404 ( .A1(n54567), .A2(n18425), .ZN(n54569) );
  XOR2_X1 U41406 ( .A1(n52621), .A2(n23221), .Z(n21962) );
  XOR2_X1 U41407 ( .A1(n51931), .A2(n51484), .Z(n52621) );
  XOR2_X1 U41408 ( .A1(n5989), .A2(n23497), .Z(n45885) );
  NOR3_X1 U41409 ( .A1(n18918), .A2(n49166), .A3(n49548), .ZN(n48272) );
  XOR2_X1 U41412 ( .A1(n21968), .A2(n21967), .Z(n38003) );
  XOR2_X1 U41413 ( .A1(n37818), .A2(n38002), .Z(n21968) );
  NAND3_X2 U41414 ( .A1(n24558), .A2(n63793), .A3(n46897), .ZN(n47261) );
  XOR2_X1 U41415 ( .A1(n21987), .A2(n18964), .Z(n31003) );
  XOR2_X1 U41416 ( .A1(n21988), .A2(n21985), .Z(n21987) );
  XOR2_X1 U41417 ( .A1(n39406), .A2(n204), .Z(n38160) );
  XOR2_X1 U41418 ( .A1(n13695), .A2(n21991), .Z(n21990) );
  XOR2_X1 U41419 ( .A1(n58827), .A2(n38129), .Z(n21991) );
  NOR2_X2 U41421 ( .A1(n22006), .A2(n22003), .ZN(n22002) );
  NAND2_X2 U41422 ( .A1(n23434), .A2(n43156), .ZN(n43151) );
  OAI21_X1 U41423 ( .A1(n47582), .A2(n47270), .B(n22549), .ZN(n22012) );
  OAI21_X1 U41424 ( .A1(n53712), .A2(n22020), .B(n22018), .ZN(n22017) );
  OAI21_X1 U41425 ( .A1(n61925), .A2(n22019), .B(n63920), .ZN(n22018) );
  NOR4_X1 U41426 ( .A1(n16489), .A2(n17286), .A3(n53732), .A4(n53726), .ZN(
        n22019) );
  NAND2_X2 U41427 ( .A1(n61925), .A2(n25116), .ZN(n53721) );
  OAI21_X1 U41430 ( .A1(n56730), .A2(n56731), .B(n22025), .ZN(n56701) );
  NAND2_X1 U41431 ( .A1(n56531), .A2(n22029), .ZN(n51348) );
  XOR2_X1 U41432 ( .A1(n51308), .A2(n20723), .Z(n22032) );
  XOR2_X1 U41433 ( .A1(n51646), .A2(n22034), .Z(n22033) );
  XOR2_X1 U41434 ( .A1(n25618), .A2(n51307), .Z(n22034) );
  XOR2_X1 U41435 ( .A1(n51645), .A2(n51374), .Z(n22035) );
  XOR2_X1 U41440 ( .A1(n17902), .A2(n44159), .Z(n44160) );
  XOR2_X1 U41441 ( .A1(n10713), .A2(n17902), .Z(n43795) );
  XOR2_X1 U41442 ( .A1(n31003), .A2(n30367), .Z(n22316) );
  XOR2_X1 U41448 ( .A1(n51661), .A2(n52505), .Z(n22057) );
  XOR2_X1 U41449 ( .A1(n51653), .A2(n51660), .Z(n22058) );
  XOR2_X1 U41452 ( .A1(n38314), .A2(n57894), .Z(n22062) );
  NAND2_X1 U41453 ( .A1(n54467), .A2(n54597), .ZN(n22065) );
  INV_X2 U41454 ( .I(n35092), .ZN(n37049) );
  INV_X2 U41457 ( .I(n22069), .ZN(n23477) );
  XOR2_X1 U41458 ( .A1(n22068), .A2(n22067), .Z(n22069) );
  INV_X1 U41461 ( .I(n22079), .ZN(n41922) );
  NOR2_X2 U41463 ( .A1(n33730), .A2(n34970), .ZN(n34546) );
  XOR2_X1 U41464 ( .A1(n6216), .A2(n51512), .Z(n51646) );
  OAI21_X1 U41466 ( .A1(n42620), .A2(n22087), .B(n43548), .ZN(n43675) );
  NOR2_X2 U41467 ( .A1(n23586), .A2(n28072), .ZN(n28239) );
  INV_X4 U41469 ( .I(n22106), .ZN(n30197) );
  NAND2_X1 U41470 ( .A1(n30193), .A2(n22091), .ZN(n28684) );
  NOR2_X2 U41474 ( .A1(n41911), .A2(n41910), .ZN(n42619) );
  XOR2_X1 U41478 ( .A1(n33079), .A2(n22104), .Z(n22103) );
  INV_X2 U41481 ( .I(n22115), .ZN(n26330) );
  INV_X1 U41483 ( .I(n24336), .ZN(n22117) );
  XOR2_X1 U41484 ( .A1(n44022), .A2(n22129), .Z(n44147) );
  NOR2_X2 U41490 ( .A1(n27446), .A2(n27445), .ZN(n30722) );
  INV_X1 U41491 ( .I(n38276), .ZN(n39002) );
  XOR2_X1 U41493 ( .A1(n19125), .A2(n22152), .Z(n50688) );
  XOR2_X1 U41494 ( .A1(n52343), .A2(n22152), .Z(n52344) );
  XOR2_X1 U41495 ( .A1(n51829), .A2(n22152), .Z(n51831) );
  XOR2_X1 U41496 ( .A1(n50566), .A2(n22152), .Z(n50567) );
  AOI21_X1 U41497 ( .A1(n22154), .A2(n39068), .B(n41168), .ZN(n38696) );
  NOR2_X1 U41498 ( .A1(n22169), .A2(n36423), .ZN(n22155) );
  NAND2_X1 U41499 ( .A1(n22156), .A2(n14729), .ZN(n29037) );
  NAND2_X1 U41502 ( .A1(n22158), .A2(n29372), .ZN(n29373) );
  XOR2_X1 U41503 ( .A1(Ciphertext[163]), .A2(Key[74]), .Z(n24481) );
  NAND2_X2 U41504 ( .A1(n9550), .A2(n55170), .ZN(n55131) );
  XOR2_X1 U41505 ( .A1(n24746), .A2(n24065), .Z(n22161) );
  XOR2_X1 U41506 ( .A1(n22163), .A2(n44061), .Z(n22291) );
  XOR2_X1 U41507 ( .A1(n43623), .A2(n45428), .Z(n22163) );
  NAND2_X1 U41516 ( .A1(n1428), .A2(n22185), .ZN(n34947) );
  XOR2_X1 U41517 ( .A1(n7199), .A2(n22187), .Z(n32270) );
  INV_X2 U41518 ( .I(n23054), .ZN(n51028) );
  XOR2_X1 U41524 ( .A1(n33033), .A2(n33171), .Z(n22195) );
  XOR2_X1 U41525 ( .A1(n37686), .A2(n37687), .Z(n37688) );
  INV_X1 U41528 ( .I(n22200), .ZN(n53706) );
  XOR2_X1 U41529 ( .A1(n15410), .A2(n22202), .Z(n37678) );
  NOR2_X2 U41530 ( .A1(n35713), .A2(n24089), .ZN(n35837) );
  NAND3_X1 U41531 ( .A1(n64187), .A2(n24321), .A3(n64719), .ZN(n24320) );
  NAND2_X1 U41534 ( .A1(n23870), .A2(n52802), .ZN(n52810) );
  XOR2_X1 U41535 ( .A1(n50459), .A2(n22778), .Z(n22209) );
  INV_X4 U41536 ( .I(n25952), .ZN(n52472) );
  NOR2_X1 U41538 ( .A1(n22110), .A2(n22115), .ZN(n26321) );
  INV_X1 U41544 ( .I(Ciphertext[25]), .ZN(n24888) );
  NAND3_X1 U41545 ( .A1(n29484), .A2(n29483), .A3(n29485), .ZN(n29486) );
  XOR2_X1 U41546 ( .A1(n51418), .A2(n22219), .Z(n52348) );
  NAND2_X1 U41548 ( .A1(n53099), .A2(n22912), .ZN(n22221) );
  AND2_X1 U41551 ( .A1(n33017), .A2(n35680), .Z(n33018) );
  BUF_X2 U41552 ( .I(n34627), .Z(n22226) );
  OAI22_X1 U41557 ( .A1(n22235), .A2(n49356), .B1(n50042), .B2(n13925), .ZN(
        n49364) );
  XOR2_X1 U41559 ( .A1(n32332), .A2(n30931), .Z(n22237) );
  NAND3_X1 U41562 ( .A1(n34609), .A2(n34608), .A3(n34610), .ZN(n34612) );
  XNOR2_X1 U41563 ( .A1(n31808), .A2(n32037), .ZN(n25700) );
  INV_X2 U41564 ( .I(n22242), .ZN(n24991) );
  NOR2_X1 U41568 ( .A1(n22630), .A2(n22628), .ZN(n25644) );
  BUF_X2 U41569 ( .I(n46282), .Z(n22247) );
  NOR2_X1 U41570 ( .A1(n22249), .A2(n22248), .ZN(n38133) );
  INV_X1 U41571 ( .I(n38136), .ZN(n22249) );
  XOR2_X1 U41572 ( .A1(n30974), .A2(n22250), .Z(n30976) );
  NAND2_X2 U41573 ( .A1(n28083), .A2(n30319), .ZN(n29278) );
  INV_X2 U41575 ( .I(n29318), .ZN(n29312) );
  AND2_X1 U41577 ( .A1(n30660), .A2(n30661), .Z(n26040) );
  OR2_X2 U41579 ( .A1(n24509), .A2(n26210), .Z(n52987) );
  XOR2_X1 U41580 ( .A1(n32066), .A2(n32067), .Z(n22265) );
  XOR2_X1 U41583 ( .A1(n39213), .A2(n39212), .Z(n39216) );
  XOR2_X1 U41584 ( .A1(n38988), .A2(n38989), .Z(n39213) );
  OAI22_X1 U41586 ( .A1(n46032), .A2(n46871), .B1(n46031), .B2(n46030), .ZN(
        n46036) );
  OR2_X1 U41587 ( .A1(n42888), .A2(n64653), .Z(n22269) );
  XOR2_X1 U41588 ( .A1(n22271), .A2(n44528), .Z(n44530) );
  XOR2_X1 U41589 ( .A1(n23553), .A2(n44527), .Z(n22271) );
  INV_X1 U41590 ( .I(n52165), .ZN(n51129) );
  INV_X1 U41594 ( .I(n56522), .ZN(n24551) );
  XOR2_X1 U41600 ( .A1(n22286), .A2(n22288), .Z(n24222) );
  OAI22_X1 U41604 ( .A1(n36897), .A2(n23765), .B1(n7103), .B2(n23764), .ZN(
        n36902) );
  AND2_X1 U41605 ( .A1(n27314), .A2(n1567), .Z(n26884) );
  AOI21_X1 U41606 ( .A1(n58303), .A2(n54503), .B(n21030), .ZN(n54504) );
  NAND3_X2 U41607 ( .A1(n33735), .A2(n33734), .A3(n33736), .ZN(n33785) );
  NOR2_X2 U41608 ( .A1(n23649), .A2(n20872), .ZN(n28460) );
  NAND3_X1 U41611 ( .A1(n45531), .A2(n22905), .A3(n45530), .ZN(n45535) );
  XOR2_X1 U41612 ( .A1(n22299), .A2(n24189), .Z(n39493) );
  OAI21_X1 U41613 ( .A1(n41390), .A2(n41391), .B(n41389), .ZN(n41396) );
  NAND3_X1 U41614 ( .A1(n28131), .A2(n28129), .A3(n28130), .ZN(n28132) );
  INV_X2 U41619 ( .I(n27837), .ZN(n26074) );
  NOR2_X2 U41622 ( .A1(n30348), .A2(n29586), .ZN(n30617) );
  XOR2_X1 U41623 ( .A1(n26924), .A2(Key[135]), .Z(n29318) );
  NOR2_X1 U41625 ( .A1(n24063), .A2(n55387), .ZN(n55388) );
  BUF_X2 U41628 ( .I(n26862), .Z(n28632) );
  NOR2_X2 U41629 ( .A1(n30820), .A2(n26506), .ZN(n29927) );
  XOR2_X1 U41630 ( .A1(n32339), .A2(n32266), .Z(n26081) );
  BUF_X2 U41632 ( .I(n51606), .Z(n54815) );
  BUF_X2 U41634 ( .I(n38910), .Z(n22321) );
  NOR2_X1 U41635 ( .A1(n29428), .A2(n29062), .ZN(n22325) );
  INV_X1 U41639 ( .I(n54254), .ZN(n54227) );
  XOR2_X1 U41640 ( .A1(n22331), .A2(n1618), .Z(n52507) );
  NAND2_X2 U41641 ( .A1(n57332), .A2(n34948), .ZN(n33757) );
  XOR2_X1 U41643 ( .A1(n33889), .A2(n31362), .Z(n22334) );
  NAND3_X1 U41646 ( .A1(n42345), .A2(n41778), .A3(n41779), .ZN(n41780) );
  BUF_X2 U41647 ( .I(n46392), .Z(n22340) );
  NAND2_X2 U41649 ( .A1(n25527), .A2(n24402), .ZN(n29814) );
  XOR2_X1 U41650 ( .A1(n12153), .A2(n23618), .Z(n44757) );
  XOR2_X1 U41651 ( .A1(Key[43]), .A2(Ciphertext[90]), .Z(n22349) );
  INV_X2 U41655 ( .I(n22355), .ZN(n34355) );
  BUF_X4 U41657 ( .I(n48818), .Z(n23156) );
  XOR2_X1 U41659 ( .A1(n32387), .A2(n111), .Z(n32389) );
  NAND2_X2 U41661 ( .A1(n26092), .A2(n26558), .ZN(n28049) );
  OR2_X1 U41663 ( .A1(n56882), .A2(n56861), .Z(n22365) );
  BUF_X2 U41668 ( .I(n3888), .Z(n22372) );
  AND2_X1 U41669 ( .A1(n26477), .A2(n26476), .Z(n25453) );
  XOR2_X1 U41671 ( .A1(n54888), .A2(n53174), .Z(n22377) );
  NAND3_X2 U41672 ( .A1(n37171), .A2(n37170), .A3(n37169), .ZN(n38659) );
  XOR2_X1 U41673 ( .A1(n22383), .A2(n54735), .Z(Plaintext[81]) );
  OAI21_X1 U41674 ( .A1(n54732), .A2(n54733), .B(n54731), .ZN(n22383) );
  NOR3_X1 U41676 ( .A1(n22388), .A2(n56405), .A3(n22387), .ZN(n56406) );
  XNOR2_X1 U41681 ( .A1(n24152), .A2(n30829), .ZN(n25667) );
  INV_X2 U41683 ( .I(n51444), .ZN(n56989) );
  NOR2_X2 U41684 ( .A1(n46982), .A2(n47472), .ZN(n47465) );
  NAND2_X2 U41687 ( .A1(n22398), .A2(n22450), .ZN(n22683) );
  NAND2_X2 U41691 ( .A1(n6979), .A2(n23179), .ZN(n33820) );
  XOR2_X1 U41692 ( .A1(n50838), .A2(n50839), .Z(n22406) );
  NOR2_X2 U41695 ( .A1(n19255), .A2(n31247), .ZN(n30888) );
  AOI21_X1 U41696 ( .A1(n57025), .A2(n57026), .B(n57024), .ZN(n57027) );
  NAND4_X2 U41697 ( .A1(n34050), .A2(n34049), .A3(n34048), .A4(n34047), .ZN(
        n35071) );
  NOR2_X1 U41698 ( .A1(n56890), .A2(n56885), .ZN(n22415) );
  NOR2_X1 U41702 ( .A1(n54195), .A2(n54196), .ZN(n54200) );
  XOR2_X1 U41704 ( .A1(n22421), .A2(n50393), .Z(n50415) );
  XOR2_X1 U41705 ( .A1(n51959), .A2(n50795), .Z(n22421) );
  NOR2_X1 U41708 ( .A1(n49034), .A2(n49033), .ZN(n25937) );
  NAND2_X1 U41709 ( .A1(n58828), .A2(n55339), .ZN(n22423) );
  NAND3_X2 U41710 ( .A1(n16063), .A2(n48746), .A3(n22424), .ZN(n52192) );
  NOR2_X2 U41712 ( .A1(n35834), .A2(n33807), .ZN(n35224) );
  XOR2_X1 U41714 ( .A1(n22429), .A2(n52017), .Z(n52032) );
  XOR2_X1 U41715 ( .A1(n51086), .A2(n19349), .Z(n22666) );
  NAND3_X1 U41716 ( .A1(n45747), .A2(n3368), .A3(n19305), .ZN(n44683) );
  BUF_X2 U41717 ( .I(n56323), .Z(n22430) );
  XOR2_X1 U41718 ( .A1(n22432), .A2(n1679), .Z(n24247) );
  XOR2_X1 U41719 ( .A1(n23548), .A2(n44043), .Z(n22432) );
  XOR2_X1 U41720 ( .A1(n22433), .A2(n23547), .Z(n24161) );
  NAND2_X2 U41721 ( .A1(n43916), .A2(n61164), .ZN(n43923) );
  XOR2_X1 U41722 ( .A1(n61665), .A2(n46297), .Z(n22434) );
  CLKBUF_X1 U41725 ( .I(n52594), .Z(n22439) );
  NAND3_X1 U41726 ( .A1(n30234), .A2(n10431), .A3(n30683), .ZN(n30236) );
  AND2_X1 U41727 ( .A1(n35931), .A2(n8520), .Z(n23545) );
  NOR2_X1 U41731 ( .A1(n55302), .A2(n65283), .ZN(n22447) );
  NAND2_X1 U41732 ( .A1(n56392), .A2(n56573), .ZN(n22453) );
  BUF_X4 U41737 ( .I(n32110), .Z(n35775) );
  NAND3_X1 U41738 ( .A1(n56201), .A2(n56199), .A3(n56200), .ZN(n56203) );
  OAI21_X1 U41740 ( .A1(n50144), .A2(n25113), .B(n50305), .ZN(n50145) );
  AOI21_X1 U41742 ( .A1(n24363), .A2(n63422), .B(n1386), .ZN(n23276) );
  AOI21_X1 U41743 ( .A1(n23276), .A2(n48547), .B(n48548), .ZN(n26027) );
  OR2_X1 U41746 ( .A1(n29631), .A2(n29284), .Z(n28131) );
  NAND2_X1 U41747 ( .A1(n31604), .A2(n33685), .ZN(n31605) );
  XNOR2_X1 U41748 ( .A1(n46705), .A2(n46704), .ZN(n25958) );
  NAND2_X2 U41749 ( .A1(n24801), .A2(n47534), .ZN(n47013) );
  XOR2_X1 U41752 ( .A1(n24547), .A2(n22471), .Z(n22470) );
  OR2_X1 U41759 ( .A1(n23331), .A2(n19361), .Z(n22484) );
  INV_X4 U41761 ( .I(n56182), .ZN(n56196) );
  INV_X1 U41762 ( .I(n22846), .ZN(n50414) );
  XOR2_X1 U41766 ( .A1(n31900), .A2(n33883), .Z(n31901) );
  OAI21_X1 U41768 ( .A1(n46825), .A2(n46826), .B(n1654), .ZN(n46830) );
  NAND2_X2 U41769 ( .A1(n42854), .A2(n42853), .ZN(n44182) );
  AOI21_X1 U41771 ( .A1(n29822), .A2(n29996), .B(n29821), .ZN(n29828) );
  NAND2_X1 U41774 ( .A1(n28064), .A2(n28063), .ZN(n25774) );
  NAND2_X2 U41775 ( .A1(n24669), .A2(n56541), .ZN(n56542) );
  XOR2_X1 U41776 ( .A1(n7679), .A2(n44049), .Z(n22512) );
  XOR2_X1 U41779 ( .A1(n22515), .A2(n15888), .Z(n22937) );
  NAND3_X1 U41780 ( .A1(n40852), .A2(n64475), .A3(n40592), .ZN(n40389) );
  OR2_X1 U41781 ( .A1(n41703), .A2(n41704), .Z(n22519) );
  BUF_X4 U41786 ( .I(n53204), .Z(n53294) );
  NOR2_X2 U41788 ( .A1(n45643), .A2(n47304), .ZN(n46013) );
  NOR2_X2 U41793 ( .A1(n22809), .A2(n25118), .ZN(n40472) );
  AOI22_X1 U41794 ( .A1(n27578), .A2(n27577), .B1(n27576), .B2(n1354), .ZN(
        n27589) );
  AND3_X1 U41795 ( .A1(n55197), .A2(n1587), .A3(n55217), .Z(n55199) );
  XOR2_X1 U41799 ( .A1(n32244), .A2(n32243), .Z(n32246) );
  NAND2_X1 U41803 ( .A1(n47196), .A2(n47490), .ZN(n22534) );
  AOI22_X1 U41804 ( .A1(n35231), .A2(n35230), .B1(n35712), .B2(n15018), .ZN(
        n35232) );
  NOR2_X1 U41805 ( .A1(n52796), .A2(n52795), .ZN(n22581) );
  BUF_X4 U41806 ( .I(n50983), .Z(n56268) );
  INV_X2 U41810 ( .I(n60293), .ZN(n28943) );
  XOR2_X1 U41812 ( .A1(n23467), .A2(n17940), .Z(n51837) );
  NAND2_X1 U41820 ( .A1(n53809), .A2(n58825), .ZN(n53824) );
  XOR2_X1 U41824 ( .A1(n15714), .A2(n15725), .Z(n22558) );
  NAND3_X2 U41825 ( .A1(n25756), .A2(n16113), .A3(n22560), .ZN(n29003) );
  OAI22_X1 U41827 ( .A1(n59961), .A2(n64308), .B1(n24649), .B2(n40756), .ZN(
        n40758) );
  AND2_X1 U41829 ( .A1(n49059), .A2(n25931), .Z(n22569) );
  INV_X1 U41831 ( .I(n22839), .ZN(n22838) );
  AND2_X1 U41832 ( .A1(n40416), .A2(n40749), .Z(n39810) );
  BUF_X2 U41837 ( .I(n11472), .Z(n23780) );
  NAND2_X1 U41840 ( .A1(n28698), .A2(n24896), .ZN(n23395) );
  MUX2_X1 U41843 ( .I0(n45711), .I1(n45712), .S(n45715), .Z(n45729) );
  INV_X2 U41844 ( .I(n22589), .ZN(n52211) );
  BUF_X4 U41845 ( .I(n26387), .Z(n27841) );
  NOR2_X2 U41847 ( .A1(n28492), .A2(n28483), .ZN(n28490) );
  XOR2_X1 U41851 ( .A1(n31970), .A2(n31679), .Z(n51968) );
  XOR2_X1 U41852 ( .A1(n37691), .A2(n39635), .Z(n31970) );
  NOR3_X1 U41853 ( .A1(n7802), .A2(n23584), .A3(n35894), .ZN(n35895) );
  AND2_X1 U41855 ( .A1(n44207), .A2(n44206), .Z(n22602) );
  NAND2_X1 U41857 ( .A1(n48659), .A2(n48653), .ZN(n22605) );
  INV_X4 U41860 ( .I(n24244), .ZN(n53672) );
  AOI22_X1 U41861 ( .A1(n48055), .A2(n1468), .B1(n48292), .B2(n65135), .ZN(
        n48056) );
  AND2_X1 U41865 ( .A1(n32901), .A2(n34159), .Z(n22613) );
  NOR2_X2 U41868 ( .A1(n23303), .A2(n26431), .ZN(n28525) );
  XOR2_X1 U41869 ( .A1(Ciphertext[166]), .A2(Key[191]), .Z(n25129) );
  NOR2_X2 U41875 ( .A1(n22626), .A2(n22625), .ZN(n23486) );
  NAND2_X1 U41876 ( .A1(n54352), .A2(n54030), .ZN(n22625) );
  INV_X2 U41877 ( .I(n25828), .ZN(n52321) );
  NOR2_X2 U41881 ( .A1(n23164), .A2(n54035), .ZN(n53561) );
  NOR2_X1 U41882 ( .A1(n53405), .A2(n53406), .ZN(n22637) );
  NAND3_X1 U41883 ( .A1(n48961), .A2(n48963), .A3(n48962), .ZN(n48965) );
  AND2_X1 U41885 ( .A1(n54261), .A2(n54260), .Z(n22641) );
  NAND2_X1 U41887 ( .A1(n24838), .A2(n24835), .ZN(n27021) );
  INV_X4 U41889 ( .I(n53109), .ZN(n23595) );
  XOR2_X1 U41890 ( .A1(Ciphertext[7]), .A2(Key[134]), .Z(n24406) );
  NOR2_X1 U41891 ( .A1(n24722), .A2(n24724), .ZN(n24717) );
  BUF_X2 U41892 ( .I(n28633), .Z(n22648) );
  AND2_X1 U41894 ( .A1(n49838), .A2(n49839), .Z(n22651) );
  NAND2_X2 U41897 ( .A1(n21915), .A2(n15805), .ZN(n36001) );
  NOR2_X2 U41899 ( .A1(n28137), .A2(n28125), .ZN(n28124) );
  BUF_X4 U41902 ( .I(n51105), .Z(n56631) );
  NAND2_X1 U41906 ( .A1(n28332), .A2(n28327), .ZN(n22671) );
  XOR2_X1 U41908 ( .A1(n17060), .A2(n49414), .Z(n49415) );
  NAND2_X2 U41909 ( .A1(n9601), .A2(n25849), .ZN(n34622) );
  AND3_X1 U41910 ( .A1(n27613), .A2(n57412), .A3(n27612), .Z(n23703) );
  XOR2_X1 U41911 ( .A1(n22675), .A2(n20302), .Z(n49413) );
  AND2_X1 U41914 ( .A1(n49653), .A2(n50053), .Z(n22682) );
  INV_X2 U41915 ( .I(n34045), .ZN(n34615) );
  NOR3_X1 U41917 ( .A1(n26696), .A2(n26694), .A3(n26695), .ZN(n26702) );
  AOI22_X1 U41921 ( .A1(n43244), .A2(n43245), .B1(n43246), .B2(n43247), .ZN(
        n43248) );
  NAND2_X1 U41923 ( .A1(n65262), .A2(n43517), .ZN(n22705) );
  NOR2_X2 U41924 ( .A1(n22703), .A2(n47181), .ZN(n47550) );
  NOR2_X2 U41925 ( .A1(n47550), .A2(n47545), .ZN(n47175) );
  XOR2_X1 U41927 ( .A1(Ciphertext[96]), .A2(Key[85]), .Z(n22709) );
  NOR2_X2 U41928 ( .A1(n5980), .A2(n12735), .ZN(n41945) );
  INV_X2 U41929 ( .I(n43549), .ZN(n43415) );
  BUF_X2 U41931 ( .I(n28211), .Z(n22714) );
  NAND3_X2 U41932 ( .A1(n53320), .A2(n53345), .A3(n53351), .ZN(n53373) );
  AOI22_X1 U41933 ( .A1(n29656), .A2(n29657), .B1(n29655), .B2(n29654), .ZN(
        n29680) );
  XOR2_X1 U41934 ( .A1(n22719), .A2(n39404), .Z(n25743) );
  NOR3_X1 U41936 ( .A1(n53747), .A2(n53745), .A3(n53746), .ZN(n53750) );
  INV_X1 U41937 ( .I(n34795), .ZN(n25900) );
  NOR2_X2 U41938 ( .A1(n28872), .A2(n29671), .ZN(n29383) );
  AOI22_X1 U41941 ( .A1(n49344), .A2(n61362), .B1(n58648), .B2(n49343), .ZN(
        n49347) );
  NOR2_X1 U41942 ( .A1(n54253), .A2(n54286), .ZN(n54263) );
  OAI21_X1 U41944 ( .A1(n28123), .A2(n28124), .B(n28122), .ZN(n28134) );
  NAND2_X1 U41947 ( .A1(n40384), .A2(n40386), .ZN(n24844) );
  XOR2_X1 U41951 ( .A1(n32634), .A2(n22732), .Z(n25826) );
  XOR2_X1 U41955 ( .A1(n23152), .A2(n31292), .Z(n22734) );
  BUF_X2 U41956 ( .I(n28362), .Z(n22735) );
  XOR2_X1 U41957 ( .A1(n37472), .A2(n37471), .Z(n23329) );
  NAND2_X1 U41958 ( .A1(n47419), .A2(n47418), .ZN(n24708) );
  XOR2_X1 U41959 ( .A1(n22743), .A2(n17668), .Z(n31464) );
  XOR2_X1 U41960 ( .A1(n9636), .A2(n56849), .Z(n22743) );
  XOR2_X1 U41961 ( .A1(n39001), .A2(n22750), .Z(n39005) );
  XOR2_X1 U41962 ( .A1(n39372), .A2(n39000), .Z(n22750) );
  XOR2_X1 U41963 ( .A1(n64285), .A2(n37799), .Z(n22757) );
  NAND2_X1 U41965 ( .A1(n33543), .A2(n35614), .ZN(n32991) );
  NAND2_X2 U41966 ( .A1(n41419), .A2(n41210), .ZN(n41414) );
  XOR2_X1 U41967 ( .A1(n22763), .A2(n51959), .Z(n51618) );
  AND2_X1 U41969 ( .A1(n25672), .A2(n43368), .Z(n22767) );
  BUF_X4 U41970 ( .I(n55994), .Z(n56107) );
  NAND2_X1 U41971 ( .A1(n24726), .A2(n36346), .ZN(n24719) );
  XOR2_X1 U41973 ( .A1(n32654), .A2(n22769), .Z(n30934) );
  NOR2_X2 U41974 ( .A1(n35709), .A2(n24089), .ZN(n35842) );
  XOR2_X1 U41977 ( .A1(n111), .A2(n32592), .Z(n31647) );
  OAI22_X1 U41980 ( .A1(n56485), .A2(n56486), .B1(n56484), .B2(n15238), .ZN(
        n56487) );
  XOR2_X1 U41981 ( .A1(n50680), .A2(n23149), .Z(n22778) );
  NOR4_X2 U41982 ( .A1(n49136), .A2(n49137), .A3(n49135), .A4(n49134), .ZN(
        n22779) );
  NAND2_X2 U41983 ( .A1(n25220), .A2(n5051), .ZN(n55082) );
  NAND3_X2 U41986 ( .A1(n52835), .A2(n52834), .A3(n52833), .ZN(n52878) );
  XOR2_X1 U41987 ( .A1(n22787), .A2(n21332), .Z(n32355) );
  XNOR2_X1 U41990 ( .A1(n46585), .A2(n32507), .ZN(n24704) );
  INV_X2 U41991 ( .I(n23582), .ZN(n52358) );
  XOR2_X1 U41998 ( .A1(n22792), .A2(n52349), .Z(n52381) );
  INV_X2 U42003 ( .I(n22800), .ZN(n24389) );
  NOR2_X2 U42007 ( .A1(n40617), .A2(n40959), .ZN(n40967) );
  XOR2_X1 U42008 ( .A1(n39755), .A2(n37778), .Z(n37123) );
  XOR2_X1 U42009 ( .A1(n61944), .A2(n50985), .Z(n37778) );
  XOR2_X1 U42010 ( .A1(n22811), .A2(n43743), .Z(n43746) );
  XOR2_X1 U42011 ( .A1(n19433), .A2(n44596), .Z(n22811) );
  NAND2_X2 U42012 ( .A1(n25112), .A2(n30159), .ZN(n30691) );
  NAND2_X1 U42013 ( .A1(n30146), .A2(n30147), .ZN(n30153) );
  XOR2_X1 U42014 ( .A1(n22812), .A2(n61092), .Z(n50387) );
  XOR2_X1 U42015 ( .A1(n50688), .A2(n50372), .Z(n22812) );
  NAND2_X2 U42016 ( .A1(n11179), .A2(n61475), .ZN(n43154) );
  AND2_X1 U42018 ( .A1(n55229), .A2(n7200), .Z(n22815) );
  OAI21_X1 U42020 ( .A1(n28340), .A2(n28341), .B(n28339), .ZN(n28345) );
  NAND2_X1 U42021 ( .A1(n55155), .A2(n55154), .ZN(n22818) );
  INV_X4 U42024 ( .I(n35709), .ZN(n35713) );
  NAND2_X2 U42026 ( .A1(n35762), .A2(n35318), .ZN(n35322) );
  INV_X2 U42031 ( .I(n35295), .ZN(n34746) );
  AND2_X2 U42033 ( .A1(n26264), .A2(n23193), .Z(n27380) );
  XOR2_X1 U42034 ( .A1(n39589), .A2(n39590), .Z(n39597) );
  OAI22_X1 U42035 ( .A1(n49688), .A2(n49365), .B1(n49687), .B2(n49686), .ZN(
        n49689) );
  NOR2_X1 U42036 ( .A1(n13725), .A2(n41855), .ZN(n41861) );
  NAND3_X1 U42038 ( .A1(n32431), .A2(n32432), .A3(n15830), .ZN(n22840) );
  XOR2_X1 U42039 ( .A1(n22841), .A2(n898), .Z(n34331) );
  AND2_X1 U42040 ( .A1(n49867), .A2(n64166), .Z(n49865) );
  XOR2_X1 U42042 ( .A1(n23365), .A2(n44270), .Z(n46206) );
  XOR2_X1 U42043 ( .A1(n38372), .A2(n38540), .Z(n22848) );
  XOR2_X1 U42044 ( .A1(n43797), .A2(n43664), .Z(n44038) );
  XOR2_X1 U42048 ( .A1(n37798), .A2(n39544), .Z(n37800) );
  INV_X1 U42049 ( .I(n55205), .ZN(n22879) );
  BUF_X2 U42051 ( .I(n55821), .Z(n22860) );
  XOR2_X1 U42053 ( .A1(n61092), .A2(n11071), .Z(n52205) );
  OR2_X1 U42054 ( .A1(n54921), .A2(n54867), .Z(n25706) );
  OAI21_X1 U42057 ( .A1(n22865), .A2(n22864), .B(n22863), .ZN(n54887) );
  NAND2_X1 U42058 ( .A1(n56892), .A2(n56881), .ZN(n22866) );
  NAND2_X1 U42059 ( .A1(n49778), .A2(n22868), .ZN(n49785) );
  NOR2_X1 U42060 ( .A1(n49776), .A2(n22869), .ZN(n22868) );
  XOR2_X1 U42062 ( .A1(n46608), .A2(n46609), .Z(n22876) );
  AOI21_X1 U42064 ( .A1(n55204), .A2(n55203), .B(n22879), .ZN(n24115) );
  INV_X4 U42065 ( .I(n25004), .ZN(n24558) );
  INV_X2 U42066 ( .I(n29343), .ZN(n27508) );
  XOR2_X1 U42067 ( .A1(n51358), .A2(n23878), .Z(n22887) );
  XOR2_X1 U42069 ( .A1(n31743), .A2(n31742), .Z(n32828) );
  NAND3_X1 U42070 ( .A1(n55657), .A2(n55658), .A3(n22977), .ZN(n55663) );
  BUF_X4 U42072 ( .I(n39035), .Z(n42784) );
  XOR2_X1 U42073 ( .A1(n32636), .A2(n30035), .Z(n30045) );
  AND2_X1 U42075 ( .A1(n28494), .A2(n22721), .Z(n27827) );
  NOR2_X2 U42077 ( .A1(n1715), .A2(n1335), .ZN(n43361) );
  NAND2_X1 U42078 ( .A1(n22897), .A2(n36244), .ZN(n22896) );
  NAND2_X1 U42079 ( .A1(n35186), .A2(n35185), .ZN(n22897) );
  NAND2_X2 U42081 ( .A1(n24052), .A2(n29609), .ZN(n28175) );
  NAND2_X1 U42083 ( .A1(n54540), .A2(n15863), .ZN(n54545) );
  NOR2_X1 U42084 ( .A1(n41191), .A2(n41190), .ZN(n22907) );
  NOR2_X1 U42086 ( .A1(n24512), .A2(n52986), .ZN(n24511) );
  AND2_X1 U42087 ( .A1(n46916), .A2(n45764), .Z(n22910) );
  NOR2_X2 U42088 ( .A1(n24926), .A2(n24925), .ZN(n24924) );
  XOR2_X1 U42089 ( .A1(n22911), .A2(n20302), .Z(n50574) );
  XOR2_X1 U42090 ( .A1(n26389), .A2(Key[169]), .Z(n23630) );
  NAND4_X1 U42093 ( .A1(n41651), .A2(n41650), .A3(n8290), .A4(n43736), .ZN(
        n41654) );
  NAND2_X1 U42094 ( .A1(n54064), .A2(n24509), .ZN(n22915) );
  OAI21_X1 U42099 ( .A1(n23300), .A2(n54564), .B(n54530), .ZN(n24489) );
  INV_X2 U42100 ( .I(n22918), .ZN(n38480) );
  XOR2_X1 U42101 ( .A1(n19171), .A2(n20818), .Z(n22919) );
  NAND3_X2 U42102 ( .A1(n39046), .A2(n39045), .A3(n39044), .ZN(n39082) );
  XOR2_X1 U42103 ( .A1(n22921), .A2(n23985), .Z(n26214) );
  NOR3_X2 U42104 ( .A1(n28549), .A2(n28548), .A3(n28547), .ZN(n29192) );
  NOR2_X2 U42106 ( .A1(n18651), .A2(n35283), .ZN(n35705) );
  BUF_X2 U42107 ( .I(n46224), .Z(n22923) );
  NOR2_X2 U42108 ( .A1(n17774), .A2(n55885), .ZN(n55842) );
  NAND2_X2 U42109 ( .A1(n24455), .A2(n15730), .ZN(n55966) );
  NAND3_X1 U42110 ( .A1(n35801), .A2(n1805), .A3(n35800), .ZN(n22927) );
  AOI22_X1 U42111 ( .A1(n1897), .A2(n56089), .B1(n56058), .B2(n56059), .ZN(
        n56060) );
  NAND2_X1 U42113 ( .A1(n24080), .A2(n60298), .ZN(n22928) );
  OAI22_X1 U42116 ( .A1(n26329), .A2(n26330), .B1(n26328), .B2(n26327), .ZN(
        n22932) );
  NAND2_X2 U42118 ( .A1(n1812), .A2(n21945), .ZN(n33944) );
  NOR2_X1 U42120 ( .A1(n54762), .A2(n54721), .ZN(n54722) );
  INV_X2 U42122 ( .I(n22937), .ZN(n41831) );
  INV_X1 U42127 ( .I(n29725), .ZN(n30026) );
  AND2_X1 U42128 ( .A1(n39934), .A2(n22944), .Z(n24612) );
  NAND3_X1 U42129 ( .A1(n42498), .A2(n41269), .A3(n9954), .ZN(n22944) );
  NAND2_X2 U42130 ( .A1(n41858), .A2(n23744), .ZN(n41851) );
  INV_X2 U42132 ( .I(n51638), .ZN(n38851) );
  XOR2_X1 U42133 ( .A1(Ciphertext[168]), .A2(Key[13]), .Z(n29343) );
  AOI22_X1 U42134 ( .A1(n42380), .A2(n41971), .B1(n62264), .B2(n42692), .ZN(
        n22951) );
  NOR2_X2 U42135 ( .A1(n34316), .A2(n35816), .ZN(n35821) );
  NAND2_X1 U42136 ( .A1(n24439), .A2(n26835), .ZN(n24438) );
  NAND2_X1 U42138 ( .A1(n23436), .A2(n23435), .ZN(n55764) );
  XOR2_X1 U42139 ( .A1(n39188), .A2(n22966), .Z(n36995) );
  XOR2_X1 U42140 ( .A1(n62502), .A2(n23790), .Z(n22966) );
  OR2_X1 U42146 ( .A1(n40125), .A2(n40128), .Z(n22983) );
  NOR2_X2 U42147 ( .A1(n27813), .A2(n27810), .ZN(n28466) );
  XOR2_X1 U42149 ( .A1(n31698), .A2(n31697), .Z(n22986) );
  NOR2_X1 U42151 ( .A1(n29700), .A2(n29699), .ZN(n23909) );
  NAND2_X2 U42155 ( .A1(n55494), .A2(n20849), .ZN(n55692) );
  AOI21_X1 U42157 ( .A1(n36190), .A2(n36402), .B(n36189), .ZN(n36191) );
  INV_X2 U42158 ( .I(n24703), .ZN(n28332) );
  NAND2_X2 U42159 ( .A1(n24837), .A2(n26558), .ZN(n24703) );
  NAND2_X1 U42160 ( .A1(n28336), .A2(n28338), .ZN(n22991) );
  INV_X1 U42161 ( .I(n28337), .ZN(n22992) );
  NAND3_X2 U42162 ( .A1(n25983), .A2(n24399), .A3(n24398), .ZN(n38168) );
  AOI22_X1 U42165 ( .A1(n30650), .A2(n8640), .B1(n30647), .B2(n3086), .ZN(
        n22998) );
  NAND2_X2 U42169 ( .A1(n24117), .A2(n16978), .ZN(n55197) );
  XOR2_X1 U42172 ( .A1(n45123), .A2(n59382), .Z(n23005) );
  NOR2_X2 U42174 ( .A1(n28510), .A2(n27846), .ZN(n26835) );
  NOR2_X2 U42175 ( .A1(n28048), .A2(n26280), .ZN(n28327) );
  NOR4_X2 U42177 ( .A1(n23013), .A2(n42763), .A3(n42764), .A4(n42762), .ZN(
        n42765) );
  NOR3_X1 U42181 ( .A1(n55762), .A2(n55764), .A3(n55763), .ZN(n55767) );
  NOR2_X2 U42183 ( .A1(n11987), .A2(n1352), .ZN(n29532) );
  XOR2_X1 U42187 ( .A1(n23027), .A2(n24822), .Z(n25658) );
  XOR2_X1 U42191 ( .A1(n52352), .A2(n52351), .Z(n52586) );
  NOR2_X2 U42192 ( .A1(n53212), .A2(n53214), .ZN(n57029) );
  NOR2_X2 U42196 ( .A1(n42518), .A2(n41831), .ZN(n42522) );
  XOR2_X1 U42197 ( .A1(n51945), .A2(n51951), .Z(n23040) );
  AOI22_X1 U42198 ( .A1(n49193), .A2(n24821), .B1(n49511), .B2(n49194), .ZN(
        n24144) );
  AOI21_X1 U42199 ( .A1(n26297), .A2(n26605), .B(n26296), .ZN(n23041) );
  INV_X4 U42203 ( .I(n24353), .ZN(n52786) );
  NAND2_X1 U42204 ( .A1(n37012), .A2(n23051), .ZN(n23050) );
  INV_X1 U42205 ( .I(n27307), .ZN(n27308) );
  INV_X2 U42206 ( .I(n23052), .ZN(n25188) );
  NAND2_X2 U42207 ( .A1(n48499), .A2(n1212), .ZN(n48648) );
  CLKBUF_X8 U42211 ( .I(n30706), .Z(n23056) );
  NAND2_X1 U42213 ( .A1(n54750), .A2(n59051), .ZN(n54704) );
  NAND2_X1 U42216 ( .A1(n47322), .A2(n47321), .ZN(n23408) );
  NAND2_X1 U42219 ( .A1(n27107), .A2(n28374), .ZN(n25800) );
  OR2_X1 U42221 ( .A1(n11987), .A2(n29528), .Z(n23068) );
  INV_X1 U42222 ( .I(n25695), .ZN(n46215) );
  NAND2_X2 U42223 ( .A1(n48545), .A2(n24364), .ZN(n48554) );
  NOR3_X1 U42226 ( .A1(n27631), .A2(n28704), .A3(n59658), .ZN(n27633) );
  NOR2_X2 U42227 ( .A1(n23084), .A2(n23083), .ZN(n30395) );
  BUF_X4 U42228 ( .I(n48944), .Z(n50044) );
  XOR2_X1 U42229 ( .A1(n23087), .A2(n55196), .Z(Plaintext[104]) );
  AND2_X1 U42230 ( .A1(n55193), .A2(n55236), .Z(n23088) );
  XOR2_X1 U42235 ( .A1(n23092), .A2(n37172), .Z(n37197) );
  XOR2_X1 U42236 ( .A1(n39749), .A2(n37160), .Z(n23092) );
  NOR2_X2 U42238 ( .A1(n23275), .A2(n55437), .ZN(n55317) );
  BUF_X2 U42241 ( .I(n2408), .Z(n23095) );
  AOI22_X1 U42242 ( .A1(n59662), .A2(n53980), .B1(n53981), .B2(n53982), .ZN(
        n53988) );
  NOR2_X1 U42243 ( .A1(n54007), .A2(n53983), .ZN(n53980) );
  XOR2_X1 U42244 ( .A1(n23098), .A2(n38435), .Z(n38436) );
  XOR2_X1 U42245 ( .A1(n38818), .A2(n38434), .Z(n23098) );
  AND2_X1 U42248 ( .A1(n53373), .A2(n53333), .Z(n26236) );
  INV_X2 U42251 ( .I(n38923), .ZN(n40770) );
  BUF_X2 U42252 ( .I(n24048), .Z(n23120) );
  NAND2_X1 U42253 ( .A1(n23121), .A2(n30176), .ZN(n30179) );
  XOR2_X1 U42254 ( .A1(n23123), .A2(n54231), .Z(Plaintext[62]) );
  NAND3_X1 U42255 ( .A1(n54230), .A2(n54229), .A3(n54228), .ZN(n23123) );
  NAND2_X2 U42257 ( .A1(n31051), .A2(n60111), .ZN(n30173) );
  OAI21_X1 U42258 ( .A1(n41107), .A2(n41108), .B(n41106), .ZN(n41116) );
  XOR2_X1 U42260 ( .A1(n23375), .A2(n52332), .Z(n23128) );
  OR2_X2 U42263 ( .A1(n50399), .A2(n50406), .Z(n50397) );
  XOR2_X1 U42264 ( .A1(n46300), .A2(n23131), .Z(n46189) );
  XOR2_X1 U42265 ( .A1(n65144), .A2(n46438), .Z(n46300) );
  OAI21_X1 U42266 ( .A1(n25817), .A2(n25815), .B(n40584), .ZN(n40587) );
  OAI21_X1 U42268 ( .A1(n23134), .A2(n23133), .B(n1404), .ZN(n39046) );
  XOR2_X1 U42276 ( .A1(n23147), .A2(n37744), .Z(n25367) );
  NOR2_X1 U42277 ( .A1(n34275), .A2(n61256), .ZN(n23148) );
  OAI21_X1 U42280 ( .A1(n23151), .A2(n59476), .B(n23150), .ZN(n41593) );
  NAND2_X1 U42281 ( .A1(n42750), .A2(n43874), .ZN(n23150) );
  NAND2_X1 U42282 ( .A1(n56406), .A2(n56587), .ZN(n24319) );
  NOR2_X1 U42284 ( .A1(n25905), .A2(n57155), .ZN(n25904) );
  INV_X2 U42285 ( .I(n23155), .ZN(n25874) );
  NAND2_X1 U42286 ( .A1(n36978), .A2(n24824), .ZN(n36984) );
  NOR2_X2 U42287 ( .A1(n35691), .A2(n22723), .ZN(n33599) );
  NAND2_X2 U42291 ( .A1(n30374), .A2(n1437), .ZN(n24172) );
  NAND2_X2 U42293 ( .A1(n30786), .A2(n30771), .ZN(n29957) );
  INV_X2 U42295 ( .I(n29616), .ZN(n28172) );
  BUF_X4 U42296 ( .I(n38056), .Z(n42407) );
  XOR2_X1 U42298 ( .A1(n23182), .A2(n854), .Z(n26970) );
  XOR2_X1 U42299 ( .A1(n54143), .A2(n24109), .Z(n23182) );
  NOR2_X2 U42300 ( .A1(n42327), .A2(n15557), .ZN(n42319) );
  INV_X1 U42301 ( .I(n43061), .ZN(n43062) );
  NOR4_X2 U42302 ( .A1(n29309), .A2(n29308), .A3(n29321), .A4(n29307), .ZN(
        n29315) );
  NAND4_X1 U42303 ( .A1(n34501), .A2(n34634), .A3(n34637), .A4(n34500), .ZN(
        n34506) );
  NAND3_X2 U42304 ( .A1(n23187), .A2(n24755), .A3(n29447), .ZN(n32289) );
  XOR2_X1 U42307 ( .A1(n51991), .A2(n58824), .Z(n23192) );
  INV_X2 U42308 ( .I(n23193), .ZN(n24853) );
  XOR2_X1 U42309 ( .A1(n24854), .A2(Key[58]), .Z(n23193) );
  INV_X2 U42310 ( .I(n56522), .ZN(n56502) );
  XOR2_X1 U42311 ( .A1(n21985), .A2(n31393), .Z(n31395) );
  NOR2_X1 U42312 ( .A1(n43658), .A2(n3696), .ZN(n23195) );
  XOR2_X1 U42316 ( .A1(n46093), .A2(n23208), .Z(n23207) );
  NAND3_X2 U42318 ( .A1(n46046), .A2(n46045), .A3(n46044), .ZN(n46047) );
  INV_X2 U42320 ( .I(n54507), .ZN(n54560) );
  BUF_X2 U42321 ( .I(n28135), .Z(n23549) );
  NAND2_X1 U42322 ( .A1(n49243), .A2(n49255), .ZN(n49248) );
  INV_X4 U42324 ( .I(n54197), .ZN(n26008) );
  INV_X1 U42325 ( .I(n39805), .ZN(n24272) );
  XOR2_X1 U42326 ( .A1(Ciphertext[12]), .A2(Key[73]), .Z(n23979) );
  NOR2_X1 U42327 ( .A1(n53407), .A2(n52977), .ZN(n52973) );
  XOR2_X1 U42328 ( .A1(n23219), .A2(n23574), .Z(n31905) );
  XOR2_X1 U42329 ( .A1(n31885), .A2(n31886), .Z(n23219) );
  INV_X1 U42331 ( .I(n53823), .ZN(n53042) );
  XOR2_X1 U42332 ( .A1(n51991), .A2(n50073), .Z(n24205) );
  NAND2_X2 U42333 ( .A1(n23887), .A2(n23793), .ZN(n30706) );
  AOI22_X1 U42335 ( .A1(n27455), .A2(n10236), .B1(n65186), .B2(n27457), .ZN(
        n27458) );
  AND2_X1 U42338 ( .A1(n34655), .A2(n34662), .Z(n23227) );
  INV_X2 U42341 ( .I(n29705), .ZN(n27813) );
  NAND2_X2 U42342 ( .A1(n28472), .A2(n27823), .ZN(n29705) );
  OR3_X1 U42343 ( .A1(n49019), .A2(n23738), .A3(n5629), .Z(n48327) );
  AOI21_X1 U42346 ( .A1(n54267), .A2(n54222), .B(n23236), .ZN(n54218) );
  NAND2_X2 U42347 ( .A1(n9655), .A2(n1257), .ZN(n56952) );
  OAI22_X1 U42350 ( .A1(n53093), .A2(n53092), .B1(n53091), .B2(n53109), .ZN(
        n53099) );
  NAND2_X2 U42352 ( .A1(n23250), .A2(n24387), .ZN(n24386) );
  XOR2_X1 U42354 ( .A1(n23254), .A2(n32341), .Z(n24656) );
  INV_X1 U42357 ( .I(n15729), .ZN(n23983) );
  XOR2_X1 U42358 ( .A1(n23261), .A2(n33023), .Z(n24600) );
  XOR2_X1 U42359 ( .A1(n33029), .A2(n33840), .Z(n23261) );
  NOR2_X2 U42361 ( .A1(n4613), .A2(n12739), .ZN(n27698) );
  OR2_X2 U42364 ( .A1(n46645), .A2(n46644), .Z(n49732) );
  NAND4_X1 U42365 ( .A1(n24190), .A2(n29104), .A3(n29105), .A4(n29106), .ZN(
        n29110) );
  AND2_X1 U42366 ( .A1(n29200), .A2(n29201), .Z(n29202) );
  NAND2_X1 U42368 ( .A1(n34530), .A2(n34973), .ZN(n34534) );
  XOR2_X1 U42369 ( .A1(n23273), .A2(n24183), .Z(n24182) );
  XOR2_X1 U42374 ( .A1(n1463), .A2(n52105), .Z(n52106) );
  XOR2_X1 U42375 ( .A1(n23282), .A2(n23442), .Z(n38709) );
  XOR2_X1 U42376 ( .A1(n25277), .A2(n39208), .Z(n23282) );
  NOR2_X2 U42378 ( .A1(n34719), .A2(n34355), .ZN(n34356) );
  XOR2_X1 U42379 ( .A1(n23287), .A2(n32386), .Z(n32391) );
  NAND2_X1 U42383 ( .A1(n23290), .A2(n23289), .ZN(n53089) );
  NOR2_X1 U42386 ( .A1(n53935), .A2(n53936), .ZN(n53942) );
  OR2_X1 U42389 ( .A1(n54035), .A2(n60049), .Z(n23295) );
  BUF_X2 U42390 ( .I(n50229), .Z(n23299) );
  AND2_X1 U42392 ( .A1(n54566), .A2(n54565), .Z(n23300) );
  NAND2_X1 U42404 ( .A1(n54948), .A2(n23309), .ZN(n54954) );
  XOR2_X1 U42406 ( .A1(n23312), .A2(n50623), .Z(n52563) );
  XOR2_X1 U42415 ( .A1(n23325), .A2(n31706), .Z(n31707) );
  XOR2_X1 U42416 ( .A1(n21083), .A2(n31705), .Z(n23325) );
  NAND2_X1 U42418 ( .A1(n23327), .A2(n23326), .ZN(n24207) );
  NAND2_X1 U42419 ( .A1(n47602), .A2(n47610), .ZN(n23327) );
  XOR2_X1 U42424 ( .A1(n39696), .A2(n23335), .Z(n39817) );
  XOR2_X1 U42425 ( .A1(n39695), .A2(n39694), .Z(n23335) );
  INV_X4 U42426 ( .I(n25259), .ZN(n53688) );
  NAND2_X2 U42431 ( .A1(n23346), .A2(n49629), .ZN(n53740) );
  NAND3_X2 U42432 ( .A1(n25242), .A2(n32855), .A3(n58080), .ZN(n35394) );
  NOR2_X2 U42433 ( .A1(n48472), .A2(n22574), .ZN(n48464) );
  INV_X1 U42437 ( .I(n50074), .ZN(n50401) );
  NAND2_X1 U42450 ( .A1(n24509), .A2(n3888), .ZN(n52983) );
  XOR2_X1 U42451 ( .A1(n16048), .A2(n46713), .Z(n23385) );
  INV_X2 U42452 ( .I(n23388), .ZN(n26180) );
  XOR2_X1 U42454 ( .A1(n5779), .A2(n23390), .Z(n38413) );
  AOI21_X1 U42458 ( .A1(n60894), .A2(n29284), .B(n23398), .ZN(n29289) );
  NAND2_X1 U42459 ( .A1(n29283), .A2(n19290), .ZN(n23398) );
  NAND2_X2 U42460 ( .A1(n36602), .A2(n36601), .ZN(n37979) );
  INV_X1 U42461 ( .I(n42991), .ZN(n25551) );
  BUF_X2 U42463 ( .I(n46702), .Z(n23402) );
  XOR2_X1 U42464 ( .A1(n24827), .A2(n31335), .Z(n24829) );
  NAND4_X2 U42466 ( .A1(n44568), .A2(n44567), .A3(n44566), .A4(n44565), .ZN(
        n44569) );
  XOR2_X1 U42468 ( .A1(n37611), .A2(n37610), .Z(n37612) );
  XOR2_X1 U42470 ( .A1(n32386), .A2(n31871), .Z(n23412) );
  XOR2_X1 U42471 ( .A1(n51226), .A2(n51225), .Z(n23417) );
  NAND2_X2 U42474 ( .A1(n35178), .A2(n35605), .ZN(n36259) );
  NAND2_X1 U42479 ( .A1(n53512), .A2(n23639), .ZN(n23638) );
  OR3_X1 U42480 ( .A1(n55756), .A2(n55757), .A3(n55820), .Z(n23436) );
  OR2_X1 U42481 ( .A1(n53426), .A2(n53425), .Z(n23437) );
  NAND2_X2 U42482 ( .A1(n24209), .A2(n49109), .ZN(n49799) );
  BUF_X4 U42485 ( .I(n49043), .Z(n23707) );
  NAND2_X1 U42486 ( .A1(n49368), .A2(n49369), .ZN(n25262) );
  INV_X2 U42488 ( .I(n25288), .ZN(n56599) );
  XOR2_X1 U42491 ( .A1(n38708), .A2(n51493), .Z(n23442) );
  NAND4_X2 U42492 ( .A1(n25503), .A2(n25504), .A3(n50018), .A4(n50017), .ZN(
        n50796) );
  XNOR2_X1 U42494 ( .A1(n51433), .A2(n51434), .ZN(n23443) );
  AND2_X1 U42495 ( .A1(n27131), .A2(n23997), .Z(n26563) );
  NAND3_X1 U42498 ( .A1(n39165), .A2(n40930), .A3(n40929), .ZN(n39166) );
  AND2_X1 U42502 ( .A1(n56140), .A2(n56139), .Z(n23456) );
  OAI22_X1 U42503 ( .A1(n56137), .A2(n56136), .B1(n56135), .B2(n11716), .ZN(
        n23457) );
  XOR2_X1 U42504 ( .A1(n43774), .A2(n12262), .Z(n23458) );
  NOR2_X2 U42507 ( .A1(n24102), .A2(n36553), .ZN(n35529) );
  XOR2_X1 U42508 ( .A1(n23463), .A2(n33897), .Z(n33912) );
  NOR3_X1 U42511 ( .A1(n45467), .A2(n45468), .A3(n49257), .ZN(n24607) );
  XOR2_X1 U42512 ( .A1(n50775), .A2(n23468), .Z(n50658) );
  XOR2_X1 U42513 ( .A1(n51286), .A2(n50657), .Z(n23468) );
  NOR2_X1 U42516 ( .A1(n28581), .A2(n28582), .ZN(n28586) );
  NAND3_X1 U42519 ( .A1(n53332), .A2(n53334), .A3(n53324), .ZN(n52798) );
  XOR2_X1 U42524 ( .A1(n23490), .A2(n44176), .Z(n44181) );
  XOR2_X1 U42525 ( .A1(n44177), .A2(n44180), .Z(n23490) );
  INV_X4 U42527 ( .I(n47603), .ZN(n47604) );
  INV_X1 U42528 ( .I(n36403), .ZN(n36405) );
  AND2_X1 U42529 ( .A1(n35201), .A2(n35624), .Z(n35622) );
  NAND3_X1 U42530 ( .A1(n33976), .A2(n34615), .A3(n23506), .ZN(n33983) );
  XOR2_X1 U42531 ( .A1(n44420), .A2(n24915), .Z(n23509) );
  XOR2_X1 U42532 ( .A1(n23510), .A2(n39743), .Z(n38452) );
  XOR2_X1 U42533 ( .A1(n38742), .A2(n38451), .Z(n23510) );
  XOR2_X1 U42534 ( .A1(Ciphertext[143]), .A2(Key[126]), .Z(n25054) );
  AOI22_X1 U42536 ( .A1(n54955), .A2(n54954), .B1(n54953), .B2(n22544), .ZN(
        n54959) );
  XOR2_X1 U42539 ( .A1(n39403), .A2(n23517), .Z(n39289) );
  XOR2_X1 U42540 ( .A1(n39285), .A2(n39277), .Z(n23517) );
  OAI21_X1 U42541 ( .A1(n4399), .A2(n14103), .B(n14446), .ZN(n52972) );
  AOI22_X1 U42542 ( .A1(n24515), .A2(n54227), .B1(n54276), .B2(n54226), .ZN(
        n54228) );
  INV_X1 U42543 ( .I(n23519), .ZN(n55636) );
  NAND2_X1 U42545 ( .A1(n55625), .A2(n15700), .ZN(n23520) );
  XOR2_X1 U42547 ( .A1(n32408), .A2(n32407), .Z(n23525) );
  AOI22_X1 U42548 ( .A1(n30104), .A2(n31039), .B1(n30135), .B2(n30103), .ZN(
        n30106) );
  AND2_X1 U42549 ( .A1(n54906), .A2(n54907), .Z(n23531) );
  XOR2_X1 U42552 ( .A1(n31448), .A2(n31732), .Z(n31450) );
  AOI21_X2 U42554 ( .A1(n30317), .A2(n30318), .B(n23537), .ZN(n24671) );
  BUF_X2 U42559 ( .I(n27822), .Z(n23540) );
  XOR2_X1 U42560 ( .A1(n24162), .A2(n44044), .Z(n23547) );
  NAND2_X2 U42561 ( .A1(n56092), .A2(n56071), .ZN(n56088) );
  XOR2_X1 U42562 ( .A1(Ciphertext[109]), .A2(Key[80]), .Z(n26091) );
  AND3_X1 U42563 ( .A1(n21268), .A2(n5277), .A3(n55275), .Z(n24526) );
  NAND2_X2 U42564 ( .A1(n9140), .A2(n48614), .ZN(n48219) );
  OR2_X2 U42565 ( .A1(n32853), .A2(n32854), .Z(n36020) );
  NOR2_X2 U42566 ( .A1(n10022), .A2(n39146), .ZN(n40490) );
  XOR2_X1 U42569 ( .A1(n45400), .A2(n45398), .Z(n23559) );
  XOR2_X1 U42572 ( .A1(n38859), .A2(n38593), .Z(n37462) );
  NAND2_X1 U42573 ( .A1(n55755), .A2(n23713), .ZN(n23712) );
  INV_X2 U42576 ( .I(n50594), .ZN(n57073) );
  INV_X4 U42577 ( .I(n40394), .ZN(n40591) );
  XOR2_X1 U42578 ( .A1(n31894), .A2(n31893), .Z(n23574) );
  NAND2_X2 U42581 ( .A1(n40547), .A2(n42670), .ZN(n42660) );
  NAND2_X2 U42583 ( .A1(n29353), .A2(n27507), .ZN(n26979) );
  INV_X2 U42584 ( .I(n23579), .ZN(n45402) );
  INV_X4 U42585 ( .I(n30419), .ZN(n24504) );
  NOR2_X2 U42586 ( .A1(n1433), .A2(n30817), .ZN(n30820) );
  INV_X2 U42587 ( .I(n37112), .ZN(n37352) );
  XOR2_X1 U42588 ( .A1(n52090), .A2(n52089), .Z(n52091) );
  INV_X4 U42589 ( .I(n25188), .ZN(n33807) );
  BUF_X4 U42590 ( .I(n51085), .Z(n56627) );
  XOR2_X1 U42593 ( .A1(n23592), .A2(n33861), .Z(n33893) );
  NAND3_X2 U42595 ( .A1(n55472), .A2(n2180), .A3(n61282), .ZN(n52389) );
  NAND2_X1 U42596 ( .A1(n32898), .A2(n34150), .ZN(n23599) );
  AOI22_X1 U42597 ( .A1(n43575), .A2(n41138), .B1(n41139), .B2(n43583), .ZN(
        n23602) );
  XOR2_X1 U42599 ( .A1(Key[139]), .A2(Ciphertext[186]), .Z(n24350) );
  NOR2_X1 U42600 ( .A1(n56134), .A2(n56162), .ZN(n56135) );
  AOI22_X1 U42602 ( .A1(n53470), .A2(n53503), .B1(n53468), .B2(n53469), .ZN(
        n53475) );
  XOR2_X1 U42603 ( .A1(n63548), .A2(n38941), .Z(n38779) );
  NOR2_X2 U42604 ( .A1(n63038), .A2(n9388), .ZN(n56638) );
  XOR2_X1 U42605 ( .A1(n29868), .A2(n29765), .Z(n23613) );
  NOR2_X2 U42611 ( .A1(n55442), .A2(n55440), .ZN(n55322) );
  AOI21_X1 U42614 ( .A1(n48192), .A2(n20788), .B(n48191), .ZN(n48198) );
  AOI21_X1 U42616 ( .A1(n28956), .A2(n28955), .B(n28954), .ZN(n24755) );
  XOR2_X1 U42617 ( .A1(n46656), .A2(n58807), .Z(n46658) );
  XOR2_X1 U42618 ( .A1(n23627), .A2(n61092), .Z(n50978) );
  XOR2_X1 U42619 ( .A1(n51360), .A2(n59555), .Z(n23628) );
  XOR2_X1 U42620 ( .A1(n23629), .A2(n33254), .Z(n33255) );
  XOR2_X1 U42621 ( .A1(n33253), .A2(n33252), .Z(n23629) );
  INV_X2 U42622 ( .I(n23630), .ZN(n26391) );
  XOR2_X1 U42625 ( .A1(n23633), .A2(n55792), .Z(Plaintext[129]) );
  NOR4_X2 U42626 ( .A1(n36790), .A2(n36803), .A3(n60925), .A4(n36796), .ZN(
        n36805) );
  XOR2_X1 U42629 ( .A1(n23638), .A2(n23929), .Z(Plaintext[28]) );
  BUF_X2 U42630 ( .I(n52207), .Z(n23642) );
  XOR2_X1 U42631 ( .A1(n50186), .A2(n50660), .Z(n50187) );
  NOR2_X1 U42633 ( .A1(n61261), .A2(n14111), .ZN(n23644) );
  NAND2_X2 U42634 ( .A1(n61741), .A2(n49529), .ZN(n49528) );
  NOR4_X2 U42635 ( .A1(n27542), .A2(n27541), .A3(n27540), .A4(n27539), .ZN(
        n27553) );
  NOR2_X1 U42637 ( .A1(n36743), .A2(n36748), .ZN(n23647) );
  NOR2_X2 U42638 ( .A1(n21018), .A2(n15754), .ZN(n35966) );
  INV_X2 U42639 ( .I(n57414), .ZN(n54982) );
  XOR2_X1 U42640 ( .A1(n45030), .A2(n46702), .Z(n23652) );
  NOR2_X1 U42643 ( .A1(n53972), .A2(n53980), .ZN(n53975) );
  BUF_X4 U42644 ( .I(n32610), .Z(n36483) );
  INV_X2 U42645 ( .I(n53621), .ZN(n53018) );
  NAND2_X2 U42646 ( .A1(n50462), .A2(n53861), .ZN(n53621) );
  INV_X2 U42647 ( .I(n26373), .ZN(n27397) );
  INV_X1 U42649 ( .I(n55117), .ZN(n25683) );
  BUF_X4 U42651 ( .I(n36732), .Z(n40994) );
  AOI21_X1 U42652 ( .A1(n28543), .A2(n27249), .B(n27248), .ZN(n26006) );
  XOR2_X1 U42655 ( .A1(n39769), .A2(n53958), .Z(n23680) );
  NAND2_X2 U42657 ( .A1(n1647), .A2(n16493), .ZN(n47500) );
  BUF_X2 U42665 ( .I(n43281), .Z(n23700) );
  XOR2_X1 U42666 ( .A1(n49294), .A2(n49295), .Z(n49321) );
  XOR2_X1 U42667 ( .A1(n25244), .A2(n19864), .Z(n25243) );
  BUF_X2 U42669 ( .I(n30535), .Z(n23706) );
  XOR2_X1 U42672 ( .A1(n23712), .A2(n23851), .Z(Plaintext[126]) );
  AND3_X1 U42673 ( .A1(n55754), .A2(n55758), .A3(n55753), .Z(n23713) );
  NAND2_X2 U42674 ( .A1(n55829), .A2(n22933), .ZN(n55800) );
  BUF_X2 U42675 ( .I(n34331), .Z(n23717) );
  XOR2_X1 U42679 ( .A1(Ciphertext[123]), .A2(Key[178]), .Z(n24139) );
  OR2_X1 U42687 ( .A1(n37218), .A2(n59617), .Z(n37220) );
  XOR2_X1 U42689 ( .A1(n26920), .A2(n23727), .Z(n32314) );
  XOR2_X1 U42690 ( .A1(n23719), .A2(n32312), .Z(n23727) );
  NAND2_X1 U42694 ( .A1(n39931), .A2(n41852), .ZN(n24610) );
  INV_X2 U42695 ( .I(n54662), .ZN(n54741) );
  XOR2_X1 U42696 ( .A1(n24932), .A2(n23733), .Z(n24931) );
  XOR2_X1 U42697 ( .A1(n39660), .A2(n16039), .Z(n23733) );
  NAND4_X2 U42698 ( .A1(n37912), .A2(n37911), .A3(n37910), .A4(n37909), .ZN(
        n37913) );
  INV_X4 U42699 ( .I(n24229), .ZN(n54196) );
  NAND2_X2 U42703 ( .A1(n18859), .A2(n25299), .ZN(n54170) );
  XOR2_X1 U42705 ( .A1(n23740), .A2(n44903), .Z(n23965) );
  OR3_X1 U42706 ( .A1(n49694), .A2(n48882), .A3(n22646), .Z(n45164) );
  XOR2_X1 U42709 ( .A1(n30400), .A2(n32121), .Z(n31872) );
  OR2_X1 U42710 ( .A1(n32150), .A2(n23749), .Z(n23748) );
  INV_X1 U42713 ( .I(n33131), .ZN(n24322) );
  INV_X2 U42714 ( .I(n49012), .ZN(n49006) );
  AOI21_X1 U42715 ( .A1(n55713), .A2(n61368), .B(n51902), .ZN(n51898) );
  BUF_X2 U42719 ( .I(n45726), .Z(n23759) );
  BUF_X2 U42720 ( .I(n51956), .Z(n23762) );
  XOR2_X1 U42723 ( .A1(Ciphertext[54]), .A2(Key[175]), .Z(n25300) );
  NAND2_X2 U42724 ( .A1(n28260), .A2(n28259), .ZN(n27936) );
  BUF_X2 U42725 ( .I(n31345), .Z(n23768) );
  NOR2_X2 U42726 ( .A1(n37051), .A2(n37050), .ZN(n36606) );
  XOR2_X1 U42728 ( .A1(n45393), .A2(n45392), .Z(n23783) );
  AND3_X1 U42731 ( .A1(n33324), .A2(n22428), .A3(n35611), .Z(n26224) );
  NAND2_X2 U42732 ( .A1(n29312), .A2(n26923), .ZN(n28855) );
  OAI22_X1 U42733 ( .A1(n29165), .A2(n23769), .B1(n29164), .B2(n29163), .ZN(
        n23798) );
  XOR2_X1 U42735 ( .A1(n7410), .A2(n25697), .Z(n23804) );
  XOR2_X1 U42736 ( .A1(n23808), .A2(n53499), .Z(Plaintext[27]) );
  NOR2_X1 U42737 ( .A1(n41654), .A2(n24360), .ZN(n23809) );
  NOR2_X1 U42738 ( .A1(n41653), .A2(n23811), .ZN(n23810) );
  NAND2_X1 U42739 ( .A1(n23817), .A2(n19290), .ZN(n25016) );
  OAI22_X1 U42740 ( .A1(n29625), .A2(n29624), .B1(n29622), .B2(n23578), .ZN(
        n23817) );
  NAND2_X2 U42741 ( .A1(n37949), .A2(n37948), .ZN(n39208) );
  INV_X4 U42742 ( .I(n25093), .ZN(n31074) );
  NAND2_X2 U42743 ( .A1(n27483), .A2(n27485), .ZN(n27537) );
  NOR2_X1 U42745 ( .A1(n24328), .A2(n30635), .ZN(n24327) );
  XOR2_X1 U42748 ( .A1(n38901), .A2(n38902), .Z(n23827) );
  NAND2_X2 U42749 ( .A1(n27691), .A2(n28470), .ZN(n28620) );
  NOR2_X2 U42750 ( .A1(n29372), .A2(n28811), .ZN(n23829) );
  NAND2_X1 U42753 ( .A1(n56923), .A2(n56921), .ZN(n23831) );
  BUF_X2 U42756 ( .I(n22861), .Z(n23835) );
  NAND2_X1 U42758 ( .A1(n26593), .A2(n26054), .ZN(n26053) );
  NAND2_X2 U42759 ( .A1(n26640), .A2(n23328), .ZN(n28300) );
  NAND2_X1 U42760 ( .A1(n40346), .A2(n15762), .ZN(n40347) );
  INV_X2 U42764 ( .I(n55656), .ZN(n55931) );
  OAI22_X1 U42768 ( .A1(n42406), .A2(n59394), .B1(n42405), .B2(n4723), .ZN(
        n42408) );
  NAND3_X1 U42769 ( .A1(n19982), .A2(n41934), .A3(n41933), .ZN(n41935) );
  NOR2_X2 U42771 ( .A1(n40229), .A2(n40295), .ZN(n40306) );
  INV_X2 U42773 ( .I(n27159), .ZN(n27611) );
  XOR2_X1 U42774 ( .A1(n52175), .A2(n23861), .Z(n49337) );
  XOR2_X1 U42775 ( .A1(n49321), .A2(n51991), .Z(n23861) );
  XOR2_X1 U42776 ( .A1(n6384), .A2(n51358), .Z(n49295) );
  XOR2_X1 U42777 ( .A1(n19627), .A2(n23714), .Z(n31317) );
  NOR3_X2 U42778 ( .A1(n29735), .A2(n24651), .A3(n29734), .ZN(n32383) );
  NAND2_X2 U42779 ( .A1(n54667), .A2(n54666), .ZN(n54662) );
  INV_X1 U42780 ( .I(n45747), .ZN(n46989) );
  AOI21_X1 U42782 ( .A1(n44770), .A2(n63311), .B(n23866), .ZN(n23865) );
  NOR2_X1 U42783 ( .A1(n1082), .A2(n44770), .ZN(n23866) );
  NAND2_X2 U42784 ( .A1(n28259), .A2(n23769), .ZN(n29168) );
  NAND2_X2 U42786 ( .A1(n53324), .A2(n53368), .ZN(n23871) );
  INV_X2 U42790 ( .I(n29383), .ZN(n29668) );
  INV_X2 U42792 ( .I(n27336), .ZN(n29671) );
  OR2_X1 U42793 ( .A1(n26897), .A2(n26896), .Z(n23888) );
  INV_X2 U42798 ( .I(n32529), .ZN(n32807) );
  XOR2_X1 U42800 ( .A1(n44731), .A2(n46573), .Z(n23902) );
  NAND2_X1 U42801 ( .A1(n49755), .A2(n49756), .ZN(n49758) );
  NAND2_X2 U42802 ( .A1(n29671), .A2(n29661), .ZN(n28200) );
  NAND3_X1 U42806 ( .A1(n45684), .A2(n45682), .A3(n45683), .ZN(n45685) );
  NAND2_X2 U42809 ( .A1(n49063), .A2(n20461), .ZN(n48292) );
  INV_X2 U42810 ( .I(n27185), .ZN(n26654) );
  XOR2_X1 U42813 ( .A1(n32417), .A2(n32413), .Z(n23915) );
  OR2_X1 U42814 ( .A1(n27660), .A2(n27668), .Z(n23916) );
  AND3_X1 U42819 ( .A1(n54448), .A2(n54654), .A3(n54688), .Z(n23924) );
  XOR2_X1 U42820 ( .A1(n37874), .A2(n37676), .Z(n25249) );
  XOR2_X1 U42822 ( .A1(n32470), .A2(n7264), .Z(n31866) );
  NOR2_X1 U42823 ( .A1(n28799), .A2(n23930), .ZN(n28807) );
  NAND2_X2 U42824 ( .A1(n21364), .A2(n23897), .ZN(n54321) );
  INV_X4 U42826 ( .I(n26226), .ZN(n48514) );
  INV_X4 U42830 ( .I(n52977), .ZN(n53916) );
  INV_X2 U42831 ( .I(n28537), .ZN(n27876) );
  XOR2_X1 U42833 ( .A1(n39583), .A2(n39582), .Z(n39675) );
  OAI21_X1 U42840 ( .A1(n53237), .A2(n53236), .B(n53235), .ZN(n25903) );
  NOR2_X2 U42843 ( .A1(n25115), .A2(n25116), .ZN(n53741) );
  OR2_X2 U42844 ( .A1(n53036), .A2(n54017), .Z(n24586) );
  OR2_X1 U42845 ( .A1(n27550), .A2(n27487), .Z(n23964) );
  XOR2_X1 U42846 ( .A1(n23965), .A2(n44904), .Z(n25472) );
  NOR2_X1 U42849 ( .A1(n35827), .A2(n25389), .ZN(n34715) );
  NOR2_X1 U42854 ( .A1(n36125), .A2(n22295), .ZN(n23975) );
  INV_X2 U42855 ( .I(n23979), .ZN(n26641) );
  NOR2_X2 U42859 ( .A1(n23549), .A2(n23578), .ZN(n29626) );
  XOR2_X1 U42860 ( .A1(n31386), .A2(n30853), .Z(n23985) );
  BUF_X2 U42863 ( .I(n46521), .Z(n23987) );
  NOR3_X2 U42864 ( .A1(n56600), .A2(n24647), .A3(n13920), .ZN(n56986) );
  INV_X2 U42866 ( .I(n29167), .ZN(n28260) );
  NAND2_X1 U42868 ( .A1(n23996), .A2(n23994), .ZN(n23993) );
  NOR2_X1 U42869 ( .A1(n47415), .A2(n263), .ZN(n23995) );
  XOR2_X1 U42871 ( .A1(n39205), .A2(n39204), .Z(n23998) );
  XOR2_X1 U42873 ( .A1(n24004), .A2(n54407), .Z(Plaintext[70]) );
  INV_X4 U42878 ( .I(n34355), .ZN(n34247) );
  BUF_X2 U42879 ( .I(Key[152]), .Z(n24011) );
  XOR2_X1 U42881 ( .A1(n42955), .A2(n42954), .Z(n24020) );
  AOI22_X1 U42883 ( .A1(n24022), .A2(n44068), .B1(n45519), .B2(n45749), .ZN(
        n44069) );
  NAND2_X2 U42884 ( .A1(n35031), .A2(n13982), .ZN(n34502) );
  NOR2_X2 U42885 ( .A1(n23982), .A2(n55494), .ZN(n55497) );
  NAND2_X2 U42887 ( .A1(n33557), .A2(n33558), .ZN(n36195) );
  AND2_X1 U42889 ( .A1(n1715), .A2(n43357), .Z(n40367) );
  BUF_X2 U42890 ( .I(n52013), .Z(n24025) );
  NAND3_X1 U42891 ( .A1(n24027), .A2(n42072), .A3(n13750), .ZN(n40095) );
  INV_X4 U42892 ( .I(n40416), .ZN(n41470) );
  NOR2_X2 U42897 ( .A1(n53420), .A2(n53860), .ZN(n53022) );
  XOR2_X1 U42901 ( .A1(n44257), .A2(n43963), .Z(n24034) );
  NAND2_X2 U42904 ( .A1(n61805), .A2(n48302), .ZN(n49068) );
  AND3_X1 U42905 ( .A1(n54750), .A2(n23448), .A3(n24038), .Z(n54753) );
  XOR2_X1 U42907 ( .A1(n36638), .A2(n38192), .Z(n38637) );
  BUF_X2 U42908 ( .I(n29619), .Z(n24052) );
  NAND2_X2 U42909 ( .A1(n34613), .A2(n23410), .ZN(n33984) );
  OR2_X1 U42912 ( .A1(n49854), .A2(n49856), .Z(n26108) );
  NAND2_X2 U42913 ( .A1(n41119), .A2(n62107), .ZN(n39829) );
  XOR2_X1 U42914 ( .A1(n33256), .A2(n16287), .Z(n33263) );
  NAND4_X2 U42915 ( .A1(n31547), .A2(n16108), .A3(n31546), .A4(n31545), .ZN(
        n31548) );
  INV_X4 U42917 ( .I(n35805), .ZN(n35799) );
  XOR2_X1 U42918 ( .A1(n32392), .A2(n31880), .Z(n31832) );
  XOR2_X1 U42919 ( .A1(n22187), .A2(n31831), .Z(n32392) );
  BUF_X4 U42922 ( .I(n32739), .Z(n35691) );
  NAND2_X2 U42924 ( .A1(n25128), .A2(n24394), .ZN(n24393) );
  INV_X4 U42929 ( .I(n25669), .ZN(n29586) );
  XOR2_X1 U42935 ( .A1(n56142), .A2(n56143), .Z(Plaintext[144]) );
  NAND2_X1 U42936 ( .A1(n29249), .A2(n29248), .ZN(n25881) );
  AND2_X1 U42937 ( .A1(n47864), .A2(n47863), .Z(n24096) );
  AND2_X1 U42938 ( .A1(n41780), .A2(n41781), .Z(n24101) );
  AND2_X1 U42948 ( .A1(n40325), .A2(n40327), .Z(n24387) );
  INV_X4 U42950 ( .I(n57017), .ZN(n53212) );
  BUF_X4 U42951 ( .I(n25347), .Z(n56867) );
  NAND3_X1 U42954 ( .A1(n56286), .A2(n56291), .A3(n24032), .ZN(n24120) );
  OAI21_X1 U42955 ( .A1(n32771), .A2(n32772), .B(n1782), .ZN(n24121) );
  INV_X4 U42956 ( .I(n11883), .ZN(n42666) );
  INV_X2 U42957 ( .I(n27594), .ZN(n27174) );
  NAND2_X2 U42959 ( .A1(n59180), .A2(n11841), .ZN(n56351) );
  NOR2_X2 U42960 ( .A1(n39095), .A2(n25570), .ZN(n39099) );
  XOR2_X1 U42961 ( .A1(n46598), .A2(n24126), .Z(n46418) );
  XOR2_X1 U42962 ( .A1(n44092), .A2(n16320), .Z(n24126) );
  NOR2_X2 U42963 ( .A1(n42155), .A2(n22898), .ZN(n42587) );
  XOR2_X1 U42965 ( .A1(n50187), .A2(n51619), .Z(n52743) );
  AOI21_X2 U42968 ( .A1(n32788), .A2(n32787), .B(n32786), .ZN(n36030) );
  NOR2_X1 U42969 ( .A1(n13412), .A2(n24251), .ZN(n30863) );
  INV_X2 U42971 ( .I(n24139), .ZN(n27823) );
  INV_X2 U42976 ( .I(n823), .ZN(n33243) );
  INV_X1 U42977 ( .I(n29567), .ZN(n24159) );
  XOR2_X1 U42979 ( .A1(n45386), .A2(n43260), .Z(n43664) );
  INV_X2 U42980 ( .I(n24166), .ZN(n55444) );
  NOR2_X2 U42981 ( .A1(n50123), .A2(n18608), .ZN(n50291) );
  NOR2_X1 U42982 ( .A1(n50284), .A2(n48716), .ZN(n24167) );
  XOR2_X1 U42983 ( .A1(n37646), .A2(n24169), .Z(n37842) );
  XOR2_X1 U42985 ( .A1(n37261), .A2(n24169), .Z(n37263) );
  XOR2_X1 U42987 ( .A1(n25316), .A2(n51477), .Z(n24183) );
  NOR2_X2 U42989 ( .A1(n47604), .A2(n3510), .ZN(n47610) );
  INV_X2 U42991 ( .I(n24192), .ZN(n54973) );
  OAI21_X1 U42992 ( .A1(n30384), .A2(n29488), .B(n24199), .ZN(n29489) );
  NAND3_X1 U42993 ( .A1(n29491), .A2(n29494), .A3(n24199), .ZN(n29497) );
  XOR2_X1 U42996 ( .A1(n38913), .A2(n38068), .Z(n24211) );
  XOR2_X1 U42997 ( .A1(n10531), .A2(n16305), .Z(n24212) );
  NOR2_X2 U43000 ( .A1(n25302), .A2(n25301), .ZN(n27988) );
  NAND2_X1 U43001 ( .A1(n41951), .A2(n61435), .ZN(n24217) );
  XOR2_X1 U43003 ( .A1(n16691), .A2(n24227), .Z(n50876) );
  XOR2_X1 U43004 ( .A1(n24758), .A2(n50875), .Z(n24227) );
  XOR2_X1 U43005 ( .A1(n52030), .A2(n51342), .Z(n51343) );
  XOR2_X1 U43006 ( .A1(n51931), .A2(n64825), .Z(n50148) );
  OAI21_X1 U43007 ( .A1(n57678), .A2(n29304), .B(n24233), .ZN(n24232) );
  XOR2_X1 U43008 ( .A1(n38792), .A2(n39233), .Z(n24234) );
  NAND2_X2 U43010 ( .A1(n21364), .A2(n54088), .ZN(n54087) );
  OAI21_X1 U43012 ( .A1(n24556), .A2(n31187), .B(n63394), .ZN(n28969) );
  XOR2_X1 U43014 ( .A1(n32592), .A2(n15733), .Z(n31763) );
  XOR2_X1 U43016 ( .A1(n39345), .A2(n22916), .Z(n38373) );
  INV_X2 U43018 ( .I(n55248), .ZN(n55397) );
  XOR2_X1 U43019 ( .A1(n25088), .A2(n25087), .Z(n52532) );
  INV_X1 U43020 ( .I(n8449), .ZN(n38180) );
  NAND2_X1 U43024 ( .A1(n39804), .A2(n39981), .ZN(n24271) );
  NAND2_X1 U43025 ( .A1(n24273), .A2(n33420), .ZN(n33418) );
  XOR2_X1 U43026 ( .A1(n39226), .A2(n38739), .Z(n38740) );
  XOR2_X1 U43027 ( .A1(n39585), .A2(n1520), .Z(n39226) );
  NOR2_X2 U43028 ( .A1(n26186), .A2(n41359), .ZN(n46433) );
  INV_X2 U43035 ( .I(n46165), .ZN(n46438) );
  NOR2_X1 U43036 ( .A1(n16694), .A2(n23478), .ZN(n30548) );
  INV_X4 U43042 ( .I(n39241), .ZN(n42477) );
  XOR2_X1 U43043 ( .A1(n14249), .A2(n33231), .Z(n24315) );
  NAND3_X1 U43044 ( .A1(n57559), .A2(n24316), .A3(n15689), .ZN(n28427) );
  AOI21_X1 U43045 ( .A1(n29580), .A2(n29575), .B(n24316), .ZN(n28923) );
  NAND2_X1 U43046 ( .A1(n61964), .A2(n56510), .ZN(n56511) );
  XOR2_X1 U43047 ( .A1(n31582), .A2(n31583), .Z(n31684) );
  NAND3_X1 U43048 ( .A1(n27776), .A2(n29863), .A3(n64940), .ZN(n27777) );
  INV_X1 U43050 ( .I(n39314), .ZN(n38101) );
  INV_X1 U43051 ( .I(n22781), .ZN(n32628) );
  XOR2_X1 U43052 ( .A1(n22781), .A2(n10378), .Z(n24349) );
  NAND2_X1 U43053 ( .A1(n24351), .A2(n61579), .ZN(n36300) );
  NAND2_X1 U43056 ( .A1(n15550), .A2(n20138), .ZN(n48316) );
  CLKBUF_X4 U43057 ( .I(Key[39]), .Z(n24355) );
  XOR2_X1 U43058 ( .A1(Ciphertext[62]), .A2(Key[39]), .Z(n28224) );
  XOR2_X1 U43059 ( .A1(n55624), .A2(n24355), .Z(n45816) );
  XOR2_X1 U43060 ( .A1(n53272), .A2(n24355), .Z(n44759) );
  XOR2_X1 U43061 ( .A1(n57131), .A2(n24355), .Z(n39611) );
  XOR2_X1 U43062 ( .A1(n49426), .A2(n24355), .Z(n37749) );
  XOR2_X1 U43063 ( .A1(n39361), .A2(n24355), .Z(n32078) );
  XOR2_X1 U43064 ( .A1(n27640), .A2(n24355), .Z(n37674) );
  XOR2_X1 U43065 ( .A1(n39183), .A2(n24355), .Z(n31381) );
  XOR2_X1 U43066 ( .A1(n50621), .A2(n24355), .Z(n50622) );
  NAND2_X1 U43068 ( .A1(n34927), .A2(n4151), .ZN(n24356) );
  NOR2_X2 U43070 ( .A1(n24990), .A2(n24991), .ZN(n41914) );
  XOR2_X1 U43071 ( .A1(n46161), .A2(n1268), .Z(n46610) );
  AOI21_X1 U43072 ( .A1(n24367), .A2(n45801), .B(n23099), .ZN(n45802) );
  XOR2_X1 U43078 ( .A1(n39579), .A2(n30908), .Z(n24383) );
  INV_X2 U43079 ( .I(n24391), .ZN(n25785) );
  XOR2_X1 U43082 ( .A1(n49125), .A2(n24397), .Z(n49127) );
  XOR2_X1 U43083 ( .A1(n51537), .A2(n24397), .Z(n51538) );
  INV_X2 U43085 ( .I(n24406), .ZN(n28349) );
  XOR2_X1 U43086 ( .A1(n38803), .A2(n38670), .Z(n24408) );
  NOR2_X2 U43087 ( .A1(n11207), .A2(n51860), .ZN(n54346) );
  XOR2_X1 U43088 ( .A1(n24412), .A2(n32388), .Z(n24414) );
  XOR2_X1 U43089 ( .A1(n31590), .A2(n24413), .Z(n32388) );
  XOR2_X1 U43090 ( .A1(n31765), .A2(n18296), .Z(n24412) );
  INV_X2 U43091 ( .I(n24415), .ZN(n54017) );
  XOR2_X1 U43092 ( .A1(n63005), .A2(n44548), .Z(n24416) );
  XOR2_X1 U43095 ( .A1(n24432), .A2(n31832), .Z(n31833) );
  XOR2_X1 U43098 ( .A1(n23898), .A2(n24435), .Z(n37970) );
  XOR2_X1 U43099 ( .A1(n24435), .A2(n26063), .Z(n37747) );
  NAND2_X2 U43100 ( .A1(n24442), .A2(n24438), .ZN(n26740) );
  XOR2_X1 U43103 ( .A1(Ciphertext[104]), .A2(Key[141]), .Z(n27709) );
  INV_X2 U43105 ( .I(n24447), .ZN(n38758) );
  XOR2_X1 U43106 ( .A1(n24449), .A2(n23440), .Z(n45085) );
  XOR2_X1 U43107 ( .A1(n46280), .A2(n24449), .Z(n46281) );
  NOR2_X2 U43108 ( .A1(n24452), .A2(n45084), .ZN(n49701) );
  OR2_X1 U43109 ( .A1(n40140), .A2(n40139), .Z(n24453) );
  OR2_X1 U43111 ( .A1(n55293), .A2(n55677), .Z(n24465) );
  INV_X2 U43118 ( .I(n24481), .ZN(n29370) );
  NAND2_X1 U43119 ( .A1(n53032), .A2(n54341), .ZN(n24483) );
  XOR2_X1 U43120 ( .A1(Key[190]), .A2(Ciphertext[15]), .Z(n28303) );
  NOR2_X2 U43121 ( .A1(n57462), .A2(n40626), .ZN(n41198) );
  NAND2_X1 U43122 ( .A1(n35822), .A2(n24488), .ZN(n35823) );
  OR2_X1 U43123 ( .A1(n49090), .A2(n24490), .Z(n49679) );
  NAND2_X1 U43124 ( .A1(n49676), .A2(n49677), .ZN(n24490) );
  NAND4_X2 U43126 ( .A1(n33819), .A2(n33818), .A3(n24497), .A4(n24496), .ZN(
        n33930) );
  NOR2_X2 U43130 ( .A1(n5267), .A2(n59129), .ZN(n30552) );
  NOR2_X1 U43131 ( .A1(n10554), .A2(n42441), .ZN(n24505) );
  NAND2_X1 U43134 ( .A1(n54259), .A2(n1280), .ZN(n54282) );
  XOR2_X1 U43135 ( .A1(n38729), .A2(n38530), .Z(n38310) );
  XOR2_X1 U43136 ( .A1(n61662), .A2(n46356), .Z(n24516) );
  XOR2_X1 U43137 ( .A1(n24521), .A2(n46650), .Z(n44161) );
  NOR2_X2 U43140 ( .A1(n56547), .A2(n52706), .ZN(n57012) );
  XOR2_X1 U43141 ( .A1(n24535), .A2(n24098), .Z(n33063) );
  XOR2_X1 U43142 ( .A1(n54587), .A2(n24535), .Z(n43768) );
  XOR2_X1 U43143 ( .A1(n55833), .A2(n24535), .Z(n50697) );
  XOR2_X1 U43144 ( .A1(n53375), .A2(n24535), .Z(n29892) );
  XOR2_X1 U43145 ( .A1(n56901), .A2(n24535), .Z(n38236) );
  XOR2_X1 U43146 ( .A1(n51193), .A2(n24535), .Z(n38165) );
  XOR2_X1 U43147 ( .A1(n38009), .A2(n24535), .Z(n38010) );
  XOR2_X1 U43148 ( .A1(n38994), .A2(n9956), .Z(n38890) );
  XOR2_X1 U43149 ( .A1(n22922), .A2(n47939), .Z(n47940) );
  XOR2_X1 U43152 ( .A1(n23714), .A2(n23791), .Z(n32331) );
  NAND2_X2 U43153 ( .A1(n62995), .A2(n33797), .ZN(n33801) );
  NAND2_X1 U43156 ( .A1(n35653), .A2(n62995), .ZN(n24574) );
  NAND2_X2 U43157 ( .A1(n1780), .A2(n37096), .ZN(n37322) );
  AOI21_X1 U43158 ( .A1(n56294), .A2(n56293), .B(n24584), .ZN(n56308) );
  INV_X2 U43161 ( .I(n24922), .ZN(n53036) );
  OR2_X1 U43162 ( .A1(n43323), .A2(n43324), .Z(n24591) );
  XOR2_X1 U43166 ( .A1(n52559), .A2(n50501), .Z(n52105) );
  XOR2_X1 U43167 ( .A1(n33160), .A2(n24600), .Z(n24599) );
  XOR2_X1 U43169 ( .A1(n39728), .A2(n57131), .Z(n38298) );
  INV_X2 U43171 ( .I(n24617), .ZN(n40962) );
  XOR2_X1 U43172 ( .A1(n32237), .A2(n24632), .Z(n32241) );
  XOR2_X1 U43173 ( .A1(n32236), .A2(n32235), .Z(n24632) );
  NAND2_X2 U43174 ( .A1(n26846), .A2(n26845), .ZN(n32089) );
  INV_X1 U43175 ( .I(n24633), .ZN(n40354) );
  XOR2_X1 U43177 ( .A1(n24639), .A2(n24638), .Z(n46412) );
  XOR2_X1 U43178 ( .A1(n61662), .A2(n46406), .Z(n24638) );
  AOI21_X1 U43181 ( .A1(n36748), .A2(n12863), .B(n36740), .ZN(n35857) );
  XOR2_X1 U43182 ( .A1(n1268), .A2(n44313), .Z(n44314) );
  XOR2_X1 U43183 ( .A1(n1268), .A2(n46505), .Z(n46506) );
  INV_X2 U43185 ( .I(n25580), .ZN(n47623) );
  OR2_X1 U43186 ( .A1(n37190), .A2(n37327), .Z(n24658) );
  XOR2_X1 U43188 ( .A1(n24672), .A2(n31732), .Z(n25245) );
  NAND2_X1 U43189 ( .A1(n55416), .A2(n55250), .ZN(n24676) );
  NAND2_X2 U43190 ( .A1(n43050), .A2(n43051), .ZN(n46702) );
  AND2_X1 U43191 ( .A1(n47447), .A2(n47446), .Z(n24683) );
  INV_X1 U43193 ( .I(n24684), .ZN(n40893) );
  XOR2_X1 U43197 ( .A1(n44856), .A2(n44857), .Z(n46511) );
  INV_X2 U43199 ( .I(n24697), .ZN(n45992) );
  XOR2_X1 U43201 ( .A1(n24698), .A2(n24704), .Z(n32508) );
  XOR2_X1 U43202 ( .A1(n11310), .A2(n37747), .Z(n24699) );
  XOR2_X1 U43203 ( .A1(n23429), .A2(n37754), .Z(n24700) );
  NAND2_X1 U43204 ( .A1(n24836), .A2(n24703), .ZN(n24835) );
  OAI22_X1 U43205 ( .A1(n28045), .A2(n21065), .B1(n24703), .B2(n27125), .ZN(
        n27127) );
  NAND2_X1 U43206 ( .A1(n47426), .A2(n47425), .ZN(n24706) );
  XOR2_X1 U43208 ( .A1(n51148), .A2(n51227), .Z(n51539) );
  NAND2_X1 U43210 ( .A1(n12863), .A2(n65234), .ZN(n24721) );
  NAND2_X1 U43211 ( .A1(n17720), .A2(n36742), .ZN(n24724) );
  AOI22_X1 U43216 ( .A1(n56986), .A2(n56993), .B1(n52890), .B2(n52889), .ZN(
        n52894) );
  NAND2_X2 U43217 ( .A1(n25329), .A2(n30967), .ZN(n35994) );
  NAND2_X1 U43219 ( .A1(n10452), .A2(n23634), .ZN(n24781) );
  XOR2_X1 U43222 ( .A1(n51823), .A2(n49190), .Z(n26107) );
  NAND2_X2 U43224 ( .A1(n36742), .A2(n36740), .ZN(n35423) );
  INV_X2 U43227 ( .I(n28806), .ZN(n28811) );
  INV_X2 U43229 ( .I(n16194), .ZN(n24801) );
  INV_X1 U43231 ( .I(n24806), .ZN(n24808) );
  INV_X2 U43233 ( .I(n24811), .ZN(n29727) );
  NOR3_X2 U43235 ( .A1(n27026), .A2(n25390), .A3(n16172), .ZN(n24811) );
  XNOR2_X1 U43236 ( .A1(n25888), .A2(n52192), .ZN(n50979) );
  NAND3_X1 U43238 ( .A1(n48600), .A2(n47530), .A3(n24820), .ZN(n47019) );
  NOR4_X2 U43239 ( .A1(n28164), .A2(n27452), .A3(n27453), .A4(n29307), .ZN(
        n24823) );
  INV_X4 U43240 ( .I(n61935), .ZN(n37224) );
  XOR2_X1 U43241 ( .A1(n33232), .A2(n33240), .Z(n24828) );
  INV_X2 U43242 ( .I(n24834), .ZN(n41105) );
  NAND2_X1 U43244 ( .A1(n30726), .A2(n30727), .ZN(n24842) );
  XOR2_X1 U43247 ( .A1(n24849), .A2(n18891), .Z(n52028) );
  NAND2_X1 U43248 ( .A1(n29511), .A2(n24852), .ZN(n29004) );
  INV_X1 U43249 ( .I(Ciphertext[51]), .ZN(n24854) );
  XOR2_X1 U43250 ( .A1(n24859), .A2(n39767), .Z(n24860) );
  NOR2_X1 U43251 ( .A1(n40854), .A2(n64475), .ZN(n24861) );
  AOI21_X2 U43253 ( .A1(n24867), .A2(n59192), .B(n24865), .ZN(n55768) );
  NOR2_X1 U43254 ( .A1(n26336), .A2(n28300), .ZN(n27080) );
  NAND2_X1 U43255 ( .A1(n43381), .A2(n24884), .ZN(n41698) );
  INV_X2 U43256 ( .I(n24885), .ZN(n28312) );
  XOR2_X1 U43258 ( .A1(n24888), .A2(Key[68]), .Z(n24889) );
  XOR2_X1 U43259 ( .A1(n31411), .A2(n5436), .Z(n31413) );
  XOR2_X1 U43260 ( .A1(n5436), .A2(n44164), .Z(n33868) );
  XOR2_X1 U43261 ( .A1(n32326), .A2(n5436), .Z(n31835) );
  NOR2_X1 U43262 ( .A1(n28083), .A2(n24896), .ZN(n28084) );
  AOI22_X1 U43263 ( .A1(n28307), .A2(n28310), .B1(n28306), .B2(n28312), .ZN(
        n24897) );
  NAND2_X1 U43264 ( .A1(n28314), .A2(n23324), .ZN(n24900) );
  NAND2_X1 U43265 ( .A1(n24902), .A2(n28315), .ZN(n24901) );
  OAI21_X1 U43266 ( .A1(n28310), .A2(n28311), .B(n19156), .ZN(n24902) );
  NOR2_X1 U43267 ( .A1(n47073), .A2(n11458), .ZN(n24906) );
  OR2_X1 U43268 ( .A1(n11458), .A2(n47073), .Z(n48766) );
  NAND2_X1 U43269 ( .A1(n60974), .A2(n9777), .ZN(n55383) );
  NAND2_X1 U43270 ( .A1(n36695), .A2(n57210), .ZN(n36697) );
  XOR2_X1 U43271 ( .A1(n38711), .A2(n39190), .Z(n24912) );
  XOR2_X1 U43273 ( .A1(n44418), .A2(n44419), .Z(n24915) );
  INV_X2 U43274 ( .I(n29619), .ZN(n28675) );
  XOR2_X1 U43276 ( .A1(n37736), .A2(n50475), .Z(n44257) );
  XOR2_X1 U43277 ( .A1(n9884), .A2(n53124), .Z(n49289) );
  XOR2_X1 U43278 ( .A1(n9884), .A2(n56819), .Z(n31746) );
  XOR2_X1 U43279 ( .A1(n9884), .A2(n55655), .Z(n51815) );
  XOR2_X1 U43280 ( .A1(n9884), .A2(n54587), .Z(n39685) );
  XOR2_X1 U43281 ( .A1(n37713), .A2(n9884), .Z(n32740) );
  XOR2_X1 U43282 ( .A1(n31338), .A2(n9884), .Z(n31339) );
  XOR2_X1 U43283 ( .A1(n50328), .A2(n9884), .Z(n50329) );
  XOR2_X1 U43284 ( .A1(n55395), .A2(n55903), .Z(n24920) );
  OAI21_X1 U43285 ( .A1(n24921), .A2(n21956), .B(n24080), .ZN(n29122) );
  NAND2_X2 U43286 ( .A1(n29119), .A2(n28211), .ZN(n24921) );
  XNOR2_X1 U43289 ( .A1(n32052), .A2(n32051), .ZN(n24935) );
  INV_X1 U43290 ( .I(n24942), .ZN(n34237) );
  OR2_X1 U43291 ( .A1(n40643), .A2(n10587), .Z(n24950) );
  NOR2_X2 U43293 ( .A1(n25848), .A2(n6609), .ZN(n29533) );
  INV_X2 U43298 ( .I(n24977), .ZN(n41197) );
  XOR2_X1 U43299 ( .A1(n44973), .A2(n5118), .Z(n44418) );
  MUX2_X1 U43300 ( .I0(n33895), .I1(n33915), .S(n24983), .Z(n33916) );
  NOR2_X1 U43301 ( .A1(n19102), .A2(n60422), .ZN(n24984) );
  XOR2_X1 U43304 ( .A1(n34481), .A2(n2823), .Z(n34496) );
  XOR2_X1 U43305 ( .A1(n16337), .A2(n36944), .Z(n25010) );
  XOR2_X1 U43307 ( .A1(n45021), .A2(n44342), .Z(n25012) );
  OR2_X1 U43308 ( .A1(n29627), .A2(n60990), .Z(n25017) );
  XOR2_X1 U43313 ( .A1(n25388), .A2(n32038), .Z(n25025) );
  INV_X1 U43314 ( .I(n25026), .ZN(n43596) );
  NAND2_X1 U43317 ( .A1(n30627), .A2(n30628), .ZN(n25038) );
  XOR2_X1 U43318 ( .A1(n31674), .A2(n4901), .Z(n31677) );
  NAND2_X1 U43324 ( .A1(n30752), .A2(n30760), .ZN(n25053) );
  NAND2_X1 U43326 ( .A1(n18583), .A2(n3691), .ZN(n25056) );
  INV_X2 U43327 ( .I(n25059), .ZN(n40970) );
  XOR2_X1 U43328 ( .A1(n52030), .A2(n50626), .Z(n25060) );
  NAND3_X2 U43330 ( .A1(n47071), .A2(n47072), .A3(n26066), .ZN(n51601) );
  XOR2_X1 U43332 ( .A1(n25873), .A2(n16034), .Z(n53377) );
  NAND2_X1 U43333 ( .A1(n38027), .A2(n11126), .ZN(n25073) );
  XOR2_X1 U43334 ( .A1(n36528), .A2(n23277), .Z(n25075) );
  NOR2_X2 U43335 ( .A1(n53793), .A2(n53809), .ZN(n53828) );
  XOR2_X1 U43338 ( .A1(n51805), .A2(n50575), .Z(n25087) );
  XOR2_X1 U43339 ( .A1(n50574), .A2(n51129), .Z(n25088) );
  AOI22_X1 U43340 ( .A1(n1628), .A2(n48691), .B1(n64167), .B2(n25091), .ZN(
        n48693) );
  XOR2_X1 U43342 ( .A1(Ciphertext[181]), .A2(Key[8]), .Z(n25094) );
  NAND2_X1 U43343 ( .A1(n33600), .A2(n23812), .ZN(n32763) );
  INV_X2 U43345 ( .I(n25947), .ZN(n53376) );
  XOR2_X1 U43346 ( .A1(n52520), .A2(n51548), .Z(n52522) );
  OAI21_X1 U43347 ( .A1(n25101), .A2(n33337), .B(n35690), .ZN(n25100) );
  NAND2_X2 U43348 ( .A1(n48545), .A2(n48148), .ZN(n48553) );
  XOR2_X1 U43349 ( .A1(n62966), .A2(n37260), .Z(n37261) );
  XOR2_X1 U43350 ( .A1(n25111), .A2(n31639), .Z(n25653) );
  XOR2_X1 U43351 ( .A1(n23369), .A2(n23461), .Z(n32188) );
  XOR2_X1 U43352 ( .A1(n9108), .A2(n32290), .Z(n32291) );
  CLKBUF_X4 U43357 ( .I(n53727), .Z(n25116) );
  NAND3_X1 U43363 ( .A1(n40963), .A2(n25139), .A3(n38607), .ZN(n25138) );
  NAND2_X1 U43365 ( .A1(n60543), .A2(n20782), .ZN(n25159) );
  NAND2_X1 U43370 ( .A1(n25172), .A2(n18422), .ZN(n54513) );
  OAI22_X1 U43371 ( .A1(n54523), .A2(n25172), .B1(n18422), .B2(n54560), .ZN(
        n54512) );
  NAND2_X1 U43372 ( .A1(n54575), .A2(n25172), .ZN(n54532) );
  OAI21_X1 U43374 ( .A1(n55983), .A2(n25173), .B(n55982), .ZN(n55993) );
  XOR2_X1 U43375 ( .A1(n13639), .A2(n50884), .Z(n50896) );
  XOR2_X1 U43376 ( .A1(n22781), .A2(n25176), .Z(n33068) );
  XOR2_X1 U43377 ( .A1(n33141), .A2(n25176), .Z(n33142) );
  XOR2_X1 U43378 ( .A1(n39455), .A2(n25177), .Z(n38242) );
  XOR2_X1 U43379 ( .A1(n38807), .A2(n25177), .Z(n38808) );
  XOR2_X1 U43380 ( .A1(n25177), .A2(n39598), .Z(n38513) );
  NAND2_X1 U43382 ( .A1(n28934), .A2(n25186), .ZN(n25185) );
  AOI21_X1 U43383 ( .A1(n30231), .A2(n1863), .B(n19218), .ZN(n25186) );
  XOR2_X1 U43384 ( .A1(n33232), .A2(n33164), .Z(n25190) );
  XOR2_X1 U43385 ( .A1(n52619), .A2(n14870), .Z(n52620) );
  INV_X2 U43386 ( .I(n27828), .ZN(n26898) );
  NOR2_X2 U43387 ( .A1(n27665), .A2(n27841), .ZN(n27828) );
  INV_X2 U43390 ( .I(n25211), .ZN(n39692) );
  XOR2_X1 U43391 ( .A1(n20742), .A2(n9635), .Z(n50392) );
  XOR2_X1 U43392 ( .A1(n20742), .A2(n51424), .Z(n51426) );
  XOR2_X1 U43393 ( .A1(n6216), .A2(n51517), .Z(n51518) );
  NOR2_X1 U43394 ( .A1(n23298), .A2(n25229), .ZN(n40338) );
  INV_X2 U43398 ( .I(n27494), .ZN(n29297) );
  OAI21_X1 U43399 ( .A1(n25239), .A2(n22627), .B(n495), .ZN(n25238) );
  INV_X1 U43401 ( .I(n42488), .ZN(n39408) );
  INV_X1 U43402 ( .I(n35437), .ZN(n36362) );
  XOR2_X1 U43403 ( .A1(n21340), .A2(n52144), .Z(n25254) );
  INV_X2 U43406 ( .I(n28045), .ZN(n28053) );
  INV_X2 U43407 ( .I(n52383), .ZN(n54778) );
  NAND2_X2 U43408 ( .A1(n28314), .A2(n28311), .ZN(n27592) );
  NOR2_X2 U43409 ( .A1(n57192), .A2(n15713), .ZN(n53196) );
  INV_X4 U43412 ( .I(n31059), .ZN(n30174) );
  NOR2_X2 U43414 ( .A1(n18583), .A2(n37224), .ZN(n36269) );
  NOR2_X2 U43416 ( .A1(n28119), .A2(n28127), .ZN(n29621) );
  NOR2_X2 U43418 ( .A1(n23056), .A2(n12908), .ZN(n31035) );
  INV_X1 U43420 ( .I(n30959), .ZN(n25338) );
  NAND2_X1 U43421 ( .A1(n45941), .A2(n25557), .ZN(n45944) );
  BUF_X4 U43422 ( .I(n26861), .Z(n28630) );
  NOR2_X2 U43423 ( .A1(n24039), .A2(n28410), .ZN(n28396) );
  NOR2_X2 U43424 ( .A1(n30659), .A2(n27989), .ZN(n30643) );
  BUF_X4 U43427 ( .I(n51491), .Z(n56659) );
  NAND2_X2 U43430 ( .A1(n48536), .A2(n47186), .ZN(n48232) );
  INV_X1 U43432 ( .I(n35328), .ZN(n25946) );
  NOR2_X2 U43436 ( .A1(n53729), .A2(n53740), .ZN(n53738) );
  NAND2_X2 U43438 ( .A1(n38551), .A2(n57860), .ZN(n37270) );
  NAND2_X2 U43441 ( .A1(n23298), .A2(n19990), .ZN(n40267) );
  NOR2_X2 U43446 ( .A1(n25092), .A2(n47774), .ZN(n47773) );
  NAND2_X2 U43447 ( .A1(n55569), .A2(n21272), .ZN(n55587) );
  NOR2_X2 U43450 ( .A1(n56047), .A2(n56108), .ZN(n56120) );
  INV_X4 U43451 ( .I(n55821), .ZN(n55828) );
  NAND3_X2 U43452 ( .A1(n29874), .A2(n29873), .A3(n29872), .ZN(n29875) );
  AND2_X2 U43453 ( .A1(n26956), .A2(n26955), .Z(n30558) );
  NOR2_X2 U43457 ( .A1(n54026), .A2(n51866), .ZN(n54018) );
  BUF_X4 U43459 ( .I(n52078), .Z(n55442) );
  INV_X2 U43460 ( .I(n27111), .ZN(n28378) );
  NOR2_X2 U43461 ( .A1(n42288), .A2(n21492), .ZN(n42281) );
  BUF_X2 U43463 ( .I(n52383), .Z(n54950) );
  BUF_X4 U43465 ( .I(n37725), .Z(n42259) );
  NOR2_X2 U43467 ( .A1(n14635), .A2(n54904), .ZN(n54915) );
  NAND2_X2 U43468 ( .A1(n37198), .A2(n40934), .ZN(n40939) );
  NOR2_X2 U43469 ( .A1(n45520), .A2(n45521), .ZN(n47470) );
  BUF_X4 U43471 ( .I(n37130), .Z(n26052) );
  NOR2_X2 U43472 ( .A1(n56600), .A2(n52683), .ZN(n56612) );
  INV_X4 U43474 ( .I(n65222), .ZN(n49013) );
  NOR2_X2 U43476 ( .A1(n10310), .A2(n9550), .ZN(n55153) );
  NAND2_X2 U43479 ( .A1(n55896), .A2(n22681), .ZN(n55879) );
  NAND2_X1 U43481 ( .A1(n25311), .A2(n26688), .ZN(n25310) );
  NAND2_X2 U43482 ( .A1(n41079), .A2(n40592), .ZN(n41072) );
  NAND2_X2 U43487 ( .A1(n10251), .A2(n33654), .ZN(n34137) );
  NAND2_X2 U43488 ( .A1(n40963), .A2(n61333), .ZN(n40619) );
  INV_X4 U43491 ( .I(n53078), .ZN(n53109) );
  NAND2_X1 U43494 ( .A1(n47136), .A2(n17905), .ZN(n25264) );
  XOR2_X1 U43496 ( .A1(n46658), .A2(n10443), .Z(n25273) );
  NAND2_X1 U43500 ( .A1(n37531), .A2(n60652), .ZN(n25287) );
  INV_X1 U43502 ( .I(n57128), .ZN(n57129) );
  NAND2_X1 U43503 ( .A1(n23538), .A2(n57146), .ZN(n57128) );
  XOR2_X1 U43504 ( .A1(n22478), .A2(n17336), .Z(n51506) );
  XOR2_X1 U43505 ( .A1(n22478), .A2(n50171), .Z(n50172) );
  OR2_X1 U43506 ( .A1(n37356), .A2(n22659), .Z(n25297) );
  XOR2_X1 U43507 ( .A1(Key[69]), .A2(Ciphertext[176]), .Z(n26447) );
  XOR2_X1 U43508 ( .A1(n53090), .A2(n23093), .Z(n50627) );
  XOR2_X1 U43509 ( .A1(n55368), .A2(n23093), .Z(n45404) );
  XOR2_X1 U43510 ( .A1(n56065), .A2(n23093), .Z(n35869) );
  XOR2_X1 U43511 ( .A1(n52734), .A2(n23093), .Z(n52551) );
  XOR2_X1 U43512 ( .A1(n50245), .A2(n23093), .Z(n50126) );
  XOR2_X1 U43513 ( .A1(n15712), .A2(n23093), .Z(n39360) );
  XOR2_X1 U43514 ( .A1(n46684), .A2(n23093), .Z(n33831) );
  XOR2_X1 U43515 ( .A1(n46397), .A2(n23093), .Z(n46400) );
  XOR2_X1 U43516 ( .A1(n45275), .A2(n23093), .Z(n31960) );
  XOR2_X1 U43517 ( .A1(n46245), .A2(n23093), .Z(n46248) );
  XOR2_X1 U43518 ( .A1(n44311), .A2(n23093), .Z(n51679) );
  NAND2_X1 U43519 ( .A1(n25306), .A2(n23399), .ZN(n41842) );
  XOR2_X1 U43521 ( .A1(n3499), .A2(n37460), .Z(n37461) );
  XOR2_X1 U43522 ( .A1(n32382), .A2(n32170), .Z(n30986) );
  INV_X2 U43523 ( .I(n32058), .ZN(n32170) );
  NOR2_X2 U43524 ( .A1(n25318), .A2(n25317), .ZN(n32058) );
  NOR2_X1 U43525 ( .A1(n1639), .A2(n49610), .ZN(n49594) );
  NAND2_X1 U43526 ( .A1(n1639), .A2(n17874), .ZN(n49309) );
  OAI21_X1 U43528 ( .A1(n25032), .A2(n49602), .B(n1639), .ZN(n48997) );
  AOI21_X1 U43529 ( .A1(n49608), .A2(n1639), .B(n49605), .ZN(n49311) );
  XOR2_X1 U43530 ( .A1(n4900), .A2(n43766), .Z(n45385) );
  INV_X2 U43533 ( .I(n25322), .ZN(n26182) );
  XOR2_X1 U43534 ( .A1(n31497), .A2(n30987), .Z(n25325) );
  XOR2_X1 U43537 ( .A1(n33857), .A2(n25331), .Z(n33858) );
  XOR2_X1 U43538 ( .A1(n25331), .A2(n31922), .Z(n31923) );
  NOR2_X1 U43540 ( .A1(n55292), .A2(n25336), .ZN(n55669) );
  INV_X2 U43543 ( .I(n25353), .ZN(n27494) );
  XNOR2_X1 U43544 ( .A1(Key[186]), .A2(Ciphertext[179]), .ZN(n25353) );
  INV_X2 U43545 ( .I(n22962), .ZN(n48678) );
  NAND4_X2 U43547 ( .A1(n28324), .A2(n25392), .A3(n28044), .A4(n25391), .ZN(
        n25390) );
  OR2_X1 U43550 ( .A1(n42766), .A2(n22182), .Z(n25398) );
  NOR2_X2 U43551 ( .A1(n27743), .A2(n13176), .ZN(n29729) );
  NAND4_X1 U43552 ( .A1(n27744), .A2(n28984), .A3(n4444), .A4(n25978), .ZN(
        n27746) );
  OAI22_X1 U43553 ( .A1(n28990), .A2(n25978), .B1(n23315), .B2(n30019), .ZN(
        n28991) );
  INV_X2 U43560 ( .I(n25418), .ZN(n41210) );
  XNOR2_X1 U43561 ( .A1(n25419), .A2(n25420), .ZN(n25418) );
  XOR2_X1 U43562 ( .A1(n38847), .A2(n38860), .Z(n25419) );
  XOR2_X1 U43563 ( .A1(n39673), .A2(n38855), .Z(n25422) );
  XOR2_X1 U43565 ( .A1(n25434), .A2(n26201), .Z(n25433) );
  XOR2_X1 U43566 ( .A1(n7079), .A2(n25442), .Z(n30913) );
  XOR2_X1 U43567 ( .A1(n32560), .A2(n25443), .Z(n32256) );
  XOR2_X1 U43568 ( .A1(n32325), .A2(n25443), .Z(n32328) );
  INV_X2 U43570 ( .I(n29835), .ZN(n30812) );
  XOR2_X1 U43572 ( .A1(n32587), .A2(n1823), .Z(n32588) );
  OR2_X1 U43578 ( .A1(n25456), .A2(n52847), .Z(n25462) );
  AOI21_X2 U43581 ( .A1(n45609), .A2(n45608), .B(n25474), .ZN(n45614) );
  NOR2_X1 U43582 ( .A1(n37341), .A2(n34884), .ZN(n25475) );
  INV_X2 U43584 ( .I(n47296), .ZN(n25477) );
  XOR2_X1 U43585 ( .A1(n24504), .A2(n29472), .Z(n28576) );
  NOR2_X1 U43586 ( .A1(n25494), .A2(n25493), .ZN(n25492) );
  XOR2_X1 U43590 ( .A1(n25515), .A2(n39627), .Z(n25514) );
  XOR2_X1 U43591 ( .A1(n37955), .A2(n25516), .Z(n25515) );
  XOR2_X1 U43592 ( .A1(n39208), .A2(n24058), .Z(n25516) );
  XOR2_X1 U43595 ( .A1(n32676), .A2(n31699), .Z(n25524) );
  NOR2_X1 U43596 ( .A1(n24402), .A2(n25527), .ZN(n30476) );
  OAI21_X1 U43597 ( .A1(n29528), .A2(n25527), .B(n62647), .ZN(n29529) );
  OAI21_X1 U43598 ( .A1(n29817), .A2(n30477), .B(n25527), .ZN(n25630) );
  MUX2_X1 U43599 ( .I0(n30495), .I1(n27754), .S(n19451), .Z(n27773) );
  XOR2_X1 U43601 ( .A1(n25530), .A2(n11317), .Z(n43775) );
  NOR2_X2 U43602 ( .A1(n39875), .A2(n25538), .ZN(n42993) );
  INV_X1 U43606 ( .I(n25555), .ZN(n46723) );
  INV_X2 U43607 ( .I(n25715), .ZN(n48546) );
  OR2_X2 U43609 ( .A1(n52750), .A2(n25572), .Z(n53368) );
  XOR2_X1 U43610 ( .A1(n39560), .A2(n24147), .Z(n39561) );
  NAND2_X1 U43611 ( .A1(n26714), .A2(n26717), .ZN(n25575) );
  OR2_X1 U43612 ( .A1(n36412), .A2(n36193), .Z(n25592) );
  INV_X1 U43613 ( .I(n19373), .ZN(n32993) );
  NAND3_X2 U43614 ( .A1(n46847), .A2(n46846), .A3(n46848), .ZN(n49043) );
  XOR2_X1 U43615 ( .A1(n44063), .A2(n25601), .Z(n25603) );
  XOR2_X1 U43616 ( .A1(n25602), .A2(n44062), .Z(n25601) );
  INV_X2 U43617 ( .I(n25603), .ZN(n45521) );
  INV_X2 U43618 ( .I(n15747), .ZN(n53587) );
  XOR2_X1 U43620 ( .A1(n49456), .A2(n25609), .Z(n25608) );
  XOR2_X1 U43621 ( .A1(n25610), .A2(n25061), .Z(n25609) );
  XOR2_X1 U43622 ( .A1(n22795), .A2(n49449), .Z(n25610) );
  NOR2_X2 U43624 ( .A1(n34453), .A2(n34452), .ZN(n25611) );
  NAND2_X2 U43626 ( .A1(n25616), .A2(n25620), .ZN(n30419) );
  XOR2_X1 U43628 ( .A1(n51933), .A2(n25618), .Z(n50525) );
  XOR2_X1 U43629 ( .A1(n50714), .A2(n63690), .Z(n50715) );
  XOR2_X1 U43630 ( .A1(n50108), .A2(n63690), .Z(n50109) );
  NAND3_X1 U43631 ( .A1(n7495), .A2(n23954), .A3(n25619), .ZN(n27511) );
  NOR2_X2 U43633 ( .A1(n27507), .A2(n23496), .ZN(n25619) );
  NAND2_X1 U43634 ( .A1(n826), .A2(n1956), .ZN(n49939) );
  XOR2_X1 U43635 ( .A1(n32058), .A2(n15732), .Z(n25959) );
  NOR2_X2 U43636 ( .A1(n30526), .A2(n25639), .ZN(n27922) );
  INV_X2 U43637 ( .I(n25647), .ZN(n54323) );
  NOR3_X1 U43640 ( .A1(n40034), .A2(n41844), .A3(n9627), .ZN(n42475) );
  NAND2_X1 U43641 ( .A1(n1515), .A2(n25666), .ZN(n25665) );
  NOR2_X1 U43644 ( .A1(n53493), .A2(n25675), .ZN(n53463) );
  NAND2_X1 U43645 ( .A1(n53489), .A2(n25675), .ZN(n53490) );
  NOR2_X1 U43646 ( .A1(n21922), .A2(n25675), .ZN(n53470) );
  INV_X2 U43647 ( .I(n25679), .ZN(n53905) );
  XOR2_X1 U43648 ( .A1(n25681), .A2(n55118), .Z(Plaintext[96]) );
  AND2_X1 U43649 ( .A1(n40909), .A2(n40910), .Z(n25687) );
  NAND2_X2 U43650 ( .A1(n29353), .A2(n23496), .ZN(n29340) );
  XOR2_X1 U43651 ( .A1(Key[27]), .A2(Ciphertext[170]), .Z(n27501) );
  XOR2_X1 U43653 ( .A1(n61450), .A2(n39379), .Z(n39380) );
  XOR2_X1 U43655 ( .A1(n20302), .A2(n51643), .Z(n51644) );
  XOR2_X1 U43656 ( .A1(n20302), .A2(n50609), .Z(n50610) );
  XOR2_X1 U43657 ( .A1(n25696), .A2(n25693), .Z(n25692) );
  XOR2_X1 U43658 ( .A1(n23906), .A2(n44816), .Z(n25696) );
  NAND2_X2 U43661 ( .A1(n45682), .A2(n25702), .ZN(n47590) );
  AOI21_X1 U43662 ( .A1(n22549), .A2(n47593), .B(n25702), .ZN(n45155) );
  NOR2_X1 U43663 ( .A1(n47581), .A2(n25702), .ZN(n47584) );
  OAI21_X1 U43664 ( .A1(n45680), .A2(n22549), .B(n25702), .ZN(n45681) );
  XOR2_X1 U43666 ( .A1(n25703), .A2(n56508), .Z(Plaintext[160]) );
  INV_X2 U43667 ( .I(n54793), .ZN(n55412) );
  AOI21_X1 U43668 ( .A1(n42838), .A2(n6706), .B(n42839), .ZN(n25710) );
  OR2_X1 U43669 ( .A1(n42837), .A2(n42838), .Z(n25711) );
  INV_X2 U43670 ( .I(n25714), .ZN(n48555) );
  XOR2_X1 U43673 ( .A1(n25725), .A2(n55139), .Z(Plaintext[99]) );
  NOR2_X1 U43675 ( .A1(n16042), .A2(n60020), .ZN(n25734) );
  NOR2_X1 U43676 ( .A1(n25736), .A2(n60020), .ZN(n25735) );
  INV_X1 U43677 ( .I(n28239), .ZN(n25736) );
  AND3_X1 U43678 ( .A1(n53433), .A2(n53524), .A3(n53519), .Z(n25739) );
  NOR2_X2 U43679 ( .A1(n53916), .A2(n54036), .ZN(n54049) );
  INV_X2 U43682 ( .I(n25745), .ZN(n53226) );
  INV_X1 U43683 ( .I(n53222), .ZN(n25747) );
  INV_X1 U43685 ( .I(n38677), .ZN(n41191) );
  NAND2_X2 U43687 ( .A1(n53794), .A2(n53790), .ZN(n53814) );
  NOR2_X2 U43688 ( .A1(n15928), .A2(n53823), .ZN(n53790) );
  NAND2_X2 U43689 ( .A1(n3888), .A2(n53845), .ZN(n54492) );
  NAND2_X1 U43690 ( .A1(n54640), .A2(n55017), .ZN(n25759) );
  XOR2_X1 U43693 ( .A1(n39214), .A2(n38871), .Z(n38512) );
  NAND3_X2 U43694 ( .A1(n37058), .A2(n37056), .A3(n37057), .ZN(n39214) );
  XOR2_X1 U43695 ( .A1(n22521), .A2(n10584), .Z(n51505) );
  XOR2_X1 U43696 ( .A1(n17336), .A2(n22521), .Z(n50840) );
  XOR2_X1 U43698 ( .A1(n31927), .A2(n31928), .Z(n25797) );
  INV_X4 U43699 ( .I(n14354), .ZN(n54268) );
  XOR2_X1 U43702 ( .A1(n20288), .A2(n38178), .Z(n38179) );
  XOR2_X1 U43703 ( .A1(n20288), .A2(n38477), .Z(n38478) );
  NAND2_X1 U43704 ( .A1(n34138), .A2(n32695), .ZN(n25820) );
  XOR2_X1 U43707 ( .A1(n26167), .A2(n44122), .Z(n25833) );
  XOR2_X1 U43708 ( .A1(n46621), .A2(n45327), .Z(n25835) );
  XOR2_X1 U43710 ( .A1(n44479), .A2(n44849), .Z(n44626) );
  INV_X2 U43714 ( .I(n25868), .ZN(n57017) );
  XOR2_X1 U43715 ( .A1(n50736), .A2(n51341), .Z(n50737) );
  XOR2_X1 U43716 ( .A1(n45400), .A2(n44329), .Z(n44037) );
  OAI21_X2 U43719 ( .A1(n25878), .A2(n22553), .B(n25877), .ZN(n46234) );
  AND2_X1 U43720 ( .A1(n43676), .A2(n43675), .Z(n25878) );
  XOR2_X1 U43724 ( .A1(n25887), .A2(n30042), .Z(n30043) );
  XOR2_X1 U43725 ( .A1(n25887), .A2(n32402), .Z(n32403) );
  INV_X1 U43727 ( .I(n50675), .ZN(n25894) );
  AND2_X1 U43730 ( .A1(n57149), .A2(n57159), .Z(n25906) );
  NAND2_X2 U43731 ( .A1(n25910), .A2(n25907), .ZN(n36717) );
  NAND2_X2 U43732 ( .A1(n24394), .A2(n58907), .ZN(n49566) );
  NAND2_X1 U43733 ( .A1(n31086), .A2(n31074), .ZN(n31082) );
  INV_X2 U43735 ( .I(n43453), .ZN(n44252) );
  XOR2_X1 U43736 ( .A1(n39692), .A2(n37745), .Z(n37901) );
  NOR2_X1 U43737 ( .A1(n1634), .A2(n5283), .ZN(n49037) );
  OR2_X1 U43739 ( .A1(n49061), .A2(n49060), .Z(n25931) );
  XOR2_X1 U43741 ( .A1(n50656), .A2(n23022), .Z(n51286) );
  NAND3_X2 U43742 ( .A1(n25938), .A2(n49035), .A3(n25937), .ZN(n51748) );
  NOR2_X2 U43748 ( .A1(n22939), .A2(n24024), .ZN(n43365) );
  INV_X2 U43749 ( .I(n25959), .ZN(n33898) );
  NOR2_X2 U43751 ( .A1(n38358), .A2(n38359), .ZN(n46691) );
  INV_X1 U43754 ( .I(n45110), .ZN(n25975) );
  INV_X1 U43755 ( .I(n30028), .ZN(n30031) );
  XNOR2_X1 U43756 ( .A1(n30034), .A2(n22699), .ZN(n25979) );
  INV_X2 U43757 ( .I(n61932), .ZN(n47291) );
  XOR2_X1 U43759 ( .A1(n46582), .A2(n44937), .Z(n25986) );
  XOR2_X1 U43761 ( .A1(n25991), .A2(n60514), .Z(n32735) );
  XOR2_X1 U43762 ( .A1(Ciphertext[148]), .A2(Key[65]), .Z(n28201) );
  XOR2_X1 U43763 ( .A1(n25995), .A2(n37791), .Z(n25996) );
  NAND2_X1 U43765 ( .A1(n60984), .A2(n23775), .ZN(n35033) );
  NAND2_X1 U43766 ( .A1(n25657), .A2(n23775), .ZN(n33448) );
  NAND2_X1 U43767 ( .A1(n35047), .A2(n23775), .ZN(n31300) );
  XOR2_X1 U43769 ( .A1(n56692), .A2(n61447), .Z(n30908) );
  XOR2_X1 U43770 ( .A1(n53138), .A2(n26010), .Z(n51379) );
  XOR2_X1 U43771 ( .A1(n51999), .A2(n26010), .Z(n52000) );
  XOR2_X1 U43772 ( .A1(n45348), .A2(n26010), .Z(n45350) );
  XOR2_X1 U43773 ( .A1(n50874), .A2(n26010), .Z(n38227) );
  XOR2_X1 U43774 ( .A1(n44490), .A2(n26010), .Z(n32708) );
  XOR2_X1 U43775 ( .A1(n22277), .A2(n26010), .Z(n39492) );
  XNOR2_X1 U43776 ( .A1(n43764), .A2(n19226), .ZN(n26011) );
  XOR2_X1 U43780 ( .A1(n50993), .A2(n26022), .Z(n50995) );
  XOR2_X1 U43781 ( .A1(n63018), .A2(n33162), .Z(n33163) );
  NOR2_X2 U43784 ( .A1(n34431), .A2(n34430), .ZN(n37358) );
  AND2_X1 U43785 ( .A1(n47079), .A2(n7186), .Z(n48138) );
  MUX2_X1 U43786 ( .I0(n47080), .I1(n47081), .S(n47079), .Z(n47086) );
  NOR2_X2 U43787 ( .A1(n45526), .A2(n26045), .ZN(n48411) );
  XOR2_X1 U43788 ( .A1(n26050), .A2(n26048), .Z(n33971) );
  XOR2_X1 U43789 ( .A1(n31405), .A2(n26049), .Z(n26048) );
  XOR2_X1 U43790 ( .A1(n19093), .A2(n32592), .Z(n26049) );
  NOR2_X1 U43793 ( .A1(n26591), .A2(n27530), .ZN(n26058) );
  AOI21_X1 U43794 ( .A1(n35894), .A2(n35888), .B(n35887), .ZN(n35889) );
  NAND2_X2 U43796 ( .A1(n23738), .A2(n23581), .ZN(n48445) );
  INV_X2 U43797 ( .I(n26070), .ZN(n55656) );
  AND3_X1 U43798 ( .A1(n42593), .A2(n42607), .A3(n42606), .Z(n42035) );
  NOR2_X2 U43799 ( .A1(n28492), .A2(n27841), .ZN(n28497) );
  XOR2_X1 U43800 ( .A1(n26075), .A2(n26079), .Z(n26077) );
  XOR2_X1 U43802 ( .A1(n26078), .A2(n31591), .Z(n26076) );
  XOR2_X1 U43804 ( .A1(n33192), .A2(n32592), .Z(n26080) );
  INV_X2 U43805 ( .I(n37812), .ZN(n38952) );
  XOR2_X1 U43808 ( .A1(n26087), .A2(n52466), .Z(n52467) );
  XOR2_X1 U43809 ( .A1(Ciphertext[37]), .A2(Key[152]), .Z(n26279) );
  INV_X2 U43812 ( .I(n26105), .ZN(n41162) );
  NAND2_X2 U43815 ( .A1(n31141), .A2(n30588), .ZN(n30369) );
  XOR2_X1 U43819 ( .A1(n3753), .A2(n38181), .Z(n38182) );
  XOR2_X1 U43820 ( .A1(n37556), .A2(n26121), .Z(n38181) );
  NAND2_X1 U43821 ( .A1(n41375), .A2(n22384), .ZN(n39678) );
  XOR2_X1 U43822 ( .A1(n43908), .A2(n57785), .Z(n26128) );
  XOR2_X1 U43824 ( .A1(n26134), .A2(n31461), .Z(n26133) );
  NAND2_X2 U43825 ( .A1(n30119), .A2(n30118), .ZN(n31461) );
  NAND2_X1 U43828 ( .A1(n48660), .A2(n16190), .ZN(n26139) );
  NAND2_X2 U43831 ( .A1(n41346), .A2(n41345), .ZN(n45326) );
  XOR2_X1 U43834 ( .A1(n11071), .A2(n51764), .Z(n51772) );
  XOR2_X1 U43835 ( .A1(n11071), .A2(n50979), .Z(n51159) );
  NAND2_X1 U43836 ( .A1(n26176), .A2(n45931), .ZN(n26175) );
  INV_X1 U43837 ( .I(n47292), .ZN(n26176) );
  XOR2_X1 U43838 ( .A1(Ciphertext[160]), .A2(Key[149]), .Z(n26184) );
  NOR2_X1 U43840 ( .A1(n42230), .A2(n42235), .ZN(n26196) );
  NAND2_X2 U43841 ( .A1(n39702), .A2(n39703), .ZN(n43124) );
  NOR2_X1 U43843 ( .A1(n24009), .A2(n61472), .ZN(n54454) );
  NAND3_X1 U43844 ( .A1(n54852), .A2(n1373), .A3(n61472), .ZN(n54853) );
  XOR2_X1 U43845 ( .A1(n25415), .A2(n26201), .Z(n51363) );
  OR2_X1 U43848 ( .A1(n36842), .A2(n36675), .Z(n26209) );
  INV_X2 U43850 ( .I(n26214), .ZN(n33453) );
  INV_X1 U43852 ( .I(n32234), .ZN(n31446) );
  AOI21_X1 U43853 ( .A1(n26770), .A2(n29187), .B(n26217), .ZN(n26771) );
  XOR2_X1 U43854 ( .A1(n32665), .A2(n32666), .Z(n26219) );
  NAND2_X1 U43856 ( .A1(n54807), .A2(n54806), .ZN(n54810) );
  NAND2_X2 U43860 ( .A1(n56635), .A2(n56631), .ZN(n56204) );
  NOR2_X2 U43863 ( .A1(n55170), .A2(n55165), .ZN(n55146) );
  BUF_X4 U43866 ( .I(n26922), .Z(n28858) );
  NAND2_X1 U43867 ( .A1(n27876), .A2(n28534), .ZN(n28532) );
  NOR2_X2 U43868 ( .A1(n56559), .A2(n56829), .ZN(n56660) );
  NAND2_X2 U43869 ( .A1(n52977), .A2(n53917), .ZN(n54054) );
  AOI21_X1 U43872 ( .A1(n55770), .A2(n55769), .B(n55828), .ZN(n55827) );
  INV_X1 U43873 ( .I(n55822), .ZN(n55770) );
  NAND2_X1 U43874 ( .A1(n36407), .A2(n35116), .ZN(n35120) );
  INV_X2 U43875 ( .I(n28525), .ZN(n27255) );
  NOR2_X2 U43876 ( .A1(n41042), .A2(n41041), .ZN(n41046) );
  BUF_X4 U43878 ( .I(n32691), .Z(n36494) );
  NAND4_X2 U43879 ( .A1(n32690), .A2(n32689), .A3(n32688), .A4(n32687), .ZN(
        n32691) );
  NOR2_X2 U43882 ( .A1(n26876), .A2(n26875), .ZN(n30145) );
  BUF_X4 U43884 ( .I(n53029), .Z(n53809) );
  XNOR2_X1 U43887 ( .A1(n46500), .A2(n33228), .ZN(n26237) );
  OR2_X1 U43888 ( .A1(n846), .A2(n23988), .Z(n26238) );
  AND2_X1 U43889 ( .A1(n47248), .A2(n4315), .Z(n26240) );
  OR2_X1 U43890 ( .A1(n48542), .A2(n48554), .Z(n26241) );
  AND2_X1 U43891 ( .A1(n40099), .A2(n40102), .Z(n26247) );
  OR2_X1 U43892 ( .A1(n54267), .A2(n54266), .Z(n26250) );
  OAI21_X1 U43894 ( .A1(n28518), .A2(n28517), .B(n7772), .ZN(n28519) );
  NOR2_X1 U43895 ( .A1(n27677), .A2(n27676), .ZN(n27687) );
  AOI21_X1 U43897 ( .A1(n27843), .A2(n27842), .B(n28483), .ZN(n27844) );
  OR2_X1 U43898 ( .A1(n34117), .A2(n62931), .Z(n32800) );
  NOR2_X1 U43900 ( .A1(n33798), .A2(n35653), .ZN(n35648) );
  NAND2_X1 U43901 ( .A1(n35497), .A2(n4754), .ZN(n36679) );
  INV_X1 U43902 ( .I(n38322), .ZN(n39384) );
  NAND3_X1 U43904 ( .A1(n41101), .A2(n59591), .A3(n61984), .ZN(n39503) );
  INV_X1 U43906 ( .I(n43434), .ZN(n43436) );
  NAND3_X1 U43907 ( .A1(n41297), .A2(n41296), .A3(n41295), .ZN(n41298) );
  NAND2_X1 U43908 ( .A1(n43614), .A2(n42587), .ZN(n42588) );
  NAND3_X1 U43910 ( .A1(n42609), .A2(n42608), .A3(n42607), .ZN(n42610) );
  NAND2_X1 U43912 ( .A1(n61510), .A2(n11899), .ZN(n47727) );
  NAND2_X1 U43913 ( .A1(n49760), .A2(n64), .ZN(n48888) );
  NOR2_X1 U43915 ( .A1(n49929), .A2(n49918), .ZN(n49635) );
  OAI21_X1 U43917 ( .A1(n48889), .A2(n64), .B(n48888), .ZN(n48891) );
  NAND2_X1 U43918 ( .A1(n49152), .A2(n49151), .ZN(n49157) );
  INV_X1 U43921 ( .I(n52381), .ZN(n54433) );
  OR2_X1 U43922 ( .A1(n61282), .A2(n2180), .Z(n52210) );
  OR2_X1 U43923 ( .A1(n53894), .A2(n61133), .Z(n53897) );
  NAND2_X1 U43924 ( .A1(n54606), .A2(n58994), .ZN(n54612) );
  NAND2_X1 U43928 ( .A1(n55057), .A2(n55036), .ZN(n55029) );
  OAI21_X1 U43929 ( .A1(n53493), .A2(n53514), .B(n53517), .ZN(n53468) );
  OR2_X1 U43931 ( .A1(n55816), .A2(n55801), .Z(n55809) );
  NOR2_X1 U43932 ( .A1(n53341), .A2(n53340), .ZN(n53342) );
  BUF_X2 U43935 ( .I(Key[31]), .Z(n29407) );
  OR2_X1 U43936 ( .A1(n53949), .A2(n53948), .Z(n53957) );
  NAND2_X1 U43937 ( .A1(n21154), .A2(n62128), .ZN(n26251) );
  INV_X1 U43938 ( .I(n28270), .ZN(n27402) );
  NAND3_X1 U43940 ( .A1(n60265), .A2(n28418), .A3(n14229), .ZN(n26258) );
  NOR2_X1 U43941 ( .A1(n24039), .A2(n23037), .ZN(n26260) );
  INV_X1 U43944 ( .I(Ciphertext[48]), .ZN(n26263) );
  XOR2_X1 U43945 ( .A1(n26263), .A2(Key[133]), .Z(n26264) );
  CLKBUF_X4 U43947 ( .I(Key[58]), .Z(n54185) );
  NOR2_X1 U43948 ( .A1(n28066), .A2(n28076), .ZN(n27042) );
  NAND3_X1 U43949 ( .A1(n27042), .A2(n97), .A3(n28073), .ZN(n26265) );
  INV_X1 U43950 ( .I(n27040), .ZN(n26267) );
  AOI21_X1 U43951 ( .A1(n26269), .A2(n26268), .B(n26524), .ZN(n26274) );
  NAND2_X1 U43952 ( .A1(n28239), .A2(n59102), .ZN(n26272) );
  NAND2_X1 U43953 ( .A1(n28250), .A2(n28066), .ZN(n26271) );
  XOR2_X1 U43954 ( .A1(Key[30]), .A2(Ciphertext[47]), .Z(n28040) );
  XOR2_X1 U43955 ( .A1(Key[105]), .A2(Ciphertext[44]), .Z(n26275) );
  NAND2_X2 U43956 ( .A1(n27051), .A2(n23943), .ZN(n28039) );
  INV_X1 U43958 ( .I(n27103), .ZN(n26276) );
  CLKBUF_X4 U43960 ( .I(Key[63]), .Z(n54249) );
  NAND2_X2 U43961 ( .A1(n27138), .A2(n27135), .ZN(n28318) );
  INV_X1 U43962 ( .I(n28048), .ZN(n28316) );
  NOR2_X1 U43963 ( .A1(n28316), .A2(n24837), .ZN(n26281) );
  NAND2_X1 U43964 ( .A1(n27138), .A2(n24837), .ZN(n28330) );
  INV_X1 U43965 ( .I(n28330), .ZN(n26282) );
  NOR3_X1 U43966 ( .A1(n61484), .A2(n26282), .A3(n26558), .ZN(n26283) );
  NOR2_X2 U43968 ( .A1(n26558), .A2(n26092), .ZN(n27139) );
  OAI21_X1 U43969 ( .A1(n28332), .A2(n23209), .B(n22408), .ZN(n26285) );
  MUX2_X1 U43970 ( .I0(n26557), .I1(n26285), .S(n7438), .Z(n26289) );
  AOI21_X1 U43971 ( .A1(n61317), .A2(n28043), .B(n27126), .ZN(n26288) );
  NOR2_X1 U43972 ( .A1(n26286), .A2(n27125), .ZN(n27124) );
  NOR2_X2 U43973 ( .A1(n27138), .A2(n28054), .ZN(n28321) );
  NAND2_X1 U43974 ( .A1(n27124), .A2(n28321), .ZN(n26287) );
  XOR2_X1 U43975 ( .A1(Ciphertext[24]), .A2(Ciphertext[27]), .Z(n26292) );
  XOR2_X1 U43976 ( .A1(Key[96]), .A2(Ciphertext[29]), .Z(n26293) );
  INV_X1 U43977 ( .I(Ciphertext[26]), .ZN(n26294) );
  XOR2_X1 U43978 ( .A1(n26294), .A2(Key[171]), .Z(n28362) );
  NOR2_X1 U43980 ( .A1(n28359), .A2(n58466), .ZN(n26299) );
  INV_X1 U43981 ( .I(n26614), .ZN(n26297) );
  OAI21_X1 U43982 ( .A1(n26539), .A2(n23942), .B(n26613), .ZN(n26296) );
  NOR2_X1 U43983 ( .A1(n64174), .A2(n26606), .ZN(n26301) );
  INV_X1 U43984 ( .I(n23942), .ZN(n26533) );
  INV_X1 U43986 ( .I(n26316), .ZN(n26302) );
  NAND3_X1 U43987 ( .A1(n26305), .A2(n22796), .A3(n30197), .ZN(n26307) );
  NAND2_X1 U43988 ( .A1(n30183), .A2(n1559), .ZN(n26308) );
  INV_X1 U43990 ( .I(Ciphertext[22]), .ZN(n26310) );
  NOR3_X1 U43991 ( .A1(n27565), .A2(n28378), .A3(n27109), .ZN(n26313) );
  AOI21_X1 U43993 ( .A1(n57318), .A2(n26316), .B(n27113), .ZN(n26318) );
  NOR3_X1 U43994 ( .A1(n28360), .A2(n64174), .A3(n27121), .ZN(n26317) );
  INV_X1 U43997 ( .I(n26610), .ZN(n26324) );
  NAND2_X1 U43998 ( .A1(n26540), .A2(n22604), .ZN(n26323) );
  NOR2_X1 U43999 ( .A1(n26605), .A2(n27114), .ZN(n26322) );
  NAND2_X1 U44000 ( .A1(n26539), .A2(n23942), .ZN(n26328) );
  INV_X1 U44001 ( .I(Ciphertext[16]), .ZN(n26333) );
  XOR2_X1 U44002 ( .A1(n26333), .A2(Key[101]), .Z(n26334) );
  INV_X1 U44003 ( .I(Ciphertext[14]), .ZN(n26335) );
  XOR2_X1 U44004 ( .A1(n26335), .A2(Key[87]), .Z(n26339) );
  NAND2_X1 U44005 ( .A1(n28314), .A2(n28299), .ZN(n26336) );
  INV_X2 U44006 ( .I(n27602), .ZN(n27605) );
  NAND3_X1 U44007 ( .A1(n60818), .A2(n28312), .A3(n28299), .ZN(n26337) );
  INV_X1 U44008 ( .I(Ciphertext[17]), .ZN(n26338) );
  XOR2_X1 U44009 ( .A1(n26338), .A2(Key[12]), .Z(n27172) );
  INV_X2 U44010 ( .I(n27172), .ZN(n28311) );
  INV_X1 U44011 ( .I(n27077), .ZN(n26342) );
  NOR2_X1 U44012 ( .A1(n26339), .A2(n27172), .ZN(n28313) );
  NAND2_X1 U44013 ( .A1(n28313), .A2(n28299), .ZN(n27074) );
  INV_X1 U44014 ( .I(n27074), .ZN(n26340) );
  INV_X1 U44015 ( .I(n27913), .ZN(n26370) );
  NAND2_X1 U44016 ( .A1(n27532), .A2(n28348), .ZN(n26349) );
  NOR2_X1 U44017 ( .A1(n27522), .A2(n28351), .ZN(n26353) );
  NAND2_X1 U44018 ( .A1(n27203), .A2(n27524), .ZN(n26589) );
  AOI22_X1 U44020 ( .A1(n26353), .A2(n26589), .B1(n26352), .B2(n26054), .ZN(
        n26354) );
  INV_X1 U44021 ( .I(Ciphertext[0]), .ZN(n26355) );
  INV_X1 U44022 ( .I(Ciphertext[3]), .ZN(n26356) );
  XOR2_X1 U44023 ( .A1(n26356), .A2(Key[106]), .Z(n26501) );
  INV_X1 U44024 ( .I(Ciphertext[4]), .ZN(n26357) );
  XOR2_X1 U44025 ( .A1(n26357), .A2(Key[17]), .Z(n26362) );
  INV_X1 U44026 ( .I(Ciphertext[1]), .ZN(n26358) );
  XOR2_X1 U44027 ( .A1(n26358), .A2(Key[92]), .Z(n27189) );
  NOR2_X2 U44028 ( .A1(n27567), .A2(n28106), .ZN(n26655) );
  NAND2_X1 U44029 ( .A1(n26655), .A2(n23225), .ZN(n26361) );
  XOR2_X1 U44030 ( .A1(Key[120]), .A2(Ciphertext[5]), .Z(n26360) );
  XOR2_X1 U44031 ( .A1(Key[3]), .A2(Ciphertext[2]), .Z(n27185) );
  AOI21_X1 U44032 ( .A1(n26500), .A2(n26361), .B(n22541), .ZN(n26365) );
  NOR2_X2 U44033 ( .A1(n27582), .A2(n26618), .ZN(n27568) );
  NOR2_X1 U44034 ( .A1(n27582), .A2(n23383), .ZN(n26363) );
  OAI21_X1 U44035 ( .A1(n27568), .A2(n27573), .B(n27581), .ZN(n26364) );
  INV_X1 U44036 ( .I(n26655), .ZN(n27572) );
  NAND2_X1 U44038 ( .A1(n26657), .A2(n26503), .ZN(n26366) );
  AOI21_X1 U44039 ( .A1(n26371), .A2(n29014), .B(n30082), .ZN(n26372) );
  XOR2_X1 U44040 ( .A1(Key[76]), .A2(Ciphertext[81]), .Z(n26373) );
  INV_X1 U44041 ( .I(Ciphertext[78]), .ZN(n26374) );
  XOR2_X1 U44042 ( .A1(n26374), .A2(Key[151]), .Z(n26375) );
  XOR2_X1 U44044 ( .A1(Ciphertext[86]), .A2(Key[15]), .Z(n29133) );
  CLKBUF_X4 U44045 ( .I(Key[1]), .Z(n53064) );
  NOR2_X1 U44047 ( .A1(n29132), .A2(n18231), .ZN(n26385) );
  INV_X1 U44048 ( .I(n29133), .ZN(n27298) );
  INV_X1 U44049 ( .I(n29138), .ZN(n26383) );
  INV_X1 U44050 ( .I(Ciphertext[113]), .ZN(n26386) );
  XOR2_X1 U44051 ( .A1(n26386), .A2(Key[108]), .Z(n26387) );
  XOR2_X1 U44052 ( .A1(Key[183]), .A2(Ciphertext[110]), .Z(n26388) );
  INV_X1 U44053 ( .I(Ciphertext[108]), .ZN(n26389) );
  NAND2_X1 U44054 ( .A1(n63094), .A2(n61491), .ZN(n26390) );
  AOI21_X1 U44055 ( .A1(n60542), .A2(n27839), .B(n26390), .ZN(n26396) );
  NAND2_X1 U44057 ( .A1(n61491), .A2(n60545), .ZN(n26393) );
  NOR2_X1 U44058 ( .A1(n28483), .A2(n60545), .ZN(n26400) );
  NAND2_X1 U44059 ( .A1(n27661), .A2(n1571), .ZN(n27658) );
  OAI21_X1 U44060 ( .A1(n27830), .A2(n62469), .B(n27658), .ZN(n26399) );
  AOI21_X1 U44061 ( .A1(n26400), .A2(n26399), .B(n26897), .ZN(n26401) );
  NAND3_X2 U44062 ( .A1(n26403), .A2(n26402), .A3(n26401), .ZN(n26438) );
  INV_X1 U44063 ( .I(Ciphertext[91]), .ZN(n26404) );
  XOR2_X1 U44064 ( .A1(n26404), .A2(Key[146]), .Z(n29180) );
  XOR2_X1 U44065 ( .A1(Key[57]), .A2(Ciphertext[92]), .Z(n27279) );
  INV_X2 U44066 ( .I(n29180), .ZN(n28552) );
  INV_X1 U44068 ( .I(n29189), .ZN(n26405) );
  XOR2_X1 U44069 ( .A1(Key[174]), .A2(Ciphertext[95]), .Z(n26407) );
  NAND2_X2 U44071 ( .A1(n26811), .A2(n23555), .ZN(n29187) );
  INV_X1 U44072 ( .I(n27279), .ZN(n29174) );
  NAND2_X2 U44073 ( .A1(n23555), .A2(n27283), .ZN(n28547) );
  INV_X1 U44074 ( .I(n27278), .ZN(n26408) );
  NOR2_X1 U44075 ( .A1(n29187), .A2(n4847), .ZN(n26411) );
  NAND2_X1 U44076 ( .A1(n26811), .A2(n28552), .ZN(n29175) );
  INV_X1 U44077 ( .I(n29175), .ZN(n26410) );
  NOR2_X1 U44079 ( .A1(n29191), .A2(n28550), .ZN(n26412) );
  INV_X1 U44080 ( .I(Ciphertext[107]), .ZN(n26413) );
  XOR2_X1 U44081 ( .A1(n26413), .A2(Key[66]), .Z(n26414) );
  CLKBUF_X4 U44082 ( .I(Key[52]), .Z(n53989) );
  OAI21_X1 U44084 ( .A1(n28509), .A2(n27712), .B(n26421), .ZN(n26422) );
  OAI21_X1 U44085 ( .A1(n27715), .A2(n26422), .B(n1568), .ZN(n26427) );
  NOR2_X1 U44086 ( .A1(n26423), .A2(n27717), .ZN(n26426) );
  XOR2_X1 U44088 ( .A1(Ciphertext[96]), .A2(Ciphertext[99]), .Z(n26430) );
  XOR2_X1 U44091 ( .A1(Ciphertext[100]), .A2(Key[113]), .Z(n28537) );
  INV_X1 U44092 ( .I(n26801), .ZN(n26432) );
  AOI21_X1 U44093 ( .A1(n28529), .A2(n28525), .B(n26432), .ZN(n26437) );
  XOR2_X1 U44094 ( .A1(Ciphertext[101]), .A2(Ciphertext[100]), .Z(n26434) );
  XOR2_X1 U44095 ( .A1(n23926), .A2(n55395), .Z(n26433) );
  XOR2_X1 U44096 ( .A1(n26434), .A2(n26433), .Z(n26435) );
  OAI21_X1 U44097 ( .A1(n26435), .A2(n7354), .B(n28526), .ZN(n26436) );
  NOR2_X1 U44098 ( .A1(n29957), .A2(n26439), .ZN(n26440) );
  INV_X1 U44099 ( .I(n10553), .ZN(n26444) );
  AOI21_X1 U44100 ( .A1(n7437), .A2(n26689), .B(n27219), .ZN(n26449) );
  NAND2_X1 U44101 ( .A1(n27213), .A2(n29295), .ZN(n26448) );
  INV_X1 U44102 ( .I(n26970), .ZN(n26451) );
  INV_X1 U44103 ( .I(n29296), .ZN(n26452) );
  NAND3_X1 U44104 ( .A1(n24233), .A2(n26452), .A3(n29297), .ZN(n26454) );
  NAND3_X1 U44105 ( .A1(n10324), .A2(n24947), .A3(n29297), .ZN(n26453) );
  XOR2_X1 U44106 ( .A1(Key[102]), .A2(Ciphertext[167]), .Z(n26456) );
  XOR2_X1 U44107 ( .A1(Key[163]), .A2(Ciphertext[162]), .Z(n26986) );
  INV_X1 U44108 ( .I(Ciphertext[165]), .ZN(n26455) );
  XOR2_X1 U44109 ( .A1(n26455), .A2(Key[88]), .Z(n28800) );
  INV_X1 U44111 ( .I(n26456), .ZN(n28810) );
  NOR2_X1 U44112 ( .A1(n28811), .A2(n28810), .ZN(n28804) );
  INV_X1 U44113 ( .I(n28812), .ZN(n28797) );
  INV_X1 U44115 ( .I(n27615), .ZN(n26465) );
  XOR2_X1 U44116 ( .A1(Key[153]), .A2(Ciphertext[188]), .Z(n27159) );
  MUX2_X1 U44117 ( .I0(n26597), .I1(n26460), .S(n63100), .Z(n26464) );
  INV_X1 U44118 ( .I(Ciphertext[191]), .ZN(n26458) );
  XOR2_X1 U44119 ( .A1(n26458), .A2(Key[78]), .Z(n26459) );
  NOR2_X1 U44120 ( .A1(n26670), .A2(n27619), .ZN(n26462) );
  XOR2_X1 U44121 ( .A1(Ciphertext[189]), .A2(Ciphertext[186]), .Z(n26467) );
  NOR2_X1 U44122 ( .A1(n26671), .A2(n20721), .ZN(n27429) );
  OAI22_X1 U44123 ( .A1(n26470), .A2(n57412), .B1(n27615), .B2(n22643), .ZN(
        n26471) );
  NAND2_X1 U44125 ( .A1(n27472), .A2(n23823), .ZN(n26480) );
  NAND3_X1 U44126 ( .A1(n20509), .A2(n27229), .A3(n14604), .ZN(n26479) );
  INV_X1 U44127 ( .I(n27547), .ZN(n26481) );
  NAND2_X1 U44128 ( .A1(n16788), .A2(n26481), .ZN(n26484) );
  AOI21_X1 U44129 ( .A1(n26484), .A2(n26483), .B(n20519), .ZN(n26485) );
  XOR2_X1 U44131 ( .A1(Key[144]), .A2(Ciphertext[173]), .Z(n26489) );
  INV_X1 U44132 ( .I(n27498), .ZN(n26487) );
  NAND2_X1 U44133 ( .A1(n28878), .A2(n26487), .ZN(n26491) );
  INV_X1 U44134 ( .I(Ciphertext[169]), .ZN(n26488) );
  XOR2_X1 U44135 ( .A1(n26488), .A2(Key[116]), .Z(n27499) );
  INV_X2 U44136 ( .I(n27499), .ZN(n27507) );
  INV_X2 U44137 ( .I(n26489), .ZN(n29353) );
  NAND2_X1 U44138 ( .A1(n27509), .A2(n26979), .ZN(n26490) );
  OAI22_X1 U44141 ( .A1(n26491), .A2(n26490), .B1(n29350), .B2(n26977), .ZN(
        n26496) );
  NOR2_X1 U44142 ( .A1(n14312), .A2(n19452), .ZN(n26492) );
  NAND2_X2 U44143 ( .A1(n27508), .A2(n28886), .ZN(n28884) );
  INV_X1 U44144 ( .I(n28884), .ZN(n29345) );
  INV_X1 U44145 ( .I(n29352), .ZN(n26493) );
  NAND3_X1 U44146 ( .A1(n29345), .A2(n29335), .A3(n26493), .ZN(n26494) );
  INV_X1 U44147 ( .I(n27504), .ZN(n27506) );
  NOR2_X1 U44148 ( .A1(n29352), .A2(n29340), .ZN(n26497) );
  AOI22_X1 U44150 ( .A1(n27506), .A2(n26497), .B1(n29357), .B2(n27508), .ZN(
        n26498) );
  NOR2_X1 U44151 ( .A1(n27573), .A2(n27583), .ZN(n26499) );
  OAI22_X1 U44152 ( .A1(n26653), .A2(n24001), .B1(n26618), .B2(n23071), .ZN(
        n26504) );
  NAND2_X1 U44153 ( .A1(n26504), .A2(n26503), .ZN(n26505) );
  NOR2_X1 U44154 ( .A1(n30817), .A2(n11830), .ZN(n26506) );
  NAND2_X1 U44155 ( .A1(n30812), .A2(n11830), .ZN(n26507) );
  NAND3_X1 U44156 ( .A1(n28754), .A2(n61187), .A3(n162), .ZN(n26510) );
  NAND2_X1 U44157 ( .A1(n30804), .A2(n58816), .ZN(n26509) );
  MUX2_X1 U44159 ( .I0(n26510), .I1(n26509), .S(n30807), .Z(n26511) );
  XOR2_X1 U44160 ( .A1(n31556), .A2(n50494), .Z(n31152) );
  XOR2_X1 U44161 ( .A1(n31859), .A2(n31152), .Z(n30959) );
  MUX2_X1 U44163 ( .I0(n26516), .I1(n26515), .S(n28396), .Z(n26523) );
  NOR3_X1 U44164 ( .A1(n26517), .A2(n60265), .A3(n28401), .ZN(n26521) );
  INV_X1 U44165 ( .I(n28417), .ZN(n26519) );
  AOI21_X1 U44166 ( .A1(n60768), .A2(n28073), .B(n26524), .ZN(n26526) );
  AOI22_X1 U44167 ( .A1(n27388), .A2(n27387), .B1(n26526), .B2(n26525), .ZN(
        n26530) );
  INV_X1 U44168 ( .I(n27122), .ZN(n26544) );
  NAND2_X1 U44169 ( .A1(n26536), .A2(n1895), .ZN(n26535) );
  NOR2_X1 U44170 ( .A1(n1441), .A2(n26606), .ZN(n26532) );
  OAI21_X1 U44171 ( .A1(n64174), .A2(n26533), .B(n26532), .ZN(n26534) );
  NAND3_X1 U44172 ( .A1(n26535), .A2(n1279), .A3(n26534), .ZN(n26543) );
  NOR2_X1 U44173 ( .A1(n26612), .A2(n26536), .ZN(n26537) );
  NOR2_X1 U44174 ( .A1(n28380), .A2(n22902), .ZN(n26546) );
  INV_X1 U44175 ( .I(n28384), .ZN(n26627) );
  INV_X1 U44177 ( .I(n26622), .ZN(n26548) );
  INV_X1 U44179 ( .I(n26633), .ZN(n26550) );
  NOR2_X1 U44182 ( .A1(n24836), .A2(n28049), .ZN(n27131) );
  OAI21_X1 U44183 ( .A1(n26558), .A2(n23997), .B(n26557), .ZN(n26562) );
  NOR2_X1 U44184 ( .A1(n23997), .A2(n26092), .ZN(n26559) );
  OAI21_X1 U44185 ( .A1(n27025), .A2(n26559), .B(n28333), .ZN(n26560) );
  INV_X1 U44186 ( .I(n28334), .ZN(n26564) );
  OAI21_X1 U44187 ( .A1(n61484), .A2(n28318), .B(n26564), .ZN(n26567) );
  NOR2_X1 U44188 ( .A1(n26565), .A2(n61317), .ZN(n26566) );
  NOR2_X1 U44189 ( .A1(n26568), .A2(n9685), .ZN(n26570) );
  INV_X1 U44190 ( .I(n27102), .ZN(n26574) );
  NOR2_X1 U44191 ( .A1(n26580), .A2(n27094), .ZN(n26581) );
  INV_X1 U44195 ( .I(n28344), .ZN(n26596) );
  OAI21_X1 U44196 ( .A1(n1441), .A2(n23942), .B(n22735), .ZN(n26607) );
  AOI21_X1 U44197 ( .A1(n27121), .A2(n1364), .B(n26607), .ZN(n26608) );
  NOR2_X1 U44198 ( .A1(n26608), .A2(n64174), .ZN(n26609) );
  NOR2_X1 U44199 ( .A1(n27572), .A2(n1885), .ZN(n26616) );
  OAI21_X1 U44202 ( .A1(n26629), .A2(n26628), .B(n26627), .ZN(n26630) );
  OAI21_X1 U44203 ( .A1(n26637), .A2(n26636), .B(n27560), .ZN(n26638) );
  NAND2_X1 U44204 ( .A1(n27174), .A2(n26640), .ZN(n26643) );
  AOI22_X1 U44205 ( .A1(n28313), .A2(n28306), .B1(n23840), .B2(n23324), .ZN(
        n26642) );
  OAI21_X1 U44206 ( .A1(n27598), .A2(n26643), .B(n26642), .ZN(n26649) );
  AOI21_X1 U44207 ( .A1(n27608), .A2(n26644), .B(n27594), .ZN(n26648) );
  NAND2_X1 U44208 ( .A1(n27179), .A2(n28314), .ZN(n26646) );
  AOI21_X1 U44209 ( .A1(n28311), .A2(n60818), .B(n23324), .ZN(n26645) );
  OAI22_X1 U44210 ( .A1(n26646), .A2(n22706), .B1(n26645), .B2(n19156), .ZN(
        n26647) );
  NAND2_X1 U44211 ( .A1(n29858), .A2(n29099), .ZN(n27784) );
  NOR2_X1 U44212 ( .A1(n17413), .A2(n17412), .ZN(n27782) );
  NAND3_X1 U44214 ( .A1(n27782), .A2(n29855), .A3(n740), .ZN(n26651) );
  NAND2_X1 U44215 ( .A1(n27784), .A2(n26651), .ZN(n30956) );
  INV_X1 U44216 ( .I(n27579), .ZN(n27187) );
  NAND2_X1 U44217 ( .A1(n26655), .A2(n26654), .ZN(n26658) );
  NAND3_X1 U44218 ( .A1(n24001), .A2(n10049), .A3(n23383), .ZN(n26656) );
  NOR2_X1 U44219 ( .A1(n26660), .A2(n27583), .ZN(n26663) );
  NOR2_X1 U44220 ( .A1(n1440), .A2(n23383), .ZN(n26662) );
  AOI22_X1 U44221 ( .A1(n26663), .A2(n27580), .B1(n27184), .B2(n26662), .ZN(
        n26666) );
  NOR2_X1 U44223 ( .A1(n26668), .A2(n19522), .ZN(n26677) );
  NAND2_X1 U44224 ( .A1(n26669), .A2(n27430), .ZN(n26676) );
  AOI22_X1 U44226 ( .A1(n10458), .A2(n26672), .B1(n61992), .B2(n430), .ZN(
        n26673) );
  NAND2_X1 U44227 ( .A1(n61918), .A2(n27524), .ZN(n27194) );
  NOR2_X1 U44228 ( .A1(n27194), .A2(n23835), .ZN(n26679) );
  MUX2_X1 U44229 ( .I0(n26679), .I1(n26678), .S(n28350), .Z(n26687) );
  INV_X1 U44231 ( .I(n28354), .ZN(n26685) );
  AOI21_X1 U44232 ( .A1(n20929), .A2(n296), .B(n23362), .ZN(n26683) );
  AOI21_X1 U44233 ( .A1(n26683), .A2(n27529), .B(n27204), .ZN(n26684) );
  OAI21_X1 U44235 ( .A1(n29356), .A2(n29339), .B(n29358), .ZN(n26696) );
  XOR2_X1 U44236 ( .A1(Ciphertext[171]), .A2(Ciphertext[168]), .Z(n26690) );
  INV_X1 U44237 ( .I(n29335), .ZN(n26693) );
  NOR3_X1 U44238 ( .A1(n29333), .A2(n20930), .A3(n26693), .ZN(n26695) );
  NOR2_X1 U44241 ( .A1(n27500), .A2(n29340), .ZN(n26698) );
  AOI22_X1 U44242 ( .A1(n26700), .A2(n23954), .B1(n26699), .B2(n26698), .ZN(
        n26701) );
  NOR3_X1 U44245 ( .A1(n27482), .A2(n27543), .A3(n27547), .ZN(n26704) );
  NOR2_X1 U44246 ( .A1(n27537), .A2(n27536), .ZN(n26703) );
  NOR2_X1 U44247 ( .A1(n27536), .A2(n27485), .ZN(n26706) );
  NAND2_X1 U44248 ( .A1(n29542), .A2(n26708), .ZN(n26712) );
  NAND2_X1 U44249 ( .A1(n30490), .A2(n28899), .ZN(n29541) );
  NAND2_X1 U44250 ( .A1(n27759), .A2(n62647), .ZN(n26709) );
  INV_X1 U44252 ( .I(n26714), .ZN(n26715) );
  INV_X1 U44253 ( .I(n27928), .ZN(n26721) );
  NAND2_X1 U44254 ( .A1(n26721), .A2(n60841), .ZN(n26724) );
  INV_X1 U44255 ( .I(Ciphertext[77]), .ZN(n26728) );
  XOR2_X1 U44256 ( .A1(n26728), .A2(Key[48]), .Z(n26730) );
  XOR2_X1 U44257 ( .A1(Key[123]), .A2(Ciphertext[74]), .Z(n28211) );
  INV_X1 U44258 ( .I(n22714), .ZN(n28212) );
  AOI21_X1 U44260 ( .A1(n26734), .A2(n23337), .B(n26733), .ZN(n26735) );
  NOR3_X1 U44261 ( .A1(n26735), .A2(n28504), .A3(n27853), .ZN(n26738) );
  NAND2_X1 U44262 ( .A1(n27717), .A2(n7110), .ZN(n26737) );
  NOR2_X1 U44263 ( .A1(n597), .A2(n1444), .ZN(n26741) );
  NAND2_X1 U44264 ( .A1(n65198), .A2(n26742), .ZN(n26743) );
  NAND2_X1 U44265 ( .A1(n27980), .A2(n26743), .ZN(n26744) );
  NAND2_X1 U44266 ( .A1(n26746), .A2(n26745), .ZN(n26752) );
  INV_X1 U44268 ( .I(n26764), .ZN(n26755) );
  NOR2_X1 U44269 ( .A1(n26431), .A2(n28533), .ZN(n26753) );
  OAI21_X1 U44270 ( .A1(n26755), .A2(n27869), .B(n26754), .ZN(n26760) );
  INV_X1 U44271 ( .I(n28532), .ZN(n26795) );
  NOR2_X1 U44272 ( .A1(n26764), .A2(n26795), .ZN(n26759) );
  NAND2_X1 U44273 ( .A1(n23508), .A2(n28534), .ZN(n28527) );
  INV_X1 U44274 ( .I(n28527), .ZN(n26757) );
  OAI22_X1 U44276 ( .A1(n26760), .A2(n26759), .B1(n26758), .B2(n27255), .ZN(
        n26763) );
  NAND4_X1 U44277 ( .A1(n15763), .A2(n63533), .A3(n28540), .A4(n28539), .ZN(
        n26761) );
  NAND2_X1 U44278 ( .A1(n27247), .A2(n27875), .ZN(n26769) );
  OAI21_X1 U44279 ( .A1(n27877), .A2(n28539), .B(n27871), .ZN(n26768) );
  NAND2_X1 U44280 ( .A1(n28539), .A2(n22768), .ZN(n26800) );
  NOR2_X1 U44281 ( .A1(n26800), .A2(n28533), .ZN(n26767) );
  OAI21_X1 U44282 ( .A1(n63533), .A2(n27868), .B(n28543), .ZN(n26766) );
  AOI22_X1 U44283 ( .A1(n26769), .A2(n26768), .B1(n26767), .B2(n26766), .ZN(
        n28779) );
  NOR2_X1 U44284 ( .A1(n26772), .A2(n23555), .ZN(n26773) );
  NAND2_X1 U44285 ( .A1(n26777), .A2(n61260), .ZN(n26778) );
  AOI21_X1 U44286 ( .A1(n26779), .A2(n26778), .B(n29178), .ZN(n26780) );
  NOR2_X1 U44287 ( .A1(n26781), .A2(n19461), .ZN(n26783) );
  NOR2_X1 U44288 ( .A1(n30680), .A2(n30232), .ZN(n26782) );
  INV_X1 U44289 ( .I(Ciphertext[115]), .ZN(n26784) );
  XOR2_X1 U44290 ( .A1(n26784), .A2(Key[122]), .Z(n28604) );
  NAND2_X1 U44291 ( .A1(n28615), .A2(n23649), .ZN(n27856) );
  INV_X1 U44292 ( .I(Ciphertext[118]), .ZN(n26785) );
  OAI21_X1 U44293 ( .A1(n23487), .A2(n27856), .B(n27857), .ZN(n26789) );
  INV_X1 U44295 ( .I(Ciphertext[119]), .ZN(n26786) );
  XOR2_X1 U44296 ( .A1(n26786), .A2(Key[150]), .Z(n26790) );
  INV_X1 U44297 ( .I(n26790), .ZN(n28606) );
  AOI21_X1 U44298 ( .A1(n27863), .A2(n22312), .B(n28606), .ZN(n26787) );
  NOR2_X1 U44299 ( .A1(n28616), .A2(n28607), .ZN(n26906) );
  NAND2_X1 U44301 ( .A1(n27860), .A2(n23033), .ZN(n26792) );
  NOR2_X1 U44302 ( .A1(n27857), .A2(n23649), .ZN(n28462) );
  NOR2_X1 U44303 ( .A1(n28543), .A2(n64809), .ZN(n26796) );
  NAND2_X1 U44304 ( .A1(n26797), .A2(n28540), .ZN(n27879) );
  NAND2_X1 U44305 ( .A1(n26431), .A2(n1443), .ZN(n28536) );
  INV_X1 U44306 ( .I(n28536), .ZN(n26799) );
  XOR2_X1 U44307 ( .A1(Ciphertext[86]), .A2(Ciphertext[89]), .Z(n26808) );
  CLKBUF_X4 U44308 ( .I(Key[132]), .Z(n55840) );
  XOR2_X1 U44309 ( .A1(n53272), .A2(n55840), .Z(n26807) );
  NOR2_X1 U44310 ( .A1(n29187), .A2(n28553), .ZN(n26810) );
  NOR2_X1 U44311 ( .A1(n19328), .A2(n23555), .ZN(n26813) );
  NOR2_X1 U44313 ( .A1(n28547), .A2(n21068), .ZN(n29177) );
  INV_X1 U44314 ( .I(n28557), .ZN(n26815) );
  NAND2_X1 U44315 ( .A1(n28794), .A2(n64057), .ZN(n26840) );
  INV_X1 U44316 ( .I(n26903), .ZN(n26820) );
  NAND2_X1 U44317 ( .A1(n26074), .A2(n62469), .ZN(n26819) );
  NOR3_X1 U44318 ( .A1(n26074), .A2(n27655), .A3(n27841), .ZN(n26821) );
  OAI21_X1 U44319 ( .A1(n27668), .A2(n28494), .B(n28492), .ZN(n26822) );
  OAI21_X1 U44320 ( .A1(n26822), .A2(n27832), .B(n26898), .ZN(n26833) );
  NOR2_X1 U44321 ( .A1(n28494), .A2(n27655), .ZN(n26825) );
  AOI21_X1 U44322 ( .A1(n10131), .A2(n27655), .B(n26825), .ZN(n26830) );
  INV_X1 U44323 ( .I(n27829), .ZN(n26828) );
  NOR2_X1 U44324 ( .A1(n28483), .A2(n58559), .ZN(n26827) );
  AOI21_X1 U44327 ( .A1(n26837), .A2(n26836), .B(n1568), .ZN(n26838) );
  INV_X1 U44328 ( .I(n29767), .ZN(n26841) );
  OAI21_X1 U44330 ( .A1(n28842), .A2(n23386), .B(n4812), .ZN(n26847) );
  AOI21_X1 U44331 ( .A1(n26849), .A2(n26848), .B(n26847), .ZN(n26852) );
  XOR2_X1 U44332 ( .A1(Ciphertext[141]), .A2(Ciphertext[138]), .Z(n26850) );
  AOI21_X1 U44333 ( .A1(n28594), .A2(n6513), .B(n28588), .ZN(n26851) );
  NOR2_X1 U44334 ( .A1(n26852), .A2(n26851), .ZN(n26859) );
  XOR2_X1 U44336 ( .A1(Key[61]), .A2(Ciphertext[120]), .Z(n26860) );
  XOR2_X1 U44337 ( .A1(Key[75]), .A2(Ciphertext[122]), .Z(n26861) );
  XOR2_X1 U44338 ( .A1(Key[0]), .A2(Ciphertext[125]), .Z(n26862) );
  XOR2_X1 U44339 ( .A1(Key[89]), .A2(Ciphertext[124]), .Z(n26866) );
  NOR3_X1 U44341 ( .A1(n27812), .A2(n28632), .A3(n23540), .ZN(n26863) );
  XOR2_X1 U44342 ( .A1(Key[164]), .A2(Ciphertext[121]), .Z(n28631) );
  INV_X2 U44343 ( .I(n28631), .ZN(n27691) );
  NAND2_X1 U44346 ( .A1(n28624), .A2(n27691), .ZN(n26864) );
  OAI21_X1 U44347 ( .A1(n28622), .A2(n28630), .B(n26865), .ZN(n26868) );
  NAND3_X1 U44348 ( .A1(n28471), .A2(n29712), .A3(n28624), .ZN(n26867) );
  OAI21_X1 U44350 ( .A1(n26871), .A2(n29713), .B(n29714), .ZN(n26874) );
  NOR2_X1 U44351 ( .A1(n28624), .A2(n28472), .ZN(n29710) );
  INV_X1 U44353 ( .I(n27810), .ZN(n26870) );
  AOI22_X1 U44354 ( .A1(n29712), .A2(n29710), .B1(n26870), .B2(n22648), .ZN(
        n26873) );
  NAND3_X1 U44355 ( .A1(n26874), .A2(n26873), .A3(n26872), .ZN(n26875) );
  XOR2_X1 U44356 ( .A1(Key[84]), .A2(Ciphertext[137]), .Z(n26877) );
  INV_X2 U44357 ( .I(n26877), .ZN(n29613) );
  NOR2_X2 U44358 ( .A1(n29613), .A2(n12739), .ZN(n28670) );
  NAND2_X1 U44359 ( .A1(n29618), .A2(n28670), .ZN(n26880) );
  NAND3_X1 U44360 ( .A1(n11873), .A2(n29617), .A3(n23816), .ZN(n26881) );
  AOI21_X1 U44361 ( .A1(n27693), .A2(n28176), .B(n26882), .ZN(n26892) );
  NOR2_X1 U44363 ( .A1(n28174), .A2(n11873), .ZN(n27310) );
  INV_X1 U44365 ( .I(n29614), .ZN(n26886) );
  NOR2_X1 U44366 ( .A1(n26886), .A2(n12739), .ZN(n26887) );
  AOI22_X1 U44367 ( .A1(n27310), .A2(n28172), .B1(n1567), .B2(n26887), .ZN(
        n26890) );
  NOR2_X1 U44368 ( .A1(n1567), .A2(n29610), .ZN(n26888) );
  INV_X1 U44369 ( .I(n28490), .ZN(n26895) );
  NOR3_X1 U44370 ( .A1(n10131), .A2(n27655), .A3(n26895), .ZN(n26896) );
  NOR2_X1 U44372 ( .A1(n26898), .A2(n27655), .ZN(n26900) );
  NAND2_X1 U44374 ( .A1(n28497), .A2(n61491), .ZN(n27834) );
  INV_X1 U44375 ( .I(n28436), .ZN(n28440) );
  NOR2_X2 U44376 ( .A1(n28616), .A2(n26791), .ZN(n28444) );
  INV_X1 U44377 ( .I(n26906), .ZN(n26907) );
  NOR2_X1 U44378 ( .A1(n27674), .A2(n29691), .ZN(n29683) );
  XOR2_X1 U44380 ( .A1(Ciphertext[126]), .A2(Ciphertext[129]), .Z(n26911) );
  NAND2_X1 U44381 ( .A1(n31035), .A2(n12907), .ZN(n26916) );
  NAND2_X1 U44384 ( .A1(n30705), .A2(n58430), .ZN(n26918) );
  INV_X1 U44385 ( .I(Ciphertext[157]), .ZN(n26921) );
  XOR2_X1 U44386 ( .A1(n26921), .A2(Key[32]), .Z(n26922) );
  XOR2_X1 U44387 ( .A1(Key[60]), .A2(Ciphertext[161]), .Z(n26923) );
  CLKBUF_X2 U44388 ( .I(n26923), .Z(n29321) );
  INV_X2 U44389 ( .I(n26923), .ZN(n28854) );
  INV_X1 U44390 ( .I(Ciphertext[158]), .ZN(n26924) );
  NAND2_X1 U44391 ( .A1(n28854), .A2(n29312), .ZN(n27447) );
  INV_X4 U44392 ( .I(n28858), .ZN(n29316) );
  OAI21_X1 U44393 ( .A1(n26926), .A2(n27447), .B(n26925), .ZN(n26934) );
  NAND2_X1 U44394 ( .A1(n64451), .A2(n29316), .ZN(n26927) );
  AOI21_X1 U44395 ( .A1(n26929), .A2(n26927), .B(n28854), .ZN(n26933) );
  NAND2_X1 U44396 ( .A1(n19972), .A2(n28854), .ZN(n26928) );
  AOI21_X1 U44397 ( .A1(n26929), .A2(n26928), .B(n27449), .ZN(n26932) );
  INV_X1 U44399 ( .I(n27451), .ZN(n29324) );
  NAND2_X1 U44400 ( .A1(n29324), .A2(n19972), .ZN(n26930) );
  OAI22_X1 U44401 ( .A1(n27450), .A2(n26930), .B1(n29319), .B2(n20093), .ZN(
        n26931) );
  OAI21_X1 U44402 ( .A1(n15779), .A2(n25786), .B(n27538), .ZN(n26941) );
  INV_X1 U44405 ( .I(n28571), .ZN(n26957) );
  INV_X1 U44406 ( .I(Ciphertext[154]), .ZN(n26942) );
  XOR2_X1 U44407 ( .A1(Ciphertext[153]), .A2(Key[4]), .Z(n29623) );
  INV_X1 U44409 ( .I(Ciphertext[155]), .ZN(n26944) );
  XOR2_X1 U44410 ( .A1(n26944), .A2(Key[18]), .Z(n26945) );
  NAND2_X1 U44411 ( .A1(n10198), .A2(n29628), .ZN(n28120) );
  NAND2_X2 U44412 ( .A1(n28119), .A2(n28831), .ZN(n29286) );
  NAND2_X1 U44413 ( .A1(n28120), .A2(n29286), .ZN(n26946) );
  XOR2_X1 U44416 ( .A1(Ciphertext[153]), .A2(Ciphertext[150]), .Z(n26952) );
  XOR2_X1 U44417 ( .A1(n59130), .A2(Key[79]), .Z(n26951) );
  INV_X1 U44418 ( .I(n29291), .ZN(n26954) );
  NAND2_X1 U44419 ( .A1(n28825), .A2(n28831), .ZN(n28827) );
  INV_X1 U44420 ( .I(n28827), .ZN(n26953) );
  OAI21_X1 U44421 ( .A1(n26954), .A2(n28835), .B(n26953), .ZN(n26955) );
  INV_X1 U44422 ( .I(n26965), .ZN(n26966) );
  INV_X1 U44423 ( .I(n27493), .ZN(n27224) );
  AOI21_X1 U44424 ( .A1(n26972), .A2(n27213), .B(n26971), .ZN(n26973) );
  OAI21_X1 U44425 ( .A1(n23496), .A2(n29356), .B(n29357), .ZN(n26976) );
  NAND3_X1 U44426 ( .A1(n29351), .A2(n7495), .A3(n29335), .ZN(n26975) );
  AOI21_X1 U44427 ( .A1(n26976), .A2(n26975), .B(n26974), .ZN(n26985) );
  INV_X1 U44428 ( .I(n26977), .ZN(n26978) );
  INV_X1 U44430 ( .I(n26979), .ZN(n26980) );
  OAI21_X1 U44431 ( .A1(n26980), .A2(n10403), .B(n20930), .ZN(n26981) );
  NAND3_X1 U44432 ( .A1(n26981), .A2(n23954), .A3(n29350), .ZN(n26983) );
  NOR2_X1 U44433 ( .A1(n29338), .A2(n23954), .ZN(n28879) );
  NAND2_X1 U44434 ( .A1(n28879), .A2(n7495), .ZN(n26982) );
  INV_X1 U44435 ( .I(n29474), .ZN(n27001) );
  INV_X1 U44436 ( .I(n28815), .ZN(n26987) );
  OAI21_X1 U44437 ( .A1(n26987), .A2(n28813), .B(n17633), .ZN(n26989) );
  NAND3_X1 U44438 ( .A1(n17633), .A2(n23824), .A3(n22158), .ZN(n26988) );
  AOI21_X1 U44439 ( .A1(n17879), .A2(n23479), .B(n28802), .ZN(n26993) );
  NAND2_X1 U44440 ( .A1(n26993), .A2(n26992), .ZN(n26999) );
  NOR2_X1 U44441 ( .A1(n28812), .A2(n26994), .ZN(n27436) );
  NAND2_X1 U44444 ( .A1(n31076), .A2(n31088), .ZN(n27005) );
  NAND3_X1 U44446 ( .A1(n5267), .A2(n31083), .A3(n22878), .ZN(n27004) );
  XOR2_X1 U44448 ( .A1(n32722), .A2(n63955), .Z(n31928) );
  INV_X1 U44449 ( .I(n31928), .ZN(n27007) );
  NAND2_X1 U44451 ( .A1(n27374), .A2(n23716), .ZN(n27010) );
  INV_X2 U44452 ( .I(n27378), .ZN(n28225) );
  XOR2_X1 U44453 ( .A1(Ciphertext[60]), .A2(Ciphertext[63]), .Z(n27013) );
  NOR2_X1 U44456 ( .A1(n61317), .A2(n28049), .ZN(n27024) );
  INV_X1 U44457 ( .I(Ciphertext[68]), .ZN(n27027) );
  CLKBUF_X4 U44458 ( .I(Key[81]), .Z(n54734) );
  XOR2_X1 U44459 ( .A1(n27027), .A2(Key[81]), .Z(n27033) );
  INV_X2 U44460 ( .I(n27033), .ZN(n28259) );
  XOR2_X1 U44461 ( .A1(Key[6]), .A2(Ciphertext[71]), .Z(n29167) );
  NOR3_X1 U44462 ( .A1(n27028), .A2(n64012), .A3(n23769), .ZN(n27032) );
  NAND2_X1 U44463 ( .A1(n29163), .A2(n27285), .ZN(n27029) );
  OAI22_X1 U44464 ( .A1(n21086), .A2(n6083), .B1(n27936), .B2(n29161), .ZN(
        n27030) );
  NAND2_X1 U44467 ( .A1(n27037), .A2(n28240), .ZN(n27038) );
  NOR2_X1 U44470 ( .A1(n28067), .A2(n23586), .ZN(n27043) );
  NOR3_X1 U44472 ( .A1(n27047), .A2(n27098), .A3(n14583), .ZN(n27050) );
  NAND2_X1 U44473 ( .A1(n23943), .A2(n28035), .ZN(n27048) );
  OAI22_X1 U44474 ( .A1(n61643), .A2(n27048), .B1(n28039), .B2(n22203), .ZN(
        n27049) );
  NOR2_X1 U44475 ( .A1(n27050), .A2(n27049), .ZN(n27060) );
  AOI21_X1 U44476 ( .A1(n28031), .A2(n28039), .B(n61643), .ZN(n27054) );
  AOI21_X1 U44477 ( .A1(n28033), .A2(n20753), .B(n27051), .ZN(n27052) );
  NAND2_X1 U44478 ( .A1(n27054), .A2(n27053), .ZN(n27059) );
  NAND3_X2 U44480 ( .A1(n27060), .A2(n27059), .A3(n27058), .ZN(n29726) );
  NAND3_X1 U44481 ( .A1(n28278), .A2(n62631), .A3(n27404), .ZN(n27064) );
  NAND2_X1 U44482 ( .A1(n27065), .A2(n61035), .ZN(n27066) );
  NOR3_X1 U44483 ( .A1(n28026), .A2(n21946), .A3(n60885), .ZN(n27067) );
  NAND2_X1 U44486 ( .A1(n61753), .A2(n30027), .ZN(n27072) );
  OAI22_X1 U44487 ( .A1(n27074), .A2(n27595), .B1(n27178), .B2(n27602), .ZN(
        n27075) );
  NAND2_X1 U44489 ( .A1(n27600), .A2(n27168), .ZN(n27076) );
  NAND2_X1 U44490 ( .A1(n27077), .A2(n27076), .ZN(n27083) );
  INV_X1 U44491 ( .I(n27595), .ZN(n27078) );
  NAND2_X1 U44492 ( .A1(n27174), .A2(n27078), .ZN(n27079) );
  AOI21_X1 U44493 ( .A1(n27079), .A2(n27168), .B(n27592), .ZN(n27081) );
  NOR2_X1 U44495 ( .A1(n28007), .A2(n28396), .ZN(n27091) );
  NOR3_X1 U44498 ( .A1(n28231), .A2(n27095), .A3(n27094), .ZN(n27096) );
  AOI21_X1 U44499 ( .A1(n60355), .A2(n28035), .B(n61177), .ZN(n27099) );
  NOR2_X1 U44500 ( .A1(n28379), .A2(n23007), .ZN(n27106) );
  NAND2_X1 U44501 ( .A1(n23191), .A2(n64174), .ZN(n27115) );
  OAI21_X1 U44503 ( .A1(n27124), .A2(n28335), .B(n27123), .ZN(n27129) );
  OAI21_X1 U44504 ( .A1(n27127), .A2(n27126), .B(n28321), .ZN(n27128) );
  NAND2_X1 U44505 ( .A1(n27129), .A2(n27128), .ZN(n27147) );
  AOI22_X1 U44506 ( .A1(n28053), .A2(n61484), .B1(n28332), .B2(n22408), .ZN(
        n27133) );
  NAND2_X1 U44507 ( .A1(n27138), .A2(n23997), .ZN(n27132) );
  NOR2_X1 U44508 ( .A1(n28327), .A2(n24837), .ZN(n27137) );
  NOR2_X1 U44513 ( .A1(n25096), .A2(n27150), .ZN(n27149) );
  INV_X1 U44515 ( .I(n29440), .ZN(n29435) );
  NAND2_X1 U44516 ( .A1(n29435), .A2(n29442), .ZN(n27151) );
  XOR2_X1 U44517 ( .A1(n23926), .A2(n52226), .Z(n37878) );
  XOR2_X1 U44518 ( .A1(n55335), .A2(n55840), .Z(n27154) );
  BUF_X2 U44519 ( .I(n27154), .Z(n51494) );
  XOR2_X1 U44520 ( .A1(n37878), .A2(n51494), .Z(n32040) );
  XOR2_X1 U44521 ( .A1(n32040), .A2(n52900), .Z(n36147) );
  XOR2_X1 U44522 ( .A1(n54517), .A2(n55118), .Z(n27155) );
  BUF_X2 U44523 ( .I(n27155), .Z(n39478) );
  XOR2_X1 U44524 ( .A1(n54870), .A2(n20814), .Z(n37303) );
  XOR2_X1 U44525 ( .A1(n39478), .A2(n37303), .Z(n32232) );
  INV_X1 U44526 ( .I(n238), .ZN(n27156) );
  XOR2_X1 U44527 ( .A1(n36147), .A2(n27156), .Z(n50836) );
  XOR2_X1 U44528 ( .A1(n24044), .A2(n24105), .Z(n38826) );
  XOR2_X1 U44529 ( .A1(n50836), .A2(n38826), .Z(n44751) );
  XOR2_X1 U44530 ( .A1(n54126), .A2(n54676), .Z(n44995) );
  XOR2_X1 U44532 ( .A1(n54360), .A2(n53772), .Z(n38699) );
  XOR2_X1 U44533 ( .A1(n44995), .A2(n63603), .Z(n35521) );
  XOR2_X1 U44534 ( .A1(n35521), .A2(n24014), .Z(n40919) );
  XOR2_X1 U44535 ( .A1(n52970), .A2(n51492), .Z(n39377) );
  XOR2_X1 U44536 ( .A1(n40919), .A2(n39377), .Z(n27157) );
  XOR2_X1 U44537 ( .A1(n44751), .A2(n27157), .Z(n27158) );
  XOR2_X1 U44538 ( .A1(n59546), .A2(n27158), .Z(n27309) );
  OAI22_X1 U44539 ( .A1(n57412), .A2(n27615), .B1(n11850), .B2(n27163), .ZN(
        n27164) );
  INV_X1 U44540 ( .I(n27613), .ZN(n27165) );
  NAND2_X1 U44541 ( .A1(n27168), .A2(n27606), .ZN(n27170) );
  NOR2_X1 U44542 ( .A1(n28312), .A2(n23636), .ZN(n28305) );
  NAND2_X1 U44543 ( .A1(n26339), .A2(n27172), .ZN(n27609) );
  INV_X1 U44544 ( .I(n27609), .ZN(n27173) );
  NAND3_X1 U44545 ( .A1(n27174), .A2(n28313), .A3(n27605), .ZN(n27175) );
  NOR2_X1 U44546 ( .A1(n23328), .A2(n23636), .ZN(n27177) );
  INV_X1 U44547 ( .I(n27180), .ZN(n27182) );
  NOR2_X1 U44548 ( .A1(n27577), .A2(n23071), .ZN(n27181) );
  NOR2_X1 U44549 ( .A1(n24001), .A2(n23225), .ZN(n27183) );
  NAND2_X1 U44550 ( .A1(n1572), .A2(n27183), .ZN(n28105) );
  INV_X1 U44551 ( .I(n28107), .ZN(n27190) );
  OAI21_X1 U44552 ( .A1(n27190), .A2(n10049), .B(n61320), .ZN(n27191) );
  NAND2_X1 U44553 ( .A1(n28350), .A2(n23362), .ZN(n27195) );
  AOI21_X1 U44554 ( .A1(n27532), .A2(n296), .B(n28350), .ZN(n27198) );
  NOR2_X1 U44555 ( .A1(n27198), .A2(n27197), .ZN(n27199) );
  NOR2_X1 U44556 ( .A1(n28342), .A2(n27529), .ZN(n27201) );
  NOR2_X1 U44557 ( .A1(n27203), .A2(n23835), .ZN(n28340) );
  INV_X1 U44558 ( .I(n28340), .ZN(n27205) );
  OAI22_X1 U44559 ( .A1(n27207), .A2(n27206), .B1(n27205), .B2(n27204), .ZN(
        n27212) );
  NAND2_X1 U44560 ( .A1(n27532), .A2(n27523), .ZN(n27209) );
  INV_X1 U44561 ( .I(n28351), .ZN(n27208) );
  OAI22_X1 U44562 ( .A1(n27210), .A2(n24735), .B1(n27209), .B2(n27208), .ZN(
        n27211) );
  AOI21_X1 U44563 ( .A1(n29295), .A2(n24947), .B(n27219), .ZN(n27216) );
  NAND2_X1 U44564 ( .A1(n27218), .A2(n27217), .ZN(n27221) );
  AOI21_X1 U44565 ( .A1(n27221), .A2(n27496), .B(n27220), .ZN(n27222) );
  NAND2_X1 U44566 ( .A1(n27229), .A2(n27228), .ZN(n27230) );
  INV_X1 U44567 ( .I(n29838), .ZN(n27238) );
  NAND2_X1 U44568 ( .A1(n29460), .A2(n27238), .ZN(n27239) );
  NAND2_X1 U44569 ( .A1(n7405), .A2(n29452), .ZN(n28733) );
  INV_X1 U44570 ( .I(n27240), .ZN(n27243) );
  INV_X1 U44571 ( .I(n27241), .ZN(n27242) );
  NOR2_X1 U44572 ( .A1(n28115), .A2(n12632), .ZN(n27244) );
  AOI22_X1 U44573 ( .A1(n27245), .A2(n28733), .B1(n29840), .B2(n27244), .ZN(
        n27246) );
  OAI21_X1 U44575 ( .A1(n28526), .A2(n27868), .B(n27869), .ZN(n27248) );
  NAND2_X1 U44577 ( .A1(n1443), .A2(n28533), .ZN(n27250) );
  AOI21_X1 U44581 ( .A1(n27260), .A2(n27259), .B(n29151), .ZN(n27261) );
  INV_X1 U44582 ( .I(n27985), .ZN(n27266) );
  NOR2_X1 U44583 ( .A1(n28557), .A2(n4847), .ZN(n27272) );
  INV_X1 U44585 ( .I(n27273), .ZN(n27275) );
  NOR3_X1 U44586 ( .A1(n27275), .A2(n19328), .A3(n27274), .ZN(n27276) );
  NAND2_X1 U44587 ( .A1(n28552), .A2(n23555), .ZN(n27280) );
  NAND4_X1 U44588 ( .A1(n28549), .A2(n4847), .A3(n19328), .A4(n20782), .ZN(
        n27284) );
  NAND2_X1 U44589 ( .A1(n27285), .A2(n11514), .ZN(n27939) );
  AOI21_X1 U44590 ( .A1(n27419), .A2(n27939), .B(n1878), .ZN(n27290) );
  NOR2_X1 U44592 ( .A1(n29132), .A2(n27292), .ZN(n27291) );
  AOI21_X1 U44594 ( .A1(n27299), .A2(n7371), .B(n27932), .ZN(n27300) );
  AOI21_X1 U44595 ( .A1(n27302), .A2(n27301), .B(n27300), .ZN(n27303) );
  XOR2_X1 U44597 ( .A1(n33033), .A2(n27309), .Z(n27629) );
  AOI21_X1 U44598 ( .A1(n59099), .A2(n29609), .B(n27310), .ZN(n27312) );
  NAND2_X1 U44599 ( .A1(n64145), .A2(n12739), .ZN(n27311) );
  NOR2_X1 U44600 ( .A1(n28174), .A2(n28175), .ZN(n27313) );
  NAND2_X1 U44601 ( .A1(n19290), .A2(n28127), .ZN(n27320) );
  NAND2_X1 U44602 ( .A1(n29285), .A2(n28831), .ZN(n27321) );
  NAND2_X1 U44603 ( .A1(n28810), .A2(n23773), .ZN(n27325) );
  AOI21_X1 U44604 ( .A1(n28802), .A2(n27325), .B(n23479), .ZN(n27326) );
  NAND2_X1 U44606 ( .A1(n28809), .A2(n23824), .ZN(n27332) );
  NOR2_X1 U44607 ( .A1(n27328), .A2(n28810), .ZN(n27330) );
  XOR2_X1 U44608 ( .A1(Key[51]), .A2(Ciphertext[146]), .Z(n27336) );
  NOR2_X1 U44609 ( .A1(n29671), .A2(n20240), .ZN(n28195) );
  XOR2_X1 U44610 ( .A1(Key[168]), .A2(Ciphertext[149]), .Z(n28192) );
  OAI21_X1 U44611 ( .A1(n1356), .A2(n28195), .B(n29660), .ZN(n27340) );
  NAND3_X1 U44612 ( .A1(n27340), .A2(n57781), .A3(n29658), .ZN(n27344) );
  NAND2_X1 U44613 ( .A1(n29384), .A2(n57781), .ZN(n27341) );
  NAND2_X1 U44614 ( .A1(n29643), .A2(n20907), .ZN(n28151) );
  AOI21_X1 U44615 ( .A1(n59935), .A2(n29638), .B(n27346), .ZN(n27353) );
  NAND2_X1 U44616 ( .A1(n28847), .A2(n28596), .ZN(n27348) );
  NOR2_X1 U44617 ( .A1(n61004), .A2(n20907), .ZN(n27347) );
  OAI21_X1 U44618 ( .A1(n27348), .A2(n27347), .B(n29634), .ZN(n27351) );
  NAND2_X1 U44619 ( .A1(n61004), .A2(n4812), .ZN(n27349) );
  NAND2_X1 U44621 ( .A1(n30174), .A2(n17627), .ZN(n27354) );
  INV_X1 U44624 ( .I(n27448), .ZN(n27356) );
  NAND4_X1 U44625 ( .A1(n27356), .A2(n58108), .A3(n28854), .A4(n19967), .ZN(
        n27357) );
  NOR2_X1 U44626 ( .A1(n27360), .A2(n23797), .ZN(n27358) );
  CLKBUF_X4 U44627 ( .I(Key[46]), .Z(n53833) );
  INV_X1 U44628 ( .I(n28003), .ZN(n27368) );
  NAND2_X1 U44629 ( .A1(n24060), .A2(n23166), .ZN(n27367) );
  AOI21_X1 U44630 ( .A1(n27370), .A2(n19170), .B(n5627), .ZN(n27372) );
  NAND2_X1 U44631 ( .A1(n27370), .A2(n29106), .ZN(n27371) );
  NAND3_X1 U44632 ( .A1(n28222), .A2(n63850), .A3(n10404), .ZN(n27377) );
  NAND2_X1 U44633 ( .A1(n27378), .A2(n29105), .ZN(n29109) );
  NOR2_X1 U44634 ( .A1(n28220), .A2(n28222), .ZN(n27379) );
  NAND3_X1 U44636 ( .A1(n27980), .A2(n29155), .A3(n27392), .ZN(n27395) );
  INV_X1 U44638 ( .I(n27977), .ZN(n27398) );
  INV_X1 U44639 ( .I(n28277), .ZN(n27400) );
  NOR2_X1 U44640 ( .A1(n29119), .A2(n28211), .ZN(n29124) );
  INV_X1 U44641 ( .I(n29129), .ZN(n27407) );
  NOR2_X1 U44642 ( .A1(n29124), .A2(n27410), .ZN(n27411) );
  NAND3_X1 U44643 ( .A1(n29162), .A2(n1359), .A3(n28260), .ZN(n27415) );
  NOR2_X1 U44644 ( .A1(n29168), .A2(n11514), .ZN(n27421) );
  NOR2_X1 U44645 ( .A1(n30250), .A2(n22014), .ZN(n27422) );
  NOR3_X1 U44647 ( .A1(n30252), .A2(n8602), .A3(n12164), .ZN(n27424) );
  INV_X1 U44648 ( .I(n29054), .ZN(n27425) );
  OAI21_X1 U44649 ( .A1(n19122), .A2(n22952), .B(n27431), .ZN(n27432) );
  AOI21_X1 U44652 ( .A1(n28813), .A2(n27441), .B(n29372), .ZN(n27443) );
  NOR2_X1 U44653 ( .A1(n29311), .A2(n27454), .ZN(n28850) );
  NOR2_X1 U44654 ( .A1(n28855), .A2(n28860), .ZN(n29327) );
  OAI21_X1 U44655 ( .A1(n28850), .A2(n29327), .B(n1884), .ZN(n27459) );
  INV_X1 U44658 ( .I(n27471), .ZN(n27467) );
  OAI21_X1 U44659 ( .A1(n27464), .A2(n14604), .B(n27546), .ZN(n27465) );
  INV_X1 U44661 ( .I(n27538), .ZN(n27469) );
  NAND2_X1 U44662 ( .A1(n27472), .A2(n27471), .ZN(n27473) );
  NAND3_X1 U44663 ( .A1(n23823), .A2(n25793), .A3(n27485), .ZN(n27481) );
  NAND2_X1 U44664 ( .A1(n27482), .A2(n27485), .ZN(n27484) );
  NOR3_X1 U44665 ( .A1(n27543), .A2(n27486), .A3(n27485), .ZN(n27487) );
  INV_X1 U44666 ( .I(n27491), .ZN(n27492) );
  NAND2_X1 U44667 ( .A1(n29292), .A2(n27494), .ZN(n27495) );
  NAND2_X1 U44668 ( .A1(n29303), .A2(n63883), .ZN(n27497) );
  NAND2_X1 U44670 ( .A1(n28883), .A2(n27498), .ZN(n27505) );
  AOI21_X1 U44671 ( .A1(n27500), .A2(n23822), .B(n23496), .ZN(n27503) );
  INV_X1 U44672 ( .I(n23496), .ZN(n29355) );
  OAI21_X1 U44673 ( .A1(n23954), .A2(n29355), .B(n19452), .ZN(n27502) );
  OAI22_X1 U44674 ( .A1(n27505), .A2(n27504), .B1(n27503), .B2(n27502), .ZN(
        n27514) );
  NAND4_X1 U44676 ( .A1(n28884), .A2(n27510), .A3(n27509), .A4(n19452), .ZN(
        n27512) );
  NOR2_X1 U44677 ( .A1(n28773), .A2(n29220), .ZN(n27517) );
  AOI22_X1 U44679 ( .A1(n30731), .A2(n27518), .B1(n27517), .B2(n29039), .ZN(
        n27519) );
  INV_X1 U44680 ( .I(n27520), .ZN(n27521) );
  NOR3_X1 U44681 ( .A1(n28341), .A2(n27521), .A3(n27526), .ZN(n27528) );
  OAI21_X1 U44682 ( .A1(n26054), .A2(n27523), .B(n27522), .ZN(n27527) );
  OAI21_X1 U44683 ( .A1(n27528), .A2(n27527), .B(n16101), .ZN(n27535) );
  AOI22_X1 U44685 ( .A1(n7974), .A2(n28351), .B1(n27531), .B2(n27530), .ZN(
        n27534) );
  NOR3_X1 U44686 ( .A1(n27543), .A2(n27537), .A3(n27536), .ZN(n27541) );
  NOR2_X1 U44687 ( .A1(n27543), .A2(n27547), .ZN(n27545) );
  AOI21_X1 U44688 ( .A1(n27545), .A2(n16788), .B(n27544), .ZN(n27552) );
  AOI21_X1 U44689 ( .A1(n27548), .A2(n27547), .B(n27546), .ZN(n27549) );
  INV_X1 U44690 ( .I(n27556), .ZN(n27557) );
  AOI21_X1 U44691 ( .A1(n27558), .A2(n27557), .B(n10321), .ZN(n27564) );
  NOR2_X1 U44693 ( .A1(n18751), .A2(n27560), .ZN(n27561) );
  NOR2_X1 U44694 ( .A1(n27568), .A2(n23071), .ZN(n27570) );
  OAI22_X1 U44695 ( .A1(n27573), .A2(n1354), .B1(n27572), .B2(n1440), .ZN(
        n27578) );
  NAND2_X1 U44696 ( .A1(n23225), .A2(n23071), .ZN(n27575) );
  OAI22_X1 U44697 ( .A1(n28107), .A2(n27575), .B1(n27583), .B2(n23071), .ZN(
        n27576) );
  NOR2_X1 U44699 ( .A1(n27583), .A2(n7477), .ZN(n27584) );
  AOI22_X1 U44700 ( .A1(n27594), .A2(n28314), .B1(n27609), .B2(n27593), .ZN(
        n27596) );
  NOR2_X1 U44701 ( .A1(n27596), .A2(n27595), .ZN(n27599) );
  INV_X1 U44702 ( .I(n28314), .ZN(n27607) );
  NAND2_X1 U44703 ( .A1(n14063), .A2(n29779), .ZN(n27610) );
  NAND2_X1 U44704 ( .A1(n13672), .A2(n27611), .ZN(n27612) );
  NOR2_X1 U44705 ( .A1(n27615), .A2(n27614), .ZN(n27617) );
  NAND2_X1 U44707 ( .A1(n10914), .A2(n22643), .ZN(n27623) );
  XOR2_X1 U44710 ( .A1(n27629), .A2(n32003), .Z(n27630) );
  AOI21_X1 U44711 ( .A1(n27634), .A2(n29508), .B(n29008), .ZN(n27637) );
  XOR2_X1 U44713 ( .A1(Key[189]), .A2(n58084), .Z(n27640) );
  XOR2_X1 U44714 ( .A1(n27640), .A2(n24051), .Z(n46348) );
  NOR2_X1 U44715 ( .A1(n28444), .A2(n22312), .ZN(n27641) );
  AOI21_X1 U44716 ( .A1(n27642), .A2(n27641), .B(n28436), .ZN(n27649) );
  NOR2_X1 U44718 ( .A1(n23033), .A2(n10544), .ZN(n27643) );
  NOR2_X1 U44719 ( .A1(n27644), .A2(n27643), .ZN(n27648) );
  NOR2_X1 U44720 ( .A1(n28434), .A2(n28452), .ZN(n27646) );
  AOI21_X1 U44721 ( .A1(n28605), .A2(n27646), .B(n28613), .ZN(n27647) );
  AOI21_X1 U44722 ( .A1(n28451), .A2(n28453), .B(n10085), .ZN(n27653) );
  INV_X1 U44723 ( .I(n27664), .ZN(n27656) );
  INV_X1 U44724 ( .I(n27658), .ZN(n27660) );
  NAND2_X1 U44725 ( .A1(n22721), .A2(n28483), .ZN(n28499) );
  OAI22_X1 U44726 ( .A1(n27664), .A2(n28494), .B1(n27668), .B2(n27839), .ZN(
        n27671) );
  NOR2_X1 U44727 ( .A1(n28485), .A2(n60545), .ZN(n27666) );
  NOR2_X1 U44728 ( .A1(n62270), .A2(n27666), .ZN(n27670) );
  NAND2_X1 U44729 ( .A1(n27668), .A2(n27841), .ZN(n27669) );
  NAND2_X2 U44731 ( .A1(n27673), .A2(n27672), .ZN(n29010) );
  NOR2_X1 U44732 ( .A1(n28653), .A2(n60547), .ZN(n27676) );
  NOR3_X1 U44733 ( .A1(n29694), .A2(n491), .A3(n27892), .ZN(n27681) );
  NOR3_X1 U44734 ( .A1(n27892), .A2(n27679), .A3(n10473), .ZN(n27680) );
  NAND2_X1 U44737 ( .A1(n28624), .A2(n26861), .ZN(n28469) );
  NAND2_X1 U44738 ( .A1(n63495), .A2(n28632), .ZN(n27689) );
  NAND2_X1 U44739 ( .A1(n27691), .A2(n28632), .ZN(n28623) );
  NAND2_X1 U44740 ( .A1(n28674), .A2(n27692), .ZN(n27697) );
  NOR2_X1 U44741 ( .A1(n28669), .A2(n24052), .ZN(n27704) );
  INV_X1 U44742 ( .I(n28676), .ZN(n27699) );
  OAI21_X1 U44743 ( .A1(n28669), .A2(n27699), .B(n27698), .ZN(n27703) );
  NOR2_X1 U44745 ( .A1(n29605), .A2(n29609), .ZN(n27701) );
  AOI22_X1 U44746 ( .A1(n27701), .A2(n264), .B1(n27700), .B2(n28172), .ZN(
        n27702) );
  OAI21_X1 U44747 ( .A1(n27704), .A2(n27703), .B(n27702), .ZN(n27705) );
  NOR2_X1 U44749 ( .A1(n23337), .A2(n28504), .ZN(n27852) );
  INV_X1 U44751 ( .I(n27851), .ZN(n27713) );
  AOI21_X1 U44754 ( .A1(n30588), .A2(n30375), .B(n1843), .ZN(n27725) );
  AOI21_X1 U44755 ( .A1(n29481), .A2(n30369), .B(n27727), .ZN(n27729) );
  OAI21_X1 U44759 ( .A1(n28989), .A2(n28988), .B(n61753), .ZN(n27741) );
  NOR2_X1 U44760 ( .A1(n4444), .A2(n22748), .ZN(n27740) );
  NOR2_X1 U44761 ( .A1(n29727), .A2(n1192), .ZN(n28984) );
  NAND2_X1 U44762 ( .A1(n25898), .A2(n23315), .ZN(n27744) );
  NAND2_X1 U44764 ( .A1(n27748), .A2(n4444), .ZN(n27752) );
  INV_X1 U44765 ( .I(n28988), .ZN(n27749) );
  NAND2_X1 U44766 ( .A1(n29731), .A2(n30027), .ZN(n27750) );
  OAI22_X1 U44767 ( .A1(n27752), .A2(n27751), .B1(n29733), .B2(n27750), .ZN(
        n27753) );
  NAND2_X1 U44768 ( .A1(n28907), .A2(n19451), .ZN(n27758) );
  MUX2_X1 U44770 ( .I0(n27758), .I1(n27757), .S(n28904), .Z(n27772) );
  INV_X1 U44771 ( .I(n30479), .ZN(n27762) );
  AOI21_X1 U44772 ( .A1(n30490), .A2(n27762), .B(n27761), .ZN(n27771) );
  NOR2_X1 U44773 ( .A1(n30475), .A2(n25848), .ZN(n27768) );
  OAI22_X1 U44774 ( .A1(n27766), .A2(n27765), .B1(n27764), .B2(n29814), .ZN(
        n27767) );
  NAND2_X1 U44776 ( .A1(n17414), .A2(n17412), .ZN(n28745) );
  INV_X1 U44777 ( .I(n28745), .ZN(n27780) );
  INV_X1 U44778 ( .I(n29093), .ZN(n27775) );
  NOR2_X1 U44779 ( .A1(n30954), .A2(n64565), .ZN(n27774) );
  INV_X1 U44780 ( .I(n29096), .ZN(n27776) );
  NAND3_X1 U44781 ( .A1(n27781), .A2(n27780), .A3(n28746), .ZN(n27785) );
  NAND3_X1 U44783 ( .A1(n27782), .A2(n740), .A3(n28744), .ZN(n27783) );
  NAND3_X1 U44784 ( .A1(n27785), .A2(n27784), .A3(n27783), .ZN(n27786) );
  XOR2_X1 U44785 ( .A1(n52734), .A2(n56322), .Z(n27787) );
  XOR2_X1 U44786 ( .A1(n15712), .A2(n45404), .Z(n51394) );
  XOR2_X1 U44787 ( .A1(n20623), .A2(n51394), .Z(n31323) );
  INV_X1 U44788 ( .I(n31323), .ZN(n27795) );
  NAND3_X1 U44791 ( .A1(n29246), .A2(n27790), .A3(n1849), .ZN(n27791) );
  CLKBUF_X4 U44792 ( .I(Key[3]), .Z(n53090) );
  XOR2_X1 U44793 ( .A1(n53499), .A2(n53090), .Z(n44378) );
  XOR2_X1 U44795 ( .A1(n44378), .A2(n56784), .Z(n39724) );
  XOR2_X1 U44796 ( .A1(n56702), .A2(n54734), .Z(n42790) );
  CLKBUF_X4 U44797 ( .I(Key[21]), .Z(n53344) );
  XOR2_X1 U44798 ( .A1(n42790), .A2(n53344), .Z(n27793) );
  XOR2_X1 U44799 ( .A1(n27795), .A2(n27794), .Z(n27796) );
  NAND2_X1 U44800 ( .A1(n31129), .A2(n27150), .ZN(n29914) );
  NAND3_X1 U44801 ( .A1(n29914), .A2(n29566), .A3(n29442), .ZN(n27804) );
  INV_X1 U44802 ( .I(n28957), .ZN(n27798) );
  NAND2_X1 U44803 ( .A1(n27800), .A2(n9904), .ZN(n27801) );
  NAND3_X1 U44804 ( .A1(n27801), .A2(n60886), .A3(n61426), .ZN(n27803) );
  NAND3_X1 U44805 ( .A1(n9904), .A2(n29564), .A3(n29566), .ZN(n27802) );
  OAI21_X1 U44806 ( .A1(n20743), .A2(n27812), .B(n28624), .ZN(n27805) );
  NOR2_X1 U44807 ( .A1(n27805), .A2(n29709), .ZN(n27806) );
  AOI22_X1 U44808 ( .A1(n28466), .A2(n4848), .B1(n27807), .B2(n27806), .ZN(
        n27820) );
  NOR2_X1 U44811 ( .A1(n27813), .A2(n27812), .ZN(n27816) );
  NOR2_X1 U44812 ( .A1(n27814), .A2(n7112), .ZN(n27815) );
  OAI21_X1 U44813 ( .A1(n27816), .A2(n29713), .B(n27815), .ZN(n27817) );
  AOI21_X1 U44814 ( .A1(n28619), .A2(n28623), .B(n23540), .ZN(n27825) );
  NOR2_X1 U44815 ( .A1(n27830), .A2(n27841), .ZN(n27831) );
  NOR3_X1 U44818 ( .A1(n10131), .A2(n28496), .A3(n28492), .ZN(n27840) );
  AOI22_X1 U44819 ( .A1(n27840), .A2(n27839), .B1(n27838), .B2(n28492), .ZN(
        n27842) );
  NOR2_X1 U44821 ( .A1(n28616), .A2(n28452), .ZN(n27855) );
  AOI21_X1 U44822 ( .A1(n28460), .A2(n63330), .B(n27855), .ZN(n27858) );
  AOI21_X1 U44823 ( .A1(n27861), .A2(n27860), .B(n20872), .ZN(n27866) );
  NOR2_X1 U44824 ( .A1(n63330), .A2(n10544), .ZN(n27862) );
  OAI21_X1 U44825 ( .A1(n27863), .A2(n27862), .B(n28610), .ZN(n27864) );
  NOR2_X1 U44826 ( .A1(n28532), .A2(n27868), .ZN(n27870) );
  NAND3_X1 U44828 ( .A1(n27877), .A2(n27871), .A3(n3211), .ZN(n27872) );
  NAND2_X1 U44829 ( .A1(n27873), .A2(n27872), .ZN(n27874) );
  NOR2_X1 U44830 ( .A1(n26003), .A2(n27874), .ZN(n27885) );
  OAI21_X1 U44831 ( .A1(n22498), .A2(n27876), .B(n27875), .ZN(n27878) );
  OAI21_X1 U44836 ( .A1(n31177), .A2(n17590), .B(n29901), .ZN(n27898) );
  NAND2_X1 U44837 ( .A1(n27887), .A2(n28188), .ZN(n27889) );
  INV_X1 U44838 ( .I(n22214), .ZN(n27891) );
  NAND2_X1 U44839 ( .A1(n29896), .A2(n24556), .ZN(n27900) );
  NOR4_X1 U44840 ( .A1(n25707), .A2(n29905), .A3(n24777), .A4(n27902), .ZN(
        n27903) );
  NAND2_X1 U44844 ( .A1(n23111), .A2(n30086), .ZN(n27911) );
  NAND3_X1 U44845 ( .A1(n27911), .A2(n64589), .A3(n29797), .ZN(n27912) );
  AOI21_X1 U44847 ( .A1(n27914), .A2(n30085), .B(n29794), .ZN(n27918) );
  AOI21_X1 U44848 ( .A1(n25241), .A2(n58630), .B(n30085), .ZN(n27916) );
  NOR4_X1 U44849 ( .A1(n27922), .A2(n27924), .A3(n27921), .A4(n64057), .ZN(
        n27926) );
  NAND2_X1 U44851 ( .A1(n28267), .A2(n28257), .ZN(n27935) );
  NAND2_X1 U44852 ( .A1(n18375), .A2(n27939), .ZN(n27940) );
  NAND2_X1 U44855 ( .A1(n27945), .A2(n27944), .ZN(n27946) );
  NAND2_X1 U44857 ( .A1(n2513), .A2(n23716), .ZN(n28001) );
  NOR2_X1 U44859 ( .A1(n5627), .A2(n14102), .ZN(n27954) );
  NOR2_X1 U44860 ( .A1(n28222), .A2(n5627), .ZN(n27957) );
  NOR2_X1 U44861 ( .A1(n28225), .A2(n29111), .ZN(n27956) );
  NAND2_X1 U44862 ( .A1(n28018), .A2(n22043), .ZN(n27961) );
  NAND2_X1 U44863 ( .A1(n28278), .A2(n27959), .ZN(n27960) );
  NAND4_X1 U44864 ( .A1(n27961), .A2(n61064), .A3(n27962), .A4(n27960), .ZN(
        n27965) );
  OAI21_X1 U44866 ( .A1(n27980), .A2(n1444), .B(n65198), .ZN(n27982) );
  NAND2_X1 U44867 ( .A1(n28711), .A2(n30334), .ZN(n29950) );
  NAND2_X1 U44869 ( .A1(n23901), .A2(n60202), .ZN(n27989) );
  NAND2_X1 U44870 ( .A1(n30643), .A2(n30408), .ZN(n27995) );
  NOR2_X1 U44871 ( .A1(n30331), .A2(n30639), .ZN(n27993) );
  NAND2_X1 U44874 ( .A1(n28002), .A2(n23665), .ZN(n27997) );
  NOR2_X1 U44875 ( .A1(n435), .A2(n23716), .ZN(n28000) );
  NOR2_X1 U44876 ( .A1(n28279), .A2(n23876), .ZN(n28014) );
  OAI21_X1 U44877 ( .A1(n28014), .A2(n61021), .B(n28021), .ZN(n28016) );
  INV_X1 U44879 ( .I(n28278), .ZN(n28022) );
  NAND2_X1 U44880 ( .A1(n28022), .A2(n28021), .ZN(n28023) );
  AOI22_X1 U44881 ( .A1(n28043), .A2(n61484), .B1(n28333), .B2(n28042), .ZN(
        n28058) );
  NOR2_X1 U44882 ( .A1(n28045), .A2(n7438), .ZN(n28046) );
  NOR2_X1 U44883 ( .A1(n28049), .A2(n22408), .ZN(n28050) );
  OAI21_X1 U44884 ( .A1(n7438), .A2(n28053), .B(n28052), .ZN(n28055) );
  NAND4_X2 U44885 ( .A1(n28058), .A2(n28057), .A3(n28056), .A4(n28055), .ZN(
        n28060) );
  NAND2_X1 U44886 ( .A1(n23397), .A2(n30319), .ZN(n28061) );
  NOR2_X1 U44887 ( .A1(n28061), .A2(n61052), .ZN(n28077) );
  INV_X1 U44888 ( .I(n28062), .ZN(n28063) );
  NAND2_X1 U44889 ( .A1(n60768), .A2(n28066), .ZN(n28068) );
  NAND3_X1 U44891 ( .A1(n30322), .A2(n29993), .A3(n14230), .ZN(n28078) );
  INV_X1 U44892 ( .I(n29994), .ZN(n29826) );
  NAND3_X1 U44893 ( .A1(n64154), .A2(n22556), .A3(n30319), .ZN(n28082) );
  OAI22_X1 U44894 ( .A1(n30322), .A2(n28082), .B1(n28083), .B2(n30319), .ZN(
        n28085) );
  OAI21_X1 U44895 ( .A1(n28085), .A2(n28084), .B(n61052), .ZN(n28088) );
  INV_X1 U44897 ( .I(n28699), .ZN(n28086) );
  NOR2_X1 U44898 ( .A1(n29272), .A2(n28086), .ZN(n28087) );
  INV_X1 U44899 ( .I(n28103), .ZN(n28111) );
  INV_X1 U44900 ( .I(n28104), .ZN(n28110) );
  INV_X1 U44901 ( .I(n28105), .ZN(n28109) );
  AOI21_X1 U44902 ( .A1(n28107), .A2(n23071), .B(n1440), .ZN(n28108) );
  NOR4_X1 U44903 ( .A1(n28111), .A2(n28110), .A3(n28109), .A4(n28108), .ZN(
        n28114) );
  INV_X1 U44904 ( .I(n28112), .ZN(n28113) );
  NAND3_X1 U44905 ( .A1(n28115), .A2(n22230), .A3(n28730), .ZN(n28116) );
  INV_X1 U44907 ( .I(n28120), .ZN(n28130) );
  INV_X1 U44908 ( .I(n28825), .ZN(n29280) );
  AOI21_X1 U44909 ( .A1(n29287), .A2(n28130), .B(n29280), .ZN(n28123) );
  NAND2_X1 U44910 ( .A1(n28124), .A2(n28121), .ZN(n28122) );
  INV_X1 U44911 ( .I(n28125), .ZN(n28821) );
  NOR2_X1 U44913 ( .A1(n28128), .A2(n28127), .ZN(n29631) );
  NAND2_X1 U44914 ( .A1(n29284), .A2(n29283), .ZN(n28129) );
  NOR3_X2 U44916 ( .A1(n28143), .A2(n28142), .A3(n28141), .ZN(n30580) );
  INV_X1 U44917 ( .I(n29645), .ZN(n28144) );
  NAND3_X1 U44918 ( .A1(n19566), .A2(n28144), .A3(n20907), .ZN(n28145) );
  NOR2_X1 U44919 ( .A1(n28148), .A2(n1358), .ZN(n28149) );
  AOI21_X1 U44921 ( .A1(n28860), .A2(n19967), .B(n29321), .ZN(n28155) );
  NAND3_X1 U44922 ( .A1(n28157), .A2(n28156), .A3(n28155), .ZN(n28160) );
  NAND3_X1 U44923 ( .A1(n29324), .A2(n23596), .A3(n28854), .ZN(n28159) );
  INV_X1 U44924 ( .I(n28164), .ZN(n28165) );
  OAI21_X1 U44925 ( .A1(n29323), .A2(n28166), .B(n28165), .ZN(n28167) );
  NAND2_X1 U44926 ( .A1(n28174), .A2(n61307), .ZN(n28169) );
  NOR2_X1 U44928 ( .A1(n12739), .A2(n29608), .ZN(n28171) );
  NAND2_X1 U44929 ( .A1(n28173), .A2(n28172), .ZN(n28180) );
  NOR2_X1 U44930 ( .A1(n28174), .A2(n4715), .ZN(n28178) );
  OAI22_X1 U44931 ( .A1(n23816), .A2(n28176), .B1(n28175), .B2(n28665), .ZN(
        n28177) );
  NAND2_X1 U44933 ( .A1(n28191), .A2(n19279), .ZN(n28194) );
  AOI21_X1 U44935 ( .A1(n28194), .A2(n28872), .B(n28193), .ZN(n28202) );
  INV_X1 U44936 ( .I(n28195), .ZN(n28197) );
  NAND2_X1 U44937 ( .A1(n58601), .A2(n29661), .ZN(n28196) );
  NOR2_X1 U44938 ( .A1(n29659), .A2(n29663), .ZN(n28199) );
  NOR3_X1 U44941 ( .A1(n28212), .A2(n21956), .A3(n24080), .ZN(n28213) );
  NAND3_X1 U44942 ( .A1(n28222), .A2(n10404), .A3(n14102), .ZN(n28227) );
  OAI21_X1 U44945 ( .A1(n28243), .A2(n28242), .B(n28241), .ZN(n28247) );
  NAND2_X1 U44946 ( .A1(n29170), .A2(n28254), .ZN(n28255) );
  INV_X1 U44947 ( .I(n28264), .ZN(n28265) );
  NAND2_X1 U44948 ( .A1(n23876), .A2(n61021), .ZN(n28274) );
  OAI21_X1 U44949 ( .A1(n28277), .A2(n28276), .B(n61049), .ZN(n28286) );
  NAND3_X1 U44950 ( .A1(n28279), .A2(n28278), .A3(n60885), .ZN(n28283) );
  AOI21_X1 U44951 ( .A1(n3097), .A2(n29430), .B(n28288), .ZN(n28290) );
  NAND2_X1 U44952 ( .A1(n22706), .A2(n28299), .ZN(n28304) );
  NOR2_X1 U44953 ( .A1(n28305), .A2(n23840), .ZN(n28307) );
  NAND2_X1 U44954 ( .A1(n28313), .A2(n28312), .ZN(n28315) );
  OAI22_X1 U44955 ( .A1(n28318), .A2(n21065), .B1(n28329), .B2(n28316), .ZN(
        n28319) );
  NAND2_X1 U44956 ( .A1(n28319), .A2(n23997), .ZN(n28326) );
  OAI21_X1 U44957 ( .A1(n28322), .A2(n28321), .B(n28320), .ZN(n28323) );
  INV_X1 U44958 ( .I(n28327), .ZN(n28331) );
  NAND4_X1 U44959 ( .A1(n28331), .A2(n28330), .A3(n28329), .A4(n23997), .ZN(
        n28338) );
  INV_X1 U44961 ( .I(n28335), .ZN(n28336) );
  NAND3_X1 U44962 ( .A1(n28342), .A2(n28341), .A3(n16021), .ZN(n28343) );
  AOI21_X1 U44964 ( .A1(n23362), .A2(n24734), .B(n28348), .ZN(n28355) );
  OAI21_X1 U44965 ( .A1(n28355), .A2(n28354), .B(n28353), .ZN(n28356) );
  NOR2_X1 U44966 ( .A1(n28359), .A2(n22604), .ZN(n28364) );
  NOR2_X1 U44967 ( .A1(n28364), .A2(n28363), .ZN(n28372) );
  NOR2_X1 U44968 ( .A1(n28366), .A2(n62083), .ZN(n28368) );
  OAI21_X1 U44969 ( .A1(n28368), .A2(n1279), .B(n28367), .ZN(n28369) );
  INV_X1 U44970 ( .I(n28374), .ZN(n28377) );
  INV_X1 U44973 ( .I(n29571), .ZN(n30298) );
  NOR2_X1 U44974 ( .A1(n30298), .A2(n28921), .ZN(n28422) );
  INV_X1 U44975 ( .I(n22397), .ZN(n28394) );
  NAND3_X1 U44976 ( .A1(n28397), .A2(n28396), .A3(n28409), .ZN(n28398) );
  INV_X1 U44977 ( .I(n28405), .ZN(n28407) );
  NAND2_X1 U44978 ( .A1(n28409), .A2(n3117), .ZN(n28411) );
  OAI22_X1 U44979 ( .A1(n28417), .A2(n28416), .B1(n28415), .B2(n1891), .ZN(
        n28421) );
  NOR3_X1 U44980 ( .A1(n29268), .A2(n63890), .A3(n1317), .ZN(n28424) );
  NAND2_X1 U44981 ( .A1(n28425), .A2(n28424), .ZN(n28433) );
  NAND2_X1 U44982 ( .A1(n30300), .A2(n9865), .ZN(n28927) );
  INV_X1 U44983 ( .I(n28927), .ZN(n28428) );
  INV_X1 U44985 ( .I(n30293), .ZN(n28429) );
  NAND4_X1 U44986 ( .A1(n28430), .A2(n63890), .A3(n28429), .A4(n64867), .ZN(
        n28432) );
  NOR2_X1 U44990 ( .A1(n28611), .A2(n28445), .ZN(n28450) );
  AOI21_X1 U44991 ( .A1(n22312), .A2(n28447), .B(n23487), .ZN(n28449) );
  OAI21_X1 U44992 ( .A1(n28450), .A2(n28449), .B(n63330), .ZN(n28458) );
  OAI21_X1 U44995 ( .A1(n28462), .A2(n28461), .B(n28617), .ZN(n28463) );
  NOR2_X1 U44997 ( .A1(n28472), .A2(n7112), .ZN(n28473) );
  INV_X1 U44998 ( .I(n28475), .ZN(n28479) );
  NAND2_X1 U44999 ( .A1(n62469), .A2(n28483), .ZN(n28484) );
  OAI21_X1 U45000 ( .A1(n28489), .A2(n62469), .B(n28487), .ZN(n28503) );
  NAND2_X1 U45001 ( .A1(n28491), .A2(n28490), .ZN(n28501) );
  NAND3_X1 U45002 ( .A1(n28494), .A2(n60541), .A3(n28492), .ZN(n28500) );
  NAND3_X1 U45003 ( .A1(n28497), .A2(n28496), .A3(n10125), .ZN(n28498) );
  NOR2_X2 U45004 ( .A1(n28503), .A2(n28502), .ZN(n30338) );
  NOR2_X2 U45005 ( .A1(n28524), .A2(n28523), .ZN(n30609) );
  NOR2_X1 U45006 ( .A1(n28529), .A2(n28528), .ZN(n28531) );
  NAND2_X1 U45007 ( .A1(n28534), .A2(n28533), .ZN(n28535) );
  NAND2_X1 U45008 ( .A1(n28536), .A2(n28535), .ZN(n28538) );
  NAND3_X1 U45009 ( .A1(n28538), .A2(n28543), .A3(n63533), .ZN(n28545) );
  NOR2_X1 U45010 ( .A1(n28540), .A2(n28539), .ZN(n28544) );
  OAI21_X1 U45011 ( .A1(n30617), .A2(n29078), .B(n30618), .ZN(n28562) );
  INV_X1 U45013 ( .I(n29594), .ZN(n30606) );
  NAND2_X1 U45014 ( .A1(n29187), .A2(n28557), .ZN(n28558) );
  NOR2_X1 U45016 ( .A1(n22504), .A2(n30616), .ZN(n29593) );
  NAND2_X1 U45019 ( .A1(n40), .A2(n30616), .ZN(n28564) );
  OAI21_X1 U45020 ( .A1(n31089), .A2(n60064), .B(n28570), .ZN(n28579) );
  NAND2_X1 U45022 ( .A1(n31080), .A2(n61629), .ZN(n28572) );
  NOR2_X1 U45024 ( .A1(n28576), .A2(n28575), .ZN(n28577) );
  NAND2_X1 U45025 ( .A1(n24504), .A2(n25384), .ZN(n28580) );
  OAI21_X1 U45026 ( .A1(n24504), .A2(n29472), .B(n28580), .ZN(n28581) );
  XOR2_X1 U45027 ( .A1(n56495), .A2(n22773), .Z(n39469) );
  XOR2_X1 U45028 ( .A1(n54556), .A2(n23886), .Z(n37481) );
  XOR2_X1 U45029 ( .A1(n37481), .A2(n39469), .Z(n51005) );
  XOR2_X1 U45030 ( .A1(n51005), .A2(n44759), .Z(n44112) );
  NAND2_X1 U45031 ( .A1(n28588), .A2(n28587), .ZN(n28590) );
  NAND2_X1 U45032 ( .A1(n28846), .A2(n59935), .ZN(n28591) );
  AOI22_X1 U45033 ( .A1(n61004), .A2(n29635), .B1(n434), .B2(n28843), .ZN(
        n28603) );
  NAND2_X1 U45034 ( .A1(n4812), .A2(n23386), .ZN(n28602) );
  NAND2_X1 U45035 ( .A1(n28607), .A2(n28606), .ZN(n28608) );
  NAND2_X1 U45038 ( .A1(n28623), .A2(n28630), .ZN(n28628) );
  NOR2_X1 U45039 ( .A1(n29713), .A2(n28624), .ZN(n28627) );
  OAI22_X1 U45041 ( .A1(n28635), .A2(n28634), .B1(n22648), .B2(n1970), .ZN(
        n28636) );
  OAI22_X1 U45042 ( .A1(n491), .A2(n25341), .B1(n28640), .B2(n10598), .ZN(
        n28642) );
  OAI21_X1 U45044 ( .A1(n28645), .A2(n28644), .B(n28643), .ZN(n28655) );
  NAND3_X1 U45045 ( .A1(n60547), .A2(n28651), .A3(n60603), .ZN(n28650) );
  NOR2_X1 U45046 ( .A1(n60547), .A2(n10598), .ZN(n28647) );
  AOI21_X1 U45047 ( .A1(n28648), .A2(n28647), .B(n28646), .ZN(n28649) );
  NOR2_X1 U45048 ( .A1(n29648), .A2(n29663), .ZN(n28656) );
  OAI21_X1 U45049 ( .A1(n29652), .A2(n58601), .B(n28656), .ZN(n28661) );
  NAND2_X1 U45050 ( .A1(n28873), .A2(n29663), .ZN(n28657) );
  AOI21_X1 U45051 ( .A1(n28658), .A2(n58955), .B(n57781), .ZN(n28660) );
  NOR3_X1 U45052 ( .A1(n29652), .A2(n8296), .A3(n58955), .ZN(n28659) );
  NAND2_X1 U45053 ( .A1(n28665), .A2(n29609), .ZN(n28666) );
  OAI21_X1 U45054 ( .A1(n28670), .A2(n59099), .B(n28669), .ZN(n28671) );
  INV_X1 U45055 ( .I(n28677), .ZN(n28678) );
  NAND2_X1 U45058 ( .A1(n14217), .A2(n1432), .ZN(n28682) );
  INV_X1 U45059 ( .I(n29736), .ZN(n28685) );
  INV_X1 U45060 ( .I(n28689), .ZN(n28693) );
  NAND2_X1 U45061 ( .A1(n364), .A2(n30197), .ZN(n28691) );
  AOI21_X1 U45062 ( .A1(n24712), .A2(n62585), .B(n28691), .ZN(n28692) );
  NOR2_X1 U45063 ( .A1(n28693), .A2(n28692), .ZN(n28694) );
  NAND2_X1 U45064 ( .A1(n16961), .A2(n14230), .ZN(n28695) );
  AOI21_X1 U45065 ( .A1(n29820), .A2(n29824), .B(n30321), .ZN(n28702) );
  MUX2_X1 U45066 ( .I0(n29824), .I1(n29820), .S(n30322), .Z(n28701) );
  NOR3_X1 U45071 ( .A1(n30771), .A2(n30786), .A3(n30767), .ZN(n28725) );
  NOR2_X1 U45072 ( .A1(n30786), .A2(n24206), .ZN(n28723) );
  OAI21_X1 U45076 ( .A1(n60030), .A2(n29458), .B(n29840), .ZN(n28728) );
  INV_X1 U45077 ( .I(n28730), .ZN(n29843) );
  NAND2_X1 U45080 ( .A1(n28732), .A2(n22230), .ZN(n28740) );
  INV_X1 U45081 ( .I(n28733), .ZN(n28734) );
  NAND2_X1 U45082 ( .A1(n28996), .A2(n28734), .ZN(n28739) );
  INV_X1 U45083 ( .I(n28995), .ZN(n28737) );
  NAND2_X1 U45085 ( .A1(n29835), .A2(n10820), .ZN(n28751) );
  XOR2_X1 U45086 ( .A1(n55655), .A2(n56202), .Z(n46180) );
  XOR2_X1 U45088 ( .A1(n23968), .A2(n56976), .Z(n38450) );
  XOR2_X1 U45089 ( .A1(n1190), .A2(n38450), .Z(n33134) );
  XOR2_X1 U45090 ( .A1(n23999), .A2(n54587), .Z(n50486) );
  XOR2_X1 U45092 ( .A1(n33134), .A2(n50793), .Z(n38502) );
  XOR2_X1 U45093 ( .A1(n53124), .A2(n56819), .Z(n32274) );
  XOR2_X1 U45094 ( .A1(n38502), .A2(n32274), .Z(n51133) );
  XOR2_X1 U45095 ( .A1(n51133), .A2(n52232), .Z(n37378) );
  XOR2_X1 U45097 ( .A1(n24098), .A2(n56901), .Z(n28757) );
  BUF_X2 U45098 ( .I(n28757), .Z(n50067) );
  XOR2_X1 U45099 ( .A1(n50067), .A2(n56745), .Z(n34467) );
  XOR2_X1 U45100 ( .A1(n34467), .A2(n23455), .Z(n38506) );
  XOR2_X1 U45101 ( .A1(n56124), .A2(n54208), .Z(n30568) );
  XOR2_X1 U45102 ( .A1(n38506), .A2(n30568), .Z(n45869) );
  CLKBUF_X4 U45103 ( .I(Key[41]), .Z(n50475) );
  XOR2_X1 U45104 ( .A1(n53308), .A2(n50475), .Z(n32741) );
  XOR2_X1 U45105 ( .A1(n32741), .A2(n53530), .Z(n37520) );
  XOR2_X1 U45106 ( .A1(n37520), .A2(n54289), .Z(n43485) );
  XOR2_X1 U45107 ( .A1(n45869), .A2(n43485), .Z(n28758) );
  XOR2_X1 U45108 ( .A1(n37378), .A2(n28758), .Z(n28770) );
  NAND2_X1 U45109 ( .A1(n28937), .A2(n58710), .ZN(n28761) );
  NOR2_X1 U45110 ( .A1(n29779), .A2(n13336), .ZN(n29780) );
  MUX2_X1 U45111 ( .I0(n28761), .I1(n28760), .S(n14063), .Z(n28769) );
  NAND2_X1 U45112 ( .A1(n28762), .A2(n58486), .ZN(n28764) );
  NAND2_X1 U45113 ( .A1(n63272), .A2(n29251), .ZN(n28763) );
  OAI22_X1 U45114 ( .A1(n28942), .A2(n28764), .B1(n28763), .B2(n29784), .ZN(
        n28768) );
  XOR2_X1 U45116 ( .A1(n28770), .A2(n31365), .Z(n28784) );
  NOR2_X1 U45117 ( .A1(n61734), .A2(n23772), .ZN(n28771) );
  NAND2_X1 U45118 ( .A1(n10431), .A2(n22496), .ZN(n28778) );
  NAND3_X1 U45120 ( .A1(n29798), .A2(n60262), .A3(n29794), .ZN(n28789) );
  NAND2_X1 U45121 ( .A1(n22877), .A2(n1351), .ZN(n28793) );
  OAI22_X1 U45122 ( .A1(n30121), .A2(n28794), .B1(n29766), .B2(n30525), .ZN(
        n28795) );
  OAI21_X1 U45123 ( .A1(n28798), .A2(n23824), .B(n28797), .ZN(n28799) );
  NOR2_X1 U45124 ( .A1(n29372), .A2(n23824), .ZN(n28816) );
  AOI21_X1 U45125 ( .A1(n28812), .A2(n20678), .B(n28810), .ZN(n28818) );
  NAND2_X1 U45127 ( .A1(n28821), .A2(n29285), .ZN(n28824) );
  OAI22_X1 U45129 ( .A1(n29626), .A2(n28824), .B1(n29625), .B2(n28823), .ZN(
        n28830) );
  NAND2_X1 U45130 ( .A1(n28825), .A2(n19290), .ZN(n28826) );
  OAI22_X1 U45131 ( .A1(n28828), .A2(n28827), .B1(n28826), .B2(n29281), .ZN(
        n28829) );
  NAND2_X1 U45132 ( .A1(n23732), .A2(n28831), .ZN(n28832) );
  NAND2_X1 U45133 ( .A1(n29286), .A2(n28832), .ZN(n28834) );
  NAND2_X1 U45135 ( .A1(n28836), .A2(n19290), .ZN(n28840) );
  NOR2_X1 U45136 ( .A1(n28838), .A2(n28837), .ZN(n28839) );
  NAND2_X1 U45137 ( .A1(n28850), .A2(n58108), .ZN(n28867) );
  NAND2_X1 U45138 ( .A1(n23797), .A2(n29310), .ZN(n28851) );
  OAI21_X1 U45139 ( .A1(n28852), .A2(n28851), .B(n64451), .ZN(n28859) );
  INV_X1 U45140 ( .I(n28853), .ZN(n28856) );
  OAI22_X1 U45141 ( .A1(n28856), .A2(n28855), .B1(n29316), .B2(n28854), .ZN(
        n28857) );
  AOI21_X1 U45142 ( .A1(n28859), .A2(n19967), .B(n28857), .ZN(n28866) );
  NOR2_X1 U45145 ( .A1(n28862), .A2(n29321), .ZN(n28863) );
  NOR2_X1 U45146 ( .A1(n29379), .A2(n28868), .ZN(n28869) );
  NAND2_X1 U45147 ( .A1(n29659), .A2(n28872), .ZN(n28874) );
  NAND3_X1 U45148 ( .A1(n28878), .A2(n28884), .A3(n58977), .ZN(n28882) );
  OAI21_X1 U45149 ( .A1(n28879), .A2(n29356), .B(n29344), .ZN(n28880) );
  NAND3_X1 U45150 ( .A1(n28882), .A2(n28881), .A3(n28880), .ZN(n28892) );
  AOI21_X1 U45151 ( .A1(n28883), .A2(n29334), .B(n29340), .ZN(n28891) );
  NAND4_X1 U45152 ( .A1(n28884), .A2(n7495), .A3(n62341), .A4(n29355), .ZN(
        n28889) );
  NOR2_X1 U45153 ( .A1(n28886), .A2(n19452), .ZN(n28887) );
  NOR3_X1 U45154 ( .A1(n30308), .A2(n30752), .A3(n31214), .ZN(n28896) );
  NAND2_X1 U45155 ( .A1(n7426), .A2(n30752), .ZN(n28893) );
  AOI21_X1 U45156 ( .A1(n28893), .A2(n30760), .B(n30013), .ZN(n28895) );
  NOR3_X1 U45158 ( .A1(n28896), .A2(n28895), .A3(n30005), .ZN(n28897) );
  INV_X1 U45159 ( .I(n30617), .ZN(n28909) );
  NAND4_X1 U45160 ( .A1(n28909), .A2(n30342), .A3(n29076), .A4(n59268), .ZN(
        n28913) );
  NAND2_X1 U45161 ( .A1(n16750), .A2(n30348), .ZN(n29595) );
  INV_X1 U45162 ( .I(n29595), .ZN(n28911) );
  OAI21_X1 U45163 ( .A1(n28911), .A2(n59268), .B(n30351), .ZN(n28912) );
  INV_X1 U45164 ( .I(n28918), .ZN(n28916) );
  INV_X1 U45165 ( .I(n30342), .ZN(n28915) );
  NAND3_X1 U45166 ( .A1(n28918), .A2(n22555), .A3(n29078), .ZN(n28919) );
  MUX2_X1 U45167 ( .I0(n30301), .I1(n28922), .S(n28921), .Z(n28929) );
  OAI21_X1 U45169 ( .A1(n30296), .A2(n23734), .B(n28923), .ZN(n28924) );
  AOI21_X1 U45170 ( .A1(n28927), .A2(n30302), .B(n28926), .ZN(n28928) );
  XOR2_X1 U45171 ( .A1(n7557), .A2(n28930), .Z(n28931) );
  NOR2_X1 U45172 ( .A1(n1863), .A2(n19461), .ZN(n28935) );
  OAI21_X1 U45173 ( .A1(n28938), .A2(n24097), .B(n7943), .ZN(n28939) );
  NAND3_X1 U45174 ( .A1(n29246), .A2(n29251), .A3(n28943), .ZN(n28944) );
  NAND2_X1 U45175 ( .A1(n29560), .A2(n31127), .ZN(n28955) );
  OAI22_X1 U45176 ( .A1(n59613), .A2(n28953), .B1(n28952), .B2(n28951), .ZN(
        n28954) );
  NAND2_X1 U45177 ( .A1(n29440), .A2(n24000), .ZN(n28961) );
  NAND2_X1 U45178 ( .A1(n31129), .A2(n59541), .ZN(n28960) );
  AOI21_X1 U45179 ( .A1(n28961), .A2(n28960), .B(n29560), .ZN(n28962) );
  NAND2_X1 U45180 ( .A1(n29896), .A2(n1353), .ZN(n28964) );
  NAND2_X1 U45182 ( .A1(n31187), .A2(n24556), .ZN(n28965) );
  NOR3_X1 U45183 ( .A1(n24777), .A2(n29896), .A3(n57937), .ZN(n28971) );
  OAI21_X1 U45185 ( .A1(n31182), .A2(n28971), .B(n28970), .ZN(n28975) );
  NAND2_X1 U45186 ( .A1(n30296), .A2(n13731), .ZN(n28977) );
  AOI21_X1 U45187 ( .A1(n1317), .A2(n13731), .B(n1562), .ZN(n28980) );
  NAND2_X1 U45188 ( .A1(n846), .A2(n1317), .ZN(n28979) );
  XOR2_X1 U45190 ( .A1(n54896), .A2(n54231), .Z(n51999) );
  XOR2_X1 U45191 ( .A1(n21006), .A2(n51999), .Z(n32611) );
  AOI21_X1 U45193 ( .A1(n25978), .A2(n28988), .B(n30027), .ZN(n28993) );
  NAND3_X1 U45194 ( .A1(n28996), .A2(n29460), .A3(n23224), .ZN(n28999) );
  AOI21_X1 U45195 ( .A1(n23224), .A2(n61421), .B(n29452), .ZN(n28997) );
  NAND2_X1 U45196 ( .A1(n29000), .A2(n60028), .ZN(n29001) );
  INV_X1 U45197 ( .I(n30589), .ZN(n29009) );
  NAND2_X1 U45199 ( .A1(n29016), .A2(n25241), .ZN(n29017) );
  NOR2_X1 U45202 ( .A1(n29027), .A2(n30174), .ZN(n29032) );
  INV_X1 U45203 ( .I(n58999), .ZN(n30167) );
  NAND2_X1 U45204 ( .A1(n31059), .A2(n31055), .ZN(n30163) );
  AOI21_X1 U45205 ( .A1(n30165), .A2(n30163), .B(n29029), .ZN(n29031) );
  NAND2_X2 U45206 ( .A1(n30285), .A2(n22139), .ZN(n30724) );
  NOR2_X1 U45208 ( .A1(n30725), .A2(n30276), .ZN(n29040) );
  NAND2_X1 U45210 ( .A1(n23317), .A2(n1438), .ZN(n30275) );
  NAND2_X1 U45215 ( .A1(n29063), .A2(n29422), .ZN(n29067) );
  INV_X1 U45216 ( .I(n30451), .ZN(n29064) );
  NOR2_X1 U45217 ( .A1(n29064), .A2(n60170), .ZN(n29066) );
  NAND2_X1 U45218 ( .A1(n29422), .A2(n21095), .ZN(n29065) );
  XOR2_X1 U45220 ( .A1(n29070), .A2(n51019), .Z(n31593) );
  XOR2_X1 U45221 ( .A1(n54716), .A2(n55196), .Z(n44262) );
  XOR2_X1 U45222 ( .A1(n31593), .A2(n44262), .Z(n51638) );
  XOR2_X1 U45223 ( .A1(n54386), .A2(n55060), .Z(n38733) );
  XOR2_X1 U45224 ( .A1(n38851), .A2(n38733), .Z(n38153) );
  XOR2_X1 U45226 ( .A1(n56040), .A2(n55546), .Z(n37513) );
  XOR2_X1 U45227 ( .A1(n37513), .A2(n55777), .Z(n38614) );
  BUF_X2 U45228 ( .I(Key[176]), .Z(n56859) );
  XOR2_X1 U45229 ( .A1(n24011), .A2(n56859), .Z(n29071) );
  BUF_X2 U45230 ( .I(n29071), .Z(n50955) );
  INV_X1 U45231 ( .I(n50955), .ZN(n29072) );
  XOR2_X1 U45232 ( .A1(n38614), .A2(n29072), .Z(n32396) );
  INV_X1 U45233 ( .I(n32396), .ZN(n44808) );
  XOR2_X1 U45234 ( .A1(n38153), .A2(n44808), .Z(n52527) );
  XOR2_X1 U45235 ( .A1(n56771), .A2(n54536), .Z(n51021) );
  XOR2_X1 U45236 ( .A1(n51021), .A2(n55126), .Z(n45240) );
  XNOR2_X1 U45237 ( .A1(n55610), .A2(n56915), .ZN(n29073) );
  XOR2_X1 U45238 ( .A1(n45240), .A2(n29073), .Z(n29074) );
  XOR2_X1 U45239 ( .A1(n52527), .A2(n29074), .Z(n29075) );
  NAND2_X1 U45241 ( .A1(n30618), .A2(n30617), .ZN(n29080) );
  NAND3_X1 U45242 ( .A1(n30623), .A2(n65233), .A3(n21029), .ZN(n29087) );
  NOR2_X1 U45243 ( .A1(n29085), .A2(n40), .ZN(n30619) );
  INV_X1 U45244 ( .I(n30619), .ZN(n29086) );
  INV_X1 U45246 ( .I(n29864), .ZN(n29090) );
  NAND2_X1 U45247 ( .A1(n29093), .A2(n29100), .ZN(n29094) );
  NOR2_X1 U45248 ( .A1(n29855), .A2(n29521), .ZN(n29098) );
  NOR2_X1 U45249 ( .A1(n21511), .A2(n23591), .ZN(n29135) );
  NOR2_X1 U45252 ( .A1(n12072), .A2(n23769), .ZN(n29169) );
  NOR2_X1 U45253 ( .A1(n1869), .A2(n24196), .ZN(n29193) );
  INV_X1 U45254 ( .I(n29177), .ZN(n29184) );
  AOI21_X1 U45255 ( .A1(n21068), .A2(n22351), .B(n4847), .ZN(n29181) );
  NOR3_X1 U45256 ( .A1(n29189), .A2(n4847), .A3(n29188), .ZN(n29190) );
  NOR3_X1 U45257 ( .A1(n7376), .A2(n29193), .A3(n29805), .ZN(n29199) );
  NAND2_X1 U45258 ( .A1(n22596), .A2(n24196), .ZN(n29196) );
  OAI22_X1 U45260 ( .A1(n30214), .A2(n29196), .B1(n29195), .B2(n29194), .ZN(
        n29198) );
  NAND2_X1 U45262 ( .A1(n34558), .A2(n34553), .ZN(n29558) );
  NAND2_X1 U45263 ( .A1(n29207), .A2(n19218), .ZN(n29208) );
  NOR2_X1 U45264 ( .A1(n19461), .A2(n22496), .ZN(n29210) );
  OAI21_X1 U45265 ( .A1(n10431), .A2(n57953), .B(n29210), .ZN(n29212) );
  NAND3_X1 U45270 ( .A1(n30273), .A2(n29218), .A3(n30718), .ZN(n29229) );
  INV_X1 U45271 ( .I(n30718), .ZN(n29219) );
  NAND2_X1 U45273 ( .A1(n29219), .A2(n30719), .ZN(n29228) );
  NOR2_X1 U45274 ( .A1(n29220), .A2(n30276), .ZN(n29223) );
  NOR3_X1 U45275 ( .A1(n29223), .A2(n29222), .A3(n29221), .ZN(n29227) );
  INV_X1 U45276 ( .I(n29224), .ZN(n29225) );
  NAND2_X1 U45279 ( .A1(n30815), .A2(n29933), .ZN(n29233) );
  INV_X1 U45280 ( .I(n29239), .ZN(n29240) );
  NOR3_X1 U45281 ( .A1(n25448), .A2(n29240), .A3(n30808), .ZN(n29243) );
  NOR2_X1 U45282 ( .A1(n29245), .A2(n29244), .ZN(n29247) );
  INV_X1 U45283 ( .I(n63355), .ZN(n29249) );
  NAND2_X1 U45284 ( .A1(n7943), .A2(n29779), .ZN(n29786) );
  INV_X1 U45287 ( .I(n29260), .ZN(n29265) );
  NAND2_X1 U45290 ( .A1(n2119), .A2(n64154), .ZN(n29275) );
  INV_X1 U45291 ( .I(n16026), .ZN(n29277) );
  NAND2_X1 U45292 ( .A1(n23237), .A2(n2119), .ZN(n29276) );
  NAND2_X1 U45293 ( .A1(n29631), .A2(n23732), .ZN(n29290) );
  NAND2_X1 U45294 ( .A1(n29292), .A2(n1360), .ZN(n29294) );
  NOR2_X1 U45295 ( .A1(n25532), .A2(n59552), .ZN(n29293) );
  NAND2_X1 U45297 ( .A1(n29313), .A2(n20665), .ZN(n29314) );
  NAND2_X1 U45298 ( .A1(n29323), .A2(n29322), .ZN(n29330) );
  NAND3_X1 U45299 ( .A1(n57424), .A2(n29325), .A3(n29324), .ZN(n29329) );
  INV_X1 U45300 ( .I(n29327), .ZN(n29328) );
  NAND2_X1 U45301 ( .A1(n29332), .A2(n31254), .ZN(n29395) );
  NAND3_X1 U45307 ( .A1(n29344), .A2(n23954), .A3(n62341), .ZN(n29347) );
  MUX2_X1 U45308 ( .I0(n29351), .I1(n29350), .S(n29355), .Z(n29354) );
  AOI21_X1 U45309 ( .A1(n29354), .A2(n62341), .B(n29352), .ZN(n29364) );
  NAND3_X1 U45310 ( .A1(n29357), .A2(n29356), .A3(n29355), .ZN(n29362) );
  NAND2_X1 U45312 ( .A1(n29367), .A2(n29372), .ZN(n29368) );
  AOI21_X1 U45313 ( .A1(n29372), .A2(n17460), .B(n22158), .ZN(n29374) );
  NAND2_X1 U45314 ( .A1(n1356), .A2(n8296), .ZN(n29376) );
  OAI22_X1 U45316 ( .A1(n29675), .A2(n29378), .B1(n29667), .B2(n10805), .ZN(
        n29389) );
  NAND2_X1 U45317 ( .A1(n29380), .A2(n29383), .ZN(n29387) );
  INV_X1 U45318 ( .I(n30885), .ZN(n29399) );
  INV_X1 U45319 ( .I(n30889), .ZN(n29398) );
  NAND3_X1 U45320 ( .A1(n29399), .A2(n12893), .A3(n29398), .ZN(n29401) );
  XOR2_X1 U45321 ( .A1(n620), .A2(n54219), .Z(n45064) );
  XOR2_X1 U45322 ( .A1(n53945), .A2(n51569), .Z(n29403) );
  XOR2_X1 U45323 ( .A1(n45064), .A2(n29403), .Z(n39235) );
  XOR2_X1 U45324 ( .A1(n55862), .A2(n23989), .Z(n38639) );
  INV_X1 U45325 ( .I(n38639), .ZN(n29404) );
  XOR2_X1 U45326 ( .A1(n39235), .A2(n29404), .Z(n44598) );
  XOR2_X1 U45327 ( .A1(n56683), .A2(n57113), .Z(n29405) );
  BUF_X2 U45328 ( .I(n29405), .Z(n52080) );
  XOR2_X1 U45329 ( .A1(n52080), .A2(n53064), .Z(n29406) );
  XOR2_X1 U45330 ( .A1(n44598), .A2(n29406), .Z(n29408) );
  XOR2_X1 U45331 ( .A1(n55534), .A2(n56030), .Z(n52513) );
  XOR2_X1 U45332 ( .A1(n54143), .A2(n29407), .Z(n48764) );
  XOR2_X1 U45333 ( .A1(n52513), .A2(n48764), .Z(n37691) );
  XOR2_X1 U45334 ( .A1(n24067), .A2(n56309), .Z(n32251) );
  XOR2_X1 U45335 ( .A1(n64355), .A2(n32251), .Z(n45854) );
  XOR2_X1 U45336 ( .A1(n29408), .A2(n45854), .Z(n29409) );
  XOR2_X1 U45337 ( .A1(n23683), .A2(n29409), .Z(n29410) );
  OAI22_X1 U45338 ( .A1(n29413), .A2(n29412), .B1(n30439), .B2(n30541), .ZN(
        n29414) );
  NOR2_X1 U45339 ( .A1(n29981), .A2(n58409), .ZN(n29417) );
  AOI21_X1 U45341 ( .A1(n30451), .A2(n58448), .B(n29423), .ZN(n29424) );
  OAI21_X1 U45342 ( .A1(n29434), .A2(n29433), .B(n60575), .ZN(n29446) );
  AOI21_X1 U45343 ( .A1(n29566), .A2(n29435), .B(n3267), .ZN(n29438) );
  NOR2_X1 U45344 ( .A1(n59613), .A2(n61426), .ZN(n29436) );
  AOI21_X1 U45346 ( .A1(n29442), .A2(n31124), .B(n29441), .ZN(n29443) );
  NAND4_X2 U45348 ( .A1(n29447), .A2(n29446), .A3(n29445), .A4(n29444), .ZN(
        n30034) );
  NAND2_X1 U45349 ( .A1(n29839), .A2(n29450), .ZN(n29466) );
  OAI21_X1 U45351 ( .A1(n29458), .A2(n60028), .B(n22230), .ZN(n29459) );
  NAND2_X1 U45352 ( .A1(n29461), .A2(n29460), .ZN(n29462) );
  NAND2_X1 U45353 ( .A1(n31073), .A2(n29467), .ZN(n29469) );
  OAI21_X1 U45355 ( .A1(n61629), .A2(n25384), .B(n31089), .ZN(n29471) );
  NAND2_X1 U45356 ( .A1(n61382), .A2(n24504), .ZN(n29470) );
  NAND2_X1 U45358 ( .A1(n31083), .A2(n29472), .ZN(n29473) );
  AOI21_X1 U45359 ( .A1(n30421), .A2(n30422), .B(n29473), .ZN(n29476) );
  OAI21_X1 U45360 ( .A1(n61382), .A2(n31086), .B(n29474), .ZN(n29475) );
  NAND2_X1 U45361 ( .A1(n29476), .A2(n29475), .ZN(n29477) );
  NAND2_X1 U45362 ( .A1(n31141), .A2(n5768), .ZN(n30370) );
  NOR2_X1 U45363 ( .A1(n161), .A2(n64128), .ZN(n29488) );
  NOR2_X1 U45364 ( .A1(n31098), .A2(n10734), .ZN(n29494) );
  NOR3_X1 U45365 ( .A1(n161), .A2(n1868), .A3(n1856), .ZN(n29493) );
  NOR3_X1 U45366 ( .A1(n161), .A2(n1856), .A3(n59841), .ZN(n29492) );
  AOI22_X1 U45367 ( .A1(n31117), .A2(n29493), .B1(n29492), .B2(n31119), .ZN(
        n29496) );
  NOR2_X1 U45370 ( .A1(n22596), .A2(n30211), .ZN(n29525) );
  OAI21_X1 U45371 ( .A1(n61900), .A2(n29525), .B(n22416), .ZN(n29526) );
  NAND2_X1 U45373 ( .A1(n30479), .A2(n6609), .ZN(n29534) );
  NOR2_X1 U45374 ( .A1(n62647), .A2(n25848), .ZN(n29539) );
  OAI21_X1 U45375 ( .A1(n29539), .A2(n29538), .B(n30482), .ZN(n29540) );
  AOI21_X1 U45376 ( .A1(n29542), .A2(n29541), .B(n29540), .ZN(n29543) );
  INV_X1 U45377 ( .I(n29547), .ZN(n29544) );
  OAI22_X1 U45378 ( .A1(n29545), .A2(n29963), .B1(n21886), .B2(n29544), .ZN(
        n29550) );
  NAND3_X1 U45379 ( .A1(n21886), .A2(n29959), .A3(n20179), .ZN(n29549) );
  NAND2_X1 U45380 ( .A1(n29965), .A2(n21886), .ZN(n29548) );
  NAND2_X1 U45381 ( .A1(n30785), .A2(n29551), .ZN(n29553) );
  XOR2_X1 U45383 ( .A1(n1900), .A2(n50817), .Z(n52512) );
  XOR2_X1 U45384 ( .A1(n54376), .A2(n55052), .Z(n50798) );
  XOR2_X1 U45385 ( .A1(n52512), .A2(n50798), .Z(n31757) );
  XOR2_X1 U45386 ( .A1(n32560), .A2(n31757), .Z(n29557) );
  OAI22_X1 U45388 ( .A1(n29561), .A2(n29566), .B1(n31129), .B2(n9904), .ZN(
        n29562) );
  OAI21_X1 U45389 ( .A1(n29565), .A2(n60886), .B(n29912), .ZN(n29567) );
  NOR2_X1 U45392 ( .A1(n30296), .A2(n29575), .ZN(n29572) );
  OAI21_X1 U45393 ( .A1(n29572), .A2(n29571), .B(n29570), .ZN(n29574) );
  NOR2_X1 U45394 ( .A1(n23988), .A2(n29575), .ZN(n29577) );
  AOI22_X1 U45395 ( .A1(n29579), .A2(n29578), .B1(n29577), .B2(n63890), .ZN(
        n29583) );
  OAI21_X1 U45397 ( .A1(n65233), .A2(n29585), .B(n30613), .ZN(n29590) );
  NAND2_X1 U45400 ( .A1(n29588), .A2(n29587), .ZN(n29589) );
  AOI22_X1 U45402 ( .A1(n29593), .A2(n28915), .B1(n29592), .B2(n29591), .ZN(
        n29598) );
  NAND2_X1 U45403 ( .A1(n29596), .A2(n29595), .ZN(n29597) );
  NOR3_X1 U45404 ( .A1(n29601), .A2(n59099), .A3(n29600), .ZN(n29604) );
  OAI21_X1 U45405 ( .A1(n12739), .A2(n11873), .B(n29605), .ZN(n29612) );
  NOR2_X1 U45406 ( .A1(n29610), .A2(n29609), .ZN(n29611) );
  NAND3_X1 U45407 ( .A1(n19223), .A2(n59099), .A3(n61307), .ZN(n29615) );
  NAND2_X1 U45408 ( .A1(n23816), .A2(n24052), .ZN(n29620) );
  INV_X1 U45409 ( .I(n29621), .ZN(n29622) );
  NOR2_X1 U45410 ( .A1(n29629), .A2(n60894), .ZN(n29630) );
  NOR2_X1 U45411 ( .A1(n29631), .A2(n28125), .ZN(n29633) );
  NOR3_X1 U45412 ( .A1(n29647), .A2(n57781), .A3(n29671), .ZN(n29657) );
  INV_X1 U45413 ( .I(n29648), .ZN(n29649) );
  NAND2_X1 U45414 ( .A1(n29653), .A2(n58955), .ZN(n29654) );
  OAI21_X1 U45415 ( .A1(n29660), .A2(n29659), .B(n29658), .ZN(n29666) );
  NOR2_X1 U45416 ( .A1(n29661), .A2(n29663), .ZN(n29665) );
  NAND2_X1 U45418 ( .A1(n29670), .A2(n58601), .ZN(n29674) );
  NAND2_X1 U45419 ( .A1(n8296), .A2(n29671), .ZN(n29672) );
  NOR2_X1 U45420 ( .A1(n10598), .A2(n29695), .ZN(n29681) );
  INV_X1 U45421 ( .I(n29683), .ZN(n29686) );
  NAND2_X1 U45422 ( .A1(n29686), .A2(n29685), .ZN(n29687) );
  AOI21_X1 U45423 ( .A1(n29688), .A2(n29698), .B(n29687), .ZN(n29701) );
  OAI21_X1 U45424 ( .A1(n29691), .A2(n25341), .B(n22214), .ZN(n29692) );
  NOR3_X1 U45425 ( .A1(n29698), .A2(n29697), .A3(n29696), .ZN(n29699) );
  NOR2_X1 U45426 ( .A1(n29704), .A2(n4848), .ZN(n29706) );
  OAI21_X1 U45428 ( .A1(n31277), .A2(n6317), .B(n31264), .ZN(n29718) );
  AOI22_X1 U45429 ( .A1(n30877), .A2(n29718), .B1(n31279), .B2(n6317), .ZN(
        n29719) );
  NOR2_X1 U45430 ( .A1(n12443), .A2(n23008), .ZN(n29722) );
  OAI21_X1 U45431 ( .A1(n9654), .A2(n1561), .B(n12893), .ZN(n29721) );
  OAI21_X1 U45432 ( .A1(n30496), .A2(n30890), .B(n30889), .ZN(n29724) );
  NAND2_X1 U45433 ( .A1(n30026), .A2(n22748), .ZN(n29728) );
  OAI21_X1 U45434 ( .A1(n29729), .A2(n29728), .B(n30023), .ZN(n29735) );
  AOI21_X1 U45435 ( .A1(n29733), .A2(n29732), .B(n29731), .ZN(n29734) );
  NAND2_X1 U45437 ( .A1(n10629), .A2(n1559), .ZN(n29739) );
  NAND2_X1 U45438 ( .A1(n21263), .A2(n1559), .ZN(n29740) );
  OAI21_X1 U45441 ( .A1(n29963), .A2(n18472), .B(n29744), .ZN(n29746) );
  NOR2_X1 U45442 ( .A1(n21886), .A2(n30767), .ZN(n29745) );
  OAI21_X1 U45443 ( .A1(n29746), .A2(n29745), .B(n20179), .ZN(n29752) );
  NOR2_X1 U45444 ( .A1(n29748), .A2(n29747), .ZN(n29749) );
  OAI21_X1 U45445 ( .A1(n30780), .A2(n30779), .B(n29750), .ZN(n29751) );
  XOR2_X1 U45447 ( .A1(n53685), .A2(n55580), .Z(n32053) );
  XOR2_X1 U45448 ( .A1(n55087), .A2(n53174), .Z(n31643) );
  XOR2_X1 U45449 ( .A1(n32053), .A2(n31643), .Z(n38472) );
  XOR2_X1 U45450 ( .A1(n38472), .A2(n54407), .Z(n38904) );
  XOR2_X1 U45451 ( .A1(n54185), .A2(n54748), .Z(n50943) );
  XOR2_X1 U45452 ( .A1(n56714), .A2(n56097), .Z(n51275) );
  XOR2_X1 U45453 ( .A1(n50943), .A2(n51275), .Z(n34834) );
  INV_X1 U45454 ( .I(n55810), .ZN(n50655) );
  XOR2_X1 U45455 ( .A1(n50655), .A2(n51946), .Z(n30716) );
  INV_X1 U45456 ( .I(n30716), .ZN(n50682) );
  XOR2_X1 U45457 ( .A1(n34834), .A2(n50682), .Z(n37993) );
  XOR2_X1 U45458 ( .A1(n38904), .A2(n37993), .Z(n50987) );
  CLKBUF_X4 U45459 ( .I(Key[76]), .Z(n54563) );
  XOR2_X1 U45460 ( .A1(n24109), .A2(n56508), .Z(n38752) );
  XOR2_X1 U45461 ( .A1(n39349), .A2(n38752), .Z(n52354) );
  CLKBUF_X4 U45462 ( .I(Key[88]), .Z(n54917) );
  XOR2_X1 U45463 ( .A1(n55379), .A2(n54917), .Z(n51530) );
  XOR2_X1 U45464 ( .A1(n51530), .A2(n53989), .Z(n29754) );
  XOR2_X1 U45465 ( .A1(n52354), .A2(n29754), .Z(n44746) );
  XOR2_X1 U45466 ( .A1(n50987), .A2(n44746), .Z(n29763) );
  NAND2_X1 U45471 ( .A1(n30254), .A2(n8602), .ZN(n29759) );
  XOR2_X1 U45472 ( .A1(n29763), .A2(n32338), .Z(n29764) );
  XOR2_X1 U45473 ( .A1(n30715), .A2(n29764), .Z(n29765) );
  NOR2_X1 U45474 ( .A1(n29766), .A2(n17495), .ZN(n29770) );
  NOR2_X1 U45475 ( .A1(n29767), .A2(n30124), .ZN(n29769) );
  NOR2_X1 U45476 ( .A1(n1351), .A2(n1872), .ZN(n29771) );
  NOR2_X1 U45477 ( .A1(n29772), .A2(n29771), .ZN(n29776) );
  NAND3_X2 U45478 ( .A1(n29777), .A2(n29776), .A3(n29775), .ZN(n33904) );
  NOR2_X1 U45479 ( .A1(n29778), .A2(n63272), .ZN(n29792) );
  INV_X1 U45480 ( .I(n29780), .ZN(n29781) );
  OAI21_X2 U45482 ( .A1(n29792), .A2(n29791), .B(n29790), .ZN(n32266) );
  XOR2_X1 U45483 ( .A1(n32266), .A2(n33904), .Z(n29804) );
  INV_X1 U45486 ( .I(n29800), .ZN(n29803) );
  XOR2_X1 U45487 ( .A1(n1824), .A2(n29804), .Z(n29818) );
  NAND3_X1 U45488 ( .A1(n30213), .A2(n770), .A3(n30224), .ZN(n29810) );
  NOR2_X1 U45489 ( .A1(n29805), .A2(n30841), .ZN(n29807) );
  NOR2_X1 U45490 ( .A1(n30217), .A2(n30841), .ZN(n29806) );
  NAND2_X1 U45491 ( .A1(n22596), .A2(n22416), .ZN(n29811) );
  NAND2_X1 U45492 ( .A1(n14230), .A2(n30319), .ZN(n29996) );
  NAND2_X1 U45493 ( .A1(n29995), .A2(n64154), .ZN(n29822) );
  INV_X1 U45494 ( .I(n29823), .ZN(n29825) );
  NOR3_X1 U45495 ( .A1(n16961), .A2(n29825), .A3(n29824), .ZN(n29827) );
  OAI21_X1 U45496 ( .A1(n30815), .A2(n30809), .B(n8521), .ZN(n29833) );
  OAI21_X1 U45497 ( .A1(n30816), .A2(n11830), .B(n29833), .ZN(n29837) );
  NAND2_X1 U45498 ( .A1(n29839), .A2(n29838), .ZN(n29853) );
  INV_X1 U45499 ( .I(n29844), .ZN(n29847) );
  OAI21_X1 U45500 ( .A1(n29847), .A2(n29846), .B(n29845), .ZN(n29850) );
  INV_X1 U45501 ( .I(n29848), .ZN(n29849) );
  NAND2_X1 U45502 ( .A1(n29850), .A2(n29849), .ZN(n29851) );
  NAND2_X1 U45504 ( .A1(n18736), .A2(n17412), .ZN(n29859) );
  NAND2_X1 U45505 ( .A1(n29861), .A2(n63891), .ZN(n29865) );
  NOR2_X1 U45507 ( .A1(n1538), .A2(n57774), .ZN(n29869) );
  NAND2_X1 U45508 ( .A1(n29871), .A2(n24077), .ZN(n29872) );
  INV_X1 U45509 ( .I(n29875), .ZN(n31306) );
  NOR2_X1 U45510 ( .A1(n61753), .A2(n30027), .ZN(n29883) );
  XOR2_X1 U45512 ( .A1(n30550), .A2(n54776), .Z(n29885) );
  BUF_X2 U45513 ( .I(n29892), .Z(n44533) );
  XOR2_X1 U45514 ( .A1(n53705), .A2(n52232), .Z(n38126) );
  XOR2_X1 U45515 ( .A1(n44533), .A2(n38126), .Z(n37786) );
  INV_X1 U45516 ( .I(n50067), .ZN(n29893) );
  XOR2_X1 U45517 ( .A1(n37786), .A2(n29893), .Z(n39400) );
  INV_X1 U45518 ( .I(n39400), .ZN(n29894) );
  XOR2_X1 U45519 ( .A1(n56745), .A2(n57162), .Z(n45371) );
  XOR2_X1 U45522 ( .A1(n45371), .A2(n52375), .Z(n38009) );
  XOR2_X1 U45523 ( .A1(n29894), .A2(n38009), .Z(n38662) );
  XOR2_X1 U45524 ( .A1(n38662), .A2(n23455), .Z(n51575) );
  XOR2_X1 U45525 ( .A1(n38450), .A2(n56819), .Z(n50197) );
  XOR2_X1 U45526 ( .A1(n56202), .A2(n54289), .Z(n31068) );
  XOR2_X1 U45527 ( .A1(n31068), .A2(n53308), .Z(n29895) );
  XOR2_X1 U45528 ( .A1(n50197), .A2(n29895), .Z(n44462) );
  XOR2_X1 U45529 ( .A1(n51575), .A2(n44462), .Z(n29907) );
  NAND2_X1 U45532 ( .A1(n29901), .A2(n29900), .ZN(n29903) );
  XOR2_X1 U45533 ( .A1(n29907), .A2(n11529), .Z(n29908) );
  NAND2_X1 U45534 ( .A1(n24000), .A2(n27150), .ZN(n29913) );
  NOR2_X1 U45535 ( .A1(n59613), .A2(n29914), .ZN(n29918) );
  OAI21_X1 U45536 ( .A1(n9904), .A2(n24000), .B(n59613), .ZN(n29917) );
  MUX2_X1 U45537 ( .I0(n29920), .I1(n29919), .S(n61251), .Z(n29923) );
  NOR2_X1 U45538 ( .A1(n25013), .A2(n4257), .ZN(n30511) );
  NAND2_X1 U45539 ( .A1(n31270), .A2(n31277), .ZN(n30875) );
  NAND2_X1 U45541 ( .A1(n2636), .A2(n21626), .ZN(n29924) );
  INV_X1 U45543 ( .I(n30532), .ZN(n29931) );
  NOR2_X1 U45544 ( .A1(n29931), .A2(n10821), .ZN(n29939) );
  INV_X1 U45548 ( .I(n29943), .ZN(n29945) );
  NAND2_X1 U45549 ( .A1(n3086), .A2(n30408), .ZN(n29944) );
  NOR2_X1 U45550 ( .A1(n29950), .A2(n29949), .ZN(n29951) );
  OAI21_X1 U45551 ( .A1(n29956), .A2(n24206), .B(n29955), .ZN(n29967) );
  XOR2_X1 U45553 ( .A1(n38733), .A2(n56859), .Z(n30527) );
  XOR2_X1 U45554 ( .A1(n22950), .A2(n55777), .Z(n29968) );
  XOR2_X1 U45555 ( .A1(n30527), .A2(n29968), .Z(n44339) );
  CLKBUF_X4 U45556 ( .I(Key[50]), .Z(n53958) );
  XOR2_X1 U45557 ( .A1(n54536), .A2(n53958), .Z(n29969) );
  XOR2_X1 U45558 ( .A1(n54896), .A2(n56915), .Z(n38407) );
  XOR2_X1 U45559 ( .A1(n29969), .A2(n38407), .Z(n29970) );
  XOR2_X1 U45560 ( .A1(n53076), .A2(n53487), .Z(n45379) );
  XOR2_X1 U45561 ( .A1(n29970), .A2(n45379), .Z(n29971) );
  XOR2_X1 U45562 ( .A1(n44339), .A2(n29971), .Z(n29973) );
  CLKBUF_X4 U45563 ( .I(Key[134]), .Z(n55876) );
  XOR2_X1 U45564 ( .A1(n55876), .A2(n56475), .Z(n38154) );
  XOR2_X1 U45565 ( .A1(n56165), .A2(n55610), .Z(n29972) );
  XOR2_X1 U45566 ( .A1(n38154), .A2(n15735), .Z(n39771) );
  CLKBUF_X4 U45567 ( .I(Key[110]), .Z(n55349) );
  XOR2_X1 U45568 ( .A1(n55126), .A2(n55349), .Z(n32344) );
  XOR2_X1 U45569 ( .A1(n39771), .A2(n32344), .Z(n39387) );
  XOR2_X1 U45570 ( .A1(n29973), .A2(n59680), .Z(n29974) );
  NOR2_X1 U45572 ( .A1(n23478), .A2(n1277), .ZN(n29978) );
  NOR2_X1 U45573 ( .A1(n1860), .A2(n29981), .ZN(n29983) );
  NOR2_X1 U45574 ( .A1(n1277), .A2(n30537), .ZN(n29982) );
  NAND2_X1 U45576 ( .A1(n30322), .A2(n29988), .ZN(n29989) );
  NOR3_X1 U45577 ( .A1(n29994), .A2(n29993), .A3(n23397), .ZN(n29997) );
  NOR2_X1 U45579 ( .A1(n7426), .A2(n30752), .ZN(n30007) );
  OAI21_X1 U45580 ( .A1(n30663), .A2(n30755), .B(n30007), .ZN(n30010) );
  INV_X1 U45582 ( .I(n30020), .ZN(n30022) );
  OAI21_X1 U45583 ( .A1(n30031), .A2(n30030), .B(n30029), .ZN(n30032) );
  XOR2_X1 U45584 ( .A1(n32642), .A2(n32560), .Z(n30035) );
  XOR2_X1 U45585 ( .A1(n53748), .A2(n22691), .Z(n52197) );
  XOR2_X1 U45588 ( .A1(n52294), .A2(n51569), .Z(n30036) );
  XOR2_X1 U45589 ( .A1(n36632), .A2(n30036), .Z(n37981) );
  INV_X1 U45590 ( .I(n37981), .ZN(n30039) );
  XOR2_X1 U45591 ( .A1(n50661), .A2(n24065), .Z(n31649) );
  INV_X1 U45592 ( .I(n31649), .ZN(n39631) );
  XOR2_X1 U45593 ( .A1(n39631), .A2(n54219), .Z(n44426) );
  XOR2_X1 U45594 ( .A1(n53064), .A2(n53477), .Z(n39555) );
  XOR2_X1 U45595 ( .A1(n15707), .A2(n23989), .Z(n30037) );
  XOR2_X1 U45596 ( .A1(n44426), .A2(n30037), .Z(n30038) );
  XOR2_X1 U45597 ( .A1(n30039), .A2(n30038), .Z(n30041) );
  XOR2_X1 U45598 ( .A1(n56683), .A2(n56309), .Z(n51542) );
  XOR2_X1 U45599 ( .A1(n54376), .A2(n54143), .Z(n51665) );
  XOR2_X1 U45600 ( .A1(n51542), .A2(n51665), .Z(n44427) );
  INV_X1 U45601 ( .I(n52512), .ZN(n50533) );
  XOR2_X1 U45602 ( .A1(n50533), .A2(n60797), .Z(n46593) );
  XOR2_X1 U45603 ( .A1(n44427), .A2(n46593), .Z(n30040) );
  XOR2_X1 U45604 ( .A1(n30041), .A2(n30040), .Z(n30042) );
  XOR2_X1 U45605 ( .A1(n30043), .A2(n33186), .Z(n30044) );
  XOR2_X1 U45606 ( .A1(n30045), .A2(n30044), .Z(n30070) );
  INV_X1 U45607 ( .I(n30258), .ZN(n30049) );
  AOI21_X1 U45608 ( .A1(n30058), .A2(n30057), .B(n30056), .ZN(n30069) );
  NOR2_X1 U45609 ( .A1(n31059), .A2(n58999), .ZN(n30059) );
  INV_X1 U45610 ( .I(n30161), .ZN(n30062) );
  NOR2_X1 U45611 ( .A1(n30691), .A2(n17627), .ZN(n30061) );
  INV_X1 U45614 ( .I(n30063), .ZN(n30066) );
  INV_X1 U45615 ( .I(n30064), .ZN(n30065) );
  INV_X1 U45616 ( .I(n30071), .ZN(n30072) );
  AOI21_X1 U45617 ( .A1(n30072), .A2(n60262), .B(n7423), .ZN(n30081) );
  OAI21_X1 U45618 ( .A1(n25241), .A2(n30086), .B(n30085), .ZN(n30090) );
  OAI21_X1 U45619 ( .A1(n60262), .A2(n21062), .B(n64589), .ZN(n30088) );
  NAND2_X1 U45620 ( .A1(n30195), .A2(n30192), .ZN(n30097) );
  OAI21_X1 U45621 ( .A1(n30097), .A2(n30197), .B(n30183), .ZN(n30098) );
  NOR2_X1 U45622 ( .A1(n21019), .A2(n58430), .ZN(n30102) );
  AOI22_X1 U45623 ( .A1(n30705), .A2(n30102), .B1(n30701), .B2(n58430), .ZN(
        n30107) );
  NOR2_X1 U45624 ( .A1(n31041), .A2(n31038), .ZN(n30103) );
  NAND3_X1 U45626 ( .A1(n31031), .A2(n31037), .A3(n31038), .ZN(n30105) );
  NAND3_X1 U45627 ( .A1(n30107), .A2(n30106), .A3(n30105), .ZN(n30111) );
  AOI21_X1 U45628 ( .A1(n30112), .A2(n12743), .B(n30109), .ZN(n30110) );
  NOR2_X1 U45629 ( .A1(n30111), .A2(n30110), .ZN(n30119) );
  INV_X1 U45630 ( .I(n30112), .ZN(n30117) );
  INV_X1 U45631 ( .I(n30142), .ZN(n30116) );
  INV_X1 U45632 ( .I(n31032), .ZN(n30113) );
  NAND2_X1 U45633 ( .A1(n30113), .A2(n31042), .ZN(n30114) );
  NOR2_X1 U45634 ( .A1(n30705), .A2(n30114), .ZN(n30115) );
  OAI21_X1 U45635 ( .A1(n30117), .A2(n30116), .B(n30115), .ZN(n30118) );
  MUX2_X1 U45636 ( .I0(n30121), .I1(n30120), .S(n1872), .Z(n30131) );
  AOI21_X1 U45637 ( .A1(n8982), .A2(n1351), .B(n30123), .ZN(n30129) );
  NOR3_X1 U45638 ( .A1(n21559), .A2(n30523), .A3(n30124), .ZN(n30128) );
  INV_X1 U45639 ( .I(n30149), .ZN(n30132) );
  NOR2_X1 U45640 ( .A1(n30132), .A2(n22322), .ZN(n30140) );
  NOR2_X1 U45641 ( .A1(n23056), .A2(n31038), .ZN(n30133) );
  AOI22_X1 U45642 ( .A1(n30134), .A2(n31038), .B1(n61376), .B2(n30133), .ZN(
        n30139) );
  NAND2_X1 U45643 ( .A1(n31035), .A2(n31039), .ZN(n30136) );
  AOI21_X1 U45644 ( .A1(n30140), .A2(n30139), .B(n30138), .ZN(n30156) );
  AND2_X1 U45645 ( .A1(n30141), .A2(n61376), .Z(n30144) );
  INV_X1 U45647 ( .I(n30700), .ZN(n30143) );
  NAND4_X1 U45648 ( .A1(n30704), .A2(n21019), .A3(n21176), .A4(n23056), .ZN(
        n30147) );
  NOR4_X1 U45649 ( .A1(n30150), .A2(n30149), .A3(n31038), .A4(n21176), .ZN(
        n30152) );
  XOR2_X1 U45651 ( .A1(n53154), .A2(n23858), .Z(n42812) );
  XOR2_X1 U45652 ( .A1(n24057), .A2(n4561), .Z(n30157) );
  BUF_X2 U45653 ( .I(n30157), .Z(n52095) );
  XOR2_X1 U45654 ( .A1(n42812), .A2(n30157), .Z(n44841) );
  INV_X1 U45655 ( .I(n30163), .ZN(n30164) );
  AOI21_X1 U45656 ( .A1(n30166), .A2(n30165), .B(n18839), .ZN(n30172) );
  NOR2_X1 U45659 ( .A1(n30182), .A2(n57436), .ZN(n30189) );
  OAI21_X1 U45664 ( .A1(n59798), .A2(n1559), .B(n30195), .ZN(n30199) );
  NAND3_X1 U45665 ( .A1(n30199), .A2(n30198), .A3(n30197), .ZN(n30201) );
  XOR2_X1 U45666 ( .A1(n54168), .A2(n54734), .Z(n38885) );
  CLKBUF_X4 U45667 ( .I(Key[141]), .Z(n56065) );
  XOR2_X1 U45668 ( .A1(n56702), .A2(n56065), .Z(n30205) );
  BUF_X2 U45669 ( .I(n30205), .Z(n52135) );
  XOR2_X1 U45670 ( .A1(n38885), .A2(n52135), .Z(n37630) );
  XOR2_X1 U45672 ( .A1(n37630), .A2(n52029), .Z(n50129) );
  INV_X1 U45673 ( .I(n50129), .ZN(n30206) );
  XOR2_X1 U45674 ( .A1(n30206), .A2(n52734), .Z(n44843) );
  XOR2_X1 U45675 ( .A1(n56495), .A2(n54556), .Z(n38215) );
  XOR2_X1 U45676 ( .A1(n39724), .A2(n38215), .Z(n46349) );
  XOR2_X1 U45677 ( .A1(n44843), .A2(n46349), .Z(n30207) );
  XOR2_X1 U45678 ( .A1(n30209), .A2(n32716), .Z(n30210) );
  NAND4_X1 U45679 ( .A1(n30846), .A2(n30212), .A3(n22416), .A4(n30211), .ZN(
        n30218) );
  NAND3_X1 U45680 ( .A1(n30839), .A2(n61900), .A3(n1869), .ZN(n30228) );
  AOI21_X1 U45681 ( .A1(n30238), .A2(n30237), .B(n30685), .ZN(n30241) );
  INV_X1 U45682 ( .I(n30239), .ZN(n30240) );
  OAI22_X1 U45683 ( .A1(n60146), .A2(n16631), .B1(n30255), .B2(n21626), .ZN(
        n30259) );
  AOI21_X1 U45684 ( .A1(n30266), .A2(n30265), .B(n61734), .ZN(n30269) );
  OAI21_X1 U45685 ( .A1(n30271), .A2(n23317), .B(n22139), .ZN(n30268) );
  NAND4_X1 U45686 ( .A1(n61734), .A2(n30271), .A3(n14389), .A4(n30276), .ZN(
        n30274) );
  NAND3_X1 U45690 ( .A1(n1562), .A2(n23734), .A3(n13731), .ZN(n30295) );
  NAND2_X1 U45691 ( .A1(n30301), .A2(n30300), .ZN(n30307) );
  NOR2_X1 U45692 ( .A1(n30305), .A2(n30304), .ZN(n30306) );
  INV_X1 U45693 ( .I(n30308), .ZN(n30310) );
  NAND2_X1 U45694 ( .A1(n30312), .A2(n1875), .ZN(n30309) );
  NAND2_X1 U45696 ( .A1(n1278), .A2(n31224), .ZN(n30758) );
  OAI21_X1 U45697 ( .A1(n30760), .A2(n15738), .B(n30752), .ZN(n30314) );
  AOI21_X1 U45699 ( .A1(n30330), .A2(n30333), .B(n30329), .ZN(n30337) );
  NAND2_X1 U45702 ( .A1(n30348), .A2(n10240), .ZN(n30607) );
  INV_X1 U45703 ( .I(n30607), .ZN(n30349) );
  XOR2_X1 U45705 ( .A1(n44995), .A2(n54360), .Z(n36736) );
  XOR2_X1 U45706 ( .A1(n36736), .A2(n56827), .Z(n37952) );
  XOR2_X1 U45707 ( .A1(n23851), .A2(n52970), .Z(n30355) );
  XOR2_X1 U45708 ( .A1(n55034), .A2(n55516), .Z(n37468) );
  XOR2_X1 U45709 ( .A1(n15710), .A2(n37468), .Z(n37584) );
  XOR2_X1 U45710 ( .A1(n53641), .A2(n51493), .Z(n30356) );
  BUF_X2 U45711 ( .I(n30356), .Z(n38653) );
  INV_X1 U45712 ( .I(n30356), .ZN(n31444) );
  XOR2_X1 U45713 ( .A1(n56008), .A2(n50494), .Z(n39375) );
  XOR2_X1 U45714 ( .A1(n31444), .A2(n39375), .Z(n31558) );
  INV_X1 U45715 ( .I(n31558), .ZN(n37758) );
  XOR2_X1 U45718 ( .A1(n54517), .A2(n51492), .Z(n38560) );
  XOR2_X1 U45719 ( .A1(n38826), .A2(n38560), .Z(n50998) );
  XOR2_X1 U45720 ( .A1(n50998), .A2(n37303), .Z(n44123) );
  XOR2_X1 U45721 ( .A1(n44123), .A2(n55335), .Z(n30358) );
  XOR2_X1 U45722 ( .A1(n43398), .A2(n30358), .Z(n30359) );
  XOR2_X1 U45723 ( .A1(n32089), .A2(n30359), .Z(n30365) );
  MUX2_X1 U45724 ( .I0(n30374), .I1(n30368), .S(n30585), .Z(n30381) );
  NOR2_X1 U45725 ( .A1(n24172), .A2(n31137), .ZN(n30373) );
  AOI21_X1 U45726 ( .A1(n30374), .A2(n30369), .B(n495), .ZN(n30372) );
  NOR2_X1 U45727 ( .A1(n30370), .A2(n31137), .ZN(n30371) );
  OAI22_X1 U45728 ( .A1(n30378), .A2(n30377), .B1(n61007), .B2(n30375), .ZN(
        n30379) );
  NOR2_X1 U45729 ( .A1(n57437), .A2(n64484), .ZN(n30382) );
  OAI21_X1 U45730 ( .A1(n14276), .A2(n30383), .B(n30382), .ZN(n30389) );
  NAND2_X1 U45731 ( .A1(n31110), .A2(n31115), .ZN(n30387) );
  CLKBUF_X4 U45732 ( .I(Key[100]), .Z(n55150) );
  XOR2_X1 U45733 ( .A1(n54563), .A2(n55150), .Z(n39228) );
  XOR2_X1 U45734 ( .A1(n52470), .A2(n39228), .Z(n31318) );
  XOR2_X1 U45735 ( .A1(n31397), .A2(n51530), .Z(n37635) );
  XOR2_X1 U45737 ( .A1(n53284), .A2(n56949), .Z(n37637) );
  XOR2_X1 U45738 ( .A1(n56714), .A2(n54407), .Z(n37638) );
  XOR2_X1 U45739 ( .A1(n55087), .A2(n55580), .Z(n43858) );
  XOR2_X1 U45740 ( .A1(n43858), .A2(n50943), .Z(n43262) );
  CLKBUF_X4 U45741 ( .I(Key[136]), .Z(n55889) );
  XOR2_X1 U45742 ( .A1(n43262), .A2(n55889), .Z(n30403) );
  XOR2_X1 U45743 ( .A1(n44100), .A2(n30403), .Z(n30404) );
  XOR2_X1 U45744 ( .A1(n30404), .A2(n23714), .Z(n30406) );
  XOR2_X1 U45745 ( .A1(n31487), .A2(n15733), .Z(n30405) );
  XOR2_X1 U45746 ( .A1(n30406), .A2(n30405), .Z(n30407) );
  AOI21_X1 U45747 ( .A1(n30416), .A2(n30415), .B(n30640), .ZN(n30417) );
  NOR3_X1 U45748 ( .A1(n30421), .A2(n58931), .A3(n22878), .ZN(n30427) );
  NAND2_X1 U45749 ( .A1(n5267), .A2(n31086), .ZN(n30425) );
  NAND2_X1 U45751 ( .A1(n31083), .A2(n24504), .ZN(n30423) );
  AOI21_X1 U45756 ( .A1(n30560), .A2(n31083), .B(n30430), .ZN(n30431) );
  OAI21_X1 U45757 ( .A1(n1852), .A2(n31083), .B(n30431), .ZN(n30432) );
  INV_X1 U45760 ( .I(n30438), .ZN(n30440) );
  INV_X1 U45762 ( .I(n30447), .ZN(n30448) );
  NOR2_X1 U45763 ( .A1(n61048), .A2(n30455), .ZN(n30457) );
  NOR2_X1 U45764 ( .A1(n30467), .A2(n18300), .ZN(n30460) );
  NAND2_X1 U45768 ( .A1(n30467), .A2(n18300), .ZN(n30461) );
  NOR2_X1 U45770 ( .A1(n33720), .A2(n2033), .ZN(n30468) );
  INV_X1 U45773 ( .I(n34070), .ZN(n30469) );
  NAND3_X1 U45779 ( .A1(n19451), .A2(n1352), .A3(n5070), .ZN(n30493) );
  OAI21_X1 U45780 ( .A1(n30884), .A2(n1561), .B(n30497), .ZN(n30498) );
  NOR2_X1 U45781 ( .A1(n31241), .A2(n5933), .ZN(n30502) );
  AOI22_X1 U45786 ( .A1(n30513), .A2(n65051), .B1(n30511), .B2(n61251), .ZN(
        n30514) );
  NAND2_X1 U45787 ( .A1(n1872), .A2(n7026), .ZN(n30518) );
  XOR2_X1 U45789 ( .A1(n55777), .A2(n53138), .Z(n32189) );
  XOR2_X1 U45790 ( .A1(n37513), .A2(n32189), .Z(n38962) );
  XOR2_X1 U45791 ( .A1(n38962), .A2(n22950), .Z(n32987) );
  XOR2_X1 U45792 ( .A1(n32987), .A2(n30527), .Z(n50102) );
  XOR2_X1 U45793 ( .A1(n56475), .A2(n55349), .Z(n30528) );
  XOR2_X1 U45794 ( .A1(n30528), .A2(n56771), .Z(n43759) );
  XOR2_X1 U45795 ( .A1(n54896), .A2(n54536), .Z(n30530) );
  XOR2_X1 U45796 ( .A1(n53958), .A2(n54231), .Z(n30529) );
  XOR2_X1 U45797 ( .A1(n30530), .A2(n30529), .Z(n31347) );
  INV_X1 U45798 ( .I(n31347), .ZN(n43900) );
  XOR2_X1 U45799 ( .A1(n30536), .A2(n32354), .Z(n31885) );
  NAND2_X1 U45800 ( .A1(n31076), .A2(n24504), .ZN(n30554) );
  AOI21_X1 U45801 ( .A1(n30552), .A2(n22411), .B(n30551), .ZN(n30553) );
  MUX2_X1 U45802 ( .I0(n30554), .I1(n30553), .S(n25384), .Z(n30563) );
  NOR2_X1 U45804 ( .A1(n30555), .A2(n31081), .ZN(n30557) );
  NOR3_X1 U45805 ( .A1(n31089), .A2(n31083), .A3(n30560), .ZN(n30561) );
  CLKBUF_X4 U45806 ( .I(Key[137]), .Z(n55903) );
  CLKBUF_X4 U45807 ( .I(Key[89]), .Z(n54936) );
  XOR2_X1 U45808 ( .A1(n54289), .A2(n54936), .Z(n37713) );
  XOR2_X1 U45809 ( .A1(n45371), .A2(n55833), .Z(n30565) );
  XOR2_X1 U45810 ( .A1(n46276), .A2(n30565), .Z(n30570) );
  XOR2_X1 U45811 ( .A1(n53308), .A2(n53530), .Z(n37737) );
  XOR2_X1 U45812 ( .A1(n56202), .A2(n24061), .Z(n30566) );
  XOR2_X1 U45813 ( .A1(n37737), .A2(n30566), .Z(n30567) );
  XOR2_X1 U45814 ( .A1(n30567), .A2(n38450), .Z(n30569) );
  XOR2_X1 U45815 ( .A1(n33063), .A2(n30568), .Z(n38380) );
  XOR2_X1 U45816 ( .A1(n30569), .A2(n38380), .Z(n44291) );
  XOR2_X1 U45817 ( .A1(n30570), .A2(n44291), .Z(n30571) );
  NAND2_X1 U45820 ( .A1(n30574), .A2(n31118), .ZN(n30575) );
  NAND2_X1 U45821 ( .A1(n30576), .A2(n31102), .ZN(n30582) );
  AOI22_X1 U45822 ( .A1(n22627), .A2(n30594), .B1(n30593), .B2(n31146), .ZN(
        n30595) );
  XOR2_X1 U45823 ( .A1(n30598), .A2(n30597), .Z(n30599) );
  XOR2_X1 U45825 ( .A1(n53787), .A2(n24067), .Z(n30601) );
  BUF_X2 U45826 ( .I(n30601), .Z(n52196) );
  XOR2_X1 U45827 ( .A1(n56309), .A2(n55765), .Z(n37651) );
  XOR2_X1 U45828 ( .A1(n52196), .A2(n37651), .Z(n52592) );
  INV_X1 U45829 ( .I(n52592), .ZN(n30603) );
  XOR2_X1 U45831 ( .A1(n52080), .A2(n61737), .Z(n39635) );
  XOR2_X1 U45832 ( .A1(n30603), .A2(n39635), .Z(n44602) );
  XOR2_X1 U45833 ( .A1(n46414), .A2(n46593), .Z(n45395) );
  XOR2_X1 U45834 ( .A1(n52294), .A2(n53945), .Z(n44330) );
  XOR2_X1 U45835 ( .A1(n45395), .A2(n44330), .Z(n38533) );
  XOR2_X1 U45836 ( .A1(n55862), .A2(n53748), .Z(n39445) );
  XOR2_X1 U45837 ( .A1(n39445), .A2(n51611), .Z(n39263) );
  XOR2_X1 U45838 ( .A1(n39263), .A2(n23989), .Z(n44332) );
  XOR2_X1 U45839 ( .A1(n38533), .A2(n44332), .Z(n30604) );
  NAND2_X1 U45841 ( .A1(n30607), .A2(n30606), .ZN(n30627) );
  INV_X1 U45844 ( .I(n30614), .ZN(n30622) );
  NAND2_X1 U45846 ( .A1(n30619), .A2(n30618), .ZN(n30625) );
  OAI21_X1 U45847 ( .A1(n30623), .A2(n30622), .B(n30621), .ZN(n30624) );
  NAND2_X1 U45848 ( .A1(n13280), .A2(n24564), .ZN(n30629) );
  AOI21_X1 U45849 ( .A1(n14217), .A2(n31208), .B(n30629), .ZN(n30630) );
  NAND3_X1 U45850 ( .A1(n13280), .A2(n1432), .A3(n31208), .ZN(n30636) );
  AOI21_X1 U45851 ( .A1(n31206), .A2(n30636), .B(n31209), .ZN(n30637) );
  INV_X1 U45852 ( .I(n30640), .ZN(n30642) );
  INV_X1 U45856 ( .I(n30655), .ZN(n30656) );
  NAND2_X1 U45860 ( .A1(n30668), .A2(n61215), .ZN(n30671) );
  INV_X1 U45861 ( .I(n30669), .ZN(n30670) );
  AOI21_X1 U45863 ( .A1(n30676), .A2(n18198), .B(n30675), .ZN(n30682) );
  NAND2_X1 U45864 ( .A1(n10431), .A2(n10525), .ZN(n30686) );
  OAI21_X1 U45865 ( .A1(n30688), .A2(n31049), .B(n30687), .ZN(n30693) );
  OAI22_X1 U45866 ( .A1(n30691), .A2(n58999), .B1(n20918), .B2(n30689), .ZN(
        n30692) );
  OAI21_X1 U45867 ( .A1(n30693), .A2(n30692), .B(n17627), .ZN(n30699) );
  NAND2_X1 U45868 ( .A1(n31046), .A2(n1858), .ZN(n30697) );
  NOR2_X1 U45869 ( .A1(n30702), .A2(n16279), .ZN(n30703) );
  AOI22_X1 U45870 ( .A1(n30705), .A2(n30704), .B1(n23072), .B2(n30703), .ZN(
        n30713) );
  INV_X1 U45872 ( .I(n30709), .ZN(n31034) );
  NAND3_X1 U45873 ( .A1(n30710), .A2(n31034), .A3(n1315), .ZN(n30711) );
  XOR2_X1 U45874 ( .A1(n53359), .A2(n57142), .Z(n51977) );
  XOR2_X1 U45875 ( .A1(n30716), .A2(n51977), .Z(n30932) );
  XOR2_X1 U45876 ( .A1(n1881), .A2(n56714), .Z(n52461) );
  XOR2_X1 U45877 ( .A1(n61380), .A2(n53833), .Z(n39434) );
  XOR2_X1 U45879 ( .A1(n39434), .A2(n56335), .Z(n31230) );
  XOR2_X1 U45880 ( .A1(n43262), .A2(n31230), .Z(n37836) );
  XOR2_X1 U45882 ( .A1(n31397), .A2(n56508), .Z(n42730) );
  XOR2_X1 U45883 ( .A1(n42730), .A2(n53989), .Z(n30717) );
  NOR2_X1 U45884 ( .A1(n30723), .A2(n23772), .ZN(n30729) );
  NAND2_X1 U45887 ( .A1(n21906), .A2(n30832), .ZN(n30831) );
  NAND2_X1 U45889 ( .A1(n30763), .A2(n59046), .ZN(n30765) );
  NAND2_X1 U45890 ( .A1(n30768), .A2(n30767), .ZN(n30774) );
  INV_X1 U45891 ( .I(n30769), .ZN(n30772) );
  NAND2_X1 U45892 ( .A1(n30778), .A2(n20179), .ZN(n30783) );
  INV_X1 U45894 ( .I(n30788), .ZN(n30789) );
  XOR2_X1 U45895 ( .A1(n52135), .A2(n54168), .Z(n52327) );
  XOR2_X1 U45896 ( .A1(n56495), .A2(n54249), .Z(n50245) );
  INV_X1 U45897 ( .I(n15712), .ZN(n50724) );
  CLKBUF_X4 U45898 ( .I(Key[147]), .Z(n56180) );
  XOR2_X1 U45899 ( .A1(n56784), .A2(n56180), .Z(n49426) );
  XOR2_X1 U45900 ( .A1(n44759), .A2(n49426), .Z(n38880) );
  INV_X1 U45902 ( .I(n39363), .ZN(n30793) );
  XOR2_X1 U45903 ( .A1(n38880), .A2(n30793), .Z(n38146) );
  XOR2_X1 U45904 ( .A1(n44378), .A2(n53154), .Z(n50247) );
  XOR2_X1 U45905 ( .A1(n46683), .A2(n50247), .Z(n39243) );
  XOR2_X1 U45906 ( .A1(n54556), .A2(n58084), .Z(n30794) );
  XOR2_X1 U45907 ( .A1(n39243), .A2(n30794), .Z(n30795) );
  XOR2_X1 U45908 ( .A1(n30796), .A2(n30797), .Z(n30798) );
  NOR3_X1 U45911 ( .A1(n30804), .A2(n162), .A3(n30803), .ZN(n30805) );
  MUX2_X1 U45912 ( .I0(n30806), .I1(n30805), .S(n10820), .Z(n30827) );
  XOR2_X1 U45915 ( .A1(n9609), .A2(n33839), .Z(n30829) );
  XOR2_X1 U45916 ( .A1(n31925), .A2(n14665), .Z(n30835) );
  XOR2_X1 U45917 ( .A1(n15714), .A2(n55034), .Z(n30834) );
  INV_X1 U45919 ( .I(n32574), .ZN(n30836) );
  INV_X1 U45920 ( .I(n30839), .ZN(n30842) );
  XOR2_X1 U45922 ( .A1(n53713), .A2(n52226), .Z(n38896) );
  INV_X1 U45923 ( .I(n38896), .ZN(n30849) );
  XOR2_X1 U45924 ( .A1(n238), .A2(n30849), .Z(n30947) );
  XOR2_X1 U45925 ( .A1(n30947), .A2(n56143), .Z(n38996) );
  XOR2_X1 U45926 ( .A1(n56905), .A2(n53246), .Z(n39530) );
  XOR2_X1 U45927 ( .A1(n38826), .A2(n39530), .Z(n38651) );
  XOR2_X1 U45928 ( .A1(n60799), .A2(n55335), .Z(n30850) );
  XOR2_X1 U45929 ( .A1(n38996), .A2(n30850), .Z(n46301) );
  XOR2_X1 U45930 ( .A1(n54126), .A2(n24014), .Z(n33166) );
  XOR2_X1 U45931 ( .A1(n33166), .A2(n63603), .Z(n50763) );
  XOR2_X1 U45932 ( .A1(n53641), .A2(n56008), .Z(n31510) );
  XOR2_X1 U45933 ( .A1(n50763), .A2(n31510), .Z(n44831) );
  XOR2_X1 U45934 ( .A1(n46301), .A2(n44831), .Z(n30851) );
  XOR2_X1 U45935 ( .A1(n63955), .A2(n30851), .Z(n30852) );
  XOR2_X1 U45936 ( .A1(n31924), .A2(n30852), .Z(n30853) );
  NAND2_X1 U45937 ( .A1(n30854), .A2(n13444), .ZN(n30855) );
  NOR2_X1 U45938 ( .A1(n30856), .A2(n30855), .ZN(n30861) );
  NAND2_X1 U45940 ( .A1(n25989), .A2(n31279), .ZN(n30874) );
  INV_X1 U45942 ( .I(n30875), .ZN(n30878) );
  INV_X1 U45945 ( .I(n30890), .ZN(n30892) );
  AOI21_X1 U45946 ( .A1(n31239), .A2(n30892), .B(n30891), .ZN(n30893) );
  XOR2_X1 U45947 ( .A1(n17463), .A2(n15725), .Z(n31452) );
  XOR2_X1 U45948 ( .A1(n54776), .A2(n54936), .Z(n51814) );
  XOR2_X1 U45949 ( .A1(n50475), .A2(n24061), .Z(n36998) );
  XOR2_X1 U45950 ( .A1(n37737), .A2(n36998), .Z(n39280) );
  XOR2_X1 U45951 ( .A1(n39280), .A2(n38450), .Z(n38378) );
  XOR2_X1 U45952 ( .A1(n38378), .A2(n22252), .Z(n50618) );
  XOR2_X1 U45953 ( .A1(n45371), .A2(n23455), .Z(n46371) );
  XOR2_X1 U45954 ( .A1(n46371), .A2(n50067), .Z(n30899) );
  XOR2_X1 U45955 ( .A1(n50618), .A2(n30899), .Z(n30900) );
  XOR2_X1 U45956 ( .A1(n32181), .A2(n30900), .Z(n30901) );
  XOR2_X1 U45959 ( .A1(n33068), .A2(n433), .Z(n30903) );
  XOR2_X1 U45961 ( .A1(n32710), .A2(n22390), .Z(n30906) );
  XOR2_X1 U45962 ( .A1(n22950), .A2(n55060), .Z(n38000) );
  XOR2_X1 U45963 ( .A1(n9826), .A2(n38000), .Z(n36318) );
  XOR2_X1 U45964 ( .A1(n38962), .A2(n24011), .Z(n30909) );
  XOR2_X1 U45965 ( .A1(n36318), .A2(n30909), .Z(n44489) );
  XNOR2_X1 U45966 ( .A1(n55876), .A2(n53076), .ZN(n30910) );
  XOR2_X1 U45967 ( .A1(n30910), .A2(n32344), .Z(n45349) );
  XOR2_X1 U45968 ( .A1(n44489), .A2(n45349), .Z(n30911) );
  XOR2_X1 U45969 ( .A1(n38407), .A2(n54536), .Z(n45348) );
  XOR2_X1 U45970 ( .A1(n17758), .A2(n45348), .Z(n33053) );
  XOR2_X1 U45971 ( .A1(n50533), .A2(n54376), .Z(n50969) );
  XOR2_X1 U45972 ( .A1(n29407), .A2(n22821), .Z(n30914) );
  XOR2_X1 U45973 ( .A1(n45064), .A2(n30914), .Z(n30915) );
  XOR2_X1 U45974 ( .A1(n50969), .A2(n30915), .Z(n30916) );
  XOR2_X1 U45975 ( .A1(n23989), .A2(n23306), .Z(n32728) );
  XOR2_X1 U45976 ( .A1(n30036), .A2(n32728), .Z(n45131) );
  XOR2_X1 U45977 ( .A1(n30916), .A2(n45131), .Z(n30917) );
  XOR2_X1 U45978 ( .A1(n32470), .A2(n30917), .Z(n30918) );
  XOR2_X1 U45979 ( .A1(n10057), .A2(n44602), .Z(n33043) );
  INV_X1 U45980 ( .I(n33043), .ZN(n30919) );
  XOR2_X1 U45981 ( .A1(n30920), .A2(n30919), .Z(n30922) );
  XOR2_X1 U45982 ( .A1(n23714), .A2(n32267), .Z(n30930) );
  XOR2_X1 U45983 ( .A1(n39228), .A2(n56949), .Z(n32263) );
  XOR2_X1 U45984 ( .A1(n32263), .A2(n24109), .Z(n51278) );
  XOR2_X1 U45985 ( .A1(n57989), .A2(n54917), .Z(n43857) );
  XOR2_X1 U45986 ( .A1(n43857), .A2(n55638), .Z(n30924) );
  XOR2_X1 U45987 ( .A1(n30924), .A2(n43858), .Z(n30925) );
  XOR2_X1 U45988 ( .A1(n51278), .A2(n30925), .Z(n30927) );
  XOR2_X1 U45989 ( .A1(n56879), .A2(n56335), .Z(n30926) );
  BUF_X2 U45990 ( .I(n30926), .Z(n52178) );
  XOR2_X1 U45991 ( .A1(n39434), .A2(n52178), .Z(n32519) );
  XOR2_X1 U45992 ( .A1(n32519), .A2(n9871), .Z(n43864) );
  XOR2_X1 U45993 ( .A1(n30927), .A2(n43864), .Z(n30928) );
  XOR2_X1 U45994 ( .A1(n32170), .A2(n30928), .Z(n30929) );
  XOR2_X1 U45995 ( .A1(n30930), .A2(n30929), .Z(n30931) );
  XOR2_X1 U45996 ( .A1(n24051), .A2(n54249), .Z(n50504) );
  XOR2_X1 U45997 ( .A1(n50504), .A2(n44378), .Z(n45274) );
  XNOR2_X1 U45998 ( .A1(n23886), .A2(n56702), .ZN(n30937) );
  XOR2_X1 U45999 ( .A1(n30937), .A2(n22323), .Z(n30938) );
  XOR2_X1 U46000 ( .A1(n22961), .A2(n30938), .Z(n30939) );
  XOR2_X1 U46001 ( .A1(n46683), .A2(n30939), .Z(n30940) );
  XOR2_X1 U46002 ( .A1(n27640), .A2(n54734), .Z(n44109) );
  XOR2_X1 U46003 ( .A1(n52734), .A2(n4561), .Z(n39538) );
  XOR2_X1 U46004 ( .A1(n44109), .A2(n39538), .Z(n46245) );
  XOR2_X1 U46005 ( .A1(n30940), .A2(n46245), .Z(n30941) );
  XOR2_X1 U46006 ( .A1(n33857), .A2(n30946), .Z(n30951) );
  INV_X1 U46007 ( .I(n30947), .ZN(n38441) );
  XOR2_X1 U46009 ( .A1(n38388), .A2(n51494), .Z(n38277) );
  XOR2_X1 U46010 ( .A1(n60207), .A2(n39530), .Z(n30948) );
  XOR2_X1 U46011 ( .A1(n38441), .A2(n30948), .Z(n44241) );
  XOR2_X1 U46012 ( .A1(n37952), .A2(n37468), .Z(n43936) );
  XOR2_X1 U46013 ( .A1(n44241), .A2(n43936), .Z(n30949) );
  OAI21_X1 U46014 ( .A1(n17414), .A2(n18736), .B(n30952), .ZN(n30955) );
  INV_X1 U46015 ( .I(n32917), .ZN(n30962) );
  NAND2_X1 U46016 ( .A1(n33509), .A2(n21041), .ZN(n30961) );
  AOI21_X1 U46017 ( .A1(n30962), .A2(n30961), .B(n32919), .ZN(n30963) );
  INV_X1 U46018 ( .I(n34540), .ZN(n30965) );
  NOR2_X1 U46019 ( .A1(n30965), .A2(n33506), .ZN(n30967) );
  XOR2_X1 U46021 ( .A1(n37981), .A2(n53945), .Z(n44163) );
  INV_X1 U46022 ( .I(n44163), .ZN(n30972) );
  XOR2_X1 U46023 ( .A1(n39631), .A2(n38639), .Z(n30968) );
  XOR2_X1 U46024 ( .A1(n52513), .A2(n29407), .Z(n43687) );
  XOR2_X1 U46025 ( .A1(n7264), .A2(n43687), .Z(n30970) );
  XOR2_X1 U46026 ( .A1(n37651), .A2(n53787), .Z(n51608) );
  XOR2_X1 U46027 ( .A1(n51608), .A2(n53064), .Z(n30969) );
  XOR2_X1 U46028 ( .A1(n30970), .A2(n30969), .Z(n30971) );
  XOR2_X1 U46029 ( .A1(n887), .A2(n31464), .Z(n30975) );
  XOR2_X1 U46030 ( .A1(n30980), .A2(n53989), .Z(n39549) );
  XOR2_X1 U46031 ( .A1(n39549), .A2(n56508), .Z(n46142) );
  XOR2_X1 U46032 ( .A1(n31230), .A2(n54185), .Z(n51841) );
  XOR2_X1 U46033 ( .A1(n53685), .A2(n57989), .Z(n31398) );
  XOR2_X1 U46034 ( .A1(n51841), .A2(n31398), .Z(n44971) );
  XOR2_X1 U46035 ( .A1(n44971), .A2(n55087), .Z(n30981) );
  XOR2_X1 U46036 ( .A1(n19627), .A2(n30981), .Z(n30982) );
  XOR2_X1 U46037 ( .A1(n46142), .A2(n30982), .Z(n30984) );
  XOR2_X1 U46038 ( .A1(n23791), .A2(n60372), .Z(n30983) );
  XOR2_X1 U46039 ( .A1(n30984), .A2(n30983), .Z(n30988) );
  XOR2_X1 U46040 ( .A1(n30986), .A2(n15733), .Z(n31497) );
  XOR2_X1 U46041 ( .A1(n39469), .A2(n23886), .Z(n46398) );
  XOR2_X1 U46042 ( .A1(n44841), .A2(n39360), .Z(n45819) );
  XOR2_X1 U46043 ( .A1(n45819), .A2(n53344), .Z(n52141) );
  XOR2_X1 U46044 ( .A1(n57131), .A2(n53090), .Z(n43968) );
  XOR2_X1 U46045 ( .A1(n49426), .A2(n43968), .Z(n46397) );
  XOR2_X1 U46046 ( .A1(n52141), .A2(n46397), .Z(n30989) );
  XOR2_X1 U46048 ( .A1(n24014), .A2(n56827), .Z(n39196) );
  XOR2_X1 U46050 ( .A1(n39707), .A2(n38653), .Z(n31622) );
  XOR2_X1 U46051 ( .A1(n37468), .A2(n52970), .Z(n38997) );
  XOR2_X1 U46052 ( .A1(n31622), .A2(n38997), .Z(n44999) );
  XOR2_X1 U46053 ( .A1(n44999), .A2(n23926), .Z(n51002) );
  XOR2_X1 U46054 ( .A1(n37303), .A2(n53713), .Z(n38562) );
  XOR2_X1 U46055 ( .A1(n24044), .A2(n55840), .Z(n31388) );
  XOR2_X1 U46056 ( .A1(n31388), .A2(n56143), .Z(n38898) );
  XOR2_X1 U46057 ( .A1(n38562), .A2(n38898), .Z(n46168) );
  XOR2_X1 U46058 ( .A1(n46168), .A2(n44995), .Z(n30995) );
  XOR2_X1 U46059 ( .A1(n51002), .A2(n30995), .Z(n30996) );
  XOR2_X1 U46061 ( .A1(n30999), .A2(n30998), .Z(n31001) );
  XOR2_X1 U46062 ( .A1(n20862), .A2(n56008), .Z(n32239) );
  XOR2_X1 U46063 ( .A1(n32239), .A2(n23826), .Z(n31000) );
  XOR2_X1 U46064 ( .A1(n31001), .A2(n31000), .Z(n31002) );
  XOR2_X1 U46065 ( .A1(n31003), .A2(n31002), .Z(n31026) );
  INV_X1 U46066 ( .I(n34046), .ZN(n31022) );
  XOR2_X1 U46067 ( .A1(n38154), .A2(n53487), .Z(n32397) );
  XOR2_X1 U46068 ( .A1(n56692), .A2(n55610), .Z(n45101) );
  XOR2_X1 U46069 ( .A1(n32397), .A2(n45101), .Z(n31005) );
  XOR2_X1 U46070 ( .A1(n53076), .A2(n56771), .Z(n32123) );
  XOR2_X1 U46071 ( .A1(n32123), .A2(n32344), .Z(n52399) );
  XOR2_X1 U46072 ( .A1(n31005), .A2(n52399), .Z(n43901) );
  XOR2_X1 U46073 ( .A1(n24011), .A2(n54153), .Z(n37565) );
  XOR2_X1 U46074 ( .A1(n37565), .A2(n54386), .Z(n44264) );
  XOR2_X1 U46075 ( .A1(n22950), .A2(n53805), .Z(n31006) );
  XOR2_X1 U46076 ( .A1(n44264), .A2(n31006), .Z(n31007) );
  XOR2_X1 U46077 ( .A1(n43901), .A2(n31007), .Z(n31008) );
  XOR2_X1 U46078 ( .A1(n31009), .A2(n33144), .Z(n31012) );
  XOR2_X1 U46079 ( .A1(n60525), .A2(n22244), .Z(n31010) );
  XOR2_X1 U46080 ( .A1(n54776), .A2(n54208), .Z(n39457) );
  XOR2_X1 U46081 ( .A1(n38009), .A2(n39457), .Z(n31634) );
  XOR2_X1 U46082 ( .A1(n50067), .A2(n55903), .Z(n33886) );
  XOR2_X1 U46083 ( .A1(n56124), .A2(n52232), .Z(n31014) );
  XOR2_X1 U46084 ( .A1(n44533), .A2(n31014), .Z(n31015) );
  XOR2_X1 U46085 ( .A1(n33886), .A2(n31015), .Z(n31016) );
  XOR2_X1 U46086 ( .A1(n31634), .A2(n31016), .Z(n45250) );
  XOR2_X1 U46087 ( .A1(n58928), .A2(n36998), .Z(n44138) );
  XOR2_X1 U46088 ( .A1(n45250), .A2(n44138), .Z(n31017) );
  INV_X1 U46089 ( .I(n33141), .ZN(n32498) );
  XOR2_X1 U46090 ( .A1(n31809), .A2(n32498), .Z(n33272) );
  XOR2_X1 U46091 ( .A1(n33272), .A2(n31019), .Z(n31020) );
  NAND2_X1 U46093 ( .A1(n23746), .A2(n19610), .ZN(n33422) );
  NOR2_X1 U46094 ( .A1(n33422), .A2(n34039), .ZN(n34616) );
  INV_X1 U46096 ( .I(n31029), .ZN(n31030) );
  NOR2_X1 U46097 ( .A1(n31040), .A2(n31039), .ZN(n31043) );
  INV_X1 U46099 ( .I(n20918), .ZN(n31050) );
  INV_X1 U46100 ( .I(n31053), .ZN(n31057) );
  OAI21_X1 U46101 ( .A1(n31059), .A2(n17627), .B(n31054), .ZN(n31056) );
  NOR2_X1 U46102 ( .A1(n31061), .A2(n31060), .ZN(n31062) );
  XOR2_X1 U46103 ( .A1(n55106), .A2(n23455), .Z(n46112) );
  XOR2_X1 U46104 ( .A1(n46112), .A2(n50067), .Z(n31066) );
  XOR2_X1 U46105 ( .A1(n55603), .A2(n56124), .Z(n31065) );
  BUF_X2 U46106 ( .I(n31065), .Z(n51193) );
  XOR2_X1 U46107 ( .A1(n31066), .A2(n51193), .Z(n44925) );
  XOR2_X1 U46110 ( .A1(n61550), .A2(n53375), .Z(n39210) );
  XOR2_X1 U46112 ( .A1(n23968), .A2(n24061), .Z(n32621) );
  XOR2_X1 U46113 ( .A1(n32621), .A2(n31068), .Z(n38007) );
  XOR2_X1 U46114 ( .A1(n50790), .A2(n38007), .Z(n45337) );
  XOR2_X1 U46115 ( .A1(n32274), .A2(n55903), .Z(n44534) );
  XOR2_X1 U46116 ( .A1(n44534), .A2(n54208), .Z(n31069) );
  XOR2_X1 U46117 ( .A1(n45337), .A2(n31069), .Z(n31071) );
  XOR2_X1 U46118 ( .A1(n31071), .A2(n31070), .Z(n31072) );
  OAI21_X1 U46119 ( .A1(n31088), .A2(n24504), .B(n23708), .ZN(n31091) );
  INV_X1 U46120 ( .I(n31089), .ZN(n31090) );
  NAND2_X1 U46121 ( .A1(n31093), .A2(n31092), .ZN(n31096) );
  NOR2_X1 U46122 ( .A1(n10427), .A2(n31098), .ZN(n31100) );
  NOR2_X1 U46123 ( .A1(n31098), .A2(n19590), .ZN(n31099) );
  XOR2_X1 U46124 ( .A1(n53262), .A2(n56915), .Z(n44014) );
  XOR2_X1 U46125 ( .A1(n44014), .A2(n32344), .Z(n32546) );
  XOR2_X1 U46126 ( .A1(n32546), .A2(n55876), .Z(n39665) );
  XOR2_X1 U46127 ( .A1(n51999), .A2(n50831), .Z(n38829) );
  XOR2_X1 U46128 ( .A1(n39665), .A2(n38829), .Z(n43730) );
  XOR2_X1 U46129 ( .A1(n54716), .A2(n56859), .Z(n45238) );
  XOR2_X1 U46130 ( .A1(n38733), .A2(n45238), .Z(n39773) );
  XOR2_X1 U46131 ( .A1(n39773), .A2(n54153), .Z(n44357) );
  XOR2_X1 U46132 ( .A1(n51021), .A2(n55546), .Z(n31106) );
  XOR2_X1 U46133 ( .A1(n44357), .A2(n31106), .Z(n31107) );
  XOR2_X1 U46134 ( .A1(n43730), .A2(n31107), .Z(n31108) );
  XOR2_X1 U46135 ( .A1(n23768), .A2(n31108), .Z(n31109) );
  OAI21_X1 U46136 ( .A1(n14276), .A2(n161), .B(n31111), .ZN(n31112) );
  INV_X1 U46137 ( .I(n31115), .ZN(n31116) );
  XOR2_X1 U46138 ( .A1(n38826), .A2(n56143), .Z(n50832) );
  NAND2_X1 U46140 ( .A1(n31125), .A2(n31124), .ZN(n31126) );
  NAND2_X1 U46141 ( .A1(n31132), .A2(n31131), .ZN(n31630) );
  XOR2_X1 U46142 ( .A1(n54676), .A2(n57096), .Z(n32410) );
  XOR2_X1 U46143 ( .A1(n54126), .A2(n53318), .Z(n39706) );
  XOR2_X1 U46144 ( .A1(n32410), .A2(n39706), .Z(n38280) );
  XOR2_X1 U46145 ( .A1(n38280), .A2(n63603), .Z(n44914) );
  XOR2_X1 U46146 ( .A1(n37584), .A2(n24014), .Z(n32172) );
  XOR2_X1 U46147 ( .A1(n44914), .A2(n32172), .Z(n50720) );
  XOR2_X1 U46148 ( .A1(n53713), .A2(n51881), .Z(n31133) );
  XOR2_X1 U46149 ( .A1(n39478), .A2(n31133), .Z(n46192) );
  XOR2_X1 U46150 ( .A1(n50720), .A2(n46192), .Z(n31134) );
  XOR2_X1 U46151 ( .A1(n23090), .A2(n31134), .Z(n31135) );
  INV_X1 U46152 ( .I(n31136), .ZN(n31151) );
  AOI22_X1 U46154 ( .A1(n31142), .A2(n31141), .B1(n31140), .B2(n31139), .ZN(
        n31150) );
  XOR2_X1 U46155 ( .A1(n31153), .A2(n31152), .Z(n31154) );
  NAND2_X1 U46158 ( .A1(n31269), .A2(n31277), .ZN(n31164) );
  OAI22_X1 U46159 ( .A1(n31278), .A2(n31167), .B1(n31166), .B2(n31165), .ZN(
        n31168) );
  NAND2_X1 U46160 ( .A1(n12125), .A2(n6316), .ZN(n31171) );
  NAND2_X1 U46162 ( .A1(n31173), .A2(n13444), .ZN(n31176) );
  NAND2_X1 U46163 ( .A1(n31174), .A2(n17590), .ZN(n31175) );
  MUX2_X1 U46164 ( .I0(n31176), .I1(n31175), .S(n31182), .Z(n31574) );
  INV_X1 U46165 ( .I(n31177), .ZN(n31179) );
  NAND2_X1 U46166 ( .A1(n31187), .A2(n17590), .ZN(n31178) );
  NOR2_X1 U46167 ( .A1(n13444), .A2(n31178), .ZN(n31569) );
  AOI21_X1 U46168 ( .A1(n31179), .A2(n1866), .B(n31569), .ZN(n31192) );
  OAI21_X1 U46169 ( .A1(n31182), .A2(n24556), .B(n57845), .ZN(n31185) );
  NOR2_X1 U46170 ( .A1(n1866), .A2(n1353), .ZN(n31183) );
  NOR2_X1 U46171 ( .A1(n62152), .A2(n63256), .ZN(n31188) );
  OAI21_X1 U46172 ( .A1(n1353), .A2(n24777), .B(n31188), .ZN(n31190) );
  NAND2_X1 U46173 ( .A1(n31191), .A2(n31190), .ZN(n31573) );
  NAND4_X1 U46174 ( .A1(n31574), .A2(n31192), .A3(n31572), .A4(n31573), .ZN(
        n31194) );
  XOR2_X1 U46175 ( .A1(n24103), .A2(n18596), .Z(n32648) );
  XOR2_X1 U46176 ( .A1(n54888), .A2(n54219), .Z(n32472) );
  XOR2_X1 U46177 ( .A1(n32472), .A2(n15707), .Z(n51667) );
  XOR2_X1 U46178 ( .A1(n51667), .A2(n53787), .Z(n37692) );
  XOR2_X1 U46180 ( .A1(n53945), .A2(n55340), .Z(n50025) );
  INV_X1 U46181 ( .I(n50025), .ZN(n31195) );
  XOR2_X1 U46182 ( .A1(n31195), .A2(n30036), .Z(n31311) );
  XOR2_X1 U46184 ( .A1(n38639), .A2(n620), .Z(n39558) );
  XOR2_X1 U46185 ( .A1(n38459), .A2(n39558), .Z(n31196) );
  XOR2_X1 U46186 ( .A1(n37692), .A2(n31196), .Z(n44546) );
  XOR2_X1 U46187 ( .A1(n52080), .A2(n37651), .Z(n38065) );
  XOR2_X1 U46188 ( .A1(n38065), .A2(n60797), .Z(n45322) );
  XOR2_X1 U46189 ( .A1(n45322), .A2(n22821), .Z(n31197) );
  XOR2_X1 U46190 ( .A1(n44546), .A2(n31197), .Z(n31198) );
  OAI21_X1 U46191 ( .A1(n31203), .A2(n31202), .B(n31201), .ZN(n31207) );
  NAND3_X1 U46192 ( .A1(n20378), .A2(n31204), .A3(n31208), .ZN(n31205) );
  NAND3_X1 U46193 ( .A1(n31207), .A2(n31206), .A3(n31205), .ZN(n31213) );
  NAND2_X1 U46194 ( .A1(n1847), .A2(n31208), .ZN(n31210) );
  AOI21_X1 U46195 ( .A1(n31211), .A2(n31210), .B(n31209), .ZN(n31212) );
  NAND2_X1 U46196 ( .A1(n62892), .A2(n31214), .ZN(n31219) );
  NOR2_X1 U46197 ( .A1(n1875), .A2(n31224), .ZN(n31225) );
  XOR2_X1 U46198 ( .A1(n23929), .A2(n53989), .Z(n31226) );
  BUF_X2 U46199 ( .I(n31226), .Z(n50551) );
  XOR2_X1 U46200 ( .A1(n55889), .A2(n56508), .Z(n38772) );
  XOR2_X1 U46201 ( .A1(n50551), .A2(n38772), .Z(n50650) );
  INV_X1 U46202 ( .I(n39228), .ZN(n50984) );
  XOR2_X1 U46203 ( .A1(n247), .A2(n50984), .Z(n31877) );
  INV_X1 U46204 ( .I(n31877), .ZN(n31227) );
  XOR2_X1 U46205 ( .A1(n24109), .A2(n59130), .Z(n44796) );
  XOR2_X1 U46206 ( .A1(n44796), .A2(n51530), .Z(n32658) );
  XOR2_X1 U46207 ( .A1(n32658), .A2(n31227), .Z(n46204) );
  XOR2_X1 U46208 ( .A1(n56714), .A2(n51946), .Z(n31228) );
  XOR2_X1 U46209 ( .A1(n50943), .A2(n31228), .Z(n31229) );
  XOR2_X1 U46210 ( .A1(n31230), .A2(n31229), .Z(n42711) );
  XOR2_X1 U46211 ( .A1(n42711), .A2(n55638), .Z(n31231) );
  XOR2_X1 U46212 ( .A1(n46204), .A2(n31231), .Z(n31232) );
  XOR2_X1 U46213 ( .A1(n23042), .A2(n31232), .Z(n31233) );
  NAND4_X1 U46215 ( .A1(n34639), .A2(n61452), .A3(n61449), .A4(n34632), .ZN(
        n31237) );
  NOR2_X1 U46216 ( .A1(n31241), .A2(n31240), .ZN(n31244) );
  NAND3_X1 U46218 ( .A1(n31250), .A2(n31249), .A3(n31248), .ZN(n31251) );
  INV_X1 U46219 ( .I(n31253), .ZN(n31258) );
  NAND2_X1 U46223 ( .A1(n31280), .A2(n31279), .ZN(n31286) );
  XOR2_X1 U46227 ( .A1(n24046), .A2(n55792), .Z(n50505) );
  INV_X1 U46229 ( .I(n22323), .ZN(n52448) );
  XOR2_X1 U46230 ( .A1(n38400), .A2(n52448), .Z(n50733) );
  XOR2_X1 U46231 ( .A1(n50733), .A2(n54556), .Z(n40459) );
  XOR2_X1 U46232 ( .A1(n42790), .A2(n27640), .Z(n44983) );
  XOR2_X1 U46233 ( .A1(n49426), .A2(n53272), .Z(n46601) );
  XOR2_X1 U46234 ( .A1(n44983), .A2(n46601), .Z(n31291) );
  XOR2_X1 U46235 ( .A1(n40459), .A2(n31291), .Z(n31292) );
  INV_X1 U46237 ( .I(n23774), .ZN(n31297) );
  NOR2_X1 U46238 ( .A1(n31298), .A2(n34643), .ZN(n31299) );
  NAND2_X1 U46239 ( .A1(n60984), .A2(n34634), .ZN(n31301) );
  OAI22_X1 U46240 ( .A1(n31301), .A2(n34641), .B1(n34643), .B2(n35032), .ZN(
        n31302) );
  NAND2_X2 U46241 ( .A1(n35994), .A2(n37046), .ZN(n37051) );
  INV_X1 U46243 ( .I(n35480), .ZN(n31307) );
  NAND2_X1 U46244 ( .A1(n35997), .A2(n37050), .ZN(n31308) );
  XOR2_X1 U46245 ( .A1(n50817), .A2(n24067), .Z(n38721) );
  XOR2_X1 U46246 ( .A1(n55534), .A2(n55191), .Z(n39334) );
  XOR2_X1 U46247 ( .A1(n38721), .A2(n39334), .Z(n38947) );
  XOR2_X1 U46248 ( .A1(n37651), .A2(n55052), .Z(n31679) );
  XOR2_X1 U46249 ( .A1(n38947), .A2(n31679), .Z(n43193) );
  XOR2_X1 U46250 ( .A1(n43193), .A2(n60556), .Z(n31312) );
  XOR2_X1 U46251 ( .A1(n51611), .A2(n22821), .Z(n31310) );
  XOR2_X1 U46252 ( .A1(n31312), .A2(n44094), .Z(n31313) );
  XOR2_X1 U46253 ( .A1(n65041), .A2(n31313), .Z(n31314) );
  XOR2_X1 U46254 ( .A1(n53359), .A2(n65079), .Z(n44613) );
  XOR2_X1 U46255 ( .A1(n50650), .A2(n37637), .Z(n33899) );
  XOR2_X1 U46256 ( .A1(n31318), .A2(n33899), .Z(n31642) );
  INV_X1 U46257 ( .I(n31642), .ZN(n31320) );
  XOR2_X1 U46258 ( .A1(n55638), .A2(n54917), .Z(n31319) );
  XOR2_X1 U46259 ( .A1(n31320), .A2(n31319), .Z(n46631) );
  XOR2_X1 U46260 ( .A1(n53685), .A2(n53174), .Z(n51216) );
  XOR2_X1 U46261 ( .A1(n51216), .A2(n55580), .Z(n36860) );
  XOR2_X1 U46262 ( .A1(n36860), .A2(n39434), .Z(n44415) );
  XOR2_X1 U46263 ( .A1(n46631), .A2(n44415), .Z(n31321) );
  INV_X1 U46264 ( .I(n31384), .ZN(n31324) );
  XOR2_X1 U46265 ( .A1(n49426), .A2(n53499), .Z(n52096) );
  XOR2_X1 U46266 ( .A1(n22773), .A2(n55624), .Z(n39723) );
  XOR2_X1 U46267 ( .A1(n39723), .A2(n39611), .Z(n31325) );
  XOR2_X1 U46268 ( .A1(n52096), .A2(n31325), .Z(n45405) );
  XOR2_X1 U46269 ( .A1(n45405), .A2(n52135), .Z(n31326) );
  XOR2_X1 U46271 ( .A1(n23754), .A2(n55792), .Z(n44467) );
  XOR2_X1 U46272 ( .A1(n23869), .A2(n23090), .Z(n31329) );
  XOR2_X1 U46273 ( .A1(n55335), .A2(n53246), .Z(n46615) );
  XOR2_X1 U46274 ( .A1(n32669), .A2(n46615), .Z(n31858) );
  XOR2_X1 U46275 ( .A1(n39707), .A2(n23851), .Z(n32087) );
  XOR2_X1 U46276 ( .A1(n32087), .A2(n38653), .Z(n38893) );
  XOR2_X1 U46277 ( .A1(n44995), .A2(n53318), .Z(n50999) );
  XOR2_X1 U46278 ( .A1(n50999), .A2(n37468), .Z(n31330) );
  XOR2_X1 U46279 ( .A1(n38893), .A2(n31330), .Z(n44446) );
  XOR2_X1 U46280 ( .A1(n23926), .A2(n52900), .Z(n33165) );
  XOR2_X1 U46281 ( .A1(n33165), .A2(n38896), .Z(n39373) );
  XOR2_X1 U46282 ( .A1(n39373), .A2(n51881), .Z(n46617) );
  XOR2_X1 U46283 ( .A1(n44446), .A2(n46617), .Z(n31331) );
  XOR2_X1 U46284 ( .A1(n727), .A2(n15725), .Z(n31333) );
  XOR2_X1 U46285 ( .A1(n26920), .A2(n60565), .Z(n31334) );
  XOR2_X1 U46287 ( .A1(n51193), .A2(n50067), .Z(n37710) );
  XOR2_X1 U46288 ( .A1(n31634), .A2(n37710), .Z(n43497) );
  XOR2_X1 U46289 ( .A1(n37737), .A2(n55655), .Z(n37897) );
  XNOR2_X1 U46290 ( .A1(n23968), .A2(n23999), .ZN(n31338) );
  XOR2_X1 U46291 ( .A1(n37897), .A2(n31339), .Z(n44078) );
  XOR2_X1 U46292 ( .A1(n43497), .A2(n44078), .Z(n31340) );
  XOR2_X1 U46295 ( .A1(n32123), .A2(n56165), .Z(n37512) );
  XOR2_X1 U46296 ( .A1(n37512), .A2(n32344), .Z(n38408) );
  XOR2_X1 U46297 ( .A1(n38408), .A2(n55876), .Z(n44812) );
  XOR2_X1 U46298 ( .A1(n55777), .A2(n56040), .Z(n37704) );
  INV_X1 U46299 ( .I(n31593), .ZN(n37889) );
  XOR2_X1 U46300 ( .A1(n37704), .A2(n37889), .Z(n38226) );
  XOR2_X1 U46301 ( .A1(n38226), .A2(n54716), .Z(n46284) );
  XOR2_X1 U46302 ( .A1(n50831), .A2(n53487), .Z(n37767) );
  XOR2_X1 U46303 ( .A1(n31347), .A2(n37767), .Z(n45026) );
  INV_X1 U46304 ( .I(n45026), .ZN(n50878) );
  XOR2_X1 U46305 ( .A1(n46284), .A2(n50878), .Z(n31348) );
  XOR2_X1 U46306 ( .A1(n44812), .A2(n31348), .Z(n31349) );
  XOR2_X1 U46307 ( .A1(n60525), .A2(n31349), .Z(n31350) );
  XOR2_X1 U46308 ( .A1(n31350), .A2(n33144), .Z(n31351) );
  NAND2_X2 U46309 ( .A1(n15786), .A2(n25251), .ZN(n34666) );
  OAI21_X1 U46310 ( .A1(n34518), .A2(n33454), .B(n34667), .ZN(n31359) );
  XOR2_X1 U46311 ( .A1(n31360), .A2(n61550), .Z(n43772) );
  XOR2_X1 U46312 ( .A1(n31746), .A2(n1190), .Z(n44024) );
  XOR2_X1 U46313 ( .A1(n44024), .A2(n50697), .Z(n31361) );
  XOR2_X1 U46314 ( .A1(n43772), .A2(n31361), .Z(n31362) );
  XOR2_X1 U46315 ( .A1(n32543), .A2(n53530), .Z(n31440) );
  XOR2_X1 U46316 ( .A1(n32540), .A2(n50475), .Z(n31366) );
  INV_X1 U46317 ( .I(n15735), .ZN(n51029) );
  XOR2_X1 U46318 ( .A1(n24017), .A2(n51029), .Z(n31367) );
  XOR2_X1 U46319 ( .A1(n22244), .A2(n32393), .Z(n31368) );
  XOR2_X1 U46320 ( .A1(n32546), .A2(n56475), .Z(n50777) );
  XOR2_X1 U46321 ( .A1(n38829), .A2(n29969), .Z(n39663) );
  XOR2_X1 U46322 ( .A1(n50777), .A2(n39663), .Z(n41739) );
  XOR2_X1 U46323 ( .A1(n38733), .A2(n24011), .Z(n31369) );
  XOR2_X1 U46324 ( .A1(n56040), .A2(n53805), .Z(n31370) );
  XOR2_X1 U46325 ( .A1(n32988), .A2(n31370), .Z(n44714) );
  XOR2_X1 U46326 ( .A1(n41739), .A2(n44714), .Z(n31371) );
  NOR2_X1 U46327 ( .A1(n31378), .A2(n31376), .ZN(n31373) );
  INV_X1 U46328 ( .I(n31377), .ZN(n31372) );
  XOR2_X1 U46329 ( .A1(n55624), .A2(n56180), .Z(n31374) );
  AOI21_X1 U46330 ( .A1(n31373), .A2(n31372), .B(n31374), .ZN(n31380) );
  INV_X1 U46331 ( .I(n31374), .ZN(n31375) );
  NOR4_X1 U46332 ( .A1(n31378), .A2(n31377), .A3(n31376), .A4(n31375), .ZN(
        n31379) );
  NOR2_X1 U46333 ( .A1(n31380), .A2(n31379), .ZN(n31382) );
  XOR2_X1 U46334 ( .A1(n15712), .A2(n53154), .Z(n49434) );
  XOR2_X1 U46335 ( .A1(n49434), .A2(n27640), .Z(n39183) );
  XOR2_X1 U46336 ( .A1(n38400), .A2(n37630), .Z(n44622) );
  XOR2_X1 U46337 ( .A1(n9040), .A2(n31517), .Z(n31383) );
  INV_X1 U46338 ( .I(n44914), .ZN(n31387) );
  XOR2_X1 U46339 ( .A1(n15710), .A2(n39375), .Z(n33851) );
  XOR2_X1 U46340 ( .A1(n33851), .A2(n53641), .Z(n46437) );
  XOR2_X1 U46341 ( .A1(n31387), .A2(n46437), .Z(n31390) );
  XOR2_X1 U46342 ( .A1(n38896), .A2(n23926), .Z(n51290) );
  XOR2_X1 U46343 ( .A1(n31388), .A2(n54517), .Z(n31389) );
  XOR2_X1 U46344 ( .A1(n51290), .A2(n31389), .Z(n46708) );
  XOR2_X1 U46345 ( .A1(n31390), .A2(n46708), .Z(n31391) );
  XOR2_X1 U46346 ( .A1(n23869), .A2(n31391), .Z(n31392) );
  XOR2_X1 U46347 ( .A1(n31392), .A2(n59521), .Z(n31393) );
  XOR2_X1 U46348 ( .A1(n32414), .A2(n1550), .Z(n31394) );
  XOR2_X1 U46350 ( .A1(n32658), .A2(n51261), .Z(n51656) );
  XOR2_X1 U46351 ( .A1(n31397), .A2(n51656), .Z(n34833) );
  XOR2_X1 U46352 ( .A1(n50551), .A2(n55889), .Z(n31491) );
  XOR2_X1 U46353 ( .A1(n34833), .A2(n31491), .Z(n46648) );
  XOR2_X1 U46354 ( .A1(n53833), .A2(n65079), .Z(n33901) );
  XOR2_X1 U46355 ( .A1(n31398), .A2(n33901), .Z(n51531) );
  XOR2_X1 U46356 ( .A1(n50943), .A2(n53359), .Z(n31399) );
  XOR2_X1 U46357 ( .A1(n51531), .A2(n31399), .Z(n44877) );
  XOR2_X1 U46358 ( .A1(n46648), .A2(n44877), .Z(n31401) );
  XOR2_X1 U46361 ( .A1(n33204), .A2(n32118), .Z(n31404) );
  XOR2_X1 U46362 ( .A1(n32267), .A2(n32590), .Z(n31406) );
  XOR2_X1 U46363 ( .A1(n31407), .A2(n31406), .Z(n31408) );
  XOR2_X1 U46365 ( .A1(n43687), .A2(n24067), .Z(n38064) );
  XOR2_X1 U46366 ( .A1(n38064), .A2(n55765), .Z(n50536) );
  XOR2_X1 U46367 ( .A1(n56683), .A2(n55191), .Z(n31755) );
  XOR2_X1 U46368 ( .A1(n50536), .A2(n31755), .Z(n43784) );
  XOR2_X1 U46369 ( .A1(n51667), .A2(n55340), .Z(n31409) );
  XOR2_X1 U46370 ( .A1(n38639), .A2(n51611), .Z(n37844) );
  XOR2_X1 U46371 ( .A1(n31409), .A2(n37844), .Z(n39760) );
  XOR2_X1 U46372 ( .A1(n30036), .A2(n53748), .Z(n31410) );
  XOR2_X1 U46373 ( .A1(n39760), .A2(n31410), .Z(n44032) );
  XOR2_X1 U46374 ( .A1(n43784), .A2(n44032), .Z(n31411) );
  XOR2_X1 U46375 ( .A1(n32640), .A2(n8329), .Z(n31412) );
  NOR2_X1 U46378 ( .A1(n15809), .A2(n23945), .ZN(n34598) );
  NAND3_X1 U46379 ( .A1(n31417), .A2(n34598), .A3(n118), .ZN(n31418) );
  XOR2_X1 U46380 ( .A1(n1881), .A2(n34834), .Z(n38302) );
  XOR2_X1 U46381 ( .A1(n39434), .A2(n53685), .Z(n38258) );
  XOR2_X1 U46382 ( .A1(n38302), .A2(n38258), .Z(n45061) );
  INV_X1 U46383 ( .I(n55638), .ZN(n31422) );
  XOR2_X1 U46384 ( .A1(n50551), .A2(n31422), .Z(n37636) );
  XOR2_X1 U46385 ( .A1(n37636), .A2(n55889), .Z(n50190) );
  XOR2_X1 U46386 ( .A1(n50190), .A2(n55087), .Z(n31423) );
  XOR2_X1 U46387 ( .A1(n45061), .A2(n31423), .Z(n31424) );
  XOR2_X1 U46388 ( .A1(n23791), .A2(n31424), .Z(n31426) );
  XOR2_X1 U46389 ( .A1(n31425), .A2(n1573), .Z(n31823) );
  XOR2_X1 U46390 ( .A1(n9753), .A2(n53090), .Z(n45360) );
  XOR2_X1 U46391 ( .A1(n23858), .A2(n56065), .Z(n50745) );
  XOR2_X1 U46392 ( .A1(n23754), .A2(n58084), .Z(n37868) );
  XOR2_X1 U46393 ( .A1(n50745), .A2(n37868), .Z(n52097) );
  XOR2_X1 U46394 ( .A1(n52097), .A2(n55792), .Z(n37577) );
  XOR2_X1 U46395 ( .A1(n45360), .A2(n37577), .Z(n31428) );
  XOR2_X1 U46396 ( .A1(n15712), .A2(n24057), .Z(n44526) );
  XOR2_X1 U46397 ( .A1(n38146), .A2(n44526), .Z(n31427) );
  XOR2_X1 U46398 ( .A1(n31428), .A2(n31427), .Z(n31429) );
  XOR2_X1 U46399 ( .A1(n38733), .A2(n50955), .Z(n46219) );
  XOR2_X1 U46400 ( .A1(n56165), .A2(n53958), .Z(n39570) );
  XOR2_X1 U46401 ( .A1(n39570), .A2(n22950), .Z(n31434) );
  XOR2_X1 U46402 ( .A1(n23767), .A2(n31434), .Z(n31435) );
  XOR2_X1 U46403 ( .A1(n37767), .A2(n55876), .Z(n43065) );
  XOR2_X1 U46404 ( .A1(n31435), .A2(n43065), .Z(n31436) );
  XOR2_X1 U46405 ( .A1(n37513), .A2(n53138), .Z(n32286) );
  XOR2_X1 U46406 ( .A1(n32286), .A2(n49787), .Z(n46220) );
  XOR2_X1 U46407 ( .A1(n31436), .A2(n46220), .Z(n31437) );
  XOR2_X1 U46408 ( .A1(n58928), .A2(n44290), .Z(n37736) );
  XOR2_X1 U46409 ( .A1(n52375), .A2(n56745), .Z(n37896) );
  XOR2_X1 U46410 ( .A1(n37896), .A2(n51193), .Z(n43963) );
  XOR2_X1 U46412 ( .A1(n60799), .A2(n32232), .Z(n37803) );
  XOR2_X1 U46413 ( .A1(n37803), .A2(n51290), .Z(n39622) );
  XOR2_X1 U46414 ( .A1(n39622), .A2(n55840), .Z(n46444) );
  XOR2_X1 U46415 ( .A1(n53318), .A2(n55516), .Z(n46443) );
  XOR2_X1 U46416 ( .A1(n46443), .A2(n23851), .Z(n31445) );
  XOR2_X1 U46417 ( .A1(n31445), .A2(n31444), .Z(n38438) );
  XOR2_X1 U46418 ( .A1(n38438), .A2(n63603), .Z(n45048) );
  XOR2_X1 U46419 ( .A1(n46444), .A2(n45048), .Z(n31447) );
  XOR2_X1 U46420 ( .A1(n31447), .A2(n31446), .Z(n31448) );
  XOR2_X1 U46421 ( .A1(n20862), .A2(n32085), .Z(n31449) );
  XOR2_X1 U46423 ( .A1(n31804), .A2(n31452), .Z(n31453) );
  XOR2_X1 U46424 ( .A1(n31455), .A2(n24831), .Z(n31719) );
  XOR2_X1 U46425 ( .A1(n24065), .A2(n55340), .Z(n51765) );
  XOR2_X1 U46426 ( .A1(n51765), .A2(n22821), .Z(n37730) );
  XOR2_X1 U46427 ( .A1(n60556), .A2(n52317), .Z(n39444) );
  XOR2_X1 U46428 ( .A1(n38639), .A2(n39444), .Z(n31458) );
  XOR2_X1 U46429 ( .A1(n37730), .A2(n31458), .Z(n44275) );
  XOR2_X1 U46430 ( .A1(n37651), .A2(n24067), .Z(n43882) );
  XOR2_X1 U46431 ( .A1(n44275), .A2(n43882), .Z(n31459) );
  XOR2_X1 U46432 ( .A1(n31459), .A2(n43880), .Z(n31460) );
  NOR2_X1 U46435 ( .A1(n34657), .A2(n34168), .ZN(n32887) );
  INV_X1 U46436 ( .I(n31674), .ZN(n31479) );
  XOR2_X1 U46437 ( .A1(n36998), .A2(n53308), .Z(n36357) );
  XOR2_X1 U46438 ( .A1(n51133), .A2(n36357), .Z(n44390) );
  XOR2_X1 U46439 ( .A1(n38165), .A2(n50067), .Z(n43721) );
  XOR2_X1 U46440 ( .A1(n55903), .A2(n55833), .Z(n50787) );
  XOR2_X1 U46441 ( .A1(n43721), .A2(n50787), .Z(n31477) );
  XOR2_X1 U46443 ( .A1(n56475), .A2(n54231), .Z(n51512) );
  XOR2_X1 U46444 ( .A1(n55777), .A2(n55546), .Z(n51128) );
  XOR2_X1 U46445 ( .A1(n37565), .A2(n51128), .Z(n31482) );
  XOR2_X1 U46446 ( .A1(n38153), .A2(n31482), .Z(n44087) );
  INV_X1 U46447 ( .I(n29969), .ZN(n31483) );
  XOR2_X1 U46448 ( .A1(n55126), .A2(n50831), .Z(n39488) );
  XOR2_X1 U46449 ( .A1(n31483), .A2(n39488), .Z(n32024) );
  INV_X1 U46450 ( .I(n32024), .ZN(n43330) );
  XOR2_X1 U46451 ( .A1(n43330), .A2(n30908), .Z(n31484) );
  XOR2_X1 U46452 ( .A1(n43864), .A2(n54185), .Z(n39649) );
  XOR2_X1 U46453 ( .A1(n39649), .A2(n38472), .Z(n45126) );
  INV_X1 U46456 ( .I(n23786), .ZN(n31489) );
  XOR2_X1 U46457 ( .A1(n51407), .A2(n54917), .Z(n38631) );
  XOR2_X1 U46458 ( .A1(n38631), .A2(n51261), .Z(n31492) );
  XOR2_X1 U46459 ( .A1(n31492), .A2(n31491), .Z(n46523) );
  XOR2_X1 U46460 ( .A1(n57989), .A2(n51946), .Z(n45121) );
  XOR2_X1 U46461 ( .A1(n46523), .A2(n45121), .Z(n31493) );
  XOR2_X1 U46462 ( .A1(n18314), .A2(n31493), .Z(n31495) );
  INV_X1 U46463 ( .I(n23042), .ZN(n31494) );
  XOR2_X1 U46464 ( .A1(n31495), .A2(n31494), .Z(n31496) );
  XOR2_X1 U46465 ( .A1(n31497), .A2(n31496), .Z(n31498) );
  XOR2_X1 U46467 ( .A1(n11930), .A2(n2259), .Z(n31503) );
  XOR2_X1 U46469 ( .A1(n42426), .A2(n53787), .Z(n37983) );
  XOR2_X1 U46470 ( .A1(n37983), .A2(n38065), .Z(n50666) );
  XOR2_X1 U46471 ( .A1(n39263), .A2(n51569), .Z(n44350) );
  XNOR2_X1 U46472 ( .A1(n60556), .A2(n55340), .ZN(n31504) );
  XOR2_X1 U46473 ( .A1(n43687), .A2(n31504), .Z(n31505) );
  XOR2_X1 U46474 ( .A1(n44350), .A2(n31505), .Z(n31506) );
  XOR2_X1 U46475 ( .A1(n50666), .A2(n31506), .Z(n31507) );
  XOR2_X1 U46477 ( .A1(n33164), .A2(n32574), .Z(n31734) );
  XOR2_X1 U46478 ( .A1(n32232), .A2(n24044), .Z(n39374) );
  XOR2_X1 U46479 ( .A1(n33165), .A2(n53713), .Z(n39200) );
  XOR2_X1 U46480 ( .A1(n39374), .A2(n39200), .Z(n36734) );
  XOR2_X1 U46481 ( .A1(n23851), .A2(n53772), .Z(n33167) );
  XOR2_X1 U46482 ( .A1(n31510), .A2(n33167), .Z(n37465) );
  XOR2_X1 U46483 ( .A1(n37465), .A2(n38277), .Z(n37883) );
  XOR2_X1 U46486 ( .A1(n31511), .A2(n15725), .Z(n31512) );
  XOR2_X1 U46487 ( .A1(n31925), .A2(n32572), .Z(n31513) );
  NOR2_X1 U46488 ( .A1(n34045), .A2(n33984), .ZN(n31516) );
  INV_X1 U46489 ( .I(n31535), .ZN(n31526) );
  XOR2_X1 U46490 ( .A1(n46398), .A2(n55368), .Z(n38882) );
  XOR2_X1 U46491 ( .A1(n27640), .A2(n56322), .Z(n50746) );
  XOR2_X1 U46492 ( .A1(n46601), .A2(n50746), .Z(n31520) );
  XOR2_X1 U46493 ( .A1(n38882), .A2(n31520), .Z(n31521) );
  XOR2_X1 U46494 ( .A1(n22961), .A2(n52327), .Z(n52449) );
  XOR2_X1 U46495 ( .A1(n31521), .A2(n52449), .Z(n31522) );
  NOR2_X1 U46496 ( .A1(n33963), .A2(n22226), .ZN(n31523) );
  NOR2_X1 U46497 ( .A1(n20800), .A2(n31523), .ZN(n31524) );
  NOR2_X1 U46499 ( .A1(n4075), .A2(n22226), .ZN(n31539) );
  INV_X1 U46500 ( .I(n31539), .ZN(n31529) );
  NAND2_X1 U46501 ( .A1(n31530), .A2(n34042), .ZN(n31531) );
  INV_X1 U46503 ( .I(n31538), .ZN(n31532) );
  INV_X1 U46505 ( .I(n35486), .ZN(n31542) );
  MUX2_X1 U46506 ( .I0(n7598), .I1(n22267), .S(n21010), .Z(n31544) );
  INV_X1 U46507 ( .I(n34860), .ZN(n31543) );
  NOR2_X1 U46508 ( .A1(n2699), .A2(n35903), .ZN(n34865) );
  NAND2_X1 U46510 ( .A1(n34865), .A2(n37031), .ZN(n31546) );
  NAND3_X1 U46511 ( .A1(n37031), .A2(n37030), .A3(n60659), .ZN(n31545) );
  INV_X1 U46512 ( .I(n50505), .ZN(n36008) );
  XOR2_X1 U46513 ( .A1(n37630), .A2(n36008), .Z(n49448) );
  INV_X1 U46514 ( .I(n49448), .ZN(n38628) );
  XOR2_X1 U46515 ( .A1(n38628), .A2(n23858), .Z(n38713) );
  XOR2_X1 U46516 ( .A1(n39469), .A2(n53499), .Z(n43615) );
  XOR2_X1 U46517 ( .A1(n24057), .A2(n53344), .Z(n38625) );
  XOR2_X1 U46518 ( .A1(n38625), .A2(n57131), .Z(n49445) );
  XOR2_X1 U46519 ( .A1(n43615), .A2(n49445), .Z(n31552) );
  XOR2_X1 U46520 ( .A1(n15712), .A2(n53272), .Z(n37795) );
  XOR2_X1 U46521 ( .A1(n31552), .A2(n31551), .Z(n31553) );
  XOR2_X1 U46522 ( .A1(n38713), .A2(n31553), .Z(n31554) );
  XOR2_X1 U46524 ( .A1(n44914), .A2(n31558), .Z(n51735) );
  XOR2_X1 U46525 ( .A1(n51735), .A2(n52970), .Z(n45474) );
  XOR2_X1 U46526 ( .A1(n33165), .A2(n55118), .Z(n37305) );
  XOR2_X1 U46527 ( .A1(n39530), .A2(n24044), .Z(n38995) );
  XOR2_X1 U46528 ( .A1(n37305), .A2(n38995), .Z(n45328) );
  XOR2_X1 U46529 ( .A1(n45328), .A2(n55335), .Z(n31559) );
  XOR2_X1 U46530 ( .A1(n45474), .A2(n31559), .Z(n31560) );
  XOR2_X1 U46531 ( .A1(n31561), .A2(n31560), .Z(n31562) );
  XOR2_X1 U46532 ( .A1(n31563), .A2(n31562), .Z(n31565) );
  XOR2_X1 U46533 ( .A1(n727), .A2(n55516), .Z(n31739) );
  XOR2_X1 U46535 ( .A1(n32472), .A2(n51569), .Z(n32729) );
  XOR2_X1 U46536 ( .A1(n36632), .A2(n32729), .Z(n38250) );
  XOR2_X1 U46537 ( .A1(n38639), .A2(n51765), .Z(n51609) );
  XOR2_X1 U46538 ( .A1(n51609), .A2(n53064), .Z(n31566) );
  XOR2_X1 U46539 ( .A1(n38250), .A2(n31566), .Z(n46239) );
  XOR2_X1 U46540 ( .A1(n61737), .A2(n57113), .Z(n35372) );
  XOR2_X1 U46541 ( .A1(n35372), .A2(n55052), .Z(n38723) );
  XOR2_X1 U46542 ( .A1(n38723), .A2(n52513), .Z(n42625) );
  INV_X1 U46544 ( .I(n31569), .ZN(n31570) );
  INV_X1 U46545 ( .I(n31574), .ZN(n31575) );
  NOR2_X2 U46546 ( .A1(n31576), .A2(n31575), .ZN(n33177) );
  XOR2_X1 U46547 ( .A1(n33283), .A2(n32326), .Z(n31579) );
  XOR2_X1 U46548 ( .A1(n17781), .A2(n31579), .Z(n31583) );
  XOR2_X1 U46551 ( .A1(n9722), .A2(n51946), .Z(n39352) );
  XOR2_X1 U46552 ( .A1(n36860), .A2(n39352), .Z(n44318) );
  XOR2_X1 U46553 ( .A1(n65171), .A2(n44318), .Z(n31585) );
  INV_X1 U46554 ( .I(n32595), .ZN(n31587) );
  XOR2_X1 U46555 ( .A1(n32658), .A2(n39650), .Z(n44414) );
  XOR2_X1 U46556 ( .A1(n44414), .A2(n50551), .Z(n45317) );
  XOR2_X1 U46557 ( .A1(n45317), .A2(n54185), .Z(n31588) );
  XOR2_X1 U46558 ( .A1(n15733), .A2(n31588), .Z(n31589) );
  XOR2_X1 U46559 ( .A1(n31589), .A2(n32387), .Z(n31591) );
  XOR2_X1 U46560 ( .A1(n45026), .A2(n23882), .Z(n44809) );
  XOR2_X1 U46561 ( .A1(n44014), .A2(n55126), .Z(n38111) );
  XOR2_X1 U46562 ( .A1(n38111), .A2(n38154), .Z(n37703) );
  XOR2_X1 U46563 ( .A1(n44809), .A2(n37703), .Z(n45105) );
  XOR2_X1 U46564 ( .A1(n31593), .A2(n32189), .Z(n31661) );
  INV_X1 U46565 ( .I(n31661), .ZN(n46554) );
  XOR2_X1 U46566 ( .A1(n54386), .A2(n55546), .Z(n31594) );
  XOR2_X1 U46567 ( .A1(n46554), .A2(n31594), .Z(n31595) );
  XOR2_X1 U46569 ( .A1(n44925), .A2(n44533), .Z(n32537) );
  XOR2_X1 U46570 ( .A1(n32537), .A2(n37896), .Z(n51817) );
  XOR2_X1 U46571 ( .A1(n53124), .A2(n53308), .Z(n38665) );
  XOR2_X1 U46572 ( .A1(n23999), .A2(n55395), .Z(n38238) );
  XOR2_X1 U46573 ( .A1(n38665), .A2(n38238), .Z(n38448) );
  XOR2_X1 U46574 ( .A1(n52232), .A2(n54936), .Z(n31601) );
  XOR2_X1 U46575 ( .A1(n1190), .A2(n31601), .Z(n31602) );
  NAND3_X1 U46576 ( .A1(n34152), .A2(n31608), .A3(n31607), .ZN(n31610) );
  XOR2_X1 U46577 ( .A1(n39363), .A2(n45404), .Z(n31613) );
  BUF_X2 U46578 ( .I(n31613), .Z(n51234) );
  XOR2_X1 U46579 ( .A1(n51234), .A2(n49434), .Z(n31617) );
  XOR2_X1 U46580 ( .A1(n56180), .A2(n53090), .Z(n31614) );
  XOR2_X1 U46581 ( .A1(n52135), .A2(n31614), .Z(n31615) );
  XOR2_X1 U46582 ( .A1(n24051), .A2(n53272), .Z(n43969) );
  XOR2_X1 U46583 ( .A1(n31615), .A2(n43969), .Z(n31616) );
  XOR2_X1 U46584 ( .A1(n31617), .A2(n31616), .Z(n31618) );
  XOR2_X1 U46585 ( .A1(n38400), .A2(n52095), .Z(n38430) );
  XOR2_X1 U46587 ( .A1(n31622), .A2(n15710), .Z(n32670) );
  XOR2_X1 U46588 ( .A1(n57096), .A2(n53318), .Z(n38556) );
  XOR2_X1 U46589 ( .A1(n38556), .A2(n54126), .Z(n33234) );
  XOR2_X1 U46590 ( .A1(n32670), .A2(n33234), .Z(n50578) );
  XOR2_X1 U46591 ( .A1(n52900), .A2(n55118), .Z(n35523) );
  XOR2_X1 U46592 ( .A1(n35523), .A2(n54870), .Z(n31856) );
  XNOR2_X1 U46593 ( .A1(n56905), .A2(n51492), .ZN(n31623) );
  XOR2_X1 U46594 ( .A1(n53713), .A2(n53246), .Z(n38825) );
  XOR2_X1 U46595 ( .A1(n31623), .A2(n38825), .Z(n31624) );
  XOR2_X1 U46596 ( .A1(n31856), .A2(n31624), .Z(n45255) );
  XOR2_X1 U46597 ( .A1(n45255), .A2(n55034), .Z(n31625) );
  XOR2_X1 U46598 ( .A1(n50578), .A2(n31625), .Z(n31626) );
  XOR2_X1 U46599 ( .A1(n31626), .A2(n59521), .Z(n31627) );
  XOR2_X1 U46600 ( .A1(n32573), .A2(n31627), .Z(n31628) );
  XOR2_X1 U46602 ( .A1(n51193), .A2(n54936), .Z(n50698) );
  XOR2_X1 U46603 ( .A1(n61550), .A2(n55106), .Z(n46487) );
  XOR2_X1 U46604 ( .A1(n50698), .A2(n46487), .Z(n31633) );
  XOR2_X1 U46605 ( .A1(n31634), .A2(n31633), .Z(n44949) );
  XOR2_X1 U46606 ( .A1(n49289), .A2(n50486), .Z(n46114) );
  XOR2_X1 U46607 ( .A1(n46114), .A2(n56976), .Z(n31635) );
  XOR2_X1 U46608 ( .A1(n32123), .A2(n53262), .Z(n45878) );
  XOR2_X1 U46609 ( .A1(n45026), .A2(n55349), .Z(n31638) );
  XOR2_X1 U46610 ( .A1(n55196), .A2(n55546), .Z(n39666) );
  XOR2_X1 U46611 ( .A1(n39666), .A2(n51019), .Z(n38734) );
  XOR2_X1 U46612 ( .A1(n38734), .A2(n51379), .Z(n46388) );
  XOR2_X1 U46613 ( .A1(n31638), .A2(n46388), .Z(n31639) );
  XOR2_X1 U46614 ( .A1(n31642), .A2(n53102), .Z(n45288) );
  XOR2_X1 U46615 ( .A1(n45288), .A2(n53833), .Z(n51215) );
  XOR2_X1 U46616 ( .A1(n39352), .A2(n31643), .Z(n52069) );
  XOR2_X1 U46617 ( .A1(n52069), .A2(n55379), .Z(n31644) );
  XOR2_X1 U46618 ( .A1(n65171), .A2(n31644), .Z(n31645) );
  XOR2_X1 U46619 ( .A1(n51215), .A2(n31645), .Z(n31646) );
  XOR2_X1 U46620 ( .A1(n13956), .A2(n33177), .Z(n31648) );
  XOR2_X1 U46621 ( .A1(n50798), .A2(n56849), .Z(n32558) );
  XOR2_X1 U46622 ( .A1(n32558), .A2(n35372), .Z(n44967) );
  XOR2_X1 U46623 ( .A1(n15707), .A2(n54888), .Z(n46128) );
  XOR2_X1 U46624 ( .A1(n44967), .A2(n46128), .Z(n45134) );
  XOR2_X1 U46625 ( .A1(n31649), .A2(n37844), .Z(n38949) );
  XOR2_X1 U46626 ( .A1(n38949), .A2(n55765), .Z(n31650) );
  XOR2_X1 U46627 ( .A1(n45134), .A2(n31650), .Z(n31651) );
  XOR2_X1 U46629 ( .A1(n50025), .A2(n52294), .Z(n42391) );
  XOR2_X1 U46630 ( .A1(n33185), .A2(n42391), .Z(n31653) );
  NAND3_X1 U46631 ( .A1(n31656), .A2(n33406), .A3(n7311), .ZN(n31660) );
  NOR2_X1 U46632 ( .A1(n33406), .A2(n23127), .ZN(n31658) );
  XOR2_X1 U46636 ( .A1(n37767), .A2(n53076), .Z(n36319) );
  XOR2_X1 U46637 ( .A1(n53262), .A2(n54231), .Z(n31663) );
  XOR2_X1 U46638 ( .A1(n36319), .A2(n31663), .Z(n44933) );
  XOR2_X1 U46639 ( .A1(n55546), .A2(n55349), .Z(n31664) );
  XOR2_X1 U46640 ( .A1(n44933), .A2(n31664), .Z(n31665) );
  XOR2_X1 U46641 ( .A1(n52366), .A2(n31665), .Z(n31666) );
  XOR2_X1 U46643 ( .A1(n57162), .A2(n55242), .Z(n31990) );
  XOR2_X1 U46644 ( .A1(n55106), .A2(n52232), .Z(n31745) );
  XOR2_X1 U46645 ( .A1(n31990), .A2(n31745), .Z(n39458) );
  XOR2_X1 U46646 ( .A1(n32741), .A2(n23999), .Z(n32178) );
  XOR2_X1 U46647 ( .A1(n39458), .A2(n32178), .Z(n46275) );
  XOR2_X1 U46648 ( .A1(n46275), .A2(n51193), .Z(n31670) );
  XOR2_X1 U46649 ( .A1(n1190), .A2(n23968), .Z(n51913) );
  XOR2_X1 U46650 ( .A1(n51913), .A2(n54776), .Z(n52167) );
  XOR2_X1 U46651 ( .A1(n46276), .A2(n52167), .Z(n31669) );
  XOR2_X1 U46652 ( .A1(n31670), .A2(n31669), .Z(n31671) );
  XOR2_X1 U46653 ( .A1(n32540), .A2(n31671), .Z(n31672) );
  XOR2_X1 U46654 ( .A1(n31677), .A2(n31676), .Z(n31678) );
  XOR2_X1 U46655 ( .A1(n54888), .A2(n53064), .Z(n32401) );
  XOR2_X1 U46656 ( .A1(n32401), .A2(n39631), .Z(n38532) );
  XOR2_X1 U46657 ( .A1(n38532), .A2(n52294), .Z(n46323) );
  XOR2_X1 U46658 ( .A1(n51968), .A2(n46323), .Z(n31680) );
  XOR2_X1 U46659 ( .A1(n55862), .A2(n55340), .Z(n46336) );
  XOR2_X1 U46660 ( .A1(n31685), .A2(n31684), .Z(n31710) );
  XOR2_X1 U46661 ( .A1(n33896), .A2(n32515), .Z(n32596) );
  XOR2_X1 U46662 ( .A1(n59638), .A2(n39434), .Z(n51978) );
  XOR2_X1 U46663 ( .A1(n37637), .A2(n53102), .Z(n37838) );
  XOR2_X1 U46664 ( .A1(n50551), .A2(n55379), .Z(n31689) );
  XOR2_X1 U46665 ( .A1(n37838), .A2(n31689), .Z(n45388) );
  XOR2_X1 U46666 ( .A1(n51978), .A2(n45388), .Z(n31690) );
  XOR2_X1 U46667 ( .A1(n32388), .A2(n31690), .Z(n31691) );
  XOR2_X1 U46668 ( .A1(n31692), .A2(n31691), .Z(n31693) );
  XOR2_X1 U46669 ( .A1(n60799), .A2(n39200), .Z(n38279) );
  XOR2_X1 U46670 ( .A1(n38279), .A2(n51494), .Z(n45416) );
  XOR2_X1 U46671 ( .A1(n56827), .A2(n55034), .Z(n32310) );
  XOR2_X1 U46672 ( .A1(n32310), .A2(n53772), .Z(n31694) );
  XOR2_X1 U46673 ( .A1(n31694), .A2(n38556), .Z(n44297) );
  XOR2_X1 U46674 ( .A1(n39478), .A2(n52970), .Z(n44631) );
  XOR2_X1 U46675 ( .A1(n51881), .A2(n51493), .Z(n51165) );
  XOR2_X1 U46676 ( .A1(n44631), .A2(n51165), .Z(n31695) );
  XOR2_X1 U46677 ( .A1(n44297), .A2(n31695), .Z(n31696) );
  XOR2_X1 U46678 ( .A1(n23260), .A2(n31924), .Z(n31700) );
  XOR2_X1 U46679 ( .A1(n38074), .A2(n37481), .Z(n52100) );
  XOR2_X1 U46680 ( .A1(n52100), .A2(n53499), .Z(n43803) );
  XOR2_X1 U46681 ( .A1(n52095), .A2(n53154), .Z(n44107) );
  XOR2_X1 U46682 ( .A1(n44107), .A2(n50505), .Z(n51007) );
  XNOR2_X1 U46683 ( .A1(n56322), .A2(n53344), .ZN(n31703) );
  XOR2_X1 U46684 ( .A1(n51007), .A2(n31703), .Z(n44047) );
  XOR2_X1 U46685 ( .A1(n46601), .A2(n58084), .Z(n51479) );
  XOR2_X1 U46686 ( .A1(n44047), .A2(n51479), .Z(n31704) );
  XOR2_X1 U46687 ( .A1(n43803), .A2(n31704), .Z(n31705) );
  NOR2_X1 U46688 ( .A1(n32695), .A2(n157), .ZN(n31709) );
  NAND2_X1 U46690 ( .A1(n34132), .A2(n6925), .ZN(n31711) );
  INV_X1 U46691 ( .I(n33654), .ZN(n33660) );
  INV_X1 U46694 ( .I(n34144), .ZN(n31716) );
  NOR2_X1 U46695 ( .A1(n22598), .A2(n6925), .ZN(n31715) );
  NAND2_X1 U46697 ( .A1(n60554), .A2(n24664), .ZN(n31720) );
  AOI21_X1 U46698 ( .A1(n33998), .A2(n31720), .B(n34168), .ZN(n31721) );
  INV_X1 U46699 ( .I(n34116), .ZN(n31722) );
  NOR2_X1 U46701 ( .A1(n34114), .A2(n60808), .ZN(n31725) );
  INV_X1 U46702 ( .I(n33950), .ZN(n31727) );
  AOI22_X1 U46703 ( .A1(n32862), .A2(n15783), .B1(n34118), .B2(n34114), .ZN(
        n31728) );
  XOR2_X1 U46705 ( .A1(n23869), .A2(n15725), .Z(n32091) );
  XOR2_X1 U46707 ( .A1(n39373), .A2(n50498), .Z(n38650) );
  XOR2_X1 U46708 ( .A1(n37303), .A2(n54517), .Z(n38387) );
  XOR2_X1 U46709 ( .A1(n38387), .A2(n24044), .Z(n31735) );
  XOR2_X1 U46710 ( .A1(n38650), .A2(n31735), .Z(n45827) );
  XOR2_X1 U46711 ( .A1(n33234), .A2(n38653), .Z(n44632) );
  XOR2_X1 U46712 ( .A1(n44632), .A2(n52970), .Z(n31736) );
  XOR2_X1 U46713 ( .A1(n45827), .A2(n31736), .Z(n31737) );
  XOR2_X1 U46714 ( .A1(n32001), .A2(n31737), .Z(n31738) );
  XOR2_X1 U46715 ( .A1(n31740), .A2(n31739), .Z(n31741) );
  XOR2_X1 U46716 ( .A1(n52375), .A2(n55603), .Z(n38862) );
  XOR2_X1 U46717 ( .A1(n38862), .A2(n31745), .Z(n41498) );
  XOR2_X1 U46718 ( .A1(n53530), .A2(n24061), .Z(n38743) );
  XOR2_X1 U46719 ( .A1(n38502), .A2(n38743), .Z(n32500) );
  INV_X1 U46720 ( .I(n32500), .ZN(n31747) );
  XOR2_X1 U46721 ( .A1(n31747), .A2(n31746), .Z(n50701) );
  XOR2_X1 U46722 ( .A1(n50701), .A2(n53308), .Z(n44728) );
  XOR2_X1 U46723 ( .A1(n845), .A2(n37704), .Z(n31751) );
  XOR2_X1 U46724 ( .A1(n38153), .A2(n31751), .Z(n46124) );
  XOR2_X1 U46725 ( .A1(n29969), .A2(n53262), .Z(n31752) );
  XOR2_X1 U46726 ( .A1(n43065), .A2(n31752), .Z(n44960) );
  XOR2_X1 U46727 ( .A1(n23249), .A2(n52513), .Z(n45130) );
  XOR2_X1 U46728 ( .A1(n45130), .A2(n31755), .Z(n42578) );
  XOR2_X1 U46729 ( .A1(n32401), .A2(n51611), .Z(n31756) );
  XOR2_X1 U46730 ( .A1(n37730), .A2(n31756), .Z(n44741) );
  XOR2_X1 U46731 ( .A1(n44741), .A2(n31757), .Z(n31758) );
  XOR2_X1 U46732 ( .A1(n42578), .A2(n31758), .Z(n31759) );
  XOR2_X1 U46733 ( .A1(n32408), .A2(n31760), .Z(n31761) );
  XOR2_X1 U46734 ( .A1(n4795), .A2(n33283), .Z(n32065) );
  XOR2_X1 U46735 ( .A1(n32010), .A2(n23714), .Z(n31764) );
  XOR2_X1 U46736 ( .A1(n55638), .A2(n55379), .Z(n37837) );
  XOR2_X1 U46737 ( .A1(n23929), .A2(n53284), .Z(n48967) );
  XOR2_X1 U46738 ( .A1(n37837), .A2(n48967), .Z(n50985) );
  XOR2_X1 U46739 ( .A1(n50985), .A2(n52470), .Z(n45847) );
  AOI22_X1 U46740 ( .A1(n32833), .A2(n58447), .B1(n10401), .B2(n5386), .ZN(
        n31778) );
  XOR2_X1 U46741 ( .A1(n37749), .A2(n39469), .Z(n50509) );
  XOR2_X1 U46742 ( .A1(n50509), .A2(n58084), .Z(n45278) );
  XOR2_X1 U46743 ( .A1(n50505), .A2(n38625), .Z(n50248) );
  XOR2_X1 U46744 ( .A1(n52135), .A2(n23858), .Z(n31769) );
  XOR2_X1 U46745 ( .A1(n50248), .A2(n31769), .Z(n44185) );
  INV_X1 U46746 ( .I(n22961), .ZN(n31770) );
  XOR2_X1 U46747 ( .A1(n44185), .A2(n31770), .Z(n31771) );
  XOR2_X1 U46748 ( .A1(n55368), .A2(n55624), .Z(n44046) );
  NAND2_X1 U46749 ( .A1(n31767), .A2(n34198), .ZN(n31776) );
  NAND2_X1 U46750 ( .A1(n35883), .A2(n35881), .ZN(n31780) );
  NOR2_X1 U46751 ( .A1(n35885), .A2(n7488), .ZN(n31785) );
  OAI21_X1 U46752 ( .A1(n31786), .A2(n1779), .B(n31785), .ZN(n31787) );
  OAI22_X1 U46754 ( .A1(n35901), .A2(n34878), .B1(n34491), .B2(n1779), .ZN(
        n31789) );
  XOR2_X1 U46756 ( .A1(n52029), .A2(n55792), .Z(n45276) );
  XOR2_X1 U46757 ( .A1(n45276), .A2(n38885), .Z(n45359) );
  XOR2_X1 U46758 ( .A1(n45274), .A2(n37481), .Z(n32364) );
  INV_X1 U46759 ( .I(n32364), .ZN(n31792) );
  XOR2_X1 U46760 ( .A1(n31792), .A2(n22773), .Z(n39536) );
  XOR2_X1 U46761 ( .A1(n55368), .A2(n55139), .Z(n44108) );
  XOR2_X1 U46762 ( .A1(n44108), .A2(n50745), .Z(n31793) );
  XOR2_X1 U46763 ( .A1(n37749), .A2(n31793), .Z(n31794) );
  INV_X1 U46764 ( .I(n31797), .ZN(n31798) );
  XOR2_X1 U46765 ( .A1(n33164), .A2(n31798), .Z(n31799) );
  XOR2_X1 U46767 ( .A1(n32001), .A2(n15725), .Z(n32721) );
  XOR2_X1 U46769 ( .A1(n51494), .A2(n24105), .Z(n31801) );
  XOR2_X1 U46770 ( .A1(n31801), .A2(n38388), .Z(n38440) );
  XOR2_X1 U46771 ( .A1(n38440), .A2(n37303), .Z(n32416) );
  XOR2_X1 U46772 ( .A1(n32416), .A2(n39373), .Z(n45049) );
  XOR2_X1 U46773 ( .A1(n45049), .A2(n46443), .Z(n31802) );
  XOR2_X1 U46774 ( .A1(n31803), .A2(n31855), .Z(n31808) );
  XOR2_X1 U46775 ( .A1(n23869), .A2(n17463), .Z(n31806) );
  XOR2_X1 U46777 ( .A1(n37713), .A2(n55655), .Z(n31811) );
  XOR2_X1 U46778 ( .A1(n31811), .A2(n50486), .Z(n33062) );
  XOR2_X1 U46779 ( .A1(n38378), .A2(n33062), .Z(n43962) );
  XNOR2_X1 U46780 ( .A1(n23455), .A2(n55603), .ZN(n31812) );
  XOR2_X1 U46781 ( .A1(n23789), .A2(n31812), .Z(n44255) );
  XOR2_X1 U46782 ( .A1(n44255), .A2(n50787), .Z(n31813) );
  XOR2_X1 U46783 ( .A1(n43962), .A2(n31813), .Z(n31814) );
  XOR2_X1 U46784 ( .A1(n38851), .A2(n32189), .Z(n33148) );
  XOR2_X1 U46785 ( .A1(n50955), .A2(n54153), .Z(n39217) );
  XOR2_X1 U46786 ( .A1(n30908), .A2(n56040), .Z(n36656) );
  XOR2_X1 U46787 ( .A1(n39217), .A2(n36656), .Z(n31817) );
  XOR2_X1 U46788 ( .A1(n33148), .A2(n31817), .Z(n43006) );
  XNOR2_X1 U46789 ( .A1(n53958), .A2(n50831), .ZN(n31818) );
  XOR2_X1 U46790 ( .A1(n39771), .A2(n31818), .Z(n46221) );
  XOR2_X1 U46791 ( .A1(n46221), .A2(n56915), .Z(n31819) );
  XOR2_X1 U46792 ( .A1(n43006), .A2(n31819), .Z(n31820) );
  XOR2_X1 U46793 ( .A1(n16820), .A2(n31820), .Z(n31821) );
  NOR2_X1 U46794 ( .A1(n5099), .A2(n35272), .ZN(n31834) );
  XOR2_X1 U46795 ( .A1(n32585), .A2(n31823), .Z(n32524) );
  INV_X1 U46796 ( .I(n51275), .ZN(n31824) );
  XOR2_X1 U46797 ( .A1(n32519), .A2(n31824), .Z(n49088) );
  XOR2_X1 U46798 ( .A1(n57142), .A2(n65079), .Z(n31825) );
  XOR2_X1 U46799 ( .A1(n38472), .A2(n31825), .Z(n31826) );
  XOR2_X1 U46800 ( .A1(n45389), .A2(n31826), .Z(n46425) );
  XOR2_X1 U46801 ( .A1(n55379), .A2(n24109), .Z(n31875) );
  XOR2_X1 U46802 ( .A1(n23929), .A2(n55889), .Z(n37256) );
  XOR2_X1 U46803 ( .A1(n31875), .A2(n37256), .Z(n45059) );
  XOR2_X1 U46804 ( .A1(n46425), .A2(n45059), .Z(n31827) );
  XOR2_X1 U46806 ( .A1(n33904), .A2(n30402), .Z(n31830) );
  XOR2_X1 U46807 ( .A1(n64794), .A2(n31830), .Z(n31831) );
  XOR2_X1 U46808 ( .A1(n42426), .A2(n60857), .Z(n38186) );
  XOR2_X1 U46809 ( .A1(n38186), .A2(n23249), .Z(n46324) );
  XOR2_X1 U46810 ( .A1(n46324), .A2(n54708), .Z(n49233) );
  XOR2_X1 U46811 ( .A1(n49233), .A2(n55534), .Z(n44274) );
  XOR2_X1 U46812 ( .A1(n15707), .A2(n52197), .Z(n32249) );
  XOR2_X1 U46813 ( .A1(n32249), .A2(n54219), .Z(n43884) );
  XOR2_X1 U46814 ( .A1(n55340), .A2(n52317), .Z(n31837) );
  XOR2_X1 U46815 ( .A1(n43884), .A2(n31837), .Z(n31838) );
  XOR2_X1 U46816 ( .A1(n17668), .A2(n31838), .Z(n31839) );
  NAND2_X1 U46817 ( .A1(n34221), .A2(n61458), .ZN(n31843) );
  OAI21_X1 U46818 ( .A1(n35807), .A2(n31843), .B(n34389), .ZN(n31844) );
  OAI22_X1 U46819 ( .A1(n34294), .A2(n35279), .B1(n34385), .B2(n35280), .ZN(
        n31846) );
  XOR2_X1 U46820 ( .A1(n44378), .A2(n55624), .Z(n31847) );
  XOR2_X1 U46821 ( .A1(n51394), .A2(n31847), .Z(n31848) );
  XOR2_X1 U46822 ( .A1(n14666), .A2(n52226), .Z(n31852) );
  XOR2_X1 U46823 ( .A1(n32085), .A2(n31852), .Z(n31853) );
  XOR2_X1 U46824 ( .A1(n37584), .A2(n39375), .Z(n39194) );
  XOR2_X1 U46825 ( .A1(n39194), .A2(n39707), .Z(n38824) );
  XOR2_X1 U46826 ( .A1(n38824), .A2(n53318), .Z(n45330) );
  XOR2_X1 U46827 ( .A1(n31856), .A2(n56143), .Z(n44513) );
  XOR2_X1 U46828 ( .A1(n45330), .A2(n44513), .Z(n31857) );
  XOR2_X1 U46829 ( .A1(n50533), .A2(n55052), .Z(n37729) );
  XOR2_X1 U46830 ( .A1(n37729), .A2(n52196), .Z(n46238) );
  XOR2_X1 U46831 ( .A1(n43884), .A2(n46238), .Z(n31860) );
  XOR2_X1 U46832 ( .A1(n23424), .A2(n31860), .Z(n31861) );
  XOR2_X1 U46833 ( .A1(n18838), .A2(n31862), .Z(n31865) );
  XOR2_X1 U46834 ( .A1(n55191), .A2(n57113), .Z(n46230) );
  XOR2_X1 U46835 ( .A1(n65041), .A2(n46230), .Z(n31864) );
  XOR2_X1 U46836 ( .A1(n43858), .A2(n53174), .Z(n32168) );
  XOR2_X1 U46837 ( .A1(n50682), .A2(n53359), .Z(n39752) );
  XOR2_X1 U46838 ( .A1(n32168), .A2(n39752), .Z(n45314) );
  XOR2_X1 U46839 ( .A1(n32338), .A2(n45314), .Z(n31869) );
  XOR2_X1 U46840 ( .A1(n31870), .A2(n31869), .Z(n32386) );
  XOR2_X1 U46842 ( .A1(n23791), .A2(n33242), .Z(n31874) );
  XOR2_X1 U46843 ( .A1(n31874), .A2(n23714), .Z(n32166) );
  XOR2_X1 U46844 ( .A1(n61034), .A2(n31875), .Z(n31876) );
  XOR2_X1 U46845 ( .A1(n31877), .A2(n31876), .Z(n44502) );
  XOR2_X1 U46846 ( .A1(n44502), .A2(n56335), .Z(n31878) );
  XOR2_X1 U46847 ( .A1(n23786), .A2(n31878), .Z(n31879) );
  XOR2_X1 U46848 ( .A1(n32166), .A2(n31879), .Z(n31881) );
  XOR2_X1 U46849 ( .A1(n31881), .A2(n31880), .Z(n31882) );
  XOR2_X1 U46850 ( .A1(n31883), .A2(n31882), .Z(n32430) );
  INV_X1 U46851 ( .I(n45371), .ZN(n31887) );
  XOR2_X1 U46852 ( .A1(n23789), .A2(n31887), .Z(n39682) );
  XOR2_X1 U46853 ( .A1(n39682), .A2(n38448), .Z(n37712) );
  XOR2_X1 U46854 ( .A1(n39457), .A2(n23455), .Z(n37739) );
  XOR2_X1 U46855 ( .A1(n37712), .A2(n37739), .Z(n46183) );
  XOR2_X1 U46856 ( .A1(n38743), .A2(n55242), .Z(n50196) );
  XOR2_X1 U46857 ( .A1(n51193), .A2(n56976), .Z(n31888) );
  XOR2_X1 U46858 ( .A1(n50196), .A2(n31888), .Z(n31889) );
  XOR2_X1 U46859 ( .A1(n46183), .A2(n31889), .Z(n31890) );
  XOR2_X1 U46862 ( .A1(n31892), .A2(n32747), .Z(n31894) );
  XOR2_X1 U46863 ( .A1(n32123), .A2(n56915), .Z(n38830) );
  XOR2_X1 U46864 ( .A1(n37767), .A2(n23882), .Z(n31895) );
  XOR2_X1 U46865 ( .A1(n38830), .A2(n31895), .Z(n31896) );
  XOR2_X1 U46866 ( .A1(n31896), .A2(n39771), .Z(n46555) );
  XOR2_X1 U46867 ( .A1(n38614), .A2(n55196), .Z(n45103) );
  XOR2_X1 U46868 ( .A1(n51999), .A2(n55349), .Z(n31897) );
  XOR2_X1 U46869 ( .A1(n45103), .A2(n31897), .Z(n31898) );
  XOR2_X1 U46870 ( .A1(n46555), .A2(n31898), .Z(n31899) );
  XOR2_X1 U46871 ( .A1(n20058), .A2(n31899), .Z(n31900) );
  NAND4_X2 U46875 ( .A1(n31909), .A2(n31908), .A3(n31907), .A4(n34220), .ZN(
        n31910) );
  XOR2_X1 U46876 ( .A1(n38743), .A2(n50475), .Z(n47768) );
  XOR2_X1 U46877 ( .A1(n47768), .A2(n56202), .Z(n39738) );
  XOR2_X1 U46878 ( .A1(n50793), .A2(n30564), .Z(n49273) );
  INV_X1 U46879 ( .I(n49273), .ZN(n37570) );
  XOR2_X1 U46880 ( .A1(n43720), .A2(n55833), .Z(n31914) );
  XOR2_X1 U46881 ( .A1(n44533), .A2(n53705), .Z(n38980) );
  XOR2_X1 U46882 ( .A1(n38980), .A2(n56124), .Z(n38798) );
  XOR2_X1 U46883 ( .A1(n38798), .A2(n39457), .Z(n44391) );
  XOR2_X1 U46884 ( .A1(n31914), .A2(n44391), .Z(n31915) );
  XOR2_X1 U46885 ( .A1(n5727), .A2(n31915), .Z(n31916) );
  XOR2_X1 U46886 ( .A1(n38154), .A2(n39570), .Z(n36320) );
  XOR2_X1 U46887 ( .A1(n32123), .A2(n54231), .Z(n31918) );
  XOR2_X1 U46888 ( .A1(n36320), .A2(n31918), .Z(n44085) );
  XOR2_X1 U46889 ( .A1(n39478), .A2(n52900), .Z(n39704) );
  XOR2_X1 U46890 ( .A1(n60799), .A2(n39704), .Z(n31920) );
  XOR2_X1 U46891 ( .A1(n38896), .A2(n55840), .Z(n44996) );
  XOR2_X1 U46892 ( .A1(n37465), .A2(n44996), .Z(n31919) );
  XOR2_X1 U46893 ( .A1(n31920), .A2(n31919), .Z(n45143) );
  XOR2_X1 U46894 ( .A1(n39196), .A2(n55516), .Z(n46532) );
  XOR2_X1 U46895 ( .A1(n46532), .A2(n38388), .Z(n31921) );
  XOR2_X1 U46896 ( .A1(n45143), .A2(n31921), .Z(n31922) );
  XOR2_X1 U46897 ( .A1(n31924), .A2(n31923), .Z(n31927) );
  XOR2_X1 U46898 ( .A1(n61304), .A2(n23389), .Z(n31929) );
  XOR2_X1 U46899 ( .A1(n52196), .A2(n55765), .Z(n32103) );
  XOR2_X1 U46900 ( .A1(n60857), .A2(n51610), .Z(n33281) );
  XOR2_X1 U46901 ( .A1(n32103), .A2(n33281), .Z(n33867) );
  INV_X1 U46902 ( .I(n33867), .ZN(n31931) );
  XOR2_X1 U46905 ( .A1(n52197), .A2(n39444), .Z(n51150) );
  XOR2_X1 U46906 ( .A1(n53945), .A2(n55862), .Z(n33180) );
  XOR2_X1 U46907 ( .A1(n33180), .A2(n23306), .Z(n31932) );
  XOR2_X1 U46908 ( .A1(n51150), .A2(n31932), .Z(n43682) );
  XOR2_X1 U46909 ( .A1(n44351), .A2(n43682), .Z(n31933) );
  XOR2_X1 U46911 ( .A1(n38772), .A2(n53989), .Z(n45123) );
  XOR2_X1 U46912 ( .A1(n111), .A2(n33193), .Z(n31936) );
  XOR2_X1 U46913 ( .A1(n31937), .A2(n31936), .Z(n31938) );
  XOR2_X1 U46914 ( .A1(n52178), .A2(n53174), .Z(n38301) );
  XOR2_X1 U46915 ( .A1(n38301), .A2(n53833), .Z(n31939) );
  XOR2_X1 U46916 ( .A1(n38302), .A2(n31939), .Z(n46524) );
  XOR2_X1 U46917 ( .A1(n46524), .A2(n30402), .Z(n31940) );
  XOR2_X1 U46918 ( .A1(n31940), .A2(n18314), .Z(n31941) );
  XOR2_X1 U46920 ( .A1(n23786), .A2(n33243), .Z(n32013) );
  XOR2_X1 U46922 ( .A1(n31943), .A2(n56949), .Z(n32060) );
  XOR2_X1 U46923 ( .A1(n1823), .A2(n32060), .Z(n31944) );
  XOR2_X1 U46924 ( .A1(n31945), .A2(n31944), .Z(n31946) );
  XOR2_X1 U46925 ( .A1(n50504), .A2(n37481), .Z(n39181) );
  XOR2_X1 U46926 ( .A1(n39181), .A2(n56495), .Z(n51596) );
  XOR2_X1 U46927 ( .A1(n51596), .A2(n51234), .Z(n31948) );
  XOR2_X1 U46928 ( .A1(n4561), .A2(n54168), .Z(n32224) );
  XOR2_X1 U46929 ( .A1(n32224), .A2(n56322), .Z(n31947) );
  XOR2_X1 U46930 ( .A1(n52097), .A2(n31947), .Z(n46603) );
  INV_X1 U46931 ( .I(n35255), .ZN(n35251) );
  NAND2_X1 U46932 ( .A1(n1794), .A2(n33814), .ZN(n31952) );
  NAND2_X1 U46934 ( .A1(n31954), .A2(n16203), .ZN(n31958) );
  XOR2_X1 U46935 ( .A1(n44112), .A2(n58084), .Z(n38397) );
  XOR2_X1 U46936 ( .A1(n50504), .A2(n53499), .Z(n44619) );
  XOR2_X1 U46937 ( .A1(n44619), .A2(n39363), .Z(n31959) );
  XOR2_X1 U46938 ( .A1(n38397), .A2(n31959), .Z(n44186) );
  XOR2_X1 U46939 ( .A1(n22323), .A2(n24057), .Z(n45275) );
  XOR2_X1 U46940 ( .A1(n31960), .A2(n45276), .Z(n31961) );
  XOR2_X1 U46941 ( .A1(n44186), .A2(n31961), .Z(n31962) );
  XOR2_X1 U46943 ( .A1(n15707), .A2(n22821), .Z(n42579) );
  XOR2_X1 U46944 ( .A1(n42391), .A2(n42579), .Z(n31969) );
  XOR2_X1 U46945 ( .A1(n52196), .A2(n24065), .Z(n31967) );
  XOR2_X1 U46946 ( .A1(n54376), .A2(n50817), .Z(n44739) );
  XOR2_X1 U46947 ( .A1(n31967), .A2(n44739), .Z(n31968) );
  XOR2_X1 U46948 ( .A1(n31969), .A2(n31968), .Z(n31971) );
  XOR2_X1 U46949 ( .A1(n31971), .A2(n4544), .Z(n31972) );
  XOR2_X1 U46950 ( .A1(n22162), .A2(n31973), .Z(n31974) );
  NOR2_X1 U46951 ( .A1(n35294), .A2(n31976), .ZN(n34340) );
  XOR2_X1 U46952 ( .A1(n23767), .A2(n38962), .Z(n39568) );
  XOR2_X1 U46953 ( .A1(n30908), .A2(n23882), .Z(n33147) );
  XOR2_X1 U46954 ( .A1(n39568), .A2(n33147), .Z(n48388) );
  XOR2_X1 U46955 ( .A1(n43065), .A2(n55349), .Z(n37458) );
  XOR2_X1 U46956 ( .A1(n37458), .A2(n56771), .Z(n31978) );
  XOR2_X1 U46957 ( .A1(n48388), .A2(n31978), .Z(n31979) );
  XOR2_X1 U46958 ( .A1(n32617), .A2(n31979), .Z(n31980) );
  XOR2_X1 U46959 ( .A1(n31987), .A2(n31986), .Z(n31988) );
  XOR2_X1 U46960 ( .A1(n39210), .A2(n55603), .Z(n39278) );
  XOR2_X1 U46961 ( .A1(n39278), .A2(n31990), .Z(n44727) );
  XOR2_X1 U46962 ( .A1(n44727), .A2(n54208), .Z(n31992) );
  XOR2_X1 U46963 ( .A1(n32274), .A2(n55395), .Z(n31991) );
  XOR2_X1 U46964 ( .A1(n39280), .A2(n31991), .Z(n51718) );
  XOR2_X1 U46965 ( .A1(n37713), .A2(n54587), .Z(n38326) );
  XOR2_X1 U46966 ( .A1(n38326), .A2(n1190), .Z(n38161) );
  XOR2_X1 U46967 ( .A1(n51718), .A2(n38161), .Z(n41497) );
  XOR2_X1 U46968 ( .A1(n31992), .A2(n41497), .Z(n31994) );
  XOR2_X1 U46969 ( .A1(n31993), .A2(n31994), .Z(n31995) );
  XOR2_X1 U46970 ( .A1(n32172), .A2(n53318), .Z(n45830) );
  INV_X1 U46971 ( .I(n32089), .ZN(n31996) );
  XOR2_X1 U46972 ( .A1(n31997), .A2(n31996), .Z(n31999) );
  NAND2_X1 U46973 ( .A1(n34335), .A2(n17958), .ZN(n32004) );
  OAI22_X1 U46974 ( .A1(n21056), .A2(n22278), .B1(n1802), .B2(n34268), .ZN(
        n32005) );
  NAND2_X1 U46975 ( .A1(n32005), .A2(n31976), .ZN(n32022) );
  XOR2_X1 U46977 ( .A1(n23714), .A2(n18296), .Z(n32009) );
  XOR2_X1 U46978 ( .A1(n38302), .A2(n32053), .Z(n45849) );
  XOR2_X1 U46979 ( .A1(n50985), .A2(n38772), .Z(n44615) );
  XOR2_X1 U46980 ( .A1(n44615), .A2(n52178), .Z(n32006) );
  XOR2_X1 U46981 ( .A1(n45849), .A2(n32006), .Z(n32007) );
  XOR2_X1 U46982 ( .A1(n32012), .A2(n32515), .Z(n32015) );
  XOR2_X1 U46983 ( .A1(n1823), .A2(n32013), .Z(n32014) );
  XOR2_X1 U46984 ( .A1(n32015), .A2(n32014), .Z(n32016) );
  NAND2_X1 U46986 ( .A1(n1802), .A2(n31976), .ZN(n32020) );
  INV_X1 U46987 ( .I(n37007), .ZN(n37336) );
  XOR2_X1 U46988 ( .A1(n32123), .A2(n44014), .Z(n50873) );
  XOR2_X1 U46989 ( .A1(n50873), .A2(n39771), .Z(n37143) );
  XOR2_X1 U46990 ( .A1(n37143), .A2(n32024), .Z(n46286) );
  XOR2_X1 U46991 ( .A1(n44808), .A2(n23882), .Z(n32025) );
  XOR2_X1 U46992 ( .A1(n46286), .A2(n32025), .Z(n32026) );
  XOR2_X1 U46993 ( .A1(n58077), .A2(n39457), .Z(n38981) );
  XOR2_X1 U46994 ( .A1(n38981), .A2(n55603), .Z(n39399) );
  XOR2_X1 U46995 ( .A1(n39399), .A2(n43485), .Z(n32033) );
  XOR2_X1 U46996 ( .A1(n50067), .A2(n55833), .Z(n32030) );
  XOR2_X1 U46997 ( .A1(n23789), .A2(n32030), .Z(n32031) );
  XOR2_X1 U46998 ( .A1(n55655), .A2(n55395), .Z(n37519) );
  XOR2_X1 U46999 ( .A1(n37519), .A2(n53124), .Z(n43498) );
  XOR2_X1 U47000 ( .A1(n32031), .A2(n43498), .Z(n32032) );
  XOR2_X1 U47001 ( .A1(n32033), .A2(n32032), .Z(n32034) );
  XOR2_X1 U47002 ( .A1(n55118), .A2(n24105), .Z(n32039) );
  XOR2_X1 U47003 ( .A1(n32040), .A2(n32039), .Z(n44443) );
  XOR2_X1 U47004 ( .A1(n38280), .A2(n46532), .Z(n32041) );
  XOR2_X1 U47005 ( .A1(n44443), .A2(n32041), .Z(n32042) );
  XOR2_X1 U47006 ( .A1(n22820), .A2(n32042), .Z(n32043) );
  XOR2_X1 U47007 ( .A1(n44759), .A2(n53499), .Z(n36215) );
  XOR2_X1 U47008 ( .A1(n36215), .A2(n39723), .Z(n44311) );
  XOR2_X1 U47009 ( .A1(n37481), .A2(n57131), .Z(n44309) );
  XOR2_X1 U47010 ( .A1(n51679), .A2(n44309), .Z(n32048) );
  XNOR2_X1 U47011 ( .A1(n23858), .A2(n4561), .ZN(n32047) );
  XOR2_X1 U47012 ( .A1(n44622), .A2(n32047), .Z(n45403) );
  XOR2_X1 U47013 ( .A1(n39752), .A2(n32053), .Z(n52577) );
  XOR2_X1 U47014 ( .A1(n38772), .A2(n23929), .Z(n44412) );
  XOR2_X1 U47015 ( .A1(n44412), .A2(n51275), .Z(n51947) );
  XOR2_X1 U47016 ( .A1(n52577), .A2(n51947), .Z(n32055) );
  INV_X1 U47017 ( .I(n44414), .ZN(n32054) );
  XOR2_X1 U47018 ( .A1(n32055), .A2(n32054), .Z(n32056) );
  XOR2_X1 U47019 ( .A1(n51667), .A2(n50025), .Z(n38948) );
  XOR2_X1 U47020 ( .A1(n38948), .A2(n51569), .Z(n33871) );
  INV_X1 U47021 ( .I(n36632), .ZN(n33280) );
  XOR2_X1 U47022 ( .A1(n33871), .A2(n33280), .Z(n43195) );
  XOR2_X1 U47023 ( .A1(n38947), .A2(n60857), .Z(n44093) );
  XOR2_X1 U47024 ( .A1(n57113), .A2(n23306), .Z(n52590) );
  XOR2_X1 U47025 ( .A1(n44093), .A2(n52590), .Z(n32061) );
  XOR2_X1 U47026 ( .A1(n43195), .A2(n32061), .Z(n32062) );
  XOR2_X1 U47027 ( .A1(n32062), .A2(n32640), .Z(n32063) );
  XOR2_X1 U47028 ( .A1(n32063), .A2(n1822), .Z(n32067) );
  XOR2_X1 U47029 ( .A1(n32064), .A2(n32065), .Z(n32066) );
  BUF_X2 U47030 ( .I(n32069), .Z(n34714) );
  INV_X1 U47031 ( .I(n35816), .ZN(n35306) );
  OAI22_X1 U47032 ( .A1(n34717), .A2(n34316), .B1(n35306), .B2(n57628), .ZN(
        n32074) );
  NAND2_X1 U47033 ( .A1(n32070), .A2(n35813), .ZN(n32072) );
  AOI21_X1 U47034 ( .A1(n35304), .A2(n32074), .B(n32073), .ZN(n32075) );
  XOR2_X1 U47035 ( .A1(n38885), .A2(n56065), .Z(n37869) );
  XOR2_X1 U47036 ( .A1(n44619), .A2(n37869), .Z(n32080) );
  XOR2_X1 U47037 ( .A1(n22773), .A2(n23886), .Z(n39361) );
  XOR2_X1 U47038 ( .A1(n24046), .A2(n56180), .Z(n50909) );
  XOR2_X1 U47039 ( .A1(n32078), .A2(n50909), .Z(n32079) );
  XOR2_X1 U47040 ( .A1(n32080), .A2(n32079), .Z(n32081) );
  XOR2_X1 U47041 ( .A1(n32081), .A2(n45819), .Z(n32082) );
  XOR2_X1 U47042 ( .A1(n37468), .A2(n39375), .Z(n32086) );
  XOR2_X1 U47043 ( .A1(n32086), .A2(n38653), .Z(n38555) );
  XOR2_X1 U47044 ( .A1(n32087), .A2(n38555), .Z(n46707) );
  XOR2_X1 U47045 ( .A1(n60207), .A2(n51290), .Z(n44913) );
  XOR2_X1 U47046 ( .A1(n46707), .A2(n44913), .Z(n32088) );
  XOR2_X1 U47047 ( .A1(n32089), .A2(n32088), .Z(n32090) );
  XOR2_X1 U47048 ( .A1(n32092), .A2(n32091), .Z(n32093) );
  XOR2_X1 U47049 ( .A1(n63955), .A2(n57096), .Z(n32094) );
  XOR2_X1 U47050 ( .A1(n23826), .A2(n32094), .Z(n33172) );
  XOR2_X1 U47051 ( .A1(n38009), .A2(n23020), .Z(n32096) );
  XOR2_X1 U47052 ( .A1(n38798), .A2(n32096), .Z(n44023) );
  XOR2_X1 U47053 ( .A1(n37897), .A2(n36998), .Z(n43770) );
  XOR2_X1 U47054 ( .A1(n43770), .A2(n55903), .Z(n32097) );
  XOR2_X1 U47055 ( .A1(n23389), .A2(n8329), .Z(n32100) );
  XOR2_X1 U47056 ( .A1(n30968), .A2(n44330), .Z(n37500) );
  XOR2_X1 U47057 ( .A1(n51150), .A2(n32472), .Z(n32102) );
  XOR2_X1 U47058 ( .A1(n37500), .A2(n32102), .Z(n43783) );
  INV_X1 U47059 ( .I(n32103), .ZN(n32104) );
  XOR2_X1 U47060 ( .A1(n32104), .A2(n55534), .Z(n52425) );
  XOR2_X1 U47061 ( .A1(n52425), .A2(n44739), .Z(n44030) );
  XOR2_X1 U47062 ( .A1(n43783), .A2(n44030), .Z(n32105) );
  INV_X1 U47063 ( .I(n33291), .ZN(n32108) );
  XOR2_X1 U47064 ( .A1(n32109), .A2(n32108), .Z(n32110) );
  XOR2_X1 U47065 ( .A1(n23714), .A2(n33243), .Z(n32111) );
  XOR2_X1 U47066 ( .A1(n32111), .A2(n33193), .Z(n32117) );
  INV_X1 U47067 ( .I(n44796), .ZN(n49955) );
  XOR2_X1 U47068 ( .A1(n37257), .A2(n49955), .Z(n32583) );
  XOR2_X1 U47069 ( .A1(n32112), .A2(n39228), .Z(n44876) );
  XOR2_X1 U47070 ( .A1(n51531), .A2(n55580), .Z(n32113) );
  XOR2_X1 U47071 ( .A1(n32113), .A2(n52178), .Z(n46647) );
  XOR2_X1 U47072 ( .A1(n44876), .A2(n46647), .Z(n32114) );
  XOR2_X1 U47073 ( .A1(n32661), .A2(n32115), .Z(n32116) );
  XOR2_X1 U47074 ( .A1(n32119), .A2(n32118), .Z(n32120) );
  XOR2_X1 U47075 ( .A1(n32122), .A2(n32590), .Z(n33191) );
  NAND2_X1 U47076 ( .A1(n33920), .A2(n34422), .ZN(n32137) );
  XOR2_X1 U47078 ( .A1(n32123), .A2(n53487), .Z(n33055) );
  INV_X1 U47079 ( .I(n44014), .ZN(n32124) );
  XOR2_X1 U47080 ( .A1(n33055), .A2(n32124), .Z(n32612) );
  INV_X1 U47081 ( .I(n32612), .ZN(n32125) );
  XOR2_X1 U47082 ( .A1(n38154), .A2(n55349), .Z(n39295) );
  XOR2_X1 U47083 ( .A1(n32125), .A2(n39295), .Z(n44718) );
  XOR2_X1 U47084 ( .A1(n37565), .A2(n30908), .Z(n32126) );
  XOR2_X1 U47085 ( .A1(n32126), .A2(n37704), .Z(n41738) );
  INV_X1 U47086 ( .I(n51999), .ZN(n51016) );
  XOR2_X1 U47087 ( .A1(n51016), .A2(n39570), .Z(n44715) );
  XOR2_X1 U47088 ( .A1(n41738), .A2(n44715), .Z(n32127) );
  XOR2_X1 U47089 ( .A1(n44718), .A2(n32127), .Z(n32128) );
  NAND3_X1 U47091 ( .A1(n33925), .A2(n34423), .A3(n1423), .ZN(n32134) );
  INV_X1 U47092 ( .I(n35769), .ZN(n32138) );
  AOI21_X1 U47093 ( .A1(n32139), .A2(n64984), .B(n32138), .ZN(n32140) );
  INV_X1 U47094 ( .I(n37190), .ZN(n32143) );
  NAND3_X1 U47096 ( .A1(n37334), .A2(n37329), .A3(n37333), .ZN(n32145) );
  OAI22_X1 U47099 ( .A1(n37005), .A2(n32154), .B1(n32153), .B2(n61574), .ZN(
        n32155) );
  XOR2_X1 U47100 ( .A1(n50129), .A2(n45275), .Z(n51680) );
  XOR2_X1 U47101 ( .A1(n44378), .A2(n24046), .Z(n46682) );
  XOR2_X1 U47102 ( .A1(n46682), .A2(n27640), .Z(n32302) );
  INV_X1 U47103 ( .I(n32302), .ZN(n32160) );
  XOR2_X1 U47104 ( .A1(n45404), .A2(n53272), .Z(n39725) );
  XOR2_X1 U47105 ( .A1(n55139), .A2(n23886), .Z(n44212) );
  XOR2_X1 U47106 ( .A1(n39725), .A2(n44212), .Z(n32159) );
  XOR2_X1 U47107 ( .A1(n32160), .A2(n32159), .Z(n32161) );
  XOR2_X1 U47108 ( .A1(n32166), .A2(n32165), .Z(n32171) );
  INV_X1 U47109 ( .I(n38772), .ZN(n32167) );
  XOR2_X1 U47110 ( .A1(n32168), .A2(n57142), .Z(n50770) );
  XOR2_X1 U47111 ( .A1(n45121), .A2(n9871), .Z(n32169) );
  XOR2_X1 U47112 ( .A1(n50770), .A2(n32169), .Z(n45286) );
  XOR2_X1 U47113 ( .A1(n56905), .A2(n54870), .Z(n50634) );
  XOR2_X1 U47114 ( .A1(n32172), .A2(n37758), .Z(n36145) );
  XOR2_X1 U47115 ( .A1(n36145), .A2(n44995), .Z(n45257) );
  XOR2_X1 U47116 ( .A1(n39704), .A2(n51494), .Z(n44170) );
  XOR2_X1 U47117 ( .A1(n44170), .A2(n57096), .Z(n32173) );
  XOR2_X1 U47118 ( .A1(n45257), .A2(n32173), .Z(n32174) );
  XOR2_X1 U47119 ( .A1(n23794), .A2(n32174), .Z(n32175) );
  XOR2_X1 U47120 ( .A1(n52375), .A2(n57162), .Z(n45087) );
  XOR2_X1 U47121 ( .A1(n45087), .A2(n54936), .Z(n32177) );
  XOR2_X1 U47122 ( .A1(n39400), .A2(n32177), .Z(n46111) );
  XOR2_X1 U47123 ( .A1(n32274), .A2(n56976), .Z(n38327) );
  XOR2_X1 U47124 ( .A1(n32178), .A2(n38327), .Z(n44950) );
  XOR2_X1 U47125 ( .A1(n44950), .A2(n54208), .Z(n32179) );
  XOR2_X1 U47126 ( .A1(n46111), .A2(n32179), .Z(n32180) );
  XOR2_X1 U47127 ( .A1(n32181), .A2(n32180), .Z(n32182) );
  XOR2_X1 U47128 ( .A1(n10378), .A2(n24008), .Z(n32378) );
  INV_X1 U47129 ( .I(n32355), .ZN(n32185) );
  XOR2_X1 U47131 ( .A1(n22390), .A2(n32393), .Z(n32187) );
  XOR2_X1 U47132 ( .A1(n38734), .A2(n32189), .Z(n51514) );
  XOR2_X1 U47133 ( .A1(n24011), .A2(n55060), .Z(n32190) );
  XOR2_X1 U47134 ( .A1(n51514), .A2(n32190), .Z(n45025) );
  XOR2_X1 U47135 ( .A1(n45025), .A2(n44014), .Z(n32191) );
  XOR2_X1 U47136 ( .A1(n53487), .A2(n56771), .Z(n38224) );
  XOR2_X1 U47137 ( .A1(n29969), .A2(n38224), .Z(n39219) );
  XOR2_X1 U47138 ( .A1(n39387), .A2(n39219), .Z(n46390) );
  XOR2_X1 U47139 ( .A1(n32191), .A2(n46390), .Z(n32192) );
  MUX2_X1 U47141 ( .I0(n33489), .I1(n10016), .S(n7116), .Z(n32211) );
  XOR2_X1 U47142 ( .A1(n32637), .A2(n32200), .Z(n32205) );
  XOR2_X1 U47143 ( .A1(n44163), .A2(n51667), .Z(n52594) );
  XOR2_X1 U47144 ( .A1(n52080), .A2(n54708), .Z(n39442) );
  XOR2_X1 U47145 ( .A1(n39442), .A2(n37729), .Z(n46130) );
  XOR2_X1 U47146 ( .A1(n52594), .A2(n46130), .Z(n32201) );
  XOR2_X1 U47147 ( .A1(n32202), .A2(n32203), .Z(n32204) );
  NOR3_X1 U47148 ( .A1(n3325), .A2(n63319), .A3(n34776), .ZN(n32214) );
  OAI22_X1 U47149 ( .A1(n33494), .A2(n33774), .B1(n61256), .B2(n19894), .ZN(
        n32213) );
  NOR3_X1 U47150 ( .A1(n34275), .A2(n15927), .A3(n34777), .ZN(n32212) );
  NAND2_X2 U47151 ( .A1(n32216), .A2(n32215), .ZN(n36451) );
  OAI21_X1 U47152 ( .A1(n35294), .A2(n21056), .B(n34335), .ZN(n32217) );
  NAND3_X1 U47153 ( .A1(n32217), .A2(n22278), .A3(n35301), .ZN(n32220) );
  XOR2_X1 U47154 ( .A1(n27640), .A2(n53090), .Z(n32223) );
  XOR2_X1 U47155 ( .A1(n24051), .A2(n55139), .Z(n37486) );
  XOR2_X1 U47156 ( .A1(n32223), .A2(n37486), .Z(n44761) );
  XOR2_X1 U47157 ( .A1(n44761), .A2(n32224), .Z(n40458) );
  XOR2_X1 U47159 ( .A1(n50733), .A2(n56784), .Z(n45112) );
  XOR2_X1 U47161 ( .A1(n38556), .A2(n54676), .Z(n37757) );
  XOR2_X1 U47162 ( .A1(n39707), .A2(n37757), .Z(n32231) );
  XOR2_X1 U47163 ( .A1(n32231), .A2(n22458), .Z(n43808) );
  XOR2_X1 U47164 ( .A1(n238), .A2(n51492), .Z(n44054) );
  XOR2_X1 U47165 ( .A1(n43808), .A2(n44054), .Z(n32233) );
  XOR2_X1 U47166 ( .A1(n60565), .A2(n32233), .Z(n32235) );
  INV_X1 U47168 ( .I(n32242), .ZN(n32243) );
  INV_X1 U47169 ( .I(n32563), .ZN(n32248) );
  XOR2_X1 U47170 ( .A1(n38459), .A2(n32249), .Z(n38638) );
  XOR2_X1 U47171 ( .A1(n38638), .A2(n54888), .Z(n38720) );
  XOR2_X1 U47172 ( .A1(n38639), .A2(n23306), .Z(n50534) );
  XOR2_X1 U47173 ( .A1(n38720), .A2(n50534), .Z(n44887) );
  INV_X1 U47174 ( .I(n39442), .ZN(n32250) );
  XOR2_X1 U47175 ( .A1(n32250), .A2(n54376), .Z(n50855) );
  XOR2_X1 U47176 ( .A1(n50855), .A2(n32251), .Z(n46660) );
  XOR2_X1 U47177 ( .A1(n46660), .A2(n56849), .Z(n32252) );
  XOR2_X1 U47178 ( .A1(n44887), .A2(n32252), .Z(n32253) );
  XOR2_X1 U47180 ( .A1(n32255), .A2(n887), .Z(n32259) );
  XOR2_X1 U47181 ( .A1(n61304), .A2(n9636), .Z(n32257) );
  XOR2_X1 U47182 ( .A1(n32257), .A2(n32256), .Z(n32258) );
  XOR2_X1 U47183 ( .A1(n32259), .A2(n32258), .Z(n32260) );
  XOR2_X1 U47185 ( .A1(n51530), .A2(n53102), .Z(n44323) );
  INV_X1 U47186 ( .I(n44323), .ZN(n37499) );
  XOR2_X1 U47187 ( .A1(n32263), .A2(n37499), .Z(n44345) );
  XOR2_X1 U47188 ( .A1(n247), .A2(n30402), .Z(n44041) );
  XOR2_X1 U47189 ( .A1(n57142), .A2(n56879), .Z(n37259) );
  XOR2_X1 U47190 ( .A1(n55087), .A2(n9871), .Z(n50453) );
  XOR2_X1 U47191 ( .A1(n37259), .A2(n50453), .Z(n43789) );
  XOR2_X1 U47192 ( .A1(n50682), .A2(n54407), .Z(n43788) );
  XOR2_X1 U47193 ( .A1(n43789), .A2(n43788), .Z(n32264) );
  XOR2_X1 U47194 ( .A1(n44041), .A2(n32264), .Z(n32265) );
  XOR2_X1 U47195 ( .A1(n32266), .A2(n32265), .Z(n32268) );
  XOR2_X1 U47196 ( .A1(n45371), .A2(n56901), .Z(n46488) );
  XOR2_X1 U47197 ( .A1(n46488), .A2(n55106), .Z(n32349) );
  XOR2_X1 U47198 ( .A1(n23789), .A2(n39457), .Z(n32272) );
  XOR2_X1 U47199 ( .A1(n32349), .A2(n32272), .Z(n46671) );
  XOR2_X1 U47200 ( .A1(n53530), .A2(n54587), .Z(n32273) );
  XOR2_X1 U47201 ( .A1(n50698), .A2(n32273), .Z(n32275) );
  XOR2_X1 U47202 ( .A1(n38450), .A2(n32274), .Z(n44924) );
  XOR2_X1 U47203 ( .A1(n32275), .A2(n44924), .Z(n32276) );
  XOR2_X1 U47205 ( .A1(n38000), .A2(n32286), .Z(n44589) );
  XOR2_X1 U47206 ( .A1(n44589), .A2(n38829), .Z(n32287) );
  XOR2_X1 U47207 ( .A1(n32287), .A2(n59680), .Z(n32288) );
  XOR2_X1 U47208 ( .A1(n22390), .A2(n32288), .Z(n32290) );
  XOR2_X1 U47210 ( .A1(n32302), .A2(n44108), .Z(n32303) );
  XOR2_X1 U47211 ( .A1(n39538), .A2(n53154), .Z(n51235) );
  XOR2_X1 U47212 ( .A1(n51235), .A2(n52029), .Z(n43588) );
  XOR2_X1 U47213 ( .A1(n32305), .A2(n32304), .Z(n32306) );
  XOR2_X1 U47214 ( .A1(n39478), .A2(n50634), .Z(n37881) );
  XOR2_X1 U47215 ( .A1(n37881), .A2(n50832), .Z(n32309) );
  XOR2_X1 U47216 ( .A1(n36147), .A2(n32309), .Z(n44365) );
  XOR2_X1 U47217 ( .A1(n32410), .A2(n32310), .Z(n39376) );
  XOR2_X1 U47218 ( .A1(n39376), .A2(n1887), .Z(n43641) );
  XOR2_X1 U47219 ( .A1(n43641), .A2(n54360), .Z(n32311) );
  XOR2_X1 U47220 ( .A1(n44365), .A2(n32311), .Z(n32312) );
  XOR2_X1 U47221 ( .A1(n32314), .A2(n32313), .Z(n32316) );
  XOR2_X1 U47222 ( .A1(n32317), .A2(n22820), .Z(n32319) );
  XOR2_X1 U47223 ( .A1(n32319), .A2(n20862), .Z(n32320) );
  XOR2_X1 U47224 ( .A1(n64355), .A2(n52196), .Z(n39443) );
  XOR2_X1 U47225 ( .A1(n39443), .A2(n46130), .Z(n46514) );
  XOR2_X1 U47226 ( .A1(n45131), .A2(n46128), .Z(n32322) );
  XOR2_X1 U47227 ( .A1(n46514), .A2(n32322), .Z(n32323) );
  XOR2_X1 U47228 ( .A1(n9283), .A2(n32323), .Z(n32325) );
  XOR2_X1 U47229 ( .A1(n23424), .A2(n32326), .Z(n33874) );
  XOR2_X1 U47230 ( .A1(n33874), .A2(n32328), .Z(n32329) );
  XOR2_X1 U47231 ( .A1(n20810), .A2(n32329), .Z(n32330) );
  XOR2_X1 U47232 ( .A1(n57142), .A2(n56335), .Z(n33900) );
  XOR2_X1 U47233 ( .A1(n37993), .A2(n33900), .Z(n43670) );
  XOR2_X1 U47234 ( .A1(n38472), .A2(n55889), .Z(n32333) );
  XOR2_X1 U47235 ( .A1(n43670), .A2(n32333), .Z(n32334) );
  XOR2_X1 U47236 ( .A1(n32335), .A2(n32334), .Z(n32337) );
  XOR2_X1 U47237 ( .A1(n32337), .A2(n32336), .Z(n32340) );
  XOR2_X1 U47238 ( .A1(n23786), .A2(n32338), .Z(n33909) );
  XOR2_X1 U47239 ( .A1(n33909), .A2(n32340), .Z(n32341) );
  XOR2_X1 U47240 ( .A1(n37889), .A2(n55196), .Z(n32549) );
  XOR2_X1 U47241 ( .A1(n39568), .A2(n32549), .Z(n44436) );
  XOR2_X1 U47242 ( .A1(n32344), .A2(n53262), .Z(n38588) );
  XOR2_X1 U47243 ( .A1(n53076), .A2(n54896), .Z(n38109) );
  XOR2_X1 U47244 ( .A1(n38588), .A2(n38109), .Z(n46583) );
  XOR2_X1 U47245 ( .A1(n44436), .A2(n46583), .Z(n32345) );
  XOR2_X1 U47247 ( .A1(n32349), .A2(n54776), .Z(n51132) );
  XOR2_X1 U47248 ( .A1(n51132), .A2(n61550), .Z(n32351) );
  XOR2_X1 U47249 ( .A1(n39280), .A2(n38327), .Z(n38162) );
  XOR2_X1 U47250 ( .A1(n1190), .A2(n23999), .Z(n39279) );
  XOR2_X1 U47251 ( .A1(n39279), .A2(n37713), .Z(n32350) );
  XOR2_X1 U47252 ( .A1(n38162), .A2(n32350), .Z(n45091) );
  XOR2_X1 U47253 ( .A1(n32351), .A2(n45091), .Z(n32352) );
  NAND2_X1 U47254 ( .A1(n34791), .A2(n61262), .ZN(n32360) );
  NOR2_X1 U47255 ( .A1(n60415), .A2(n9648), .ZN(n32359) );
  NAND2_X1 U47258 ( .A1(n64753), .A2(n36456), .ZN(n35164) );
  INV_X1 U47259 ( .I(n35164), .ZN(n32442) );
  XOR2_X1 U47260 ( .A1(n32364), .A2(n245), .Z(n50741) );
  XOR2_X1 U47261 ( .A1(n22323), .A2(n38625), .Z(n51926) );
  XOR2_X1 U47262 ( .A1(n24046), .A2(n54168), .Z(n32365) );
  XOR2_X1 U47263 ( .A1(n51926), .A2(n32365), .Z(n43798) );
  XOR2_X1 U47264 ( .A1(n43798), .A2(n57131), .Z(n32366) );
  XOR2_X1 U47265 ( .A1(n50741), .A2(n32366), .Z(n32367) );
  INV_X1 U47266 ( .I(n46114), .ZN(n32373) );
  XOR2_X1 U47267 ( .A1(n39458), .A2(n54289), .Z(n32372) );
  XOR2_X1 U47268 ( .A1(n32373), .A2(n32372), .Z(n32374) );
  XOR2_X1 U47269 ( .A1(n32374), .A2(n38378), .Z(n44822) );
  XOR2_X1 U47270 ( .A1(n44533), .A2(n56901), .Z(n46273) );
  XOR2_X1 U47271 ( .A1(n44822), .A2(n46273), .Z(n32375) );
  XOR2_X1 U47272 ( .A1(n32375), .A2(n33891), .Z(n32376) );
  XOR2_X1 U47273 ( .A1(n4278), .A2(n32378), .Z(n32379) );
  XOR2_X1 U47274 ( .A1(n49088), .A2(n44323), .Z(n32381) );
  XOR2_X1 U47275 ( .A1(n32382), .A2(n32381), .Z(n32384) );
  XOR2_X1 U47276 ( .A1(n32384), .A2(n23714), .Z(n32385) );
  XOR2_X1 U47277 ( .A1(n32389), .A2(n1827), .Z(n32390) );
  INV_X1 U47278 ( .I(n32394), .ZN(n32395) );
  XOR2_X1 U47279 ( .A1(n32397), .A2(n38588), .Z(n46698) );
  XOR2_X1 U47280 ( .A1(n44932), .A2(n46698), .Z(n32398) );
  XOR2_X1 U47281 ( .A1(n30036), .A2(n32401), .Z(n51766) );
  XOR2_X1 U47282 ( .A1(n51766), .A2(n52197), .Z(n44803) );
  XOR2_X1 U47283 ( .A1(n46324), .A2(n44803), .Z(n32402) );
  AOI22_X1 U47284 ( .A1(n15181), .A2(n34247), .B1(n4591), .B2(n34353), .ZN(
        n32423) );
  XOR2_X1 U47285 ( .A1(n38997), .A2(n32410), .Z(n45418) );
  XOR2_X1 U47286 ( .A1(n45418), .A2(n51493), .Z(n32411) );
  XOR2_X1 U47287 ( .A1(n32412), .A2(n32411), .Z(n32413) );
  XOR2_X1 U47288 ( .A1(n38896), .A2(n35523), .Z(n32415) );
  XOR2_X1 U47289 ( .A1(n32416), .A2(n32415), .Z(n44299) );
  XOR2_X1 U47290 ( .A1(n44299), .A2(n56008), .Z(n50764) );
  XOR2_X1 U47291 ( .A1(n50764), .A2(n33857), .Z(n32417) );
  NAND2_X1 U47293 ( .A1(n15184), .A2(n34727), .ZN(n32427) );
  NAND2_X1 U47294 ( .A1(n493), .A2(n34719), .ZN(n32927) );
  INV_X1 U47295 ( .I(n32430), .ZN(n34302) );
  NAND2_X1 U47296 ( .A1(n60970), .A2(n34309), .ZN(n32431) );
  INV_X1 U47298 ( .I(n60970), .ZN(n34219) );
  NAND2_X1 U47299 ( .A1(n32435), .A2(n60970), .ZN(n32437) );
  NOR2_X1 U47300 ( .A1(n36443), .A2(n1419), .ZN(n35592) );
  NOR2_X1 U47301 ( .A1(n60562), .A2(n36224), .ZN(n32439) );
  NOR2_X1 U47302 ( .A1(n35592), .A2(n32439), .ZN(n35163) );
  NOR2_X1 U47303 ( .A1(n32440), .A2(n35598), .ZN(n32441) );
  NOR2_X1 U47304 ( .A1(n1531), .A2(n60562), .ZN(n32445) );
  INV_X1 U47305 ( .I(n35588), .ZN(n32443) );
  NOR2_X1 U47306 ( .A1(n32443), .A2(n9633), .ZN(n32444) );
  NOR3_X1 U47307 ( .A1(n1792), .A2(n60562), .A3(n9633), .ZN(n32446) );
  OAI21_X1 U47308 ( .A1(n57171), .A2(n32446), .B(n36449), .ZN(n32449) );
  INV_X1 U47309 ( .I(n36449), .ZN(n32447) );
  NAND3_X1 U47310 ( .A1(n32447), .A2(n1419), .A3(n36437), .ZN(n32448) );
  OAI22_X1 U47311 ( .A1(n33616), .A2(n32460), .B1(n7311), .B2(n33405), .ZN(
        n32455) );
  NOR2_X1 U47312 ( .A1(n32456), .A2(n32455), .ZN(n32466) );
  NOR2_X1 U47313 ( .A1(n65256), .A2(n1542), .ZN(n32462) );
  INV_X1 U47314 ( .I(n32784), .ZN(n33000) );
  XOR2_X1 U47315 ( .A1(n32467), .A2(n52317), .Z(n32469) );
  XOR2_X1 U47316 ( .A1(n32469), .A2(n32468), .Z(n32645) );
  XOR2_X1 U47317 ( .A1(n33176), .A2(n32470), .Z(n32471) );
  XOR2_X1 U47318 ( .A1(n32472), .A2(n39631), .Z(n33279) );
  XOR2_X1 U47319 ( .A1(n33279), .A2(n30036), .Z(n46515) );
  XOR2_X1 U47320 ( .A1(n45130), .A2(n46515), .Z(n32473) );
  XOR2_X1 U47321 ( .A1(n32473), .A2(n44967), .Z(n32474) );
  XOR2_X1 U47322 ( .A1(n1825), .A2(n32474), .Z(n32476) );
  XOR2_X1 U47325 ( .A1(n38650), .A2(n38995), .Z(n37464) );
  XOR2_X1 U47326 ( .A1(n37464), .A2(n37303), .Z(n43645) );
  XOR2_X1 U47327 ( .A1(n39376), .A2(n38653), .Z(n44363) );
  XOR2_X1 U47328 ( .A1(n44363), .A2(n55118), .Z(n32481) );
  XOR2_X1 U47329 ( .A1(n43645), .A2(n32481), .Z(n32482) );
  XOR2_X1 U47330 ( .A1(n20862), .A2(n32482), .Z(n32484) );
  XOR2_X1 U47331 ( .A1(n32667), .A2(n32484), .Z(n32485) );
  XOR2_X1 U47332 ( .A1(n32488), .A2(n32487), .Z(n32489) );
  NAND2_X1 U47333 ( .A1(n33103), .A2(n33561), .ZN(n33694) );
  INV_X1 U47334 ( .I(n38074), .ZN(n32490) );
  XOR2_X1 U47335 ( .A1(n32490), .A2(n50504), .Z(n37748) );
  XOR2_X1 U47336 ( .A1(n38880), .A2(n24046), .Z(n50128) );
  XOR2_X1 U47337 ( .A1(n50128), .A2(n43968), .Z(n32491) );
  XOR2_X1 U47338 ( .A1(n37748), .A2(n32491), .Z(n43587) );
  XOR2_X1 U47339 ( .A1(n43587), .A2(n44107), .Z(n32492) );
  NAND2_X1 U47341 ( .A1(n33694), .A2(n63624), .ZN(n32511) );
  XOR2_X1 U47342 ( .A1(n32500), .A2(n49289), .Z(n46486) );
  XOR2_X1 U47343 ( .A1(n58077), .A2(n56901), .Z(n32501) );
  XOR2_X1 U47344 ( .A1(n45087), .A2(n32501), .Z(n32502) );
  XOR2_X1 U47345 ( .A1(n46486), .A2(n32502), .Z(n32503) );
  XOR2_X1 U47346 ( .A1(n45379), .A2(n53958), .Z(n32506) );
  XOR2_X1 U47347 ( .A1(n32546), .A2(n32506), .Z(n44437) );
  XOR2_X1 U47348 ( .A1(n44437), .A2(n54386), .Z(n32507) );
  INV_X1 U47350 ( .I(n33348), .ZN(n32526) );
  XOR2_X1 U47352 ( .A1(n32519), .A2(n54185), .Z(n49897) );
  XOR2_X1 U47353 ( .A1(n51216), .A2(n55087), .Z(n50646) );
  XOR2_X1 U47354 ( .A1(n49897), .A2(n50646), .Z(n44346) );
  XOR2_X1 U47355 ( .A1(n44796), .A2(n37637), .Z(n43667) );
  XOR2_X1 U47356 ( .A1(n43667), .A2(n54917), .Z(n32520) );
  XOR2_X1 U47357 ( .A1(n44346), .A2(n32520), .Z(n32521) );
  NAND2_X1 U47359 ( .A1(n32530), .A2(n32814), .ZN(n32534) );
  NOR2_X1 U47360 ( .A1(n33097), .A2(n63064), .ZN(n32532) );
  XOR2_X1 U47361 ( .A1(n56819), .A2(n56976), .Z(n32536) );
  XOR2_X1 U47362 ( .A1(n33062), .A2(n32536), .Z(n46669) );
  XOR2_X1 U47363 ( .A1(n46669), .A2(n45087), .Z(n32538) );
  XOR2_X1 U47364 ( .A1(n32538), .A2(n32537), .Z(n32539) );
  XOR2_X1 U47366 ( .A1(n32546), .A2(n36319), .Z(n32548) );
  XOR2_X1 U47367 ( .A1(n29969), .A2(n54231), .Z(n51729) );
  XOR2_X1 U47368 ( .A1(n51729), .A2(n38154), .Z(n32547) );
  XOR2_X1 U47369 ( .A1(n32548), .A2(n32547), .Z(n44588) );
  XOR2_X1 U47370 ( .A1(n32549), .A2(n56859), .Z(n32550) );
  XOR2_X1 U47371 ( .A1(n51379), .A2(n55060), .Z(n39667) );
  XOR2_X1 U47372 ( .A1(n32550), .A2(n39667), .Z(n45879) );
  XOR2_X1 U47373 ( .A1(n44588), .A2(n45879), .Z(n32551) );
  XOR2_X1 U47374 ( .A1(n32553), .A2(n32552), .Z(n32554) );
  XOR2_X1 U47375 ( .A1(n32558), .A2(n56683), .Z(n36630) );
  XOR2_X1 U47376 ( .A1(n36630), .A2(n54708), .Z(n36929) );
  XOR2_X1 U47377 ( .A1(n36929), .A2(n55534), .Z(n44888) );
  XOR2_X1 U47378 ( .A1(n37981), .A2(n33279), .Z(n46659) );
  XOR2_X1 U47379 ( .A1(n44888), .A2(n46659), .Z(n32559) );
  XOR2_X1 U47380 ( .A1(n9636), .A2(n32559), .Z(n32561) );
  XOR2_X1 U47381 ( .A1(n44841), .A2(n56322), .Z(n32566) );
  XOR2_X1 U47382 ( .A1(n32566), .A2(n49448), .Z(n44758) );
  XOR2_X1 U47383 ( .A1(n44758), .A2(n54556), .Z(n51740) );
  XOR2_X1 U47384 ( .A1(n44761), .A2(n55368), .Z(n50726) );
  XOR2_X1 U47385 ( .A1(n50726), .A2(n22773), .Z(n32567) );
  XOR2_X1 U47386 ( .A1(n51740), .A2(n32567), .Z(n32569) );
  XOR2_X1 U47387 ( .A1(n32569), .A2(n32568), .Z(n32570) );
  XOR2_X1 U47388 ( .A1(n38280), .A2(n56827), .Z(n32575) );
  XOR2_X1 U47389 ( .A1(n32575), .A2(n38555), .Z(n44056) );
  XOR2_X1 U47390 ( .A1(n24105), .A2(n51492), .Z(n37585) );
  XOR2_X1 U47391 ( .A1(n37585), .A2(n54517), .Z(n32576) );
  XOR2_X1 U47392 ( .A1(n32576), .A2(n33165), .Z(n43809) );
  XOR2_X1 U47393 ( .A1(n43809), .A2(n53772), .Z(n32577) );
  XOR2_X1 U47394 ( .A1(n44056), .A2(n32577), .Z(n32578) );
  INV_X1 U47395 ( .I(n727), .ZN(n32579) );
  XOR2_X1 U47396 ( .A1(n32580), .A2(n32579), .Z(n32581) );
  XOR2_X1 U47397 ( .A1(n32583), .A2(n50551), .Z(n52463) );
  XOR2_X1 U47398 ( .A1(n52463), .A2(n38631), .Z(n43787) );
  XOR2_X1 U47399 ( .A1(n51216), .A2(n56714), .Z(n33071) );
  XOR2_X1 U47400 ( .A1(n43789), .A2(n33071), .Z(n44040) );
  XOR2_X1 U47401 ( .A1(n43787), .A2(n44040), .Z(n32584) );
  XOR2_X1 U47402 ( .A1(n32584), .A2(n22583), .Z(n32586) );
  XOR2_X1 U47403 ( .A1(n32585), .A2(n32586), .Z(n32589) );
  XOR2_X1 U47404 ( .A1(n32591), .A2(n32590), .Z(n32593) );
  XOR2_X1 U47405 ( .A1(n32593), .A2(n32592), .Z(n32594) );
  AOI21_X1 U47406 ( .A1(n33117), .A2(n33644), .B(n32599), .ZN(n32609) );
  NOR2_X1 U47407 ( .A1(n60434), .A2(n33539), .ZN(n32600) );
  AOI22_X1 U47408 ( .A1(n33536), .A2(n33644), .B1(n33630), .B2(n32600), .ZN(
        n32608) );
  AOI22_X1 U47411 ( .A1(n33627), .A2(n33220), .B1(n33112), .B2(n33537), .ZN(
        n32602) );
  NAND2_X1 U47412 ( .A1(n13942), .A2(n25428), .ZN(n33533) );
  OAI21_X1 U47413 ( .A1(n33375), .A2(n33533), .B(n33374), .ZN(n32605) );
  NAND3_X1 U47414 ( .A1(n32605), .A2(n33539), .A3(n60434), .ZN(n32606) );
  INV_X1 U47415 ( .I(n35159), .ZN(n32692) );
  XOR2_X1 U47416 ( .A1(n32612), .A2(n39488), .Z(n33878) );
  XOR2_X1 U47417 ( .A1(n33878), .A2(n53958), .Z(n38732) );
  XOR2_X1 U47418 ( .A1(n33147), .A2(n53138), .Z(n32613) );
  XOR2_X1 U47419 ( .A1(n45238), .A2(n55060), .Z(n33056) );
  XOR2_X1 U47420 ( .A1(n32613), .A2(n33056), .Z(n45380) );
  XOR2_X1 U47421 ( .A1(n38732), .A2(n45380), .Z(n32614) );
  XOR2_X1 U47422 ( .A1(n1832), .A2(n32617), .Z(n32618) );
  XOR2_X1 U47423 ( .A1(n38326), .A2(n56819), .Z(n51915) );
  XOR2_X1 U47424 ( .A1(n32621), .A2(n55395), .Z(n32622) );
  XOR2_X1 U47425 ( .A1(n51915), .A2(n32622), .Z(n46571) );
  XOR2_X1 U47426 ( .A1(n51193), .A2(n56901), .Z(n44461) );
  XOR2_X1 U47427 ( .A1(n23020), .A2(n44461), .Z(n32624) );
  XOR2_X1 U47428 ( .A1(n37896), .A2(n61550), .Z(n32623) );
  XOR2_X1 U47429 ( .A1(n32624), .A2(n32623), .Z(n32625) );
  XOR2_X1 U47430 ( .A1(n46571), .A2(n32625), .Z(n32626) );
  XOR2_X1 U47431 ( .A1(n23950), .A2(n32626), .Z(n32627) );
  XOR2_X1 U47432 ( .A1(n1834), .A2(n32628), .Z(n32629) );
  INV_X1 U47433 ( .I(n38430), .ZN(n50621) );
  XOR2_X1 U47435 ( .A1(n46396), .A2(n52551), .Z(n37973) );
  XOR2_X1 U47436 ( .A1(n50504), .A2(n54556), .Z(n33024) );
  XOR2_X1 U47437 ( .A1(n33024), .A2(n56784), .Z(n50628) );
  XOR2_X1 U47438 ( .A1(n50628), .A2(n39363), .Z(n44844) );
  XOR2_X1 U47439 ( .A1(n44844), .A2(n44109), .Z(n32630) );
  XOR2_X1 U47440 ( .A1(n37973), .A2(n32630), .Z(n32631) );
  XOR2_X1 U47441 ( .A1(n32632), .A2(n32631), .Z(n32633) );
  XOR2_X1 U47443 ( .A1(n33871), .A2(n44427), .Z(n37808) );
  XOR2_X1 U47444 ( .A1(n61737), .A2(n53787), .Z(n32639) );
  XOR2_X1 U47445 ( .A1(n37808), .A2(n32639), .Z(n32641) );
  XOR2_X1 U47446 ( .A1(n32641), .A2(n32640), .Z(n32644) );
  INV_X1 U47447 ( .I(n32642), .ZN(n32643) );
  XOR2_X1 U47448 ( .A1(n32644), .A2(n32643), .Z(n32646) );
  XOR2_X1 U47449 ( .A1(n32658), .A2(n37638), .Z(n37255) );
  XOR2_X1 U47450 ( .A1(n33899), .A2(n37255), .Z(n43263) );
  XOR2_X1 U47451 ( .A1(n9722), .A2(n52178), .Z(n37497) );
  XOR2_X1 U47452 ( .A1(n37497), .A2(n9871), .Z(n44099) );
  XOR2_X1 U47453 ( .A1(n44099), .A2(n54563), .Z(n32659) );
  XOR2_X1 U47454 ( .A1(n43263), .A2(n32659), .Z(n32660) );
  XOR2_X1 U47455 ( .A1(n32661), .A2(n32662), .Z(n32664) );
  XOR2_X1 U47456 ( .A1(n22583), .A2(n32663), .Z(n33194) );
  XOR2_X1 U47457 ( .A1(n32670), .A2(n37757), .Z(n44124) );
  XOR2_X1 U47458 ( .A1(n39530), .A2(n24105), .Z(n52565) );
  XOR2_X1 U47459 ( .A1(n52565), .A2(n54517), .Z(n32671) );
  XOR2_X1 U47460 ( .A1(n38388), .A2(n51881), .Z(n45470) );
  XOR2_X1 U47461 ( .A1(n32671), .A2(n45470), .Z(n43399) );
  XOR2_X1 U47462 ( .A1(n44124), .A2(n43399), .Z(n32672) );
  XOR2_X1 U47463 ( .A1(n32673), .A2(n32672), .Z(n32674) );
  OAI22_X1 U47464 ( .A1(n33316), .A2(n32678), .B1(n35611), .B2(n32677), .ZN(
        n32679) );
  OAI21_X1 U47465 ( .A1(n8365), .A2(n32680), .B(n33550), .ZN(n32689) );
  NOR2_X1 U47466 ( .A1(n32681), .A2(n35630), .ZN(n32682) );
  AOI21_X1 U47467 ( .A1(n32993), .A2(n7342), .B(n32685), .ZN(n32686) );
  OAI21_X1 U47468 ( .A1(n35622), .A2(n35203), .B(n32686), .ZN(n32687) );
  NAND2_X1 U47470 ( .A1(n33396), .A2(n32694), .ZN(n32697) );
  AOI21_X1 U47471 ( .A1(n33649), .A2(n19416), .B(n22598), .ZN(n32696) );
  NAND3_X1 U47472 ( .A1(n34138), .A2(n34143), .A3(n33397), .ZN(n32702) );
  XOR2_X1 U47473 ( .A1(n32706), .A2(n55196), .Z(n45347) );
  XOR2_X1 U47474 ( .A1(n39488), .A2(n54896), .Z(n32707) );
  XOR2_X1 U47475 ( .A1(n50873), .A2(n32707), .Z(n44490) );
  XOR2_X1 U47476 ( .A1(n45347), .A2(n32708), .Z(n32709) );
  XOR2_X1 U47477 ( .A1(n32710), .A2(n32711), .Z(n32713) );
  XOR2_X1 U47478 ( .A1(n32712), .A2(n32713), .Z(n32714) );
  XOR2_X1 U47479 ( .A1(n9753), .A2(n31613), .Z(n52614) );
  XOR2_X1 U47480 ( .A1(n39538), .A2(n44378), .Z(n42814) );
  XOR2_X1 U47481 ( .A1(n42814), .A2(n50505), .Z(n32717) );
  XOR2_X1 U47482 ( .A1(n52614), .A2(n32717), .Z(n32718) );
  XOR2_X1 U47483 ( .A1(n45416), .A2(n38560), .Z(n50903) );
  XOR2_X1 U47484 ( .A1(n50903), .A2(n54870), .Z(n43937) );
  XOR2_X1 U47485 ( .A1(n39196), .A2(n54360), .Z(n38558) );
  XOR2_X1 U47486 ( .A1(n38558), .A2(n37757), .Z(n44240) );
  XOR2_X1 U47487 ( .A1(n44240), .A2(n50494), .Z(n32723) );
  XOR2_X1 U47489 ( .A1(n37691), .A2(n61737), .Z(n33179) );
  XOR2_X1 U47490 ( .A1(n33179), .A2(n56683), .Z(n45067) );
  XOR2_X1 U47491 ( .A1(n32729), .A2(n32728), .Z(n46415) );
  XOR2_X1 U47492 ( .A1(n50025), .A2(n55765), .Z(n32730) );
  XOR2_X1 U47493 ( .A1(n46415), .A2(n32730), .Z(n32731) );
  XOR2_X1 U47494 ( .A1(n45067), .A2(n32731), .Z(n32732) );
  XOR2_X1 U47495 ( .A1(n23465), .A2(n32736), .Z(n32737) );
  XOR2_X1 U47496 ( .A1(n32740), .A2(n50486), .Z(n36356) );
  XOR2_X1 U47497 ( .A1(n32741), .A2(n56819), .Z(n50924) );
  XOR2_X1 U47498 ( .A1(n36356), .A2(n50924), .Z(n52169) );
  XOR2_X1 U47499 ( .A1(n1190), .A2(n56976), .Z(n51194) );
  XOR2_X1 U47500 ( .A1(n52169), .A2(n51194), .Z(n32743) );
  XNOR2_X1 U47501 ( .A1(n56901), .A2(n56745), .ZN(n32742) );
  XOR2_X1 U47502 ( .A1(n39399), .A2(n32742), .Z(n45011) );
  XOR2_X1 U47503 ( .A1(n32745), .A2(n11529), .Z(n32746) );
  XOR2_X1 U47504 ( .A1(n38472), .A2(n54917), .Z(n51071) );
  XOR2_X1 U47505 ( .A1(n9722), .A2(n53833), .Z(n32750) );
  XOR2_X1 U47506 ( .A1(n59638), .A2(n32750), .Z(n32751) );
  XOR2_X1 U47507 ( .A1(n51071), .A2(n32751), .Z(n44271) );
  XOR2_X1 U47508 ( .A1(n44796), .A2(n54563), .Z(n38632) );
  XOR2_X1 U47509 ( .A1(n23929), .A2(n56508), .Z(n32752) );
  XOR2_X1 U47510 ( .A1(n38632), .A2(n32752), .Z(n43860) );
  XOR2_X1 U47511 ( .A1(n44271), .A2(n43860), .Z(n32753) );
  XOR2_X1 U47512 ( .A1(n33194), .A2(n32755), .Z(n32756) );
  XOR2_X1 U47513 ( .A1(n32757), .A2(n32756), .Z(n32758) );
  INV_X2 U47515 ( .I(n33336), .ZN(n33600) );
  NAND2_X1 U47516 ( .A1(n60456), .A2(n35688), .ZN(n32767) );
  NAND3_X1 U47518 ( .A1(n32770), .A2(n32769), .A3(n36485), .ZN(n32779) );
  INV_X1 U47519 ( .I(n35154), .ZN(n32771) );
  NAND2_X1 U47520 ( .A1(n36238), .A2(n36483), .ZN(n32773) );
  NOR3_X1 U47521 ( .A1(n35154), .A2(n35153), .A3(n22527), .ZN(n32776) );
  NOR2_X1 U47522 ( .A1(n34488), .A2(n32776), .ZN(n32777) );
  AOI21_X1 U47526 ( .A1(n32781), .A2(n64838), .B(n64417), .ZN(n32787) );
  NAND2_X1 U47528 ( .A1(n32784), .A2(n23127), .ZN(n32785) );
  NOR2_X1 U47532 ( .A1(n32796), .A2(n60892), .ZN(n32797) );
  NOR2_X1 U47533 ( .A1(n32798), .A2(n32797), .ZN(n32799) );
  AOI21_X1 U47534 ( .A1(n32800), .A2(n32799), .B(n34114), .ZN(n32801) );
  INV_X1 U47535 ( .I(n32802), .ZN(n32805) );
  NAND2_X1 U47536 ( .A1(n33097), .A2(n7273), .ZN(n32803) );
  NAND2_X1 U47538 ( .A1(n32807), .A2(n61483), .ZN(n32806) );
  NOR2_X1 U47539 ( .A1(n33349), .A2(n33342), .ZN(n32808) );
  NOR2_X1 U47541 ( .A1(n33564), .A2(n33559), .ZN(n32809) );
  NAND2_X1 U47545 ( .A1(n32820), .A2(n32819), .ZN(n32827) );
  NAND4_X1 U47546 ( .A1(n33652), .A2(n32821), .A3(n33654), .A4(n34132), .ZN(
        n32823) );
  NAND2_X1 U47550 ( .A1(n32891), .A2(n32834), .ZN(n33990) );
  NAND2_X1 U47551 ( .A1(n34197), .A2(n33990), .ZN(n32832) );
  NAND2_X1 U47552 ( .A1(n32835), .A2(n32834), .ZN(n32837) );
  NAND3_X1 U47553 ( .A1(n32899), .A2(n33670), .A3(n65052), .ZN(n32844) );
  INV_X1 U47554 ( .I(n33674), .ZN(n32843) );
  NAND2_X1 U47555 ( .A1(n32844), .A2(n32843), .ZN(n32854) );
  NOR2_X1 U47556 ( .A1(n59626), .A2(n32845), .ZN(n32847) );
  OAI21_X1 U47557 ( .A1(n61197), .A2(n34155), .B(n23757), .ZN(n32848) );
  NAND2_X1 U47558 ( .A1(n32848), .A2(n12412), .ZN(n32851) );
  NAND3_X1 U47559 ( .A1(n24287), .A2(n33685), .A3(n65052), .ZN(n32849) );
  INV_X1 U47564 ( .I(n35582), .ZN(n32858) );
  NOR2_X1 U47566 ( .A1(n34460), .A2(n63484), .ZN(n32860) );
  AOI21_X1 U47567 ( .A1(n32864), .A2(n62931), .B(n32862), .ZN(n32867) );
  NAND3_X1 U47568 ( .A1(n34116), .A2(n32870), .A3(n62931), .ZN(n32871) );
  NAND2_X2 U47569 ( .A1(n57165), .A2(n7453), .ZN(n33432) );
  NOR2_X1 U47570 ( .A1(n20835), .A2(n7453), .ZN(n34187) );
  NAND2_X1 U47572 ( .A1(n33966), .A2(n118), .ZN(n32879) );
  NOR2_X1 U47573 ( .A1(n32882), .A2(n34002), .ZN(n32883) );
  INV_X1 U47574 ( .I(n32900), .ZN(n32896) );
  NAND3_X1 U47575 ( .A1(n33356), .A2(n33684), .A3(n32896), .ZN(n32904) );
  NOR2_X1 U47577 ( .A1(n34150), .A2(n61197), .ZN(n33677) );
  NAND3_X1 U47578 ( .A1(n33677), .A2(n33676), .A3(n34146), .ZN(n32902) );
  MUX2_X1 U47579 ( .I0(n32906), .I1(n32905), .S(n24198), .Z(n32913) );
  NAND2_X1 U47580 ( .A1(n62041), .A2(n24198), .ZN(n36928) );
  INV_X1 U47581 ( .I(n36928), .ZN(n32908) );
  NAND3_X1 U47582 ( .A1(n34924), .A2(n35506), .A3(n35949), .ZN(n32911) );
  INV_X1 U47583 ( .I(n38414), .ZN(n33335) );
  NAND2_X1 U47584 ( .A1(n33509), .A2(n34542), .ZN(n32916) );
  OAI21_X1 U47587 ( .A1(n63581), .A2(n34247), .B(n34719), .ZN(n32923) );
  NAND2_X1 U47588 ( .A1(n34352), .A2(n32923), .ZN(n32926) );
  INV_X1 U47590 ( .I(n32934), .ZN(n34252) );
  OAI22_X1 U47591 ( .A1(n32928), .A2(n32927), .B1(n34254), .B2(n34252), .ZN(
        n32929) );
  MUX2_X1 U47595 ( .I0(n32932), .I1(n32931), .S(n32933), .Z(n32938) );
  OAI22_X1 U47596 ( .A1(n32933), .A2(n33747), .B1(n34720), .B2(n64965), .ZN(
        n32936) );
  NAND2_X1 U47599 ( .A1(n34771), .A2(n23567), .ZN(n32942) );
  AOI21_X1 U47600 ( .A1(n34213), .A2(n32942), .B(n21388), .ZN(n32943) );
  NOR2_X1 U47602 ( .A1(n23761), .A2(n560), .ZN(n32953) );
  AOI21_X1 U47603 ( .A1(n32951), .A2(n23761), .B(n32950), .ZN(n32952) );
  NAND2_X1 U47607 ( .A1(n34948), .A2(n58713), .ZN(n32963) );
  OAI21_X1 U47609 ( .A1(n34956), .A2(n33752), .B(n1545), .ZN(n32966) );
  INV_X1 U47610 ( .I(n35533), .ZN(n32977) );
  NOR2_X1 U47611 ( .A1(n34777), .A2(n61028), .ZN(n32974) );
  NAND4_X1 U47614 ( .A1(n32985), .A2(n35529), .A3(n36558), .A4(n35534), .ZN(
        n32986) );
  INV_X1 U47615 ( .I(n32987), .ZN(n39218) );
  XOR2_X1 U47616 ( .A1(n39218), .A2(n32988), .Z(n50608) );
  XOR2_X1 U47617 ( .A1(n53487), .A2(n55349), .Z(n37142) );
  XOR2_X1 U47618 ( .A1(n45878), .A2(n37142), .Z(n52160) );
  XOR2_X1 U47619 ( .A1(n50608), .A2(n52160), .Z(n32989) );
  XOR2_X1 U47620 ( .A1(n37511), .A2(n32989), .Z(n33127) );
  NAND2_X1 U47622 ( .A1(n35629), .A2(n59134), .ZN(n35614) );
  NAND2_X1 U47623 ( .A1(n35624), .A2(n32684), .ZN(n32994) );
  AOI21_X1 U47624 ( .A1(n35207), .A2(n32994), .B(n35612), .ZN(n32995) );
  NOR2_X1 U47625 ( .A1(n33006), .A2(n33611), .ZN(n33007) );
  NOR2_X1 U47626 ( .A1(n1808), .A2(n35688), .ZN(n36541) );
  NOR2_X1 U47627 ( .A1(n33017), .A2(n11061), .ZN(n36542) );
  INV_X1 U47632 ( .I(n33024), .ZN(n33025) );
  XOR2_X1 U47633 ( .A1(n245), .A2(n33025), .Z(n38073) );
  XOR2_X1 U47634 ( .A1(n38073), .A2(n22773), .Z(n44981) );
  XOR2_X1 U47635 ( .A1(n52734), .A2(n58084), .Z(n46501) );
  XOR2_X1 U47636 ( .A1(n52095), .A2(n46501), .Z(n33026) );
  XOR2_X1 U47637 ( .A1(n51234), .A2(n33026), .Z(n33027) );
  XOR2_X1 U47638 ( .A1(n44981), .A2(n33027), .Z(n33028) );
  XOR2_X1 U47639 ( .A1(n33158), .A2(n33028), .Z(n33029) );
  XOR2_X1 U47640 ( .A1(n38885), .A2(n56702), .Z(n46684) );
  XOR2_X1 U47641 ( .A1(n727), .A2(n33034), .Z(n33040) );
  XOR2_X1 U47642 ( .A1(n38650), .A2(n52565), .Z(n38698) );
  XOR2_X1 U47643 ( .A1(n39375), .A2(n54126), .Z(n33036) );
  XOR2_X1 U47644 ( .A1(n38558), .A2(n33036), .Z(n44749) );
  XOR2_X1 U47645 ( .A1(n39478), .A2(n51165), .Z(n45417) );
  XOR2_X1 U47646 ( .A1(n44749), .A2(n45417), .Z(n33037) );
  XOR2_X1 U47647 ( .A1(n38698), .A2(n33037), .Z(n33038) );
  XOR2_X1 U47648 ( .A1(n10553), .A2(n33038), .Z(n33039) );
  XOR2_X1 U47649 ( .A1(n33040), .A2(n33039), .Z(n33041) );
  XOR2_X1 U47650 ( .A1(n33044), .A2(n33043), .Z(n33050) );
  XOR2_X1 U47651 ( .A1(n39631), .A2(n620), .Z(n37809) );
  XNOR2_X1 U47652 ( .A1(n23989), .A2(n54219), .ZN(n33045) );
  XOR2_X1 U47653 ( .A1(n53945), .A2(n53748), .Z(n39556) );
  XOR2_X1 U47654 ( .A1(n33045), .A2(n39556), .Z(n33046) );
  XOR2_X1 U47655 ( .A1(n37809), .A2(n33046), .Z(n45853) );
  XOR2_X1 U47656 ( .A1(n50798), .A2(n55534), .Z(n44599) );
  XOR2_X1 U47657 ( .A1(n45853), .A2(n44599), .Z(n33047) );
  XOR2_X1 U47658 ( .A1(n33049), .A2(n33050), .Z(n33052) );
  XOR2_X1 U47659 ( .A1(n33055), .A2(n56475), .Z(n44148) );
  XOR2_X1 U47660 ( .A1(n44148), .A2(n33056), .Z(n33057) );
  INV_X1 U47661 ( .I(n22252), .ZN(n33061) );
  XOR2_X1 U47662 ( .A1(n33062), .A2(n33061), .Z(n47937) );
  XOR2_X1 U47663 ( .A1(n47937), .A2(n23968), .Z(n45867) );
  XOR2_X1 U47664 ( .A1(n37739), .A2(n56745), .Z(n51310) );
  XOR2_X1 U47665 ( .A1(n51310), .A2(n33063), .Z(n44579) );
  XOR2_X1 U47666 ( .A1(n44579), .A2(n50196), .Z(n33064) );
  XOR2_X1 U47667 ( .A1(n45867), .A2(n33064), .Z(n33065) );
  INV_X1 U47668 ( .I(n23667), .ZN(n33067) );
  XOR2_X1 U47669 ( .A1(n52354), .A2(n37637), .Z(n42021) );
  XOR2_X1 U47670 ( .A1(n42021), .A2(n43864), .Z(n33072) );
  XOR2_X1 U47671 ( .A1(n1881), .A2(n33071), .Z(n49957) );
  XOR2_X1 U47672 ( .A1(n33072), .A2(n49957), .Z(n33073) );
  NAND2_X1 U47674 ( .A1(n33820), .A2(n57986), .ZN(n33081) );
  NOR2_X1 U47676 ( .A1(n35663), .A2(n7321), .ZN(n33130) );
  NOR2_X1 U47678 ( .A1(n35663), .A2(n1341), .ZN(n33084) );
  NOR2_X1 U47693 ( .A1(n19206), .A2(n36385), .ZN(n33121) );
  AOI21_X1 U47695 ( .A1(n33130), .A2(n62322), .B(n35217), .ZN(n33131) );
  XOR2_X1 U47696 ( .A1(n36357), .A2(n55395), .Z(n33133) );
  XOR2_X1 U47697 ( .A1(n33133), .A2(n49273), .Z(n33136) );
  XOR2_X1 U47698 ( .A1(n58928), .A2(n38380), .Z(n33135) );
  XOR2_X1 U47699 ( .A1(n33136), .A2(n33135), .Z(n45370) );
  XOR2_X1 U47700 ( .A1(n21531), .A2(n45370), .Z(n33137) );
  XOR2_X1 U47701 ( .A1(n33148), .A2(n33147), .Z(n38107) );
  XOR2_X1 U47702 ( .A1(n50955), .A2(n54386), .Z(n37764) );
  XOR2_X1 U47703 ( .A1(n38107), .A2(n37764), .Z(n43758) );
  XOR2_X1 U47704 ( .A1(n51021), .A2(n44014), .Z(n33149) );
  XOR2_X1 U47705 ( .A1(n43758), .A2(n33149), .Z(n33151) );
  XOR2_X1 U47706 ( .A1(n33150), .A2(n33151), .Z(n33152) );
  XOR2_X1 U47707 ( .A1(n52614), .A2(n22961), .Z(n50912) );
  XOR2_X1 U47708 ( .A1(n24046), .A2(n56784), .Z(n52018) );
  XOR2_X1 U47709 ( .A1(n52018), .A2(n56322), .Z(n33156) );
  XOR2_X1 U47710 ( .A1(n50912), .A2(n33156), .Z(n33157) );
  XOR2_X1 U47711 ( .A1(n33165), .A2(n37303), .Z(n37950) );
  XOR2_X1 U47712 ( .A1(n39705), .A2(n37950), .Z(n44830) );
  XOR2_X1 U47713 ( .A1(n33166), .A2(n39375), .Z(n37073) );
  XOR2_X1 U47714 ( .A1(n37073), .A2(n33167), .Z(n46302) );
  XOR2_X1 U47715 ( .A1(n44830), .A2(n46302), .Z(n33168) );
  XOR2_X1 U47716 ( .A1(n16884), .A2(n33169), .Z(n33170) );
  XOR2_X1 U47718 ( .A1(n33174), .A2(n17616), .Z(n33175) );
  XOR2_X1 U47719 ( .A1(n33176), .A2(n33177), .Z(n33286) );
  XOR2_X1 U47720 ( .A1(n33286), .A2(n23465), .Z(n33189) );
  XOR2_X1 U47721 ( .A1(n33179), .A2(n37983), .Z(n44331) );
  XOR2_X1 U47722 ( .A1(n54888), .A2(n60556), .Z(n38460) );
  XOR2_X1 U47723 ( .A1(n33180), .A2(n38460), .Z(n33181) );
  XOR2_X1 U47724 ( .A1(n53748), .A2(n54219), .Z(n37847) );
  XOR2_X1 U47725 ( .A1(n33181), .A2(n37847), .Z(n45396) );
  XOR2_X1 U47726 ( .A1(n620), .A2(n56309), .Z(n33182) );
  XOR2_X1 U47727 ( .A1(n45396), .A2(n33182), .Z(n33183) );
  XOR2_X1 U47728 ( .A1(n44331), .A2(n33183), .Z(n33184) );
  XOR2_X1 U47729 ( .A1(n23683), .A2(n33184), .Z(n33187) );
  XOR2_X1 U47730 ( .A1(n33187), .A2(n33186), .Z(n33188) );
  XOR2_X1 U47731 ( .A1(n33194), .A2(n33193), .Z(n33200) );
  XOR2_X1 U47732 ( .A1(n38904), .A2(n37497), .Z(n51280) );
  XOR2_X1 U47733 ( .A1(n51275), .A2(n54185), .Z(n51218) );
  XOR2_X1 U47734 ( .A1(n51218), .A2(n33195), .Z(n33196) );
  XOR2_X1 U47735 ( .A1(n51280), .A2(n33196), .Z(n33197) );
  XOR2_X1 U47736 ( .A1(n20838), .A2(n33197), .Z(n33198) );
  XOR2_X1 U47737 ( .A1(n33200), .A2(n33199), .Z(n33201) );
  XOR2_X1 U47738 ( .A1(n33202), .A2(n33201), .Z(n33209) );
  XOR2_X1 U47739 ( .A1(n33205), .A2(n33204), .Z(n33206) );
  XOR2_X1 U47740 ( .A1(n33207), .A2(n33206), .Z(n33208) );
  XOR2_X1 U47741 ( .A1(n33209), .A2(n33208), .Z(n35710) );
  NOR2_X1 U47744 ( .A1(n59824), .A2(n33212), .ZN(n33213) );
  INV_X1 U47745 ( .I(n33219), .ZN(n33541) );
  OAI21_X1 U47746 ( .A1(n33224), .A2(n33375), .B(n33627), .ZN(n33222) );
  INV_X1 U47747 ( .I(n33220), .ZN(n33221) );
  NAND3_X1 U47748 ( .A1(n60434), .A2(n33537), .A3(n14329), .ZN(n33223) );
  XOR2_X1 U47751 ( .A1(n38628), .A2(n33226), .Z(n46500) );
  XOR2_X1 U47752 ( .A1(n45404), .A2(n52734), .Z(n39613) );
  XOR2_X1 U47753 ( .A1(n39613), .A2(n56784), .Z(n33227) );
  XOR2_X1 U47754 ( .A1(n51596), .A2(n33227), .Z(n33228) );
  XOR2_X1 U47755 ( .A1(n38555), .A2(n33234), .Z(n52566) );
  XOR2_X1 U47756 ( .A1(n52566), .A2(n38558), .Z(n46191) );
  XOR2_X1 U47757 ( .A1(n52900), .A2(n55840), .Z(n33235) );
  XOR2_X1 U47758 ( .A1(n38826), .A2(n33235), .Z(n33236) );
  XOR2_X1 U47759 ( .A1(n45470), .A2(n33236), .Z(n42950) );
  XOR2_X1 U47760 ( .A1(n46191), .A2(n42950), .Z(n33237) );
  XOR2_X1 U47762 ( .A1(n33857), .A2(n20673), .Z(n33240) );
  XOR2_X1 U47763 ( .A1(n33242), .A2(n33243), .Z(n33244) );
  XOR2_X1 U47764 ( .A1(n33898), .A2(n33244), .Z(n33251) );
  XOR2_X1 U47765 ( .A1(n38301), .A2(n54407), .Z(n46203) );
  XOR2_X1 U47766 ( .A1(n46203), .A2(n51218), .Z(n33245) );
  XOR2_X1 U47767 ( .A1(n33245), .A2(n42730), .Z(n33246) );
  XOR2_X1 U47768 ( .A1(n61034), .A2(n23929), .Z(n39753) );
  XOR2_X1 U47769 ( .A1(n39753), .A2(n49955), .Z(n42710) );
  XOR2_X1 U47770 ( .A1(n33246), .A2(n42710), .Z(n33247) );
  XOR2_X1 U47771 ( .A1(n33247), .A2(n20838), .Z(n33249) );
  XOR2_X1 U47772 ( .A1(n33248), .A2(n33249), .Z(n33250) );
  XOR2_X1 U47773 ( .A1(n33251), .A2(n33250), .Z(n33252) );
  NAND2_X1 U47775 ( .A1(n34448), .A2(n35247), .ZN(n33275) );
  XOR2_X1 U47776 ( .A1(n30908), .A2(n54716), .Z(n33257) );
  XOR2_X1 U47777 ( .A1(n37764), .A2(n33257), .Z(n43728) );
  XOR2_X1 U47778 ( .A1(n602), .A2(n43728), .Z(n33260) );
  XOR2_X1 U47779 ( .A1(n39295), .A2(n37767), .Z(n33259) );
  XOR2_X1 U47780 ( .A1(n33259), .A2(n50873), .Z(n51801) );
  XOR2_X1 U47781 ( .A1(n51801), .A2(n54896), .Z(n37999) );
  XOR2_X1 U47782 ( .A1(n37999), .A2(n29969), .Z(n44358) );
  XOR2_X1 U47783 ( .A1(n33260), .A2(n44358), .Z(n33262) );
  XOR2_X1 U47784 ( .A1(n23667), .A2(n22363), .Z(n33265) );
  XOR2_X1 U47785 ( .A1(n38007), .A2(n23020), .Z(n39684) );
  XOR2_X1 U47786 ( .A1(n38862), .A2(n45371), .Z(n51992) );
  XOR2_X1 U47787 ( .A1(n39684), .A2(n51992), .Z(n44536) );
  XOR2_X1 U47788 ( .A1(n44533), .A2(n50486), .Z(n33267) );
  XOR2_X1 U47789 ( .A1(n44536), .A2(n33267), .Z(n33268) );
  XOR2_X1 U47790 ( .A1(n33269), .A2(n33268), .Z(n33270) );
  XOR2_X1 U47791 ( .A1(n33271), .A2(n33270), .Z(n33273) );
  NAND2_X1 U47792 ( .A1(n35655), .A2(n35247), .ZN(n33274) );
  NAND2_X1 U47793 ( .A1(n35659), .A2(n35241), .ZN(n33278) );
  XOR2_X1 U47794 ( .A1(n33279), .A2(n42391), .Z(n36930) );
  XOR2_X1 U47795 ( .A1(n36930), .A2(n33280), .Z(n39332) );
  XOR2_X1 U47796 ( .A1(n53787), .A2(n23989), .Z(n44424) );
  XOR2_X1 U47797 ( .A1(n39332), .A2(n44424), .Z(n45321) );
  INV_X1 U47798 ( .I(n33281), .ZN(n37852) );
  XOR2_X1 U47799 ( .A1(n50798), .A2(n56309), .Z(n33282) );
  XOR2_X1 U47800 ( .A1(n37852), .A2(n33282), .Z(n44543) );
  XOR2_X1 U47801 ( .A1(n45321), .A2(n44543), .Z(n33284) );
  XOR2_X1 U47802 ( .A1(n33284), .A2(n33283), .Z(n33285) );
  INV_X1 U47803 ( .I(n33286), .ZN(n33287) );
  NAND2_X1 U47805 ( .A1(n35645), .A2(n35656), .ZN(n33295) );
  NAND3_X1 U47806 ( .A1(n34374), .A2(n4969), .A3(n37376), .ZN(n33326) );
  NOR2_X1 U47807 ( .A1(n22723), .A2(n10682), .ZN(n33301) );
  OAI21_X1 U47808 ( .A1(n33306), .A2(n33305), .B(n33304), .ZN(n33309) );
  NAND3_X1 U47809 ( .A1(n61699), .A2(n32684), .A3(n33542), .ZN(n33314) );
  OAI21_X1 U47810 ( .A1(n33315), .A2(n35611), .B(n33314), .ZN(n33317) );
  INV_X1 U47811 ( .I(n35199), .ZN(n33320) );
  OAI22_X1 U47812 ( .A1(n6527), .A2(n35614), .B1(n33320), .B2(n33319), .ZN(
        n33322) );
  NAND2_X1 U47814 ( .A1(n36520), .A2(n37369), .ZN(n33327) );
  NAND3_X1 U47816 ( .A1(n36589), .A2(n37376), .A3(n2594), .ZN(n33328) );
  INV_X1 U47817 ( .I(n36511), .ZN(n33330) );
  NAND3_X1 U47819 ( .A1(n60456), .A2(n33601), .A3(n35687), .ZN(n33339) );
  OAI21_X1 U47823 ( .A1(n33359), .A2(n33358), .B(n33357), .ZN(n33360) );
  NAND2_X1 U47827 ( .A1(n33374), .A2(n33540), .ZN(n33377) );
  NAND2_X1 U47828 ( .A1(n33375), .A2(n33537), .ZN(n33376) );
  NAND3_X1 U47829 ( .A1(n63866), .A2(n33627), .A3(n5250), .ZN(n33378) );
  NOR2_X1 U47830 ( .A1(n34132), .A2(n34137), .ZN(n33384) );
  NAND3_X1 U47831 ( .A1(n34134), .A2(n34142), .A3(n33654), .ZN(n33386) );
  NOR2_X1 U47833 ( .A1(n22598), .A2(n34128), .ZN(n33393) );
  NOR2_X1 U47835 ( .A1(n22598), .A2(n157), .ZN(n33395) );
  AOI21_X1 U47836 ( .A1(n19663), .A2(n157), .B(n34137), .ZN(n33400) );
  NAND3_X1 U47837 ( .A1(n33616), .A2(n33614), .A3(n63085), .ZN(n33403) );
  NAND2_X1 U47838 ( .A1(n33405), .A2(n1796), .ZN(n33407) );
  INV_X1 U47839 ( .I(n36259), .ZN(n33411) );
  INV_X1 U47840 ( .I(n36257), .ZN(n33409) );
  INV_X1 U47843 ( .I(n33422), .ZN(n33423) );
  INV_X1 U47845 ( .I(n34020), .ZN(n33428) );
  NAND2_X1 U47846 ( .A1(n35026), .A2(n64708), .ZN(n33426) );
  OAI22_X1 U47847 ( .A1(n33428), .A2(n33427), .B1(n35020), .B2(n33426), .ZN(
        n33429) );
  INV_X1 U47848 ( .I(n34908), .ZN(n34482) );
  INV_X1 U47849 ( .I(n34621), .ZN(n33438) );
  INV_X1 U47851 ( .I(n34641), .ZN(n33446) );
  NOR2_X1 U47856 ( .A1(n36944), .A2(n22993), .ZN(n35428) );
  OAI21_X1 U47857 ( .A1(n1789), .A2(n64101), .B(n35428), .ZN(n33457) );
  AOI21_X1 U47858 ( .A1(n36892), .A2(n35433), .B(n1789), .ZN(n33459) );
  NOR2_X1 U47862 ( .A1(n560), .A2(n9766), .ZN(n33466) );
  MUX2_X1 U47863 ( .I0(n33466), .I1(n34787), .S(n64158), .Z(n33475) );
  NAND2_X1 U47864 ( .A1(n34797), .A2(n33467), .ZN(n33471) );
  NAND2_X1 U47865 ( .A1(n12405), .A2(n60926), .ZN(n33476) );
  NAND2_X1 U47866 ( .A1(n20660), .A2(n58713), .ZN(n33478) );
  INV_X1 U47868 ( .I(n34570), .ZN(n33482) );
  NOR2_X1 U47870 ( .A1(n57710), .A2(n61256), .ZN(n33488) );
  NOR4_X1 U47871 ( .A1(n34784), .A2(n57710), .A3(n61108), .A4(n1430), .ZN(
        n33487) );
  AOI21_X1 U47872 ( .A1(n33489), .A2(n33488), .B(n33487), .ZN(n33492) );
  OAI21_X1 U47873 ( .A1(n33777), .A2(n33776), .B(n34786), .ZN(n33490) );
  AOI22_X1 U47875 ( .A1(n10175), .A2(n3325), .B1(n33770), .B2(n63319), .ZN(
        n33495) );
  NOR2_X1 U47876 ( .A1(n34534), .A2(n33729), .ZN(n33728) );
  NOR2_X1 U47877 ( .A1(n34972), .A2(n34529), .ZN(n33723) );
  NOR2_X1 U47878 ( .A1(n33723), .A2(n33496), .ZN(n33498) );
  NOR2_X1 U47880 ( .A1(n34969), .A2(n34538), .ZN(n33497) );
  INV_X1 U47881 ( .I(n33725), .ZN(n33505) );
  INV_X1 U47882 ( .I(n33500), .ZN(n33501) );
  NOR2_X1 U47884 ( .A1(n25404), .A2(n34970), .ZN(n33502) );
  AOI22_X1 U47885 ( .A1(n33505), .A2(n33504), .B1(n33503), .B2(n33502), .ZN(
        n33508) );
  INV_X1 U47887 ( .I(n34544), .ZN(n34968) );
  NAND2_X1 U47888 ( .A1(n57423), .A2(n22419), .ZN(n33510) );
  NAND2_X1 U47889 ( .A1(n34968), .A2(n33510), .ZN(n33514) );
  NAND2_X1 U47891 ( .A1(n33511), .A2(n25404), .ZN(n33512) );
  NAND2_X1 U47892 ( .A1(n24077), .A2(n34025), .ZN(n34021) );
  NAND2_X1 U47893 ( .A1(n34021), .A2(n2207), .ZN(n33517) );
  NOR2_X1 U47894 ( .A1(n10340), .A2(n2207), .ZN(n33521) );
  NAND2_X1 U47897 ( .A1(n36150), .A2(n33523), .ZN(n33524) );
  AOI21_X1 U47898 ( .A1(n798), .A2(n64087), .B(n33526), .ZN(n33525) );
  NOR2_X1 U47899 ( .A1(n36584), .A2(n33525), .ZN(n33528) );
  NAND2_X1 U47900 ( .A1(n36154), .A2(n11272), .ZN(n33527) );
  INV_X1 U47901 ( .I(n45101), .ZN(n50606) );
  INV_X1 U47902 ( .I(n37820), .ZN(n33529) );
  NOR2_X1 U47903 ( .A1(n33539), .A2(n61350), .ZN(n33530) );
  NAND2_X1 U47904 ( .A1(n33547), .A2(n35618), .ZN(n33545) );
  NAND3_X1 U47905 ( .A1(n33543), .A2(n33550), .A3(n35206), .ZN(n33544) );
  MUX2_X1 U47906 ( .I0(n33545), .I1(n33544), .S(n35612), .Z(n33558) );
  NAND2_X1 U47908 ( .A1(n35198), .A2(n33550), .ZN(n33552) );
  INV_X1 U47909 ( .I(n35622), .ZN(n33553) );
  OAI21_X1 U47910 ( .A1(n33554), .A2(n35206), .B(n33553), .ZN(n33555) );
  OAI21_X1 U47911 ( .A1(n33575), .A2(n33574), .B(n57200), .ZN(n33582) );
  NAND2_X1 U47912 ( .A1(n24286), .A2(n23179), .ZN(n33576) );
  NAND2_X1 U47915 ( .A1(n35650), .A2(n35247), .ZN(n33585) );
  NAND4_X1 U47916 ( .A1(n33585), .A2(n35249), .A3(n22909), .A4(n33801), .ZN(
        n33593) );
  NOR2_X1 U47917 ( .A1(n35651), .A2(n35241), .ZN(n35660) );
  AOI21_X1 U47919 ( .A1(n35654), .A2(n35647), .B(n33587), .ZN(n33588) );
  NAND4_X1 U47920 ( .A1(n35642), .A2(n35656), .A3(n33589), .A4(n35643), .ZN(
        n33590) );
  OAI21_X1 U47921 ( .A1(n11061), .A2(n24688), .B(n35688), .ZN(n33594) );
  OAI21_X1 U47922 ( .A1(n33595), .A2(n33594), .B(n9679), .ZN(n33603) );
  NAND3_X1 U47924 ( .A1(n33601), .A2(n33600), .A3(n63273), .ZN(n33602) );
  NOR2_X1 U47929 ( .A1(n23127), .A2(n1542), .ZN(n33620) );
  INV_X1 U47930 ( .I(n33639), .ZN(n33626) );
  NOR2_X1 U47931 ( .A1(n24093), .A2(n33627), .ZN(n33631) );
  INV_X1 U47933 ( .I(n33634), .ZN(n33641) );
  NAND2_X1 U47934 ( .A1(n63103), .A2(n33635), .ZN(n33640) );
  AOI22_X1 U47936 ( .A1(n33641), .A2(n33640), .B1(n33639), .B2(n33638), .ZN(
        n33647) );
  NAND2_X1 U47937 ( .A1(n33663), .A2(n33654), .ZN(n33651) );
  NOR2_X1 U47939 ( .A1(n34132), .A2(n33654), .ZN(n33656) );
  OAI21_X1 U47940 ( .A1(n33657), .A2(n33656), .B(n33655), .ZN(n33658) );
  NAND2_X1 U47944 ( .A1(n33677), .A2(n33676), .ZN(n33678) );
  AOI22_X1 U47945 ( .A1(n33682), .A2(n33681), .B1(n34152), .B2(n33680), .ZN(
        n33687) );
  NOR2_X1 U47947 ( .A1(n33689), .A2(n33702), .ZN(n33692) );
  OAI22_X1 U47949 ( .A1(n33695), .A2(n33694), .B1(n33701), .B2(n33693), .ZN(
        n33696) );
  AOI21_X1 U47950 ( .A1(n33698), .A2(n7273), .B(n33696), .ZN(n33707) );
  INV_X1 U47951 ( .I(n33699), .ZN(n33700) );
  NAND2_X1 U47952 ( .A1(n33704), .A2(n33703), .ZN(n33705) );
  NAND2_X1 U47953 ( .A1(n34194), .A2(n60684), .ZN(n33713) );
  NOR2_X1 U47955 ( .A1(n35964), .A2(n35962), .ZN(n35148) );
  NAND3_X1 U47956 ( .A1(n34544), .A2(n34546), .A3(n33722), .ZN(n33736) );
  NAND2_X1 U47958 ( .A1(n7883), .A2(n60579), .ZN(n33724) );
  NOR2_X1 U47960 ( .A1(n33729), .A2(n34970), .ZN(n33731) );
  OAI21_X1 U47961 ( .A1(n33731), .A2(n34971), .B(n33730), .ZN(n33733) );
  NAND2_X1 U47962 ( .A1(n34546), .A2(n22419), .ZN(n33732) );
  NAND3_X1 U47963 ( .A1(n33733), .A2(n57423), .A3(n33732), .ZN(n33734) );
  NAND3_X1 U47965 ( .A1(n34727), .A2(n4591), .A3(n34355), .ZN(n33739) );
  AOI21_X1 U47966 ( .A1(n34725), .A2(n33739), .B(n33747), .ZN(n33740) );
  NAND2_X1 U47968 ( .A1(n34719), .A2(n34247), .ZN(n33742) );
  AOI21_X1 U47969 ( .A1(n34720), .A2(n64965), .B(n33742), .ZN(n33745) );
  NOR2_X1 U47970 ( .A1(n34358), .A2(n33743), .ZN(n33744) );
  AOI21_X1 U47971 ( .A1(n15184), .A2(n4591), .B(n1536), .ZN(n33746) );
  NAND2_X1 U47972 ( .A1(n23761), .A2(n33762), .ZN(n33764) );
  NAND3_X1 U47973 ( .A1(n33767), .A2(n61028), .A3(n34273), .ZN(n33773) );
  OAI21_X1 U47977 ( .A1(n33777), .A2(n61108), .B(n33776), .ZN(n33778) );
  NAND2_X1 U47978 ( .A1(n65160), .A2(n1227), .ZN(n36418) );
  AOI21_X1 U47979 ( .A1(n35130), .A2(n59468), .B(n36418), .ZN(n33781) );
  NAND2_X1 U47980 ( .A1(n36427), .A2(n3458), .ZN(n33783) );
  NOR2_X1 U47981 ( .A1(n35130), .A2(n59468), .ZN(n33787) );
  INV_X1 U47982 ( .I(n36179), .ZN(n33789) );
  NOR2_X1 U47983 ( .A1(n36432), .A2(n36121), .ZN(n33790) );
  NOR2_X1 U47985 ( .A1(n35656), .A2(n35247), .ZN(n33791) );
  NOR2_X1 U47987 ( .A1(n35656), .A2(n58598), .ZN(n33795) );
  NOR2_X1 U47989 ( .A1(n33798), .A2(n9030), .ZN(n33799) );
  NOR2_X1 U47991 ( .A1(n35651), .A2(n35247), .ZN(n34444) );
  NAND3_X1 U47992 ( .A1(n34444), .A2(n33802), .A3(n33801), .ZN(n33803) );
  NAND2_X1 U47993 ( .A1(n34392), .A2(n15018), .ZN(n35717) );
  NOR2_X1 U47996 ( .A1(n33811), .A2(n35759), .ZN(n33812) );
  NOR3_X1 U47997 ( .A1(n63220), .A2(n35322), .A3(n34438), .ZN(n33817) );
  NAND2_X1 U47998 ( .A1(n21096), .A2(n35318), .ZN(n33815) );
  NAND2_X1 U47999 ( .A1(n37090), .A2(n37319), .ZN(n37316) );
  NAND2_X1 U48000 ( .A1(n59825), .A2(n37316), .ZN(n33917) );
  INV_X1 U48002 ( .I(n33820), .ZN(n35668) );
  OAI21_X1 U48003 ( .A1(n35668), .A2(n35662), .B(n57200), .ZN(n33821) );
  NOR2_X1 U48004 ( .A1(n6979), .A2(n57986), .ZN(n33826) );
  XOR2_X1 U48007 ( .A1(n39611), .A2(n56180), .Z(n39362) );
  XOR2_X1 U48008 ( .A1(n39362), .A2(n55139), .Z(n33830) );
  XOR2_X1 U48009 ( .A1(n37481), .A2(n50245), .Z(n52020) );
  XOR2_X1 U48010 ( .A1(n33830), .A2(n52020), .Z(n45036) );
  XOR2_X1 U48011 ( .A1(n45036), .A2(n33831), .Z(n33832) );
  XOR2_X1 U48013 ( .A1(n33835), .A2(n33834), .Z(n33836) );
  INV_X1 U48014 ( .I(n33837), .ZN(n33844) );
  XOR2_X1 U48015 ( .A1(n33838), .A2(n33839), .Z(n33842) );
  XOR2_X1 U48016 ( .A1(n9609), .A2(n33840), .Z(n33841) );
  XOR2_X1 U48017 ( .A1(n33842), .A2(n33841), .Z(n33843) );
  XOR2_X1 U48018 ( .A1(n33844), .A2(n33843), .Z(n33845) );
  XOR2_X1 U48019 ( .A1(n33846), .A2(n33845), .Z(n33847) );
  XOR2_X1 U48020 ( .A1(n1550), .A2(n64968), .Z(n33850) );
  XOR2_X1 U48021 ( .A1(n33849), .A2(n33850), .Z(n33861) );
  XOR2_X1 U48022 ( .A1(n38280), .A2(n39196), .Z(n46616) );
  INV_X1 U48023 ( .I(n33851), .ZN(n33852) );
  XOR2_X1 U48024 ( .A1(n46616), .A2(n33852), .Z(n49967) );
  XOR2_X1 U48025 ( .A1(n56905), .A2(n53772), .Z(n44052) );
  XOR2_X1 U48026 ( .A1(n44052), .A2(n51493), .Z(n33853) );
  XOR2_X1 U48027 ( .A1(n44996), .A2(n33853), .Z(n33854) );
  XOR2_X1 U48028 ( .A1(n49967), .A2(n33854), .Z(n33855) );
  XOR2_X1 U48029 ( .A1(n23869), .A2(n33855), .Z(n33859) );
  XOR2_X1 U48030 ( .A1(n33858), .A2(n33859), .Z(n33860) );
  XOR2_X1 U48031 ( .A1(n23719), .A2(n23690), .Z(n33864) );
  XOR2_X1 U48032 ( .A1(n10363), .A2(n33864), .Z(n33865) );
  XOR2_X1 U48033 ( .A1(n33867), .A2(n54708), .Z(n44164) );
  XOR2_X1 U48034 ( .A1(n33871), .A2(n39445), .Z(n39633) );
  XOR2_X1 U48035 ( .A1(n39633), .A2(n37809), .Z(n45295) );
  INV_X1 U48036 ( .I(n8329), .ZN(n33873) );
  XOR2_X1 U48038 ( .A1(n33878), .A2(n54536), .Z(n39770) );
  XOR2_X1 U48039 ( .A1(n39770), .A2(n51512), .Z(n44263) );
  XOR2_X1 U48041 ( .A1(n37764), .A2(n54153), .Z(n37890) );
  XOR2_X1 U48042 ( .A1(n56040), .A2(n53138), .Z(n39294) );
  XOR2_X1 U48043 ( .A1(n37890), .A2(n39294), .Z(n43902) );
  XOR2_X1 U48044 ( .A1(n33886), .A2(n55242), .Z(n33887) );
  XOR2_X1 U48045 ( .A1(n33887), .A2(n38165), .Z(n44139) );
  XOR2_X1 U48046 ( .A1(n38981), .A2(n61550), .Z(n38235) );
  XOR2_X1 U48047 ( .A1(n44139), .A2(n38235), .Z(n33888) );
  XOR2_X1 U48048 ( .A1(n39738), .A2(n37713), .Z(n45251) );
  XOR2_X1 U48049 ( .A1(n33888), .A2(n45251), .Z(n33890) );
  XOR2_X1 U48050 ( .A1(n33891), .A2(n19069), .Z(n33892) );
  INV_X1 U48051 ( .I(n35286), .ZN(n33894) );
  XOR2_X1 U48052 ( .A1(n51656), .A2(n38177), .Z(n50772) );
  XOR2_X1 U48053 ( .A1(n33901), .A2(n33900), .Z(n33902) );
  XOR2_X1 U48054 ( .A1(n51218), .A2(n33902), .Z(n46141) );
  XOR2_X1 U48055 ( .A1(n50772), .A2(n46141), .Z(n33903) );
  XOR2_X1 U48056 ( .A1(n33903), .A2(n20838), .Z(n33908) );
  XOR2_X1 U48057 ( .A1(n22583), .A2(n18314), .Z(n33907) );
  AOI21_X1 U48061 ( .A1(n33917), .A2(n19252), .B(n65236), .ZN(n33943) );
  OAI21_X1 U48062 ( .A1(n33920), .A2(n33925), .B(n33919), .ZN(n33923) );
  NAND2_X1 U48063 ( .A1(n34427), .A2(n34421), .ZN(n35773) );
  NAND3_X1 U48064 ( .A1(n33925), .A2(n34423), .A3(n35770), .ZN(n33922) );
  AOI21_X1 U48065 ( .A1(n35782), .A2(n33926), .B(n35783), .ZN(n33928) );
  INV_X1 U48068 ( .I(n35081), .ZN(n37023) );
  NOR2_X1 U48069 ( .A1(n22223), .A2(n37096), .ZN(n33935) );
  NOR3_X1 U48071 ( .A1(n37085), .A2(n37319), .A3(n37096), .ZN(n33937) );
  NOR2_X1 U48072 ( .A1(n37945), .A2(n22223), .ZN(n33936) );
  AOI22_X1 U48073 ( .A1(n37023), .A2(n33937), .B1(n33936), .B2(n4745), .ZN(
        n33939) );
  NAND2_X1 U48074 ( .A1(n33953), .A2(n60808), .ZN(n33946) );
  AOI22_X1 U48075 ( .A1(n33950), .A2(n33949), .B1(n34118), .B2(n60892), .ZN(
        n33951) );
  NOR2_X1 U48077 ( .A1(n15819), .A2(n33963), .ZN(n33964) );
  NAND2_X1 U48078 ( .A1(n1312), .A2(n20835), .ZN(n33967) );
  NOR2_X1 U48079 ( .A1(n20607), .A2(n7453), .ZN(n33970) );
  NAND3_X1 U48080 ( .A1(n34042), .A2(n19610), .A3(n23746), .ZN(n33974) );
  NAND3_X1 U48081 ( .A1(n34610), .A2(n34603), .A3(n33974), .ZN(n33976) );
  INV_X1 U48082 ( .I(n34610), .ZN(n33985) );
  NOR2_X1 U48083 ( .A1(n19823), .A2(n10401), .ZN(n33988) );
  NAND2_X1 U48084 ( .A1(n58447), .A2(n34201), .ZN(n33991) );
  INV_X1 U48086 ( .I(n33998), .ZN(n33999) );
  NAND2_X1 U48088 ( .A1(n17096), .A2(n20060), .ZN(n34004) );
  NAND2_X1 U48089 ( .A1(n34008), .A2(n36777), .ZN(n34011) );
  NOR2_X1 U48092 ( .A1(n25657), .A2(n34640), .ZN(n34015) );
  OAI21_X1 U48093 ( .A1(n60984), .A2(n34015), .B(n35039), .ZN(n34016) );
  NAND2_X1 U48094 ( .A1(n34023), .A2(n34022), .ZN(n34024) );
  NAND2_X1 U48095 ( .A1(n64954), .A2(n10340), .ZN(n34027) );
  NAND2_X1 U48096 ( .A1(n34042), .A2(n20507), .ZN(n34036) );
  NAND2_X1 U48098 ( .A1(n34614), .A2(n23746), .ZN(n34043) );
  NAND3_X1 U48099 ( .A1(n34044), .A2(n34602), .A3(n34043), .ZN(n34048) );
  NAND2_X1 U48100 ( .A1(n34046), .A2(n34045), .ZN(n34047) );
  NAND3_X1 U48101 ( .A1(n34680), .A2(n34670), .A3(n34679), .ZN(n34059) );
  INV_X1 U48103 ( .I(n34069), .ZN(n34068) );
  NAND4_X1 U48104 ( .A1(n34071), .A2(n34070), .A3(n63444), .A4(n34069), .ZN(
        n34075) );
  NAND3_X1 U48105 ( .A1(n34073), .A2(n34982), .A3(n34072), .ZN(n34074) );
  NAND3_X1 U48106 ( .A1(n17595), .A2(n36742), .A3(n34077), .ZN(n34094) );
  NOR2_X1 U48107 ( .A1(n34083), .A2(n12039), .ZN(n34085) );
  NAND2_X1 U48108 ( .A1(n23119), .A2(n58421), .ZN(n34089) );
  INV_X1 U48109 ( .I(n36343), .ZN(n34093) );
  NOR2_X1 U48110 ( .A1(n36748), .A2(n1417), .ZN(n35065) );
  NAND2_X1 U48111 ( .A1(n11272), .A2(n60462), .ZN(n34097) );
  NAND2_X1 U48112 ( .A1(n25842), .A2(n60462), .ZN(n34099) );
  MUX2_X1 U48113 ( .I0(n36583), .I1(n34099), .S(n36472), .Z(n34104) );
  NOR2_X1 U48114 ( .A1(n34101), .A2(n34100), .ZN(n34102) );
  OAI21_X1 U48115 ( .A1(n34102), .A2(n10498), .B(n36584), .ZN(n34103) );
  NAND3_X1 U48116 ( .A1(n36262), .A2(n19231), .A3(n3856), .ZN(n34106) );
  NAND2_X1 U48118 ( .A1(n34120), .A2(n62931), .ZN(n34121) );
  NOR2_X1 U48119 ( .A1(n34137), .A2(n34136), .ZN(n34139) );
  NAND2_X1 U48120 ( .A1(n34146), .A2(n23351), .ZN(n34147) );
  NAND2_X1 U48121 ( .A1(n34156), .A2(n34155), .ZN(n34158) );
  NOR2_X1 U48122 ( .A1(n34168), .A2(n34658), .ZN(n34169) );
  NOR2_X1 U48123 ( .A1(n5411), .A2(n60628), .ZN(n34171) );
  NOR2_X1 U48124 ( .A1(n34185), .A2(n118), .ZN(n34192) );
  NAND2_X1 U48126 ( .A1(n15720), .A2(n20147), .ZN(n36700) );
  INV_X1 U48127 ( .I(n36700), .ZN(n34204) );
  INV_X1 U48128 ( .I(n35463), .ZN(n34205) );
  INV_X1 U48129 ( .I(n34208), .ZN(n34211) );
  OAI21_X1 U48130 ( .A1(n34771), .A2(n21388), .B(n65194), .ZN(n34210) );
  AOI21_X1 U48131 ( .A1(n60738), .A2(n34211), .B(n34210), .ZN(n34216) );
  NOR3_X1 U48132 ( .A1(n34760), .A2(n23366), .A3(n60738), .ZN(n34215) );
  NOR3_X1 U48134 ( .A1(n35806), .A2(n35805), .A3(n34385), .ZN(n34228) );
  OAI21_X1 U48138 ( .A1(n34237), .A2(n35827), .B(n34714), .ZN(n34244) );
  NAND4_X1 U48140 ( .A1(n34241), .A2(n34240), .A3(n22633), .A4(n34239), .ZN(
        n34242) );
  NAND2_X1 U48141 ( .A1(n34250), .A2(n4591), .ZN(n34258) );
  NAND2_X1 U48142 ( .A1(n34360), .A2(n23281), .ZN(n34257) );
  NOR2_X1 U48146 ( .A1(n17958), .A2(n35301), .ZN(n34263) );
  NOR2_X1 U48147 ( .A1(n34269), .A2(n20989), .ZN(n34271) );
  NAND2_X1 U48148 ( .A1(n34278), .A2(n19457), .ZN(n34282) );
  NOR2_X1 U48149 ( .A1(n61028), .A2(n57710), .ZN(n34281) );
  NAND2_X1 U48150 ( .A1(n34779), .A2(n1815), .ZN(n34280) );
  NOR2_X1 U48151 ( .A1(n36914), .A2(n36904), .ZN(n34286) );
  NOR2_X1 U48152 ( .A1(n64967), .A2(n37426), .ZN(n34290) );
  AOI21_X1 U48153 ( .A1(n34290), .A2(n36916), .B(n37437), .ZN(n34292) );
  NAND2_X1 U48154 ( .A1(n35941), .A2(n37422), .ZN(n34291) );
  NAND2_X1 U48155 ( .A1(n36916), .A2(n37436), .ZN(n37432) );
  NOR2_X1 U48160 ( .A1(n21388), .A2(n23567), .ZN(n34310) );
  NOR2_X1 U48161 ( .A1(n34311), .A2(n34310), .ZN(n34313) );
  NAND2_X1 U48164 ( .A1(n35822), .A2(n34321), .ZN(n34320) );
  NAND2_X1 U48165 ( .A1(n732), .A2(n34714), .ZN(n34323) );
  NOR2_X1 U48166 ( .A1(n34321), .A2(n34714), .ZN(n34322) );
  AOI21_X1 U48167 ( .A1(n26242), .A2(n23556), .B(n22797), .ZN(n34326) );
  NOR3_X1 U48168 ( .A1(n35820), .A2(n35817), .A3(n34324), .ZN(n34325) );
  NAND4_X1 U48170 ( .A1(n35769), .A2(n58231), .A3(n35775), .A4(n10769), .ZN(
        n34332) );
  INV_X1 U48171 ( .I(n34340), .ZN(n34345) );
  OAI22_X1 U48172 ( .A1(n34345), .A2(n23354), .B1(n34344), .B2(n34343), .ZN(
        n34348) );
  OAI21_X1 U48173 ( .A1(n34356), .A2(n34355), .B(n63581), .ZN(n34357) );
  INV_X1 U48174 ( .I(n37131), .ZN(n34361) );
  INV_X1 U48175 ( .I(n34853), .ZN(n34364) );
  AOI21_X1 U48176 ( .A1(n15794), .A2(n20060), .B(n35416), .ZN(n34363) );
  OAI21_X1 U48177 ( .A1(n34364), .A2(n15794), .B(n34363), .ZN(n34366) );
  AOI21_X1 U48178 ( .A1(n34369), .A2(n36046), .B(n34368), .ZN(n34370) );
  NAND2_X1 U48179 ( .A1(n34377), .A2(n10087), .ZN(n34373) );
  INV_X1 U48180 ( .I(n34374), .ZN(n34375) );
  NOR2_X1 U48181 ( .A1(n34375), .A2(n592), .ZN(n34376) );
  NOR3_X1 U48183 ( .A1(n10087), .A2(n34378), .A3(n37376), .ZN(n34379) );
  NOR3_X1 U48184 ( .A1(n34389), .A2(n34388), .A3(n34387), .ZN(n34390) );
  NAND2_X1 U48185 ( .A1(n34392), .A2(n59824), .ZN(n34393) );
  NOR2_X1 U48186 ( .A1(n35713), .A2(n15018), .ZN(n34394) );
  NAND2_X1 U48190 ( .A1(n35229), .A2(n34404), .ZN(n34403) );
  OAI22_X1 U48191 ( .A1(n34405), .A2(n34404), .B1(n34403), .B2(n58048), .ZN(
        n34406) );
  NAND2_X1 U48192 ( .A1(n34412), .A2(n35283), .ZN(n34419) );
  NAND3_X1 U48193 ( .A1(n35740), .A2(n35743), .A3(n10608), .ZN(n34416) );
  OAI21_X1 U48194 ( .A1(n64984), .A2(n34421), .B(n34420), .ZN(n34426) );
  NAND2_X1 U48195 ( .A1(n34426), .A2(n34425), .ZN(n34431) );
  NOR2_X1 U48196 ( .A1(n34427), .A2(n1544), .ZN(n34429) );
  OAI22_X1 U48197 ( .A1(n34429), .A2(n34428), .B1(n1806), .B2(n35783), .ZN(
        n34430) );
  NAND2_X1 U48198 ( .A1(n34432), .A2(n37355), .ZN(n34454) );
  OAI21_X1 U48199 ( .A1(n35255), .A2(n35759), .B(n59930), .ZN(n34436) );
  NAND2_X1 U48201 ( .A1(n34437), .A2(n35316), .ZN(n35257) );
  OAI21_X1 U48202 ( .A1(n34439), .A2(n34438), .B(n35257), .ZN(n34440) );
  NAND2_X1 U48203 ( .A1(n16402), .A2(n35762), .ZN(n35259) );
  NOR2_X1 U48204 ( .A1(n34443), .A2(n35646), .ZN(n34445) );
  NOR2_X1 U48205 ( .A1(n59005), .A2(n35643), .ZN(n34450) );
  AOI21_X1 U48206 ( .A1(n62995), .A2(n35652), .B(n34451), .ZN(n34452) );
  NOR2_X1 U48207 ( .A1(n37288), .A2(n4541), .ZN(n36756) );
  AOI21_X1 U48208 ( .A1(n34456), .A2(n34455), .B(n36755), .ZN(n34458) );
  NOR2_X1 U48209 ( .A1(n34828), .A2(n23626), .ZN(n34461) );
  INV_X1 U48211 ( .I(n34822), .ZN(n34465) );
  NAND2_X1 U48212 ( .A1(n37613), .A2(n37617), .ZN(n34466) );
  XOR2_X1 U48213 ( .A1(n43962), .A2(n55395), .Z(n51059) );
  XOR2_X1 U48214 ( .A1(n58077), .A2(n54776), .Z(n45088) );
  XOR2_X1 U48215 ( .A1(n34467), .A2(n45088), .Z(n51648) );
  XOR2_X1 U48216 ( .A1(n51059), .A2(n51648), .Z(n34468) );
  XOR2_X1 U48217 ( .A1(n37525), .A2(n34468), .Z(n34481) );
  INV_X1 U48219 ( .I(n34924), .ZN(n34470) );
  NAND2_X1 U48220 ( .A1(n34475), .A2(n21018), .ZN(n34476) );
  OAI22_X1 U48221 ( .A1(n35353), .A2(n34476), .B1(n35964), .B2(n35974), .ZN(
        n34477) );
  OAI22_X1 U48222 ( .A1(n34478), .A2(n35964), .B1(n35965), .B2(n35971), .ZN(
        n34479) );
  NAND2_X1 U48223 ( .A1(n34479), .A2(n1770), .ZN(n34480) );
  NAND2_X1 U48224 ( .A1(n34482), .A2(n36892), .ZN(n34483) );
  INV_X1 U48225 ( .I(n36946), .ZN(n34485) );
  XOR2_X1 U48226 ( .A1(n38168), .A2(n55833), .Z(n38333) );
  INV_X1 U48227 ( .I(n34878), .ZN(n34493) );
  XOR2_X1 U48228 ( .A1(n34495), .A2(n34496), .Z(n34809) );
  NOR2_X1 U48229 ( .A1(n34497), .A2(n34502), .ZN(n34498) );
  NAND3_X1 U48231 ( .A1(n60984), .A2(n24485), .A3(n35047), .ZN(n34637) );
  NAND4_X1 U48232 ( .A1(n34503), .A2(n35039), .A3(n34632), .A4(n34502), .ZN(
        n34505) );
  NOR2_X1 U48233 ( .A1(n34507), .A2(n1424), .ZN(n34508) );
  OAI21_X1 U48234 ( .A1(n1424), .A2(n63421), .B(n10091), .ZN(n34511) );
  NAND3_X1 U48235 ( .A1(n34513), .A2(n21008), .A3(n63444), .ZN(n34514) );
  INV_X1 U48236 ( .I(n34667), .ZN(n34519) );
  MUX2_X1 U48238 ( .I0(n36803), .I1(n36308), .S(n21605), .Z(n34574) );
  INV_X1 U48240 ( .I(n34526), .ZN(n34527) );
  NAND3_X1 U48242 ( .A1(n34539), .A2(n22419), .A3(n34538), .ZN(n34541) );
  NOR2_X1 U48245 ( .A1(n34558), .A2(n1543), .ZN(n34560) );
  OAI21_X1 U48246 ( .A1(n34571), .A2(n34570), .B(n34569), .ZN(n34573) );
  OAI21_X1 U48247 ( .A1(n34574), .A2(n36790), .B(n36309), .ZN(n34582) );
  NAND2_X2 U48249 ( .A1(n34582), .A2(n34581), .ZN(n39733) );
  NOR2_X1 U48250 ( .A1(n64234), .A2(n7453), .ZN(n34592) );
  OAI21_X1 U48251 ( .A1(n34596), .A2(n34590), .B(n34589), .ZN(n34591) );
  OAI21_X1 U48252 ( .A1(n34593), .A2(n34592), .B(n34591), .ZN(n34600) );
  NAND2_X1 U48253 ( .A1(n64618), .A2(n34604), .ZN(n34609) );
  NAND2_X1 U48254 ( .A1(n34607), .A2(n20946), .ZN(n34608) );
  AOI21_X1 U48255 ( .A1(n34626), .A2(n34618), .B(n12039), .ZN(n34620) );
  NAND3_X1 U48256 ( .A1(n9130), .A2(n34632), .A3(n34643), .ZN(n34633) );
  AOI21_X1 U48257 ( .A1(n34634), .A2(n34633), .B(n35038), .ZN(n34635) );
  NAND2_X1 U48258 ( .A1(n34637), .A2(n34636), .ZN(n34638) );
  AOI21_X1 U48259 ( .A1(n34642), .A2(n13068), .B(n34641), .ZN(n34645) );
  NAND2_X1 U48260 ( .A1(n60984), .A2(n34643), .ZN(n34644) );
  INV_X1 U48261 ( .I(n36858), .ZN(n34694) );
  NAND2_X1 U48262 ( .A1(n34665), .A2(n34664), .ZN(n34691) );
  NAND3_X1 U48263 ( .A1(n34667), .A2(n34670), .A3(n34666), .ZN(n34674) );
  NAND3_X1 U48264 ( .A1(n34668), .A2(n34670), .A3(n64461), .ZN(n34673) );
  NAND3_X1 U48265 ( .A1(n3467), .A2(n24083), .A3(n34679), .ZN(n34671) );
  NAND3_X1 U48267 ( .A1(n34680), .A2(n23400), .A3(n34679), .ZN(n34681) );
  NAND2_X1 U48268 ( .A1(n34682), .A2(n34681), .ZN(n34683) );
  INV_X1 U48271 ( .I(n36679), .ZN(n34697) );
  NAND2_X1 U48272 ( .A1(n60374), .A2(n61747), .ZN(n34696) );
  OAI21_X1 U48273 ( .A1(n34697), .A2(n34696), .B(n36850), .ZN(n34698) );
  INV_X1 U48274 ( .I(n35595), .ZN(n34701) );
  NAND3_X1 U48275 ( .A1(n34701), .A2(n36449), .A3(n34700), .ZN(n34706) );
  INV_X1 U48276 ( .I(n35162), .ZN(n34702) );
  NOR2_X1 U48277 ( .A1(n34702), .A2(n15038), .ZN(n34703) );
  AOI21_X1 U48278 ( .A1(n36454), .A2(n34703), .B(n57171), .ZN(n34705) );
  NAND2_X1 U48280 ( .A1(n34708), .A2(n35816), .ZN(n34709) );
  NAND3_X1 U48281 ( .A1(n34710), .A2(n35304), .A3(n34709), .ZN(n34711) );
  NAND2_X1 U48282 ( .A1(n15181), .A2(n34727), .ZN(n34723) );
  MUX2_X1 U48283 ( .I0(n15184), .I1(n34720), .S(n34719), .Z(n34722) );
  MUX2_X1 U48284 ( .I0(n34723), .I1(n34722), .S(n34721), .Z(n34732) );
  NAND2_X1 U48285 ( .A1(n34725), .A2(n15184), .ZN(n34724) );
  MUX2_X1 U48287 ( .I0(n34734), .I1(n23354), .S(n35301), .Z(n34735) );
  NOR2_X1 U48288 ( .A1(n34735), .A2(n35297), .ZN(n34738) );
  NAND4_X1 U48290 ( .A1(n35299), .A2(n21056), .A3(n35294), .A4(n31976), .ZN(
        n34744) );
  NOR2_X1 U48291 ( .A1(n34740), .A2(n64812), .ZN(n34742) );
  INV_X1 U48292 ( .I(n34748), .ZN(n34749) );
  OAI22_X1 U48294 ( .A1(n34760), .A2(n34759), .B1(n34758), .B2(n34764), .ZN(
        n34769) );
  AOI21_X1 U48295 ( .A1(n57619), .A2(n34761), .B(n34771), .ZN(n34767) );
  NAND2_X1 U48296 ( .A1(n34763), .A2(n64304), .ZN(n34765) );
  OAI22_X1 U48297 ( .A1(n34767), .A2(n60738), .B1(n34765), .B2(n34764), .ZN(
        n34768) );
  NAND2_X1 U48298 ( .A1(n57619), .A2(n34771), .ZN(n34773) );
  AOI21_X1 U48299 ( .A1(n34783), .A2(n61256), .B(n34781), .ZN(n34785) );
  NAND4_X1 U48300 ( .A1(n34790), .A2(n34798), .A3(n35001), .A4(n34789), .ZN(
        n34793) );
  NAND3_X1 U48301 ( .A1(n34795), .A2(n65119), .A3(n34796), .ZN(n34802) );
  NAND2_X1 U48303 ( .A1(n34804), .A2(n59147), .ZN(n34805) );
  NAND2_X1 U48304 ( .A1(n21489), .A2(n2418), .ZN(n34934) );
  NAND2_X1 U48308 ( .A1(n34823), .A2(n5317), .ZN(n34820) );
  INV_X1 U48309 ( .I(n35571), .ZN(n34826) );
  OAI21_X1 U48312 ( .A1(n35387), .A2(n60891), .B(n34828), .ZN(n34830) );
  NOR3_X1 U48313 ( .A1(n36040), .A2(n576), .A3(n4802), .ZN(n34829) );
  XOR2_X1 U48314 ( .A1(n34833), .A2(n50551), .Z(n49877) );
  XOR2_X1 U48315 ( .A1(n54407), .A2(n59638), .Z(n50885) );
  XOR2_X1 U48316 ( .A1(n50885), .A2(n56335), .Z(n34835) );
  MUX2_X1 U48317 ( .I0(n34838), .I1(n34837), .S(n7270), .Z(n34840) );
  NOR3_X1 U48319 ( .A1(n36778), .A2(n18496), .A3(n63838), .ZN(n34839) );
  NAND2_X1 U48320 ( .A1(n37271), .A2(n57860), .ZN(n34845) );
  NOR2_X1 U48321 ( .A1(n58580), .A2(n37268), .ZN(n34842) );
  NOR2_X1 U48322 ( .A1(n37490), .A2(n23842), .ZN(n34848) );
  AOI22_X1 U48323 ( .A1(n18983), .A2(n23471), .B1(n34848), .B2(n37270), .ZN(
        n34850) );
  NOR3_X1 U48324 ( .A1(n36050), .A2(n17096), .A3(n34854), .ZN(n34856) );
  MUX2_X1 U48325 ( .I0(n34857), .I1(n36050), .S(n7028), .Z(n34858) );
  INV_X1 U48327 ( .I(n35489), .ZN(n34864) );
  NAND2_X1 U48329 ( .A1(n1779), .A2(n1788), .ZN(n34869) );
  NOR2_X1 U48330 ( .A1(n34874), .A2(n35888), .ZN(n34870) );
  NAND2_X1 U48332 ( .A1(n35885), .A2(n10596), .ZN(n34879) );
  NOR3_X1 U48335 ( .A1(n36252), .A2(n19231), .A3(n35182), .ZN(n34890) );
  INV_X1 U48336 ( .I(n59396), .ZN(n34887) );
  NAND4_X1 U48338 ( .A1(n10067), .A2(n61223), .A3(n34887), .A4(n36249), .ZN(
        n34888) );
  INV_X1 U48340 ( .I(n35984), .ZN(n34892) );
  OAI21_X1 U48341 ( .A1(n34892), .A2(n35350), .B(n34891), .ZN(n34894) );
  NAND2_X1 U48344 ( .A1(n36698), .A2(n10849), .ZN(n34897) );
  NAND2_X1 U48345 ( .A1(n35426), .A2(n64101), .ZN(n34902) );
  NAND2_X1 U48346 ( .A1(n34907), .A2(n64101), .ZN(n34909) );
  NOR2_X1 U48347 ( .A1(n34912), .A2(n35432), .ZN(n34919) );
  NOR2_X1 U48348 ( .A1(n16337), .A2(n22993), .ZN(n34913) );
  NOR2_X1 U48349 ( .A1(n35430), .A2(n34913), .ZN(n34917) );
  NAND2_X1 U48350 ( .A1(n35427), .A2(n36944), .ZN(n36937) );
  INV_X1 U48351 ( .I(n36937), .ZN(n34916) );
  NAND2_X1 U48352 ( .A1(n34914), .A2(n35431), .ZN(n34915) );
  NAND2_X1 U48353 ( .A1(n35506), .A2(n34926), .ZN(n34923) );
  NAND2_X1 U48355 ( .A1(n1418), .A2(n1310), .ZN(n34932) );
  NAND2_X1 U48356 ( .A1(n26243), .A2(n21467), .ZN(n34931) );
  NAND3_X1 U48357 ( .A1(n34932), .A2(n64679), .A3(n34931), .ZN(n34933) );
  AOI21_X1 U48358 ( .A1(n26243), .A2(n34934), .B(n34933), .ZN(n34940) );
  NOR2_X1 U48362 ( .A1(n34947), .A2(n34952), .ZN(n34949) );
  OAI21_X1 U48363 ( .A1(n34971), .A2(n34970), .B(n34969), .ZN(n34978) );
  INV_X1 U48364 ( .I(n57423), .ZN(n34977) );
  NAND3_X1 U48365 ( .A1(n34981), .A2(n1424), .A3(n34980), .ZN(n34984) );
  INV_X1 U48367 ( .I(n35004), .ZN(n34999) );
  OAI21_X1 U48373 ( .A1(n35047), .A2(n35046), .B(n35045), .ZN(n35048) );
  NAND2_X1 U48374 ( .A1(n35049), .A2(n35048), .ZN(n35050) );
  XOR2_X1 U48376 ( .A1(n57448), .A2(n35075), .Z(n35076) );
  MUX2_X1 U48377 ( .I0(n35077), .I1(n37313), .S(n65236), .Z(n35085) );
  NAND2_X1 U48379 ( .A1(n35086), .A2(n22936), .ZN(n37311) );
  NOR4_X1 U48382 ( .A1(n22223), .A2(n37085), .A3(n4745), .A4(n37084), .ZN(
        n35082) );
  NOR2_X1 U48384 ( .A1(n35994), .A2(n37049), .ZN(n35093) );
  NOR3_X1 U48385 ( .A1(n35093), .A2(n63469), .A3(n37050), .ZN(n35094) );
  INV_X1 U48386 ( .I(n35991), .ZN(n35099) );
  NAND2_X1 U48387 ( .A1(n35095), .A2(n35096), .ZN(n35098) );
  NAND3_X1 U48388 ( .A1(n62010), .A2(n63469), .A3(n35096), .ZN(n35097) );
  OAI22_X1 U48389 ( .A1(n35099), .A2(n35098), .B1(n35482), .B2(n35097), .ZN(
        n35102) );
  NAND3_X1 U48390 ( .A1(n1793), .A2(n35994), .A3(n37049), .ZN(n37964) );
  OAI21_X1 U48391 ( .A1(n37044), .A2(n35482), .B(n37964), .ZN(n35101) );
  NOR2_X1 U48392 ( .A1(n35102), .A2(n35101), .ZN(n35108) );
  NAND2_X1 U48394 ( .A1(n37050), .A2(n63469), .ZN(n35989) );
  INV_X1 U48395 ( .I(n35989), .ZN(n35104) );
  INV_X1 U48397 ( .I(n35109), .ZN(n35110) );
  NAND4_X1 U48398 ( .A1(n36412), .A2(n35111), .A3(n35110), .A4(n10601), .ZN(
        n35112) );
  NAND2_X1 U48399 ( .A1(n36404), .A2(n16851), .ZN(n35116) );
  NOR2_X1 U48400 ( .A1(n36413), .A2(n35361), .ZN(n35119) );
  NAND3_X1 U48401 ( .A1(n36412), .A2(n36110), .A3(n35361), .ZN(n35117) );
  NAND2_X1 U48402 ( .A1(n23503), .A2(n22474), .ZN(n35121) );
  NAND2_X1 U48406 ( .A1(n1227), .A2(n35130), .ZN(n35131) );
  NAND3_X1 U48407 ( .A1(n59468), .A2(n3458), .A3(n22169), .ZN(n35132) );
  NAND4_X1 U48408 ( .A1(n35134), .A2(n35133), .A3(n21801), .A4(n35132), .ZN(
        n35135) );
  NAND2_X1 U48409 ( .A1(n35548), .A2(n35965), .ZN(n35137) );
  NAND3_X1 U48413 ( .A1(n35543), .A2(n35966), .A3(n35974), .ZN(n35149) );
  NOR2_X1 U48417 ( .A1(n36221), .A2(n1531), .ZN(n35161) );
  MUX2_X1 U48421 ( .I0(n35180), .I1(n35179), .S(n36262), .Z(n35187) );
  OAI21_X1 U48422 ( .A1(n948), .A2(n63897), .B(n36259), .ZN(n35186) );
  INV_X1 U48423 ( .I(n35181), .ZN(n35185) );
  INV_X1 U48424 ( .I(n36261), .ZN(n35184) );
  NOR2_X1 U48425 ( .A1(n36554), .A2(n36098), .ZN(n35190) );
  INV_X1 U48426 ( .I(n36092), .ZN(n35189) );
  AOI22_X1 U48427 ( .A1(n35190), .A2(n36561), .B1(n35189), .B2(n8356), .ZN(
        n35192) );
  NAND4_X1 U48428 ( .A1(n36574), .A2(n36565), .A3(n22785), .A4(n36566), .ZN(
        n35191) );
  XOR2_X1 U48429 ( .A1(n24147), .A2(n38784), .Z(n35194) );
  NAND3_X1 U48432 ( .A1(n7342), .A2(n19373), .A3(n35204), .ZN(n35205) );
  NAND2_X1 U48435 ( .A1(n35225), .A2(n35224), .ZN(n35226) );
  NAND2_X1 U48436 ( .A1(n35834), .A2(n35833), .ZN(n35231) );
  AOI21_X1 U48437 ( .A1(n57492), .A2(n35229), .B(n15018), .ZN(n35230) );
  OAI21_X1 U48439 ( .A1(n35712), .A2(n35833), .B(n15018), .ZN(n35233) );
  NAND2_X1 U48441 ( .A1(n35654), .A2(n60835), .ZN(n35243) );
  NOR2_X1 U48442 ( .A1(n62683), .A2(n58598), .ZN(n35242) );
  NAND2_X1 U48446 ( .A1(n63220), .A2(n35255), .ZN(n35256) );
  NAND3_X1 U48447 ( .A1(n35260), .A2(n59930), .A3(n35322), .ZN(n35261) );
  INV_X1 U48448 ( .I(n36332), .ZN(n36325) );
  NAND4_X1 U48449 ( .A1(n35794), .A2(n11182), .A3(n35272), .A4(n35799), .ZN(
        n35275) );
  OAI21_X1 U48451 ( .A1(n35807), .A2(n20736), .B(n35802), .ZN(n35277) );
  NAND2_X1 U48452 ( .A1(n35287), .A2(n904), .ZN(n35288) );
  NAND3_X1 U48453 ( .A1(n35288), .A2(n63329), .A3(n10608), .ZN(n35289) );
  NOR2_X1 U48454 ( .A1(n35316), .A2(n35758), .ZN(n35313) );
  NAND2_X1 U48455 ( .A1(n10503), .A2(n35316), .ZN(n35317) );
  NOR2_X1 U48456 ( .A1(n35320), .A2(n35755), .ZN(n35319) );
  OAI22_X1 U48457 ( .A1(n35324), .A2(n35778), .B1(n35775), .B2(n60152), .ZN(
        n35328) );
  OAI21_X1 U48458 ( .A1(n35331), .A2(n35330), .B(n64984), .ZN(n35334) );
  NAND3_X1 U48460 ( .A1(n36864), .A2(n1413), .A3(n62720), .ZN(n35337) );
  NAND2_X1 U48462 ( .A1(n35930), .A2(n1413), .ZN(n35336) );
  INV_X1 U48469 ( .I(n50798), .ZN(n35358) );
  AOI22_X1 U48470 ( .A1(n35360), .A2(n9984), .B1(n36196), .B2(n36413), .ZN(
        n35366) );
  INV_X1 U48471 ( .I(n36119), .ZN(n35362) );
  NAND2_X1 U48472 ( .A1(n36185), .A2(n9984), .ZN(n35364) );
  INV_X1 U48473 ( .I(n38309), .ZN(n35367) );
  XOR2_X1 U48474 ( .A1(n37730), .A2(n35372), .Z(n35373) );
  XOR2_X1 U48475 ( .A1(n45130), .A2(n35373), .Z(n51669) );
  XNOR2_X1 U48476 ( .A1(n23989), .A2(n52317), .ZN(n35375) );
  XOR2_X1 U48477 ( .A1(n52294), .A2(n53064), .Z(n35374) );
  XOR2_X1 U48478 ( .A1(n35375), .A2(n35374), .Z(n51088) );
  XOR2_X1 U48479 ( .A1(n51669), .A2(n51088), .Z(n35376) );
  XOR2_X1 U48480 ( .A1(n38916), .A2(n35376), .Z(n35377) );
  NAND2_X1 U48481 ( .A1(n18144), .A2(n65075), .ZN(n35378) );
  NOR2_X1 U48482 ( .A1(n36548), .A2(n35382), .ZN(n35380) );
  NAND2_X1 U48483 ( .A1(n35382), .A2(n36384), .ZN(n36894) );
  NAND4_X1 U48484 ( .A1(n36894), .A2(n36895), .A3(n35384), .A4(n7103), .ZN(
        n35385) );
  NOR2_X1 U48485 ( .A1(n35581), .A2(n576), .ZN(n35390) );
  NAND2_X1 U48486 ( .A1(n35569), .A2(n35391), .ZN(n35392) );
  NAND3_X2 U48487 ( .A1(n35394), .A2(n35393), .A3(n35392), .ZN(n38535) );
  INV_X1 U48488 ( .I(n36794), .ZN(n35400) );
  NAND2_X1 U48489 ( .A1(n36133), .A2(n35400), .ZN(n35402) );
  INV_X1 U48490 ( .I(n36131), .ZN(n35401) );
  INV_X1 U48494 ( .I(n35497), .ZN(n35409) );
  NOR3_X1 U48495 ( .A1(n35494), .A2(n61747), .A3(n36673), .ZN(n35410) );
  INV_X1 U48496 ( .I(n36774), .ZN(n36771) );
  NOR2_X1 U48497 ( .A1(n35422), .A2(n1417), .ZN(n35424) );
  INV_X1 U48498 ( .I(n35433), .ZN(n35434) );
  INV_X1 U48499 ( .I(n36279), .ZN(n35436) );
  NAND2_X1 U48501 ( .A1(n35437), .A2(n59852), .ZN(n35438) );
  NOR2_X1 U48505 ( .A1(n36534), .A2(n35455), .ZN(n35458) );
  NOR2_X1 U48506 ( .A1(n36386), .A2(n65075), .ZN(n35456) );
  AOI21_X1 U48507 ( .A1(n19206), .A2(n36535), .B(n36532), .ZN(n35459) );
  NOR2_X1 U48508 ( .A1(n35460), .A2(n35459), .ZN(n35461) );
  NOR2_X1 U48510 ( .A1(n36705), .A2(n35472), .ZN(n35473) );
  OAI21_X1 U48516 ( .A1(n35908), .A2(n35486), .B(n7598), .ZN(n35487) );
  MUX2_X1 U48518 ( .I0(n36850), .I1(n35493), .S(n61747), .Z(n35496) );
  NOR2_X1 U48519 ( .A1(n23146), .A2(n4754), .ZN(n35495) );
  XOR2_X1 U48520 ( .A1(n36851), .A2(n26213), .Z(n35499) );
  NOR2_X1 U48521 ( .A1(n35499), .A2(n61747), .ZN(n35500) );
  INV_X1 U48522 ( .I(n35511), .ZN(n35514) );
  INV_X1 U48524 ( .I(n36910), .ZN(n35513) );
  NAND3_X1 U48525 ( .A1(n35514), .A2(n35513), .A3(n35512), .ZN(n35519) );
  NOR2_X1 U48526 ( .A1(n22461), .A2(n37424), .ZN(n35515) );
  AOI22_X1 U48527 ( .A1(n37423), .A2(n35517), .B1(n35516), .B2(n35515), .ZN(
        n35518) );
  XOR2_X1 U48528 ( .A1(n22458), .A2(n38653), .Z(n35522) );
  XOR2_X1 U48529 ( .A1(n35522), .A2(n35521), .Z(n52152) );
  XOR2_X1 U48530 ( .A1(n35523), .A2(n55335), .Z(n50641) );
  XOR2_X1 U48531 ( .A1(n56827), .A2(n54870), .Z(n52149) );
  XOR2_X1 U48532 ( .A1(n52149), .A2(n132), .Z(n35524) );
  XOR2_X1 U48533 ( .A1(n50641), .A2(n35524), .Z(n35525) );
  XOR2_X1 U48534 ( .A1(n52152), .A2(n35525), .Z(n35541) );
  AOI22_X1 U48538 ( .A1(n35528), .A2(n57443), .B1(n35526), .B2(n9273), .ZN(
        n35530) );
  NAND2_X1 U48541 ( .A1(n35965), .A2(n15754), .ZN(n35546) );
  AOI21_X1 U48542 ( .A1(n35561), .A2(n35883), .B(n1779), .ZN(n35562) );
  NOR2_X1 U48543 ( .A1(n685), .A2(n35564), .ZN(n35566) );
  NAND2_X1 U48547 ( .A1(n35576), .A2(n36021), .ZN(n35577) );
  INV_X1 U48550 ( .I(n35591), .ZN(n35593) );
  OAI21_X1 U48551 ( .A1(n35593), .A2(n35592), .B(n9633), .ZN(n35594) );
  NOR2_X1 U48552 ( .A1(n23257), .A2(n36436), .ZN(n36225) );
  NOR2_X1 U48554 ( .A1(n19231), .A2(n35602), .ZN(n35603) );
  AOI21_X1 U48555 ( .A1(n35608), .A2(n1310), .B(n2418), .ZN(n35609) );
  NAND2_X1 U48557 ( .A1(n35612), .A2(n32684), .ZN(n35613) );
  NAND3_X1 U48558 ( .A1(n35619), .A2(n35614), .A3(n35613), .ZN(n35615) );
  OAI22_X1 U48560 ( .A1(n35619), .A2(n35618), .B1(n1811), .B2(n35617), .ZN(
        n35621) );
  OAI21_X1 U48561 ( .A1(n35622), .A2(n35621), .B(n35620), .ZN(n35639) );
  AOI21_X1 U48562 ( .A1(n35624), .A2(n59134), .B(n22428), .ZN(n35626) );
  NOR2_X1 U48563 ( .A1(n35626), .A2(n35625), .ZN(n35627) );
  NOR2_X1 U48564 ( .A1(n7342), .A2(n35628), .ZN(n35634) );
  INV_X1 U48566 ( .I(n35648), .ZN(n35649) );
  NAND2_X1 U48567 ( .A1(n35654), .A2(n35653), .ZN(n35657) );
  NAND3_X1 U48568 ( .A1(n35660), .A2(n35659), .A3(n35658), .ZN(n35661) );
  OAI22_X1 U48569 ( .A1(n35664), .A2(n35663), .B1(n6979), .B2(n35662), .ZN(
        n35665) );
  NOR3_X1 U48572 ( .A1(n35688), .A2(n10682), .A3(n35687), .ZN(n35689) );
  NOR2_X1 U48573 ( .A1(n35690), .A2(n35689), .ZN(n35697) );
  NAND3_X1 U48574 ( .A1(n63273), .A2(n11061), .A3(n24688), .ZN(n35696) );
  AOI22_X1 U48575 ( .A1(n35697), .A2(n35696), .B1(n35695), .B2(n35694), .ZN(
        n35698) );
  NAND2_X1 U48577 ( .A1(n35842), .A2(n35712), .ZN(n35718) );
  NAND2_X1 U48578 ( .A1(n35713), .A2(n15018), .ZN(n35714) );
  NAND3_X1 U48582 ( .A1(n36991), .A2(n23357), .A3(n37211), .ZN(n35726) );
  INV_X1 U48583 ( .I(n36613), .ZN(n35724) );
  NAND2_X1 U48584 ( .A1(n35724), .A2(n37212), .ZN(n35725) );
  NOR2_X1 U48585 ( .A1(n36618), .A2(n60431), .ZN(n35728) );
  INV_X1 U48586 ( .I(n35729), .ZN(n35734) );
  NAND2_X1 U48588 ( .A1(n35731), .A2(n60819), .ZN(n35732) );
  NOR2_X1 U48590 ( .A1(n10566), .A2(n35738), .ZN(n35739) );
  OAI22_X1 U48594 ( .A1(n10503), .A2(n35759), .B1(n59930), .B2(n35758), .ZN(
        n35760) );
  NAND2_X1 U48595 ( .A1(n35761), .A2(n35760), .ZN(n35767) );
  NAND2_X1 U48596 ( .A1(n35769), .A2(n1544), .ZN(n35772) );
  NAND3_X1 U48597 ( .A1(n35769), .A2(n58231), .A3(n64984), .ZN(n35771) );
  INV_X1 U48598 ( .I(n35773), .ZN(n35781) );
  OAI21_X1 U48599 ( .A1(n35781), .A2(n35780), .B(n35779), .ZN(n35791) );
  OAI22_X1 U48600 ( .A1(n35787), .A2(n35786), .B1(n60152), .B2(n35785), .ZN(
        n35788) );
  NAND2_X1 U48601 ( .A1(n10448), .A2(n18489), .ZN(n35797) );
  INV_X1 U48602 ( .I(n35795), .ZN(n35796) );
  NAND2_X1 U48603 ( .A1(n10448), .A2(n5099), .ZN(n35800) );
  NAND2_X1 U48604 ( .A1(n35803), .A2(n35802), .ZN(n35804) );
  NAND2_X1 U48605 ( .A1(n35807), .A2(n1805), .ZN(n35808) );
  NAND2_X1 U48608 ( .A1(n35817), .A2(n35816), .ZN(n35819) );
  NOR2_X1 U48611 ( .A1(n1309), .A2(n461), .ZN(n35832) );
  OAI21_X1 U48613 ( .A1(n35835), .A2(n35834), .B(n15018), .ZN(n35836) );
  AND2_X1 U48614 ( .A1(n35840), .A2(n35839), .Z(n35850) );
  INV_X1 U48615 ( .I(n35841), .ZN(n35845) );
  NAND2_X1 U48619 ( .A1(n36340), .A2(n36749), .ZN(n35856) );
  OAI21_X1 U48621 ( .A1(n36740), .A2(n20720), .B(n36340), .ZN(n35862) );
  NOR2_X1 U48622 ( .A1(n1417), .A2(n36749), .ZN(n35861) );
  XOR2_X1 U48624 ( .A1(n37868), .A2(n56322), .Z(n50502) );
  XOR2_X1 U48625 ( .A1(n44112), .A2(n50502), .Z(n52451) );
  XOR2_X1 U48626 ( .A1(n52451), .A2(n35869), .Z(n35870) );
  XOR2_X1 U48627 ( .A1(n38433), .A2(n35870), .Z(n35879) );
  NOR2_X1 U48628 ( .A1(n37190), .A2(n6779), .ZN(n35874) );
  NAND2_X1 U48629 ( .A1(n10226), .A2(n37327), .ZN(n35871) );
  XOR2_X1 U48630 ( .A1(n38577), .A2(n35879), .Z(n35912) );
  NAND2_X1 U48633 ( .A1(n35885), .A2(n35887), .ZN(n35890) );
  XOR2_X1 U48634 ( .A1(n21010), .A2(n25671), .Z(n35902) );
  NOR3_X1 U48635 ( .A1(n36825), .A2(n8195), .A3(n24041), .ZN(n35917) );
  AOI21_X1 U48638 ( .A1(n21881), .A2(n5873), .B(n35925), .ZN(n35926) );
  NAND3_X1 U48640 ( .A1(n35932), .A2(n5873), .A3(n25964), .ZN(n35933) );
  NAND2_X1 U48641 ( .A1(n21921), .A2(n8520), .ZN(n35934) );
  NOR2_X1 U48642 ( .A1(n37436), .A2(n35937), .ZN(n35940) );
  NAND2_X1 U48643 ( .A1(n35938), .A2(n37424), .ZN(n35939) );
  NAND2_X1 U48645 ( .A1(n35945), .A2(n35944), .ZN(n35948) );
  MUX2_X1 U48646 ( .I0(n35952), .I1(n35951), .S(n63406), .Z(n35955) );
  XOR2_X1 U48647 ( .A1(n23790), .A2(n61949), .Z(n35956) );
  INV_X1 U48648 ( .I(n35961), .ZN(n35963) );
  NOR2_X1 U48649 ( .A1(n35963), .A2(n35962), .ZN(n35969) );
  OAI22_X1 U48650 ( .A1(n35969), .A2(n35968), .B1(n62026), .B2(n35967), .ZN(
        n35978) );
  OAI22_X1 U48651 ( .A1(n35991), .A2(n22892), .B1(n35989), .B2(n15582), .ZN(
        n35992) );
  NAND2_X1 U48652 ( .A1(n35993), .A2(n35992), .ZN(n36007) );
  NOR2_X1 U48655 ( .A1(n37052), .A2(n37055), .ZN(n36004) );
  NAND2_X1 U48656 ( .A1(n36001), .A2(n37049), .ZN(n36003) );
  NOR3_X1 U48657 ( .A1(n37051), .A2(n23778), .A3(n37050), .ZN(n36002) );
  XOR2_X1 U48658 ( .A1(n22961), .A2(n36008), .Z(n46246) );
  XOR2_X1 U48659 ( .A1(n38145), .A2(n46246), .Z(n36018) );
  NAND2_X1 U48660 ( .A1(n36013), .A2(n7092), .ZN(n36011) );
  INV_X1 U48661 ( .I(n36019), .ZN(n36025) );
  NAND2_X1 U48662 ( .A1(n36027), .A2(n60891), .ZN(n36028) );
  NOR3_X1 U48663 ( .A1(n36031), .A2(n63484), .A3(n36040), .ZN(n36032) );
  NAND2_X1 U48664 ( .A1(n36038), .A2(n36037), .ZN(n36043) );
  OAI21_X1 U48665 ( .A1(n36043), .A2(n36042), .B(n36041), .ZN(n36044) );
  INV_X1 U48669 ( .I(n36531), .ZN(n36058) );
  NOR2_X1 U48671 ( .A1(n36394), .A2(n6440), .ZN(n36062) );
  NOR2_X1 U48676 ( .A1(n36308), .A2(n36138), .ZN(n36074) );
  MUX2_X1 U48678 ( .I0(n36076), .I1(n38550), .S(n37133), .Z(n36079) );
  NAND2_X1 U48680 ( .A1(n36082), .A2(n22733), .ZN(n36086) );
  NAND2_X1 U48683 ( .A1(n19364), .A2(n22785), .ZN(n36097) );
  NOR2_X1 U48685 ( .A1(n36098), .A2(n25261), .ZN(n36099) );
  OAI22_X1 U48686 ( .A1(n36101), .A2(n36100), .B1(n36099), .B2(n36566), .ZN(
        n36102) );
  NAND2_X1 U48687 ( .A1(n25570), .A2(n21736), .ZN(n38497) );
  NAND2_X1 U48690 ( .A1(n36119), .A2(n36118), .ZN(n36120) );
  NAND2_X1 U48692 ( .A1(n36124), .A2(n36169), .ZN(n36127) );
  NAND3_X1 U48693 ( .A1(n36135), .A2(n36804), .A3(n36134), .ZN(n36136) );
  XOR2_X1 U48696 ( .A1(n36145), .A2(n36736), .Z(n52320) );
  XOR2_X1 U48697 ( .A1(n51492), .A2(n53246), .Z(n36146) );
  XOR2_X1 U48698 ( .A1(n36147), .A2(n36146), .Z(n50577) );
  XOR2_X1 U48699 ( .A1(n52320), .A2(n50577), .Z(n36148) );
  INV_X1 U48700 ( .I(n36151), .ZN(n36149) );
  NAND2_X1 U48701 ( .A1(n36584), .A2(n36472), .ZN(n36153) );
  NAND2_X1 U48704 ( .A1(n36161), .A2(n36589), .ZN(n36162) );
  INV_X1 U48707 ( .I(n36508), .ZN(n36166) );
  INV_X1 U48708 ( .I(n36506), .ZN(n36165) );
  AOI21_X1 U48709 ( .A1(n36167), .A2(n36166), .B(n36165), .ZN(n36168) );
  AOI21_X1 U48710 ( .A1(n36423), .A2(n36170), .B(n36169), .ZN(n36174) );
  NAND2_X1 U48711 ( .A1(n36179), .A2(n3458), .ZN(n36181) );
  OAI21_X1 U48712 ( .A1(n36181), .A2(n36180), .B(n36420), .ZN(n36182) );
  NAND2_X1 U48713 ( .A1(n61936), .A2(n22474), .ZN(n36184) );
  NAND2_X1 U48714 ( .A1(n36188), .A2(n10601), .ZN(n36189) );
  NOR2_X1 U48715 ( .A1(n36404), .A2(n36193), .ZN(n36194) );
  NAND2_X1 U48716 ( .A1(n36201), .A2(n21467), .ZN(n36204) );
  NAND2_X1 U48717 ( .A1(n20867), .A2(n2418), .ZN(n36203) );
  NOR2_X1 U48718 ( .A1(n36207), .A2(n21467), .ZN(n36210) );
  XOR2_X1 U48720 ( .A1(n51234), .A2(n36215), .Z(n51604) );
  XOR2_X1 U48721 ( .A1(n55792), .A2(n4561), .Z(n36216) );
  XOR2_X1 U48722 ( .A1(n42790), .A2(n36216), .Z(n51485) );
  XOR2_X1 U48723 ( .A1(n46501), .A2(n56322), .Z(n36217) );
  XOR2_X1 U48724 ( .A1(n51485), .A2(n36217), .Z(n36218) );
  NOR2_X1 U48725 ( .A1(n36444), .A2(n36437), .ZN(n36228) );
  NOR3_X1 U48726 ( .A1(n36229), .A2(n22527), .A3(n36483), .ZN(n36231) );
  AOI21_X1 U48727 ( .A1(n36235), .A2(n36234), .B(n36494), .ZN(n36237) );
  NOR2_X1 U48728 ( .A1(n36238), .A2(n10829), .ZN(n36239) );
  NOR2_X1 U48729 ( .A1(n36244), .A2(n61770), .ZN(n36255) );
  AOI21_X1 U48730 ( .A1(n59396), .A2(n36246), .B(n36245), .ZN(n36248) );
  AOI21_X1 U48732 ( .A1(n36259), .A2(n62794), .B(n36258), .ZN(n36260) );
  OAI21_X1 U48734 ( .A1(n36265), .A2(n37218), .B(n37212), .ZN(n36268) );
  NAND2_X1 U48735 ( .A1(n37222), .A2(n37225), .ZN(n36266) );
  NAND4_X1 U48736 ( .A1(n36266), .A2(n37210), .A3(n37219), .A4(n23357), .ZN(
        n36267) );
  NOR2_X1 U48738 ( .A1(n57209), .A2(n1527), .ZN(n36272) );
  OAI21_X1 U48739 ( .A1(n36272), .A2(n36271), .B(n36628), .ZN(n36274) );
  NAND2_X1 U48741 ( .A1(n36275), .A2(n36365), .ZN(n36276) );
  OAI22_X1 U48743 ( .A1(n36627), .A2(n36279), .B1(n63643), .B2(n36962), .ZN(
        n36283) );
  NAND3_X1 U48744 ( .A1(n1530), .A2(n36959), .A3(n1781), .ZN(n36280) );
  AOI21_X1 U48745 ( .A1(n36281), .A2(n36280), .B(n60694), .ZN(n36282) );
  XOR2_X1 U48746 ( .A1(n38848), .A2(n58235), .Z(n36660) );
  XOR2_X1 U48747 ( .A1(n36660), .A2(n22698), .Z(n37147) );
  INV_X1 U48748 ( .I(n37115), .ZN(n36287) );
  INV_X1 U48749 ( .I(n37113), .ZN(n36290) );
  NOR2_X1 U48751 ( .A1(n37111), .A2(n22659), .ZN(n36293) );
  NAND2_X1 U48752 ( .A1(n36794), .A2(n21605), .ZN(n36303) );
  INV_X1 U48753 ( .I(n36300), .ZN(n36302) );
  XOR2_X1 U48758 ( .A1(n36318), .A2(n44808), .Z(n50573) );
  XOR2_X1 U48759 ( .A1(n36320), .A2(n36319), .Z(n52365) );
  XOR2_X1 U48760 ( .A1(n50573), .A2(n52365), .Z(n36321) );
  OAI21_X1 U48761 ( .A1(n36325), .A2(n37400), .B(n36834), .ZN(n36326) );
  NAND3_X1 U48762 ( .A1(n36327), .A2(n17660), .A3(n37404), .ZN(n36328) );
  NAND2_X1 U48764 ( .A1(n36345), .A2(n36344), .ZN(n36346) );
  NOR2_X1 U48765 ( .A1(n37222), .A2(n59617), .ZN(n36350) );
  OAI21_X1 U48766 ( .A1(n37210), .A2(n58250), .B(n37225), .ZN(n36351) );
  NAND3_X1 U48767 ( .A1(n36352), .A2(n37219), .A3(n36351), .ZN(n36353) );
  XOR2_X1 U48768 ( .A1(n39458), .A2(n55603), .Z(n50068) );
  XOR2_X1 U48769 ( .A1(n51194), .A2(n50067), .Z(n46373) );
  XOR2_X1 U48770 ( .A1(n50068), .A2(n46373), .Z(n36359) );
  INV_X1 U48771 ( .I(n36356), .ZN(n36358) );
  XOR2_X1 U48772 ( .A1(n36358), .A2(n36357), .Z(n50961) );
  XOR2_X1 U48773 ( .A1(n36359), .A2(n50961), .Z(n36360) );
  NOR2_X1 U48775 ( .A1(n59852), .A2(n1338), .ZN(n36361) );
  NAND2_X1 U48776 ( .A1(n36363), .A2(n57209), .ZN(n36364) );
  INV_X1 U48777 ( .I(n36628), .ZN(n36366) );
  INV_X1 U48779 ( .I(n62864), .ZN(n36368) );
  XOR2_X1 U48780 ( .A1(n36368), .A2(n39460), .Z(n38170) );
  NOR2_X1 U48782 ( .A1(n36384), .A2(n58888), .ZN(n36390) );
  NOR2_X1 U48788 ( .A1(n36395), .A2(n22454), .ZN(n36396) );
  NOR2_X1 U48790 ( .A1(n36402), .A2(n10601), .ZN(n36406) );
  AOI22_X1 U48791 ( .A1(n36407), .A2(n36406), .B1(n36405), .B2(n9984), .ZN(
        n36417) );
  NOR2_X1 U48792 ( .A1(n36412), .A2(n22474), .ZN(n36414) );
  OAI21_X1 U48793 ( .A1(n36415), .A2(n36414), .B(n36413), .ZN(n36416) );
  INV_X1 U48794 ( .I(n36418), .ZN(n36421) );
  OAI21_X1 U48795 ( .A1(n36421), .A2(n36420), .B(n36419), .ZN(n36425) );
  OAI21_X1 U48796 ( .A1(n36430), .A2(n36429), .B(n36428), .ZN(n36433) );
  NOR2_X1 U48797 ( .A1(n1531), .A2(n36434), .ZN(n36440) );
  NOR2_X1 U48798 ( .A1(n1531), .A2(n36441), .ZN(n36439) );
  NOR2_X1 U48799 ( .A1(n36441), .A2(n36444), .ZN(n36448) );
  OAI21_X1 U48800 ( .A1(n23257), .A2(n36446), .B(n36445), .ZN(n36447) );
  NOR2_X1 U48802 ( .A1(n36460), .A2(n36459), .ZN(n36461) );
  NAND4_X1 U48803 ( .A1(n36472), .A2(n36471), .A3(n11272), .A4(n22113), .ZN(
        n36464) );
  OAI21_X1 U48804 ( .A1(n63247), .A2(n36465), .B(n7933), .ZN(n36467) );
  INV_X1 U48805 ( .I(n36469), .ZN(n36475) );
  AOI22_X1 U48806 ( .A1(n932), .A2(n36478), .B1(n59379), .B2(n36476), .ZN(
        n36482) );
  INV_X1 U48807 ( .I(n36487), .ZN(n36488) );
  NOR2_X1 U48808 ( .A1(n36495), .A2(n36494), .ZN(n36497) );
  XOR2_X1 U48809 ( .A1(n23115), .A2(n50190), .Z(n36859) );
  NOR2_X1 U48810 ( .A1(n18525), .A2(n37376), .ZN(n36510) );
  NAND3_X1 U48812 ( .A1(n36515), .A2(n36514), .A3(n2589), .ZN(n36524) );
  NOR2_X1 U48813 ( .A1(n36587), .A2(n592), .ZN(n36519) );
  OAI21_X1 U48814 ( .A1(n36519), .A2(n36518), .B(n61704), .ZN(n36522) );
  XOR2_X1 U48815 ( .A1(n43789), .A2(n44796), .Z(n36525) );
  XOR2_X1 U48816 ( .A1(n37635), .A2(n36525), .Z(n50192) );
  XOR2_X1 U48817 ( .A1(n51275), .A2(n51946), .Z(n36526) );
  XOR2_X1 U48818 ( .A1(n50192), .A2(n36526), .Z(n36527) );
  XOR2_X1 U48819 ( .A1(n39307), .A2(n36527), .Z(n36528) );
  NOR2_X1 U48820 ( .A1(n18144), .A2(n59912), .ZN(n36530) );
  NOR2_X1 U48821 ( .A1(n36531), .A2(n36530), .ZN(n36552) );
  NOR2_X1 U48822 ( .A1(n36548), .A2(n36535), .ZN(n36537) );
  INV_X1 U48823 ( .I(n36539), .ZN(n36546) );
  AOI22_X1 U48824 ( .A1(n36543), .A2(n36542), .B1(n36541), .B2(n63273), .ZN(
        n36544) );
  XOR2_X1 U48826 ( .A1(n22785), .A2(n36555), .Z(n36556) );
  INV_X1 U48828 ( .I(n36564), .ZN(n36570) );
  NAND4_X1 U48829 ( .A1(n36568), .A2(n24102), .A3(n8356), .A4(n36566), .ZN(
        n36569) );
  OAI21_X1 U48831 ( .A1(n36574), .A2(n22785), .B(n36573), .ZN(n36578) );
  INV_X1 U48832 ( .I(n36575), .ZN(n36577) );
  INV_X1 U48834 ( .I(n36586), .ZN(n36593) );
  NOR2_X1 U48835 ( .A1(n36590), .A2(n36589), .ZN(n36591) );
  NOR3_X1 U48836 ( .A1(n10087), .A2(n22632), .A3(n60980), .ZN(n36599) );
  NOR3_X1 U48837 ( .A1(n36597), .A2(n36596), .A3(n60980), .ZN(n36598) );
  XOR2_X1 U48838 ( .A1(n37979), .A2(n24151), .Z(n39562) );
  NOR2_X1 U48839 ( .A1(n37212), .A2(n59617), .ZN(n36611) );
  OAI21_X1 U48840 ( .A1(n36611), .A2(n36610), .B(n18583), .ZN(n36614) );
  NOR2_X1 U48841 ( .A1(n37222), .A2(n37224), .ZN(n36617) );
  INV_X1 U48842 ( .I(n36620), .ZN(n36621) );
  NOR2_X1 U48843 ( .A1(n36959), .A2(n36623), .ZN(n36625) );
  XOR2_X1 U48845 ( .A1(n45130), .A2(n36630), .Z(n50028) );
  XNOR2_X1 U48846 ( .A1(n55862), .A2(n52294), .ZN(n36631) );
  XOR2_X1 U48847 ( .A1(n36632), .A2(n36631), .Z(n50970) );
  XOR2_X1 U48848 ( .A1(n61737), .A2(n60556), .Z(n36633) );
  XOR2_X1 U48849 ( .A1(n50970), .A2(n36633), .Z(n36634) );
  XOR2_X1 U48850 ( .A1(n50028), .A2(n36634), .Z(n36635) );
  XOR2_X1 U48851 ( .A1(n23280), .A2(n36635), .Z(n36636) );
  NOR2_X1 U48852 ( .A1(n4745), .A2(n37319), .ZN(n36641) );
  NOR2_X2 U48853 ( .A1(n36646), .A2(n36645), .ZN(n37556) );
  NAND3_X1 U48854 ( .A1(n38026), .A2(n13166), .A3(n9215), .ZN(n40237) );
  INV_X1 U48855 ( .I(n40237), .ZN(n36651) );
  NOR2_X1 U48856 ( .A1(n59199), .A2(n39415), .ZN(n36650) );
  XOR2_X1 U48857 ( .A1(n36656), .A2(n56859), .Z(n36657) );
  XOR2_X1 U48858 ( .A1(n36657), .A2(n38000), .Z(n50526) );
  XOR2_X1 U48859 ( .A1(n50878), .A2(n52399), .Z(n36658) );
  XOR2_X1 U48860 ( .A1(n18115), .A2(n36659), .Z(n36661) );
  INV_X1 U48861 ( .I(n36660), .ZN(n39767) );
  XOR2_X1 U48862 ( .A1(n36661), .A2(n39767), .Z(n36662) );
  XOR2_X1 U48863 ( .A1(n37418), .A2(n36662), .Z(n36686) );
  OAI21_X1 U48864 ( .A1(n36671), .A2(n36665), .B(n4754), .ZN(n36666) );
  NAND2_X1 U48865 ( .A1(n36852), .A2(n62920), .ZN(n36675) );
  INV_X1 U48866 ( .I(n36669), .ZN(n36670) );
  NAND2_X1 U48867 ( .A1(n36677), .A2(n61747), .ZN(n36678) );
  OAI21_X1 U48868 ( .A1(n36680), .A2(n36679), .B(n36678), .ZN(n36681) );
  NAND2_X1 U48871 ( .A1(n36689), .A2(n37395), .ZN(n36690) );
  INV_X1 U48872 ( .I(n37389), .ZN(n36692) );
  NAND3_X1 U48873 ( .A1(n36692), .A2(n1416), .A3(n8520), .ZN(n36693) );
  AOI21_X1 U48874 ( .A1(n60022), .A2(n652), .B(n15720), .ZN(n36696) );
  AOI21_X1 U48875 ( .A1(n36697), .A2(n36696), .B(n21584), .ZN(n36703) );
  OAI21_X1 U48876 ( .A1(n36698), .A2(n652), .B(n36706), .ZN(n36701) );
  OAI21_X1 U48877 ( .A1(n21584), .A2(n652), .B(n61517), .ZN(n36710) );
  NAND2_X1 U48878 ( .A1(n36710), .A2(n36709), .ZN(n36711) );
  NAND2_X1 U48879 ( .A1(n1766), .A2(n26243), .ZN(n36731) );
  NOR2_X1 U48880 ( .A1(n20867), .A2(n36716), .ZN(n36718) );
  NAND2_X1 U48881 ( .A1(n36725), .A2(n36724), .ZN(n36726) );
  INV_X1 U48882 ( .I(n46615), .ZN(n45829) );
  XOR2_X1 U48883 ( .A1(n36734), .A2(n45829), .Z(n50496) );
  XOR2_X1 U48884 ( .A1(n39375), .A2(n24014), .Z(n36735) );
  XOR2_X1 U48885 ( .A1(n36736), .A2(n36735), .Z(n52437) );
  XOR2_X1 U48886 ( .A1(n38388), .A2(n55516), .Z(n36737) );
  XOR2_X1 U48887 ( .A1(n52437), .A2(n36737), .Z(n36738) );
  XOR2_X1 U48888 ( .A1(n50496), .A2(n36738), .Z(n36739) );
  INV_X1 U48892 ( .I(n37291), .ZN(n36761) );
  INV_X1 U48893 ( .I(n36758), .ZN(n36759) );
  NOR2_X1 U48894 ( .A1(n17096), .A2(n3622), .ZN(n36767) );
  NOR2_X1 U48895 ( .A1(n36769), .A2(n20060), .ZN(n36770) );
  NAND2_X1 U48896 ( .A1(n63838), .A2(n38550), .ZN(n36779) );
  NOR2_X1 U48899 ( .A1(n26052), .A2(n38550), .ZN(n36785) );
  NAND2_X1 U48900 ( .A1(n38552), .A2(n36785), .ZN(n37477) );
  NOR2_X1 U48901 ( .A1(n37278), .A2(n16027), .ZN(n36788) );
  NAND2_X1 U48902 ( .A1(n36789), .A2(n36809), .ZN(n36791) );
  MUX2_X1 U48903 ( .I0(n36792), .I1(n36791), .S(n36790), .Z(n36817) );
  NOR4_X1 U48904 ( .A1(n36794), .A2(n57278), .A3(n60925), .A4(n36793), .ZN(
        n36799) );
  INV_X1 U48906 ( .I(n36808), .ZN(n36811) );
  INV_X1 U48907 ( .I(n36809), .ZN(n36810) );
  OAI21_X1 U48910 ( .A1(n36829), .A2(n8195), .B(n37400), .ZN(n36830) );
  AOI21_X1 U48914 ( .A1(n61747), .A2(n62942), .B(n60374), .ZN(n36857) );
  NOR2_X1 U48915 ( .A1(n7092), .A2(n26213), .ZN(n36854) );
  NAND4_X1 U48916 ( .A1(n36854), .A2(n7208), .A3(n36852), .A4(n61207), .ZN(
        n36855) );
  XOR2_X1 U48917 ( .A1(n57458), .A2(n36859), .Z(n36863) );
  INV_X1 U48918 ( .I(n51978), .ZN(n44325) );
  XOR2_X1 U48919 ( .A1(n9722), .A2(n51530), .Z(n38095) );
  XOR2_X1 U48920 ( .A1(n44325), .A2(n38095), .Z(n36861) );
  XOR2_X1 U48921 ( .A1(n36860), .A2(n56879), .Z(n51979) );
  XOR2_X1 U48922 ( .A1(n36861), .A2(n51979), .Z(n36862) );
  NAND2_X1 U48923 ( .A1(n36866), .A2(n36865), .ZN(n36867) );
  MUX2_X1 U48924 ( .I0(n36868), .I1(n36867), .S(n59924), .Z(n36881) );
  NOR2_X1 U48925 ( .A1(n25396), .A2(n4798), .ZN(n36871) );
  INV_X1 U48926 ( .I(n37064), .ZN(n36874) );
  NAND2_X1 U48933 ( .A1(n36939), .A2(n36946), .ZN(n36891) );
  INV_X1 U48934 ( .I(n36894), .ZN(n36897) );
  INV_X1 U48935 ( .I(n36900), .ZN(n36901) );
  INV_X1 U48936 ( .I(n36916), .ZN(n36906) );
  NOR2_X1 U48937 ( .A1(n36908), .A2(n37435), .ZN(n36912) );
  INV_X1 U48941 ( .I(n36923), .ZN(n36927) );
  XOR2_X1 U48942 ( .A1(n36929), .A2(n37651), .Z(n49822) );
  XOR2_X1 U48943 ( .A1(n36930), .A2(n23989), .Z(n50857) );
  XOR2_X1 U48944 ( .A1(n50857), .A2(n51150), .Z(n36931) );
  XOR2_X1 U48945 ( .A1(n49822), .A2(n36931), .Z(n36932) );
  XOR2_X1 U48946 ( .A1(n11534), .A2(n36932), .Z(n36933) );
  XOR2_X1 U48947 ( .A1(n36935), .A2(n36934), .Z(n36936) );
  NAND2_X1 U48949 ( .A1(n36967), .A2(n7074), .ZN(n36968) );
  INV_X1 U48950 ( .I(n36971), .ZN(n36972) );
  OAI21_X1 U48951 ( .A1(n37249), .A2(n461), .B(n36972), .ZN(n36974) );
  AOI21_X1 U48953 ( .A1(n37212), .A2(n37210), .B(n36990), .ZN(n36982) );
  NAND2_X1 U48954 ( .A1(n36980), .A2(n37225), .ZN(n36981) );
  XOR2_X1 U48957 ( .A1(n56702), .A2(n54168), .Z(n51392) );
  XOR2_X1 U48958 ( .A1(n51392), .A2(n15712), .Z(n37348) );
  XOR2_X1 U48960 ( .A1(n39275), .A2(n57162), .Z(n37382) );
  XOR2_X1 U48961 ( .A1(n38866), .A2(n54289), .Z(n39286) );
  XOR2_X1 U48962 ( .A1(n23020), .A2(n50787), .Z(n36997) );
  XOR2_X1 U48963 ( .A1(n39400), .A2(n36997), .Z(n49736) );
  XOR2_X1 U48964 ( .A1(n39279), .A2(n36998), .Z(n50866) );
  XOR2_X1 U48965 ( .A1(n49736), .A2(n50866), .Z(n36999) );
  XOR2_X1 U48966 ( .A1(n38168), .A2(n36999), .Z(n37000) );
  XOR2_X1 U48967 ( .A1(n39286), .A2(n37000), .Z(n37001) );
  INV_X1 U48968 ( .I(n37010), .ZN(n37013) );
  NOR2_X1 U48969 ( .A1(n37011), .A2(n37327), .ZN(n37012) );
  NOR2_X1 U48970 ( .A1(n37023), .A2(n37016), .ZN(n37021) );
  AOI22_X1 U48971 ( .A1(n37023), .A2(n37084), .B1(n23651), .B2(n37022), .ZN(
        n37024) );
  NOR2_X1 U48972 ( .A1(n37024), .A2(n37319), .ZN(n37025) );
  NAND2_X1 U48973 ( .A1(n37031), .A2(n37030), .ZN(n37032) );
  AOI21_X1 U48974 ( .A1(n37033), .A2(n37032), .B(n2699), .ZN(n37041) );
  NAND2_X1 U48975 ( .A1(n1773), .A2(n60659), .ZN(n37039) );
  NAND2_X1 U48977 ( .A1(n7598), .A2(n14904), .ZN(n37037) );
  OAI22_X1 U48978 ( .A1(n37039), .A2(n37038), .B1(n37037), .B2(n2699), .ZN(
        n37040) );
  NOR2_X1 U48979 ( .A1(n37041), .A2(n37040), .ZN(n37042) );
  NAND2_X1 U48980 ( .A1(n37050), .A2(n37049), .ZN(n37054) );
  AOI21_X1 U48981 ( .A1(n37052), .A2(n2483), .B(n37051), .ZN(n37053) );
  OAI21_X1 U48982 ( .A1(n37055), .A2(n37054), .B(n37053), .ZN(n37056) );
  NOR2_X1 U48984 ( .A1(n23752), .A2(n62681), .ZN(n37061) );
  XOR2_X1 U48986 ( .A1(n37073), .A2(n38653), .Z(n52109) );
  XOR2_X1 U48987 ( .A1(n52109), .A2(n44052), .Z(n37074) );
  XOR2_X1 U48988 ( .A1(n44299), .A2(n37074), .Z(n37075) );
  XOR2_X1 U48989 ( .A1(n22435), .A2(n37075), .Z(n37076) );
  XOR2_X1 U48990 ( .A1(n38903), .A2(n37076), .Z(n37077) );
  XOR2_X1 U48991 ( .A1(n37077), .A2(n23120), .Z(n37078) );
  XOR2_X1 U48992 ( .A1(n38430), .A2(n53272), .Z(n44211) );
  XOR2_X1 U48993 ( .A1(n44211), .A2(n37869), .Z(n50587) );
  XOR2_X1 U48994 ( .A1(n50746), .A2(n56495), .Z(n37079) );
  INV_X1 U48995 ( .I(n51234), .ZN(n43971) );
  XOR2_X1 U48996 ( .A1(n37079), .A2(n43971), .Z(n37080) );
  XOR2_X1 U48997 ( .A1(n50587), .A2(n37080), .Z(n37081) );
  XOR2_X1 U48998 ( .A1(n23062), .A2(n37081), .Z(n37082) );
  NAND3_X1 U49000 ( .A1(n1780), .A2(n37084), .A3(n37945), .ZN(n37087) );
  NOR2_X1 U49002 ( .A1(n37091), .A2(n37311), .ZN(n37093) );
  AOI21_X1 U49003 ( .A1(n37319), .A2(n37096), .B(n37095), .ZN(n37097) );
  XOR2_X1 U49005 ( .A1(n57836), .A2(n23898), .Z(n37101) );
  XOR2_X1 U49006 ( .A1(n37101), .A2(n37100), .Z(n37102) );
  INV_X1 U49007 ( .I(n37107), .ZN(n37108) );
  OAI21_X1 U49008 ( .A1(n37109), .A2(n37108), .B(n36288), .ZN(n37110) );
  XOR2_X1 U49009 ( .A1(n23115), .A2(n55889), .Z(n39755) );
  INV_X1 U49010 ( .I(n50987), .ZN(n37119) );
  XOR2_X1 U49011 ( .A1(n37119), .A2(n44796), .Z(n37120) );
  NAND2_X1 U49012 ( .A1(n37125), .A2(n37268), .ZN(n37127) );
  AOI21_X1 U49013 ( .A1(n37127), .A2(n37270), .B(n37126), .ZN(n37128) );
  NOR2_X1 U49014 ( .A1(n37129), .A2(n37128), .ZN(n37141) );
  NOR2_X1 U49015 ( .A1(n37277), .A2(n37131), .ZN(n37281) );
  OAI22_X1 U49018 ( .A1(n37136), .A2(n38550), .B1(n7270), .B2(n37135), .ZN(
        n37137) );
  XOR2_X1 U49020 ( .A1(n37143), .A2(n37142), .Z(n52051) );
  XOR2_X1 U49021 ( .A1(n45238), .A2(n54386), .Z(n50709) );
  XOR2_X1 U49022 ( .A1(n9826), .A2(n50709), .Z(n50776) );
  XOR2_X1 U49023 ( .A1(n52051), .A2(n50776), .Z(n37144) );
  XOR2_X1 U49024 ( .A1(n18049), .A2(n37144), .Z(n37145) );
  XOR2_X1 U49025 ( .A1(n51999), .A2(n37511), .Z(n37148) );
  XOR2_X1 U49026 ( .A1(n37148), .A2(n23493), .Z(n37150) );
  XOR2_X1 U49027 ( .A1(n39299), .A2(n17347), .Z(n37149) );
  XOR2_X1 U49028 ( .A1(n38596), .A2(n24927), .Z(n37151) );
  NAND2_X1 U49030 ( .A1(n61159), .A2(n40263), .ZN(n37196) );
  XOR2_X1 U49031 ( .A1(n39214), .A2(n54776), .Z(n38873) );
  XOR2_X1 U49032 ( .A1(n39406), .A2(n38873), .Z(n37157) );
  INV_X1 U49033 ( .I(n51817), .ZN(n37153) );
  XOR2_X1 U49034 ( .A1(n37520), .A2(n55903), .Z(n51137) );
  XOR2_X1 U49035 ( .A1(n51137), .A2(n51194), .Z(n37152) );
  XOR2_X1 U49036 ( .A1(n37153), .A2(n37152), .Z(n37154) );
  XOR2_X1 U49037 ( .A1(n62864), .A2(n37154), .Z(n37155) );
  XOR2_X1 U49038 ( .A1(n37155), .A2(n204), .Z(n37156) );
  XOR2_X1 U49039 ( .A1(n37157), .A2(n37156), .Z(n37160) );
  XOR2_X1 U49040 ( .A1(n37159), .A2(n58827), .Z(n39749) );
  NOR2_X1 U49041 ( .A1(n37455), .A2(n12797), .ZN(n37164) );
  NAND2_X1 U49042 ( .A1(n61438), .A2(n22801), .ZN(n37163) );
  OAI21_X1 U49043 ( .A1(n37164), .A2(n37163), .B(n24033), .ZN(n37167) );
  NAND2_X1 U49044 ( .A1(n37234), .A2(n12797), .ZN(n37445) );
  NAND3_X1 U49045 ( .A1(n37445), .A2(n37249), .A3(n37233), .ZN(n37166) );
  AOI22_X1 U49046 ( .A1(n37249), .A2(n9869), .B1(n24033), .B2(n37233), .ZN(
        n37165) );
  NAND2_X1 U49048 ( .A1(n909), .A2(n37168), .ZN(n37169) );
  XOR2_X1 U49049 ( .A1(n38457), .A2(n37385), .Z(n37172) );
  XOR2_X1 U49050 ( .A1(n37979), .A2(n37174), .Z(n37175) );
  XOR2_X1 U49052 ( .A1(n44427), .A2(n53064), .Z(n37176) );
  XOR2_X1 U49053 ( .A1(n44094), .A2(n37176), .Z(n51205) );
  XOR2_X1 U49054 ( .A1(n52196), .A2(n56849), .Z(n37177) );
  XOR2_X1 U49055 ( .A1(n51205), .A2(n37177), .Z(n37178) );
  XOR2_X1 U49056 ( .A1(n38916), .A2(n37178), .Z(n37179) );
  XOR2_X1 U49057 ( .A1(n37179), .A2(n23927), .Z(n37180) );
  NAND3_X1 U49059 ( .A1(n37183), .A2(n37182), .A3(n62734), .ZN(n37185) );
  XOR2_X1 U49061 ( .A1(n37556), .A2(n22988), .Z(n38253) );
  NOR3_X1 U49062 ( .A1(n40471), .A2(n9969), .A3(n40463), .ZN(n37203) );
  NOR2_X1 U49064 ( .A1(n40257), .A2(n9969), .ZN(n37200) );
  INV_X1 U49069 ( .I(n37209), .ZN(n37214) );
  NOR2_X1 U49071 ( .A1(n23357), .A2(n3691), .ZN(n37229) );
  NAND2_X1 U49074 ( .A1(n461), .A2(n37233), .ZN(n37235) );
  NAND4_X1 U49075 ( .A1(n37235), .A2(n37249), .A3(n12797), .A4(n22801), .ZN(
        n37239) );
  MUX2_X1 U49077 ( .I0(n37239), .I1(n37238), .S(n37237), .Z(n37246) );
  NAND4_X1 U49081 ( .A1(n909), .A2(n1309), .A3(n24033), .A4(n61438), .ZN(
        n37253) );
  INV_X1 U49082 ( .I(n50943), .ZN(n52068) );
  XOR2_X1 U49083 ( .A1(n37255), .A2(n37254), .Z(n37258) );
  XOR2_X1 U49084 ( .A1(n61034), .A2(n37256), .Z(n51980) );
  XOR2_X1 U49085 ( .A1(n37258), .A2(n51980), .Z(n50456) );
  XOR2_X1 U49086 ( .A1(n37259), .A2(n53685), .Z(n50944) );
  XOR2_X1 U49087 ( .A1(n50456), .A2(n50944), .Z(n37260) );
  XOR2_X1 U49088 ( .A1(n38909), .A2(n39437), .Z(n37262) );
  XOR2_X1 U49089 ( .A1(n37263), .A2(n37262), .Z(n37264) );
  XOR2_X1 U49090 ( .A1(n60039), .A2(n37264), .Z(n37265) );
  INV_X1 U49091 ( .I(n37277), .ZN(n37279) );
  INV_X1 U49092 ( .I(n37281), .ZN(n37282) );
  XOR2_X1 U49093 ( .A1(n38307), .A2(n55191), .Z(n39234) );
  XOR2_X1 U49095 ( .A1(n39631), .A2(n55340), .Z(n51149) );
  XOR2_X1 U49096 ( .A1(n52080), .A2(n60857), .Z(n37294) );
  XOR2_X1 U49097 ( .A1(n51149), .A2(n37294), .Z(n37295) );
  XOR2_X1 U49098 ( .A1(n37295), .A2(n51150), .Z(n37296) );
  XOR2_X1 U49099 ( .A1(n23249), .A2(n50969), .Z(n48748) );
  XOR2_X1 U49100 ( .A1(n37296), .A2(n48748), .Z(n37297) );
  XOR2_X1 U49101 ( .A1(n38916), .A2(n37297), .Z(n37298) );
  XOR2_X1 U49102 ( .A1(n37298), .A2(n24147), .Z(n37299) );
  INV_X1 U49104 ( .I(n52566), .ZN(n37306) );
  XOR2_X1 U49105 ( .A1(n46615), .A2(n37303), .Z(n37304) );
  XOR2_X1 U49106 ( .A1(n37305), .A2(n37304), .Z(n50719) );
  XOR2_X1 U49107 ( .A1(n37306), .A2(n50719), .Z(n37307) );
  XOR2_X1 U49108 ( .A1(n39004), .A2(n37308), .Z(n37309) );
  NAND2_X1 U49109 ( .A1(n37311), .A2(n37310), .ZN(n37941) );
  NAND2_X1 U49110 ( .A1(n37941), .A2(n37940), .ZN(n37312) );
  NAND3_X1 U49111 ( .A1(n4745), .A2(n13666), .A3(n37319), .ZN(n37321) );
  NAND2_X1 U49112 ( .A1(n37322), .A2(n37321), .ZN(n37944) );
  NAND3_X1 U49113 ( .A1(n37944), .A2(n19252), .A3(n37943), .ZN(n37323) );
  NAND2_X1 U49114 ( .A1(n37324), .A2(n37327), .ZN(n37325) );
  INV_X1 U49115 ( .I(n37339), .ZN(n37343) );
  INV_X1 U49116 ( .I(n37340), .ZN(n37342) );
  XOR2_X1 U49117 ( .A1(n39196), .A2(n53772), .Z(n50640) );
  XOR2_X1 U49118 ( .A1(n50640), .A2(n24058), .Z(n37347) );
  XOR2_X1 U49120 ( .A1(n39186), .A2(n52029), .Z(n37799) );
  XOR2_X1 U49121 ( .A1(n51479), .A2(n37348), .Z(n37349) );
  OAI21_X1 U49122 ( .A1(n2594), .A2(n37365), .B(n37364), .ZN(n37366) );
  AOI21_X1 U49123 ( .A1(n37369), .A2(n9783), .B(n37376), .ZN(n37370) );
  INV_X1 U49124 ( .I(n37378), .ZN(n37380) );
  XOR2_X1 U49125 ( .A1(n45088), .A2(n38236), .Z(n47936) );
  XOR2_X1 U49126 ( .A1(n51137), .A2(n47936), .Z(n37379) );
  XOR2_X1 U49127 ( .A1(n37380), .A2(n37379), .Z(n37381) );
  XOR2_X1 U49128 ( .A1(n37383), .A2(n37382), .Z(n37384) );
  XOR2_X1 U49129 ( .A1(n38878), .A2(n4691), .Z(n37386) );
  AOI21_X1 U49130 ( .A1(n37392), .A2(n37391), .B(n37390), .ZN(n37396) );
  NAND2_X1 U49131 ( .A1(n37398), .A2(n6540), .ZN(n37403) );
  INV_X1 U49132 ( .I(n37399), .ZN(n37401) );
  NAND2_X1 U49133 ( .A1(n37401), .A2(n37400), .ZN(n37402) );
  INV_X1 U49135 ( .I(n37406), .ZN(n37407) );
  INV_X1 U49136 ( .I(n37410), .ZN(n37413) );
  INV_X1 U49140 ( .I(n37419), .ZN(n37421) );
  OAI21_X1 U49141 ( .A1(n37421), .A2(n37420), .B(n37424), .ZN(n37433) );
  NAND3_X1 U49143 ( .A1(n22461), .A2(n37427), .A3(n37426), .ZN(n37429) );
  NAND2_X1 U49144 ( .A1(n37436), .A2(n37435), .ZN(n37439) );
  INV_X1 U49147 ( .I(n50712), .ZN(n45243) );
  XOR2_X1 U49148 ( .A1(n21967), .A2(n45243), .Z(n38593) );
  NOR3_X1 U49149 ( .A1(n37442), .A2(n12797), .A3(n22801), .ZN(n37443) );
  NOR2_X1 U49150 ( .A1(n37444), .A2(n37454), .ZN(n37449) );
  INV_X1 U49151 ( .I(n37445), .ZN(n37448) );
  NAND2_X1 U49154 ( .A1(n24033), .A2(n9869), .ZN(n37456) );
  XOR2_X1 U49156 ( .A1(n37458), .A2(n54896), .Z(n52526) );
  XOR2_X1 U49157 ( .A1(n52526), .A2(n50709), .Z(n37459) );
  XOR2_X1 U49158 ( .A1(n22480), .A2(n37459), .Z(n37460) );
  XOR2_X1 U49159 ( .A1(n38276), .A2(n63000), .Z(n37472) );
  INV_X1 U49160 ( .I(n37464), .ZN(n37467) );
  XOR2_X1 U49161 ( .A1(n37465), .A2(n38387), .Z(n37466) );
  XOR2_X1 U49162 ( .A1(n37467), .A2(n37466), .Z(n50169) );
  XOR2_X1 U49163 ( .A1(n37468), .A2(n54126), .Z(n51920) );
  XOR2_X1 U49164 ( .A1(n50169), .A2(n51920), .Z(n37469) );
  XOR2_X1 U49165 ( .A1(n23199), .A2(n37469), .Z(n37470) );
  XOR2_X1 U49166 ( .A1(n59882), .A2(n37470), .Z(n37471) );
  NAND2_X1 U49167 ( .A1(n37473), .A2(n63838), .ZN(n37474) );
  NAND2_X1 U49168 ( .A1(n37475), .A2(n37474), .ZN(n38549) );
  AOI21_X1 U49169 ( .A1(n38549), .A2(n38550), .B(n37478), .ZN(n37479) );
  NAND2_X1 U49170 ( .A1(n37479), .A2(n38548), .ZN(n37673) );
  XOR2_X1 U49171 ( .A1(n52135), .A2(n54734), .Z(n51045) );
  XOR2_X1 U49172 ( .A1(n15712), .A2(n53090), .Z(n37480) );
  XOR2_X1 U49173 ( .A1(n51045), .A2(n37480), .Z(n37482) );
  XOR2_X1 U49174 ( .A1(n37481), .A2(n53272), .Z(n52553) );
  XOR2_X1 U49175 ( .A1(n37482), .A2(n52553), .Z(n37484) );
  INV_X1 U49176 ( .I(n50733), .ZN(n37483) );
  XOR2_X1 U49177 ( .A1(n37484), .A2(n37483), .Z(n37485) );
  XOR2_X1 U49178 ( .A1(n37486), .A2(n27640), .Z(n52138) );
  XOR2_X1 U49179 ( .A1(n23931), .A2(n52138), .Z(n38428) );
  XOR2_X1 U49180 ( .A1(n37487), .A2(n38428), .Z(n37488) );
  NOR2_X1 U49181 ( .A1(n37491), .A2(n37490), .ZN(n37493) );
  INV_X1 U49182 ( .I(n51218), .ZN(n46207) );
  XOR2_X1 U49183 ( .A1(n53833), .A2(n55150), .Z(n51654) );
  XOR2_X1 U49184 ( .A1(n46207), .A2(n51654), .Z(n38517) );
  XOR2_X1 U49185 ( .A1(n38472), .A2(n37497), .Z(n37498) );
  XOR2_X1 U49186 ( .A1(n38517), .A2(n37498), .Z(n51142) );
  XOR2_X1 U49187 ( .A1(n37692), .A2(n37500), .Z(n51545) );
  XOR2_X1 U49188 ( .A1(n51665), .A2(n52197), .Z(n37503) );
  XNOR2_X1 U49189 ( .A1(n55191), .A2(n60797), .ZN(n37501) );
  XOR2_X1 U49190 ( .A1(n37501), .A2(n37651), .Z(n37502) );
  XOR2_X1 U49191 ( .A1(n37503), .A2(n37502), .Z(n37504) );
  XOR2_X1 U49192 ( .A1(n51545), .A2(n37504), .Z(n37505) );
  XOR2_X1 U49193 ( .A1(n38912), .A2(n37505), .Z(n37506) );
  XOR2_X1 U49194 ( .A1(n38373), .A2(n38946), .Z(n37508) );
  AOI22_X1 U49195 ( .A1(n37510), .A2(n37529), .B1(n7649), .B2(n1512), .ZN(
        n37528) );
  XOR2_X1 U49196 ( .A1(n37512), .A2(n38588), .Z(n51934) );
  XOR2_X1 U49197 ( .A1(n37513), .A2(n54716), .Z(n37514) );
  XOR2_X1 U49198 ( .A1(n44264), .A2(n37514), .Z(n50161) );
  XOR2_X1 U49199 ( .A1(n51934), .A2(n50161), .Z(n37515) );
  XOR2_X1 U49200 ( .A1(n58926), .A2(n37888), .Z(n37516) );
  XOR2_X1 U49201 ( .A1(n38988), .A2(n23695), .Z(n37517) );
  INV_X1 U49202 ( .I(n51575), .ZN(n37522) );
  XOR2_X1 U49203 ( .A1(n37520), .A2(n37519), .Z(n51524) );
  XOR2_X1 U49204 ( .A1(n50486), .A2(n54208), .Z(n45338) );
  XOR2_X1 U49205 ( .A1(n51524), .A2(n45338), .Z(n37521) );
  XOR2_X1 U49206 ( .A1(n37522), .A2(n37521), .Z(n37523) );
  XOR2_X1 U49207 ( .A1(n39284), .A2(n37523), .Z(n37524) );
  NOR2_X1 U49208 ( .A1(n1512), .A2(n23355), .ZN(n37530) );
  INV_X1 U49209 ( .I(n37535), .ZN(n37537) );
  INV_X1 U49210 ( .I(n41795), .ZN(n37542) );
  NAND2_X1 U49211 ( .A1(n429), .A2(n5126), .ZN(n37541) );
  OAI21_X1 U49212 ( .A1(n41796), .A2(n37541), .B(n42031), .ZN(n43585) );
  AOI21_X1 U49213 ( .A1(n37542), .A2(n41794), .B(n43585), .ZN(n37543) );
  INV_X1 U49214 ( .I(n45288), .ZN(n37546) );
  XOR2_X1 U49215 ( .A1(n45121), .A2(n65079), .Z(n37544) );
  XOR2_X1 U49216 ( .A1(n51841), .A2(n37544), .Z(n37545) );
  XOR2_X1 U49217 ( .A1(n37546), .A2(n37545), .Z(n37547) );
  INV_X1 U49220 ( .I(n37721), .ZN(n37550) );
  XOR2_X1 U49221 ( .A1(n23330), .A2(n55765), .Z(n38957) );
  XOR2_X1 U49222 ( .A1(n51765), .A2(n620), .Z(n37557) );
  XOR2_X1 U49223 ( .A1(n51766), .A2(n37557), .Z(n37558) );
  XOR2_X1 U49224 ( .A1(n44331), .A2(n37558), .Z(n37559) );
  XOR2_X1 U49225 ( .A1(n39259), .A2(n37559), .Z(n37560) );
  XOR2_X1 U49226 ( .A1(n7619), .A2(n37560), .Z(n37561) );
  INV_X1 U49227 ( .I(n38117), .ZN(n37564) );
  XOR2_X1 U49228 ( .A1(n38614), .A2(n37565), .Z(n37566) );
  XOR2_X1 U49229 ( .A1(n38153), .A2(n37566), .Z(n52003) );
  XOR2_X1 U49230 ( .A1(n50777), .A2(n53076), .Z(n49403) );
  XOR2_X1 U49231 ( .A1(n39492), .A2(n37567), .Z(n37568) );
  XOR2_X1 U49232 ( .A1(n22487), .A2(n55610), .Z(n37770) );
  XOR2_X1 U49233 ( .A1(n37698), .A2(n37770), .Z(n37569) );
  XOR2_X1 U49234 ( .A1(n51193), .A2(n24098), .Z(n51319) );
  XOR2_X1 U49235 ( .A1(n37570), .A2(n51319), .Z(n37571) );
  XOR2_X1 U49236 ( .A1(n51310), .A2(n37571), .Z(n37572) );
  XOR2_X1 U49237 ( .A1(n37572), .A2(n51718), .Z(n37573) );
  XOR2_X1 U49238 ( .A1(n60597), .A2(n37573), .Z(n37574) );
  XOR2_X1 U49239 ( .A1(n37745), .A2(n37574), .Z(n37575) );
  XOR2_X1 U49240 ( .A1(n23790), .A2(n50741), .Z(n37579) );
  XOR2_X1 U49241 ( .A1(n44914), .A2(n22458), .Z(n49589) );
  XOR2_X1 U49242 ( .A1(n37881), .A2(n37585), .Z(n37586) );
  XOR2_X1 U49243 ( .A1(n37586), .A2(n55840), .Z(n52010) );
  XOR2_X1 U49244 ( .A1(n49589), .A2(n52010), .Z(n37587) );
  XOR2_X1 U49245 ( .A1(n39625), .A2(n37587), .Z(n37588) );
  NAND2_X1 U49250 ( .A1(n41248), .A2(n22713), .ZN(n37594) );
  XOR2_X1 U49251 ( .A1(n43065), .A2(n44014), .Z(n50710) );
  XOR2_X1 U49252 ( .A1(n52527), .A2(n50710), .Z(n37602) );
  AOI21_X1 U49253 ( .A1(n37600), .A2(n37601), .B(n37602), .ZN(n37607) );
  INV_X1 U49254 ( .I(n37600), .ZN(n37605) );
  INV_X1 U49255 ( .I(n37601), .ZN(n37604) );
  INV_X1 U49256 ( .I(n37602), .ZN(n37603) );
  NOR3_X1 U49257 ( .A1(n37605), .A2(n37604), .A3(n37603), .ZN(n37606) );
  NOR2_X1 U49258 ( .A1(n37607), .A2(n37606), .ZN(n37608) );
  XOR2_X1 U49259 ( .A1(n23493), .A2(n38411), .Z(n37823) );
  NAND3_X1 U49260 ( .A1(n37613), .A2(n37617), .A3(n47768), .ZN(n37614) );
  OAI22_X1 U49261 ( .A1(n37615), .A2(n37614), .B1(n47768), .B2(n37613), .ZN(
        n37623) );
  INV_X1 U49262 ( .I(n37616), .ZN(n37619) );
  INV_X1 U49263 ( .I(n37617), .ZN(n37618) );
  NOR2_X1 U49264 ( .A1(n37619), .A2(n37618), .ZN(n37621) );
  AOI21_X1 U49265 ( .A1(n37621), .A2(n37620), .B(n47768), .ZN(n37622) );
  XOR2_X1 U49267 ( .A1(n38741), .A2(n38120), .Z(n37627) );
  XOR2_X1 U49268 ( .A1(n56124), .A2(n55242), .Z(n51131) );
  XOR2_X1 U49269 ( .A1(n4762), .A2(n51131), .Z(n37626) );
  XOR2_X1 U49270 ( .A1(n37626), .A2(n37627), .Z(n39681) );
  XOR2_X1 U49272 ( .A1(n24057), .A2(n56322), .Z(n37629) );
  XOR2_X1 U49273 ( .A1(n37630), .A2(n37629), .Z(n52613) );
  XOR2_X1 U49274 ( .A1(n37631), .A2(n52613), .Z(n37632) );
  INV_X1 U49275 ( .I(n37635), .ZN(n38774) );
  INV_X1 U49276 ( .I(n37636), .ZN(n37640) );
  XOR2_X1 U49277 ( .A1(n37638), .A2(n37637), .Z(n37639) );
  XOR2_X1 U49278 ( .A1(n37640), .A2(n37639), .Z(n37641) );
  XOR2_X1 U49279 ( .A1(n38774), .A2(n37641), .Z(n50945) );
  XOR2_X1 U49280 ( .A1(n65079), .A2(n56508), .Z(n37642) );
  XOR2_X1 U49281 ( .A1(n52178), .A2(n37642), .Z(n37643) );
  XOR2_X1 U49282 ( .A1(n37643), .A2(n50453), .Z(n37644) );
  XOR2_X1 U49283 ( .A1(n50945), .A2(n37644), .Z(n37645) );
  INV_X1 U49284 ( .I(n24276), .ZN(n37646) );
  XOR2_X1 U49285 ( .A1(n37651), .A2(n50817), .Z(n37652) );
  XOR2_X1 U49286 ( .A1(n37652), .A2(n50798), .Z(n37653) );
  XOR2_X1 U49287 ( .A1(n45067), .A2(n37653), .Z(n51152) );
  XNOR2_X1 U49288 ( .A1(n52317), .A2(n51569), .ZN(n37654) );
  XOR2_X1 U49289 ( .A1(n37654), .A2(n46336), .Z(n37655) );
  XOR2_X1 U49290 ( .A1(n42579), .A2(n37655), .Z(n48747) );
  XOR2_X1 U49291 ( .A1(n51152), .A2(n48747), .Z(n37656) );
  INV_X1 U49293 ( .I(n50720), .ZN(n37660) );
  XOR2_X1 U49294 ( .A1(n50641), .A2(n52565), .Z(n37659) );
  XOR2_X1 U49295 ( .A1(n37660), .A2(n37659), .Z(n37661) );
  XOR2_X1 U49296 ( .A1(n39628), .A2(n16449), .Z(n37662) );
  NAND2_X1 U49298 ( .A1(n18338), .A2(n40826), .ZN(n37664) );
  AOI22_X1 U49299 ( .A1(n39516), .A2(n37664), .B1(n39508), .B2(n23890), .ZN(
        n37665) );
  INV_X1 U49300 ( .I(n50903), .ZN(n37668) );
  XOR2_X1 U49301 ( .A1(n54676), .A2(n53772), .Z(n37666) );
  XOR2_X1 U49302 ( .A1(n46443), .A2(n37666), .Z(n50227) );
  XOR2_X1 U49303 ( .A1(n50227), .A2(n15710), .Z(n37667) );
  XOR2_X1 U49304 ( .A1(n37668), .A2(n37667), .Z(n37669) );
  INV_X1 U49306 ( .I(n52141), .ZN(n45037) );
  XOR2_X1 U49307 ( .A1(n50628), .A2(n37674), .Z(n37675) );
  XOR2_X1 U49308 ( .A1(n45037), .A2(n37675), .Z(n37676) );
  INV_X1 U49309 ( .I(n52135), .ZN(n37679) );
  XOR2_X1 U49310 ( .A1(n11751), .A2(n37679), .Z(n37680) );
  XOR2_X1 U49311 ( .A1(n52178), .A2(n57989), .Z(n37683) );
  XOR2_X1 U49312 ( .A1(n49957), .A2(n37683), .Z(n51658) );
  XOR2_X1 U49313 ( .A1(n37838), .A2(n53989), .Z(n51070) );
  XOR2_X1 U49314 ( .A1(n51658), .A2(n51070), .Z(n37684) );
  XOR2_X1 U49315 ( .A1(n9871), .A2(n53833), .Z(n52575) );
  XOR2_X1 U49316 ( .A1(n25161), .A2(n20087), .Z(n37687) );
  XOR2_X1 U49317 ( .A1(n10017), .A2(n23330), .Z(n37689) );
  XOR2_X1 U49318 ( .A1(n24257), .A2(n23306), .Z(n38913) );
  XNOR2_X1 U49319 ( .A1(n55765), .A2(n55052), .ZN(n37690) );
  XOR2_X1 U49320 ( .A1(n64355), .A2(n37690), .Z(n51419) );
  XOR2_X1 U49321 ( .A1(n37692), .A2(n51419), .Z(n37693) );
  XOR2_X1 U49322 ( .A1(n10304), .A2(n37693), .Z(n37694) );
  XOR2_X1 U49323 ( .A1(n37695), .A2(n9398), .Z(n37696) );
  XOR2_X1 U49324 ( .A1(n57452), .A2(n50878), .Z(n37701) );
  XOR2_X1 U49325 ( .A1(n37703), .A2(n53076), .Z(n50320) );
  XOR2_X1 U49326 ( .A1(n55196), .A2(n53805), .Z(n39567) );
  XOR2_X1 U49327 ( .A1(n37704), .A2(n39567), .Z(n37705) );
  XOR2_X1 U49328 ( .A1(n44264), .A2(n37705), .Z(n50917) );
  XOR2_X1 U49329 ( .A1(n50320), .A2(n50917), .Z(n37706) );
  XOR2_X1 U49332 ( .A1(n59688), .A2(n39460), .Z(n37717) );
  XOR2_X1 U49333 ( .A1(n37710), .A2(n55106), .Z(n37711) );
  XOR2_X1 U49334 ( .A1(n37712), .A2(n37711), .Z(n51354) );
  XOR2_X1 U49335 ( .A1(n37713), .A2(n53530), .Z(n52633) );
  XOR2_X1 U49336 ( .A1(n52633), .A2(n54208), .Z(n37714) );
  XOR2_X1 U49337 ( .A1(n51354), .A2(n37714), .Z(n37715) );
  XOR2_X1 U49338 ( .A1(n39284), .A2(n37715), .Z(n37716) );
  XOR2_X1 U49339 ( .A1(n37717), .A2(n37716), .Z(n37718) );
  INV_X1 U49340 ( .I(n39439), .ZN(n37722) );
  XOR2_X1 U49341 ( .A1(n45123), .A2(n55379), .Z(n39350) );
  XOR2_X1 U49342 ( .A1(n44876), .A2(n39350), .Z(n50887) );
  XOR2_X1 U49343 ( .A1(n56714), .A2(n53359), .Z(n49875) );
  XOR2_X1 U49344 ( .A1(n50887), .A2(n49875), .Z(n37723) );
  XOR2_X1 U49345 ( .A1(n37729), .A2(n56309), .Z(n39335) );
  XOR2_X1 U49346 ( .A1(n39335), .A2(n37730), .Z(n37731) );
  XOR2_X1 U49347 ( .A1(n37731), .A2(n39443), .Z(n51091) );
  XOR2_X1 U49348 ( .A1(n51667), .A2(n52080), .Z(n37732) );
  XOR2_X1 U49349 ( .A1(n51091), .A2(n37732), .Z(n37733) );
  XOR2_X1 U49350 ( .A1(n10017), .A2(n37733), .Z(n37734) );
  INV_X1 U49351 ( .I(n37736), .ZN(n37738) );
  XOR2_X1 U49352 ( .A1(n37738), .A2(n37737), .Z(n51649) );
  XOR2_X1 U49353 ( .A1(n37739), .A2(n46488), .Z(n37788) );
  XOR2_X1 U49354 ( .A1(n37788), .A2(n53705), .Z(n51060) );
  XOR2_X1 U49355 ( .A1(n51649), .A2(n51060), .Z(n37740) );
  XOR2_X1 U49356 ( .A1(n18057), .A2(n37740), .Z(n37741) );
  XOR2_X1 U49357 ( .A1(n37742), .A2(n37741), .Z(n37743) );
  XOR2_X1 U49358 ( .A1(n59688), .A2(n22485), .Z(n37899) );
  XOR2_X1 U49359 ( .A1(n38500), .A2(n37899), .Z(n37744) );
  XOR2_X1 U49360 ( .A1(n12669), .A2(n23332), .Z(n38173) );
  XOR2_X1 U49361 ( .A1(n38173), .A2(n37901), .Z(n37746) );
  INV_X1 U49362 ( .I(n37748), .ZN(n37753) );
  XOR2_X1 U49363 ( .A1(n52327), .A2(n50502), .Z(n37751) );
  XOR2_X1 U49364 ( .A1(n37749), .A2(n22323), .Z(n37750) );
  XOR2_X1 U49365 ( .A1(n37751), .A2(n37750), .Z(n37752) );
  XOR2_X1 U49366 ( .A1(n37753), .A2(n37752), .Z(n37754) );
  XOR2_X1 U49367 ( .A1(n37758), .A2(n37757), .Z(n50636) );
  XOR2_X1 U49368 ( .A1(n15710), .A2(n54870), .Z(n37759) );
  XOR2_X1 U49369 ( .A1(n50636), .A2(n37759), .Z(n37760) );
  XOR2_X1 U49370 ( .A1(n39704), .A2(n38995), .Z(n52150) );
  NAND2_X1 U49372 ( .A1(n42264), .A2(n11677), .ZN(n37762) );
  NAND3_X1 U49373 ( .A1(n42265), .A2(n41098), .A3(n37762), .ZN(n37772) );
  XOR2_X1 U49374 ( .A1(n37763), .A2(n38966), .Z(n39225) );
  XOR2_X1 U49375 ( .A1(n9826), .A2(n46554), .Z(n37766) );
  XOR2_X1 U49376 ( .A1(n37764), .A2(n55196), .Z(n37765) );
  XOR2_X1 U49377 ( .A1(n37766), .A2(n37765), .Z(n52162) );
  XOR2_X1 U49378 ( .A1(n37767), .A2(n54536), .Z(n37768) );
  XOR2_X1 U49379 ( .A1(n38588), .A2(n37768), .Z(n50607) );
  XOR2_X1 U49380 ( .A1(n52162), .A2(n50607), .Z(n37769) );
  INV_X1 U49382 ( .I(n37778), .ZN(n37781) );
  XOR2_X1 U49383 ( .A1(n49957), .A2(n53764), .Z(n37779) );
  XOR2_X1 U49384 ( .A1(n12356), .A2(n37779), .Z(n37780) );
  XOR2_X1 U49385 ( .A1(n37781), .A2(n37780), .Z(n37782) );
  XOR2_X1 U49387 ( .A1(n61105), .A2(n22485), .Z(n37785) );
  INV_X1 U49388 ( .I(n23789), .ZN(n37787) );
  XOR2_X1 U49389 ( .A1(n37788), .A2(n37787), .Z(n51192) );
  XOR2_X1 U49390 ( .A1(n50698), .A2(n51815), .Z(n37789) );
  XOR2_X1 U49391 ( .A1(n51192), .A2(n37789), .Z(n37790) );
  INV_X1 U49392 ( .I(n52449), .ZN(n37794) );
  XOR2_X1 U49393 ( .A1(n37794), .A2(n44108), .Z(n37796) );
  XOR2_X1 U49394 ( .A1(n44841), .A2(n37795), .Z(n52329) );
  XOR2_X1 U49395 ( .A1(n37796), .A2(n52329), .Z(n37797) );
  XOR2_X1 U49396 ( .A1(n23931), .A2(n37797), .Z(n37798) );
  XOR2_X1 U49397 ( .A1(n37803), .A2(n39200), .Z(n52111) );
  XOR2_X1 U49398 ( .A1(n50763), .A2(n15710), .Z(n37804) );
  XOR2_X1 U49399 ( .A1(n52111), .A2(n37804), .Z(n37805) );
  XOR2_X1 U49400 ( .A1(n24300), .A2(n37805), .Z(n37806) );
  INV_X1 U49401 ( .I(n37808), .ZN(n46595) );
  XOR2_X1 U49402 ( .A1(n46595), .A2(n37809), .Z(n51826) );
  XOR2_X1 U49403 ( .A1(n52513), .A2(n54708), .Z(n51204) );
  XOR2_X1 U49404 ( .A1(n51826), .A2(n51204), .Z(n37810) );
  XOR2_X1 U49405 ( .A1(n38784), .A2(n37810), .Z(n37811) );
  INV_X1 U49406 ( .I(n52197), .ZN(n51543) );
  XOR2_X1 U49407 ( .A1(n15704), .A2(n22988), .Z(n37813) );
  XOR2_X1 U49408 ( .A1(n39450), .A2(n37813), .Z(n37814) );
  XOR2_X1 U49410 ( .A1(n37818), .A2(n9896), .Z(n37819) );
  XNOR2_X1 U49411 ( .A1(n55777), .A2(n54716), .ZN(n37822) );
  XOR2_X1 U49412 ( .A1(n23767), .A2(n37822), .Z(n52050) );
  NAND2_X1 U49413 ( .A1(n59583), .A2(n41051), .ZN(n37827) );
  NAND2_X1 U49415 ( .A1(n41873), .A2(n41064), .ZN(n37829) );
  NAND2_X1 U49416 ( .A1(n39795), .A2(n41876), .ZN(n37830) );
  NOR2_X1 U49417 ( .A1(n37833), .A2(n37832), .ZN(n37923) );
  XOR2_X1 U49418 ( .A1(n57989), .A2(n55150), .Z(n51840) );
  XOR2_X1 U49419 ( .A1(n1881), .A2(n51840), .Z(n37835) );
  XOR2_X1 U49420 ( .A1(n37836), .A2(n37835), .Z(n48968) );
  XOR2_X1 U49421 ( .A1(n37838), .A2(n37837), .Z(n51141) );
  XOR2_X1 U49422 ( .A1(n51141), .A2(n56508), .Z(n37839) );
  XOR2_X1 U49423 ( .A1(n48968), .A2(n37839), .Z(n37840) );
  XOR2_X1 U49425 ( .A1(n51765), .A2(n53787), .Z(n37843) );
  XOR2_X1 U49426 ( .A1(n37843), .A2(n51542), .Z(n37845) );
  XOR2_X1 U49427 ( .A1(n37845), .A2(n37844), .Z(n37846) );
  XOR2_X1 U49428 ( .A1(n38530), .A2(n37846), .Z(n37848) );
  XOR2_X1 U49429 ( .A1(n51766), .A2(n37847), .Z(n51607) );
  XOR2_X1 U49430 ( .A1(n19261), .A2(n51607), .Z(n38062) );
  NOR2_X1 U49431 ( .A1(n37851), .A2(n37850), .ZN(n37854) );
  INV_X1 U49432 ( .I(n37856), .ZN(n37853) );
  XOR2_X1 U49433 ( .A1(n37852), .A2(n50817), .Z(n37855) );
  NAND4_X1 U49434 ( .A1(n37854), .A2(n37853), .A3(n37858), .A4(n37855), .ZN(
        n37862) );
  INV_X1 U49435 ( .I(n37854), .ZN(n37857) );
  INV_X1 U49436 ( .I(n37855), .ZN(n51551) );
  OAI21_X1 U49437 ( .A1(n37857), .A2(n37856), .B(n51551), .ZN(n37861) );
  INV_X1 U49438 ( .I(n37858), .ZN(n37859) );
  NAND2_X1 U49439 ( .A1(n37859), .A2(n51551), .ZN(n37860) );
  NAND3_X1 U49440 ( .A1(n37862), .A2(n37861), .A3(n37860), .ZN(n38920) );
  XOR2_X1 U49441 ( .A1(n37863), .A2(n38920), .Z(n37864) );
  XOR2_X1 U49442 ( .A1(n37869), .A2(n37868), .Z(n45818) );
  XOR2_X1 U49443 ( .A1(n44841), .A2(n50505), .Z(n37870) );
  XOR2_X1 U49444 ( .A1(n45818), .A2(n37870), .Z(n52555) );
  XOR2_X1 U49445 ( .A1(n39613), .A2(n24051), .Z(n46152) );
  XOR2_X1 U49446 ( .A1(n46152), .A2(n55139), .Z(n37871) );
  XOR2_X1 U49447 ( .A1(n52555), .A2(n37871), .Z(n37872) );
  XOR2_X1 U49448 ( .A1(n38575), .A2(n59882), .Z(n38447) );
  XOR2_X1 U49449 ( .A1(n39528), .A2(n38447), .Z(n37877) );
  XOR2_X1 U49450 ( .A1(n37876), .A2(n37877), .Z(n37887) );
  INV_X1 U49451 ( .I(n38826), .ZN(n37879) );
  XOR2_X1 U49452 ( .A1(n37879), .A2(n37878), .Z(n37880) );
  XOR2_X1 U49453 ( .A1(n37881), .A2(n37880), .Z(n37882) );
  XOR2_X1 U49454 ( .A1(n37883), .A2(n37882), .Z(n51921) );
  XOR2_X1 U49455 ( .A1(n38556), .A2(n24014), .Z(n50168) );
  XOR2_X1 U49456 ( .A1(n51921), .A2(n50168), .Z(n37884) );
  XOR2_X1 U49457 ( .A1(n39625), .A2(n37884), .Z(n37885) );
  XOR2_X1 U49458 ( .A1(n59680), .A2(n29969), .Z(n38223) );
  XOR2_X1 U49459 ( .A1(n38223), .A2(n50873), .Z(n50162) );
  XOR2_X1 U49460 ( .A1(n37890), .A2(n37889), .Z(n51935) );
  XOR2_X1 U49461 ( .A1(n50162), .A2(n51935), .Z(n37891) );
  XOR2_X1 U49462 ( .A1(n38411), .A2(n37891), .Z(n37892) );
  XOR2_X1 U49463 ( .A1(n37894), .A2(n9896), .Z(n39779) );
  XOR2_X1 U49464 ( .A1(n38235), .A2(n37896), .Z(n51523) );
  XOR2_X1 U49465 ( .A1(n22252), .A2(n37897), .Z(n51573) );
  XOR2_X1 U49466 ( .A1(n51523), .A2(n51573), .Z(n37898) );
  XOR2_X1 U49467 ( .A1(n60597), .A2(n51319), .Z(n38456) );
  XOR2_X1 U49468 ( .A1(n38456), .A2(n37899), .Z(n37900) );
  INV_X1 U49469 ( .I(n22855), .ZN(n38121) );
  XOR2_X1 U49470 ( .A1(n7418), .A2(n38121), .Z(n38245) );
  NOR3_X1 U49473 ( .A1(n41924), .A2(n64768), .A3(n61785), .ZN(n37904) );
  INV_X1 U49475 ( .I(n40786), .ZN(n37906) );
  NOR2_X1 U49476 ( .A1(n37907), .A2(n37906), .ZN(n37910) );
  INV_X1 U49477 ( .I(n40559), .ZN(n37908) );
  NAND2_X1 U49478 ( .A1(n37908), .A2(n41255), .ZN(n37909) );
  INV_X1 U49479 ( .I(n43703), .ZN(n37914) );
  NAND2_X1 U49486 ( .A1(n40250), .A2(n40464), .ZN(n37928) );
  MUX2_X1 U49489 ( .I0(n37942), .I1(n37941), .S(n37940), .Z(n37947) );
  NAND2_X1 U49490 ( .A1(n37944), .A2(n37943), .ZN(n37946) );
  MUX2_X1 U49491 ( .I0(n37947), .I1(n37946), .S(n19252), .Z(n37949) );
  XOR2_X1 U49492 ( .A1(n60207), .A2(n52565), .Z(n37951) );
  XOR2_X1 U49493 ( .A1(n37951), .A2(n37950), .Z(n51381) );
  XOR2_X1 U49494 ( .A1(n51381), .A2(n52226), .Z(n37953) );
  XOR2_X1 U49495 ( .A1(n53641), .A2(n57096), .Z(n39195) );
  XOR2_X1 U49496 ( .A1(n37952), .A2(n39195), .Z(n52605) );
  XOR2_X1 U49497 ( .A1(n37953), .A2(n52605), .Z(n37954) );
  INV_X1 U49498 ( .I(n37956), .ZN(n39523) );
  INV_X1 U49499 ( .I(n37958), .ZN(n37959) );
  NAND2_X1 U49500 ( .A1(n37960), .A2(n37959), .ZN(n37961) );
  INV_X1 U49501 ( .I(n37962), .ZN(n37963) );
  XOR2_X1 U49503 ( .A1(n39206), .A2(n16594), .Z(n39627) );
  XOR2_X1 U49504 ( .A1(n2334), .A2(n9931), .Z(n37969) );
  XOR2_X1 U49505 ( .A1(n37973), .A2(n54734), .Z(n46351) );
  XOR2_X1 U49506 ( .A1(n52135), .A2(n56180), .Z(n51004) );
  XOR2_X1 U49507 ( .A1(n44311), .A2(n51004), .Z(n37974) );
  XOR2_X1 U49508 ( .A1(n46351), .A2(n37974), .Z(n37975) );
  XOR2_X1 U49510 ( .A1(n37981), .A2(n15707), .Z(n44430) );
  INV_X1 U49511 ( .I(n7264), .ZN(n37982) );
  XOR2_X1 U49512 ( .A1(n44430), .A2(n37982), .Z(n50935) );
  XOR2_X1 U49513 ( .A1(n37983), .A2(n54708), .Z(n50388) );
  XOR2_X1 U49514 ( .A1(n50388), .A2(n57113), .Z(n37984) );
  XOR2_X1 U49515 ( .A1(n50935), .A2(n37984), .Z(n37985) );
  XOR2_X1 U49516 ( .A1(n9397), .A2(n37985), .Z(n37986) );
  XOR2_X1 U49518 ( .A1(n1755), .A2(n39267), .Z(n37990) );
  XOR2_X1 U49519 ( .A1(n53685), .A2(n57142), .Z(n37991) );
  XOR2_X1 U49520 ( .A1(n43858), .A2(n37991), .Z(n37992) );
  XOR2_X1 U49521 ( .A1(n37993), .A2(n37992), .Z(n52182) );
  XOR2_X1 U49522 ( .A1(n52178), .A2(n53102), .Z(n45846) );
  XOR2_X1 U49523 ( .A1(n45846), .A2(n51261), .Z(n37994) );
  XOR2_X1 U49524 ( .A1(n37994), .A2(n247), .Z(n37995) );
  XOR2_X1 U49525 ( .A1(n4563), .A2(n39582), .Z(n37997) );
  INV_X1 U49526 ( .I(n58235), .ZN(n37998) );
  XOR2_X1 U49527 ( .A1(n37999), .A2(n39570), .Z(n52625) );
  XOR2_X1 U49528 ( .A1(n38000), .A2(n54153), .Z(n51371) );
  XOR2_X1 U49529 ( .A1(n51371), .A2(n51379), .Z(n38001) );
  XOR2_X1 U49530 ( .A1(n52625), .A2(n38001), .Z(n38002) );
  INV_X1 U49531 ( .I(n39733), .ZN(n38005) );
  XOR2_X1 U49532 ( .A1(n38006), .A2(n38005), .Z(n39680) );
  INV_X1 U49533 ( .I(n44925), .ZN(n38008) );
  XOR2_X1 U49534 ( .A1(n38008), .A2(n38007), .Z(n38011) );
  XOR2_X1 U49535 ( .A1(n38011), .A2(n38010), .Z(n50328) );
  XOR2_X1 U49536 ( .A1(n50924), .A2(n52232), .Z(n38012) );
  XOR2_X1 U49537 ( .A1(n50328), .A2(n38012), .Z(n38013) );
  XOR2_X1 U49538 ( .A1(n38989), .A2(n38013), .Z(n38014) );
  XOR2_X1 U49539 ( .A1(n38014), .A2(n204), .Z(n38015) );
  INV_X1 U49540 ( .I(n40051), .ZN(n40055) );
  NAND2_X1 U49542 ( .A1(n23711), .A2(n4581), .ZN(n38018) );
  NOR2_X1 U49543 ( .A1(n40056), .A2(n40267), .ZN(n38017) );
  NOR2_X1 U49544 ( .A1(n12285), .A2(n19990), .ZN(n38022) );
  INV_X1 U49547 ( .I(n40236), .ZN(n38029) );
  INV_X1 U49548 ( .I(n40232), .ZN(n38028) );
  OAI22_X1 U49549 ( .A1(n38029), .A2(n38028), .B1(n39414), .B2(n39419), .ZN(
        n38034) );
  OAI21_X1 U49550 ( .A1(n24188), .A2(n40070), .B(n36648), .ZN(n38030) );
  OAI21_X1 U49551 ( .A1(n39418), .A2(n2234), .B(n38030), .ZN(n38033) );
  NAND2_X1 U49552 ( .A1(n24188), .A2(n40070), .ZN(n38031) );
  NOR2_X1 U49555 ( .A1(n40996), .A2(n23752), .ZN(n38037) );
  NAND3_X1 U49556 ( .A1(n40146), .A2(n40143), .A3(n23833), .ZN(n38043) );
  NAND3_X1 U49557 ( .A1(n40147), .A2(n40215), .A3(n1509), .ZN(n38042) );
  NAND3_X1 U49559 ( .A1(n38046), .A2(n15558), .A3(n58941), .ZN(n38047) );
  NAND3_X1 U49560 ( .A1(n18612), .A2(n40944), .A3(n40200), .ZN(n38050) );
  AOI21_X1 U49561 ( .A1(n40204), .A2(n40202), .B(n38050), .ZN(n38051) );
  OAI21_X1 U49563 ( .A1(n38055), .A2(n42392), .B(n64492), .ZN(n38057) );
  NAND2_X1 U49564 ( .A1(n38057), .A2(n41708), .ZN(n38060) );
  MUX2_X1 U49565 ( .I0(n38058), .I1(n41694), .S(n41692), .Z(n38059) );
  INV_X1 U49566 ( .I(n38064), .ZN(n38067) );
  XOR2_X1 U49567 ( .A1(n38065), .A2(n42426), .Z(n38066) );
  XOR2_X1 U49568 ( .A1(n38067), .A2(n38066), .Z(n50564) );
  XOR2_X1 U49569 ( .A1(n38645), .A2(n50564), .Z(n38068) );
  INV_X1 U49570 ( .I(n38073), .ZN(n38075) );
  XOR2_X1 U49571 ( .A1(n38074), .A2(n38075), .Z(n50174) );
  XOR2_X1 U49572 ( .A1(n52734), .A2(n56065), .Z(n38076) );
  XOR2_X1 U49573 ( .A1(n51926), .A2(n38076), .Z(n38077) );
  XOR2_X1 U49574 ( .A1(n50174), .A2(n38077), .Z(n38078) );
  XOR2_X1 U49575 ( .A1(n23898), .A2(n38078), .Z(n38079) );
  INV_X1 U49576 ( .I(n49967), .ZN(n38085) );
  XOR2_X1 U49577 ( .A1(n38085), .A2(n23926), .Z(n46170) );
  XOR2_X1 U49578 ( .A1(n50998), .A2(n56905), .Z(n38086) );
  XOR2_X1 U49579 ( .A1(n39625), .A2(n16594), .Z(n38087) );
  XOR2_X1 U49580 ( .A1(n38087), .A2(n38386), .Z(n38089) );
  XOR2_X1 U49582 ( .A1(n39258), .A2(n38089), .Z(n38090) );
  INV_X1 U49583 ( .I(n51165), .ZN(n38091) );
  BUF_X2 U49584 ( .I(n38093), .Z(n42518) );
  INV_X1 U49585 ( .I(n44041), .ZN(n38094) );
  XOR2_X1 U49586 ( .A1(n38094), .A2(n51278), .Z(n51535) );
  XOR2_X1 U49587 ( .A1(n38095), .A2(n56335), .Z(n38096) );
  XOR2_X1 U49588 ( .A1(n38096), .A2(n51531), .Z(n38097) );
  XOR2_X1 U49589 ( .A1(n51535), .A2(n38097), .Z(n38098) );
  XOR2_X1 U49590 ( .A1(n24018), .A2(n38098), .Z(n38100) );
  XOR2_X1 U49591 ( .A1(n24468), .A2(n38101), .Z(n38102) );
  INV_X1 U49592 ( .I(n38107), .ZN(n38108) );
  XOR2_X1 U49593 ( .A1(n38108), .A2(n56040), .Z(n50958) );
  XOR2_X1 U49594 ( .A1(n29969), .A2(n38109), .Z(n38110) );
  XOR2_X1 U49595 ( .A1(n38111), .A2(n38110), .Z(n50101) );
  XOR2_X1 U49596 ( .A1(n50101), .A2(n50955), .Z(n38112) );
  XOR2_X1 U49597 ( .A1(n50958), .A2(n38112), .Z(n38113) );
  XOR2_X1 U49598 ( .A1(n38158), .A2(n38115), .Z(n38118) );
  XOR2_X1 U49599 ( .A1(n15729), .A2(n15711), .Z(n38119) );
  XOR2_X1 U49600 ( .A1(n60597), .A2(n38120), .Z(n38374) );
  INV_X1 U49601 ( .I(n38374), .ZN(n38122) );
  XOR2_X1 U49602 ( .A1(n38122), .A2(n38121), .Z(n38124) );
  XOR2_X1 U49603 ( .A1(n23332), .A2(n38124), .Z(n38130) );
  INV_X1 U49604 ( .I(n44257), .ZN(n38125) );
  XOR2_X1 U49605 ( .A1(n38125), .A2(n23999), .Z(n52378) );
  XOR2_X1 U49606 ( .A1(n61550), .A2(n56745), .Z(n38127) );
  XOR2_X1 U49607 ( .A1(n38380), .A2(n38127), .Z(n50595) );
  XOR2_X1 U49608 ( .A1(n52378), .A2(n50595), .Z(n38128) );
  XOR2_X1 U49609 ( .A1(n38325), .A2(n38128), .Z(n38129) );
  MUX2_X1 U49611 ( .I0(n38133), .I1(n38132), .S(n41294), .Z(n38137) );
  OAI21_X1 U49612 ( .A1(n64353), .A2(n42199), .B(n42215), .ZN(n38135) );
  INV_X1 U49613 ( .I(n45474), .ZN(n44515) );
  XOR2_X1 U49614 ( .A1(n51494), .A2(n54517), .Z(n51167) );
  XOR2_X1 U49615 ( .A1(n51167), .A2(n51881), .Z(n38138) );
  XOR2_X1 U49616 ( .A1(n44515), .A2(n38138), .Z(n38139) );
  XOR2_X1 U49618 ( .A1(n38146), .A2(n23886), .Z(n50251) );
  XOR2_X1 U49619 ( .A1(n44841), .A2(n53344), .Z(n50910) );
  XOR2_X1 U49620 ( .A1(n50126), .A2(n46682), .Z(n38147) );
  XOR2_X1 U49621 ( .A1(n50910), .A2(n38147), .Z(n38148) );
  XOR2_X1 U49622 ( .A1(n50251), .A2(n38148), .Z(n38149) );
  XOR2_X1 U49623 ( .A1(n20948), .A2(n38149), .Z(n38150) );
  XOR2_X1 U49624 ( .A1(n25769), .A2(n38150), .Z(n38151) );
  INV_X1 U49625 ( .I(n9826), .ZN(n38152) );
  XOR2_X1 U49626 ( .A1(n38153), .A2(n38152), .Z(n51122) );
  INV_X1 U49627 ( .I(n51122), .ZN(n38156) );
  XOR2_X1 U49628 ( .A1(n38154), .A2(n38407), .Z(n38155) );
  XOR2_X1 U49629 ( .A1(n45240), .A2(n38155), .Z(n48387) );
  XOR2_X1 U49631 ( .A1(n38162), .A2(n38161), .Z(n52534) );
  XNOR2_X1 U49632 ( .A1(n54208), .A2(n55833), .ZN(n38163) );
  XOR2_X1 U49633 ( .A1(n55106), .A2(n53705), .Z(n50864) );
  XOR2_X1 U49634 ( .A1(n38163), .A2(n50864), .Z(n38164) );
  XOR2_X1 U49635 ( .A1(n38165), .A2(n38164), .Z(n38166) );
  XOR2_X1 U49636 ( .A1(n52534), .A2(n38166), .Z(n38167) );
  XOR2_X1 U49637 ( .A1(n39284), .A2(n38167), .Z(n38169) );
  XOR2_X1 U49638 ( .A1(n38168), .A2(n38169), .Z(n38172) );
  INV_X1 U49639 ( .I(n38170), .ZN(n38171) );
  XOR2_X1 U49640 ( .A1(n38172), .A2(n38171), .Z(n38174) );
  XOR2_X1 U49641 ( .A1(n38632), .A2(n55379), .Z(n38176) );
  XOR2_X1 U49642 ( .A1(n38177), .A2(n38176), .Z(n51411) );
  XOR2_X1 U49643 ( .A1(n51411), .A2(n52577), .Z(n38178) );
  XOR2_X1 U49644 ( .A1(n24223), .A2(n38182), .Z(n38183) );
  XOR2_X1 U49645 ( .A1(n55534), .A2(n56309), .Z(n38184) );
  XOR2_X1 U49646 ( .A1(n52196), .A2(n38184), .Z(n38185) );
  XOR2_X1 U49647 ( .A1(n38186), .A2(n38185), .Z(n50691) );
  XOR2_X1 U49648 ( .A1(n46415), .A2(n51611), .Z(n52518) );
  XOR2_X1 U49649 ( .A1(n50691), .A2(n52518), .Z(n38187) );
  XOR2_X1 U49650 ( .A1(n22916), .A2(n38187), .Z(n38189) );
  XOR2_X1 U49651 ( .A1(n38189), .A2(n24147), .Z(n38190) );
  XOR2_X1 U49653 ( .A1(n10402), .A2(n61737), .Z(n38192) );
  NOR2_X1 U49656 ( .A1(n41306), .A2(n664), .ZN(n38197) );
  INV_X1 U49659 ( .I(n38203), .ZN(n38204) );
  XOR2_X1 U49660 ( .A1(n1750), .A2(n38207), .Z(n38213) );
  XOR2_X1 U49661 ( .A1(n15710), .A2(n38556), .Z(n49667) );
  XOR2_X1 U49662 ( .A1(n49667), .A2(n51493), .Z(n38208) );
  XOR2_X1 U49663 ( .A1(n50836), .A2(n38208), .Z(n38209) );
  XOR2_X1 U49664 ( .A1(n25277), .A2(n38209), .Z(n38211) );
  XOR2_X1 U49665 ( .A1(n38211), .A2(n38210), .Z(n38212) );
  XOR2_X1 U49666 ( .A1(n45819), .A2(n38885), .Z(n52022) );
  XOR2_X1 U49667 ( .A1(n38215), .A2(n50504), .Z(n49446) );
  XOR2_X1 U49668 ( .A1(n49446), .A2(n24046), .Z(n38216) );
  XOR2_X1 U49669 ( .A1(n52022), .A2(n38216), .Z(n38217) );
  XOR2_X1 U49670 ( .A1(n20948), .A2(n38217), .Z(n38218) );
  XOR2_X1 U49671 ( .A1(n38223), .A2(n38407), .Z(n45378) );
  XOR2_X1 U49672 ( .A1(n45378), .A2(n38224), .Z(n49807) );
  XOR2_X1 U49673 ( .A1(n24011), .A2(n23882), .Z(n38225) );
  XOR2_X1 U49674 ( .A1(n38226), .A2(n38225), .Z(n50874) );
  XOR2_X1 U49675 ( .A1(n49807), .A2(n38227), .Z(n38228) );
  XOR2_X1 U49676 ( .A1(n7713), .A2(n38228), .Z(n38230) );
  INV_X1 U49677 ( .I(n23493), .ZN(n38229) );
  XOR2_X1 U49678 ( .A1(n38230), .A2(n38229), .Z(n38231) );
  XOR2_X1 U49679 ( .A1(n38232), .A2(n38231), .Z(n38233) );
  XOR2_X1 U49681 ( .A1(n38330), .A2(n38806), .Z(n38668) );
  INV_X1 U49682 ( .I(n38235), .ZN(n44137) );
  XOR2_X1 U49683 ( .A1(n50698), .A2(n38236), .Z(n38237) );
  XOR2_X1 U49684 ( .A1(n44137), .A2(n38237), .Z(n50490) );
  XOR2_X1 U49685 ( .A1(n38327), .A2(n38238), .Z(n52410) );
  XOR2_X1 U49686 ( .A1(n50490), .A2(n52410), .Z(n38239) );
  XOR2_X1 U49687 ( .A1(n38668), .A2(n38240), .Z(n38241) );
  XOR2_X1 U49688 ( .A1(n38242), .A2(n38241), .Z(n38243) );
  XOR2_X1 U49689 ( .A1(n39750), .A2(n38243), .Z(n38248) );
  XOR2_X1 U49690 ( .A1(n38871), .A2(n52375), .Z(n38384) );
  INV_X1 U49691 ( .I(n38384), .ZN(n38244) );
  XOR2_X1 U49692 ( .A1(n38990), .A2(n38244), .Z(n38246) );
  XOR2_X1 U49693 ( .A1(n38246), .A2(n38245), .Z(n38247) );
  XOR2_X1 U49694 ( .A1(n38248), .A2(n38247), .Z(n42504) );
  XOR2_X1 U49696 ( .A1(n38952), .A2(n50533), .Z(n38791) );
  XOR2_X1 U49697 ( .A1(n50534), .A2(n51765), .Z(n38249) );
  XOR2_X1 U49698 ( .A1(n38250), .A2(n38249), .Z(n52427) );
  XOR2_X1 U49699 ( .A1(n50536), .A2(n52427), .Z(n38251) );
  XOR2_X1 U49700 ( .A1(n10402), .A2(n38251), .Z(n38252) );
  XOR2_X1 U49701 ( .A1(n233), .A2(n38645), .Z(n38254) );
  XOR2_X1 U49702 ( .A1(n38253), .A2(n38254), .Z(n38255) );
  INV_X1 U49703 ( .I(n39227), .ZN(n38257) );
  XOR2_X1 U49704 ( .A1(n38772), .A2(n54917), .Z(n51276) );
  XOR2_X1 U49705 ( .A1(n51278), .A2(n51276), .Z(n38259) );
  XOR2_X1 U49706 ( .A1(n43262), .A2(n38258), .Z(n51752) );
  XOR2_X1 U49707 ( .A1(n38259), .A2(n51752), .Z(n38260) );
  NAND2_X1 U49710 ( .A1(n41858), .A2(n3534), .ZN(n38266) );
  NAND3_X1 U49711 ( .A1(n22448), .A2(n23744), .A3(n41859), .ZN(n38265) );
  XOR2_X1 U49712 ( .A1(n60207), .A2(n54870), .Z(n38278) );
  XOR2_X1 U49713 ( .A1(n38279), .A2(n38278), .Z(n51247) );
  XOR2_X1 U49714 ( .A1(n38280), .A2(n55034), .Z(n38894) );
  XNOR2_X1 U49715 ( .A1(n51493), .A2(n52970), .ZN(n38281) );
  XOR2_X1 U49716 ( .A1(n38894), .A2(n38281), .Z(n51781) );
  XOR2_X1 U49717 ( .A1(n51247), .A2(n51781), .Z(n38282) );
  XOR2_X1 U49718 ( .A1(n38283), .A2(n38282), .Z(n38284) );
  XOR2_X1 U49719 ( .A1(n38288), .A2(n38287), .Z(n38290) );
  XOR2_X1 U49720 ( .A1(n245), .A2(n23886), .Z(n38293) );
  XOR2_X1 U49721 ( .A1(n756), .A2(n38293), .Z(n38294) );
  XOR2_X1 U49722 ( .A1(n38294), .A2(n51007), .Z(n38295) );
  XOR2_X1 U49723 ( .A1(n38298), .A2(n38297), .Z(n38299) );
  XOR2_X1 U49724 ( .A1(n38302), .A2(n38301), .Z(n52356) );
  XOR2_X1 U49725 ( .A1(n52356), .A2(n50551), .Z(n38303) );
  XOR2_X1 U49726 ( .A1(n20087), .A2(n38303), .Z(n38305) );
  XOR2_X1 U49727 ( .A1(n53945), .A2(n54219), .Z(n38787) );
  XOR2_X1 U49728 ( .A1(n38787), .A2(n24065), .Z(n39262) );
  XOR2_X1 U49729 ( .A1(n39262), .A2(n23989), .Z(n38311) );
  XOR2_X1 U49730 ( .A1(n38311), .A2(n38947), .Z(n38312) );
  XOR2_X1 U49731 ( .A1(n44430), .A2(n38312), .Z(n52082) );
  INV_X1 U49732 ( .I(n51801), .ZN(n38316) );
  XOR2_X1 U49733 ( .A1(n38851), .A2(n51729), .Z(n38315) );
  XOR2_X1 U49734 ( .A1(n38316), .A2(n38315), .Z(n38317) );
  XOR2_X1 U49735 ( .A1(n21098), .A2(n38317), .Z(n38318) );
  INV_X1 U49737 ( .I(n39214), .ZN(n38324) );
  XOR2_X1 U49738 ( .A1(n38325), .A2(n38324), .Z(n38332) );
  XOR2_X1 U49739 ( .A1(n38326), .A2(n50475), .Z(n38328) );
  XOR2_X1 U49740 ( .A1(n38328), .A2(n38327), .Z(n52060) );
  XOR2_X1 U49741 ( .A1(n50790), .A2(n52060), .Z(n38329) );
  XOR2_X1 U49742 ( .A1(n62864), .A2(n38329), .Z(n38331) );
  XOR2_X1 U49743 ( .A1(n63922), .A2(n38333), .Z(n38793) );
  XOR2_X1 U49744 ( .A1(n63081), .A2(n38793), .Z(n38335) );
  OAI22_X1 U49745 ( .A1(n42439), .A2(n11994), .B1(n57208), .B2(n10479), .ZN(
        n38342) );
  AOI22_X1 U49746 ( .A1(n38337), .A2(n41817), .B1(n42431), .B2(n7057), .ZN(
        n38341) );
  NAND3_X1 U49747 ( .A1(n41816), .A2(n42427), .A3(n62291), .ZN(n38340) );
  NOR2_X1 U49748 ( .A1(n43869), .A2(n59476), .ZN(n38347) );
  NAND2_X1 U49749 ( .A1(n6412), .A2(n58262), .ZN(n38343) );
  MUX2_X1 U49750 ( .I0(n41596), .I1(n38347), .S(n65147), .Z(n38359) );
  INV_X1 U49751 ( .I(n38349), .ZN(n38348) );
  NAND2_X1 U49752 ( .A1(n38349), .A2(n59476), .ZN(n38351) );
  INV_X1 U49753 ( .I(n43351), .ZN(n38350) );
  XOR2_X1 U49755 ( .A1(n51531), .A2(n54563), .Z(n38362) );
  XOR2_X1 U49756 ( .A1(n43787), .A2(n38362), .Z(n51623) );
  XOR2_X1 U49757 ( .A1(n43858), .A2(n54185), .Z(n51532) );
  XOR2_X1 U49758 ( .A1(n51623), .A2(n51532), .Z(n38363) );
  XOR2_X1 U49759 ( .A1(n38364), .A2(n38363), .Z(n38365) );
  XOR2_X1 U49760 ( .A1(n38365), .A2(n59895), .Z(n38366) );
  INV_X1 U49761 ( .I(n52425), .ZN(n38369) );
  XOR2_X1 U49762 ( .A1(n30036), .A2(n60857), .Z(n39761) );
  XOR2_X1 U49763 ( .A1(n39761), .A2(n7264), .Z(n38368) );
  XOR2_X1 U49764 ( .A1(n38369), .A2(n38368), .Z(n38370) );
  XOR2_X1 U49765 ( .A1(n25376), .A2(n12669), .Z(n38375) );
  INV_X1 U49766 ( .I(n38378), .ZN(n38379) );
  XOR2_X1 U49767 ( .A1(n53124), .A2(n55903), .Z(n39739) );
  XOR2_X1 U49768 ( .A1(n38379), .A2(n39739), .Z(n50596) );
  XOR2_X1 U49769 ( .A1(n38380), .A2(n23455), .Z(n52376) );
  XOR2_X1 U49770 ( .A1(n50596), .A2(n52376), .Z(n38381) );
  XOR2_X1 U49771 ( .A1(n39275), .A2(n38381), .Z(n38383) );
  XOR2_X1 U49772 ( .A1(n38382), .A2(n38383), .Z(n38385) );
  XOR2_X1 U49773 ( .A1(n38387), .A2(n52226), .Z(n49965) );
  XOR2_X1 U49774 ( .A1(n49965), .A2(n24105), .Z(n38389) );
  XOR2_X1 U49775 ( .A1(n50999), .A2(n38388), .Z(n45141) );
  XOR2_X1 U49776 ( .A1(n38389), .A2(n45141), .Z(n38391) );
  INV_X1 U49777 ( .I(n44999), .ZN(n38390) );
  XOR2_X1 U49778 ( .A1(n38391), .A2(n38390), .Z(n38392) );
  XOR2_X1 U49779 ( .A1(n39253), .A2(n38392), .Z(n38394) );
  INV_X1 U49780 ( .I(n38649), .ZN(n38393) );
  XOR2_X1 U49781 ( .A1(n38393), .A2(n38394), .Z(n38395) );
  XOR2_X1 U49783 ( .A1(n38397), .A2(n39724), .Z(n46154) );
  XOR2_X1 U49784 ( .A1(n46154), .A2(n55368), .Z(n51928) );
  XOR2_X1 U49785 ( .A1(n23858), .A2(n54734), .Z(n38398) );
  XOR2_X1 U49786 ( .A1(n38398), .A2(n24057), .Z(n38399) );
  XOR2_X1 U49787 ( .A1(n38400), .A2(n38399), .Z(n50173) );
  XOR2_X1 U49788 ( .A1(n50173), .A2(n54249), .Z(n38401) );
  XOR2_X1 U49789 ( .A1(n50102), .A2(n49787), .Z(n38409) );
  XOR2_X1 U49790 ( .A1(n38408), .A2(n38407), .Z(n50956) );
  XOR2_X1 U49791 ( .A1(n38409), .A2(n50956), .Z(n38410) );
  XOR2_X1 U49792 ( .A1(n17583), .A2(n15711), .Z(n38412) );
  MUX2_X1 U49795 ( .I0(n38418), .I1(n38417), .S(n39066), .Z(n38419) );
  NAND2_X1 U49796 ( .A1(n38421), .A2(n23355), .ZN(n38424) );
  NAND3_X1 U49797 ( .A1(n7649), .A2(n60928), .A3(n23355), .ZN(n38423) );
  NAND2_X1 U49798 ( .A1(n16601), .A2(n1275), .ZN(n38422) );
  INV_X1 U49799 ( .I(n38428), .ZN(n38435) );
  XOR2_X1 U49800 ( .A1(n46684), .A2(n23858), .Z(n50624) );
  XOR2_X1 U49801 ( .A1(n39469), .A2(n54556), .Z(n52137) );
  XOR2_X1 U49802 ( .A1(n52137), .A2(n56784), .Z(n38429) );
  XOR2_X1 U49803 ( .A1(n50624), .A2(n38429), .Z(n38431) );
  XOR2_X1 U49804 ( .A1(n38431), .A2(n38430), .Z(n38432) );
  XOR2_X1 U49805 ( .A1(n23062), .A2(n38432), .Z(n38434) );
  XOR2_X1 U49806 ( .A1(n8539), .A2(n38436), .Z(n38437) );
  INV_X1 U49807 ( .I(n38438), .ZN(n38439) );
  XOR2_X1 U49808 ( .A1(n38439), .A2(n56827), .Z(n50901) );
  XOR2_X1 U49809 ( .A1(n50901), .A2(n56008), .Z(n38443) );
  XOR2_X1 U49810 ( .A1(n38440), .A2(n53246), .Z(n38442) );
  XOR2_X1 U49811 ( .A1(n38442), .A2(n38441), .Z(n50228) );
  XOR2_X1 U49812 ( .A1(n38443), .A2(n50228), .Z(n38444) );
  XOR2_X1 U49813 ( .A1(n38444), .A2(n20234), .Z(n38445) );
  XOR2_X1 U49814 ( .A1(n45087), .A2(n44533), .Z(n44927) );
  XOR2_X1 U49815 ( .A1(n38448), .A2(n23020), .Z(n38449) );
  XOR2_X1 U49816 ( .A1(n44927), .A2(n38449), .Z(n52634) );
  XOR2_X1 U49817 ( .A1(n38450), .A2(n55655), .Z(n51355) );
  XOR2_X1 U49818 ( .A1(n52634), .A2(n51355), .Z(n38451) );
  INV_X1 U49819 ( .I(n59688), .ZN(n38454) );
  XOR2_X1 U49820 ( .A1(n38453), .A2(n38454), .Z(n38455) );
  INV_X1 U49821 ( .I(n38512), .ZN(n38807) );
  INV_X1 U49823 ( .I(n38949), .ZN(n46129) );
  XOR2_X1 U49824 ( .A1(n46129), .A2(n38459), .Z(n51423) );
  XOR2_X1 U49825 ( .A1(n38460), .A2(n60797), .Z(n38461) );
  XOR2_X1 U49826 ( .A1(n23249), .A2(n38461), .Z(n38462) );
  XOR2_X1 U49827 ( .A1(n51423), .A2(n38462), .Z(n38463) );
  XOR2_X1 U49828 ( .A1(n38530), .A2(n38463), .Z(n38464) );
  XOR2_X1 U49829 ( .A1(n15699), .A2(n38786), .Z(n38467) );
  XOR2_X1 U49830 ( .A1(n50943), .A2(n56949), .Z(n38471) );
  XOR2_X1 U49831 ( .A1(n38472), .A2(n38471), .Z(n38475) );
  XOR2_X1 U49832 ( .A1(n39434), .A2(n51840), .Z(n38474) );
  XOR2_X1 U49833 ( .A1(n50682), .A2(n56879), .Z(n38473) );
  XOR2_X1 U49834 ( .A1(n38474), .A2(n38473), .Z(n51072) );
  XOR2_X1 U49835 ( .A1(n38475), .A2(n51072), .Z(n38476) );
  XOR2_X1 U49836 ( .A1(n38476), .A2(n51656), .Z(n38477) );
  XOR2_X1 U49837 ( .A1(n59680), .A2(n38829), .Z(n38961) );
  INV_X1 U49838 ( .I(n38961), .ZN(n45880) );
  XOR2_X1 U49839 ( .A1(n45880), .A2(n38830), .Z(n50918) );
  XOR2_X1 U49840 ( .A1(n39294), .A2(n24011), .Z(n38481) );
  XOR2_X1 U49841 ( .A1(n49787), .A2(n38481), .Z(n50319) );
  XOR2_X1 U49842 ( .A1(n50918), .A2(n50319), .Z(n38482) );
  XOR2_X1 U49843 ( .A1(n23019), .A2(n38482), .Z(n38483) );
  XOR2_X1 U49844 ( .A1(n2355), .A2(n38483), .Z(n38485) );
  XOR2_X1 U49845 ( .A1(n38485), .A2(n38484), .Z(n38489) );
  XOR2_X1 U49846 ( .A1(n38487), .A2(n38486), .Z(n38488) );
  XOR2_X1 U49847 ( .A1(n38489), .A2(n38488), .Z(n38490) );
  XOR2_X1 U49848 ( .A1(n38491), .A2(n38490), .Z(n38493) );
  INV_X1 U49849 ( .I(n38497), .ZN(n38499) );
  INV_X1 U49850 ( .I(n38502), .ZN(n38504) );
  XOR2_X1 U49851 ( .A1(n22252), .A2(n53308), .Z(n38503) );
  XOR2_X1 U49852 ( .A1(n38504), .A2(n38503), .Z(n51309) );
  XOR2_X1 U49853 ( .A1(n44533), .A2(n54208), .Z(n38505) );
  XOR2_X1 U49854 ( .A1(n38506), .A2(n38505), .Z(n51719) );
  XOR2_X1 U49855 ( .A1(n51309), .A2(n51719), .Z(n38507) );
  XOR2_X1 U49856 ( .A1(n59688), .A2(n24061), .Z(n38511) );
  XOR2_X1 U49857 ( .A1(n38512), .A2(n38511), .Z(n38670) );
  XOR2_X1 U49858 ( .A1(n38670), .A2(n38513), .Z(n38514) );
  INV_X1 U49860 ( .I(n16299), .ZN(n38521) );
  INV_X1 U49861 ( .I(n38517), .ZN(n38519) );
  XOR2_X1 U49862 ( .A1(n51216), .A2(n56949), .Z(n38518) );
  XOR2_X1 U49863 ( .A1(n38519), .A2(n38518), .Z(n38520) );
  XOR2_X1 U49864 ( .A1(n38521), .A2(n38520), .Z(n38522) );
  XOR2_X1 U49865 ( .A1(n38523), .A2(n38522), .Z(n38524) );
  XOR2_X1 U49867 ( .A1(n38532), .A2(n22821), .Z(n51321) );
  XOR2_X1 U49868 ( .A1(n38533), .A2(n51321), .Z(n38534) );
  XOR2_X1 U49869 ( .A1(n10017), .A2(n38534), .Z(n38536) );
  XOR2_X1 U49870 ( .A1(n233), .A2(n38536), .Z(n38538) );
  XOR2_X1 U49871 ( .A1(n38541), .A2(n38540), .Z(n38542) );
  INV_X1 U49872 ( .I(n38544), .ZN(n38545) );
  NOR2_X1 U49873 ( .A1(n38546), .A2(n38545), .ZN(n38547) );
  NAND2_X1 U49874 ( .A1(n38548), .A2(n38547), .ZN(n38564) );
  INV_X1 U49875 ( .I(n38549), .ZN(n38554) );
  AOI21_X1 U49876 ( .A1(n38552), .A2(n7270), .B(n38550), .ZN(n38553) );
  NOR2_X1 U49877 ( .A1(n38554), .A2(n38553), .ZN(n38566) );
  INV_X1 U49878 ( .I(n38555), .ZN(n38557) );
  XOR2_X1 U49879 ( .A1(n38557), .A2(n38556), .Z(n38559) );
  XOR2_X1 U49880 ( .A1(n38558), .A2(n23851), .Z(n39623) );
  XOR2_X1 U49881 ( .A1(n38559), .A2(n39623), .Z(n52011) );
  XOR2_X1 U49882 ( .A1(n38560), .A2(n52900), .Z(n38561) );
  XOR2_X1 U49883 ( .A1(n38562), .A2(n38561), .Z(n49588) );
  XOR2_X1 U49884 ( .A1(n49588), .A2(n56905), .Z(n38563) );
  XOR2_X1 U49885 ( .A1(n52011), .A2(n38563), .Z(n38565) );
  OAI21_X1 U49886 ( .A1(n38564), .A2(n38566), .B(n38565), .ZN(n38571) );
  INV_X1 U49887 ( .I(n38564), .ZN(n38569) );
  INV_X1 U49888 ( .I(n38565), .ZN(n38568) );
  INV_X1 U49889 ( .I(n38566), .ZN(n38567) );
  NAND3_X1 U49890 ( .A1(n38569), .A2(n38568), .A3(n38567), .ZN(n38570) );
  NAND2_X1 U49891 ( .A1(n38571), .A2(n38570), .ZN(n38572) );
  XOR2_X1 U49892 ( .A1(n38577), .A2(n38578), .Z(n38579) );
  INV_X1 U49893 ( .I(n52100), .ZN(n38581) );
  XOR2_X1 U49894 ( .A1(n38581), .A2(n46348), .Z(n42816) );
  XOR2_X1 U49895 ( .A1(n50745), .A2(n56322), .Z(n38582) );
  XOR2_X1 U49896 ( .A1(n52096), .A2(n38582), .Z(n38583) );
  XOR2_X1 U49897 ( .A1(n38583), .A2(n45276), .Z(n38584) );
  XOR2_X1 U49898 ( .A1(n42816), .A2(n38584), .Z(n38585) );
  XOR2_X1 U49899 ( .A1(n10898), .A2(n38585), .Z(n38586) );
  XOR2_X1 U49900 ( .A1(n38588), .A2(n45379), .Z(n52001) );
  XOR2_X1 U49901 ( .A1(n50955), .A2(n55060), .Z(n38589) );
  XOR2_X1 U49902 ( .A1(n52001), .A2(n38589), .Z(n38590) );
  XOR2_X1 U49903 ( .A1(n64241), .A2(n38590), .Z(n38592) );
  XOR2_X1 U49904 ( .A1(n38593), .A2(n38592), .Z(n38595) );
  NAND3_X1 U49905 ( .A1(n38597), .A2(n39123), .A3(n40968), .ZN(n38599) );
  INV_X1 U49906 ( .I(n39058), .ZN(n39139) );
  NAND2_X1 U49908 ( .A1(n39129), .A2(n40523), .ZN(n38601) );
  NAND2_X1 U49909 ( .A1(n40967), .A2(n40619), .ZN(n38602) );
  NAND2_X1 U49910 ( .A1(n25139), .A2(n40613), .ZN(n38606) );
  INV_X1 U49911 ( .I(n40957), .ZN(n38605) );
  OAI21_X1 U49912 ( .A1(n39127), .A2(n38606), .B(n38605), .ZN(n38609) );
  NOR2_X1 U49913 ( .A1(n39130), .A2(n25139), .ZN(n40974) );
  NAND4_X1 U49914 ( .A1(n38612), .A2(n42554), .A3(n1718), .A4(n38611), .ZN(
        n38613) );
  XOR2_X1 U49915 ( .A1(n38614), .A2(n55060), .Z(n49806) );
  XOR2_X1 U49916 ( .A1(n50873), .A2(n49787), .Z(n38615) );
  XOR2_X1 U49917 ( .A1(n49806), .A2(n38615), .Z(n38616) );
  XOR2_X1 U49918 ( .A1(n38617), .A2(n22698), .Z(n38618) );
  XOR2_X1 U49919 ( .A1(n53499), .A2(n56784), .Z(n38624) );
  XOR2_X1 U49920 ( .A1(n38625), .A2(n38624), .Z(n38626) );
  XOR2_X1 U49921 ( .A1(n52020), .A2(n38626), .Z(n38627) );
  XOR2_X1 U49922 ( .A1(n38628), .A2(n38627), .Z(n38629) );
  INV_X1 U49924 ( .I(n51280), .ZN(n46316) );
  XOR2_X1 U49925 ( .A1(n38632), .A2(n38631), .Z(n51751) );
  XOR2_X1 U49926 ( .A1(n51751), .A2(n51275), .Z(n38633) );
  XOR2_X1 U49927 ( .A1(n46316), .A2(n38633), .Z(n38634) );
  XOR2_X1 U49928 ( .A1(n38638), .A2(n54219), .Z(n50537) );
  XOR2_X1 U49929 ( .A1(n38639), .A2(n29407), .Z(n38640) );
  XOR2_X1 U49930 ( .A1(n52425), .A2(n38640), .Z(n38641) );
  XOR2_X1 U49931 ( .A1(n50537), .A2(n38641), .Z(n38642) );
  XOR2_X1 U49932 ( .A1(n38916), .A2(n38642), .Z(n38644) );
  XOR2_X1 U49933 ( .A1(n38643), .A2(n38644), .Z(n38647) );
  XOR2_X1 U49934 ( .A1(n38645), .A2(n9398), .Z(n38646) );
  INV_X1 U49935 ( .I(n38650), .ZN(n38652) );
  XOR2_X1 U49936 ( .A1(n38652), .A2(n60799), .Z(n49669) );
  XOR2_X1 U49937 ( .A1(n38653), .A2(n53318), .Z(n38654) );
  XOR2_X1 U49938 ( .A1(n38997), .A2(n38654), .Z(n50834) );
  XOR2_X1 U49939 ( .A1(n54360), .A2(n55118), .Z(n43642) );
  XOR2_X1 U49940 ( .A1(n50834), .A2(n43642), .Z(n38655) );
  XOR2_X1 U49942 ( .A1(n4762), .A2(n38659), .Z(n38660) );
  XOR2_X1 U49943 ( .A1(n38660), .A2(n38741), .Z(n38803) );
  INV_X1 U49944 ( .I(n38662), .ZN(n38664) );
  XOR2_X1 U49945 ( .A1(n51814), .A2(n56124), .Z(n38663) );
  XOR2_X1 U49946 ( .A1(n38664), .A2(n38663), .Z(n52411) );
  XOR2_X1 U49947 ( .A1(n38665), .A2(n56976), .Z(n50488) );
  XOR2_X1 U49948 ( .A1(n52411), .A2(n50488), .Z(n38666) );
  XOR2_X1 U49949 ( .A1(n63922), .A2(n38667), .Z(n38669) );
  XOR2_X1 U49950 ( .A1(n38669), .A2(n38668), .Z(n38671) );
  NOR2_X1 U49951 ( .A1(n41198), .A2(n60567), .ZN(n38676) );
  NOR2_X1 U49952 ( .A1(n40628), .A2(n40728), .ZN(n38674) );
  INV_X1 U49955 ( .I(n61407), .ZN(n38678) );
  NOR2_X1 U49958 ( .A1(n42555), .A2(n1269), .ZN(n38686) );
  NAND2_X1 U49961 ( .A1(n41198), .A2(n40634), .ZN(n38689) );
  INV_X1 U49962 ( .I(n41188), .ZN(n38690) );
  OAI21_X1 U49964 ( .A1(n14462), .A2(n10587), .B(n41167), .ZN(n38693) );
  AOI21_X1 U49965 ( .A1(n40542), .A2(n40645), .B(n39074), .ZN(n38695) );
  INV_X1 U49966 ( .I(n38698), .ZN(n40918) );
  XOR2_X1 U49967 ( .A1(n39376), .A2(n63603), .Z(n51497) );
  XOR2_X1 U49968 ( .A1(n51497), .A2(n39478), .Z(n38700) );
  XOR2_X1 U49969 ( .A1(n40918), .A2(n38700), .Z(n38701) );
  XOR2_X1 U49970 ( .A1(n23199), .A2(n38701), .Z(n38703) );
  XOR2_X1 U49971 ( .A1(n38704), .A2(n38703), .Z(n38705) );
  XOR2_X1 U49972 ( .A1(n38705), .A2(n39528), .Z(n38706) );
  INV_X1 U49973 ( .I(n23949), .ZN(n38710) );
  XOR2_X1 U49974 ( .A1(n38713), .A2(n15712), .Z(n47341) );
  XOR2_X1 U49975 ( .A1(n39362), .A2(n44378), .Z(n38714) );
  XOR2_X1 U49976 ( .A1(n38714), .A2(n46398), .Z(n51173) );
  XOR2_X1 U49977 ( .A1(n47341), .A2(n51173), .Z(n38715) );
  XOR2_X1 U49979 ( .A1(n38720), .A2(n39558), .Z(n50182) );
  XOR2_X1 U49980 ( .A1(n38721), .A2(n13114), .Z(n38722) );
  XOR2_X1 U49981 ( .A1(n38723), .A2(n38722), .Z(n51953) );
  XOR2_X1 U49982 ( .A1(n50182), .A2(n51953), .Z(n38724) );
  XOR2_X1 U49983 ( .A1(n11534), .A2(n38724), .Z(n38725) );
  INV_X1 U49984 ( .I(n38727), .ZN(n38728) );
  XOR2_X1 U49986 ( .A1(n24189), .A2(n22698), .Z(n38738) );
  INV_X1 U49987 ( .I(n38732), .ZN(n51516) );
  XOR2_X1 U49988 ( .A1(n38734), .A2(n38733), .Z(n38735) );
  XOR2_X1 U49989 ( .A1(n38735), .A2(n53138), .Z(n51578) );
  XOR2_X1 U49990 ( .A1(n51516), .A2(n51578), .Z(n38736) );
  XOR2_X1 U49991 ( .A1(n23019), .A2(n38736), .Z(n38737) );
  XOR2_X1 U49992 ( .A1(n38738), .A2(n38737), .Z(n38739) );
  XOR2_X1 U49993 ( .A1(n64786), .A2(n38741), .Z(n39466) );
  XOR2_X1 U49994 ( .A1(n39214), .A2(n53375), .Z(n39454) );
  XOR2_X1 U49995 ( .A1(n38743), .A2(n52232), .Z(n45868) );
  XOR2_X1 U49996 ( .A1(n39454), .A2(n45868), .Z(n39595) );
  XOR2_X1 U49998 ( .A1(n50197), .A2(n54587), .Z(n38746) );
  XOR2_X1 U49999 ( .A1(n43497), .A2(n38746), .Z(n38747) );
  XOR2_X1 U50000 ( .A1(n4762), .A2(n38747), .Z(n38748) );
  INV_X1 U50001 ( .I(n38989), .ZN(n38795) );
  XOR2_X1 U50002 ( .A1(n38748), .A2(n38795), .Z(n38749) );
  XOR2_X1 U50004 ( .A1(n53989), .A2(n51261), .Z(n46315) );
  XOR2_X1 U50005 ( .A1(n46315), .A2(n38752), .Z(n52500) );
  XOR2_X1 U50006 ( .A1(n52470), .A2(n50682), .Z(n38753) );
  XOR2_X1 U50007 ( .A1(n52500), .A2(n38753), .Z(n38754) );
  NAND2_X1 U50008 ( .A1(n25131), .A2(n62611), .ZN(n38760) );
  OAI22_X1 U50009 ( .A1(n64308), .A2(n8942), .B1(n61561), .B2(n38760), .ZN(
        n38761) );
  NAND2_X1 U50010 ( .A1(n40748), .A2(n24982), .ZN(n38763) );
  NAND3_X1 U50012 ( .A1(n38764), .A2(n41470), .A3(n7165), .ZN(n38768) );
  NAND3_X1 U50013 ( .A1(n40761), .A2(n25131), .A3(n24649), .ZN(n38767) );
  XOR2_X1 U50014 ( .A1(n38772), .A2(n24109), .Z(n38773) );
  XOR2_X1 U50015 ( .A1(n38774), .A2(n38773), .Z(n52579) );
  XOR2_X1 U50016 ( .A1(n44613), .A2(n57989), .Z(n51408) );
  XOR2_X1 U50017 ( .A1(n51979), .A2(n51408), .Z(n38775) );
  XOR2_X1 U50018 ( .A1(n52579), .A2(n38775), .Z(n38776) );
  XOR2_X1 U50019 ( .A1(n38777), .A2(n38776), .Z(n38778) );
  XOR2_X1 U50020 ( .A1(n24151), .A2(n52513), .Z(n38782) );
  XOR2_X1 U50021 ( .A1(n61238), .A2(n43882), .Z(n52516) );
  XOR2_X1 U50022 ( .A1(n60556), .A2(n52516), .Z(n38788) );
  XOR2_X1 U50023 ( .A1(n45131), .A2(n38787), .Z(n50690) );
  XOR2_X1 U50024 ( .A1(n38788), .A2(n50690), .Z(n38789) );
  XOR2_X1 U50025 ( .A1(n1337), .A2(n38789), .Z(n38790) );
  XOR2_X1 U50026 ( .A1(n38791), .A2(n38790), .Z(n38792) );
  XOR2_X1 U50027 ( .A1(n60597), .A2(n38795), .Z(n38802) );
  XOR2_X1 U50028 ( .A1(n24098), .A2(n57162), .Z(n38797) );
  XOR2_X1 U50029 ( .A1(n38798), .A2(n38797), .Z(n52533) );
  XOR2_X1 U50030 ( .A1(n52533), .A2(n54936), .Z(n38799) );
  XOR2_X1 U50031 ( .A1(n50701), .A2(n38799), .Z(n38800) );
  XOR2_X1 U50032 ( .A1(n39284), .A2(n38800), .Z(n38801) );
  XOR2_X1 U50033 ( .A1(n38802), .A2(n38801), .Z(n38804) );
  XOR2_X1 U50034 ( .A1(n38804), .A2(n38803), .Z(n38805) );
  XOR2_X1 U50035 ( .A1(n38805), .A2(n39209), .Z(n38810) );
  XOR2_X1 U50036 ( .A1(n38986), .A2(n38808), .Z(n38809) );
  XOR2_X1 U50037 ( .A1(n38810), .A2(n38809), .Z(n38811) );
  XOR2_X1 U50039 ( .A1(n56702), .A2(n56180), .Z(n38813) );
  XOR2_X1 U50040 ( .A1(n38813), .A2(n53154), .Z(n38814) );
  XOR2_X1 U50041 ( .A1(n49445), .A2(n38814), .Z(n38815) );
  XOR2_X1 U50042 ( .A1(n52100), .A2(n38815), .Z(n38816) );
  XOR2_X1 U50043 ( .A1(n23429), .A2(n38816), .Z(n38817) );
  XOR2_X1 U50044 ( .A1(n38821), .A2(n39208), .Z(n38823) );
  INV_X1 U50045 ( .I(n38824), .ZN(n51169) );
  XOR2_X1 U50046 ( .A1(n38826), .A2(n38825), .Z(n45471) );
  XOR2_X1 U50047 ( .A1(n38829), .A2(n54536), .Z(n38831) );
  XOR2_X1 U50048 ( .A1(n38831), .A2(n38830), .Z(n51121) );
  XOR2_X1 U50049 ( .A1(n51121), .A2(n51019), .Z(n38832) );
  INV_X1 U50050 ( .I(n48388), .ZN(n44962) );
  XOR2_X1 U50051 ( .A1(n38832), .A2(n44962), .Z(n38833) );
  XOR2_X1 U50052 ( .A1(n17347), .A2(n9896), .Z(n38837) );
  NAND3_X1 U50053 ( .A1(n41462), .A2(n60810), .A3(n39019), .ZN(n38840) );
  OAI22_X1 U50054 ( .A1(n39019), .A2(n25777), .B1(n38841), .B2(n41455), .ZN(
        n38842) );
  NAND2_X1 U50055 ( .A1(n38842), .A2(n41149), .ZN(n38846) );
  NAND3_X1 U50057 ( .A1(n25777), .A2(n1516), .A3(n40713), .ZN(n38844) );
  NAND2_X1 U50058 ( .A1(n41457), .A2(n38844), .ZN(n38845) );
  XOR2_X1 U50059 ( .A1(n38849), .A2(n23019), .Z(n39673) );
  XOR2_X1 U50060 ( .A1(n38850), .A2(n55546), .Z(n51642) );
  XOR2_X1 U50061 ( .A1(n38851), .A2(n51021), .Z(n51187) );
  XOR2_X1 U50062 ( .A1(n56475), .A2(n53138), .Z(n38852) );
  XOR2_X1 U50063 ( .A1(n51999), .A2(n38852), .Z(n38853) );
  XOR2_X1 U50064 ( .A1(n51187), .A2(n38853), .Z(n38854) );
  XOR2_X1 U50065 ( .A1(n39299), .A2(n38857), .Z(n38858) );
  XOR2_X1 U50066 ( .A1(n38859), .A2(n38858), .Z(n38860) );
  XOR2_X1 U50067 ( .A1(n38980), .A2(n38862), .Z(n52168) );
  XOR2_X1 U50068 ( .A1(n54289), .A2(n54587), .Z(n38863) );
  XOR2_X1 U50069 ( .A1(n52168), .A2(n38863), .Z(n38864) );
  XOR2_X1 U50070 ( .A1(n50618), .A2(n38864), .Z(n38865) );
  XOR2_X1 U50071 ( .A1(n23573), .A2(n38865), .Z(n38869) );
  XOR2_X1 U50072 ( .A1(n38866), .A2(n38867), .Z(n38868) );
  XOR2_X1 U50073 ( .A1(n22485), .A2(n204), .Z(n38872) );
  XOR2_X1 U50074 ( .A1(n38873), .A2(n38872), .Z(n38874) );
  XOR2_X1 U50076 ( .A1(n245), .A2(n46348), .Z(n38881) );
  XOR2_X1 U50077 ( .A1(n38881), .A2(n46682), .Z(n38883) );
  XOR2_X1 U50078 ( .A1(n38883), .A2(n38882), .Z(n50845) );
  XOR2_X1 U50079 ( .A1(n53154), .A2(n53344), .Z(n38884) );
  XOR2_X1 U50080 ( .A1(n38884), .A2(n4561), .Z(n38886) );
  XOR2_X1 U50081 ( .A1(n38886), .A2(n38885), .Z(n49691) );
  XOR2_X1 U50082 ( .A1(n50845), .A2(n49691), .Z(n38887) );
  XOR2_X1 U50083 ( .A1(n23429), .A2(n38887), .Z(n38888) );
  INV_X1 U50084 ( .I(n38893), .ZN(n38895) );
  XOR2_X1 U50085 ( .A1(n38895), .A2(n38894), .Z(n51037) );
  XOR2_X1 U50086 ( .A1(n38896), .A2(n55118), .Z(n38897) );
  XOR2_X1 U50087 ( .A1(n38898), .A2(n38897), .Z(n51694) );
  XOR2_X1 U50088 ( .A1(n51037), .A2(n51694), .Z(n38899) );
  XOR2_X1 U50089 ( .A1(n39626), .A2(n38899), .Z(n38900) );
  XOR2_X1 U50090 ( .A1(n38900), .A2(n21348), .Z(n38902) );
  XOR2_X1 U50091 ( .A1(n52463), .A2(n56508), .Z(n38905) );
  XOR2_X1 U50092 ( .A1(n38904), .A2(n53359), .Z(n50513) );
  XOR2_X1 U50093 ( .A1(n38905), .A2(n50513), .Z(n38906) );
  XOR2_X1 U50094 ( .A1(n24276), .A2(n38906), .Z(n38908) );
  XOR2_X1 U50095 ( .A1(n1337), .A2(n8984), .Z(n38954) );
  XOR2_X1 U50096 ( .A1(n50025), .A2(n54219), .Z(n38914) );
  XOR2_X1 U50097 ( .A1(n39558), .A2(n38914), .Z(n50664) );
  XOR2_X1 U50098 ( .A1(n50664), .A2(n52196), .Z(n38915) );
  XOR2_X1 U50099 ( .A1(n38916), .A2(n38915), .Z(n38917) );
  XOR2_X1 U50100 ( .A1(n38954), .A2(n38917), .Z(n38918) );
  NOR2_X2 U50101 ( .A1(n1743), .A2(n40770), .ZN(n41425) );
  INV_X1 U50102 ( .I(n40401), .ZN(n38925) );
  NAND2_X1 U50103 ( .A1(n40400), .A2(n10173), .ZN(n38927) );
  NAND2_X1 U50104 ( .A1(n38935), .A2(n65184), .ZN(n39863) );
  AOI21_X1 U50105 ( .A1(n38928), .A2(n38927), .B(n39863), .ZN(n38929) );
  NOR2_X1 U50106 ( .A1(n38930), .A2(n38929), .ZN(n38940) );
  NOR2_X1 U50108 ( .A1(n65184), .A2(n64364), .ZN(n38938) );
  NAND2_X1 U50109 ( .A1(n61094), .A2(n40403), .ZN(n38936) );
  INV_X1 U50110 ( .I(n45126), .ZN(n44617) );
  XOR2_X1 U50111 ( .A1(n44617), .A2(n53359), .Z(n50554) );
  XOR2_X1 U50112 ( .A1(n50554), .A2(n54917), .Z(n38944) );
  XOR2_X1 U50113 ( .A1(n38948), .A2(n38947), .Z(n38950) );
  XOR2_X1 U50114 ( .A1(n38950), .A2(n38949), .Z(n50800) );
  XOR2_X1 U50115 ( .A1(n50800), .A2(n52080), .Z(n38951) );
  XOR2_X1 U50116 ( .A1(n38952), .A2(n38951), .Z(n38953) );
  XOR2_X1 U50117 ( .A1(n38954), .A2(n38953), .Z(n38955) );
  INV_X1 U50118 ( .I(n11142), .ZN(n38956) );
  XOR2_X1 U50119 ( .A1(n38958), .A2(n38957), .Z(n38959) );
  XOR2_X1 U50120 ( .A1(n38961), .A2(n53262), .Z(n51188) );
  XOR2_X1 U50121 ( .A1(n38962), .A2(n56859), .Z(n51800) );
  XOR2_X1 U50122 ( .A1(n51021), .A2(n51019), .Z(n38963) );
  XOR2_X1 U50123 ( .A1(n51800), .A2(n38963), .Z(n38964) );
  XOR2_X1 U50124 ( .A1(n4563), .A2(n38966), .Z(n38967) );
  XOR2_X1 U50125 ( .A1(n50909), .A2(n57131), .Z(n38969) );
  XOR2_X1 U50126 ( .A1(n9753), .A2(n38969), .Z(n38970) );
  XOR2_X1 U50127 ( .A1(n50129), .A2(n38970), .Z(n38971) );
  XOR2_X1 U50128 ( .A1(n23429), .A2(n38971), .Z(n38974) );
  XOR2_X1 U50129 ( .A1(n38974), .A2(n38973), .Z(n38975) );
  XOR2_X1 U50130 ( .A1(n22323), .A2(n4561), .Z(n50125) );
  XOR2_X1 U50131 ( .A1(n50125), .A2(n54249), .Z(n38978) );
  XOR2_X1 U50132 ( .A1(n23020), .A2(n38980), .Z(n38982) );
  XOR2_X1 U50133 ( .A1(n51992), .A2(n38982), .Z(n52061) );
  XOR2_X1 U50134 ( .A1(n50197), .A2(n54936), .Z(n50788) );
  XOR2_X1 U50135 ( .A1(n50788), .A2(n55903), .Z(n38983) );
  XOR2_X1 U50136 ( .A1(n52061), .A2(n38983), .Z(n38984) );
  XOR2_X1 U50137 ( .A1(n23573), .A2(n38984), .Z(n38985) );
  INV_X1 U50138 ( .I(n51494), .ZN(n38993) );
  XOR2_X1 U50139 ( .A1(n38996), .A2(n38995), .Z(n51782) );
  XOR2_X1 U50140 ( .A1(n38997), .A2(n39196), .Z(n51244) );
  XOR2_X1 U50141 ( .A1(n51782), .A2(n51244), .Z(n38998) );
  XOR2_X1 U50142 ( .A1(n38999), .A2(n38998), .Z(n39000) );
  XOR2_X1 U50143 ( .A1(n39002), .A2(n39625), .Z(n39003) );
  OAI21_X1 U50144 ( .A1(n60132), .A2(n41397), .B(n21471), .ZN(n39008) );
  NAND2_X1 U50145 ( .A1(n41239), .A2(n17063), .ZN(n39053) );
  OAI22_X1 U50146 ( .A1(n41399), .A2(n39008), .B1(n23780), .B2(n39053), .ZN(
        n39010) );
  OAI21_X1 U50147 ( .A1(n42542), .A2(n42931), .B(n57557), .ZN(n39013) );
  INV_X1 U50148 ( .I(n41454), .ZN(n39017) );
  NOR2_X1 U50149 ( .A1(n64366), .A2(n41453), .ZN(n39016) );
  INV_X1 U50150 ( .I(n41451), .ZN(n39023) );
  INV_X1 U50152 ( .I(n39025), .ZN(n39026) );
  NAND2_X1 U50153 ( .A1(n40723), .A2(n39026), .ZN(n39034) );
  AOI22_X1 U50155 ( .A1(n61407), .A2(n40633), .B1(n38675), .B2(n39028), .ZN(
        n39032) );
  NOR2_X1 U50159 ( .A1(n1404), .A2(n39040), .ZN(n39043) );
  NOR2_X1 U50161 ( .A1(n5774), .A2(n15723), .ZN(n39041) );
  NAND2_X1 U50164 ( .A1(n11472), .A2(n39007), .ZN(n39047) );
  OAI21_X1 U50165 ( .A1(n41236), .A2(n23780), .B(n41411), .ZN(n39049) );
  NAND2_X1 U50167 ( .A1(n39050), .A2(n24523), .ZN(n39051) );
  INV_X1 U50170 ( .I(n40522), .ZN(n39059) );
  NOR2_X1 U50173 ( .A1(n41670), .A2(n42788), .ZN(n39080) );
  NAND3_X1 U50174 ( .A1(n41159), .A2(n7012), .A3(n39066), .ZN(n39079) );
  NOR2_X1 U50175 ( .A1(n39072), .A2(n59252), .ZN(n39071) );
  INV_X1 U50176 ( .I(n41167), .ZN(n39067) );
  NAND2_X1 U50183 ( .A1(n39086), .A2(n61344), .ZN(n39083) );
  OAI21_X1 U50185 ( .A1(n42775), .A2(n40912), .B(n40914), .ZN(n39089) );
  NAND3_X1 U50186 ( .A1(n42788), .A2(n39087), .A3(n41660), .ZN(n39088) );
  NOR2_X1 U50189 ( .A1(n39100), .A2(n19148), .ZN(n39101) );
  INV_X1 U50193 ( .I(n39106), .ZN(n40117) );
  NOR2_X1 U50194 ( .A1(n40117), .A2(n10341), .ZN(n39107) );
  NOR2_X1 U50196 ( .A1(n19277), .A2(n39111), .ZN(n39114) );
  INV_X1 U50197 ( .I(n40205), .ZN(n39112) );
  NAND2_X1 U50198 ( .A1(n19148), .A2(n39112), .ZN(n39113) );
  OAI21_X1 U50200 ( .A1(n1275), .A2(n25201), .B(n37532), .ZN(n39120) );
  NAND3_X1 U50202 ( .A1(n39129), .A2(n39123), .A3(n40968), .ZN(n39125) );
  NAND2_X1 U50203 ( .A1(n40617), .A2(n38607), .ZN(n39128) );
  INV_X1 U50205 ( .I(n40532), .ZN(n39126) );
  OAI22_X1 U50206 ( .A1(n40622), .A2(n39128), .B1(n39127), .B2(n39126), .ZN(
        n39135) );
  INV_X1 U50207 ( .I(n40619), .ZN(n40531) );
  NAND3_X1 U50208 ( .A1(n64571), .A2(n40523), .A3(n40617), .ZN(n39133) );
  INV_X1 U50209 ( .I(n39129), .ZN(n39131) );
  NAND3_X1 U50210 ( .A1(n39131), .A2(n39130), .A3(n40523), .ZN(n39132) );
  OAI21_X1 U50211 ( .A1(n40619), .A2(n39133), .B(n39132), .ZN(n39134) );
  NOR2_X1 U50212 ( .A1(n39135), .A2(n39134), .ZN(n39140) );
  INV_X1 U50213 ( .I(n39141), .ZN(n39142) );
  OAI21_X1 U50216 ( .A1(n40494), .A2(n9915), .B(n9711), .ZN(n39151) );
  NOR2_X1 U50217 ( .A1(n39146), .A2(n41182), .ZN(n40658) );
  NAND2_X1 U50218 ( .A1(n40658), .A2(n23616), .ZN(n39150) );
  NAND2_X1 U50219 ( .A1(n40656), .A2(n39147), .ZN(n39148) );
  NAND4_X1 U50221 ( .A1(n39152), .A2(n39151), .A3(n39150), .A4(n39149), .ZN(
        n39153) );
  NAND3_X1 U50222 ( .A1(n40939), .A2(n40470), .A3(n9969), .ZN(n39161) );
  NOR2_X1 U50223 ( .A1(n40923), .A2(n9969), .ZN(n40256) );
  NAND2_X1 U50224 ( .A1(n39158), .A2(n40256), .ZN(n39160) );
  NAND2_X1 U50225 ( .A1(n39164), .A2(n40923), .ZN(n39159) );
  NAND2_X1 U50226 ( .A1(n39163), .A2(n62157), .ZN(n39168) );
  NAND3_X1 U50227 ( .A1(n61159), .A2(n40472), .A3(n40477), .ZN(n39167) );
  NOR2_X1 U50229 ( .A1(n43015), .A2(n43017), .ZN(n39173) );
  NAND3_X1 U50230 ( .A1(n43016), .A2(n42001), .A3(n60792), .ZN(n39171) );
  NAND2_X1 U50231 ( .A1(n43016), .A2(n42329), .ZN(n39170) );
  MUX2_X1 U50233 ( .I0(n23184), .I1(n42324), .S(n42327), .Z(n39177) );
  NOR2_X1 U50234 ( .A1(n42327), .A2(n23425), .ZN(n41677) );
  INV_X1 U50235 ( .I(n41677), .ZN(n39176) );
  NAND4_X1 U50236 ( .A1(n39177), .A2(n42328), .A3(n39176), .A4(n42332), .ZN(
        n39178) );
  XOR2_X1 U50237 ( .A1(n50909), .A2(n22773), .Z(n39180) );
  XOR2_X1 U50238 ( .A1(n39181), .A2(n39180), .Z(n39182) );
  XOR2_X1 U50239 ( .A1(n44470), .A2(n39182), .Z(n49693) );
  XOR2_X1 U50240 ( .A1(n39183), .A2(n52095), .Z(n39184) );
  XOR2_X1 U50241 ( .A1(n49693), .A2(n39184), .Z(n39185) );
  XOR2_X1 U50242 ( .A1(n61489), .A2(n39185), .Z(n39187) );
  INV_X1 U50243 ( .I(n39194), .ZN(n39199) );
  XOR2_X1 U50244 ( .A1(n39196), .A2(n39195), .Z(n39197) );
  XOR2_X1 U50245 ( .A1(n39197), .A2(n44995), .Z(n39198) );
  XOR2_X1 U50246 ( .A1(n39199), .A2(n39198), .Z(n51696) );
  XOR2_X1 U50247 ( .A1(n39200), .A2(n55840), .Z(n51038) );
  XOR2_X1 U50248 ( .A1(n51038), .A2(n50832), .Z(n39201) );
  XOR2_X1 U50249 ( .A1(n51696), .A2(n39201), .Z(n39202) );
  XOR2_X1 U50250 ( .A1(n9956), .A2(n39202), .Z(n39203) );
  INV_X1 U50251 ( .I(n52169), .ZN(n46375) );
  XOR2_X1 U50252 ( .A1(n44461), .A2(n39210), .Z(n50617) );
  XOR2_X1 U50253 ( .A1(n46375), .A2(n50617), .Z(n39211) );
  XOR2_X1 U50254 ( .A1(n39214), .A2(n22855), .Z(n39287) );
  INV_X1 U50255 ( .I(n39287), .ZN(n39215) );
  XOR2_X1 U50256 ( .A1(n39733), .A2(n51913), .Z(n39405) );
  XOR2_X1 U50257 ( .A1(n39218), .A2(n39217), .Z(n51020) );
  XOR2_X1 U50258 ( .A1(n39219), .A2(n56915), .Z(n51640) );
  XOR2_X1 U50259 ( .A1(n51020), .A2(n51640), .Z(n39220) );
  XOR2_X1 U50260 ( .A1(n44041), .A2(n39228), .Z(n50514) );
  INV_X1 U50261 ( .I(n50666), .ZN(n43683) );
  XOR2_X1 U50262 ( .A1(n39235), .A2(n23989), .Z(n52199) );
  INV_X1 U50264 ( .I(n39243), .ZN(n39244) );
  XOR2_X1 U50265 ( .A1(n46245), .A2(n52137), .Z(n51794) );
  XOR2_X1 U50266 ( .A1(n39244), .A2(n51794), .Z(n39245) );
  INV_X1 U50267 ( .I(n51735), .ZN(n39251) );
  XOR2_X1 U50268 ( .A1(n52149), .A2(n24044), .Z(n39250) );
  XOR2_X1 U50269 ( .A1(n39251), .A2(n39250), .Z(n39252) );
  XOR2_X1 U50270 ( .A1(n39253), .A2(n39252), .Z(n39256) );
  INV_X1 U50271 ( .I(n49233), .ZN(n39264) );
  XOR2_X1 U50272 ( .A1(n39263), .A2(n39262), .Z(n51967) );
  XOR2_X1 U50273 ( .A1(n39264), .A2(n51967), .Z(n39265) );
  XOR2_X1 U50276 ( .A1(n39268), .A2(n39267), .Z(n39269) );
  XOR2_X1 U50277 ( .A1(n39348), .A2(n39269), .Z(n39271) );
  XOR2_X1 U50279 ( .A1(n63922), .A2(n39275), .Z(n39277) );
  XOR2_X1 U50280 ( .A1(n39278), .A2(n58077), .Z(n49292) );
  XOR2_X1 U50281 ( .A1(n39280), .A2(n39279), .Z(n39282) );
  INV_X1 U50282 ( .I(n44924), .ZN(n39281) );
  XOR2_X1 U50283 ( .A1(n39282), .A2(n39281), .Z(n51993) );
  XOR2_X1 U50284 ( .A1(n49292), .A2(n51993), .Z(n39283) );
  XOR2_X1 U50285 ( .A1(n39284), .A2(n39283), .Z(n39285) );
  XOR2_X1 U50286 ( .A1(n39286), .A2(n39287), .Z(n39288) );
  XOR2_X1 U50287 ( .A1(n51122), .A2(n39294), .Z(n51304) );
  XOR2_X1 U50288 ( .A1(n39295), .A2(n56165), .Z(n51723) );
  XOR2_X1 U50289 ( .A1(n51723), .A2(n51729), .Z(n39296) );
  XOR2_X1 U50290 ( .A1(n51304), .A2(n39296), .Z(n39297) );
  XOR2_X1 U50291 ( .A1(n39298), .A2(n39299), .Z(n39301) );
  XOR2_X1 U50292 ( .A1(n39301), .A2(n39300), .Z(n39302) );
  XOR2_X1 U50293 ( .A1(n39303), .A2(n39302), .Z(n39304) );
  XOR2_X1 U50294 ( .A1(n39305), .A2(n39304), .Z(n39306) );
  INV_X1 U50295 ( .I(n50772), .ZN(n39308) );
  XOR2_X1 U50296 ( .A1(n39308), .A2(n52069), .Z(n39309) );
  XOR2_X1 U50297 ( .A1(n7370), .A2(n39309), .Z(n39311) );
  XOR2_X1 U50298 ( .A1(n39357), .A2(n39311), .Z(n39313) );
  NOR3_X1 U50299 ( .A1(n40139), .A2(n40133), .A3(n64613), .ZN(n39318) );
  NAND2_X1 U50301 ( .A1(n4364), .A2(n40028), .ZN(n39319) );
  NOR2_X1 U50302 ( .A1(n40297), .A2(n57955), .ZN(n39320) );
  NAND2_X1 U50303 ( .A1(n40306), .A2(n40133), .ZN(n40140) );
  NAND3_X1 U50306 ( .A1(n40147), .A2(n40150), .A3(n6768), .ZN(n39328) );
  INV_X1 U50307 ( .I(n39332), .ZN(n39333) );
  XOR2_X1 U50308 ( .A1(n39333), .A2(n55862), .Z(n51954) );
  XOR2_X1 U50309 ( .A1(n39335), .A2(n39334), .Z(n50181) );
  XOR2_X1 U50310 ( .A1(n51954), .A2(n50181), .Z(n39336) );
  INV_X1 U50311 ( .I(n39337), .ZN(n39338) );
  XOR2_X1 U50312 ( .A1(n39339), .A2(n39338), .Z(n39341) );
  XOR2_X1 U50313 ( .A1(n23927), .A2(n15704), .Z(n39347) );
  XOR2_X1 U50314 ( .A1(n39350), .A2(n39349), .Z(n50684) );
  XOR2_X1 U50315 ( .A1(n50646), .A2(n51261), .Z(n39351) );
  XOR2_X1 U50316 ( .A1(n50684), .A2(n39351), .Z(n39353) );
  XOR2_X1 U50317 ( .A1(n51978), .A2(n39352), .Z(n52502) );
  XOR2_X1 U50318 ( .A1(n39353), .A2(n52502), .Z(n39354) );
  XOR2_X1 U50319 ( .A1(n45359), .A2(n39360), .Z(n51174) );
  XOR2_X1 U50320 ( .A1(n39362), .A2(n39361), .Z(n44621) );
  XOR2_X1 U50321 ( .A1(n44621), .A2(n39363), .Z(n47340) );
  XOR2_X1 U50322 ( .A1(n51174), .A2(n47340), .Z(n39364) );
  XOR2_X1 U50323 ( .A1(n2334), .A2(n39364), .Z(n39366) );
  XOR2_X1 U50324 ( .A1(n39366), .A2(n23790), .Z(n39367) );
  XOR2_X1 U50325 ( .A1(n39374), .A2(n39373), .Z(n51499) );
  XOR2_X1 U50326 ( .A1(n39376), .A2(n39375), .Z(n51585) );
  XOR2_X1 U50327 ( .A1(n51585), .A2(n39377), .Z(n39378) );
  XOR2_X1 U50328 ( .A1(n51499), .A2(n39378), .Z(n39379) );
  INV_X1 U50329 ( .I(n59680), .ZN(n39389) );
  XOR2_X1 U50330 ( .A1(n31347), .A2(n45379), .Z(n39388) );
  XOR2_X1 U50331 ( .A1(n39389), .A2(n39388), .Z(n51579) );
  XOR2_X1 U50332 ( .A1(n51579), .A2(n51514), .Z(n39390) );
  XOR2_X1 U50333 ( .A1(n18049), .A2(n39390), .Z(n39392) );
  XOR2_X1 U50334 ( .A1(n39393), .A2(n39392), .Z(n39394) );
  MUX2_X1 U50335 ( .I0(n39398), .I1(n39397), .S(n40091), .Z(n39413) );
  XOR2_X1 U50336 ( .A1(n39399), .A2(n39400), .Z(n50199) );
  XOR2_X1 U50337 ( .A1(n50199), .A2(n51915), .Z(n39401) );
  XOR2_X1 U50338 ( .A1(n22855), .A2(n39401), .Z(n39402) );
  XOR2_X1 U50339 ( .A1(n39403), .A2(n39402), .Z(n39404) );
  INV_X1 U50340 ( .I(n39894), .ZN(n39410) );
  NAND2_X1 U50341 ( .A1(n6576), .A2(n40069), .ZN(n39421) );
  INV_X1 U50342 ( .I(n40106), .ZN(n39423) );
  NOR2_X1 U50344 ( .A1(n40328), .A2(n64566), .ZN(n39424) );
  NAND2_X1 U50345 ( .A1(n40103), .A2(n19611), .ZN(n39425) );
  NAND2_X1 U50346 ( .A1(n40047), .A2(n4581), .ZN(n40054) );
  OAI21_X1 U50347 ( .A1(n23700), .A2(n7349), .B(n43117), .ZN(n39428) );
  NAND2_X1 U50348 ( .A1(n43111), .A2(n39429), .ZN(n39430) );
  XOR2_X1 U50349 ( .A1(n44876), .A2(n43789), .Z(n51949) );
  XOR2_X1 U50350 ( .A1(n53174), .A2(n39434), .Z(n50189) );
  XOR2_X1 U50351 ( .A1(n50189), .A2(n44412), .Z(n39435) );
  XOR2_X1 U50352 ( .A1(n51949), .A2(n39435), .Z(n39436) );
  XOR2_X1 U50353 ( .A1(n58252), .A2(n58972), .Z(n39441) );
  XOR2_X1 U50354 ( .A1(n39443), .A2(n39442), .Z(n50972) );
  XOR2_X1 U50355 ( .A1(n50969), .A2(n50025), .Z(n46413) );
  XOR2_X1 U50356 ( .A1(n39445), .A2(n39444), .Z(n50026) );
  XOR2_X1 U50357 ( .A1(n46413), .A2(n50026), .Z(n39446) );
  XOR2_X1 U50358 ( .A1(n50972), .A2(n39446), .Z(n39447) );
  XOR2_X1 U50359 ( .A1(n39451), .A2(n39450), .Z(n39452) );
  XOR2_X1 U50360 ( .A1(n39455), .A2(n39454), .Z(n39463) );
  INV_X1 U50361 ( .I(n50618), .ZN(n39456) );
  XOR2_X1 U50362 ( .A1(n39456), .A2(n54936), .Z(n50070) );
  XOR2_X1 U50363 ( .A1(n39458), .A2(n39457), .Z(n50960) );
  XOR2_X1 U50364 ( .A1(n50070), .A2(n50960), .Z(n39459) );
  XOR2_X1 U50365 ( .A1(n39460), .A2(n39459), .Z(n39461) );
  XOR2_X1 U50366 ( .A1(n39461), .A2(n39690), .Z(n39462) );
  XOR2_X1 U50367 ( .A1(n39463), .A2(n39462), .Z(n39464) );
  XOR2_X1 U50368 ( .A1(n22953), .A2(n39466), .Z(n39467) );
  XOR2_X1 U50369 ( .A1(n22961), .A2(n39469), .Z(n51487) );
  XOR2_X1 U50370 ( .A1(n51487), .A2(n50624), .Z(n39471) );
  INV_X1 U50371 ( .I(n27640), .ZN(n51686) );
  XOR2_X1 U50372 ( .A1(n46601), .A2(n51686), .Z(n43799) );
  XOR2_X1 U50373 ( .A1(n43799), .A2(n39613), .Z(n39470) );
  XOR2_X1 U50374 ( .A1(n39472), .A2(n22344), .Z(n39473) );
  XOR2_X1 U50376 ( .A1(n39478), .A2(n46615), .Z(n52319) );
  XOR2_X1 U50377 ( .A1(n50578), .A2(n52319), .Z(n39479) );
  OAI21_X1 U50379 ( .A1(n23046), .A2(n40568), .B(n41109), .ZN(n39487) );
  INV_X1 U50380 ( .I(n52366), .ZN(n39489) );
  XOR2_X1 U50381 ( .A1(n39488), .A2(n54231), .Z(n50571) );
  XOR2_X1 U50382 ( .A1(n39489), .A2(n50571), .Z(n39490) );
  XOR2_X1 U50383 ( .A1(n39493), .A2(n39492), .Z(n39496) );
  INV_X1 U50384 ( .I(n39494), .ZN(n39495) );
  NAND2_X1 U50387 ( .A1(n5241), .A2(n39957), .ZN(n39504) );
  NAND4_X1 U50388 ( .A1(n60091), .A2(n39512), .A3(n61233), .A4(n39511), .ZN(
        n39513) );
  INV_X1 U50389 ( .I(n39516), .ZN(n39520) );
  NAND2_X1 U50391 ( .A1(n39523), .A2(n16112), .ZN(n39526) );
  AOI21_X1 U50392 ( .A1(n39526), .A2(n39525), .B(n39524), .ZN(n39527) );
  INV_X1 U50393 ( .I(n45330), .ZN(n39529) );
  XOR2_X1 U50394 ( .A1(n39529), .A2(n54676), .Z(n51294) );
  XOR2_X1 U50395 ( .A1(n39530), .A2(n56143), .Z(n39531) );
  XOR2_X1 U50396 ( .A1(n51290), .A2(n39531), .Z(n51733) );
  XOR2_X1 U50397 ( .A1(n51733), .A2(n55840), .Z(n39532) );
  XOR2_X1 U50398 ( .A1(n51294), .A2(n39532), .Z(n39533) );
  XOR2_X1 U50399 ( .A1(n39625), .A2(n39533), .Z(n39535) );
  INV_X1 U50400 ( .I(n39536), .ZN(n39537) );
  XOR2_X1 U50401 ( .A1(n39537), .A2(n39611), .Z(n51238) );
  XOR2_X1 U50402 ( .A1(n39538), .A2(n52018), .Z(n39539) );
  XOR2_X1 U50403 ( .A1(n39540), .A2(n51045), .Z(n39541) );
  XOR2_X1 U50404 ( .A1(n51238), .A2(n39541), .Z(n39542) );
  XOR2_X1 U50405 ( .A1(n23655), .A2(n39542), .Z(n39545) );
  XOR2_X1 U50406 ( .A1(n39549), .A2(n55889), .Z(n52071) );
  XOR2_X1 U50407 ( .A1(n52071), .A2(n52178), .Z(n39550) );
  XOR2_X1 U50408 ( .A1(n23115), .A2(n39550), .Z(n39552) );
  XOR2_X1 U50409 ( .A1(n39556), .A2(n15707), .Z(n39557) );
  XOR2_X1 U50410 ( .A1(n39558), .A2(n39557), .Z(n49232) );
  XOR2_X1 U50411 ( .A1(n49232), .A2(n56849), .Z(n39559) );
  XOR2_X1 U50413 ( .A1(n15711), .A2(n23181), .Z(n39576) );
  XOR2_X1 U50414 ( .A1(n39568), .A2(n39567), .Z(n51724) );
  XOR2_X1 U50415 ( .A1(n53262), .A2(n56771), .Z(n39569) );
  XOR2_X1 U50416 ( .A1(n39569), .A2(n50831), .Z(n39571) );
  XOR2_X1 U50417 ( .A1(n39571), .A2(n39570), .Z(n51305) );
  INV_X1 U50418 ( .I(n30908), .ZN(n39572) );
  XOR2_X1 U50419 ( .A1(n51305), .A2(n39572), .Z(n39573) );
  XOR2_X1 U50420 ( .A1(n51724), .A2(n39573), .Z(n39574) );
  XOR2_X1 U50421 ( .A1(n17583), .A2(n39574), .Z(n39575) );
  XOR2_X1 U50422 ( .A1(n39576), .A2(n39575), .Z(n39577) );
  XOR2_X1 U50423 ( .A1(n25914), .A2(n39577), .Z(n39584) );
  XOR2_X1 U50424 ( .A1(n58235), .A2(n15729), .Z(n39581) );
  XOR2_X1 U50426 ( .A1(n39585), .A2(n39586), .Z(n39587) );
  XOR2_X1 U50427 ( .A1(n51992), .A2(n49289), .Z(n39591) );
  XOR2_X1 U50428 ( .A1(n23573), .A2(n39591), .Z(n39593) );
  XOR2_X1 U50429 ( .A1(n39692), .A2(n39593), .Z(n39594) );
  XOR2_X1 U50430 ( .A1(n39595), .A2(n39594), .Z(n39596) );
  XOR2_X1 U50431 ( .A1(n39597), .A2(n39596), .Z(n39600) );
  XOR2_X1 U50432 ( .A1(n23962), .A2(n39598), .Z(n39599) );
  NAND2_X2 U50433 ( .A1(n41430), .A2(n24302), .ZN(n41432) );
  NAND2_X1 U50434 ( .A1(n15439), .A2(n22832), .ZN(n39606) );
  NAND2_X1 U50435 ( .A1(n22638), .A2(n41433), .ZN(n39605) );
  NAND3_X1 U50436 ( .A1(n39606), .A2(n64773), .A3(n39605), .ZN(n39607) );
  AOI21_X1 U50437 ( .A1(n39609), .A2(n39608), .B(n39607), .ZN(n39610) );
  XOR2_X1 U50438 ( .A1(n39611), .A2(n53499), .Z(n39612) );
  XOR2_X1 U50439 ( .A1(n39613), .A2(n39612), .Z(n39615) );
  XOR2_X1 U50440 ( .A1(n24051), .A2(n23886), .Z(n39614) );
  XOR2_X1 U50441 ( .A1(n39723), .A2(n39614), .Z(n51046) );
  XOR2_X1 U50442 ( .A1(n39615), .A2(n51046), .Z(n39616) );
  XOR2_X1 U50443 ( .A1(n51680), .A2(n39616), .Z(n39617) );
  XOR2_X1 U50444 ( .A1(n39618), .A2(n39617), .Z(n39619) );
  XOR2_X1 U50446 ( .A1(n39622), .A2(n55335), .Z(n52606) );
  XOR2_X1 U50447 ( .A1(n39623), .A2(n54676), .Z(n51382) );
  XOR2_X1 U50448 ( .A1(n52606), .A2(n51382), .Z(n39624) );
  XOR2_X1 U50449 ( .A1(n39631), .A2(n52317), .Z(n39632) );
  XOR2_X1 U50450 ( .A1(n39633), .A2(n39632), .Z(n50389) );
  XOR2_X1 U50451 ( .A1(n55052), .A2(n60797), .Z(n39634) );
  XOR2_X1 U50452 ( .A1(n61238), .A2(n39634), .Z(n50934) );
  XOR2_X1 U50453 ( .A1(n50389), .A2(n50934), .Z(n39636) );
  XOR2_X1 U50454 ( .A1(n39639), .A2(n39640), .Z(n39759) );
  XOR2_X1 U50455 ( .A1(n9398), .A2(n23330), .Z(n39645) );
  NAND2_X1 U50456 ( .A1(n25760), .A2(n473), .ZN(n39648) );
  XOR2_X1 U50458 ( .A1(n39649), .A2(n9722), .Z(n50652) );
  XOR2_X1 U50459 ( .A1(n39650), .A2(n53989), .Z(n52180) );
  XOR2_X1 U50460 ( .A1(n52180), .A2(n50646), .Z(n39651) );
  XOR2_X1 U50461 ( .A1(n50652), .A2(n39651), .Z(n39652) );
  XOR2_X1 U50463 ( .A1(n39656), .A2(n39655), .Z(n39657) );
  INV_X1 U50464 ( .I(n39663), .ZN(n39664) );
  XOR2_X1 U50465 ( .A1(n39665), .A2(n39664), .Z(n51370) );
  XOR2_X1 U50466 ( .A1(n39667), .A2(n39666), .Z(n39668) );
  XOR2_X1 U50467 ( .A1(n39668), .A2(n50955), .Z(n52624) );
  XOR2_X1 U50468 ( .A1(n51370), .A2(n52624), .Z(n39669) );
  XOR2_X1 U50469 ( .A1(n22480), .A2(n39669), .Z(n39671) );
  XOR2_X1 U50470 ( .A1(n39673), .A2(n39672), .Z(n39674) );
  XOR2_X1 U50471 ( .A1(n39675), .A2(n39674), .Z(n39676) );
  XOR2_X1 U50473 ( .A1(n39680), .A2(n39681), .Z(n39695) );
  INV_X1 U50474 ( .I(n39682), .ZN(n39683) );
  XOR2_X1 U50475 ( .A1(n39684), .A2(n39683), .Z(n50926) );
  XOR2_X1 U50477 ( .A1(n39690), .A2(n22485), .Z(n39691) );
  INV_X1 U50479 ( .I(n40004), .ZN(n39700) );
  INV_X1 U50480 ( .I(n41126), .ZN(n40003) );
  XOR2_X1 U50482 ( .A1(n39705), .A2(n39704), .Z(n52438) );
  XOR2_X1 U50483 ( .A1(n39707), .A2(n39706), .Z(n50495) );
  XOR2_X1 U50484 ( .A1(n52438), .A2(n50495), .Z(n39708) );
  XOR2_X1 U50485 ( .A1(n21348), .A2(n39708), .Z(n39711) );
  XOR2_X1 U50486 ( .A1(n39711), .A2(n39710), .Z(n39712) );
  XOR2_X1 U50489 ( .A1(n39724), .A2(n39723), .Z(n51339) );
  XOR2_X1 U50490 ( .A1(n51339), .A2(n39725), .Z(n39726) );
  XOR2_X1 U50491 ( .A1(n44758), .A2(n39726), .Z(n39727) );
  XOR2_X1 U50492 ( .A1(n23898), .A2(n39727), .Z(n39729) );
  XOR2_X1 U50493 ( .A1(n59788), .A2(n39733), .Z(n39734) );
  XOR2_X1 U50494 ( .A1(n39735), .A2(n39734), .Z(n39747) );
  XOR2_X1 U50495 ( .A1(n39738), .A2(n23968), .Z(n49735) );
  XOR2_X1 U50496 ( .A1(n50864), .A2(n39739), .Z(n39740) );
  XOR2_X1 U50497 ( .A1(n49735), .A2(n39740), .Z(n39741) );
  XOR2_X1 U50498 ( .A1(n39741), .A2(n43497), .Z(n39742) );
  XOR2_X1 U50499 ( .A1(n39743), .A2(n39742), .Z(n39744) );
  XOR2_X1 U50500 ( .A1(n39745), .A2(n39744), .Z(n39746) );
  XOR2_X1 U50502 ( .A1(n43858), .A2(n9871), .Z(n39751) );
  XOR2_X1 U50503 ( .A1(n39752), .A2(n39751), .Z(n49122) );
  XOR2_X1 U50505 ( .A1(n39760), .A2(n22821), .Z(n49821) );
  INV_X1 U50506 ( .I(n50855), .ZN(n39762) );
  XOR2_X1 U50507 ( .A1(n39762), .A2(n39761), .Z(n39763) );
  XOR2_X1 U50508 ( .A1(n49821), .A2(n39763), .Z(n39764) );
  INV_X1 U50509 ( .I(n39770), .ZN(n39772) );
  XOR2_X1 U50510 ( .A1(n39772), .A2(n39771), .Z(n50527) );
  XOR2_X1 U50511 ( .A1(n39773), .A2(n53805), .Z(n52401) );
  XOR2_X1 U50512 ( .A1(n52401), .A2(n51379), .Z(n39774) );
  XOR2_X1 U50513 ( .A1(n50527), .A2(n39774), .Z(n39775) );
  NAND4_X1 U50516 ( .A1(n39782), .A2(n40857), .A3(n41073), .A4(n984), .ZN(
        n39785) );
  NAND2_X1 U50518 ( .A1(n41083), .A2(n39783), .ZN(n39784) );
  INV_X1 U50519 ( .I(n40390), .ZN(n39788) );
  NAND2_X1 U50520 ( .A1(n984), .A2(n40591), .ZN(n39787) );
  AOI21_X1 U50521 ( .A1(n40849), .A2(n39788), .B(n39787), .ZN(n39789) );
  NOR2_X1 U50523 ( .A1(n39792), .A2(n39791), .ZN(n39794) );
  NOR2_X1 U50527 ( .A1(n41325), .A2(n39798), .ZN(n39799) );
  INV_X1 U50528 ( .I(n43129), .ZN(n39801) );
  NOR2_X1 U50529 ( .A1(n22606), .A2(n43130), .ZN(n39800) );
  INV_X1 U50530 ( .I(n40747), .ZN(n39803) );
  OAI21_X1 U50531 ( .A1(n39803), .A2(n39810), .B(n40412), .ZN(n39805) );
  NAND2_X1 U50532 ( .A1(n40413), .A2(n59961), .ZN(n39804) );
  INV_X1 U50535 ( .I(n41466), .ZN(n39808) );
  INV_X1 U50536 ( .I(n41473), .ZN(n39811) );
  AOI21_X1 U50537 ( .A1(n39811), .A2(n41470), .B(n39810), .ZN(n39813) );
  OAI21_X1 U50538 ( .A1(n40755), .A2(n25131), .B(n41473), .ZN(n39812) );
  NAND2_X1 U50539 ( .A1(n39994), .A2(n41384), .ZN(n40421) );
  INV_X1 U50540 ( .I(n41127), .ZN(n39827) );
  NAND2_X1 U50543 ( .A1(n1748), .A2(n40568), .ZN(n39832) );
  OAI22_X1 U50544 ( .A1(n40571), .A2(n41106), .B1(n40443), .B2(n39832), .ZN(
        n39833) );
  AOI21_X1 U50545 ( .A1(n40568), .A2(n41101), .B(n39833), .ZN(n39839) );
  NAND2_X1 U50546 ( .A1(n39834), .A2(n40441), .ZN(n39837) );
  INV_X1 U50547 ( .I(n41449), .ZN(n39843) );
  OAI22_X1 U50548 ( .A1(n39848), .A2(n23406), .B1(n40380), .B2(n40702), .ZN(
        n39849) );
  NOR3_X1 U50549 ( .A1(n1303), .A2(n39852), .A3(n40737), .ZN(n39854) );
  NOR3_X1 U50550 ( .A1(n23108), .A2(n17063), .A3(n41397), .ZN(n39853) );
  NOR2_X1 U50551 ( .A1(n41402), .A2(n17063), .ZN(n39857) );
  INV_X1 U50552 ( .I(n42013), .ZN(n39877) );
  INV_X1 U50553 ( .I(n39862), .ZN(n39866) );
  INV_X1 U50554 ( .I(n39863), .ZN(n41209) );
  NAND2_X1 U50555 ( .A1(n41209), .A2(n997), .ZN(n39865) );
  NAND2_X1 U50556 ( .A1(n41223), .A2(n9935), .ZN(n39864) );
  INV_X1 U50557 ( .I(n41425), .ZN(n39867) );
  NAND2_X1 U50558 ( .A1(n40405), .A2(n39868), .ZN(n39874) );
  INV_X1 U50559 ( .I(n39869), .ZN(n39873) );
  NAND2_X1 U50560 ( .A1(n38935), .A2(n41415), .ZN(n39871) );
  NAND3_X1 U50561 ( .A1(n39871), .A2(n61316), .A3(n39870), .ZN(n39872) );
  NOR4_X1 U50562 ( .A1(n39877), .A2(n39876), .A3(n60472), .A4(n59381), .ZN(
        n39879) );
  OAI21_X1 U50563 ( .A1(n42014), .A2(n59381), .B(n43100), .ZN(n39881) );
  NOR2_X1 U50566 ( .A1(n19102), .A2(n42488), .ZN(n40093) );
  NAND3_X1 U50567 ( .A1(n40320), .A2(n60422), .A3(n61264), .ZN(n39891) );
  INV_X1 U50569 ( .I(n40349), .ZN(n39900) );
  NAND2_X1 U50571 ( .A1(n41810), .A2(n10593), .ZN(n39903) );
  OAI21_X1 U50572 ( .A1(n22759), .A2(n9808), .B(n753), .ZN(n39906) );
  NAND2_X1 U50573 ( .A1(n39906), .A2(n41308), .ZN(n39908) );
  NAND2_X1 U50574 ( .A1(n41307), .A2(n42453), .ZN(n39907) );
  MUX2_X1 U50575 ( .I0(n39908), .I1(n39907), .S(n63795), .Z(n39909) );
  NAND3_X1 U50576 ( .A1(n40135), .A2(n58970), .A3(n40296), .ZN(n39911) );
  NOR2_X1 U50577 ( .A1(n23904), .A2(n14018), .ZN(n40300) );
  OAI21_X1 U50578 ( .A1(n40295), .A2(n14014), .B(n23855), .ZN(n39912) );
  OAI21_X1 U50581 ( .A1(n64613), .A2(n4364), .B(n40296), .ZN(n39914) );
  INV_X1 U50583 ( .I(n40312), .ZN(n39921) );
  NAND2_X1 U50584 ( .A1(n42439), .A2(n39921), .ZN(n39923) );
  NAND3_X1 U50586 ( .A1(n41816), .A2(n41820), .A3(n21207), .ZN(n39930) );
  NAND2_X1 U50587 ( .A1(n13169), .A2(n20277), .ZN(n41272) );
  AOI21_X1 U50588 ( .A1(n41276), .A2(n41272), .B(n41280), .ZN(n39932) );
  NOR2_X1 U50590 ( .A1(n19487), .A2(n41350), .ZN(n39940) );
  NAND2_X1 U50591 ( .A1(n43206), .A2(n41347), .ZN(n39939) );
  OAI21_X1 U50592 ( .A1(n24002), .A2(n43058), .B(n22673), .ZN(n39941) );
  OAI21_X1 U50594 ( .A1(n7237), .A2(n62123), .B(n39949), .ZN(n39951) );
  NOR2_X1 U50595 ( .A1(n41428), .A2(n41439), .ZN(n39954) );
  INV_X1 U50596 ( .I(n40703), .ZN(n39955) );
  NAND2_X1 U50601 ( .A1(n40858), .A2(n39973), .ZN(n39964) );
  NAND4_X1 U50602 ( .A1(n39967), .A2(n39966), .A3(n39965), .A4(n39964), .ZN(
        n39980) );
  NAND2_X1 U50606 ( .A1(n39971), .A2(n40393), .ZN(n39978) );
  INV_X1 U50607 ( .I(n40593), .ZN(n39975) );
  NAND2_X1 U50608 ( .A1(n984), .A2(n40854), .ZN(n39974) );
  NAND3_X1 U50609 ( .A1(n41072), .A2(n39975), .A3(n39974), .ZN(n39976) );
  NAND3_X1 U50610 ( .A1(n39978), .A2(n39977), .A3(n39976), .ZN(n39979) );
  OAI21_X1 U50615 ( .A1(n40759), .A2(n25131), .B(n39986), .ZN(n39990) );
  NAND2_X1 U50622 ( .A1(n39999), .A2(n41122), .ZN(n40001) );
  NAND4_X1 U50623 ( .A1(n40002), .A2(n40001), .A3(n10294), .A4(n40000), .ZN(
        n40009) );
  NAND2_X1 U50624 ( .A1(n40004), .A2(n40003), .ZN(n40008) );
  INV_X1 U50625 ( .I(n41124), .ZN(n40006) );
  NOR3_X1 U50626 ( .A1(n43434), .A2(n43444), .A3(n43437), .ZN(n40012) );
  INV_X1 U50628 ( .I(n42372), .ZN(n40018) );
  NOR2_X1 U50629 ( .A1(n40018), .A2(n62001), .ZN(n40019) );
  NOR3_X1 U50631 ( .A1(n41744), .A2(n41743), .A3(n43439), .ZN(n40022) );
  NOR2_X1 U50632 ( .A1(n42051), .A2(n42944), .ZN(n40021) );
  AOI21_X1 U50633 ( .A1(n57955), .A2(n40295), .B(n40224), .ZN(n40027) );
  NOR2_X1 U50634 ( .A1(n40034), .A2(n22943), .ZN(n40036) );
  MUX2_X1 U50635 ( .I0(n40036), .I1(n40035), .S(n9627), .Z(n40046) );
  NAND2_X1 U50636 ( .A1(n42468), .A2(n25666), .ZN(n40041) );
  NAND2_X1 U50637 ( .A1(n40350), .A2(n1515), .ZN(n40040) );
  NAND3_X1 U50638 ( .A1(n40041), .A2(n41844), .A3(n40040), .ZN(n40042) );
  NOR2_X1 U50639 ( .A1(n40056), .A2(n40337), .ZN(n40058) );
  INV_X1 U50640 ( .I(n42417), .ZN(n40085) );
  NAND2_X1 U50641 ( .A1(n65128), .A2(n14863), .ZN(n40060) );
  NAND2_X1 U50643 ( .A1(n63952), .A2(n1721), .ZN(n40067) );
  OR2_X1 U50647 ( .A1(n40081), .A2(n1193), .Z(n40084) );
  OAI21_X1 U50649 ( .A1(n60422), .A2(n60929), .B(n60971), .ZN(n40088) );
  NAND2_X1 U50650 ( .A1(n40094), .A2(n40093), .ZN(n40126) );
  NAND2_X1 U50651 ( .A1(n43464), .A2(n26020), .ZN(n43474) );
  OAI21_X1 U50652 ( .A1(n42966), .A2(n43457), .B(n1193), .ZN(n40098) );
  NAND4_X1 U50653 ( .A1(n40102), .A2(n40101), .A3(n57536), .A4(n12285), .ZN(
        n40105) );
  NAND3_X1 U50656 ( .A1(n40946), .A2(n58941), .A3(n40196), .ZN(n40114) );
  OAI21_X1 U50658 ( .A1(n23986), .A2(n40952), .B(n40116), .ZN(n40119) );
  AOI21_X1 U50659 ( .A1(n58941), .A2(n40200), .B(n10341), .ZN(n40118) );
  OAI22_X1 U50660 ( .A1(n40120), .A2(n40119), .B1(n40118), .B2(n40117), .ZN(
        n40121) );
  NAND3_X1 U50661 ( .A1(n40123), .A2(n23654), .A3(n60422), .ZN(n40124) );
  OAI21_X1 U50662 ( .A1(n40133), .A2(n40304), .B(n22746), .ZN(n40134) );
  NOR2_X1 U50663 ( .A1(n60153), .A2(n40296), .ZN(n40137) );
  OAI21_X1 U50664 ( .A1(n40299), .A2(n40137), .B(n40136), .ZN(n40138) );
  NOR2_X1 U50666 ( .A1(n40162), .A2(n64948), .ZN(n40159) );
  NAND2_X1 U50669 ( .A1(n40166), .A2(n40238), .ZN(n40170) );
  INV_X1 U50671 ( .I(n41977), .ZN(n40187) );
  NOR2_X1 U50673 ( .A1(n4805), .A2(n42383), .ZN(n40179) );
  NOR2_X1 U50675 ( .A1(n42697), .A2(n42703), .ZN(n40176) );
  AOI21_X1 U50676 ( .A1(n40176), .A2(n41972), .B(n40175), .ZN(n40177) );
  NAND3_X1 U50678 ( .A1(n42689), .A2(n41522), .A3(n42694), .ZN(n40183) );
  NOR2_X1 U50679 ( .A1(n41972), .A2(n5939), .ZN(n40181) );
  NOR3_X1 U50680 ( .A1(n42383), .A2(n9672), .A3(n42703), .ZN(n40180) );
  AOI21_X1 U50681 ( .A1(n40181), .A2(n42704), .B(n40180), .ZN(n40182) );
  OAI21_X1 U50683 ( .A1(n40200), .A2(n40199), .B(n40944), .ZN(n40201) );
  NAND2_X1 U50684 ( .A1(n40205), .A2(n40943), .ZN(n40206) );
  NOR2_X1 U50686 ( .A1(n23855), .A2(n14014), .ZN(n40219) );
  NOR2_X1 U50687 ( .A1(n6932), .A2(n40219), .ZN(n40222) );
  NAND2_X1 U50689 ( .A1(n40288), .A2(n40224), .ZN(n40225) );
  NOR2_X1 U50691 ( .A1(n40233), .A2(n40238), .ZN(n40234) );
  NOR2_X1 U50692 ( .A1(n40235), .A2(n40234), .ZN(n40247) );
  NAND3_X1 U50693 ( .A1(n40237), .A2(n40236), .A3(n11126), .ZN(n40245) );
  NOR2_X1 U50695 ( .A1(n40250), .A2(n60172), .ZN(n40254) );
  NAND2_X1 U50696 ( .A1(n4968), .A2(n40470), .ZN(n40253) );
  NAND2_X1 U50697 ( .A1(n40923), .A2(n7201), .ZN(n40473) );
  AOI21_X1 U50698 ( .A1(n40930), .A2(n40473), .B(n40465), .ZN(n40252) );
  NAND2_X1 U50699 ( .A1(n40930), .A2(n40924), .ZN(n40251) );
  NAND2_X1 U50702 ( .A1(n40923), .A2(n40257), .ZN(n40260) );
  NOR2_X1 U50706 ( .A1(n40263), .A2(n40470), .ZN(n40264) );
  INV_X1 U50707 ( .I(n40272), .ZN(n40273) );
  AOI21_X1 U50708 ( .A1(n22999), .A2(n40276), .B(n1694), .ZN(n40277) );
  NAND2_X1 U50709 ( .A1(n41980), .A2(n40893), .ZN(n40279) );
  INV_X1 U50711 ( .I(n42362), .ZN(n40281) );
  NAND3_X1 U50713 ( .A1(n64961), .A2(n9801), .A3(n42355), .ZN(n40284) );
  NAND2_X1 U50716 ( .A1(n64613), .A2(n4364), .ZN(n40298) );
  NOR2_X1 U50718 ( .A1(n42427), .A2(n57208), .ZN(n40313) );
  OAI22_X1 U50719 ( .A1(n40317), .A2(n40316), .B1(n60422), .B2(n42495), .ZN(
        n40318) );
  AOI21_X1 U50720 ( .A1(n61264), .A2(n40320), .B(n40319), .ZN(n40327) );
  NOR2_X1 U50721 ( .A1(n9980), .A2(n60971), .ZN(n40323) );
  AOI22_X1 U50722 ( .A1(n57327), .A2(n19102), .B1(n40323), .B2(n40322), .ZN(
        n40326) );
  OAI21_X1 U50723 ( .A1(n40324), .A2(n42486), .B(n64077), .ZN(n40325) );
  NAND3_X1 U50724 ( .A1(n40331), .A2(n40330), .A3(n40329), .ZN(n40332) );
  NAND2_X1 U50725 ( .A1(n40333), .A2(n40332), .ZN(n40345) );
  NAND2_X1 U50726 ( .A1(n22282), .A2(n4322), .ZN(n42652) );
  INV_X1 U50727 ( .I(n42652), .ZN(n40365) );
  NAND2_X1 U50728 ( .A1(n42479), .A2(n18473), .ZN(n40352) );
  INV_X1 U50729 ( .I(n58307), .ZN(n40353) );
  NAND2_X1 U50730 ( .A1(n753), .A2(n42451), .ZN(n40357) );
  NOR2_X1 U50732 ( .A1(n59674), .A2(n664), .ZN(n40359) );
  AOI21_X1 U50734 ( .A1(n40361), .A2(n64359), .B(n40360), .ZN(n40362) );
  AOI21_X1 U50735 ( .A1(n40366), .A2(n40365), .B(n43358), .ZN(n40373) );
  NAND2_X1 U50736 ( .A1(n22282), .A2(n21644), .ZN(n40369) );
  NAND4_X1 U50737 ( .A1(n42648), .A2(n42655), .A3(n40369), .A4(n40368), .ZN(
        n40370) );
  MUX2_X1 U50738 ( .I0(n357), .I1(n25976), .S(n41432), .Z(n40375) );
  NAND2_X1 U50739 ( .A1(n40375), .A2(n40374), .ZN(n40386) );
  NOR3_X1 U50740 ( .A1(n41432), .A2(n41428), .A3(n60653), .ZN(n40377) );
  OAI21_X1 U50743 ( .A1(n14132), .A2(n63914), .B(n40854), .ZN(n40388) );
  NAND2_X1 U50746 ( .A1(n41084), .A2(n41073), .ZN(n40396) );
  AOI21_X1 U50749 ( .A1(n9935), .A2(n10173), .B(n20652), .ZN(n40410) );
  AOI21_X1 U50750 ( .A1(n64826), .A2(n13049), .B(n59203), .ZN(n40409) );
  NAND2_X1 U50751 ( .A1(n40748), .A2(n7165), .ZN(n40411) );
  NAND2_X1 U50752 ( .A1(n40413), .A2(n41466), .ZN(n40415) );
  AOI22_X1 U50756 ( .A1(n40421), .A2(n41122), .B1(n10294), .B2(n61638), .ZN(
        n40423) );
  NAND2_X1 U50757 ( .A1(n61417), .A2(n41382), .ZN(n40422) );
  NAND3_X1 U50758 ( .A1(n40424), .A2(n40423), .A3(n40422), .ZN(n40430) );
  NAND3_X1 U50759 ( .A1(n57309), .A2(n41377), .A3(n40425), .ZN(n40429) );
  NAND2_X1 U50760 ( .A1(n1724), .A2(n41118), .ZN(n40428) );
  NAND4_X2 U50761 ( .A1(n40430), .A2(n40429), .A3(n40428), .A4(n40427), .ZN(
        n40448) );
  NOR2_X1 U50762 ( .A1(n40431), .A2(n57651), .ZN(n40447) );
  OAI21_X1 U50764 ( .A1(n40568), .A2(n25358), .B(n61710), .ZN(n40433) );
  AOI21_X1 U50769 ( .A1(n42759), .A2(n1691), .B(n42757), .ZN(n40449) );
  INV_X1 U50770 ( .I(n40449), .ZN(n40450) );
  NAND3_X1 U50772 ( .A1(n42754), .A2(n22182), .A3(n11198), .ZN(n40454) );
  XOR2_X1 U50773 ( .A1(n40458), .A2(n22773), .Z(n40461) );
  INV_X1 U50774 ( .I(n40459), .ZN(n40460) );
  XOR2_X1 U50775 ( .A1(n40461), .A2(n40460), .Z(n40462) );
  XOR2_X1 U50776 ( .A1(n22731), .A2(n40462), .Z(n40554) );
  INV_X1 U50781 ( .I(n40473), .ZN(n40474) );
  NOR2_X1 U50786 ( .A1(n40653), .A2(n23616), .ZN(n40492) );
  NAND3_X1 U50788 ( .A1(n40670), .A2(n40494), .A3(n40663), .ZN(n40495) );
  NAND2_X1 U50790 ( .A1(n40500), .A2(n60652), .ZN(n40501) );
  NOR2_X1 U50793 ( .A1(n22738), .A2(n37532), .ZN(n40508) );
  BUF_X4 U50795 ( .I(n40511), .Z(n42127) );
  NOR2_X1 U50796 ( .A1(n22617), .A2(n23319), .ZN(n40513) );
  NAND2_X1 U50797 ( .A1(n1747), .A2(n41034), .ZN(n40512) );
  NOR2_X1 U50798 ( .A1(n40958), .A2(n61333), .ZN(n40521) );
  OAI21_X1 U50799 ( .A1(n40522), .A2(n40521), .B(n23787), .ZN(n40536) );
  NAND2_X1 U50800 ( .A1(n40617), .A2(n40963), .ZN(n40524) );
  NOR2_X1 U50802 ( .A1(n40619), .A2(n40968), .ZN(n40529) );
  OAI21_X1 U50803 ( .A1(n40530), .A2(n40529), .B(n64571), .ZN(n40534) );
  OAI21_X1 U50804 ( .A1(n40967), .A2(n40532), .B(n40531), .ZN(n40533) );
  NAND2_X1 U50806 ( .A1(n42143), .A2(n10004), .ZN(n41555) );
  NAND2_X1 U50807 ( .A1(n42140), .A2(n42670), .ZN(n41335) );
  AOI21_X1 U50808 ( .A1(n41555), .A2(n41335), .B(n42666), .ZN(n40544) );
  NAND2_X1 U50811 ( .A1(n41785), .A2(n42849), .ZN(n40552) );
  NOR2_X1 U50812 ( .A1(n42670), .A2(n21376), .ZN(n40549) );
  INV_X1 U50813 ( .I(n40547), .ZN(n40548) );
  AOI21_X1 U50814 ( .A1(n40549), .A2(n40548), .B(n41562), .ZN(n42852) );
  NAND2_X1 U50815 ( .A1(n42667), .A2(n10004), .ZN(n40551) );
  AOI21_X1 U50816 ( .A1(n40552), .A2(n42852), .B(n42850), .ZN(n40553) );
  NAND2_X1 U50820 ( .A1(n24644), .A2(n25837), .ZN(n40575) );
  NAND2_X1 U50822 ( .A1(n41873), .A2(n40585), .ZN(n40586) );
  INV_X1 U50823 ( .I(n43335), .ZN(n40596) );
  NAND2_X1 U50824 ( .A1(n40597), .A2(n40596), .ZN(n40600) );
  INV_X1 U50825 ( .I(n42587), .ZN(n40598) );
  NAND4_X1 U50826 ( .A1(n40598), .A2(n43341), .A3(n43601), .A4(n41627), .ZN(
        n40599) );
  NOR2_X1 U50827 ( .A1(n38675), .A2(n60567), .ZN(n40625) );
  INV_X1 U50828 ( .I(n40720), .ZN(n40635) );
  NOR3_X1 U50829 ( .A1(n65021), .A2(n7012), .A3(n40641), .ZN(n40649) );
  NAND2_X1 U50830 ( .A1(n7012), .A2(n40650), .ZN(n40646) );
  OAI21_X1 U50831 ( .A1(n40646), .A2(n40645), .B(n23884), .ZN(n40647) );
  NOR2_X2 U50832 ( .A1(n23709), .A2(n22002), .ZN(n42892) );
  NAND2_X1 U50833 ( .A1(n40654), .A2(n40653), .ZN(n40655) );
  OAI22_X1 U50835 ( .A1(n41178), .A2(n23616), .B1(n10022), .B2(n9915), .ZN(
        n40665) );
  NOR2_X1 U50837 ( .A1(n41178), .A2(n41173), .ZN(n40669) );
  NOR2_X1 U50838 ( .A1(n40667), .A2(n23616), .ZN(n40668) );
  AOI22_X1 U50839 ( .A1(n40670), .A2(n40669), .B1(n41172), .B2(n40668), .ZN(
        n40671) );
  NAND3_X1 U50840 ( .A1(n64366), .A2(n41453), .A3(n40713), .ZN(n40675) );
  NOR2_X1 U50841 ( .A1(n41155), .A2(n20984), .ZN(n40678) );
  OAI21_X1 U50842 ( .A1(n4819), .A2(n20994), .B(n1516), .ZN(n40677) );
  NAND2_X1 U50846 ( .A1(n42054), .A2(n43155), .ZN(n40686) );
  NOR2_X1 U50847 ( .A1(n40686), .A2(n42572), .ZN(n40688) );
  XOR2_X1 U50849 ( .A1(n45145), .A2(n50494), .Z(n40785) );
  INV_X1 U50850 ( .I(n40691), .ZN(n40692) );
  NAND3_X1 U50851 ( .A1(n40692), .A2(n41437), .A3(n41445), .ZN(n40693) );
  NAND2_X1 U50852 ( .A1(n41444), .A2(n40695), .ZN(n40696) );
  INV_X1 U50853 ( .I(n40699), .ZN(n40700) );
  NAND2_X1 U50854 ( .A1(n40701), .A2(n40700), .ZN(n40704) );
  INV_X1 U50855 ( .I(n40707), .ZN(n40709) );
  NAND2_X1 U50862 ( .A1(n41232), .A2(n41236), .ZN(n40741) );
  AOI22_X1 U50864 ( .A1(n41231), .A2(n40745), .B1(n23780), .B2(n41411), .ZN(
        n40746) );
  NAND2_X1 U50865 ( .A1(n42038), .A2(n20888), .ZN(n40784) );
  NAND2_X1 U50868 ( .A1(n40766), .A2(n38935), .ZN(n40767) );
  NOR2_X1 U50869 ( .A1(n41419), .A2(n64364), .ZN(n41211) );
  INV_X1 U50870 ( .I(n41211), .ZN(n41216) );
  AOI21_X1 U50871 ( .A1(n40767), .A2(n41216), .B(n64826), .ZN(n40768) );
  NAND2_X1 U50872 ( .A1(n12806), .A2(n57615), .ZN(n40772) );
  OAI22_X1 U50873 ( .A1(n40772), .A2(n41414), .B1(n40771), .B2(n61316), .ZN(
        n40773) );
  INV_X1 U50874 ( .I(n40773), .ZN(n40774) );
  INV_X1 U50875 ( .I(n43511), .ZN(n40780) );
  OAI21_X1 U50876 ( .A1(n65262), .A2(n40777), .B(n43513), .ZN(n40778) );
  AOI22_X1 U50877 ( .A1(n40781), .A2(n40780), .B1(n40779), .B2(n40778), .ZN(
        n40783) );
  INV_X1 U50880 ( .I(n41097), .ZN(n40801) );
  NAND2_X1 U50881 ( .A1(n42263), .A2(n22502), .ZN(n40800) );
  NAND2_X1 U50882 ( .A1(n40802), .A2(n41894), .ZN(n40803) );
  NAND2_X1 U50883 ( .A1(n41906), .A2(n40805), .ZN(n40806) );
  AOI21_X1 U50887 ( .A1(n40814), .A2(n40813), .B(n22713), .ZN(n40815) );
  OAI21_X1 U50890 ( .A1(n13465), .A2(n40826), .B(n40825), .ZN(n40837) );
  INV_X1 U50893 ( .I(n40829), .ZN(n40830) );
  INV_X1 U50894 ( .I(n40833), .ZN(n40834) );
  NAND2_X1 U50895 ( .A1(n40834), .A2(n7237), .ZN(n40835) );
  NOR2_X1 U50896 ( .A1(n60006), .A2(n62461), .ZN(n40867) );
  NOR2_X1 U50899 ( .A1(n41072), .A2(n9790), .ZN(n40856) );
  NAND2_X1 U50901 ( .A1(n41883), .A2(n40862), .ZN(n41639) );
  NAND2_X1 U50902 ( .A1(n61008), .A2(n25817), .ZN(n40863) );
  NAND3_X1 U50903 ( .A1(n41642), .A2(n40864), .A3(n40863), .ZN(n40865) );
  NOR3_X1 U50904 ( .A1(n41641), .A2(n41639), .A3(n40865), .ZN(n40866) );
  NAND2_X1 U50905 ( .A1(n58210), .A2(n42118), .ZN(n40869) );
  OAI22_X1 U50906 ( .A1(n40869), .A2(n43212), .B1(n41637), .B2(n40868), .ZN(
        n40870) );
  AOI21_X1 U50907 ( .A1(n57788), .A2(n12073), .B(n58343), .ZN(n40873) );
  AOI21_X1 U50908 ( .A1(n41692), .A2(n40873), .B(n42401), .ZN(n40875) );
  NAND2_X1 U50909 ( .A1(n25534), .A2(n42399), .ZN(n40874) );
  OAI21_X1 U50910 ( .A1(n42607), .A2(n57454), .B(n64629), .ZN(n40876) );
  NOR2_X1 U50911 ( .A1(n8799), .A2(n9200), .ZN(n40878) );
  NOR2_X1 U50912 ( .A1(n429), .A2(n59771), .ZN(n40877) );
  NAND2_X1 U50913 ( .A1(n41797), .A2(n60657), .ZN(n40879) );
  INV_X1 U50914 ( .I(n40885), .ZN(n40889) );
  INV_X1 U50916 ( .I(n40896), .ZN(n40898) );
  INV_X1 U50917 ( .I(n43016), .ZN(n40905) );
  INV_X1 U50918 ( .I(n42329), .ZN(n40904) );
  NAND3_X1 U50920 ( .A1(n42319), .A2(n5261), .A3(n41996), .ZN(n40906) );
  NAND3_X1 U50922 ( .A1(n42314), .A2(n41684), .A3(n42324), .ZN(n40910) );
  OAI21_X1 U50923 ( .A1(n40908), .A2(n43015), .B(n41682), .ZN(n40909) );
  AOI21_X1 U50924 ( .A1(n43024), .A2(n43027), .B(n43028), .ZN(n40913) );
  NOR2_X1 U50925 ( .A1(n41666), .A2(n42180), .ZN(n40916) );
  NAND2_X1 U50926 ( .A1(n41670), .A2(n61344), .ZN(n40915) );
  OAI21_X1 U50927 ( .A1(n40916), .A2(n40915), .B(n40914), .ZN(n40917) );
  XOR2_X1 U50928 ( .A1(n40918), .A2(n44631), .Z(n51587) );
  XOR2_X1 U50929 ( .A1(n40919), .A2(n51881), .Z(n40920) );
  XOR2_X1 U50930 ( .A1(n51587), .A2(n40920), .Z(n40921) );
  XOR2_X1 U50931 ( .A1(n22376), .A2(n40921), .Z(n40922) );
  NAND2_X1 U50934 ( .A1(n40939), .A2(n22809), .ZN(n40931) );
  NAND3_X1 U50935 ( .A1(n40933), .A2(n65206), .A3(n40932), .ZN(n41516) );
  INV_X1 U50937 ( .I(n40936), .ZN(n40937) );
  NOR2_X1 U50938 ( .A1(n40942), .A2(n40941), .ZN(n41510) );
  AOI22_X1 U50939 ( .A1(n18612), .A2(n15558), .B1(n58941), .B2(n40952), .ZN(
        n40955) );
  NOR2_X1 U50941 ( .A1(n38607), .A2(n40968), .ZN(n40966) );
  NAND2_X1 U50942 ( .A1(n61333), .A2(n23787), .ZN(n40969) );
  INV_X1 U50943 ( .I(n40969), .ZN(n40965) );
  AOI22_X1 U50944 ( .A1(n40967), .A2(n40966), .B1(n40965), .B2(n40964), .ZN(
        n40977) );
  AOI21_X1 U50945 ( .A1(n40969), .A2(n18704), .B(n40968), .ZN(n40973) );
  NAND2_X1 U50946 ( .A1(n61000), .A2(n23833), .ZN(n40982) );
  NAND2_X1 U50949 ( .A1(n40996), .A2(n23833), .ZN(n40985) );
  INV_X1 U50950 ( .I(n40990), .ZN(n40992) );
  NOR2_X1 U50951 ( .A1(n63721), .A2(n295), .ZN(n41045) );
  NOR2_X1 U50955 ( .A1(n41020), .A2(n12523), .ZN(n41021) );
  OAI21_X1 U50956 ( .A1(n14306), .A2(n23355), .B(n1275), .ZN(n41023) );
  NAND2_X1 U50957 ( .A1(n41023), .A2(n1728), .ZN(n41024) );
  NAND2_X1 U50958 ( .A1(n41030), .A2(n41034), .ZN(n41028) );
  AOI21_X1 U50959 ( .A1(n41029), .A2(n41028), .B(n41027), .ZN(n41033) );
  NOR2_X1 U50960 ( .A1(n41035), .A2(n21736), .ZN(n41036) );
  INV_X1 U50961 ( .I(n42870), .ZN(n41044) );
  OAI21_X1 U50962 ( .A1(n60952), .A2(n42866), .B(n42171), .ZN(n43819) );
  INV_X1 U50964 ( .I(n43816), .ZN(n41047) );
  NAND2_X1 U50965 ( .A1(n43817), .A2(n41048), .ZN(n41049) );
  AOI21_X1 U50966 ( .A1(n41885), .A2(n41876), .B(n41877), .ZN(n41055) );
  NOR2_X1 U50967 ( .A1(n20598), .A2(n64592), .ZN(n41058) );
  OAI22_X1 U50968 ( .A1(n41066), .A2(n64592), .B1(n41065), .B2(n41064), .ZN(
        n41067) );
  NOR2_X1 U50970 ( .A1(n41083), .A2(n9790), .ZN(n41086) );
  NAND2_X1 U50973 ( .A1(n41109), .A2(n59591), .ZN(n41110) );
  NAND2_X1 U50976 ( .A1(n60091), .A2(n23420), .ZN(n41133) );
  NOR2_X1 U50977 ( .A1(n25328), .A2(n43572), .ZN(n41138) );
  INV_X1 U50978 ( .I(n6967), .ZN(n45052) );
  AOI21_X1 U50980 ( .A1(n41453), .A2(n41148), .B(n59871), .ZN(n41150) );
  NAND3_X1 U50981 ( .A1(n64366), .A2(n58996), .A3(n1516), .ZN(n41154) );
  NAND2_X1 U50983 ( .A1(n41462), .A2(n1516), .ZN(n41452) );
  NOR2_X1 U50984 ( .A1(n41452), .A2(n41155), .ZN(n41156) );
  NAND3_X1 U50985 ( .A1(n41159), .A2(n7012), .A3(n22380), .ZN(n41170) );
  AOI22_X1 U50986 ( .A1(n41166), .A2(n14462), .B1(n64277), .B2(n7011), .ZN(
        n41169) );
  NAND2_X1 U50987 ( .A1(n41177), .A2(n41183), .ZN(n41179) );
  NAND2_X1 U50988 ( .A1(n41183), .A2(n15723), .ZN(n41184) );
  NAND3_X1 U50991 ( .A1(n12805), .A2(n41209), .A3(n41420), .ZN(n41228) );
  INV_X1 U50994 ( .I(n12806), .ZN(n41224) );
  INV_X1 U50997 ( .I(n16103), .ZN(n41244) );
  NAND3_X1 U50999 ( .A1(n1303), .A2(n41234), .A3(n61013), .ZN(n41238) );
  NAND2_X1 U51001 ( .A1(n41249), .A2(n42287), .ZN(n41253) );
  NAND3_X2 U51002 ( .A1(n41253), .A2(n41252), .A3(n41251), .ZN(n41254) );
  NAND2_X1 U51005 ( .A1(n42249), .A2(n60826), .ZN(n41267) );
  NAND2_X1 U51006 ( .A1(n43889), .A2(n7516), .ZN(n41314) );
  NOR2_X1 U51007 ( .A1(n41858), .A2(n41270), .ZN(n42300) );
  NOR2_X1 U51008 ( .A1(n41280), .A2(n23744), .ZN(n41277) );
  NOR2_X1 U51009 ( .A1(n42509), .A2(n41270), .ZN(n41271) );
  OAI21_X1 U51010 ( .A1(n41277), .A2(n41271), .B(n42503), .ZN(n41275) );
  AOI22_X1 U51011 ( .A1(n41275), .A2(n41274), .B1(n41273), .B2(n1403), .ZN(
        n41286) );
  INV_X1 U51012 ( .I(n41277), .ZN(n41278) );
  NAND3_X1 U51013 ( .A1(n41279), .A2(n9954), .A3(n23744), .ZN(n41282) );
  NAND3_X1 U51014 ( .A1(n42498), .A2(n41280), .A3(n9954), .ZN(n41281) );
  INV_X1 U51017 ( .I(n42211), .ZN(n42520) );
  OAI21_X1 U51018 ( .A1(n41288), .A2(n63233), .B(n42520), .ZN(n41292) );
  NAND2_X1 U51019 ( .A1(n41832), .A2(n60947), .ZN(n41290) );
  NAND3_X1 U51020 ( .A1(n41292), .A2(n41291), .A3(n41290), .ZN(n41299) );
  NAND2_X1 U51021 ( .A1(n41867), .A2(n23501), .ZN(n41297) );
  NAND3_X1 U51024 ( .A1(n41303), .A2(n41954), .A3(n42237), .ZN(n41305) );
  INV_X1 U51025 ( .I(n41310), .ZN(n41311) );
  MUX2_X1 U51026 ( .I0(n41314), .I1(n43142), .S(n20685), .Z(n41319) );
  NOR2_X1 U51028 ( .A1(n43140), .A2(n61951), .ZN(n41316) );
  NOR2_X2 U51029 ( .A1(n43890), .A2(n43241), .ZN(n43655) );
  NAND2_X1 U51032 ( .A1(n41322), .A2(n2330), .ZN(n41323) );
  INV_X1 U51034 ( .I(n43272), .ZN(n41326) );
  OAI21_X1 U51035 ( .A1(n41791), .A2(n41326), .B(n43131), .ZN(n41327) );
  NOR2_X1 U51036 ( .A1(n42377), .A2(n42383), .ZN(n41328) );
  NAND2_X1 U51038 ( .A1(n41532), .A2(n41969), .ZN(n41331) );
  XOR2_X1 U51039 ( .A1(n24278), .A2(n45261), .Z(n41333) );
  OAI21_X1 U51040 ( .A1(n42140), .A2(n41334), .B(n42660), .ZN(n41338) );
  AOI21_X1 U51041 ( .A1(n41335), .A2(n9914), .B(n64105), .ZN(n41337) );
  OAI21_X1 U51042 ( .A1(n42660), .A2(n64105), .B(n64532), .ZN(n41336) );
  OAI21_X1 U51043 ( .A1(n41338), .A2(n41337), .B(n41336), .ZN(n41346) );
  NOR2_X1 U51045 ( .A1(n41562), .A2(n41560), .ZN(n41343) );
  NAND2_X1 U51047 ( .A1(n43202), .A2(n24002), .ZN(n41349) );
  INV_X1 U51048 ( .I(n41354), .ZN(n41356) );
  NOR2_X1 U51049 ( .A1(n24981), .A2(n43225), .ZN(n41355) );
  OAI21_X1 U51050 ( .A1(n43220), .A2(n41356), .B(n41355), .ZN(n41357) );
  NOR2_X1 U51051 ( .A1(n42674), .A2(n41369), .ZN(n41361) );
  NAND2_X1 U51053 ( .A1(n6705), .A2(n42827), .ZN(n41362) );
  NAND2_X1 U51054 ( .A1(n17467), .A2(n42835), .ZN(n41368) );
  NOR2_X1 U51055 ( .A1(n42824), .A2(n42672), .ZN(n41370) );
  NAND2_X1 U51056 ( .A1(n41392), .A2(n473), .ZN(n41390) );
  NAND2_X1 U51057 ( .A1(n10294), .A2(n41385), .ZN(n41387) );
  AOI21_X1 U51058 ( .A1(n41388), .A2(n41387), .B(n10074), .ZN(n41389) );
  INV_X1 U51059 ( .I(n41392), .ZN(n41393) );
  NOR2_X1 U51060 ( .A1(n41394), .A2(n41393), .ZN(n41395) );
  INV_X1 U51062 ( .I(n41399), .ZN(n41404) );
  OAI21_X1 U51066 ( .A1(n23108), .A2(n41411), .B(n41410), .ZN(n41413) );
  INV_X1 U51069 ( .I(n41424), .ZN(n41426) );
  NAND2_X1 U51070 ( .A1(n277), .A2(n357), .ZN(n41431) );
  AOI21_X1 U51071 ( .A1(n41432), .A2(n41431), .B(n15441), .ZN(n41434) );
  INV_X1 U51072 ( .I(n43320), .ZN(n41465) );
  NOR2_X1 U51073 ( .A1(n41454), .A2(n41453), .ZN(n41456) );
  AOI21_X1 U51074 ( .A1(n41470), .A2(n24649), .B(n8942), .ZN(n41471) );
  NAND2_X1 U51077 ( .A1(n41478), .A2(n62565), .ZN(n41479) );
  AOI21_X1 U51079 ( .A1(n41485), .A2(n61186), .B(n41484), .ZN(n41487) );
  INV_X1 U51084 ( .I(n41497), .ZN(n41499) );
  XOR2_X1 U51085 ( .A1(n41499), .A2(n41498), .Z(n41500) );
  XOR2_X1 U51086 ( .A1(n46279), .A2(n41500), .Z(n41501) );
  NOR2_X1 U51087 ( .A1(n1502), .A2(n42868), .ZN(n41509) );
  INV_X1 U51088 ( .I(n41510), .ZN(n41517) );
  NAND4_X1 U51089 ( .A1(n41514), .A2(n41513), .A3(n41511), .A4(n41512), .ZN(
        n41515) );
  OAI21_X1 U51090 ( .A1(n41517), .A2(n41516), .B(n41515), .ZN(n41518) );
  NAND2_X1 U51092 ( .A1(n41522), .A2(n19928), .ZN(n41523) );
  MUX2_X1 U51093 ( .I0(n41524), .I1(n41523), .S(n1700), .Z(n41536) );
  NAND3_X1 U51098 ( .A1(n42022), .A2(n61372), .A3(n41538), .ZN(n41537) );
  INV_X1 U51100 ( .I(n41796), .ZN(n41543) );
  INV_X1 U51102 ( .I(n42656), .ZN(n41548) );
  NOR2_X1 U51103 ( .A1(n41557), .A2(n42127), .ZN(n41558) );
  NAND2_X1 U51104 ( .A1(n42139), .A2(n10004), .ZN(n41561) );
  NAND2_X1 U51105 ( .A1(n24884), .A2(n42634), .ZN(n41564) );
  NOR2_X1 U51107 ( .A1(n42635), .A2(n11198), .ZN(n41565) );
  NAND2_X1 U51108 ( .A1(n43042), .A2(n61107), .ZN(n41576) );
  NAND2_X1 U51110 ( .A1(n1492), .A2(n1709), .ZN(n41589) );
  NAND2_X1 U51111 ( .A1(n11606), .A2(n8305), .ZN(n43346) );
  NAND2_X1 U51112 ( .A1(n11606), .A2(n59476), .ZN(n41594) );
  NAND2_X1 U51115 ( .A1(n42559), .A2(n20180), .ZN(n41600) );
  OAI22_X1 U51117 ( .A1(n6338), .A2(n64363), .B1(n41600), .B2(n42557), .ZN(
        n41603) );
  NAND3_X1 U51118 ( .A1(n5773), .A2(n42554), .A3(n64363), .ZN(n41601) );
  OAI22_X1 U51119 ( .A1(n41601), .A2(n42551), .B1(n1718), .B2(n42912), .ZN(
        n41602) );
  INV_X1 U51121 ( .I(n41717), .ZN(n41607) );
  NOR2_X1 U51124 ( .A1(n22999), .A2(n9801), .ZN(n41724) );
  OAI21_X1 U51125 ( .A1(n41724), .A2(n1697), .B(n20817), .ZN(n41619) );
  NAND2_X1 U51126 ( .A1(n41619), .A2(n41984), .ZN(n41620) );
  NAND2_X1 U51130 ( .A1(n41629), .A2(n41628), .ZN(n41633) );
  OAI21_X1 U51132 ( .A1(n41631), .A2(n41630), .B(n42158), .ZN(n41632) );
  NOR2_X1 U51133 ( .A1(n41639), .A2(n41638), .ZN(n41646) );
  INV_X1 U51134 ( .I(n41641), .ZN(n41643) );
  NAND2_X1 U51135 ( .A1(n41643), .A2(n41642), .ZN(n41648) );
  INV_X1 U51136 ( .I(n41645), .ZN(n41647) );
  NAND3_X1 U51137 ( .A1(n41652), .A2(n43736), .A3(n15091), .ZN(n41653) );
  NAND2_X1 U51142 ( .A1(n41661), .A2(n42786), .ZN(n41663) );
  NAND3_X1 U51145 ( .A1(n57196), .A2(n9792), .A3(n42784), .ZN(n41668) );
  INV_X1 U51147 ( .I(n41670), .ZN(n42780) );
  NAND2_X1 U51148 ( .A1(n42327), .A2(n42328), .ZN(n41672) );
  MUX2_X1 U51149 ( .I0(n43012), .I1(n41672), .S(n57873), .Z(n41674) );
  OAI21_X1 U51150 ( .A1(n10652), .A2(n5261), .B(n42317), .ZN(n41673) );
  NOR2_X1 U51151 ( .A1(n41674), .A2(n41673), .ZN(n41688) );
  NOR2_X1 U51152 ( .A1(n1252), .A2(n42324), .ZN(n42333) );
  NOR2_X1 U51153 ( .A1(n42325), .A2(n42333), .ZN(n41678) );
  OAI21_X1 U51154 ( .A1(n63036), .A2(n5261), .B(n1252), .ZN(n41676) );
  INV_X1 U51156 ( .I(n41679), .ZN(n41680) );
  INV_X1 U51157 ( .I(n41996), .ZN(n41683) );
  INV_X1 U51158 ( .I(n41684), .ZN(n41685) );
  OAI21_X1 U51160 ( .A1(n59067), .A2(n41695), .B(n42655), .ZN(n41696) );
  AOI21_X1 U51161 ( .A1(n41699), .A2(n11198), .B(n18398), .ZN(n41700) );
  OAI21_X1 U51162 ( .A1(n41701), .A2(n42629), .B(n41700), .ZN(n41707) );
  INV_X1 U51163 ( .I(n42630), .ZN(n41703) );
  OAI21_X1 U51164 ( .A1(n43380), .A2(n43381), .B(n11198), .ZN(n41705) );
  NAND2_X1 U51165 ( .A1(n41720), .A2(n41719), .ZN(n41722) );
  NAND2_X1 U51166 ( .A1(n41722), .A2(n41721), .ZN(n41727) );
  NAND3_X1 U51167 ( .A1(n41724), .A2(n41984), .A3(n64961), .ZN(n41725) );
  OAI22_X1 U51168 ( .A1(n41729), .A2(n17467), .B1(n6705), .B2(n42835), .ZN(
        n41730) );
  NOR2_X1 U51169 ( .A1(n6705), .A2(n42672), .ZN(n42683) );
  NOR2_X1 U51170 ( .A1(n41730), .A2(n42683), .ZN(n41737) );
  NAND2_X1 U51171 ( .A1(n6705), .A2(n42839), .ZN(n41736) );
  NAND3_X1 U51172 ( .A1(n42827), .A2(n1713), .A3(n65185), .ZN(n41734) );
  XOR2_X1 U51173 ( .A1(n41739), .A2(n41738), .Z(n41740) );
  XOR2_X1 U51174 ( .A1(n23210), .A2(n41740), .Z(n41741) );
  NOR2_X1 U51175 ( .A1(n42371), .A2(n43449), .ZN(n41748) );
  NAND2_X1 U51177 ( .A1(n43449), .A2(n43433), .ZN(n41745) );
  INV_X1 U51180 ( .I(n42373), .ZN(n41749) );
  XOR2_X1 U51181 ( .A1(n15735), .A2(n53805), .Z(n41754) );
  NAND2_X1 U51182 ( .A1(n42962), .A2(n42412), .ZN(n41756) );
  AOI21_X1 U51183 ( .A1(n41757), .A2(n13750), .B(n41756), .ZN(n41759) );
  INV_X1 U51185 ( .I(n43167), .ZN(n41768) );
  OAI21_X1 U51186 ( .A1(n42058), .A2(n41768), .B(n42572), .ZN(n41770) );
  NAND3_X1 U51187 ( .A1(n43163), .A2(n42890), .A3(n43169), .ZN(n41769) );
  NOR2_X1 U51189 ( .A1(n42659), .A2(n42139), .ZN(n41782) );
  NOR2_X1 U51190 ( .A1(n41783), .A2(n41782), .ZN(n41786) );
  NOR4_X1 U51191 ( .A1(n8962), .A2(n43130), .A3(n43268), .A4(n1398), .ZN(
        n41787) );
  NAND2_X1 U51192 ( .A1(n41944), .A2(n20227), .ZN(n41798) );
  OAI21_X1 U51193 ( .A1(n664), .A2(n24066), .B(n41805), .ZN(n41807) );
  INV_X1 U51194 ( .I(n42446), .ZN(n41814) );
  OAI21_X1 U51195 ( .A1(n21206), .A2(n41817), .B(n42434), .ZN(n41819) );
  OAI21_X1 U51196 ( .A1(n41819), .A2(n41818), .B(n57208), .ZN(n41822) );
  OAI21_X1 U51198 ( .A1(n42199), .A2(n18717), .B(n42211), .ZN(n41830) );
  NOR2_X1 U51199 ( .A1(n42516), .A2(n42209), .ZN(n41834) );
  NAND2_X1 U51200 ( .A1(n59976), .A2(n42199), .ZN(n41838) );
  INV_X1 U51201 ( .I(n41843), .ZN(n41845) );
  NOR2_X1 U51202 ( .A1(n42304), .A2(n20277), .ZN(n41862) );
  INV_X1 U51203 ( .I(n41853), .ZN(n41855) );
  NAND2_X1 U51204 ( .A1(n43925), .A2(n23488), .ZN(n41865) );
  NAND2_X1 U51205 ( .A1(n9875), .A2(n42526), .ZN(n41866) );
  NAND3_X1 U51206 ( .A1(n42213), .A2(n60947), .A3(n41866), .ZN(n41869) );
  NAND3_X1 U51207 ( .A1(n41871), .A2(n14280), .A3(n64986), .ZN(n41872) );
  INV_X1 U51208 ( .I(n41873), .ZN(n41880) );
  NAND3_X1 U51210 ( .A1(n41886), .A2(n41885), .A3(n41884), .ZN(n41892) );
  NAND3_X1 U51214 ( .A1(n42264), .A2(n11677), .A3(n41904), .ZN(n41909) );
  NAND2_X1 U51215 ( .A1(n42266), .A2(n22502), .ZN(n41908) );
  NAND2_X1 U51216 ( .A1(n42263), .A2(n41906), .ZN(n41907) );
  NAND3_X1 U51217 ( .A1(n41909), .A2(n41908), .A3(n41907), .ZN(n41910) );
  NOR2_X1 U51218 ( .A1(n41918), .A2(n60709), .ZN(n41919) );
  NOR2_X1 U51219 ( .A1(n60709), .A2(n21529), .ZN(n41921) );
  AOI22_X1 U51220 ( .A1(n41924), .A2(n41923), .B1(n41922), .B2(n41921), .ZN(
        n41926) );
  AOI22_X1 U51222 ( .A1(n41929), .A2(n41928), .B1(n42288), .B2(n22713), .ZN(
        n41931) );
  INV_X1 U51223 ( .I(n41945), .ZN(n41940) );
  NOR2_X1 U51225 ( .A1(n59577), .A2(n41949), .ZN(n41948) );
  NAND3_X1 U51227 ( .A1(n41951), .A2(n7519), .A3(n20190), .ZN(n41952) );
  INV_X1 U51228 ( .I(n43624), .ZN(n41958) );
  NAND2_X1 U51229 ( .A1(n41958), .A2(n42097), .ZN(n41959) );
  NOR2_X1 U51230 ( .A1(n43582), .A2(n43569), .ZN(n41961) );
  OAI21_X1 U51231 ( .A1(n41964), .A2(n41963), .B(n41962), .ZN(n41968) );
  NOR2_X1 U51232 ( .A1(n42686), .A2(n42703), .ZN(n41975) );
  NAND2_X1 U51233 ( .A1(n42694), .A2(n19928), .ZN(n41973) );
  AOI21_X1 U51234 ( .A1(n5939), .A2(n41973), .B(n1393), .ZN(n41974) );
  OAI21_X1 U51235 ( .A1(n41975), .A2(n1394), .B(n41974), .ZN(n41976) );
  INV_X1 U51239 ( .I(n43010), .ZN(n41991) );
  NAND3_X1 U51241 ( .A1(n60792), .A2(n42328), .A3(n41996), .ZN(n41998) );
  NAND3_X1 U51242 ( .A1(n8343), .A2(n10203), .A3(n59381), .ZN(n42009) );
  AOI21_X1 U51243 ( .A1(n43000), .A2(n24981), .B(n42009), .ZN(n42010) );
  INV_X1 U51244 ( .I(n43393), .ZN(n42020) );
  INV_X1 U51245 ( .I(n42024), .ZN(n42025) );
  NOR2_X1 U51247 ( .A1(n42607), .A2(n42027), .ZN(n42028) );
  OAI21_X1 U51248 ( .A1(n59898), .A2(n42600), .B(n42605), .ZN(n42030) );
  AOI21_X1 U51249 ( .A1(n60657), .A2(n42032), .B(n42030), .ZN(n42034) );
  NOR3_X1 U51250 ( .A1(n42032), .A2(n8799), .A3(n13825), .ZN(n42033) );
  NAND2_X1 U51251 ( .A1(n20888), .A2(n43516), .ZN(n42036) );
  NOR2_X1 U51252 ( .A1(n43437), .A2(n43433), .ZN(n42050) );
  NAND3_X1 U51253 ( .A1(n43154), .A2(n43150), .A3(n42054), .ZN(n42055) );
  NOR2_X1 U51254 ( .A1(n43156), .A2(n11179), .ZN(n42057) );
  NOR2_X1 U51255 ( .A1(n42968), .A2(n13478), .ZN(n42068) );
  INV_X1 U51256 ( .I(n42070), .ZN(n42069) );
  NAND2_X1 U51257 ( .A1(n42069), .A2(n1336), .ZN(n42071) );
  INV_X1 U51258 ( .I(n43464), .ZN(n42072) );
  NOR2_X1 U51260 ( .A1(n42404), .A2(n42080), .ZN(n42085) );
  INV_X1 U51261 ( .I(n42085), .ZN(n42081) );
  NOR3_X1 U51262 ( .A1(n42082), .A2(n19793), .A3(n42081), .ZN(n42089) );
  NAND2_X1 U51263 ( .A1(n59394), .A2(n59263), .ZN(n42086) );
  OAI22_X1 U51264 ( .A1(n42087), .A2(n42086), .B1(n42085), .B2(n42084), .ZN(
        n42088) );
  INV_X1 U51266 ( .I(n43417), .ZN(n42094) );
  NAND2_X1 U51267 ( .A1(n5001), .A2(n43415), .ZN(n42093) );
  NAND2_X1 U51268 ( .A1(n5001), .A2(n43548), .ZN(n42098) );
  INV_X1 U51269 ( .I(n43410), .ZN(n43565) );
  INV_X1 U51272 ( .I(n42120), .ZN(n42121) );
  AOI21_X1 U51273 ( .A1(n15091), .A2(n43735), .B(n42121), .ZN(n42122) );
  INV_X1 U51274 ( .I(n42659), .ZN(n42126) );
  NOR3_X1 U51276 ( .A1(n42139), .A2(n42670), .A3(n11883), .ZN(n42133) );
  NOR2_X1 U51278 ( .A1(n42139), .A2(n43254), .ZN(n42131) );
  INV_X1 U51281 ( .I(n42146), .ZN(n42147) );
  INV_X1 U51283 ( .I(n42149), .ZN(n42150) );
  NAND3_X1 U51284 ( .A1(n42150), .A2(n1497), .A3(n42152), .ZN(n42153) );
  NAND3_X1 U51285 ( .A1(n43602), .A2(n42585), .A3(n11229), .ZN(n42157) );
  MUX2_X1 U51286 ( .I0(n42157), .I1(n42156), .S(n41624), .Z(n42165) );
  NOR2_X1 U51290 ( .A1(n16850), .A2(n64346), .ZN(n42168) );
  NOR2_X1 U51292 ( .A1(n42171), .A2(n42871), .ZN(n42172) );
  NAND2_X1 U51293 ( .A1(n17848), .A2(n42180), .ZN(n42181) );
  NAND2_X1 U51297 ( .A1(n1689), .A2(n42788), .ZN(n42190) );
  NOR2_X1 U51298 ( .A1(n14605), .A2(n24779), .ZN(n42197) );
  NAND2_X1 U51299 ( .A1(n42199), .A2(n18717), .ZN(n42201) );
  AOI21_X1 U51300 ( .A1(n42202), .A2(n42201), .B(n42200), .ZN(n42204) );
  MUX2_X1 U51301 ( .I0(n42204), .I1(n42203), .S(n57545), .Z(n42223) );
  NOR3_X1 U51302 ( .A1(n42207), .A2(n23501), .A3(n59976), .ZN(n42208) );
  NOR2_X1 U51303 ( .A1(n42209), .A2(n18717), .ZN(n42210) );
  NOR2_X1 U51304 ( .A1(n42215), .A2(n42526), .ZN(n42216) );
  NAND3_X1 U51306 ( .A1(n61394), .A2(n42235), .A3(n22290), .ZN(n42227) );
  NOR2_X1 U51307 ( .A1(n7519), .A2(n42230), .ZN(n42233) );
  OAI22_X1 U51308 ( .A1(n42231), .A2(n22289), .B1(n42237), .B2(n42230), .ZN(
        n42232) );
  AOI21_X1 U51309 ( .A1(n42234), .A2(n42233), .B(n42232), .ZN(n42238) );
  NOR2_X1 U51310 ( .A1(n59531), .A2(n42239), .ZN(n42244) );
  MUX2_X1 U51311 ( .I0(n42244), .I1(n42243), .S(n42242), .Z(n42257) );
  NAND3_X1 U51313 ( .A1(n42252), .A2(n42251), .A3(n61047), .ZN(n42253) );
  NAND3_X1 U51314 ( .A1(n11677), .A2(n9716), .A3(n19938), .ZN(n42270) );
  NOR2_X1 U51315 ( .A1(n1495), .A2(n23314), .ZN(n42291) );
  INV_X1 U51316 ( .I(n42280), .ZN(n42282) );
  NAND2_X1 U51318 ( .A1(n1734), .A2(n42499), .ZN(n42295) );
  NOR2_X1 U51319 ( .A1(n42299), .A2(n42502), .ZN(n42301) );
  NAND3_X1 U51321 ( .A1(n44226), .A2(n43309), .A3(n22716), .ZN(n42312) );
  INV_X1 U51322 ( .I(n42317), .ZN(n42318) );
  NAND2_X1 U51323 ( .A1(n42318), .A2(n42328), .ZN(n42321) );
  NAND2_X1 U51324 ( .A1(n42319), .A2(n42328), .ZN(n42320) );
  OAI21_X1 U51325 ( .A1(n42326), .A2(n43017), .B(n43016), .ZN(n42336) );
  NOR2_X1 U51326 ( .A1(n42327), .A2(n42328), .ZN(n42331) );
  NOR2_X1 U51327 ( .A1(n10652), .A2(n42328), .ZN(n42330) );
  NAND3_X1 U51328 ( .A1(n43014), .A2(n42333), .A3(n42332), .ZN(n42334) );
  AOI21_X1 U51329 ( .A1(n42870), .A2(n42878), .B(n295), .ZN(n42348) );
  NAND3_X1 U51330 ( .A1(n42362), .A2(n64663), .A3(n42360), .ZN(n42363) );
  NOR2_X1 U51335 ( .A1(n43429), .A2(n42373), .ZN(n42374) );
  NAND2_X1 U51337 ( .A1(n42383), .A2(n42697), .ZN(n42384) );
  AOI21_X1 U51338 ( .A1(n42385), .A2(n42384), .B(n42687), .ZN(n42390) );
  NAND2_X1 U51339 ( .A1(n42388), .A2(n42703), .ZN(n42389) );
  NAND2_X1 U51340 ( .A1(n42413), .A2(n42968), .ZN(n42416) );
  NAND2_X1 U51341 ( .A1(n42419), .A2(n43460), .ZN(n42420) );
  AOI22_X1 U51342 ( .A1(n42428), .A2(n22285), .B1(n42427), .B2(n10554), .ZN(
        n42430) );
  NOR2_X1 U51344 ( .A1(n42433), .A2(n42432), .ZN(n42437) );
  AOI21_X1 U51345 ( .A1(n42437), .A2(n42436), .B(n42435), .ZN(n42444) );
  NAND3_X1 U51346 ( .A1(n42439), .A2(n42438), .A3(n22285), .ZN(n42443) );
  NAND3_X1 U51347 ( .A1(n15542), .A2(n42441), .A3(n62018), .ZN(n42442) );
  AOI21_X1 U51349 ( .A1(n6170), .A2(n22759), .B(n664), .ZN(n42457) );
  AOI21_X1 U51350 ( .A1(n42458), .A2(n42457), .B(n24066), .ZN(n42463) );
  AOI22_X1 U51352 ( .A1(n42463), .A2(n61838), .B1(n63795), .B2(n42461), .ZN(
        n42464) );
  NAND2_X1 U51353 ( .A1(n11278), .A2(n42465), .ZN(n42467) );
  MUX2_X1 U51354 ( .I0(n42467), .I1(n42466), .S(n23399), .Z(n42472) );
  INV_X1 U51355 ( .I(n42470), .ZN(n42471) );
  NAND2_X1 U51356 ( .A1(n64914), .A2(n19331), .ZN(n42473) );
  AOI21_X1 U51358 ( .A1(n42478), .A2(n22943), .B(n42477), .ZN(n42482) );
  NAND3_X1 U51359 ( .A1(n64914), .A2(n42480), .A3(n42479), .ZN(n42481) );
  NAND2_X1 U51360 ( .A1(n43299), .A2(n16890), .ZN(n42531) );
  AOI21_X1 U51361 ( .A1(n42486), .A2(n19102), .B(n1738), .ZN(n42492) );
  AOI21_X1 U51362 ( .A1(n20751), .A2(n23654), .B(n42488), .ZN(n42490) );
  INV_X1 U51363 ( .I(n42494), .ZN(n42497) );
  INV_X1 U51364 ( .I(n42495), .ZN(n42496) );
  NAND2_X1 U51365 ( .A1(n42498), .A2(n1505), .ZN(n42501) );
  NAND2_X1 U51366 ( .A1(n1403), .A2(n42499), .ZN(n42500) );
  AOI21_X1 U51367 ( .A1(n42501), .A2(n42500), .B(n988), .ZN(n42515) );
  NAND2_X1 U51368 ( .A1(n42503), .A2(n42502), .ZN(n42505) );
  NAND3_X1 U51369 ( .A1(n42505), .A2(n3534), .A3(n23744), .ZN(n42506) );
  INV_X1 U51370 ( .I(n42510), .ZN(n42511) );
  OAI21_X1 U51371 ( .A1(n42523), .A2(n42522), .B(n14280), .ZN(n42524) );
  OAI21_X1 U51372 ( .A1(n42526), .A2(n9875), .B(n14280), .ZN(n42529) );
  AOI21_X1 U51373 ( .A1(n1299), .A2(n43947), .B(n12864), .ZN(n42530) );
  NAND3_X1 U51374 ( .A1(n42531), .A2(n43300), .A3(n42530), .ZN(n42536) );
  INV_X1 U51375 ( .I(n43958), .ZN(n42532) );
  OAI21_X1 U51376 ( .A1(n43301), .A2(n42532), .B(n59709), .ZN(n42535) );
  NAND3_X1 U51377 ( .A1(n42533), .A2(n59709), .A3(n12864), .ZN(n42534) );
  INV_X1 U51378 ( .I(n42989), .ZN(n42537) );
  NAND2_X1 U51379 ( .A1(n23702), .A2(n63392), .ZN(n42552) );
  NAND2_X1 U51384 ( .A1(n42901), .A2(n64653), .ZN(n42573) );
  INV_X1 U51386 ( .I(n42578), .ZN(n42580) );
  XOR2_X1 U51387 ( .A1(n42580), .A2(n42579), .Z(n42581) );
  XOR2_X1 U51388 ( .A1(n23641), .A2(n42581), .Z(n42591) );
  OAI22_X1 U51389 ( .A1(n43336), .A2(n42584), .B1(n62299), .B2(n43339), .ZN(
        n42586) );
  INV_X1 U51391 ( .I(n42598), .ZN(n42599) );
  NOR2_X1 U51392 ( .A1(n42599), .A2(n42600), .ZN(n42604) );
  NAND2_X1 U51393 ( .A1(n1701), .A2(n2330), .ZN(n42613) );
  NAND2_X1 U51395 ( .A1(n43633), .A2(n62997), .ZN(n43678) );
  NAND3_X1 U51396 ( .A1(n43678), .A2(n43677), .A3(n22553), .ZN(n42623) );
  XOR2_X1 U51397 ( .A1(n43884), .A2(n7264), .Z(n42624) );
  XOR2_X1 U51398 ( .A1(n42625), .A2(n42624), .Z(n42626) );
  NAND2_X1 U51400 ( .A1(n18398), .A2(n11198), .ZN(n42633) );
  INV_X1 U51401 ( .I(n43185), .ZN(n42640) );
  NAND2_X1 U51402 ( .A1(n43196), .A2(n43178), .ZN(n42644) );
  NOR2_X1 U51403 ( .A1(n20351), .A2(n43924), .ZN(n43527) );
  NAND2_X1 U51404 ( .A1(n43923), .A2(n43922), .ZN(n42645) );
  NOR2_X1 U51405 ( .A1(n43925), .A2(n43922), .ZN(n43534) );
  NAND2_X1 U51406 ( .A1(n42654), .A2(n42653), .ZN(n42657) );
  INV_X1 U51407 ( .I(n42848), .ZN(n42663) );
  NAND2_X1 U51408 ( .A1(n42669), .A2(n10004), .ZN(n43251) );
  INV_X1 U51409 ( .I(n42669), .ZN(n42671) );
  NAND2_X1 U51410 ( .A1(n42838), .A2(n42672), .ZN(n42673) );
  NAND2_X1 U51411 ( .A1(n6705), .A2(n42673), .ZN(n42675) );
  NAND2_X1 U51412 ( .A1(n42677), .A2(n65185), .ZN(n42678) );
  NOR2_X1 U51413 ( .A1(n16103), .A2(n42821), .ZN(n42682) );
  AOI21_X1 U51415 ( .A1(n1394), .A2(n42694), .B(n1686), .ZN(n42691) );
  NOR2_X1 U51416 ( .A1(n42697), .A2(n42694), .ZN(n42688) );
  NOR2_X1 U51418 ( .A1(n42696), .A2(n23350), .ZN(n42702) );
  NAND4_X1 U51420 ( .A1(n42704), .A2(n20244), .A3(n42703), .A4(n5939), .ZN(
        n42705) );
  INV_X1 U51421 ( .I(n42710), .ZN(n42713) );
  INV_X1 U51422 ( .I(n42711), .ZN(n42712) );
  XOR2_X1 U51423 ( .A1(n42713), .A2(n42712), .Z(n42714) );
  XOR2_X1 U51424 ( .A1(n24262), .A2(n42714), .Z(n42715) );
  INV_X1 U51428 ( .I(n42730), .ZN(n42731) );
  OAI22_X1 U51429 ( .A1(n43359), .A2(n42740), .B1(n42739), .B2(n23838), .ZN(
        n42741) );
  NOR3_X1 U51430 ( .A1(n43869), .A2(n42750), .A3(n11606), .ZN(n42748) );
  AOI22_X1 U51431 ( .A1(n42755), .A2(n42754), .B1(n42753), .B2(n24715), .ZN(
        n42766) );
  AOI21_X1 U51432 ( .A1(n18398), .A2(n3785), .B(n42757), .ZN(n42758) );
  NAND2_X1 U51434 ( .A1(n42760), .A2(n57651), .ZN(n42761) );
  NAND2_X1 U51435 ( .A1(n42804), .A2(n42807), .ZN(n42768) );
  NAND2_X1 U51439 ( .A1(n42788), .A2(n42785), .ZN(n42783) );
  NAND3_X1 U51441 ( .A1(n1299), .A2(n12864), .A3(n1503), .ZN(n42792) );
  NAND2_X1 U51443 ( .A1(n43297), .A2(n11986), .ZN(n42796) );
  OAI21_X1 U51444 ( .A1(n42808), .A2(n42807), .B(n42806), .ZN(n42809) );
  XOR2_X1 U51445 ( .A1(n22323), .A2(n56180), .Z(n42813) );
  XOR2_X1 U51446 ( .A1(n42814), .A2(n42813), .Z(n42815) );
  INV_X1 U51448 ( .I(n42834), .ZN(n42833) );
  NAND4_X1 U51449 ( .A1(n6705), .A2(n17467), .A3(n65181), .A4(n42821), .ZN(
        n42832) );
  OAI21_X1 U51452 ( .A1(n42833), .A2(n42832), .B(n42831), .ZN(n42841) );
  NOR2_X1 U51455 ( .A1(n24195), .A2(n43657), .ZN(n42855) );
  NAND2_X1 U51457 ( .A1(n42857), .A2(n43234), .ZN(n42863) );
  NAND3_X1 U51458 ( .A1(n60593), .A2(n3696), .A3(n42860), .ZN(n42861) );
  NAND2_X1 U51459 ( .A1(n42871), .A2(n42868), .ZN(n42875) );
  NOR2_X1 U51460 ( .A1(n42876), .A2(n42871), .ZN(n42874) );
  INV_X1 U51461 ( .I(n42875), .ZN(n42879) );
  INV_X1 U51462 ( .I(n42876), .ZN(n42877) );
  NAND3_X1 U51463 ( .A1(n42879), .A2(n63721), .A3(n42877), .ZN(n42883) );
  NAND3_X1 U51464 ( .A1(n42881), .A2(n60952), .A3(n775), .ZN(n42882) );
  NAND2_X1 U51465 ( .A1(n43155), .A2(n15214), .ZN(n42893) );
  NOR2_X1 U51466 ( .A1(n42892), .A2(n42891), .ZN(n42898) );
  AOI21_X1 U51467 ( .A1(n64653), .A2(n42893), .B(n43150), .ZN(n42895) );
  INV_X1 U51469 ( .I(n43157), .ZN(n42899) );
  NAND3_X1 U51471 ( .A1(n42904), .A2(n42903), .A3(n42902), .ZN(n42905) );
  INV_X1 U51473 ( .I(n42925), .ZN(n42928) );
  INV_X1 U51474 ( .I(n43430), .ZN(n42938) );
  NAND2_X1 U51475 ( .A1(n65179), .A2(n43433), .ZN(n42934) );
  NAND2_X1 U51476 ( .A1(n42935), .A2(n42934), .ZN(n42937) );
  AOI21_X1 U51477 ( .A1(n42938), .A2(n42937), .B(n42936), .ZN(n42949) );
  INV_X1 U51478 ( .I(n42939), .ZN(n42943) );
  NAND3_X1 U51480 ( .A1(n42944), .A2(n43437), .A3(n65179), .ZN(n42945) );
  MUX2_X1 U51481 ( .I0(n42945), .I1(n43449), .S(n43444), .Z(n42946) );
  INV_X1 U51482 ( .I(n42950), .ZN(n42951) );
  XOR2_X1 U51483 ( .A1(n50720), .A2(n42951), .Z(n42952) );
  XOR2_X1 U51484 ( .A1(n46164), .A2(n42952), .Z(n42953) );
  XOR2_X1 U51485 ( .A1(n42953), .A2(n1489), .Z(n42954) );
  NOR2_X1 U51487 ( .A1(n44229), .A2(n20526), .ZN(n42958) );
  NOR2_X1 U51488 ( .A1(n43984), .A2(n62462), .ZN(n42957) );
  AOI21_X1 U51489 ( .A1(n42962), .A2(n13750), .B(n42968), .ZN(n42963) );
  NOR2_X1 U51490 ( .A1(n57198), .A2(n13478), .ZN(n42970) );
  NOR2_X1 U51491 ( .A1(n43464), .A2(n42968), .ZN(n42969) );
  OAI21_X1 U51492 ( .A1(n42971), .A2(n42970), .B(n42969), .ZN(n42972) );
  NOR2_X1 U51493 ( .A1(n43302), .A2(n42985), .ZN(n42987) );
  NAND2_X1 U51494 ( .A1(n42987), .A2(n22228), .ZN(n42990) );
  NOR2_X1 U51495 ( .A1(n42995), .A2(n42994), .ZN(n42997) );
  AND2_X1 U51496 ( .A1(n43227), .A2(n43085), .Z(n43004) );
  NOR2_X1 U51497 ( .A1(n43001), .A2(n43222), .ZN(n43002) );
  XOR2_X1 U51498 ( .A1(n23722), .A2(n22923), .Z(n43009) );
  XOR2_X1 U51499 ( .A1(n43006), .A2(n44715), .Z(n43007) );
  XOR2_X1 U51500 ( .A1(n23905), .A2(n43007), .Z(n43008) );
  NAND2_X1 U51501 ( .A1(n43010), .A2(n43011), .ZN(n43020) );
  AOI22_X1 U51502 ( .A1(n43015), .A2(n23184), .B1(n43014), .B2(n43013), .ZN(
        n43019) );
  NOR2_X1 U51503 ( .A1(n43026), .A2(n43025), .ZN(n43032) );
  NAND2_X1 U51504 ( .A1(n43028), .A2(n43027), .ZN(n43030) );
  INV_X1 U51509 ( .I(n43072), .ZN(n43056) );
  NAND2_X1 U51510 ( .A1(n63792), .A2(n43056), .ZN(n43057) );
  NOR2_X1 U51511 ( .A1(n22695), .A2(n22112), .ZN(n43060) );
  XOR2_X1 U51512 ( .A1(n43065), .A2(n22340), .Z(n43066) );
  XOR2_X1 U51513 ( .A1(n46385), .A2(n43066), .Z(n43067) );
  NAND2_X1 U51514 ( .A1(n43205), .A2(n43068), .ZN(n43070) );
  NAND2_X1 U51515 ( .A1(n41350), .A2(n43845), .ZN(n43074) );
  NAND2_X1 U51519 ( .A1(n43080), .A2(n43837), .ZN(n43081) );
  NAND2_X1 U51521 ( .A1(n23700), .A2(n20844), .ZN(n43278) );
  OAI21_X1 U51522 ( .A1(n43290), .A2(n43286), .B(n43278), .ZN(n43113) );
  INV_X1 U51523 ( .I(n43111), .ZN(n43112) );
  NAND2_X1 U51524 ( .A1(n43113), .A2(n43112), .ZN(n43115) );
  NAND2_X1 U51525 ( .A1(n1712), .A2(n7349), .ZN(n43114) );
  INV_X1 U51526 ( .I(n43269), .ZN(n43132) );
  INV_X1 U51527 ( .I(n43135), .ZN(n43137) );
  XOR2_X1 U51528 ( .A1(n45868), .A2(n56976), .Z(n43136) );
  XOR2_X1 U51529 ( .A1(n43137), .A2(n43136), .Z(n43138) );
  NOR3_X1 U51530 ( .A1(n23279), .A2(n43897), .A3(n13037), .ZN(n43139) );
  NAND2_X1 U51531 ( .A1(n23279), .A2(n43655), .ZN(n43141) );
  NOR2_X1 U51532 ( .A1(n2824), .A2(n3696), .ZN(n43651) );
  OAI21_X1 U51533 ( .A1(n43651), .A2(n20183), .B(n61951), .ZN(n43146) );
  NOR3_X1 U51535 ( .A1(n43161), .A2(n15214), .A3(n20601), .ZN(n43162) );
  NAND2_X1 U51537 ( .A1(n43517), .A2(n43504), .ZN(n43175) );
  NOR2_X1 U51539 ( .A1(n43183), .A2(n61744), .ZN(n43187) );
  XOR2_X1 U51540 ( .A1(n43193), .A2(n23306), .Z(n43194) );
  NAND2_X1 U51541 ( .A1(n43196), .A2(n43513), .ZN(n46333) );
  XOR2_X1 U51545 ( .A1(n45325), .A2(n57892), .Z(n43209) );
  NAND2_X1 U51548 ( .A1(n21851), .A2(n15091), .ZN(n43213) );
  OAI21_X1 U51549 ( .A1(n58874), .A2(n43226), .B(n43225), .ZN(n43230) );
  NAND2_X1 U51550 ( .A1(n58874), .A2(n43227), .ZN(n43229) );
  INV_X1 U51551 ( .I(n43231), .ZN(n43232) );
  INV_X1 U51552 ( .I(n43243), .ZN(n43233) );
  NOR2_X1 U51554 ( .A1(n43243), .A2(n43889), .ZN(n43244) );
  XOR2_X1 U51555 ( .A1(n43263), .A2(n43262), .Z(n43264) );
  XOR2_X1 U51556 ( .A1(n23365), .A2(n43264), .Z(n43265) );
  INV_X1 U51558 ( .I(n43278), .ZN(n43279) );
  NAND3_X1 U51559 ( .A1(n43280), .A2(n43290), .A3(n43279), .ZN(n43285) );
  NAND3_X1 U51560 ( .A1(n1712), .A2(n43290), .A3(n7349), .ZN(n43291) );
  INV_X1 U51561 ( .I(n43305), .ZN(n43308) );
  INV_X1 U51562 ( .I(n43990), .ZN(n43310) );
  AOI22_X1 U51563 ( .A1(n43984), .A2(n43311), .B1(n43310), .B2(n43309), .ZN(
        n43315) );
  NAND2_X1 U51564 ( .A1(n43991), .A2(n44226), .ZN(n43313) );
  NOR3_X1 U51565 ( .A1(n43318), .A2(n19428), .A3(n1298), .ZN(n43323) );
  NOR2_X1 U51566 ( .A1(n14605), .A2(n61186), .ZN(n43321) );
  AOI22_X1 U51567 ( .A1(n43321), .A2(n43320), .B1(n14605), .B2(n24779), .ZN(
        n43322) );
  XOR2_X1 U51568 ( .A1(n23767), .A2(n51019), .Z(n43331) );
  XOR2_X1 U51569 ( .A1(n43331), .A2(n43330), .Z(n43333) );
  XOR2_X1 U51570 ( .A1(n21724), .A2(n46282), .Z(n46384) );
  NOR2_X1 U51571 ( .A1(n43873), .A2(n60843), .ZN(n43349) );
  NAND2_X1 U51573 ( .A1(n43346), .A2(n43345), .ZN(n43347) );
  OAI21_X1 U51574 ( .A1(n43349), .A2(n43348), .B(n43347), .ZN(n43356) );
  AOI21_X1 U51575 ( .A1(n43359), .A2(n43358), .B(n13453), .ZN(n43360) );
  INV_X1 U51576 ( .I(n43360), .ZN(n43369) );
  XOR2_X1 U51578 ( .A1(n43370), .A2(n1489), .Z(n43371) );
  XOR2_X1 U51579 ( .A1(n44829), .A2(n43371), .Z(n43372) );
  XOR2_X1 U51580 ( .A1(n1039), .A2(n43372), .Z(n43407) );
  AOI21_X1 U51581 ( .A1(n43375), .A2(n43374), .B(n43373), .ZN(n43379) );
  NAND2_X1 U51582 ( .A1(n43380), .A2(n577), .ZN(n43387) );
  NAND2_X1 U51583 ( .A1(n18398), .A2(n43381), .ZN(n43384) );
  OAI22_X1 U51584 ( .A1(n59288), .A2(n43384), .B1(n65228), .B2(n577), .ZN(
        n43386) );
  AOI21_X1 U51585 ( .A1(n59517), .A2(n43387), .B(n43386), .ZN(n43389) );
  XOR2_X1 U51586 ( .A1(n63448), .A2(n22376), .Z(n43403) );
  INV_X1 U51588 ( .I(n43395), .ZN(n43396) );
  INV_X1 U51589 ( .I(n43398), .ZN(n43400) );
  XOR2_X1 U51590 ( .A1(n43400), .A2(n43399), .Z(n43401) );
  XOR2_X1 U51591 ( .A1(n43403), .A2(n43402), .Z(n43404) );
  XOR2_X1 U51592 ( .A1(n43405), .A2(n43404), .Z(n43406) );
  NOR2_X1 U51595 ( .A1(n43553), .A2(n43624), .ZN(n43423) );
  NOR3_X1 U51596 ( .A1(n65179), .A2(n43438), .A3(n43437), .ZN(n43427) );
  NAND3_X1 U51598 ( .A1(n43430), .A2(n43435), .A3(n43429), .ZN(n43431) );
  MUX2_X1 U51599 ( .I0(n43432), .I1(n43431), .S(n62001), .Z(n43452) );
  NAND2_X1 U51600 ( .A1(n43436), .A2(n43435), .ZN(n43443) );
  OAI21_X1 U51601 ( .A1(n43438), .A2(n43437), .B(n65179), .ZN(n43440) );
  NAND4_X1 U51602 ( .A1(n43440), .A2(n43439), .A3(n25806), .A4(n43447), .ZN(
        n43441) );
  NOR3_X1 U51604 ( .A1(n58530), .A2(n43454), .A3(n43467), .ZN(n43455) );
  NAND3_X1 U51606 ( .A1(n43459), .A2(n1193), .A3(n43458), .ZN(n43466) );
  AOI22_X1 U51607 ( .A1(n43462), .A2(n13750), .B1(n43460), .B2(n13478), .ZN(
        n43465) );
  INV_X1 U51609 ( .I(n43467), .ZN(n43470) );
  NOR2_X1 U51610 ( .A1(n43470), .A2(n43469), .ZN(n43473) );
  INV_X1 U51611 ( .I(n43471), .ZN(n43472) );
  NAND4_X2 U51613 ( .A1(n43482), .A2(n43481), .A3(n43480), .A4(n43479), .ZN(
        n45015) );
  XOR2_X1 U51614 ( .A1(n46674), .A2(n3750), .Z(n43483) );
  XOR2_X1 U51615 ( .A1(n46271), .A2(n43483), .Z(n43484) );
  NAND2_X1 U51616 ( .A1(n43490), .A2(n16864), .ZN(n43492) );
  NAND2_X1 U51617 ( .A1(n43531), .A2(n21073), .ZN(n43494) );
  INV_X1 U51619 ( .I(n43497), .ZN(n50870) );
  XOR2_X1 U51620 ( .A1(n50870), .A2(n43498), .Z(n43499) );
  NAND2_X1 U51621 ( .A1(n43504), .A2(n61442), .ZN(n43505) );
  NAND2_X1 U51622 ( .A1(n43510), .A2(n43517), .ZN(n43525) );
  INV_X1 U51629 ( .I(n43527), .ZN(n43530) );
  NOR2_X1 U51630 ( .A1(n23488), .A2(n61743), .ZN(n43528) );
  INV_X1 U51631 ( .I(n43531), .ZN(n43533) );
  AOI22_X1 U51632 ( .A1(n43535), .A2(n43534), .B1(n43533), .B2(n43532), .ZN(
        n43547) );
  NAND2_X1 U51633 ( .A1(n15695), .A2(n21073), .ZN(n43537) );
  AOI21_X1 U51634 ( .A1(n43537), .A2(n43536), .B(n279), .ZN(n43545) );
  NAND3_X1 U51636 ( .A1(n43540), .A2(n43912), .A3(n43539), .ZN(n43543) );
  NAND2_X1 U51637 ( .A1(n43541), .A2(n15695), .ZN(n43542) );
  OAI21_X1 U51639 ( .A1(n59682), .A2(n43548), .B(n16447), .ZN(n43550) );
  NOR2_X1 U51640 ( .A1(n62997), .A2(n43550), .ZN(n43551) );
  NAND2_X1 U51641 ( .A1(n43552), .A2(n43551), .ZN(n43555) );
  INV_X1 U51642 ( .I(n43556), .ZN(n43563) );
  INV_X1 U51643 ( .I(n43627), .ZN(n43557) );
  NAND2_X1 U51644 ( .A1(n1296), .A2(n43557), .ZN(n43560) );
  NAND2_X1 U51645 ( .A1(n5972), .A2(n22087), .ZN(n43558) );
  OAI21_X1 U51646 ( .A1(n43565), .A2(n5972), .B(n43564), .ZN(n43567) );
  NAND2_X1 U51647 ( .A1(n43567), .A2(n43566), .ZN(n43568) );
  INV_X1 U51649 ( .I(n43579), .ZN(n43580) );
  INV_X1 U51650 ( .I(n43587), .ZN(n43589) );
  XOR2_X1 U51651 ( .A1(n43589), .A2(n43588), .Z(n43590) );
  XOR2_X1 U51652 ( .A1(n22731), .A2(n43590), .Z(n43591) );
  XOR2_X1 U51653 ( .A1(n43591), .A2(n44480), .Z(n43592) );
  XOR2_X1 U51655 ( .A1(n45811), .A2(n45823), .Z(n45365) );
  XOR2_X1 U51656 ( .A1(n45365), .A2(n43592), .Z(n43593) );
  XOR2_X1 U51660 ( .A1(n51234), .A2(n43615), .Z(n43616) );
  XOR2_X1 U51661 ( .A1(n52329), .A2(n43616), .Z(n43617) );
  XOR2_X1 U51662 ( .A1(n43617), .A2(n45359), .Z(n43618) );
  XOR2_X1 U51664 ( .A1(n61363), .A2(n20919), .Z(n43620) );
  XOR2_X1 U51665 ( .A1(n44465), .A2(n43620), .Z(n43621) );
  XOR2_X1 U51666 ( .A1(n46442), .A2(n44238), .Z(n43622) );
  XOR2_X1 U51667 ( .A1(n44639), .A2(n43622), .Z(n45428) );
  NOR2_X1 U51668 ( .A1(n43627), .A2(n5972), .ZN(n43630) );
  AOI22_X1 U51670 ( .A1(n43635), .A2(n43631), .B1(n43630), .B2(n43629), .ZN(
        n43638) );
  NAND2_X1 U51671 ( .A1(n62072), .A2(n63983), .ZN(n43637) );
  AOI21_X1 U51672 ( .A1(n43635), .A2(n43634), .B(n43633), .ZN(n43636) );
  XOR2_X1 U51673 ( .A1(n6967), .A2(n43640), .Z(n44061) );
  INV_X1 U51674 ( .I(n43641), .ZN(n43643) );
  XOR2_X1 U51675 ( .A1(n43643), .A2(n43642), .Z(n43644) );
  XOR2_X1 U51676 ( .A1(n43645), .A2(n43644), .Z(n43646) );
  XOR2_X1 U51677 ( .A1(n61142), .A2(n43646), .Z(n43647) );
  XOR2_X1 U51678 ( .A1(n43647), .A2(n46621), .Z(n43648) );
  NAND3_X1 U51679 ( .A1(n43658), .A2(n20183), .A3(n43657), .ZN(n43659) );
  INV_X1 U51680 ( .I(n24521), .ZN(n43665) );
  XOR2_X1 U51681 ( .A1(n55150), .A2(n53764), .Z(n43666) );
  XOR2_X1 U51682 ( .A1(n43667), .A2(n43666), .Z(n43668) );
  XOR2_X1 U51683 ( .A1(n51071), .A2(n43668), .Z(n43669) );
  XOR2_X1 U51684 ( .A1(n43670), .A2(n43669), .Z(n43671) );
  NAND2_X1 U51685 ( .A1(n43678), .A2(n43677), .ZN(n43680) );
  XOR2_X1 U51686 ( .A1(n43683), .A2(n43682), .Z(n43684) );
  XOR2_X1 U51688 ( .A1(n43687), .A2(n46520), .Z(n45299) );
  INV_X1 U51689 ( .I(n45299), .ZN(n43688) );
  NAND2_X1 U51693 ( .A1(n24071), .A2(n1334), .ZN(n43713) );
  XOR2_X1 U51694 ( .A1(n43960), .A2(n24094), .Z(n43725) );
  INV_X1 U51695 ( .I(n43720), .ZN(n43722) );
  XOR2_X1 U51696 ( .A1(n43722), .A2(n43721), .Z(n43723) );
  XOR2_X1 U51697 ( .A1(n44442), .A2(n46587), .Z(n43727) );
  XOR2_X1 U51698 ( .A1(n43727), .A2(n22247), .Z(n45099) );
  XOR2_X1 U51701 ( .A1(n43728), .A2(n51021), .Z(n43729) );
  XOR2_X1 U51702 ( .A1(n43730), .A2(n43729), .Z(n43731) );
  XOR2_X1 U51704 ( .A1(n44940), .A2(n43732), .Z(n43743) );
  NAND2_X1 U51705 ( .A1(n43734), .A2(n43733), .ZN(n43737) );
  XOR2_X1 U51707 ( .A1(n45021), .A2(n46212), .Z(n43745) );
  NOR2_X1 U51708 ( .A1(n46744), .A2(n43747), .ZN(n43756) );
  OAI21_X1 U51709 ( .A1(n47431), .A2(n64096), .B(n43752), .ZN(n43753) );
  INV_X1 U51711 ( .I(n43758), .ZN(n43761) );
  XOR2_X1 U51712 ( .A1(n31347), .A2(n43759), .Z(n43760) );
  XOR2_X1 U51713 ( .A1(n43761), .A2(n43760), .Z(n43762) );
  XOR2_X1 U51714 ( .A1(n23210), .A2(n43762), .Z(n43763) );
  XOR2_X1 U51716 ( .A1(n50787), .A2(n43768), .Z(n43769) );
  XOR2_X1 U51717 ( .A1(n43770), .A2(n43769), .Z(n43771) );
  XOR2_X1 U51718 ( .A1(n43772), .A2(n43771), .Z(n43773) );
  XOR2_X1 U51719 ( .A1(n43784), .A2(n43783), .Z(n43785) );
  XOR2_X1 U51720 ( .A1(n46343), .A2(n43785), .Z(n43786) );
  INV_X1 U51721 ( .I(n43787), .ZN(n43792) );
  XOR2_X1 U51722 ( .A1(n43788), .A2(n55150), .Z(n43790) );
  XOR2_X1 U51723 ( .A1(n43790), .A2(n43789), .Z(n43791) );
  XOR2_X1 U51724 ( .A1(n43792), .A2(n43791), .Z(n43793) );
  XOR2_X1 U51725 ( .A1(n6872), .A2(n43793), .Z(n43794) );
  INV_X1 U51726 ( .I(n43798), .ZN(n43801) );
  INV_X1 U51727 ( .I(n43799), .ZN(n43800) );
  XOR2_X1 U51728 ( .A1(n43801), .A2(n43800), .Z(n43802) );
  XOR2_X1 U51729 ( .A1(n43803), .A2(n43802), .Z(n43804) );
  XOR2_X1 U51730 ( .A1(n23818), .A2(n43804), .Z(n43805) );
  XOR2_X1 U51731 ( .A1(n43805), .A2(n44480), .Z(n43806) );
  INV_X1 U51734 ( .I(n43808), .ZN(n43810) );
  XOR2_X1 U51735 ( .A1(n43810), .A2(n43809), .Z(n43811) );
  NAND3_X1 U51736 ( .A1(n43817), .A2(n43816), .A3(n43815), .ZN(n43818) );
  XOR2_X1 U51737 ( .A1(n44911), .A2(n22207), .Z(n45263) );
  XOR2_X1 U51739 ( .A1(n46538), .A2(n56008), .Z(n45423) );
  XOR2_X1 U51740 ( .A1(n44639), .A2(n23828), .Z(n43822) );
  XOR2_X1 U51741 ( .A1(n45423), .A2(n43822), .Z(n43823) );
  NAND2_X1 U51743 ( .A1(n637), .A2(n47858), .ZN(n43830) );
  OAI22_X1 U51745 ( .A1(n43848), .A2(n43847), .B1(n41350), .B2(n43846), .ZN(
        n43849) );
  INV_X1 U51746 ( .I(n21170), .ZN(n43856) );
  XOR2_X1 U51747 ( .A1(n43858), .A2(n43857), .Z(n43859) );
  XOR2_X1 U51748 ( .A1(n43860), .A2(n43859), .Z(n43861) );
  XOR2_X1 U51749 ( .A1(n6872), .A2(n43861), .Z(n43862) );
  INV_X1 U51750 ( .I(n43864), .ZN(n43865) );
  XOR2_X1 U51751 ( .A1(n23365), .A2(n43865), .Z(n43866) );
  XOR2_X1 U51755 ( .A1(n44897), .A2(n43880), .Z(n44738) );
  XNOR2_X1 U51756 ( .A1(n56849), .A2(n52317), .ZN(n43881) );
  XOR2_X1 U51757 ( .A1(n43882), .A2(n43881), .Z(n43883) );
  XOR2_X1 U51758 ( .A1(n43884), .A2(n43883), .Z(n43885) );
  XOR2_X1 U51759 ( .A1(n21142), .A2(n43885), .Z(n43886) );
  XOR2_X1 U51760 ( .A1(n43886), .A2(n44738), .Z(n43887) );
  NAND4_X1 U51762 ( .A1(n23279), .A2(n13037), .A3(n63818), .A4(n43889), .ZN(
        n43895) );
  OAI21_X1 U51764 ( .A1(n43893), .A2(n43892), .B(n43891), .ZN(n43894) );
  XOR2_X1 U51765 ( .A1(n43901), .A2(n43900), .Z(n43903) );
  XOR2_X1 U51766 ( .A1(n43903), .A2(n43902), .Z(n43904) );
  XOR2_X1 U51767 ( .A1(n43906), .A2(n43905), .Z(n43907) );
  XOR2_X1 U51768 ( .A1(n43907), .A2(n45376), .Z(n43908) );
  INV_X1 U51769 ( .I(n43910), .ZN(n43911) );
  INV_X1 U51770 ( .I(n43913), .ZN(n43920) );
  INV_X1 U51771 ( .I(n43914), .ZN(n43919) );
  NOR2_X1 U51772 ( .A1(n43923), .A2(n43922), .ZN(n43928) );
  AOI21_X1 U51773 ( .A1(n43928), .A2(n43927), .B(n43926), .ZN(n43931) );
  NAND2_X1 U51774 ( .A1(n4467), .A2(n23488), .ZN(n43930) );
  INV_X1 U51776 ( .I(n43933), .ZN(n43934) );
  XOR2_X1 U51778 ( .A1(n43937), .A2(n43936), .Z(n43938) );
  XOR2_X1 U51779 ( .A1(n45333), .A2(n43939), .Z(n43942) );
  XOR2_X1 U51780 ( .A1(n43940), .A2(n43941), .Z(n44247) );
  INV_X1 U51781 ( .I(n44911), .ZN(n43945) );
  XOR2_X1 U51782 ( .A1(n62873), .A2(n43945), .Z(n43946) );
  INV_X1 U51783 ( .I(n43962), .ZN(n43965) );
  XOR2_X1 U51784 ( .A1(n43963), .A2(n55903), .Z(n43964) );
  XOR2_X1 U51785 ( .A1(n43965), .A2(n43964), .Z(n43966) );
  XOR2_X1 U51786 ( .A1(n43967), .A2(n44480), .Z(n45271) );
  XOR2_X1 U51787 ( .A1(n50909), .A2(n43968), .Z(n43970) );
  XOR2_X1 U51788 ( .A1(n43970), .A2(n43969), .Z(n43972) );
  XOR2_X1 U51789 ( .A1(n43972), .A2(n43971), .Z(n43973) );
  XOR2_X1 U51790 ( .A1(n51680), .A2(n43973), .Z(n43974) );
  INV_X1 U51791 ( .I(n43975), .ZN(n43976) );
  AOI21_X1 U51792 ( .A1(n44230), .A2(n43981), .B(n44228), .ZN(n43982) );
  NAND2_X1 U51793 ( .A1(n45203), .A2(n25896), .ZN(n45201) );
  NAND3_X1 U51796 ( .A1(n1375), .A2(n57949), .A3(n44003), .ZN(n44008) );
  NAND3_X1 U51797 ( .A1(n48869), .A2(n49389), .A3(n44003), .ZN(n44007) );
  NAND2_X1 U51798 ( .A1(n44005), .A2(n49395), .ZN(n44006) );
  XOR2_X1 U51802 ( .A1(n46387), .A2(n51021), .Z(n44015) );
  XOR2_X1 U51803 ( .A1(n50102), .A2(n44015), .Z(n44016) );
  XOR2_X1 U51806 ( .A1(n46211), .A2(n56692), .Z(n44360) );
  XOR2_X1 U51807 ( .A1(n25638), .A2(n53530), .Z(n44254) );
  INV_X1 U51808 ( .I(n44023), .ZN(n44026) );
  XOR2_X1 U51809 ( .A1(n44024), .A2(n50475), .Z(n44025) );
  XOR2_X1 U51810 ( .A1(n44026), .A2(n44025), .Z(n44027) );
  INV_X1 U51811 ( .I(n46135), .ZN(n44036) );
  INV_X1 U51812 ( .I(n44030), .ZN(n44031) );
  XOR2_X1 U51813 ( .A1(n44032), .A2(n44031), .Z(n44033) );
  XOR2_X1 U51814 ( .A1(n44034), .A2(n46136), .Z(n44035) );
  XOR2_X1 U51815 ( .A1(n23987), .A2(n46208), .Z(n44039) );
  XOR2_X1 U51816 ( .A1(n44039), .A2(n44501), .Z(n44044) );
  XOR2_X1 U51817 ( .A1(n44040), .A2(n23253), .Z(n44042) );
  XOR2_X1 U51818 ( .A1(n44042), .A2(n44041), .Z(n44043) );
  XOR2_X1 U51819 ( .A1(n5011), .A2(n44223), .Z(n44050) );
  INV_X1 U51820 ( .I(n44047), .ZN(n44048) );
  XOR2_X1 U51821 ( .A1(n50741), .A2(n44048), .Z(n44049) );
  XOR2_X1 U51822 ( .A1(n4529), .A2(n20950), .Z(n44051) );
  XOR2_X1 U51823 ( .A1(n44052), .A2(n52226), .Z(n44053) );
  XOR2_X1 U51824 ( .A1(n44054), .A2(n44053), .Z(n44055) );
  XOR2_X1 U51825 ( .A1(n44056), .A2(n44055), .Z(n44057) );
  XOR2_X1 U51826 ( .A1(n44057), .A2(n23828), .Z(n44058) );
  XOR2_X1 U51827 ( .A1(n44120), .A2(n44058), .Z(n44059) );
  XOR2_X1 U51828 ( .A1(n44060), .A2(n44920), .Z(n44063) );
  INV_X1 U51829 ( .I(n44061), .ZN(n44062) );
  NOR2_X1 U51830 ( .A1(n47468), .A2(n20917), .ZN(n44068) );
  INV_X1 U51834 ( .I(n2826), .ZN(n44073) );
  INV_X1 U51835 ( .I(n46984), .ZN(n44072) );
  NAND2_X1 U51836 ( .A1(n45740), .A2(n20917), .ZN(n44071) );
  INV_X1 U51838 ( .I(n50199), .ZN(n44080) );
  XOR2_X1 U51839 ( .A1(n44078), .A2(n55833), .Z(n44079) );
  XOR2_X1 U51840 ( .A1(n44080), .A2(n44079), .Z(n44081) );
  XOR2_X1 U51841 ( .A1(n44082), .A2(n44252), .Z(n44083) );
  XOR2_X1 U51842 ( .A1(n23722), .A2(n23078), .Z(n44090) );
  XOR2_X1 U51843 ( .A1(n44085), .A2(n30908), .Z(n44086) );
  XOR2_X1 U51844 ( .A1(n44087), .A2(n44086), .Z(n44088) );
  XOR2_X1 U51845 ( .A1(n44093), .A2(n57113), .Z(n44096) );
  INV_X1 U51846 ( .I(n44094), .ZN(n44095) );
  XOR2_X1 U51847 ( .A1(n44096), .A2(n44095), .Z(n44097) );
  INV_X1 U51848 ( .I(n44356), .ZN(n45859) );
  XOR2_X1 U51849 ( .A1(n44100), .A2(n44099), .Z(n44101) );
  XOR2_X1 U51850 ( .A1(n44103), .A2(n44102), .Z(n44105) );
  XOR2_X1 U51852 ( .A1(n44107), .A2(n46682), .Z(n44111) );
  XOR2_X1 U51853 ( .A1(n44109), .A2(n44108), .Z(n44110) );
  XOR2_X1 U51854 ( .A1(n44111), .A2(n44110), .Z(n44113) );
  XOR2_X1 U51855 ( .A1(n44112), .A2(n44113), .Z(n44114) );
  XOR2_X1 U51856 ( .A1(n44115), .A2(n44465), .Z(n44117) );
  XOR2_X1 U51858 ( .A1(n44121), .A2(n23445), .Z(n44122) );
  XOR2_X1 U51859 ( .A1(n44124), .A2(n44123), .Z(n44125) );
  XOR2_X1 U51860 ( .A1(n44125), .A2(n65144), .Z(n44126) );
  XOR2_X1 U51861 ( .A1(n44127), .A2(n45428), .Z(n44128) );
  XOR2_X1 U51862 ( .A1(n46436), .A2(n44130), .Z(n44131) );
  XOR2_X1 U51863 ( .A1(n44225), .A2(n44131), .Z(n44132) );
  XOR2_X1 U51864 ( .A1(n44138), .A2(n44137), .Z(n44140) );
  XOR2_X1 U51865 ( .A1(n44140), .A2(n44139), .Z(n44141) );
  XOR2_X1 U51866 ( .A1(n46279), .A2(n44141), .Z(n44142) );
  INV_X1 U51867 ( .I(n52527), .ZN(n44150) );
  XOR2_X1 U51868 ( .A1(n44148), .A2(n45348), .Z(n44149) );
  XOR2_X1 U51869 ( .A1(n44150), .A2(n44149), .Z(n44151) );
  XOR2_X1 U51870 ( .A1(n46557), .A2(n44151), .Z(n44152) );
  XOR2_X1 U51871 ( .A1(n10043), .A2(n44152), .Z(n44153) );
  XOR2_X1 U51872 ( .A1(n51654), .A2(n56879), .Z(n44157) );
  XOR2_X1 U51873 ( .A1(n52069), .A2(n44157), .Z(n44158) );
  XOR2_X1 U51874 ( .A1(n16299), .A2(n44158), .Z(n44159) );
  XOR2_X1 U51875 ( .A1(n10304), .A2(n7264), .Z(n44166) );
  INV_X1 U51876 ( .I(n44164), .ZN(n44165) );
  XOR2_X1 U51877 ( .A1(n44166), .A2(n44165), .Z(n44167) );
  XOR2_X1 U51878 ( .A1(n11317), .A2(n44167), .Z(n44168) );
  XOR2_X1 U51879 ( .A1(n46307), .A2(n46188), .Z(n44175) );
  INV_X1 U51880 ( .I(n50578), .ZN(n44171) );
  XOR2_X1 U51881 ( .A1(n44171), .A2(n44170), .Z(n44172) );
  XOR2_X1 U51882 ( .A1(n23426), .A2(n44172), .Z(n44173) );
  XOR2_X1 U51883 ( .A1(n44175), .A2(n44174), .Z(n44176) );
  XOR2_X1 U51884 ( .A1(n24021), .A2(n55034), .Z(n44906) );
  XOR2_X1 U51885 ( .A1(n44909), .A2(n23828), .Z(n44178) );
  XOR2_X1 U51886 ( .A1(n44906), .A2(n44178), .Z(n44179) );
  XOR2_X1 U51887 ( .A1(n60227), .A2(n44179), .Z(n44180) );
  XOR2_X1 U51888 ( .A1(n44182), .A2(n4686), .Z(n44183) );
  XOR2_X1 U51889 ( .A1(n44186), .A2(n44185), .Z(n44187) );
  XOR2_X1 U51890 ( .A1(n65082), .A2(n44187), .Z(n44188) );
  INV_X1 U51891 ( .I(n45366), .ZN(n44192) );
  XOR2_X1 U51892 ( .A1(n44191), .A2(n44192), .Z(n44193) );
  NAND2_X2 U51895 ( .A1(n45765), .A2(n46913), .ZN(n46906) );
  NAND3_X1 U51898 ( .A1(n1388), .A2(n22326), .A3(n1267), .ZN(n44201) );
  NOR2_X1 U51899 ( .A1(n1267), .A2(n10512), .ZN(n44202) );
  AOI21_X1 U51900 ( .A1(n44202), .A2(n23990), .B(n46905), .ZN(n44203) );
  NAND2_X1 U51901 ( .A1(n15666), .A2(n45765), .ZN(n44661) );
  NAND3_X1 U51902 ( .A1(n44205), .A2(n46913), .A3(n44661), .ZN(n44208) );
  NAND3_X1 U51904 ( .A1(n9972), .A2(n57731), .A3(n45766), .ZN(n44206) );
  INV_X1 U51905 ( .I(n44211), .ZN(n44216) );
  XOR2_X1 U51906 ( .A1(n44212), .A2(n58084), .Z(n44213) );
  XOR2_X1 U51907 ( .A1(n44213), .A2(n52135), .Z(n44214) );
  XOR2_X1 U51908 ( .A1(n44214), .A2(n50247), .Z(n44215) );
  XOR2_X1 U51909 ( .A1(n44216), .A2(n44215), .Z(n44217) );
  XOR2_X1 U51910 ( .A1(n44219), .A2(n44218), .Z(n44222) );
  INV_X1 U51911 ( .I(n12153), .ZN(n44220) );
  XOR2_X1 U51913 ( .A1(n46451), .A2(n44225), .Z(n44250) );
  NOR3_X1 U51914 ( .A1(n44230), .A2(n62462), .A3(n44226), .ZN(n44233) );
  AOI21_X1 U51915 ( .A1(n44230), .A2(n44229), .B(n44228), .ZN(n44231) );
  NOR3_X1 U51916 ( .A1(n44233), .A2(n44232), .A3(n44231), .ZN(n44236) );
  INV_X1 U51917 ( .I(n44234), .ZN(n44235) );
  NAND3_X1 U51918 ( .A1(n44237), .A2(n44236), .A3(n44235), .ZN(n44239) );
  XOR2_X1 U51919 ( .A1(n44238), .A2(n44239), .Z(n44367) );
  XOR2_X1 U51920 ( .A1(n44241), .A2(n44240), .Z(n44243) );
  XOR2_X1 U51921 ( .A1(n44243), .A2(n23828), .Z(n44244) );
  XOR2_X1 U51922 ( .A1(n44367), .A2(n44244), .Z(n44245) );
  XOR2_X1 U51923 ( .A1(n44909), .A2(n24278), .Z(n46163) );
  XOR2_X1 U51924 ( .A1(n44247), .A2(n44246), .Z(n44248) );
  XOR2_X1 U51925 ( .A1(n44249), .A2(n44250), .Z(n44670) );
  INV_X1 U51926 ( .I(n45865), .ZN(n44253) );
  INV_X1 U51927 ( .I(n44255), .ZN(n44256) );
  XOR2_X1 U51928 ( .A1(n44257), .A2(n44256), .Z(n44258) );
  XOR2_X1 U51930 ( .A1(n7544), .A2(n22950), .Z(n46218) );
  INV_X1 U51931 ( .I(n44263), .ZN(n44265) );
  XOR2_X1 U51932 ( .A1(n44265), .A2(n44264), .Z(n44266) );
  XOR2_X1 U51933 ( .A1(n46218), .A2(n44266), .Z(n44267) );
  INV_X1 U51934 ( .I(n44274), .ZN(n44276) );
  XOR2_X1 U51935 ( .A1(n44276), .A2(n44275), .Z(n44277) );
  XOR2_X1 U51936 ( .A1(n11317), .A2(n44277), .Z(n44278) );
  XOR2_X1 U51937 ( .A1(n44278), .A2(n44329), .Z(n44279) );
  OAI21_X1 U51938 ( .A1(n65275), .A2(n12850), .B(n61980), .ZN(n44282) );
  NAND3_X1 U51941 ( .A1(n1086), .A2(n47517), .A3(n47503), .ZN(n44287) );
  XOR2_X1 U51942 ( .A1(n44290), .A2(n58077), .Z(n44292) );
  XOR2_X1 U51943 ( .A1(n44292), .A2(n44291), .Z(n44293) );
  XOR2_X1 U51944 ( .A1(n52970), .A2(n53246), .Z(n44296) );
  XOR2_X1 U51945 ( .A1(n44297), .A2(n44296), .Z(n44298) );
  XOR2_X1 U51946 ( .A1(n44299), .A2(n44298), .Z(n44300) );
  XOR2_X1 U51947 ( .A1(n44301), .A2(n46197), .Z(n44303) );
  XOR2_X1 U51948 ( .A1(n61142), .A2(n22639), .Z(n44302) );
  XOR2_X1 U51949 ( .A1(n46166), .A2(n51493), .Z(n44304) );
  XOR2_X1 U51953 ( .A1(n44309), .A2(n52135), .Z(n44310) );
  XOR2_X1 U51954 ( .A1(n44311), .A2(n44310), .Z(n44312) );
  XOR2_X1 U51955 ( .A1(n44312), .A2(n45819), .Z(n44313) );
  XOR2_X1 U51956 ( .A1(n44314), .A2(n20919), .Z(n44315) );
  XOR2_X1 U51957 ( .A1(n65082), .A2(n44467), .Z(n44316) );
  XOR2_X1 U51959 ( .A1(n30402), .A2(n55150), .Z(n44322) );
  XOR2_X1 U51960 ( .A1(n44323), .A2(n44322), .Z(n44324) );
  XOR2_X1 U51961 ( .A1(n44325), .A2(n44324), .Z(n44326) );
  XOR2_X1 U51964 ( .A1(n44331), .A2(n44330), .Z(n51323) );
  XOR2_X1 U51965 ( .A1(n44332), .A2(n56309), .Z(n44333) );
  XOR2_X1 U51966 ( .A1(n18098), .A2(n44334), .Z(n44336) );
  XOR2_X1 U51967 ( .A1(n24090), .A2(n21141), .Z(n44337) );
  XOR2_X1 U51968 ( .A1(n51516), .A2(n44339), .Z(n44340) );
  XOR2_X1 U51969 ( .A1(n10255), .A2(n44340), .Z(n44341) );
  OAI21_X1 U51971 ( .A1(n10563), .A2(n23738), .B(n48324), .ZN(n44407) );
  XOR2_X1 U51972 ( .A1(n44346), .A2(n44345), .Z(n44347) );
  XOR2_X1 U51973 ( .A1(n24521), .A2(n44347), .Z(n44348) );
  XOR2_X1 U51974 ( .A1(n44351), .A2(n44350), .Z(n44352) );
  XOR2_X1 U51975 ( .A1(n44358), .A2(n44357), .Z(n44359) );
  INV_X1 U51977 ( .I(n44363), .ZN(n44364) );
  XOR2_X1 U51978 ( .A1(n44365), .A2(n44364), .Z(n44366) );
  XOR2_X1 U51979 ( .A1(n44368), .A2(n44367), .Z(n44370) );
  INV_X1 U51981 ( .I(n45429), .ZN(n44373) );
  XOR2_X1 U51982 ( .A1(n44373), .A2(n44372), .Z(n44374) );
  XOR2_X1 U51983 ( .A1(n44375), .A2(n44374), .Z(n44376) );
  INV_X1 U51984 ( .I(n4686), .ZN(n44847) );
  INV_X1 U51985 ( .I(n47341), .ZN(n44381) );
  XOR2_X1 U51986 ( .A1(n44759), .A2(n44378), .Z(n44379) );
  XOR2_X1 U51987 ( .A1(n49445), .A2(n44379), .Z(n44380) );
  XOR2_X1 U51988 ( .A1(n44381), .A2(n44380), .Z(n44382) );
  XOR2_X1 U51989 ( .A1(n45040), .A2(n44382), .Z(n44383) );
  INV_X1 U51991 ( .I(n44390), .ZN(n44393) );
  XOR2_X1 U51992 ( .A1(n44391), .A2(n50787), .Z(n44392) );
  XOR2_X1 U51993 ( .A1(n44393), .A2(n44392), .Z(n44394) );
  NAND3_X1 U51995 ( .A1(n45779), .A2(n61563), .A3(n1294), .ZN(n44398) );
  INV_X1 U51997 ( .I(n44401), .ZN(n44402) );
  NAND2_X1 U51999 ( .A1(n49013), .A2(n64823), .ZN(n44408) );
  XOR2_X1 U52000 ( .A1(n44613), .A2(n56949), .Z(n44411) );
  XOR2_X1 U52001 ( .A1(n44412), .A2(n44411), .Z(n44413) );
  XOR2_X1 U52002 ( .A1(n44414), .A2(n44413), .Z(n44416) );
  XOR2_X1 U52003 ( .A1(n44416), .A2(n44415), .Z(n44417) );
  XOR2_X1 U52004 ( .A1(n44424), .A2(n61737), .Z(n44425) );
  XOR2_X1 U52005 ( .A1(n44426), .A2(n44425), .Z(n44428) );
  XOR2_X1 U52006 ( .A1(n44428), .A2(n44427), .Z(n44429) );
  XOR2_X1 U52007 ( .A1(n44430), .A2(n44429), .Z(n44431) );
  INV_X1 U52009 ( .I(n44436), .ZN(n44439) );
  XOR2_X1 U52010 ( .A1(n44437), .A2(n56692), .Z(n44438) );
  XOR2_X1 U52011 ( .A1(n44439), .A2(n44438), .Z(n44440) );
  XOR2_X1 U52012 ( .A1(n45875), .A2(n44440), .Z(n44441) );
  XOR2_X1 U52013 ( .A1(n44442), .A2(n22923), .Z(n44964) );
  INV_X1 U52014 ( .I(n44443), .ZN(n44444) );
  XOR2_X1 U52015 ( .A1(n44444), .A2(n53246), .Z(n44445) );
  XOR2_X1 U52016 ( .A1(n44446), .A2(n44445), .Z(n44447) );
  INV_X1 U52019 ( .I(n44483), .ZN(n44484) );
  INV_X1 U52020 ( .I(n44451), .ZN(n44452) );
  INV_X1 U52021 ( .I(n44453), .ZN(n44454) );
  AOI21_X1 U52022 ( .A1(n44457), .A2(n44456), .B(n54587), .ZN(n44458) );
  NOR2_X1 U52023 ( .A1(n44459), .A2(n44458), .ZN(n44460) );
  XOR2_X1 U52024 ( .A1(n44462), .A2(n44461), .Z(n44463) );
  XOR2_X1 U52026 ( .A1(n44467), .A2(n56180), .Z(n44468) );
  XOR2_X1 U52027 ( .A1(n50746), .A2(n44468), .Z(n44469) );
  XOR2_X1 U52028 ( .A1(n44469), .A2(n52327), .Z(n44472) );
  INV_X1 U52029 ( .I(n44470), .ZN(n44471) );
  XOR2_X1 U52030 ( .A1(n44472), .A2(n44471), .Z(n44473) );
  XOR2_X1 U52031 ( .A1(n46688), .A2(n44473), .Z(n44474) );
  XOR2_X1 U52032 ( .A1(n44475), .A2(n44474), .Z(n44476) );
  XOR2_X1 U52033 ( .A1(n44476), .A2(n44980), .Z(n44477) );
  XOR2_X1 U52034 ( .A1(n44478), .A2(n24030), .Z(n44849) );
  NAND2_X1 U52036 ( .A1(n21793), .A2(n59707), .ZN(n44486) );
  INV_X1 U52037 ( .I(n46122), .ZN(n44488) );
  INV_X1 U52038 ( .I(n44489), .ZN(n44491) );
  XOR2_X1 U52039 ( .A1(n44491), .A2(n44490), .Z(n44492) );
  XOR2_X1 U52040 ( .A1(n23905), .A2(n44492), .Z(n44493) );
  XOR2_X1 U52041 ( .A1(n44494), .A2(n44493), .Z(n44495) );
  XOR2_X1 U52042 ( .A1(n44496), .A2(n44495), .Z(n44497) );
  XOR2_X1 U52043 ( .A1(n44498), .A2(n4761), .Z(n44499) );
  XOR2_X1 U52045 ( .A1(n44502), .A2(n54185), .Z(n44503) );
  XOR2_X1 U52046 ( .A1(n12507), .A2(n44503), .Z(n44505) );
  XOR2_X1 U52047 ( .A1(n45063), .A2(n1671), .Z(n44508) );
  XOR2_X1 U52048 ( .A1(n44509), .A2(n44508), .Z(n44510) );
  XOR2_X1 U52051 ( .A1(n46615), .A2(n52226), .Z(n44512) );
  XOR2_X1 U52052 ( .A1(n44513), .A2(n44512), .Z(n44514) );
  XOR2_X1 U52053 ( .A1(n44515), .A2(n44514), .Z(n44516) );
  XOR2_X1 U52054 ( .A1(n44517), .A2(n23270), .Z(n44520) );
  XOR2_X1 U52055 ( .A1(n46535), .A2(n55516), .Z(n44629) );
  XOR2_X1 U52056 ( .A1(n44629), .A2(n46197), .Z(n44519) );
  XOR2_X1 U52058 ( .A1(n16324), .A2(n44526), .Z(n44527) );
  XOR2_X1 U52059 ( .A1(n45811), .A2(n23893), .Z(n44529) );
  INV_X1 U52060 ( .I(n44531), .ZN(n44532) );
  INV_X1 U52061 ( .I(n45487), .ZN(n44553) );
  XOR2_X1 U52062 ( .A1(n44534), .A2(n44533), .Z(n44535) );
  XOR2_X1 U52063 ( .A1(n44536), .A2(n44535), .Z(n44537) );
  XOR2_X1 U52064 ( .A1(n22650), .A2(n44537), .Z(n44538) );
  INV_X1 U52065 ( .I(n44543), .ZN(n44544) );
  XOR2_X1 U52066 ( .A1(n44544), .A2(n22821), .Z(n44545) );
  XOR2_X1 U52067 ( .A1(n44546), .A2(n44545), .Z(n44547) );
  XOR2_X1 U52068 ( .A1(n46598), .A2(n44547), .Z(n44548) );
  MUX2_X1 U52072 ( .I0(n44557), .I1(n44556), .S(n20426), .Z(n47779) );
  INV_X1 U52074 ( .I(n46949), .ZN(n44560) );
  OAI22_X1 U52076 ( .A1(n46958), .A2(n1328), .B1(n6786), .B2(n46950), .ZN(
        n44564) );
  OAI21_X1 U52078 ( .A1(n48341), .A2(n14314), .B(n44663), .ZN(n44662) );
  AOI21_X1 U52080 ( .A1(n44702), .A2(n44572), .B(n25066), .ZN(n44573) );
  NAND2_X1 U52081 ( .A1(n44706), .A2(n44577), .ZN(n44711) );
  INV_X1 U52082 ( .I(n45785), .ZN(n44575) );
  NOR2_X1 U52083 ( .A1(n44575), .A2(n45530), .ZN(n44576) );
  XOR2_X1 U52084 ( .A1(n44579), .A2(n55242), .Z(n44581) );
  INV_X1 U52085 ( .I(n51133), .ZN(n44580) );
  XOR2_X1 U52086 ( .A1(n44581), .A2(n44580), .Z(n44582) );
  XOR2_X1 U52087 ( .A1(n23267), .A2(n44582), .Z(n44583) );
  INV_X1 U52088 ( .I(n44588), .ZN(n44590) );
  XOR2_X1 U52089 ( .A1(n44590), .A2(n44589), .Z(n44591) );
  XOR2_X1 U52090 ( .A1(n44592), .A2(n44591), .Z(n44593) );
  XOR2_X1 U52091 ( .A1(n45019), .A2(n44594), .Z(n44595) );
  XOR2_X1 U52092 ( .A1(n44595), .A2(n22923), .Z(n44597) );
  INV_X1 U52093 ( .I(n44598), .ZN(n44601) );
  XOR2_X1 U52094 ( .A1(n44599), .A2(n54143), .Z(n44600) );
  XOR2_X1 U52095 ( .A1(n44601), .A2(n44600), .Z(n44603) );
  XOR2_X1 U52096 ( .A1(n44603), .A2(n44602), .Z(n44604) );
  INV_X1 U52097 ( .I(n44607), .ZN(n44610) );
  XOR2_X1 U52098 ( .A1(n23641), .A2(n44608), .Z(n46133) );
  INV_X1 U52099 ( .I(n46133), .ZN(n44609) );
  XOR2_X1 U52100 ( .A1(n44613), .A2(n55150), .Z(n44614) );
  XOR2_X1 U52101 ( .A1(n44615), .A2(n44614), .Z(n44616) );
  XOR2_X1 U52102 ( .A1(n44617), .A2(n44616), .Z(n44618) );
  XOR2_X1 U52103 ( .A1(n44619), .A2(n49434), .Z(n44620) );
  XOR2_X1 U52104 ( .A1(n44621), .A2(n44620), .Z(n44623) );
  XOR2_X1 U52105 ( .A1(n44623), .A2(n44622), .Z(n44624) );
  XOR2_X1 U52106 ( .A1(n19985), .A2(n44624), .Z(n44625) );
  XOR2_X1 U52108 ( .A1(n44911), .A2(n46197), .Z(n44628) );
  XOR2_X1 U52110 ( .A1(n44629), .A2(n65022), .Z(n46624) );
  XOR2_X1 U52111 ( .A1(n46624), .A2(n44630), .Z(n44638) );
  XOR2_X1 U52112 ( .A1(n44632), .A2(n44631), .Z(n44633) );
  XOR2_X1 U52113 ( .A1(n44634), .A2(n44633), .Z(n44635) );
  XOR2_X1 U52114 ( .A1(n24055), .A2(n44635), .Z(n44636) );
  INV_X1 U52115 ( .I(n22376), .ZN(n44640) );
  XOR2_X1 U52116 ( .A1(n44919), .A2(n18726), .Z(n44641) );
  XOR2_X1 U52117 ( .A1(n46451), .A2(n44641), .Z(n44642) );
  NOR2_X1 U52118 ( .A1(n59861), .A2(n44645), .ZN(n44646) );
  NAND2_X1 U52119 ( .A1(n22852), .A2(n47985), .ZN(n44649) );
  NAND2_X1 U52122 ( .A1(n19715), .A2(n15697), .ZN(n44652) );
  NOR2_X1 U52124 ( .A1(n44663), .A2(n25812), .ZN(n44666) );
  INV_X1 U52125 ( .I(n48737), .ZN(n44665) );
  NAND2_X1 U52127 ( .A1(n44663), .A2(n19243), .ZN(n44664) );
  INV_X1 U52128 ( .I(n48734), .ZN(n44667) );
  INV_X1 U52129 ( .I(n49914), .ZN(n44669) );
  INV_X1 U52130 ( .I(n45479), .ZN(n47513) );
  AOI21_X1 U52131 ( .A1(n47495), .A2(n12850), .B(n16493), .ZN(n44672) );
  OAI22_X1 U52132 ( .A1(n44674), .A2(n12687), .B1(n44672), .B2(n47494), .ZN(
        n44675) );
  NAND2_X1 U52133 ( .A1(n8152), .A2(n65224), .ZN(n44679) );
  MUX2_X1 U52135 ( .I0(n44679), .I1(n44678), .S(n46979), .Z(n44690) );
  NOR2_X1 U52136 ( .A1(n58174), .A2(n1660), .ZN(n44681) );
  NOR2_X1 U52141 ( .A1(n44684), .A2(n44065), .ZN(n44686) );
  NAND2_X2 U52142 ( .A1(n44690), .A2(n44689), .ZN(n49281) );
  AOI21_X1 U52145 ( .A1(n57194), .A2(n19107), .B(n22457), .ZN(n44787) );
  INV_X1 U52148 ( .I(n44703), .ZN(n44709) );
  NAND2_X1 U52149 ( .A1(n45532), .A2(n21755), .ZN(n45539) );
  NAND2_X1 U52150 ( .A1(n45539), .A2(n44706), .ZN(n44707) );
  OAI22_X1 U52151 ( .A1(n44709), .A2(n45536), .B1(n44708), .B2(n44707), .ZN(
        n44713) );
  INV_X1 U52152 ( .I(n45529), .ZN(n44710) );
  INV_X1 U52154 ( .I(n44714), .ZN(n44717) );
  INV_X1 U52155 ( .I(n44715), .ZN(n44716) );
  XOR2_X1 U52156 ( .A1(n44717), .A2(n44716), .Z(n44719) );
  XOR2_X1 U52157 ( .A1(n44719), .A2(n44718), .Z(n44720) );
  XOR2_X1 U52158 ( .A1(n7544), .A2(n44720), .Z(n44721) );
  XOR2_X1 U52159 ( .A1(n44722), .A2(n44721), .Z(n44724) );
  XOR2_X1 U52160 ( .A1(n44724), .A2(n46383), .Z(n44725) );
  XOR2_X1 U52161 ( .A1(n46120), .A2(n44725), .Z(n44726) );
  XOR2_X1 U52162 ( .A1(n44728), .A2(n44727), .Z(n44729) );
  XOR2_X1 U52163 ( .A1(n44739), .A2(n52196), .Z(n44740) );
  XOR2_X1 U52164 ( .A1(n44741), .A2(n44740), .Z(n44742) );
  INV_X1 U52165 ( .I(n49957), .ZN(n44745) );
  INV_X1 U52166 ( .I(n44747), .ZN(n44748) );
  XOR2_X1 U52167 ( .A1(n44749), .A2(n51492), .Z(n44750) );
  XOR2_X1 U52168 ( .A1(n44751), .A2(n44750), .Z(n44752) );
  XOR2_X1 U52169 ( .A1(n46188), .A2(n44753), .Z(n44755) );
  INV_X1 U52171 ( .I(n44758), .ZN(n44763) );
  XOR2_X1 U52172 ( .A1(n44759), .A2(n56784), .Z(n44760) );
  XOR2_X1 U52173 ( .A1(n44761), .A2(n44760), .Z(n44762) );
  XOR2_X1 U52174 ( .A1(n44763), .A2(n44762), .Z(n44764) );
  XOR2_X1 U52175 ( .A1(n8021), .A2(n44764), .Z(n44766) );
  XOR2_X1 U52176 ( .A1(n5011), .A2(n44766), .Z(n44767) );
  XOR2_X1 U52177 ( .A1(n44768), .A2(n44767), .Z(n44769) );
  INV_X1 U52178 ( .I(n44773), .ZN(n44777) );
  NAND4_X1 U52180 ( .A1(n45766), .A2(n46913), .A3(n23480), .A4(n44780), .ZN(
        n44783) );
  AOI21_X1 U52181 ( .A1(n45766), .A2(n15666), .B(n44781), .ZN(n44782) );
  OAI21_X1 U52183 ( .A1(n44787), .A2(n48923), .B(n49288), .ZN(n44792) );
  NAND2_X1 U52184 ( .A1(n57194), .A2(n49276), .ZN(n44789) );
  NAND2_X1 U52185 ( .A1(n48931), .A2(n64488), .ZN(n44795) );
  XOR2_X1 U52186 ( .A1(n44797), .A2(n44796), .Z(n44798) );
  XOR2_X1 U52187 ( .A1(n51968), .A2(n44803), .Z(n44804) );
  XOR2_X1 U52188 ( .A1(n44808), .A2(n53805), .Z(n44811) );
  INV_X1 U52189 ( .I(n44809), .ZN(n44810) );
  XOR2_X1 U52190 ( .A1(n44811), .A2(n44810), .Z(n44813) );
  XOR2_X1 U52191 ( .A1(n44813), .A2(n44812), .Z(n44814) );
  XOR2_X1 U52192 ( .A1(n23210), .A2(n44814), .Z(n44815) );
  XOR2_X1 U52193 ( .A1(n44815), .A2(n23722), .Z(n44816) );
  INV_X1 U52194 ( .I(n44822), .ZN(n44824) );
  XOR2_X1 U52195 ( .A1(n51193), .A2(n54776), .Z(n44823) );
  XOR2_X1 U52196 ( .A1(n44824), .A2(n44823), .Z(n44825) );
  XOR2_X1 U52197 ( .A1(n44826), .A2(n44825), .Z(n44827) );
  XOR2_X1 U52198 ( .A1(n46272), .A2(n44827), .Z(n44828) );
  XOR2_X1 U52199 ( .A1(n59218), .A2(n46164), .Z(n44837) );
  INV_X1 U52200 ( .I(n44830), .ZN(n44832) );
  XOR2_X1 U52201 ( .A1(n44832), .A2(n44831), .Z(n44833) );
  XOR2_X1 U52202 ( .A1(n58027), .A2(n44833), .Z(n44835) );
  XOR2_X1 U52203 ( .A1(n46621), .A2(n44835), .Z(n44836) );
  XOR2_X1 U52204 ( .A1(n44836), .A2(n44837), .Z(n44838) );
  NOR2_X1 U52206 ( .A1(n47570), .A2(n47900), .ZN(n44860) );
  XOR2_X1 U52208 ( .A1(n44841), .A2(n27640), .Z(n44842) );
  XOR2_X1 U52209 ( .A1(n44843), .A2(n44842), .Z(n44845) );
  XOR2_X1 U52210 ( .A1(n44845), .A2(n44844), .Z(n44846) );
  XOR2_X1 U52211 ( .A1(n44847), .A2(n44846), .Z(n44848) );
  INV_X1 U52212 ( .I(n44850), .ZN(n44852) );
  XOR2_X1 U52213 ( .A1(n44852), .A2(n60918), .Z(n44853) );
  XOR2_X1 U52214 ( .A1(n44853), .A2(n23893), .Z(n44854) );
  AOI21_X1 U52217 ( .A1(n47905), .A2(n45592), .B(n45594), .ZN(n44862) );
  NOR2_X2 U52218 ( .A1(n44866), .A2(n44865), .ZN(n48883) );
  INV_X2 U52220 ( .I(n44868), .ZN(n46893) );
  NAND2_X1 U52221 ( .A1(n46893), .A2(n47259), .ZN(n44871) );
  OAI21_X1 U52223 ( .A1(n21976), .A2(n9730), .B(n46891), .ZN(n44874) );
  INV_X1 U52226 ( .I(n44876), .ZN(n44879) );
  XOR2_X1 U52227 ( .A1(n44877), .A2(n53764), .Z(n44878) );
  XOR2_X1 U52228 ( .A1(n44879), .A2(n44878), .Z(n44880) );
  XOR2_X1 U52230 ( .A1(n22551), .A2(n10713), .Z(n44883) );
  XOR2_X1 U52231 ( .A1(n44887), .A2(n54143), .Z(n44890) );
  INV_X1 U52232 ( .I(n44888), .ZN(n44889) );
  XOR2_X1 U52233 ( .A1(n44890), .A2(n44889), .Z(n44891) );
  XOR2_X1 U52234 ( .A1(n65177), .A2(n64610), .Z(n44894) );
  XOR2_X1 U52235 ( .A1(n49434), .A2(n56784), .Z(n44899) );
  XOR2_X1 U52236 ( .A1(n52614), .A2(n44899), .Z(n44900) );
  XOR2_X1 U52237 ( .A1(n44900), .A2(n52449), .Z(n44901) );
  XOR2_X1 U52238 ( .A1(n44901), .A2(n46688), .Z(n44902) );
  XOR2_X1 U52239 ( .A1(n44902), .A2(n23893), .Z(n44903) );
  XOR2_X1 U52240 ( .A1(n65022), .A2(n44911), .Z(n44918) );
  XOR2_X1 U52241 ( .A1(n44913), .A2(n46437), .Z(n44915) );
  XOR2_X1 U52242 ( .A1(n44915), .A2(n44914), .Z(n44916) );
  XOR2_X1 U52243 ( .A1(n23872), .A2(n44916), .Z(n44917) );
  XOR2_X1 U52244 ( .A1(n44924), .A2(n51814), .Z(n44926) );
  XOR2_X1 U52245 ( .A1(n44926), .A2(n44925), .Z(n44928) );
  XOR2_X1 U52246 ( .A1(n44928), .A2(n44927), .Z(n44929) );
  XOR2_X1 U52247 ( .A1(n23953), .A2(n44929), .Z(n44930) );
  INV_X1 U52248 ( .I(n44932), .ZN(n44936) );
  INV_X1 U52249 ( .I(n44933), .ZN(n44934) );
  XOR2_X1 U52250 ( .A1(n44934), .A2(n55610), .Z(n44935) );
  XOR2_X1 U52251 ( .A1(n44936), .A2(n44935), .Z(n44937) );
  NAND2_X1 U52256 ( .A1(n44942), .A2(n45932), .ZN(n44946) );
  NAND2_X1 U52258 ( .A1(n47302), .A2(n46025), .ZN(n44945) );
  INV_X1 U52259 ( .I(n44949), .ZN(n44951) );
  XOR2_X1 U52260 ( .A1(n44951), .A2(n44950), .Z(n44952) );
  XOR2_X1 U52261 ( .A1(n23953), .A2(n44952), .Z(n44953) );
  XOR2_X1 U52263 ( .A1(n17301), .A2(n55610), .Z(n44959) );
  XOR2_X1 U52264 ( .A1(n44960), .A2(n53805), .Z(n44961) );
  XOR2_X1 U52265 ( .A1(n44962), .A2(n44961), .Z(n44963) );
  XOR2_X1 U52266 ( .A1(n15354), .A2(n55765), .Z(n45070) );
  XOR2_X1 U52267 ( .A1(n22439), .A2(n44967), .Z(n44968) );
  XOR2_X1 U52268 ( .A1(n50772), .A2(n44971), .Z(n44972) );
  XOR2_X1 U52269 ( .A1(n44973), .A2(n44972), .Z(n44974) );
  XOR2_X1 U52270 ( .A1(n44978), .A2(n10552), .Z(n44979) );
  INV_X1 U52271 ( .I(n44981), .ZN(n44986) );
  XOR2_X1 U52272 ( .A1(n15712), .A2(n53344), .Z(n44982) );
  XOR2_X1 U52273 ( .A1(n51234), .A2(n44982), .Z(n44984) );
  XOR2_X1 U52274 ( .A1(n44984), .A2(n44983), .Z(n44985) );
  XOR2_X1 U52275 ( .A1(n44986), .A2(n44985), .Z(n44987) );
  XOR2_X1 U52276 ( .A1(n24030), .A2(n44987), .Z(n44988) );
  XOR2_X1 U52277 ( .A1(n44988), .A2(n45823), .Z(n44989) );
  XOR2_X1 U52278 ( .A1(n44992), .A2(n61010), .Z(n46159) );
  XOR2_X1 U52279 ( .A1(n50832), .A2(n44995), .Z(n44997) );
  XOR2_X1 U52280 ( .A1(n44997), .A2(n44996), .Z(n44998) );
  XOR2_X1 U52281 ( .A1(n44999), .A2(n44998), .Z(n45000) );
  XOR2_X1 U52282 ( .A1(n22376), .A2(n45000), .Z(n45001) );
  XOR2_X1 U52283 ( .A1(n45001), .A2(n46164), .Z(n45002) );
  NAND2_X1 U52285 ( .A1(n47244), .A2(n45988), .ZN(n47618) );
  NOR2_X1 U52286 ( .A1(n45990), .A2(n15360), .ZN(n45007) );
  INV_X1 U52287 ( .I(n47239), .ZN(n45006) );
  NOR2_X1 U52288 ( .A1(n45008), .A2(n47244), .ZN(n45009) );
  OAI21_X1 U52289 ( .A1(n45206), .A2(n45009), .B(n58155), .ZN(n45010) );
  INV_X1 U52290 ( .I(n50070), .ZN(n45012) );
  XOR2_X1 U52291 ( .A1(n45011), .A2(n45012), .Z(n45013) );
  XOR2_X1 U52292 ( .A1(n46493), .A2(n45013), .Z(n45014) );
  XOR2_X1 U52293 ( .A1(n46550), .A2(n23078), .Z(n45020) );
  XOR2_X1 U52294 ( .A1(n46385), .A2(n45020), .Z(n45022) );
  INV_X1 U52295 ( .I(n45025), .ZN(n45028) );
  XOR2_X1 U52296 ( .A1(n45026), .A2(n45878), .Z(n45027) );
  XOR2_X1 U52297 ( .A1(n45028), .A2(n45027), .Z(n45029) );
  XOR2_X1 U52298 ( .A1(n23210), .A2(n45029), .Z(n45031) );
  XOR2_X1 U52299 ( .A1(n46553), .A2(n45032), .Z(n45033) );
  XOR2_X1 U52301 ( .A1(n45036), .A2(n52327), .Z(n45038) );
  XOR2_X1 U52302 ( .A1(n45038), .A2(n45037), .Z(n45039) );
  XOR2_X1 U52303 ( .A1(n45040), .A2(n45039), .Z(n45042) );
  XOR2_X1 U52304 ( .A1(n45042), .A2(n24062), .Z(n45043) );
  XOR2_X1 U52305 ( .A1(n45049), .A2(n45048), .Z(n45050) );
  XOR2_X1 U52306 ( .A1(n63789), .A2(n45050), .Z(n45051) );
  XOR2_X1 U52308 ( .A1(n45059), .A2(n52350), .Z(n45060) );
  XOR2_X1 U52309 ( .A1(n45061), .A2(n45060), .Z(n45062) );
  XOR2_X1 U52310 ( .A1(n45064), .A2(n22821), .Z(n45065) );
  XOR2_X1 U52311 ( .A1(n45131), .A2(n45065), .Z(n45066) );
  XOR2_X1 U52312 ( .A1(n45067), .A2(n45066), .Z(n45068) );
  XOR2_X1 U52313 ( .A1(n12178), .A2(n45068), .Z(n45069) );
  NAND2_X1 U52315 ( .A1(n45958), .A2(n47328), .ZN(n45079) );
  NAND3_X1 U52316 ( .A1(n46066), .A2(n47310), .A3(n47312), .ZN(n45078) );
  NAND2_X1 U52317 ( .A1(n59670), .A2(n47329), .ZN(n45081) );
  INV_X1 U52318 ( .I(n47310), .ZN(n46921) );
  NAND3_X1 U52319 ( .A1(n45081), .A2(n46921), .A3(n45080), .ZN(n45082) );
  XOR2_X1 U52320 ( .A1(n64837), .A2(n45085), .Z(n45086) );
  XOR2_X1 U52321 ( .A1(n45087), .A2(n56901), .Z(n45089) );
  XOR2_X1 U52322 ( .A1(n45089), .A2(n45088), .Z(n45090) );
  XOR2_X1 U52323 ( .A1(n45091), .A2(n45090), .Z(n45092) );
  XOR2_X1 U52324 ( .A1(n23264), .A2(n45092), .Z(n45094) );
  XOR2_X1 U52325 ( .A1(n10255), .A2(n23722), .Z(n45097) );
  XOR2_X1 U52326 ( .A1(n1676), .A2(n45097), .Z(n45098) );
  XOR2_X1 U52327 ( .A1(n45101), .A2(n51019), .Z(n45102) );
  XOR2_X1 U52328 ( .A1(n45103), .A2(n45102), .Z(n45104) );
  XOR2_X1 U52329 ( .A1(n45105), .A2(n45104), .Z(n45106) );
  INV_X1 U52332 ( .I(n45112), .ZN(n45113) );
  XOR2_X1 U52333 ( .A1(n45113), .A2(n57131), .Z(n45114) );
  XOR2_X1 U52334 ( .A1(n24030), .A2(n45116), .Z(n45117) );
  XOR2_X1 U52336 ( .A1(n45121), .A2(n53764), .Z(n45122) );
  XOR2_X1 U52337 ( .A1(n45122), .A2(n30402), .Z(n45124) );
  XOR2_X1 U52338 ( .A1(n45124), .A2(n45123), .Z(n45125) );
  XOR2_X1 U52339 ( .A1(n45126), .A2(n45125), .Z(n45127) );
  INV_X1 U52340 ( .I(n45130), .ZN(n45132) );
  XOR2_X1 U52341 ( .A1(n45132), .A2(n45131), .Z(n45133) );
  XOR2_X1 U52342 ( .A1(n45134), .A2(n45133), .Z(n45135) );
  XOR2_X1 U52343 ( .A1(n64373), .A2(n45135), .Z(n45137) );
  XOR2_X1 U52344 ( .A1(n45137), .A2(n45136), .Z(n45138) );
  INV_X1 U52345 ( .I(n45141), .ZN(n45142) );
  XOR2_X1 U52346 ( .A1(n45143), .A2(n45142), .Z(n45144) );
  XOR2_X1 U52347 ( .A1(n45145), .A2(n45144), .Z(n45146) );
  XOR2_X1 U52348 ( .A1(n45146), .A2(n22639), .Z(n45148) );
  XOR2_X1 U52349 ( .A1(n45148), .A2(n45147), .Z(n45149) );
  XOR2_X1 U52350 ( .A1(n45149), .A2(n46440), .Z(n45150) );
  XOR2_X1 U52351 ( .A1(n45151), .A2(n45150), .Z(n45152) );
  NAND2_X1 U52352 ( .A1(n45682), .A2(n14888), .ZN(n45153) );
  NAND2_X1 U52353 ( .A1(n45154), .A2(n47592), .ZN(n45158) );
  NOR2_X1 U52355 ( .A1(n47280), .A2(n47281), .ZN(n45156) );
  AOI22_X1 U52356 ( .A1(n45156), .A2(n47590), .B1(n45155), .B2(n47580), .ZN(
        n45157) );
  NAND2_X1 U52358 ( .A1(n15737), .A2(n22157), .ZN(n45162) );
  NAND2_X1 U52361 ( .A1(n49697), .A2(n48894), .ZN(n49755) );
  NOR3_X1 U52362 ( .A1(n9863), .A2(n24049), .A3(n45171), .ZN(n45175) );
  NOR2_X1 U52363 ( .A1(n48883), .A2(n48349), .ZN(n49703) );
  INV_X1 U52364 ( .I(n49703), .ZN(n49761) );
  NAND4_X1 U52365 ( .A1(n45172), .A2(n9863), .A3(n22157), .A4(n49698), .ZN(
        n45173) );
  OAI21_X1 U52366 ( .A1(n49761), .A2(n48885), .B(n45173), .ZN(n45174) );
  NAND2_X1 U52372 ( .A1(n47885), .A2(n14121), .ZN(n45184) );
  OAI22_X1 U52373 ( .A1(n45184), .A2(n61510), .B1(n47879), .B2(n47721), .ZN(
        n45186) );
  NOR2_X1 U52374 ( .A1(n47896), .A2(n47900), .ZN(n45195) );
  NAND2_X1 U52375 ( .A1(n23969), .A2(n47900), .ZN(n45192) );
  NOR2_X1 U52376 ( .A1(n47902), .A2(n47901), .ZN(n45946) );
  NAND2_X1 U52377 ( .A1(n47894), .A2(n47572), .ZN(n45194) );
  INV_X1 U52378 ( .I(n47385), .ZN(n45197) );
  NAND2_X1 U52379 ( .A1(n47803), .A2(n25895), .ZN(n45196) );
  INV_X1 U52380 ( .I(n47706), .ZN(n45198) );
  NAND3_X1 U52381 ( .A1(n47699), .A2(n25841), .A3(n8048), .ZN(n45200) );
  AOI21_X1 U52382 ( .A1(n62739), .A2(n47622), .B(n45204), .ZN(n45205) );
  NOR2_X1 U52383 ( .A1(n45207), .A2(n47621), .ZN(n45210) );
  NOR2_X1 U52384 ( .A1(n45208), .A2(n64470), .ZN(n45209) );
  OAI21_X1 U52385 ( .A1(n10420), .A2(n60881), .B(n47845), .ZN(n45214) );
  NAND2_X1 U52386 ( .A1(n10420), .A2(n62952), .ZN(n45212) );
  OAI22_X1 U52387 ( .A1(n2641), .A2(n45212), .B1(n47828), .B2(n24114), .ZN(
        n45213) );
  AOI21_X1 U52388 ( .A1(n45215), .A2(n45214), .B(n45213), .ZN(n45221) );
  OAI21_X1 U52390 ( .A1(n47828), .A2(n62952), .B(n24114), .ZN(n45216) );
  NAND2_X1 U52392 ( .A1(n47655), .A2(n62424), .ZN(n45219) );
  NOR3_X1 U52394 ( .A1(n45223), .A2(n45225), .A3(n47817), .ZN(n45224) );
  NAND2_X1 U52395 ( .A1(n47610), .A2(n59629), .ZN(n45226) );
  NOR2_X1 U52398 ( .A1(n49222), .A2(n1205), .ZN(n49158) );
  XOR2_X1 U52399 ( .A1(n55060), .A2(n55610), .Z(n49401) );
  XOR2_X1 U52400 ( .A1(n51999), .A2(n49401), .Z(n45239) );
  XOR2_X1 U52401 ( .A1(n45239), .A2(n45238), .Z(n45241) );
  XOR2_X1 U52402 ( .A1(n45241), .A2(n45240), .Z(n45242) );
  XOR2_X1 U52403 ( .A1(n45243), .A2(n45242), .Z(n45244) );
  XOR2_X1 U52404 ( .A1(n23402), .A2(n45244), .Z(n45245) );
  XOR2_X1 U52405 ( .A1(n45246), .A2(n7544), .Z(n45247) );
  INV_X1 U52407 ( .I(n45250), .ZN(n45252) );
  XOR2_X1 U52408 ( .A1(n45252), .A2(n45251), .Z(n45253) );
  INV_X1 U52409 ( .I(n45255), .ZN(n45256) );
  XOR2_X1 U52410 ( .A1(n45257), .A2(n45256), .Z(n45258) );
  XOR2_X1 U52411 ( .A1(n23426), .A2(n45258), .Z(n45259) );
  XOR2_X1 U52412 ( .A1(n46312), .A2(n45259), .Z(n45260) );
  XOR2_X1 U52413 ( .A1(n45261), .A2(n20900), .Z(n45262) );
  XOR2_X1 U52414 ( .A1(n45262), .A2(n45263), .Z(n45264) );
  XOR2_X1 U52418 ( .A1(n23553), .A2(n61457), .Z(n45270) );
  XOR2_X1 U52420 ( .A1(n22961), .A2(n17129), .Z(n50585) );
  XOR2_X1 U52421 ( .A1(n50585), .A2(n45275), .Z(n45277) );
  XOR2_X1 U52422 ( .A1(n45276), .A2(n55624), .Z(n50748) );
  XOR2_X1 U52423 ( .A1(n45277), .A2(n50748), .Z(n45279) );
  XOR2_X1 U52424 ( .A1(n45279), .A2(n45278), .Z(n45280) );
  XOR2_X1 U52425 ( .A1(n12002), .A2(n10713), .Z(n45291) );
  XOR2_X1 U52426 ( .A1(n45286), .A2(n55379), .Z(n45287) );
  XOR2_X1 U52427 ( .A1(n45288), .A2(n45287), .Z(n45289) );
  XOR2_X1 U52428 ( .A1(n4990), .A2(n45289), .Z(n45290) );
  XOR2_X1 U52430 ( .A1(n51608), .A2(n56849), .Z(n45294) );
  XOR2_X1 U52431 ( .A1(n45295), .A2(n45294), .Z(n45296) );
  XOR2_X1 U52432 ( .A1(n11515), .A2(n45297), .Z(n45298) );
  NAND2_X1 U52433 ( .A1(n61720), .A2(n45267), .ZN(n45301) );
  OAI21_X1 U52434 ( .A1(n1263), .A2(n59528), .B(n1649), .ZN(n45302) );
  BUF_X4 U52435 ( .I(n45304), .Z(n50426) );
  NAND2_X1 U52437 ( .A1(n47797), .A2(n25896), .ZN(n45308) );
  NOR2_X1 U52440 ( .A1(n47386), .A2(n25895), .ZN(n47391) );
  NOR2_X1 U52441 ( .A1(n14323), .A2(n47699), .ZN(n45311) );
  OAI21_X1 U52442 ( .A1(n47391), .A2(n45311), .B(n1385), .ZN(n45312) );
  INV_X1 U52443 ( .I(n45314), .ZN(n45315) );
  INV_X1 U52444 ( .I(n45321), .ZN(n45323) );
  XOR2_X1 U52445 ( .A1(n45323), .A2(n45322), .Z(n45324) );
  XOR2_X1 U52446 ( .A1(n23426), .A2(n23059), .Z(n45327) );
  XOR2_X1 U52447 ( .A1(n45328), .A2(n51493), .Z(n45329) );
  XOR2_X1 U52448 ( .A1(n45330), .A2(n45329), .Z(n45331) );
  XOR2_X1 U52449 ( .A1(n46442), .A2(n45331), .Z(n45332) );
  XOR2_X1 U52450 ( .A1(n45332), .A2(n46164), .Z(n45334) );
  XOR2_X1 U52451 ( .A1(n45333), .A2(n45334), .Z(n45335) );
  XOR2_X1 U52452 ( .A1(n45425), .A2(n45335), .Z(n45336) );
  INV_X1 U52453 ( .I(n45337), .ZN(n45340) );
  XOR2_X1 U52454 ( .A1(n45338), .A2(n50475), .Z(n45339) );
  INV_X1 U52455 ( .I(n64443), .ZN(n45344) );
  XOR2_X1 U52456 ( .A1(n23687), .A2(n45344), .Z(n45345) );
  XOR2_X1 U52457 ( .A1(n63745), .A2(n45345), .Z(n45346) );
  INV_X1 U52458 ( .I(n45347), .ZN(n45352) );
  XOR2_X1 U52459 ( .A1(n45350), .A2(n45349), .Z(n45351) );
  XOR2_X1 U52460 ( .A1(n1331), .A2(n45353), .Z(n45354) );
  XOR2_X1 U52461 ( .A1(n5989), .A2(n45354), .Z(n45355) );
  XOR2_X1 U52462 ( .A1(n45360), .A2(n45359), .Z(n45363) );
  XOR2_X1 U52463 ( .A1(n50745), .A2(n58084), .Z(n45361) );
  XOR2_X1 U52464 ( .A1(n46683), .A2(n45361), .Z(n45362) );
  XOR2_X1 U52465 ( .A1(n45363), .A2(n45362), .Z(n45364) );
  INV_X1 U52466 ( .I(n45370), .ZN(n45372) );
  INV_X1 U52467 ( .I(n45378), .ZN(n45382) );
  XOR2_X1 U52468 ( .A1(n45380), .A2(n45379), .Z(n45381) );
  XOR2_X1 U52469 ( .A1(n45382), .A2(n45381), .Z(n45383) );
  XOR2_X1 U52470 ( .A1(n45388), .A2(n55150), .Z(n45390) );
  XOR2_X1 U52471 ( .A1(n45390), .A2(n45389), .Z(n45391) );
  XOR2_X1 U52472 ( .A1(n46522), .A2(n45391), .Z(n45392) );
  XOR2_X1 U52473 ( .A1(n45395), .A2(n620), .Z(n51768) );
  XOR2_X1 U52474 ( .A1(n51768), .A2(n45396), .Z(n45397) );
  XOR2_X1 U52475 ( .A1(n19232), .A2(n45397), .Z(n45398) );
  AOI21_X1 U52476 ( .A1(n15825), .A2(n65161), .B(n47144), .ZN(n45413) );
  INV_X1 U52477 ( .I(n45403), .ZN(n45407) );
  XOR2_X1 U52478 ( .A1(n45405), .A2(n45404), .Z(n45406) );
  XOR2_X1 U52479 ( .A1(n45407), .A2(n45406), .Z(n45408) );
  AOI21_X1 U52480 ( .A1(n45413), .A2(n45809), .B(n47140), .ZN(n45434) );
  NAND4_X1 U52481 ( .A1(n10172), .A2(n10475), .A3(n45437), .A4(n22736), .ZN(
        n45414) );
  INV_X1 U52483 ( .I(n45416), .ZN(n45420) );
  XOR2_X1 U52484 ( .A1(n45418), .A2(n45417), .Z(n45419) );
  XOR2_X1 U52485 ( .A1(n45420), .A2(n45419), .Z(n45421) );
  XOR2_X1 U52486 ( .A1(n23059), .A2(n45421), .Z(n45422) );
  XOR2_X1 U52487 ( .A1(n45423), .A2(n45422), .Z(n45424) );
  XOR2_X1 U52488 ( .A1(n46438), .A2(n20900), .Z(n45427) );
  XOR2_X1 U52489 ( .A1(n45428), .A2(n45427), .Z(n45430) );
  XOR2_X1 U52490 ( .A1(n45429), .A2(n45430), .Z(n45431) );
  NAND3_X1 U52492 ( .A1(n47372), .A2(n47377), .A3(n47367), .ZN(n45438) );
  MUX2_X1 U52494 ( .I0(n45444), .I1(n45443), .S(n50427), .Z(n45463) );
  OAI22_X1 U52495 ( .A1(n47857), .A2(n62990), .B1(n47398), .B2(n47852), .ZN(
        n45445) );
  NAND2_X1 U52496 ( .A1(n20912), .A2(n7395), .ZN(n45446) );
  NAND2_X1 U52497 ( .A1(n47868), .A2(n45905), .ZN(n45447) );
  NOR3_X1 U52498 ( .A1(n47671), .A2(n47407), .A3(n11627), .ZN(n45448) );
  NAND2_X1 U52499 ( .A1(n22700), .A2(n47728), .ZN(n45449) );
  MUX2_X1 U52501 ( .I0(n45449), .I1(n45452), .S(n47735), .Z(n45455) );
  MUX2_X1 U52502 ( .I0(n24252), .I1(n45450), .S(n47735), .Z(n45451) );
  NAND2_X1 U52503 ( .A1(n45913), .A2(n47744), .ZN(n45453) );
  AOI21_X1 U52504 ( .A1(n46739), .A2(n46736), .B(n59008), .ZN(n45456) );
  INV_X1 U52505 ( .I(n48287), .ZN(n45458) );
  NAND2_X1 U52506 ( .A1(n48757), .A2(n78), .ZN(n45457) );
  NOR2_X1 U52508 ( .A1(n23063), .A2(n2736), .ZN(n49249) );
  NOR2_X1 U52510 ( .A1(n25680), .A2(n78), .ZN(n45465) );
  NOR2_X1 U52511 ( .A1(n50427), .A2(n45464), .ZN(n49258) );
  AOI22_X1 U52512 ( .A1(n47458), .A2(n45465), .B1(n50430), .B2(n49258), .ZN(
        n45469) );
  XOR2_X1 U52514 ( .A1(n45470), .A2(n55034), .Z(n45472) );
  XOR2_X1 U52515 ( .A1(n45472), .A2(n45471), .Z(n45473) );
  XOR2_X1 U52516 ( .A1(n45474), .A2(n45473), .Z(n45475) );
  NOR2_X1 U52518 ( .A1(n45479), .A2(n47516), .ZN(n45481) );
  NAND2_X1 U52519 ( .A1(n47511), .A2(n22899), .ZN(n45480) );
  NOR2_X1 U52520 ( .A1(n65275), .A2(n45482), .ZN(n45483) );
  XOR2_X1 U52522 ( .A1(n63501), .A2(n45724), .Z(n45490) );
  NAND2_X1 U52523 ( .A1(n23759), .A2(n46033), .ZN(n45489) );
  NAND2_X1 U52524 ( .A1(n20426), .A2(n7161), .ZN(n45491) );
  NOR3_X1 U52525 ( .A1(n9988), .A2(n64888), .A3(n1666), .ZN(n45492) );
  NAND3_X1 U52527 ( .A1(n62247), .A2(n13258), .A3(n45498), .ZN(n45499) );
  NOR2_X1 U52530 ( .A1(n46949), .A2(n45505), .ZN(n45508) );
  AOI22_X1 U52532 ( .A1(n16238), .A2(n9972), .B1(n45765), .B2(n1388), .ZN(
        n45515) );
  NAND2_X1 U52533 ( .A1(n46978), .A2(n20917), .ZN(n45523) );
  NAND2_X1 U52534 ( .A1(n44065), .A2(n45521), .ZN(n45522) );
  NAND2_X1 U52535 ( .A1(n64061), .A2(n65224), .ZN(n45524) );
  OAI21_X1 U52536 ( .A1(n47020), .A2(n22905), .B(n18321), .ZN(n45528) );
  AOI21_X1 U52538 ( .A1(n20299), .A2(n1294), .B(n64274), .ZN(n45534) );
  NAND3_X1 U52539 ( .A1(n21755), .A2(n13655), .A3(n45538), .ZN(n45533) );
  NAND2_X1 U52544 ( .A1(n838), .A2(n47838), .ZN(n45549) );
  NAND2_X1 U52545 ( .A1(n45551), .A2(n47281), .ZN(n47289) );
  NOR2_X1 U52546 ( .A1(n47280), .A2(n47289), .ZN(n47591) );
  NAND2_X1 U52547 ( .A1(n47591), .A2(n45979), .ZN(n45557) );
  NAND2_X1 U52549 ( .A1(n45554), .A2(n23186), .ZN(n45555) );
  NAND2_X1 U52550 ( .A1(n47818), .A2(n47827), .ZN(n45559) );
  NAND2_X1 U52552 ( .A1(n45968), .A2(n47827), .ZN(n45562) );
  NOR2_X1 U52553 ( .A1(n1295), .A2(n23894), .ZN(n45567) );
  NAND2_X1 U52555 ( .A1(n45990), .A2(n22239), .ZN(n45572) );
  NAND2_X1 U52556 ( .A1(n45573), .A2(n45572), .ZN(n45574) );
  AOI22_X1 U52558 ( .A1(n47238), .A2(n45577), .B1(n45576), .B2(n45988), .ZN(
        n45581) );
  OAI21_X1 U52559 ( .A1(n412), .A2(n47902), .B(n47575), .ZN(n45584) );
  NAND2_X1 U52560 ( .A1(n45584), .A2(n7298), .ZN(n45588) );
  NAND2_X1 U52565 ( .A1(n47899), .A2(n1483), .ZN(n45597) );
  NAND2_X1 U52566 ( .A1(n46025), .A2(n59859), .ZN(n45599) );
  INV_X1 U52569 ( .I(n45602), .ZN(n47293) );
  AOI22_X1 U52570 ( .A1(n47293), .A2(n65095), .B1(n46013), .B2(n46025), .ZN(
        n45603) );
  NAND2_X1 U52571 ( .A1(n45609), .A2(n45608), .ZN(n48976) );
  NOR2_X1 U52572 ( .A1(n45607), .A2(n48374), .ZN(n45611) );
  NOR2_X1 U52573 ( .A1(n48058), .A2(n22756), .ZN(n45610) );
  NOR3_X1 U52574 ( .A1(n49849), .A2(n22756), .A3(n48977), .ZN(n45612) );
  NAND2_X1 U52576 ( .A1(n46923), .A2(n45957), .ZN(n45617) );
  INV_X1 U52578 ( .I(n45619), .ZN(n45954) );
  INV_X1 U52580 ( .I(n47312), .ZN(n45621) );
  NOR2_X1 U52581 ( .A1(n47308), .A2(n47329), .ZN(n45623) );
  NOR2_X1 U52582 ( .A1(n45639), .A2(n47299), .ZN(n45631) );
  NOR2_X1 U52584 ( .A1(n47296), .A2(n26180), .ZN(n45642) );
  NAND3_X1 U52585 ( .A1(n45634), .A2(n47305), .A3(n45642), .ZN(n45638) );
  NAND2_X1 U52587 ( .A1(n45635), .A2(n45932), .ZN(n45636) );
  NAND3_X1 U52589 ( .A1(n47297), .A2(n47295), .A3(n45642), .ZN(n45646) );
  INV_X1 U52590 ( .I(n1078), .ZN(n45644) );
  NAND3_X1 U52591 ( .A1(n45644), .A2(n45932), .A3(n59859), .ZN(n45645) );
  INV_X1 U52595 ( .I(n45723), .ZN(n47775) );
  INV_X1 U52597 ( .I(n46859), .ZN(n45655) );
  AOI21_X1 U52598 ( .A1(n47775), .A2(n64878), .B(n45655), .ZN(n45660) );
  NOR2_X1 U52599 ( .A1(n9988), .A2(n4569), .ZN(n45657) );
  NAND3_X1 U52600 ( .A1(n20426), .A2(n7161), .A3(n62571), .ZN(n45656) );
  OAI22_X1 U52602 ( .A1(n45657), .A2(n45656), .B1(n46038), .B2(n46864), .ZN(
        n45658) );
  NAND2_X1 U52603 ( .A1(n45658), .A2(n64849), .ZN(n45659) );
  NAND3_X2 U52604 ( .A1(n45661), .A2(n45660), .A3(n45659), .ZN(n45662) );
  NAND4_X1 U52606 ( .A1(n45675), .A2(n46882), .A3(n47251), .A4(n47256), .ZN(
        n45676) );
  NAND2_X1 U52607 ( .A1(n47590), .A2(n47281), .ZN(n45678) );
  NOR2_X1 U52608 ( .A1(n23186), .A2(n47270), .ZN(n47277) );
  NAND2_X1 U52610 ( .A1(n47270), .A2(n47592), .ZN(n45680) );
  NAND3_X1 U52612 ( .A1(n47228), .A2(n47232), .A3(n19715), .ZN(n45690) );
  NAND2_X1 U52613 ( .A1(n47233), .A2(n46946), .ZN(n45689) );
  OAI21_X1 U52614 ( .A1(n22391), .A2(n23643), .B(n46943), .ZN(n45696) );
  NAND2_X1 U52615 ( .A1(n46049), .A2(n64899), .ZN(n45694) );
  NOR2_X1 U52616 ( .A1(n48294), .A2(n21071), .ZN(n49835) );
  NAND2_X1 U52617 ( .A1(n47451), .A2(n49074), .ZN(n45699) );
  NOR2_X1 U52618 ( .A1(n49063), .A2(n65135), .ZN(n47450) );
  MUX2_X1 U52619 ( .I0(n45700), .I1(n45699), .S(n47450), .Z(n45709) );
  NOR4_X1 U52620 ( .A1(n49831), .A2(n45703), .A3(n45701), .A4(n45702), .ZN(
        n45708) );
  NOR2_X1 U52621 ( .A1(n11950), .A2(n49074), .ZN(n45704) );
  OAI21_X1 U52622 ( .A1(n45705), .A2(n49063), .B(n45704), .ZN(n45706) );
  NAND3_X1 U52623 ( .A1(n24578), .A2(n45725), .A3(n64888), .ZN(n45712) );
  NAND2_X1 U52625 ( .A1(n46026), .A2(n4569), .ZN(n45714) );
  NAND2_X1 U52626 ( .A1(n46858), .A2(n46863), .ZN(n45713) );
  NAND2_X1 U52628 ( .A1(n46026), .A2(n46875), .ZN(n45719) );
  NOR2_X1 U52629 ( .A1(n45716), .A2(n47774), .ZN(n45717) );
  NAND2_X1 U52630 ( .A1(n9988), .A2(n45717), .ZN(n46873) );
  NAND4_X1 U52631 ( .A1(n45720), .A2(n45719), .A3(n45718), .A4(n46873), .ZN(
        n45721) );
  OAI22_X1 U52633 ( .A1(n19715), .A2(n15697), .B1(n46946), .B2(n23643), .ZN(
        n45736) );
  NAND3_X1 U52634 ( .A1(n45736), .A2(n64899), .A3(n24359), .ZN(n45737) );
  INV_X1 U52638 ( .I(n46987), .ZN(n45748) );
  NAND2_X1 U52639 ( .A1(n45750), .A2(n1328), .ZN(n45754) );
  INV_X1 U52642 ( .I(n45758), .ZN(n45756) );
  NAND3_X1 U52643 ( .A1(n45756), .A2(n46948), .A3(n62490), .ZN(n45761) );
  NAND2_X1 U52644 ( .A1(n45757), .A2(n46948), .ZN(n45759) );
  NAND3_X1 U52645 ( .A1(n45759), .A2(n58705), .A3(n45758), .ZN(n45760) );
  NAND2_X1 U52646 ( .A1(n45766), .A2(n45765), .ZN(n45774) );
  AOI22_X1 U52647 ( .A1(n6081), .A2(n45774), .B1(n45767), .B2(n15666), .ZN(
        n45772) );
  AOI21_X1 U52648 ( .A1(n45770), .A2(n45769), .B(n46905), .ZN(n45771) );
  INV_X1 U52649 ( .I(n45774), .ZN(n45777) );
  AOI21_X1 U52650 ( .A1(n46911), .A2(n45775), .B(n23990), .ZN(n45776) );
  NOR3_X1 U52651 ( .A1(n45779), .A2(n47035), .A3(n1294), .ZN(n45780) );
  NAND2_X1 U52652 ( .A1(n47028), .A2(n45781), .ZN(n45782) );
  OAI22_X1 U52653 ( .A1(n20299), .A2(n47035), .B1(n13655), .B2(n23903), .ZN(
        n45786) );
  INV_X1 U52654 ( .I(n45787), .ZN(n45788) );
  NAND2_X1 U52655 ( .A1(n3971), .A2(n1474), .ZN(n45791) );
  NAND3_X1 U52656 ( .A1(n49057), .A2(n49046), .A3(n48067), .ZN(n45793) );
  NOR3_X1 U52657 ( .A1(n64167), .A2(n47920), .A3(n1474), .ZN(n45792) );
  NAND2_X1 U52661 ( .A1(n47688), .A2(n46835), .ZN(n45798) );
  NAND2_X1 U52663 ( .A1(n24099), .A2(n15728), .ZN(n45801) );
  NOR2_X1 U52664 ( .A1(n58018), .A2(n2955), .ZN(n45806) );
  NAND2_X1 U52665 ( .A1(n47378), .A2(n10475), .ZN(n45808) );
  XOR2_X1 U52666 ( .A1(n45811), .A2(n45812), .Z(n46609) );
  XOR2_X1 U52667 ( .A1(n50909), .A2(n45816), .Z(n45817) );
  XOR2_X1 U52668 ( .A1(n45818), .A2(n45817), .Z(n45820) );
  XOR2_X1 U52670 ( .A1(n46507), .A2(n45823), .Z(n46408) );
  INV_X1 U52673 ( .I(n45827), .ZN(n45828) );
  XOR2_X1 U52674 ( .A1(n22376), .A2(n45828), .Z(n45840) );
  INV_X1 U52675 ( .I(n45836), .ZN(n45832) );
  INV_X1 U52676 ( .I(n45835), .ZN(n45831) );
  XOR2_X1 U52677 ( .A1(n45830), .A2(n45829), .Z(n45833) );
  OAI21_X1 U52678 ( .A1(n45832), .A2(n45831), .B(n45833), .ZN(n45838) );
  INV_X1 U52679 ( .I(n45833), .ZN(n45834) );
  NAND3_X1 U52680 ( .A1(n45836), .A2(n45835), .A3(n45834), .ZN(n45837) );
  NAND2_X1 U52681 ( .A1(n45838), .A2(n45837), .ZN(n45839) );
  XOR2_X1 U52682 ( .A1(n45840), .A2(n45839), .Z(n45841) );
  XOR2_X1 U52683 ( .A1(n45841), .A2(n46440), .Z(n45842) );
  NAND2_X1 U52684 ( .A1(n48085), .A2(n64859), .ZN(n46763) );
  XOR2_X1 U52685 ( .A1(n45847), .A2(n45846), .Z(n45848) );
  XOR2_X1 U52686 ( .A1(n45849), .A2(n45848), .Z(n45850) );
  XOR2_X1 U52687 ( .A1(n45853), .A2(n52080), .Z(n45855) );
  XOR2_X1 U52688 ( .A1(n45855), .A2(n45854), .Z(n45856) );
  XOR2_X1 U52689 ( .A1(n23641), .A2(n45857), .Z(n45858) );
  XOR2_X1 U52690 ( .A1(n5093), .A2(n45865), .Z(n45866) );
  INV_X1 U52691 ( .I(n45867), .ZN(n45871) );
  XOR2_X1 U52692 ( .A1(n45869), .A2(n45868), .Z(n45870) );
  XOR2_X1 U52693 ( .A1(n45871), .A2(n45870), .Z(n45872) );
  XOR2_X1 U52694 ( .A1(n45873), .A2(n8813), .Z(n45874) );
  INV_X1 U52695 ( .I(n45876), .ZN(n45877) );
  XOR2_X1 U52696 ( .A1(n45879), .A2(n45878), .Z(n45881) );
  XOR2_X1 U52697 ( .A1(n45881), .A2(n45880), .Z(n45882) );
  XOR2_X1 U52698 ( .A1(n7544), .A2(n45882), .Z(n45883) );
  XOR2_X1 U52699 ( .A1(n45883), .A2(n1331), .Z(n45884) );
  NAND2_X1 U52706 ( .A1(n45897), .A2(n7395), .ZN(n45898) );
  MUX2_X1 U52710 ( .I0(n1486), .I1(n47434), .S(n47435), .Z(n45911) );
  NOR2_X1 U52711 ( .A1(n47437), .A2(n45907), .ZN(n45910) );
  NAND2_X1 U52712 ( .A1(n15421), .A2(n47728), .ZN(n45912) );
  NAND2_X1 U52713 ( .A1(n24374), .A2(n49948), .ZN(n45916) );
  NOR2_X1 U52714 ( .A1(n13614), .A2(n57543), .ZN(n45921) );
  NOR3_X1 U52715 ( .A1(n45923), .A2(n61624), .A3(n48317), .ZN(n45926) );
  NAND2_X1 U52716 ( .A1(n48026), .A2(n24374), .ZN(n45925) );
  NOR3_X1 U52717 ( .A1(n13614), .A2(n15550), .A3(n50268), .ZN(n45924) );
  NOR2_X1 U52718 ( .A1(n45929), .A2(n26180), .ZN(n46018) );
  NAND2_X1 U52719 ( .A1(n46018), .A2(n46017), .ZN(n45930) );
  NAND2_X1 U52720 ( .A1(n45932), .A2(n46024), .ZN(n45933) );
  MUX2_X1 U52721 ( .I0(n45934), .I1(n45933), .S(n47297), .Z(n45940) );
  NAND2_X1 U52725 ( .A1(n47894), .A2(n47900), .ZN(n45948) );
  NAND2_X1 U52726 ( .A1(n61889), .A2(n45946), .ZN(n45947) );
  AOI21_X1 U52727 ( .A1(n45949), .A2(n24290), .B(n47896), .ZN(n45950) );
  NAND2_X1 U52728 ( .A1(n46066), .A2(n7389), .ZN(n45952) );
  NAND2_X1 U52729 ( .A1(n7389), .A2(n20832), .ZN(n45955) );
  OAI22_X1 U52731 ( .A1(n8603), .A2(n61961), .B1(n45962), .B2(n45961), .ZN(
        n45965) );
  INV_X1 U52733 ( .I(n47289), .ZN(n45975) );
  AOI22_X1 U52734 ( .A1(n47282), .A2(n45975), .B1(n47594), .B2(n45979), .ZN(
        n45977) );
  NAND2_X1 U52735 ( .A1(n45978), .A2(n45976), .ZN(n47597) );
  INV_X1 U52736 ( .I(n47273), .ZN(n45983) );
  NAND2_X1 U52738 ( .A1(n49109), .A2(n20708), .ZN(n45997) );
  NAND2_X1 U52739 ( .A1(n47616), .A2(n58155), .ZN(n45987) );
  AOI21_X1 U52741 ( .A1(n22239), .A2(n45988), .B(n1069), .ZN(n45989) );
  OAI21_X1 U52742 ( .A1(n22468), .A2(n22239), .B(n45989), .ZN(n45995) );
  NAND3_X1 U52743 ( .A1(n1663), .A2(n47615), .A3(n59059), .ZN(n45994) );
  NAND2_X1 U52744 ( .A1(n47343), .A2(n7146), .ZN(n48443) );
  AOI22_X1 U52747 ( .A1(n46000), .A2(n49793), .B1(n19646), .B2(n48436), .ZN(
        n46003) );
  NOR2_X1 U52748 ( .A1(n47346), .A2(n49115), .ZN(n46001) );
  NAND2_X1 U52749 ( .A1(n46004), .A2(n47947), .ZN(n46007) );
  INV_X1 U52750 ( .I(n47941), .ZN(n46006) );
  AOI22_X1 U52752 ( .A1(n46008), .A2(n46007), .B1(n46006), .B2(n46005), .ZN(
        n46009) );
  NAND2_X1 U52753 ( .A1(n1078), .A2(n46013), .ZN(n46015) );
  NAND3_X1 U52755 ( .A1(n46018), .A2(n46017), .A3(n25477), .ZN(n46019) );
  OAI22_X1 U52756 ( .A1(n24578), .A2(n46866), .B1(n46871), .B2(n46027), .ZN(
        n46029) );
  NAND2_X1 U52757 ( .A1(n46029), .A2(n46028), .ZN(n46046) );
  NAND2_X1 U52758 ( .A1(n20426), .A2(n1666), .ZN(n46032) );
  NAND2_X1 U52759 ( .A1(n9988), .A2(n46039), .ZN(n46030) );
  AOI21_X1 U52760 ( .A1(n46871), .A2(n20426), .B(n46034), .ZN(n46035) );
  NOR2_X1 U52761 ( .A1(n46036), .A2(n46035), .ZN(n46045) );
  NOR2_X1 U52763 ( .A1(n46038), .A2(n63501), .ZN(n46042) );
  NOR2_X1 U52764 ( .A1(n46040), .A2(n64888), .ZN(n46041) );
  NOR2_X1 U52766 ( .A1(n49777), .A2(n49767), .ZN(n46068) );
  NAND2_X1 U52768 ( .A1(n58009), .A2(n47227), .ZN(n46057) );
  OAI21_X1 U52769 ( .A1(n19715), .A2(n46946), .B(n22852), .ZN(n46054) );
  NAND2_X1 U52770 ( .A1(n47233), .A2(n46054), .ZN(n46055) );
  NAND2_X1 U52771 ( .A1(n47329), .A2(n20832), .ZN(n46928) );
  INV_X1 U52772 ( .I(n46928), .ZN(n46063) );
  AOI21_X1 U52774 ( .A1(n46068), .A2(n149), .B(n63724), .ZN(n46086) );
  NOR2_X1 U52775 ( .A1(n46075), .A2(n57234), .ZN(n46073) );
  OAI21_X1 U52776 ( .A1(n58705), .A2(n46070), .B(n46069), .ZN(n46072) );
  NAND2_X1 U52778 ( .A1(n46082), .A2(n49774), .ZN(n46085) );
  INV_X1 U52779 ( .I(n47249), .ZN(n46081) );
  NOR2_X1 U52780 ( .A1(n46077), .A2(n21793), .ZN(n46080) );
  NOR2_X1 U52781 ( .A1(n49770), .A2(n21550), .ZN(n46083) );
  NAND2_X1 U52782 ( .A1(n49780), .A2(n48949), .ZN(n46088) );
  OAI22_X1 U52783 ( .A1(n46088), .A2(n48947), .B1(n48950), .B2(n46087), .ZN(
        n46091) );
  NAND3_X1 U52784 ( .A1(n4017), .A2(n63724), .A3(n47972), .ZN(n46089) );
  NAND2_X1 U52785 ( .A1(n46096), .A2(n20090), .ZN(n47003) );
  OAI21_X1 U52786 ( .A1(n8012), .A2(n61212), .B(n47003), .ZN(n46094) );
  NOR2_X1 U52788 ( .A1(n20162), .A2(n44770), .ZN(n46104) );
  INV_X1 U52789 ( .I(n46111), .ZN(n46116) );
  XOR2_X1 U52790 ( .A1(n56976), .A2(n58077), .Z(n46113) );
  XOR2_X1 U52791 ( .A1(n46114), .A2(n46113), .Z(n46115) );
  XOR2_X1 U52792 ( .A1(n46116), .A2(n46115), .Z(n46117) );
  XOR2_X1 U52793 ( .A1(n46125), .A2(n46553), .Z(n46126) );
  XOR2_X1 U52794 ( .A1(n46129), .A2(n46128), .Z(n46131) );
  XOR2_X1 U52795 ( .A1(n46131), .A2(n46130), .Z(n46132) );
  XOR2_X1 U52798 ( .A1(n46142), .A2(n46141), .Z(n46143) );
  XOR2_X1 U52799 ( .A1(n46145), .A2(n46144), .Z(n46146) );
  XOR2_X1 U52800 ( .A1(n7202), .A2(n23818), .Z(n46157) );
  XOR2_X1 U52801 ( .A1(n46684), .A2(n52095), .Z(n46151) );
  XOR2_X1 U52802 ( .A1(n46152), .A2(n46151), .Z(n46153) );
  XOR2_X1 U52803 ( .A1(n46154), .A2(n46153), .Z(n46155) );
  XOR2_X1 U52804 ( .A1(n64258), .A2(n46155), .Z(n46156) );
  XOR2_X1 U52807 ( .A1(n63448), .A2(n23059), .Z(n46173) );
  XNOR2_X1 U52808 ( .A1(n51493), .A2(n53772), .ZN(n46167) );
  XOR2_X1 U52809 ( .A1(n46168), .A2(n46167), .Z(n46169) );
  XOR2_X1 U52810 ( .A1(n46170), .A2(n46169), .Z(n46171) );
  XOR2_X1 U52811 ( .A1(n22207), .A2(n46171), .Z(n46172) );
  XOR2_X1 U52812 ( .A1(n46173), .A2(n46172), .Z(n46174) );
  NAND3_X1 U52814 ( .A1(n46176), .A2(n10621), .A3(n59071), .ZN(n48180) );
  XOR2_X1 U52815 ( .A1(n1190), .A2(n55242), .Z(n46181) );
  XOR2_X1 U52816 ( .A1(n50698), .A2(n46181), .Z(n46182) );
  XOR2_X1 U52817 ( .A1(n46183), .A2(n46182), .Z(n46184) );
  XOR2_X1 U52818 ( .A1(n23953), .A2(n46184), .Z(n46185) );
  INV_X1 U52819 ( .I(n46191), .ZN(n46194) );
  XOR2_X1 U52820 ( .A1(n46192), .A2(n50832), .Z(n46193) );
  XOR2_X1 U52821 ( .A1(n46194), .A2(n46193), .Z(n46195) );
  XOR2_X1 U52822 ( .A1(n46198), .A2(n46197), .Z(n46199) );
  XOR2_X1 U52824 ( .A1(n46211), .A2(n64443), .Z(n46697) );
  XOR2_X1 U52825 ( .A1(n19226), .A2(n23722), .Z(n46214) );
  XOR2_X1 U52826 ( .A1(n46218), .A2(n46217), .Z(n46227) );
  XOR2_X1 U52827 ( .A1(n46220), .A2(n23767), .Z(n46222) );
  XOR2_X1 U52828 ( .A1(n46222), .A2(n46221), .Z(n46223) );
  XOR2_X1 U52829 ( .A1(n46557), .A2(n46223), .Z(n46225) );
  XOR2_X1 U52830 ( .A1(n46225), .A2(n22923), .Z(n46226) );
  XOR2_X1 U52832 ( .A1(n19232), .A2(n46230), .Z(n46232) );
  XOR2_X1 U52833 ( .A1(n46234), .A2(n46233), .Z(n46655) );
  XOR2_X1 U52834 ( .A1(n46239), .A2(n46238), .Z(n46240) );
  XOR2_X1 U52835 ( .A1(n12178), .A2(n46240), .Z(n46241) );
  INV_X1 U52836 ( .I(n46246), .ZN(n46247) );
  XOR2_X1 U52837 ( .A1(n46248), .A2(n46247), .Z(n46249) );
  XOR2_X1 U52838 ( .A1(n46249), .A2(n50251), .Z(n46250) );
  INV_X1 U52839 ( .I(n46252), .ZN(n46256) );
  XOR2_X1 U52840 ( .A1(n61457), .A2(n22731), .Z(n46612) );
  XOR2_X1 U52841 ( .A1(n46612), .A2(n46254), .Z(n46255) );
  XOR2_X1 U52842 ( .A1(n46256), .A2(n46255), .Z(n46257) );
  OAI21_X1 U52843 ( .A1(n46259), .A2(n48213), .B(n46997), .ZN(n46260) );
  NAND2_X1 U52846 ( .A1(n12850), .A2(n23035), .ZN(n46264) );
  NAND2_X1 U52848 ( .A1(n47042), .A2(n12850), .ZN(n46265) );
  XOR2_X1 U52849 ( .A1(n51913), .A2(n46273), .Z(n46274) );
  XOR2_X1 U52850 ( .A1(n46275), .A2(n46274), .Z(n46277) );
  XOR2_X1 U52851 ( .A1(n46277), .A2(n46276), .Z(n46278) );
  XOR2_X1 U52852 ( .A1(n46279), .A2(n46278), .Z(n46280) );
  XOR2_X1 U52853 ( .A1(n22247), .A2(n23687), .Z(n46290) );
  XOR2_X1 U52854 ( .A1(n46286), .A2(n46285), .Z(n46287) );
  XOR2_X1 U52856 ( .A1(n10043), .A2(n23722), .Z(n46293) );
  XOR2_X1 U52858 ( .A1(n46296), .A2(n46697), .Z(n46297) );
  INV_X1 U52859 ( .I(n46301), .ZN(n46303) );
  XOR2_X1 U52860 ( .A1(n46303), .A2(n46302), .Z(n46304) );
  XOR2_X1 U52861 ( .A1(n22639), .A2(n46304), .Z(n46306) );
  XOR2_X1 U52862 ( .A1(n46307), .A2(n46306), .Z(n46308) );
  XOR2_X1 U52864 ( .A1(n46316), .A2(n46315), .Z(n46317) );
  NAND2_X1 U52865 ( .A1(n10487), .A2(n46336), .ZN(n46327) );
  NAND2_X1 U52866 ( .A1(n13680), .A2(n46336), .ZN(n46325) );
  OAI22_X1 U52867 ( .A1(n46328), .A2(n46327), .B1(n46326), .B2(n46325), .ZN(
        n46330) );
  INV_X1 U52868 ( .I(n46337), .ZN(n46329) );
  NAND2_X1 U52869 ( .A1(n46330), .A2(n46329), .ZN(n46342) );
  NAND3_X1 U52870 ( .A1(n46333), .A2(n46332), .A3(n10487), .ZN(n46340) );
  AOI21_X1 U52871 ( .A1(n57525), .A2(n13680), .B(n46336), .ZN(n46339) );
  INV_X1 U52872 ( .I(n46336), .ZN(n46338) );
  AOI22_X1 U52873 ( .A1(n46340), .A2(n46339), .B1(n46338), .B2(n46337), .ZN(
        n46341) );
  XOR2_X1 U52874 ( .A1(n46349), .A2(n46348), .Z(n46350) );
  XOR2_X1 U52875 ( .A1(n46351), .A2(n46350), .Z(n46352) );
  XOR2_X1 U52876 ( .A1(n46355), .A2(n46354), .Z(n46356) );
  NAND2_X2 U52878 ( .A1(n47541), .A2(n25855), .ZN(n47545) );
  NAND4_X1 U52879 ( .A1(n48623), .A2(n3341), .A3(n47545), .A4(n58675), .ZN(
        n46360) );
  NAND3_X1 U52880 ( .A1(n46358), .A2(n3340), .A3(n46357), .ZN(n46359) );
  NAND3_X1 U52881 ( .A1(n47542), .A2(n22635), .A3(n65059), .ZN(n46363) );
  INV_X1 U52882 ( .I(n49412), .ZN(n46369) );
  XOR2_X1 U52883 ( .A1(n46371), .A2(n53375), .Z(n46372) );
  XOR2_X1 U52884 ( .A1(n46373), .A2(n46372), .Z(n46374) );
  XOR2_X1 U52885 ( .A1(n46375), .A2(n46374), .Z(n46376) );
  INV_X1 U52886 ( .I(n24094), .ZN(n46378) );
  XOR2_X1 U52887 ( .A1(n46379), .A2(n46378), .Z(n46380) );
  XOR2_X1 U52888 ( .A1(n46388), .A2(n46387), .Z(n46389) );
  XOR2_X1 U52889 ( .A1(n46390), .A2(n46389), .Z(n46391) );
  XOR2_X1 U52890 ( .A1(n46393), .A2(n22340), .Z(n46394) );
  INV_X1 U52891 ( .I(n46396), .ZN(n46402) );
  XOR2_X1 U52892 ( .A1(n46398), .A2(n46684), .Z(n46399) );
  XOR2_X1 U52893 ( .A1(n46400), .A2(n46399), .Z(n46401) );
  XOR2_X1 U52894 ( .A1(n46402), .A2(n46401), .Z(n46404) );
  XOR2_X1 U52895 ( .A1(n46404), .A2(n46403), .Z(n46405) );
  XOR2_X1 U52896 ( .A1(n19994), .A2(n46405), .Z(n46406) );
  XOR2_X1 U52897 ( .A1(n46409), .A2(n46408), .Z(n46410) );
  NAND2_X1 U52898 ( .A1(n48462), .A2(n7186), .ZN(n46431) );
  NOR2_X1 U52899 ( .A1(n47084), .A2(n48472), .ZN(n48471) );
  XOR2_X1 U52900 ( .A1(n46414), .A2(n46413), .Z(n46417) );
  XOR2_X1 U52901 ( .A1(n46415), .A2(n29407), .Z(n46416) );
  INV_X1 U52902 ( .I(n50190), .ZN(n46423) );
  XNOR2_X1 U52903 ( .A1(n53764), .A2(n54563), .ZN(n46422) );
  XOR2_X1 U52904 ( .A1(n46423), .A2(n46422), .Z(n46424) );
  XOR2_X1 U52905 ( .A1(n46425), .A2(n46424), .Z(n46426) );
  XOR2_X1 U52906 ( .A1(n24055), .A2(n20900), .Z(n46434) );
  XOR2_X1 U52907 ( .A1(n46529), .A2(n46437), .Z(n46439) );
  XOR2_X1 U52908 ( .A1(n46439), .A2(n46438), .Z(n46441) );
  XOR2_X1 U52909 ( .A1(n63789), .A2(n22376), .Z(n46448) );
  XOR2_X1 U52910 ( .A1(n46444), .A2(n46443), .Z(n46445) );
  XOR2_X1 U52911 ( .A1(n22207), .A2(n46445), .Z(n46447) );
  XOR2_X1 U52912 ( .A1(n46448), .A2(n46447), .Z(n46449) );
  XOR2_X1 U52913 ( .A1(n18726), .A2(n46449), .Z(n46450) );
  XOR2_X1 U52914 ( .A1(n46451), .A2(n46450), .Z(n46452) );
  XOR2_X1 U52915 ( .A1(n46453), .A2(n46452), .Z(n48130) );
  NOR2_X2 U52916 ( .A1(n48134), .A2(n24545), .ZN(n48475) );
  AOI22_X1 U52918 ( .A1(n46454), .A2(n48459), .B1(n47079), .B2(n60398), .ZN(
        n46457) );
  NOR2_X1 U52919 ( .A1(n48219), .A2(n62308), .ZN(n46465) );
  NAND2_X1 U52920 ( .A1(n48614), .A2(n8639), .ZN(n46461) );
  OAI22_X1 U52921 ( .A1(n48218), .A2(n46461), .B1(n46460), .B2(n48620), .ZN(
        n46464) );
  NAND3_X1 U52922 ( .A1(n62308), .A2(n47180), .A3(n58675), .ZN(n46462) );
  NOR2_X1 U52924 ( .A1(n47545), .A2(n22703), .ZN(n48220) );
  OAI21_X1 U52925 ( .A1(n48220), .A2(n3341), .B(n48626), .ZN(n46466) );
  NOR2_X1 U52929 ( .A1(n2403), .A2(n48484), .ZN(n46475) );
  INV_X1 U52930 ( .I(n48176), .ZN(n46473) );
  NAND2_X1 U52932 ( .A1(n48174), .A2(n46475), .ZN(n46476) );
  NOR2_X1 U52935 ( .A1(n19200), .A2(n48177), .ZN(n46484) );
  INV_X1 U52936 ( .I(n46486), .ZN(n46491) );
  XOR2_X1 U52937 ( .A1(n46487), .A2(n51814), .Z(n46489) );
  XOR2_X1 U52938 ( .A1(n46489), .A2(n46488), .Z(n46490) );
  XOR2_X1 U52939 ( .A1(n46491), .A2(n46490), .Z(n46492) );
  XOR2_X1 U52940 ( .A1(n23953), .A2(n46492), .Z(n46494) );
  XOR2_X1 U52941 ( .A1(n64349), .A2(n58532), .Z(n46498) );
  INV_X1 U52942 ( .I(n46500), .ZN(n46504) );
  XOR2_X1 U52943 ( .A1(n50126), .A2(n54556), .Z(n46686) );
  XOR2_X1 U52944 ( .A1(n46601), .A2(n46501), .Z(n46502) );
  XOR2_X1 U52945 ( .A1(n46686), .A2(n46502), .Z(n46503) );
  XOR2_X1 U52946 ( .A1(n46504), .A2(n46503), .Z(n46505) );
  XOR2_X1 U52947 ( .A1(n61363), .A2(n46506), .Z(n46508) );
  INV_X1 U52948 ( .I(n46514), .ZN(n46516) );
  XOR2_X1 U52949 ( .A1(n46516), .A2(n46515), .Z(n46517) );
  XOR2_X1 U52950 ( .A1(n21141), .A2(n46517), .Z(n46518) );
  XOR2_X1 U52951 ( .A1(n46524), .A2(n46523), .Z(n46525) );
  XOR2_X1 U52952 ( .A1(n23872), .A2(n61071), .Z(n46537) );
  INV_X1 U52953 ( .I(n46531), .ZN(n46533) );
  XOR2_X1 U52954 ( .A1(n46533), .A2(n46532), .Z(n46534) );
  XOR2_X1 U52955 ( .A1(n46535), .A2(n46534), .Z(n46536) );
  XOR2_X1 U52956 ( .A1(n46537), .A2(n46536), .Z(n46540) );
  XOR2_X1 U52957 ( .A1(n64971), .A2(n23445), .Z(n46539) );
  INV_X1 U52960 ( .I(n46543), .ZN(n46544) );
  XOR2_X1 U52961 ( .A1(n46545), .A2(n46544), .Z(n48161) );
  XOR2_X1 U52962 ( .A1(n46549), .A2(n54386), .Z(n46551) );
  XOR2_X1 U52963 ( .A1(n46555), .A2(n46554), .Z(n46556) );
  XOR2_X1 U52964 ( .A1(n46557), .A2(n46556), .Z(n46559) );
  XOR2_X1 U52965 ( .A1(n46558), .A2(n46559), .Z(n46560) );
  NAND2_X1 U52966 ( .A1(n48166), .A2(n48514), .ZN(n46563) );
  AOI21_X1 U52968 ( .A1(n46564), .A2(n46563), .B(n46562), .ZN(n46568) );
  INV_X4 U52969 ( .I(n20937), .ZN(n48511) );
  NOR2_X1 U52970 ( .A1(n48636), .A2(n48504), .ZN(n46565) );
  XOR2_X1 U52971 ( .A1(n51575), .A2(n46571), .Z(n46572) );
  XOR2_X1 U52973 ( .A1(n46583), .A2(n15735), .Z(n46584) );
  XOR2_X1 U52974 ( .A1(n46585), .A2(n46584), .Z(n46586) );
  XOR2_X1 U52975 ( .A1(n23905), .A2(n46586), .Z(n46588) );
  XOR2_X1 U52976 ( .A1(n7264), .A2(n46593), .Z(n46594) );
  XOR2_X1 U52977 ( .A1(n46595), .A2(n46594), .Z(n46596) );
  INV_X1 U52978 ( .I(n50585), .ZN(n46602) );
  XOR2_X1 U52979 ( .A1(n46602), .A2(n46601), .Z(n46604) );
  XOR2_X1 U52980 ( .A1(n46604), .A2(n46603), .Z(n46606) );
  XOR2_X1 U52981 ( .A1(n46606), .A2(n23553), .Z(n46607) );
  XOR2_X1 U52982 ( .A1(n46611), .A2(n13069), .Z(n46614) );
  XOR2_X1 U52983 ( .A1(n46616), .A2(n46615), .Z(n46618) );
  XOR2_X1 U52984 ( .A1(n46618), .A2(n46617), .Z(n46619) );
  XOR2_X1 U52985 ( .A1(n46621), .A2(n46622), .Z(n46623) );
  INV_X1 U52987 ( .I(n46631), .ZN(n46633) );
  XOR2_X1 U52988 ( .A1(n52577), .A2(n51275), .Z(n46632) );
  XOR2_X1 U52989 ( .A1(n46633), .A2(n46632), .Z(n46634) );
  XOR2_X1 U52990 ( .A1(n16518), .A2(n46635), .Z(n46636) );
  NOR2_X1 U52991 ( .A1(n24364), .A2(n46751), .ZN(n46638) );
  NOR2_X1 U52993 ( .A1(n48553), .A2(n46751), .ZN(n46641) );
  NAND2_X1 U52994 ( .A1(n47097), .A2(n21820), .ZN(n46642) );
  NAND2_X1 U52995 ( .A1(n46643), .A2(n46642), .ZN(n46644) );
  XOR2_X1 U52996 ( .A1(n46648), .A2(n46647), .Z(n46649) );
  XOR2_X1 U52997 ( .A1(n46650), .A2(n46649), .Z(n46651) );
  XOR2_X1 U52998 ( .A1(n46653), .A2(n46652), .Z(n46654) );
  XOR2_X1 U52999 ( .A1(n46659), .A2(n56849), .Z(n46662) );
  INV_X1 U53000 ( .I(n46660), .ZN(n46661) );
  XOR2_X1 U53001 ( .A1(n46662), .A2(n46661), .Z(n46663) );
  XOR2_X1 U53002 ( .A1(n57892), .A2(n46663), .Z(n46665) );
  INV_X1 U53004 ( .I(n46669), .ZN(n46670) );
  XOR2_X1 U53005 ( .A1(n46670), .A2(n51193), .Z(n46672) );
  XOR2_X1 U53006 ( .A1(n46672), .A2(n46671), .Z(n46673) );
  XOR2_X1 U53008 ( .A1(n46680), .A2(n46681), .Z(n46695) );
  XOR2_X1 U53009 ( .A1(n46683), .A2(n46682), .Z(n51793) );
  XOR2_X1 U53010 ( .A1(n46684), .A2(n50502), .Z(n46685) );
  XOR2_X1 U53011 ( .A1(n46686), .A2(n46685), .Z(n46687) );
  XOR2_X1 U53012 ( .A1(n51793), .A2(n46687), .Z(n46689) );
  XOR2_X1 U53013 ( .A1(n23618), .A2(n58532), .Z(n46692) );
  XOR2_X1 U53014 ( .A1(n46693), .A2(n46692), .Z(n46694) );
  XOR2_X1 U53015 ( .A1(n46698), .A2(n55546), .Z(n46699) );
  XOR2_X1 U53016 ( .A1(n52366), .A2(n46699), .Z(n46700) );
  XOR2_X1 U53017 ( .A1(n22212), .A2(n46700), .Z(n46703) );
  XOR2_X1 U53018 ( .A1(n46703), .A2(n23402), .Z(n46704) );
  INV_X1 U53019 ( .I(n46707), .ZN(n46710) );
  XOR2_X1 U53020 ( .A1(n46708), .A2(n53246), .Z(n46709) );
  XOR2_X1 U53021 ( .A1(n46710), .A2(n46709), .Z(n46711) );
  XOR2_X1 U53022 ( .A1(n23270), .A2(n46711), .Z(n46712) );
  OAI22_X1 U53023 ( .A1(n47192), .A2(n47185), .B1(n47194), .B2(n46715), .ZN(
        n46718) );
  NAND2_X1 U53025 ( .A1(n48232), .A2(n48540), .ZN(n46717) );
  INV_X1 U53026 ( .I(n49420), .ZN(n46721) );
  AOI21_X1 U53027 ( .A1(n50081), .A2(n46723), .B(n21183), .ZN(n46720) );
  NAND2_X1 U53029 ( .A1(n50407), .A2(n22764), .ZN(n46728) );
  NOR2_X1 U53030 ( .A1(n47730), .A2(n46731), .ZN(n47747) );
  INV_X1 U53031 ( .I(n47747), .ZN(n46732) );
  NAND2_X1 U53033 ( .A1(n24252), .A2(n47736), .ZN(n46738) );
  NAND3_X1 U53036 ( .A1(n23934), .A2(n47368), .A3(n21451), .ZN(n46747) );
  NOR2_X1 U53037 ( .A1(n47370), .A2(n23718), .ZN(n46749) );
  NOR2_X1 U53039 ( .A1(n22874), .A2(n46751), .ZN(n46752) );
  OAI21_X1 U53041 ( .A1(n57740), .A2(n63465), .B(n47415), .ZN(n46754) );
  INV_X1 U53045 ( .I(n48566), .ZN(n46767) );
  INV_X1 U53049 ( .I(n64036), .ZN(n47122) );
  NAND2_X1 U53051 ( .A1(n48571), .A2(n57398), .ZN(n46773) );
  MUX2_X1 U53055 ( .I0(n48087), .I1(n46782), .S(n64859), .Z(n46786) );
  MUX2_X1 U53056 ( .I0(n48076), .I1(n48572), .S(n48085), .Z(n46784) );
  OAI21_X1 U53057 ( .A1(n47123), .A2(n23617), .B(n47128), .ZN(n46783) );
  NOR2_X1 U53058 ( .A1(n48144), .A2(n48552), .ZN(n46789) );
  NOR2_X1 U53059 ( .A1(n47100), .A2(n24364), .ZN(n46793) );
  OAI21_X1 U53060 ( .A1(n18099), .A2(n59160), .B(n48544), .ZN(n46792) );
  OAI21_X1 U53061 ( .A1(n46793), .A2(n46792), .B(n48154), .ZN(n46796) );
  NAND3_X1 U53062 ( .A1(n48155), .A2(n60138), .A3(n46798), .ZN(n46801) );
  NAND2_X1 U53063 ( .A1(n47209), .A2(n48136), .ZN(n46803) );
  NAND3_X1 U53064 ( .A1(n48475), .A2(n10626), .A3(n7186), .ZN(n46807) );
  NAND3_X1 U53065 ( .A1(n47209), .A2(n63105), .A3(n47087), .ZN(n46806) );
  NOR2_X1 U53066 ( .A1(n47204), .A2(n48472), .ZN(n46804) );
  NAND2_X1 U53067 ( .A1(n24354), .A2(n24099), .ZN(n46810) );
  NAND3_X1 U53070 ( .A1(n23850), .A2(n15728), .A3(n12698), .ZN(n46818) );
  NAND3_X1 U53071 ( .A1(n48098), .A2(n46819), .A3(n46818), .ZN(n46820) );
  OAI21_X1 U53073 ( .A1(n23934), .A2(n10172), .B(n46824), .ZN(n46825) );
  AOI22_X1 U53074 ( .A1(n47378), .A2(n17951), .B1(n47382), .B2(n10475), .ZN(
        n46829) );
  NOR2_X1 U53076 ( .A1(n49620), .A2(n46833), .ZN(n46849) );
  NAND2_X1 U53077 ( .A1(n47418), .A2(n46835), .ZN(n46836) );
  NAND3_X1 U53078 ( .A1(n47413), .A2(n47686), .A3(n46836), .ZN(n46837) );
  NAND2_X1 U53079 ( .A1(n46837), .A2(n47688), .ZN(n46848) );
  NAND2_X1 U53080 ( .A1(n47682), .A2(n263), .ZN(n46838) );
  AOI21_X1 U53081 ( .A1(n47427), .A2(n46838), .B(n1263), .ZN(n46842) );
  INV_X1 U53082 ( .I(n47687), .ZN(n46839) );
  AOI21_X1 U53083 ( .A1(n46839), .A2(n45267), .B(n59205), .ZN(n46841) );
  OAI21_X1 U53084 ( .A1(n47687), .A2(n46843), .B(n47427), .ZN(n46844) );
  NAND2_X1 U53085 ( .A1(n46845), .A2(n46844), .ZN(n46846) );
  NOR2_X1 U53087 ( .A1(n47924), .A2(n50376), .ZN(n46852) );
  INV_X1 U53088 ( .I(n49721), .ZN(n50382) );
  AOI21_X1 U53089 ( .A1(n49619), .A2(n50382), .B(n49039), .ZN(n46855) );
  NAND2_X1 U53090 ( .A1(n47933), .A2(n23707), .ZN(n46854) );
  NOR2_X1 U53091 ( .A1(n46855), .A2(n46854), .ZN(n49617) );
  INV_X1 U53092 ( .I(n46858), .ZN(n46860) );
  INV_X1 U53094 ( .I(n46862), .ZN(n46870) );
  NAND2_X1 U53096 ( .A1(n46872), .A2(n46871), .ZN(n46878) );
  INV_X1 U53097 ( .I(n46873), .ZN(n46877) );
  NOR2_X1 U53098 ( .A1(n46875), .A2(n20426), .ZN(n46876) );
  OAI21_X1 U53099 ( .A1(n46878), .A2(n46877), .B(n46876), .ZN(n46879) );
  INV_X1 U53100 ( .I(n46882), .ZN(n46896) );
  OAI21_X1 U53101 ( .A1(n46896), .A2(n47262), .B(n46883), .ZN(n46889) );
  NAND4_X1 U53105 ( .A1(n46896), .A2(n59418), .A3(n21793), .A4(n16212), .ZN(
        n46903) );
  NAND3_X1 U53106 ( .A1(n47267), .A2(n59707), .A3(n60753), .ZN(n46902) );
  AOI21_X1 U53107 ( .A1(n47250), .A2(n59707), .B(n47259), .ZN(n46899) );
  NAND2_X1 U53108 ( .A1(n21976), .A2(n47250), .ZN(n46898) );
  NAND4_X1 U53109 ( .A1(n46900), .A2(n46899), .A3(n47252), .A4(n46898), .ZN(
        n46901) );
  NOR3_X1 U53110 ( .A1(n23990), .A2(n46913), .A3(n23480), .ZN(n46915) );
  NAND2_X1 U53111 ( .A1(n46920), .A2(n63700), .ZN(n46935) );
  AOI21_X1 U53112 ( .A1(n46930), .A2(n46929), .B(n46928), .ZN(n46931) );
  INV_X1 U53114 ( .I(n46936), .ZN(n46937) );
  OAI21_X1 U53115 ( .A1(n47984), .A2(n47986), .B(n47985), .ZN(n46945) );
  AOI21_X1 U53119 ( .A1(n48808), .A2(n48422), .B(n48421), .ZN(n46972) );
  NAND2_X1 U53120 ( .A1(n47923), .A2(n48690), .ZN(n50754) );
  NAND3_X1 U53121 ( .A1(n50754), .A2(n64167), .A3(n48683), .ZN(n46975) );
  NAND2_X1 U53122 ( .A1(n46982), .A2(n44065), .ZN(n47466) );
  NOR2_X1 U53123 ( .A1(n47466), .A2(n58174), .ZN(n46983) );
  NAND2_X1 U53124 ( .A1(n46985), .A2(n10055), .ZN(n46986) );
  OAI21_X1 U53125 ( .A1(n46989), .A2(n46988), .B(n46987), .ZN(n46990) );
  NAND2_X1 U53126 ( .A1(n48199), .A2(n48208), .ZN(n46991) );
  NAND4_X1 U53127 ( .A1(n46993), .A2(n48209), .A3(n48212), .A4(n47197), .ZN(
        n46994) );
  INV_X1 U53128 ( .I(n46995), .ZN(n46999) );
  INV_X1 U53129 ( .I(n46996), .ZN(n46998) );
  NAND2_X1 U53130 ( .A1(n22684), .A2(n5771), .ZN(n47002) );
  AOI21_X1 U53131 ( .A1(n47003), .A2(n61993), .B(n47002), .ZN(n47010) );
  INV_X1 U53134 ( .I(n47016), .ZN(n47012) );
  NAND3_X1 U53135 ( .A1(n47013), .A2(n47012), .A3(n20090), .ZN(n47015) );
  OAI21_X1 U53136 ( .A1(n22872), .A2(n20238), .B(n47022), .ZN(n47024) );
  NAND3_X1 U53138 ( .A1(n47029), .A2(n64063), .A3(n47028), .ZN(n47031) );
  NOR2_X1 U53141 ( .A1(n9594), .A2(n64341), .ZN(n49502) );
  NAND4_X1 U53145 ( .A1(n48038), .A2(n49013), .A3(n48323), .A4(n23738), .ZN(
        n47051) );
  NAND3_X1 U53146 ( .A1(n47059), .A2(n49266), .A3(n49412), .ZN(n47060) );
  NAND2_X1 U53147 ( .A1(n7078), .A2(n61513), .ZN(n47061) );
  MUX2_X1 U53148 ( .I0(n47063), .I1(n47062), .S(n359), .Z(n47064) );
  NAND2_X1 U53149 ( .A1(n49784), .A2(n49776), .ZN(n47072) );
  NAND2_X1 U53152 ( .A1(n47972), .A2(n57735), .ZN(n47069) );
  AOI21_X1 U53153 ( .A1(n47977), .A2(n21737), .B(n47069), .ZN(n47070) );
  XOR2_X1 U53154 ( .A1(n20874), .A2(n51601), .Z(n52610) );
  NAND2_X1 U53158 ( .A1(n47083), .A2(n48472), .ZN(n47081) );
  NOR2_X1 U53159 ( .A1(n48472), .A2(n60358), .ZN(n47085) );
  NAND2_X1 U53160 ( .A1(n47088), .A2(n47211), .ZN(n47090) );
  NAND2_X1 U53161 ( .A1(n47088), .A2(n48459), .ZN(n47089) );
  OAI21_X1 U53165 ( .A1(n23185), .A2(n47099), .B(n47098), .ZN(n47105) );
  NOR2_X1 U53166 ( .A1(n63547), .A2(n60138), .ZN(n47104) );
  NAND2_X1 U53168 ( .A1(n22874), .A2(n63422), .ZN(n47102) );
  NAND2_X1 U53169 ( .A1(n19144), .A2(n23299), .ZN(n47763) );
  NOR2_X1 U53170 ( .A1(n10624), .A2(n48566), .ZN(n47118) );
  NAND2_X1 U53171 ( .A1(n48561), .A2(n697), .ZN(n47126) );
  AOI22_X1 U53172 ( .A1(n47124), .A2(n48577), .B1(n48559), .B2(n47123), .ZN(
        n47125) );
  NAND3_X1 U53175 ( .A1(n17905), .A2(n49862), .A3(n48530), .ZN(n47133) );
  NOR2_X1 U53177 ( .A1(n16227), .A2(n48538), .ZN(n47136) );
  AOI21_X1 U53178 ( .A1(n23934), .A2(n47367), .B(n47144), .ZN(n47143) );
  MUX2_X1 U53179 ( .I0(n47763), .I1(n47148), .S(n50444), .Z(n47151) );
  AOI21_X1 U53180 ( .A1(n47149), .A2(n50239), .B(n59621), .ZN(n47150) );
  INV_X1 U53181 ( .I(n47153), .ZN(n47155) );
  NOR2_X1 U53182 ( .A1(n47155), .A2(n4655), .ZN(n47159) );
  NAND2_X1 U53183 ( .A1(n48482), .A2(n9851), .ZN(n47157) );
  OAI22_X1 U53184 ( .A1(n47157), .A2(n48587), .B1(n23542), .B2(n48588), .ZN(
        n47158) );
  NOR2_X1 U53185 ( .A1(n48487), .A2(n10621), .ZN(n47160) );
  NAND2_X1 U53186 ( .A1(n47167), .A2(n47163), .ZN(n47164) );
  INV_X1 U53187 ( .I(n47550), .ZN(n47168) );
  INV_X1 U53188 ( .I(n48623), .ZN(n47170) );
  NAND2_X1 U53189 ( .A1(n47170), .A2(n48620), .ZN(n47171) );
  INV_X1 U53190 ( .I(n47175), .ZN(n47176) );
  NOR2_X1 U53191 ( .A1(n3341), .A2(n65059), .ZN(n47179) );
  NOR2_X1 U53192 ( .A1(n62308), .A2(n47546), .ZN(n47178) );
  NOR2_X1 U53193 ( .A1(n47546), .A2(n8639), .ZN(n47177) );
  NAND2_X1 U53194 ( .A1(n58675), .A2(n65059), .ZN(n47182) );
  NAND4_X1 U53195 ( .A1(n48623), .A2(n3340), .A3(n48619), .A4(n47182), .ZN(
        n47183) );
  NOR2_X1 U53196 ( .A1(n47194), .A2(n47193), .ZN(n47195) );
  NOR2_X1 U53197 ( .A1(n48665), .A2(n48667), .ZN(n48196) );
  NAND2_X1 U53201 ( .A1(n48166), .A2(n64922), .ZN(n47214) );
  AOI21_X1 U53202 ( .A1(n47215), .A2(n47214), .B(n47213), .ZN(n47221) );
  NAND2_X1 U53204 ( .A1(n48518), .A2(n48521), .ZN(n47216) );
  OAI21_X1 U53205 ( .A1(n48254), .A2(n47216), .B(n48632), .ZN(n47217) );
  NOR2_X1 U53207 ( .A1(n50207), .A2(n47222), .ZN(n47224) );
  NAND2_X1 U53208 ( .A1(n47228), .A2(n58009), .ZN(n47230) );
  NOR2_X1 U53212 ( .A1(n47256), .A2(n47255), .ZN(n47257) );
  NOR3_X1 U53213 ( .A1(n47261), .A2(n47260), .A3(n47259), .ZN(n47265) );
  NAND3_X1 U53214 ( .A1(n47592), .A2(n47275), .A3(n47274), .ZN(n47276) );
  NOR2_X1 U53215 ( .A1(n47593), .A2(n47276), .ZN(n47278) );
  OAI21_X1 U53216 ( .A1(n47279), .A2(n47278), .B(n47277), .ZN(n47286) );
  INV_X1 U53217 ( .I(n47280), .ZN(n47585) );
  NAND3_X1 U53218 ( .A1(n47585), .A2(n47281), .A3(n47590), .ZN(n47285) );
  NAND3_X1 U53219 ( .A1(n47283), .A2(n47282), .A3(n22908), .ZN(n47284) );
  NAND3_X1 U53220 ( .A1(n47293), .A2(n47292), .A3(n20666), .ZN(n47300) );
  NOR2_X1 U53221 ( .A1(n47301), .A2(n47296), .ZN(n47294) );
  AOI21_X1 U53223 ( .A1(n47305), .A2(n25477), .B(n47303), .ZN(n47306) );
  AOI21_X1 U53224 ( .A1(n24692), .A2(n49641), .B(n61867), .ZN(n47339) );
  NOR2_X1 U53225 ( .A1(n47312), .A2(n47307), .ZN(n47321) );
  OAI21_X1 U53226 ( .A1(n47310), .A2(n47309), .B(n47308), .ZN(n47311) );
  NAND2_X1 U53227 ( .A1(n47317), .A2(n47329), .ZN(n47318) );
  AOI21_X1 U53230 ( .A1(n47327), .A2(n47326), .B(n47325), .ZN(n47332) );
  NOR3_X1 U53231 ( .A1(n59670), .A2(n47329), .A3(n47328), .ZN(n47331) );
  NOR3_X1 U53232 ( .A1(n2786), .A2(n47332), .A3(n47331), .ZN(n47333) );
  NAND2_X1 U53233 ( .A1(n48726), .A2(n49926), .ZN(n47338) );
  XOR2_X1 U53235 ( .A1(n47341), .A2(n47340), .Z(n47342) );
  XOR2_X1 U53236 ( .A1(n51741), .A2(n47342), .Z(n47352) );
  INV_X1 U53237 ( .I(n49115), .ZN(n47345) );
  NOR2_X1 U53239 ( .A1(n10015), .A2(n23802), .ZN(n49116) );
  NAND3_X1 U53241 ( .A1(n11058), .A2(n60510), .A3(n24788), .ZN(n47353) );
  NAND2_X1 U53242 ( .A1(n7113), .A2(n48064), .ZN(n47357) );
  NAND2_X1 U53246 ( .A1(n47797), .A2(n1481), .ZN(n47384) );
  NOR2_X1 U53248 ( .A1(n47700), .A2(n1657), .ZN(n47387) );
  NOR2_X1 U53250 ( .A1(n47806), .A2(n47797), .ZN(n47390) );
  NAND2_X1 U53252 ( .A1(n47693), .A2(n47706), .ZN(n47392) );
  NOR2_X1 U53255 ( .A1(n47422), .A2(n263), .ZN(n47424) );
  NOR2_X1 U53257 ( .A1(n59205), .A2(n4760), .ZN(n47430) );
  OAI21_X1 U53258 ( .A1(n47433), .A2(n47736), .B(n47432), .ZN(n47441) );
  NAND2_X1 U53260 ( .A1(n47746), .A2(n47434), .ZN(n47439) );
  XOR2_X1 U53262 ( .A1(n23697), .A2(n52617), .Z(n47448) );
  NAND3_X1 U53264 ( .A1(n48301), .A2(n47451), .A3(n47450), .ZN(n47452) );
  OAI22_X1 U53265 ( .A1(n50421), .A2(n57572), .B1(n49244), .B2(n23063), .ZN(
        n47455) );
  AOI21_X1 U53266 ( .A1(n50421), .A2(n57572), .B(n63876), .ZN(n47454) );
  XOR2_X1 U53269 ( .A1(n20332), .A2(n63021), .Z(n47461) );
  XOR2_X1 U53270 ( .A1(n47462), .A2(n47461), .Z(n47757) );
  AOI21_X1 U53272 ( .A1(n10055), .A2(n44065), .B(n47471), .ZN(n47475) );
  INV_X1 U53273 ( .I(n48242), .ZN(n47486) );
  INV_X1 U53274 ( .I(n47493), .ZN(n47497) );
  MUX2_X1 U53275 ( .I0(n47497), .I1(n47496), .S(n10333), .Z(n47523) );
  NAND2_X1 U53276 ( .A1(n47502), .A2(n61146), .ZN(n47498) );
  AOI21_X1 U53277 ( .A1(n47500), .A2(n22899), .B(n47498), .ZN(n47509) );
  NAND2_X1 U53278 ( .A1(n47500), .A2(n47499), .ZN(n47508) );
  NAND2_X1 U53279 ( .A1(n1086), .A2(n47501), .ZN(n47506) );
  NAND2_X1 U53280 ( .A1(n47503), .A2(n47502), .ZN(n47504) );
  MUX2_X1 U53283 ( .I0(n47516), .I1(n47515), .S(n61146), .Z(n47519) );
  OAI21_X1 U53284 ( .A1(n47519), .A2(n61980), .B(n47517), .ZN(n47520) );
  NAND3_X1 U53286 ( .A1(n47535), .A2(n59056), .A3(n47536), .ZN(n47538) );
  NAND3_X1 U53287 ( .A1(n47542), .A2(n22703), .A3(n25481), .ZN(n48629) );
  NAND2_X1 U53288 ( .A1(n48626), .A2(n3340), .ZN(n47539) );
  NAND2_X1 U53290 ( .A1(n47541), .A2(n48625), .ZN(n48607) );
  AOI22_X1 U53291 ( .A1(n47544), .A2(n47543), .B1(n47542), .B2(n48622), .ZN(
        n47551) );
  NOR2_X1 U53293 ( .A1(n3340), .A2(n47546), .ZN(n47547) );
  OAI21_X1 U53294 ( .A1(n47548), .A2(n47547), .B(n48623), .ZN(n47549) );
  OAI21_X1 U53295 ( .A1(n47551), .A2(n47550), .B(n47549), .ZN(n47552) );
  NOR2_X1 U53298 ( .A1(n49508), .A2(n48847), .ZN(n47555) );
  AOI22_X1 U53299 ( .A1(n48283), .A2(n49521), .B1(n61833), .B2(n47555), .ZN(
        n47558) );
  XOR2_X1 U53301 ( .A1(n51788), .A2(n52095), .Z(n47652) );
  INV_X1 U53302 ( .I(n47663), .ZN(n47563) );
  OAI22_X1 U53303 ( .A1(n47564), .A2(n47563), .B1(n47659), .B2(n47562), .ZN(
        n47566) );
  MUX2_X1 U53304 ( .I0(n47570), .I1(n177), .S(n47576), .Z(n47571) );
  NOR2_X1 U53305 ( .A1(n47572), .A2(n1669), .ZN(n47573) );
  NOR2_X2 U53306 ( .A1(n47572), .A2(n47578), .ZN(n47898) );
  INV_X1 U53307 ( .I(n47582), .ZN(n47583) );
  NAND2_X1 U53308 ( .A1(n47586), .A2(n47585), .ZN(n47587) );
  NAND2_X1 U53310 ( .A1(n47591), .A2(n47590), .ZN(n47599) );
  NOR2_X1 U53311 ( .A1(n47593), .A2(n47592), .ZN(n47595) );
  NAND2_X1 U53312 ( .A1(n47606), .A2(n47605), .ZN(n47607) );
  INV_X1 U53314 ( .I(n47608), .ZN(n47613) );
  OAI22_X1 U53316 ( .A1(n64470), .A2(n15360), .B1(n22303), .B2(n1069), .ZN(
        n47620) );
  INV_X1 U53317 ( .I(n47618), .ZN(n47619) );
  OAI21_X1 U53319 ( .A1(n47623), .A2(n13746), .B(n47622), .ZN(n47624) );
  NAND2_X1 U53320 ( .A1(n47625), .A2(n47624), .ZN(n47626) );
  AOI21_X1 U53321 ( .A1(n47879), .A2(n47631), .B(n47721), .ZN(n47632) );
  INV_X1 U53323 ( .I(n47634), .ZN(n47635) );
  NAND2_X1 U53324 ( .A1(n10225), .A2(n14121), .ZN(n47637) );
  NAND2_X1 U53325 ( .A1(n47881), .A2(n47874), .ZN(n47636) );
  INV_X1 U53327 ( .I(n20911), .ZN(n47643) );
  NOR2_X1 U53328 ( .A1(n49096), .A2(n47643), .ZN(n47644) );
  AOI22_X1 U53331 ( .A1(n47648), .A2(n49674), .B1(n49096), .B2(n47647), .ZN(
        n47649) );
  OAI21_X1 U53332 ( .A1(n48707), .A2(n49686), .B(n47649), .ZN(n47650) );
  NOR2_X1 U53333 ( .A1(n57603), .A2(n64944), .ZN(n47654) );
  AOI21_X1 U53334 ( .A1(n47664), .A2(n47838), .B(n22537), .ZN(n47665) );
  OAI21_X1 U53335 ( .A1(n47670), .A2(n7395), .B(n47669), .ZN(n47673) );
  NAND2_X1 U53336 ( .A1(n20912), .A2(n47674), .ZN(n47676) );
  OAI21_X1 U53337 ( .A1(n63465), .A2(n57852), .B(n45267), .ZN(n47681) );
  OAI21_X1 U53338 ( .A1(n47687), .A2(n47691), .B(n47686), .ZN(n47689) );
  NAND2_X1 U53339 ( .A1(n47689), .A2(n47688), .ZN(n47692) );
  NAND2_X1 U53340 ( .A1(n47695), .A2(n47694), .ZN(n47698) );
  OAI21_X1 U53341 ( .A1(n47696), .A2(n47699), .B(n47802), .ZN(n47697) );
  MUX2_X1 U53342 ( .I0(n47698), .I1(n47697), .S(n47811), .Z(n47713) );
  NOR2_X1 U53343 ( .A1(n47700), .A2(n47699), .ZN(n47701) );
  NAND3_X1 U53344 ( .A1(n47703), .A2(n47809), .A3(n47811), .ZN(n47710) );
  OAI22_X1 U53345 ( .A1(n47809), .A2(n47705), .B1(n47798), .B2(n14323), .ZN(
        n47707) );
  INV_X1 U53346 ( .I(n47708), .ZN(n47709) );
  NOR2_X1 U53348 ( .A1(n47714), .A2(n47880), .ZN(n47719) );
  INV_X1 U53349 ( .I(n47726), .ZN(n47878) );
  NOR2_X1 U53350 ( .A1(n47746), .A2(n59008), .ZN(n47733) );
  NOR2_X1 U53351 ( .A1(n47730), .A2(n24081), .ZN(n47731) );
  MUX2_X1 U53352 ( .I0(n47733), .I1(n47732), .S(n47731), .Z(n47734) );
  MUX2_X1 U53356 ( .I0(n49566), .I1(n47753), .S(n18975), .Z(n47756) );
  NAND3_X1 U53358 ( .A1(n24393), .A2(n49172), .A3(n49551), .ZN(n47754) );
  AOI21_X1 U53359 ( .A1(n49547), .A2(n47754), .B(n49570), .ZN(n47755) );
  NAND2_X2 U53360 ( .A1(n47756), .A2(n47755), .ZN(n52334) );
  INV_X1 U53362 ( .I(n47761), .ZN(n47762) );
  INV_X1 U53363 ( .I(n47763), .ZN(n47766) );
  INV_X1 U53364 ( .I(n50437), .ZN(n47765) );
  INV_X1 U53365 ( .I(n47768), .ZN(n47769) );
  NAND2_X1 U53366 ( .A1(n14315), .A2(n24069), .ZN(n48732) );
  NAND2_X1 U53367 ( .A1(n48732), .A2(n63546), .ZN(n47771) );
  MUX2_X1 U53368 ( .I0(n47771), .I1(n47770), .S(n48341), .Z(n47794) );
  OAI21_X1 U53369 ( .A1(n47776), .A2(n47775), .B(n7161), .ZN(n47777) );
  NAND3_X1 U53370 ( .A1(n47779), .A2(n47778), .A3(n47777), .ZN(n47780) );
  AOI21_X1 U53371 ( .A1(n47780), .A2(n24069), .B(n49910), .ZN(n47783) );
  NOR2_X1 U53373 ( .A1(n47787), .A2(n14314), .ZN(n47788) );
  NAND2_X1 U53378 ( .A1(n47837), .A2(n59119), .ZN(n47841) );
  NAND3_X1 U53379 ( .A1(n47839), .A2(n5532), .A3(n47838), .ZN(n47840) );
  NOR2_X1 U53380 ( .A1(n47844), .A2(n60881), .ZN(n47847) );
  NOR2_X1 U53381 ( .A1(n47845), .A2(n24114), .ZN(n47846) );
  NOR2_X1 U53383 ( .A1(n59216), .A2(n47858), .ZN(n47861) );
  INV_X1 U53384 ( .I(n47867), .ZN(n47871) );
  OAI21_X1 U53387 ( .A1(n47879), .A2(n47878), .B(n47877), .ZN(n47891) );
  NAND2_X1 U53388 ( .A1(n10225), .A2(n1387), .ZN(n47888) );
  NAND3_X1 U53389 ( .A1(n47889), .A2(n47888), .A3(n47887), .ZN(n47890) );
  INV_X1 U53391 ( .I(n47896), .ZN(n47897) );
  NOR3_X1 U53392 ( .A1(n47902), .A2(n47901), .A3(n47900), .ZN(n47903) );
  NAND2_X1 U53393 ( .A1(n47906), .A2(n47905), .ZN(n47907) );
  NAND2_X1 U53398 ( .A1(n5283), .A2(n47924), .ZN(n47927) );
  INV_X1 U53399 ( .I(n47925), .ZN(n47926) );
  NAND2_X1 U53400 ( .A1(n15386), .A2(n61355), .ZN(n47929) );
  NAND3_X1 U53401 ( .A1(n47929), .A2(n50373), .A3(n12580), .ZN(n47930) );
  XOR2_X1 U53402 ( .A1(n47936), .A2(n57162), .Z(n47938) );
  XOR2_X1 U53403 ( .A1(n47938), .A2(n47937), .Z(n47939) );
  INV_X1 U53407 ( .I(n49793), .ZN(n47946) );
  AOI21_X1 U53408 ( .A1(n858), .A2(n47946), .B(n47945), .ZN(n47951) );
  NOR2_X1 U53409 ( .A1(n49788), .A2(n1642), .ZN(n47949) );
  NOR2_X1 U53412 ( .A1(n50287), .A2(n18608), .ZN(n50122) );
  INV_X1 U53413 ( .I(n50288), .ZN(n47956) );
  NAND3_X1 U53414 ( .A1(n49890), .A2(n60487), .A3(n58861), .ZN(n47957) );
  NAND2_X1 U53415 ( .A1(n18608), .A2(n60487), .ZN(n48718) );
  MUX2_X1 U53416 ( .I0(n21822), .I1(n47961), .S(n50284), .Z(n47962) );
  OAI21_X1 U53420 ( .A1(n48953), .A2(n22869), .B(n47972), .ZN(n47975) );
  NOR2_X1 U53422 ( .A1(n49777), .A2(n47977), .ZN(n47978) );
  INV_X1 U53423 ( .I(n48423), .ZN(n47980) );
  XOR2_X1 U53424 ( .A1(n48803), .A2(n48421), .Z(n47979) );
  NAND2_X1 U53425 ( .A1(n47982), .A2(n47981), .ZN(n47989) );
  NAND2_X1 U53426 ( .A1(n47986), .A2(n47985), .ZN(n47987) );
  INV_X1 U53427 ( .I(n48346), .ZN(n47991) );
  MUX2_X1 U53428 ( .I0(n1383), .I1(n61362), .S(n1262), .Z(n47993) );
  INV_X1 U53431 ( .I(n49526), .ZN(n48003) );
  NAND2_X1 U53432 ( .A1(n49524), .A2(n48845), .ZN(n48005) );
  NAND2_X1 U53436 ( .A1(n49685), .A2(n49092), .ZN(n48012) );
  NAND2_X1 U53441 ( .A1(n24394), .A2(n49556), .ZN(n48828) );
  OAI21_X1 U53442 ( .A1(n49013), .A2(n64823), .B(n10563), .ZN(n48029) );
  NOR2_X1 U53443 ( .A1(n11641), .A2(n48029), .ZN(n48034) );
  NOR2_X1 U53444 ( .A1(n49014), .A2(n49006), .ZN(n48035) );
  OAI21_X1 U53445 ( .A1(n5629), .A2(n49013), .B(n49019), .ZN(n48037) );
  NOR2_X1 U53447 ( .A1(n48038), .A2(n23738), .ZN(n48041) );
  INV_X1 U53450 ( .I(n48054), .ZN(n48055) );
  NAND2_X1 U53451 ( .A1(n49055), .A2(n49056), .ZN(n48072) );
  MUX2_X1 U53452 ( .I0(n48077), .I1(n10981), .S(n64036), .Z(n48079) );
  AOI21_X1 U53456 ( .A1(n48089), .A2(n57398), .B(n48088), .ZN(n48090) );
  NAND3_X1 U53457 ( .A1(n48104), .A2(n23850), .A3(n48102), .ZN(n48105) );
  NOR2_X1 U53458 ( .A1(n48232), .A2(n64605), .ZN(n49860) );
  INV_X1 U53459 ( .I(n48108), .ZN(n48111) );
  NAND2_X1 U53460 ( .A1(n21178), .A2(n22464), .ZN(n48110) );
  INV_X1 U53461 ( .I(n48113), .ZN(n48114) );
  INV_X1 U53463 ( .I(n48126), .ZN(n48129) );
  NAND2_X1 U53464 ( .A1(n63105), .A2(n60398), .ZN(n48128) );
  AOI21_X1 U53465 ( .A1(n48129), .A2(n48128), .B(n58620), .ZN(n48133) );
  OAI22_X1 U53466 ( .A1(n48462), .A2(n48131), .B1(n48134), .B2(n7186), .ZN(
        n48132) );
  NOR2_X1 U53467 ( .A1(n48133), .A2(n48132), .ZN(n48140) );
  OAI21_X1 U53469 ( .A1(n48138), .A2(n48137), .B(n48136), .ZN(n48139) );
  MUX2_X1 U53470 ( .I0(n49868), .I1(n48142), .S(n50254), .Z(n48173) );
  INV_X1 U53478 ( .I(n49979), .ZN(n48171) );
  OAI21_X1 U53480 ( .A1(n21052), .A2(n64166), .B(n13024), .ZN(n48169) );
  INV_X1 U53481 ( .I(n48174), .ZN(n48175) );
  INV_X1 U53482 ( .I(n48482), .ZN(n48178) );
  AOI21_X1 U53483 ( .A1(n48175), .A2(n48587), .B(n48178), .ZN(n48183) );
  NAND3_X1 U53486 ( .A1(n24185), .A2(n8794), .A3(n48484), .ZN(n48185) );
  NAND3_X1 U53488 ( .A1(n23661), .A2(n22436), .A3(n48667), .ZN(n48192) );
  OAI22_X1 U53489 ( .A1(n48210), .A2(n48200), .B1(n48205), .B2(n48199), .ZN(
        n48201) );
  NAND2_X1 U53490 ( .A1(n48201), .A2(n48665), .ZN(n48202) );
  NOR3_X1 U53492 ( .A1(n48205), .A2(n48667), .A3(n48204), .ZN(n48206) );
  NAND2_X1 U53493 ( .A1(n48209), .A2(n48208), .ZN(n48666) );
  NAND2_X1 U53494 ( .A1(n18757), .A2(n22436), .ZN(n48211) );
  NAND2_X1 U53496 ( .A1(n48219), .A2(n48218), .ZN(n48222) );
  INV_X1 U53497 ( .I(n48220), .ZN(n48221) );
  AOI21_X1 U53498 ( .A1(n48222), .A2(n48221), .B(n48606), .ZN(n48223) );
  NAND2_X1 U53499 ( .A1(n48529), .A2(n48239), .ZN(n48240) );
  NAND3_X1 U53501 ( .A1(n48248), .A2(n48654), .A3(n48659), .ZN(n48250) );
  NAND2_X1 U53507 ( .A1(n48259), .A2(n48511), .ZN(n48262) );
  NAND3_X1 U53508 ( .A1(n48637), .A2(n48631), .A3(n48641), .ZN(n48260) );
  NOR2_X1 U53510 ( .A1(n49131), .A2(n49473), .ZN(n48265) );
  NAND2_X1 U53511 ( .A1(n16336), .A2(n50360), .ZN(n49472) );
  INV_X1 U53512 ( .I(n49472), .ZN(n48268) );
  INV_X1 U53513 ( .I(n48273), .ZN(n48277) );
  NAND2_X1 U53514 ( .A1(n50427), .A2(n48757), .ZN(n48759) );
  INV_X1 U53515 ( .I(n48759), .ZN(n48290) );
  MUX2_X1 U53516 ( .I0(n48292), .I1(n48299), .S(n23238), .Z(n48298) );
  INV_X1 U53518 ( .I(n48302), .ZN(n48303) );
  NAND2_X1 U53520 ( .A1(n49315), .A2(n49308), .ZN(n48312) );
  INV_X1 U53524 ( .I(n48332), .ZN(n48739) );
  INV_X1 U53531 ( .I(n7485), .ZN(n48345) );
  NAND2_X1 U53532 ( .A1(n49760), .A2(n49702), .ZN(n48353) );
  NOR2_X1 U53533 ( .A1(n48349), .A2(n49757), .ZN(n48350) );
  MUX2_X1 U53535 ( .I0(n48353), .I1(n48352), .S(n48885), .Z(n48359) );
  INV_X1 U53539 ( .I(n11458), .ZN(n48914) );
  NOR2_X1 U53541 ( .A1(n11458), .A2(n49276), .ZN(n48365) );
  NAND2_X1 U53542 ( .A1(n57194), .A2(n22457), .ZN(n48363) );
  INV_X1 U53543 ( .I(n48374), .ZN(n48375) );
  NAND2_X1 U53544 ( .A1(n2433), .A2(n25253), .ZN(n48377) );
  NOR2_X1 U53545 ( .A1(n22756), .A2(n58205), .ZN(n48379) );
  XOR2_X1 U53549 ( .A1(n48388), .A2(n48387), .Z(n48389) );
  XOR2_X1 U53550 ( .A1(n21905), .A2(n48389), .Z(n48390) );
  XOR2_X1 U53551 ( .A1(n48390), .A2(n52406), .Z(n48401) );
  NAND2_X1 U53552 ( .A1(n16595), .A2(n6313), .ZN(n48398) );
  XOR2_X1 U53554 ( .A1(n48401), .A2(n9752), .Z(n48402) );
  NAND2_X2 U53556 ( .A1(n54347), .A2(n51863), .ZN(n54349) );
  OAI21_X1 U53559 ( .A1(n48424), .A2(n48423), .B(n48422), .ZN(n48430) );
  INV_X1 U53560 ( .I(n48425), .ZN(n48426) );
  INV_X1 U53561 ( .I(n48792), .ZN(n48429) );
  NAND3_X1 U53562 ( .A1(n49111), .A2(n48434), .A3(n48433), .ZN(n48435) );
  NAND2_X1 U53563 ( .A1(n7271), .A2(n59493), .ZN(n48437) );
  NAND3_X1 U53564 ( .A1(n48439), .A2(n48438), .A3(n48437), .ZN(n48444) );
  NOR3_X1 U53566 ( .A1(n9853), .A2(n48445), .A3(n49013), .ZN(n48447) );
  NOR2_X1 U53567 ( .A1(n48447), .A2(n48446), .ZN(n48452) );
  OAI21_X1 U53568 ( .A1(n48449), .A2(n49007), .B(n48448), .ZN(n48451) );
  AND3_X1 U53569 ( .A1(n48452), .A2(n48451), .A3(n48450), .Z(n48458) );
  NAND2_X1 U53570 ( .A1(n48456), .A2(n48455), .ZN(n48457) );
  NOR2_X1 U53571 ( .A1(n48459), .A2(n60386), .ZN(n48478) );
  NAND2_X1 U53572 ( .A1(n48460), .A2(n60358), .ZN(n48461) );
  INV_X1 U53573 ( .I(n48464), .ZN(n48465) );
  NAND2_X1 U53574 ( .A1(n48468), .A2(n48467), .ZN(n48469) );
  NOR2_X1 U53575 ( .A1(n58620), .A2(n60398), .ZN(n48474) );
  OAI21_X1 U53576 ( .A1(n48484), .A2(n23301), .B(n48482), .ZN(n48485) );
  NAND2_X1 U53577 ( .A1(n48489), .A2(n1659), .ZN(n48493) );
  NAND2_X1 U53579 ( .A1(n48495), .A2(n48642), .ZN(n48497) );
  INV_X1 U53584 ( .I(n48507), .ZN(n48508) );
  NOR2_X1 U53585 ( .A1(n23263), .A2(n48512), .ZN(n48517) );
  NOR2_X1 U53587 ( .A1(n48636), .A2(n48514), .ZN(n48515) );
  OAI22_X1 U53590 ( .A1(n48535), .A2(n48534), .B1(n48533), .B2(n22255), .ZN(
        n48537) );
  NAND2_X1 U53591 ( .A1(n48537), .A2(n22464), .ZN(n48541) );
  NAND2_X1 U53592 ( .A1(n12100), .A2(n19361), .ZN(n48539) );
  OAI21_X1 U53593 ( .A1(n48553), .A2(n48552), .B(n48551), .ZN(n48556) );
  AOI22_X1 U53594 ( .A1(n48561), .A2(n63871), .B1(n697), .B2(n48559), .ZN(
        n48563) );
  NOR2_X1 U53595 ( .A1(n48563), .A2(n48562), .ZN(n48569) );
  NAND2_X1 U53596 ( .A1(n697), .A2(n64859), .ZN(n48565) );
  NAND2_X1 U53597 ( .A1(n48573), .A2(n48572), .ZN(n48574) );
  NAND4_X1 U53598 ( .A1(n1650), .A2(n48576), .A3(n48575), .A4(n48574), .ZN(
        n48578) );
  AOI22_X1 U53600 ( .A1(n178), .A2(n23542), .B1(n48585), .B2(n48584), .ZN(
        n48593) );
  NAND2_X1 U53601 ( .A1(n48587), .A2(n48588), .ZN(n48591) );
  NAND3_X1 U53602 ( .A1(n48589), .A2(n9851), .A3(n23813), .ZN(n48590) );
  INV_X1 U53604 ( .I(n48607), .ZN(n48609) );
  NAND3_X1 U53605 ( .A1(n48610), .A2(n48609), .A3(n48608), .ZN(n48618) );
  NAND3_X1 U53606 ( .A1(n48623), .A2(n3341), .A3(n22635), .ZN(n48615) );
  INV_X1 U53607 ( .I(n48619), .ZN(n48621) );
  NAND4_X1 U53608 ( .A1(n48623), .A2(n48622), .A3(n48621), .A4(n48620), .ZN(
        n48628) );
  NAND3_X1 U53609 ( .A1(n48626), .A2(n22635), .A3(n48624), .ZN(n48627) );
  INV_X1 U53610 ( .I(n48666), .ZN(n48671) );
  OAI21_X1 U53611 ( .A1(n49759), .A2(n49697), .B(n49757), .ZN(n48679) );
  AOI22_X1 U53612 ( .A1(n49700), .A2(n48680), .B1(n22157), .B2(n19302), .ZN(
        n48681) );
  AOI21_X1 U53613 ( .A1(n48684), .A2(n16024), .B(n48688), .ZN(n48686) );
  OAI21_X1 U53614 ( .A1(n49057), .A2(n48689), .B(n13554), .ZN(n48694) );
  NAND2_X1 U53615 ( .A1(n49050), .A2(n48691), .ZN(n48692) );
  NAND2_X1 U53616 ( .A1(n17334), .A2(n17335), .ZN(n48858) );
  NAND2_X1 U53617 ( .A1(n49491), .A2(n17335), .ZN(n48698) );
  NAND2_X1 U53618 ( .A1(n9177), .A2(n48701), .ZN(n48702) );
  AOI21_X1 U53619 ( .A1(n48863), .A2(n48702), .B(n23500), .ZN(n49236) );
  NOR2_X1 U53621 ( .A1(n48711), .A2(n49676), .ZN(n49675) );
  OAI21_X1 U53622 ( .A1(n49673), .A2(n16922), .B(n49684), .ZN(n48712) );
  OAI21_X1 U53623 ( .A1(n48713), .A2(n20971), .B(n49370), .ZN(n48714) );
  INV_X1 U53626 ( .I(n50121), .ZN(n48722) );
  NAND2_X1 U53630 ( .A1(n1641), .A2(n6130), .ZN(n48727) );
  INV_X1 U53631 ( .I(n49909), .ZN(n48731) );
  NOR2_X1 U53632 ( .A1(n13839), .A2(n25812), .ZN(n48738) );
  NOR2_X1 U53633 ( .A1(n13614), .A2(n22694), .ZN(n49950) );
  NAND3_X1 U53634 ( .A1(n11623), .A2(n24374), .A3(n61624), .ZN(n48740) );
  XOR2_X1 U53635 ( .A1(n48747), .A2(n52080), .Z(n48749) );
  XOR2_X1 U53636 ( .A1(n48749), .A2(n48748), .Z(n48750) );
  XOR2_X1 U53637 ( .A1(n52420), .A2(n48750), .Z(n48751) );
  XOR2_X1 U53638 ( .A1(n51762), .A2(n48751), .Z(n48752) );
  NAND3_X1 U53641 ( .A1(n63876), .A2(n57572), .A3(n22533), .ZN(n48758) );
  INV_X1 U53645 ( .I(n48768), .ZN(n48769) );
  NOR2_X1 U53646 ( .A1(n18185), .A2(n48771), .ZN(n48772) );
  INV_X1 U53647 ( .I(n48919), .ZN(n48775) );
  INV_X1 U53649 ( .I(n48779), .ZN(n48780) );
  NAND2_X1 U53652 ( .A1(n49377), .A2(n9983), .ZN(n49429) );
  OAI21_X1 U53653 ( .A1(n48906), .A2(n49429), .B(n49376), .ZN(n48785) );
  NAND2_X1 U53654 ( .A1(n49528), .A2(n49538), .ZN(n48783) );
  NOR2_X1 U53656 ( .A1(n48785), .A2(n48784), .ZN(n48786) );
  NOR3_X1 U53660 ( .A1(n48794), .A2(n48793), .A3(n48792), .ZN(n48795) );
  INV_X1 U53661 ( .I(n48798), .ZN(n48800) );
  NOR3_X1 U53663 ( .A1(n48804), .A2(n48803), .A3(n48811), .ZN(n48805) );
  INV_X1 U53665 ( .I(n48808), .ZN(n48814) );
  NOR2_X1 U53667 ( .A1(n48823), .A2(n48822), .ZN(n48824) );
  NAND2_X1 U53668 ( .A1(n48828), .A2(n49547), .ZN(n48830) );
  INV_X1 U53670 ( .I(n49555), .ZN(n48833) );
  NAND2_X1 U53671 ( .A1(n48833), .A2(n48832), .ZN(n48834) );
  INV_X1 U53672 ( .I(n48838), .ZN(n48839) );
  NAND2_X1 U53673 ( .A1(n48840), .A2(n49525), .ZN(n48842) );
  OAI21_X1 U53676 ( .A1(n58975), .A2(n49195), .B(n48848), .ZN(n48850) );
  OAI22_X1 U53677 ( .A1(n48855), .A2(n17334), .B1(n64335), .B2(n48854), .ZN(
        n48856) );
  NOR2_X1 U53678 ( .A1(n48858), .A2(n6704), .ZN(n48860) );
  NAND2_X1 U53679 ( .A1(n48863), .A2(n17335), .ZN(n48864) );
  AOI21_X1 U53680 ( .A1(n48864), .A2(n49488), .B(n49300), .ZN(n48865) );
  OAI21_X1 U53681 ( .A1(n49389), .A2(n49325), .B(n48870), .ZN(n48867) );
  NOR2_X1 U53682 ( .A1(n48867), .A2(n48873), .ZN(n48881) );
  OAI21_X1 U53683 ( .A1(n48869), .A2(n49398), .B(n49395), .ZN(n48872) );
  OAI21_X1 U53684 ( .A1(n49331), .A2(n63725), .B(n48875), .ZN(n48879) );
  INV_X1 U53685 ( .I(n7078), .ZN(n48877) );
  NOR2_X1 U53688 ( .A1(n48898), .A2(n49698), .ZN(n48884) );
  NAND2_X1 U53689 ( .A1(n49759), .A2(n49702), .ZN(n49756) );
  INV_X1 U53690 ( .I(n49756), .ZN(n48887) );
  INV_X1 U53691 ( .I(n48885), .ZN(n48886) );
  INV_X1 U53692 ( .I(n48892), .ZN(n48896) );
  NOR2_X1 U53693 ( .A1(n48893), .A2(n49702), .ZN(n48895) );
  AOI22_X1 U53694 ( .A1(n48896), .A2(n58306), .B1(n48895), .B2(n48894), .ZN(
        n48900) );
  OAI21_X1 U53696 ( .A1(n49533), .A2(n48902), .B(n7358), .ZN(n48903) );
  NOR2_X1 U53697 ( .A1(n18769), .A2(n49374), .ZN(n48909) );
  NAND2_X1 U53698 ( .A1(n48907), .A2(n49377), .ZN(n48908) );
  INV_X1 U53699 ( .I(n48923), .ZN(n48915) );
  NAND3_X1 U53700 ( .A1(n48916), .A2(n48915), .A3(n48914), .ZN(n48937) );
  INV_X1 U53701 ( .I(n48917), .ZN(n48918) );
  OAI22_X1 U53702 ( .A1(n49278), .A2(n48919), .B1(n48918), .B2(n1633), .ZN(
        n48922) );
  NAND2_X1 U53703 ( .A1(n57194), .A2(n16986), .ZN(n48920) );
  AOI21_X1 U53704 ( .A1(n62200), .A2(n48925), .B(n48920), .ZN(n48921) );
  NOR2_X1 U53705 ( .A1(n48922), .A2(n48921), .ZN(n48936) );
  NOR2_X1 U53706 ( .A1(n11458), .A2(n48930), .ZN(n48933) );
  INV_X1 U53707 ( .I(n48931), .ZN(n48932) );
  NAND2_X1 U53709 ( .A1(n50039), .A2(n3335), .ZN(n48943) );
  NAND2_X1 U53710 ( .A1(n50049), .A2(n50044), .ZN(n48942) );
  XOR2_X1 U53712 ( .A1(n4311), .A2(n48954), .Z(n48955) );
  OAI21_X1 U53713 ( .A1(n48958), .A2(n49409), .B(n49176), .ZN(n48959) );
  XOR2_X1 U53714 ( .A1(n48968), .A2(n48967), .Z(n48969) );
  INV_X1 U53716 ( .I(n49854), .ZN(n48971) );
  MUX2_X1 U53717 ( .I0(n48972), .I1(n48971), .S(n61070), .Z(n48990) );
  INV_X1 U53718 ( .I(n49856), .ZN(n48974) );
  AOI21_X1 U53719 ( .A1(n48974), .A2(n48973), .B(n49843), .ZN(n48989) );
  NAND3_X1 U53720 ( .A1(n48976), .A2(n25253), .A3(n48975), .ZN(n48978) );
  INV_X1 U53722 ( .I(n48984), .ZN(n48985) );
  NOR2_X1 U53723 ( .A1(n49602), .A2(n49318), .ZN(n48991) );
  AOI21_X1 U53724 ( .A1(n48992), .A2(n48991), .B(n49314), .ZN(n49002) );
  NOR3_X1 U53725 ( .A1(n49313), .A2(n8129), .A3(n25032), .ZN(n48995) );
  INV_X1 U53728 ( .I(n49000), .ZN(n49001) );
  NAND2_X1 U53729 ( .A1(n49006), .A2(n64823), .ZN(n49008) );
  NAND2_X1 U53730 ( .A1(n23581), .A2(n49014), .ZN(n49016) );
  INV_X1 U53731 ( .I(n49729), .ZN(n49023) );
  INV_X1 U53732 ( .I(n49419), .ZN(n49024) );
  NOR2_X1 U53733 ( .A1(n21183), .A2(n7494), .ZN(n49027) );
  OAI22_X1 U53734 ( .A1(n49030), .A2(n49425), .B1(n50408), .B2(n50083), .ZN(
        n49026) );
  INV_X1 U53735 ( .I(n49029), .ZN(n49031) );
  OAI21_X1 U53736 ( .A1(n49031), .A2(n49030), .B(n50075), .ZN(n49034) );
  AOI21_X1 U53737 ( .A1(n25944), .A2(n59021), .B(n50079), .ZN(n49032) );
  NAND2_X1 U53738 ( .A1(n50407), .A2(n50394), .ZN(n50080) );
  OAI22_X1 U53739 ( .A1(n49032), .A2(n50080), .B1(n50408), .B2(n50412), .ZN(
        n49033) );
  INV_X1 U53740 ( .I(n50097), .ZN(n49036) );
  INV_X1 U53741 ( .I(n49038), .ZN(n49042) );
  NAND2_X1 U53744 ( .A1(n23707), .A2(n50093), .ZN(n49044) );
  NOR2_X1 U53745 ( .A1(n49055), .A2(n1474), .ZN(n49058) );
  INV_X1 U53747 ( .I(n49062), .ZN(n49828) );
  NOR2_X1 U53749 ( .A1(n49071), .A2(n63954), .ZN(n49082) );
  NOR2_X1 U53750 ( .A1(n49073), .A2(n11950), .ZN(n49081) );
  NAND2_X2 U53752 ( .A1(n49084), .A2(n49083), .ZN(n52465) );
  OAI21_X1 U53753 ( .A1(n54026), .A2(n4564), .B(n54028), .ZN(n49085) );
  NAND2_X1 U53754 ( .A1(n54348), .A2(n51863), .ZN(n49087) );
  NAND2_X1 U53755 ( .A1(n51860), .A2(n11207), .ZN(n53030) );
  INV_X1 U53756 ( .I(n53030), .ZN(n53037) );
  NAND2_X1 U53757 ( .A1(n53037), .A2(n53881), .ZN(n49086) );
  OAI22_X1 U53758 ( .A1(n49093), .A2(n49682), .B1(n49677), .B2(n49092), .ZN(
        n49094) );
  AOI21_X1 U53760 ( .A1(n49677), .A2(n49674), .B(n49673), .ZN(n49097) );
  NAND2_X1 U53762 ( .A1(n13537), .A2(n7588), .ZN(n49104) );
  NAND4_X1 U53763 ( .A1(n20708), .A2(n49107), .A3(n49106), .A4(n49803), .ZN(
        n49108) );
  OAI22_X1 U53764 ( .A1(n49116), .A2(n49115), .B1(n59493), .B2(n7146), .ZN(
        n49118) );
  XOR2_X1 U53765 ( .A1(n50769), .A2(n1573), .Z(n51941) );
  XOR2_X1 U53766 ( .A1(n49122), .A2(n51530), .Z(n49123) );
  XOR2_X1 U53767 ( .A1(n49123), .A2(n50190), .Z(n49124) );
  XOR2_X1 U53768 ( .A1(n65143), .A2(n49124), .Z(n49125) );
  OAI21_X1 U53770 ( .A1(n50002), .A2(n49476), .B(n49139), .ZN(n49140) );
  NOR2_X1 U53772 ( .A1(n50296), .A2(n22717), .ZN(n50140) );
  INV_X1 U53773 ( .I(n50140), .ZN(n49144) );
  INV_X1 U53774 ( .I(n49145), .ZN(n49146) );
  AND2_X1 U53776 ( .A1(n49155), .A2(n49154), .Z(n49156) );
  NAND2_X1 U53777 ( .A1(n49158), .A2(n49751), .ZN(n49164) );
  INV_X1 U53778 ( .I(n49225), .ZN(n49161) );
  NAND2_X1 U53779 ( .A1(n49161), .A2(n49221), .ZN(n49162) );
  NAND4_X2 U53780 ( .A1(n49165), .A2(n49164), .A3(n49163), .A4(n49162), .ZN(
        n51214) );
  NAND2_X1 U53784 ( .A1(n49266), .A2(n49177), .ZN(n49178) );
  INV_X1 U53786 ( .I(n49268), .ZN(n49182) );
  AOI21_X1 U53787 ( .A1(n49182), .A2(n49181), .B(n65208), .ZN(n49183) );
  NOR2_X1 U53788 ( .A1(n49184), .A2(n49183), .ZN(n49187) );
  INV_X1 U53789 ( .I(n10461), .ZN(n49188) );
  XOR2_X1 U53791 ( .A1(n57644), .A2(n51203), .Z(n49190) );
  NOR2_X1 U53792 ( .A1(n49195), .A2(n64170), .ZN(n49196) );
  INV_X1 U53793 ( .I(n49197), .ZN(n49198) );
  OAI21_X1 U53795 ( .A1(n7078), .A2(n49211), .B(n49330), .ZN(n49220) );
  OAI21_X1 U53796 ( .A1(n10456), .A2(n617), .B(n49215), .ZN(n49219) );
  NOR2_X1 U53797 ( .A1(n49213), .A2(n57949), .ZN(n49214) );
  NAND3_X1 U53799 ( .A1(n49216), .A2(n49215), .A3(n49323), .ZN(n49217) );
  XOR2_X1 U53800 ( .A1(n51615), .A2(n52429), .Z(n49231) );
  NAND2_X1 U53802 ( .A1(n59966), .A2(n49741), .ZN(n49228) );
  XOR2_X1 U53803 ( .A1(n49233), .A2(n49232), .Z(n49235) );
  AOI21_X1 U53804 ( .A1(n49237), .A2(n49236), .B(n49235), .ZN(n49234) );
  INV_X1 U53805 ( .I(n49234), .ZN(n49239) );
  NAND3_X1 U53806 ( .A1(n49237), .A2(n49236), .A3(n49235), .ZN(n49238) );
  NAND2_X1 U53807 ( .A1(n49239), .A2(n49238), .ZN(n49240) );
  NAND3_X1 U53810 ( .A1(n2878), .A2(n49244), .A3(n50427), .ZN(n49247) );
  INV_X1 U53813 ( .I(n49249), .ZN(n49250) );
  NOR2_X1 U53814 ( .A1(n49256), .A2(n49250), .ZN(n49251) );
  NOR2_X1 U53815 ( .A1(n49252), .A2(n49251), .ZN(n49259) );
  INV_X1 U53816 ( .I(n49260), .ZN(n49261) );
  NAND3_X1 U53817 ( .A1(n49283), .A2(n49286), .A3(n49281), .ZN(n49282) );
  XOR2_X1 U53819 ( .A1(n50196), .A2(n49289), .Z(n49290) );
  XOR2_X1 U53820 ( .A1(n49290), .A2(n51913), .Z(n49291) );
  XOR2_X1 U53821 ( .A1(n49292), .A2(n49291), .Z(n49293) );
  XOR2_X1 U53822 ( .A1(n51313), .A2(n49293), .Z(n49294) );
  NAND2_X1 U53824 ( .A1(n49308), .A2(n49610), .ZN(n49605) );
  NOR2_X1 U53825 ( .A1(n49613), .A2(n49309), .ZN(n49310) );
  NAND2_X1 U53826 ( .A1(n49319), .A2(n49318), .ZN(n49320) );
  NOR2_X1 U53828 ( .A1(n49325), .A2(n49395), .ZN(n49327) );
  NOR2_X1 U53829 ( .A1(n61513), .A2(n15753), .ZN(n49328) );
  AOI22_X1 U53830 ( .A1(n49330), .A2(n49329), .B1(n49394), .B2(n49328), .ZN(
        n49334) );
  NAND2_X1 U53831 ( .A1(n49331), .A2(n63725), .ZN(n49333) );
  AOI22_X1 U53833 ( .A1(n49339), .A2(n61846), .B1(n18249), .B2(n49338), .ZN(
        n49342) );
  NAND2_X1 U53834 ( .A1(n49340), .A2(n58648), .ZN(n49341) );
  NAND2_X1 U53836 ( .A1(n49347), .A2(n49346), .ZN(n49352) );
  NAND3_X1 U53837 ( .A1(n50221), .A2(n50216), .A3(n14931), .ZN(n49349) );
  AOI21_X1 U53838 ( .A1(n49350), .A2(n49349), .B(n64751), .ZN(n49351) );
  NAND2_X1 U53839 ( .A1(n50044), .A2(n3348), .ZN(n49357) );
  NOR2_X1 U53840 ( .A1(n49371), .A2(n49671), .ZN(n49373) );
  OAI21_X1 U53842 ( .A1(n61513), .A2(n49382), .B(n63725), .ZN(n49387) );
  AOI21_X1 U53843 ( .A1(n49383), .A2(n49389), .B(n49393), .ZN(n49386) );
  NOR3_X1 U53846 ( .A1(n22509), .A2(n49393), .A3(n8604), .ZN(n49399) );
  NOR2_X1 U53847 ( .A1(n15753), .A2(n49395), .ZN(n49396) );
  XOR2_X1 U53848 ( .A1(n50955), .A2(n49401), .Z(n49402) );
  XOR2_X1 U53849 ( .A1(n50712), .A2(n49402), .Z(n49404) );
  XOR2_X1 U53850 ( .A1(n49404), .A2(n49403), .Z(n49405) );
  XOR2_X1 U53851 ( .A1(n9752), .A2(n49413), .Z(n49414) );
  XOR2_X1 U53852 ( .A1(n49415), .A2(n49416), .Z(n53222) );
  NAND2_X1 U53853 ( .A1(n60833), .A2(n533), .ZN(n49628) );
  NAND2_X1 U53856 ( .A1(n19773), .A2(n3335), .ZN(n49576) );
  INV_X1 U53857 ( .I(n49576), .ZN(n49438) );
  INV_X1 U53858 ( .I(n49440), .ZN(n49443) );
  NAND2_X1 U53859 ( .A1(n50049), .A2(n20199), .ZN(n49442) );
  OAI22_X1 U53860 ( .A1(n49443), .A2(n49442), .B1(n49581), .B2(n50040), .ZN(
        n49444) );
  XOR2_X1 U53861 ( .A1(n49446), .A2(n49445), .Z(n49447) );
  XOR2_X1 U53862 ( .A1(n49448), .A2(n49447), .Z(n49449) );
  NOR2_X1 U53863 ( .A1(n61716), .A2(n2433), .ZN(n49845) );
  INV_X1 U53864 ( .I(n49845), .ZN(n49455) );
  NAND2_X1 U53869 ( .A1(n49472), .A2(n49471), .ZN(n49475) );
  INV_X1 U53871 ( .I(n65245), .ZN(n49483) );
  OAI22_X1 U53872 ( .A1(n49483), .A2(n49482), .B1(n6704), .B2(n64341), .ZN(
        n49485) );
  INV_X1 U53873 ( .I(n49487), .ZN(n49489) );
  NOR3_X1 U53874 ( .A1(n49489), .A2(n17334), .A3(n49488), .ZN(n49492) );
  NAND2_X1 U53875 ( .A1(n49501), .A2(n6704), .ZN(n49505) );
  INV_X1 U53876 ( .I(n49502), .ZN(n49503) );
  OAI21_X1 U53880 ( .A1(n49534), .A2(n49533), .B(n49532), .ZN(n49535) );
  NAND2_X1 U53881 ( .A1(n49543), .A2(n49542), .ZN(n49544) );
  NOR4_X1 U53882 ( .A1(n49551), .A2(n22571), .A3(n24394), .A4(n49547), .ZN(
        n49554) );
  AOI21_X1 U53883 ( .A1(n49567), .A2(n25128), .B(n49566), .ZN(n49568) );
  XOR2_X1 U53884 ( .A1(n52154), .A2(n24025), .Z(n49571) );
  NAND2_X1 U53887 ( .A1(n50049), .A2(n50043), .ZN(n49579) );
  AOI21_X1 U53888 ( .A1(n49581), .A2(n49580), .B(n49579), .ZN(n49585) );
  NAND2_X1 U53889 ( .A1(n19773), .A2(n1637), .ZN(n49583) );
  OAI22_X1 U53890 ( .A1(n50044), .A2(n50046), .B1(n3347), .B2(n49583), .ZN(
        n49584) );
  XOR2_X1 U53891 ( .A1(n49589), .A2(n49588), .Z(n49590) );
  XOR2_X1 U53892 ( .A1(n15096), .A2(n49590), .Z(n49591) );
  XOR2_X1 U53893 ( .A1(n49591), .A2(n10584), .Z(n49623) );
  XOR2_X1 U53897 ( .A1(n49625), .A2(n49624), .Z(n49626) );
  NAND3_X1 U53898 ( .A1(n49628), .A2(n52998), .A3(n49627), .ZN(n49629) );
  AND2_X2 U53900 ( .A1(n9616), .A2(n53740), .Z(n53709) );
  MUX2_X1 U53901 ( .I0(n49633), .I1(n49632), .S(n10958), .Z(n49646) );
  XOR2_X1 U53902 ( .A1(n49635), .A2(n1636), .Z(n49640) );
  XOR2_X1 U53904 ( .A1(n10958), .A2(n502), .Z(n49638) );
  NAND3_X1 U53905 ( .A1(n49640), .A2(n49639), .A3(n49638), .ZN(n49645) );
  NAND2_X1 U53906 ( .A1(n49642), .A2(n49641), .ZN(n49643) );
  NAND2_X1 U53907 ( .A1(n49659), .A2(n50143), .ZN(n49647) );
  MUX2_X1 U53908 ( .I0(n49647), .I1(n50313), .S(n4699), .Z(n49654) );
  INV_X1 U53909 ( .I(n50059), .ZN(n49648) );
  NOR4_X1 U53910 ( .A1(n50309), .A2(n1643), .A3(n3054), .A4(n9646), .ZN(n49651) );
  OAI21_X1 U53911 ( .A1(n49651), .A2(n49650), .B(n50304), .ZN(n49652) );
  OAI21_X1 U53912 ( .A1(n49657), .A2(n9646), .B(n49656), .ZN(n49665) );
  OAI21_X1 U53913 ( .A1(n50304), .A2(n3055), .B(n50297), .ZN(n49664) );
  NOR2_X1 U53914 ( .A1(n50308), .A2(n50142), .ZN(n49658) );
  OAI22_X1 U53915 ( .A1(n49659), .A2(n49658), .B1(n60397), .B2(n50143), .ZN(
        n49662) );
  XOR2_X1 U53918 ( .A1(n51165), .A2(n55118), .Z(n49666) );
  XOR2_X1 U53919 ( .A1(n49667), .A2(n49666), .Z(n49668) );
  XOR2_X1 U53920 ( .A1(n49669), .A2(n49668), .Z(n49670) );
  NAND2_X1 U53921 ( .A1(n49685), .A2(n49684), .ZN(n49688) );
  XOR2_X1 U53922 ( .A1(n49691), .A2(n51686), .Z(n49692) );
  OAI21_X1 U53923 ( .A1(n22646), .A2(n24073), .B(n49694), .ZN(n49696) );
  NOR2_X1 U53924 ( .A1(n49762), .A2(n49702), .ZN(n49695) );
  XOR2_X1 U53925 ( .A1(n49708), .A2(n23670), .Z(n49716) );
  NAND3_X1 U53926 ( .A1(n49712), .A2(n49711), .A3(n14561), .ZN(n49713) );
  XOR2_X1 U53927 ( .A1(n51744), .A2(n49716), .Z(n49719) );
  XOR2_X1 U53928 ( .A1(n50582), .A2(n16984), .Z(n49717) );
  XOR2_X1 U53929 ( .A1(n49717), .A2(n24076), .Z(n49718) );
  NOR2_X1 U53930 ( .A1(n49729), .A2(n50074), .ZN(n49730) );
  XNOR2_X1 U53931 ( .A1(n57162), .A2(n53124), .ZN(n49734) );
  XOR2_X1 U53932 ( .A1(n49735), .A2(n49734), .Z(n49737) );
  XOR2_X1 U53933 ( .A1(n49737), .A2(n49736), .Z(n49738) );
  XOR2_X1 U53934 ( .A1(n52630), .A2(n49738), .Z(n49753) );
  OAI21_X1 U53935 ( .A1(n49743), .A2(n16595), .B(n49742), .ZN(n49744) );
  XOR2_X1 U53936 ( .A1(n49753), .A2(n22577), .Z(n49754) );
  NOR2_X1 U53937 ( .A1(n49762), .A2(n2357), .ZN(n49763) );
  XOR2_X1 U53938 ( .A1(n49767), .A2(n49783), .Z(n49769) );
  NAND2_X1 U53939 ( .A1(n49770), .A2(n21550), .ZN(n49771) );
  NAND2_X1 U53940 ( .A1(n49775), .A2(n49774), .ZN(n49778) );
  MUX2_X1 U53941 ( .I0(n49781), .I1(n49780), .S(n21550), .Z(n49782) );
  XOR2_X1 U53944 ( .A1(n49807), .A2(n49806), .Z(n49808) );
  XOR2_X1 U53945 ( .A1(n64102), .A2(n49808), .Z(n49809) );
  NAND2_X1 U53947 ( .A1(n15929), .A2(n51711), .ZN(n49818) );
  NAND3_X1 U53948 ( .A1(n53880), .A2(n51710), .A3(n49818), .ZN(n49874) );
  NAND3_X1 U53949 ( .A1(n49820), .A2(n49819), .A3(n53868), .ZN(n49873) );
  XOR2_X1 U53950 ( .A1(n49821), .A2(n30036), .Z(n49823) );
  XOR2_X1 U53951 ( .A1(n49823), .A2(n49822), .Z(n49824) );
  XOR2_X1 U53952 ( .A1(n51615), .A2(n49824), .Z(n49825) );
  NOR3_X1 U53953 ( .A1(n49827), .A2(n63954), .A3(n65135), .ZN(n49830) );
  INV_X1 U53954 ( .I(n49831), .ZN(n49834) );
  OAI21_X1 U53955 ( .A1(n61805), .A2(n49836), .B(n49835), .ZN(n49838) );
  XOR2_X1 U53957 ( .A1(n22790), .A2(n12985), .Z(n51830) );
  INV_X1 U53958 ( .I(n49860), .ZN(n49861) );
  NAND2_X1 U53959 ( .A1(n49969), .A2(n50345), .ZN(n49870) );
  AOI21_X1 U53960 ( .A1(n50333), .A2(n13024), .B(n49868), .ZN(n49869) );
  AOI22_X1 U53961 ( .A1(n49870), .A2(n50334), .B1(n22506), .B2(n49869), .ZN(
        n49871) );
  XOR2_X1 U53962 ( .A1(n49875), .A2(n53284), .Z(n49876) );
  XOR2_X1 U53963 ( .A1(n49877), .A2(n49876), .Z(n49878) );
  XOR2_X1 U53964 ( .A1(n4846), .A2(n49878), .Z(n49879) );
  INV_X1 U53965 ( .I(n1471), .ZN(n49886) );
  NOR2_X1 U53966 ( .A1(n49881), .A2(n18607), .ZN(n49883) );
  INV_X1 U53968 ( .I(n49891), .ZN(n49894) );
  NAND2_X1 U53969 ( .A1(n61759), .A2(n18608), .ZN(n49893) );
  NAND2_X1 U53970 ( .A1(n49900), .A2(n49899), .ZN(n49902) );
  NAND4_X1 U53971 ( .A1(n49905), .A2(n63923), .A3(n63546), .A4(n19243), .ZN(
        n49906) );
  MUX2_X1 U53972 ( .I0(n49910), .I1(n22263), .S(n64990), .Z(n49915) );
  NOR2_X1 U53973 ( .A1(n22263), .A2(n49909), .ZN(n49912) );
  NOR2_X1 U53974 ( .A1(n14315), .A2(n49910), .ZN(n49911) );
  OAI21_X1 U53975 ( .A1(n49915), .A2(n49914), .B(n49913), .ZN(n49916) );
  MUX2_X1 U53976 ( .I0(n61867), .I1(n3738), .S(n49918), .Z(n49920) );
  OAI21_X1 U53977 ( .A1(n3065), .A2(n61835), .B(n49924), .ZN(n49928) );
  NAND2_X1 U53978 ( .A1(n3065), .A2(n49926), .ZN(n49927) );
  NAND2_X1 U53981 ( .A1(n53876), .A2(n1158), .ZN(n49932) );
  INV_X1 U53982 ( .I(n49934), .ZN(n49935) );
  NAND2_X1 U53983 ( .A1(n50277), .A2(n13614), .ZN(n49944) );
  INV_X1 U53984 ( .I(n49939), .ZN(n49941) );
  OAI21_X1 U53985 ( .A1(n49942), .A2(n49941), .B(n61624), .ZN(n49943) );
  MUX2_X1 U53986 ( .I0(n49944), .I1(n49943), .S(n57543), .Z(n49954) );
  NAND2_X1 U53987 ( .A1(n22694), .A2(n49948), .ZN(n50276) );
  INV_X1 U53988 ( .I(n50276), .ZN(n49945) );
  INV_X1 U53989 ( .I(n49947), .ZN(n49949) );
  NAND3_X1 U53990 ( .A1(n49950), .A2(n49949), .A3(n61170), .ZN(n49952) );
  XOR2_X1 U53991 ( .A1(n50985), .A2(n49955), .Z(n49956) );
  XOR2_X1 U53992 ( .A1(n49957), .A2(n49956), .Z(n49958) );
  XOR2_X1 U53993 ( .A1(n51625), .A2(n49958), .Z(n49959) );
  XOR2_X1 U53994 ( .A1(n49959), .A2(n52465), .Z(n49961) );
  XOR2_X1 U53995 ( .A1(n24105), .A2(n55516), .Z(n49963) );
  XOR2_X1 U53996 ( .A1(n50498), .A2(n49963), .Z(n49964) );
  XOR2_X1 U53997 ( .A1(n49965), .A2(n49964), .Z(n49966) );
  NAND3_X1 U54000 ( .A1(n50336), .A2(n23414), .A3(n50333), .ZN(n49973) );
  NOR3_X1 U54002 ( .A1(n7098), .A2(n13024), .A3(n13684), .ZN(n49978) );
  XOR2_X1 U54003 ( .A1(n51298), .A2(n16709), .Z(n49985) );
  INV_X1 U54005 ( .I(n49991), .ZN(n49994) );
  NOR3_X1 U54007 ( .A1(n50005), .A2(n50360), .A3(n26208), .ZN(n50007) );
  INV_X1 U54008 ( .I(n61737), .ZN(n50009) );
  XOR2_X1 U54009 ( .A1(n12985), .A2(n50009), .Z(n50010) );
  INV_X1 U54010 ( .I(n50211), .ZN(n50014) );
  OAI21_X1 U54011 ( .A1(n50014), .A2(n62413), .B(n1383), .ZN(n50015) );
  NAND2_X1 U54012 ( .A1(n50015), .A2(n50215), .ZN(n50018) );
  NAND2_X1 U54013 ( .A1(n50016), .A2(n16107), .ZN(n50017) );
  XOR2_X1 U54015 ( .A1(n50026), .A2(n50025), .Z(n50027) );
  XOR2_X1 U54018 ( .A1(n50030), .A2(n23069), .Z(n50031) );
  XOR2_X1 U54019 ( .A1(n50032), .A2(n50660), .Z(n50033) );
  NOR3_X1 U54021 ( .A1(n50047), .A2(n20428), .A3(n50046), .ZN(n50052) );
  INV_X1 U54022 ( .I(n50049), .ZN(n50050) );
  NOR2_X1 U54023 ( .A1(n50050), .A2(n3347), .ZN(n50051) );
  OAI21_X1 U54024 ( .A1(n50056), .A2(n22717), .B(n50055), .ZN(n50057) );
  NOR2_X1 U54025 ( .A1(n50140), .A2(n50141), .ZN(n50062) );
  AOI22_X1 U54026 ( .A1(n60397), .A2(n50307), .B1(n50308), .B2(n9646), .ZN(
        n50063) );
  NAND2_X1 U54027 ( .A1(n50064), .A2(n50063), .ZN(n50065) );
  INV_X1 U54028 ( .I(n62616), .ZN(n50066) );
  XOR2_X1 U54029 ( .A1(n18645), .A2(n51358), .Z(n50072) );
  XOR2_X1 U54030 ( .A1(n50068), .A2(n50067), .Z(n50069) );
  XOR2_X1 U54031 ( .A1(n50072), .A2(n50071), .Z(n50073) );
  MUX2_X1 U54032 ( .I0(n52974), .I1(n57700), .S(n4399), .Z(n50155) );
  INV_X1 U54033 ( .I(n53566), .ZN(n50112) );
  INV_X1 U54034 ( .I(n50410), .ZN(n50078) );
  AOI21_X1 U54035 ( .A1(n21183), .A2(n50397), .B(n50080), .ZN(n50086) );
  NAND2_X1 U54036 ( .A1(n50081), .A2(n50398), .ZN(n50084) );
  INV_X1 U54037 ( .I(n50375), .ZN(n50091) );
  XOR2_X1 U54038 ( .A1(n50102), .A2(n50101), .Z(n50103) );
  XOR2_X1 U54039 ( .A1(n50103), .A2(n10594), .Z(n50104) );
  XOR2_X1 U54040 ( .A1(n50104), .A2(n52165), .Z(n50105) );
  INV_X1 U54041 ( .I(n50107), .ZN(n50108) );
  XOR2_X1 U54042 ( .A1(n24757), .A2(n50109), .Z(n50110) );
  NOR2_X2 U54043 ( .A1(n54058), .A2(n54035), .ZN(n53907) );
  NAND2_X1 U54044 ( .A1(n50112), .A2(n54045), .ZN(n50154) );
  INV_X1 U54045 ( .I(n54046), .ZN(n50152) );
  XOR2_X1 U54046 ( .A1(n20774), .A2(n57131), .Z(n50113) );
  XOR2_X1 U54047 ( .A1(n51790), .A2(n51744), .Z(n50115) );
  OAI21_X1 U54049 ( .A1(n18607), .A2(n21092), .B(n50122), .ZN(n50124) );
  XOR2_X1 U54050 ( .A1(n50126), .A2(n23886), .Z(n50127) );
  XOR2_X1 U54051 ( .A1(n50128), .A2(n50127), .Z(n50130) );
  XOR2_X1 U54052 ( .A1(n50130), .A2(n50129), .Z(n50131) );
  XOR2_X1 U54053 ( .A1(n51788), .A2(n50131), .Z(n50132) );
  XOR2_X1 U54054 ( .A1(n50132), .A2(n62589), .Z(n50133) );
  XOR2_X1 U54055 ( .A1(n51181), .A2(n50133), .Z(n50134) );
  NOR2_X1 U54056 ( .A1(n4699), .A2(n50304), .ZN(n50137) );
  NOR2_X1 U54058 ( .A1(n20763), .A2(n50142), .ZN(n50144) );
  AND2_X1 U54059 ( .A1(n50146), .A2(n50145), .Z(n50147) );
  XOR2_X1 U54060 ( .A1(n50150), .A2(n50149), .Z(n50151) );
  NAND2_X1 U54061 ( .A1(n50152), .A2(n60049), .ZN(n53565) );
  INV_X1 U54062 ( .I(n53565), .ZN(n50153) );
  OAI21_X1 U54063 ( .A1(n50155), .A2(n50154), .B(n50153), .ZN(n50160) );
  NAND2_X1 U54067 ( .A1(n54052), .A2(n53916), .ZN(n53913) );
  NOR2_X1 U54068 ( .A1(n53410), .A2(n53913), .ZN(n50157) );
  NAND2_X2 U54070 ( .A1(n50160), .A2(n50159), .ZN(n53728) );
  INV_X1 U54071 ( .I(n53728), .ZN(n53724) );
  XOR2_X1 U54072 ( .A1(n50162), .A2(n50161), .Z(n50163) );
  XOR2_X1 U54073 ( .A1(n9230), .A2(n56692), .Z(n51932) );
  INV_X1 U54074 ( .I(n24758), .ZN(n50165) );
  XOR2_X1 U54075 ( .A1(n50169), .A2(n50168), .Z(n50170) );
  XOR2_X1 U54076 ( .A1(n22584), .A2(n50170), .Z(n50171) );
  XOR2_X1 U54077 ( .A1(n50174), .A2(n50173), .Z(n50175) );
  XOR2_X1 U54078 ( .A1(n50175), .A2(n52103), .Z(n50176) );
  XOR2_X1 U54079 ( .A1(n50177), .A2(n50176), .Z(n50178) );
  XOR2_X1 U54081 ( .A1(n52587), .A2(n23344), .Z(n50180) );
  XOR2_X1 U54082 ( .A1(n50979), .A2(n50180), .Z(n50185) );
  XOR2_X1 U54083 ( .A1(n50182), .A2(n50181), .Z(n50183) );
  INV_X2 U54084 ( .I(n52743), .ZN(n53532) );
  XOR2_X1 U54085 ( .A1(n23016), .A2(n23022), .Z(n50188) );
  XOR2_X1 U54086 ( .A1(n50190), .A2(n50189), .Z(n50191) );
  XOR2_X1 U54087 ( .A1(n50192), .A2(n50191), .Z(n50193) );
  XNOR2_X1 U54089 ( .A1(n50197), .A2(n50196), .ZN(n50198) );
  XOR2_X1 U54090 ( .A1(n50199), .A2(n50198), .Z(n50200) );
  XOR2_X1 U54091 ( .A1(n4265), .A2(n50200), .Z(n50201) );
  XOR2_X1 U54092 ( .A1(n50202), .A2(n50201), .Z(n50203) );
  XOR2_X1 U54093 ( .A1(n52630), .A2(n51313), .Z(n50204) );
  NAND2_X1 U54094 ( .A1(n53535), .A2(n53178), .ZN(n50205) );
  NOR2_X1 U54095 ( .A1(n50219), .A2(n1383), .ZN(n50225) );
  NOR4_X1 U54096 ( .A1(n50222), .A2(n50221), .A3(n7824), .A4(n50220), .ZN(
        n50223) );
  NAND2_X1 U54097 ( .A1(n50239), .A2(n50238), .ZN(n50241) );
  XOR2_X1 U54098 ( .A1(n63352), .A2(n22747), .Z(n50243) );
  XOR2_X1 U54099 ( .A1(n51590), .A2(n50243), .Z(n50244) );
  XOR2_X1 U54100 ( .A1(n50245), .A2(n56702), .Z(n50246) );
  XOR2_X1 U54101 ( .A1(n50247), .A2(n50246), .Z(n50249) );
  XOR2_X1 U54102 ( .A1(n50249), .A2(n50248), .Z(n50250) );
  XOR2_X1 U54103 ( .A1(n50251), .A2(n50250), .Z(n50252) );
  XOR2_X1 U54104 ( .A1(n52103), .A2(n50252), .Z(n50253) );
  XOR2_X1 U54105 ( .A1(n50625), .A2(n50253), .Z(n50265) );
  NAND2_X1 U54106 ( .A1(n7098), .A2(n23414), .ZN(n50255) );
  OAI21_X1 U54107 ( .A1(n50258), .A2(n50338), .B(n64166), .ZN(n50260) );
  NAND3_X1 U54108 ( .A1(n50263), .A2(n50262), .A3(n50261), .ZN(n50264) );
  NOR2_X1 U54110 ( .A1(n50272), .A2(n22694), .ZN(n50273) );
  XOR2_X1 U54113 ( .A1(n65016), .A2(n50878), .Z(n50317) );
  MUX2_X1 U54114 ( .I0(n22717), .I1(n50294), .S(n50309), .Z(n50300) );
  NAND2_X1 U54116 ( .A1(n50301), .A2(n50304), .ZN(n50302) );
  INV_X1 U54117 ( .I(n50312), .ZN(n50314) );
  XOR2_X1 U54118 ( .A1(n50320), .A2(n50319), .Z(n50321) );
  XOR2_X1 U54119 ( .A1(n50323), .A2(n50322), .Z(n50324) );
  XOR2_X1 U54120 ( .A1(n51313), .A2(n50329), .Z(n50352) );
  AOI21_X1 U54126 ( .A1(n50348), .A2(n13684), .B(n50346), .ZN(n50350) );
  NAND2_X1 U54127 ( .A1(n50354), .A2(n50353), .ZN(n50357) );
  NOR2_X1 U54128 ( .A1(n260), .A2(n23394), .ZN(n50355) );
  XOR2_X1 U54130 ( .A1(n57644), .A2(n52086), .Z(n50386) );
  XOR2_X1 U54131 ( .A1(n50387), .A2(n50386), .Z(n50416) );
  XOR2_X1 U54132 ( .A1(n50389), .A2(n50388), .Z(n50390) );
  XOR2_X1 U54133 ( .A1(n52429), .A2(n50390), .Z(n50391) );
  XOR2_X1 U54134 ( .A1(n50392), .A2(n50391), .Z(n50393) );
  NOR2_X1 U54135 ( .A1(n21183), .A2(n50394), .ZN(n50396) );
  NOR2_X1 U54136 ( .A1(n50397), .A2(n50396), .ZN(n50405) );
  NAND3_X1 U54137 ( .A1(n1381), .A2(n50398), .A3(n7494), .ZN(n50404) );
  NAND2_X1 U54138 ( .A1(n50407), .A2(n7494), .ZN(n50411) );
  INV_X1 U54139 ( .I(n50408), .ZN(n50409) );
  INV_X1 U54140 ( .I(n50414), .ZN(n51092) );
  XOR2_X1 U54141 ( .A1(n50850), .A2(n51092), .Z(n50795) );
  XOR2_X1 U54142 ( .A1(n50416), .A2(n50415), .Z(n53612) );
  NAND2_X1 U54144 ( .A1(n50423), .A2(n23063), .ZN(n50433) );
  NAND2_X1 U54148 ( .A1(n50438), .A2(n50437), .ZN(n50439) );
  AOI22_X1 U54149 ( .A1(n50442), .A2(n50441), .B1(n50440), .B2(n50439), .ZN(
        n50451) );
  NOR3_X1 U54150 ( .A1(n59621), .A2(n60622), .A3(n50444), .ZN(n50449) );
  XOR2_X1 U54151 ( .A1(n52178), .A2(n50655), .Z(n50454) );
  XOR2_X1 U54152 ( .A1(n50454), .A2(n50453), .Z(n50455) );
  XOR2_X1 U54153 ( .A1(n50456), .A2(n50455), .Z(n50457) );
  XOR2_X1 U54154 ( .A1(n52472), .A2(n50457), .Z(n50458) );
  NOR2_X2 U54155 ( .A1(n53860), .A2(n53861), .ZN(n53616) );
  INV_X1 U54156 ( .I(n50461), .ZN(n53428) );
  INV_X1 U54157 ( .I(n53857), .ZN(n50463) );
  INV_X1 U54158 ( .I(n50829), .ZN(n50464) );
  AOI22_X1 U54159 ( .A1(n53709), .A2(n1579), .B1(n17287), .B2(n50464), .ZN(
        n50474) );
  NAND2_X1 U54160 ( .A1(n25117), .A2(n53726), .ZN(n50465) );
  NAND3_X1 U54163 ( .A1(n25117), .A2(n53726), .A3(n63920), .ZN(n50466) );
  NAND3_X1 U54164 ( .A1(n50467), .A2(n50830), .A3(n50466), .ZN(n50473) );
  NOR2_X1 U54165 ( .A1(n53731), .A2(n53716), .ZN(n50469) );
  NOR2_X1 U54166 ( .A1(n17286), .A2(n63920), .ZN(n50468) );
  AOI22_X1 U54167 ( .A1(n50469), .A2(n50829), .B1(n50468), .B2(n53709), .ZN(
        n50472) );
  NAND3_X1 U54169 ( .A1(n17286), .A2(n7240), .A3(n63920), .ZN(n50470) );
  NOR3_X1 U54171 ( .A1(n53532), .A2(n23784), .A3(n58763), .ZN(n50478) );
  XOR2_X1 U54175 ( .A1(n52375), .A2(n50486), .Z(n50487) );
  XOR2_X1 U54176 ( .A1(n50488), .A2(n50487), .Z(n50489) );
  XOR2_X1 U54177 ( .A1(n50490), .A2(n50489), .Z(n50491) );
  XOR2_X1 U54178 ( .A1(n18645), .A2(n50491), .Z(n50492) );
  XOR2_X1 U54179 ( .A1(n50496), .A2(n50495), .Z(n50497) );
  XOR2_X1 U54180 ( .A1(n51035), .A2(n50498), .Z(n50499) );
  XOR2_X1 U54181 ( .A1(n50500), .A2(n25061), .Z(n50501) );
  XOR2_X1 U54182 ( .A1(n51234), .A2(n50502), .Z(n50508) );
  XOR2_X1 U54183 ( .A1(n56065), .A2(n53090), .Z(n50503) );
  XOR2_X1 U54184 ( .A1(n50504), .A2(n50503), .Z(n50506) );
  XOR2_X1 U54185 ( .A1(n50506), .A2(n50505), .Z(n50507) );
  XOR2_X1 U54186 ( .A1(n50508), .A2(n50507), .Z(n50510) );
  XOR2_X1 U54187 ( .A1(n50510), .A2(n50509), .Z(n50511) );
  XOR2_X1 U54188 ( .A1(n21425), .A2(n50511), .Z(n50512) );
  XOR2_X1 U54189 ( .A1(n50513), .A2(n1902), .Z(n50515) );
  XOR2_X1 U54190 ( .A1(n50515), .A2(n50514), .Z(n50516) );
  XOR2_X1 U54191 ( .A1(n50517), .A2(n23288), .Z(n50518) );
  XOR2_X1 U54192 ( .A1(n50523), .A2(n1289), .Z(n50524) );
  XOR2_X1 U54193 ( .A1(n50524), .A2(n50525), .Z(n50532) );
  XOR2_X1 U54194 ( .A1(n50527), .A2(n50526), .Z(n50528) );
  XOR2_X1 U54195 ( .A1(n21905), .A2(n50528), .Z(n50529) );
  NAND2_X1 U54196 ( .A1(n23110), .A2(n20921), .ZN(n50546) );
  XOR2_X1 U54197 ( .A1(n50534), .A2(n50533), .Z(n50535) );
  XOR2_X1 U54198 ( .A1(n50536), .A2(n50535), .Z(n50538) );
  XOR2_X1 U54199 ( .A1(n50538), .A2(n50537), .Z(n50539) );
  XOR2_X1 U54200 ( .A1(n58738), .A2(n50539), .Z(n50540) );
  XOR2_X1 U54201 ( .A1(n50979), .A2(n50670), .Z(n50545) );
  MUX2_X1 U54204 ( .I0(n64657), .I1(n57390), .S(n20982), .Z(n50548) );
  XOR2_X1 U54206 ( .A1(n50551), .A2(n56949), .Z(n50552) );
  XOR2_X1 U54207 ( .A1(n52354), .A2(n50552), .Z(n50553) );
  XOR2_X1 U54208 ( .A1(n50554), .A2(n50553), .Z(n50555) );
  XOR2_X1 U54209 ( .A1(n50948), .A2(n50555), .Z(n50556) );
  XOR2_X1 U54210 ( .A1(n50557), .A2(n50556), .Z(n50558) );
  XOR2_X1 U54211 ( .A1(n5272), .A2(n23022), .Z(n50561) );
  XOR2_X1 U54212 ( .A1(n30036), .A2(n54888), .Z(n50562) );
  XOR2_X1 U54213 ( .A1(n7264), .A2(n50562), .Z(n50563) );
  XOR2_X1 U54214 ( .A1(n50564), .A2(n50563), .Z(n50565) );
  XOR2_X1 U54215 ( .A1(n61423), .A2(n50565), .Z(n50566) );
  XOR2_X1 U54216 ( .A1(n51418), .A2(n50567), .Z(n50568) );
  XOR2_X1 U54219 ( .A1(n7343), .A2(n23762), .Z(n51099) );
  XOR2_X1 U54220 ( .A1(n51541), .A2(n51099), .Z(n50569) );
  XOR2_X1 U54221 ( .A1(n51102), .A2(n50569), .Z(n50570) );
  XOR2_X1 U54222 ( .A1(n50571), .A2(n55876), .Z(n50572) );
  XOR2_X1 U54223 ( .A1(n50578), .A2(n50577), .Z(n50579) );
  XOR2_X1 U54224 ( .A1(n23678), .A2(n50579), .Z(n50580) );
  XOR2_X1 U54226 ( .A1(n57131), .A2(n56322), .Z(n50584) );
  XOR2_X1 U54227 ( .A1(n50585), .A2(n50584), .Z(n50586) );
  XOR2_X1 U54228 ( .A1(n50587), .A2(n50586), .Z(n50588) );
  XOR2_X1 U54229 ( .A1(n20774), .A2(n50588), .Z(n50589) );
  XOR2_X1 U54230 ( .A1(n50589), .A2(n20332), .Z(n50591) );
  XOR2_X1 U54231 ( .A1(n50591), .A2(n50590), .Z(n50592) );
  XOR2_X1 U54232 ( .A1(n50593), .A2(n52563), .Z(n50594) );
  XOR2_X1 U54233 ( .A1(n50596), .A2(n50595), .Z(n50597) );
  XOR2_X1 U54234 ( .A1(n51358), .A2(n50597), .Z(n50598) );
  XOR2_X1 U54235 ( .A1(n50598), .A2(n52630), .Z(n50599) );
  NAND2_X1 U54236 ( .A1(n57070), .A2(n57074), .ZN(n52673) );
  INV_X1 U54238 ( .I(n50602), .ZN(n50604) );
  XOR2_X1 U54240 ( .A1(n50608), .A2(n50607), .Z(n50609) );
  XOR2_X1 U54241 ( .A1(n50618), .A2(n50617), .Z(n50619) );
  XOR2_X1 U54242 ( .A1(n51358), .A2(n50619), .Z(n50620) );
  XOR2_X1 U54243 ( .A1(n50628), .A2(n50627), .Z(n50629) );
  XOR2_X1 U54244 ( .A1(n50629), .A2(n52103), .Z(n50630) );
  XOR2_X1 U54245 ( .A1(n50630), .A2(n22795), .Z(n50631) );
  XOR2_X1 U54246 ( .A1(n24040), .A2(n51298), .Z(n50632) );
  XNOR2_X1 U54247 ( .A1(n50634), .A2(n15710), .ZN(n50635) );
  XOR2_X1 U54248 ( .A1(n50636), .A2(n50635), .Z(n50637) );
  XNOR2_X1 U54249 ( .A1(n50641), .A2(n50640), .ZN(n50642) );
  NAND2_X1 U54250 ( .A1(n53381), .A2(n57192), .ZN(n50671) );
  XOR2_X1 U54251 ( .A1(n23288), .A2(n51261), .Z(n50679) );
  XOR2_X1 U54256 ( .A1(n247), .A2(n53102), .Z(n50651) );
  XOR2_X1 U54257 ( .A1(n50652), .A2(n50651), .Z(n50653) );
  XOR2_X1 U54258 ( .A1(n51625), .A2(n50653), .Z(n50654) );
  XOR2_X1 U54259 ( .A1(n10502), .A2(n50654), .Z(n50657) );
  XOR2_X1 U54260 ( .A1(n22658), .A2(n50655), .Z(n50656) );
  XOR2_X1 U54261 ( .A1(n50661), .A2(n55191), .Z(n50662) );
  XOR2_X1 U54262 ( .A1(n50662), .A2(n52513), .Z(n50663) );
  XOR2_X1 U54263 ( .A1(n50664), .A2(n50663), .Z(n50665) );
  XOR2_X1 U54264 ( .A1(n50666), .A2(n50665), .Z(n50667) );
  INV_X1 U54265 ( .I(n58738), .ZN(n51207) );
  XOR2_X1 U54266 ( .A1(n50668), .A2(n51207), .Z(n50669) );
  AOI21_X1 U54267 ( .A1(n52843), .A2(n50671), .B(n53601), .ZN(n50673) );
  INV_X1 U54270 ( .I(n50676), .ZN(n52847) );
  XOR2_X1 U54271 ( .A1(n50680), .A2(n50679), .Z(n50681) );
  XOR2_X1 U54272 ( .A1(n50684), .A2(n50770), .Z(n50685) );
  XOR2_X1 U54273 ( .A1(n23344), .A2(n1898), .Z(n50687) );
  XOR2_X1 U54274 ( .A1(n50687), .A2(n23762), .Z(n50975) );
  XOR2_X1 U54275 ( .A1(n50688), .A2(n50975), .Z(n50689) );
  XOR2_X1 U54276 ( .A1(n50691), .A2(n50690), .Z(n50692) );
  XOR2_X1 U54277 ( .A1(n18645), .A2(n52537), .Z(n50696) );
  XOR2_X1 U54278 ( .A1(n50696), .A2(n52630), .Z(n50706) );
  XNOR2_X1 U54279 ( .A1(n50697), .A2(n50864), .ZN(n50699) );
  XOR2_X1 U54280 ( .A1(n50699), .A2(n50698), .Z(n50700) );
  XOR2_X1 U54281 ( .A1(n50701), .A2(n50700), .Z(n50702) );
  XOR2_X1 U54282 ( .A1(n51313), .A2(n50702), .Z(n50703) );
  XOR2_X1 U54283 ( .A1(n50704), .A2(n50703), .Z(n50705) );
  XOR2_X1 U54284 ( .A1(n50706), .A2(n50705), .Z(n50707) );
  XOR2_X1 U54285 ( .A1(n6336), .A2(n54208), .Z(n51361) );
  XOR2_X1 U54286 ( .A1(n50710), .A2(n50709), .Z(n50711) );
  XOR2_X1 U54287 ( .A1(n50712), .A2(n50711), .Z(n50713) );
  XOR2_X1 U54288 ( .A1(n21905), .A2(n50713), .Z(n50714) );
  XOR2_X1 U54289 ( .A1(n50720), .A2(n50719), .Z(n50721) );
  XOR2_X1 U54290 ( .A1(n51045), .A2(n50724), .Z(n50725) );
  XOR2_X1 U54291 ( .A1(n50726), .A2(n50725), .Z(n50727) );
  XOR2_X1 U54292 ( .A1(n21425), .A2(n50727), .Z(n50728) );
  XOR2_X1 U54293 ( .A1(n50729), .A2(n50728), .Z(n50731) );
  XOR2_X1 U54294 ( .A1(n50731), .A2(n50730), .Z(n50732) );
  XOR2_X1 U54295 ( .A1(n51788), .A2(n50733), .Z(n50735) );
  XOR2_X1 U54296 ( .A1(n50735), .A2(n50734), .Z(n51341) );
  XOR2_X1 U54297 ( .A1(n50742), .A2(n7744), .Z(n50743) );
  XOR2_X1 U54299 ( .A1(n50746), .A2(n50745), .Z(n50747) );
  XOR2_X1 U54300 ( .A1(n50748), .A2(n50747), .Z(n50749) );
  NAND2_X1 U54301 ( .A1(n50751), .A2(n4908), .ZN(n50760) );
  NAND2_X1 U54302 ( .A1(n50754), .A2(n64167), .ZN(n50757) );
  NAND2_X2 U54303 ( .A1(n50760), .A2(n50759), .ZN(n52335) );
  XOR2_X1 U54304 ( .A1(n50764), .A2(n50763), .Z(n50765) );
  XOR2_X1 U54305 ( .A1(n65143), .A2(n22658), .Z(n50766) );
  XOR2_X1 U54306 ( .A1(n50770), .A2(n52178), .Z(n50771) );
  XOR2_X1 U54307 ( .A1(n50772), .A2(n50771), .Z(n50773) );
  XOR2_X1 U54310 ( .A1(n50776), .A2(n55610), .Z(n50778) );
  XOR2_X1 U54311 ( .A1(n50778), .A2(n50777), .Z(n50779) );
  XOR2_X1 U54312 ( .A1(n17597), .A2(n50779), .Z(n50781) );
  XOR2_X1 U54313 ( .A1(n50782), .A2(n50781), .Z(n50784) );
  XOR2_X1 U54314 ( .A1(n50785), .A2(n50954), .Z(n50786) );
  XOR2_X1 U54315 ( .A1(n50788), .A2(n50787), .Z(n50789) );
  XOR2_X1 U54316 ( .A1(n50790), .A2(n50789), .Z(n50791) );
  XOR2_X1 U54317 ( .A1(n6384), .A2(n50793), .Z(n50794) );
  XOR2_X1 U54319 ( .A1(n50798), .A2(n29407), .Z(n50799) );
  XOR2_X1 U54320 ( .A1(n50800), .A2(n50799), .Z(n50801) );
  XOR2_X1 U54321 ( .A1(n51211), .A2(n50801), .Z(n50802) );
  NOR2_X1 U54323 ( .A1(n23248), .A2(n52786), .ZN(n53206) );
  AOI21_X1 U54324 ( .A1(n53437), .A2(n57050), .B(n53206), .ZN(n50809) );
  NAND2_X1 U54325 ( .A1(n53167), .A2(n53147), .ZN(n50810) );
  NOR2_X1 U54327 ( .A1(n1579), .A2(n25117), .ZN(n50821) );
  NAND2_X1 U54328 ( .A1(n53731), .A2(n53728), .ZN(n53717) );
  NAND2_X1 U54330 ( .A1(n53727), .A2(n53728), .ZN(n53751) );
  AOI22_X1 U54332 ( .A1(n53741), .A2(n17287), .B1(n1579), .B2(n53709), .ZN(
        n50825) );
  OAI21_X1 U54334 ( .A1(n53757), .A2(n53756), .B(n25116), .ZN(n50824) );
  AOI21_X1 U54336 ( .A1(n53731), .A2(n25117), .B(n53752), .ZN(n50822) );
  NAND2_X1 U54337 ( .A1(n53754), .A2(n50822), .ZN(n50823) );
  OAI21_X1 U54338 ( .A1(n53731), .A2(n25011), .B(n50830), .ZN(n50828) );
  XOR2_X1 U54339 ( .A1(n50834), .A2(n54360), .Z(n50835) );
  XOR2_X1 U54340 ( .A1(n50836), .A2(n50835), .Z(n50837) );
  XOR2_X1 U54341 ( .A1(n15096), .A2(n50837), .Z(n50838) );
  XOR2_X1 U54342 ( .A1(n50840), .A2(n51043), .Z(n50841) );
  XOR2_X1 U54343 ( .A1(n50842), .A2(n50841), .Z(n50843) );
  XOR2_X1 U54344 ( .A1(n61518), .A2(n50845), .Z(n50846) );
  XOR2_X1 U54345 ( .A1(n50847), .A2(n50846), .Z(n50848) );
  XOR2_X1 U54346 ( .A1(n51086), .A2(n1625), .Z(n50852) );
  XOR2_X1 U54347 ( .A1(n51154), .A2(n50852), .Z(n50853) );
  XOR2_X1 U54349 ( .A1(n50855), .A2(n51150), .Z(n50856) );
  XOR2_X1 U54350 ( .A1(n50857), .A2(n50856), .Z(n50858) );
  XOR2_X1 U54351 ( .A1(n50859), .A2(n23762), .Z(n50860) );
  XOR2_X1 U54352 ( .A1(n15719), .A2(n50860), .Z(n50861) );
  XOR2_X1 U54353 ( .A1(n50864), .A2(n55903), .Z(n50865) );
  XOR2_X1 U54354 ( .A1(n50866), .A2(n50865), .Z(n50867) );
  XOR2_X1 U54355 ( .A1(n50867), .A2(n52537), .Z(n50868) );
  XOR2_X1 U54356 ( .A1(n63009), .A2(n50870), .Z(n50871) );
  XOR2_X1 U54357 ( .A1(n50871), .A2(n23878), .Z(n51912) );
  XOR2_X1 U54358 ( .A1(n50968), .A2(n51912), .Z(n50872) );
  XOR2_X1 U54359 ( .A1(n50874), .A2(n50873), .Z(n50875) );
  OAI21_X1 U54361 ( .A1(n61213), .A2(n14884), .B(n56225), .ZN(n50880) );
  INV_X1 U54363 ( .I(n55709), .ZN(n50883) );
  XOR2_X1 U54364 ( .A1(n50885), .A2(n55580), .Z(n50886) );
  XOR2_X1 U54365 ( .A1(n50887), .A2(n50886), .Z(n50888) );
  INV_X1 U54367 ( .I(n51629), .ZN(n50890) );
  XOR2_X1 U54368 ( .A1(n50890), .A2(n56335), .Z(n51229) );
  XOR2_X1 U54370 ( .A1(n23991), .A2(n50893), .Z(n51146) );
  XOR2_X1 U54371 ( .A1(n51146), .A2(n50894), .Z(n50895) );
  XOR2_X1 U54372 ( .A1(n56008), .A2(n51881), .Z(n50900) );
  XOR2_X1 U54373 ( .A1(n50901), .A2(n50900), .Z(n50902) );
  XOR2_X1 U54374 ( .A1(n50903), .A2(n50902), .Z(n50904) );
  XOR2_X1 U54375 ( .A1(n52154), .A2(n50904), .Z(n50905) );
  XOR2_X1 U54376 ( .A1(n64316), .A2(n50907), .Z(n50908) );
  XOR2_X1 U54377 ( .A1(n50910), .A2(n50909), .Z(n50911) );
  XOR2_X1 U54378 ( .A1(n50912), .A2(n50911), .Z(n50913) );
  XOR2_X1 U54379 ( .A1(n21425), .A2(n50913), .Z(n50914) );
  XOR2_X1 U54380 ( .A1(n50914), .A2(n22783), .Z(n50915) );
  XOR2_X1 U54381 ( .A1(n50918), .A2(n50917), .Z(n50919) );
  XOR2_X1 U54382 ( .A1(n50924), .A2(n51131), .Z(n50925) );
  XOR2_X1 U54383 ( .A1(n50926), .A2(n50925), .Z(n50927) );
  XOR2_X1 U54384 ( .A1(n62616), .A2(n50929), .Z(n50930) );
  INV_X1 U54385 ( .I(n55910), .ZN(n50931) );
  NAND2_X1 U54386 ( .A1(n55915), .A2(n50932), .ZN(n50933) );
  XOR2_X1 U54387 ( .A1(n50935), .A2(n50934), .Z(n50936) );
  XOR2_X1 U54388 ( .A1(n58738), .A2(n52420), .Z(n50939) );
  XOR2_X1 U54389 ( .A1(n50945), .A2(n50944), .Z(n50946) );
  XOR2_X1 U54390 ( .A1(n52073), .A2(n50946), .Z(n50947) );
  XOR2_X1 U54391 ( .A1(n50956), .A2(n50955), .Z(n50957) );
  XOR2_X1 U54392 ( .A1(n50958), .A2(n50957), .Z(n50959) );
  XOR2_X1 U54393 ( .A1(n50960), .A2(n51194), .Z(n50962) );
  XOR2_X1 U54394 ( .A1(n50962), .A2(n50961), .Z(n50963) );
  XOR2_X1 U54395 ( .A1(n50964), .A2(n50963), .Z(n50965) );
  XOR2_X1 U54396 ( .A1(n52630), .A2(n50965), .Z(n50966) );
  XOR2_X1 U54397 ( .A1(n50970), .A2(n50969), .Z(n50971) );
  XOR2_X1 U54398 ( .A1(n50972), .A2(n50971), .Z(n50973) );
  XOR2_X1 U54399 ( .A1(n50976), .A2(n50975), .Z(n50977) );
  XOR2_X1 U54400 ( .A1(n50978), .A2(n50977), .Z(n50982) );
  XOR2_X1 U54402 ( .A1(n50985), .A2(n50984), .Z(n50986) );
  XOR2_X1 U54403 ( .A1(n50987), .A2(n50986), .Z(n50988) );
  XOR2_X1 U54404 ( .A1(n50990), .A2(n50989), .Z(n50991) );
  XOR2_X1 U54406 ( .A1(n50998), .A2(n51881), .Z(n51000) );
  XOR2_X1 U54407 ( .A1(n51000), .A2(n50999), .Z(n51001) );
  XOR2_X1 U54408 ( .A1(n9753), .A2(n51004), .Z(n51006) );
  XOR2_X1 U54409 ( .A1(n51007), .A2(n51006), .Z(n51008) );
  XOR2_X1 U54410 ( .A1(n51008), .A2(n22783), .Z(n51009) );
  XOR2_X1 U54411 ( .A1(n51009), .A2(n51232), .Z(n51010) );
  XOR2_X1 U54412 ( .A1(n22795), .A2(n52334), .Z(n51013) );
  OAI22_X1 U54413 ( .A1(n10040), .A2(n58050), .B1(n56264), .B2(n3616), .ZN(
        n51015) );
  XOR2_X1 U54415 ( .A1(n51581), .A2(n51019), .Z(n51365) );
  INV_X1 U54416 ( .I(n51020), .ZN(n51023) );
  XOR2_X1 U54417 ( .A1(n51021), .A2(n56475), .Z(n51022) );
  XOR2_X1 U54418 ( .A1(n51023), .A2(n51022), .Z(n51024) );
  XOR2_X1 U54419 ( .A1(n51365), .A2(n51025), .Z(n51026) );
  XOR2_X1 U54420 ( .A1(n52055), .A2(n51026), .Z(n51027) );
  XOR2_X1 U54421 ( .A1(n51030), .A2(n51029), .Z(n51031) );
  XOR2_X1 U54422 ( .A1(n51933), .A2(n51031), .Z(n51520) );
  XOR2_X1 U54423 ( .A1(n51190), .A2(n51520), .Z(n51032) );
  INV_X1 U54424 ( .I(n51033), .ZN(n51034) );
  INV_X1 U54426 ( .I(n51037), .ZN(n51039) );
  XOR2_X1 U54427 ( .A1(n51039), .A2(n51038), .Z(n51040) );
  XOR2_X1 U54428 ( .A1(n15096), .A2(n51040), .Z(n51041) );
  XOR2_X1 U54430 ( .A1(n51046), .A2(n51045), .Z(n51047) );
  XOR2_X1 U54431 ( .A1(n61518), .A2(n51047), .Z(n51049) );
  XOR2_X1 U54433 ( .A1(n51049), .A2(n51048), .Z(n51050) );
  XOR2_X1 U54434 ( .A1(n51797), .A2(n53499), .Z(n51051) );
  INV_X1 U54435 ( .I(n20874), .ZN(n51594) );
  XOR2_X1 U54436 ( .A1(n51051), .A2(n51594), .Z(n52025) );
  XOR2_X1 U54437 ( .A1(n51053), .A2(n51052), .Z(n51054) );
  XOR2_X1 U54439 ( .A1(n51358), .A2(n52537), .Z(n51058) );
  XOR2_X1 U54440 ( .A1(n63041), .A2(n51058), .Z(n51066) );
  INV_X1 U54441 ( .I(n51059), .ZN(n51061) );
  XOR2_X1 U54442 ( .A1(n51061), .A2(n51060), .Z(n51062) );
  XOR2_X1 U54443 ( .A1(n8076), .A2(n51062), .Z(n51063) );
  XOR2_X1 U54444 ( .A1(n51064), .A2(n51063), .Z(n51065) );
  XOR2_X1 U54445 ( .A1(n51066), .A2(n51065), .Z(n51067) );
  XOR2_X1 U54447 ( .A1(n1094), .A2(n51069), .Z(n51078) );
  XOR2_X1 U54448 ( .A1(n51071), .A2(n51070), .Z(n51074) );
  XOR2_X1 U54449 ( .A1(n51072), .A2(n54563), .Z(n51073) );
  XOR2_X1 U54450 ( .A1(n51074), .A2(n51073), .Z(n51075) );
  XOR2_X1 U54451 ( .A1(n52073), .A2(n51075), .Z(n51076) );
  XOR2_X1 U54452 ( .A1(n51076), .A2(n51757), .Z(n51077) );
  INV_X1 U54454 ( .I(n51228), .ZN(n51082) );
  NOR2_X1 U54455 ( .A1(n64345), .A2(n56420), .ZN(n51107) );
  AOI21_X1 U54456 ( .A1(n23165), .A2(n56417), .B(n56635), .ZN(n51106) );
  XOR2_X1 U54457 ( .A1(n22666), .A2(n23069), .Z(n51156) );
  XOR2_X1 U54458 ( .A1(n51087), .A2(n52420), .Z(n51095) );
  INV_X1 U54459 ( .I(n51088), .ZN(n51089) );
  XOR2_X1 U54460 ( .A1(n51089), .A2(n52080), .Z(n51090) );
  XOR2_X1 U54461 ( .A1(n51091), .A2(n51090), .Z(n51093) );
  XOR2_X1 U54462 ( .A1(n51093), .A2(n51092), .Z(n51094) );
  XOR2_X1 U54463 ( .A1(n51095), .A2(n51094), .Z(n51096) );
  INV_X1 U54466 ( .I(n51554), .ZN(n51100) );
  XOR2_X1 U54467 ( .A1(n51100), .A2(n51099), .Z(n51101) );
  XOR2_X1 U54468 ( .A1(n51102), .A2(n51101), .Z(n51103) );
  XOR2_X1 U54469 ( .A1(n51104), .A2(n51103), .Z(n51105) );
  INV_X1 U54471 ( .I(n56214), .ZN(n51114) );
  NAND3_X1 U54472 ( .A1(n51114), .A2(n56205), .A3(n61914), .ZN(n51115) );
  NAND2_X1 U54473 ( .A1(n56213), .A2(n51115), .ZN(n51116) );
  XOR2_X1 U54475 ( .A1(n51122), .A2(n51121), .Z(n51123) );
  XOR2_X1 U54476 ( .A1(n51125), .A2(n51937), .Z(n51126) );
  XOR2_X1 U54477 ( .A1(n51132), .A2(n51131), .Z(n51134) );
  XOR2_X1 U54478 ( .A1(n51133), .A2(n51134), .Z(n51135) );
  XOR2_X1 U54479 ( .A1(n51138), .A2(n51137), .Z(n51139) );
  XOR2_X1 U54481 ( .A1(n51142), .A2(n51141), .Z(n51143) );
  XOR2_X1 U54482 ( .A1(n23288), .A2(n51143), .Z(n51145) );
  XOR2_X1 U54483 ( .A1(n51150), .A2(n51149), .Z(n51151) );
  XOR2_X1 U54484 ( .A1(n51152), .A2(n51151), .Z(n51153) );
  XOR2_X1 U54485 ( .A1(n51154), .A2(n51153), .Z(n51155) );
  XOR2_X1 U54487 ( .A1(n51159), .A2(n51160), .Z(n51161) );
  XOR2_X1 U54488 ( .A1(n51165), .A2(n57096), .Z(n51166) );
  XOR2_X1 U54489 ( .A1(n51167), .A2(n51166), .Z(n51168) );
  XOR2_X1 U54490 ( .A1(n51169), .A2(n51168), .Z(n51170) );
  XOR2_X1 U54491 ( .A1(n9044), .A2(n51170), .Z(n51171) );
  XOR2_X1 U54492 ( .A1(n10344), .A2(n64825), .Z(n51172) );
  XOR2_X1 U54493 ( .A1(n51174), .A2(n51173), .Z(n51175) );
  XOR2_X1 U54494 ( .A1(n21425), .A2(n51175), .Z(n51176) );
  XOR2_X1 U54495 ( .A1(n51177), .A2(n51176), .Z(n51178) );
  XOR2_X1 U54497 ( .A1(n51180), .A2(n52617), .Z(n51792) );
  INV_X1 U54501 ( .I(n51192), .ZN(n51196) );
  XOR2_X1 U54502 ( .A1(n51194), .A2(n51193), .Z(n51195) );
  XOR2_X1 U54503 ( .A1(n51196), .A2(n51195), .Z(n51197) );
  XOR2_X1 U54505 ( .A1(n51205), .A2(n51204), .Z(n51206) );
  XOR2_X1 U54506 ( .A1(n52420), .A2(n51206), .Z(n51208) );
  XOR2_X1 U54507 ( .A1(n51208), .A2(n51207), .Z(n51210) );
  XOR2_X1 U54508 ( .A1(n23991), .A2(n724), .Z(n51225) );
  XOR2_X1 U54509 ( .A1(n22658), .A2(n19202), .Z(n51223) );
  INV_X1 U54510 ( .I(n51215), .ZN(n51220) );
  XOR2_X1 U54511 ( .A1(n51216), .A2(n54917), .Z(n51217) );
  XOR2_X1 U54512 ( .A1(n51218), .A2(n51217), .Z(n51219) );
  XOR2_X1 U54513 ( .A1(n51220), .A2(n51219), .Z(n51221) );
  XOR2_X1 U54514 ( .A1(n52471), .A2(n51221), .Z(n51222) );
  XOR2_X1 U54515 ( .A1(n51223), .A2(n51222), .Z(n51224) );
  XOR2_X1 U54516 ( .A1(n52335), .A2(n21425), .Z(n51334) );
  XOR2_X1 U54517 ( .A1(n51232), .A2(n51231), .Z(n51242) );
  XOR2_X1 U54518 ( .A1(n54734), .A2(n56784), .Z(n51233) );
  XOR2_X1 U54519 ( .A1(n51234), .A2(n51233), .Z(n51236) );
  XOR2_X1 U54520 ( .A1(n51236), .A2(n51235), .Z(n51237) );
  XOR2_X1 U54521 ( .A1(n51238), .A2(n51237), .Z(n51239) );
  XOR2_X1 U54522 ( .A1(n51240), .A2(n24076), .Z(n51241) );
  XOR2_X1 U54523 ( .A1(n51242), .A2(n51241), .Z(n51243) );
  INV_X1 U54524 ( .I(n51244), .ZN(n51245) );
  XOR2_X1 U54525 ( .A1(n51245), .A2(n57096), .Z(n51246) );
  XOR2_X1 U54526 ( .A1(n51247), .A2(n51246), .Z(n51248) );
  XOR2_X1 U54527 ( .A1(n22845), .A2(n51248), .Z(n51249) );
  NAND4_X1 U54530 ( .A1(n56188), .A2(n64438), .A3(n56184), .A4(n56149), .ZN(
        n51260) );
  NAND2_X1 U54531 ( .A1(n56564), .A2(n56567), .ZN(n51262) );
  OAI21_X1 U54533 ( .A1(n56564), .A2(n10183), .B(n51265), .ZN(n51266) );
  NAND2_X1 U54534 ( .A1(n56397), .A2(n56389), .ZN(n51269) );
  XOR2_X1 U54535 ( .A1(n13325), .A2(n52073), .Z(n51283) );
  XOR2_X1 U54536 ( .A1(n51276), .A2(n51275), .Z(n51277) );
  XOR2_X1 U54537 ( .A1(n51278), .A2(n51277), .Z(n51279) );
  XOR2_X1 U54538 ( .A1(n51280), .A2(n51279), .Z(n51281) );
  XOR2_X1 U54539 ( .A1(n52358), .A2(n51281), .Z(n51282) );
  XOR2_X1 U54540 ( .A1(n51283), .A2(n51282), .Z(n51285) );
  XOR2_X1 U54541 ( .A1(n51284), .A2(n51285), .Z(n51287) );
  XOR2_X1 U54542 ( .A1(n51287), .A2(n51286), .Z(n51288) );
  INV_X1 U54543 ( .I(n51290), .ZN(n51291) );
  INV_X1 U54544 ( .I(n23758), .ZN(n51292) );
  INV_X1 U54545 ( .I(n51294), .ZN(n51296) );
  XOR2_X1 U54546 ( .A1(n24044), .A2(n54870), .Z(n51295) );
  XOR2_X1 U54547 ( .A1(n51296), .A2(n51295), .Z(n51297) );
  XOR2_X1 U54548 ( .A1(n51385), .A2(n51297), .Z(n51300) );
  XOR2_X1 U54549 ( .A1(n22845), .A2(n51298), .Z(n51299) );
  XOR2_X1 U54550 ( .A1(n51300), .A2(n51299), .Z(n51301) );
  INV_X1 U54551 ( .I(n51304), .ZN(n51306) );
  XOR2_X1 U54552 ( .A1(n51306), .A2(n51305), .Z(n51307) );
  INV_X1 U54554 ( .I(n51309), .ZN(n51311) );
  XOR2_X1 U54555 ( .A1(n51310), .A2(n51311), .Z(n51312) );
  XOR2_X1 U54556 ( .A1(n51313), .A2(n51312), .Z(n51314) );
  XOR2_X1 U54557 ( .A1(n25415), .A2(n51314), .Z(n51315) );
  XOR2_X1 U54558 ( .A1(n52420), .A2(n12985), .Z(n51326) );
  XOR2_X1 U54559 ( .A1(n51321), .A2(n55765), .Z(n51322) );
  XOR2_X1 U54560 ( .A1(n51323), .A2(n51322), .Z(n51324) );
  XOR2_X1 U54561 ( .A1(n9416), .A2(n51324), .Z(n51325) );
  XOR2_X1 U54562 ( .A1(n51326), .A2(n51325), .Z(n51329) );
  XOR2_X1 U54563 ( .A1(n51329), .A2(n51328), .Z(n51330) );
  XOR2_X1 U54564 ( .A1(n52348), .A2(n51330), .Z(n51332) );
  NAND3_X1 U54566 ( .A1(n52701), .A2(n56547), .A3(n56544), .ZN(n56386) );
  XOR2_X1 U54569 ( .A1(n53272), .A2(n57131), .Z(n51337) );
  XOR2_X1 U54570 ( .A1(n51392), .A2(n51337), .Z(n51338) );
  XOR2_X1 U54571 ( .A1(n51339), .A2(n51338), .Z(n51340) );
  INV_X1 U54572 ( .I(n23213), .ZN(n51342) );
  NAND3_X1 U54573 ( .A1(n51346), .A2(n22229), .A3(n51345), .ZN(n51350) );
  NAND4_X1 U54574 ( .A1(n51350), .A2(n52708), .A3(n51349), .A4(n51348), .ZN(
        n51353) );
  INV_X1 U54575 ( .I(n51354), .ZN(n51356) );
  XOR2_X1 U54576 ( .A1(n51356), .A2(n51355), .Z(n51357) );
  XOR2_X1 U54577 ( .A1(n50195), .A2(n51357), .Z(n51360) );
  INV_X1 U54578 ( .I(n51521), .ZN(n51577) );
  XOR2_X1 U54579 ( .A1(n51364), .A2(n51365), .Z(n51367) );
  XOR2_X1 U54580 ( .A1(n51369), .A2(n51368), .Z(n51377) );
  INV_X1 U54581 ( .I(n51370), .ZN(n51372) );
  XOR2_X1 U54582 ( .A1(n51372), .A2(n51371), .Z(n51373) );
  XOR2_X1 U54583 ( .A1(n51374), .A2(n51373), .Z(n51375) );
  XOR2_X1 U54584 ( .A1(n51375), .A2(n1289), .Z(n51376) );
  XOR2_X1 U54586 ( .A1(n51381), .A2(n55034), .Z(n51383) );
  XOR2_X1 U54587 ( .A1(n51383), .A2(n51382), .Z(n51384) );
  XOR2_X1 U54588 ( .A1(n51687), .A2(n52331), .Z(n52611) );
  XOR2_X1 U54589 ( .A1(n51390), .A2(n52457), .Z(n51402) );
  XOR2_X1 U54591 ( .A1(n52029), .A2(n51392), .Z(n51393) );
  XOR2_X1 U54592 ( .A1(n51394), .A2(n51393), .Z(n51395) );
  XOR2_X1 U54593 ( .A1(n51397), .A2(n51396), .Z(n51398) );
  XOR2_X1 U54594 ( .A1(n51398), .A2(n14870), .Z(n51399) );
  NAND2_X1 U54597 ( .A1(n56612), .A2(n61902), .ZN(n51403) );
  XOR2_X1 U54599 ( .A1(n51408), .A2(n51407), .Z(n51409) );
  XOR2_X1 U54600 ( .A1(n51979), .A2(n51409), .Z(n51410) );
  XOR2_X1 U54601 ( .A1(n51411), .A2(n51410), .Z(n51412) );
  XOR2_X1 U54602 ( .A1(n52471), .A2(n51412), .Z(n51413) );
  XOR2_X1 U54603 ( .A1(n22614), .A2(n51413), .Z(n51414) );
  XOR2_X1 U54604 ( .A1(n8273), .A2(n51414), .Z(n51416) );
  XOR2_X1 U54605 ( .A1(n51945), .A2(n23885), .Z(n51415) );
  XOR2_X1 U54606 ( .A1(n51416), .A2(n51415), .Z(n51417) );
  INV_X1 U54608 ( .I(n51419), .ZN(n51421) );
  XNOR2_X1 U54609 ( .A1(n60556), .A2(n53787), .ZN(n51420) );
  XOR2_X1 U54610 ( .A1(n51421), .A2(n51420), .Z(n51422) );
  XOR2_X1 U54611 ( .A1(n51423), .A2(n51422), .Z(n51424) );
  XOR2_X1 U54612 ( .A1(n1625), .A2(n10335), .Z(n51425) );
  XOR2_X1 U54613 ( .A1(n51426), .A2(n51425), .Z(n51429) );
  XOR2_X1 U54614 ( .A1(n60964), .A2(n23762), .Z(n51428) );
  XOR2_X1 U54615 ( .A1(n51429), .A2(n51428), .Z(n51432) );
  XOR2_X1 U54616 ( .A1(n51554), .A2(n51430), .Z(n51431) );
  XOR2_X1 U54617 ( .A1(n51432), .A2(n51431), .Z(n51433) );
  OR2_X2 U54618 ( .A1(n13920), .A2(n52270), .Z(n56980) );
  INV_X1 U54619 ( .I(n56980), .ZN(n51435) );
  AOI21_X1 U54621 ( .A1(n51438), .A2(n52682), .B(n56978), .ZN(n51441) );
  AOI21_X1 U54623 ( .A1(n52688), .A2(n61528), .B(n13920), .ZN(n51442) );
  NOR2_X1 U54624 ( .A1(n51442), .A2(n52890), .ZN(n51446) );
  NAND2_X1 U54625 ( .A1(n61902), .A2(n56978), .ZN(n51443) );
  NAND2_X1 U54627 ( .A1(n21066), .A2(n56631), .ZN(n51450) );
  NAND2_X1 U54628 ( .A1(n52717), .A2(n56623), .ZN(n51455) );
  NAND2_X1 U54630 ( .A1(n56217), .A2(n23165), .ZN(n51451) );
  INV_X1 U54633 ( .I(n56204), .ZN(n51456) );
  NOR2_X1 U54634 ( .A1(n56630), .A2(n51457), .ZN(n51458) );
  NAND2_X1 U54635 ( .A1(n56413), .A2(n51458), .ZN(n51459) );
  NAND2_X2 U54636 ( .A1(n51460), .A2(n51459), .ZN(n56803) );
  NAND3_X1 U54639 ( .A1(n57063), .A2(n21079), .A3(n60934), .ZN(n51462) );
  INV_X1 U54643 ( .I(n52854), .ZN(n51465) );
  NAND2_X1 U54645 ( .A1(n57062), .A2(n57070), .ZN(n51466) );
  NAND3_X1 U54646 ( .A1(n51466), .A2(n63743), .A3(n507), .ZN(n51467) );
  AOI21_X1 U54647 ( .A1(n56747), .A2(n51473), .B(n56806), .ZN(n51562) );
  NAND2_X1 U54648 ( .A1(n56808), .A2(n56803), .ZN(n51560) );
  XOR2_X1 U54649 ( .A1(n23670), .A2(n63021), .Z(n51476) );
  XOR2_X1 U54650 ( .A1(n51476), .A2(n51475), .Z(n51477) );
  INV_X1 U54651 ( .I(n51479), .ZN(n51480) );
  XOR2_X1 U54652 ( .A1(n51481), .A2(n51480), .Z(n51483) );
  INV_X1 U54653 ( .I(n51485), .ZN(n51486) );
  XOR2_X1 U54654 ( .A1(n51487), .A2(n51486), .Z(n51488) );
  XOR2_X1 U54655 ( .A1(n23213), .A2(n51488), .Z(n51489) );
  XNOR2_X1 U54656 ( .A1(n51493), .A2(n51492), .ZN(n51495) );
  XOR2_X1 U54657 ( .A1(n51495), .A2(n51494), .Z(n51496) );
  XOR2_X1 U54658 ( .A1(n51497), .A2(n51496), .Z(n51498) );
  XOR2_X1 U54659 ( .A1(n51499), .A2(n51498), .Z(n51500) );
  XOR2_X1 U54660 ( .A1(n15096), .A2(n51500), .Z(n51501) );
  XOR2_X1 U54661 ( .A1(n9854), .A2(n24758), .Z(n51511) );
  XOR2_X1 U54662 ( .A1(n30908), .A2(n51512), .Z(n51513) );
  XOR2_X1 U54663 ( .A1(n51514), .A2(n51513), .Z(n51515) );
  XOR2_X1 U54664 ( .A1(n51516), .A2(n51515), .Z(n51517) );
  XOR2_X1 U54665 ( .A1(n51518), .A2(n59891), .Z(n51519) );
  INV_X1 U54666 ( .I(n51523), .ZN(n51525) );
  XOR2_X1 U54667 ( .A1(n51525), .A2(n51524), .Z(n51526) );
  XOR2_X1 U54668 ( .A1(n51530), .A2(n51531), .Z(n51533) );
  XOR2_X1 U54669 ( .A1(n51533), .A2(n51532), .Z(n51534) );
  XOR2_X1 U54670 ( .A1(n51535), .A2(n51534), .Z(n51536) );
  XOR2_X1 U54671 ( .A1(n52073), .A2(n51536), .Z(n51537) );
  XOR2_X1 U54672 ( .A1(n51543), .A2(n51542), .Z(n51544) );
  XOR2_X1 U54673 ( .A1(n51545), .A2(n51544), .Z(n51546) );
  XOR2_X1 U54674 ( .A1(n10335), .A2(n51546), .Z(n51547) );
  XOR2_X1 U54675 ( .A1(n51548), .A2(n51547), .Z(n51549) );
  XOR2_X1 U54676 ( .A1(n51554), .A2(n51553), .Z(n51555) );
  XOR2_X1 U54677 ( .A1(n52195), .A2(n51555), .Z(n51556) );
  INV_X1 U54679 ( .I(n56659), .ZN(n56369) );
  NAND2_X1 U54681 ( .A1(n51560), .A2(n23879), .ZN(n51561) );
  XOR2_X1 U54683 ( .A1(n51573), .A2(n54208), .Z(n51574) );
  XOR2_X1 U54684 ( .A1(n51575), .A2(n51574), .Z(n51576) );
  XOR2_X1 U54685 ( .A1(n51579), .A2(n51578), .Z(n51580) );
  XOR2_X1 U54686 ( .A1(n59891), .A2(n1289), .Z(n51582) );
  XOR2_X1 U54687 ( .A1(n51585), .A2(n55840), .Z(n51586) );
  XOR2_X1 U54688 ( .A1(n51587), .A2(n51586), .Z(n51588) );
  XOR2_X1 U54689 ( .A1(n51797), .A2(n52734), .Z(n51595) );
  XOR2_X1 U54690 ( .A1(n63021), .A2(n51596), .Z(n51598) );
  INV_X1 U54691 ( .I(n22783), .ZN(n51597) );
  XOR2_X1 U54692 ( .A1(n51598), .A2(n51597), .Z(n51599) );
  XOR2_X1 U54693 ( .A1(n20332), .A2(n25061), .Z(n51602) );
  XOR2_X1 U54694 ( .A1(n51609), .A2(n51608), .Z(n51614) );
  XOR2_X1 U54695 ( .A1(n51611), .A2(n51610), .Z(n51612) );
  XOR2_X1 U54696 ( .A1(n51612), .A2(n51665), .Z(n51613) );
  XOR2_X1 U54697 ( .A1(n51620), .A2(n51619), .Z(n51633) );
  XOR2_X1 U54698 ( .A1(n9722), .A2(n56335), .Z(n51622) );
  XOR2_X1 U54699 ( .A1(n51623), .A2(n51622), .Z(n51624) );
  XOR2_X1 U54700 ( .A1(n51625), .A2(n51624), .Z(n51626) );
  XOR2_X1 U54701 ( .A1(n51653), .A2(n51630), .Z(n51631) );
  NAND2_X1 U54703 ( .A1(n5227), .A2(n54814), .ZN(n51635) );
  XOR2_X1 U54705 ( .A1(n51638), .A2(n53138), .Z(n51639) );
  XOR2_X1 U54706 ( .A1(n51640), .A2(n51639), .Z(n51641) );
  XOR2_X1 U54707 ( .A1(n51642), .A2(n51641), .Z(n51643) );
  XOR2_X1 U54708 ( .A1(n51646), .A2(n20304), .Z(n51647) );
  XOR2_X1 U54709 ( .A1(n51649), .A2(n51648), .Z(n51650) );
  XOR2_X1 U54710 ( .A1(n4265), .A2(n51650), .Z(n51651) );
  XOR2_X1 U54711 ( .A1(n51654), .A2(n9871), .Z(n51655) );
  XOR2_X1 U54712 ( .A1(n51656), .A2(n51655), .Z(n51657) );
  XOR2_X1 U54713 ( .A1(n51658), .A2(n51657), .Z(n51659) );
  XOR2_X1 U54714 ( .A1(n52472), .A2(n51659), .Z(n51660) );
  XOR2_X1 U54715 ( .A1(n52073), .A2(n56949), .Z(n51661) );
  INV_X1 U54716 ( .I(n51703), .ZN(n54470) );
  XOR2_X1 U54717 ( .A1(n52420), .A2(n23642), .Z(n51663) );
  XOR2_X1 U54718 ( .A1(n19125), .A2(n51663), .Z(n51664) );
  XOR2_X1 U54719 ( .A1(n51665), .A2(n55052), .Z(n51666) );
  XOR2_X1 U54720 ( .A1(n51667), .A2(n51666), .Z(n51668) );
  XOR2_X1 U54721 ( .A1(n51669), .A2(n51668), .Z(n51670) );
  XOR2_X1 U54722 ( .A1(n7229), .A2(n51670), .Z(n51672) );
  XOR2_X1 U54723 ( .A1(n51960), .A2(n51673), .Z(n51675) );
  XOR2_X1 U54724 ( .A1(n15719), .A2(n22666), .Z(n51674) );
  XNOR2_X1 U54725 ( .A1(n56180), .A2(n52734), .ZN(n51678) );
  XOR2_X1 U54726 ( .A1(n51679), .A2(n51678), .Z(n51681) );
  XOR2_X1 U54727 ( .A1(n51681), .A2(n51680), .Z(n51682) );
  XOR2_X1 U54728 ( .A1(n52325), .A2(n51682), .Z(n51683) );
  XOR2_X1 U54729 ( .A1(n51684), .A2(n51683), .Z(n51685) );
  XOR2_X1 U54730 ( .A1(n51687), .A2(n51686), .Z(n51688) );
  XOR2_X1 U54731 ( .A1(n4470), .A2(n23758), .Z(n51692) );
  XOR2_X1 U54732 ( .A1(n51694), .A2(n51881), .Z(n51695) );
  XOR2_X1 U54733 ( .A1(n51696), .A2(n51695), .Z(n51697) );
  MUX2_X1 U54735 ( .I0(n61133), .I1(n51704), .S(n64307), .Z(n51709) );
  NOR2_X1 U54736 ( .A1(n54597), .A2(n54088), .ZN(n51705) );
  NAND2_X1 U54737 ( .A1(n54599), .A2(n54596), .ZN(n51707) );
  OAI22_X1 U54739 ( .A1(n53016), .A2(n13815), .B1(n53876), .B2(n53548), .ZN(
        n51717) );
  XOR2_X1 U54740 ( .A1(n51719), .A2(n51718), .Z(n51720) );
  XOR2_X1 U54741 ( .A1(n51724), .A2(n51723), .Z(n51725) );
  XOR2_X1 U54742 ( .A1(n52406), .A2(n51726), .Z(n51727) );
  XOR2_X1 U54744 ( .A1(n56827), .A2(n55840), .Z(n51732) );
  XOR2_X1 U54745 ( .A1(n51733), .A2(n51732), .Z(n51734) );
  XOR2_X1 U54746 ( .A1(n51735), .A2(n51734), .Z(n51736) );
  XOR2_X1 U54747 ( .A1(n20774), .A2(n51740), .Z(n51742) );
  XOR2_X1 U54748 ( .A1(n23213), .A2(n62589), .Z(n51743) );
  XOR2_X1 U54749 ( .A1(n51744), .A2(n51743), .Z(n51745) );
  XOR2_X1 U54750 ( .A1(n51986), .A2(n23022), .Z(n51750) );
  XOR2_X1 U54751 ( .A1(n51752), .A2(n51751), .Z(n51754) );
  XOR2_X1 U54752 ( .A1(n52461), .A2(n56949), .Z(n51753) );
  XOR2_X1 U54753 ( .A1(n51754), .A2(n51753), .Z(n51755) );
  XOR2_X1 U54754 ( .A1(n52073), .A2(n51757), .Z(n51758) );
  XOR2_X1 U54755 ( .A1(n51759), .A2(n51758), .Z(n51760) );
  XOR2_X1 U54756 ( .A1(n51766), .A2(n51765), .Z(n51767) );
  XOR2_X1 U54757 ( .A1(n51768), .A2(n51767), .Z(n51769) );
  XOR2_X1 U54758 ( .A1(n22666), .A2(n51770), .Z(n51771) );
  NOR2_X1 U54761 ( .A1(n7518), .A2(n54481), .ZN(n51777) );
  NAND2_X1 U54762 ( .A1(n51775), .A2(n63569), .ZN(n51776) );
  NAND2_X1 U54763 ( .A1(n54622), .A2(n54966), .ZN(n51780) );
  XOR2_X1 U54764 ( .A1(n51782), .A2(n51781), .Z(n51783) );
  XOR2_X1 U54766 ( .A1(n51788), .A2(n63021), .Z(n51789) );
  XOR2_X1 U54768 ( .A1(n51793), .A2(n52135), .Z(n51795) );
  XOR2_X1 U54769 ( .A1(n51795), .A2(n51794), .Z(n51796) );
  XOR2_X1 U54770 ( .A1(n23213), .A2(n51796), .Z(n51798) );
  XOR2_X1 U54771 ( .A1(n51798), .A2(n24076), .Z(n51799) );
  XOR2_X1 U54773 ( .A1(n51800), .A2(n23882), .Z(n51802) );
  XOR2_X1 U54774 ( .A1(n51802), .A2(n51801), .Z(n51803) );
  XOR2_X1 U54776 ( .A1(n51815), .A2(n51814), .Z(n51816) );
  XOR2_X1 U54777 ( .A1(n22979), .A2(n51819), .Z(n51820) );
  XOR2_X1 U54779 ( .A1(n52197), .A2(n1900), .Z(n51824) );
  XOR2_X1 U54780 ( .A1(n51824), .A2(n52196), .Z(n51825) );
  XOR2_X1 U54781 ( .A1(n51826), .A2(n51825), .Z(n51827) );
  XOR2_X1 U54782 ( .A1(n51828), .A2(n51827), .Z(n51829) );
  XOR2_X1 U54783 ( .A1(n51830), .A2(n51831), .Z(n51835) );
  XOR2_X1 U54784 ( .A1(n22666), .A2(n51833), .Z(n51834) );
  INV_X2 U54786 ( .I(n51837), .ZN(n53848) );
  INV_X1 U54787 ( .I(n52983), .ZN(n51838) );
  XOR2_X1 U54788 ( .A1(n51841), .A2(n51840), .Z(n51842) );
  XOR2_X1 U54789 ( .A1(n16299), .A2(n51842), .Z(n51843) );
  XOR2_X1 U54790 ( .A1(n52472), .A2(n51843), .Z(n51844) );
  XOR2_X1 U54791 ( .A1(n51845), .A2(n51844), .Z(n51848) );
  XOR2_X1 U54792 ( .A1(n51846), .A2(n52465), .Z(n51847) );
  XOR2_X1 U54793 ( .A1(n51848), .A2(n51847), .Z(n51849) );
  XOR2_X1 U54795 ( .A1(n22660), .A2(n51851), .Z(n51852) );
  XOR2_X1 U54796 ( .A1(n51853), .A2(n51852), .Z(n51855) );
  NAND2_X1 U54800 ( .A1(n53850), .A2(n4473), .ZN(n51859) );
  INV_X1 U54804 ( .I(n54018), .ZN(n51862) );
  NAND2_X1 U54805 ( .A1(n54015), .A2(n59970), .ZN(n51861) );
  NAND3_X1 U54806 ( .A1(n51862), .A2(n54349), .A3(n51861), .ZN(n51873) );
  NAND2_X1 U54808 ( .A1(n51865), .A2(n53881), .ZN(n51869) );
  INV_X1 U54809 ( .I(n54344), .ZN(n51867) );
  NAND2_X1 U54810 ( .A1(n51867), .A2(n65155), .ZN(n51868) );
  NAND3_X1 U54811 ( .A1(n51869), .A2(n51868), .A3(n54348), .ZN(n51872) );
  NAND2_X1 U54812 ( .A1(n53885), .A2(n23482), .ZN(n51871) );
  NAND3_X1 U54813 ( .A1(n54242), .A2(n22545), .A3(n57202), .ZN(n51874) );
  NAND2_X1 U54814 ( .A1(n54272), .A2(n57202), .ZN(n54270) );
  INV_X1 U54815 ( .I(n54270), .ZN(n51876) );
  INV_X1 U54816 ( .I(n54232), .ZN(n51879) );
  NOR2_X1 U54817 ( .A1(n1256), .A2(n54277), .ZN(n54273) );
  NAND2_X1 U54818 ( .A1(n54273), .A2(n54271), .ZN(n51880) );
  INV_X1 U54819 ( .I(n55911), .ZN(n51882) );
  NAND2_X1 U54820 ( .A1(n56248), .A2(n22473), .ZN(n51889) );
  NAND2_X1 U54821 ( .A1(n52222), .A2(n56264), .ZN(n51892) );
  NAND2_X1 U54822 ( .A1(n52219), .A2(n9003), .ZN(n51893) );
  INV_X1 U54823 ( .I(n55660), .ZN(n51895) );
  INV_X1 U54824 ( .I(n1616), .ZN(n56227) );
  NOR2_X1 U54825 ( .A1(n56425), .A2(n61368), .ZN(n51897) );
  INV_X1 U54826 ( .I(n56433), .ZN(n51903) );
  NOR2_X1 U54827 ( .A1(n14884), .A2(n56436), .ZN(n55987) );
  AND2_X1 U54828 ( .A1(n55987), .A2(n56229), .Z(n51899) );
  NOR2_X1 U54830 ( .A1(n51904), .A2(n56430), .ZN(n51907) );
  XOR2_X1 U54831 ( .A1(n15649), .A2(n52232), .Z(n51908) );
  XOR2_X1 U54832 ( .A1(n52538), .A2(n51908), .Z(n51909) );
  XOR2_X1 U54833 ( .A1(n51913), .A2(n53375), .Z(n51914) );
  XOR2_X1 U54834 ( .A1(n51915), .A2(n51914), .Z(n51916) );
  XOR2_X1 U54835 ( .A1(n17336), .A2(n22747), .Z(n51919) );
  XOR2_X1 U54836 ( .A1(n51921), .A2(n51920), .Z(n51922) );
  XOR2_X1 U54838 ( .A1(n54249), .A2(n56065), .Z(n51925) );
  XOR2_X1 U54839 ( .A1(n51926), .A2(n51925), .Z(n51927) );
  XOR2_X1 U54840 ( .A1(n51928), .A2(n51927), .Z(n51929) );
  XOR2_X1 U54841 ( .A1(n52325), .A2(n55792), .Z(n52092) );
  XOR2_X1 U54844 ( .A1(n23991), .A2(n13325), .Z(n51944) );
  XOR2_X1 U54845 ( .A1(n51947), .A2(n51946), .Z(n51948) );
  XOR2_X1 U54846 ( .A1(n51949), .A2(n51948), .Z(n51950) );
  XOR2_X1 U54847 ( .A1(n23016), .A2(n51950), .Z(n51951) );
  XOR2_X1 U54848 ( .A1(n51954), .A2(n51953), .Z(n51955) );
  XOR2_X1 U54849 ( .A1(n51957), .A2(n23762), .Z(n51958) );
  XOR2_X1 U54850 ( .A1(n52421), .A2(n23642), .Z(n52589) );
  XOR2_X1 U54852 ( .A1(n51968), .A2(n51967), .Z(n51969) );
  XOR2_X1 U54853 ( .A1(n52429), .A2(n51969), .Z(n51970) );
  XOR2_X1 U54854 ( .A1(n51970), .A2(n1625), .Z(n51971) );
  XOR2_X1 U54855 ( .A1(n51972), .A2(n51971), .Z(n51974) );
  XOR2_X1 U54856 ( .A1(n51974), .A2(n51973), .Z(n51976) );
  XOR2_X1 U54857 ( .A1(n51978), .A2(n9722), .Z(n51982) );
  XOR2_X1 U54858 ( .A1(n51980), .A2(n51979), .Z(n51981) );
  XOR2_X1 U54859 ( .A1(n51982), .A2(n51981), .Z(n51983) );
  XOR2_X1 U54860 ( .A1(n23991), .A2(n51984), .Z(n51985) );
  XOR2_X1 U54861 ( .A1(n724), .A2(n51985), .Z(n51988) );
  XOR2_X1 U54863 ( .A1(n51993), .A2(n51992), .Z(n51994) );
  XOR2_X1 U54864 ( .A1(n7528), .A2(n51994), .Z(n51995) );
  XNOR2_X1 U54865 ( .A1(n9231), .A2(n10594), .ZN(n51998) );
  XOR2_X1 U54866 ( .A1(n17598), .A2(n51998), .Z(n52006) );
  XOR2_X1 U54867 ( .A1(n52001), .A2(n52000), .Z(n52002) );
  XOR2_X1 U54868 ( .A1(n52003), .A2(n52002), .Z(n52004) );
  NAND2_X1 U54870 ( .A1(n52009), .A2(n52008), .ZN(n52035) );
  XOR2_X1 U54871 ( .A1(n52011), .A2(n52010), .Z(n52012) );
  XOR2_X1 U54872 ( .A1(n24025), .A2(n52012), .Z(n52014) );
  XOR2_X1 U54873 ( .A1(n52323), .A2(n52014), .Z(n52015) );
  XOR2_X1 U54874 ( .A1(n22373), .A2(n52015), .Z(n52016) );
  XOR2_X1 U54875 ( .A1(n52114), .A2(n52016), .Z(n52017) );
  XOR2_X1 U54876 ( .A1(n52018), .A2(n58084), .Z(n52019) );
  XOR2_X1 U54877 ( .A1(n52020), .A2(n52019), .Z(n52021) );
  XOR2_X1 U54878 ( .A1(n52022), .A2(n52021), .Z(n52023) );
  XOR2_X1 U54879 ( .A1(n52617), .A2(n52023), .Z(n52024) );
  OAI22_X1 U54881 ( .A1(n55966), .A2(n20891), .B1(n58626), .B2(n14142), .ZN(
        n52034) );
  AOI22_X1 U54882 ( .A1(n52035), .A2(n55975), .B1(n52034), .B2(n52033), .ZN(
        n52040) );
  INV_X1 U54883 ( .I(n24091), .ZN(n52036) );
  NAND2_X1 U54884 ( .A1(n55680), .A2(n52036), .ZN(n52037) );
  NAND3_X1 U54885 ( .A1(n52130), .A2(n55967), .A3(n52037), .ZN(n52038) );
  AOI22_X1 U54886 ( .A1(n52038), .A2(n4830), .B1(n55294), .B2(n23900), .ZN(
        n52039) );
  NOR2_X1 U54888 ( .A1(n55896), .A2(n55885), .ZN(n55837) );
  NOR3_X1 U54889 ( .A1(n55896), .A2(n19307), .A3(n55885), .ZN(n55835) );
  OAI21_X1 U54890 ( .A1(n15716), .A2(n55893), .B(n55854), .ZN(n52042) );
  MUX2_X1 U54891 ( .I0(n13858), .I1(n55898), .S(n60203), .Z(n52043) );
  NAND4_X1 U54892 ( .A1(n55295), .A2(n10362), .A3(n55690), .A4(n51961), .ZN(
        n52045) );
  XOR2_X1 U54893 ( .A1(n52051), .A2(n52050), .Z(n52052) );
  XOR2_X1 U54894 ( .A1(n8006), .A2(n52052), .Z(n52054) );
  XOR2_X1 U54895 ( .A1(n52061), .A2(n52060), .Z(n52062) );
  XOR2_X1 U54896 ( .A1(n52062), .A2(n52537), .Z(n52063) );
  XOR2_X1 U54897 ( .A1(n23173), .A2(n52063), .Z(n52064) );
  XOR2_X1 U54898 ( .A1(n52069), .A2(n52068), .Z(n52070) );
  XOR2_X1 U54899 ( .A1(n52071), .A2(n52070), .Z(n52072) );
  XOR2_X1 U54900 ( .A1(n52076), .A2(n52075), .Z(n52077) );
  XOR2_X1 U54901 ( .A1(n52080), .A2(n55765), .Z(n52081) );
  XOR2_X1 U54902 ( .A1(n52082), .A2(n52081), .Z(n52083) );
  XOR2_X1 U54903 ( .A1(n23642), .A2(n52083), .Z(n52084) );
  XOR2_X1 U54905 ( .A1(n52088), .A2(n10896), .Z(n52089) );
  XOR2_X1 U54906 ( .A1(n52096), .A2(n52095), .Z(n52098) );
  XOR2_X1 U54907 ( .A1(n52098), .A2(n52097), .Z(n52099) );
  XOR2_X1 U54908 ( .A1(n52100), .A2(n52099), .Z(n52101) );
  XOR2_X1 U54909 ( .A1(n52101), .A2(n19847), .Z(n52102) );
  XOR2_X1 U54910 ( .A1(n52609), .A2(n52102), .Z(n52104) );
  XOR2_X1 U54911 ( .A1(n53772), .A2(n55840), .Z(n52108) );
  XOR2_X1 U54912 ( .A1(n52109), .A2(n52108), .Z(n52110) );
  XOR2_X1 U54913 ( .A1(n52111), .A2(n52110), .Z(n52112) );
  XOR2_X1 U54914 ( .A1(n52321), .A2(n52112), .Z(n52113) );
  XOR2_X1 U54915 ( .A1(n535), .A2(n22747), .Z(n52115) );
  INV_X1 U54916 ( .I(n55317), .ZN(n52493) );
  NAND3_X1 U54917 ( .A1(n58626), .A2(n20891), .A3(n64970), .ZN(n52129) );
  XOR2_X1 U54919 ( .A1(n52135), .A2(n56784), .Z(n52136) );
  XOR2_X1 U54920 ( .A1(n52137), .A2(n52136), .Z(n52139) );
  XOR2_X1 U54921 ( .A1(n52139), .A2(n52138), .Z(n52140) );
  XOR2_X1 U54922 ( .A1(n52141), .A2(n52140), .Z(n52142) );
  XOR2_X1 U54923 ( .A1(n52453), .A2(n52142), .Z(n52143) );
  XOR2_X1 U54924 ( .A1(n52334), .A2(n52143), .Z(n52144) );
  XOR2_X1 U54925 ( .A1(n52150), .A2(n52149), .Z(n52151) );
  XOR2_X1 U54926 ( .A1(n52152), .A2(n52151), .Z(n52153) );
  XOR2_X1 U54927 ( .A1(n55876), .A2(n55610), .Z(n52398) );
  XOR2_X1 U54928 ( .A1(n52160), .A2(n52398), .Z(n52161) );
  XOR2_X1 U54931 ( .A1(n52164), .A2(n52165), .Z(n52166) );
  XNOR2_X1 U54932 ( .A1(n52168), .A2(n52167), .ZN(n52170) );
  XOR2_X1 U54933 ( .A1(n52170), .A2(n52169), .Z(n52171) );
  XOR2_X1 U54934 ( .A1(n52172), .A2(n52171), .Z(n52173) );
  XOR2_X1 U54935 ( .A1(n23016), .A2(n13325), .Z(n52185) );
  XOR2_X1 U54936 ( .A1(n52178), .A2(n55150), .Z(n52179) );
  XOR2_X1 U54937 ( .A1(n52180), .A2(n52179), .Z(n52181) );
  XOR2_X1 U54938 ( .A1(n52182), .A2(n52181), .Z(n52183) );
  XOR2_X1 U54939 ( .A1(n52358), .A2(n52183), .Z(n52184) );
  XOR2_X1 U54940 ( .A1(n52185), .A2(n52184), .Z(n52186) );
  XNOR2_X1 U54946 ( .A1(n52197), .A2(n52196), .ZN(n52198) );
  XOR2_X1 U54947 ( .A1(n52199), .A2(n52198), .Z(n52200) );
  XOR2_X1 U54948 ( .A1(n23642), .A2(n52206), .Z(n52208) );
  XOR2_X1 U54949 ( .A1(n7343), .A2(n52208), .Z(n52209) );
  NAND2_X1 U54951 ( .A1(n55735), .A2(n55475), .ZN(n52212) );
  NAND2_X1 U54952 ( .A1(n22817), .A2(n56268), .ZN(n52217) );
  INV_X1 U54953 ( .I(n55924), .ZN(n52220) );
  NOR2_X1 U54954 ( .A1(n55639), .A2(n55644), .ZN(n52225) );
  INV_X1 U54955 ( .I(n52302), .ZN(n52224) );
  NAND2_X1 U54957 ( .A1(n2820), .A2(n53129), .ZN(n52229) );
  NAND2_X1 U54959 ( .A1(n59020), .A2(n53212), .ZN(n52236) );
  NAND3_X1 U54961 ( .A1(n53219), .A2(n57031), .A3(n52238), .ZN(n52239) );
  NAND2_X1 U54963 ( .A1(n57063), .A2(n60934), .ZN(n52249) );
  NOR2_X1 U54964 ( .A1(n15498), .A2(n59951), .ZN(n52253) );
  INV_X1 U54967 ( .I(n52256), .ZN(n52258) );
  AOI21_X1 U54968 ( .A1(n52256), .A2(n52255), .B(n59951), .ZN(n52257) );
  OAI21_X1 U54969 ( .A1(n52258), .A2(n52670), .B(n52257), .ZN(n52259) );
  NAND2_X1 U54970 ( .A1(n10237), .A2(n22114), .ZN(n57008) );
  OR2_X1 U54972 ( .A1(n56612), .A2(n52888), .Z(n52268) );
  NAND4_X1 U54973 ( .A1(n52268), .A2(n56977), .A3(n19151), .A4(n56980), .ZN(
        n52277) );
  OAI22_X1 U54974 ( .A1(n13920), .A2(n7835), .B1(n61902), .B2(n52888), .ZN(
        n52269) );
  INV_X1 U54975 ( .I(n56612), .ZN(n52272) );
  AOI21_X1 U54976 ( .A1(n56598), .A2(n61405), .B(n52687), .ZN(n52271) );
  AOI21_X1 U54977 ( .A1(n52272), .A2(n52687), .B(n52271), .ZN(n52273) );
  AOI21_X1 U54979 ( .A1(n56374), .A2(n60809), .B(n52281), .ZN(n52280) );
  NOR2_X1 U54981 ( .A1(n52280), .A2(n56365), .ZN(n52284) );
  NAND2_X1 U54983 ( .A1(n56942), .A2(n1583), .ZN(n56924) );
  NAND2_X1 U54984 ( .A1(n52248), .A2(n56935), .ZN(n56959) );
  XOR2_X1 U54985 ( .A1(n1583), .A2(n1257), .Z(n52289) );
  NAND2_X2 U54987 ( .A1(n55627), .A2(n59610), .ZN(n55619) );
  NOR3_X1 U54990 ( .A1(n52297), .A2(n52296), .A3(n58701), .ZN(n52305) );
  NOR4_X1 U54992 ( .A1(n58701), .A2(n52302), .A3(n52301), .A4(n63520), .ZN(
        n52303) );
  XOR2_X1 U55001 ( .A1(n52328), .A2(n52327), .Z(n52330) );
  XOR2_X1 U55002 ( .A1(n22783), .A2(n52334), .Z(n52337) );
  XOR2_X1 U55003 ( .A1(n52337), .A2(n52336), .Z(n52338) );
  XOR2_X1 U55004 ( .A1(n52425), .A2(n23306), .Z(n52342) );
  XOR2_X1 U55005 ( .A1(n52596), .A2(n52342), .Z(n52343) );
  XOR2_X1 U55007 ( .A1(n52472), .A2(n52350), .Z(n52351) );
  XNOR2_X1 U55008 ( .A1(n54917), .A2(n55580), .ZN(n52353) );
  XOR2_X1 U55009 ( .A1(n52354), .A2(n52353), .Z(n52355) );
  XOR2_X1 U55010 ( .A1(n52356), .A2(n52355), .Z(n52357) );
  XOR2_X1 U55012 ( .A1(n52362), .A2(n52361), .Z(n52363) );
  XOR2_X1 U55013 ( .A1(n52586), .A2(n52363), .Z(n52364) );
  XOR2_X1 U55014 ( .A1(n52366), .A2(n52365), .Z(n52367) );
  XOR2_X1 U55015 ( .A1(n52367), .A2(n24053), .Z(n52368) );
  XOR2_X1 U55016 ( .A1(n52376), .A2(n52375), .Z(n52377) );
  XOR2_X1 U55017 ( .A1(n52378), .A2(n52377), .Z(n52379) );
  OAI21_X1 U55019 ( .A1(n52958), .A2(n22231), .B(n1604), .ZN(n52384) );
  NAND3_X1 U55020 ( .A1(n52384), .A2(n58994), .A3(n54614), .ZN(n52387) );
  INV_X1 U55022 ( .I(n52389), .ZN(n52390) );
  INV_X1 U55023 ( .I(n55279), .ZN(n52394) );
  NOR2_X1 U55026 ( .A1(n55472), .A2(n55475), .ZN(n52396) );
  INV_X1 U55027 ( .I(n55280), .ZN(n55728) );
  NAND2_X1 U55028 ( .A1(n55479), .A2(n22592), .ZN(n52397) );
  XOR2_X1 U55029 ( .A1(n52399), .A2(n52398), .Z(n52400) );
  XOR2_X1 U55030 ( .A1(n52401), .A2(n52400), .Z(n52402) );
  XOR2_X1 U55031 ( .A1(n52411), .A2(n52410), .Z(n52412) );
  XOR2_X1 U55032 ( .A1(n7343), .A2(n52420), .Z(n52422) );
  XOR2_X1 U55033 ( .A1(n52423), .A2(n52422), .Z(n52433) );
  XOR2_X1 U55034 ( .A1(n9635), .A2(n1625), .Z(n52431) );
  XOR2_X1 U55035 ( .A1(n52425), .A2(n61737), .Z(n52426) );
  XOR2_X1 U55036 ( .A1(n52427), .A2(n52426), .Z(n52428) );
  XOR2_X1 U55037 ( .A1(n52429), .A2(n52428), .Z(n52430) );
  XOR2_X1 U55038 ( .A1(n52431), .A2(n52430), .Z(n52432) );
  XOR2_X1 U55039 ( .A1(n52433), .A2(n52432), .Z(n52434) );
  XOR2_X1 U55040 ( .A1(n17738), .A2(n52434), .Z(n52435) );
  XOR2_X1 U55041 ( .A1(n52438), .A2(n52437), .Z(n52439) );
  XOR2_X1 U55042 ( .A1(n52446), .A2(n22783), .Z(n52455) );
  XOR2_X1 U55043 ( .A1(n52449), .A2(n52448), .Z(n52450) );
  XOR2_X1 U55044 ( .A1(n52451), .A2(n52450), .Z(n52452) );
  XOR2_X1 U55045 ( .A1(n23697), .A2(n52452), .Z(n52454) );
  XOR2_X1 U55046 ( .A1(n52455), .A2(n52454), .Z(n52456) );
  XOR2_X1 U55047 ( .A1(n53174), .A2(n55150), .Z(n52459) );
  XOR2_X1 U55048 ( .A1(n52459), .A2(n55580), .Z(n52460) );
  XOR2_X1 U55049 ( .A1(n52461), .A2(n52460), .Z(n52462) );
  XOR2_X1 U55050 ( .A1(n52463), .A2(n52462), .Z(n52464) );
  XOR2_X1 U55051 ( .A1(n52465), .A2(n52464), .Z(n52466) );
  XOR2_X1 U55052 ( .A1(n52468), .A2(n52467), .Z(n52469) );
  NAND4_X1 U55053 ( .A1(n1613), .A2(n5279), .A3(n55275), .A4(n5277), .ZN(
        n52478) );
  AOI21_X1 U55054 ( .A1(n52943), .A2(n52478), .B(n55265), .ZN(n52482) );
  INV_X1 U55056 ( .I(n54647), .ZN(n52486) );
  NOR2_X1 U55057 ( .A1(n61081), .A2(n58283), .ZN(n52485) );
  NOR2_X1 U55059 ( .A1(n12074), .A2(n58283), .ZN(n52483) );
  NAND2_X1 U55060 ( .A1(n52488), .A2(n55322), .ZN(n52489) );
  XOR2_X1 U55061 ( .A1(n52500), .A2(n53284), .Z(n52501) );
  XOR2_X1 U55062 ( .A1(n52502), .A2(n52501), .Z(n52503) );
  XOR2_X1 U55063 ( .A1(n724), .A2(n52504), .Z(n52506) );
  XOR2_X1 U55064 ( .A1(n52507), .A2(n52506), .Z(n52508) );
  BUF_X4 U55065 ( .I(n52509), .Z(n55416) );
  XOR2_X1 U55066 ( .A1(n52512), .A2(n52511), .Z(n52514) );
  XOR2_X1 U55067 ( .A1(n52514), .A2(n52513), .Z(n52515) );
  XOR2_X1 U55068 ( .A1(n52516), .A2(n52515), .Z(n52517) );
  XOR2_X1 U55069 ( .A1(n52518), .A2(n52517), .Z(n52519) );
  XOR2_X1 U55070 ( .A1(n11070), .A2(n52519), .Z(n52520) );
  XOR2_X1 U55071 ( .A1(n52521), .A2(n52522), .Z(n52524) );
  XOR2_X1 U55074 ( .A1(n52533), .A2(n55833), .Z(n52535) );
  XOR2_X1 U55075 ( .A1(n52535), .A2(n52534), .Z(n52536) );
  XOR2_X1 U55076 ( .A1(n6004), .A2(n52536), .Z(n52540) );
  XOR2_X1 U55077 ( .A1(n52538), .A2(n52537), .Z(n52539) );
  XOR2_X1 U55080 ( .A1(n52544), .A2(n52543), .Z(n52546) );
  INV_X1 U55082 ( .I(n52547), .ZN(n55250) );
  XOR2_X1 U55084 ( .A1(n52551), .A2(n53090), .Z(n52552) );
  XOR2_X1 U55085 ( .A1(n52553), .A2(n52552), .Z(n52554) );
  XOR2_X1 U55086 ( .A1(n52555), .A2(n52554), .Z(n52556) );
  XOR2_X1 U55087 ( .A1(n20874), .A2(n52556), .Z(n52557) );
  XOR2_X1 U55088 ( .A1(n52558), .A2(n52557), .Z(n52561) );
  INV_X1 U55089 ( .I(n52559), .ZN(n52560) );
  XOR2_X1 U55090 ( .A1(n52561), .A2(n52560), .Z(n52562) );
  XOR2_X1 U55091 ( .A1(n52566), .A2(n52565), .Z(n52567) );
  NAND2_X1 U55092 ( .A1(n54793), .A2(n55250), .ZN(n52572) );
  NAND2_X2 U55094 ( .A1(n55397), .A2(n55400), .ZN(n55404) );
  XOR2_X1 U55095 ( .A1(n52575), .A2(n53284), .Z(n52576) );
  XOR2_X1 U55096 ( .A1(n52577), .A2(n52576), .Z(n52578) );
  XOR2_X1 U55097 ( .A1(n52579), .A2(n52578), .Z(n52580) );
  XOR2_X1 U55098 ( .A1(n63010), .A2(n52582), .Z(n52583) );
  XOR2_X1 U55099 ( .A1(n52589), .A2(n52588), .Z(n52599) );
  XOR2_X1 U55100 ( .A1(n52590), .A2(n60797), .Z(n52591) );
  XOR2_X1 U55101 ( .A1(n23249), .A2(n52591), .Z(n52593) );
  XOR2_X1 U55102 ( .A1(n22439), .A2(n52593), .Z(n52595) );
  XOR2_X1 U55103 ( .A1(n1625), .A2(n52595), .Z(n52597) );
  XOR2_X1 U55104 ( .A1(n52599), .A2(n52598), .Z(n52600) );
  XOR2_X1 U55105 ( .A1(n52606), .A2(n52605), .Z(n52607) );
  XOR2_X1 U55106 ( .A1(n52614), .A2(n52613), .Z(n52615) );
  XOR2_X1 U55107 ( .A1(n52618), .A2(n62589), .Z(n52619) );
  XOR2_X1 U55108 ( .A1(n52625), .A2(n52624), .Z(n52626) );
  XOR2_X1 U55110 ( .A1(n52634), .A2(n52633), .Z(n52635) );
  XOR2_X1 U55111 ( .A1(n52636), .A2(n52635), .Z(n52638) );
  OAI21_X1 U55112 ( .A1(n17499), .A2(n4504), .B(n54862), .ZN(n52641) );
  INV_X1 U55114 ( .I(n54862), .ZN(n52643) );
  INV_X4 U55117 ( .I(n8325), .ZN(n55168) );
  AOI22_X1 U55118 ( .A1(n55111), .A2(n1593), .B1(n52647), .B2(n52646), .ZN(
        n52658) );
  NOR2_X2 U55120 ( .A1(n55156), .A2(n26094), .ZN(n55145) );
  INV_X1 U55121 ( .I(n55145), .ZN(n52650) );
  AOI21_X1 U55122 ( .A1(n52652), .A2(n55146), .B(n52651), .ZN(n52656) );
  OAI21_X1 U55123 ( .A1(n55156), .A2(n11353), .B(n8027), .ZN(n52654) );
  AOI21_X1 U55124 ( .A1(n55157), .A2(n55168), .B(n1593), .ZN(n52653) );
  NAND3_X1 U55125 ( .A1(n55153), .A2(n52654), .A3(n52653), .ZN(n52655) );
  NAND3_X1 U55132 ( .A1(n52670), .A2(n59951), .A3(n57067), .ZN(n52678) );
  INV_X1 U55134 ( .I(n52673), .ZN(n52675) );
  INV_X4 U55136 ( .I(n56897), .ZN(n56885) );
  NOR2_X1 U55138 ( .A1(n13921), .A2(n24647), .ZN(n52689) );
  NOR2_X1 U55140 ( .A1(n56885), .A2(n56890), .ZN(n52725) );
  OAI21_X1 U55141 ( .A1(n56530), .A2(n56542), .B(n57013), .ZN(n52702) );
  NOR2_X1 U55143 ( .A1(n22229), .A2(n23334), .ZN(n52707) );
  AND2_X1 U55144 ( .A1(n56639), .A2(n56211), .Z(n52715) );
  NOR2_X1 U55146 ( .A1(n56622), .A2(n56630), .ZN(n52714) );
  NAND2_X1 U55149 ( .A1(n21066), .A2(n63038), .ZN(n52720) );
  NAND2_X1 U55151 ( .A1(n56882), .A2(n56880), .ZN(n52727) );
  NAND2_X1 U55152 ( .A1(n56885), .A2(n56892), .ZN(n56865) );
  NAND2_X1 U55154 ( .A1(n56865), .A2(n52729), .ZN(n52732) );
  INV_X1 U55157 ( .I(n52737), .ZN(n52738) );
  NOR2_X1 U55160 ( .A1(n53533), .A2(n13370), .ZN(n52744) );
  OAI21_X1 U55161 ( .A1(n52746), .A2(n52745), .B(n62090), .ZN(n52747) );
  NAND2_X1 U55162 ( .A1(n52753), .A2(n23169), .ZN(n52754) );
  OAI21_X1 U55163 ( .A1(n52755), .A2(n23169), .B(n52754), .ZN(n52761) );
  AOI21_X1 U55167 ( .A1(n52759), .A2(n52836), .B(n52758), .ZN(n52760) );
  NAND2_X1 U55168 ( .A1(n53000), .A2(n15747), .ZN(n52766) );
  NAND2_X2 U55172 ( .A1(n53580), .A2(n53009), .ZN(n53588) );
  NAND3_X1 U55177 ( .A1(n53590), .A2(n53580), .A3(n58300), .ZN(n52774) );
  NAND2_X1 U55181 ( .A1(n22105), .A2(n53860), .ZN(n52778) );
  OAI22_X1 U55182 ( .A1(n52778), .A2(n53621), .B1(n53417), .B2(n53859), .ZN(
        n52779) );
  OAI21_X1 U55186 ( .A1(n57047), .A2(n23248), .B(n833), .ZN(n52788) );
  NOR2_X1 U55187 ( .A1(n58218), .A2(n58225), .ZN(n52787) );
  INV_X1 U55188 ( .I(n53209), .ZN(n52789) );
  OAI22_X1 U55189 ( .A1(n52789), .A2(n57050), .B1(n57046), .B2(n57037), .ZN(
        n52790) );
  NAND4_X1 U55191 ( .A1(n57040), .A2(n52816), .A3(n57039), .A4(n23248), .ZN(
        n52792) );
  INV_X4 U55192 ( .I(n52762), .ZN(n53324) );
  AOI21_X1 U55193 ( .A1(n53312), .A2(n53324), .B(n53351), .ZN(n52795) );
  NAND2_X1 U55194 ( .A1(n53315), .A2(n53348), .ZN(n52801) );
  NOR2_X1 U55195 ( .A1(n1450), .A2(n53351), .ZN(n52800) );
  AOI21_X1 U55196 ( .A1(n53369), .A2(n53347), .B(n53346), .ZN(n52799) );
  AOI21_X1 U55197 ( .A1(n52801), .A2(n52800), .B(n52799), .ZN(n52812) );
  AOI21_X1 U55198 ( .A1(n53355), .A2(n17012), .B(n53369), .ZN(n52802) );
  NOR2_X1 U55199 ( .A1(n52804), .A2(n52803), .ZN(n52807) );
  INV_X1 U55200 ( .I(n52805), .ZN(n52806) );
  INV_X1 U55202 ( .I(n57050), .ZN(n52822) );
  NAND3_X1 U55203 ( .A1(n52822), .A2(n57042), .A3(n53444), .ZN(n52824) );
  NOR2_X1 U55205 ( .A1(n57029), .A2(n15434), .ZN(n52832) );
  NOR2_X1 U55206 ( .A1(n57030), .A2(n15434), .ZN(n52831) );
  OAI22_X1 U55207 ( .A1(n52832), .A2(n4658), .B1(n63339), .B2(n52831), .ZN(
        n52833) );
  OAI21_X1 U55209 ( .A1(n52837), .A2(n53198), .B(n52836), .ZN(n52838) );
  NOR2_X1 U55210 ( .A1(n52839), .A2(n52838), .ZN(n52841) );
  NAND3_X1 U55214 ( .A1(n52852), .A2(n52851), .A3(n52850), .ZN(n52856) );
  OAI21_X1 U55215 ( .A1(n57073), .A2(n57070), .B(n58815), .ZN(n52853) );
  OAI21_X1 U55216 ( .A1(n52854), .A2(n52853), .B(n21079), .ZN(n52855) );
  NOR2_X1 U55217 ( .A1(n59951), .A2(n57070), .ZN(n52859) );
  AOI21_X1 U55218 ( .A1(n58326), .A2(n60498), .B(n507), .ZN(n52864) );
  NAND2_X1 U55219 ( .A1(n52864), .A2(n52863), .ZN(n52865) );
  NOR3_X1 U55220 ( .A1(n64424), .A2(n61730), .A3(n62515), .ZN(n52869) );
  INV_X1 U55221 ( .I(n52870), .ZN(n52871) );
  NOR3_X1 U55222 ( .A1(n57008), .A2(n57390), .A3(n52871), .ZN(n52872) );
  NAND2_X1 U55223 ( .A1(n52878), .A2(n53077), .ZN(n52896) );
  NOR2_X1 U55224 ( .A1(n13757), .A2(n56978), .ZN(n52882) );
  AOI22_X1 U55225 ( .A1(n56991), .A2(n52882), .B1(n56612), .B2(n7835), .ZN(
        n52886) );
  INV_X1 U55226 ( .I(n56610), .ZN(n52885) );
  NOR3_X1 U55228 ( .A1(n4033), .A2(n22980), .A3(n23243), .ZN(n52897) );
  INV_X1 U55229 ( .I(n53119), .ZN(n53086) );
  OAI22_X1 U55230 ( .A1(n53116), .A2(n52897), .B1(n53086), .B2(n53108), .ZN(
        n52899) );
  OAI21_X1 U55231 ( .A1(n53114), .A2(n53108), .B(n53070), .ZN(n52898) );
  NOR2_X1 U55232 ( .A1(n55416), .A2(n22807), .ZN(n55245) );
  INV_X1 U55233 ( .I(n55246), .ZN(n52901) );
  INV_X1 U55235 ( .I(n55419), .ZN(n52905) );
  NAND2_X1 U55236 ( .A1(n55404), .A2(n55401), .ZN(n52903) );
  NAND2_X1 U55240 ( .A1(n55255), .A2(n55416), .ZN(n54796) );
  NOR3_X1 U55241 ( .A1(n54796), .A2(n65011), .A3(n54990), .ZN(n52906) );
  NAND2_X1 U55242 ( .A1(n52908), .A2(n55416), .ZN(n52913) );
  NOR2_X1 U55245 ( .A1(n55244), .A2(n55398), .ZN(n52911) );
  NOR2_X1 U55246 ( .A1(n55300), .A2(n55690), .ZN(n55304) );
  NAND2_X1 U55247 ( .A1(n52920), .A2(n52919), .ZN(n52921) );
  NAND2_X1 U55249 ( .A1(n55287), .A2(n55474), .ZN(n52922) );
  OAI21_X1 U55250 ( .A1(n61282), .A2(n52922), .B(n55740), .ZN(n52924) );
  INV_X1 U55251 ( .I(n55465), .ZN(n52930) );
  INV_X1 U55252 ( .I(n52927), .ZN(n52929) );
  AOI21_X1 U55254 ( .A1(n52930), .A2(n52929), .B(n52928), .ZN(n52940) );
  NOR2_X1 U55255 ( .A1(n52933), .A2(n55472), .ZN(n52938) );
  NAND2_X1 U55257 ( .A1(n12074), .A2(n21268), .ZN(n52945) );
  NOR2_X1 U55260 ( .A1(n58283), .A2(n54997), .ZN(n52948) );
  NOR2_X1 U55261 ( .A1(n55316), .A2(n55306), .ZN(n52951) );
  NAND2_X1 U55262 ( .A1(n55442), .A2(n55433), .ZN(n52953) );
  NAND2_X1 U55263 ( .A1(n54618), .A2(n1604), .ZN(n52959) );
  NAND3_X1 U55264 ( .A1(n52959), .A2(n54955), .A3(n64879), .ZN(n52962) );
  NAND3_X1 U55265 ( .A1(n64879), .A2(n54616), .A3(n59879), .ZN(n52961) );
  NAND2_X1 U55267 ( .A1(n16978), .A2(n17155), .ZN(n52965) );
  AOI21_X1 U55268 ( .A1(n52966), .A2(n55222), .B(n20839), .ZN(n55202) );
  NAND2_X1 U55269 ( .A1(n55237), .A2(n16383), .ZN(n52967) );
  NAND2_X1 U55270 ( .A1(n55202), .A2(n52967), .ZN(n52968) );
  NOR2_X1 U55272 ( .A1(n21919), .A2(n52972), .ZN(n53552) );
  NAND2_X1 U55273 ( .A1(n52974), .A2(n14446), .ZN(n52976) );
  NAND3_X1 U55274 ( .A1(n53907), .A2(n21919), .A3(n54033), .ZN(n52979) );
  NAND3_X1 U55275 ( .A1(n550), .A2(n54033), .A3(n53407), .ZN(n52978) );
  NAND2_X1 U55276 ( .A1(n52979), .A2(n52978), .ZN(n52980) );
  NAND2_X1 U55278 ( .A1(n52983), .A2(n17057), .ZN(n52984) );
  NAND3_X1 U55279 ( .A1(n52984), .A2(n61371), .A3(n54067), .ZN(n52985) );
  MUX2_X1 U55280 ( .I0(n7532), .I1(n52985), .S(n52987), .Z(n52992) );
  AOI21_X1 U55281 ( .A1(n64832), .A2(n54073), .B(n52986), .ZN(n52990) );
  OAI21_X1 U55284 ( .A1(n52993), .A2(n54063), .B(n54496), .ZN(n52994) );
  INV_X1 U55285 ( .I(n52996), .ZN(n52997) );
  NAND2_X1 U55286 ( .A1(n23025), .A2(n52997), .ZN(n53581) );
  INV_X1 U55287 ( .I(n53581), .ZN(n52999) );
  INV_X1 U55288 ( .I(n53588), .ZN(n53004) );
  NAND2_X1 U55291 ( .A1(n53005), .A2(n21082), .ZN(n53008) );
  NAND2_X1 U55292 ( .A1(n53455), .A2(n5008), .ZN(n53007) );
  OAI22_X1 U55294 ( .A1(n22105), .A2(n53427), .B1(n4481), .B2(n62664), .ZN(
        n53021) );
  AOI21_X1 U55295 ( .A1(n53860), .A2(n53427), .B(n1259), .ZN(n53020) );
  OAI21_X1 U55296 ( .A1(n4480), .A2(n53421), .B(n53018), .ZN(n53019) );
  NAND2_X1 U55298 ( .A1(n53022), .A2(n7303), .ZN(n53027) );
  AOI22_X1 U55299 ( .A1(n53025), .A2(n53024), .B1(n53616), .B2(n61147), .ZN(
        n53026) );
  OAI21_X1 U55303 ( .A1(n54022), .A2(n54343), .B(n54028), .ZN(n53040) );
  NAND2_X1 U55305 ( .A1(n53820), .A2(n53809), .ZN(n53798) );
  NAND2_X1 U55306 ( .A1(n53814), .A2(n53808), .ZN(n53043) );
  AOI21_X1 U55308 ( .A1(n53113), .A2(n23243), .B(n53049), .ZN(n53063) );
  OAI21_X1 U55309 ( .A1(n62412), .A2(n53108), .B(n22980), .ZN(n53052) );
  OAI21_X1 U55310 ( .A1(n53100), .A2(n23212), .B(n53082), .ZN(n53051) );
  NOR3_X1 U55311 ( .A1(n23595), .A2(n63767), .A3(n53108), .ZN(n53050) );
  NOR2_X1 U55314 ( .A1(n53097), .A2(n53094), .ZN(n53055) );
  INV_X1 U55316 ( .I(n53082), .ZN(n53057) );
  NOR3_X1 U55317 ( .A1(n53057), .A2(n23243), .A3(n23212), .ZN(n53059) );
  OAI21_X1 U55318 ( .A1(n53059), .A2(n23595), .B(n53058), .ZN(n53060) );
  AOI21_X1 U55321 ( .A1(n53097), .A2(n53096), .B(n53117), .ZN(n53074) );
  AOI21_X1 U55322 ( .A1(n4033), .A2(n53110), .B(n53111), .ZN(n53073) );
  NOR2_X1 U55324 ( .A1(n53070), .A2(n53109), .ZN(n53071) );
  OAI21_X1 U55325 ( .A1(n53110), .A2(n53092), .B(n53071), .ZN(n53072) );
  OAI21_X1 U55326 ( .A1(n53083), .A2(n22980), .B(n53094), .ZN(n53079) );
  NOR3_X1 U55328 ( .A1(n53117), .A2(n53091), .A3(n53093), .ZN(n53088) );
  NOR2_X1 U55329 ( .A1(n53110), .A2(n53108), .ZN(n53085) );
  NAND2_X1 U55330 ( .A1(n4033), .A2(n53107), .ZN(n53084) );
  NOR2_X1 U55331 ( .A1(n53094), .A2(n53109), .ZN(n53095) );
  NAND2_X1 U55332 ( .A1(n53097), .A2(n53108), .ZN(n53098) );
  NAND3_X1 U55333 ( .A1(n53100), .A2(n53109), .A3(n23212), .ZN(n53101) );
  NOR2_X1 U55334 ( .A1(n53109), .A2(n53108), .ZN(n53112) );
  AOI21_X1 U55335 ( .A1(n53119), .A2(n23212), .B(n53117), .ZN(n53120) );
  NOR3_X1 U55337 ( .A1(n26135), .A2(n53167), .A3(n53160), .ZN(n53132) );
  NAND3_X1 U55338 ( .A1(n15415), .A2(n5614), .A3(n20735), .ZN(n53127) );
  NAND2_X1 U55339 ( .A1(n53166), .A2(n25484), .ZN(n53133) );
  NAND3_X1 U55340 ( .A1(n53133), .A2(n53135), .A3(n53160), .ZN(n53137) );
  XOR2_X1 U55342 ( .A1(n53139), .A2(n53138), .Z(Plaintext[8]) );
  NAND2_X1 U55343 ( .A1(n53145), .A2(n23856), .ZN(n53149) );
  XOR2_X1 U55344 ( .A1(n53156), .A2(n53155), .Z(Plaintext[9]) );
  NOR2_X1 U55345 ( .A1(n53162), .A2(n2037), .ZN(n53164) );
  NAND4_X1 U55346 ( .A1(n53164), .A2(n12111), .A3(n15415), .A4(n23856), .ZN(
        n53170) );
  NAND2_X1 U55347 ( .A1(n53166), .A2(n53165), .ZN(n53169) );
  NAND3_X1 U55348 ( .A1(n53170), .A2(n53169), .A3(n53168), .ZN(n53171) );
  INV_X1 U55349 ( .I(n53185), .ZN(n53176) );
  NAND2_X1 U55351 ( .A1(n53533), .A2(n23047), .ZN(n53186) );
  NOR2_X1 U55352 ( .A1(n53198), .A2(n23974), .ZN(n53190) );
  INV_X1 U55354 ( .I(n53195), .ZN(n53202) );
  NOR2_X1 U55355 ( .A1(n53198), .A2(n23169), .ZN(n53199) );
  NAND2_X1 U55356 ( .A1(n53206), .A2(n57050), .ZN(n53208) );
  NAND2_X1 U55358 ( .A1(n4658), .A2(n12777), .ZN(n53215) );
  NAND3_X1 U55359 ( .A1(n53275), .A2(n61361), .A3(n19735), .ZN(n53244) );
  NAND4_X1 U55360 ( .A1(n53258), .A2(n53265), .A3(n19735), .A4(n22889), .ZN(
        n53249) );
  NOR2_X1 U55361 ( .A1(n9338), .A2(n19735), .ZN(n53253) );
  NOR2_X1 U55362 ( .A1(n6789), .A2(n53269), .ZN(n53254) );
  AOI21_X1 U55363 ( .A1(n53257), .A2(n53267), .B(n23411), .ZN(n53260) );
  OAI21_X1 U55364 ( .A1(n53258), .A2(n53279), .B(n53288), .ZN(n53259) );
  INV_X1 U55366 ( .I(n53272), .ZN(n53273) );
  NOR3_X1 U55367 ( .A1(n59907), .A2(n53284), .A3(n53288), .ZN(n53278) );
  NOR3_X1 U55368 ( .A1(n53275), .A2(n53302), .A3(n53285), .ZN(n53277) );
  NAND2_X1 U55369 ( .A1(n22889), .A2(n1574), .ZN(n53281) );
  NOR4_X1 U55370 ( .A1(n15771), .A2(n53278), .A3(n53277), .A4(n53276), .ZN(
        n53292) );
  INV_X1 U55371 ( .I(n53281), .ZN(n53282) );
  NAND2_X1 U55372 ( .A1(n53283), .A2(n53282), .ZN(n53291) );
  NOR2_X1 U55373 ( .A1(n53286), .A2(n53285), .ZN(n53287) );
  OAI21_X1 U55374 ( .A1(n53288), .A2(n59907), .B(n53287), .ZN(n53289) );
  OAI22_X1 U55376 ( .A1(n6789), .A2(n53303), .B1(n53302), .B2(n13239), .ZN(
        n53304) );
  NOR2_X1 U55377 ( .A1(n53322), .A2(n53345), .ZN(n53309) );
  NOR2_X1 U55378 ( .A1(n11963), .A2(n53346), .ZN(n53311) );
  OAI21_X1 U55379 ( .A1(n17012), .A2(n25604), .B(n52762), .ZN(n53310) );
  NAND3_X1 U55380 ( .A1(n53312), .A2(n53369), .A3(n53324), .ZN(n53313) );
  NAND2_X1 U55381 ( .A1(n53334), .A2(n53324), .ZN(n53316) );
  AOI22_X1 U55383 ( .A1(n60517), .A2(n53316), .B1(n53315), .B2(n53314), .ZN(
        n53317) );
  NAND3_X1 U55384 ( .A1(n53323), .A2(n53324), .A3(n53345), .ZN(n53327) );
  NAND2_X1 U55385 ( .A1(n53334), .A2(n53351), .ZN(n53338) );
  AOI21_X1 U55386 ( .A1(n60115), .A2(n7093), .B(n52762), .ZN(n53337) );
  NAND2_X1 U55387 ( .A1(n11963), .A2(n53335), .ZN(n53336) );
  AOI21_X1 U55388 ( .A1(n53338), .A2(n53337), .B(n53336), .ZN(n53341) );
  AOI21_X1 U55390 ( .A1(n53339), .A2(n1450), .B(n53348), .ZN(n53340) );
  XOR2_X1 U55391 ( .A1(n9731), .A2(n25604), .Z(n53350) );
  NAND2_X1 U55392 ( .A1(n53348), .A2(n7093), .ZN(n53349) );
  NAND4_X1 U55393 ( .A1(n53350), .A2(n53349), .A3(n60517), .A4(n1450), .ZN(
        n53357) );
  NAND2_X1 U55394 ( .A1(n53355), .A2(n53368), .ZN(n53352) );
  AOI22_X1 U55395 ( .A1(n53352), .A2(n53351), .B1(n1450), .B2(n7093), .ZN(
        n53353) );
  OAI21_X1 U55396 ( .A1(n53355), .A2(n53354), .B(n53353), .ZN(n53356) );
  NAND2_X1 U55400 ( .A1(n23401), .A2(n53383), .ZN(n53378) );
  OAI21_X1 U55402 ( .A1(n53384), .A2(n23169), .B(n53382), .ZN(n53388) );
  NAND2_X1 U55403 ( .A1(n53598), .A2(n23157), .ZN(n53385) );
  NAND2_X1 U55404 ( .A1(n53386), .A2(n53385), .ZN(n53387) );
  NAND2_X2 U55405 ( .A1(n53390), .A2(n53389), .ZN(n53483) );
  AOI21_X1 U55407 ( .A1(n53541), .A2(n53540), .B(n53391), .ZN(n53395) );
  XOR2_X1 U55408 ( .A1(n22708), .A2(n23047), .Z(n53393) );
  NOR2_X1 U55409 ( .A1(n54036), .A2(n54039), .ZN(n53399) );
  MUX2_X1 U55410 ( .I0(n53403), .I1(n53399), .S(n4399), .Z(n53406) );
  INV_X1 U55411 ( .I(n53410), .ZN(n53400) );
  NOR2_X1 U55415 ( .A1(n54041), .A2(n54039), .ZN(n53408) );
  INV_X1 U55416 ( .I(n53616), .ZN(n53425) );
  NAND2_X1 U55417 ( .A1(n53859), .A2(n4226), .ZN(n53414) );
  NAND2_X1 U55419 ( .A1(n22885), .A2(n53624), .ZN(n53422) );
  INV_X1 U55420 ( .I(n65282), .ZN(n53862) );
  INV_X1 U55422 ( .I(n53852), .ZN(n53430) );
  AOI22_X1 U55423 ( .A1(n53430), .A2(n53429), .B1(n53620), .B2(n53614), .ZN(
        n53431) );
  NAND2_X1 U55424 ( .A1(n25789), .A2(n53516), .ZN(n53524) );
  NAND2_X1 U55425 ( .A1(n53492), .A2(n23611), .ZN(n53478) );
  INV_X1 U55426 ( .I(n53478), .ZN(n53460) );
  XOR2_X1 U55428 ( .A1(n26089), .A2(n15747), .Z(n53452) );
  NOR2_X1 U55431 ( .A1(n53576), .A2(n10748), .ZN(n53456) );
  INV_X4 U55432 ( .I(n53492), .ZN(n53506) );
  INV_X1 U55434 ( .I(n23926), .ZN(n53464) );
  NOR2_X1 U55435 ( .A1(n53480), .A2(n53506), .ZN(n53465) );
  AOI21_X1 U55436 ( .A1(n53492), .A2(n53519), .B(n53467), .ZN(n53469) );
  AOI21_X1 U55437 ( .A1(n53493), .A2(n53514), .B(n53480), .ZN(n53473) );
  OAI21_X1 U55438 ( .A1(n53473), .A2(n53528), .B(n53491), .ZN(n53474) );
  INV_X1 U55439 ( .I(n53489), .ZN(n53479) );
  NAND4_X1 U55440 ( .A1(n1581), .A2(n53479), .A3(n53519), .A4(n53478), .ZN(
        n53481) );
  NAND2_X1 U55441 ( .A1(n53481), .A2(n53515), .ZN(n53486) );
  INV_X1 U55442 ( .I(n53501), .ZN(n53482) );
  OAI21_X1 U55443 ( .A1(n53528), .A2(n53507), .B(n53482), .ZN(n53485) );
  NAND3_X1 U55444 ( .A1(n53524), .A2(n53505), .A3(n23611), .ZN(n53484) );
  INV_X1 U55447 ( .I(n53491), .ZN(n53500) );
  NAND2_X1 U55448 ( .A1(n53527), .A2(n53514), .ZN(n53496) );
  NAND3_X1 U55449 ( .A1(n53494), .A2(n53516), .A3(n53493), .ZN(n53495) );
  AOI21_X1 U55450 ( .A1(n53496), .A2(n53495), .B(n25789), .ZN(n53498) );
  NOR2_X1 U55451 ( .A1(n53505), .A2(n53501), .ZN(n53502) );
  NOR3_X1 U55452 ( .A1(n53504), .A2(n53503), .A3(n53502), .ZN(n53512) );
  OAI21_X1 U55453 ( .A1(n53508), .A2(n53507), .B(n53506), .ZN(n53510) );
  NAND2_X1 U55454 ( .A1(n53528), .A2(n1161), .ZN(n53509) );
  NAND2_X1 U55455 ( .A1(n53517), .A2(n53516), .ZN(n53520) );
  NAND3_X1 U55456 ( .A1(n53520), .A2(n53519), .A3(n25789), .ZN(n53522) );
  NAND2_X1 U55457 ( .A1(n53533), .A2(n23784), .ZN(n53536) );
  NAND2_X1 U55458 ( .A1(n53540), .A2(n53539), .ZN(n53542) );
  AOI21_X1 U55459 ( .A1(n53543), .A2(n53542), .B(n17264), .ZN(n53544) );
  OAI21_X1 U55461 ( .A1(n53552), .A2(n53551), .B(n53907), .ZN(n53556) );
  NAND3_X1 U55462 ( .A1(n57700), .A2(n54057), .A3(n54054), .ZN(n53554) );
  NAND3_X1 U55463 ( .A1(n53556), .A2(n53555), .A3(n53554), .ZN(n53570) );
  NOR2_X1 U55464 ( .A1(n53916), .A2(n58656), .ZN(n53558) );
  NAND2_X1 U55466 ( .A1(n54046), .A2(n54052), .ZN(n53562) );
  NAND2_X1 U55467 ( .A1(n53562), .A2(n53561), .ZN(n53564) );
  NAND2_X1 U55468 ( .A1(n53562), .A2(n54057), .ZN(n53563) );
  NAND3_X1 U55469 ( .A1(n53564), .A2(n53563), .A3(n54033), .ZN(n53568) );
  NAND3_X1 U55470 ( .A1(n53566), .A2(n54057), .A3(n53565), .ZN(n53567) );
  NAND2_X1 U55472 ( .A1(n53582), .A2(n53581), .ZN(n53583) );
  NOR3_X1 U55473 ( .A1(n53588), .A2(n53587), .A3(n53586), .ZN(n53593) );
  AOI21_X1 U55475 ( .A1(n57192), .A2(n25067), .B(n53598), .ZN(n53600) );
  NAND2_X1 U55476 ( .A1(n53672), .A2(n53688), .ZN(n53610) );
  NAND2_X1 U55477 ( .A1(n53610), .A2(n53700), .ZN(n53679) );
  INV_X1 U55478 ( .I(n53679), .ZN(n53630) );
  NOR2_X1 U55479 ( .A1(n1259), .A2(n22201), .ZN(n53611) );
  NOR3_X1 U55480 ( .A1(n53611), .A2(n4481), .A3(n53624), .ZN(n53618) );
  NOR2_X1 U55481 ( .A1(n53860), .A2(n22201), .ZN(n53613) );
  NAND2_X1 U55482 ( .A1(n53616), .A2(n18522), .ZN(n53617) );
  NOR2_X1 U55483 ( .A1(n53620), .A2(n61560), .ZN(n53623) );
  OAI22_X1 U55484 ( .A1(n53623), .A2(n53622), .B1(n4480), .B2(n53621), .ZN(
        n53626) );
  AOI22_X1 U55485 ( .A1(n53626), .A2(n53625), .B1(n61560), .B2(n53624), .ZN(
        n53627) );
  NAND2_X1 U55487 ( .A1(n53673), .A2(n53695), .ZN(n53629) );
  NOR2_X1 U55488 ( .A1(n53688), .A2(n53676), .ZN(n53628) );
  NAND2_X1 U55489 ( .A1(n53628), .A2(n53700), .ZN(n53704) );
  OAI22_X1 U55490 ( .A1(n53630), .A2(n53629), .B1(n53695), .B2(n53704), .ZN(
        n53640) );
  INV_X1 U55491 ( .I(n53667), .ZN(n53631) );
  NAND2_X1 U55492 ( .A1(n53631), .A2(n53700), .ZN(n53634) );
  NAND2_X1 U55493 ( .A1(n19475), .A2(n53699), .ZN(n53633) );
  NOR2_X1 U55494 ( .A1(n53694), .A2(n53699), .ZN(n53637) );
  NAND2_X1 U55495 ( .A1(n53678), .A2(n53691), .ZN(n53636) );
  INV_X1 U55496 ( .I(n53700), .ZN(n53689) );
  NAND3_X1 U55497 ( .A1(n53689), .A2(n53675), .A3(n53690), .ZN(n53635) );
  OAI21_X1 U55498 ( .A1(n53637), .A2(n53636), .B(n53635), .ZN(n53638) );
  NAND2_X1 U55499 ( .A1(n53699), .A2(n53676), .ZN(n53643) );
  NOR2_X1 U55500 ( .A1(n53700), .A2(n53692), .ZN(n53650) );
  MUX2_X1 U55502 ( .I0(n53652), .I1(n53651), .S(n23935), .Z(n53653) );
  NAND2_X1 U55503 ( .A1(n53657), .A2(n53656), .ZN(n53661) );
  NAND2_X1 U55504 ( .A1(n53659), .A2(n53667), .ZN(n53660) );
  AOI21_X1 U55505 ( .A1(n53661), .A2(n19475), .B(n53660), .ZN(n53663) );
  XOR2_X1 U55506 ( .A1(n53663), .A2(n53662), .Z(Plaintext[32]) );
  OAI21_X1 U55508 ( .A1(n53673), .A2(n53700), .B(n53672), .ZN(n53674) );
  AOI21_X1 U55510 ( .A1(n53682), .A2(n25859), .B(n53680), .ZN(n53683) );
  OAI21_X1 U55514 ( .A1(n53694), .A2(n53700), .B(n53693), .ZN(n53698) );
  NOR2_X1 U55515 ( .A1(n53699), .A2(n53695), .ZN(n53696) );
  NAND3_X1 U55516 ( .A1(n53756), .A2(n16489), .A3(n9616), .ZN(n53708) );
  NAND3_X1 U55517 ( .A1(n1579), .A2(n17286), .A3(n53732), .ZN(n53707) );
  NOR2_X1 U55519 ( .A1(n53756), .A2(n53718), .ZN(n53719) );
  NOR2_X1 U55521 ( .A1(n53724), .A2(n53732), .ZN(n53725) );
  NOR2_X1 U55522 ( .A1(n53738), .A2(n53725), .ZN(n53735) );
  NAND2_X1 U55523 ( .A1(n25116), .A2(n53726), .ZN(n53730) );
  NAND3_X1 U55524 ( .A1(n53730), .A2(n17286), .A3(n63920), .ZN(n53734) );
  OAI21_X1 U55525 ( .A1(n53732), .A2(n25011), .B(n53731), .ZN(n53733) );
  AOI21_X1 U55526 ( .A1(n53735), .A2(n53734), .B(n53733), .ZN(n53746) );
  INV_X1 U55527 ( .I(n53751), .ZN(n53739) );
  NAND2_X1 U55528 ( .A1(n53739), .A2(n25011), .ZN(n53743) );
  XOR2_X1 U55530 ( .A1(n53750), .A2(n53749), .Z(Plaintext[37]) );
  NOR2_X1 U55531 ( .A1(n53752), .A2(n53751), .ZN(n53753) );
  AOI21_X1 U55532 ( .A1(n25117), .A2(n25011), .B(n16489), .ZN(n53758) );
  INV_X1 U55533 ( .I(n53759), .ZN(n53761) );
  NAND2_X1 U55534 ( .A1(n53761), .A2(n61933), .ZN(n53762) );
  AOI21_X1 U55535 ( .A1(n53807), .A2(n53797), .B(n53774), .ZN(n53768) );
  NOR3_X1 U55536 ( .A1(n53797), .A2(n53826), .A3(n53809), .ZN(n53767) );
  NAND2_X1 U55537 ( .A1(n53795), .A2(n53809), .ZN(n53765) );
  NAND2_X1 U55539 ( .A1(n9161), .A2(n23206), .ZN(n53779) );
  MUX2_X1 U55542 ( .I0(n53773), .I1(n53814), .S(n21), .Z(n53786) );
  AOI21_X1 U55544 ( .A1(n53780), .A2(n53809), .B(n53811), .ZN(n53777) );
  AOI21_X1 U55546 ( .A1(n53779), .A2(n53809), .B(n4540), .ZN(n53783) );
  OAI21_X1 U55547 ( .A1(n53820), .A2(n53780), .B(n53797), .ZN(n53782) );
  INV_X1 U55549 ( .I(n53790), .ZN(n53792) );
  NAND2_X1 U55550 ( .A1(n53817), .A2(n53809), .ZN(n53791) );
  INV_X1 U55551 ( .I(n53793), .ZN(n53796) );
  NAND3_X1 U55553 ( .A1(n53796), .A2(n53815), .A3(n53821), .ZN(n53802) );
  INV_X1 U55554 ( .I(n53798), .ZN(n53799) );
  OAI21_X1 U55555 ( .A1(n53825), .A2(n53800), .B(n53799), .ZN(n53801) );
  NOR2_X1 U55556 ( .A1(n53814), .A2(n53813), .ZN(n53819) );
  NOR3_X1 U55557 ( .A1(n53817), .A2(n53826), .A3(n53042), .ZN(n53818) );
  NAND2_X1 U55558 ( .A1(n53822), .A2(n53821), .ZN(n53832) );
  NOR2_X1 U55559 ( .A1(n53824), .A2(n4540), .ZN(n53827) );
  AOI22_X1 U55560 ( .A1(n53827), .A2(n53826), .B1(n53825), .B2(n21), .ZN(
        n53831) );
  NAND2_X1 U55561 ( .A1(n53829), .A2(n53828), .ZN(n53830) );
  XOR2_X1 U55563 ( .A1(n53834), .A2(n53833), .Z(Plaintext[46]) );
  NAND2_X1 U55569 ( .A1(n54073), .A2(n53847), .ZN(n54310) );
  NAND2_X1 U55570 ( .A1(n53850), .A2(n22372), .ZN(n53851) );
  OAI21_X1 U55572 ( .A1(n4480), .A2(n62186), .B(n53858), .ZN(n53864) );
  XOR2_X1 U55573 ( .A1(n53861), .A2(n53860), .Z(n53863) );
  NAND3_X1 U55574 ( .A1(n53864), .A2(n53863), .A3(n53862), .ZN(n53865) );
  OAI21_X1 U55576 ( .A1(n53882), .A2(n54340), .B(n54349), .ZN(n53883) );
  OAI21_X1 U55577 ( .A1(n53885), .A2(n53884), .B(n53883), .ZN(n53887) );
  INV_X1 U55580 ( .I(n54321), .ZN(n54588) );
  NAND2_X1 U55581 ( .A1(n54321), .A2(n54594), .ZN(n54079) );
  NOR2_X1 U55582 ( .A1(n54088), .A2(n54594), .ZN(n53895) );
  OAI21_X1 U55583 ( .A1(n61133), .A2(n54598), .B(n53895), .ZN(n53896) );
  NAND2_X1 U55586 ( .A1(n58656), .A2(n54035), .ZN(n53906) );
  NOR2_X1 U55587 ( .A1(n53906), .A2(n23164), .ZN(n53908) );
  OAI21_X1 U55588 ( .A1(n53908), .A2(n53907), .B(n54033), .ZN(n53910) );
  NOR2_X1 U55589 ( .A1(n53908), .A2(n23217), .ZN(n53909) );
  INV_X1 U55590 ( .I(n54049), .ZN(n53921) );
  NAND3_X1 U55591 ( .A1(n53914), .A2(n54041), .A3(n53913), .ZN(n53920) );
  OR2_X1 U55592 ( .A1(n53916), .A2(n4399), .Z(n53918) );
  NAND4_X1 U55593 ( .A1(n550), .A2(n53918), .A3(n54055), .A4(n60049), .ZN(
        n53919) );
  NAND3_X1 U55594 ( .A1(n53921), .A2(n53920), .A3(n53919), .ZN(n53922) );
  NOR2_X2 U55595 ( .A1(n53923), .A2(n53922), .ZN(n54000) );
  NAND2_X1 U55597 ( .A1(n53927), .A2(n53996), .ZN(n53924) );
  NOR2_X1 U55598 ( .A1(n54001), .A2(n7492), .ZN(n53929) );
  NOR3_X1 U55601 ( .A1(n53946), .A2(n53947), .A3(n53931), .ZN(n53936) );
  NAND3_X1 U55602 ( .A1(n23292), .A2(n12915), .A3(n54012), .ZN(n53938) );
  OAI22_X1 U55603 ( .A1(n53938), .A2(n53960), .B1(n54006), .B2(n53937), .ZN(
        n53940) );
  NAND2_X1 U55604 ( .A1(n53983), .A2(n22669), .ZN(n53939) );
  NAND2_X1 U55605 ( .A1(n53940), .A2(n53939), .ZN(n53941) );
  OAI21_X1 U55606 ( .A1(n53946), .A2(n53953), .B(n53983), .ZN(n53949) );
  NOR2_X1 U55607 ( .A1(n53947), .A2(n53969), .ZN(n53948) );
  INV_X1 U55608 ( .I(n54007), .ZN(n53951) );
  OAI21_X1 U55609 ( .A1(n53952), .A2(n53951), .B(n53966), .ZN(n53956) );
  NAND2_X1 U55610 ( .A1(n58817), .A2(n53953), .ZN(n53982) );
  NAND3_X1 U55611 ( .A1(n53982), .A2(n22669), .A3(n9715), .ZN(n53955) );
  XOR2_X1 U55612 ( .A1(n53959), .A2(n53958), .Z(Plaintext[50]) );
  INV_X1 U55613 ( .I(n53960), .ZN(n53961) );
  NOR2_X1 U55614 ( .A1(n53961), .A2(n53996), .ZN(n53965) );
  INV_X1 U55615 ( .I(n53962), .ZN(n53964) );
  INV_X1 U55617 ( .I(n53983), .ZN(n53968) );
  NOR2_X1 U55618 ( .A1(n54006), .A2(n53966), .ZN(n53967) );
  AOI22_X1 U55620 ( .A1(n53968), .A2(n53967), .B1(n53979), .B2(n53999), .ZN(
        n53976) );
  NAND3_X1 U55621 ( .A1(n23292), .A2(n53969), .A3(n53992), .ZN(n53970) );
  NAND2_X1 U55622 ( .A1(n53971), .A2(n53970), .ZN(n53972) );
  NAND2_X1 U55623 ( .A1(n54001), .A2(n60426), .ZN(n53973) );
  NAND4_X1 U55624 ( .A1(n53973), .A2(n23292), .A3(n53995), .A4(n54012), .ZN(
        n53974) );
  NOR2_X1 U55626 ( .A1(n53979), .A2(n60426), .ZN(n53981) );
  NAND3_X1 U55627 ( .A1(n53983), .A2(n53995), .A3(n22669), .ZN(n53987) );
  NAND3_X1 U55628 ( .A1(n53985), .A2(n54006), .A3(n53984), .ZN(n53986) );
  NAND2_X1 U55629 ( .A1(n9715), .A2(n54006), .ZN(n53991) );
  NAND3_X1 U55630 ( .A1(n54001), .A2(n22669), .A3(n23292), .ZN(n54002) );
  INV_X1 U55634 ( .I(n54348), .ZN(n54019) );
  OAI21_X1 U55635 ( .A1(n54019), .A2(n65155), .B(n54351), .ZN(n54020) );
  INV_X1 U55636 ( .I(n54349), .ZN(n54024) );
  NAND3_X1 U55637 ( .A1(n54348), .A2(n54029), .A3(n54344), .ZN(n54030) );
  INV_X1 U55642 ( .I(n54045), .ZN(n54051) );
  INV_X1 U55644 ( .I(n54053), .ZN(n54048) );
  NAND2_X1 U55646 ( .A1(n54053), .A2(n54052), .ZN(n54059) );
  OAI21_X1 U55647 ( .A1(n54055), .A2(n14446), .B(n54054), .ZN(n54056) );
  NAND3_X1 U55651 ( .A1(n54068), .A2(n64978), .A3(n54067), .ZN(n54069) );
  INV_X1 U55652 ( .I(n54320), .ZN(n54077) );
  NAND3_X1 U55653 ( .A1(n61443), .A2(n61133), .A3(n54074), .ZN(n54075) );
  NAND3_X1 U55656 ( .A1(n61443), .A2(n54597), .A3(n54594), .ZN(n54082) );
  XOR2_X1 U55658 ( .A1(n54087), .A2(n54598), .Z(n54093) );
  NAND2_X1 U55659 ( .A1(n54466), .A2(n54088), .ZN(n54089) );
  NAND2_X1 U55660 ( .A1(n54090), .A2(n54596), .ZN(n54091) );
  NAND2_X1 U55661 ( .A1(n54091), .A2(n54470), .ZN(n54092) );
  AOI21_X1 U55662 ( .A1(n23736), .A2(n54093), .B(n54092), .ZN(n54094) );
  NAND2_X1 U55664 ( .A1(n15040), .A2(n23849), .ZN(n54100) );
  OAI21_X1 U55665 ( .A1(n54102), .A2(n24111), .B(n9137), .ZN(n54103) );
  NAND3_X1 U55666 ( .A1(n54109), .A2(n23704), .A3(n54108), .ZN(n54115) );
  NAND2_X1 U55667 ( .A1(n10425), .A2(n23704), .ZN(n54111) );
  NAND2_X1 U55668 ( .A1(n1158), .A2(n10425), .ZN(n54113) );
  NAND2_X2 U55670 ( .A1(n54199), .A2(n18859), .ZN(n54194) );
  NAND2_X1 U55672 ( .A1(n14643), .A2(n18859), .ZN(n54118) );
  NAND2_X1 U55673 ( .A1(n26008), .A2(n2984), .ZN(n54136) );
  AOI21_X1 U55674 ( .A1(n54201), .A2(n54207), .B(n54136), .ZN(n54119) );
  OAI21_X1 U55675 ( .A1(n54187), .A2(n63726), .B(n54192), .ZN(n54121) );
  OAI21_X1 U55676 ( .A1(n54189), .A2(n54198), .B(n54196), .ZN(n54120) );
  NAND2_X1 U55677 ( .A1(n54121), .A2(n54120), .ZN(n54123) );
  NOR2_X1 U55678 ( .A1(n54189), .A2(n54170), .ZN(n54161) );
  NAND2_X1 U55679 ( .A1(n54161), .A2(n10480), .ZN(n54122) );
  NAND2_X1 U55681 ( .A1(n54158), .A2(n18859), .ZN(n54128) );
  NAND2_X1 U55682 ( .A1(n54128), .A2(n63726), .ZN(n54132) );
  OAI21_X1 U55683 ( .A1(n54199), .A2(n54158), .B(n14643), .ZN(n54131) );
  INV_X1 U55684 ( .I(n54194), .ZN(n54150) );
  AOI22_X1 U55688 ( .A1(n54150), .A2(n54135), .B1(n54134), .B2(n54175), .ZN(
        n54140) );
  XOR2_X1 U55689 ( .A1(n54207), .A2(n25299), .Z(n54137) );
  NAND4_X1 U55690 ( .A1(n9968), .A2(n54137), .A3(n10480), .A4(n54136), .ZN(
        n54139) );
  NAND2_X1 U55691 ( .A1(n54175), .A2(n54192), .ZN(n54138) );
  NAND2_X1 U55693 ( .A1(n54172), .A2(n54201), .ZN(n54147) );
  NAND2_X1 U55694 ( .A1(n2984), .A2(n54207), .ZN(n54171) );
  INV_X1 U55695 ( .I(n54171), .ZN(n54146) );
  INV_X1 U55696 ( .I(n54186), .ZN(n54145) );
  AOI22_X1 U55697 ( .A1(n54147), .A2(n54146), .B1(n54145), .B2(n54144), .ZN(
        n54152) );
  NAND3_X1 U55698 ( .A1(n63726), .A2(n54197), .A3(n2984), .ZN(n54149) );
  NAND3_X1 U55700 ( .A1(n54150), .A2(n54149), .A3(n54148), .ZN(n54151) );
  NAND2_X1 U55703 ( .A1(n54189), .A2(n2984), .ZN(n54179) );
  AOI21_X1 U55705 ( .A1(n54198), .A2(n25299), .B(n54207), .ZN(n54156) );
  NAND3_X1 U55706 ( .A1(n9968), .A2(n26008), .A3(n63726), .ZN(n54155) );
  NAND3_X1 U55707 ( .A1(n54157), .A2(n54156), .A3(n54155), .ZN(n54167) );
  NAND2_X1 U55708 ( .A1(n54158), .A2(n54198), .ZN(n54160) );
  AOI22_X1 U55709 ( .A1(n54161), .A2(n54160), .B1(n54175), .B2(n54159), .ZN(
        n54166) );
  NAND4_X1 U55710 ( .A1(n54172), .A2(n54192), .A3(n54162), .A4(n54207), .ZN(
        n54165) );
  NAND2_X1 U55711 ( .A1(n54189), .A2(n26008), .ZN(n54202) );
  XOR2_X1 U55714 ( .A1(n54169), .A2(n54168), .Z(Plaintext[57]) );
  NAND2_X1 U55716 ( .A1(n54197), .A2(n54207), .ZN(n54177) );
  NAND3_X1 U55717 ( .A1(n54172), .A2(n54171), .A3(n54177), .ZN(n54173) );
  OAI22_X1 U55718 ( .A1(n54174), .A2(n54173), .B1(n10480), .B2(n63726), .ZN(
        n54183) );
  OAI22_X1 U55719 ( .A1(n9968), .A2(n54176), .B1(n54201), .B2(n26008), .ZN(
        n54181) );
  NAND2_X1 U55720 ( .A1(n54177), .A2(n54192), .ZN(n54178) );
  NOR2_X1 U55721 ( .A1(n54179), .A2(n54178), .ZN(n54180) );
  NOR2_X1 U55722 ( .A1(n54181), .A2(n54180), .ZN(n54182) );
  NAND2_X1 U55723 ( .A1(n54183), .A2(n54182), .ZN(n54184) );
  XOR2_X1 U55724 ( .A1(n54184), .A2(n54185), .Z(Plaintext[58]) );
  NAND2_X1 U55727 ( .A1(n54259), .A2(n1256), .ZN(n54251) );
  INV_X1 U55729 ( .I(n54213), .ZN(n54212) );
  OAI21_X1 U55732 ( .A1(n54277), .A2(n23731), .B(n54221), .ZN(n54224) );
  NAND3_X1 U55733 ( .A1(n54224), .A2(n54251), .A3(n54223), .ZN(n54230) );
  OAI21_X1 U55734 ( .A1(n54225), .A2(n54268), .B(n19404), .ZN(n54229) );
  NOR2_X1 U55735 ( .A1(n54277), .A2(n19404), .ZN(n54226) );
  NAND2_X1 U55736 ( .A1(n54232), .A2(n22315), .ZN(n54237) );
  INV_X1 U55737 ( .I(n54233), .ZN(n54236) );
  NAND2_X1 U55739 ( .A1(n54281), .A2(n54271), .ZN(n54241) );
  NAND2_X1 U55740 ( .A1(n1256), .A2(n1280), .ZN(n54258) );
  NAND2_X1 U55741 ( .A1(n54258), .A2(n54280), .ZN(n54240) );
  NAND4_X1 U55742 ( .A1(n54242), .A2(n54282), .A3(n54241), .A4(n54240), .ZN(
        n54247) );
  NAND2_X1 U55743 ( .A1(n54266), .A2(n54285), .ZN(n54244) );
  NAND2_X1 U55744 ( .A1(n54244), .A2(n54273), .ZN(n54245) );
  XOR2_X1 U55745 ( .A1(n54250), .A2(n54249), .Z(Plaintext[63]) );
  NAND3_X1 U55746 ( .A1(n54282), .A2(n54254), .A3(n54258), .ZN(n54255) );
  NAND2_X1 U55747 ( .A1(n54255), .A2(n54285), .ZN(n54262) );
  NAND4_X1 U55748 ( .A1(n22545), .A2(n54258), .A3(n54268), .A4(n57202), .ZN(
        n54260) );
  AOI21_X1 U55750 ( .A1(n54271), .A2(n54270), .B(n54269), .ZN(n54275) );
  AOI22_X1 U55752 ( .A1(n54276), .A2(n54275), .B1(n54274), .B2(n54273), .ZN(
        n54288) );
  OAI21_X1 U55755 ( .A1(n54286), .A2(n54285), .B(n54284), .ZN(n54287) );
  NOR2_X1 U55759 ( .A1(n54963), .A2(n54625), .ZN(n54298) );
  AOI22_X1 U55760 ( .A1(n54972), .A2(n54971), .B1(n54298), .B2(n54970), .ZN(
        n54304) );
  INV_X1 U55761 ( .I(n54961), .ZN(n54299) );
  NAND2_X1 U55765 ( .A1(n4504), .A2(n10523), .ZN(n54328) );
  NAND2_X1 U55766 ( .A1(n54366), .A2(n54362), .ZN(n54332) );
  NAND2_X1 U55767 ( .A1(n54822), .A2(n54440), .ZN(n54333) );
  MUX2_X1 U55769 ( .I0(n54657), .I1(n54437), .S(n54659), .Z(n54338) );
  NAND3_X1 U55770 ( .A1(n19137), .A2(n23849), .A3(n1607), .ZN(n54334) );
  NAND2_X1 U55771 ( .A1(n54383), .A2(n271), .ZN(n54355) );
  NAND2_X1 U55772 ( .A1(n61829), .A2(n1367), .ZN(n54356) );
  NOR2_X1 U55774 ( .A1(n54383), .A2(n54390), .ZN(n54365) );
  INV_X1 U55776 ( .I(n54363), .ZN(n54361) );
  NAND2_X1 U55777 ( .A1(n54361), .A2(n54417), .ZN(n54364) );
  AOI22_X1 U55778 ( .A1(n54365), .A2(n54364), .B1(n54393), .B2(n54363), .ZN(
        n54375) );
  NAND2_X1 U55779 ( .A1(n54366), .A2(n54400), .ZN(n54367) );
  NAND3_X1 U55780 ( .A1(n54387), .A2(n54367), .A3(n54390), .ZN(n54374) );
  NAND4_X1 U55782 ( .A1(n54372), .A2(n54371), .A3(n54370), .A4(n54408), .ZN(
        n54373) );
  AOI21_X1 U55783 ( .A1(n54375), .A2(n54374), .B(n54373), .ZN(n54378) );
  XOR2_X1 U55784 ( .A1(n54378), .A2(n54377), .Z(Plaintext[67]) );
  AOI21_X1 U55785 ( .A1(n54390), .A2(n54380), .B(n1367), .ZN(n54382) );
  NAND3_X1 U55787 ( .A1(n4688), .A2(n20985), .A3(n271), .ZN(n54381) );
  NAND4_X1 U55788 ( .A1(n54384), .A2(n54382), .A3(n54415), .A4(n54381), .ZN(
        n54385) );
  AOI21_X1 U55789 ( .A1(n271), .A2(n15202), .B(n54400), .ZN(n54396) );
  INV_X1 U55791 ( .I(n54400), .ZN(n54401) );
  NAND3_X1 U55792 ( .A1(n54401), .A2(n7138), .A3(n4688), .ZN(n54405) );
  NOR2_X1 U55793 ( .A1(n54419), .A2(n54418), .ZN(n54420) );
  NAND2_X1 U55794 ( .A1(n54425), .A2(n54424), .ZN(n54426) );
  NAND4_X1 U55795 ( .A1(n54427), .A2(n4688), .A3(n54392), .A4(n54426), .ZN(
        n54428) );
  INV_X1 U55796 ( .I(n54785), .ZN(n54432) );
  NOR3_X1 U55797 ( .A1(n59081), .A2(n21877), .A3(n54433), .ZN(n54434) );
  AOI21_X1 U55798 ( .A1(n54438), .A2(n62768), .B(n23849), .ZN(n54439) );
  MUX2_X1 U55799 ( .I0(n20095), .I1(n54439), .S(n54825), .Z(n54450) );
  NAND3_X1 U55802 ( .A1(n6312), .A2(n6311), .A3(n54659), .ZN(n54442) );
  NOR2_X1 U55804 ( .A1(n54445), .A2(n54444), .ZN(n54448) );
  OAI21_X1 U55805 ( .A1(n54455), .A2(n54454), .B(n55022), .ZN(n54456) );
  NOR2_X1 U55806 ( .A1(n54466), .A2(n23897), .ZN(n54467) );
  NOR2_X1 U55807 ( .A1(n54598), .A2(n64129), .ZN(n54468) );
  NAND2_X1 U55808 ( .A1(n54471), .A2(n54470), .ZN(n54475) );
  NOR2_X1 U55810 ( .A1(n54530), .A2(n54531), .ZN(n54510) );
  NOR2_X1 U55812 ( .A1(n7518), .A2(n54625), .ZN(n54478) );
  AOI21_X1 U55813 ( .A1(n54965), .A2(n54970), .B(n54478), .ZN(n54488) );
  XOR2_X1 U55814 ( .A1(n54802), .A2(n54487), .Z(n54479) );
  AOI21_X1 U55815 ( .A1(n54479), .A2(n54481), .B(n1146), .ZN(n54485) );
  NAND2_X1 U55816 ( .A1(n54626), .A2(n54963), .ZN(n54480) );
  NOR2_X1 U55817 ( .A1(n54480), .A2(n61736), .ZN(n54484) );
  AOI21_X1 U55818 ( .A1(n54482), .A2(n54806), .B(n54481), .ZN(n54483) );
  NAND2_X1 U55819 ( .A1(n54493), .A2(n7532), .ZN(n54494) );
  NAND2_X1 U55821 ( .A1(n4232), .A2(n65013), .ZN(n54511) );
  NAND2_X1 U55822 ( .A1(n54513), .A2(n54566), .ZN(n54514) );
  NAND2_X1 U55825 ( .A1(n54525), .A2(n54581), .ZN(n54526) );
  NAND2_X1 U55826 ( .A1(n54561), .A2(n22572), .ZN(n54576) );
  NAND2_X1 U55829 ( .A1(n54573), .A2(n54565), .ZN(n54529) );
  NAND3_X1 U55830 ( .A1(n54530), .A2(n54548), .A3(n54529), .ZN(n54535) );
  INV_X1 U55833 ( .I(n54567), .ZN(n54533) );
  NAND2_X1 U55834 ( .A1(n54533), .A2(n54532), .ZN(n54534) );
  AOI21_X1 U55835 ( .A1(n54564), .A2(n58810), .B(n54538), .ZN(n54555) );
  NAND2_X1 U55836 ( .A1(n60433), .A2(n54565), .ZN(n54539) );
  OAI21_X1 U55837 ( .A1(n60433), .A2(n58810), .B(n54541), .ZN(n54544) );
  OAI21_X1 U55838 ( .A1(n54545), .A2(n54544), .B(n54548), .ZN(n54554) );
  NOR2_X1 U55839 ( .A1(n54568), .A2(n22572), .ZN(n54552) );
  AOI21_X1 U55841 ( .A1(n54552), .A2(n54551), .B(n54550), .ZN(n54553) );
  NAND2_X1 U55842 ( .A1(n54561), .A2(n54560), .ZN(n54579) );
  OAI21_X1 U55844 ( .A1(n54580), .A2(n54579), .B(n54578), .ZN(n54585) );
  NAND3_X1 U55845 ( .A1(n54583), .A2(n54582), .A3(n54581), .ZN(n54584) );
  XOR2_X1 U55846 ( .A1(n54597), .A2(n54594), .Z(n54604) );
  NAND2_X1 U55847 ( .A1(n54601), .A2(n54595), .ZN(n54603) );
  NAND3_X1 U55849 ( .A1(n54601), .A2(n54600), .A3(n54599), .ZN(n54602) );
  NOR2_X1 U55851 ( .A1(n54614), .A2(n21877), .ZN(n54609) );
  OAI21_X1 U55852 ( .A1(n54609), .A2(n54608), .B(n54607), .ZN(n54610) );
  NAND2_X1 U55853 ( .A1(n54973), .A2(n58978), .ZN(n54621) );
  NAND2_X1 U55854 ( .A1(n54619), .A2(n54626), .ZN(n54620) );
  MUX2_X1 U55855 ( .I0(n54621), .I1(n54620), .S(n54970), .Z(n54666) );
  AOI21_X1 U55857 ( .A1(n54624), .A2(n54623), .B(n58978), .ZN(n54633) );
  INV_X1 U55858 ( .I(n54974), .ZN(n54628) );
  AOI21_X1 U55860 ( .A1(n54630), .A2(n54807), .B(n54629), .ZN(n54631) );
  NOR2_X1 U55861 ( .A1(n54728), .A2(n54741), .ZN(n54757) );
  NAND2_X1 U55862 ( .A1(n55024), .A2(n4504), .ZN(n54635) );
  AOI21_X1 U55864 ( .A1(n54647), .A2(n63194), .B(n55265), .ZN(n54686) );
  NAND2_X1 U55866 ( .A1(n2489), .A2(n15023), .ZN(n54656) );
  NAND3_X1 U55868 ( .A1(n54660), .A2(n54659), .A3(n54658), .ZN(n54694) );
  OAI21_X1 U55871 ( .A1(n65124), .A2(n54757), .B(n54661), .ZN(n54675) );
  NOR2_X1 U55872 ( .A1(n54769), .A2(n54762), .ZN(n54664) );
  OAI21_X1 U55873 ( .A1(n54668), .A2(n54738), .B(n19492), .ZN(n54673) );
  NOR2_X1 U55874 ( .A1(n57201), .A2(n59051), .ZN(n54671) );
  NAND2_X1 U55875 ( .A1(n54769), .A2(n14848), .ZN(n54752) );
  NAND2_X1 U55876 ( .A1(n54741), .A2(n57201), .ZN(n54677) );
  AOI21_X1 U55878 ( .A1(n54718), .A2(n54677), .B(n54736), .ZN(n54678) );
  NOR2_X1 U55879 ( .A1(n54679), .A2(n54678), .ZN(n54707) );
  NAND3_X1 U55880 ( .A1(n63473), .A2(n22385), .A3(n54727), .ZN(n54680) );
  OAI22_X1 U55881 ( .A1(n54682), .A2(n54680), .B1(n19492), .B2(n54759), .ZN(
        n54681) );
  NOR2_X1 U55882 ( .A1(n54681), .A2(n54737), .ZN(n54706) );
  INV_X1 U55883 ( .I(n54682), .ZN(n54702) );
  NAND2_X1 U55884 ( .A1(n54683), .A2(n64255), .ZN(n54685) );
  AOI21_X1 U55885 ( .A1(n54686), .A2(n54685), .B(n54684), .ZN(n54687) );
  NAND2_X1 U55886 ( .A1(n54768), .A2(n54687), .ZN(n54699) );
  INV_X1 U55887 ( .I(n54688), .ZN(n54690) );
  NAND2_X1 U55888 ( .A1(n54690), .A2(n15040), .ZN(n54693) );
  NAND4_X1 U55889 ( .A1(n54694), .A2(n54693), .A3(n54692), .A4(n54691), .ZN(
        n54696) );
  OAI21_X1 U55890 ( .A1(n54697), .A2(n54696), .B(n54695), .ZN(n54698) );
  NAND2_X1 U55892 ( .A1(n54741), .A2(n65124), .ZN(n54703) );
  NAND3_X1 U55893 ( .A1(n57201), .A2(n22122), .A3(n54769), .ZN(n54711) );
  INV_X1 U55895 ( .I(n54724), .ZN(n54713) );
  AOI21_X1 U55896 ( .A1(n54728), .A2(n14848), .B(n22122), .ZN(n54720) );
  NAND2_X1 U55897 ( .A1(n19492), .A2(n54768), .ZN(n54751) );
  INV_X1 U55898 ( .I(n54718), .ZN(n54719) );
  AOI21_X1 U55899 ( .A1(n54720), .A2(n54751), .B(n54719), .ZN(n54733) );
  NAND4_X1 U55900 ( .A1(n54725), .A2(n54724), .A3(n23448), .A4(n54723), .ZN(
        n54732) );
  NAND3_X1 U55901 ( .A1(n54728), .A2(n54741), .A3(n54768), .ZN(n54729) );
  NAND4_X1 U55902 ( .A1(n54730), .A2(n61057), .A3(n54736), .A4(n54729), .ZN(
        n54731) );
  INV_X1 U55903 ( .I(n54736), .ZN(n54739) );
  AOI21_X1 U55904 ( .A1(n54739), .A2(n54738), .B(n54737), .ZN(n54747) );
  NAND2_X1 U55906 ( .A1(n54742), .A2(n54741), .ZN(n54743) );
  NAND3_X1 U55907 ( .A1(n54743), .A2(n54768), .A3(n54771), .ZN(n54745) );
  NAND3_X1 U55908 ( .A1(n54771), .A2(n61057), .A3(n54750), .ZN(n54744) );
  XOR2_X1 U55909 ( .A1(n54749), .A2(n9871), .Z(Plaintext[82]) );
  OR2_X1 U55910 ( .A1(n54754), .A2(n63473), .Z(n54756) );
  AOI22_X1 U55911 ( .A1(n54757), .A2(n54756), .B1(n54755), .B2(n61057), .ZN(
        n54774) );
  NOR2_X1 U55912 ( .A1(n54759), .A2(n14848), .ZN(n54763) );
  NOR2_X1 U55913 ( .A1(n57201), .A2(n54767), .ZN(n54761) );
  OAI21_X1 U55915 ( .A1(n19492), .A2(n54767), .B(n54766), .ZN(n54770) );
  NAND4_X1 U55916 ( .A1(n54771), .A2(n54770), .A3(n54769), .A4(n54768), .ZN(
        n54772) );
  NAND4_X1 U55917 ( .A1(n54775), .A2(n54774), .A3(n54773), .A4(n54772), .ZN(
        n54777) );
  XOR2_X1 U55918 ( .A1(n54777), .A2(n54776), .Z(Plaintext[83]) );
  NAND2_X1 U55919 ( .A1(n54783), .A2(n54782), .ZN(n54784) );
  OAI22_X1 U55920 ( .A1(n65010), .A2(n54982), .B1(n54990), .B2(n55398), .ZN(
        n54789) );
  NAND2_X1 U55921 ( .A1(n61895), .A2(n54786), .ZN(n54788) );
  NOR2_X1 U55922 ( .A1(n55244), .A2(n55415), .ZN(n54787) );
  NAND2_X1 U55924 ( .A1(n55416), .A2(n24075), .ZN(n54794) );
  OAI22_X1 U55926 ( .A1(n55246), .A2(n54796), .B1(n54982), .B2(n55404), .ZN(
        n54797) );
  NAND2_X1 U55927 ( .A1(n1146), .A2(n54961), .ZN(n54799) );
  NOR2_X1 U55928 ( .A1(n54802), .A2(n54801), .ZN(n54803) );
  OAI21_X1 U55929 ( .A1(n61736), .A2(n54803), .B(n54971), .ZN(n54804) );
  NAND2_X1 U55930 ( .A1(n23122), .A2(n58491), .ZN(n54809) );
  NAND2_X1 U55931 ( .A1(n54963), .A2(n61509), .ZN(n54811) );
  NOR2_X1 U55934 ( .A1(n62768), .A2(n62986), .ZN(n54821) );
  NAND2_X1 U55936 ( .A1(n54824), .A2(n18629), .ZN(n54830) );
  OAI21_X1 U55937 ( .A1(n18629), .A2(n54827), .B(n54826), .ZN(n54829) );
  NAND2_X1 U55940 ( .A1(n61870), .A2(n16846), .ZN(n54838) );
  OAI21_X1 U55941 ( .A1(n55275), .A2(n19167), .B(n58283), .ZN(n54839) );
  NAND2_X1 U55942 ( .A1(n21268), .A2(n54839), .ZN(n54840) );
  AOI22_X1 U55943 ( .A1(n55266), .A2(n61081), .B1(n12074), .B2(n5570), .ZN(
        n54845) );
  NOR2_X1 U55944 ( .A1(n14635), .A2(n54892), .ZN(n54847) );
  AOI22_X1 U55945 ( .A1(n7956), .A2(n54846), .B1(n15937), .B2(n54847), .ZN(
        n54868) );
  NAND2_X1 U55947 ( .A1(n1373), .A2(n22760), .ZN(n54857) );
  OAI21_X1 U55948 ( .A1(n10523), .A2(n54857), .B(n55020), .ZN(n54859) );
  NAND3_X1 U55950 ( .A1(n55016), .A2(n55022), .A3(n3916), .ZN(n54861) );
  NAND2_X1 U55951 ( .A1(n13671), .A2(n54904), .ZN(n54866) );
  INV_X1 U55952 ( .I(n54871), .ZN(n54872) );
  INV_X1 U55953 ( .I(n54874), .ZN(n54875) );
  NOR2_X1 U55954 ( .A1(n54915), .A2(n63022), .ZN(n54879) );
  NOR4_X1 U55955 ( .A1(n54880), .A2(n2049), .A3(n63022), .A4(n20752), .ZN(
        n54881) );
  NOR3_X1 U55956 ( .A1(n54882), .A2(n54920), .A3(n54881), .ZN(n54885) );
  NAND2_X1 U55957 ( .A1(n2049), .A2(n63022), .ZN(n54925) );
  OAI21_X1 U55958 ( .A1(n54925), .A2(n736), .B(n54892), .ZN(n54883) );
  INV_X1 U55959 ( .I(n54929), .ZN(n54890) );
  INV_X1 U55961 ( .I(n54911), .ZN(n54891) );
  AOI22_X1 U55962 ( .A1(n54929), .A2(n54893), .B1(n4152), .B2(n2329), .ZN(
        n54895) );
  NAND2_X1 U55964 ( .A1(n54914), .A2(n63022), .ZN(n54899) );
  MUX2_X1 U55965 ( .I0(n54900), .I1(n54899), .S(n4152), .Z(n54909) );
  NAND3_X1 U55966 ( .A1(n54905), .A2(n54929), .A3(n54904), .ZN(n54906) );
  NOR3_X1 U55967 ( .A1(n54921), .A2(n54914), .A3(n63022), .ZN(n54916) );
  INV_X1 U55968 ( .I(n54915), .ZN(n54930) );
  XOR2_X1 U55969 ( .A1(n54919), .A2(n54918), .Z(Plaintext[88]) );
  NOR2_X1 U55970 ( .A1(n54925), .A2(n2329), .ZN(n54927) );
  OAI22_X1 U55971 ( .A1(n54929), .A2(n4152), .B1(n2049), .B2(n54928), .ZN(
        n54931) );
  NAND2_X1 U55972 ( .A1(n54931), .A2(n54930), .ZN(n54932) );
  NOR2_X1 U55973 ( .A1(n57404), .A2(n60439), .ZN(n54942) );
  MUX2_X1 U55978 ( .I0(n55244), .I1(n54990), .S(n55415), .Z(n54989) );
  NAND3_X1 U55979 ( .A1(n55407), .A2(n54990), .A3(n55406), .ZN(n54987) );
  INV_X1 U55980 ( .I(n55012), .ZN(n54994) );
  MUX2_X1 U55981 ( .I0(n65010), .I1(n54990), .S(n55412), .Z(n54992) );
  NOR2_X1 U55982 ( .A1(n65011), .A2(n61065), .ZN(n54991) );
  OAI21_X1 U55983 ( .A1(n54992), .A2(n55252), .B(n54991), .ZN(n54993) );
  NAND2_X1 U55984 ( .A1(n55042), .A2(n55075), .ZN(n55030) );
  NAND2_X1 U55985 ( .A1(n23275), .A2(n55440), .ZN(n55000) );
  XOR2_X1 U55987 ( .A1(n55433), .A2(n55440), .Z(n55001) );
  INV_X1 U55988 ( .I(n55002), .ZN(n55003) );
  INV_X1 U55989 ( .I(n55322), .ZN(n55005) );
  AOI21_X1 U55990 ( .A1(n18247), .A2(n55020), .B(n55019), .ZN(n55021) );
  NAND2_X1 U55991 ( .A1(n55024), .A2(n59713), .ZN(n55025) );
  NAND2_X1 U55993 ( .A1(n55031), .A2(n55076), .ZN(n55033) );
  NAND3_X1 U55996 ( .A1(n55042), .A2(n9067), .A3(n62822), .ZN(n55044) );
  AOI21_X1 U55998 ( .A1(n55044), .A2(n55043), .B(n55089), .ZN(n55050) );
  NAND2_X1 U56000 ( .A1(n55056), .A2(n55089), .ZN(n55046) );
  NOR3_X1 U56001 ( .A1(n55051), .A2(n55050), .A3(n55049), .ZN(n55054) );
  XOR2_X1 U56002 ( .A1(n55054), .A2(n55053), .Z(Plaintext[91]) );
  NAND3_X1 U56004 ( .A1(n59533), .A2(n55075), .A3(n591), .ZN(n55059) );
  NOR2_X1 U56005 ( .A1(n55089), .A2(n55061), .ZN(n55063) );
  INV_X1 U56006 ( .I(n55082), .ZN(n55062) );
  INV_X1 U56007 ( .I(n55065), .ZN(n55067) );
  NOR2_X1 U56008 ( .A1(n55067), .A2(n55066), .ZN(n55071) );
  OAI22_X1 U56009 ( .A1(n55068), .A2(n55077), .B1(n9067), .B2(n674), .ZN(
        n55069) );
  NAND2_X1 U56010 ( .A1(n55074), .A2(n55069), .ZN(n55070) );
  INV_X1 U56012 ( .I(n55074), .ZN(n55081) );
  NOR2_X1 U56013 ( .A1(n55075), .A2(n55101), .ZN(n55080) );
  NOR2_X1 U56014 ( .A1(n55077), .A2(n55076), .ZN(n55078) );
  AOI22_X1 U56015 ( .A1(n55081), .A2(n55080), .B1(n55079), .B2(n55078), .ZN(
        n55086) );
  AOI21_X1 U56020 ( .A1(n8027), .A2(n55140), .B(n55110), .ZN(n55117) );
  INV_X1 U56021 ( .I(n55146), .ZN(n55121) );
  NOR2_X1 U56022 ( .A1(n55119), .A2(n55168), .ZN(n55113) );
  OAI21_X1 U56023 ( .A1(n55132), .A2(n55168), .B(n1593), .ZN(n55114) );
  NAND4_X1 U56024 ( .A1(n55115), .A2(n55114), .A3(n55140), .A4(n55165), .ZN(
        n55116) );
  NOR2_X1 U56025 ( .A1(n55144), .A2(n55171), .ZN(n55125) );
  NOR3_X1 U56027 ( .A1(n55159), .A2(n55145), .A3(n11353), .ZN(n55124) );
  NAND2_X1 U56028 ( .A1(n55119), .A2(n55165), .ZN(n55120) );
  AOI21_X1 U56029 ( .A1(n55121), .A2(n55120), .B(n55166), .ZN(n55123) );
  INV_X1 U56031 ( .I(n55126), .ZN(n55127) );
  XOR2_X1 U56032 ( .A1(n55128), .A2(n55127), .Z(Plaintext[98]) );
  NAND2_X1 U56033 ( .A1(n55163), .A2(n55131), .ZN(n55130) );
  NAND2_X1 U56034 ( .A1(n55156), .A2(n10310), .ZN(n55129) );
  AOI21_X1 U56035 ( .A1(n55130), .A2(n55157), .B(n55129), .ZN(n55138) );
  NAND2_X1 U56036 ( .A1(n55143), .A2(n8027), .ZN(n55137) );
  NOR2_X1 U56037 ( .A1(n10310), .A2(n55170), .ZN(n55152) );
  OAI21_X1 U56038 ( .A1(n55153), .A2(n55152), .B(n55161), .ZN(n55155) );
  NOR2_X1 U56039 ( .A1(n55157), .A2(n55156), .ZN(n55158) );
  OAI21_X1 U56041 ( .A1(n55163), .A2(n55166), .B(n55162), .ZN(n55172) );
  NAND2_X1 U56042 ( .A1(n55165), .A2(n11353), .ZN(n55167) );
  AOI22_X1 U56043 ( .A1(n55172), .A2(n55171), .B1(n7986), .B2(n55169), .ZN(
        n55173) );
  INV_X1 U56044 ( .I(n55216), .ZN(n55209) );
  NOR2_X1 U56046 ( .A1(n55208), .A2(n20839), .ZN(n55181) );
  INV_X1 U56048 ( .I(n55197), .ZN(n55186) );
  NAND2_X1 U56049 ( .A1(n55222), .A2(n55225), .ZN(n55183) );
  NOR2_X1 U56050 ( .A1(n55183), .A2(n20839), .ZN(n55184) );
  OAI22_X1 U56051 ( .A1(n55186), .A2(n55185), .B1(n55184), .B2(n55218), .ZN(
        n55187) );
  MUX2_X1 U56052 ( .I0(n58813), .I1(n55218), .S(n55203), .Z(n55192) );
  NAND2_X1 U56053 ( .A1(n55192), .A2(n17155), .ZN(n55195) );
  NAND3_X1 U56054 ( .A1(n55233), .A2(n62711), .A3(n17155), .ZN(n55193) );
  NOR2_X1 U56055 ( .A1(n55236), .A2(n20839), .ZN(n55201) );
  NAND2_X1 U56057 ( .A1(n55202), .A2(n55208), .ZN(n55206) );
  XOR2_X1 U56058 ( .A1(n55207), .A2(n24046), .Z(Plaintext[105]) );
  NAND3_X1 U56059 ( .A1(n55210), .A2(n55209), .A3(n55208), .ZN(n55215) );
  NAND2_X1 U56061 ( .A1(n16978), .A2(n1587), .ZN(n55211) );
  NAND3_X1 U56062 ( .A1(n55211), .A2(n62711), .A3(n55217), .ZN(n55212) );
  XOR2_X1 U56064 ( .A1(n55221), .A2(n1902), .Z(Plaintext[106]) );
  MUX2_X1 U56065 ( .I0(n55228), .I1(n55227), .S(n55226), .Z(n55241) );
  NAND2_X1 U56066 ( .A1(n1587), .A2(n16383), .ZN(n55229) );
  MUX2_X1 U56067 ( .I0(n55237), .I1(n55236), .S(n55235), .Z(n55238) );
  NAND2_X1 U56069 ( .A1(n55245), .A2(n55244), .ZN(n55254) );
  NAND2_X1 U56071 ( .A1(n23763), .A2(n22807), .ZN(n55249) );
  OAI22_X1 U56073 ( .A1(n64813), .A2(n55403), .B1(n55257), .B2(n55256), .ZN(
        n55258) );
  NAND2_X1 U56074 ( .A1(n58283), .A2(n65101), .ZN(n55268) );
  NOR2_X1 U56076 ( .A1(n58283), .A2(n1613), .ZN(n55276) );
  NAND3_X1 U56078 ( .A1(n55279), .A2(n55472), .A3(n55475), .ZN(n55283) );
  NAND2_X1 U56079 ( .A1(n55474), .A2(n2180), .ZN(n55281) );
  NAND2_X1 U56080 ( .A1(n55287), .A2(n61282), .ZN(n55288) );
  NOR2_X1 U56081 ( .A1(n15730), .A2(n64970), .ZN(n55290) );
  MUX2_X1 U56082 ( .I0(n59040), .I1(n55295), .S(n65283), .Z(n55297) );
  NOR2_X1 U56083 ( .A1(n55300), .A2(n55299), .ZN(n55301) );
  NAND2_X1 U56084 ( .A1(n55345), .A2(n55362), .ZN(n55327) );
  NAND3_X1 U56085 ( .A1(n55310), .A2(n55317), .A3(n55442), .ZN(n55311) );
  NAND2_X1 U56086 ( .A1(n55317), .A2(n23522), .ZN(n55319) );
  AOI21_X1 U56087 ( .A1(n55320), .A2(n55319), .B(n55318), .ZN(n55326) );
  NAND3_X1 U56089 ( .A1(n55327), .A2(n21210), .A3(n58828), .ZN(n55329) );
  OAI21_X1 U56091 ( .A1(n55386), .A2(n55332), .B(n14428), .ZN(n55333) );
  NAND2_X1 U56092 ( .A1(n55334), .A2(n55333), .ZN(n55336) );
  XOR2_X1 U56093 ( .A1(n55336), .A2(n55335), .Z(Plaintext[108]) );
  NAND2_X1 U56094 ( .A1(n19973), .A2(n24063), .ZN(n55347) );
  AOI21_X1 U56096 ( .A1(n58828), .A2(n9777), .B(n55382), .ZN(n55346) );
  NAND2_X1 U56097 ( .A1(n55355), .A2(n15936), .ZN(n55354) );
  NAND3_X1 U56098 ( .A1(n55350), .A2(n15703), .A3(n21210), .ZN(n55353) );
  INV_X1 U56099 ( .I(n55355), .ZN(n55358) );
  NOR2_X1 U56101 ( .A1(n55361), .A2(n55360), .ZN(n55367) );
  OAI22_X1 U56102 ( .A1(n55364), .A2(n19973), .B1(n55363), .B2(n55362), .ZN(
        n55365) );
  NAND2_X1 U56103 ( .A1(n55365), .A2(n55389), .ZN(n55366) );
  NAND2_X1 U56104 ( .A1(n55367), .A2(n55366), .ZN(n55369) );
  XOR2_X1 U56105 ( .A1(n55369), .A2(n55368), .Z(Plaintext[111]) );
  INV_X1 U56106 ( .I(n55372), .ZN(n55370) );
  NAND2_X1 U56107 ( .A1(n55370), .A2(n9777), .ZN(n55371) );
  OAI21_X1 U56108 ( .A1(n55382), .A2(n64598), .B(n55372), .ZN(n55374) );
  INV_X1 U56109 ( .I(n55377), .ZN(n55378) );
  XOR2_X1 U56110 ( .A1(n55380), .A2(n55379), .Z(Plaintext[112]) );
  OAI21_X1 U56111 ( .A1(n18135), .A2(n55383), .B(n55382), .ZN(n55394) );
  XOR2_X1 U56115 ( .A1(n55396), .A2(n55395), .Z(Plaintext[113]) );
  NOR2_X1 U56116 ( .A1(n55398), .A2(n64813), .ZN(n55399) );
  OAI21_X1 U56117 ( .A1(n55413), .A2(n55399), .B(n62988), .ZN(n55411) );
  NAND3_X1 U56118 ( .A1(n62988), .A2(n55401), .A3(n197), .ZN(n55410) );
  AOI21_X1 U56121 ( .A1(n1615), .A2(n55721), .B(n1324), .ZN(n55426) );
  OAI21_X1 U56122 ( .A1(n1324), .A2(n23360), .B(n55915), .ZN(n55428) );
  NAND3_X1 U56123 ( .A1(n55718), .A2(n55428), .A3(n50932), .ZN(n55432) );
  NAND3_X1 U56124 ( .A1(n55430), .A2(n55429), .A3(n20653), .ZN(n55431) );
  NAND2_X1 U56125 ( .A1(n55569), .A2(n1592), .ZN(n55518) );
  NAND2_X1 U56126 ( .A1(n55434), .A2(n55435), .ZN(n55439) );
  NOR2_X1 U56127 ( .A1(n24454), .A2(n23522), .ZN(n55446) );
  NAND2_X1 U56128 ( .A1(n55565), .A2(n21272), .ZN(n55461) );
  INV_X1 U56129 ( .I(n55965), .ZN(n55447) );
  NAND3_X1 U56130 ( .A1(n55450), .A2(n55449), .A3(n55448), .ZN(n55460) );
  INV_X1 U56131 ( .I(n4830), .ZN(n55451) );
  NAND2_X1 U56132 ( .A1(n55453), .A2(n55967), .ZN(n55454) );
  NAND3_X1 U56133 ( .A1(n55454), .A2(n55968), .A3(n55975), .ZN(n55459) );
  NAND2_X1 U56134 ( .A1(n14142), .A2(n55680), .ZN(n55455) );
  NAND4_X1 U56135 ( .A1(n55966), .A2(n55456), .A3(n55973), .A4(n55455), .ZN(
        n55457) );
  AOI21_X1 U56137 ( .A1(n55518), .A2(n55461), .B(n55549), .ZN(n55508) );
  AOI22_X1 U56138 ( .A1(n55739), .A2(n248), .B1(n55740), .B2(n55473), .ZN(
        n55462) );
  NAND2_X1 U56140 ( .A1(n55462), .A2(n55733), .ZN(n55468) );
  NOR2_X1 U56141 ( .A1(n55478), .A2(n55463), .ZN(n55466) );
  NOR2_X1 U56144 ( .A1(n55473), .A2(n57720), .ZN(n55477) );
  NAND3_X1 U56147 ( .A1(n55480), .A2(n55479), .A3(n22588), .ZN(n55481) );
  NAND3_X1 U56149 ( .A1(n55489), .A2(n55488), .A3(n55487), .ZN(n55493) );
  NAND2_X1 U56150 ( .A1(n55689), .A2(n55690), .ZN(n55491) );
  NAND2_X1 U56151 ( .A1(n55491), .A2(n1609), .ZN(n55492) );
  NAND2_X1 U56152 ( .A1(n55496), .A2(n55495), .ZN(n55501) );
  NOR2_X1 U56153 ( .A1(n10414), .A2(n51961), .ZN(n55500) );
  OAI22_X1 U56154 ( .A1(n55498), .A2(n55690), .B1(n55695), .B2(n64019), .ZN(
        n55499) );
  AOI22_X1 U56155 ( .A1(n55595), .A2(n55550), .B1(n55587), .B2(n19183), .ZN(
        n55507) );
  NAND2_X1 U56156 ( .A1(n19183), .A2(n55569), .ZN(n55502) );
  AOI21_X1 U56157 ( .A1(n55575), .A2(n55502), .B(n55592), .ZN(n55506) );
  OAI21_X1 U56158 ( .A1(n1592), .A2(n55597), .B(n21273), .ZN(n55504) );
  AOI22_X1 U56160 ( .A1(n55508), .A2(n55507), .B1(n55506), .B2(n55505), .ZN(
        n55515) );
  INV_X1 U56161 ( .I(n55587), .ZN(n55538) );
  NOR2_X1 U56162 ( .A1(n55575), .A2(n55550), .ZN(n55593) );
  NOR2_X1 U56163 ( .A1(n55595), .A2(n21273), .ZN(n55509) );
  AOI22_X1 U56164 ( .A1(n55566), .A2(n55538), .B1(n55593), .B2(n55509), .ZN(
        n55514) );
  AOI21_X1 U56165 ( .A1(n55584), .A2(n55570), .B(n55509), .ZN(n55512) );
  NAND2_X1 U56166 ( .A1(n55565), .A2(n55550), .ZN(n55510) );
  AOI21_X1 U56167 ( .A1(n55570), .A2(n55510), .B(n55575), .ZN(n55511) );
  NAND2_X1 U56168 ( .A1(n55512), .A2(n55511), .ZN(n55513) );
  NOR2_X1 U56171 ( .A1(n55590), .A2(n55547), .ZN(n55539) );
  NOR2_X1 U56172 ( .A1(n55539), .A2(n55567), .ZN(n55524) );
  OAI21_X1 U56173 ( .A1(n55569), .A2(n55567), .B(n55568), .ZN(n55523) );
  NOR2_X1 U56174 ( .A1(n55518), .A2(n55597), .ZN(n55520) );
  NOR2_X1 U56175 ( .A1(n55592), .A2(n55575), .ZN(n55519) );
  OAI21_X1 U56176 ( .A1(n55521), .A2(n55520), .B(n55519), .ZN(n55522) );
  OAI21_X1 U56177 ( .A1(n55524), .A2(n55523), .B(n55522), .ZN(n55533) );
  OAI21_X1 U56178 ( .A1(n55569), .A2(n55575), .B(n55592), .ZN(n55526) );
  OAI22_X1 U56179 ( .A1(n55574), .A2(n55597), .B1(n55587), .B2(n1592), .ZN(
        n55525) );
  NAND3_X1 U56180 ( .A1(n55556), .A2(n4801), .A3(n55569), .ZN(n55529) );
  NOR2_X1 U56181 ( .A1(n55550), .A2(n55569), .ZN(n55527) );
  AOI22_X1 U56182 ( .A1(n55527), .A2(n55597), .B1(n55567), .B2(n55575), .ZN(
        n55528) );
  OAI21_X1 U56183 ( .A1(n55530), .A2(n55529), .B(n55528), .ZN(n55531) );
  INV_X1 U56186 ( .I(n55570), .ZN(n55537) );
  OAI21_X1 U56187 ( .A1(n55566), .A2(n55585), .B(n55537), .ZN(n55545) );
  INV_X1 U56188 ( .I(n55568), .ZN(n55540) );
  INV_X1 U56189 ( .I(n55571), .ZN(n55588) );
  AOI22_X1 U56190 ( .A1(n55540), .A2(n55539), .B1(n55588), .B2(n55538), .ZN(
        n55544) );
  NAND2_X1 U56191 ( .A1(n55586), .A2(n55571), .ZN(n55542) );
  NAND3_X1 U56192 ( .A1(n55590), .A2(n55582), .A3(n55597), .ZN(n55541) );
  NAND3_X1 U56193 ( .A1(n55542), .A2(n55596), .A3(n55541), .ZN(n55543) );
  OAI22_X1 U56194 ( .A1(n55598), .A2(n55573), .B1(n55575), .B2(n55547), .ZN(
        n55548) );
  NAND2_X1 U56195 ( .A1(n55548), .A2(n4801), .ZN(n55554) );
  AOI21_X1 U56196 ( .A1(n15933), .A2(n55574), .B(n55549), .ZN(n55553) );
  NAND3_X1 U56197 ( .A1(n55590), .A2(n55569), .A3(n21273), .ZN(n55555) );
  NAND2_X1 U56198 ( .A1(n55595), .A2(n55565), .ZN(n55551) );
  NAND3_X1 U56199 ( .A1(n55551), .A2(n55573), .A3(n55550), .ZN(n55552) );
  NAND4_X1 U56200 ( .A1(n55554), .A2(n55553), .A3(n55555), .A4(n55552), .ZN(
        n55561) );
  INV_X1 U56201 ( .I(n55555), .ZN(n55559) );
  AOI21_X1 U56202 ( .A1(n19183), .A2(n55590), .B(n55592), .ZN(n55558) );
  NOR2_X1 U56203 ( .A1(n55556), .A2(n55565), .ZN(n55557) );
  AOI22_X1 U56204 ( .A1(n55568), .A2(n55559), .B1(n55558), .B2(n55557), .ZN(
        n55560) );
  NAND2_X1 U56205 ( .A1(n55561), .A2(n55560), .ZN(n55562) );
  XOR2_X1 U56206 ( .A1(n55562), .A2(n24057), .Z(Plaintext[117]) );
  NOR2_X1 U56207 ( .A1(n55590), .A2(n55595), .ZN(n55564) );
  NAND2_X1 U56208 ( .A1(n55587), .A2(n55598), .ZN(n55563) );
  AOI22_X1 U56209 ( .A1(n55566), .A2(n55565), .B1(n55564), .B2(n55563), .ZN(
        n55579) );
  NAND2_X1 U56210 ( .A1(n55572), .A2(n55571), .ZN(n55578) );
  INV_X1 U56211 ( .I(n55573), .ZN(n55576) );
  NAND4_X1 U56212 ( .A1(n55576), .A2(n55575), .A3(n55574), .A4(n4801), .ZN(
        n55577) );
  XOR2_X1 U56213 ( .A1(n55581), .A2(n55580), .Z(Plaintext[118]) );
  NOR2_X1 U56214 ( .A1(n1592), .A2(n21272), .ZN(n55591) );
  NAND2_X1 U56215 ( .A1(n55591), .A2(n55597), .ZN(n55583) );
  OAI21_X1 U56216 ( .A1(n19183), .A2(n55587), .B(n55586), .ZN(n55589) );
  NAND2_X1 U56217 ( .A1(n55589), .A2(n55588), .ZN(n55602) );
  AOI22_X1 U56218 ( .A1(n55593), .A2(n55592), .B1(n55591), .B2(n55590), .ZN(
        n55601) );
  OAI21_X1 U56219 ( .A1(n55625), .A2(n55611), .B(n55640), .ZN(n55609) );
  NAND3_X1 U56220 ( .A1(n55607), .A2(n55651), .A3(n55619), .ZN(n55608) );
  NAND2_X1 U56222 ( .A1(n55613), .A2(n58701), .ZN(n55616) );
  NAND2_X1 U56224 ( .A1(n55631), .A2(n63520), .ZN(n55614) );
  NAND4_X1 U56225 ( .A1(n55616), .A2(n55644), .A3(n55615), .A4(n55614), .ZN(
        n55622) );
  NOR2_X1 U56226 ( .A1(n55643), .A2(n19021), .ZN(n55618) );
  NAND3_X1 U56228 ( .A1(n55632), .A2(n55651), .A3(n19020), .ZN(n55620) );
  AOI21_X1 U56229 ( .A1(n55628), .A2(n55627), .B(n55631), .ZN(n55629) );
  INV_X1 U56230 ( .I(n55649), .ZN(n55635) );
  NAND3_X1 U56231 ( .A1(n55630), .A2(n19020), .A3(n55643), .ZN(n55634) );
  NAND4_X1 U56232 ( .A1(n55632), .A2(n19020), .A3(n55651), .A4(n55631), .ZN(
        n55633) );
  NAND4_X1 U56235 ( .A1(n55645), .A2(n19021), .A3(n55644), .A4(n55643), .ZN(
        n55646) );
  NAND2_X1 U56236 ( .A1(n55649), .A2(n19021), .ZN(n55653) );
  NAND2_X1 U56237 ( .A1(n55926), .A2(n3616), .ZN(n55657) );
  NAND2_X1 U56238 ( .A1(n55661), .A2(n55660), .ZN(n55662) );
  INV_X1 U56239 ( .I(n55926), .ZN(n55664) );
  NAND3_X1 U56240 ( .A1(n55969), .A2(n55674), .A3(n55673), .ZN(n55675) );
  NOR2_X1 U56242 ( .A1(n55677), .A2(n15730), .ZN(n55678) );
  NOR2_X1 U56243 ( .A1(n55694), .A2(n55695), .ZN(n55688) );
  NAND2_X1 U56244 ( .A1(n55686), .A2(n55685), .ZN(n55687) );
  OAI21_X1 U56245 ( .A1(n55689), .A2(n55688), .B(n55687), .ZN(n55702) );
  NOR2_X1 U56246 ( .A1(n59040), .A2(n55695), .ZN(n55693) );
  NAND2_X1 U56247 ( .A1(n52044), .A2(n20849), .ZN(n55697) );
  NAND2_X1 U56248 ( .A1(n55697), .A2(n55696), .ZN(n55698) );
  NAND3_X1 U56249 ( .A1(n24472), .A2(n56229), .A3(n61213), .ZN(n55705) );
  NAND2_X1 U56250 ( .A1(n55706), .A2(n55705), .ZN(n55707) );
  NAND2_X1 U56251 ( .A1(n56225), .A2(n55982), .ZN(n55710) );
  AOI21_X1 U56252 ( .A1(n55710), .A2(n56434), .B(n61368), .ZN(n55711) );
  OAI21_X1 U56253 ( .A1(n55714), .A2(n1369), .B(n55713), .ZN(n55715) );
  INV_X1 U56255 ( .I(n55724), .ZN(n55725) );
  NAND3_X1 U56256 ( .A1(n55726), .A2(n55725), .A3(n55740), .ZN(n55732) );
  AOI21_X1 U56257 ( .A1(n57901), .A2(n55728), .B(n55727), .ZN(n55729) );
  NAND2_X1 U56258 ( .A1(n55730), .A2(n55729), .ZN(n55731) );
  OAI21_X1 U56259 ( .A1(n55737), .A2(n6531), .B(n55735), .ZN(n55744) );
  NAND2_X1 U56260 ( .A1(n55741), .A2(n55740), .ZN(n55742) );
  AOI21_X1 U56261 ( .A1(n55816), .A2(n55831), .B(n55811), .ZN(n55749) );
  OAI22_X1 U56263 ( .A1(n55747), .A2(n14890), .B1(n55800), .B2(n55757), .ZN(
        n55748) );
  NAND3_X1 U56265 ( .A1(n55750), .A2(n22860), .A3(n21403), .ZN(n55754) );
  NAND2_X1 U56266 ( .A1(n55784), .A2(n55759), .ZN(n55751) );
  NAND3_X1 U56267 ( .A1(n55751), .A2(n55752), .A3(n55820), .ZN(n55753) );
  NAND3_X1 U56268 ( .A1(n55820), .A2(n55752), .A3(n55802), .ZN(n55758) );
  NAND2_X1 U56269 ( .A1(n55812), .A2(n55759), .ZN(n55756) );
  AOI21_X1 U56270 ( .A1(n55793), .A2(n55758), .B(n22860), .ZN(n55763) );
  NAND2_X1 U56271 ( .A1(n24958), .A2(n55821), .ZN(n55788) );
  NAND3_X1 U56272 ( .A1(n55812), .A2(n60855), .A3(n55828), .ZN(n55761) );
  XOR2_X1 U56273 ( .A1(n55767), .A2(n55766), .Z(Plaintext[127]) );
  NOR2_X1 U56274 ( .A1(n55827), .A2(n55820), .ZN(n55776) );
  INV_X1 U56275 ( .I(n55802), .ZN(n55771) );
  AOI21_X1 U56276 ( .A1(n55817), .A2(n55796), .B(n55771), .ZN(n55775) );
  OAI22_X1 U56277 ( .A1(n55773), .A2(n55826), .B1(n55795), .B2(n55820), .ZN(
        n55774) );
  NOR3_X1 U56278 ( .A1(n55776), .A2(n55775), .A3(n55774), .ZN(n55779) );
  XOR2_X1 U56279 ( .A1(n55779), .A2(n55778), .Z(Plaintext[128]) );
  NAND2_X1 U56280 ( .A1(n55811), .A2(n55781), .ZN(n55782) );
  OAI21_X1 U56281 ( .A1(n55783), .A2(n55782), .B(n60855), .ZN(n55791) );
  OAI21_X1 U56282 ( .A1(n55793), .A2(n55828), .B(n55784), .ZN(n55790) );
  INV_X1 U56284 ( .I(n55793), .ZN(n55799) );
  INV_X1 U56286 ( .I(n55796), .ZN(n55797) );
  OAI21_X1 U56287 ( .A1(n55802), .A2(n55801), .B(n55800), .ZN(n55807) );
  INV_X1 U56288 ( .I(n55811), .ZN(n55805) );
  AOI21_X1 U56289 ( .A1(n55805), .A2(n55820), .B(n55804), .ZN(n55806) );
  NAND2_X1 U56291 ( .A1(n55817), .A2(n22860), .ZN(n55832) );
  OAI21_X1 U56292 ( .A1(n55822), .A2(n55820), .B(n55819), .ZN(n55825) );
  OAI21_X1 U56294 ( .A1(n55881), .A2(n55835), .B(n15716), .ZN(n55839) );
  NOR2_X1 U56296 ( .A1(n55891), .A2(n55842), .ZN(n55836) );
  NOR2_X1 U56297 ( .A1(n55896), .A2(n55854), .ZN(n55852) );
  NAND4_X1 U56300 ( .A1(n55842), .A2(n60203), .A3(n15716), .A4(n55893), .ZN(
        n55844) );
  NOR2_X1 U56304 ( .A1(n55898), .A2(n22681), .ZN(n55853) );
  AOI22_X1 U56305 ( .A1(n55853), .A2(n55899), .B1(n55852), .B2(n55893), .ZN(
        n55859) );
  NAND2_X1 U56307 ( .A1(n55867), .A2(n55856), .ZN(n55857) );
  NAND4_X1 U56308 ( .A1(n55857), .A2(n17774), .A3(n55871), .A4(n55879), .ZN(
        n55858) );
  XOR2_X1 U56310 ( .A1(n55863), .A2(n55862), .Z(Plaintext[133]) );
  NAND3_X1 U56311 ( .A1(n18561), .A2(n60092), .A3(n55871), .ZN(n55866) );
  NAND2_X1 U56312 ( .A1(n55864), .A2(n60092), .ZN(n55865) );
  NAND3_X1 U56313 ( .A1(n55866), .A2(n55898), .A3(n55865), .ZN(n55875) );
  OAI21_X1 U56314 ( .A1(n55887), .A2(n11782), .B(n55900), .ZN(n55874) );
  NAND2_X1 U56315 ( .A1(n60092), .A2(n22681), .ZN(n55869) );
  NAND3_X1 U56316 ( .A1(n55871), .A2(n55870), .A3(n55869), .ZN(n55872) );
  NAND2_X1 U56317 ( .A1(n55872), .A2(n55899), .ZN(n55873) );
  NAND3_X1 U56318 ( .A1(n55875), .A2(n55874), .A3(n55873), .ZN(n55877) );
  XOR2_X1 U56319 ( .A1(n55877), .A2(n55876), .Z(Plaintext[134]) );
  NOR2_X1 U56320 ( .A1(n55885), .A2(n15716), .ZN(n55890) );
  NAND3_X1 U56321 ( .A1(n55886), .A2(n55890), .A3(n17774), .ZN(n55888) );
  NOR2_X1 U56322 ( .A1(n55891), .A2(n55890), .ZN(n55902) );
  NAND2_X1 U56323 ( .A1(n17774), .A2(n13858), .ZN(n55894) );
  XOR2_X1 U56324 ( .A1(n55904), .A2(n55903), .Z(Plaintext[137]) );
  OAI22_X1 U56326 ( .A1(n55910), .A2(n13025), .B1(n23360), .B2(n55908), .ZN(
        n55913) );
  NOR2_X1 U56327 ( .A1(n13025), .A2(n1324), .ZN(n55917) );
  OAI21_X1 U56328 ( .A1(n55917), .A2(n55916), .B(n55915), .ZN(n55918) );
  AOI21_X1 U56329 ( .A1(n56273), .A2(n55921), .B(n55920), .ZN(n55923) );
  NOR3_X1 U56331 ( .A1(n56264), .A2(n22817), .A3(n55931), .ZN(n55932) );
  NAND2_X1 U56333 ( .A1(n56396), .A2(n55935), .ZN(n55940) );
  NAND2_X1 U56334 ( .A1(n55937), .A2(n55936), .ZN(n55938) );
  INV_X1 U56335 ( .I(n56389), .ZN(n55941) );
  NAND2_X1 U56337 ( .A1(n56389), .A2(n56563), .ZN(n55942) );
  INV_X2 U56341 ( .I(n56092), .ZN(n56045) );
  MUX2_X1 U56342 ( .I0(n56255), .I1(n56254), .S(n65175), .Z(n55948) );
  INV_X1 U56343 ( .I(n56404), .ZN(n56409) );
  INV_X1 U56345 ( .I(n55952), .ZN(n55949) );
  OAI21_X1 U56346 ( .A1(n7274), .A2(n55949), .B(n56579), .ZN(n55955) );
  NAND2_X1 U56347 ( .A1(n56593), .A2(n57691), .ZN(n55953) );
  NAND2_X1 U56348 ( .A1(n23952), .A2(n21957), .ZN(n55951) );
  OAI21_X1 U56351 ( .A1(n55957), .A2(n55956), .B(n56580), .ZN(n55961) );
  INV_X1 U56352 ( .I(n56256), .ZN(n55958) );
  NOR2_X1 U56354 ( .A1(n56035), .A2(n9568), .ZN(n55996) );
  NOR2_X2 U56355 ( .A1(n56047), .A2(n56071), .ZN(n56105) );
  NOR2_X1 U56357 ( .A1(n56227), .A2(n56229), .ZN(n55984) );
  NOR2_X1 U56358 ( .A1(n55985), .A2(n55984), .ZN(n55992) );
  NOR2_X1 U56359 ( .A1(n55988), .A2(n55987), .ZN(n55989) );
  NOR2_X1 U56360 ( .A1(n56080), .A2(n9567), .ZN(n55995) );
  NAND2_X1 U56361 ( .A1(n56071), .A2(n56084), .ZN(n56010) );
  NOR2_X1 U56362 ( .A1(n56108), .A2(n56010), .ZN(n55999) );
  AOI21_X1 U56364 ( .A1(n56071), .A2(n24092), .B(n56009), .ZN(n55998) );
  NOR2_X1 U56366 ( .A1(n56120), .A2(n56092), .ZN(n56001) );
  NOR2_X1 U56368 ( .A1(n24092), .A2(n56071), .ZN(n56002) );
  OAI21_X1 U56370 ( .A1(n56045), .A2(n56010), .B(n56009), .ZN(n56011) );
  OAI21_X1 U56371 ( .A1(n56100), .A2(n24092), .B(n56011), .ZN(n56029) );
  NAND2_X1 U56372 ( .A1(n56047), .A2(n56045), .ZN(n56063) );
  INV_X1 U56373 ( .I(n56063), .ZN(n56017) );
  NAND2_X1 U56375 ( .A1(n63012), .A2(n56106), .ZN(n56020) );
  NAND2_X1 U56378 ( .A1(n56013), .A2(n56012), .ZN(n56015) );
  INV_X1 U56381 ( .I(n56018), .ZN(n56019) );
  NAND3_X1 U56382 ( .A1(n56105), .A2(n56035), .A3(n56019), .ZN(n56027) );
  NOR2_X1 U56383 ( .A1(n56020), .A2(n63023), .ZN(n56023) );
  INV_X1 U56386 ( .I(n56115), .ZN(n56031) );
  AOI21_X1 U56387 ( .A1(n56082), .A2(n56080), .B(n56031), .ZN(n56033) );
  NOR3_X1 U56388 ( .A1(n56033), .A2(n56120), .A3(n56032), .ZN(n56039) );
  NAND2_X1 U56389 ( .A1(n56047), .A2(n56071), .ZN(n56034) );
  NAND2_X1 U56390 ( .A1(n24092), .A2(n61740), .ZN(n56067) );
  NAND3_X1 U56391 ( .A1(n56034), .A2(n56117), .A3(n56067), .ZN(n56038) );
  INV_X1 U56392 ( .I(n56035), .ZN(n56036) );
  NAND3_X1 U56393 ( .A1(n56036), .A2(n56105), .A3(n9567), .ZN(n56037) );
  NAND3_X1 U56394 ( .A1(n56039), .A2(n56038), .A3(n56037), .ZN(n56041) );
  XOR2_X1 U56395 ( .A1(n56041), .A2(n56040), .Z(Plaintext[140]) );
  NOR2_X1 U56396 ( .A1(n56042), .A2(n60672), .ZN(n56044) );
  NOR3_X1 U56397 ( .A1(n56072), .A2(n63699), .A3(n56088), .ZN(n56043) );
  AOI21_X1 U56398 ( .A1(n56044), .A2(n56063), .B(n56043), .ZN(n56057) );
  NAND2_X1 U56399 ( .A1(n56120), .A2(n56045), .ZN(n56062) );
  INV_X1 U56400 ( .I(n56062), .ZN(n56046) );
  NAND2_X1 U56401 ( .A1(n56046), .A2(n60672), .ZN(n56056) );
  NOR2_X1 U56402 ( .A1(n56047), .A2(n24092), .ZN(n56090) );
  INV_X1 U56403 ( .I(n56048), .ZN(n56049) );
  INV_X1 U56404 ( .I(n56089), .ZN(n56051) );
  NAND2_X1 U56405 ( .A1(n56051), .A2(n56065), .ZN(n56052) );
  OAI21_X1 U56407 ( .A1(n56081), .A2(n56106), .B(n56067), .ZN(n56053) );
  NAND3_X1 U56408 ( .A1(n56053), .A2(n63699), .A3(n56072), .ZN(n56054) );
  NAND2_X1 U56410 ( .A1(n60672), .A2(n1897), .ZN(n56061) );
  NOR2_X1 U56411 ( .A1(n56088), .A2(n56061), .ZN(n56059) );
  NAND2_X1 U56412 ( .A1(n56064), .A2(n56063), .ZN(n56068) );
  NOR2_X1 U56413 ( .A1(n60672), .A2(n56065), .ZN(n56070) );
  INV_X1 U56414 ( .I(n56070), .ZN(n56066) );
  AOI21_X1 U56415 ( .A1(n56068), .A2(n56067), .B(n56066), .ZN(n56076) );
  NAND3_X1 U56416 ( .A1(n56069), .A2(n56090), .A3(n1897), .ZN(n56074) );
  NAND4_X1 U56418 ( .A1(n64875), .A2(n56072), .A3(n56071), .A4(n56070), .ZN(
        n56073) );
  NAND2_X1 U56419 ( .A1(n56074), .A2(n56073), .ZN(n56075) );
  NOR3_X1 U56420 ( .A1(n56077), .A2(n56076), .A3(n56075), .ZN(n56078) );
  NOR2_X1 U56421 ( .A1(n56082), .A2(n56108), .ZN(n56083) );
  NOR2_X1 U56422 ( .A1(n56102), .A2(n56083), .ZN(n56096) );
  INV_X1 U56424 ( .I(n56091), .ZN(n56087) );
  OAI21_X1 U56425 ( .A1(n56115), .A2(n56087), .B(n64875), .ZN(n56095) );
  NAND3_X1 U56427 ( .A1(n56105), .A2(n63023), .A3(n56091), .ZN(n56093) );
  XOR2_X1 U56429 ( .A1(n56098), .A2(n57989), .Z(Plaintext[142]) );
  NOR2_X1 U56430 ( .A1(n56099), .A2(n61740), .ZN(n56101) );
  NAND4_X1 U56433 ( .A1(n56117), .A2(n56108), .A3(n61740), .A4(n56106), .ZN(
        n56112) );
  NOR2_X1 U56436 ( .A1(n9568), .A2(n56115), .ZN(n56119) );
  INV_X1 U56437 ( .I(n56117), .ZN(n56118) );
  XOR2_X1 U56438 ( .A1(n56126), .A2(n56125), .Z(Plaintext[143]) );
  OAI21_X1 U56439 ( .A1(n56128), .A2(n56127), .B(n5172), .ZN(n56132) );
  OAI21_X1 U56440 ( .A1(n56132), .A2(n56150), .B(n56131), .ZN(n56137) );
  XOR2_X1 U56441 ( .A1(n56182), .A2(n56146), .Z(n56133) );
  NAND2_X1 U56442 ( .A1(n56171), .A2(n61228), .ZN(n56134) );
  NAND2_X1 U56443 ( .A1(n56174), .A2(n56191), .ZN(n56138) );
  NAND2_X1 U56444 ( .A1(n56138), .A2(n56185), .ZN(n56166) );
  NAND3_X1 U56445 ( .A1(n19853), .A2(n56150), .A3(n56166), .ZN(n56141) );
  NAND3_X1 U56446 ( .A1(n56158), .A2(n23258), .A3(n56196), .ZN(n56139) );
  NAND4_X1 U56448 ( .A1(n56149), .A2(n19853), .A3(n61228), .A4(n56184), .ZN(
        n56154) );
  INV_X1 U56451 ( .I(n56150), .ZN(n56151) );
  NAND2_X1 U56452 ( .A1(n56152), .A2(n56151), .ZN(n56153) );
  NAND2_X1 U56454 ( .A1(n56171), .A2(n64438), .ZN(n56161) );
  NAND3_X1 U56455 ( .A1(n56188), .A2(n56162), .A3(n56161), .ZN(n56164) );
  NAND3_X1 U56456 ( .A1(n56192), .A2(n23258), .A3(n56171), .ZN(n56163) );
  NAND3_X1 U56457 ( .A1(n56188), .A2(n64438), .A3(n56166), .ZN(n56179) );
  INV_X1 U56458 ( .I(n56168), .ZN(n56170) );
  NAND2_X1 U56459 ( .A1(n56185), .A2(n56174), .ZN(n56175) );
  XOR2_X1 U56460 ( .A1(n56181), .A2(n56180), .Z(Plaintext[147]) );
  NAND2_X1 U56461 ( .A1(n56191), .A2(n11716), .ZN(n56194) );
  NAND3_X1 U56462 ( .A1(n23258), .A2(n56194), .A3(n61228), .ZN(n56183) );
  OAI21_X1 U56463 ( .A1(n56186), .A2(n56185), .B(n56184), .ZN(n56187) );
  NAND2_X1 U56464 ( .A1(n56188), .A2(n56187), .ZN(n56200) );
  XOR2_X1 U56466 ( .A1(n56203), .A2(n56202), .Z(Plaintext[149]) );
  NOR2_X1 U56467 ( .A1(n56204), .A2(n56417), .ZN(n56208) );
  INV_X1 U56468 ( .I(n56205), .ZN(n56620) );
  OAI22_X1 U56469 ( .A1(n56620), .A2(n56217), .B1(n58846), .B2(n56214), .ZN(
        n56207) );
  NOR2_X1 U56471 ( .A1(n1598), .A2(n56420), .ZN(n56221) );
  NOR2_X1 U56472 ( .A1(n56221), .A2(n56220), .ZN(n56222) );
  NAND3_X1 U56473 ( .A1(n56231), .A2(n62263), .A3(n56230), .ZN(n56232) );
  OAI21_X1 U56474 ( .A1(n56234), .A2(n56554), .B(n56233), .ZN(n56235) );
  NAND2_X1 U56475 ( .A1(n57239), .A2(n60809), .ZN(n56243) );
  INV_X1 U56476 ( .I(n56359), .ZN(n56240) );
  OAI21_X1 U56477 ( .A1(n56407), .A2(n56248), .B(n56408), .ZN(n56247) );
  NAND3_X1 U56478 ( .A1(n22473), .A2(n56245), .A3(n61554), .ZN(n56246) );
  NAND2_X1 U56479 ( .A1(n56247), .A2(n56246), .ZN(n56252) );
  INV_X1 U56481 ( .I(n56579), .ZN(n56253) );
  INV_X1 U56482 ( .I(n56590), .ZN(n56259) );
  NAND2_X1 U56483 ( .A1(n56257), .A2(n56412), .ZN(n56258) );
  INV_X1 U56484 ( .I(n56267), .ZN(n56272) );
  NOR2_X1 U56485 ( .A1(n56269), .A2(n56268), .ZN(n56270) );
  AOI21_X1 U56487 ( .A1(n24032), .A2(n56328), .B(n56347), .ZN(n56284) );
  OAI21_X1 U56488 ( .A1(n56284), .A2(n56296), .B(n56283), .ZN(n56288) );
  NAND2_X1 U56489 ( .A1(n1591), .A2(n56351), .ZN(n56285) );
  OAI21_X1 U56490 ( .A1(n56293), .A2(n23318), .B(n56351), .ZN(n56286) );
  XOR2_X1 U56491 ( .A1(n56289), .A2(n24014), .Z(Plaintext[150]) );
  INV_X1 U56492 ( .I(n56347), .ZN(n56298) );
  NOR2_X1 U56493 ( .A1(n59180), .A2(n12058), .ZN(n56295) );
  AOI22_X1 U56494 ( .A1(n56298), .A2(n56320), .B1(n56297), .B2(n56296), .ZN(
        n56307) );
  NOR2_X1 U56495 ( .A1(n22891), .A2(n1591), .ZN(n56326) );
  NAND3_X1 U56496 ( .A1(n56313), .A2(n61627), .A3(n23318), .ZN(n56299) );
  NOR2_X1 U56497 ( .A1(n24032), .A2(n56299), .ZN(n56302) );
  AOI21_X1 U56499 ( .A1(n56326), .A2(n56302), .B(n56301), .ZN(n56306) );
  NAND2_X1 U56500 ( .A1(n20957), .A2(n59180), .ZN(n56303) );
  NAND4_X1 U56501 ( .A1(n61727), .A2(n24032), .A3(n56304), .A4(n56303), .ZN(
        n56305) );
  INV_X1 U56504 ( .I(n56328), .ZN(n56312) );
  INV_X1 U56505 ( .I(n56318), .ZN(n56315) );
  NAND3_X1 U56506 ( .A1(n56315), .A2(n56350), .A3(n20957), .ZN(n56316) );
  XOR2_X1 U56507 ( .A1(n56317), .A2(n24011), .Z(Plaintext[152]) );
  NOR2_X1 U56508 ( .A1(n20957), .A2(n22430), .ZN(n56321) );
  NAND3_X1 U56509 ( .A1(n56324), .A2(n22430), .A3(n56330), .ZN(n56334) );
  NOR2_X1 U56510 ( .A1(n1580), .A2(n24032), .ZN(n56325) );
  NAND2_X1 U56511 ( .A1(n56328), .A2(n56327), .ZN(n56329) );
  NAND2_X1 U56512 ( .A1(n56330), .A2(n56329), .ZN(n56332) );
  AOI21_X1 U56513 ( .A1(n56342), .A2(n58755), .B(n23318), .ZN(n56348) );
  AOI22_X1 U56514 ( .A1(n56348), .A2(n56347), .B1(n56346), .B2(n24032), .ZN(
        n56357) );
  INV_X1 U56515 ( .I(n56351), .ZN(n56353) );
  NAND3_X1 U56516 ( .A1(n61727), .A2(n56353), .A3(n20957), .ZN(n56355) );
  NAND2_X1 U56520 ( .A1(n56534), .A2(n22229), .ZN(n56385) );
  OAI21_X1 U56521 ( .A1(n56385), .A2(n56381), .B(n56384), .ZN(n56388) );
  OAI22_X1 U56524 ( .A1(n51264), .A2(n56565), .B1(n56572), .B2(n56568), .ZN(
        n56392) );
  INV_X1 U56526 ( .I(n56402), .ZN(n56405) );
  NAND2_X1 U56529 ( .A1(n56425), .A2(n56424), .ZN(n56426) );
  AOI21_X1 U56530 ( .A1(n56428), .A2(n62261), .B(n56426), .ZN(n56443) );
  INV_X1 U56531 ( .I(n56430), .ZN(n56431) );
  AOI21_X1 U56532 ( .A1(n1616), .A2(n24473), .B(n64808), .ZN(n56438) );
  NAND2_X1 U56534 ( .A1(n20587), .A2(n56502), .ZN(n56445) );
  NAND2_X1 U56535 ( .A1(n56453), .A2(n56502), .ZN(n56444) );
  NAND2_X1 U56538 ( .A1(n26162), .A2(n19999), .ZN(n56446) );
  AOI21_X1 U56548 ( .A1(n15238), .A2(n56489), .B(n56510), .ZN(n56461) );
  NOR2_X1 U56549 ( .A1(n56463), .A2(n20587), .ZN(n56464) );
  INV_X1 U56550 ( .I(n56466), .ZN(n56467) );
  NOR2_X1 U56554 ( .A1(n56473), .A2(n23920), .ZN(n56472) );
  NAND3_X1 U56555 ( .A1(n15238), .A2(n56473), .A3(n10286), .ZN(n56474) );
  INV_X1 U56557 ( .I(n26162), .ZN(n56491) );
  NOR2_X1 U56558 ( .A1(n24551), .A2(n56489), .ZN(n56490) );
  AOI22_X1 U56559 ( .A1(n56491), .A2(n56490), .B1(n56523), .B2(n15765), .ZN(
        n56494) );
  NAND2_X1 U56560 ( .A1(n56492), .A2(n56496), .ZN(n56493) );
  NAND2_X1 U56561 ( .A1(n56502), .A2(n19999), .ZN(n56497) );
  INV_X1 U56562 ( .I(n56498), .ZN(n56501) );
  NOR2_X1 U56563 ( .A1(n65216), .A2(n20587), .ZN(n56521) );
  NOR2_X1 U56564 ( .A1(n56499), .A2(n1366), .ZN(n56500) );
  AOI22_X1 U56565 ( .A1(n56501), .A2(n56521), .B1(n20587), .B2(n56500), .ZN(
        n56507) );
  INV_X1 U56568 ( .I(n56505), .ZN(n56506) );
  NOR2_X1 U56570 ( .A1(n26162), .A2(n9311), .ZN(n56514) );
  NAND2_X1 U56572 ( .A1(n20587), .A2(n10286), .ZN(n56518) );
  AOI21_X1 U56573 ( .A1(n15765), .A2(n56518), .B(n56517), .ZN(n56519) );
  NOR2_X1 U56575 ( .A1(n23920), .A2(n19999), .ZN(n56524) );
  OAI21_X1 U56576 ( .A1(n15765), .A2(n56524), .B(n56523), .ZN(n56525) );
  NAND3_X1 U56580 ( .A1(n56531), .A2(n56530), .A3(n56381), .ZN(n56536) );
  OAI21_X1 U56583 ( .A1(n56543), .A2(n1153), .B(n57012), .ZN(n56550) );
  NAND2_X1 U56585 ( .A1(n56555), .A2(n15875), .ZN(n56556) );
  NAND2_X1 U56587 ( .A1(n56572), .A2(n11121), .ZN(n56566) );
  NOR2_X1 U56592 ( .A1(n56586), .A2(n57691), .ZN(n56588) );
  OAI21_X1 U56594 ( .A1(n19151), .A2(n56978), .B(n56598), .ZN(n56602) );
  INV_X1 U56597 ( .I(n56985), .ZN(n56609) );
  OAI21_X1 U56598 ( .A1(n56993), .A2(n56609), .B(n7835), .ZN(n56611) );
  NAND3_X1 U56602 ( .A1(n56716), .A2(n56719), .A3(n56697), .ZN(n56647) );
  INV_X1 U56606 ( .I(n56623), .ZN(n56628) );
  OAI21_X1 U56607 ( .A1(n60129), .A2(n56632), .B(n59449), .ZN(n56626) );
  NAND3_X1 U56608 ( .A1(n56628), .A2(n56627), .A3(n56626), .ZN(n56642) );
  NOR2_X1 U56609 ( .A1(n56629), .A2(n56635), .ZN(n56634) );
  OAI21_X1 U56610 ( .A1(n56632), .A2(n58846), .B(n56630), .ZN(n56633) );
  AOI22_X1 U56611 ( .A1(n56636), .A2(n56635), .B1(n56634), .B2(n56633), .ZN(
        n56641) );
  AOI21_X1 U56612 ( .A1(n56639), .A2(n56638), .B(n56637), .ZN(n56640) );
  NAND3_X1 U56613 ( .A1(n56645), .A2(n56703), .A3(n56719), .ZN(n56646) );
  NAND3_X1 U56616 ( .A1(n56732), .A2(n56697), .A3(n56731), .ZN(n56654) );
  NAND2_X1 U56617 ( .A1(n56677), .A2(n56703), .ZN(n56652) );
  NAND2_X1 U56621 ( .A1(n56658), .A2(n59461), .ZN(n56664) );
  NAND3_X1 U56622 ( .A1(n56661), .A2(n56660), .A3(n59461), .ZN(n56662) );
  NAND3_X1 U56623 ( .A1(n56664), .A2(n56663), .A3(n56662), .ZN(n56665) );
  NOR2_X1 U56624 ( .A1(n56666), .A2(n56665), .ZN(n56669) );
  NAND2_X1 U56625 ( .A1(n56669), .A2(n56717), .ZN(n56724) );
  NOR2_X1 U56626 ( .A1(n56724), .A2(n20269), .ZN(n56668) );
  OAI21_X1 U56627 ( .A1(n56668), .A2(n56667), .B(n56719), .ZN(n56672) );
  INV_X1 U56628 ( .I(n56669), .ZN(n56670) );
  INV_X1 U56629 ( .I(n56724), .ZN(n56673) );
  NOR2_X1 U56630 ( .A1(n56708), .A2(n56731), .ZN(n56676) );
  NOR2_X1 U56632 ( .A1(n20269), .A2(n56722), .ZN(n56678) );
  XOR2_X1 U56636 ( .A1(n56685), .A2(n56684), .Z(Plaintext[163]) );
  NAND2_X1 U56637 ( .A1(n20269), .A2(n56697), .ZN(n56723) );
  OAI21_X1 U56638 ( .A1(n56707), .A2(n56723), .B(n56703), .ZN(n56686) );
  NOR2_X1 U56639 ( .A1(n56696), .A2(n56686), .ZN(n56691) );
  NAND2_X1 U56640 ( .A1(n20269), .A2(n56731), .ZN(n56736) );
  XOR2_X1 U56641 ( .A1(n56694), .A2(n56693), .Z(Plaintext[164]) );
  NOR3_X1 U56642 ( .A1(n56734), .A2(n56697), .A3(n56644), .ZN(n56698) );
  INV_X1 U56643 ( .I(n56738), .ZN(n56706) );
  NOR2_X1 U56644 ( .A1(n56704), .A2(n56703), .ZN(n56705) );
  NOR2_X1 U56647 ( .A1(n56734), .A2(n56731), .ZN(n56729) );
  NAND4_X1 U56648 ( .A1(n56716), .A2(n56725), .A3(n56722), .A4(n56729), .ZN(
        n56710) );
  INV_X1 U56650 ( .I(n56716), .ZN(n56721) );
  NAND2_X1 U56653 ( .A1(n56734), .A2(n56722), .ZN(n56737) );
  OAI22_X1 U56654 ( .A1(n56725), .A2(n56737), .B1(n56724), .B2(n56723), .ZN(
        n56726) );
  NOR3_X1 U56655 ( .A1(n56728), .A2(n56727), .A3(n56726), .ZN(n56744) );
  AOI22_X1 U56656 ( .A1(n56732), .A2(n56731), .B1(n56730), .B2(n56729), .ZN(
        n56743) );
  NAND3_X1 U56657 ( .A1(n56735), .A2(n56734), .A3(n56733), .ZN(n56741) );
  INV_X1 U56658 ( .I(n56736), .ZN(n56740) );
  NAND2_X1 U56659 ( .A1(n56738), .A2(n56737), .ZN(n56739) );
  NAND3_X1 U56660 ( .A1(n56741), .A2(n56740), .A3(n56739), .ZN(n56742) );
  XOR2_X1 U56661 ( .A1(n56746), .A2(n56745), .Z(Plaintext[167]) );
  NAND3_X1 U56663 ( .A1(n56755), .A2(n23879), .A3(n56816), .ZN(n56754) );
  NAND3_X1 U56666 ( .A1(n56788), .A2(n56775), .A3(n56809), .ZN(n56752) );
  NAND3_X1 U56669 ( .A1(n7209), .A2(n56806), .A3(n56775), .ZN(n56758) );
  NAND3_X1 U56670 ( .A1(n56760), .A2(n56759), .A3(n56758), .ZN(n56761) );
  AOI21_X1 U56672 ( .A1(n56763), .A2(n56815), .B(n56814), .ZN(n56770) );
  NAND2_X1 U56673 ( .A1(n56804), .A2(n56795), .ZN(n56765) );
  AOI21_X1 U56674 ( .A1(n23030), .A2(n23879), .B(n56791), .ZN(n56764) );
  NAND2_X1 U56675 ( .A1(n56765), .A2(n56764), .ZN(n56769) );
  INV_X1 U56676 ( .I(n56786), .ZN(n56767) );
  OAI21_X1 U56677 ( .A1(n56797), .A2(n56767), .B(n56766), .ZN(n56768) );
  NAND3_X1 U56678 ( .A1(n56770), .A2(n56769), .A3(n56768), .ZN(n56772) );
  XOR2_X1 U56679 ( .A1(n56772), .A2(n56771), .Z(Plaintext[170]) );
  NAND2_X1 U56680 ( .A1(n56775), .A2(n56791), .ZN(n56793) );
  OAI21_X1 U56682 ( .A1(n61971), .A2(n56788), .B(n56791), .ZN(n56780) );
  INV_X1 U56685 ( .I(n56785), .ZN(n56789) );
  NAND3_X1 U56688 ( .A1(n56795), .A2(n23030), .A3(n56793), .ZN(n56799) );
  XOR2_X1 U56690 ( .A1(n56802), .A2(n24109), .Z(Plaintext[172]) );
  NOR2_X1 U56691 ( .A1(n56809), .A2(n56808), .ZN(n56810) );
  AOI22_X1 U56692 ( .A1(n61971), .A2(n56810), .B1(n56815), .B2(n56814), .ZN(
        n56818) );
  AOI21_X1 U56693 ( .A1(n22667), .A2(n56890), .B(n56853), .ZN(n56821) );
  NAND2_X1 U56695 ( .A1(n56821), .A2(n56820), .ZN(n56826) );
  NOR3_X1 U56696 ( .A1(n56881), .A2(n23074), .A3(n56838), .ZN(n56823) );
  NAND4_X1 U56697 ( .A1(n56885), .A2(n56844), .A3(n56881), .A4(n56867), .ZN(
        n56825) );
  NAND2_X1 U56699 ( .A1(n56830), .A2(n59827), .ZN(n56833) );
  NAND2_X1 U56700 ( .A1(n10507), .A2(n56834), .ZN(n56836) );
  INV_X1 U56702 ( .I(n56853), .ZN(n56866) );
  NOR2_X1 U56703 ( .A1(n23682), .A2(n64230), .ZN(n56855) );
  INV_X1 U56704 ( .I(n56862), .ZN(n56854) );
  OAI21_X1 U56705 ( .A1(n56866), .A2(n56855), .B(n56854), .ZN(n56858) );
  NAND2_X1 U56706 ( .A1(n56888), .A2(n56856), .ZN(n56857) );
  XOR2_X1 U56707 ( .A1(n56860), .A2(n56859), .Z(Plaintext[176]) );
  AOI21_X1 U56708 ( .A1(n64230), .A2(n56862), .B(n56861), .ZN(n56864) );
  NAND2_X1 U56710 ( .A1(n56868), .A2(n56867), .ZN(n56869) );
  INV_X1 U56711 ( .I(n56869), .ZN(n56871) );
  OAI21_X1 U56712 ( .A1(n56871), .A2(n56870), .B(n56885), .ZN(n56877) );
  INV_X1 U56713 ( .I(n56872), .ZN(n56875) );
  AOI21_X1 U56714 ( .A1(n56875), .A2(n56874), .B(n56873), .ZN(n56876) );
  INV_X1 U56715 ( .I(n56883), .ZN(n56884) );
  OAI21_X1 U56716 ( .A1(n56885), .A2(n23682), .B(n56884), .ZN(n56889) );
  AOI21_X1 U56719 ( .A1(n56895), .A2(n23682), .B(n56893), .ZN(n56896) );
  OAI21_X1 U56720 ( .A1(n59273), .A2(n64833), .B(n56896), .ZN(n56899) );
  NOR2_X1 U56722 ( .A1(n9655), .A2(n1583), .ZN(n56903) );
  NOR3_X1 U56723 ( .A1(n56906), .A2(n64845), .A3(n14708), .ZN(n56907) );
  INV_X1 U56724 ( .I(n56908), .ZN(n56910) );
  OAI21_X1 U56725 ( .A1(n56910), .A2(n56909), .B(n56957), .ZN(n56913) );
  NAND4_X1 U56726 ( .A1(n56916), .A2(n56958), .A3(n25987), .A4(n1583), .ZN(
        n56923) );
  NOR2_X1 U56727 ( .A1(n25988), .A2(n1257), .ZN(n56918) );
  NOR2_X1 U56728 ( .A1(n56953), .A2(n56961), .ZN(n56917) );
  NAND2_X1 U56732 ( .A1(n56953), .A2(n1583), .ZN(n56941) );
  NAND3_X1 U56733 ( .A1(n56941), .A2(n56940), .A3(n25987), .ZN(n56946) );
  INV_X1 U56734 ( .I(n56941), .ZN(n56943) );
  NAND3_X1 U56736 ( .A1(n56946), .A2(n56945), .A3(n56944), .ZN(n56947) );
  NOR3_X1 U56739 ( .A1(n25987), .A2(n14708), .A3(n1257), .ZN(n56954) );
  INV_X1 U56740 ( .I(n56957), .ZN(n56960) );
  INV_X1 U56741 ( .I(n56964), .ZN(n56971) );
  AOI22_X1 U56750 ( .A1(n1601), .A2(n15718), .B1(n23102), .B2(n57030), .ZN(
        n57020) );
  AOI21_X1 U56753 ( .A1(n23563), .A2(n24353), .B(n57046), .ZN(n57049) );
  OAI21_X1 U56754 ( .A1(n57051), .A2(n57050), .B(n57049), .ZN(n57052) );
  NAND2_X1 U56755 ( .A1(n57064), .A2(n57063), .ZN(n57065) );
  NAND4_X1 U56761 ( .A1(n57088), .A2(n57087), .A3(n57138), .A4(n57086), .ZN(
        n57095) );
  AOI21_X1 U56762 ( .A1(n57433), .A2(n57099), .B(n57089), .ZN(n57094) );
  NAND2_X1 U56763 ( .A1(n23538), .A2(n21829), .ZN(n57090) );
  AOI22_X1 U56764 ( .A1(n57092), .A2(n23302), .B1(n57120), .B2(n57091), .ZN(
        n57093) );
  NAND3_X1 U56766 ( .A1(n4030), .A2(n57015), .A3(n23538), .ZN(n57097) );
  NOR2_X1 U56773 ( .A1(n57123), .A2(n57124), .ZN(n57107) );
  NAND2_X1 U56774 ( .A1(n57015), .A2(n21829), .ZN(n57121) );
  NOR2_X1 U56775 ( .A1(n57105), .A2(n57121), .ZN(n57106) );
  NOR2_X1 U56776 ( .A1(n57128), .A2(n21569), .ZN(n57158) );
  NAND3_X1 U56778 ( .A1(n57132), .A2(n57148), .A3(n23302), .ZN(n57119) );
  INV_X1 U56779 ( .I(n57123), .ZN(n57127) );
  NAND2_X1 U56782 ( .A1(n57127), .A2(n57157), .ZN(n57130) );
  NAND2_X1 U56783 ( .A1(n57132), .A2(n63784), .ZN(n57135) );
  NAND3_X1 U56785 ( .A1(n57233), .A2(n15877), .A3(n57144), .ZN(n57150) );
  NAND3_X1 U56786 ( .A1(n57148), .A2(n61760), .A3(n23302), .ZN(n57149) );
  NAND2_X1 U56787 ( .A1(n61687), .A2(n4030), .ZN(n57153) );
  OAI21_X1 U56788 ( .A1(n57158), .A2(n57157), .B(n57156), .ZN(n57161) );
  NOR2_X2 U1993 ( .A1(n41856), .A2(n42502), .ZN(n41280) );
  BUF_X4 U3005 ( .I(n22444), .Z(n17590) );
  NAND2_X2 U1225 ( .A1(n46985), .A2(n45521), .ZN(n11250) );
  NOR2_X2 U177 ( .A1(n9777), .A2(n58828), .ZN(n9065) );
  NOR3_X2 U44810 ( .A1(n29705), .A2(n1970), .A3(n28624), .ZN(n27811) );
  INV_X2 U1865 ( .I(n2787), .ZN(n42294) );
  BUF_X2 U19901 ( .I(n28631), .Z(n23825) );
  NOR2_X2 U3138 ( .A1(n29915), .A2(n31129), .ZN(n29565) );
  BUF_X4 U7509 ( .I(n60930), .Z(n5126) );
  INV_X2 U10046 ( .I(n43458), .ZN(n43457) );
  INV_X4 U42804 ( .I(n26391), .ZN(n28495) );
  INV_X2 U1231 ( .I(n16742), .ZN(n45639) );
  NOR2_X2 U968 ( .A1(n9177), .A2(n49300), .ZN(n49499) );
  INV_X2 U1385 ( .I(n44897), .ZN(n25531) );
  NAND2_X2 U16370 ( .A1(n4049), .A2(n25426), .ZN(n4048) );
  NAND2_X2 U19222 ( .A1(n6680), .A2(n59046), .ZN(n17631) );
  INV_X2 U37588 ( .I(n25426), .ZN(n44973) );
  INV_X2 U11688 ( .I(n4189), .ZN(n15085) );
  AOI21_X2 U1453 ( .A1(n41245), .A2(n41244), .B(n41243), .ZN(n45836) );
  BUF_X4 U19361 ( .I(n27988), .Z(n23901) );
  INV_X4 U3119 ( .I(n10585), .ZN(n31264) );
  INV_X2 U2675 ( .I(n12479), .ZN(n33752) );
  NAND2_X2 U4075 ( .A1(n45606), .A2(n61582), .ZN(n48975) );
  NAND2_X2 U24913 ( .A1(n22817), .A2(n58373), .ZN(n55658) );
  NOR3_X2 U10783 ( .A1(n14068), .A2(n14067), .A3(n14070), .ZN(n4785) );
  INV_X2 U1714 ( .I(n39082), .ZN(n42180) );
  NOR2_X2 U153 ( .A1(n53351), .A2(n53345), .ZN(n53321) );
  INV_X2 U1134 ( .I(n10333), .ZN(n22899) );
  INV_X4 U2673 ( .I(n33), .ZN(n7047) );
  NOR2_X2 U2611 ( .A1(n35629), .A2(n33319), .ZN(n35201) );
  INV_X2 U2119 ( .I(n26146), .ZN(n23518) );
  NOR3_X2 U9526 ( .A1(n26224), .A2(n33321), .A3(n33322), .ZN(n24634) );
  INV_X2 U2309 ( .I(n36769), .ZN(n35414) );
  BUF_X4 U25289 ( .I(n51482), .Z(n5603) );
  INV_X2 U2146 ( .I(n57313), .ZN(n18057) );
  AOI21_X2 U1452 ( .A1(n39939), .A2(n39940), .B(n5030), .ZN(n39943) );
  NAND3_X2 U27520 ( .A1(n39894), .A2(n40090), .A3(n20751), .ZN(n42483) );
  INV_X2 U31728 ( .I(n30450), .ZN(n11425) );
  NOR2_X2 U1713 ( .A1(n16850), .A2(n42347), .ZN(n42171) );
  INV_X2 U4262 ( .I(n23162), .ZN(n43960) );
  INV_X2 U12040 ( .I(n26834), .ZN(n8302) );
  NOR2_X2 U9490 ( .A1(n2117), .A2(n798), .ZN(n36478) );
  INV_X4 U8874 ( .I(n32972), .ZN(n2618) );
  NAND2_X2 U16543 ( .A1(n42007), .A2(n60472), .ZN(n7400) );
  NOR2_X2 U3367 ( .A1(n27374), .A2(n23568), .ZN(n3626) );
  INV_X2 U251 ( .I(n22755), .ZN(n53147) );
  INV_X4 U1992 ( .I(n21701), .ZN(n1721) );
  NOR2_X2 U8373 ( .A1(n58888), .A2(n36538), .ZN(n36393) );
  INV_X2 U10435 ( .I(n2310), .ZN(n1842) );
  OAI21_X2 U11620 ( .A1(n33299), .A2(n35692), .B(n35690), .ZN(n33021) );
  NOR2_X2 U2751 ( .A1(n5411), .A2(n5410), .ZN(n5409) );
  BUF_X2 U16408 ( .I(n43261), .Z(n23365) );
  INV_X2 U1203 ( .I(n16882), .ZN(n48653) );
  INV_X2 U1265 ( .I(n7318), .ZN(n47536) );
  NOR2_X2 U8011 ( .A1(n7282), .A2(n42019), .ZN(n10806) );
  NOR2_X2 U2298 ( .A1(n1782), .A2(n36483), .ZN(n6329) );
  BUF_X2 U17617 ( .I(n39551), .Z(n23115) );
  BUF_X4 U10614 ( .I(n26034), .Z(n5371) );
  INV_X4 U2002 ( .I(n41306), .ZN(n42453) );
  INV_X4 U11534 ( .I(n22936), .ZN(n1780) );
  NOR2_X2 U4371 ( .A1(n13071), .A2(n1889), .ZN(n27896) );
  AOI22_X2 U10549 ( .A1(n27178), .A2(n27605), .B1(n28306), .B2(n27177), .ZN(
        n14028) );
  NOR3_X2 U10517 ( .A1(n12281), .A2(n27599), .A3(n12278), .ZN(n12277) );
  AOI21_X2 U2195 ( .A1(n36480), .A2(n35958), .B(n2092), .ZN(n11493) );
  NAND2_X2 U7160 ( .A1(n12806), .A2(n38932), .ZN(n12805) );
  INV_X2 U2213 ( .I(n35529), .ZN(n19560) );
  NOR2_X2 U421 ( .A1(n8122), .A2(n24944), .ZN(n9111) );
  INV_X2 U2133 ( .I(n57458), .ZN(n1752) );
  NAND3_X2 U13228 ( .A1(n19630), .A2(n19633), .A3(n35170), .ZN(n8495) );
  INV_X4 U3347 ( .I(n27178), .ZN(n19156) );
  NAND2_X2 U8988 ( .A1(n28466), .A2(n29714), .ZN(n8087) );
  INV_X2 U11735 ( .I(n21083), .ZN(n21707) );
  NAND2_X2 U3418 ( .A1(n29317), .A2(n28858), .ZN(n27360) );
  NAND2_X2 U860 ( .A1(n1639), .A2(n49610), .ZN(n49607) );
  INV_X2 U14085 ( .I(n1439), .ZN(n5290) );
  INV_X2 U2602 ( .I(n33613), .ZN(n1796) );
  INV_X4 U2478 ( .I(n15045), .ZN(n2059) );
  NAND2_X2 U86 ( .A1(n56191), .A2(n5193), .ZN(n56150) );
  NAND2_X2 U2445 ( .A1(n37233), .A2(n61438), .ZN(n20007) );
  NOR2_X2 U9635 ( .A1(n30641), .A2(n30651), .ZN(n29952) );
  INV_X2 U2801 ( .I(n9166), .ZN(n33176) );
  INV_X2 U39206 ( .I(n23683), .ZN(n32101) );
  NAND2_X2 U1977 ( .A1(n41082), .A2(n40592), .ZN(n41077) );
  NOR2_X2 U4356 ( .A1(n2958), .A2(n9830), .ZN(n12301) );
  BUF_X4 U1325 ( .I(n44376), .Z(n47034) );
  NAND2_X2 U9671 ( .A1(n2921), .A2(n30767), .ZN(n30770) );
  INV_X4 U3414 ( .I(n27841), .ZN(n28483) );
  NAND2_X2 U4036 ( .A1(n12074), .A2(n21248), .ZN(n17138) );
  NAND2_X2 U2300 ( .A1(n37049), .A2(n22892), .ZN(n37044) );
  INV_X2 U9593 ( .I(n33975), .ZN(n34602) );
  NAND2_X2 U4362 ( .A1(n3618), .A2(n41506), .ZN(n42867) );
  NOR2_X2 U7094 ( .A1(n1793), .A2(n35096), .ZN(n35997) );
  NAND2_X2 U1960 ( .A1(n40936), .A2(n40464), .ZN(n40925) );
  NAND2_X2 U729 ( .A1(n49211), .A2(n49383), .ZN(n48870) );
  NOR3_X2 U8484 ( .A1(n6011), .A2(n6010), .A3(n6009), .ZN(n6008) );
  NOR3_X2 U15436 ( .A1(n49168), .A2(n48282), .A3(n48281), .ZN(n22656) );
  INV_X2 U14927 ( .I(n56604), .ZN(n52688) );
  NAND3_X2 U1106 ( .A1(n15666), .A2(n1267), .A3(n45765), .ZN(n45510) );
  NOR2_X2 U828 ( .A1(n50059), .A2(n1643), .ZN(n50312) );
  BUF_X4 U945 ( .I(n49888), .Z(n1224) );
  INV_X2 U1980 ( .I(n40850), .ZN(n14132) );
  NAND2_X2 U7220 ( .A1(n3729), .A2(n8373), .ZN(n41321) );
  BUF_X4 U9075 ( .I(Key[90]), .Z(n55034) );
  INV_X4 U5294 ( .I(n40469), .ZN(n40464) );
  NAND2_X2 U3387 ( .A1(n27691), .A2(n27822), .ZN(n29709) );
  NOR2_X2 U8228 ( .A1(n20391), .A2(n30632), .ZN(n31201) );
  NAND3_X2 U2179 ( .A1(n3316), .A2(n36481), .A3(n3315), .ZN(n3314) );
  NAND2_X2 U17348 ( .A1(n9091), .A2(n321), .ZN(n9090) );
  NOR2_X2 U3152 ( .A1(n29860), .A2(n58424), .ZN(n29099) );
  INV_X2 U526 ( .I(n55017), .ZN(n54461) );
  INV_X4 U3425 ( .I(n24951), .ZN(n28400) );
  OAI21_X2 U1777 ( .A1(n41176), .A2(n39141), .B(n10022), .ZN(n38611) );
  NAND2_X2 U719 ( .A1(n22717), .A2(n1643), .ZN(n50143) );
  BUF_X4 U529 ( .I(n7055), .Z(n5129) );
  INV_X2 U3220 ( .I(n27389), .ZN(n27388) );
  NAND2_X2 U1526 ( .A1(n17467), .A2(n42672), .ZN(n42677) );
  NOR2_X2 U9094 ( .A1(n56088), .A2(n56091), .ZN(n56110) );
  NOR2_X2 U12777 ( .A1(n11607), .A2(n11606), .ZN(n13832) );
  AOI22_X2 U24103 ( .A1(n35370), .A2(n35369), .B1(n36170), .B2(n36420), .ZN(
        n12500) );
  NOR2_X2 U2734 ( .A1(n3082), .A2(n24077), .ZN(n34550) );
  OAI21_X2 U10254 ( .A1(n20085), .A2(n57209), .B(n7230), .ZN(n36961) );
  INV_X2 U1217 ( .I(n9140), .ZN(n3341) );
  NAND3_X2 U316 ( .A1(n54841), .A2(n54842), .A3(n54840), .ZN(n3207) );
  NAND3_X2 U10086 ( .A1(n39865), .A2(n39866), .A3(n39864), .ZN(n25538) );
  NAND2_X2 U3161 ( .A1(n7918), .A2(n7913), .ZN(n30267) );
  INV_X4 U39133 ( .I(n23343), .ZN(n33269) );
  BUF_X4 U8816 ( .I(n36020), .Z(n4802) );
  INV_X2 U3283 ( .I(n25619), .ZN(n27509) );
  INV_X4 U37587 ( .I(n21158), .ZN(n28073) );
  BUF_X4 U19924 ( .I(Key[55]), .Z(n54143) );
  BUF_X4 U2134 ( .I(n39670), .Z(n16404) );
  NOR3_X2 U44465 ( .A1(n27032), .A2(n27031), .A3(n27030), .ZN(n27035) );
  NAND2_X2 U18874 ( .A1(n7179), .A2(n7180), .ZN(n25980) );
  INV_X4 U33438 ( .I(n35086), .ZN(n13666) );
  NOR2_X2 U3398 ( .A1(n11617), .A2(n13079), .ZN(n27414) );
  INV_X4 U3056 ( .I(n5070), .ZN(n25848) );
  NAND2_X2 U2939 ( .A1(n29532), .A2(n29533), .ZN(n30495) );
  INV_X4 U42267 ( .I(n18751), .ZN(n27109) );
  NOR2_X2 U1955 ( .A1(n25306), .A2(n39242), .ZN(n39899) );
  OAI21_X2 U1055 ( .A1(n48238), .A2(n48237), .B(n48236), .ZN(n14769) );
  NAND3_X2 U9399 ( .A1(n40032), .A2(n40031), .A3(n40030), .ZN(n40033) );
  OAI21_X2 U1056 ( .A1(n47621), .A2(n1069), .B(n1663), .ZN(n47627) );
  NOR2_X2 U75 ( .A1(n55068), .A2(n15520), .ZN(n55079) );
  NAND2_X2 U3142 ( .A1(n18129), .A2(n1319), .ZN(n29748) );
  INV_X2 U3066 ( .I(n30844), .ZN(n23055) );
  INV_X2 U3403 ( .I(n28542), .ZN(n28534) );
  NOR2_X2 U10530 ( .A1(n23798), .A2(n15197), .ZN(n12131) );
  NAND3_X2 U14054 ( .A1(n28480), .A2(n28479), .A3(n28478), .ZN(n28481) );
  BUF_X4 U21385 ( .I(n5312), .Z(n2952) );
  BUF_X4 U10065 ( .I(n43382), .Z(n18398) );
  AOI21_X2 U3584 ( .A1(n42020), .A2(n20283), .B(n2148), .ZN(n8193) );
  INV_X4 U3344 ( .I(n29317), .ZN(n29310) );
  INV_X2 U1380 ( .I(n15401), .ZN(n46343) );
  BUF_X4 U18841 ( .I(n17700), .Z(n12591) );
  NOR3_X2 U18284 ( .A1(n21812), .A2(n21810), .A3(n21809), .ZN(n21808) );
  INV_X4 U1719 ( .I(n21377), .ZN(n11883) );
  INV_X2 U2026 ( .I(n39414), .ZN(n40076) );
  AND2_X2 U8691 ( .A1(n462), .A2(n4714), .Z(n40903) );
  NAND2_X2 U19437 ( .A1(n27021), .A2(n27020), .ZN(n27026) );
  INV_X4 U34101 ( .I(n27233), .ZN(n14869) );
  INV_X2 U2165 ( .I(n14550), .ZN(n38468) );
  INV_X2 U2799 ( .I(n31823), .ZN(n32661) );
  NAND2_X2 U1593 ( .A1(n13478), .A2(n57198), .ZN(n43467) );
  INV_X2 U2079 ( .I(n5868), .ZN(n41289) );
  NOR2_X2 U1589 ( .A1(n1495), .A2(n44226), .ZN(n4282) );
  INV_X2 U4283 ( .I(n15457), .ZN(n47603) );
  NOR2_X2 U725 ( .A1(n19523), .A2(n61530), .ZN(n49926) );
  NAND2_X2 U2515 ( .A1(n61795), .A2(n7016), .ZN(n33987) );
  NAND2_X2 U44398 ( .A1(n23797), .A2(n28858), .ZN(n27451) );
  INV_X4 U1665 ( .I(n8589), .ZN(n41350) );
  BUF_X2 U10629 ( .I(Key[65]), .Z(n54289) );
  INV_X2 U2380 ( .I(n36026), .ZN(n21329) );
  NAND2_X2 U1157 ( .A1(n45746), .A2(n47470), .ZN(n46987) );
  NOR2_X2 U1942 ( .A1(n25666), .A2(n64914), .ZN(n40349) );
  INV_X4 U3415 ( .I(n14633), .ZN(n23474) );
  NAND2_X2 U11423 ( .A1(n5734), .A2(n37393), .ZN(n2918) );
  BUF_X4 U1283 ( .I(n44551), .Z(n46033) );
  INV_X4 U539 ( .I(n53917), .ZN(n14446) );
  NOR3_X2 U28558 ( .A1(n34825), .A2(n36040), .A3(n8474), .ZN(n35391) );
  NOR3_X2 U18151 ( .A1(n32996), .A2(n35197), .A3(n32995), .ZN(n32997) );
  NAND2_X2 U1671 ( .A1(n41660), .A2(n42180), .ZN(n41670) );
  NOR2_X2 U3377 ( .A1(n28615), .A2(n28616), .ZN(n28617) );
  INV_X2 U2792 ( .I(n12014), .ZN(n32591) );
  INV_X4 U2476 ( .I(n12830), .ZN(n22559) );
  OAI21_X2 U36973 ( .A1(n40545), .A2(n40544), .B(n21376), .ZN(n42854) );
  OAI21_X2 U3216 ( .A1(n22706), .A2(n9251), .B(n27073), .ZN(n27176) );
  INV_X2 U9053 ( .I(n26501), .ZN(n26618) );
  NAND3_X2 U44251 ( .A1(n26710), .A2(n29541), .A3(n26709), .ZN(n26711) );
  INV_X2 U11881 ( .I(n27756), .ZN(n6609) );
  INV_X2 U11992 ( .I(n20860), .ZN(n5659) );
  NOR2_X2 U1621 ( .A1(n43735), .A2(n8290), .ZN(n42845) );
  INV_X8 U24077 ( .I(n37536), .ZN(n42607) );
  NAND2_X2 U129 ( .A1(n17012), .A2(n25604), .ZN(n53346) );
  INV_X2 U1214 ( .I(n8632), .ZN(n17573) );
  INV_X2 U37810 ( .I(n18174), .ZN(n56146) );
  NAND2_X2 U889 ( .A1(n19646), .A2(n49792), .ZN(n13878) );
  NAND2_X2 U3078 ( .A1(n4270), .A2(n10068), .ZN(n29502) );
  NAND4_X2 U35604 ( .A1(n54628), .A2(n54975), .A3(n54627), .A4(n54967), .ZN(
        n54632) );
  OAI21_X2 U264 ( .A1(n21843), .A2(n21842), .B(n52692), .ZN(n56832) );
  INV_X4 U2012 ( .I(n24389), .ZN(n4171) );
  INV_X2 U2472 ( .I(n37397), .ZN(n36821) );
  NAND3_X2 U11919 ( .A1(n5290), .A2(n12030), .A3(n5292), .ZN(n5289) );
  BUF_X4 U4996 ( .I(n30817), .Z(n162) );
  NOR2_X2 U4192 ( .A1(n54285), .A2(n54254), .ZN(n54211) );
  NAND4_X1 U43442 ( .A1(n54336), .A2(n54335), .A3(n54447), .A4(n54334), .ZN(
        n54337) );
  INV_X2 U46468 ( .I(n31757), .ZN(n42426) );
  NOR2_X2 U369 ( .A1(n54814), .A2(n5226), .ZN(n54824) );
  BUF_X4 U228 ( .I(n54411), .Z(n5324) );
  BUF_X4 U12114 ( .I(Key[91]), .Z(n55052) );
  NAND2_X2 U22363 ( .A1(n29824), .A2(n1208), .ZN(n28083) );
  NOR3_X1 U11740 ( .A1(n2283), .A2(n2281), .A3(n2280), .ZN(n2297) );
  NOR3_X1 U27562 ( .A1(n49113), .A2(n49112), .A3(n49795), .ZN(n49120) );
  INV_X2 U8933 ( .I(n31138), .ZN(n31146) );
  NAND2_X2 U1222 ( .A1(n1294), .A2(n10428), .ZN(n16974) );
  INV_X2 U8756 ( .I(n9606), .ZN(n11959) );
  NOR2_X2 U12766 ( .A1(n1686), .A2(n1394), .ZN(n11926) );
  BUF_X4 U1723 ( .I(n42695), .Z(n2160) );
  INV_X2 U8616 ( .I(n47664), .ZN(n47844) );
  OAI21_X2 U2944 ( .A1(n30370), .A2(n18810), .B(n29480), .ZN(n31136) );
  NAND2_X2 U4600 ( .A1(n30538), .A2(n24298), .ZN(n30439) );
  INV_X4 U2606 ( .I(n17538), .ZN(n35294) );
  AND2_X2 U10146 ( .A1(n6853), .A2(n57615), .Z(n6852) );
  NAND2_X2 U14104 ( .A1(n6826), .A2(n6827), .ZN(n6825) );
  BUF_X4 U12954 ( .I(n42822), .Z(n17467) );
  INV_X2 U1258 ( .I(n24759), .ZN(n45576) );
  NAND2_X2 U4277 ( .A1(n53077), .A2(n53115), .ZN(n53107) );
  NOR2_X2 U4156 ( .A1(n48594), .A2(n1265), .ZN(n46096) );
  NAND2_X2 U3082 ( .A1(n18839), .A2(n17627), .ZN(n7683) );
  NOR2_X2 U3940 ( .A1(n54625), .A2(n61509), .ZN(n54974) );
  INV_X8 U234 ( .I(n55627), .ZN(n55643) );
  INV_X2 U9889 ( .I(n50000), .ZN(n50006) );
  NAND2_X2 U191 ( .A1(n5051), .A2(n1233), .ZN(n55096) );
  NOR2_X2 U3019 ( .A1(n30786), .A2(n17745), .ZN(n11465) );
  AND2_X2 U12088 ( .A1(n23303), .A2(n26431), .Z(n3211) );
  NAND2_X2 U1809 ( .A1(n42302), .A2(n42510), .ZN(n42298) );
  NAND2_X2 U3058 ( .A1(n1352), .A2(n30492), .ZN(n25526) );
  NAND2_X2 U3096 ( .A1(n22877), .A2(n19830), .ZN(n30126) );
  INV_X2 U4349 ( .I(n20763), .ZN(n49659) );
  NOR2_X2 U4151 ( .A1(n43150), .A2(n20602), .ZN(n43163) );
  OAI21_X2 U11600 ( .A1(n34170), .A2(n11874), .B(n34169), .ZN(n34174) );
  NOR2_X2 U1068 ( .A1(n46985), .A2(n4380), .ZN(n46980) );
  INV_X4 U43033 ( .I(n1623), .ZN(n51313) );
  BUF_X4 U16944 ( .I(n43166), .Z(n23709) );
  NAND2_X2 U812 ( .A1(n19544), .A2(n62700), .ZN(n26102) );
  NOR2_X2 U22263 ( .A1(n20507), .A2(n34606), .ZN(n33975) );
  INV_X4 U1148 ( .I(n19142), .ZN(n48552) );
  INV_X2 U143 ( .I(n58808), .ZN(n55218) );
  NAND2_X2 U8322 ( .A1(n16869), .A2(n21008), .ZN(n33718) );
  NAND2_X2 U11577 ( .A1(n12913), .A2(n12952), .ZN(n12912) );
  OAI21_X2 U10314 ( .A1(n34509), .A2(n34508), .B(n63421), .ZN(n12913) );
  INV_X4 U39351 ( .I(n30743), .ZN(n30736) );
  NOR2_X2 U996 ( .A1(n25486), .A2(n15145), .ZN(n12829) );
  INV_X2 U498 ( .I(n55672), .ZN(n55456) );
  INV_X2 U11511 ( .I(n36393), .ZN(n18566) );
  INV_X4 U11329 ( .I(n24302), .ZN(n40695) );
  INV_X2 U47597 ( .I(n34730), .ZN(n33741) );
  INV_X2 U858 ( .I(n47923), .ZN(n1628) );
  NOR2_X2 U8870 ( .A1(n35688), .A2(n22597), .ZN(n35692) );
  NAND3_X2 U3981 ( .A1(n23226), .A2(n36288), .A3(n6831), .ZN(n2220) );
  NOR2_X2 U6842 ( .A1(n2168), .A2(n21252), .ZN(n20260) );
  OR2_X1 U37557 ( .A1(n21127), .A2(n18918), .Z(n15961) );
  INV_X2 U7002 ( .I(n28920), .ZN(n24316) );
  NAND2_X2 U2972 ( .A1(n23446), .A2(n4270), .ZN(n29007) );
  NAND2_X2 U31535 ( .A1(n27040), .A2(n4443), .ZN(n16902) );
  INV_X4 U727 ( .I(n18882), .ZN(n50444) );
  NAND2_X2 U2034 ( .A1(n40617), .A2(n61333), .ZN(n39129) );
  INV_X2 U1103 ( .I(n4660), .ZN(n48144) );
  NOR2_X2 U1251 ( .A1(n47087), .A2(n14518), .ZN(n14517) );
  INV_X2 U10511 ( .I(n23024), .ZN(n25639) );
  NOR2_X2 U2460 ( .A1(n36926), .A2(n34926), .ZN(n36923) );
  INV_X2 U4073 ( .I(n6016), .ZN(n42499) );
  INV_X4 U20330 ( .I(n2636), .ZN(n2267) );
  NOR2_X2 U14060 ( .A1(n28613), .A2(n13010), .ZN(n13009) );
  INV_X2 U11927 ( .I(n28441), .ZN(n28613) );
  BUF_X4 U549 ( .I(n52622), .Z(n54640) );
  NOR2_X2 U91 ( .A1(n7680), .A2(n1919), .ZN(n54912) );
  INV_X2 U37474 ( .I(n40651), .ZN(n23434) );
  INV_X2 U8693 ( .I(n43151), .ZN(n42901) );
  NOR2_X2 U40124 ( .A1(n28862), .A2(n27454), .ZN(n27457) );
  NOR3_X2 U5548 ( .A1(n15992), .A2(n26398), .A3(n26397), .ZN(n27843) );
  INV_X4 U7675 ( .I(n36262), .ZN(n9041) );
  NOR2_X2 U500 ( .A1(n5907), .A2(n55440), .ZN(n55316) );
  NAND3_X2 U37289 ( .A1(n54971), .A2(n7518), .A3(n58491), .ZN(n54967) );
  INV_X1 U5825 ( .I(n1146), .ZN(n54622) );
  NAND2_X2 U2655 ( .A1(n35273), .A2(n34385), .ZN(n34300) );
  INV_X2 U23654 ( .I(n54952), .ZN(n14468) );
  BUF_X2 U19743 ( .I(n27837), .Z(n10131) );
  NOR2_X2 U1419 ( .A1(n41587), .A2(n5928), .ZN(n12563) );
  INV_X8 U43320 ( .I(n23056), .ZN(n30702) );
  BUF_X8 U52493 ( .I(n45442), .Z(n50427) );
  NOR2_X2 U3395 ( .A1(n23737), .A2(n27574), .ZN(n26653) );
  INV_X2 U594 ( .I(n24537), .ZN(n21481) );
  NOR3_X1 U33671 ( .A1(n14036), .A2(n23459), .A3(n48319), .ZN(n48320) );
  BUF_X4 U973 ( .I(n50271), .Z(n22694) );
  NAND2_X2 U14021 ( .A1(n17307), .A2(n19678), .ZN(n9959) );
  AOI22_X2 U4001 ( .A1(n14209), .A2(n49526), .B1(n1374), .B2(n65005), .ZN(
        n14208) );
  NOR2_X2 U901 ( .A1(n25857), .A2(n49195), .ZN(n49526) );
  NAND2_X2 U9577 ( .A1(n35037), .A2(n60984), .ZN(n34500) );
  NAND2_X2 U68 ( .A1(n55893), .A2(n60203), .ZN(n55886) );
  NAND2_X2 U906 ( .A1(n50340), .A2(n50346), .ZN(n23414) );
  NAND2_X2 U7275 ( .A1(n50394), .A2(n50406), .ZN(n50082) );
  OAI21_X2 U1611 ( .A1(n64363), .A2(n63392), .B(n1269), .ZN(n42560) );
  NOR2_X2 U3392 ( .A1(n23997), .A2(n23209), .ZN(n27123) );
  NAND2_X2 U8650 ( .A1(n46333), .A2(n46332), .ZN(n46328) );
  NOR2_X1 U25031 ( .A1(n5337), .A2(n5336), .ZN(n5335) );
  INV_X2 U3207 ( .I(n26665), .ZN(n27580) );
  BUF_X4 U6466 ( .I(n35570), .Z(n576) );
  NAND2_X2 U714 ( .A1(n1643), .A2(n3054), .ZN(n50307) );
  NOR2_X1 U23513 ( .A1(n42645), .A2(n43532), .ZN(n43777) );
  NAND2_X2 U8878 ( .A1(n34627), .A2(n31509), .ZN(n34618) );
  NOR2_X2 U13806 ( .A1(n60030), .A2(n8804), .ZN(n28994) );
  INV_X4 U5176 ( .I(n35508), .ZN(n3561) );
  INV_X4 U23635 ( .I(n10830), .ZN(n10821) );
  NOR2_X2 U3379 ( .A1(n28040), .A2(n2941), .ZN(n28036) );
  NAND2_X2 U2904 ( .A1(n27362), .A2(n30063), .ZN(n30058) );
  NAND3_X2 U3223 ( .A1(n27338), .A2(n29385), .A3(n27339), .ZN(n10642) );
  INV_X2 U19249 ( .I(n14944), .ZN(n16979) );
  AND2_X2 U216 ( .A1(n15928), .A2(n53014), .Z(n53781) );
  INV_X2 U7128 ( .I(n41887), .ZN(n41876) );
  NAND2_X2 U2413 ( .A1(n5734), .A2(n8808), .ZN(n8816) );
  INV_X4 U2748 ( .I(n34714), .ZN(n23556) );
  INV_X1 U32944 ( .I(n15777), .ZN(n56586) );
  INV_X2 U53047 ( .I(n47128), .ZN(n48078) );
  NOR2_X2 U8913 ( .A1(n57952), .A2(n15136), .ZN(n16116) );
  INV_X2 U2839 ( .I(n22751), .ZN(n16625) );
  OAI21_X2 U1798 ( .A1(n41036), .A2(n41037), .B(n1747), .ZN(n41040) );
  NAND2_X2 U3306 ( .A1(n28459), .A2(n28610), .ZN(n5268) );
  NOR2_X2 U2431 ( .A1(n35965), .A2(n35962), .ZN(n35972) );
  NOR2_X2 U11957 ( .A1(n26905), .A2(n10544), .ZN(n28605) );
  INV_X2 U19735 ( .I(n28444), .ZN(n26905) );
  INV_X4 U3436 ( .I(n13399), .ZN(n23033) );
  NOR2_X2 U10441 ( .A1(n21964), .A2(n30046), .ZN(n30260) );
  INV_X2 U3686 ( .I(n32892), .ZN(n34198) );
  INV_X2 U211 ( .I(n15928), .ZN(n53820) );
  NAND2_X2 U2405 ( .A1(n6540), .A2(n8195), .ZN(n36828) );
  INV_X4 U2011 ( .I(n39028), .ZN(n20555) );
  NOR2_X2 U2667 ( .A1(n33568), .A2(n4034), .ZN(n33096) );
  INV_X4 U29658 ( .I(n24195), .ZN(n20183) );
  NAND2_X2 U1608 ( .A1(n15539), .A2(n42985), .ZN(n16911) );
  INV_X2 U1378 ( .I(n44594), .ZN(n46557) );
  INV_X4 U130 ( .I(n56803), .ZN(n56791) );
  INV_X2 U14146 ( .I(n29339), .ZN(n29344) );
  NOR2_X2 U3439 ( .A1(n29636), .A2(n29641), .ZN(n28587) );
  NAND2_X2 U4133 ( .A1(n56422), .A2(n56204), .ZN(n52717) );
  NAND2_X2 U2411 ( .A1(n35965), .A2(n35971), .ZN(n22116) );
  NAND3_X2 U14018 ( .A1(n13381), .A2(n26505), .A3(n13380), .ZN(n7062) );
  NOR2_X2 U7283 ( .A1(n5629), .A2(n49014), .ZN(n5628) );
  NOR2_X2 U9325 ( .A1(n43913), .A2(n21073), .ZN(n43929) );
  INV_X2 U7039 ( .I(n9319), .ZN(n32036) );
  NOR2_X2 U3092 ( .A1(n5768), .A2(n30588), .ZN(n5285) );
  NOR2_X2 U2392 ( .A1(n13983), .A2(n57209), .ZN(n36626) );
  AOI21_X2 U12389 ( .A1(n49607), .A2(n49308), .B(n23656), .ZN(n26031) );
  INV_X2 U2760 ( .I(n60937), .ZN(n25465) );
  NAND2_X2 U3993 ( .A1(n3029), .A2(n10939), .ZN(n2749) );
  NOR2_X2 U9841 ( .A1(n56204), .A2(n56630), .ZN(n56639) );
  NOR2_X2 U14039 ( .A1(n27555), .A2(n21000), .ZN(n14650) );
  INV_X4 U2452 ( .I(n19231), .ZN(n1415) );
  BUF_X4 U942 ( .I(n45895), .Z(n49940) );
  NOR3_X2 U4346 ( .A1(n27096), .A2(n6047), .A3(n10729), .ZN(n6120) );
  NAND2_X2 U12898 ( .A1(n10897), .A2(n24779), .ZN(n9377) );
  INV_X2 U10745 ( .I(n10441), .ZN(n54801) );
  NAND2_X2 U4011 ( .A1(n64166), .A2(n4594), .ZN(n50339) );
  NOR2_X2 U15732 ( .A1(n47677), .A2(n7491), .ZN(n10490) );
  NAND3_X2 U12547 ( .A1(n18264), .A2(n47676), .A3(n47675), .ZN(n7491) );
  OR2_X2 U24008 ( .A1(n11416), .A2(n195), .Z(n45527) );
  OAI21_X2 U38024 ( .A1(n17278), .A2(n16707), .B(n28551), .ZN(n17277) );
  NAND2_X2 U1562 ( .A1(n43975), .A2(n21360), .ZN(n43715) );
  NOR2_X2 U3397 ( .A1(n22352), .A2(n28552), .ZN(n28551) );
  INV_X2 U9261 ( .I(n18321), .ZN(n20938) );
  NAND2_X2 U36164 ( .A1(n20971), .A2(n65061), .ZN(n49369) );
  INV_X4 U428 ( .I(n25215), .ZN(n54970) );
  NAND2_X2 U4384 ( .A1(n19102), .A2(n9143), .ZN(n40090) );
  NAND3_X2 U1543 ( .A1(n42420), .A2(n43478), .A3(n42968), .ZN(n16569) );
  BUF_X4 U12101 ( .I(n26877), .Z(n29609) );
  INV_X2 U410 ( .I(n21893), .ZN(n56632) );
  INV_X4 U2078 ( .I(n38264), .ZN(n42299) );
  NAND2_X2 U8669 ( .A1(n43929), .A2(n43912), .ZN(n43495) );
  INV_X2 U2109 ( .I(n17365), .ZN(n38731) );
  INV_X4 U32476 ( .I(n12477), .ZN(n12739) );
  NOR2_X2 U8858 ( .A1(n22342), .A2(n5529), .ZN(n33758) );
  NAND2_X2 U6994 ( .A1(n6349), .A2(n21176), .ZN(n6509) );
  OAI21_X2 U2901 ( .A1(n31265), .A2(n31266), .B(n61251), .ZN(n9782) );
  INV_X8 U41455 ( .I(n15805), .ZN(n37050) );
  NAND2_X2 U2333 ( .A1(n35965), .A2(n35964), .ZN(n13769) );
  NOR2_X2 U2015 ( .A1(n1743), .A2(n38932), .ZN(n40400) );
  INV_X1 U42421 ( .I(n28201), .ZN(n25222) );
  INV_X1 U25384 ( .I(n8026), .ZN(n9444) );
  BUF_X2 U14258 ( .I(n26501), .Z(n23737) );
  NAND2_X2 U1417 ( .A1(n10199), .A2(n43663), .ZN(n16519) );
  INV_X2 U10523 ( .I(n44602), .ZN(n46414) );
  INV_X4 U1924 ( .I(n42251), .ZN(n42242) );
  NAND2_X2 U8409 ( .A1(n16798), .A2(n15757), .ZN(n47197) );
  INV_X2 U24285 ( .I(n43468), .ZN(n13750) );
  BUF_X4 U38919 ( .I(n23024), .Z(n18075) );
  NAND2_X2 U36651 ( .A1(n40850), .A2(n64459), .ZN(n40593) );
  NOR2_X2 U2603 ( .A1(n34993), .A2(n21008), .ZN(n34982) );
  NAND3_X2 U26927 ( .A1(n34154), .A2(n26122), .A3(n34153), .ZN(n23353) );
  INV_X1 U509 ( .I(n54459), .ZN(n3916) );
  INV_X4 U8249 ( .I(n25449), .ZN(n29835) );
  INV_X2 U46476 ( .I(n31508), .ZN(n31509) );
  INV_X4 U4433 ( .I(n43764), .ZN(n46550) );
  INV_X2 U527 ( .I(n6095), .ZN(n54634) );
  NAND2_X2 U2327 ( .A1(n23584), .A2(n10596), .ZN(n34877) );
  NOR2_X2 U3118 ( .A1(n22411), .A2(n24504), .ZN(n7130) );
  NAND4_X2 U48932 ( .A1(n36889), .A2(n5936), .A3(n36888), .A4(n9456), .ZN(
        n36890) );
  NAND2_X2 U10564 ( .A1(n4324), .A2(n26363), .ZN(n27581) );
  INV_X2 U1318 ( .I(n13438), .ZN(n46106) );
  NOR2_X2 U3014 ( .A1(n29523), .A2(n17414), .ZN(n29858) );
  NAND2_X2 U10933 ( .A1(n48244), .A2(n3364), .ZN(n48242) );
  NAND3_X1 U42501 ( .A1(n23457), .A2(n56141), .A3(n23456), .ZN(n56142) );
  NAND3_X2 U24209 ( .A1(n33714), .A2(n33713), .A3(n33710), .ZN(n19949) );
  AND2_X2 U1263 ( .A1(n22283), .A2(n13029), .Z(n1082) );
  INV_X2 U4457 ( .I(n10806), .ZN(n18363) );
  NAND2_X2 U20344 ( .A1(n2177), .A2(n14944), .ZN(n18476) );
  INV_X2 U39012 ( .I(n22617), .ZN(n18241) );
  INV_X2 U2294 ( .I(n21801), .ZN(n36175) );
  NOR2_X2 U11784 ( .A1(n28099), .A2(n29460), .ZN(n28735) );
  NOR2_X2 U1211 ( .A1(n22386), .A2(n47603), .ZN(n45568) );
  NAND2_X2 U12636 ( .A1(n3203), .A2(n47317), .ZN(n5297) );
  INV_X2 U8515 ( .I(n24586), .ZN(n54350) );
  NAND3_X2 U9669 ( .A1(n20755), .A2(n25466), .A3(n8803), .ZN(n29841) );
  OR2_X2 U2047 ( .A1(n39994), .A2(n41383), .Z(n14616) );
  INV_X2 U14259 ( .I(n26730), .ZN(n29119) );
  NAND3_X2 U13301 ( .A1(n3768), .A2(n3767), .A3(n3766), .ZN(n3765) );
  INV_X2 U10830 ( .I(n47787), .ZN(n48337) );
  NAND2_X2 U1580 ( .A1(n20180), .A2(n1718), .ZN(n42551) );
  NAND2_X2 U50182 ( .A1(n42788), .A2(n41665), .ZN(n39086) );
  INV_X4 U2057 ( .I(n41401), .ZN(n15548) );
  INV_X2 U9519 ( .I(n36335), .ZN(n36334) );
  NAND2_X2 U7369 ( .A1(n25116), .A2(n53732), .ZN(n50829) );
  INV_X2 U10203 ( .I(n11700), .ZN(n20408) );
  INV_X2 U10437 ( .I(n30324), .ZN(n2120) );
  BUF_X4 U21569 ( .I(n7854), .Z(n3091) );
  INV_X2 U3446 ( .I(n4394), .ZN(n14604) );
  NAND3_X2 U8649 ( .A1(n18673), .A2(n42644), .A3(n43200), .ZN(n16568) );
  NOR2_X1 U19435 ( .A1(n26342), .A2(n27597), .ZN(n14679) );
  NAND2_X2 U1233 ( .A1(n9331), .A2(n47502), .ZN(n44284) );
  NAND2_X2 U1104 ( .A1(n18227), .A2(n70), .ZN(n47671) );
  INV_X2 U523 ( .I(n24318), .ZN(n52819) );
  AND2_X2 U26871 ( .A1(n6100), .A2(n42008), .Z(n43085) );
  NAND2_X2 U385 ( .A1(n52235), .A2(n12818), .ZN(n52739) );
  OR2_X2 U3063 ( .A1(n30748), .A2(n30632), .Z(n20378) );
  NOR3_X2 U6431 ( .A1(n28978), .A2(n2098), .A3(n29260), .ZN(n2097) );
  AOI22_X2 U3187 ( .A1(n13564), .A2(n21804), .B1(n13565), .B2(n3555), .ZN(
        n13563) );
  NAND2_X2 U1286 ( .A1(n1293), .A2(n48103), .ZN(n6805) );
  NAND2_X2 U2920 ( .A1(n30766), .A2(n10926), .ZN(n30666) );
  INV_X2 U2790 ( .I(n31998), .ZN(n31732) );
  NAND2_X2 U10244 ( .A1(n18677), .A2(n15720), .ZN(n35472) );
  INV_X4 U3128 ( .I(n1868), .ZN(n24199) );
  NOR3_X2 U11928 ( .A1(n23703), .A2(n27625), .A3(n27624), .ZN(n22422) );
  NOR2_X2 U2932 ( .A1(n31113), .A2(n64128), .ZN(n14274) );
  BUF_X2 U14282 ( .I(n20716), .Z(n23007) );
  NOR2_X2 U4373 ( .A1(n1889), .A2(n60547), .ZN(n11352) );
  NOR2_X2 U52847 ( .A1(n16493), .A2(n61146), .ZN(n47042) );
  NAND2_X2 U27600 ( .A1(n52690), .A2(n52682), .ZN(n17540) );
  NAND2_X2 U30244 ( .A1(n10023), .A2(n27365), .ZN(n33035) );
  NAND3_X2 U3210 ( .A1(n28012), .A2(n62663), .A3(n7452), .ZN(n28015) );
  NOR2_X2 U2878 ( .A1(n2840), .A2(n2841), .ZN(n73) );
  NAND2_X2 U2254 ( .A1(n15488), .A2(n35903), .ZN(n37029) );
  NAND2_X2 U10536 ( .A1(n28267), .A2(n17103), .ZN(n27419) );
  NOR2_X2 U3081 ( .A1(n31241), .A2(n23008), .ZN(n31253) );
  NAND2_X2 U19697 ( .A1(n26692), .A2(n23504), .ZN(n29333) );
  INV_X2 U1710 ( .I(n42175), .ZN(n42868) );
  NOR2_X2 U3393 ( .A1(n10544), .A2(n28452), .ZN(n28459) );
  NOR3_X2 U9630 ( .A1(n30373), .A2(n30372), .A3(n30371), .ZN(n30380) );
  AOI21_X2 U10692 ( .A1(n18010), .A2(n56360), .B(n56371), .ZN(n18009) );
  NAND4_X2 U15938 ( .A1(n10031), .A2(n44671), .A3(n1087), .A4(n47512), .ZN(
        n19258) );
  INV_X2 U6584 ( .I(n18121), .ZN(n56362) );
  NAND2_X2 U25086 ( .A1(n32831), .A2(n5389), .ZN(n34197) );
  NOR2_X2 U2442 ( .A1(n61703), .A2(n36220), .ZN(n36434) );
  NAND2_X2 U916 ( .A1(n50407), .A2(n50398), .ZN(n49420) );
  NOR2_X2 U7183 ( .A1(n43695), .A2(n42019), .ZN(n42018) );
  NOR2_X2 U45578 ( .A1(n61215), .A2(n31224), .ZN(n30755) );
  INV_X4 U2455 ( .I(n11413), .ZN(n1776) );
  NAND3_X2 U35101 ( .A1(n14202), .A2(n24000), .A3(n60575), .ZN(n29910) );
  NOR4_X2 U38933 ( .A1(n29940), .A2(n29938), .A3(n18120), .A4(n29939), .ZN(
        n29941) );
  INV_X1 U16233 ( .I(n47380), .ZN(n1654) );
  INV_X4 U2090 ( .I(n20552), .ZN(n287) );
  NOR2_X2 U2017 ( .A1(n42267), .A2(n3566), .ZN(n37773) );
  NAND2_X2 U872 ( .A1(n687), .A2(n49698), .ZN(n49762) );
  NAND2_X2 U4107 ( .A1(n29148), .A2(n6888), .ZN(n26376) );
  AND3_X1 U37690 ( .A1(n35735), .A2(n61496), .A3(n35743), .Z(n16215) );
  NAND4_X2 U2868 ( .A1(n29809), .A2(n29810), .A3(n29808), .A4(n29884), .ZN(
        n25318) );
  AND2_X2 U37863 ( .A1(n36953), .A2(n22587), .Z(n36888) );
  BUF_X4 U28946 ( .I(n9427), .Z(n8912) );
  NAND3_X2 U24170 ( .A1(n13651), .A2(n24462), .A3(n13652), .ZN(n24461) );
  INV_X2 U34659 ( .I(n191), .ZN(n32158) );
  INV_X4 U10605 ( .I(n28548), .ZN(n1355) );
  BUF_X4 U8637 ( .I(n47323), .Z(n23588) );
  NOR2_X1 U7301 ( .A1(n4298), .A2(n4296), .ZN(n4295) );
  NOR3_X1 U24335 ( .A1(n61792), .A2(n20245), .A3(n20246), .ZN(n4884) );
  AOI22_X1 U13813 ( .A1(n28773), .A2(n28774), .B1(n8357), .B2(n30723), .ZN(
        n14387) );
  INV_X2 U12700 ( .I(n23114), .ZN(n21231) );
  INV_X2 U8353 ( .I(n6744), .ZN(n25314) );
  INV_X2 U12562 ( .I(n48123), .ZN(n48125) );
  INV_X2 U2688 ( .I(n33453), .ZN(n34679) );
  NAND2_X2 U8790 ( .A1(n25339), .A2(n24041), .ZN(n36820) );
  NOR2_X2 U1854 ( .A1(n19466), .A2(n41054), .ZN(n41873) );
  NAND3_X2 U8365 ( .A1(n33786), .A2(n3057), .A3(n21802), .ZN(n5641) );
  NAND2_X2 U10402 ( .A1(n6318), .A2(n20365), .ZN(n31377) );
  INV_X2 U588 ( .I(n50582), .ZN(n1290) );
  INV_X2 U3409 ( .I(n21656), .ZN(n23568) );
  NOR3_X2 U283 ( .A1(n20003), .A2(n20002), .A3(n20001), .ZN(n20000) );
  NAND2_X2 U47895 ( .A1(n2362), .A2(n36471), .ZN(n34100) );
  NOR2_X2 U13129 ( .A1(n61850), .A2(n59203), .ZN(n39869) );
  NOR2_X2 U48688 ( .A1(n22786), .A2(n23319), .ZN(n38024) );
  BUF_X4 U3080 ( .I(n30492), .Z(n19451) );
  OR3_X2 U22663 ( .A1(n12955), .A2(n42543), .A3(n1714), .Z(n3963) );
  INV_X2 U1415 ( .I(n43878), .ZN(n15354) );
  INV_X1 U2967 ( .I(n28772), .ZN(n29218) );
  INV_X4 U9761 ( .I(n29684), .ZN(n17274) );
  INV_X2 U1902 ( .I(n5362), .ZN(n40150) );
  BUF_X4 U31081 ( .I(n29684), .Z(n10598) );
  NOR2_X2 U37158 ( .A1(n20458), .A2(n49074), .ZN(n48054) );
  NOR2_X2 U1207 ( .A1(n3510), .A2(n47603), .ZN(n45972) );
  NAND2_X2 U799 ( .A1(n15220), .A2(n49803), .ZN(n47941) );
  NAND2_X2 U4220 ( .A1(n54951), .A2(n54778), .ZN(n54430) );
  AOI21_X2 U3769 ( .A1(n17750), .A2(n5847), .B(n14499), .ZN(n14495) );
  NAND2_X2 U9680 ( .A1(n9392), .A2(n24402), .ZN(n29528) );
  AOI21_X1 U23874 ( .A1(n47379), .A2(n47378), .B(n47145), .ZN(n18883) );
  NOR2_X2 U7103 ( .A1(n37957), .A2(n2483), .ZN(n36608) );
  INV_X2 U1983 ( .I(n22304), .ZN(n40732) );
  NOR2_X2 U2876 ( .A1(n14270), .A2(n14274), .ZN(n31121) );
  NAND2_X2 U30124 ( .A1(n17546), .A2(n17913), .ZN(n17545) );
  NAND2_X2 U3015 ( .A1(n30343), .A2(n59268), .ZN(n30610) );
  INV_X4 U14269 ( .I(n28448), .ZN(n28607) );
  NAND2_X2 U8008 ( .A1(n13242), .A2(n42019), .ZN(n22802) );
  INV_X4 U3410 ( .I(n23033), .ZN(n28610) );
  AOI21_X2 U13225 ( .A1(n10707), .A2(n34858), .B(n4769), .ZN(n10706) );
  OAI22_X2 U16654 ( .A1(n16448), .A2(n43414), .B1(n42096), .B2(n42095), .ZN(
        n13080) );
  NAND2_X2 U11860 ( .A1(n29076), .A2(n10240), .ZN(n7252) );
  INV_X2 U1216 ( .I(n45957), .ZN(n47324) );
  INV_X2 U1921 ( .I(n40029), .ZN(n40297) );
  NAND2_X2 U5790 ( .A1(n33453), .A2(n25668), .ZN(n1813) );
  INV_X4 U2477 ( .I(n24934), .ZN(n26243) );
  NAND2_X2 U2269 ( .A1(n25842), .A2(n798), .ZN(n3649) );
  INV_X4 U13712 ( .I(n19868), .ZN(n20326) );
  AOI21_X1 U34912 ( .A1(n34717), .A2(n22797), .B(n17163), .ZN(n17162) );
  INV_X4 U225 ( .I(n56106), .ZN(n56071) );
  INV_X2 U14138 ( .I(n21854), .ZN(n28435) );
  BUF_X4 U31745 ( .I(n52616), .Z(n11448) );
  BUF_X2 U13800 ( .I(n33058), .Z(n21006) );
  BUF_X4 U3156 ( .I(n24334), .Z(n2005) );
  NAND2_X2 U26962 ( .A1(n11621), .A2(n30033), .ZN(n7179) );
  BUF_X2 U10641 ( .I(Key[133]), .Z(n55862) );
  BUF_X4 U12110 ( .I(Key[150]), .Z(n24014) );
  NAND2_X2 U6114 ( .A1(n16902), .A2(n16903), .ZN(n28065) );
  NOR2_X2 U218 ( .A1(n518), .A2(n53294), .ZN(n53306) );
  INV_X2 U27452 ( .I(n8260), .ZN(n25976) );
  NAND2_X2 U2619 ( .A1(n34766), .A2(n34309), .ZN(n14156) );
  NOR3_X2 U13457 ( .A1(n16679), .A2(n16678), .A3(n908), .ZN(n11543) );
  NOR2_X2 U2682 ( .A1(n33375), .A2(n5250), .ZN(n33630) );
  NAND2_X2 U9353 ( .A1(n43561), .A2(n42619), .ZN(n42095) );
  INV_X2 U10350 ( .I(n35653), .ZN(n9028) );
  NAND2_X2 U3103 ( .A1(n17496), .A2(n19830), .ZN(n20315) );
  OAI21_X2 U37202 ( .A1(n19305), .A2(n64061), .B(n63098), .ZN(n22319) );
  INV_X2 U8632 ( .I(n11250), .ZN(n19305) );
  NOR3_X2 U53664 ( .A1(n48807), .A2(n48806), .A3(n48805), .ZN(n48816) );
  INV_X2 U10603 ( .I(n28200), .ZN(n29670) );
  AOI22_X2 U55730 ( .A1(n54265), .A2(n15923), .B1(n54212), .B2(n54211), .ZN(
        n54217) );
  INV_X2 U10829 ( .I(n8459), .ZN(n49370) );
  NOR2_X2 U822 ( .A1(n49089), .A2(n57473), .ZN(n8459) );
  INV_X2 U10242 ( .I(n5233), .ZN(n34488) );
  NAND3_X2 U11763 ( .A1(n27792), .A2(n28949), .A3(n28945), .ZN(n15529) );
  AOI21_X2 U13802 ( .A1(n29840), .A2(n7979), .B(n28735), .ZN(n25399) );
  OR2_X2 U12084 ( .A1(n59604), .A2(n11329), .Z(n27674) );
  INV_X1 U514 ( .I(n63038), .ZN(n51457) );
  BUF_X2 U11732 ( .I(n31984), .Z(n5489) );
  NAND2_X2 U758 ( .A1(n48977), .A2(n22756), .ZN(n49844) );
  INV_X2 U3435 ( .I(n9556), .ZN(n13955) );
  INV_X2 U2444 ( .I(n35990), .ZN(n37046) );
  INV_X2 U2778 ( .I(n24485), .ZN(n13068) );
  NOR3_X2 U35599 ( .A1(n12074), .A2(n55270), .A3(n54996), .ZN(n54835) );
  AOI21_X1 U25032 ( .A1(n6754), .A2(n37062), .B(n6581), .ZN(n5337) );
  OAI21_X2 U11088 ( .A1(n42078), .A2(n42077), .B(n12073), .ZN(n6451) );
  NOR2_X2 U1276 ( .A1(n6417), .A2(n15697), .ZN(n3080) );
  INV_X2 U1659 ( .I(n43014), .ZN(n42314) );
  NOR2_X2 U467 ( .A1(n54053), .A2(n53916), .ZN(n53409) );
  NOR3_X2 U1171 ( .A1(n22391), .A2(n59922), .A3(n46049), .ZN(n9064) );
  BUF_X4 U14589 ( .I(n11557), .Z(n20985) );
  INV_X2 U46183 ( .I(n31311), .ZN(n38459) );
  INV_X2 U8866 ( .I(n12354), .ZN(n12405) );
  NOR2_X2 U2942 ( .A1(n9426), .A2(n23317), .ZN(n28773) );
  INV_X2 U11339 ( .I(n40995), .ZN(n18706) );
  NAND4_X2 U9189 ( .A1(n49460), .A2(n5947), .A3(n48395), .A4(n49152), .ZN(
        n8581) );
  BUF_X2 U40963 ( .I(Key[169]), .Z(n51569) );
  NOR2_X2 U1771 ( .A1(n21966), .A2(n21965), .ZN(n6601) );
  NAND2_X2 U1855 ( .A1(n25511), .A2(n4581), .ZN(n40107) );
  NAND2_X2 U9573 ( .A1(n34604), .A2(n20443), .ZN(n33419) );
  INV_X4 U21932 ( .I(n13029), .ZN(n6957) );
  AOI22_X2 U35423 ( .A1(n26812), .A2(n58971), .B1(n28551), .B2(n26810), .ZN(
        n23598) );
  OAI22_X2 U35069 ( .A1(n60543), .A2(n27274), .B1(n28548), .B2(n22351), .ZN(
        n26812) );
  AOI21_X2 U19116 ( .A1(n7087), .A2(n26840), .B(n26839), .ZN(n26842) );
  NOR2_X2 U38259 ( .A1(n48427), .A2(n48811), .ZN(n48809) );
  NAND2_X2 U2323 ( .A1(n2483), .A2(n1793), .ZN(n37055) );
  INV_X1 U16253 ( .I(n14323), .ZN(n1657) );
  INV_X2 U3288 ( .I(n10236), .ZN(n28860) );
  NOR2_X2 U4274 ( .A1(n40924), .A2(n40470), .ZN(n40248) );
  NOR2_X2 U8093 ( .A1(n34308), .A2(n19005), .ZN(n15830) );
  NOR3_X2 U2891 ( .A1(n20990), .A2(n30178), .A3(n30179), .ZN(n17491) );
  INV_X2 U2617 ( .I(n34622), .ZN(n34628) );
  NOR2_X2 U1087 ( .A1(n48163), .A2(n48511), .ZN(n48507) );
  NAND3_X2 U11595 ( .A1(n3559), .A2(n33965), .A3(n61809), .ZN(n25194) );
  NAND2_X2 U2985 ( .A1(n23799), .A2(n59046), .ZN(n30313) );
  BUF_X2 U3590 ( .I(n56282), .Z(n187) );
  INV_X2 U33599 ( .I(n19438), .ZN(n40094) );
  INV_X8 U3100 ( .I(n16971), .ZN(n30455) );
  NOR4_X2 U4345 ( .A1(n28234), .A2(n14581), .A3(n14582), .A4(n10729), .ZN(
        n6018) );
  NOR3_X2 U6996 ( .A1(n5982), .A2(n28031), .A3(n28039), .ZN(n10729) );
  NAND2_X2 U9003 ( .A1(n17633), .A2(n17522), .ZN(n17634) );
  INV_X2 U9608 ( .I(n31984), .ZN(n23461) );
  INV_X2 U587 ( .I(n49817), .ZN(n51933) );
  INV_X4 U895 ( .I(n24966), .ZN(n19144) );
  NAND3_X1 U3519 ( .A1(n12162), .A2(n30053), .A3(n16630), .ZN(n12161) );
  NAND3_X2 U53162 ( .A1(n47090), .A2(n47089), .A3(n58620), .ZN(n47094) );
  NAND2_X2 U10970 ( .A1(n48475), .A2(n47091), .ZN(n47088) );
  NOR2_X2 U18310 ( .A1(n24036), .A2(n34166), .ZN(n34175) );
  INV_X4 U23129 ( .I(n52476), .ZN(n5569) );
  NAND2_X2 U9674 ( .A1(n9476), .A2(n29778), .ZN(n28949) );
  NAND2_X2 U28162 ( .A1(n1218), .A2(n7426), .ZN(n30754) );
  NOR2_X2 U2943 ( .A1(n30752), .A2(n25052), .ZN(n31217) );
  BUF_X2 U5700 ( .I(n14714), .Z(n13982) );
  INV_X2 U1201 ( .I(n47186), .ZN(n48530) );
  NAND2_X2 U4081 ( .A1(n57199), .A2(n5531), .ZN(n40602) );
  BUF_X8 U41542 ( .I(n1218), .Z(n23799) );
  NAND2_X2 U4110 ( .A1(n6540), .A2(n12521), .ZN(n18877) );
  NOR2_X2 U693 ( .A1(n49602), .A2(n8129), .ZN(n49316) );
  INV_X2 U3313 ( .I(n27698), .ZN(n29610) );
  NAND2_X2 U35114 ( .A1(n43548), .A2(n59682), .ZN(n43627) );
  INV_X4 U2670 ( .I(n34308), .ZN(n34771) );
  INV_X2 U12356 ( .I(n47068), .ZN(n25451) );
  BUF_X2 U14280 ( .I(n29180), .Z(n23608) );
  BUF_X4 U24709 ( .I(n55099), .Z(n5051) );
  AOI22_X2 U4098 ( .A1(n35295), .A2(n21751), .B1(n35296), .B2(n35294), .ZN(
        n20108) );
  AOI21_X2 U40050 ( .A1(n28599), .A2(n59903), .B(n28598), .ZN(n19788) );
  NOR2_X2 U38904 ( .A1(n28127), .A2(n18062), .ZN(n28825) );
  NOR3_X2 U43871 ( .A1(n40667), .A2(n709), .A3(n10126), .ZN(n41171) );
  NAND2_X2 U1212 ( .A1(n44770), .A2(n26145), .ZN(n47487) );
  NAND3_X2 U8535 ( .A1(n19851), .A2(n49439), .A3(n49572), .ZN(n19850) );
  NAND3_X2 U50220 ( .A1(n39148), .A2(n40494), .A3(n9915), .ZN(n39149) );
  INV_X1 U38867 ( .I(n60894), .ZN(n28136) );
  NOR4_X2 U44415 ( .A1(n26950), .A2(n29632), .A3(n26949), .A4(n28838), .ZN(
        n26956) );
  NOR3_X2 U10212 ( .A1(n25753), .A2(n34098), .A3(n25752), .ZN(n25751) );
  INV_X2 U396 ( .I(n56637), .ZN(n52721) );
  OAI21_X2 U10014 ( .A1(n9163), .A2(n9162), .B(n19346), .ZN(n43719) );
  INV_X2 U418 ( .I(n12692), .ZN(n20740) );
  INV_X2 U5735 ( .I(n40591), .ZN(n1272) );
  AND2_X2 U1218 ( .A1(n24475), .A2(n45218), .Z(n838) );
  NOR2_X2 U2671 ( .A1(n25849), .A2(n64603), .ZN(n33960) );
  NAND3_X1 U12497 ( .A1(n47008), .A2(n57205), .A3(n47007), .ZN(n47009) );
  NOR2_X2 U28542 ( .A1(n12898), .A2(n14050), .ZN(n12414) );
  AOI21_X2 U2204 ( .A1(n35552), .A2(n9513), .B(n10730), .ZN(n13303) );
  NAND2_X2 U4556 ( .A1(n5233), .A2(n35554), .ZN(n10730) );
  NAND2_X2 U3374 ( .A1(n11655), .A2(n24197), .ZN(n29697) );
  INV_X2 U2813 ( .I(n19282), .ZN(n12781) );
  NAND2_X2 U7055 ( .A1(n33737), .A2(n21196), .ZN(n34731) );
  BUF_X4 U2809 ( .I(n24064), .Z(n14818) );
  NOR2_X2 U7050 ( .A1(n33600), .A2(n10682), .ZN(n35690) );
  NOR2_X2 U9745 ( .A1(n29284), .A2(n29283), .ZN(n28838) );
  NOR3_X2 U12265 ( .A1(n21893), .A2(n56624), .A3(n1286), .ZN(n8828) );
  NAND2_X2 U93 ( .A1(n53527), .A2(n53506), .ZN(n53497) );
  OAI21_X2 U2188 ( .A1(n34827), .A2(n35583), .B(n34464), .ZN(n37613) );
  OR2_X2 U16550 ( .A1(n41625), .A2(n41632), .Z(n4347) );
  NOR2_X2 U897 ( .A1(n49410), .A2(n11314), .ZN(n10872) );
  NAND3_X2 U7127 ( .A1(n22348), .A2(n40197), .A3(n40198), .ZN(n26160) );
  BUF_X4 U19377 ( .I(n30580), .Z(n23955) );
  INV_X4 U20443 ( .I(n49379), .ZN(n49432) );
  INV_X1 U41522 ( .I(n48527), .ZN(n50308) );
  NOR2_X2 U20575 ( .A1(n19302), .A2(n2357), .ZN(n45172) );
  NAND2_X2 U7690 ( .A1(n3090), .A2(n12735), .ZN(n2814) );
  CLKBUF_X4 U4638 ( .I(n12051), .Z(n65) );
  NOR2_X2 U1812 ( .A1(n64672), .A2(n18441), .ZN(n39516) );
  INV_X4 U25070 ( .I(n5377), .ZN(n32892) );
  NOR2_X2 U2564 ( .A1(n30467), .A2(n16869), .ZN(n34992) );
  INV_X4 U9691 ( .I(n30547), .ZN(n15205) );
  NOR2_X2 U15569 ( .A1(n18769), .A2(n47916), .ZN(n47917) );
  NOR2_X2 U3076 ( .A1(n16279), .A2(n19598), .ZN(n30704) );
  INV_X4 U10198 ( .I(n2355), .ZN(n39299) );
  NOR2_X2 U25017 ( .A1(n36442), .A2(n36443), .ZN(n35588) );
  AOI21_X2 U11982 ( .A1(n28648), .A2(n29695), .B(n28639), .ZN(n27683) );
  INV_X2 U19286 ( .I(n24467), .ZN(n10888) );
  INV_X2 U34404 ( .I(n15078), .ZN(n40850) );
  NOR2_X2 U43957 ( .A1(n28039), .A2(n61177), .ZN(n27103) );
  NAND3_X2 U4426 ( .A1(n48115), .A2(n49859), .A3(n49864), .ZN(n25352) );
  NAND2_X2 U51382 ( .A1(n42567), .A2(n42566), .ZN(n42903) );
  INV_X4 U13666 ( .I(n6914), .ZN(n35674) );
  INV_X2 U47209 ( .I(n33481), .ZN(n34950) );
  NOR2_X2 U2732 ( .A1(n1545), .A2(n22185), .ZN(n33481) );
  INV_X1 U41068 ( .I(n49075), .ZN(n49833) );
  NAND4_X2 U2563 ( .A1(n33345), .A2(n7273), .A3(n33568), .A4(n33561), .ZN(
        n19095) );
  NOR2_X2 U3077 ( .A1(n23446), .A2(n58829), .ZN(n23502) );
  OR2_X2 U1527 ( .A1(n43995), .A2(n22716), .Z(n43256) );
  NAND3_X2 U14052 ( .A1(n27225), .A2(n24785), .A3(n24784), .ZN(n4941) );
  NAND2_X2 U10329 ( .A1(n34787), .A2(n34797), .ZN(n35013) );
  INV_X2 U3345 ( .I(n22352), .ZN(n29178) );
  INV_X4 U41365 ( .I(n37699), .ZN(n24859) );
  NAND2_X2 U18237 ( .A1(n35246), .A2(n35245), .ZN(n35920) );
  INV_X4 U29686 ( .I(n14448), .ZN(n13258) );
  INV_X1 U2927 ( .I(n4037), .ZN(n30393) );
  INV_X2 U22087 ( .I(n65160), .ZN(n36427) );
  INV_X2 U3234 ( .I(n60020), .ZN(n28237) );
  OAI21_X2 U2498 ( .A1(n34509), .A2(n34991), .B(n34995), .ZN(n3511) );
  NOR3_X2 U2514 ( .A1(n35704), .A2(n12937), .A3(n35751), .ZN(n12936) );
  INV_X2 U10137 ( .I(n9189), .ZN(n1504) );
  INV_X2 U32849 ( .I(n12810), .ZN(n56559) );
  NAND2_X2 U7309 ( .A1(n12601), .A2(n50948), .ZN(n12602) );
  AOI21_X2 U50214 ( .A1(n39142), .A2(n59179), .B(n40653), .ZN(n39156) );
  NAND2_X1 U27384 ( .A1(n7421), .A2(n12630), .ZN(n53243) );
  NAND2_X2 U2215 ( .A1(n36987), .A2(n37227), .ZN(n37230) );
  OR3_X2 U5845 ( .A1(n40421), .A2(n39821), .A3(n41122), .Z(n41381) );
  INV_X2 U10501 ( .I(n1319), .ZN(n24206) );
  INV_X2 U1757 ( .I(n42636), .ZN(n43383) );
  NAND2_X2 U50745 ( .A1(n18741), .A2(n40592), .ZN(n41084) );
  NAND2_X2 U2740 ( .A1(n34324), .A2(n35816), .ZN(n35305) );
  AOI22_X2 U9413 ( .A1(n4489), .A2(n40291), .B1(n14018), .B2(n22746), .ZN(
        n40031) );
  INV_X2 U11129 ( .I(n43302), .ZN(n25600) );
  NOR2_X2 U35188 ( .A1(n21655), .A2(n21330), .ZN(n52705) );
  NAND2_X2 U10917 ( .A1(n47405), .A2(n47669), .ZN(n47869) );
  INV_X2 U10951 ( .I(n61909), .ZN(n47405) );
  BUF_X4 U20485 ( .I(n8443), .Z(n2269) );
  NOR2_X2 U3390 ( .A1(n29120), .A2(n22714), .ZN(n29127) );
  NAND2_X2 U34982 ( .A1(n34335), .A2(n64812), .ZN(n21538) );
  INV_X2 U408 ( .I(n56591), .ZN(n56255) );
  NAND2_X2 U1794 ( .A1(n11016), .A2(n20974), .ZN(n40558) );
  NOR2_X2 U3371 ( .A1(n6345), .A2(n6370), .ZN(n19581) );
  NAND2_X2 U2991 ( .A1(n15407), .A2(n31055), .ZN(n15333) );
  INV_X2 U34785 ( .I(n18335), .ZN(n56565) );
  AOI21_X2 U6840 ( .A1(n45891), .A2(n60848), .B(n64869), .ZN(n695) );
  NAND2_X2 U4118 ( .A1(n18969), .A2(n17030), .ZN(n37278) );
  BUF_X4 U4977 ( .I(n33661), .Z(n157) );
  NOR2_X2 U7057 ( .A1(n3467), .A2(n9687), .ZN(n34667) );
  AOI21_X1 U30346 ( .A1(n49796), .A2(n49797), .B(n49795), .ZN(n49798) );
  NAND2_X2 U14056 ( .A1(n19700), .A2(n6293), .ZN(n10206) );
  OAI21_X2 U1410 ( .A1(n43133), .A2(n43134), .B(n12502), .ZN(n25495) );
  INV_X2 U1525 ( .I(n42572), .ZN(n42567) );
  NAND2_X2 U9484 ( .A1(n18857), .A2(n37044), .ZN(n37960) );
  OAI21_X2 U50785 ( .A1(n41174), .A2(n40484), .B(n40488), .ZN(n40485) );
  NAND2_X2 U18405 ( .A1(n19570), .A2(n34423), .ZN(n35327) );
  NAND2_X2 U10941 ( .A1(n25728), .A2(n48246), .ZN(n4620) );
  NAND4_X2 U7227 ( .A1(n20162), .A2(n3364), .A3(n48659), .A4(n48248), .ZN(
        n25728) );
  NOR2_X2 U2008 ( .A1(n1745), .A2(n41132), .ZN(n40833) );
  NAND3_X2 U4019 ( .A1(n58645), .A2(n64006), .A3(n49674), .ZN(n49091) );
  OAI22_X2 U13355 ( .A1(n23739), .A2(n34484), .B1(n35426), .B2(n36943), .ZN(
        n36893) );
  INV_X2 U791 ( .I(n49365), .ZN(n49099) );
  OAI21_X2 U36257 ( .A1(n56986), .A2(n52689), .B(n52688), .ZN(n52690) );
  INV_X2 U12994 ( .I(n42985), .ZN(n1503) );
  NAND2_X2 U35170 ( .A1(n1781), .A2(n36959), .ZN(n36279) );
  INV_X1 U10825 ( .I(n2608), .ZN(n49203) );
  NOR2_X2 U51336 ( .A1(n42376), .A2(n42703), .ZN(n42378) );
  NAND2_X2 U12060 ( .A1(n19359), .A2(n64337), .ZN(n26805) );
  BUF_X4 U44090 ( .I(Key[85]), .Z(n54888) );
  INV_X4 U29754 ( .I(n36533), .ZN(n20530) );
  NAND2_X2 U9906 ( .A1(n1468), .A2(n20458), .ZN(n17816) );
  OR2_X1 U15831 ( .A1(n45629), .A2(n46064), .Z(n10078) );
  INV_X2 U6988 ( .I(n28609), .ZN(n28453) );
  INV_X2 U5370 ( .I(n248), .ZN(n2104) );
  INV_X2 U887 ( .I(n19544), .ZN(n47972) );
  INV_X4 U30364 ( .I(n1664), .ZN(n47876) );
  INV_X4 U19296 ( .I(n5070), .ZN(n5192) );
  NOR2_X2 U47690 ( .A1(n33112), .A2(n33375), .ZN(n33634) );
  BUF_X4 U14297 ( .I(Key[59]), .Z(n54208) );
  NOR2_X2 U2638 ( .A1(n16402), .A2(n60669), .ZN(n35255) );
  NOR2_X2 U2519 ( .A1(n13818), .A2(n57423), .ZN(n34966) );
  INV_X2 U19812 ( .I(n29643), .ZN(n6370) );
  NAND2_X2 U2370 ( .A1(n36831), .A2(n6540), .ZN(n36835) );
  NOR2_X2 U2993 ( .A1(n30492), .A2(n5070), .ZN(n30490) );
  INV_X2 U2816 ( .I(n7079), .ZN(n25443) );
  NAND3_X2 U9569 ( .A1(n35294), .A2(n21730), .A3(n34335), .ZN(n34755) );
  NAND2_X2 U50228 ( .A1(n39164), .A2(n40470), .ZN(n40929) );
  NAND3_X2 U1486 ( .A1(n10196), .A2(n3855), .A3(n42174), .ZN(n3852) );
  NAND2_X2 U337 ( .A1(n1596), .A2(n56374), .ZN(n24729) );
  NOR2_X2 U20245 ( .A1(n24712), .A2(n364), .ZN(n28688) );
  INV_X2 U9014 ( .I(n12070), .ZN(n13097) );
  INV_X1 U9857 ( .I(n51557), .ZN(n56371) );
  INV_X2 U23036 ( .I(n16907), .ZN(n24933) );
  AOI22_X2 U18344 ( .A1(n33100), .A2(n33559), .B1(n11024), .B2(n33099), .ZN(
        n33107) );
  INV_X2 U7654 ( .I(n39604), .ZN(n22638) );
  NAND2_X2 U768 ( .A1(n14561), .A2(n6633), .ZN(n7289) );
  NAND2_X2 U31987 ( .A1(n11793), .A2(n11790), .ZN(n36158) );
  BUF_X4 U8148 ( .I(n22107), .Z(n1208) );
  NAND4_X2 U10083 ( .A1(n40975), .A2(n39063), .A3(n39137), .A4(n39062), .ZN(
        n39064) );
  NAND2_X2 U2950 ( .A1(n875), .A2(n4999), .ZN(n30363) );
  INV_X4 U14248 ( .I(n5982), .ZN(n21301) );
  NOR3_X2 U16600 ( .A1(n5365), .A2(n4409), .A3(n5367), .ZN(n41622) );
  NOR2_X2 U847 ( .A1(n49411), .A2(n10872), .ZN(n48956) );
  NAND2_X2 U10348 ( .A1(n1537), .A2(n33756), .ZN(n34946) );
  INV_X2 U1581 ( .I(n24360), .ZN(n23811) );
  AOI22_X2 U35961 ( .A1(n42074), .A2(n42407), .B1(n19793), .B2(n42404), .ZN(
        n42075) );
  BUF_X4 U9079 ( .I(Key[144]), .Z(n56143) );
  NOR2_X2 U33932 ( .A1(n23732), .A2(n28119), .ZN(n14433) );
  BUF_X4 U9442 ( .I(n38021), .Z(n16962) );
  INV_X4 U41342 ( .I(n21831), .ZN(n26092) );
  INV_X8 U28161 ( .I(n1218), .ZN(n30752) );
  NAND2_X1 U36910 ( .A1(n17429), .A2(n20526), .ZN(n42311) );
  INV_X2 U383 ( .I(n54657), .ZN(n18629) );
  NOR2_X2 U11822 ( .A1(n30753), .A2(n61215), .ZN(n30669) );
  NOR2_X2 U8597 ( .A1(n47327), .A2(n46919), .ZN(n21246) );
  NAND2_X2 U13531 ( .A1(n33802), .A2(n33584), .ZN(n35249) );
  NAND2_X2 U13282 ( .A1(n36765), .A2(n35414), .ZN(n18705) );
  NAND3_X2 U7365 ( .A1(n55611), .A2(n55650), .A3(n19020), .ZN(n19845) );
  NAND2_X2 U19443 ( .A1(n23880), .A2(n19912), .ZN(n19911) );
  NAND4_X1 U55166 ( .A1(n52757), .A2(n52843), .A3(n53603), .A4(n53608), .ZN(
        n52758) );
  NAND4_X2 U50805 ( .A1(n40536), .A2(n40535), .A3(n40534), .A4(n40533), .ZN(
        n40537) );
  NAND2_X2 U6974 ( .A1(n28667), .A2(n28666), .ZN(n12636) );
  INV_X4 U2690 ( .I(n15028), .ZN(n1535) );
  INV_X2 U2815 ( .I(n8667), .ZN(n22146) );
  NAND4_X2 U4943 ( .A1(n147), .A2(n21216), .A3(n14291), .A4(n21181), .ZN(
        n14290) );
  NAND2_X1 U30864 ( .A1(n22510), .A2(n52703), .ZN(n52712) );
  NAND2_X2 U2525 ( .A1(n35003), .A2(n24799), .ZN(n32958) );
  INV_X1 U464 ( .I(n52845), .ZN(n19062) );
  INV_X1 U12267 ( .I(n53605), .ZN(n53380) );
  NAND2_X2 U10458 ( .A1(n6609), .A2(n5070), .ZN(n28902) );
  INV_X2 U7297 ( .I(n23414), .ZN(n50334) );
  AOI21_X2 U18292 ( .A1(n31730), .A2(n31729), .B(n17828), .ZN(n17827) );
  OAI22_X2 U35033 ( .A1(n17377), .A2(n60700), .B1(n34126), .B2(n34127), .ZN(
        n17828) );
  BUF_X4 U42190 ( .I(n30943), .Z(n34973) );
  INV_X2 U13995 ( .I(n14522), .ZN(n16764) );
  NOR2_X2 U29733 ( .A1(n6440), .A2(n36533), .ZN(n36053) );
  NAND2_X2 U12983 ( .A1(n41094), .A2(n42266), .ZN(n22479) );
  OR2_X1 U8323 ( .A1(n16869), .A2(n33486), .Z(n34071) );
  NAND2_X2 U27154 ( .A1(n7297), .A2(n10412), .ZN(n10411) );
  INV_X2 U1766 ( .I(n62353), .ZN(n3785) );
  BUF_X4 U9701 ( .I(n23569), .Z(n1352) );
  BUF_X4 U1255 ( .I(n13029), .Z(n3364) );
  INV_X4 U32520 ( .I(n20391), .ZN(n31208) );
  BUF_X4 U19913 ( .I(Key[61]), .Z(n54219) );
  INV_X4 U2681 ( .I(n15588), .ZN(n32951) );
  INV_X2 U1381 ( .I(n19155), .ZN(n5630) );
  OAI21_X2 U17377 ( .A1(n2760), .A2(n63119), .B(n41084), .ZN(n41085) );
  INV_X2 U3054 ( .I(n14276), .ZN(n31117) );
  NAND2_X2 U4170 ( .A1(n15157), .A2(n5145), .ZN(n3807) );
  BUF_X4 U14517 ( .I(n52762), .Z(n9731) );
  INV_X2 U349 ( .I(n54943), .ZN(n54611) );
  NOR2_X2 U8046 ( .A1(n1393), .A2(n9672), .ZN(n42376) );
  AOI22_X2 U48620 ( .A1(n35859), .A2(n35858), .B1(n35857), .B2(n35856), .ZN(
        n35868) );
  AOI21_X2 U36498 ( .A1(n12004), .A2(n1417), .B(n65234), .ZN(n35858) );
  INV_X2 U2817 ( .I(n21025), .ZN(n25822) );
  BUF_X4 U1949 ( .I(n24389), .Z(n40091) );
  INV_X2 U3012 ( .I(n8522), .ZN(n3901) );
  INV_X1 U36139 ( .I(n35013), .ZN(n35014) );
  INV_X2 U6969 ( .I(n29626), .ZN(n29281) );
  OAI21_X2 U55184 ( .A1(n61147), .A2(n62664), .B(n53024), .ZN(n52780) );
  NAND2_X1 U11629 ( .A1(n64706), .A2(n64708), .ZN(n35022) );
  INV_X1 U27630 ( .I(n7564), .ZN(n10908) );
  INV_X2 U11856 ( .I(n30055), .ZN(n30054) );
  NAND2_X2 U37179 ( .A1(n617), .A2(n15693), .ZN(n48875) );
  NAND2_X2 U9697 ( .A1(n30743), .A2(n58273), .ZN(n18880) );
  NOR3_X2 U3174 ( .A1(n23964), .A2(n27488), .A3(n27489), .ZN(n188) );
  NOR3_X2 U27766 ( .A1(n7683), .A2(n31049), .A3(n30177), .ZN(n30178) );
  INV_X2 U6411 ( .I(n62353), .ZN(n43380) );
  INV_X1 U956 ( .I(n10636), .ZN(n25091) );
  NAND2_X2 U8229 ( .A1(n5833), .A2(n6241), .ZN(n6497) );
  NAND2_X2 U11259 ( .A1(n14558), .A2(n40228), .ZN(n3896) );
  OR2_X2 U3511 ( .A1(n10353), .A2(n6027), .Z(n5961) );
  INV_X2 U3232 ( .I(n28002), .ZN(n29105) );
  AOI21_X2 U11815 ( .A1(n29266), .A2(n29580), .B(n10129), .ZN(n2098) );
  BUF_X2 U1241 ( .I(n1265), .Z(n8820) );
  INV_X4 U2739 ( .I(n22185), .ZN(n1345) );
  INV_X1 U10131 ( .I(n42252), .ZN(n42245) );
  INV_X4 U38168 ( .I(n16938), .ZN(n21755) );
  NOR2_X1 U23641 ( .A1(n42866), .A2(n4574), .ZN(n42881) );
  INV_X4 U10864 ( .I(n1224), .ZN(n1377) );
  NAND3_X2 U22121 ( .A1(n29069), .A2(n18356), .A3(n29068), .ZN(n3533) );
  INV_X4 U10360 ( .I(n20978), .ZN(n6760) );
  NAND2_X2 U2218 ( .A1(n36512), .A2(n36511), .ZN(n36585) );
  BUF_X2 U19811 ( .I(n29282), .Z(n23732) );
  INV_X2 U3353 ( .I(n28311), .ZN(n24878) );
  INV_X4 U2755 ( .I(n30895), .ZN(n3467) );
  NAND2_X2 U44362 ( .A1(n28675), .A2(n29609), .ZN(n28673) );
  NOR2_X2 U2319 ( .A1(n37050), .A2(n35096), .ZN(n35995) );
  NOR2_X2 U12061 ( .A1(n22312), .A2(n26791), .ZN(n28611) );
  INV_X4 U3157 ( .I(n25698), .ZN(n22014) );
  NAND2_X2 U2520 ( .A1(n31528), .A2(n7849), .ZN(n33417) );
  AOI22_X2 U13279 ( .A1(n35390), .A2(n35389), .B1(n35388), .B2(n36040), .ZN(
        n35393) );
  INV_X4 U3444 ( .I(n815), .ZN(n29608) );
  AOI21_X2 U9121 ( .A1(n52830), .A2(n57029), .B(n52829), .ZN(n52834) );
  OAI21_X2 U8503 ( .A1(n57019), .A2(n23102), .B(n53220), .ZN(n52830) );
  INV_X2 U138 ( .I(n55595), .ZN(n55592) );
  INV_X4 U8351 ( .I(n1562), .ZN(n8218) );
  NAND2_X2 U1678 ( .A1(n4275), .A2(n42019), .ZN(n43395) );
  INV_X1 U5463 ( .I(n34666), .ZN(n34677) );
  CLKBUF_X4 U7434 ( .I(n21014), .Z(n1559) );
  CLKBUF_X4 U14288 ( .I(n28446), .Z(n14019) );
  NOR2_X2 U9658 ( .A1(n30501), .A2(n31241), .ZN(n30887) );
  NAND2_X2 U10239 ( .A1(n34365), .A2(n3622), .ZN(n36772) );
  NAND4_X2 U3029 ( .A1(n30752), .A2(n59046), .A3(n19929), .A4(n31224), .ZN(
        n30764) );
  INV_X4 U14277 ( .I(n29370), .ZN(n23479) );
  BUF_X4 U4442 ( .I(n35341), .Z(n22528) );
  INV_X2 U82 ( .I(n55556), .ZN(n55574) );
  BUF_X2 U16302 ( .I(n45074), .Z(n47314) );
  NAND2_X2 U31004 ( .A1(n28067), .A2(n24853), .ZN(n27037) );
  BUF_X4 U5365 ( .I(n33697), .Z(n7273) );
  INV_X4 U27780 ( .I(n26126), .ZN(n10236) );
  INV_X2 U10185 ( .I(n39502), .ZN(n15139) );
  INV_X2 U8965 ( .I(n21838), .ZN(n5933) );
  INV_X4 U7857 ( .I(n25857), .ZN(n48845) );
  BUF_X2 U14600 ( .I(n53727), .Z(n9616) );
  NAND2_X2 U7026 ( .A1(n8891), .A2(n30124), .ZN(n30525) );
  OAI21_X2 U15514 ( .A1(n48580), .A2(n49650), .B(n62035), .ZN(n9501) );
  INV_X4 U931 ( .I(n50360), .ZN(n24134) );
  NAND2_X2 U10451 ( .A1(n31174), .A2(n29905), .ZN(n30858) );
  NAND3_X2 U18419 ( .A1(n35248), .A2(n22909), .A3(n35249), .ZN(n19661) );
  NOR2_X2 U9299 ( .A1(n41728), .A2(n14240), .ZN(n13180) );
  INV_X2 U37748 ( .I(n20812), .ZN(n36748) );
  INV_X4 U31197 ( .I(n23812), .ZN(n35688) );
  INV_X2 U8116 ( .I(n19085), .ZN(n13504) );
  AOI21_X2 U10249 ( .A1(n36484), .A2(n36483), .B(n19539), .ZN(n36486) );
  NOR2_X2 U36537 ( .A1(n36206), .A2(n36205), .ZN(n23333) );
  BUF_X2 U11875 ( .I(n5242), .Z(n3180) );
  CLKBUF_X4 U6652 ( .I(n13826), .Z(n9548) );
  INV_X2 U6993 ( .I(n29727), .ZN(n28986) );
  AOI21_X1 U48637 ( .A1(n6984), .A2(n35920), .B(n35919), .ZN(n35921) );
  INV_X4 U2449 ( .I(n1235), .ZN(n8223) );
  NAND2_X2 U740 ( .A1(n48680), .A2(n22157), .ZN(n48892) );
  NOR2_X2 U8374 ( .A1(n6440), .A2(n36538), .ZN(n35452) );
  INV_X2 U13726 ( .I(n32461), .ZN(n9205) );
  NAND3_X2 U2191 ( .A1(n17912), .A2(n4450), .A3(n4449), .ZN(n16627) );
  BUF_X4 U24150 ( .I(n6410), .Z(n6411) );
  AOI21_X2 U17860 ( .A1(n4679), .A2(n36813), .B(n25771), .ZN(n25770) );
  INV_X1 U4248 ( .I(n25972), .ZN(n32794) );
  NOR2_X2 U998 ( .A1(n1636), .A2(n49929), .ZN(n49922) );
  NOR2_X2 U16961 ( .A1(n13419), .A2(n39828), .ZN(n6102) );
  OAI21_X2 U12527 ( .A1(n46062), .A2(n60893), .B(n21245), .ZN(n21552) );
  NAND3_X2 U19304 ( .A1(n8182), .A2(n6316), .A3(n31277), .ZN(n29919) );
  NAND4_X1 U38757 ( .A1(n28136), .A2(n17993), .A3(n29287), .A4(n19290), .ZN(
        n17992) );
  NAND2_X2 U76 ( .A1(n54001), .A2(n53992), .ZN(n53953) );
  NAND2_X2 U2552 ( .A1(n23313), .A2(n23812), .ZN(n33012) );
  NOR2_X2 U11598 ( .A1(n33676), .A2(n17283), .ZN(n12737) );
  NAND2_X2 U2553 ( .A1(n19435), .A2(n17759), .ZN(n33676) );
  BUF_X4 U7426 ( .I(n26414), .Z(n28510) );
  NAND3_X1 U33907 ( .A1(n28782), .A2(n30231), .A3(n14393), .ZN(n14392) );
  NAND2_X2 U16827 ( .A1(n43205), .A2(n22695), .ZN(n10937) );
  NAND2_X1 U29380 ( .A1(n55008), .A2(n9418), .ZN(n55009) );
  NOR2_X2 U2258 ( .A1(n35916), .A2(n35917), .ZN(n19130) );
  NOR2_X2 U37178 ( .A1(n61513), .A2(n617), .ZN(n48869) );
  NAND2_X2 U9386 ( .A1(n42275), .A2(n1001), .ZN(n40820) );
  NAND2_X2 U4091 ( .A1(n5299), .A2(n45075), .ZN(n47316) );
  OR2_X2 U19355 ( .A1(n7127), .A2(n1192), .Z(n27743) );
  INV_X2 U2093 ( .I(n12887), .ZN(n38023) );
  NOR2_X2 U3384 ( .A1(n23469), .A2(n14834), .ZN(n27056) );
  NAND2_X2 U9507 ( .A1(n63583), .A2(n35452), .ZN(n36551) );
  INV_X2 U33382 ( .I(n15047), .ZN(n26150) );
  NAND2_X2 U2278 ( .A1(n36512), .A2(n36508), .ZN(n37368) );
  INV_X2 U10184 ( .I(n60587), .ZN(n12735) );
  INV_X2 U44752 ( .I(n27717), .ZN(n28514) );
  NAND2_X2 U7090 ( .A1(n35604), .A2(n1311), .ZN(n36263) );
  INV_X2 U551 ( .I(n10969), .ZN(n10968) );
  OAI22_X2 U41317 ( .A1(n34264), .A2(n35294), .B1(n34265), .B2(n59676), .ZN(
        n34266) );
  INV_X1 U18770 ( .I(n32556), .ZN(n4949) );
  NAND2_X2 U7097 ( .A1(n7028), .A2(n35416), .ZN(n36776) );
  NAND2_X2 U35561 ( .A1(n49410), .A2(n10874), .ZN(n48962) );
  NAND3_X2 U35479 ( .A1(n16526), .A2(n38346), .A3(n8017), .ZN(n37595) );
  BUF_X4 U37780 ( .I(Key[122]), .Z(n55610) );
  NAND2_X2 U37046 ( .A1(n47250), .A2(n65145), .ZN(n46891) );
  BUF_X2 U9161 ( .I(n53222), .Z(n23701) );
  NAND4_X1 U27248 ( .A1(n7348), .A2(n38351), .A3(n7720), .A4(n38350), .ZN(
        n38357) );
  BUF_X4 U14295 ( .I(Key[73]), .Z(n23306) );
  INV_X1 U1409 ( .I(n46547), .ZN(n8164) );
  INV_X2 U37162 ( .I(n48875), .ZN(n49397) );
  NAND2_X2 U11133 ( .A1(n19283), .A2(n42667), .ZN(n43253) );
  NOR2_X2 U16822 ( .A1(n42665), .A2(n65141), .ZN(n19283) );
  OAI21_X2 U18372 ( .A1(n11024), .A2(n33693), .B(n33097), .ZN(n33089) );
  NAND3_X2 U13490 ( .A1(n35682), .A2(n35684), .A3(n35683), .ZN(n4577) );
  INV_X4 U23143 ( .I(n21030), .ZN(n54307) );
  NAND4_X2 U8715 ( .A1(n40929), .A2(n40931), .A3(n40930), .A4(n60172), .ZN(
        n41512) );
  AOI21_X1 U27127 ( .A1(n21118), .A2(n21125), .B(n21120), .ZN(n21117) );
  INV_X2 U3072 ( .I(n28060), .ZN(n29988) );
  NOR3_X2 U8660 ( .A1(n9886), .A2(n7049), .A3(n15878), .ZN(n25438) );
  NAND2_X2 U1519 ( .A1(n2557), .A2(n11727), .ZN(n41325) );
  INV_X2 U10575 ( .I(n28321), .ZN(n3022) );
  NAND4_X2 U41935 ( .A1(n34271), .A2(n35300), .A3(n34733), .A4(n34270), .ZN(
        n34272) );
  OAI21_X2 U15927 ( .A1(n46108), .A2(n46107), .B(n48248), .ZN(n16520) );
  NAND2_X2 U1946 ( .A1(n40664), .A2(n41182), .ZN(n13909) );
  BUF_X2 U12118 ( .I(Key[166]), .Z(n56714) );
  BUF_X2 U37496 ( .I(n32828), .Z(n17199) );
  AOI21_X2 U35036 ( .A1(n20260), .A2(n23859), .B(n20259), .ZN(n20258) );
  INV_X4 U26393 ( .I(n6726), .ZN(n29295) );
  NAND2_X2 U8304 ( .A1(n46951), .A2(n6034), .ZN(n45506) );
  NAND2_X2 U12888 ( .A1(n14496), .A2(n23557), .ZN(n14408) );
  OR2_X2 U988 ( .A1(n19175), .A2(n17334), .Z(n49300) );
  AOI22_X2 U19493 ( .A1(n28474), .A2(n15986), .B1(n28473), .B2(n17688), .ZN(
        n28480) );
  NOR2_X2 U1279 ( .A1(n1387), .A2(n47874), .ZN(n47885) );
  NOR2_X2 U2059 ( .A1(n36648), .A2(n9215), .ZN(n39414) );
  NOR2_X2 U8437 ( .A1(n64183), .A2(n59637), .ZN(n41103) );
  INV_X2 U10334 ( .I(n34156), .ZN(n33683) );
  NOR2_X2 U39928 ( .A1(n16224), .A2(n19532), .ZN(n21622) );
  NAND2_X2 U10420 ( .A1(n29560), .A2(n27149), .ZN(n31128) );
  OAI21_X2 U12556 ( .A1(n15164), .A2(n15163), .B(n49862), .ZN(n18630) );
  INV_X2 U7259 ( .I(n47059), .ZN(n46261) );
  NAND2_X2 U2572 ( .A1(n18488), .A2(n35806), .ZN(n31841) );
  NOR3_X2 U14022 ( .A1(n15880), .A2(n19371), .A3(n26738), .ZN(n24442) );
  NOR2_X2 U17647 ( .A1(n949), .A2(n35978), .ZN(n5109) );
  INV_X4 U27353 ( .I(n56107), .ZN(n9567) );
  INV_X2 U36177 ( .I(n18598), .ZN(n25103) );
  NOR2_X2 U840 ( .A1(n18975), .A2(n49556), .ZN(n19866) );
  OAI21_X2 U48459 ( .A1(n1806), .A2(n1544), .B(n35331), .ZN(n35333) );
  INV_X2 U13684 ( .I(n60152), .ZN(n1806) );
  NAND2_X2 U1872 ( .A1(n982), .A2(n41951), .ZN(n41799) );
  INV_X4 U11628 ( .I(n10503), .ZN(n35320) );
  INV_X2 U3432 ( .I(n23699), .ZN(n26446) );
  NOR3_X2 U33083 ( .A1(n13172), .A2(n13171), .A3(n35889), .ZN(n13170) );
  NAND2_X2 U3385 ( .A1(n23504), .A2(n23822), .ZN(n29352) );
  INV_X2 U4363 ( .I(n41506), .ZN(n42878) );
  AOI21_X2 U18407 ( .A1(n5357), .A2(n5356), .B(n5354), .ZN(n5534) );
  OAI22_X2 U18523 ( .A1(n5355), .A2(n1540), .B1(n11061), .B2(n35688), .ZN(
        n5354) );
  AOI22_X2 U3182 ( .A1(n22576), .A2(n28182), .B1(n27684), .B2(n29689), .ZN(
        n27685) );
  NAND3_X2 U19533 ( .A1(n18825), .A2(n18824), .A3(n18823), .ZN(n22576) );
  NAND2_X2 U38647 ( .A1(n36057), .A2(n60196), .ZN(n36531) );
  NOR2_X2 U1155 ( .A1(n9331), .A2(n1480), .ZN(n47517) );
  INV_X4 U3126 ( .I(n19118), .ZN(n31269) );
  NAND3_X2 U8239 ( .A1(n30885), .A2(n12893), .A3(n23008), .ZN(n31252) );
  NOR2_X2 U2641 ( .A1(n35713), .A2(n34404), .ZN(n35841) );
  NAND2_X2 U13267 ( .A1(n36970), .A2(n37446), .ZN(n37252) );
  NOR2_X2 U3388 ( .A1(n14876), .A2(n7129), .ZN(n26626) );
  INV_X2 U2922 ( .I(n30820), .ZN(n30808) );
  OAI21_X2 U13569 ( .A1(n12023), .A2(n9679), .B(n59534), .ZN(n35684) );
  BUF_X4 U14311 ( .I(Key[127]), .Z(n55765) );
  INV_X2 U1618 ( .I(n43104), .ZN(n42425) );
  NOR3_X2 U1438 ( .A1(n15175), .A2(n15064), .A3(n15063), .ZN(n15062) );
  OR2_X1 U16504 ( .A1(n40889), .A2(n40888), .Z(n40902) );
  NOR2_X2 U9374 ( .A1(n15481), .A2(n18611), .ZN(n10752) );
  BUF_X4 U9073 ( .I(Key[121]), .Z(n52317) );
  INV_X2 U8814 ( .I(n14331), .ZN(n36956) );
  INV_X4 U2749 ( .I(n32425), .ZN(n15184) );
  NAND2_X2 U2587 ( .A1(n34042), .A2(n2635), .ZN(n34601) );
  AOI21_X2 U19061 ( .A1(n29471), .A2(n60064), .B(n14193), .ZN(n29478) );
  NAND2_X2 U2004 ( .A1(n42225), .A2(n42235), .ZN(n41949) );
  NAND3_X2 U36926 ( .A1(n43491), .A2(n4467), .A3(n61743), .ZN(n20217) );
  NAND2_X2 U47613 ( .A1(n8356), .A2(n19364), .ZN(n36575) );
  NAND2_X2 U2305 ( .A1(n36338), .A2(n36740), .ZN(n34077) );
  NAND2_X2 U9769 ( .A1(n20907), .A2(n6345), .ZN(n19712) );
  INV_X2 U1270 ( .I(n47291), .ZN(n47298) );
  NAND2_X2 U4402 ( .A1(n45618), .A2(n59687), .ZN(n45953) );
  OAI21_X2 U14075 ( .A1(n26415), .A2(n28507), .B(n26736), .ZN(n26419) );
  NAND2_X2 U8589 ( .A1(n46058), .A2(n46057), .ZN(n21620) );
  BUF_X2 U13779 ( .I(n16820), .Z(n24017) );
  NAND2_X2 U35221 ( .A1(n18549), .A2(n24614), .ZN(n19790) );
  NAND3_X2 U9717 ( .A1(n28513), .A2(n28511), .A3(n28512), .ZN(n28524) );
  INV_X2 U1413 ( .I(n42984), .ZN(n46196) );
  NOR2_X2 U9489 ( .A1(n21615), .A2(n36170), .ZN(n36124) );
  NAND2_X2 U9296 ( .A1(n43780), .A2(n6233), .ZN(n20209) );
  NOR2_X2 U26834 ( .A1(n1432), .A2(n3761), .ZN(n31202) );
  BUF_X4 U19849 ( .I(n24885), .Z(n23328) );
  NAND2_X2 U40347 ( .A1(n20338), .A2(n2824), .ZN(n43237) );
  INV_X2 U41405 ( .I(n25823), .ZN(n48076) );
  NAND2_X2 U160 ( .A1(n56048), .A2(n56045), .ZN(n13960) );
  AOI21_X2 U11989 ( .A1(n28037), .A2(n28036), .B(n28228), .ZN(n6826) );
  NAND2_X2 U13593 ( .A1(n18199), .A2(n16179), .ZN(n16919) );
  INV_X1 U35646 ( .I(n56520), .ZN(n56476) );
  NAND2_X2 U317 ( .A1(n54312), .A2(n51838), .ZN(n54495) );
  INV_X2 U475 ( .I(n56572), .ZN(n51265) );
  OAI21_X1 U14642 ( .A1(n51254), .A2(n4740), .B(n6393), .ZN(n6392) );
  INV_X4 U13717 ( .I(n16736), .ZN(n1816) );
  INV_X1 U241 ( .I(n61361), .ZN(n2014) );
  INV_X4 U2322 ( .I(n36494), .ZN(n1525) );
  INV_X2 U43112 ( .I(n30311), .ZN(n24467) );
  NAND3_X2 U19419 ( .A1(n28840), .A2(n28839), .A3(n28841), .ZN(n23058) );
  NAND3_X2 U3856 ( .A1(n46361), .A2(n46360), .A3(n46359), .ZN(n46366) );
  NOR2_X2 U2955 ( .A1(n29954), .A2(n30771), .ZN(n30784) );
  NAND2_X2 U4144 ( .A1(n43364), .A2(n995), .ZN(n41551) );
  NAND2_X2 U36705 ( .A1(n41858), .A2(n41270), .ZN(n39933) );
  NAND2_X1 U20171 ( .A1(n2052), .A2(n2051), .ZN(n12688) );
  NOR2_X1 U20172 ( .A1(n2053), .A2(n54920), .ZN(n2052) );
  INV_X2 U2116 ( .I(n15701), .ZN(n38786) );
  NOR2_X2 U13364 ( .A1(n8132), .A2(n1416), .ZN(n37387) );
  NAND2_X2 U3980 ( .A1(n23226), .A2(n37351), .ZN(n37115) );
  INV_X2 U17231 ( .I(n38692), .ZN(n2089) );
  NAND3_X2 U39879 ( .A1(n22927), .A2(n22586), .A3(n35804), .ZN(n20597) );
  INV_X2 U4360 ( .I(n900), .ZN(n34530) );
  NOR2_X2 U7273 ( .A1(n49430), .A2(n49377), .ZN(n49541) );
  INV_X4 U7785 ( .I(n59866), .ZN(n46271) );
  INV_X4 U11174 ( .I(n10970), .ZN(n42697) );
  NOR2_X2 U7284 ( .A1(n23707), .A2(n61355), .ZN(n50097) );
  NOR2_X2 U33783 ( .A1(n23522), .A2(n14226), .ZN(n52949) );
  NOR2_X2 U52255 ( .A1(n344), .A2(n47291), .ZN(n45932) );
  INV_X2 U3407 ( .I(n14834), .ZN(n15650) );
  BUF_X4 U37760 ( .I(n46813), .Z(n23099) );
  BUF_X4 U28046 ( .I(n14759), .Z(n7979) );
  INV_X1 U6673 ( .I(n5348), .ZN(n19811) );
  NOR2_X2 U10354 ( .A1(n32684), .A2(n22428), .ZN(n32990) );
  INV_X2 U11717 ( .I(n35685), .ZN(n24688) );
  BUF_X2 U17465 ( .I(n39781), .Z(n40387) );
  NOR2_X2 U21246 ( .A1(n1713), .A2(n42838), .ZN(n42674) );
  OR2_X1 U30442 ( .A1(n35563), .A2(n15870), .Z(n35176) );
  OR2_X2 U10061 ( .A1(n12962), .A2(n1714), .Z(n12961) );
  NAND2_X1 U2584 ( .A1(n34144), .A2(n19662), .ZN(n19664) );
  INV_X1 U3740 ( .I(n42405), .ZN(n42402) );
  NAND2_X2 U36026 ( .A1(n43089), .A2(n43088), .ZN(n43090) );
  BUF_X4 U9370 ( .I(n61388), .Z(n24981) );
  INV_X4 U10355 ( .I(n13043), .ZN(n18488) );
  NAND2_X2 U44758 ( .A1(n28986), .A2(n1192), .ZN(n28988) );
  NOR2_X2 U8946 ( .A1(n30585), .A2(n1316), .ZN(n29482) );
  INV_X2 U794 ( .I(n61742), .ZN(n22570) );
  BUF_X4 U10862 ( .I(n7738), .Z(n9177) );
  NAND2_X1 U26563 ( .A1(n6956), .A2(n6955), .ZN(n6881) );
  NAND2_X2 U10442 ( .A1(n29239), .A2(n29835), .ZN(n6769) );
  NAND2_X2 U3315 ( .A1(n28004), .A2(n25992), .ZN(n11226) );
  CLKBUF_X4 U3440 ( .I(n23286), .Z(n23037) );
  BUF_X4 U45096 ( .I(Key[179]), .Z(n56901) );
  CLKBUF_X4 U17556 ( .I(n6927), .Z(n3717) );
  INV_X2 U42994 ( .I(n24200), .ZN(n57079) );
  INV_X2 U39748 ( .I(n23533), .ZN(n48717) );
  INV_X2 U570 ( .I(n4470), .ZN(n51385) );
  NAND2_X2 U39904 ( .A1(n1516), .A2(n59871), .ZN(n40707) );
  NOR2_X2 U11052 ( .A1(n43133), .A2(n43134), .ZN(n16954) );
  NAND3_X2 U11910 ( .A1(n18530), .A2(n18529), .A3(n18528), .ZN(n7081) );
  NAND3_X1 U6013 ( .A1(n34965), .A2(n34963), .A3(n34964), .ZN(n34967) );
  NOR2_X2 U1773 ( .A1(n41299), .A2(n41298), .ZN(n43241) );
  INV_X2 U43883 ( .I(n15775), .ZN(n48665) );
  INV_X2 U556 ( .I(n9011), .ZN(n8821) );
  NAND2_X1 U2360 ( .A1(n36454), .A2(n1419), .ZN(n36455) );
  INV_X4 U1304 ( .I(n16616), .ZN(n44770) );
  INV_X4 U2054 ( .I(n26113), .ZN(n41306) );
  BUF_X2 U13214 ( .I(n23049), .Z(n4105) );
  INV_X2 U22354 ( .I(n3716), .ZN(n5298) );
  INV_X2 U1084 ( .I(n48553), .ZN(n48154) );
  INV_X2 U3285 ( .I(n5124), .ZN(n27522) );
  NOR2_X2 U8455 ( .A1(n11578), .A2(n53163), .ZN(n53165) );
  INV_X2 U10412 ( .I(n28735), .ZN(n28738) );
  OAI22_X2 U9715 ( .A1(n29651), .A2(n10148), .B1(n29383), .B2(n28662), .ZN(
        n20170) );
  NAND4_X2 U5249 ( .A1(n10759), .A2(n10757), .A3(n10758), .A4(n34087), .ZN(
        n10075) );
  BUF_X4 U24011 ( .I(n23194), .Z(n4734) );
  NOR2_X2 U18176 ( .A1(n10104), .A2(n10103), .ZN(n20798) );
  INV_X2 U44934 ( .I(n28192), .ZN(n28872) );
  NOR2_X2 U8010 ( .A1(n12034), .A2(n42019), .ZN(n13229) );
  OAI21_X1 U5484 ( .A1(n48523), .A2(n48522), .B(n48521), .ZN(n588) );
  NAND2_X1 U49080 ( .A1(n37242), .A2(n9869), .ZN(n37244) );
  INV_X4 U25840 ( .I(n36691), .ZN(n25964) );
  INV_X2 U8506 ( .I(n15244), .ZN(n55292) );
  NAND2_X2 U9199 ( .A1(n47061), .A2(n48870), .ZN(n7756) );
  INV_X1 U6940 ( .I(n30076), .ZN(n1845) );
  INV_X4 U34727 ( .I(n15507), .ZN(n21099) );
  CLKBUF_X8 U8246 ( .I(n31221), .Z(n1218) );
  INV_X4 U8122 ( .I(n48536), .ZN(n19361) );
  NOR2_X2 U8861 ( .A1(n15303), .A2(n33012), .ZN(n33019) );
  AOI21_X1 U19 ( .A1(n54702), .A2(n54701), .B(n54700), .ZN(n19383) );
  NOR2_X2 U9546 ( .A1(n17282), .A2(n31609), .ZN(n33675) );
  INV_X2 U39509 ( .I(n26127), .ZN(n34155) );
  INV_X2 U18661 ( .I(n33012), .ZN(n33304) );
  NAND2_X2 U960 ( .A1(n18252), .A2(n49673), .ZN(n49367) );
  NAND3_X1 U43497 ( .A1(n50451), .A2(n50450), .A3(n25274), .ZN(n51144) );
  NAND2_X2 U38385 ( .A1(n29191), .A2(n27282), .ZN(n17307) );
  AOI21_X1 U9877 ( .A1(n12536), .A2(n17929), .B(n1632), .ZN(n4362) );
  INV_X1 U1843 ( .I(n13525), .ZN(n40563) );
  NOR2_X2 U53771 ( .A1(n4699), .A2(n50142), .ZN(n50139) );
  INV_X4 U902 ( .I(n8727), .ZN(n7868) );
  NAND2_X2 U2433 ( .A1(n4541), .A2(n37361), .ZN(n37293) );
  INV_X2 U11507 ( .I(n35452), .ZN(n36054) );
  NAND2_X2 U11666 ( .A1(n33445), .A2(n35047), .ZN(n34497) );
  INV_X4 U2393 ( .I(n22524), .ZN(n35909) );
  OAI22_X2 U1569 ( .A1(n22802), .A2(n12503), .B1(n41489), .B2(n16677), .ZN(
        n41494) );
  NOR2_X1 U14693 ( .A1(n5496), .A2(n5495), .ZN(n6669) );
  NAND2_X2 U3318 ( .A1(n27523), .A2(n24734), .ZN(n27206) );
  NAND3_X2 U5338 ( .A1(n9327), .A2(n9326), .A3(n28790), .ZN(n2668) );
  INV_X1 U13670 ( .I(n61108), .ZN(n34781) );
  NOR3_X2 U5966 ( .A1(n52907), .A2(n52906), .A3(n55413), .ZN(n52916) );
  INV_X2 U7945 ( .I(n65283), .ZN(n19968) );
  NOR2_X2 U2342 ( .A1(n3864), .A2(n21605), .ZN(n36130) );
  INV_X4 U992 ( .I(n50218), .ZN(n7588) );
  INV_X1 U10368 ( .I(n34447), .ZN(n9030) );
  AOI21_X2 U55865 ( .A1(n54822), .A2(n54814), .B(n54653), .ZN(n54655) );
  NAND2_X2 U9185 ( .A1(n16829), .A2(n48843), .ZN(n49524) );
  INV_X2 U8387 ( .I(n24911), .ZN(n9602) );
  BUF_X2 U11402 ( .I(n38433), .Z(n23062) );
  AOI21_X2 U15806 ( .A1(n46842), .A2(n46841), .B(n14268), .ZN(n46847) );
  NAND2_X2 U19409 ( .A1(n11859), .A2(n13415), .ZN(n11814) );
  OAI21_X2 U14086 ( .A1(n28644), .A2(n60603), .B(n28182), .ZN(n13415) );
  OAI21_X2 U5451 ( .A1(n19193), .A2(n7404), .B(n43005), .ZN(n46291) );
  NOR2_X2 U1244 ( .A1(n47874), .A2(n12647), .ZN(n47883) );
  NAND2_X2 U8542 ( .A1(n50752), .A2(n48683), .ZN(n21602) );
  AOI22_X2 U45345 ( .A1(n29439), .A2(n29438), .B1(n29437), .B2(n29436), .ZN(
        n29445) );
  NAND3_X2 U8985 ( .A1(n13414), .A2(n27894), .A3(n13416), .ZN(n11815) );
  NOR2_X2 U30055 ( .A1(n30084), .A2(n1318), .ZN(n28788) );
  INV_X4 U41550 ( .I(n36536), .ZN(n36533) );
  BUF_X4 U45087 ( .I(Key[185]), .Z(n56976) );
  NOR2_X2 U1670 ( .A1(n61744), .A2(n13678), .ZN(n43178) );
  NAND4_X1 U52707 ( .A1(n45899), .A2(n70), .A3(n45901), .A4(n45898), .ZN(
        n45904) );
  NAND4_X1 U23937 ( .A1(n54747), .A2(n54746), .A3(n54745), .A4(n54744), .ZN(
        n54749) );
  NOR3_X1 U3992 ( .A1(n9489), .A2(n17607), .A3(n9490), .ZN(n5178) );
  INV_X2 U24219 ( .I(n54798), .ZN(n54626) );
  NAND2_X2 U1617 ( .A1(n17848), .A2(n42785), .ZN(n43022) );
  NAND4_X2 U13240 ( .A1(n33941), .A2(n33940), .A3(n33939), .A4(n33938), .ZN(
        n33942) );
  BUF_X2 U12494 ( .I(n50395), .Z(n21183) );
  INV_X2 U2032 ( .I(n14616), .ZN(n41125) );
  NAND2_X2 U9239 ( .A1(n16437), .A2(n47382), .ZN(n47376) );
  NOR2_X2 U3102 ( .A1(n25241), .A2(n21222), .ZN(n29019) );
  AOI22_X2 U18298 ( .A1(n21651), .A2(n33637), .B1(n33642), .B2(n33536), .ZN(
        n12747) );
  INV_X4 U7361 ( .I(n55643), .ZN(n8259) );
  AOI22_X2 U11941 ( .A1(n8628), .A2(n8626), .B1(n27983), .B2(n1320), .ZN(
        n18529) );
  NAND3_X2 U2230 ( .A1(n36973), .A2(n909), .A3(n1309), .ZN(n12460) );
  NAND2_X2 U2014 ( .A1(n21492), .A2(n42285), .ZN(n17349) );
  NOR2_X2 U3358 ( .A1(n19269), .A2(n7322), .ZN(n22482) );
  NAND2_X1 U23131 ( .A1(n41633), .A2(n43612), .ZN(n4344) );
  NOR2_X2 U35530 ( .A1(n58648), .A2(n50221), .ZN(n49348) );
  NAND2_X2 U7568 ( .A1(n2369), .A2(n2267), .ZN(n30263) );
  NAND2_X1 U42601 ( .A1(n48182), .A2(n48588), .ZN(n24654) );
  BUF_X4 U53007 ( .I(n46679), .Z(n47186) );
  NAND2_X2 U14775 ( .A1(n58380), .A2(n8828), .ZN(n56621) );
  INV_X2 U9015 ( .I(n27392), .ZN(n18780) );
  NAND2_X1 U10942 ( .A1(n46915), .A2(n46916), .ZN(n16877) );
  INV_X4 U22841 ( .I(n61710), .ZN(n41113) );
  BUF_X2 U17533 ( .I(n15932), .Z(n23962) );
  NAND2_X2 U53155 ( .A1(n64488), .A2(n19107), .ZN(n48925) );
  NAND2_X2 U13580 ( .A1(n19053), .A2(n34646), .ZN(n5186) );
  NOR2_X2 U9649 ( .A1(n29511), .A2(n29506), .ZN(n29509) );
  OAI21_X1 U17821 ( .A1(n35906), .A2(n3589), .B(n1911), .ZN(n3583) );
  OAI22_X2 U11593 ( .A1(n34619), .A2(n34082), .B1(n34081), .B2(n6360), .ZN(
        n10759) );
  INV_X2 U19626 ( .I(n27974), .ZN(n8628) );
  NOR2_X2 U38446 ( .A1(n1793), .A2(n23778), .ZN(n35991) );
  NAND3_X1 U49502 ( .A1(n37965), .A2(n37964), .A3(n37963), .ZN(n39524) );
  AOI21_X2 U35150 ( .A1(n20687), .A2(n48154), .B(n46788), .ZN(n23076) );
  NAND4_X2 U21672 ( .A1(n34911), .A2(n34910), .A3(n35435), .A4(n34909), .ZN(
        n3155) );
  AOI22_X1 U51470 ( .A1(n42900), .A2(n43169), .B1(n42899), .B2(n43150), .ZN(
        n42904) );
  INV_X4 U20058 ( .I(n1967), .ZN(n24117) );
  INV_X1 U12261 ( .I(n55403), .ZN(n52914) );
  NOR2_X2 U1206 ( .A1(n64548), .A2(n12647), .ZN(n47718) );
  NOR3_X2 U2493 ( .A1(n3581), .A2(n19240), .A3(n31540), .ZN(n20436) );
  INV_X1 U14273 ( .I(n25992), .ZN(n2569) );
  AOI21_X1 U51624 ( .A1(n25210), .A2(n43515), .B(n43514), .ZN(n43523) );
  OAI21_X1 U14886 ( .A1(n15706), .A2(n5668), .B(n24404), .ZN(n5667) );
  INV_X2 U1098 ( .I(n47101), .ZN(n48147) );
  INV_X2 U2148 ( .I(n36158), .ZN(n1750) );
  INV_X1 U41381 ( .I(n53462), .ZN(n53519) );
  BUF_X4 U7972 ( .I(n20399), .Z(n19735) );
  NOR2_X2 U3265 ( .A1(n20540), .A2(n28384), .ZN(n28387) );
  INV_X2 U13191 ( .I(n3053), .ZN(n37699) );
  INV_X1 U7348 ( .I(n23411), .ZN(n25199) );
  INV_X1 U37384 ( .I(n56454), .ZN(n56453) );
  AND2_X2 U10373 ( .A1(n35027), .A2(n1427), .Z(n34019) );
  NAND2_X2 U8927 ( .A1(n8336), .A2(n29019), .ZN(n29793) );
  NOR2_X2 U15240 ( .A1(n48715), .A2(n48714), .ZN(n11270) );
  AND3_X2 U42910 ( .A1(n19156), .A2(n23324), .A3(n28308), .Z(n26341) );
  NOR2_X2 U3366 ( .A1(n24431), .A2(n23753), .ZN(n27849) );
  INV_X2 U534 ( .I(n54112), .ZN(n13940) );
  NAND2_X1 U9236 ( .A1(n9101), .A2(n9100), .ZN(n9099) );
  INV_X4 U491 ( .I(n19434), .ZN(n1457) );
  INV_X2 U9541 ( .I(n62322), .ZN(n24317) );
  NAND3_X2 U12515 ( .A1(n47479), .A2(n47478), .A3(n47477), .ZN(n47480) );
  NAND2_X2 U1248 ( .A1(n48209), .A2(n48199), .ZN(n47201) );
  INV_X1 U15068 ( .I(n55722), .ZN(n1615) );
  BUF_X2 U14278 ( .I(n26802), .Z(n23303) );
  NOR2_X1 U50975 ( .A1(n41124), .A2(n41123), .ZN(n41129) );
  NAND3_X2 U53433 ( .A1(n49677), .A2(n49671), .A3(n49676), .ZN(n48006) );
  AOI22_X1 U3799 ( .A1(n33327), .A2(n34377), .B1(n34372), .B2(n36590), .ZN(
        n33332) );
  BUF_X4 U14315 ( .I(Key[165]), .Z(n56702) );
  NAND2_X1 U2907 ( .A1(n682), .A2(n7944), .ZN(n15528) );
  AOI21_X1 U22951 ( .A1(n43689), .A2(n7282), .B(n4229), .ZN(n12447) );
  INV_X1 U10049 ( .I(n57177), .ZN(n1332) );
  OR2_X2 U3237 ( .A1(n21720), .A2(n3617), .Z(n820) );
  NOR2_X2 U2237 ( .A1(n1786), .A2(n60694), .ZN(n36628) );
  NOR2_X2 U11778 ( .A1(n30742), .A2(n30739), .ZN(n10711) );
  NAND2_X2 U4002 ( .A1(n34972), .A2(n34970), .ZN(n32919) );
  INV_X2 U11948 ( .I(n28229), .ZN(n26277) );
  NOR2_X2 U9870 ( .A1(n5701), .A2(n5699), .ZN(n4528) );
  INV_X2 U37751 ( .I(n22427), .ZN(n36886) );
  INV_X2 U45545 ( .I(n30531), .ZN(n29937) );
  NAND3_X1 U44651 ( .A1(n27440), .A2(n27439), .A3(n27438), .ZN(n27446) );
  INV_X2 U50525 ( .I(n40845), .ZN(n40843) );
  NAND2_X2 U3253 ( .A1(n27337), .A2(n1356), .ZN(n29385) );
  OR2_X2 U22401 ( .A1(n30736), .A2(n30748), .Z(n30738) );
  AOI22_X1 U55645 ( .A1(n54051), .A2(n54050), .B1(n54049), .B2(n54048), .ZN(
        n54061) );
  AOI22_X2 U41943 ( .A1(n28749), .A2(n17413), .B1(n29860), .B2(n17414), .ZN(
        n28750) );
  INV_X1 U35436 ( .I(n38056), .ZN(n18051) );
  NAND3_X2 U2505 ( .A1(n34996), .A2(n13899), .A3(n13898), .ZN(n13358) );
  NOR3_X2 U8079 ( .A1(n11582), .A2(n11581), .A3(n11580), .ZN(n11579) );
  NAND2_X2 U22651 ( .A1(n11608), .A2(n7950), .ZN(n11607) );
  NAND3_X1 U49610 ( .A1(n41833), .A2(n41293), .A3(n59976), .ZN(n38132) );
  INV_X2 U13993 ( .I(n29766), .ZN(n1551) );
  NAND2_X1 U4740 ( .A1(n49482), .A2(n48854), .ZN(n49304) );
  NOR2_X2 U11773 ( .A1(n6321), .A2(n6319), .ZN(n6318) );
  OAI21_X2 U47834 ( .A1(n33394), .A2(n34140), .B(n33393), .ZN(n33402) );
  NOR3_X2 U9626 ( .A1(n28928), .A2(n9689), .A3(n9688), .ZN(n20731) );
  NOR3_X2 U15421 ( .A1(n49094), .A2(n49095), .A3(n8459), .ZN(n2631) );
  NAND2_X2 U8803 ( .A1(n1772), .A2(n35482), .ZN(n18857) );
  INV_X1 U26554 ( .I(n6867), .ZN(n30463) );
  BUF_X2 U9074 ( .I(Key[94]), .Z(n55087) );
  CLKBUF_X2 U3022 ( .I(Key[181]), .Z(n52294) );
  NAND2_X1 U32711 ( .A1(n34967), .A2(n34968), .ZN(n12633) );
  INV_X2 U23271 ( .I(n12072), .ZN(n13764) );
  NAND2_X2 U16087 ( .A1(n47301), .A2(n47292), .ZN(n12359) );
  INV_X4 U23546 ( .I(n24948), .ZN(n30396) );
  INV_X4 U22514 ( .I(n3935), .ZN(n5322) );
  BUF_X2 U16293 ( .I(n48103), .Z(n23850) );
  AND2_X2 U3357 ( .A1(n27114), .A2(n22735), .Z(n26540) );
  OAI22_X2 U53866 ( .A1(n49464), .A2(n49463), .B1(n49462), .B2(n49739), .ZN(
        n49470) );
  NAND3_X2 U29778 ( .A1(n49461), .A2(n49460), .A3(n10831), .ZN(n49464) );
  INV_X2 U52568 ( .I(n45932), .ZN(n45936) );
  INV_X2 U42847 ( .I(n44627), .ZN(n46688) );
  OAI21_X2 U10343 ( .A1(n26242), .A2(n35306), .B(n34708), .ZN(n32070) );
  INV_X2 U13122 ( .I(n22502), .ZN(n19938) );
  AOI22_X2 U44730 ( .A1(n27671), .A2(n27828), .B1(n27670), .B2(n27669), .ZN(
        n27672) );
  INV_X2 U16900 ( .I(n23984), .ZN(n14496) );
  BUF_X2 U2031 ( .I(n42288), .Z(n6412) );
  NOR2_X1 U48412 ( .A1(n35357), .A2(n35141), .ZN(n35143) );
  NAND2_X2 U9055 ( .A1(n19279), .A2(n28872), .ZN(n29673) );
  INV_X2 U8182 ( .I(n49923), .ZN(n24362) );
  NAND2_X2 U13024 ( .A1(n2340), .A2(n41381), .ZN(n2339) );
  BUF_X2 U12196 ( .I(n55595), .Z(n4801) );
  OR2_X1 U29071 ( .A1(n11215), .A2(n11216), .Z(n9069) );
  BUF_X4 U19911 ( .I(Key[77]), .Z(n54587) );
  BUF_X2 U24437 ( .I(n33277), .Z(n33797) );
  BUF_X2 U18840 ( .I(n33178), .Z(n23465) );
  INV_X4 U16223 ( .I(n59216), .ZN(n3597) );
  AOI21_X1 U50731 ( .A1(n42448), .A2(n41306), .B(n40357), .ZN(n40358) );
  NOR2_X2 U34896 ( .A1(n33115), .A2(n59125), .ZN(n33536) );
  NAND2_X2 U35248 ( .A1(n23215), .A2(n32984), .ZN(n35532) );
  NOR2_X2 U17975 ( .A1(n36883), .A2(n37233), .ZN(n37161) );
  NOR2_X2 U11058 ( .A1(n3957), .A2(n3955), .ZN(n3954) );
  OAI21_X2 U14492 ( .A1(n55645), .A2(n55631), .B(n17500), .ZN(n52307) );
  INV_X4 U43729 ( .I(n30029), .ZN(n29732) );
  BUF_X4 U18128 ( .I(n35899), .Z(n24118) );
  BUF_X4 U30304 ( .I(n1557), .Z(n10068) );
  INV_X4 U1302 ( .I(n47881), .ZN(n14473) );
  NAND3_X2 U16396 ( .A1(n40184), .A2(n40183), .A3(n40182), .ZN(n40185) );
  INV_X2 U2738 ( .I(n34606), .ZN(n17922) );
  NOR2_X2 U32720 ( .A1(n12647), .A2(n45183), .ZN(n47726) );
  NOR2_X2 U7025 ( .A1(n25927), .A2(n29729), .ZN(n5632) );
  NOR2_X2 U12413 ( .A1(n48309), .A2(n1639), .ZN(n12496) );
  OR2_X1 U43833 ( .A1(n34739), .A2(n34737), .Z(n26168) );
  OAI21_X1 U19446 ( .A1(n28006), .A2(n11226), .B(n3382), .ZN(n28011) );
  NOR2_X2 U11392 ( .A1(n35381), .A2(n35380), .ZN(n36900) );
  NOR2_X2 U9257 ( .A1(n1656), .A2(n9860), .ZN(n47655) );
  NOR3_X2 U27634 ( .A1(n17352), .A2(n17353), .A3(n17351), .ZN(n7567) );
  INV_X4 U9708 ( .I(n29010), .ZN(n30588) );
  NAND2_X1 U2522 ( .A1(n13576), .A2(n9757), .ZN(n30465) );
  INV_X4 U30841 ( .I(n61743), .ZN(n16864) );
  NOR2_X2 U7091 ( .A1(n37333), .A2(n37010), .ZN(n37341) );
  INV_X4 U9585 ( .I(n34233), .ZN(n26242) );
  OAI21_X1 U47598 ( .A1(n32936), .A2(n33741), .B(n34726), .ZN(n32937) );
  NOR2_X2 U813 ( .A1(n18585), .A2(n6977), .ZN(n50363) );
  OAI22_X2 U13890 ( .A1(n29470), .A2(n30421), .B1(n31084), .B2(n18060), .ZN(
        n14193) );
  INV_X2 U28930 ( .I(n49471), .ZN(n49999) );
  NAND3_X2 U766 ( .A1(n57425), .A2(n16986), .A3(n48366), .ZN(n49288) );
  NAND3_X1 U3667 ( .A1(n10106), .A2(n17185), .A3(n42455), .ZN(n17184) );
  INV_X2 U8813 ( .I(n37048), .ZN(n1772) );
  INV_X2 U9204 ( .I(n17816), .ZN(n47451) );
  AOI21_X2 U11632 ( .A1(n34946), .A2(n10528), .B(n1345), .ZN(n11581) );
  NOR2_X1 U15693 ( .A1(n3096), .A2(n23597), .ZN(n3095) );
  NOR2_X2 U4278 ( .A1(n6313), .A2(n25162), .ZN(n45231) );
  AOI22_X2 U35454 ( .A1(n40738), .A2(n20889), .B1(n19992), .B2(n41400), .ZN(
        n24176) );
  INV_X1 U26169 ( .I(n23849), .ZN(n6510) );
  INV_X2 U3413 ( .I(n1447), .ZN(n24734) );
  BUF_X4 U23723 ( .I(n31470), .Z(n34168) );
  NOR2_X2 U1517 ( .A1(n42697), .A2(n41970), .ZN(n42704) );
  INV_X4 U3903 ( .I(n53212), .ZN(n25160) );
  NAND3_X2 U10102 ( .A1(n12286), .A2(n39423), .A3(n994), .ZN(n21965) );
  NAND2_X2 U8451 ( .A1(n60297), .A2(n592), .ZN(n15011) );
  NAND2_X2 U18037 ( .A1(n35508), .A2(n35507), .ZN(n35505) );
  OAI21_X2 U2503 ( .A1(n35209), .A2(n35208), .B(n35207), .ZN(n35264) );
  BUF_X4 U9592 ( .I(n6530), .Z(n22428) );
  NAND2_X1 U10204 ( .A1(n14342), .A2(n14341), .ZN(n9992) );
  AOI21_X2 U15356 ( .A1(n4733), .A2(n4208), .B(n4206), .ZN(n4205) );
  OAI21_X2 U12830 ( .A1(n63983), .A2(n20650), .B(n43627), .ZN(n43631) );
  INV_X2 U43686 ( .I(n57183), .ZN(n53451) );
  INV_X2 U30593 ( .I(n50359), .ZN(n50004) );
  AOI21_X2 U11853 ( .A1(n59481), .A2(n17745), .B(n24206), .ZN(n29961) );
  INV_X2 U29036 ( .I(n34149), .ZN(n34146) );
  OAI21_X2 U17672 ( .A1(n34895), .A2(n35464), .B(n3012), .ZN(n3011) );
  NAND3_X1 U56385 ( .A1(n56025), .A2(n9568), .A3(n56024), .ZN(n56026) );
  INV_X2 U3370 ( .I(n28273), .ZN(n21946) );
  NOR2_X2 U55414 ( .A1(n54057), .A2(n54054), .ZN(n53551) );
  NOR3_X2 U16486 ( .A1(n6071), .A2(n6073), .A3(n6072), .ZN(n6068) );
  NOR2_X1 U16648 ( .A1(n42342), .A2(n16740), .ZN(n16739) );
  OAI21_X2 U3179 ( .A1(n28229), .A2(n28228), .B(n6222), .ZN(n15609) );
  INV_X2 U10578 ( .I(n21301), .ZN(n18224) );
  OAI22_X1 U22950 ( .A1(n5816), .A2(n40363), .B1(n38200), .B2(n4227), .ZN(
        n4424) );
  INV_X1 U757 ( .I(n4212), .ZN(n3044) );
  AND2_X2 U32934 ( .A1(n27184), .A2(n12929), .Z(n28112) );
  OAI21_X1 U9632 ( .A1(n30701), .A2(n3985), .B(n31035), .ZN(n3984) );
  OAI22_X2 U8986 ( .A1(n27383), .A2(n16069), .B1(n4059), .B2(n21151), .ZN(
        n7142) );
  BUF_X4 U23025 ( .I(n4294), .Z(n4265) );
  NAND3_X2 U7074 ( .A1(n31537), .A2(n31536), .A3(n14319), .ZN(n20445) );
  BUF_X4 U14316 ( .I(Key[129]), .Z(n55792) );
  NAND2_X2 U17237 ( .A1(n38404), .A2(n41166), .ZN(n39070) );
  INV_X1 U17283 ( .I(n6841), .ZN(n41391) );
  INV_X2 U6347 ( .I(n41376), .ZN(n41378) );
  INV_X1 U6847 ( .I(n26856), .ZN(n6382) );
  NAND2_X1 U2856 ( .A1(n24282), .A2(n31122), .ZN(n120) );
  NOR2_X2 U45765 ( .A1(n33718), .A2(n63421), .ZN(n30459) );
  INV_X1 U8911 ( .I(n5688), .ZN(n30477) );
  INV_X1 U32124 ( .I(n26667), .ZN(n30480) );
  INV_X2 U2166 ( .I(n58203), .ZN(n38575) );
  NAND3_X2 U35389 ( .A1(n23884), .A2(n40650), .A3(n10452), .ZN(n38404) );
  INV_X4 U26677 ( .I(n6996), .ZN(n38273) );
  OAI22_X2 U18963 ( .A1(n26914), .A2(n57392), .B1(n31036), .B2(n26916), .ZN(
        n19465) );
  INV_X1 U5093 ( .I(n22498), .ZN(n18203) );
  INV_X2 U11874 ( .I(n22579), .ZN(n1861) );
  INV_X2 U13944 ( .I(n29565), .ZN(n27797) );
  OAI21_X2 U44735 ( .A1(n29695), .A2(n27887), .B(n27683), .ZN(n27684) );
  NOR2_X2 U2582 ( .A1(n33465), .A2(n61748), .ZN(n34790) );
  BUF_X4 U5840 ( .I(n43867), .Z(n45199) );
  BUF_X2 U12042 ( .I(n12070), .Z(n10309) );
  BUF_X2 U12090 ( .I(n28488), .Z(n17589) );
  NOR4_X2 U10512 ( .A1(n17604), .A2(n26821), .A3(n17603), .A4(n28486), .ZN(
        n17602) );
  INV_X4 U9276 ( .I(n47797), .ZN(n47699) );
  BUF_X2 U9252 ( .I(n47826), .Z(n7050) );
  INV_X2 U43728 ( .I(n1865), .ZN(n30027) );
  BUF_X4 U12113 ( .I(Key[151]), .Z(n56309) );
  AOI22_X1 U13325 ( .A1(n57266), .A2(n2002), .B1(n15794), .B2(n16191), .ZN(
        n17687) );
  INV_X1 U22480 ( .I(n25166), .ZN(n47832) );
  INV_X2 U934 ( .I(n58269), .ZN(n48979) );
  AND2_X2 U26870 ( .A1(n28426), .A2(n9865), .Z(n29571) );
  INV_X4 U32313 ( .I(n26791), .ZN(n28615) );
  NAND2_X2 U9270 ( .A1(n47370), .A2(n23718), .ZN(n16438) );
  INV_X2 U6976 ( .I(n29316), .ZN(n19967) );
  OAI21_X2 U1023 ( .A1(n45761), .A2(n46076), .B(n45760), .ZN(n48070) );
  AOI22_X2 U637 ( .A1(n50138), .A2(n50139), .B1(n50136), .B2(n50137), .ZN(
        n23640) );
  OAI21_X2 U40130 ( .A1(n41971), .A2(n41525), .B(n42707), .ZN(n41530) );
  INV_X4 U12093 ( .I(n7651), .ZN(n1443) );
  AOI21_X1 U12546 ( .A1(n10763), .A2(n21200), .B(n1649), .ZN(n10762) );
  INV_X2 U47543 ( .I(n33567), .ZN(n32810) );
  INV_X1 U11321 ( .I(n39992), .ZN(n41377) );
  NAND3_X1 U31144 ( .A1(n38041), .A2(n58364), .A3(n61986), .ZN(n12876) );
  NAND4_X2 U2203 ( .A1(n34898), .A2(n36699), .A3(n34896), .A4(n34897), .ZN(
        n34899) );
  INV_X2 U28012 ( .I(n29779), .ZN(n29251) );
  NAND3_X2 U1509 ( .A1(n43850), .A2(n43078), .A3(n60052), .ZN(n43082) );
  NOR2_X2 U12025 ( .A1(n1358), .A2(n28843), .ZN(n19620) );
  NAND4_X1 U34654 ( .A1(n30175), .A2(n30174), .A3(n58999), .A4(n15407), .ZN(
        n23121) );
  OR2_X1 U19108 ( .A1(n14399), .A2(n8802), .Z(n8804) );
  INV_X1 U12077 ( .I(n25785), .ZN(n27536) );
  INV_X2 U18926 ( .I(n28994), .ZN(n14854) );
  NAND2_X2 U4355 ( .A1(n37328), .A2(n9830), .ZN(n37339) );
  BUF_X2 U13749 ( .I(n33030), .Z(n14249) );
  OAI22_X2 U11834 ( .A1(n29266), .A2(n24316), .B1(n13817), .B2(n2429), .ZN(
        n2430) );
  INV_X2 U17747 ( .I(n20502), .ZN(n10816) );
  NAND3_X2 U8984 ( .A1(n26369), .A2(n26368), .A3(n26367), .ZN(n29795) );
  INV_X2 U20107 ( .I(n61735), .ZN(n26163) );
  AOI21_X2 U8774 ( .A1(n4831), .A2(n36687), .B(n62720), .ZN(n5033) );
  INV_X2 U7918 ( .I(n21597), .ZN(n55286) );
  CLKBUF_X2 U14294 ( .I(Key[97]), .Z(n24065) );
  AOI21_X2 U1775 ( .A1(n40851), .A2(n2760), .B(n2759), .ZN(n25929) );
  NAND2_X2 U45910 ( .A1(n30802), .A2(n30801), .ZN(n30806) );
  INV_X1 U13164 ( .I(n16601), .ZN(n40607) );
  INV_X4 U31580 ( .I(n13731), .ZN(n11205) );
  NAND2_X1 U52077 ( .A1(n44564), .A2(n59384), .ZN(n44565) );
  INV_X2 U13996 ( .I(n1437), .ZN(n8584) );
  INV_X2 U11835 ( .I(n29085), .ZN(n29078) );
  NOR2_X2 U4423 ( .A1(n24586), .A2(n53881), .ZN(n24923) );
  NAND3_X2 U4571 ( .A1(n14852), .A2(n14851), .A3(n14850), .ZN(n14849) );
  OR2_X1 U17658 ( .A1(n26221), .A2(n5462), .Z(n5461) );
  INV_X2 U9812 ( .I(n53816), .ZN(n53823) );
  NAND2_X2 U1011 ( .A1(n45604), .A2(n45603), .ZN(n45608) );
  INV_X2 U9148 ( .I(n15362), .ZN(n53024) );
  AOI22_X1 U47537 ( .A1(n33570), .A2(n32805), .B1(n32804), .B2(n32803), .ZN(
        n32813) );
  BUF_X2 U45446 ( .I(Key[118]), .Z(n55580) );
  NAND2_X2 U1013 ( .A1(n45604), .A2(n45936), .ZN(n45609) );
  INV_X2 U21477 ( .I(n3027), .ZN(n23209) );
  OAI21_X2 U14047 ( .A1(n28047), .A2(n28046), .B(n21065), .ZN(n28057) );
  NOR2_X2 U4152 ( .A1(n60855), .A2(n22860), .ZN(n55801) );
  NOR3_X2 U15210 ( .A1(n49082), .A2(n49081), .A3(n49080), .ZN(n49083) );
  NAND2_X2 U37989 ( .A1(n17410), .A2(n16631), .ZN(n21626) );
  NAND3_X1 U39613 ( .A1(n52769), .A2(n53588), .A3(n52998), .ZN(n19201) );
  INV_X2 U5959 ( .I(n13297), .ZN(n1420) );
  NAND4_X1 U7292 ( .A1(n49606), .A2(n48314), .A3(n49613), .A4(n49318), .ZN(
        n9385) );
  INV_X2 U8998 ( .I(n28243), .ZN(n28069) );
  NOR4_X2 U48938 ( .A1(n36910), .A2(n64967), .A3(n22461), .A4(n22595), .ZN(
        n36911) );
  BUF_X4 U7583 ( .I(n34238), .Z(n23743) );
  OAI21_X1 U10916 ( .A1(n14437), .A2(n48236), .B(n48112), .ZN(n49864) );
  NOR2_X2 U9492 ( .A1(n37329), .A2(n24661), .ZN(n37009) );
  BUF_X8 U24589 ( .I(n37428), .Z(n22461) );
  INV_X4 U3291 ( .I(n4081), .ZN(n28648) );
  NOR2_X2 U7017 ( .A1(n30211), .A2(n22416), .ZN(n30843) );
  NAND2_X1 U42105 ( .A1(n35746), .A2(n35745), .ZN(n24462) );
  AOI21_X2 U10095 ( .A1(n16173), .A2(n14017), .B(n14012), .ZN(n20216) );
  BUF_X2 U45511 ( .I(Key[83]), .Z(n54776) );
  NAND2_X2 U17636 ( .A1(n37414), .A2(n5005), .ZN(n5004) );
  NOR2_X2 U10096 ( .A1(n11080), .A2(n11079), .ZN(n11078) );
  BUF_X4 U14306 ( .I(Key[164]), .Z(n56692) );
  NOR2_X2 U7013 ( .A1(n7979), .A2(n14399), .ZN(n28996) );
  NAND3_X2 U9938 ( .A1(n8137), .A2(n8136), .A3(n8134), .ZN(n8133) );
  NAND3_X2 U54 ( .A1(n18287), .A2(n55351), .A3(n55373), .ZN(n18286) );
  NOR2_X2 U1547 ( .A1(n41624), .A2(n22446), .ZN(n43605) );
  INV_X2 U31493 ( .I(n11041), .ZN(n53192) );
  NAND3_X2 U9230 ( .A1(n44400), .A2(n44398), .A3(n44399), .ZN(n44406) );
  INV_X2 U34721 ( .I(n15503), .ZN(n41820) );
  INV_X2 U1707 ( .I(n15540), .ZN(n1299) );
  INV_X2 U13178 ( .I(n10554), .ZN(n1517) );
  NAND4_X1 U21209 ( .A1(n36133), .A2(n36132), .A3(n36131), .A4(n2857), .ZN(
        n36137) );
  INV_X2 U28690 ( .I(n22146), .ZN(n32206) );
  INV_X1 U18812 ( .I(n8463), .ZN(n9570) );
  NAND3_X2 U35184 ( .A1(n54018), .A2(n4564), .A3(n61123), .ZN(n54351) );
  NAND2_X2 U21249 ( .A1(n17467), .A2(n541), .ZN(n17501) );
  NOR2_X1 U11085 ( .A1(n9080), .A2(n43896), .ZN(n3425) );
  NAND2_X1 U4717 ( .A1(n26776), .A2(n89), .ZN(n13935) );
  INV_X2 U3300 ( .I(n29148), .ZN(n29153) );
  NAND2_X1 U9673 ( .A1(n24448), .A2(n30302), .ZN(n28425) );
  INV_X1 U1344 ( .I(n22142), .ZN(n44980) );
  INV_X2 U20963 ( .I(n2670), .ZN(n23941) );
  NOR2_X1 U10645 ( .A1(n11936), .A2(n11937), .ZN(n53654) );
  INV_X2 U29246 ( .I(n24964), .ZN(n24091) );
  INV_X2 U13687 ( .I(n33978), .ZN(n34034) );
  INV_X2 U19365 ( .I(n24896), .ZN(n2119) );
  NOR3_X1 U39806 ( .A1(n53271), .A2(n53270), .A3(n20980), .ZN(n19453) );
  INV_X2 U9732 ( .I(n820), .ZN(n27981) );
  OAI21_X2 U37434 ( .A1(n55631), .A2(n15700), .B(n19020), .ZN(n55612) );
  NAND3_X2 U2175 ( .A1(n37346), .A2(n37344), .A3(n37345), .ZN(n20470) );
  NAND2_X2 U2386 ( .A1(n14904), .A2(n22524), .ZN(n34863) );
  INV_X1 U26653 ( .I(n49990), .ZN(n20894) );
  INV_X1 U8117 ( .I(n45411), .ZN(n23718) );
  INV_X2 U2994 ( .I(n29019), .ZN(n29797) );
  INV_X4 U26094 ( .I(n24418), .ZN(n28842) );
  NOR2_X2 U45772 ( .A1(n18300), .A2(n34993), .ZN(n34070) );
  INV_X2 U2841 ( .I(n63050), .ZN(n33905) );
  BUF_X4 U14013 ( .I(n28690), .Z(n30192) );
  NOR2_X2 U9756 ( .A1(n19156), .A2(n27595), .ZN(n28309) );
  OAI22_X2 U50982 ( .A1(n41459), .A2(n41455), .B1(n41454), .B2(n41154), .ZN(
        n41157) );
  NAND2_X2 U13615 ( .A1(n33737), .A2(n34719), .ZN(n34251) );
  NAND2_X2 U28861 ( .A1(n22230), .A2(n29457), .ZN(n28736) );
  INV_X2 U11653 ( .I(n33737), .ZN(n34248) );
  INV_X1 U43574 ( .I(n33628), .ZN(n33537) );
  INV_X2 U3041 ( .I(n28898), .ZN(n30481) );
  INV_X2 U23094 ( .I(n4320), .ZN(n33540) );
  NAND2_X1 U15408 ( .A1(n50007), .A2(n50006), .ZN(n16672) );
  NAND3_X2 U53502 ( .A1(n48253), .A2(n64922), .A3(n48251), .ZN(n48258) );
  BUF_X2 U10639 ( .I(Key[146]), .Z(n56165) );
  CLKBUF_X4 U29818 ( .I(Key[51]), .Z(n23886) );
  CLKBUF_X2 U5683 ( .I(Key[139]), .Z(n56030) );
  CLKBUF_X2 U10632 ( .I(Key[142]), .Z(n56097) );
  BUF_X2 U2945 ( .I(Key[75]), .Z(n54556) );
  BUF_X2 U9072 ( .I(Key[45]), .Z(n23754) );
  BUF_X2 U19916 ( .I(Key[87]), .Z(n24051) );
  CLKBUF_X2 U6035 ( .I(n21656), .Z(n435) );
  CLKBUF_X2 U12099 ( .I(n28589), .Z(n19593) );
  CLKBUF_X4 U19890 ( .I(n28192), .Z(n29661) );
  CLKBUF_X4 U19858 ( .I(n26456), .Z(n29372) );
  INV_X1 U19897 ( .I(n56692), .ZN(n56693) );
  INV_X2 U44344 ( .I(n26862), .ZN(n28624) );
  CLKBUF_X4 U19866 ( .I(n26388), .Z(n27665) );
  BUF_X2 U19875 ( .I(n28537), .Z(n23508) );
  BUF_X2 U19874 ( .I(n22691), .Z(n22821) );
  INV_X2 U29899 ( .I(n21264), .ZN(n21265) );
  BUF_X2 U9066 ( .I(n54748), .Z(n9871) );
  INV_X2 U45091 ( .I(n50486), .ZN(n50793) );
  BUF_X2 U19835 ( .I(n44262), .Z(n22950) );
  INV_X4 U3445 ( .I(n14604), .ZN(n27485) );
  CLKBUF_X2 U14267 ( .I(n29317), .Z(n9987) );
  BUF_X2 U19807 ( .I(n28328), .Z(n23997) );
  BUF_X2 U19846 ( .I(n42812), .Z(n22323) );
  INV_X2 U3482 ( .I(n20753), .ZN(n27097) );
  INV_X1 U19816 ( .I(n26010), .ZN(n22129) );
  CLKBUF_X2 U3335 ( .I(n8478), .Z(n8613) );
  CLKBUF_X2 U5351 ( .I(n38880), .Z(n245) );
  INV_X2 U28087 ( .I(n60816), .ZN(n27567) );
  CLKBUF_X2 U14231 ( .I(n51005), .Z(n9753) );
  BUF_X2 U3254 ( .I(n10403), .Z(n7495) );
  CLKBUF_X2 U5261 ( .I(n37786), .Z(n23789) );
  INV_X1 U5213 ( .I(n27854), .ZN(n211) );
  OR2_X1 U34321 ( .A1(n29118), .A2(n14947), .Z(n21804) );
  NAND2_X1 U14152 ( .A1(n1886), .A2(n820), .ZN(n3827) );
  CLKBUF_X2 U5363 ( .I(n50650), .Z(n247) );
  NAND2_X1 U19747 ( .A1(n14434), .A2(n14433), .ZN(n26948) );
  CLKBUF_X4 U4727 ( .I(n28250), .Z(n93) );
  CLKBUF_X1 U14120 ( .I(n44163), .Z(n10304) );
  NAND2_X1 U45144 ( .A1(n64451), .A2(n28861), .ZN(n28864) );
  OR2_X1 U37563 ( .A1(n27402), .A2(n27401), .Z(n15976) );
  INV_X1 U19539 ( .I(n28191), .ZN(n10305) );
  NAND2_X1 U19639 ( .A1(n29125), .A2(n29124), .ZN(n15025) );
  OAI21_X1 U25722 ( .A1(n27103), .A2(n61643), .B(n28231), .ZN(n6048) );
  CLKBUF_X1 U36560 ( .I(n52461), .Z(n19862) );
  CLKBUF_X1 U14064 ( .I(n31970), .Z(n4544) );
  INV_X1 U4546 ( .I(n2547), .ZN(n2546) );
  CLKBUF_X4 U3147 ( .I(n30087), .Z(n22903) );
  CLKBUF_X4 U19385 ( .I(n30844), .Z(n22596) );
  CLKBUF_X4 U10500 ( .I(n28920), .Z(n9865) );
  INV_X4 U11907 ( .I(n31247), .ZN(n1436) );
  CLKBUF_X1 U10502 ( .I(n31270), .Z(n22934) );
  CLKBUF_X4 U19380 ( .I(n28059), .Z(n30322) );
  INV_X2 U14009 ( .I(n18129), .ZN(n24335) );
  CLKBUF_X4 U42872 ( .I(n27085), .Z(n24000) );
  CLKBUF_X1 U13965 ( .I(n28683), .Z(n30001) );
  CLKBUF_X2 U4986 ( .I(n20747), .Z(n161) );
  INV_X1 U11840 ( .I(n22696), .ZN(n30750) );
  CLKBUF_X8 U9683 ( .I(n5163), .Z(n5070) );
  INV_X1 U19314 ( .I(n3908), .ZN(n29508) );
  INV_X1 U44843 ( .I(n28788), .ZN(n30086) );
  INV_X2 U2979 ( .I(n30046), .ZN(n1349) );
  INV_X1 U35463 ( .I(n30651), .ZN(n30653) );
  NAND2_X1 U7015 ( .A1(n29482), .A2(n1437), .ZN(n12858) );
  INV_X1 U44782 ( .I(n29855), .ZN(n28744) );
  INV_X1 U3768 ( .I(n30173), .ZN(n30175) );
  INV_X1 U19255 ( .I(n30704), .ZN(n6256) );
  NAND2_X1 U46153 ( .A1(n7461), .A2(n31137), .ZN(n31139) );
  INV_X1 U45070 ( .I(n29551), .ZN(n28721) );
  INV_X1 U8910 ( .I(n29545), .ZN(n29964) );
  NAND2_X1 U24161 ( .A1(n20282), .A2(n29891), .ZN(n5691) );
  NOR2_X1 U26974 ( .A1(n30297), .A2(n21313), .ZN(n21312) );
  AOI21_X1 U45184 ( .A1(n29906), .A2(n31182), .B(n28969), .ZN(n28970) );
  INV_X1 U19037 ( .I(n29434), .ZN(n3262) );
  AOI21_X1 U19102 ( .A1(n3445), .A2(n18880), .B(n6428), .ZN(n3444) );
  NAND2_X1 U20941 ( .A1(n5985), .A2(n5984), .ZN(n2651) );
  NAND3_X1 U13817 ( .A1(n28913), .A2(n28912), .A3(n28919), .ZN(n25506) );
  INV_X1 U3071 ( .I(n19721), .ZN(n6343) );
  BUF_X2 U18865 ( .I(n33185), .Z(n23683) );
  BUF_X2 U18923 ( .I(n33906), .Z(n22583) );
  CLKBUF_X8 U10396 ( .I(n22540), .Z(n17463) );
  CLKBUF_X4 U2830 ( .I(n25174), .Z(n21172) );
  INV_X1 U35224 ( .I(n496), .ZN(n21581) );
  CLKBUF_X2 U18758 ( .I(n31719), .Z(n7323) );
  CLKBUF_X4 U10379 ( .I(n31315), .Z(n34119) );
  CLKBUF_X2 U6836 ( .I(n9330), .Z(n4685) );
  BUF_X2 U10384 ( .I(n34341), .Z(n20989) );
  CLKBUF_X4 U21560 ( .I(n35025), .Z(n3082) );
  INV_X2 U2741 ( .I(n25849), .ZN(n34088) );
  CLKBUF_X4 U11718 ( .I(n32133), .Z(n1426) );
  BUF_X2 U18765 ( .I(n23781), .Z(n19457) );
  NAND2_X1 U18471 ( .A1(n5927), .A2(n61449), .ZN(n34501) );
  INV_X4 U7593 ( .I(n15756), .ZN(n34640) );
  INV_X2 U5106 ( .I(n61699), .ZN(n35612) );
  CLKBUF_X1 U10375 ( .I(n25372), .Z(n23567) );
  NOR2_X1 U13667 ( .A1(n2695), .A2(n34114), .ZN(n31724) );
  INV_X2 U10357 ( .I(n34623), .ZN(n34084) );
  CLKBUF_X4 U18654 ( .I(n34149), .Z(n23757) );
  NAND2_X1 U21925 ( .A1(n32869), .A2(n3363), .ZN(n14291) );
  INV_X2 U13658 ( .I(n33984), .ZN(n34607) );
  INV_X2 U18481 ( .I(n20443), .ZN(n34041) );
  CLKBUF_X2 U6286 ( .I(n6205), .Z(n10608) );
  NOR2_X1 U25593 ( .A1(n5927), .A2(n31300), .ZN(n35036) );
  INV_X1 U47907 ( .I(n35207), .ZN(n33546) );
  CLKBUF_X4 U2635 ( .I(n7797), .Z(n5529) );
  INV_X1 U18573 ( .I(n32700), .ZN(n7537) );
  NOR2_X1 U3676 ( .A1(n34246), .A2(n34721), .ZN(n32928) );
  NAND2_X1 U40798 ( .A1(n33118), .A2(n24093), .ZN(n20913) );
  INV_X1 U4481 ( .I(n33307), .ZN(n33595) );
  NAND4_X1 U48266 ( .A1(n34674), .A2(n34673), .A3(n34672), .A4(n34671), .ZN(
        n34684) );
  NAND2_X1 U13548 ( .A1(n18773), .A2(n1805), .ZN(n15453) );
  INV_X2 U9570 ( .I(n14913), .ZN(n14954) );
  INV_X1 U18420 ( .I(n33347), .ZN(n3995) );
  NAND2_X1 U18472 ( .A1(n33006), .A2(n32785), .ZN(n4892) );
  OAI21_X1 U47990 ( .A1(n33800), .A2(n33799), .B(n35659), .ZN(n33804) );
  INV_X1 U6724 ( .I(n33494), .ZN(n33770) );
  NAND3_X1 U22360 ( .A1(n34966), .A2(n25404), .A3(n127), .ZN(n3721) );
  AOI22_X1 U48565 ( .A1(n35634), .A2(n35633), .B1(n35632), .B2(n35631), .ZN(
        n35637) );
  INV_X1 U48144 ( .I(n35298), .ZN(n34261) );
  NAND2_X1 U18397 ( .A1(n32925), .A2(n32926), .ZN(n25290) );
  AOI22_X1 U40842 ( .A1(n35838), .A2(n35842), .B1(n35836), .B2(n35837), .ZN(
        n35840) );
  NAND3_X1 U18279 ( .A1(n33514), .A2(n58076), .A3(n33512), .ZN(n33515) );
  INV_X1 U47886 ( .I(n33506), .ZN(n33507) );
  NAND2_X1 U18276 ( .A1(n35211), .A2(n35210), .ZN(n4161) );
  NAND4_X1 U13518 ( .A1(n17040), .A2(n19824), .A3(n31776), .A4(n17039), .ZN(
        n19822) );
  NAND2_X1 U18406 ( .A1(n9889), .A2(n12166), .ZN(n11580) );
  AOI21_X1 U48370 ( .A1(n35008), .A2(n35007), .B(n35006), .ZN(n35018) );
  INV_X1 U42799 ( .I(n34160), .ZN(n26122) );
  CLKBUF_X2 U4617 ( .I(n36410), .Z(n55) );
  INV_X2 U4351 ( .I(n15742), .ZN(n18205) );
  CLKBUF_X4 U17914 ( .I(n36195), .Z(n23503) );
  CLKBUF_X2 U10257 ( .I(n9830), .Z(n5807) );
  INV_X1 U49079 ( .I(n62992), .ZN(n37242) );
  INV_X2 U29168 ( .I(n35173), .ZN(n9721) );
  CLKBUF_X4 U38348 ( .I(n34836), .Z(n17243) );
  BUF_X4 U18118 ( .I(n37269), .Z(n22733) );
  CLKBUF_X1 U6808 ( .I(n13297), .Z(n685) );
  INV_X1 U48218 ( .I(n35949), .ZN(n36920) );
  INV_X1 U18077 ( .I(n35483), .ZN(n37052) );
  NAND2_X1 U49016 ( .A1(n23842), .A2(n22733), .ZN(n37134) );
  INV_X1 U18083 ( .I(n36130), .ZN(n36138) );
  NAND3_X1 U11398 ( .A1(n36612), .A2(n60431), .A3(n36613), .ZN(n18672) );
  AOI22_X1 U5919 ( .A1(n10963), .A2(n35982), .B1(n20712), .B2(n24994), .ZN(
        n10962) );
  INV_X1 U25640 ( .I(n36786), .ZN(n36787) );
  INV_X1 U48830 ( .I(n36572), .ZN(n36573) );
  NAND2_X1 U17955 ( .A1(n35064), .A2(n35063), .ZN(n26019) );
  NAND3_X1 U6863 ( .A1(n34105), .A2(n34106), .A3(n12116), .ZN(n699) );
  AOI22_X1 U36468 ( .A1(n37019), .A2(n37940), .B1(n37018), .B2(n37017), .ZN(
        n20419) );
  INV_X1 U10253 ( .I(n36580), .ZN(n1767) );
  NOR2_X1 U34165 ( .A1(n31781), .A2(n31784), .ZN(n14723) );
  NAND2_X1 U17727 ( .A1(n25297), .A2(n25296), .ZN(n6833) );
  OAI22_X1 U25550 ( .A1(n36361), .A2(n36362), .B1(n5900), .B2(n36962), .ZN(
        n7724) );
  OAI21_X1 U21037 ( .A1(n13209), .A2(n2715), .B(n36582), .ZN(n2716) );
  NOR2_X1 U13231 ( .A1(n35115), .A2(n35114), .ZN(n35126) );
  INV_X1 U41204 ( .I(n24962), .ZN(n21502) );
  NOR2_X1 U11408 ( .A1(n35405), .A2(n19380), .ZN(n35413) );
  INV_X2 U37493 ( .I(n25155), .ZN(n37174) );
  BUF_X2 U2153 ( .I(n19314), .Z(n14) );
  INV_X2 U10199 ( .I(n39315), .ZN(n1757) );
  CLKBUF_X4 U11373 ( .I(n39579), .Z(n15729) );
  INV_X1 U50003 ( .I(n39554), .ZN(n38756) );
  BUF_X2 U13177 ( .I(n36649), .Z(n40070) );
  INV_X2 U2050 ( .I(n17382), .ZN(n41152) );
  INV_X2 U31768 ( .I(n15590), .ZN(n17966) );
  CLKBUF_X2 U5367 ( .I(n37173), .Z(n40258) );
  CLKBUF_X2 U8755 ( .I(n13050), .Z(n9935) );
  INV_X2 U9452 ( .I(n41160), .ZN(n1306) );
  CLKBUF_X2 U6889 ( .I(n40661), .Z(n709) );
  INV_X1 U38651 ( .I(n40039), .ZN(n42468) );
  INV_X2 U33189 ( .I(n36106), .ZN(n41031) );
  NOR2_X1 U10134 ( .A1(n39509), .A2(n1407), .ZN(n8131) );
  INV_X2 U42718 ( .I(n40490), .ZN(n41178) );
  INV_X2 U1839 ( .I(n60971), .ZN(n40123) );
  NAND2_X1 U17315 ( .A1(n5581), .A2(n42261), .ZN(n41096) );
  NAND2_X1 U36633 ( .A1(n41101), .A2(n61984), .ZN(n40445) );
  NOR3_X1 U49956 ( .A1(n40732), .A2(n40729), .A3(n38678), .ZN(n38679) );
  INV_X2 U5031 ( .I(n41294), .ZN(n42528) );
  AND2_X1 U7725 ( .A1(n41425), .A2(n40766), .Z(n997) );
  INV_X1 U35053 ( .I(n40609), .ZN(n20054) );
  INV_X1 U8711 ( .I(n40606), .ZN(n16465) );
  OAI21_X1 U17341 ( .A1(n42293), .A2(n42292), .B(n42507), .ZN(n15369) );
  NAND2_X1 U17314 ( .A1(n41205), .A2(n41204), .ZN(n9788) );
  INV_X2 U5374 ( .I(n11704), .ZN(n20974) );
  INV_X1 U1874 ( .I(n4227), .ZN(n41804) );
  NAND2_X1 U12999 ( .A1(n9788), .A2(n41206), .ZN(n41207) );
  NAND3_X1 U12945 ( .A1(n41305), .A2(n41304), .A3(n41803), .ZN(n9081) );
  NAND3_X1 U9385 ( .A1(n42513), .A2(n42512), .A3(n42511), .ZN(n42514) );
  CLKBUF_X4 U10079 ( .I(n21665), .Z(n19591) );
  NOR2_X1 U17023 ( .A1(n16395), .A2(n16394), .ZN(n16393) );
  BUF_X2 U16984 ( .I(n40537), .Z(n42668) );
  BUF_X2 U16992 ( .I(n40537), .Z(n10004) );
  CLKBUF_X4 U10048 ( .I(n20086), .Z(n1494) );
  INV_X4 U7170 ( .I(n43156), .ZN(n15214) );
  CLKBUF_X4 U16915 ( .I(n43319), .Z(n24779) );
  BUF_X4 U16974 ( .I(n41242), .Z(n42676) );
  NAND2_X1 U42017 ( .A1(n40673), .A2(n40671), .ZN(n22813) );
  BUF_X4 U16929 ( .I(n43717), .Z(n23314) );
  BUF_X2 U12872 ( .I(n12089), .Z(n12091) );
  CLKBUF_X4 U7717 ( .I(n41131), .Z(n2994) );
  INV_X2 U21334 ( .I(n42716), .ZN(n43583) );
  INV_X1 U29930 ( .I(n16473), .ZN(n42900) );
  OR2_X1 U12913 ( .A1(n1709), .A2(n59292), .Z(n42751) );
  INV_X1 U22478 ( .I(n42393), .ZN(n42392) );
  NOR2_X1 U16815 ( .A1(n6144), .A2(n61198), .ZN(n43870) );
  INV_X2 U7199 ( .I(n43092), .ZN(n42006) );
  INV_X2 U11205 ( .I(n42726), .ZN(n1397) );
  NAND2_X1 U12915 ( .A1(n41559), .A2(n42139), .ZN(n3630) );
  AOI21_X1 U51425 ( .A1(n2994), .A2(n43569), .B(n59746), .ZN(n42718) );
  NOR2_X1 U9332 ( .A1(n41716), .A2(n42112), .ZN(n41599) );
  NAND2_X1 U36942 ( .A1(n43506), .A2(n43505), .ZN(n17560) );
  INV_X1 U12924 ( .I(n41715), .ZN(n42559) );
  INV_X1 U6153 ( .I(n42346), .ZN(n472) );
  NAND2_X1 U38653 ( .A1(n17755), .A2(n43948), .ZN(n42988) );
  OAI21_X1 U21285 ( .A1(n43583), .A2(n42339), .B(n2898), .ZN(n41141) );
  INV_X1 U16738 ( .I(n41322), .ZN(n43266) );
  INV_X1 U7184 ( .I(n43578), .ZN(n13547) );
  NOR2_X1 U26752 ( .A1(n57255), .A2(n43914), .ZN(n12642) );
  NAND3_X1 U1572 ( .A1(n13730), .A2(n12089), .A3(n23488), .ZN(n43541) );
  NAND2_X1 U1701 ( .A1(n1269), .A2(n57808), .ZN(n42105) );
  NOR2_X1 U51394 ( .A1(n43266), .A2(n43122), .ZN(n42615) );
  NOR3_X1 U50670 ( .A1(n41972), .A2(n41969), .A3(n42383), .ZN(n40171) );
  NAND2_X1 U4145 ( .A1(n43364), .A2(n4322), .ZN(n42740) );
  OAI21_X1 U11116 ( .A1(n13167), .A2(n11635), .B(n43144), .ZN(n9080) );
  NAND2_X1 U43753 ( .A1(n43000), .A2(n43100), .ZN(n43001) );
  OAI21_X1 U16507 ( .A1(n41324), .A2(n4672), .B(n63205), .ZN(n7677) );
  NAND2_X1 U20676 ( .A1(n42656), .A2(n2450), .ZN(n25672) );
  AND2_X1 U50648 ( .A1(n25851), .A2(n42968), .Z(n40082) );
  NAND2_X1 U9994 ( .A1(n39936), .A2(n10998), .ZN(n39937) );
  OR2_X1 U25883 ( .A1(n43779), .A2(n12091), .Z(n6232) );
  NOR2_X1 U16450 ( .A1(n8321), .A2(n17859), .ZN(n8320) );
  CLKBUF_X4 U27602 ( .I(n46121), .Z(n7544) );
  NAND2_X1 U12738 ( .A1(n10159), .A2(n18153), .ZN(n21759) );
  NAND3_X1 U16518 ( .A1(n40098), .A2(n42965), .A3(n40097), .ZN(n18575) );
  CLKBUF_X2 U6795 ( .I(n44098), .Z(n672) );
  NAND2_X1 U16414 ( .A1(n6421), .A2(n13450), .ZN(n6419) );
  BUF_X2 U12725 ( .I(n46253), .Z(n22731) );
  CLKBUF_X4 U1366 ( .I(n46605), .Z(n23553) );
  CLKBUF_X2 U42163 ( .I(n26248), .Z(n22994) );
  INV_X1 U16342 ( .I(n14514), .ZN(n8385) );
  INV_X2 U16359 ( .I(n45045), .ZN(n46403) );
  CLKBUF_X1 U51472 ( .I(n45409), .Z(n42909) );
  CLKBUF_X2 U36104 ( .I(n11380), .Z(n23316) );
  INV_X2 U1317 ( .I(n43597), .ZN(n45183) );
  BUF_X2 U16267 ( .I(n47774), .Z(n7161) );
  INV_X2 U7814 ( .I(n47680), .ZN(n47421) );
  CLKBUF_X4 U27335 ( .I(n47851), .Z(n7395) );
  INV_X1 U37104 ( .I(n48641), .ZN(n48500) );
  CLKBUF_X2 U5452 ( .I(n47421), .Z(n263) );
  BUF_X2 U10996 ( .I(n16194), .Z(n8666) );
  INV_X2 U34747 ( .I(n47510), .ZN(n47516) );
  INV_X2 U1132 ( .I(n22468), .ZN(n47616) );
  NOR2_X1 U53176 ( .A1(n21178), .A2(n48538), .ZN(n47137) );
  INV_X1 U9955 ( .I(n48194), .ZN(n48664) );
  NOR2_X1 U12670 ( .A1(n47259), .A2(n47250), .ZN(n46884) );
  INV_X2 U20201 ( .I(n8152), .ZN(n47468) );
  INV_X2 U7471 ( .I(n11708), .ZN(n48577) );
  NAND2_X1 U41620 ( .A1(n47153), .A2(n46469), .ZN(n46471) );
  INV_X1 U5879 ( .I(n8043), .ZN(n48479) );
  INV_X1 U9259 ( .I(n4213), .ZN(n48523) );
  OR3_X1 U8346 ( .A1(n13356), .A2(n45590), .A3(n44840), .Z(n45943) );
  CLKBUF_X2 U12638 ( .I(n48567), .Z(n10250) );
  AOI21_X1 U10977 ( .A1(n62853), .A2(n16882), .B(n48654), .ZN(n12620) );
  INV_X1 U52140 ( .I(n46988), .ZN(n44684) );
  NAND2_X1 U52705 ( .A1(n47853), .A2(n1266), .ZN(n45896) );
  NOR2_X1 U52640 ( .A1(n45751), .A2(n62490), .ZN(n45752) );
  INV_X1 U53475 ( .I(n48261), .ZN(n48160) );
  OAI22_X1 U5464 ( .A1(n47427), .A2(n47690), .B1(n61216), .B2(n47428), .ZN(
        n11838) );
  NAND2_X1 U12622 ( .A1(n48653), .A2(n5717), .ZN(n44771) );
  INV_X1 U15950 ( .I(n46980), .ZN(n44685) );
  NAND2_X1 U52134 ( .A1(n46980), .A2(n46977), .ZN(n44678) );
  AOI21_X1 U12640 ( .A1(n47431), .A2(n47736), .B(n5132), .ZN(n5131) );
  NAND2_X1 U53484 ( .A1(n1659), .A2(n48178), .ZN(n48179) );
  NAND2_X1 U30199 ( .A1(n12687), .A2(n65275), .ZN(n44285) );
  NAND2_X1 U15924 ( .A1(n24339), .A2(n3081), .ZN(n24338) );
  AOI22_X1 U12551 ( .A1(n7051), .A2(n48641), .B1(n12997), .B2(n48160), .ZN(
        n12996) );
  OAI21_X1 U15863 ( .A1(n47981), .A2(n46946), .B(n46945), .ZN(n18465) );
  INV_X1 U15866 ( .I(n47152), .ZN(n13527) );
  INV_X1 U37066 ( .I(n47022), .ZN(n47021) );
  NAND4_X1 U26779 ( .A1(n47165), .A2(n47164), .A3(n25481), .A4(n22635), .ZN(
        n47173) );
  INV_X1 U52605 ( .I(n45663), .ZN(n45664) );
  OAI21_X1 U35148 ( .A1(n16225), .A2(n22093), .B(n46948), .ZN(n45755) );
  NOR3_X1 U9922 ( .A1(n22206), .A2(n46073), .A3(n46072), .ZN(n4584) );
  AOI21_X1 U15789 ( .A1(n24338), .A2(n47230), .B(n47229), .ZN(n6574) );
  CLKBUF_X4 U5084 ( .I(n45229), .Z(n49739) );
  NAND2_X1 U52730 ( .A1(n45958), .A2(n5298), .ZN(n45959) );
  BUF_X2 U15696 ( .I(n49803), .Z(n7146) );
  CLKBUF_X4 U3857 ( .I(n49263), .Z(n7086) );
  NOR2_X1 U53113 ( .A1(n46932), .A2(n46931), .ZN(n46933) );
  CLKBUF_X4 U3744 ( .I(n16539), .Z(n6977) );
  INV_X1 U15498 ( .I(n49508), .ZN(n14205) );
  NAND2_X1 U53946 ( .A1(n19144), .A2(n5258), .ZN(n49813) );
  NAND2_X1 U31777 ( .A1(n64631), .A2(n49538), .ZN(n18814) );
  INV_X1 U8563 ( .I(n49723), .ZN(n1634) );
  NAND2_X1 U40905 ( .A1(n50074), .A2(n63084), .ZN(n21017) );
  CLKBUF_X4 U915 ( .I(n8727), .Z(n7866) );
  NOR2_X1 U15698 ( .A1(n47009), .A2(n19786), .ZN(n18511) );
  INV_X2 U28435 ( .I(n49171), .ZN(n49556) );
  NOR2_X1 U40834 ( .A1(n49205), .A2(n50004), .ZN(n49137) );
  OAI22_X1 U53418 ( .A1(n23156), .A2(n48413), .B1(n47967), .B2(n1630), .ZN(
        n47968) );
  NOR2_X1 U769 ( .A1(n49914), .A2(n13839), .ZN(n6030) );
  NOR2_X1 U15378 ( .A1(n48840), .A2(n49525), .ZN(n12337) );
  CLKBUF_X2 U4569 ( .I(n49564), .Z(n42) );
  INV_X1 U5103 ( .I(n49130), .ZN(n49136) );
  INV_X1 U53751 ( .I(n49829), .ZN(n49079) );
  INV_X1 U52751 ( .I(n48434), .ZN(n46005) );
  NAND2_X1 U53521 ( .A1(n48312), .A2(n49593), .ZN(n48313) );
  NAND2_X1 U41662 ( .A1(n50039), .A2(n13440), .ZN(n49437) );
  OAI21_X1 U9195 ( .A1(n7156), .A2(n50405), .B(n63084), .ZN(n50413) );
  OAI21_X1 U15219 ( .A1(n15301), .A2(n49937), .B(n17884), .ZN(n15300) );
  INV_X1 U22913 ( .I(n49619), .ZN(n4193) );
  NAND3_X1 U41330 ( .A1(n50293), .A2(n21790), .A3(n50292), .ZN(n21789) );
  INV_X2 U15373 ( .I(n14265), .ZN(n50383) );
  NAND3_X1 U22691 ( .A1(n49776), .A2(n49777), .A3(n149), .ZN(n4019) );
  NAND2_X1 U52397 ( .A1(n45233), .A2(n49467), .ZN(n45234) );
  NAND3_X1 U53238 ( .A1(n858), .A2(n47346), .A3(n47345), .ZN(n47350) );
  AOI21_X1 U53798 ( .A1(n49214), .A2(n49394), .B(n49397), .ZN(n49218) );
  NOR2_X1 U53329 ( .A1(n47645), .A2(n47644), .ZN(n47651) );
  CLKBUF_X4 U606 ( .I(n52623), .Z(n22338) );
  CLKBUF_X4 U8532 ( .I(n3333), .Z(n3334) );
  CLKBUF_X4 U15143 ( .I(n15066), .Z(n22478) );
  INV_X1 U12328 ( .I(n8065), .ZN(n52440) );
  CLKBUF_X4 U5288 ( .I(n52340), .Z(n19125) );
  INV_X2 U564 ( .I(n24929), .ZN(n18891) );
  CLKBUF_X2 U10767 ( .I(n55672), .Z(n24003) );
  BUF_X2 U15051 ( .I(n18230), .Z(n17935) );
  INV_X2 U30309 ( .I(n57032), .ZN(n15304) );
  CLKBUF_X2 U15054 ( .I(n53612), .Z(n22201) );
  INV_X2 U4343 ( .I(n52704), .ZN(n56540) );
  CLKBUF_X2 U7916 ( .I(n23982), .Z(n10362) );
  INV_X2 U6412 ( .I(n50601), .ZN(n52862) );
  CLKBUF_X2 U6352 ( .I(n25746), .Z(n533) );
  INV_X1 U55283 ( .I(n53847), .ZN(n54068) );
  INV_X2 U12286 ( .I(n5236), .ZN(n15706) );
  CLKBUF_X2 U8512 ( .I(n16948), .Z(n10551) );
  CLKBUF_X4 U505 ( .I(n52866), .Z(n20982) );
  OR2_X1 U32989 ( .A1(n56269), .A2(n15804), .Z(n13020) );
  INV_X1 U14759 ( .I(n51440), .ZN(n56608) );
  NAND2_X1 U23788 ( .A1(n53441), .A2(n53442), .ZN(n13401) );
  NAND2_X1 U14673 ( .A1(n56413), .A2(n56632), .ZN(n56423) );
  NAND2_X1 U3941 ( .A1(n54974), .A2(n54973), .ZN(n54976) );
  NOR2_X1 U14869 ( .A1(n1455), .A2(n17257), .ZN(n15897) );
  OAI21_X1 U9115 ( .A1(n1149), .A2(n6459), .B(n6220), .ZN(n6219) );
  BUF_X2 U14577 ( .I(n56352), .Z(n20957) );
  CLKBUF_X4 U28414 ( .I(n55135), .Z(n8325) );
  CLKBUF_X8 U259 ( .I(n23862), .Z(n4283) );
  CLKBUF_X4 U5667 ( .I(n54662), .Z(n54769) );
  INV_X1 U42858 ( .I(n55781), .ZN(n55760) );
  CLKBUF_X4 U3542 ( .I(n8325), .Z(n8027) );
  INV_X1 U111 ( .I(n55879), .ZN(n55900) );
  OR2_X1 U42972 ( .A1(n16978), .A2(n55209), .Z(n24146) );
  NAND2_X1 U9095 ( .A1(n53158), .A2(n53140), .ZN(n53144) );
  NAND2_X1 U113 ( .A1(n8307), .A2(n1919), .ZN(n54905) );
  INV_X1 U56662 ( .I(n56747), .ZN(n56755) );
  INV_X1 U110 ( .I(n56773), .ZN(n56756) );
  NAND3_X1 U6257 ( .A1(n22364), .A2(n56857), .A3(n56858), .ZN(n56860) );
  NAND3_X1 U43858 ( .A1(n53957), .A2(n53956), .A3(n53955), .ZN(n53959) );
  CLKBUF_X4 U42414 ( .I(Key[123]), .Z(n55624) );
  CLKBUF_X4 U19907 ( .I(Key[92]), .Z(n55060) );
  CLKBUF_X2 U14299 ( .I(Key[95]), .Z(n55106) );
  CLKBUF_X2 U12106 ( .I(Key[9]), .Z(n53154) );
  CLKBUF_X2 U12107 ( .I(Key[33]), .Z(n23858) );
  BUF_X2 U45901 ( .I(Key[99]), .Z(n55139) );
  BUF_X2 U19861 ( .I(n29167), .Z(n23769) );
  BUF_X2 U12085 ( .I(n28811), .Z(n20678) );
  CLKBUF_X2 U19873 ( .I(n28542), .Z(n22768) );
  BUF_X2 U19841 ( .I(n23469), .Z(n22203) );
  INV_X1 U20430 ( .I(n29104), .ZN(n2513) );
  AND3_X1 U37723 ( .A1(n29120), .A2(n22714), .A3(n60298), .Z(n16272) );
  CLKBUF_X1 U6019 ( .I(n13672), .Z(n430) );
  CLKBUF_X2 U9036 ( .I(n24124), .Z(n10049) );
  BUF_X2 U19774 ( .I(n45274), .Z(n22961) );
  INV_X2 U6540 ( .I(n29659), .ZN(n1356) );
  AND2_X1 U44858 ( .A1(n29105), .A2(n23665), .Z(n27950) );
  AND2_X1 U8994 ( .A1(n29108), .A2(n10404), .Z(n2123) );
  NAND2_X1 U14118 ( .A1(n29111), .A2(n19170), .ZN(n27951) );
  NAND2_X1 U20834 ( .A1(n27087), .A2(n58792), .ZN(n26345) );
  AOI21_X1 U19547 ( .A1(n17489), .A2(n26719), .B(n12706), .ZN(n22680) );
  NAND2_X1 U43992 ( .A1(n26315), .A2(n26314), .ZN(n30087) );
  CLKBUF_X4 U3162 ( .I(n24056), .Z(n12907) );
  CLKBUF_X4 U3817 ( .I(n61729), .Z(n8336) );
  OAI21_X1 U44763 ( .A1(n28986), .A2(n23315), .B(n28989), .ZN(n27748) );
  AOI22_X1 U19082 ( .A1(n28941), .A2(n28940), .B1(n28939), .B2(n14064), .ZN(
        n28947) );
  AOI21_X1 U34653 ( .A1(n1858), .A2(n30167), .B(n60112), .ZN(n29033) );
  INV_X1 U45012 ( .I(n29591), .ZN(n28917) );
  INV_X1 U33086 ( .I(n13175), .ZN(n20028) );
  NAND2_X1 U21073 ( .A1(n29802), .A2(n3150), .ZN(n9280) );
  NAND3_X1 U4747 ( .A1(n30052), .A2(n2252), .A3(n63140), .ZN(n100) );
  BUF_X4 U31814 ( .I(n23341), .Z(n11529) );
  CLKBUF_X1 U11746 ( .I(n18295), .Z(n10622) );
  INV_X1 U3545 ( .I(n32335), .ZN(n24413) );
  INV_X2 U9597 ( .I(n25891), .ZN(n35651) );
  BUF_X2 U13733 ( .I(n31465), .Z(n1547) );
  CLKBUF_X2 U11681 ( .I(n9971), .Z(n23179) );
  BUF_X2 U13714 ( .I(n25999), .Z(n23775) );
  INV_X1 U18611 ( .I(n35694), .ZN(n5355) );
  INV_X1 U40796 ( .I(n33118), .ZN(n33629) );
  NOR2_X1 U10316 ( .A1(n34747), .A2(n34740), .ZN(n35298) );
  INV_X1 U13572 ( .I(n32460), .ZN(n33612) );
  INV_X1 U13662 ( .I(n34646), .ZN(n35044) );
  INV_X1 U48369 ( .I(n35005), .ZN(n35006) );
  AOI21_X1 U35030 ( .A1(n33470), .A2(n33471), .B(n21317), .ZN(n33474) );
  NOR2_X1 U18277 ( .A1(n18801), .A2(n22642), .ZN(n18800) );
  NOR2_X1 U18137 ( .A1(n34124), .A2(n34123), .ZN(n14470) );
  NOR2_X1 U35006 ( .A1(n33007), .A2(n18568), .ZN(n33011) );
  BUF_X4 U27818 ( .I(n19473), .Z(n7729) );
  OR2_X1 U8043 ( .A1(n36443), .A2(n36435), .Z(n36441) );
  INV_X2 U5608 ( .I(n37492), .ZN(n37125) );
  CLKBUF_X2 U8245 ( .I(n4893), .Z(n1217) );
  CLKBUF_X2 U18094 ( .I(n35173), .Z(n7488) );
  INV_X2 U8821 ( .I(n1792), .ZN(n15038) );
  NAND2_X1 U30209 ( .A1(n23449), .A2(n36610), .ZN(n13656) );
  NAND2_X1 U25016 ( .A1(n35588), .A2(n36444), .ZN(n35590) );
  INV_X1 U18043 ( .I(n37293), .ZN(n37357) );
  OAI21_X1 U36538 ( .A1(n36721), .A2(n36212), .B(n36211), .ZN(n36213) );
  INV_X1 U6857 ( .I(n37111), .ZN(n36754) );
  INV_X1 U40216 ( .I(n36278), .ZN(n36962) );
  INV_X1 U13319 ( .I(n37168), .ZN(n37243) );
  NOR2_X1 U17989 ( .A1(n11272), .A2(n22113), .ZN(n34101) );
  NAND2_X1 U27010 ( .A1(n7732), .A2(n31782), .ZN(n31781) );
  AOI22_X1 U48311 ( .A1(n34827), .A2(n34826), .B1(n35391), .B2(n34828), .ZN(
        n34832) );
  INV_X1 U11427 ( .I(n36667), .ZN(n19380) );
  NAND2_X1 U40284 ( .A1(n36015), .A2(n36847), .ZN(n36016) );
  NOR2_X1 U17692 ( .A1(n22520), .A2(n34371), .ZN(n17924) );
  BUF_X2 U13236 ( .I(n39391), .Z(n18049) );
  CLKBUF_X4 U13200 ( .I(n19008), .Z(n18797) );
  INV_X1 U17560 ( .I(n36859), .ZN(n36505) );
  CLKBUF_X4 U49680 ( .I(n38234), .Z(n41858) );
  BUF_X2 U17491 ( .I(n40644), .Z(n10587) );
  CLKBUF_X4 U30314 ( .I(n41386), .Z(n10074) );
  BUF_X2 U17454 ( .I(n39099), .Z(n21381) );
  AND2_X1 U2024 ( .A1(n41020), .A2(n5531), .Z(n38421) );
  INV_X1 U23473 ( .I(n41854), .ZN(n22448) );
  INV_X1 U37758 ( .I(n19458), .ZN(n40604) );
  CLKBUF_X4 U5653 ( .I(n40303), .Z(n321) );
  INV_X4 U31243 ( .I(n40943), .ZN(n40952) );
  BUF_X2 U8712 ( .I(n6689), .Z(n22943) );
  NAND2_X1 U39865 ( .A1(n40027), .A2(n9091), .ZN(n22359) );
  OAI21_X1 U50993 ( .A1(n38935), .A2(n41216), .B(n61316), .ZN(n41217) );
  NOR3_X1 U1970 ( .A1(n6412), .A2(n11525), .A3(n42287), .ZN(n16870) );
  INV_X2 U32087 ( .I(n61658), .ZN(n40998) );
  OAI21_X1 U17010 ( .A1(n39899), .A2(n41843), .B(n5837), .ZN(n39902) );
  BUF_X2 U10178 ( .I(n1408), .Z(n9802) );
  AND2_X1 U1894 ( .A1(n40051), .A2(n19611), .Z(n13877) );
  NAND4_X1 U32530 ( .A1(n24122), .A2(n38695), .A3(n39069), .A4(n40543), .ZN(
        n38697) );
  AOI21_X1 U17052 ( .A1(n2337), .A2(n2336), .B(n41126), .ZN(n2335) );
  INV_X1 U17343 ( .I(n40489), .ZN(n40488) );
  NOR2_X1 U35842 ( .A1(n57303), .A2(n41174), .ZN(n41175) );
  NOR3_X1 U13012 ( .A1(n7326), .A2(n41174), .A3(n10517), .ZN(n40673) );
  BUF_X2 U1637 ( .I(n2995), .Z(n6865) );
  CLKBUF_X2 U16981 ( .I(n39841), .Z(n8676) );
  BUF_X4 U16918 ( .I(n24386), .Z(n22282) );
  CLKBUF_X2 U39594 ( .I(n3619), .Z(n19174) );
  NOR2_X1 U34786 ( .A1(n43290), .A2(n23700), .ZN(n24575) );
  NOR2_X1 U8112 ( .A1(n40334), .A2(n12353), .ZN(n40343) );
  INV_X2 U1674 ( .I(n1499), .ZN(n1694) );
  INV_X1 U1698 ( .I(n39175), .ZN(n43015) );
  INV_X4 U30150 ( .I(n26020), .ZN(n13478) );
  BUF_X4 U1725 ( .I(n39082), .Z(n42785) );
  NOR2_X1 U16611 ( .A1(n43316), .A2(n2496), .ZN(n42979) );
  AOI22_X1 U51692 ( .A1(n43709), .A2(n64156), .B1(n16880), .B2(n43708), .ZN(
        n43711) );
  INV_X1 U11179 ( .I(n21360), .ZN(n43985) );
  NAND2_X1 U29340 ( .A1(n9377), .A2(n61858), .ZN(n20904) );
  NOR2_X1 U11108 ( .A1(n9634), .A2(n43027), .ZN(n9858) );
  NAND3_X1 U36900 ( .A1(n21326), .A2(n10004), .A3(n9914), .ZN(n41341) );
  AOI22_X1 U12746 ( .A1(n42809), .A2(n7048), .B1(n15250), .B2(n42973), .ZN(
        n7386) );
  CLKBUF_X1 U11190 ( .I(n42387), .Z(n4805) );
  INV_X1 U51536 ( .I(n43173), .ZN(n43176) );
  CLKBUF_X4 U16437 ( .I(n46587), .Z(n23905) );
  BUF_X2 U9297 ( .I(n13180), .Z(n13179) );
  CLKBUF_X2 U9984 ( .I(n44098), .Z(n6204) );
  INV_X1 U16417 ( .I(n13884), .ZN(n4556) );
  INV_X1 U16386 ( .I(n46305), .ZN(n2723) );
  CLKBUF_X4 U1365 ( .I(n46674), .Z(n5180) );
  BUF_X2 U16329 ( .I(n20854), .Z(n7506) );
  INV_X2 U21939 ( .I(n47467), .ZN(n3368) );
  INV_X2 U11003 ( .I(n48564), .ZN(n47127) );
  INV_X2 U4129 ( .I(n48612), .ZN(n14419) );
  BUF_X2 U12690 ( .I(n48145), .Z(n23185) );
  BUF_X2 U16275 ( .I(n44435), .Z(n47266) );
  CLKBUF_X2 U6457 ( .I(n48612), .Z(n571) );
  OAI21_X1 U53468 ( .A1(n7186), .A2(n60390), .B(n48134), .ZN(n48137) );
  NOR3_X1 U12625 ( .A1(n23407), .A2(n45493), .A3(n13258), .ZN(n7191) );
  INV_X2 U1133 ( .I(n62308), .ZN(n47544) );
  INV_X1 U16249 ( .I(n11627), .ZN(n10653) );
  INV_X1 U1187 ( .I(n45779), .ZN(n47029) );
  NOR2_X1 U29467 ( .A1(n47289), .A2(n9505), .ZN(n45553) );
  NAND2_X1 U10950 ( .A1(n47544), .A2(n47180), .ZN(n46362) );
  OR3_X1 U7847 ( .A1(n45479), .A2(n9331), .A3(n65275), .Z(n1087) );
  NAND2_X1 U52529 ( .A1(n45504), .A2(n46070), .ZN(n45509) );
  NOR2_X1 U16080 ( .A1(n46105), .A2(n17318), .ZN(n4448) );
  INV_X1 U37038 ( .I(n45527), .ZN(n47026) );
  NAND2_X1 U10926 ( .A1(n45741), .A2(n47476), .ZN(n2069) );
  AOI21_X1 U12656 ( .A1(n64791), .A2(n48642), .B(n64922), .ZN(n46564) );
  OAI21_X1 U33974 ( .A1(n47207), .A2(n48124), .B(n60386), .ZN(n14487) );
  AOI21_X1 U15895 ( .A1(n5298), .A2(n5297), .B(n59687), .ZN(n46932) );
  NAND2_X1 U53132 ( .A1(n47536), .A2(n48594), .ZN(n47006) );
  BUF_X4 U944 ( .I(n47444), .Z(n49610) );
  AND4_X2 U12514 ( .A1(n9332), .A2(n9227), .A3(n9226), .A4(n47722), .Z(n9225)
         );
  CLKBUF_X2 U12490 ( .I(n48868), .Z(n4815) );
  BUF_X4 U8576 ( .I(n46850), .Z(n12580) );
  CLKBUF_X4 U15600 ( .I(n17994), .Z(n13038) );
  INV_X1 U15711 ( .I(n49923), .ZN(n6575) );
  INV_X1 U12462 ( .I(n24613), .ZN(n13122) );
  AOI21_X1 U53479 ( .A1(n1291), .A2(n13024), .B(n50334), .ZN(n48170) );
  INV_X1 U15446 ( .I(n19096), .ZN(n20595) );
  AOI22_X1 U8543 ( .A1(n47993), .A2(n50011), .B1(n47992), .B2(n49339), .ZN(
        n48001) );
  OAI22_X1 U15473 ( .A1(n49696), .A2(n49695), .B1(n64), .B2(n49698), .ZN(
        n49707) );
  AOI21_X1 U53410 ( .A1(n48721), .A2(n58861), .B(n1471), .ZN(n47954) );
  AND3_X1 U7917 ( .A1(n49527), .A2(n2956), .A3(n10637), .Z(n1136) );
  CLKBUF_X4 U4382 ( .I(n22678), .Z(n12985) );
  BUF_X2 U15175 ( .I(n51671), .Z(n7229) );
  INV_X1 U12323 ( .I(n50550), .ZN(n12874) );
  INV_X2 U12343 ( .I(n52360), .ZN(n8569) );
  CLKBUF_X2 U15153 ( .I(n18715), .Z(n10594) );
  BUF_X4 U9167 ( .I(n50436), .Z(n15447) );
  BUF_X4 U27803 ( .I(n10502), .Z(n7711) );
  INV_X1 U42995 ( .I(n50111), .ZN(n54037) );
  INV_X1 U12309 ( .I(n19639), .ZN(n53232) );
  CLKBUF_X2 U6450 ( .I(n53377), .Z(n23401) );
  INV_X1 U34283 ( .I(n19716), .ZN(n51529) );
  BUF_X4 U12305 ( .I(n13232), .Z(n23248) );
  CLKBUF_X2 U9155 ( .I(n24455), .Z(n4194) );
  CLKBUF_X2 U12287 ( .I(n56593), .Z(n7274) );
  BUF_X2 U5644 ( .I(n53859), .Z(n4480) );
  CLKBUF_X4 U8508 ( .I(n53858), .Z(n4481) );
  CLKBUF_X2 U6410 ( .I(n54058), .Z(n550) );
  NAND2_X1 U56523 ( .A1(n56390), .A2(n51264), .ZN(n56391) );
  NAND2_X1 U35580 ( .A1(n56359), .A2(n56370), .ZN(n20599) );
  NAND2_X1 U14879 ( .A1(n53241), .A2(n1325), .ZN(n53234) );
  INV_X2 U423 ( .I(n54047), .ZN(n54033) );
  CLKBUF_X2 U14798 ( .I(n9136), .Z(n7159) );
  AOI21_X1 U267 ( .A1(n1150), .A2(n51889), .B(n57203), .ZN(n4863) );
  AOI21_X1 U55293 ( .A1(n53008), .A2(n53007), .B(n53006), .ZN(n53010) );
  NAND2_X1 U36246 ( .A1(n54692), .A2(n54694), .ZN(n22124) );
  CLKBUF_X4 U8253 ( .I(n56341), .Z(n23318) );
  NAND2_X1 U21467 ( .A1(n3021), .A2(n14708), .ZN(n23631) );
  NAND2_X1 U4034 ( .A1(n54742), .A2(n54771), .ZN(n54665) );
  INV_X1 U12131 ( .I(n3937), .ZN(n57110) );
  NOR2_X2 U4105 ( .A1(n43889), .A2(n7516), .ZN(n43140) );
  INV_X2 U3424 ( .I(n27661), .ZN(n28485) );
  BUF_X4 U4910 ( .I(n34119), .Z(n139) );
  BUF_X4 U41006 ( .I(n28244), .Z(n21158) );
  AOI22_X2 U10896 ( .A1(n46822), .A2(n16004), .B1(n12268), .B2(n21451), .ZN(
        n21450) );
  NAND2_X2 U25865 ( .A1(n21301), .A2(n6215), .ZN(n26573) );
  NOR2_X2 U175 ( .A1(n13504), .A2(n25267), .ZN(n13503) );
  INV_X2 U3433 ( .I(n25202), .ZN(n29142) );
  INV_X2 U3437 ( .I(n61918), .ZN(n1894) );
  INV_X1 U42117 ( .I(n28362), .ZN(n26606) );
  INV_X2 U3319 ( .I(n3617), .ZN(n29152) );
  BUF_X2 U9750 ( .I(n29154), .Z(n7499) );
  NAND2_X1 U39846 ( .A1(n28639), .A2(n26912), .ZN(n20070) );
  NOR2_X1 U42612 ( .A1(n23568), .A2(n3697), .ZN(n27378) );
  NAND2_X1 U44244 ( .A1(n24391), .A2(n27478), .ZN(n27482) );
  INV_X1 U3369 ( .I(n5218), .ZN(n27217) );
  NAND2_X1 U42816 ( .A1(n28811), .A2(n26456), .ZN(n26994) );
  BUF_X2 U42592 ( .I(n29133), .Z(n23591) );
  INV_X1 U44110 ( .I(n29371), .ZN(n28808) );
  INV_X1 U44070 ( .I(n26407), .ZN(n26811) );
  BUF_X2 U19857 ( .I(n26791), .Z(n28447) );
  NAND2_X1 U3411 ( .A1(n23649), .A2(n26791), .ZN(n4869) );
  INV_X1 U10556 ( .I(n28067), .ZN(n24498) );
  OAI21_X1 U44717 ( .A1(n28610), .A2(n28452), .B(n28436), .ZN(n27644) );
  INV_X2 U6053 ( .I(n7110), .ZN(n25858) );
  INV_X1 U44404 ( .I(n27482), .ZN(n27546) );
  INV_X1 U7486 ( .I(n28224), .ZN(n14102) );
  INV_X1 U5743 ( .I(n29306), .ZN(n1439) );
  INV_X2 U33760 ( .I(n22514), .ZN(n15358) );
  NAND2_X1 U12029 ( .A1(n28587), .A2(n26061), .ZN(n19643) );
  NAND2_X1 U44744 ( .A1(n28675), .A2(n12739), .ZN(n29605) );
  BUF_X2 U9035 ( .I(n60816), .Z(n24001) );
  BUF_X2 U3423 ( .I(n26278), .Z(n22408) );
  NAND2_X1 U29506 ( .A1(n13955), .A2(n7760), .ZN(n27851) );
  NOR2_X1 U39477 ( .A1(n28025), .A2(n22044), .ZN(n28275) );
  NOR2_X1 U9038 ( .A1(n27232), .A2(n27479), .ZN(n25090) );
  INV_X2 U24560 ( .I(n29660), .ZN(n29652) );
  NOR2_X1 U41473 ( .A1(n60505), .A2(n28240), .ZN(n28070) );
  OR2_X1 U4734 ( .A1(n27381), .A2(n28067), .Z(n16042) );
  INV_X1 U32026 ( .I(n14439), .ZN(n19122) );
  INV_X1 U29419 ( .I(n9473), .ZN(n25786) );
  NOR2_X1 U44364 ( .A1(n28675), .A2(n29608), .ZN(n29614) );
  NOR2_X1 U6973 ( .A1(n28517), .A2(n27851), .ZN(n28508) );
  NAND2_X1 U6960 ( .A1(n62406), .A2(n28217), .ZN(n29117) );
  NAND2_X1 U8419 ( .A1(n28279), .A2(n28270), .ZN(n8777) );
  NOR2_X1 U6992 ( .A1(n27451), .A2(n27450), .ZN(n29307) );
  INV_X1 U12009 ( .I(n28540), .ZN(n1883) );
  OAI21_X1 U40125 ( .A1(n28852), .A2(n9987), .B(n23797), .ZN(n28156) );
  NOR2_X1 U19651 ( .A1(n28648), .A2(n28651), .ZN(n28184) );
  NAND2_X1 U14220 ( .A1(n27123), .A2(n15156), .ZN(n26565) );
  INV_X1 U22902 ( .I(n21086), .ZN(n28257) );
  INV_X1 U11999 ( .I(n28301), .ZN(n28306) );
  NOR2_X1 U44502 ( .A1(n27142), .A2(n28049), .ZN(n28335) );
  NAND2_X1 U14182 ( .A1(n29381), .A2(n2066), .ZN(n29658) );
  NAND2_X1 U9018 ( .A1(n20678), .A2(n28813), .ZN(n6759) );
  NOR2_X1 U14235 ( .A1(n10754), .A2(n29661), .ZN(n8072) );
  NAND2_X1 U27643 ( .A1(n29174), .A2(n26407), .ZN(n28557) );
  NOR2_X1 U6965 ( .A1(n28534), .A2(n23508), .ZN(n27869) );
  NAND2_X1 U31587 ( .A1(n23352), .A2(n24350), .ZN(n11225) );
  INV_X1 U44083 ( .I(n26835), .ZN(n27712) );
  INV_X1 U3208 ( .I(n28275), .ZN(n7719) );
  NOR2_X1 U3316 ( .A1(n26339), .A2(n28311), .ZN(n28308) );
  INV_X1 U10540 ( .I(n27931), .ZN(n29137) );
  INV_X1 U3228 ( .I(n28855), .ZN(n28163) );
  NAND3_X1 U3209 ( .A1(n29643), .A2(n29644), .A3(n6345), .ZN(n21203) );
  NOR2_X1 U3569 ( .A1(n1567), .A2(n28175), .ZN(n27693) );
  INV_X1 U3360 ( .I(n29662), .ZN(n29382) );
  INV_X1 U21362 ( .I(n28036), .ZN(n27098) );
  INV_X1 U3332 ( .I(n28410), .ZN(n28401) );
  INV_X1 U10589 ( .I(n29356), .ZN(n28878) );
  INV_X1 U34052 ( .I(n61643), .ZN(n14583) );
  INV_X1 U20914 ( .I(n27374), .ZN(n23665) );
  NOR2_X1 U44509 ( .A1(n27142), .A2(n27138), .ZN(n27140) );
  NOR2_X1 U14189 ( .A1(n28174), .A2(n29609), .ZN(n26878) );
  AOI21_X1 U8990 ( .A1(n28509), .A2(n28508), .B(n28507), .ZN(n28512) );
  INV_X1 U19616 ( .I(n28188), .ZN(n27679) );
  NOR2_X1 U35300 ( .A1(n28673), .A2(n28176), .ZN(n27314) );
  NAND3_X1 U26593 ( .A1(n12705), .A2(n26714), .A3(n6913), .ZN(n12706) );
  NOR2_X1 U38552 ( .A1(n18006), .A2(n27664), .ZN(n26397) );
  INV_X1 U19754 ( .I(n27126), .ZN(n25392) );
  AOI21_X1 U4610 ( .A1(n25735), .A2(n27389), .B(n25734), .ZN(n25737) );
  INV_X1 U45311 ( .I(n29358), .ZN(n29361) );
  INV_X1 U19700 ( .I(n26217), .ZN(n16811) );
  NAND2_X1 U14176 ( .A1(n2342), .A2(n29178), .ZN(n29183) );
  NOR2_X1 U3269 ( .A1(n21956), .A2(n29118), .ZN(n29125) );
  NAND2_X1 U5375 ( .A1(n3087), .A2(n8613), .ZN(n29130) );
  INV_X2 U28564 ( .I(n29118), .ZN(n27970) );
  INV_X1 U12030 ( .I(n18848), .ZN(n26736) );
  NOR2_X1 U6957 ( .A1(n22351), .A2(n29178), .ZN(n27273) );
  INV_X1 U19685 ( .I(n28137), .ZN(n28828) );
  AOI22_X1 U6596 ( .A1(n29602), .A2(n29618), .B1(n27313), .B2(n29603), .ZN(
        n27317) );
  AOI21_X1 U36588 ( .A1(n27255), .A2(n19359), .B(n27875), .ZN(n26002) );
  NAND3_X1 U44915 ( .A1(n28828), .A2(n28138), .A3(n60894), .ZN(n28139) );
  NOR2_X1 U14053 ( .A1(n11066), .A2(n11065), .ZN(n20476) );
  NOR3_X1 U44963 ( .A1(n28347), .A2(n296), .A3(n28346), .ZN(n28357) );
  NOR2_X1 U29693 ( .A1(n27970), .A2(n24080), .ZN(n27271) );
  INV_X1 U11950 ( .I(n28015), .ZN(n21947) );
  NAND2_X1 U3274 ( .A1(n555), .A2(n61004), .ZN(n19565) );
  NOR2_X1 U44312 ( .A1(n61169), .A2(n26813), .ZN(n26814) );
  NOR2_X1 U44809 ( .A1(n27808), .A2(n27812), .ZN(n27809) );
  OAI21_X1 U25270 ( .A1(n61820), .A2(n26445), .B(n15684), .ZN(n26450) );
  NAND2_X1 U19687 ( .A1(n29714), .A2(n28625), .ZN(n28626) );
  NOR2_X1 U19479 ( .A1(n17882), .A2(n17881), .ZN(n17880) );
  INV_X1 U12004 ( .I(n6519), .ZN(n7023) );
  NAND2_X1 U19421 ( .A1(n24816), .A2(n28237), .ZN(n24812) );
  NAND2_X1 U4979 ( .A1(n28885), .A2(n28884), .ZN(n8362) );
  OAI22_X1 U8999 ( .A1(n29652), .A2(n58955), .B1(n29382), .B2(n20126), .ZN(
        n10148) );
  OAI22_X1 U19495 ( .A1(n26814), .A2(n29177), .B1(n1355), .B2(n20782), .ZN(
        n26818) );
  INV_X1 U6698 ( .I(n28347), .ZN(n27202) );
  NAND3_X1 U3533 ( .A1(n2656), .A2(n2655), .A3(n26809), .ZN(n2654) );
  OAI21_X1 U6060 ( .A1(n27708), .A2(n26416), .B(n28509), .ZN(n26417) );
  NOR3_X1 U3173 ( .A1(n29190), .A2(n29185), .A3(n23892), .ZN(n24970) );
  OAI21_X1 U14045 ( .A1(n27202), .A2(n27201), .B(n16021), .ZN(n24774) );
  OAI21_X1 U3165 ( .A1(n29646), .A2(n29645), .B(n434), .ZN(n31156) );
  BUF_X2 U40718 ( .I(n27003), .Z(n30430) );
  AOI21_X1 U44834 ( .A1(n27883), .A2(n7354), .B(n27882), .ZN(n27884) );
  BUF_X4 U25464 ( .I(n14767), .Z(n5768) );
  BUF_X2 U3708 ( .I(n19624), .Z(n19590) );
  BUF_X2 U3150 ( .I(n31051), .Z(n18839) );
  INV_X2 U30884 ( .I(n29232), .ZN(n30817) );
  INV_X1 U8206 ( .I(n21713), .ZN(n13176) );
  INV_X1 U37633 ( .I(n27003), .ZN(n31086) );
  INV_X1 U10504 ( .I(n28932), .ZN(n22496) );
  BUF_X4 U21141 ( .I(n6149), .Z(n2795) );
  INV_X1 U3069 ( .I(n29862), .ZN(n29523) );
  INV_X1 U11817 ( .I(n30252), .ZN(n1848) );
  INV_X1 U8948 ( .I(n18880), .ZN(n30747) );
  OR2_X1 U8163 ( .A1(n25669), .A2(n30347), .Z(n29585) );
  CLKBUF_X2 U10466 ( .I(n29232), .Z(n24123) );
  INV_X4 U3168 ( .I(n19701), .ZN(n14217) );
  CLKBUF_X2 U3021 ( .I(Key[111]), .Z(n55368) );
  NAND2_X1 U25975 ( .A1(n6317), .A2(n31261), .ZN(n31159) );
  INV_X2 U8321 ( .I(n29457), .ZN(n20755) );
  CLKBUF_X2 U4866 ( .I(n29801), .Z(n131) );
  BUF_X2 U8981 ( .I(n29795), .Z(n23370) );
  INV_X2 U9684 ( .I(n19624), .ZN(n20747) );
  INV_X1 U3084 ( .I(n26740), .ZN(n30242) );
  INV_X2 U3057 ( .I(n30664), .ZN(n25052) );
  INV_X2 U3141 ( .I(n24056), .ZN(n31038) );
  INV_X1 U5497 ( .I(n29748), .ZN(n18128) );
  NOR2_X1 U8342 ( .A1(n29794), .A2(n25241), .ZN(n29014) );
  INV_X2 U3125 ( .I(n25051), .ZN(n30760) );
  INV_X1 U32457 ( .I(n12443), .ZN(n30501) );
  NAND2_X1 U3060 ( .A1(n25051), .A2(n30761), .ZN(n22696) );
  BUF_X2 U3122 ( .I(n31247), .Z(n9654) );
  NAND2_X1 U9654 ( .A1(n29034), .A2(n17872), .ZN(n30176) );
  INV_X1 U3090 ( .I(n31159), .ZN(n1853) );
  INV_X1 U19192 ( .I(n21964), .ZN(n18326) );
  INV_X1 U11842 ( .I(n31127), .ZN(n1844) );
  NOR2_X1 U5492 ( .A1(n23397), .A2(n30322), .ZN(n29984) );
  NAND2_X1 U19274 ( .A1(n26957), .A2(n60895), .ZN(n28582) );
  INV_X1 U35934 ( .I(n31041), .ZN(n30707) );
  NAND2_X1 U41950 ( .A1(n31045), .A2(n30059), .ZN(n30161) );
  NOR2_X1 U45057 ( .A1(n28683), .A2(n58273), .ZN(n30739) );
  NOR2_X1 U3116 ( .A1(n15808), .A2(n27305), .ZN(n11565) );
  INV_X2 U3148 ( .I(n19830), .ZN(n1872) );
  NAND2_X1 U7009 ( .A1(n9197), .A2(n25241), .ZN(n27915) );
  NOR2_X1 U3105 ( .A1(n24564), .A2(n20391), .ZN(n30631) );
  NOR2_X1 U3035 ( .A1(n1436), .A2(n23008), .ZN(n2042) );
  INV_X2 U33418 ( .I(n23168), .ZN(n15126) );
  NAND2_X1 U29970 ( .A1(n30311), .A2(n7426), .ZN(n30004) );
  INV_X4 U9681 ( .I(n29773), .ZN(n1351) );
  NOR2_X1 U9678 ( .A1(n57437), .A2(n23955), .ZN(n31093) );
  INV_X2 U5988 ( .I(n20025), .ZN(n25978) );
  INV_X1 U2926 ( .I(n29442), .ZN(n29909) );
  NOR2_X1 U2999 ( .A1(n18198), .A2(n30680), .ZN(n29205) );
  NAND2_X1 U21594 ( .A1(n8218), .A2(n13731), .ZN(n12612) );
  NOR2_X1 U22058 ( .A1(n9654), .A2(n12893), .ZN(n3486) );
  NOR2_X1 U26105 ( .A1(n30760), .A2(n10888), .ZN(n31216) );
  NAND2_X1 U2975 ( .A1(n17745), .A2(n30781), .ZN(n29545) );
  NOR2_X1 U45646 ( .A1(n21176), .A2(n30702), .ZN(n30700) );
  NAND2_X1 U32621 ( .A1(n1316), .A2(n23918), .ZN(n31137) );
  NAND2_X1 U19313 ( .A1(n31224), .A2(n15738), .ZN(n28894) );
  NOR2_X1 U31393 ( .A1(n59046), .A2(n25052), .ZN(n30663) );
  NAND2_X1 U44940 ( .A1(n19590), .A2(n31105), .ZN(n31118) );
  INV_X1 U10483 ( .I(n17872), .ZN(n30689) );
  NOR2_X1 U2997 ( .A1(n19701), .A2(n1432), .ZN(n19535) );
  NOR2_X1 U39549 ( .A1(n1433), .A2(n29835), .ZN(n28754) );
  INV_X2 U10490 ( .I(n15727), .ZN(n1558) );
  NOR3_X1 U45168 ( .A1(n30294), .A2(n57559), .A3(n1317), .ZN(n28925) );
  NOR2_X1 U3730 ( .A1(n30663), .A2(n61215), .ZN(n10923) );
  NAND2_X1 U2953 ( .A1(n25978), .A2(n58560), .ZN(n30023) );
  NAND2_X1 U6999 ( .A1(n15126), .A2(n20859), .ZN(n3098) );
  NAND2_X1 U45581 ( .A1(n23799), .A2(n25052), .ZN(n30008) );
  NAND2_X1 U8917 ( .A1(n30887), .A2(n30883), .ZN(n30500) );
  INV_X1 U3009 ( .I(n17495), .ZN(n28794) );
  NAND2_X1 U44445 ( .A1(n31080), .A2(n58931), .ZN(n28570) );
  INV_X1 U3011 ( .I(n11565), .ZN(n13766) );
  INV_X1 U5040 ( .I(n29863), .ZN(n173) );
  INV_X1 U6504 ( .I(n14350), .ZN(n4993) );
  AOI21_X1 U9670 ( .A1(n20378), .A2(n1432), .B(n19701), .ZN(n13032) );
  NAND2_X1 U3479 ( .A1(n6090), .A2(n30396), .ZN(n6089) );
  INV_X1 U3007 ( .I(n29490), .ZN(n31102) );
  NAND2_X1 U2952 ( .A1(n20025), .A2(n13087), .ZN(n30019) );
  NAND2_X1 U32268 ( .A1(n8602), .A2(n22014), .ZN(n12165) );
  NAND2_X1 U38644 ( .A1(n21886), .A2(n17745), .ZN(n20178) );
  NAND2_X1 U3025 ( .A1(n30679), .A2(n22496), .ZN(n30678) );
  NOR2_X1 U38555 ( .A1(n29905), .A2(n17590), .ZN(n28972) );
  NOR2_X1 U21691 ( .A1(n30455), .A2(n11425), .ZN(n30361) );
  NOR2_X1 U34180 ( .A1(n14739), .A2(n15205), .ZN(n30545) );
  NOR2_X1 U3038 ( .A1(n8218), .A2(n9865), .ZN(n11206) );
  NOR2_X1 U29969 ( .A1(n1875), .A2(n30004), .ZN(n30006) );
  NAND2_X1 U13904 ( .A1(n30757), .A2(n59046), .ZN(n31223) );
  NAND2_X1 U21692 ( .A1(n30455), .A2(n21095), .ZN(n29430) );
  BUF_X2 U10624 ( .I(n61447), .Z(n26010) );
  NAND2_X1 U29144 ( .A1(n9153), .A2(n30430), .ZN(n31089) );
  NAND2_X1 U2924 ( .A1(n20025), .A2(n21478), .ZN(n29733) );
  NAND2_X1 U45484 ( .A1(n29794), .A2(n131), .ZN(n29800) );
  INV_X1 U10460 ( .I(n27922), .ZN(n30524) );
  INV_X1 U7391 ( .I(n27905), .ZN(n31182) );
  NAND2_X1 U45858 ( .A1(n23799), .A2(n31224), .ZN(n30665) );
  NOR2_X1 U27310 ( .A1(n59046), .A2(n1875), .ZN(n31220) );
  INV_X1 U19347 ( .I(n20859), .ZN(n8378) );
  AOI22_X1 U40653 ( .A1(n28942), .A2(n29780), .B1(n28943), .B2(n29778), .ZN(
        n28760) );
  OAI22_X1 U11800 ( .A1(n1847), .A2(n30634), .B1(n9979), .B2(n28681), .ZN(
        n3443) );
  OAI21_X1 U13790 ( .A1(n29840), .A2(n28995), .B(n7979), .ZN(n14850) );
  AOI22_X1 U11796 ( .A1(n19697), .A2(n31120), .B1(n31119), .B2(n57437), .ZN(
        n14275) );
  OAI21_X1 U41191 ( .A1(n29879), .A2(n21478), .B(n29878), .ZN(n21703) );
  OAI21_X1 U9638 ( .A1(n61162), .A2(n6714), .B(n24728), .ZN(n5861) );
  AOI21_X1 U44841 ( .A1(n24777), .A2(n29904), .B(n27906), .ZN(n27909) );
  NAND2_X1 U35417 ( .A1(n28772), .A2(n23317), .ZN(n30721) );
  NAND3_X1 U44447 ( .A1(n27005), .A2(n28570), .A3(n27004), .ZN(n27006) );
  NAND2_X1 U36780 ( .A1(n23111), .A2(n23370), .ZN(n29013) );
  AOI21_X1 U4387 ( .A1(n29098), .A2(n173), .B(n29096), .ZN(n29103) );
  OAI21_X1 U13946 ( .A1(n31110), .A2(n26084), .B(n1868), .ZN(n31095) );
  NAND2_X1 U19231 ( .A1(n16504), .A2(n1552), .ZN(n8959) );
  NAND2_X1 U2897 ( .A1(n770), .A2(n7040), .ZN(n30222) );
  NAND2_X1 U45289 ( .A1(n30294), .A2(n29579), .ZN(n29573) );
  INV_X1 U4564 ( .I(n61048), .ZN(n29428) );
  INV_X1 U3003 ( .I(n30077), .ZN(n1554) );
  INV_X1 U9636 ( .I(n30545), .ZN(n15147) );
  INV_X1 U6163 ( .I(n4196), .ZN(n30442) );
  INV_X1 U36016 ( .I(n30126), .ZN(n29774) );
  NAND3_X1 U29824 ( .A1(n16388), .A2(n19697), .A3(n14350), .ZN(n19696) );
  NAND2_X1 U19135 ( .A1(n30327), .A2(n30326), .ZN(n23537) );
  OAI21_X1 U45871 ( .A1(n30708), .A2(n31029), .B(n30707), .ZN(n30712) );
  NOR3_X1 U45650 ( .A1(n30153), .A2(n30152), .A3(n30151), .ZN(n30154) );
  NAND2_X1 U13977 ( .A1(n30680), .A2(n30679), .ZN(n6537) );
  OAI21_X1 U11782 ( .A1(n3934), .A2(n29733), .B(n3933), .ZN(n5493) );
  AOI21_X1 U36791 ( .A1(n26844), .A2(n9618), .B(n17605), .ZN(n20316) );
  OAI21_X1 U19034 ( .A1(n15138), .A2(n6038), .B(n30676), .ZN(n15137) );
  NAND2_X1 U45436 ( .A1(n22799), .A2(n5631), .ZN(n29737) );
  NOR3_X1 U11767 ( .A1(n17626), .A2(n17628), .A3(n29035), .ZN(n4439) );
  NAND2_X1 U18898 ( .A1(n14745), .A2(n25399), .ZN(n8708) );
  NAND2_X1 U13827 ( .A1(n6178), .A2(n6585), .ZN(n6584) );
  AOI22_X1 U45440 ( .A1(n29743), .A2(n29748), .B1(n21886), .B2(n30782), .ZN(
        n29753) );
  NOR2_X1 U45347 ( .A1(n29911), .A2(n29443), .ZN(n29444) );
  NAND3_X1 U19178 ( .A1(n31223), .A2(n57806), .A3(n23799), .ZN(n24221) );
  AOI21_X1 U3456 ( .A1(n27424), .A2(n30261), .B(n30260), .ZN(n27427) );
  NAND2_X1 U13771 ( .A1(n10235), .A2(n31121), .ZN(n6405) );
  NAND3_X1 U11779 ( .A1(n6178), .A2(n22513), .A3(n4051), .ZN(n29510) );
  AOI22_X1 U2869 ( .A1(n3820), .A2(n30362), .B1(n13628), .B2(n29061), .ZN(
        n29068) );
  NOR3_X1 U4628 ( .A1(n30435), .A2(n30437), .A3(n30436), .ZN(n4585) );
  NAND3_X1 U40516 ( .A1(n30874), .A2(n30873), .A3(n25013), .ZN(n30881) );
  INV_X1 U25014 ( .I(n5726), .ZN(n32542) );
  INV_X2 U2819 ( .I(n15982), .ZN(n21094) );
  OAI21_X1 U35458 ( .A1(n18634), .A2(n18637), .B(n33239), .ZN(n17544) );
  INV_X1 U5662 ( .I(n61152), .ZN(n31917) );
  BUF_X2 U2836 ( .I(n32542), .Z(n5727) );
  BUF_X2 U8078 ( .I(n30034), .Z(n11265) );
  BUF_X2 U33606 ( .I(n24746), .Z(n13956) );
  BUF_X2 U13761 ( .I(n32301), .Z(n21083) );
  BUF_X2 U8895 ( .I(n21885), .Z(n21884) );
  BUF_X2 U18879 ( .I(n32044), .Z(n23090) );
  INV_X1 U18867 ( .I(n32267), .ZN(n1824) );
  INV_X1 U9607 ( .I(n31439), .ZN(n31365) );
  BUF_X2 U26345 ( .I(n33139), .Z(n6701) );
  INV_X2 U29868 ( .I(n24471), .ZN(n33158) );
  INV_X1 U2829 ( .I(n30229), .ZN(n31706) );
  INV_X1 U7564 ( .I(n30833), .ZN(n31925) );
  INV_X1 U28306 ( .I(n31863), .ZN(n32640) );
  INV_X1 U8090 ( .I(n24839), .ZN(n32540) );
  BUF_X2 U13744 ( .I(n31336), .Z(n16884) );
  BUF_X2 U34262 ( .I(n14867), .Z(n14866) );
  INV_X1 U21686 ( .I(n31385), .ZN(n17914) );
  INV_X1 U2811 ( .I(n15725), .ZN(n30946) );
  INV_X2 U22310 ( .I(n24258), .ZN(n32354) );
  INV_X1 U18872 ( .I(n32388), .ZN(n1827) );
  INV_X1 U2784 ( .I(n6611), .ZN(n7814) );
  INV_X1 U2787 ( .I(n33914), .ZN(n24822) );
  INV_X1 U24746 ( .I(n64417), .ZN(n5086) );
  INV_X2 U2759 ( .I(n21592), .ZN(n13942) );
  INV_X2 U34483 ( .I(n18524), .ZN(n18879) );
  INV_X2 U11689 ( .I(n24331), .ZN(n5472) );
  NOR2_X1 U25404 ( .A1(n32892), .A2(n32829), .ZN(n32891) );
  INV_X1 U7045 ( .I(n262), .ZN(n34130) );
  NAND2_X1 U34984 ( .A1(n25256), .A2(n20989), .ZN(n21731) );
  BUF_X2 U3882 ( .I(n34521), .Z(n2891) );
  INV_X2 U2668 ( .I(n35218), .ZN(n17401) );
  NOR2_X1 U47923 ( .A1(n33600), .A2(n33596), .ZN(n35694) );
  INV_X1 U29191 ( .I(n9330), .ZN(n17255) );
  NAND2_X1 U32388 ( .A1(n34950), .A2(n12354), .ZN(n32298) );
  INV_X2 U2678 ( .I(n13487), .ZN(n15018) );
  NOR2_X1 U43132 ( .A1(n65194), .A2(n34302), .ZN(n32945) );
  INV_X1 U4850 ( .I(n5250), .ZN(n33370) );
  INV_X1 U40441 ( .I(n34035), .ZN(n20507) );
  INV_X1 U31359 ( .I(n22333), .ZN(n25625) );
  INV_X1 U18704 ( .I(n34753), .ZN(n1802) );
  INV_X2 U11682 ( .I(n32435), .ZN(n34305) );
  NAND2_X1 U48289 ( .A1(n23354), .A2(n35301), .ZN(n35299) );
  INV_X1 U22615 ( .I(n5322), .ZN(n25632) );
  INV_X1 U2683 ( .I(n35229), .ZN(n35833) );
  INV_X1 U2712 ( .I(n7932), .ZN(n33465) );
  INV_X1 U10356 ( .I(n18077), .ZN(n1425) );
  INV_X2 U2679 ( .I(n61249), .ZN(n3023) );
  NAND2_X1 U5925 ( .A1(n21945), .A2(n15783), .ZN(n32796) );
  INV_X2 U5970 ( .I(n21945), .ZN(n33949) );
  NAND3_X1 U37972 ( .A1(n34766), .A2(n59724), .A3(n34302), .ZN(n32432) );
  OAI22_X1 U37872 ( .A1(n57200), .A2(n25563), .B1(n24286), .B2(n35674), .ZN(
        n33579) );
  NOR2_X1 U29037 ( .A1(n33362), .A2(n60633), .ZN(n33681) );
  NAND2_X1 U13688 ( .A1(n34623), .A2(n34622), .ZN(n25175) );
  AOI22_X1 U13537 ( .A1(n33778), .A2(n10016), .B1(n34273), .B2(n10175), .ZN(
        n12266) );
  INV_X2 U2615 ( .I(n33583), .ZN(n33802) );
  INV_X1 U47544 ( .I(n34137), .ZN(n34133) );
  INV_X1 U8854 ( .I(n34448), .ZN(n35659) );
  INV_X2 U21656 ( .I(n34188), .ZN(n20607) );
  NOR2_X1 U8279 ( .A1(n34634), .A2(n9130), .ZN(n23774) );
  BUF_X2 U2707 ( .I(n24522), .Z(n7534) );
  NAND2_X1 U20827 ( .A1(n139), .A2(n2695), .ZN(n33947) );
  NAND2_X1 U3949 ( .A1(n25657), .A2(n34632), .ZN(n34641) );
  BUF_X2 U4664 ( .I(n16402), .Z(n77) );
  NAND2_X1 U3575 ( .A1(n15184), .A2(n34253), .ZN(n34254) );
  INV_X1 U13560 ( .I(n14156), .ZN(n34217) );
  NOR2_X1 U2628 ( .A1(n1545), .A2(n3947), .ZN(n32965) );
  NAND2_X1 U2613 ( .A1(n15545), .A2(n35241), .ZN(n35654) );
  INV_X1 U5892 ( .I(n2122), .ZN(n34276) );
  INV_X1 U29194 ( .I(n9329), .ZN(n35200) );
  INV_X1 U18690 ( .I(n34056), .ZN(n7173) );
  NAND3_X1 U47826 ( .A1(n57172), .A2(n33372), .A3(n33371), .ZN(n33381) );
  NAND2_X1 U13582 ( .A1(n9030), .A2(n15815), .ZN(n33793) );
  NOR2_X1 U9576 ( .A1(n31358), .A2(n1813), .ZN(n8401) );
  NAND2_X1 U8276 ( .A1(n33624), .A2(n23086), .ZN(n33379) );
  AOI21_X1 U18325 ( .A1(n12266), .A2(n33779), .B(n12776), .ZN(n12816) );
  OR2_X1 U26900 ( .A1(n33096), .A2(n15298), .Z(n33347) );
  NOR2_X1 U18597 ( .A1(n262), .A2(n18908), .ZN(n18907) );
  NAND2_X1 U37146 ( .A1(n60579), .A2(n34962), .ZN(n34963) );
  INV_X1 U18446 ( .I(n32948), .ZN(n16678) );
  NAND2_X1 U2539 ( .A1(n34248), .A2(n34719), .ZN(n34249) );
  OAI21_X1 U4616 ( .A1(n33674), .A2(n33673), .B(n23351), .ZN(n33679) );
  INV_X1 U13683 ( .I(n4231), .ZN(n35679) );
  INV_X1 U41084 ( .I(n33993), .ZN(n32890) );
  NAND2_X1 U2535 ( .A1(n33499), .A2(n33730), .ZN(n34979) );
  AOI21_X1 U48434 ( .A1(n57986), .A2(n24286), .B(n35212), .ZN(n35213) );
  INV_X1 U18549 ( .I(n33117), .ZN(n33369) );
  NOR2_X1 U2558 ( .A1(n21020), .A2(n59626), .ZN(n32899) );
  NOR2_X1 U13691 ( .A1(n31358), .A2(n61249), .ZN(n33454) );
  NOR2_X1 U46498 ( .A1(n34613), .A2(n19512), .ZN(n33981) );
  NOR2_X1 U21473 ( .A1(n15786), .A2(n25251), .ZN(n34669) );
  NOR2_X1 U37145 ( .A1(n33448), .A2(n35038), .ZN(n24296) );
  INV_X1 U47586 ( .I(n34254), .ZN(n34352) );
  INV_X1 U18686 ( .I(n34164), .ZN(n34657) );
  INV_X1 U2662 ( .I(n10448), .ZN(n35807) );
  NOR2_X1 U36471 ( .A1(n16939), .A2(n7273), .ZN(n33101) );
  INV_X1 U47688 ( .I(n33342), .ZN(n33104) );
  NAND2_X1 U18586 ( .A1(n33454), .A2(n9687), .ZN(n9459) );
  NAND3_X1 U27799 ( .A1(n7710), .A2(n35842), .A3(n58048), .ZN(n16505) );
  BUF_X2 U13530 ( .I(n10866), .Z(n5874) );
  INV_X1 U18637 ( .I(n61896), .ZN(n18680) );
  NOR2_X1 U47853 ( .A1(n3467), .A2(n24083), .ZN(n33451) );
  AOI22_X1 U18354 ( .A1(n33400), .A2(n33399), .B1(n33657), .B2(n33398), .ZN(
        n25230) );
  NAND2_X1 U46095 ( .A1(n34041), .A2(n1798), .ZN(n33424) );
  NOR2_X1 U48612 ( .A1(n35847), .A2(n58048), .ZN(n35838) );
  NOR2_X1 U21927 ( .A1(n31725), .A2(n3363), .ZN(n4701) );
  INV_X1 U8838 ( .I(n18440), .ZN(n34304) );
  NAND2_X1 U13634 ( .A1(n34607), .A2(n60763), .ZN(n11762) );
  NAND2_X1 U2647 ( .A1(n34779), .A2(n19457), .ZN(n18508) );
  NAND2_X1 U2569 ( .A1(n8401), .A2(n34666), .ZN(n34516) );
  NOR2_X1 U9545 ( .A1(n10699), .A2(n24664), .ZN(n34180) );
  NAND2_X1 U36410 ( .A1(n33683), .A2(n34155), .ZN(n34148) );
  NOR2_X1 U21926 ( .A1(n1809), .A2(n3363), .ZN(n21322) );
  NOR2_X1 U47687 ( .A1(n33342), .A2(n61483), .ZN(n33099) );
  NAND4_X1 U48302 ( .A1(n34795), .A2(n23645), .A3(n60415), .A4(n560), .ZN(
        n34801) );
  NAND2_X1 U24099 ( .A1(n34218), .A2(n34217), .ZN(n18895) );
  NAND3_X1 U9564 ( .A1(n34797), .A2(n34796), .A3(n14112), .ZN(n34800) );
  NAND2_X1 U28173 ( .A1(n34179), .A2(n34178), .ZN(n8095) );
  INV_X1 U7051 ( .I(n33385), .ZN(n32703) );
  INV_X1 U4746 ( .I(n34516), .ZN(n99) );
  NOR2_X1 U41177 ( .A1(n34358), .A2(n34353), .ZN(n21461) );
  NOR2_X1 U25214 ( .A1(n63273), .A2(n4496), .ZN(n33302) );
  NAND2_X1 U18312 ( .A1(n11763), .A2(n11762), .ZN(n21111) );
  NOR2_X1 U13644 ( .A1(n35783), .A2(n11659), .ZN(n19996) );
  NAND3_X1 U13460 ( .A1(n32916), .A2(n32915), .A3(n19246), .ZN(n9279) );
  NAND2_X1 U47608 ( .A1(n33758), .A2(n12405), .ZN(n32969) );
  NAND2_X1 U13595 ( .A1(n34763), .A2(n34305), .ZN(n8114) );
  NAND2_X1 U18334 ( .A1(n25309), .A2(n35741), .ZN(n24460) );
  OR2_X1 U2499 ( .A1(n21217), .A2(n2695), .Z(n21216) );
  OAI21_X1 U10322 ( .A1(n35655), .A2(n35646), .B(n35654), .ZN(n35652) );
  NAND3_X1 U31939 ( .A1(n33757), .A2(n32964), .A3(n32963), .ZN(n32971) );
  NAND3_X1 U5204 ( .A1(n32703), .A2(n34135), .A3(n32702), .ZN(n32704) );
  NOR2_X1 U2507 ( .A1(n6526), .A2(n35627), .ZN(n35638) );
  NAND2_X1 U31347 ( .A1(n34334), .A2(n10866), .ZN(n33921) );
  OAI22_X1 U13455 ( .A1(n5388), .A2(n5386), .B1(n33988), .B2(n24160), .ZN(
        n7030) );
  NAND2_X1 U46502 ( .A1(n31531), .A2(n33980), .ZN(n31538) );
  INV_X4 U2448 ( .I(n35962), .ZN(n35548) );
  INV_X2 U4732 ( .I(n17202), .ZN(n36740) );
  NAND2_X1 U24112 ( .A1(n23503), .A2(n10601), .ZN(n35122) );
  BUF_X2 U3447 ( .I(n36377), .Z(n1785) );
  NAND2_X1 U17891 ( .A1(n36923), .A2(n35508), .ZN(n11561) );
  NAND2_X1 U48911 ( .A1(n36851), .A2(n36846), .ZN(n36837) );
  NAND2_X1 U11493 ( .A1(n37435), .A2(n8177), .ZN(n18427) );
  NAND2_X1 U7082 ( .A1(n25124), .A2(n36959), .ZN(n13557) );
  NOR2_X1 U29005 ( .A1(n10485), .A2(n36742), .ZN(n9013) );
  BUF_X2 U2410 ( .I(n36493), .Z(n22527) );
  INV_X1 U2391 ( .I(n1528), .ZN(n20147) );
  INV_X1 U21526 ( .I(n3057), .ZN(n36424) );
  INV_X2 U2295 ( .I(n32984), .ZN(n36553) );
  INV_X2 U11546 ( .I(n20908), .ZN(n37030) );
  INV_X2 U29457 ( .I(n24358), .ZN(n11558) );
  INV_X2 U13439 ( .I(n36483), .ZN(n18048) );
  INV_X2 U6750 ( .I(n33930), .ZN(n37319) );
  NOR2_X1 U41670 ( .A1(n36191), .A2(n36192), .ZN(n23387) );
  CLKBUF_X2 U18126 ( .I(n20571), .Z(n10254) );
  INV_X1 U8130 ( .I(n36207), .ZN(n36198) );
  INV_X1 U8823 ( .I(n36719), .ZN(n36721) );
  INV_X2 U2296 ( .I(n22254), .ZN(n36584) );
  NAND3_X1 U2321 ( .A1(n12652), .A2(n1338), .A3(n8438), .ZN(n18076) );
  NAND2_X1 U2344 ( .A1(n37455), .A2(n22801), .ZN(n37236) );
  NAND2_X1 U48339 ( .A1(n61517), .A2(n10849), .ZN(n35984) );
  NAND2_X1 U47601 ( .A1(n36574), .A2(n19364), .ZN(n32978) );
  INV_X1 U49078 ( .I(n37240), .ZN(n37245) );
  NAND2_X1 U22192 ( .A1(n14138), .A2(n25571), .ZN(n3590) );
  NOR2_X1 U2267 ( .A1(n36013), .A2(n36846), .ZN(n19553) );
  NOR2_X1 U10252 ( .A1(n10317), .A2(n10829), .ZN(n15940) );
  NOR2_X1 U18089 ( .A1(n35986), .A2(n652), .ZN(n35987) );
  INV_X1 U8798 ( .I(n35983), .ZN(n36708) );
  NAND2_X1 U36454 ( .A1(n61747), .A2(n36847), .ZN(n36856) );
  NAND2_X1 U38648 ( .A1(n36898), .A2(n60196), .ZN(n33124) );
  NAND2_X1 U47927 ( .A1(n36404), .A2(n35361), .ZN(n33606) );
  NAND2_X1 U38120 ( .A1(n16851), .A2(n36412), .ZN(n18602) );
  NOR2_X1 U7067 ( .A1(n36846), .A2(n4754), .ZN(n36669) );
  NAND2_X1 U2251 ( .A1(n32984), .A2(n1339), .ZN(n36092) );
  NOR2_X1 U25201 ( .A1(n15034), .A2(n7705), .ZN(n36221) );
  INV_X1 U5713 ( .I(n35396), .ZN(n36305) );
  NAND2_X1 U36474 ( .A1(n18496), .A2(n17243), .ZN(n37131) );
  NAND2_X1 U35046 ( .A1(n7933), .A2(n1217), .ZN(n36460) );
  NAND2_X1 U2328 ( .A1(n37181), .A2(n37335), .ZN(n37003) );
  OAI21_X1 U35794 ( .A1(n2589), .A2(n20779), .B(n37363), .ZN(n37367) );
  NAND2_X1 U13382 ( .A1(n24358), .A2(n36926), .ZN(n11835) );
  NOR2_X1 U2234 ( .A1(n18583), .A2(n37212), .ZN(n37221) );
  OAI21_X1 U8792 ( .A1(n36494), .A2(n36483), .B(n21058), .ZN(n35555) );
  NAND2_X1 U13274 ( .A1(n36664), .A2(n36672), .ZN(n36667) );
  NOR3_X1 U46504 ( .A1(n1773), .A2(n21010), .A3(n35909), .ZN(n31533) );
  NOR3_X1 U31313 ( .A1(n22527), .A2(n10829), .A3(n36494), .ZN(n36498) );
  NAND2_X1 U40478 ( .A1(n23626), .A2(n10254), .ZN(n35573) );
  NOR2_X1 U36467 ( .A1(n36072), .A2(n35396), .ZN(n25771) );
  NAND2_X1 U48342 ( .A1(n35985), .A2(n61180), .ZN(n34893) );
  NAND2_X1 U42911 ( .A1(n35383), .A2(n18144), .ZN(n35384) );
  NAND3_X1 U36459 ( .A1(n26052), .A2(n63430), .A3(n18496), .ZN(n37273) );
  INV_X1 U42377 ( .I(n37271), .ZN(n38552) );
  NOR2_X1 U27346 ( .A1(n36786), .A2(n22733), .ZN(n37129) );
  NOR2_X1 U41112 ( .A1(n576), .A2(n21329), .ZN(n32857) );
  NAND2_X1 U17921 ( .A1(n35896), .A2(n31786), .ZN(n31782) );
  INV_X1 U18001 ( .I(n15488), .ZN(n35368) );
  NAND2_X1 U35023 ( .A1(n34484), .A2(n36940), .ZN(n34486) );
  OAI21_X1 U48756 ( .A1(n36311), .A2(n36310), .B(n36309), .ZN(n36315) );
  NOR2_X1 U2225 ( .A1(n36663), .A2(n62942), .ZN(n7966) );
  NOR2_X1 U32326 ( .A1(n36176), .A2(n12288), .ZN(n35370) );
  OAI21_X1 U48617 ( .A1(n36886), .A2(n36973), .B(n61937), .ZN(n35855) );
  INV_X1 U17991 ( .I(n35897), .ZN(n34491) );
  OAI21_X1 U17817 ( .A1(n3171), .A2(n23449), .B(n18583), .ZN(n36352) );
  NOR2_X1 U11471 ( .A1(n11558), .A2(n36928), .ZN(n7430) );
  NAND2_X1 U37480 ( .A1(n18208), .A2(n35351), .ZN(n18206) );
  NAND2_X1 U8770 ( .A1(n24961), .A2(n24962), .ZN(n24050) );
  NAND4_X1 U48844 ( .A1(n36626), .A2(n36625), .A3(n36624), .A4(n63643), .ZN(
        n36629) );
  NAND3_X1 U49047 ( .A1(n37167), .A2(n37166), .A3(n37165), .ZN(n37170) );
  NAND4_X1 U4415 ( .A1(n34917), .A2(n34916), .A3(n35429), .A4(n34915), .ZN(
        n34918) );
  NOR2_X1 U6380 ( .A1(n36609), .A2(n25334), .ZN(n25565) );
  OAI21_X1 U34164 ( .A1(n31783), .A2(n31784), .B(n24118), .ZN(n14722) );
  OAI21_X1 U35296 ( .A1(n36674), .A2(n35407), .B(n26209), .ZN(n24381) );
  NAND3_X1 U23068 ( .A1(n4308), .A2(n34480), .A3(n25385), .ZN(n20042) );
  CLKBUF_X2 U2159 ( .I(n14738), .Z(n14737) );
  INV_X1 U30050 ( .I(n37799), .ZN(n38219) );
  INV_X1 U17577 ( .I(n18057), .ZN(n14143) );
  BUF_X2 U41919 ( .I(n38835), .Z(n22698) );
  INV_X2 U9461 ( .I(n1762), .ZN(n1337) );
  INV_X1 U33816 ( .I(n14259), .ZN(n38892) );
  INV_X1 U25058 ( .I(n18115), .ZN(n5363) );
  INV_X1 U2124 ( .I(n25721), .ZN(n18832) );
  INV_X2 U2058 ( .I(n19611), .ZN(n40104) );
  INV_X2 U17492 ( .I(n38023), .ZN(n1747) );
  INV_X2 U11353 ( .I(n39507), .ZN(n1407) );
  INV_X2 U2040 ( .I(n1410), .ZN(n12285) );
  INV_X1 U2056 ( .I(n39817), .ZN(n41382) );
  INV_X2 U8408 ( .I(n24991), .ZN(n1744) );
  NOR2_X1 U32387 ( .A1(n40056), .A2(n40047), .ZN(n12353) );
  INV_X1 U2075 ( .I(n1408), .ZN(n25921) );
  NOR2_X1 U5129 ( .A1(n12082), .A2(n25118), .ZN(n37926) );
  NAND2_X1 U2016 ( .A1(n12609), .A2(n14165), .ZN(n40737) );
  BUF_X2 U11346 ( .I(n14317), .Z(n24066) );
  BUF_X2 U11355 ( .I(n38923), .Z(n38932) );
  INV_X1 U7136 ( .I(n18623), .ZN(n18661) );
  INV_X2 U41954 ( .I(n25258), .ZN(n42479) );
  INV_X2 U1919 ( .I(n41210), .ZN(n38935) );
  INV_X1 U1904 ( .I(n22525), .ZN(n40766) );
  INV_X1 U28575 ( .I(n39094), .ZN(n13307) );
  INV_X2 U8761 ( .I(n26110), .ZN(n1274) );
  INV_X2 U1916 ( .I(n39959), .ZN(n16980) );
  NAND2_X1 U13095 ( .A1(n12384), .A2(n21171), .ZN(n21717) );
  INV_X2 U9433 ( .I(n40666), .ZN(n41183) );
  INV_X1 U2030 ( .I(n17212), .ZN(n1731) );
  NOR2_X1 U10141 ( .A1(n7257), .A2(n38035), .ZN(n40991) );
  INV_X1 U10173 ( .I(n41949), .ZN(n20227) );
  INV_X1 U1906 ( .I(n40857), .ZN(n40852) );
  NAND2_X1 U7710 ( .A1(n41854), .A2(n42503), .ZN(n13725) );
  NAND2_X1 U13146 ( .A1(n64793), .A2(n38675), .ZN(n40727) );
  CLKBUF_X2 U40635 ( .I(n42489), .Z(n20751) );
  NOR2_X1 U2003 ( .A1(n1306), .A2(n41161), .ZN(n40641) );
  INV_X2 U33339 ( .I(n25247), .ZN(n41257) );
  NAND2_X1 U1899 ( .A1(n41122), .A2(n473), .ZN(n40000) );
  INV_X2 U11286 ( .I(n41059), .ZN(n6855) );
  BUF_X2 U6767 ( .I(n1733), .Z(n664) );
  NAND3_X1 U30882 ( .A1(n40047), .A2(n19611), .A3(n12285), .ZN(n40099) );
  NAND2_X1 U7114 ( .A1(n1307), .A2(n42432), .ZN(n40312) );
  INV_X1 U9440 ( .I(n1741), .ZN(n41255) );
  AOI21_X1 U3564 ( .A1(n64793), .A2(n3246), .B(n11959), .ZN(n6891) );
  NAND2_X1 U32474 ( .A1(n12466), .A2(n9980), .ZN(n42491) );
  NOR2_X1 U9416 ( .A1(n61308), .A2(n40603), .ZN(n17769) );
  INV_X1 U1958 ( .I(n41951), .ZN(n41943) );
  NOR2_X1 U27671 ( .A1(n21295), .A2(n60928), .ZN(n41009) );
  NAND2_X1 U1922 ( .A1(n42299), .A2(n41270), .ZN(n42292) );
  CLKBUF_X2 U17440 ( .I(n15378), .Z(n22746) );
  NAND2_X1 U1858 ( .A1(n40100), .A2(n19990), .ZN(n40337) );
  INV_X2 U1912 ( .I(n1743), .ZN(n12895) );
  INV_X2 U1991 ( .I(n20925), .ZN(n40541) );
  INV_X1 U26270 ( .I(n10542), .ZN(n22459) );
  INV_X1 U8746 ( .I(n40605), .ZN(n1511) );
  INV_X2 U10152 ( .I(n40491), .ZN(n40659) );
  INV_X1 U9429 ( .I(n41469), .ZN(n14512) );
  NAND2_X1 U9410 ( .A1(n12466), .A2(n13984), .ZN(n42494) );
  NOR2_X1 U35054 ( .A1(n40602), .A2(n1512), .ZN(n41022) );
  NAND2_X1 U1844 ( .A1(n14462), .A2(n40644), .ZN(n41167) );
  INV_X1 U7168 ( .I(n40441), .ZN(n41101) );
  INV_X1 U31497 ( .I(n4968), .ZN(n40930) );
  INV_X1 U42734 ( .I(n40224), .ZN(n40133) );
  NAND2_X1 U22871 ( .A1(n13984), .A2(n4171), .ZN(n40129) );
  NAND2_X1 U11326 ( .A1(n41906), .A2(n42263), .ZN(n10668) );
  NAND2_X1 U7163 ( .A1(n60971), .A2(n40091), .ZN(n40086) );
  NAND2_X1 U1834 ( .A1(n39072), .A2(n40542), .ZN(n40540) );
  NAND3_X1 U13112 ( .A1(n11787), .A2(n40490), .A3(n40659), .ZN(n39036) );
  AOI22_X1 U50733 ( .A1(n40363), .A2(n40359), .B1(n41312), .B2(n10593), .ZN(
        n40364) );
  NOR2_X1 U50597 ( .A1(n61710), .A2(n40568), .ZN(n39958) );
  NOR2_X1 U10120 ( .A1(n1401), .A2(n753), .ZN(n6262) );
  NAND2_X1 U6924 ( .A1(n37774), .A2(n5319), .ZN(n40583) );
  OAI21_X1 U33647 ( .A1(n14004), .A2(n37935), .B(n37934), .ZN(n37936) );
  NOR2_X1 U28199 ( .A1(n22713), .A2(n8303), .ZN(n8116) );
  NAND2_X1 U50156 ( .A1(n23492), .A2(n38675), .ZN(n39030) );
  NOR2_X1 U49923 ( .A1(n38675), .A2(n40726), .ZN(n41200) );
  NAND2_X1 U9404 ( .A1(n17769), .A2(n40607), .ZN(n40606) );
  NAND2_X1 U3793 ( .A1(n40051), .A2(n16852), .ZN(n40275) );
  NAND2_X1 U28159 ( .A1(n1510), .A2(n42448), .ZN(n42455) );
  NOR2_X1 U1864 ( .A1(n17964), .A2(n22913), .ZN(n40516) );
  NAND2_X1 U13115 ( .A1(n13985), .A2(n40094), .ZN(n40125) );
  INV_X1 U9432 ( .I(n41885), .ZN(n39795) );
  NAND2_X1 U41462 ( .A1(n1741), .A2(n1744), .ZN(n22079) );
  NAND2_X1 U21856 ( .A1(n3306), .A2(n6276), .ZN(n40468) );
  AND2_X1 U8290 ( .A1(n40315), .A2(n24389), .Z(n16118) );
  AOI22_X1 U50971 ( .A1(n41102), .A2(n41101), .B1(n41100), .B2(n25358), .ZN(
        n41117) );
  OAI21_X1 U6055 ( .A1(n40515), .A2(n40516), .B(n41030), .ZN(n40520) );
  OAI21_X1 U29450 ( .A1(n41002), .A2(n22738), .B(n40611), .ZN(n16464) );
  NAND3_X1 U26246 ( .A1(n6598), .A2(n40054), .A3(n19611), .ZN(n19105) );
  AOI22_X1 U9392 ( .A1(n24742), .A2(n17450), .B1(n41021), .B2(n41022), .ZN(
        n19173) );
  NOR3_X1 U50948 ( .A1(n61005), .A2(n40997), .A3(n7257), .ZN(n40989) );
  OAI21_X1 U17195 ( .A1(n6801), .A2(n6800), .B(n60693), .ZN(n6799) );
  NAND3_X1 U51022 ( .A1(n42200), .A2(n42528), .A3(n42209), .ZN(n41296) );
  NAND3_X1 U1799 ( .A1(n66), .A2(n61850), .A3(n40406), .ZN(n6875) );
  NAND2_X1 U13071 ( .A1(n40363), .A2(n6200), .ZN(n5815) );
  NAND2_X1 U20446 ( .A1(n2247), .A2(n42263), .ZN(n24400) );
  OAI21_X1 U50160 ( .A1(n40656), .A2(n9915), .B(n5774), .ZN(n39042) );
  INV_X1 U50657 ( .I(n40190), .ZN(n40112) );
  AND2_X1 U13034 ( .A1(n41868), .A2(n41293), .Z(n15776) );
  NOR2_X1 U50717 ( .A1(n42427), .A2(n22285), .ZN(n40311) );
  NAND2_X1 U11285 ( .A1(n8853), .A2(n40954), .ZN(n10373) );
  AOI21_X1 U13015 ( .A1(n12805), .A2(n41420), .B(n20652), .ZN(n13124) );
  NAND2_X1 U23014 ( .A1(n18338), .A2(n4259), .ZN(n18328) );
  NAND2_X1 U13005 ( .A1(n14288), .A2(n41239), .ZN(n8914) );
  AOI21_X1 U34149 ( .A1(n41171), .A2(n11787), .B(n14704), .ZN(n40486) );
  NAND3_X1 U1779 ( .A1(n18016), .A2(n40105), .A3(n25923), .ZN(n25922) );
  NAND2_X1 U13000 ( .A1(n41241), .A2(n58046), .ZN(n5062) );
  AOI22_X1 U50162 ( .A1(n39043), .A2(n39042), .B1(n59554), .B2(n39041), .ZN(
        n39044) );
  NAND3_X1 U8701 ( .A1(n39330), .A2(n39329), .A3(n39328), .ZN(n39331) );
  OAI21_X1 U17021 ( .A1(n22259), .A2(n22260), .B(n42427), .ZN(n15513) );
  OAI22_X1 U49695 ( .A1(n42294), .A2(n41851), .B1(n57207), .B2(n39933), .ZN(
        n38269) );
  AOI22_X1 U11217 ( .A1(n16055), .A2(n42290), .B1(n22713), .B2(n42283), .ZN(
        n16802) );
  INV_X1 U35445 ( .I(n61442), .ZN(n20619) );
  INV_X2 U39059 ( .I(n18742), .ZN(n22606) );
  NOR2_X1 U1730 ( .A1(n42407), .A2(n19517), .ZN(n42394) );
  INV_X2 U1681 ( .I(n1704), .ZN(n43582) );
  INV_X1 U37733 ( .I(n40448), .ZN(n42634) );
  NOR2_X1 U1716 ( .A1(n43517), .A2(n19000), .ZN(n46326) );
  BUF_X4 U1684 ( .I(n42347), .Z(n295) );
  NOR2_X1 U27388 ( .A1(n23364), .A2(n39082), .ZN(n18847) );
  CLKBUF_X2 U9373 ( .I(n40448), .Z(n43381) );
  INV_X2 U33840 ( .I(n20602), .ZN(n14305) );
  BUF_X2 U40531 ( .I(n42619), .Z(n20650) );
  NAND2_X1 U34885 ( .A1(n41043), .A2(n41046), .ZN(n41773) );
  INV_X2 U23831 ( .I(n20844), .ZN(n43286) );
  NAND2_X1 U50163 ( .A1(n42180), .A2(n42784), .ZN(n42776) );
  NOR2_X1 U8680 ( .A1(n43181), .A2(n61744), .ZN(n43182) );
  OAI21_X1 U16747 ( .A1(n43527), .A2(n14364), .B(n16864), .ZN(n14363) );
  NOR4_X1 U36882 ( .A1(n4789), .A2(n43154), .A3(n20602), .A4(n64251), .ZN(
        n43159) );
  INV_X1 U36043 ( .I(n43735), .ZN(n21850) );
  NAND2_X1 U10063 ( .A1(n1501), .A2(n20922), .ZN(n41721) );
  NAND3_X1 U1540 ( .A1(n10990), .A2(n43839), .A3(n23730), .ZN(n43206) );
  NAND2_X1 U23577 ( .A1(n1717), .A2(n25210), .ZN(n40777) );
  NAND2_X1 U39628 ( .A1(n62535), .A2(n5971), .ZN(n43418) );
  CLKBUF_X2 U8666 ( .I(n43929), .Z(n4467) );
  NOR2_X1 U1623 ( .A1(n42140), .A2(n42127), .ZN(n42143) );
  INV_X2 U1664 ( .I(n22657), .ZN(n43100) );
  INV_X2 U36932 ( .I(n43154), .ZN(n43169) );
  INV_X2 U1658 ( .I(n42016), .ZN(n43043) );
  INV_X1 U43426 ( .I(n43357), .ZN(n41550) );
  NOR2_X1 U7130 ( .A1(n4322), .A2(n11039), .ZN(n6900) );
  INV_X2 U11196 ( .I(n16880), .ZN(n1706) );
  INV_X1 U32571 ( .I(n40096), .ZN(n13751) );
  INV_X1 U9305 ( .I(n42341), .ZN(n42340) );
  INV_X2 U1583 ( .I(n42672), .ZN(n1713) );
  INV_X1 U6703 ( .I(n41719), .ZN(n1699) );
  NAND2_X1 U36984 ( .A1(n1687), .A2(n24191), .ZN(n20848) );
  NAND3_X1 U16563 ( .A1(n42901), .A2(n43169), .A3(n43155), .ZN(n42902) );
  NOR2_X1 U35474 ( .A1(n43376), .A2(n43383), .ZN(n22186) );
  NOR2_X1 U1640 ( .A1(n62600), .A2(n59746), .ZN(n11019) );
  NOR2_X1 U4189 ( .A1(n42807), .A2(n61739), .ZN(n42978) );
  NOR2_X1 U8688 ( .A1(n63036), .A2(n62389), .ZN(n42316) );
  NAND2_X1 U11102 ( .A1(n21850), .A2(n8986), .ZN(n42847) );
  NAND2_X1 U51140 ( .A1(n2994), .A2(n43572), .ZN(n43579) );
  NAND2_X1 U1588 ( .A1(n15539), .A2(n43947), .ZN(n43948) );
  OR2_X1 U5725 ( .A1(n16473), .A2(n43165), .Z(n24895) );
  OAI21_X1 U50768 ( .A1(n43377), .A2(n41567), .B(n42753), .ZN(n40451) );
  NOR2_X1 U24235 ( .A1(n41757), .A2(n41755), .ZN(n43456) );
  NAND2_X1 U51094 ( .A1(n42704), .A2(n4805), .ZN(n41525) );
  NOR2_X1 U1528 ( .A1(n13478), .A2(n12312), .ZN(n43471) );
  AOI21_X1 U27673 ( .A1(n43713), .A2(n43714), .B(n1706), .ZN(n43716) );
  NOR2_X1 U28016 ( .A1(n43352), .A2(n7950), .ZN(n43353) );
  NAND4_X1 U51091 ( .A1(n41519), .A2(n42865), .A3(n295), .A4(n41518), .ZN(
        n41520) );
  NAND2_X1 U32391 ( .A1(n42355), .A2(n41980), .ZN(n12355) );
  NAND2_X1 U9342 ( .A1(n22606), .A2(n3302), .ZN(n42614) );
  NAND2_X1 U1496 ( .A1(n43339), .A2(n1708), .ZN(n8874) );
  INV_X1 U7171 ( .I(n42177), .ZN(n42174) );
  NOR2_X1 U27412 ( .A1(n15090), .A2(n42845), .ZN(n7435) );
  INV_X1 U11177 ( .I(n43039), .ZN(n42929) );
  INV_X1 U6308 ( .I(n41713), .ZN(n42919) );
  NAND2_X1 U21247 ( .A1(n42676), .A2(n2879), .ZN(n42146) );
  NAND2_X1 U4317 ( .A1(n42871), .A2(n6764), .ZN(n19319) );
  NAND2_X1 U1622 ( .A1(n8247), .A2(n43438), .ZN(n43430) );
  NAND2_X1 U1538 ( .A1(n1495), .A2(n43995), .ZN(n43986) );
  NAND2_X1 U16548 ( .A1(n20632), .A2(n16134), .ZN(n41246) );
  INV_X1 U39369 ( .I(n18919), .ZN(n43491) );
  INV_X1 U7761 ( .I(n43709), .ZN(n44229) );
  INV_X1 U1476 ( .I(n24071), .ZN(n44230) );
  NAND3_X1 U7185 ( .A1(n8185), .A2(n42155), .A3(n1708), .ZN(n43342) );
  OAI21_X1 U51113 ( .A1(n8305), .A2(n59292), .B(n59476), .ZN(n41597) );
  OAI21_X1 U28015 ( .A1(n1709), .A2(n7950), .B(n7451), .ZN(n38355) );
  NOR3_X1 U38739 ( .A1(n21935), .A2(n43290), .A3(n24179), .ZN(n21934) );
  NOR3_X1 U6154 ( .A1(n19319), .A2(n42345), .A3(n472), .ZN(n3853) );
  NAND3_X1 U40239 ( .A1(n19882), .A2(n43043), .A3(n42926), .ZN(n42549) );
  NAND2_X1 U51176 ( .A1(n60866), .A2(n57528), .ZN(n41747) );
  NOR2_X1 U1494 ( .A1(n43306), .A2(n22881), .ZN(n12064) );
  NAND3_X1 U16837 ( .A1(n43163), .A2(n15214), .A3(n42896), .ZN(n42059) );
  NOR2_X1 U25878 ( .A1(n43912), .A2(n6225), .ZN(n43926) );
  NAND2_X1 U51669 ( .A1(n22087), .A2(n22553), .ZN(n43629) );
  OAI21_X1 U51414 ( .A1(n20784), .A2(n6705), .B(n1497), .ZN(n42685) );
  OAI21_X1 U51037 ( .A1(n20244), .A2(n5939), .B(n9672), .ZN(n42381) );
  NOR4_X1 U7208 ( .A1(n41605), .A2(n5026), .A3(n41606), .A4(n42103), .ZN(n5313) );
  AOI21_X1 U28925 ( .A1(n42586), .A2(n42585), .B(n8873), .ZN(n8872) );
  NOR3_X1 U29810 ( .A1(n9749), .A2(n43109), .A3(n9748), .ZN(n12272) );
  NAND3_X1 U20013 ( .A1(n42646), .A2(n43489), .A3(n13730), .ZN(n1935) );
  BUF_X4 U1389 ( .I(n46291), .Z(n23722) );
  BUF_X2 U16398 ( .I(n26246), .Z(n4990) );
  INV_X1 U5982 ( .I(n46538), .ZN(n419) );
  BUF_X2 U1395 ( .I(n44242), .Z(n23828) );
  INV_X1 U1384 ( .I(n11113), .ZN(n44501) );
  INV_X1 U37515 ( .I(n21516), .ZN(n46582) );
  INV_X1 U1386 ( .I(n7302), .ZN(n44389) );
  INV_X1 U36894 ( .I(n22883), .ZN(n44319) );
  INV_X1 U5893 ( .I(n7410), .ZN(n1683) );
  INV_X1 U4246 ( .I(n46269), .ZN(n9079) );
  INV_X1 U12713 ( .I(n44965), .ZN(n1670) );
  INV_X1 U29881 ( .I(n26212), .ZN(n46386) );
  INV_X1 U7229 ( .I(n22994), .ZN(n1679) );
  INV_X2 U8226 ( .I(n45992), .ZN(n45988) );
  NOR2_X1 U34688 ( .A1(n47605), .A2(n45967), .ZN(n47611) );
  INV_X2 U9283 ( .I(n25841), .ZN(n45203) );
  INV_X2 U1300 ( .I(n863), .ZN(n12850) );
  INV_X4 U4475 ( .I(n15728), .ZN(n2955) );
  BUF_X2 U12693 ( .I(n24579), .Z(n1666) );
  INV_X1 U12692 ( .I(n24579), .ZN(n45724) );
  INV_X1 U1221 ( .I(n58232), .ZN(n45493) );
  INV_X2 U11008 ( .I(n44770), .ZN(n48248) );
  INV_X1 U16151 ( .I(n9907), .ZN(n11810) );
  INV_X1 U37040 ( .I(n47328), .ZN(n47317) );
  BUF_X2 U8630 ( .I(n2024), .Z(n23606) );
  BUF_X4 U4715 ( .I(n17128), .Z(n24114) );
  INV_X2 U43579 ( .I(n47304), .ZN(n47296) );
  NOR2_X1 U1254 ( .A1(n22508), .A2(n25896), .ZN(n47706) );
  INV_X1 U25647 ( .I(n9758), .ZN(n24340) );
  INV_X2 U1309 ( .I(n48533), .ZN(n21178) );
  NAND2_X1 U8621 ( .A1(n22574), .A2(n20897), .ZN(n47204) );
  NAND2_X1 U53044 ( .A1(n48082), .A2(n48076), .ZN(n48566) );
  INV_X2 U27159 ( .I(n59418), .ZN(n47251) );
  INV_X2 U23084 ( .I(n16020), .ZN(n47250) );
  NOR2_X1 U25700 ( .A1(n13258), .A2(n6034), .ZN(n45494) );
  NOR2_X1 U8620 ( .A1(n48248), .A2(n1082), .ZN(n48651) );
  INV_X1 U38151 ( .I(n48654), .ZN(n47488) );
  NAND2_X1 U16185 ( .A1(n3510), .A2(n61025), .ZN(n45962) );
  NAND3_X1 U31876 ( .A1(n637), .A2(n7395), .A3(n11627), .ZN(n47396) );
  NOR3_X1 U53203 ( .A1(n48511), .A2(n48521), .A3(n48514), .ZN(n47218) );
  NAND2_X1 U37099 ( .A1(n19361), .A2(n46716), .ZN(n47185) );
  INV_X2 U29161 ( .I(n44781), .ZN(n23990) );
  NAND2_X1 U1119 ( .A1(n21894), .A2(n19361), .ZN(n48113) );
  INV_X2 U1146 ( .I(n65224), .ZN(n46978) );
  NOR2_X1 U1118 ( .A1(n47180), .A2(n48622), .ZN(n48224) );
  CLKBUF_X2 U1150 ( .I(n48625), .Z(n22635) );
  NOR2_X1 U37047 ( .A1(n21976), .A2(n60753), .ZN(n46890) );
  NAND2_X1 U25812 ( .A1(n14289), .A2(n64548), .ZN(n47879) );
  INV_X1 U16110 ( .I(n61720), .ZN(n47428) );
  NOR2_X1 U9970 ( .A1(n48612), .A2(n47181), .ZN(n14418) );
  NAND2_X1 U8225 ( .A1(n7541), .A2(n59059), .ZN(n45984) );
  NAND2_X1 U9264 ( .A1(n48199), .A2(n48667), .ZN(n16538) );
  INV_X1 U16174 ( .I(n10626), .ZN(n14520) );
  INV_X1 U1137 ( .I(n45437), .ZN(n47368) );
  NAND2_X1 U35138 ( .A1(n48213), .A2(n16538), .ZN(n48197) );
  NOR3_X1 U1252 ( .A1(n47361), .A2(n47360), .A3(n64548), .ZN(n45185) );
  NAND2_X1 U16091 ( .A1(n1479), .A2(n60398), .ZN(n9101) );
  NAND2_X1 U53229 ( .A1(n47324), .A2(n60504), .ZN(n47326) );
  NOR2_X1 U52928 ( .A1(n48587), .A2(n48482), .ZN(n46474) );
  NAND2_X1 U35499 ( .A1(n60848), .A2(n48572), .ZN(n48087) );
  INV_X1 U1066 ( .I(n6034), .ZN(n45505) );
  NOR2_X1 U8622 ( .A1(n4090), .A2(n47144), .ZN(n47379) );
  NAND2_X1 U52146 ( .A1(n1294), .A2(n64063), .ZN(n44700) );
  INV_X1 U15972 ( .I(n44704), .ZN(n20725) );
  NAND2_X1 U20200 ( .A1(n47473), .A2(n47468), .ZN(n47476) );
  INV_X1 U5836 ( .I(n23263), .ZN(n48640) );
  NOR2_X1 U3773 ( .A1(n13722), .A2(n2743), .ZN(n11698) );
  INV_X1 U16224 ( .I(n45900), .ZN(n47398) );
  NAND2_X1 U52139 ( .A1(n46985), .A2(n58174), .ZN(n46988) );
  NAND2_X1 U7257 ( .A1(n46469), .A2(n2403), .ZN(n46481) );
  NAND3_X1 U22557 ( .A1(n65224), .A2(n44680), .A3(n45521), .ZN(n45741) );
  INV_X1 U8076 ( .I(n59695), .ZN(n22537) );
  NAND2_X1 U1070 ( .A1(n57731), .A2(n23990), .ZN(n45512) );
  NOR2_X1 U34950 ( .A1(n46949), .A2(n2026), .ZN(n17147) );
  NAND2_X1 U51896 ( .A1(n44194), .A2(n23480), .ZN(n44195) );
  NAND2_X1 U35512 ( .A1(n46050), .A2(n22389), .ZN(n45692) );
  NAND4_X1 U38545 ( .A1(n21953), .A2(n60946), .A3(n17573), .A4(n59616), .ZN(
        n48241) );
  NAND2_X1 U40348 ( .A1(n20340), .A2(n48544), .ZN(n21719) );
  INV_X1 U53586 ( .I(n48513), .ZN(n48516) );
  NOR2_X1 U53117 ( .A1(n46958), .A2(n13258), .ZN(n46961) );
  NOR2_X1 U12612 ( .A1(n45527), .A2(n25066), .ZN(n44703) );
  NAND2_X1 U39260 ( .A1(n18688), .A2(n16230), .ZN(n47685) );
  AOI22_X1 U34949 ( .A1(n17147), .A2(n62247), .B1(n46951), .B2(n46950), .ZN(
        n46952) );
  NAND4_X1 U22797 ( .A1(n43830), .A2(n47406), .A3(n43829), .A4(n7395), .ZN(
        n4092) );
  NAND2_X1 U10921 ( .A1(n57463), .A2(n48105), .ZN(n14623) );
  NAND2_X1 U53163 ( .A1(n48123), .A2(n48464), .ZN(n47093) );
  INV_X2 U958 ( .I(n48682), .ZN(n1644) );
  OAI22_X1 U3628 ( .A1(n10132), .A2(n48147), .B1(n21399), .B2(n21398), .ZN(
        n48159) );
  BUF_X4 U4887 ( .I(n9532), .Z(n687) );
  INV_X2 U24615 ( .I(n21269), .ZN(n49075) );
  INV_X2 U894 ( .I(n50422), .ZN(n48757) );
  BUF_X4 U23702 ( .I(n50123), .Z(n18607) );
  CLKBUF_X2 U41792 ( .I(n49466), .Z(n22526) );
  INV_X2 U967 ( .I(n49263), .ZN(n9395) );
  BUF_X2 U15735 ( .I(n25857), .Z(n24821) );
  INV_X2 U910 ( .I(n9229), .ZN(n18585) );
  NAND2_X1 U53417 ( .A1(n19681), .A2(n8044), .ZN(n47967) );
  NOR2_X1 U43914 ( .A1(n15708), .A2(n25857), .ZN(n49508) );
  INV_X1 U53263 ( .I(n49835), .ZN(n49069) );
  NAND2_X1 U920 ( .A1(n15021), .A2(n1641), .ZN(n14809) );
  NOR2_X1 U923 ( .A1(n9395), .A2(n11314), .ZN(n49412) );
  INV_X2 U893 ( .I(n57194), .ZN(n48366) );
  INV_X1 U870 ( .I(n23738), .ZN(n1472) );
  NOR2_X1 U27919 ( .A1(n14931), .A2(n1262), .ZN(n49345) );
  INV_X2 U809 ( .I(n18364), .ZN(n18469) );
  INV_X1 U26058 ( .I(n6410), .ZN(n48803) );
  INV_X1 U24653 ( .I(n22098), .ZN(n25018) );
  NAND2_X1 U38365 ( .A1(n6977), .A2(n60975), .ZN(n50005) );
  OAI21_X1 U15565 ( .A1(n45236), .A2(n49158), .B(n49459), .ZN(n3241) );
  NAND2_X1 U4505 ( .A1(n16107), .A2(n50216), .ZN(n49339) );
  NOR2_X1 U859 ( .A1(n49265), .A2(n20004), .ZN(n49407) );
  AOI21_X1 U20609 ( .A1(n23912), .A2(n9164), .B(n9455), .ZN(n2380) );
  NAND2_X1 U15654 ( .A1(n60397), .A2(n50312), .ZN(n49147) );
  NOR2_X1 U41615 ( .A1(n48006), .A2(n49090), .ZN(n49095) );
  NOR2_X1 U7265 ( .A1(n60209), .A2(n18585), .ZN(n16335) );
  NAND2_X1 U12486 ( .A1(n49323), .A2(n1292), .ZN(n49398) );
  INV_X1 U35551 ( .I(n65005), .ZN(n18683) );
  INV_X1 U9201 ( .I(n48391), .ZN(n48853) );
  NAND2_X1 U845 ( .A1(n9853), .A2(n49006), .ZN(n48324) );
  NAND2_X1 U898 ( .A1(n20428), .A2(n13440), .ZN(n18565) );
  NAND2_X1 U25968 ( .A1(n10030), .A2(n6314), .ZN(n49741) );
  NOR2_X1 U846 ( .A1(n49610), .A2(n49308), .ZN(n49612) );
  NAND2_X1 U788 ( .A1(n23738), .A2(n6654), .ZN(n49017) );
  INV_X1 U7300 ( .I(n50397), .ZN(n50079) );
  NOR2_X1 U35572 ( .A1(n50044), .A2(n19773), .ZN(n20427) );
  NOR2_X1 U53477 ( .A1(n1291), .A2(n4594), .ZN(n49979) );
  NAND3_X1 U52357 ( .A1(n9863), .A2(n15737), .A3(n2357), .ZN(n45163) );
  OAI21_X1 U22063 ( .A1(n48907), .A2(n49379), .B(n3497), .ZN(n10228) );
  NAND2_X1 U15577 ( .A1(n4017), .A2(n22869), .ZN(n4015) );
  AOI21_X1 U37118 ( .A1(n17422), .A2(n49842), .B(n49846), .ZN(n48378) );
  NAND2_X1 U10819 ( .A1(n57267), .A2(n48845), .ZN(n49197) );
  OAI21_X1 U37215 ( .A1(n48036), .A2(n48035), .B(n23738), .ZN(n48044) );
  NOR2_X1 U32238 ( .A1(n16986), .A2(n64764), .ZN(n12108) );
  INV_X1 U814 ( .I(n49383), .ZN(n49394) );
  NOR3_X1 U23267 ( .A1(n49075), .A2(n49063), .A3(n63954), .ZN(n49829) );
  NAND2_X1 U53529 ( .A1(n49910), .A2(n58037), .ZN(n48339) );
  NAND2_X1 U15475 ( .A1(n21373), .A2(n21371), .ZN(n23242) );
  NAND2_X1 U673 ( .A1(n21183), .A2(n50394), .ZN(n50408) );
  NAND2_X1 U23275 ( .A1(n8729), .A2(n17885), .ZN(n47761) );
  NOR2_X1 U28929 ( .A1(n19144), .A2(n7866), .ZN(n8878) );
  NAND3_X1 U53330 ( .A1(n49677), .A2(n20971), .A3(n49671), .ZN(n47648) );
  AOI21_X1 U665 ( .A1(n25459), .A2(n48453), .B(n49017), .ZN(n5812) );
  NAND2_X1 U10796 ( .A1(n49775), .A2(n48949), .ZN(n4299) );
  NOR3_X1 U9880 ( .A1(n14642), .A2(n49258), .A3(n25680), .ZN(n19831) );
  OAI21_X1 U53406 ( .A1(n49112), .A2(n47942), .B(n48441), .ZN(n47952) );
  NAND2_X1 U4269 ( .A1(n48450), .A2(n49011), .ZN(n23421) );
  AOI21_X1 U9182 ( .A1(n49020), .A2(n5219), .B(n63389), .ZN(n49021) );
  OAI21_X1 U34043 ( .A1(n48346), .A2(n48798), .B(n14561), .ZN(n48348) );
  NOR3_X1 U33422 ( .A1(n13632), .A2(n49553), .A3(n13631), .ZN(n48023) );
  OAI21_X1 U8552 ( .A1(n49699), .A2(n49698), .B(n49697), .ZN(n49706) );
  INV_X1 U12351 ( .I(n6583), .ZN(n48796) );
  NAND2_X1 U691 ( .A1(n7779), .A2(n11314), .ZN(n5208) );
  NOR2_X1 U15575 ( .A1(n49743), .A2(n49458), .ZN(n13363) );
  NAND2_X1 U743 ( .A1(n23650), .A2(n61355), .ZN(n9409) );
  AOI21_X1 U15516 ( .A1(n48738), .A2(n48737), .B(n48736), .ZN(n12292) );
  NOR2_X1 U31746 ( .A1(n50120), .A2(n50121), .ZN(n11449) );
  INV_X1 U15525 ( .I(n49359), .ZN(n8502) );
  BUF_X2 U43329 ( .I(n51601), .Z(n25061) );
  INV_X2 U41291 ( .I(n1622), .ZN(n21700) );
  BUF_X2 U15146 ( .I(n52331), .Z(n23375) );
  BUF_X2 U34270 ( .I(n25192), .Z(n14870) );
  BUF_X2 U9168 ( .I(n12800), .Z(n12799) );
  CLKBUF_X2 U28348 ( .I(n19540), .Z(n8273) );
  INV_X1 U54014 ( .I(n23344), .ZN(n51087) );
  INV_X1 U558 ( .I(n14870), .ZN(n9847) );
  INV_X1 U584 ( .I(n1189), .ZN(n24379) );
  INV_X1 U38101 ( .I(n65280), .ZN(n51990) );
  INV_X1 U540 ( .I(n55950), .ZN(n20125) );
  INV_X1 U538 ( .I(n52686), .ZN(n52683) );
  BUF_X2 U495 ( .I(n53915), .Z(n4399) );
  INV_X1 U15033 ( .I(n54815), .ZN(n1607) );
  BUF_X2 U23764 ( .I(n55950), .Z(n4634) );
  INV_X1 U14878 ( .I(n51529), .ZN(n25359) );
  NOR2_X1 U39894 ( .A1(n13370), .A2(n19555), .ZN(n53185) );
  CLKBUF_X2 U5150 ( .I(n55400), .Z(n197) );
  INV_X1 U42623 ( .I(n2408), .ZN(n52701) );
  INV_X2 U41075 ( .I(n55909), .ZN(n55721) );
  NAND2_X1 U22232 ( .A1(n3616), .A2(n56268), .ZN(n5668) );
  NOR2_X1 U9156 ( .A1(n23763), .A2(n22807), .ZN(n55255) );
  NAND2_X1 U32759 ( .A1(n5536), .A2(n52866), .ZN(n52696) );
  INV_X2 U536 ( .I(n55671), .ZN(n55677) );
  INV_X1 U42334 ( .I(n53407), .ZN(n54041) );
  OAI21_X1 U29577 ( .A1(n25522), .A2(n53576), .B(n23476), .ZN(n53227) );
  NAND2_X1 U458 ( .A1(n53861), .A2(n53860), .ZN(n53417) );
  NAND2_X1 U55578 ( .A1(n54594), .A2(n54074), .ZN(n53890) );
  NOR2_X1 U449 ( .A1(n55433), .A2(n23275), .ZN(n55323) );
  INV_X1 U12295 ( .I(n22807), .ZN(n54980) );
  NAND2_X1 U20710 ( .A1(n22544), .A2(n54949), .ZN(n54785) );
  NAND2_X1 U54971 ( .A1(n20156), .A2(n20982), .ZN(n52870) );
  INV_X4 U406 ( .I(n54594), .ZN(n54596) );
  INV_X1 U41031 ( .I(n65281), .ZN(n56441) );
  NAND3_X1 U4407 ( .A1(n8597), .A2(n52890), .A3(n56985), .ZN(n51440) );
  NAND2_X1 U56075 ( .A1(n55271), .A2(n63194), .ZN(n55272) );
  NOR2_X1 U4135 ( .A1(n3567), .A2(n55679), .ZN(n9263) );
  INV_X2 U5372 ( .I(n61725), .ZN(n54601) );
  NAND2_X1 U364 ( .A1(n1157), .A2(n13940), .ZN(n53880) );
  INV_X1 U14969 ( .I(n54955), .ZN(n1597) );
  NAND2_X1 U31906 ( .A1(n1370), .A2(n14324), .ZN(n13022) );
  NOR2_X1 U371 ( .A1(n54814), .A2(n1371), .ZN(n54096) );
  INV_X1 U54980 ( .I(n56234), .ZN(n56365) );
  NOR2_X1 U54798 ( .A1(n52987), .A2(n60794), .ZN(n53850) );
  NOR2_X1 U55083 ( .A1(n61895), .A2(n197), .ZN(n52564) );
  OAI21_X1 U55128 ( .A1(n52863), .A2(n62434), .B(n62886), .ZN(n52661) );
  NAND3_X1 U56470 ( .A1(n56211), .A2(n56635), .A3(n21893), .ZN(n56212) );
  INV_X1 U28463 ( .I(n8375), .ZN(n20933) );
  NOR2_X1 U27418 ( .A1(n56593), .A2(n57691), .ZN(n56254) );
  INV_X1 U309 ( .I(n53577), .ZN(n52998) );
  NAND2_X1 U27859 ( .A1(n54601), .A2(n7789), .ZN(n54593) );
  AOI21_X1 U33874 ( .A1(n55288), .A2(n22588), .B(n61247), .ZN(n55289) );
  NOR2_X1 U55239 ( .A1(n61895), .A2(n55250), .ZN(n52907) );
  NAND2_X1 U35213 ( .A1(n61213), .A2(n56434), .ZN(n56230) );
  NAND3_X1 U54680 ( .A1(n56374), .A2(n56660), .A3(n52282), .ZN(n51559) );
  INV_X1 U30152 ( .I(n52120), .ZN(n9975) );
  NOR2_X1 U34577 ( .A1(n15317), .A2(n15314), .ZN(n15313) );
  OAI21_X1 U37812 ( .A1(n50899), .A2(n56230), .B(n16331), .ZN(n56127) );
  OAI21_X1 U300 ( .A1(n53000), .A2(n52999), .B(n52998), .ZN(n53013) );
  NAND2_X1 U10684 ( .A1(n52694), .A2(n23526), .ZN(n56831) );
  NOR3_X1 U274 ( .A1(n50672), .A2(n50673), .A3(n52842), .ZN(n50678) );
  NAND2_X1 U8309 ( .A1(n54863), .A2(n671), .ZN(n5216) );
  OAI21_X1 U14752 ( .A1(n19321), .A2(n19320), .B(n25160), .ZN(n52835) );
  NOR3_X1 U30239 ( .A1(n53583), .A2(n53584), .A3(n53585), .ZN(n53595) );
  OAI21_X1 U26771 ( .A1(n54989), .A2(n61895), .B(n54987), .ZN(n55012) );
  BUF_X4 U14614 ( .I(n8966), .Z(n1592) );
  INV_X1 U256 ( .I(n1232), .ZN(n12959) );
  INV_X1 U55406 ( .I(n53483), .ZN(n53514) );
  INV_X1 U14495 ( .I(n53807), .ZN(n53808) );
  NAND2_X1 U149 ( .A1(n2329), .A2(n2049), .ZN(n54913) );
  NOR2_X1 U8307 ( .A1(n53129), .A2(n4808), .ZN(n53140) );
  NAND2_X1 U185 ( .A1(n56697), .A2(n56734), .ZN(n6954) );
  NAND2_X1 U43433 ( .A1(n57122), .A2(n23538), .ZN(n57115) );
  NAND2_X1 U34610 ( .A1(n19491), .A2(n54758), .ZN(n54742) );
  INV_X2 U7961 ( .I(n54542), .ZN(n54581) );
  INV_X1 U36301 ( .I(n54272), .ZN(n54280) );
  NOR2_X1 U55433 ( .A1(n53492), .A2(n23611), .ZN(n53489) );
  INV_X1 U142 ( .I(n21922), .ZN(n53505) );
  NAND2_X1 U26964 ( .A1(n17795), .A2(n21860), .ZN(n56489) );
  NAND2_X1 U37420 ( .A1(n55166), .A2(n62699), .ZN(n55162) );
  NAND4_X1 U55399 ( .A1(n53369), .A2(n1450), .A3(n60115), .A4(n52762), .ZN(
        n53370) );
  NAND3_X1 U56306 ( .A1(n55855), .A2(n11789), .A3(n55854), .ZN(n55856) );
  NAND2_X1 U55995 ( .A1(n55102), .A2(n25170), .ZN(n55037) );
  NAND2_X1 U4082 ( .A1(n9550), .A2(n26094), .ZN(n26093) );
  NAND2_X1 U4025 ( .A1(n54769), .A2(n54767), .ZN(n24038) );
  INV_X1 U26576 ( .I(n6902), .ZN(n13775) );
  NAND2_X1 U30892 ( .A1(n1257), .A2(n14708), .ZN(n56968) );
  CLKBUF_X2 U40728 ( .I(n16943), .Z(n20839) );
  NAND2_X1 U3530 ( .A1(n19491), .A2(n54741), .ZN(n54682) );
  INV_X1 U70 ( .I(n19735), .ZN(n53302) );
  INV_X1 U34393 ( .I(n15237), .ZN(n19827) );
  AOI21_X1 U3832 ( .A1(n2820), .A2(n9187), .B(n53130), .ZN(n12209) );
  NAND3_X1 U55994 ( .A1(n55079), .A2(n55057), .A3(n1233), .ZN(n55040) );
  NOR2_X1 U55751 ( .A1(n22315), .A2(n23731), .ZN(n54274) );
  NAND2_X1 U14539 ( .A1(n53351), .A2(n53334), .ZN(n17013) );
  NAND2_X1 U41 ( .A1(n8412), .A2(n55097), .ZN(n55048) );
  NOR2_X1 U56185 ( .A1(n4801), .A2(n55569), .ZN(n55585) );
  OAI21_X1 U28496 ( .A1(n8411), .A2(n8410), .B(n55068), .ZN(n55094) );
  AOI21_X1 U42 ( .A1(n5649), .A2(n53904), .B(n5651), .ZN(n2568) );
  AND2_X1 U37486 ( .A1(n55880), .A2(n60203), .Z(n15800) );
  NAND2_X1 U14394 ( .A1(n2820), .A2(n3195), .ZN(n4644) );
  NOR3_X1 U39501 ( .A1(n56956), .A2(n56955), .A3(n56954), .ZN(n56975) );
  OAI21_X1 U5650 ( .A1(n320), .A2(n1181), .B(n53700), .ZN(n22707) );
  NOR2_X1 U14360 ( .A1(n13708), .A2(n13707), .ZN(n13706) );
  NAND4_X1 U56428 ( .A1(n56096), .A2(n56095), .A3(n56094), .A4(n56093), .ZN(
        n56098) );
  NAND2_X1 U14 ( .A1(n60240), .A2(n12395), .ZN(n12394) );
  NAND2_X1 U15 ( .A1(n59537), .A2(n9096), .ZN(n9700) );
  NAND2_X1 U16 ( .A1(n59920), .A2(n57099), .ZN(n57112) );
  AND2_X1 U23 ( .A1(n518), .A2(n53294), .Z(n16097) );
  NOR3_X1 U34 ( .A1(n1582), .A2(n56295), .A3(n60353), .ZN(n56320) );
  OAI21_X1 U45 ( .A1(n15238), .A2(n56502), .B(n21859), .ZN(n56492) );
  NAND2_X1 U49 ( .A1(n7209), .A2(n23030), .ZN(n61688) );
  NOR2_X1 U52 ( .A1(n9093), .A2(n9094), .ZN(n59537) );
  NAND2_X1 U58 ( .A1(n1578), .A2(n56967), .ZN(n21504) );
  OAI21_X1 U61 ( .A1(n13775), .A2(n56955), .B(n56940), .ZN(n60240) );
  INV_X1 U89 ( .I(n56290), .ZN(n56296) );
  NAND2_X1 U90 ( .A1(n57129), .A2(n19054), .ZN(n57160) );
  INV_X1 U119 ( .I(n55899), .ZN(n18561) );
  NOR2_X1 U128 ( .A1(n6061), .A2(n6168), .ZN(n53996) );
  NAND2_X1 U152 ( .A1(n61058), .A2(n16503), .ZN(n15293) );
  BUF_X2 U173 ( .I(n59610), .Z(n10381) );
  NAND2_X1 U197 ( .A1(n56725), .A2(n56674), .ZN(n60563) );
  INV_X2 U248 ( .I(n56965), .ZN(n56953) );
  NAND2_X1 U269 ( .A1(n57675), .A2(n57672), .ZN(n55485) );
  AOI21_X1 U280 ( .A1(n51454), .A2(n51455), .B(n58060), .ZN(n51460) );
  AOI21_X1 U281 ( .A1(n60045), .A2(n22447), .B(n17754), .ZN(n22450) );
  NAND3_X1 U286 ( .A1(n55408), .A2(n58333), .A3(n55403), .ZN(n20822) );
  NAND2_X1 U307 ( .A1(n10190), .A2(n61907), .ZN(n59791) );
  AND2_X1 U311 ( .A1(n52247), .A2(n13489), .Z(n15988) );
  AOI22_X1 U313 ( .A1(n57035), .A2(n57034), .B1(n2742), .B2(n57027), .ZN(
        n21574) );
  NOR2_X1 U314 ( .A1(n22592), .A2(n248), .ZN(n57673) );
  AND2_X1 U331 ( .A1(n13489), .A2(n16645), .Z(n56380) );
  NOR2_X1 U334 ( .A1(n55720), .A2(n1324), .ZN(n60103) );
  INV_X1 U339 ( .I(n12729), .ZN(n61476) );
  NOR2_X1 U344 ( .A1(n55905), .A2(n55908), .ZN(n60102) );
  NOR2_X1 U348 ( .A1(n53181), .A2(n62090), .ZN(n53189) );
  NAND2_X1 U370 ( .A1(n540), .A2(n58978), .ZN(n54629) );
  NAND3_X1 U374 ( .A1(n1597), .A2(n2467), .A3(n22749), .ZN(n2466) );
  NOR2_X1 U379 ( .A1(n57083), .A2(n10191), .ZN(n10190) );
  NAND2_X1 U380 ( .A1(n9765), .A2(n9296), .ZN(n53230) );
  OR2_X1 U386 ( .A1(n5569), .A2(n58283), .Z(n57235) );
  NAND2_X1 U412 ( .A1(n55270), .A2(n61081), .ZN(n57695) );
  NOR2_X1 U434 ( .A1(n61247), .A2(n55726), .ZN(n58552) );
  NAND2_X1 U438 ( .A1(n9111), .A2(n56268), .ZN(n58784) );
  NAND2_X1 U446 ( .A1(n53835), .A2(n60794), .ZN(n57744) );
  NAND2_X1 U454 ( .A1(n7148), .A2(n22760), .ZN(n54462) );
  NAND2_X1 U459 ( .A1(n55476), .A2(n55474), .ZN(n52927) );
  NOR2_X1 U460 ( .A1(n54034), .A2(n54035), .ZN(n58006) );
  NOR2_X1 U470 ( .A1(n53916), .A2(n23164), .ZN(n52974) );
  INV_X1 U476 ( .I(n3708), .ZN(n54822) );
  CLKBUF_X2 U478 ( .I(n1616), .Z(n61213) );
  BUF_X2 U494 ( .I(n21957), .Z(n61554) );
  NAND2_X1 U502 ( .A1(n24003), .A2(n55680), .ZN(n55452) );
  INV_X1 U506 ( .I(n56412), .ZN(n57191) );
  INV_X1 U519 ( .I(n55456), .ZN(n60553) );
  NAND2_X1 U544 ( .A1(n57073), .A2(n21669), .ZN(n52674) );
  INV_X1 U552 ( .I(n6351), .ZN(n17257) );
  NOR2_X1 U559 ( .A1(n54798), .A2(n10441), .ZN(n54972) );
  NOR2_X1 U560 ( .A1(n54034), .A2(n21919), .ZN(n57699) );
  INV_X1 U566 ( .I(n3376), .ZN(n7518) );
  INV_X1 U592 ( .I(n54292), .ZN(n58491) );
  BUF_X4 U622 ( .I(n52475), .Z(n58283) );
  NAND2_X1 U628 ( .A1(n26041), .A2(n53917), .ZN(n54034) );
  BUF_X2 U636 ( .I(n55248), .Z(n23763) );
  INV_X1 U643 ( .I(n1463), .ZN(n15079) );
  NAND2_X1 U676 ( .A1(n49237), .A2(n49236), .ZN(n50942) );
  OAI21_X1 U752 ( .A1(n57816), .A2(n57815), .B(n57610), .ZN(n49469) );
  NAND3_X1 U775 ( .A1(n58322), .A2(n50375), .A3(n3031), .ZN(n12581) );
  NAND2_X1 U786 ( .A1(n49475), .A2(n60209), .ZN(n59717) );
  AOI21_X1 U787 ( .A1(n60515), .A2(n47949), .B(n47948), .ZN(n47950) );
  NOR2_X1 U797 ( .A1(n49150), .A2(n57609), .ZN(n1115) );
  INV_X1 U807 ( .I(n48450), .ZN(n2075) );
  NOR2_X1 U815 ( .A1(n48691), .A2(n47921), .ZN(n17675) );
  NOR2_X1 U816 ( .A1(n49272), .A2(n9455), .ZN(n12556) );
  NOR3_X1 U820 ( .A1(n3738), .A2(n19523), .A3(n1641), .ZN(n3737) );
  NAND2_X1 U823 ( .A1(n49452), .A2(n49844), .ZN(n58271) );
  AOI21_X1 U824 ( .A1(n14561), .A2(n48811), .B(n48810), .ZN(n48812) );
  NAND2_X1 U826 ( .A1(n50374), .A2(n12580), .ZN(n58322) );
  NAND3_X1 U838 ( .A1(n23992), .A2(n60853), .A3(n60041), .ZN(n3681) );
  NAND2_X1 U864 ( .A1(n2878), .A2(n23063), .ZN(n60041) );
  NOR3_X1 U876 ( .A1(n14315), .A2(n63546), .A3(n49910), .ZN(n48735) );
  OR2_X1 U903 ( .A1(n14315), .A2(n21406), .Z(n15832) );
  NAND2_X1 U917 ( .A1(n2810), .A2(n47920), .ZN(n61525) );
  NOR2_X1 U929 ( .A1(n20004), .A2(n9395), .ZN(n12558) );
  NOR2_X1 U932 ( .A1(n59621), .A2(n17885), .ZN(n10080) );
  AOI21_X1 U933 ( .A1(n11154), .A2(n11155), .B(n49674), .ZN(n61248) );
  NOR3_X1 U936 ( .A1(n50438), .A2(n18882), .A3(n17885), .ZN(n8725) );
  NOR3_X1 U941 ( .A1(n50079), .A2(n20174), .A3(n50078), .ZN(n58198) );
  NOR3_X1 U943 ( .A1(n24821), .A2(n406), .A3(n48847), .ZN(n14779) );
  NAND3_X1 U947 ( .A1(n49301), .A2(n49300), .A3(n9594), .ZN(n58657) );
  NAND2_X1 U961 ( .A1(n7271), .A2(n23802), .ZN(n49110) );
  OR2_X1 U970 ( .A1(n58856), .A2(n5743), .Z(n57465) );
  INV_X1 U1001 ( .I(n13118), .ZN(n59884) );
  INV_X1 U1003 ( .I(n2754), .ZN(n58336) );
  NOR2_X1 U1004 ( .A1(n64631), .A2(n49538), .ZN(n10637) );
  AOI22_X1 U1029 ( .A1(n48041), .A2(n48449), .B1(n48448), .B2(n48040), .ZN(
        n59207) );
  OAI22_X1 U1031 ( .A1(n50211), .A2(n16766), .B1(n50212), .B2(n50213), .ZN(
        n5190) );
  AND2_X1 U1048 ( .A1(n44788), .A2(n48362), .Z(n57425) );
  NOR2_X1 U1053 ( .A1(n49630), .A2(n19489), .ZN(n49631) );
  NAND2_X1 U1057 ( .A1(n7824), .A2(n16765), .ZN(n50219) );
  NOR2_X1 U1074 ( .A1(n49701), .A2(n45160), .ZN(n48680) );
  INV_X1 U1120 ( .I(n5146), .ZN(n60719) );
  BUF_X2 U1130 ( .I(n49720), .Z(n61355) );
  NAND2_X1 U1174 ( .A1(n17629), .A2(n44002), .ZN(n61157) );
  NAND2_X1 U1176 ( .A1(n60850), .A2(n47023), .ZN(n10368) );
  NAND2_X1 U1242 ( .A1(n59384), .A2(n1328), .ZN(n58353) );
  OAI21_X1 U1278 ( .A1(n47800), .A2(n47699), .B(n59611), .ZN(n47805) );
  AOI21_X1 U1284 ( .A1(n58974), .A2(n48480), .B(n57238), .ZN(n1066) );
  NAND3_X1 U1307 ( .A1(n48184), .A2(n13587), .A3(n48484), .ZN(n46470) );
  OAI21_X1 U1311 ( .A1(n46814), .A2(n1477), .B(n48104), .ZN(n46815) );
  AOI21_X1 U1313 ( .A1(n21178), .A2(n20878), .B(n47190), .ZN(n7674) );
  NAND2_X1 U1319 ( .A1(n47688), .A2(n63686), .ZN(n57739) );
  INV_X1 U1329 ( .I(n47473), .ZN(n47464) );
  NAND2_X1 U1334 ( .A1(n62247), .A2(n45494), .ZN(n59651) );
  NAND3_X1 U1335 ( .A1(n44649), .A2(n46946), .A3(n23643), .ZN(n58124) );
  INV_X1 U1341 ( .I(n18138), .ZN(n47744) );
  AND2_X1 U1362 ( .A1(n21793), .A2(n65145), .Z(n57248) );
  NAND2_X1 U1363 ( .A1(n1656), .A2(n22536), .ZN(n57531) );
  NAND2_X1 U1370 ( .A1(n60557), .A2(n46890), .ZN(n58095) );
  AND2_X1 U1393 ( .A1(n20937), .A2(n23416), .Z(n48641) );
  NAND2_X1 U1408 ( .A1(n47429), .A2(n47425), .ZN(n21200) );
  NOR2_X1 U1458 ( .A1(n23542), .A2(n9851), .ZN(n8043) );
  NAND2_X1 U1466 ( .A1(n47181), .A2(n8639), .ZN(n47163) );
  CLKBUF_X2 U1467 ( .I(n11416), .Z(n57670) );
  INV_X1 U1474 ( .I(n11899), .ZN(n57635) );
  INV_X1 U1544 ( .I(n10241), .ZN(n6904) );
  INV_X1 U1559 ( .I(n9628), .ZN(n46637) );
  BUF_X2 U1645 ( .I(n22108), .Z(n21141) );
  INV_X1 U1651 ( .I(n58867), .ZN(n3504) );
  INV_X1 U1661 ( .I(n46546), .ZN(n5448) );
  OAI21_X1 U1662 ( .A1(n5059), .A2(n4386), .B(n44156), .ZN(n4047) );
  NOR2_X1 U1717 ( .A1(n8936), .A2(n42629), .ZN(n59628) );
  NOR2_X1 U1742 ( .A1(n57251), .A2(n5543), .ZN(n58017) );
  NOR2_X1 U1743 ( .A1(n58032), .A2(n61593), .ZN(n18586) );
  OAI22_X1 U1746 ( .A1(n42037), .A2(n43506), .B1(n42641), .B2(n42036), .ZN(
        n22880) );
  NOR3_X1 U1752 ( .A1(n57178), .A2(n23811), .A3(n8290), .ZN(n24999) );
  AOI21_X1 U1753 ( .A1(n291), .A2(n43416), .B(n22553), .ZN(n60474) );
  NOR2_X1 U1754 ( .A1(n1698), .A2(n42923), .ZN(n42107) );
  AND2_X1 U1758 ( .A1(n43602), .A2(n43601), .Z(n57335) );
  NOR2_X1 U1764 ( .A1(n43694), .A2(n43698), .ZN(n58274) );
  NAND3_X1 U1789 ( .A1(n59345), .A2(n59356), .A3(n1715), .ZN(n59344) );
  AND2_X1 U1792 ( .A1(n40020), .A2(n25458), .Z(n42366) );
  NAND3_X1 U1818 ( .A1(n42878), .A2(n6764), .A3(n21336), .ZN(n3855) );
  INV_X1 U1824 ( .I(n43177), .ZN(n61348) );
  NAND3_X1 U1826 ( .A1(n20848), .A2(n20847), .A3(n42989), .ZN(n60862) );
  NAND2_X1 U1828 ( .A1(n22999), .A2(n42354), .ZN(n12402) );
  NOR3_X1 U1847 ( .A1(n41657), .A2(n43579), .A3(n41656), .ZN(n41658) );
  OR2_X1 U1860 ( .A1(n25851), .A2(n65129), .Z(n57261) );
  NAND2_X1 U1869 ( .A1(n11019), .A2(n43571), .ZN(n59415) );
  NOR2_X1 U1881 ( .A1(n42108), .A2(n42551), .ZN(n58613) );
  NOR2_X1 U1890 ( .A1(n43364), .A2(n43366), .ZN(n59345) );
  NAND4_X1 U1900 ( .A1(n42848), .A2(n21326), .A3(n42667), .A4(n64532), .ZN(
        n20705) );
  NOR2_X1 U1905 ( .A1(n43848), .A2(n24002), .ZN(n521) );
  OAI21_X1 U1907 ( .A1(n42806), .A2(n1298), .B(n61858), .ZN(n15250) );
  AND2_X1 U1934 ( .A1(n42398), .A2(n42402), .Z(n57385) );
  INV_X1 U1937 ( .I(n61894), .ZN(n59517) );
  INV_X1 U1967 ( .I(n41704), .ZN(n59288) );
  OAI21_X1 U1976 ( .A1(n58872), .A2(n11229), .B(n58871), .ZN(n41629) );
  NOR2_X1 U1979 ( .A1(n43839), .A2(n60706), .ZN(n19702) );
  INV_X2 U1986 ( .I(n23702), .ZN(n1269) );
  NAND2_X1 U1995 ( .A1(n11229), .A2(n8185), .ZN(n58871) );
  CLKBUF_X2 U2013 ( .I(n9663), .Z(n59139) );
  NAND2_X1 U2019 ( .A1(n42355), .A2(n42361), .ZN(n15283) );
  NAND2_X1 U2020 ( .A1(n18398), .A2(n41568), .ZN(n19271) );
  NAND2_X1 U2042 ( .A1(n10827), .A2(n41773), .ZN(n58171) );
  NOR2_X1 U2049 ( .A1(n13730), .A2(n43912), .ZN(n14364) );
  NAND2_X1 U2065 ( .A1(n42640), .A2(n43518), .ZN(n43198) );
  BUF_X2 U2066 ( .I(n43069), .Z(n23730) );
  AND2_X1 U2073 ( .A1(n14498), .A2(n42986), .Z(n43959) );
  BUF_X2 U2076 ( .I(n41046), .Z(n42865) );
  AOI22_X1 U2102 ( .A1(n41217), .A2(n41422), .B1(n60333), .B2(n41219), .ZN(
        n57910) );
  NOR2_X1 U2104 ( .A1(n16805), .A2(n57345), .ZN(n16804) );
  NAND3_X1 U2105 ( .A1(n38267), .A2(n38265), .A3(n38266), .ZN(n59985) );
  NAND2_X1 U2106 ( .A1(n40558), .A2(n4259), .ZN(n58584) );
  OAI21_X1 U2111 ( .A1(n41198), .A2(n41199), .B(n41200), .ZN(n17468) );
  AND2_X1 U2112 ( .A1(n7571), .A2(n4918), .Z(n57387) );
  NOR2_X1 U2137 ( .A1(n60101), .A2(n12679), .ZN(n61280) );
  NAND2_X1 U2151 ( .A1(n41215), .A2(n41214), .ZN(n60333) );
  AOI21_X1 U2152 ( .A1(n17476), .A2(n41889), .B(n13551), .ZN(n57717) );
  INV_X1 U2162 ( .I(n40211), .ZN(n59285) );
  AOI21_X1 U2171 ( .A1(n3048), .A2(n41882), .B(n39793), .ZN(n8746) );
  NAND2_X1 U2180 ( .A1(n40543), .A2(n3642), .ZN(n58981) );
  AOI21_X1 U2184 ( .A1(n21928), .A2(n40271), .B(n60223), .ZN(n21925) );
  AOI22_X1 U2190 ( .A1(n41199), .A2(n41194), .B1(n40634), .B2(n57406), .ZN(
        n39033) );
  NAND2_X1 U2194 ( .A1(n42276), .A2(n16072), .ZN(n16805) );
  OR2_X1 U2197 ( .A1(n40091), .A2(n9980), .Z(n57244) );
  NOR2_X1 U2208 ( .A1(n7511), .A2(n41060), .ZN(n60690) );
  NAND3_X1 U2217 ( .A1(n60612), .A2(n42249), .A3(n41255), .ZN(n40790) );
  AOI21_X1 U2248 ( .A1(n41861), .A2(n41862), .B(n59190), .ZN(n41863) );
  OAI21_X1 U2250 ( .A1(n58139), .A2(n57382), .B(n62157), .ZN(n40266) );
  INV_X1 U2252 ( .I(n42483), .ZN(n60101) );
  NAND2_X1 U2256 ( .A1(n41806), .A2(n22759), .ZN(n38200) );
  NAND2_X1 U2270 ( .A1(n6768), .A2(n6767), .ZN(n60218) );
  NAND2_X1 U2281 ( .A1(n21927), .A2(n40275), .ZN(n60223) );
  NAND3_X1 U2287 ( .A1(n42275), .A2(n19982), .A3(n41928), .ZN(n18358) );
  AND2_X1 U2312 ( .A1(n60075), .A2(n42288), .Z(n1001) );
  NAND2_X1 U2351 ( .A1(n40946), .A2(n22593), .ZN(n59238) );
  AND2_X1 U2354 ( .A1(n57791), .A2(n12384), .Z(n39098) );
  NAND2_X1 U2363 ( .A1(n39028), .A2(n40728), .ZN(n12922) );
  INV_X1 U2364 ( .I(n40721), .ZN(n40634) );
  OAI21_X1 U2365 ( .A1(n7237), .A2(n7501), .B(n8394), .ZN(n41134) );
  NAND3_X1 U2366 ( .A1(n42450), .A2(n753), .A3(n42451), .ZN(n59155) );
  NAND3_X1 U2369 ( .A1(n16749), .A2(n40349), .A3(n17945), .ZN(n58305) );
  BUF_X2 U2394 ( .I(n60075), .Z(n22776) );
  BUF_X2 U2397 ( .I(n1402), .Z(n58262) );
  INV_X1 U2417 ( .I(n40663), .ZN(n39143) );
  NAND2_X1 U2432 ( .A1(n7011), .A2(n23634), .ZN(n59016) );
  CLKBUF_X2 U2437 ( .I(n5980), .Z(n61394) );
  NAND3_X1 U2450 ( .A1(n61000), .A2(n6581), .A3(n40211), .ZN(n59860) );
  NOR2_X1 U2457 ( .A1(n58798), .A2(n41460), .ZN(n59026) );
  INV_X1 U2469 ( .I(n37199), .ZN(n40938) );
  NAND2_X1 U2513 ( .A1(n22638), .A2(n22832), .ZN(n41439) );
  INV_X1 U2527 ( .I(n42489), .ZN(n59851) );
  BUF_X4 U2536 ( .I(n39507), .Z(n60693) );
  NAND2_X1 U2546 ( .A1(n18706), .A2(n40998), .ZN(n40149) );
  INV_X1 U2565 ( .I(n1307), .ZN(n22285) );
  NAND2_X1 U2575 ( .A1(n16102), .A2(n25020), .ZN(n40721) );
  CLKBUF_X2 U2580 ( .I(n21050), .Z(n60929) );
  INV_X1 U2594 ( .I(n40980), .ZN(n38035) );
  NOR2_X1 U2620 ( .A1(n11188), .A2(n11187), .ZN(n9711) );
  BUF_X2 U2649 ( .I(n19184), .Z(n2355) );
  INV_X2 U2666 ( .I(n24677), .ZN(n38300) );
  NAND2_X1 U2680 ( .A1(n59291), .A2(n35903), .ZN(n14909) );
  AOI22_X1 U2699 ( .A1(n59135), .A2(n59137), .B1(n15831), .B2(n35903), .ZN(
        n7859) );
  OAI21_X1 U2714 ( .A1(n12116), .A2(n3856), .B(n22559), .ZN(n34111) );
  NOR2_X1 U2720 ( .A1(n35122), .A2(n36408), .ZN(n57616) );
  NOR3_X1 U2728 ( .A1(n37274), .A2(n58257), .A3(n37272), .ZN(n37284) );
  NOR2_X1 U2774 ( .A1(n58335), .A2(n35895), .ZN(n26064) );
  NAND3_X1 U2775 ( .A1(n25339), .A2(n37404), .A3(n35268), .ZN(n35269) );
  NAND3_X1 U2779 ( .A1(n37368), .A2(n37367), .A3(n37366), .ZN(n26222) );
  OAI21_X1 U2783 ( .A1(n13768), .A2(n59645), .B(n22116), .ZN(n34474) );
  NOR2_X1 U2797 ( .A1(n36940), .A2(n504), .ZN(n59325) );
  NOR3_X1 U2808 ( .A1(n32982), .A2(n58161), .A3(n36091), .ZN(n9744) );
  NAND2_X1 U2810 ( .A1(n21467), .A2(n64679), .ZN(n34937) );
  NAND3_X1 U2814 ( .A1(n36969), .A2(n37240), .A3(n36968), .ZN(n12461) );
  NAND2_X1 U2825 ( .A1(n35964), .A2(n57444), .ZN(n59645) );
  INV_X1 U2827 ( .I(n7103), .ZN(n58924) );
  OAI22_X1 U2831 ( .A1(n36575), .A2(n24102), .B1(n32981), .B2(n18850), .ZN(
        n58161) );
  INV_X1 U2842 ( .I(n36072), .ZN(n58772) );
  NOR2_X1 U2858 ( .A1(n33609), .A2(n59562), .ZN(n17396) );
  OAI21_X1 U2864 ( .A1(n10254), .A2(n35583), .B(n35582), .ZN(n35584) );
  NOR2_X1 U2913 ( .A1(n12652), .A2(n36959), .ZN(n36278) );
  NAND3_X1 U2930 ( .A1(n35439), .A2(n35438), .A3(n35443), .ZN(n58594) );
  NOR2_X1 U2933 ( .A1(n23503), .A2(n35363), .ZN(n59562) );
  NAND2_X1 U2934 ( .A1(n57443), .A2(n8356), .ZN(n36093) );
  NAND2_X1 U2936 ( .A1(n22595), .A2(n22461), .ZN(n57573) );
  NAND2_X1 U2951 ( .A1(n24118), .A2(n35885), .ZN(n57768) );
  NOR2_X1 U2954 ( .A1(n21584), .A2(n58062), .ZN(n3012) );
  NAND3_X1 U2968 ( .A1(n4305), .A2(n59229), .A3(n3561), .ZN(n35502) );
  NAND2_X1 U2973 ( .A1(n35352), .A2(n21018), .ZN(n20134) );
  NOR3_X1 U2974 ( .A1(n1781), .A2(n1530), .A3(n60694), .ZN(n11593) );
  NOR2_X1 U2977 ( .A1(n35059), .A2(n57209), .ZN(n60440) );
  OAI22_X1 U3024 ( .A1(n35056), .A2(n35057), .B1(n36966), .B2(n36620), .ZN(
        n59657) );
  NAND3_X1 U3031 ( .A1(n21467), .A2(n35346), .A3(n36198), .ZN(n35349) );
  NOR2_X1 U3033 ( .A1(n24198), .A2(n24358), .ZN(n11893) );
  NAND2_X1 U3037 ( .A1(n6440), .A2(n60325), .ZN(n36547) );
  INV_X1 U3046 ( .I(n19507), .ZN(n58026) );
  AND2_X1 U3047 ( .A1(n25261), .A2(n36377), .Z(n57443) );
  NAND2_X1 U3074 ( .A1(n10601), .A2(n24924), .ZN(n33609) );
  NAND3_X1 U3113 ( .A1(n14904), .A2(n35909), .A3(n37030), .ZN(n13247) );
  BUF_X2 U3153 ( .I(n37441), .Z(n22801) );
  NAND2_X1 U3189 ( .A1(n37425), .A2(n22503), .ZN(n35935) );
  OAI21_X1 U3191 ( .A1(n37420), .A2(n35937), .B(n22461), .ZN(n34818) );
  NOR2_X1 U3212 ( .A1(n37404), .A2(n16501), .ZN(n58933) );
  NAND2_X1 U3221 ( .A1(n35936), .A2(n35943), .ZN(n3768) );
  NOR2_X1 U3230 ( .A1(n4798), .A2(n21921), .ZN(n35932) );
  NOR2_X1 U3240 ( .A1(n37428), .A2(n37425), .ZN(n35936) );
  INV_X2 U3286 ( .I(n36451), .ZN(n1531) );
  AOI21_X1 U3299 ( .A1(n16556), .A2(n34391), .B(n34390), .ZN(n37106) );
  OAI21_X1 U3321 ( .A1(n32946), .A2(n57619), .B(n57618), .ZN(n31907) );
  NAND3_X1 U3401 ( .A1(n58105), .A2(n35611), .A3(n58533), .ZN(n22976) );
  NAND2_X1 U3402 ( .A1(n60685), .A2(n60683), .ZN(n32841) );
  NOR3_X1 U3404 ( .A1(n32214), .A2(n32213), .A3(n60404), .ZN(n32215) );
  NAND2_X1 U3406 ( .A1(n33456), .A2(n9459), .ZN(n60872) );
  AOI22_X1 U3452 ( .A1(n32838), .A2(n32837), .B1(n32836), .B2(n61795), .ZN(
        n32839) );
  NAND3_X1 U3459 ( .A1(n61648), .A2(n33462), .A3(n60413), .ZN(n32956) );
  NOR2_X1 U3467 ( .A1(n14156), .A2(n32435), .ZN(n34770) );
  NAND4_X1 U3476 ( .A1(n33421), .A2(n2635), .A3(n34614), .A4(n33420), .ZN(
        n14285) );
  OR2_X1 U3477 ( .A1(n33995), .A2(n19825), .Z(n19824) );
  NAND2_X1 U3478 ( .A1(n59676), .A2(n34752), .ZN(n34270) );
  NAND3_X1 U3483 ( .A1(n33794), .A2(n33793), .A3(n35646), .ZN(n7610) );
  NAND3_X1 U3487 ( .A1(n7183), .A2(n22598), .A3(n33649), .ZN(n32822) );
  NOR2_X1 U3488 ( .A1(n14269), .A2(n33635), .ZN(n57991) );
  AOI21_X1 U3489 ( .A1(n33433), .A2(n33432), .B(n20835), .ZN(n57535) );
  OAI21_X1 U3490 ( .A1(n21969), .A2(n33977), .B(n34607), .ZN(n59847) );
  NAND3_X1 U3492 ( .A1(n60295), .A2(n35320), .A3(n35252), .ZN(n60294) );
  BUF_X2 U3504 ( .I(n7932), .Z(n560) );
  NAND2_X1 U3505 ( .A1(n19246), .A2(n34546), .ZN(n34965) );
  OR2_X1 U3506 ( .A1(n34198), .A2(n33995), .Z(n17342) );
  NAND2_X1 U3518 ( .A1(n32900), .A2(n61195), .ZN(n34159) );
  NAND2_X1 U3525 ( .A1(n35254), .A2(n16402), .ZN(n60295) );
  NAND2_X1 U3526 ( .A1(n32917), .A2(n34962), .ZN(n3670) );
  OAI22_X1 U3529 ( .A1(n2122), .A2(n33494), .B1(n34275), .B2(n57338), .ZN(
        n13088) );
  NAND2_X1 U3536 ( .A1(n34998), .A2(n34997), .ZN(n61287) );
  INV_X2 U3549 ( .I(n34640), .ZN(n61452) );
  NAND2_X1 U3552 ( .A1(n6867), .A2(n1424), .ZN(n1532) );
  INV_X1 U3554 ( .I(n35735), .ZN(n60175) );
  INV_X1 U3556 ( .I(n34763), .ZN(n57571) );
  NOR2_X1 U3562 ( .A1(n34640), .A2(n25999), .ZN(n34642) );
  NAND2_X1 U3570 ( .A1(n57940), .A2(n61795), .ZN(n33714) );
  NAND3_X1 U3576 ( .A1(n35031), .A2(n24485), .A3(n34640), .ZN(n57907) );
  NOR2_X1 U3583 ( .A1(n33561), .A2(n32807), .ZN(n33699) );
  NOR2_X1 U3591 ( .A1(n127), .A2(n34972), .ZN(n33513) );
  NAND2_X1 U3592 ( .A1(n33319), .A2(n18180), .ZN(n35207) );
  NAND2_X1 U3595 ( .A1(n32975), .A2(n33776), .ZN(n32976) );
  INV_X2 U3605 ( .I(n25658), .ZN(n34632) );
  INV_X1 U3617 ( .I(n32357), .ZN(n60654) );
  BUF_X2 U3622 ( .I(n26023), .Z(n59701) );
  INV_X1 U3625 ( .I(n32617), .ZN(n60173) );
  INV_X1 U3626 ( .I(n8073), .ZN(n20719) );
  NOR2_X1 U3632 ( .A1(n26652), .A2(n30956), .ZN(n32242) );
  INV_X1 U3646 ( .I(n23768), .ZN(n60580) );
  INV_X1 U3651 ( .I(n38388), .ZN(n50498) );
  NAND2_X1 U3661 ( .A1(n30559), .A2(n60627), .ZN(n60626) );
  AOI21_X1 U3662 ( .A1(n29451), .A2(n60031), .B(n60030), .ZN(n7981) );
  OAI21_X1 U3664 ( .A1(n65120), .A2(n28994), .B(n8706), .ZN(n8704) );
  OAI21_X1 U3682 ( .A1(n27635), .A2(n30396), .B(n2795), .ZN(n4062) );
  NOR2_X1 U3685 ( .A1(n57271), .A2(n59735), .ZN(n59734) );
  NAND2_X1 U3694 ( .A1(n7736), .A2(n7737), .ZN(n57499) );
  NAND3_X1 U3695 ( .A1(n59770), .A2(n30016), .A3(n30014), .ZN(n30017) );
  NOR2_X1 U3696 ( .A1(n57796), .A2(n57558), .ZN(n348) );
  NOR2_X1 U3700 ( .A1(n8960), .A2(n8959), .ZN(n58681) );
  NOR2_X1 U3701 ( .A1(n16631), .A2(n30252), .ZN(n60849) );
  NAND4_X1 U3702 ( .A1(n29004), .A2(n23446), .A3(n10068), .A4(n57381), .ZN(
        n59684) );
  INV_X1 U3706 ( .I(n61629), .ZN(n60627) );
  INV_X1 U3713 ( .I(n30759), .ZN(n31214) );
  NAND2_X1 U3716 ( .A1(n30876), .A2(n30875), .ZN(n30508) );
  NAND2_X1 U3717 ( .A1(n61229), .A2(n30812), .ZN(n58387) );
  OAI22_X1 U3724 ( .A1(n28685), .A2(n57436), .B1(n28687), .B2(n30181), .ZN(
        n58019) );
  OAI22_X1 U3726 ( .A1(n29927), .A2(n26508), .B1(n26507), .B2(n61187), .ZN(
        n58092) );
  NAND2_X1 U3733 ( .A1(n27724), .A2(n31146), .ZN(n60110) );
  AND2_X1 U3746 ( .A1(n6343), .A2(n30740), .Z(n57328) );
  NOR2_X1 U3762 ( .A1(n28703), .A2(n30396), .ZN(n24851) );
  OAI21_X1 U3763 ( .A1(n29552), .A2(n29553), .B(n30767), .ZN(n29554) );
  OAI21_X1 U3770 ( .A1(n30005), .A2(n30006), .B(n23799), .ZN(n30011) );
  AOI21_X1 U3771 ( .A1(n30780), .A2(n30782), .B(n61335), .ZN(n17482) );
  OAI21_X1 U3774 ( .A1(n24172), .A2(n60109), .B(n7461), .ZN(n60108) );
  OAI22_X1 U3775 ( .A1(n58422), .A2(n495), .B1(n31146), .B2(n31145), .ZN(
        n31148) );
  INV_X1 U3777 ( .I(n29841), .ZN(n29840) );
  INV_X1 U3778 ( .I(n26441), .ZN(n61335) );
  NOR2_X1 U3779 ( .A1(n30702), .A2(n6349), .ZN(n19887) );
  AND2_X1 U3780 ( .A1(n1866), .A2(n63906), .Z(n29906) );
  OR2_X1 U3784 ( .A1(n29516), .A2(n17413), .Z(n29096) );
  INV_X1 U3785 ( .I(n30739), .ZN(n59365) );
  NAND2_X1 U3789 ( .A1(n60895), .A2(n31085), .ZN(n5594) );
  NAND2_X1 U3795 ( .A1(n6149), .A2(n23446), .ZN(n30394) );
  NAND2_X1 U3798 ( .A1(n31137), .A2(n5768), .ZN(n60109) );
  NAND4_X1 U3804 ( .A1(n30293), .A2(n8218), .A3(n23988), .A4(n1317), .ZN(
        n57566) );
  NOR2_X1 U3806 ( .A1(n64565), .A2(n29858), .ZN(n58766) );
  AOI21_X1 U3812 ( .A1(n30659), .A2(n62285), .B(n30333), .ZN(n21676) );
  BUF_X2 U3815 ( .I(n26084), .Z(n59841) );
  NOR3_X1 U3820 ( .A1(n4567), .A2(n1433), .A3(n24123), .ZN(n29935) );
  AND2_X1 U3822 ( .A1(n27516), .A2(n30722), .Z(n28772) );
  INV_X1 U3826 ( .I(n22513), .ZN(n6090) );
  BUF_X2 U3829 ( .I(n31144), .Z(n495) );
  NOR2_X1 U3834 ( .A1(n25698), .A2(n30252), .ZN(n30258) );
  NAND2_X1 U3836 ( .A1(n31049), .A2(n31053), .ZN(n30063) );
  AND2_X1 U3839 ( .A1(n59798), .A2(n64950), .Z(n29043) );
  INV_X1 U3842 ( .I(n29879), .ZN(n27739) );
  BUF_X2 U3846 ( .I(n31147), .Z(n59810) );
  NAND3_X1 U3852 ( .A1(n31044), .A2(n30167), .A3(n31059), .ZN(n30169) );
  NOR2_X1 U3867 ( .A1(n27516), .A2(n30730), .ZN(n30266) );
  NAND2_X1 U3870 ( .A1(n15407), .A2(n60111), .ZN(n31044) );
  BUF_X2 U3876 ( .I(n30845), .Z(n23589) );
  NAND2_X1 U3880 ( .A1(n28347), .A2(n57368), .ZN(n58654) );
  NOR2_X1 U3887 ( .A1(n19565), .A2(n28148), .ZN(n28848) );
  AOI21_X1 U3891 ( .A1(n58596), .A2(n26737), .B(n27853), .ZN(n19371) );
  OAI22_X1 U3895 ( .A1(n10239), .A2(n27717), .B1(n25858), .B2(n18848), .ZN(
        n15880) );
  OR4_X1 U3896 ( .A1(n15763), .A2(n64809), .A3(n28533), .A4(n64337), .Z(n57259) );
  INV_X1 U3898 ( .I(n28477), .ZN(n57915) );
  NAND2_X1 U3899 ( .A1(n26736), .A2(n15896), .ZN(n58596) );
  NOR3_X1 U3908 ( .A1(n27255), .A2(n7354), .A3(n15763), .ZN(n57648) );
  NOR3_X1 U3920 ( .A1(n9751), .A2(n28401), .A3(n2569), .ZN(n16222) );
  OR2_X1 U3928 ( .A1(n1362), .A2(n29662), .Z(n57270) );
  AND2_X1 U3931 ( .A1(n28178), .A2(n28676), .Z(n57411) );
  NAND2_X1 U3932 ( .A1(n60541), .A2(n26827), .ZN(n26901) );
  NOR2_X1 U3936 ( .A1(n29291), .A2(n29290), .ZN(n60198) );
  NOR2_X1 U3937 ( .A1(n27250), .A2(n64809), .ZN(n57576) );
  NAND2_X1 U3938 ( .A1(n26977), .A2(n57429), .ZN(n26700) );
  NOR2_X1 U3939 ( .A1(n29630), .A2(n29632), .ZN(n60479) );
  NOR2_X1 U3944 ( .A1(n10399), .A2(n28216), .ZN(n60457) );
  INV_X1 U3951 ( .I(n26926), .ZN(n29309) );
  NAND3_X1 U3952 ( .A1(n16523), .A2(n27470), .A3(n27486), .ZN(n61179) );
  INV_X1 U3959 ( .I(n27249), .ZN(n28541) );
  NOR2_X1 U3970 ( .A1(n29286), .A2(n28128), .ZN(n29627) );
  INV_X1 U3974 ( .I(n555), .ZN(n60767) );
  OR2_X1 U3975 ( .A1(n29352), .A2(n29338), .Z(n57429) );
  OR2_X1 U3977 ( .A1(n29372), .A2(n28813), .Z(n57306) );
  NAND3_X1 U3978 ( .A1(n28842), .A2(n19593), .A3(n20907), .ZN(n19783) );
  CLKBUF_X2 U3999 ( .I(n3256), .Z(n2789) );
  BUF_X2 U4007 ( .I(n21154), .Z(n60885) );
  BUF_X2 U4012 ( .I(n27033), .Z(n29171) );
  NOR2_X2 U4017 ( .A1(n54447), .A2(n54441), .ZN(n54818) );
  BUF_X4 U4018 ( .I(n51891), .Z(n55896) );
  AOI22_X2 U4024 ( .A1(n54819), .A2(n54818), .B1(n54817), .B2(n54816), .ZN(
        n54832) );
  NOR2_X2 U4031 ( .A1(n56936), .A2(n14708), .ZN(n17850) );
  NAND2_X1 U4039 ( .A1(n37206), .A2(n37219), .ZN(n57541) );
  NAND2_X2 U4053 ( .A1(n9111), .A2(n23447), .ZN(n56267) );
  NAND3_X1 U4054 ( .A1(n58104), .A2(n41915), .A3(n11316), .ZN(n13091) );
  INV_X2 U4058 ( .I(n16525), .ZN(n57876) );
  CLKBUF_X2 U4076 ( .I(n22900), .Z(n59713) );
  OAI22_X1 U4083 ( .A1(n57201), .A2(n22122), .B1(n54699), .B2(n54698), .ZN(
        n54701) );
  NAND3_X1 U4096 ( .A1(n55416), .A2(n55255), .A3(n55401), .ZN(n55257) );
  NAND2_X1 U4102 ( .A1(n55412), .A2(n55401), .ZN(n52910) );
  OR2_X1 U4113 ( .A1(n46824), .A2(n10475), .Z(n47139) );
  CLKBUF_X2 U4124 ( .I(n25170), .Z(n4985) );
  NOR2_X1 U4136 ( .A1(n14056), .A2(n15454), .ZN(n59792) );
  NAND2_X1 U4137 ( .A1(n54379), .A2(n15202), .ZN(n4154) );
  NOR2_X1 U4143 ( .A1(n13757), .A2(n13920), .ZN(n51437) );
  NAND2_X1 U4154 ( .A1(n56789), .A2(n56790), .ZN(n61613) );
  NAND2_X1 U4161 ( .A1(n21860), .A2(n23163), .ZN(n56520) );
  BUF_X2 U4168 ( .I(n21860), .Z(n10286) );
  AOI22_X1 U4169 ( .A1(n16995), .A2(n55232), .B1(n55233), .B2(n55234), .ZN(
        n55239) );
  INV_X2 U4187 ( .I(n53056), .ZN(n1281) );
  NOR2_X1 U4190 ( .A1(n16342), .A2(n22925), .ZN(n55813) );
  NAND2_X1 U4193 ( .A1(n16342), .A2(n20447), .ZN(n55759) );
  OAI21_X1 U4207 ( .A1(n57183), .A2(n60310), .B(n52763), .ZN(n52765) );
  AOI21_X1 U4230 ( .A1(n54333), .A2(n61463), .B(n59422), .ZN(n59421) );
  NAND2_X1 U4249 ( .A1(n56817), .A2(n23030), .ZN(n60811) );
  CLKBUF_X1 U4250 ( .I(n16935), .Z(n59370) );
  NOR3_X1 U4254 ( .A1(n36558), .A2(n64405), .A3(n24102), .ZN(n32982) );
  NOR3_X1 U4258 ( .A1(n48472), .A2(n60390), .A3(n2499), .ZN(n48473) );
  NAND2_X1 U4272 ( .A1(n54983), .A2(n16948), .ZN(n55418) );
  NOR2_X1 U4284 ( .A1(n34841), .A2(n37492), .ZN(n7269) );
  NAND2_X1 U4302 ( .A1(n4617), .A2(n27229), .ZN(n60033) );
  NAND3_X1 U4310 ( .A1(n51452), .A2(n51451), .A3(n56627), .ZN(n51454) );
  NAND2_X1 U4313 ( .A1(n55575), .A2(n55597), .ZN(n55530) );
  NAND2_X1 U4320 ( .A1(n48688), .A2(n10636), .ZN(n49060) );
  CLKBUF_X4 U4327 ( .I(n52032), .Z(n24455) );
  AND2_X1 U4330 ( .A1(n56407), .A2(n7274), .Z(n57347) );
  CLKBUF_X2 U4338 ( .I(n55768), .Z(n22933) );
  INV_X2 U4340 ( .I(n25510), .ZN(n54409) );
  NOR2_X1 U4353 ( .A1(n49467), .A2(n49742), .ZN(n57816) );
  OAI21_X1 U4359 ( .A1(n10030), .A2(n49459), .B(n16239), .ZN(n49742) );
  CLKBUF_X4 U4367 ( .I(n26200), .Z(n61472) );
  NOR2_X1 U4389 ( .A1(n53083), .A2(n53094), .ZN(n53096) );
  NOR2_X1 U4397 ( .A1(n10033), .A2(n10032), .ZN(n22752) );
  NAND3_X1 U4401 ( .A1(n55322), .A2(n52488), .A3(n14927), .ZN(n5049) );
  NAND2_X1 U4408 ( .A1(n1580), .A2(n1582), .ZN(n12045) );
  NOR2_X1 U4411 ( .A1(n7138), .A2(n54424), .ZN(n54419) );
  BUF_X2 U4418 ( .I(n6747), .Z(n508) );
  NAND2_X1 U4429 ( .A1(n47501), .A2(n863), .ZN(n45482) );
  INV_X2 U4436 ( .I(n57182), .ZN(n50284) );
  NAND2_X1 U4438 ( .A1(n50292), .A2(n57182), .ZN(n50119) );
  AOI21_X1 U4443 ( .A1(n57182), .A2(n60487), .B(n50286), .ZN(n16494) );
  NAND2_X1 U4451 ( .A1(n20601), .A2(n43161), .ZN(n20603) );
  INV_X1 U4454 ( .I(n36299), .ZN(n23432) );
  NAND2_X1 U4455 ( .A1(n35403), .A2(n36299), .ZN(n11636) );
  CLKBUF_X2 U4456 ( .I(n12930), .Z(n2905) );
  INV_X2 U4466 ( .I(n55235), .ZN(n16995) );
  AOI21_X1 U4468 ( .A1(n35045), .A2(n35033), .B(n35032), .ZN(n35034) );
  OAI21_X1 U4472 ( .A1(n54205), .A2(n54204), .B(n54203), .ZN(n13708) );
  NAND2_X1 U4473 ( .A1(n7148), .A2(n54459), .ZN(n23562) );
  OAI21_X1 U4494 ( .A1(n15853), .A2(n55225), .B(n22466), .ZN(n52969) );
  INV_X2 U4496 ( .I(n41007), .ZN(n1275) );
  CLKBUF_X4 U4501 ( .I(n7955), .Z(n7680) );
  NAND2_X1 U4509 ( .A1(n29516), .A2(n29521), .ZN(n16665) );
  NOR2_X1 U4512 ( .A1(n10286), .A2(n19999), .ZN(n56484) );
  OAI21_X1 U4515 ( .A1(n47696), .A2(n47809), .B(n23180), .ZN(n2901) );
  INV_X1 U4520 ( .I(n20547), .ZN(n53396) );
  OR2_X1 U4525 ( .A1(n52738), .A2(n12573), .Z(n57407) );
  INV_X1 U4533 ( .I(n33467), .ZN(n24589) );
  AOI21_X1 U4538 ( .A1(n31780), .A2(n1420), .B(n35887), .ZN(n31784) );
  OAI21_X1 U4552 ( .A1(n1765), .A2(n13928), .B(n5105), .ZN(n7957) );
  NOR3_X1 U4567 ( .A1(n54916), .A2(n12689), .A3(n12688), .ZN(n54919) );
  NOR2_X1 U4576 ( .A1(n18196), .A2(n22852), .ZN(n6173) );
  NOR2_X1 U4577 ( .A1(n18196), .A2(n47985), .ZN(n47231) );
  INV_X2 U4578 ( .I(n18196), .ZN(n46946) );
  NAND4_X1 U4580 ( .A1(n54056), .A2(n54059), .A3(n54057), .A4(n550), .ZN(
        n54060) );
  INV_X1 U4595 ( .I(n5550), .ZN(n55925) );
  OAI22_X1 U4601 ( .A1(n42431), .A2(n40061), .B1(n42433), .B2(n40060), .ZN(
        n40062) );
  NAND2_X1 U4606 ( .A1(n57876), .A2(n18006), .ZN(n25043) );
  NAND2_X1 U4611 ( .A1(n57876), .A2(n28497), .ZN(n57875) );
  NOR2_X1 U4613 ( .A1(n24207), .A2(n45970), .ZN(n59044) );
  OAI22_X1 U4614 ( .A1(n13881), .A2(n3663), .B1(n45967), .B2(n13879), .ZN(
        n45970) );
  INV_X2 U4623 ( .I(n45614), .ZN(n16379) );
  BUF_X2 U4625 ( .I(n45614), .Z(n49843) );
  NOR2_X1 U4626 ( .A1(n55575), .A2(n1592), .ZN(n55549) );
  INV_X2 U4645 ( .I(n55503), .ZN(n55590) );
  BUF_X4 U4646 ( .I(n55503), .Z(n55575) );
  NOR3_X1 U4656 ( .A1(n46014), .A2(n46016), .A3(n47296), .ZN(n24597) );
  NAND2_X1 U4659 ( .A1(n49903), .A2(n4417), .ZN(n4664) );
  NAND2_X1 U4661 ( .A1(n49903), .A2(n19243), .ZN(n47793) );
  NAND3_X1 U4676 ( .A1(n48760), .A2(n48759), .A3(n48758), .ZN(n48761) );
  NOR2_X1 U4685 ( .A1(n2005), .A2(n29747), .ZN(n29547) );
  NOR2_X1 U4687 ( .A1(n50397), .A2(n49419), .ZN(n60464) );
  NAND2_X1 U4688 ( .A1(n50397), .A2(n22764), .ZN(n49030) );
  NAND2_X1 U4694 ( .A1(n20351), .A2(n43924), .ZN(n43915) );
  NOR2_X1 U4699 ( .A1(n30332), .A2(n23901), .ZN(n3898) );
  NAND2_X1 U4700 ( .A1(n57037), .A2(n8850), .ZN(n25490) );
  AOI21_X1 U4702 ( .A1(n53440), .A2(n57037), .B(n7095), .ZN(n53441) );
  NAND2_X1 U4722 ( .A1(n54338), .A2(n59052), .ZN(n59422) );
  NAND3_X1 U4724 ( .A1(n5569), .A2(n54996), .A3(n5279), .ZN(n54844) );
  AOI21_X1 U4726 ( .A1(n55727), .A2(n2104), .B(n55278), .ZN(n52190) );
  BUF_X4 U4741 ( .I(n52794), .Z(n53351) );
  INV_X1 U4742 ( .I(n52794), .ZN(n53369) );
  NAND3_X1 U4762 ( .A1(n57414), .A2(n55244), .A3(n55416), .ZN(n57805) );
  INV_X2 U4763 ( .I(n7007), .ZN(n24181) );
  AOI21_X1 U4769 ( .A1(n34382), .A2(n34386), .B(n15453), .ZN(n15452) );
  INV_X1 U4770 ( .I(n34386), .ZN(n35282) );
  NOR2_X1 U4782 ( .A1(n23708), .A2(n5267), .ZN(n30429) );
  NAND2_X1 U4784 ( .A1(n5267), .A2(n29472), .ZN(n31084) );
  NAND2_X1 U4790 ( .A1(n30606), .A2(n30623), .ZN(n59202) );
  NAND2_X1 U4802 ( .A1(n13038), .A2(n61673), .ZN(n12752) );
  INV_X1 U4806 ( .I(n28018), .ZN(n61055) );
  AOI22_X1 U4809 ( .A1(n54823), .A2(n6311), .B1(n54822), .B2(n54821), .ZN(
        n54831) );
  OAI21_X1 U4811 ( .A1(n36090), .A2(n8356), .B(n59105), .ZN(n59104) );
  NAND2_X1 U4813 ( .A1(n19707), .A2(n1583), .ZN(n56973) );
  NOR2_X1 U4824 ( .A1(n40943), .A2(n39102), .ZN(n39106) );
  CLKBUF_X2 U4825 ( .I(n39102), .Z(n58351) );
  INV_X1 U4829 ( .I(n52380), .ZN(n54938) );
  INV_X1 U4830 ( .I(n49549), .ZN(n8347) );
  AOI21_X1 U4835 ( .A1(n9914), .A2(n42667), .B(n11883), .ZN(n42664) );
  INV_X1 U4845 ( .I(n47013), .ZN(n48600) );
  BUF_X2 U4846 ( .I(n33879), .Z(n22476) );
  INV_X1 U4847 ( .I(n46916), .ZN(n60632) );
  NAND2_X1 U4854 ( .A1(n24353), .A2(n52819), .ZN(n57040) );
  NAND4_X1 U4856 ( .A1(n31598), .A2(n34148), .A3(n32845), .A4(n34151), .ZN(
        n31606) );
  NAND2_X1 U4861 ( .A1(n15040), .A2(n54815), .ZN(n54443) );
  NAND2_X1 U4874 ( .A1(n43844), .A2(n43069), .ZN(n23485) );
  INV_X2 U4876 ( .I(n43069), .ZN(n43845) );
  NAND2_X1 U4885 ( .A1(n57845), .A2(n27907), .ZN(n57679) );
  OAI21_X1 U4886 ( .A1(n46727), .A2(n59200), .B(n46729), .ZN(n8990) );
  NAND3_X1 U4890 ( .A1(n54402), .A2(n7138), .A3(n54414), .ZN(n54404) );
  CLKBUF_X4 U4902 ( .I(n33863), .Z(n23719) );
  NAND4_X1 U4907 ( .A1(n56652), .A2(n56653), .A3(n56654), .A4(n56651), .ZN(
        n60419) );
  INV_X1 U4912 ( .I(n34000), .ZN(n34654) );
  OAI21_X1 U4913 ( .A1(n34000), .A2(n34179), .B(n23947), .ZN(n31474) );
  AOI21_X1 U4917 ( .A1(n33999), .A2(n34180), .B(n34000), .ZN(n4548) );
  NOR2_X1 U4923 ( .A1(n53505), .A2(n25789), .ZN(n6080) );
  INV_X2 U4931 ( .I(n24405), .ZN(n59309) );
  NAND2_X1 U4932 ( .A1(n27529), .A2(n28342), .ZN(n27210) );
  NOR2_X1 U4939 ( .A1(n60232), .A2(n2403), .ZN(n47153) );
  INV_X1 U4942 ( .I(n60232), .ZN(n46177) );
  NAND2_X1 U5002 ( .A1(n40842), .A2(n59409), .ZN(n40588) );
  NAND2_X1 U5009 ( .A1(n35145), .A2(n35355), .ZN(n60691) );
  CLKBUF_X2 U5022 ( .I(n51035), .Z(n22584) );
  AOI21_X1 U5027 ( .A1(n17958), .A2(n20989), .B(n17538), .ZN(n34265) );
  AOI21_X1 U5036 ( .A1(n35533), .A2(n22785), .B(n36564), .ZN(n35538) );
  INV_X1 U5067 ( .I(n1237), .ZN(n60601) );
  OAI21_X1 U5071 ( .A1(n48757), .A2(n63876), .B(n50421), .ZN(n48760) );
  NAND2_X1 U5072 ( .A1(n50427), .A2(n58336), .ZN(n19367) );
  OAI21_X1 U5077 ( .A1(n53384), .A2(n11041), .B(n23169), .ZN(n50675) );
  CLKBUF_X1 U5107 ( .I(n37939), .Z(n14971) );
  CLKBUF_X1 U5111 ( .I(n62027), .Z(n24927) );
  BUF_X2 U5113 ( .I(n28406), .Z(n9751) );
  INV_X2 U5114 ( .I(n28406), .ZN(n28007) );
  INV_X1 U5115 ( .I(n6780), .ZN(n17533) );
  INV_X1 U5124 ( .I(n60839), .ZN(n48662) );
  NAND3_X1 U5125 ( .A1(n60839), .A2(n48246), .A3(n60838), .ZN(n16703) );
  NOR2_X1 U5127 ( .A1(n10364), .A2(n16757), .ZN(n18757) );
  INV_X2 U5144 ( .I(n7846), .ZN(n14931) );
  CLKBUF_X4 U5149 ( .I(n33862), .Z(n23690) );
  INV_X1 U5151 ( .I(n34119), .ZN(n34114) );
  OR2_X2 U5152 ( .A1(n4591), .A2(n9369), .Z(n57164) );
  INV_X2 U5155 ( .I(n13126), .ZN(n37425) );
  OR2_X2 U5156 ( .A1(n8178), .A2(n15046), .Z(n34358) );
  NAND2_X1 U5157 ( .A1(n35031), .A2(n15756), .ZN(n5123) );
  OR2_X2 U5171 ( .A1(n12480), .A2(n1428), .Z(n57166) );
  XNOR2_X1 U5174 ( .A1(n46671), .A2(n32276), .ZN(n57167) );
  AND2_X1 U5177 ( .A1(n35286), .A2(n35750), .Z(n57168) );
  OR2_X1 U5178 ( .A1(n35307), .A2(n21487), .Z(n57169) );
  NAND2_X2 U5191 ( .A1(n13699), .A2(n20060), .ZN(n34852) );
  INV_X2 U5195 ( .I(n37197), .ZN(n40923) );
  NAND2_X2 U5196 ( .A1(n57207), .A2(n6058), .ZN(n41857) );
  INV_X2 U5199 ( .I(n10044), .ZN(n61477) );
  BUF_X2 U5200 ( .I(n38264), .Z(n3534) );
  AND2_X2 U5203 ( .A1(n2469), .A2(n59495), .Z(n41234) );
  INV_X2 U5208 ( .I(n61653), .ZN(n5531) );
  BUF_X2 U5209 ( .I(n16755), .Z(n21050) );
  XNOR2_X1 U5210 ( .A1(n39190), .A2(n39191), .ZN(n57174) );
  AND2_X1 U5211 ( .A1(n3090), .A2(n42230), .Z(n57175) );
  INV_X1 U5215 ( .I(n43844), .ZN(n4689) );
  CLKBUF_X12 U5219 ( .I(n23003), .Z(n60657) );
  NAND2_X2 U5225 ( .A1(n15478), .A2(n41793), .ZN(n3656) );
  OR2_X2 U5229 ( .A1(n42846), .A2(n24361), .Z(n57178) );
  OR2_X1 U5232 ( .A1(n41544), .A2(n59771), .Z(n57179) );
  BUF_X4 U5234 ( .I(n6564), .Z(n2036) );
  NOR2_X1 U5235 ( .A1(n13871), .A2(n13872), .ZN(n21650) );
  INV_X2 U5246 ( .I(n24475), .ZN(n47843) );
  NAND2_X2 U5252 ( .A1(n9907), .A2(n47502), .ZN(n12687) );
  BUF_X2 U5253 ( .I(n47653), .Z(n23405) );
  INV_X2 U5257 ( .I(n2025), .ZN(n58232) );
  INV_X1 U5263 ( .I(n22780), .ZN(n49501) );
  AND2_X2 U5281 ( .A1(n23533), .A2(n15741), .Z(n57182) );
  AND2_X2 U5286 ( .A1(n15777), .A2(n12944), .Z(n56412) );
  OR2_X2 U5290 ( .A1(n53226), .A2(n25747), .Z(n57183) );
  INV_X2 U5296 ( .I(n56341), .ZN(n25393) );
  INV_X4 U5299 ( .I(n23756), .ZN(n14354) );
  OR2_X1 U5302 ( .A1(n7200), .A2(n55228), .Z(n57186) );
  OAI22_X1 U5310 ( .A1(n26823), .A2(n57875), .B1(n27655), .B2(n26074), .ZN(
        n26395) );
  NAND2_X1 U5315 ( .A1(n23017), .A2(n23863), .ZN(n42716) );
  INV_X2 U5317 ( .I(n23017), .ZN(n25328) );
  NOR2_X1 U5322 ( .A1(n25261), .A2(n36377), .ZN(n35533) );
  CLKBUF_X12 U5327 ( .I(n1313), .Z(n60118) );
  NAND2_X1 U5329 ( .A1(n42651), .A2(n24024), .ZN(n43357) );
  AOI22_X2 U5343 ( .A1(n28819), .A2(n28818), .B1(n28817), .B2(n28816), .ZN(
        n28820) );
  OR2_X1 U5346 ( .A1(n61728), .A2(n48074), .Z(n48067) );
  CLKBUF_X1 U5347 ( .I(n13548), .Z(n9491) );
  OR2_X2 U5354 ( .A1(n57197), .A2(n25458), .Z(n18407) );
  NAND3_X1 U5355 ( .A1(n42944), .A2(n25458), .A3(n42049), .ZN(n58678) );
  INV_X2 U5358 ( .I(n11056), .ZN(n4370) );
  AOI21_X1 U5369 ( .A1(n57735), .A2(n49779), .B(n4271), .ZN(n22172) );
  NAND2_X1 U5376 ( .A1(n23334), .A2(n56545), .ZN(n58510) );
  BUF_X2 U5378 ( .I(n38796), .Z(n60597) );
  AND2_X2 U5400 ( .A1(n9880), .A2(n14733), .Z(n12412) );
  BUF_X4 U5402 ( .I(n15723), .Z(n41182) );
  NAND2_X1 U5410 ( .A1(n37441), .A2(n7074), .ZN(n36971) );
  INV_X2 U5411 ( .I(n37441), .ZN(n37454) );
  NAND2_X1 U5421 ( .A1(n138), .A2(n61567), .ZN(n10038) );
  NAND2_X1 U5432 ( .A1(n56888), .A2(n60708), .ZN(n60781) );
  BUF_X4 U5438 ( .I(n23603), .Z(n2984) );
  CLKBUF_X2 U5439 ( .I(n25393), .Z(n60353) );
  INV_X1 U5441 ( .I(n22864), .ZN(n58812) );
  AND2_X1 U5442 ( .A1(n2037), .A2(n20735), .Z(n61690) );
  CLKBUF_X2 U5456 ( .I(n11841), .Z(n61627) );
  NOR2_X1 U5466 ( .A1(n61412), .A2(n52980), .ZN(n61411) );
  AOI21_X1 U5469 ( .A1(n61559), .A2(n61558), .B(n7303), .ZN(n23921) );
  NAND2_X1 U5470 ( .A1(n485), .A2(n61413), .ZN(n61412) );
  AND3_X1 U5475 ( .A1(n52573), .A2(n55415), .A3(n54786), .Z(n57468) );
  INV_X1 U5479 ( .I(n53409), .ZN(n61413) );
  NOR3_X1 U5481 ( .A1(n20802), .A2(n19499), .A3(n57325), .ZN(n60530) );
  NAND2_X1 U5483 ( .A1(n56391), .A2(n56567), .ZN(n58040) );
  NAND2_X1 U5485 ( .A1(n54079), .A2(n54471), .ZN(n59928) );
  NOR2_X1 U5486 ( .A1(n54597), .A2(n54325), .ZN(n7789) );
  NOR2_X1 U5495 ( .A1(n54047), .A2(n54036), .ZN(n58005) );
  NAND2_X1 U5499 ( .A1(n56571), .A2(n11121), .ZN(n58039) );
  NOR2_X1 U5500 ( .A1(n56592), .A2(n56408), .ZN(n57948) );
  CLKBUF_X2 U5501 ( .I(n53537), .Z(n60105) );
  NAND2_X1 U5505 ( .A1(n22775), .A2(n53848), .ZN(n59812) );
  NAND3_X1 U5506 ( .A1(n59951), .A2(n507), .A3(n57070), .ZN(n52850) );
  CLKBUF_X1 U5515 ( .I(n55966), .Z(n61182) );
  CLKBUF_X2 U5516 ( .I(n55692), .Z(n59040) );
  CLKBUF_X2 U5521 ( .I(n52281), .Z(n7213) );
  CLKBUF_X2 U5529 ( .I(n22550), .Z(n61502) );
  CLKBUF_X2 U5530 ( .I(n1139), .Z(n59879) );
  CLKBUF_X2 U5533 ( .I(n5236), .Z(n58373) );
  CLKBUF_X2 U5539 ( .I(n56624), .Z(n59449) );
  CLKBUF_X2 U5550 ( .I(n56544), .Z(n23334) );
  BUF_X2 U5551 ( .I(n51855), .Z(n54072) );
  INV_X2 U5556 ( .I(n53377), .ZN(n57192) );
  CLKBUF_X2 U5558 ( .I(n19890), .Z(n60448) );
  CLKBUF_X2 U5561 ( .I(n50385), .Z(n57644) );
  INV_X1 U5568 ( .I(n9044), .ZN(n59464) );
  CLKBUF_X2 U5569 ( .I(n50949), .Z(n58341) );
  AND2_X1 U5574 ( .A1(n15471), .A2(n14007), .Z(n57419) );
  NAND2_X1 U5578 ( .A1(n48951), .A2(n49777), .ZN(n61069) );
  OAI22_X1 U5583 ( .A1(n12629), .A2(n50099), .B1(n49044), .B2(n49619), .ZN(
        n58880) );
  AOI21_X1 U5607 ( .A1(n3737), .A2(n57296), .B(n48385), .ZN(n17693) );
  NAND2_X1 U5612 ( .A1(n47994), .A2(n18833), .ZN(n23373) );
  INV_X1 U5613 ( .I(n50354), .ZN(n60539) );
  OR2_X1 U5614 ( .A1(n1205), .A2(n49459), .Z(n57312) );
  NAND2_X1 U5616 ( .A1(n9240), .A2(n24362), .ZN(n58377) );
  AND2_X1 U5618 ( .A1(n24692), .A2(n1636), .Z(n57296) );
  CLKBUF_X2 U5630 ( .I(n47075), .Z(n60730) );
  BUF_X2 U5635 ( .I(n8044), .Z(n59808) );
  OR2_X1 U5645 ( .A1(n58297), .A2(n21362), .Z(n48952) );
  NOR2_X1 U5663 ( .A1(n57945), .A2(n44713), .ZN(n10376) );
  CLKBUF_X8 U5665 ( .I(n44793), .Z(n57194) );
  CLKBUF_X2 U5671 ( .I(n7318), .Z(n61422) );
  NAND3_X1 U5672 ( .A1(n47531), .A2(n9152), .A3(n60343), .ZN(n60342) );
  AOI21_X1 U5684 ( .A1(n45179), .A2(n47723), .B(n57635), .ZN(n57634) );
  AOI21_X1 U5689 ( .A1(n45752), .A2(n60727), .B(n5979), .ZN(n58845) );
  NAND2_X1 U5696 ( .A1(n23617), .A2(n46762), .ZN(n46764) );
  NAND2_X1 U5708 ( .A1(n46755), .A2(n57739), .ZN(n46756) );
  OAI21_X1 U5712 ( .A1(n47428), .A2(n59205), .B(n46840), .ZN(n12069) );
  INV_X1 U5716 ( .I(n47014), .ZN(n18510) );
  NOR2_X1 U5734 ( .A1(n61543), .A2(n59698), .ZN(n59697) );
  NAND2_X1 U5738 ( .A1(n48194), .A2(n48208), .ZN(n59775) );
  CLKBUF_X2 U5740 ( .I(n3942), .Z(n61166) );
  CLKBUF_X2 U5742 ( .I(n47154), .Z(n4655) );
  CLKBUF_X1 U5745 ( .I(n6034), .Z(n57839) );
  INV_X2 U5746 ( .I(n48232), .ZN(n57195) );
  CLKBUF_X1 U5776 ( .I(n47429), .Z(n61216) );
  CLKBUF_X2 U5781 ( .I(n46753), .Z(n57973) );
  BUF_X2 U5785 ( .I(n46314), .Z(n47541) );
  CLKBUF_X2 U5800 ( .I(n46507), .Z(n61363) );
  CLKBUF_X2 U5817 ( .I(n44851), .Z(n60918) );
  NAND2_X1 U5824 ( .A1(n59737), .A2(n57788), .ZN(n57827) );
  OAI21_X1 U5826 ( .A1(n57282), .A2(n43851), .B(n59655), .ZN(n43084) );
  NOR2_X1 U5831 ( .A1(n57178), .A2(n23811), .ZN(n59232) );
  NOR2_X1 U5837 ( .A1(n42345), .A2(n17706), .ZN(n6043) );
  NAND2_X1 U5847 ( .A1(n43661), .A2(n59889), .ZN(n59888) );
  NOR3_X1 U5851 ( .A1(n43603), .A2(n57335), .A3(n13107), .ZN(n43609) );
  INV_X1 U5854 ( .I(n42824), .ZN(n58086) );
  OAI21_X1 U5860 ( .A1(n13036), .A2(n2824), .B(n43655), .ZN(n59889) );
  NOR2_X1 U5863 ( .A1(n18958), .A2(n57283), .ZN(n60916) );
  NAND2_X1 U5865 ( .A1(n41676), .A2(n42319), .ZN(n59703) );
  NOR2_X1 U5869 ( .A1(n21138), .A2(n12064), .ZN(n21137) );
  INV_X1 U5872 ( .I(n42385), .ZN(n1700) );
  AOI21_X1 U5873 ( .A1(n59416), .A2(n59415), .B(n43573), .ZN(n2626) );
  CLKBUF_X4 U5884 ( .I(n24024), .Z(n4322) );
  NAND2_X1 U5899 ( .A1(n57974), .A2(n18126), .ZN(n13385) );
  OR2_X1 U5900 ( .A1(n42985), .A2(n42986), .Z(n43958) );
  AOI21_X1 U5916 ( .A1(n20277), .A2(n38269), .B(n59985), .ZN(n38272) );
  NAND2_X1 U5918 ( .A1(n37931), .A2(n40470), .ZN(n59885) );
  AOI21_X1 U5923 ( .A1(n40540), .A2(n40539), .B(n58981), .ZN(n3871) );
  OAI22_X1 U5927 ( .A1(n59281), .A2(n59280), .B1(n7928), .B2(n41301), .ZN(
        n7923) );
  OAI21_X1 U5932 ( .A1(n42299), .A2(n57207), .B(n41857), .ZN(n3536) );
  AND2_X1 U5944 ( .A1(n40491), .A2(n40484), .Z(n57303) );
  AOI21_X1 U5946 ( .A1(n59195), .A2(n59199), .B(n59193), .ZN(n2164) );
  NAND2_X1 U5950 ( .A1(n57389), .A2(n12453), .ZN(n58771) );
  NOR2_X1 U5958 ( .A1(n7927), .A2(n7926), .ZN(n59281) );
  AOI21_X1 U5962 ( .A1(n39698), .A2(n41122), .B(n39697), .ZN(n61125) );
  NAND2_X1 U5963 ( .A1(n57309), .A2(n39995), .ZN(n59730) );
  INV_X1 U5964 ( .I(n40983), .ZN(n10307) );
  OR2_X1 U5965 ( .A1(n24606), .A2(n40840), .Z(n57389) );
  NAND2_X1 U5968 ( .A1(n41888), .A2(n41887), .ZN(n41890) );
  NAND2_X1 U5969 ( .A1(n41294), .A2(n60947), .ZN(n16079) );
  NAND3_X1 U5972 ( .A1(n61000), .A2(n40154), .A3(n1509), .ZN(n59120) );
  INV_X1 U5973 ( .I(n12057), .ZN(n18341) );
  NOR2_X1 U5977 ( .A1(n41168), .A2(n40645), .ZN(n61183) );
  NAND3_X1 U5979 ( .A1(n40996), .A2(n40213), .A3(n40146), .ZN(n5395) );
  NOR2_X1 U5987 ( .A1(n11126), .A2(n24188), .ZN(n59193) );
  INV_X2 U5998 ( .I(n40484), .ZN(n40653) );
  NOR2_X1 U5999 ( .A1(n41017), .A2(n61308), .ZN(n24742) );
  AND2_X1 U6001 ( .A1(n23492), .A2(n22304), .Z(n57406) );
  OR2_X1 U6007 ( .A1(n41376), .A2(n10074), .Z(n57309) );
  OR2_X1 U6008 ( .A1(n17212), .A2(n12158), .Z(n57257) );
  CLKBUF_X2 U6032 ( .I(n40770), .Z(n57615) );
  BUF_X2 U6033 ( .I(n17594), .Z(n58926) );
  INV_X1 U6034 ( .I(n16476), .ZN(n60221) );
  CLKBUF_X2 U6036 ( .I(n39732), .Z(n59788) );
  NOR2_X1 U6038 ( .A1(n60161), .A2(n17195), .ZN(n17194) );
  AOI21_X1 U6039 ( .A1(n58925), .A2(n35384), .B(n58924), .ZN(n17195) );
  INV_X1 U6041 ( .I(n36559), .ZN(n59037) );
  NOR2_X1 U6042 ( .A1(n36192), .A2(n17390), .ZN(n17389) );
  OAI21_X1 U6044 ( .A1(n35530), .A2(n35529), .B(n59104), .ZN(n35540) );
  NOR2_X1 U6048 ( .A1(n59117), .A2(n57391), .ZN(n11466) );
  NAND2_X1 U6051 ( .A1(n14925), .A2(n19245), .ZN(n58335) );
  NAND2_X1 U6059 ( .A1(n17243), .A2(n38550), .ZN(n37135) );
  NOR2_X1 U6066 ( .A1(n1788), .A2(n35883), .ZN(n60954) );
  INV_X1 U6067 ( .I(n35932), .ZN(n36873) );
  NAND2_X1 U6069 ( .A1(n11020), .A2(n15720), .ZN(n57838) );
  CLKBUF_X2 U6080 ( .I(n25124), .Z(n59852) );
  BUF_X2 U6086 ( .I(n35086), .Z(n22223) );
  CLKBUF_X4 U6087 ( .I(n17775), .Z(n2002) );
  INV_X1 U6088 ( .I(n16886), .ZN(n9178) );
  NAND2_X1 U6091 ( .A1(n15984), .A2(n18800), .ZN(n57947) );
  OAI21_X1 U6095 ( .A1(n31022), .A2(n33419), .B(n59847), .ZN(n31028) );
  NOR2_X1 U6109 ( .A1(n33368), .A2(n33369), .ZN(n57990) );
  NOR2_X1 U6112 ( .A1(n32864), .A2(n139), .ZN(n60245) );
  NAND2_X1 U6113 ( .A1(n35045), .A2(n57907), .ZN(n9132) );
  NAND3_X1 U6116 ( .A1(n32924), .A2(n34356), .A3(n64965), .ZN(n32925) );
  AOI21_X1 U6117 ( .A1(n33364), .A2(n22601), .B(n34151), .ZN(n57696) );
  OAI21_X1 U6119 ( .A1(n34140), .A2(n34139), .B(n34138), .ZN(n58860) );
  NOR2_X1 U6130 ( .A1(n35214), .A2(n57986), .ZN(n4163) );
  BUF_X4 U6133 ( .I(n35667), .Z(n57200) );
  INV_X1 U6141 ( .I(n33359), .ZN(n61195) );
  BUF_X2 U6158 ( .I(n35241), .Z(n58598) );
  CLKBUF_X1 U6160 ( .I(n34018), .Z(n57774) );
  BUF_X2 U6164 ( .I(n35218), .Z(n57986) );
  CLKBUF_X2 U6165 ( .I(n15807), .Z(n59134) );
  BUF_X2 U6166 ( .I(n1342), .Z(n118) );
  CLKBUF_X1 U6174 ( .I(n31815), .Z(n59773) );
  BUF_X2 U6179 ( .I(n25856), .Z(n59163) );
  NAND4_X1 U6181 ( .A1(n19696), .A2(n28210), .A3(n61272), .A4(n9819), .ZN(
        n19695) );
  NOR2_X1 U6186 ( .A1(n57769), .A2(n29511), .ZN(n26587) );
  NAND4_X1 U6188 ( .A1(n30248), .A2(n30246), .A3(n30245), .A4(n30247), .ZN(
        n61244) );
  NAND3_X1 U6191 ( .A1(n19471), .A2(n30720), .A3(n30721), .ZN(n12661) );
  NOR2_X1 U6198 ( .A1(n29469), .A2(n31083), .ZN(n61385) );
  NOR2_X1 U6200 ( .A1(n1553), .A2(n2119), .ZN(n61043) );
  NAND2_X1 U6202 ( .A1(n29418), .A2(n30437), .ZN(n60614) );
  NAND2_X1 U6203 ( .A1(n31216), .A2(n8364), .ZN(n25120) );
  NAND2_X1 U6204 ( .A1(n8811), .A2(n60665), .ZN(n30327) );
  OAI21_X1 U6205 ( .A1(n60112), .A2(n58999), .B(n30173), .ZN(n23144) );
  CLKBUF_X4 U6207 ( .I(n30695), .Z(n60142) );
  CLKBUF_X2 U6210 ( .I(n30728), .Z(n57733) );
  BUF_X4 U6216 ( .I(n25755), .Z(n4270) );
  CLKBUF_X2 U6219 ( .I(n21222), .Z(n58630) );
  OAI21_X1 U6225 ( .A1(n1931), .A2(n60457), .B(n28217), .ZN(n2547) );
  NOR2_X1 U6226 ( .A1(n7023), .A2(n7024), .ZN(n2659) );
  AOI22_X1 U6229 ( .A1(n60183), .A2(n27951), .B1(n27955), .B2(n27954), .ZN(
        n11094) );
  BUF_X1 U6230 ( .I(n39635), .Z(n61238) );
  NAND2_X1 U6232 ( .A1(n1877), .A2(n27087), .ZN(n58588) );
  BUF_X2 U6233 ( .I(n39387), .Z(n59680) );
  NOR2_X1 U6236 ( .A1(n29108), .A2(n27949), .ZN(n60183) );
  NOR2_X1 U6237 ( .A1(n27251), .A2(n1883), .ZN(n57577) );
  INV_X1 U6238 ( .I(n60324), .ZN(n60323) );
  NAND2_X1 U6239 ( .A1(n15358), .A2(n28855), .ZN(n28158) );
  NAND3_X1 U6241 ( .A1(n23386), .A2(n61004), .A3(n6369), .ZN(n19462) );
  CLKBUF_X1 U6242 ( .I(n33134), .Z(n58928) );
  BUF_X2 U6249 ( .I(n28280), .Z(n61049) );
  BUF_X2 U6254 ( .I(n20070), .Z(n60547) );
  CLKBUF_X2 U6255 ( .I(n27171), .Z(n60818) );
  INV_X2 U6264 ( .I(n6913), .ZN(n27932) );
  CLKBUF_X2 U6269 ( .I(n29613), .Z(n61307) );
  CLKBUF_X2 U6270 ( .I(n20292), .Z(n58601) );
  BUF_X2 U6277 ( .I(n56097), .Z(n57989) );
  CLKBUF_X2 U6280 ( .I(Key[25]), .Z(n53477) );
  CLKBUF_X2 U6281 ( .I(Key[188]), .Z(n61447) );
  AOI22_X1 U6287 ( .A1(n58869), .A2(n58868), .B1(n53817), .B2(n53828), .ZN(
        n53770) );
  NAND2_X1 U6296 ( .A1(n15972), .A2(n21973), .ZN(n50820) );
  NOR3_X1 U6297 ( .A1(n7982), .A2(n7987), .A3(n7985), .ZN(n25724) );
  NAND2_X1 U6298 ( .A1(n56795), .A2(n56778), .ZN(n56779) );
  INV_X1 U6299 ( .I(n53779), .ZN(n58869) );
  INV_X1 U6301 ( .I(n21922), .ZN(n61193) );
  NAND2_X1 U6302 ( .A1(n54907), .A2(n22864), .ZN(n22863) );
  NAND2_X1 U6309 ( .A1(n55817), .A2(n14890), .ZN(n55750) );
  NAND2_X1 U6311 ( .A1(n58812), .A2(n54911), .ZN(n54900) );
  AND2_X1 U6313 ( .A1(n54571), .A2(n54572), .Z(n57334) );
  INV_X2 U6314 ( .I(n55036), .ZN(n25170) );
  CLKBUF_X2 U6316 ( .I(n53992), .Z(n59662) );
  NAND3_X1 U6317 ( .A1(n55772), .A2(n14890), .A3(n55820), .ZN(n11686) );
  CLKBUF_X8 U6318 ( .I(n55088), .Z(n25220) );
  CLKBUF_X2 U6327 ( .I(n54543), .Z(n60433) );
  BUF_X4 U6334 ( .I(n52878), .Z(n53108) );
  NAND2_X1 U6338 ( .A1(n54061), .A2(n54060), .ZN(n57698) );
  CLKBUF_X4 U6341 ( .I(n54257), .Z(n57202) );
  NAND2_X1 U6344 ( .A1(n55468), .A2(n22592), .ZN(n57675) );
  AOI21_X1 U6345 ( .A1(n13021), .A2(n1284), .B(n13018), .ZN(n56276) );
  NAND2_X1 U6354 ( .A1(n9253), .A2(n8851), .ZN(n9252) );
  NAND2_X1 U6357 ( .A1(n25447), .A2(n25446), .ZN(n59006) );
  NOR2_X1 U6362 ( .A1(n55708), .A2(n55707), .ZN(n16343) );
  NOR2_X1 U6364 ( .A1(n57985), .A2(n57372), .ZN(n14644) );
  AOI22_X1 U6366 ( .A1(n53019), .A2(n53020), .B1(n53860), .B2(n53021), .ZN(
        n59739) );
  NAND2_X1 U6368 ( .A1(n54456), .A2(n54453), .ZN(n61340) );
  NAND2_X1 U6372 ( .A1(n57191), .A2(n61492), .ZN(n5199) );
  OAI21_X1 U6373 ( .A1(n58005), .A2(n58006), .B(n58656), .ZN(n54043) );
  OAI21_X1 U6386 ( .A1(n52903), .A2(n54790), .B(n57805), .ZN(n52904) );
  OAI21_X1 U6387 ( .A1(n57347), .A2(n57948), .B(n56409), .ZN(n24311) );
  NAND2_X1 U6396 ( .A1(n54070), .A2(n57319), .ZN(n57985) );
  NAND2_X1 U6399 ( .A1(n58511), .A2(n58510), .ZN(n56548) );
  INV_X1 U6403 ( .I(n52873), .ZN(n60336) );
  OAI21_X1 U6405 ( .A1(n54945), .A2(n54605), .B(n58650), .ZN(n54606) );
  OAI21_X1 U6406 ( .A1(n52282), .A2(n56371), .B(n56372), .ZN(n52279) );
  NOR3_X1 U6417 ( .A1(n55922), .A2(n55664), .A3(n58050), .ZN(n11679) );
  OR3_X1 U6418 ( .A1(n833), .A2(n57051), .A3(n60475), .Z(n52823) );
  OR2_X1 U6420 ( .A1(n53578), .A2(n60310), .Z(n52775) );
  NAND2_X1 U6422 ( .A1(n57354), .A2(n54849), .ZN(n61698) );
  NOR2_X1 U6430 ( .A1(n2742), .A2(n16767), .ZN(n60573) );
  OAI21_X1 U6439 ( .A1(n6311), .A2(n54659), .B(n59142), .ZN(n54438) );
  AND3_X1 U6442 ( .A1(n55269), .A2(n58283), .A3(n55271), .Z(n57231) );
  NAND2_X1 U6446 ( .A1(n54780), .A2(n54605), .ZN(n58650) );
  AND2_X1 U6449 ( .A1(n24510), .A2(n54067), .Z(n57316) );
  NAND3_X1 U6453 ( .A1(n54996), .A2(n1613), .A3(n55265), .ZN(n52480) );
  AND2_X1 U6454 ( .A1(n55927), .A2(n60370), .Z(n57361) );
  OR2_X1 U6467 ( .A1(n2951), .A2(n1459), .Z(n11938) );
  CLKBUF_X2 U6475 ( .I(n54938), .Z(n60439) );
  CLKBUF_X2 U6476 ( .I(n23701), .Z(n58300) );
  BUF_X4 U6479 ( .I(n50460), .Z(n53860) );
  CLKBUF_X2 U6483 ( .I(n2199), .Z(n22231) );
  BUF_X2 U6484 ( .I(n19639), .Z(n23836) );
  CLKBUF_X2 U6485 ( .I(n56659), .Z(n59461) );
  INV_X1 U6493 ( .I(n51577), .ZN(n61464) );
  INV_X1 U6494 ( .I(n52441), .ZN(n60760) );
  INV_X1 U6495 ( .I(n51125), .ZN(n59706) );
  INV_X1 U6501 ( .I(n51997), .ZN(n58787) );
  NAND2_X1 U6508 ( .A1(n12874), .A2(n50436), .ZN(n61565) );
  BUF_X2 U6517 ( .I(n51797), .Z(n23213) );
  NOR2_X1 U6542 ( .A1(n25048), .A2(n61069), .ZN(n4825) );
  NOR2_X1 U6564 ( .A1(n16089), .A2(n48858), .ZN(n57640) );
  NAND2_X1 U6572 ( .A1(n49604), .A2(n59084), .ZN(n58461) );
  NAND3_X1 U6582 ( .A1(n59076), .A2(n49993), .A3(n49994), .ZN(n20999) );
  NAND2_X1 U6591 ( .A1(n58377), .A2(n9241), .ZN(n49644) );
  AOI22_X1 U6592 ( .A1(n48171), .A2(n58676), .B1(n48169), .B2(n48170), .ZN(
        n21465) );
  NOR2_X1 U6599 ( .A1(n10637), .A2(n60591), .ZN(n60590) );
  NOR2_X1 U6602 ( .A1(n48697), .A2(n1631), .ZN(n57639) );
  AOI22_X1 U6604 ( .A1(n49887), .A2(n50286), .B1(n49889), .B2(n49886), .ZN(
        n49895) );
  NAND2_X1 U6606 ( .A1(n60485), .A2(n60484), .ZN(n3320) );
  INV_X1 U6608 ( .I(n49002), .ZN(n58261) );
  NOR2_X1 U6610 ( .A1(n59777), .A2(n59167), .ZN(n19897) );
  NOR2_X1 U6612 ( .A1(n49741), .A2(n22526), .ZN(n57815) );
  NAND3_X1 U6617 ( .A1(n57302), .A2(n49515), .A3(n16483), .ZN(n9233) );
  NOR2_X1 U6618 ( .A1(n12838), .A2(n48417), .ZN(n59714) );
  NAND2_X1 U6620 ( .A1(n19900), .A2(n19899), .ZN(n59777) );
  OR2_X1 U6621 ( .A1(n48374), .A2(n48058), .Z(n57474) );
  NAND2_X1 U6624 ( .A1(n47760), .A2(n16211), .ZN(n60696) );
  INV_X1 U6626 ( .I(n49245), .ZN(n61235) );
  INV_X1 U6628 ( .I(n10768), .ZN(n60485) );
  NAND2_X1 U6629 ( .A1(n50012), .A2(n50214), .ZN(n60484) );
  NOR2_X1 U6630 ( .A1(n61016), .A2(n11058), .ZN(n58298) );
  NAND2_X1 U6636 ( .A1(n47966), .A2(n25018), .ZN(n61150) );
  NOR2_X1 U6638 ( .A1(n59545), .A2(n48718), .ZN(n47961) );
  NOR2_X1 U6642 ( .A1(n10080), .A2(n17446), .ZN(n61487) );
  OAI21_X1 U6643 ( .A1(n60719), .A2(n60718), .B(n57608), .ZN(n49750) );
  NAND2_X1 U6650 ( .A1(n50084), .A2(n62405), .ZN(n61540) );
  NAND2_X1 U6653 ( .A1(n21189), .A2(n1384), .ZN(n17957) );
  INV_X1 U6654 ( .I(n60378), .ZN(n50349) );
  INV_X2 U6656 ( .I(n50345), .ZN(n50336) );
  INV_X1 U6657 ( .I(n1630), .ZN(n13645) );
  INV_X1 U6666 ( .I(n49491), .ZN(n58443) );
  NAND2_X1 U6672 ( .A1(n49377), .A2(n49538), .ZN(n60592) );
  OR2_X1 U6674 ( .A1(n21183), .A2(n4174), .Z(n57224) );
  CLKBUF_X2 U6679 ( .I(n21406), .Z(n58037) );
  CLKBUF_X2 U6682 ( .I(n8994), .Z(n59200) );
  CLKBUF_X2 U6687 ( .I(n25162), .Z(n57608) );
  BUF_X2 U6691 ( .I(n50361), .Z(n23394) );
  CLKBUF_X2 U6702 ( .I(n21320), .Z(n13120) );
  CLKBUF_X2 U6709 ( .I(n24966), .Z(n60163) );
  NAND2_X1 U6725 ( .A1(n45181), .A2(n57635), .ZN(n57632) );
  NAND2_X1 U6740 ( .A1(n60631), .A2(n59447), .ZN(n59446) );
  INV_X1 U6741 ( .I(n57634), .ZN(n57633) );
  NAND2_X1 U6744 ( .A1(n45227), .A2(n45226), .ZN(n61139) );
  NAND2_X1 U6747 ( .A1(n45597), .A2(n57654), .ZN(n25637) );
  AND2_X1 U6749 ( .A1(n45653), .A2(n64878), .Z(n57369) );
  NAND2_X1 U6755 ( .A1(n2538), .A2(n4353), .ZN(n60348) );
  INV_X1 U6757 ( .I(n45667), .ZN(n45666) );
  OAI22_X1 U6762 ( .A1(n12826), .A2(n47502), .B1(n12823), .B2(n12824), .ZN(
        n44677) );
  NAND3_X1 U6770 ( .A1(n47246), .A2(n8648), .A3(n8650), .ZN(n58666) );
  NAND2_X1 U6777 ( .A1(n45646), .A2(n45647), .ZN(n58528) );
  OAI21_X1 U6780 ( .A1(n58134), .A2(n58133), .B(n23061), .ZN(n25179) );
  NAND2_X1 U6781 ( .A1(n47200), .A2(n47199), .ZN(n59557) );
  NAND2_X1 U6788 ( .A1(n46566), .A2(n4213), .ZN(n61204) );
  AOI21_X1 U6789 ( .A1(n57243), .A2(n19041), .B(n4623), .ZN(n25790) );
  OR3_X1 U6790 ( .A1(n47115), .A2(n12698), .A3(n58018), .Z(n47117) );
  NAND2_X1 U6793 ( .A1(n46765), .A2(n46770), .ZN(n60411) );
  NAND2_X1 U6799 ( .A1(n45574), .A2(n22303), .ZN(n60005) );
  INV_X1 U6803 ( .I(n46805), .ZN(n58728) );
  INV_X1 U6816 ( .I(n45495), .ZN(n57487) );
  NAND2_X1 U6817 ( .A1(n47029), .A2(n60465), .ZN(n44404) );
  INV_X1 U6824 ( .I(n59383), .ZN(n58352) );
  NAND3_X1 U6826 ( .A1(n13759), .A2(n48651), .A3(n48653), .ZN(n59153) );
  NOR2_X1 U6827 ( .A1(n57532), .A2(n57531), .ZN(n57530) );
  OAI21_X1 U6829 ( .A1(n19804), .A2(n59775), .B(n20404), .ZN(n11490) );
  NOR2_X1 U6832 ( .A1(n10005), .A2(n47809), .ZN(n59611) );
  NAND2_X1 U6833 ( .A1(n48237), .A2(n57305), .ZN(n48121) );
  CLKBUF_X2 U6834 ( .I(n48234), .Z(n59616) );
  AND2_X1 U6835 ( .A1(n8043), .A2(n48584), .Z(n57238) );
  AND2_X1 U6838 ( .A1(n44284), .A2(n21044), .Z(n57262) );
  NOR2_X1 U6846 ( .A1(n45674), .A2(n44868), .ZN(n59127) );
  OAI22_X1 U6850 ( .A1(n48519), .A2(n48645), .B1(n48514), .B2(n7834), .ZN(
        n48259) );
  AND2_X1 U6851 ( .A1(n4428), .A2(n64605), .Z(n57305) );
  AND2_X1 U6860 ( .A1(n8820), .A2(n8666), .Z(n57333) );
  CLKBUF_X2 U6865 ( .I(n47683), .Z(n59205) );
  CLKBUF_X2 U6869 ( .I(n46897), .Z(n59707) );
  CLKBUF_X2 U6872 ( .I(n8632), .Z(n60560) );
  CLKBUF_X2 U6879 ( .I(n508), .Z(n60038) );
  CLKBUF_X2 U6881 ( .I(n47308), .Z(n60893) );
  CLKBUF_X2 U6883 ( .I(n47495), .Z(n61014) );
  CLKBUF_X2 U6884 ( .I(n47725), .Z(n61510) );
  INV_X1 U6885 ( .I(n47163), .ZN(n47166) );
  NOR2_X1 U6886 ( .A1(n63547), .A2(n46794), .ZN(n57766) );
  CLKBUF_X2 U6888 ( .I(n47245), .Z(n58155) );
  INV_X1 U6894 ( .I(n47115), .ZN(n47110) );
  CLKBUF_X2 U6899 ( .I(n21090), .Z(n59861) );
  CLKBUF_X2 U6900 ( .I(n47121), .Z(n60651) );
  CLKBUF_X2 U6905 ( .I(n25580), .Z(n59802) );
  INV_X2 U6908 ( .I(n26180), .ZN(n45643) );
  BUF_X2 U6910 ( .I(n48483), .Z(n23301) );
  INV_X1 U6916 ( .I(n13658), .ZN(n60073) );
  INV_X1 U6917 ( .I(n9249), .ZN(n59228) );
  INV_X1 U6926 ( .I(n46200), .ZN(n58802) );
  CLKBUF_X2 U6932 ( .I(n46690), .Z(n58532) );
  NAND2_X1 U6933 ( .A1(n61071), .A2(n43909), .ZN(n14899) );
  CLKBUF_X2 U6937 ( .I(n10776), .Z(n60458) );
  OR2_X2 U6943 ( .A1(n25009), .A2(n22831), .Z(n5029) );
  INV_X1 U6947 ( .I(n44851), .ZN(n60999) );
  OAI22_X1 U6954 ( .A1(n40872), .A2(n57827), .B1(n57385), .B2(n57788), .ZN(
        n38061) );
  CLKBUF_X2 U6980 ( .I(n46231), .Z(n19232) );
  NAND2_X1 U6989 ( .A1(n59197), .A2(n59196), .ZN(n41535) );
  NAND2_X1 U7024 ( .A1(n41534), .A2(n5939), .ZN(n59197) );
  NAND2_X1 U7032 ( .A1(n41533), .A2(n42383), .ZN(n59196) );
  OAI21_X1 U7043 ( .A1(n6764), .A2(n42871), .B(n42343), .ZN(n59833) );
  NAND2_X1 U7052 ( .A1(n41551), .A2(n59066), .ZN(n59065) );
  NAND2_X1 U7064 ( .A1(n42887), .A2(n60952), .ZN(n60951) );
  AOI21_X1 U7065 ( .A1(n16992), .A2(n1034), .B(n58288), .ZN(n3453) );
  NAND2_X1 U7075 ( .A1(n60363), .A2(n60361), .ZN(n20851) );
  NAND2_X1 U7077 ( .A1(n42125), .A2(n42126), .ZN(n42136) );
  NOR2_X1 U7084 ( .A1(n10487), .A2(n57525), .ZN(n59276) );
  NOR3_X1 U7085 ( .A1(n41360), .A2(n58086), .A3(n41361), .ZN(n41366) );
  INV_X1 U7095 ( .I(n41775), .ZN(n59948) );
  NAND2_X1 U7104 ( .A1(n19214), .A2(n43172), .ZN(n58032) );
  NAND2_X1 U7108 ( .A1(n42735), .A2(n59067), .ZN(n42737) );
  AOI21_X1 U7116 ( .A1(n24250), .A2(n63095), .B(n42007), .ZN(n26187) );
  NAND2_X1 U7119 ( .A1(n43076), .A2(n60706), .ZN(n59655) );
  NAND2_X1 U7123 ( .A1(n61120), .A2(n61119), .ZN(n4672) );
  AND2_X1 U7141 ( .A1(n295), .A2(n42867), .Z(n57315) );
  NOR2_X1 U7147 ( .A1(n42382), .A2(n42381), .ZN(n59048) );
  OR2_X1 U7154 ( .A1(n43074), .A2(n60706), .Z(n57282) );
  NAND2_X1 U7172 ( .A1(n42848), .A2(n42849), .ZN(n59412) );
  NAND3_X1 U7173 ( .A1(n2625), .A2(n43576), .A3(n5238), .ZN(n58199) );
  NAND3_X1 U7181 ( .A1(n59288), .A2(n41567), .A3(n57651), .ZN(n41570) );
  NOR2_X1 U7182 ( .A1(n9212), .A2(n61372), .ZN(n61397) );
  INV_X1 U7197 ( .I(n7620), .ZN(n61120) );
  AOI21_X1 U7198 ( .A1(n42973), .A2(n23188), .B(n19428), .ZN(n641) );
  NOR2_X1 U7213 ( .A1(n58180), .A2(n42896), .ZN(n58179) );
  NAND2_X1 U7228 ( .A1(n43659), .A2(n43662), .ZN(n59887) );
  NAND2_X1 U7230 ( .A1(n59288), .A2(n41567), .ZN(n43378) );
  NOR2_X1 U7240 ( .A1(n41546), .A2(n42600), .ZN(n59998) );
  INV_X1 U7241 ( .I(n19271), .ZN(n42628) );
  NAND2_X1 U7244 ( .A1(n59440), .A2(n59439), .ZN(n5026) );
  CLKBUF_X2 U7247 ( .I(n7285), .Z(n60472) );
  INV_X1 U7255 ( .I(n41627), .ZN(n58872) );
  CLKBUF_X1 U7256 ( .I(n42598), .Z(n59898) );
  BUF_X4 U7260 ( .I(n43099), .Z(n24250) );
  NAND2_X1 U7263 ( .A1(n295), .A2(n42871), .ZN(n59946) );
  NAND2_X1 U7270 ( .A1(n42911), .A2(n42923), .ZN(n59440) );
  NOR2_X1 U7278 ( .A1(n23488), .A2(n43925), .ZN(n59491) );
  CLKBUF_X2 U7279 ( .I(n6995), .Z(n60593) );
  CLKBUF_X2 U7290 ( .I(n43844), .Z(n57591) );
  INV_X1 U7299 ( .I(n43448), .ZN(n58850) );
  BUF_X4 U7305 ( .I(n40020), .Z(n43439) );
  INV_X1 U7326 ( .I(n39824), .ZN(n60471) );
  INV_X1 U7329 ( .I(n41648), .ZN(n60948) );
  NAND2_X1 U7336 ( .A1(n59885), .A2(n59375), .ZN(n37933) );
  CLKBUF_X2 U7337 ( .I(n4077), .Z(n57808) );
  BUF_X4 U7340 ( .I(n40096), .Z(n42968) );
  CLKBUF_X2 U7347 ( .I(n42008), .Z(n59381) );
  INV_X1 U7351 ( .I(n6799), .ZN(n60216) );
  NOR2_X1 U7372 ( .A1(n58584), .A2(n58583), .ZN(n13468) );
  CLKBUF_X2 U7377 ( .I(n40651), .Z(n57886) );
  NAND2_X1 U7389 ( .A1(n19276), .A2(n2800), .ZN(n59190) );
  NAND2_X1 U7407 ( .A1(n61626), .A2(n2164), .ZN(n2162) );
  NAND2_X1 U7462 ( .A1(n59376), .A2(n40923), .ZN(n59375) );
  OAI21_X1 U7466 ( .A1(n41919), .A2(n5642), .B(n12057), .ZN(n60619) );
  NAND2_X1 U7494 ( .A1(n16400), .A2(n16391), .ZN(n61292) );
  OAI21_X1 U7498 ( .A1(n39997), .A2(n39995), .B(n59730), .ZN(n11588) );
  NAND2_X1 U7501 ( .A1(n9954), .A2(n41279), .ZN(n38267) );
  NAND2_X1 U7503 ( .A1(n9184), .A2(n36652), .ZN(n59093) );
  NAND2_X1 U7519 ( .A1(n42270), .A2(n42271), .ZN(n57890) );
  AOI22_X1 U7525 ( .A1(n41150), .A2(n60810), .B1(n41149), .B2(n11631), .ZN(
        n15943) );
  NOR2_X1 U7538 ( .A1(n57244), .A2(n61291), .ZN(n61290) );
  NOR2_X1 U7548 ( .A1(n40088), .A2(n40089), .ZN(n61291) );
  NAND2_X1 U7551 ( .A1(n41060), .A2(n41061), .ZN(n17479) );
  INV_X1 U7556 ( .I(n8201), .ZN(n59982) );
  NOR2_X1 U7557 ( .A1(n8017), .A2(n3078), .ZN(n57655) );
  NAND2_X1 U7561 ( .A1(n42268), .A2(n42269), .ZN(n57889) );
  NAND2_X1 U7563 ( .A1(n40993), .A2(n6766), .ZN(n60219) );
  INV_X4 U7580 ( .I(n42507), .ZN(n57207) );
  NOR2_X1 U7582 ( .A1(n222), .A2(n59583), .ZN(n41053) );
  CLKBUF_X2 U7599 ( .I(n3356), .Z(n59062) );
  INV_X1 U7601 ( .I(n40163), .ZN(n59195) );
  INV_X1 U7603 ( .I(n39111), .ZN(n40116) );
  INV_X2 U7606 ( .I(n22738), .ZN(n21295) );
  NAND2_X1 U7610 ( .A1(n41466), .A2(n41467), .ZN(n61519) );
  CLKBUF_X2 U7621 ( .I(n19458), .Z(n60166) );
  CLKBUF_X2 U7630 ( .I(n42484), .Z(n61264) );
  CLKBUF_X2 U7636 ( .I(n40315), .Z(n60422) );
  INV_X1 U7642 ( .I(n41439), .ZN(n40374) );
  CLKBUF_X2 U7652 ( .I(n20871), .Z(n60172) );
  CLKBUF_X2 U7656 ( .I(n40229), .Z(n60153) );
  CLKBUF_X2 U7662 ( .I(n40995), .Z(n61005) );
  CLKBUF_X2 U7666 ( .I(n40132), .Z(n57955) );
  CLKBUF_X2 U7667 ( .I(n21920), .Z(n59674) );
  CLKBUF_X2 U7668 ( .I(n41152), .Z(n58996) );
  CLKBUF_X4 U7673 ( .I(n37199), .Z(n40924) );
  BUF_X4 U7683 ( .I(n1307), .Z(n57208) );
  INV_X1 U7689 ( .I(n38820), .ZN(n57606) );
  INV_X1 U7692 ( .I(n26021), .ZN(n58293) );
  INV_X1 U7694 ( .I(n1753), .ZN(n59284) );
  CLKBUF_X2 U7704 ( .I(n39659), .Z(n58972) );
  BUF_X2 U7705 ( .I(n2788), .Z(n2191) );
  CLKBUF_X2 U7712 ( .I(n37866), .Z(n57836) );
  CLKBUF_X2 U7714 ( .I(n11636), .Z(n60141) );
  CLKBUF_X2 U7724 ( .I(n21239), .Z(n57755) );
  CLKBUF_X2 U7728 ( .I(n38510), .Z(n59688) );
  OAI21_X1 U7739 ( .A1(n18602), .A2(n36415), .B(n59631), .ZN(n20791) );
  OAI21_X1 U7748 ( .A1(n60823), .A2(n25919), .B(n36731), .ZN(n25918) );
  NOR2_X1 U7758 ( .A1(n22474), .A2(n59632), .ZN(n59631) );
  NAND2_X1 U7760 ( .A1(n35138), .A2(n35137), .ZN(n35139) );
  NAND2_X1 U7764 ( .A1(n31788), .A2(n31787), .ZN(n58557) );
  NAND2_X1 U7781 ( .A1(n33326), .A2(n2594), .ZN(n59123) );
  INV_X1 U7789 ( .I(n59117), .ZN(n16112) );
  NAND2_X1 U7792 ( .A1(n34885), .A2(n36259), .ZN(n60636) );
  NAND2_X1 U7796 ( .A1(n11593), .A2(n36278), .ZN(n60084) );
  OAI21_X1 U7803 ( .A1(n37437), .A2(n37425), .B(n57944), .ZN(n37440) );
  INV_X1 U7804 ( .I(n18207), .ZN(n59208) );
  NOR3_X1 U7807 ( .A1(n36873), .A2(n36874), .A3(n21881), .ZN(n59244) );
  INV_X1 U7813 ( .I(n33121), .ZN(n58925) );
  NOR2_X1 U7815 ( .A1(n36884), .A2(n36883), .ZN(n57972) );
  NAND2_X1 U7819 ( .A1(n35547), .A2(n35964), .ZN(n58898) );
  INV_X1 U7820 ( .I(n36196), .ZN(n59632) );
  NOR2_X1 U7821 ( .A1(n60953), .A2(n35884), .ZN(n13171) );
  NOR2_X1 U7828 ( .A1(n20504), .A2(n36947), .ZN(n59326) );
  AOI22_X1 U7834 ( .A1(n35469), .A2(n35465), .B1(n58267), .B2(n35476), .ZN(
        n60771) );
  NAND2_X1 U7837 ( .A1(n35890), .A2(n60954), .ZN(n60953) );
  NOR2_X1 U7838 ( .A1(n35350), .A2(n57838), .ZN(n57837) );
  NAND2_X1 U7841 ( .A1(n37439), .A2(n37425), .ZN(n57944) );
  INV_X1 U7843 ( .I(n37324), .ZN(n32149) );
  NAND2_X1 U7846 ( .A1(n37069), .A2(n37070), .ZN(n61631) );
  NAND2_X1 U7848 ( .A1(n37457), .A2(n461), .ZN(n57960) );
  NAND2_X1 U7850 ( .A1(n37456), .A2(n37455), .ZN(n57962) );
  INV_X1 U7852 ( .I(n35560), .ZN(n21131) );
  INV_X1 U7854 ( .I(n36964), .ZN(n9675) );
  NAND2_X1 U7855 ( .A1(n35450), .A2(n1786), .ZN(n35057) );
  NOR2_X1 U7858 ( .A1(n37457), .A2(n36882), .ZN(n57971) );
  NAND2_X1 U7870 ( .A1(n35995), .A2(n23778), .ZN(n58400) );
  INV_X1 U7878 ( .I(n36673), .ZN(n60824) );
  INV_X1 U7879 ( .I(n57656), .ZN(n36129) );
  INV_X1 U7880 ( .I(n63742), .ZN(n58162) );
  INV_X1 U7881 ( .I(n58062), .ZN(n36695) );
  NAND2_X1 U7882 ( .A1(n36252), .A2(n22431), .ZN(n57828) );
  BUF_X4 U7908 ( .I(n37035), .Z(n21010) );
  CLKBUF_X2 U7910 ( .I(n13734), .Z(n60507) );
  INV_X1 U7926 ( .I(n59147), .ZN(n34942) );
  CLKBUF_X8 U7934 ( .I(n14054), .Z(n57209) );
  CLKBUF_X2 U7941 ( .I(n60014), .Z(n59912) );
  CLKBUF_X8 U7943 ( .I(n11160), .Z(n57210) );
  NOR2_X1 U7946 ( .A1(n59462), .A2(n25909), .ZN(n25907) );
  NOR2_X1 U7948 ( .A1(n19794), .A2(n31718), .ZN(n58172) );
  CLKBUF_X8 U7950 ( .I(n8697), .Z(n57211) );
  NAND2_X1 U7951 ( .A1(n57729), .A2(n21046), .ZN(n33297) );
  NAND2_X1 U7962 ( .A1(n34774), .A2(n34773), .ZN(n59462) );
  NOR2_X1 U7973 ( .A1(n60024), .A2(n4493), .ZN(n59057) );
  NOR2_X1 U7980 ( .A1(n35255), .A2(n60294), .ZN(n35262) );
  NAND2_X1 U7987 ( .A1(n32768), .A2(n59711), .ZN(n4493) );
  NAND2_X1 U7988 ( .A1(n33615), .A2(n33616), .ZN(n60275) );
  NAND2_X1 U7990 ( .A1(n34645), .A2(n34644), .ZN(n58001) );
  INV_X1 U7991 ( .I(n59874), .ZN(n59873) );
  OAI22_X1 U7992 ( .A1(n34715), .A2(n23556), .B1(n34716), .B2(n34714), .ZN(
        n61337) );
  INV_X1 U7999 ( .I(n58860), .ZN(n6920) );
  OAI21_X1 U8006 ( .A1(n57571), .A2(n32946), .B(n34216), .ZN(n2390) );
  INV_X1 U8026 ( .I(n11403), .ZN(n33436) );
  AND3_X1 U8032 ( .A1(n34195), .A2(n58447), .A3(n34201), .Z(n57388) );
  AOI21_X1 U8033 ( .A1(n34130), .A2(n34131), .B(n59347), .ZN(n59346) );
  NAND2_X1 U8034 ( .A1(n5732), .A2(n5733), .ZN(n57940) );
  AOI21_X1 U8036 ( .A1(n1345), .A2(n34571), .B(n8552), .ZN(n15088) );
  NAND2_X1 U8037 ( .A1(n32766), .A2(n32767), .ZN(n60024) );
  INV_X1 U8040 ( .I(n33638), .ZN(n33637) );
  INV_X1 U8042 ( .I(n35618), .ZN(n58533) );
  INV_X1 U8044 ( .I(n1532), .ZN(n34986) );
  INV_X1 U8049 ( .I(n33791), .ZN(n58186) );
  CLKBUF_X4 U8059 ( .I(n34167), .Z(n60554) );
  INV_X1 U8060 ( .I(n33537), .ZN(n59121) );
  BUF_X2 U8063 ( .I(n4097), .Z(n60700) );
  CLKBUF_X2 U8067 ( .I(n32955), .Z(n60413) );
  CLKBUF_X2 U8069 ( .I(n34088), .Z(n58421) );
  INV_X1 U8070 ( .I(n21849), .ZN(n61500) );
  BUF_X2 U8082 ( .I(n6686), .Z(n2674) );
  CLKBUF_X2 U8085 ( .I(n17255), .Z(n57546) );
  BUF_X2 U8086 ( .I(n12954), .Z(n12953) );
  AND2_X1 U8087 ( .A1(n34980), .A2(n2033), .Z(n57304) );
  CLKBUF_X2 U8088 ( .I(n13559), .Z(n9648) );
  CLKBUF_X2 U8091 ( .I(n23945), .Z(n59328) );
  NAND2_X1 U8096 ( .A1(n10504), .A2(n35755), .ZN(n61532) );
  INV_X1 U8105 ( .I(n32496), .ZN(n60302) );
  INV_X1 U8110 ( .I(n32645), .ZN(n58718) );
  INV_X1 U8113 ( .I(n24254), .ZN(n24255) );
  INV_X1 U8120 ( .I(n32237), .ZN(n60023) );
  INV_X1 U8121 ( .I(n30354), .ZN(n58775) );
  CLKBUF_X2 U8125 ( .I(n33869), .Z(n708) );
  CLKBUF_X2 U8134 ( .I(n33283), .Z(n60514) );
  CLKBUF_X2 U8136 ( .I(n33173), .Z(n61304) );
  NAND2_X1 U8137 ( .A1(n23135), .A2(n59589), .ZN(n30826) );
  NAND2_X1 U8146 ( .A1(n27770), .A2(n27773), .ZN(n59790) );
  CLKBUF_X2 U8150 ( .I(n32234), .Z(n60565) );
  CLKBUF_X2 U8153 ( .I(n22978), .Z(n60372) );
  AND2_X1 U8154 ( .A1(n14272), .A2(n14275), .Z(n10235) );
  NAND2_X1 U8159 ( .A1(n61044), .A2(n61043), .ZN(n6796) );
  NAND2_X1 U8160 ( .A1(n60626), .A2(n60625), .ZN(n30433) );
  NAND2_X1 U8168 ( .A1(n29535), .A2(n29534), .ZN(n61314) );
  INV_X1 U8170 ( .I(n30327), .ZN(n61044) );
  AND2_X1 U8175 ( .A1(n30074), .A2(n7735), .Z(n57219) );
  NAND2_X1 U8176 ( .A1(n822), .A2(n60185), .ZN(n2376) );
  NAND3_X1 U8180 ( .A1(n59151), .A2(n64962), .A3(n29800), .ZN(n2731) );
  INV_X1 U8181 ( .I(n29743), .ZN(n30773) );
  NAND2_X1 U8187 ( .A1(n61534), .A2(n30286), .ZN(n61533) );
  INV_X1 U8194 ( .I(n29047), .ZN(n57796) );
  INV_X1 U8195 ( .I(n27634), .ZN(n57769) );
  NOR2_X1 U8213 ( .A1(n29997), .A2(n2101), .ZN(n60249) );
  INV_X1 U8214 ( .I(n29485), .ZN(n5860) );
  NOR2_X1 U8215 ( .A1(n30424), .A2(n30425), .ZN(n57721) );
  NOR2_X1 U8216 ( .A1(n13339), .A2(n13338), .ZN(n59561) );
  NAND2_X1 U8222 ( .A1(n31204), .A2(n30631), .ZN(n59366) );
  INV_X1 U8232 ( .I(n30345), .ZN(n61131) );
  OAI21_X1 U8237 ( .A1(n31222), .A2(n24221), .B(n31225), .ZN(n59558) );
  NAND2_X1 U8240 ( .A1(n58423), .A2(n1437), .ZN(n58422) );
  AND2_X1 U8244 ( .A1(n30878), .A2(n31271), .Z(n57417) );
  NAND2_X1 U8251 ( .A1(n31268), .A2(n59755), .ZN(n59754) );
  NAND2_X1 U8254 ( .A1(n31209), .A2(n20378), .ZN(n3445) );
  INV_X1 U8260 ( .I(n27886), .ZN(n18005) );
  CLKBUF_X2 U8261 ( .I(n30376), .Z(n61007) );
  CLKBUF_X2 U8266 ( .I(n22696), .Z(n57806) );
  INV_X1 U8269 ( .I(n8364), .ZN(n30762) );
  CLKBUF_X2 U8270 ( .I(n25269), .Z(n60886) );
  BUF_X4 U8271 ( .I(n27626), .Z(n29779) );
  CLKBUF_X2 U8273 ( .I(n60125), .Z(n57537) );
  NOR2_X1 U8284 ( .A1(n4602), .A2(n57363), .ZN(n17175) );
  NAND2_X1 U8286 ( .A1(n26702), .A2(n26701), .ZN(n57620) );
  CLKBUF_X2 U8289 ( .I(n28959), .Z(n59541) );
  NOR2_X1 U8295 ( .A1(n20049), .A2(n7280), .ZN(n20053) );
  CLKBUF_X2 U8298 ( .I(n30125), .Z(n60009) );
  INV_X1 U8301 ( .I(n26747), .ZN(n57684) );
  AOI21_X1 U8303 ( .A1(n26773), .A2(n1355), .B(n61239), .ZN(n89) );
  NAND2_X1 U8305 ( .A1(n26616), .A2(n61320), .ZN(n61324) );
  NOR2_X1 U8306 ( .A1(n28284), .A2(n61055), .ZN(n61054) );
  NAND3_X2 U8311 ( .A1(n60537), .A2(n27254), .A3(n57259), .ZN(n26004) );
  NAND2_X1 U8314 ( .A1(n26412), .A2(n21890), .ZN(n59878) );
  NAND2_X1 U8320 ( .A1(n60155), .A2(n60154), .ZN(n27882) );
  NAND3_X1 U8325 ( .A1(n28006), .A2(n8340), .A3(n58588), .ZN(n27088) );
  NOR2_X1 U8326 ( .A1(n28848), .A2(n61006), .ZN(n26857) );
  NOR2_X1 U8329 ( .A1(n27227), .A2(n9473), .ZN(n60056) );
  AOI21_X1 U8332 ( .A1(n17878), .A2(n29366), .B(n58667), .ZN(n17876) );
  INV_X1 U8334 ( .I(n58215), .ZN(n27289) );
  NAND3_X1 U8336 ( .A1(n26480), .A2(n26479), .A3(n61179), .ZN(n20760) );
  OAI22_X1 U8337 ( .A1(n27017), .A2(n29106), .B1(n23466), .B2(n24190), .ZN(
        n4986) );
  OAI22_X1 U8344 ( .A1(n17931), .A2(n24190), .B1(n14150), .B2(n28003), .ZN(
        n2110) );
  NOR2_X1 U8349 ( .A1(n5627), .A2(n29106), .ZN(n432) );
  OAI21_X1 U8358 ( .A1(n27373), .A2(n23568), .B(n28001), .ZN(n7125) );
  NAND2_X1 U8361 ( .A1(n16272), .A2(n29130), .ZN(n58332) );
  NAND3_X1 U8368 ( .A1(n27878), .A2(n27877), .A3(n28525), .ZN(n60155) );
  NAND2_X1 U8372 ( .A1(n28590), .A2(n555), .ZN(n59089) );
  NOR2_X1 U8375 ( .A1(n5908), .A2(n5291), .ZN(n59990) );
  INV_X1 U8376 ( .I(n61491), .ZN(n61544) );
  INV_X1 U8378 ( .I(n17451), .ZN(n61599) );
  CLKBUF_X2 U8380 ( .I(n29614), .Z(n59099) );
  NAND2_X1 U8384 ( .A1(n10946), .A2(n26540), .ZN(n26329) );
  NOR2_X1 U8386 ( .A1(n6083), .A2(n29170), .ZN(n27286) );
  CLKBUF_X2 U8388 ( .I(n38277), .Z(n60207) );
  NAND2_X1 U8389 ( .A1(n61064), .A2(n28275), .ZN(n61053) );
  NOR2_X1 U8390 ( .A1(n18213), .A2(n28609), .ZN(n28438) );
  CLKBUF_X2 U8396 ( .I(n38651), .Z(n60799) );
  OR2_X1 U8403 ( .A1(n23732), .A2(n23578), .Z(n57289) );
  CLKBUF_X2 U8411 ( .I(n17339), .Z(n61045) );
  CLKBUF_X2 U8414 ( .I(n37257), .Z(n61034) );
  CLKBUF_X2 U8421 ( .I(n26362), .Z(n60816) );
  CLKBUF_X2 U8422 ( .I(n26270), .Z(n59102) );
  INV_X1 U8426 ( .I(n17221), .ZN(n60500) );
  BUF_X2 U8427 ( .I(n837), .Z(n23586) );
  CLKBUF_X2 U8429 ( .I(n29343), .Z(n23954) );
  INV_X1 U8438 ( .I(n54716), .ZN(n61401) );
  CLKBUF_X2 U8439 ( .I(Key[4]), .Z(n59130) );
  NOR2_X1 U8441 ( .A1(n10131), .A2(n60545), .ZN(n61155) );
  INV_X1 U8444 ( .I(n27573), .ZN(n9671) );
  AND2_X1 U8457 ( .A1(n8528), .A2(n4687), .Z(n26377) );
  OAI21_X1 U8470 ( .A1(n26900), .A2(n27838), .B(n61155), .ZN(n25044) );
  CLKBUF_X4 U8471 ( .I(n28870), .Z(n20240) );
  NAND2_X1 U8474 ( .A1(n28333), .A2(n28045), .ZN(n24838) );
  NAND2_X1 U8476 ( .A1(n23170), .A2(n23166), .ZN(n27998) );
  AOI22_X1 U8480 ( .A1(n29162), .A2(n29161), .B1(n12072), .B2(n64012), .ZN(
        n29165) );
  CLKBUF_X1 U8481 ( .I(n14439), .Z(n22810) );
  NOR3_X1 U8500 ( .A1(n27036), .A2(n28241), .A3(n27044), .ZN(n27039) );
  INV_X1 U8516 ( .I(n27470), .ZN(n27548) );
  OAI21_X1 U8518 ( .A1(n28838), .A2(n28126), .B(n28821), .ZN(n28133) );
  NAND2_X1 U8521 ( .A1(n26936), .A2(n25793), .ZN(n26937) );
  CLKBUF_X1 U8526 ( .I(n29641), .Z(n4812) );
  NOR2_X1 U8530 ( .A1(n26901), .A2(n61544), .ZN(n15842) );
  CLKBUF_X2 U8531 ( .I(n29691), .Z(n60603) );
  OAI21_X1 U8536 ( .A1(n60767), .A2(n60766), .B(n4988), .ZN(n6377) );
  AOI21_X1 U8545 ( .A1(n26320), .A2(n26321), .B(n26319), .ZN(n26326) );
  INV_X1 U8550 ( .I(n27419), .ZN(n12183) );
  NAND2_X1 U8578 ( .A1(n28341), .A2(n27532), .ZN(n28344) );
  CLKBUF_X2 U8581 ( .I(n3580), .Z(n60298) );
  INV_X1 U8590 ( .I(n29639), .ZN(n22443) );
  NAND2_X1 U8591 ( .A1(n8113), .A2(n29662), .ZN(n29675) );
  AND2_X1 U8606 ( .A1(n63525), .A2(n23540), .Z(n57249) );
  OAI21_X1 U8607 ( .A1(n18177), .A2(n26718), .B(n29138), .ZN(n60746) );
  NAND2_X1 U8611 ( .A1(n27690), .A2(n27812), .ZN(n27807) );
  INV_X1 U8612 ( .I(n29644), .ZN(n28847) );
  OAI21_X1 U8618 ( .A1(n28440), .A2(n5268), .B(n6257), .ZN(n7280) );
  INV_X1 U8619 ( .I(n27896), .ZN(n13416) );
  NAND2_X1 U8633 ( .A1(n23797), .A2(n29321), .ZN(n27454) );
  INV_X1 U8638 ( .I(n21281), .ZN(n27168) );
  OAI21_X1 U8645 ( .A1(n26816), .A2(n2343), .B(n26815), .ZN(n26817) );
  OAI21_X1 U8651 ( .A1(n27327), .A2(n27326), .B(n27329), .ZN(n27333) );
  NOR2_X1 U8658 ( .A1(n28805), .A2(n29372), .ZN(n29366) );
  INV_X1 U8661 ( .I(n19287), .ZN(n17688) );
  OAI21_X1 U8679 ( .A1(n31245), .A2(n1435), .B(n31247), .ZN(n31250) );
  INV_X1 U8683 ( .I(n19700), .ZN(n23564) );
  INV_X1 U8695 ( .I(n30883), .ZN(n31256) );
  NOR2_X1 U8704 ( .A1(n6859), .A2(n6862), .ZN(n6858) );
  INV_X2 U8705 ( .I(n28989), .ZN(n25898) );
  INV_X1 U8709 ( .I(n30764), .ZN(n30012) );
  OR2_X1 U8717 ( .A1(n58829), .A2(n4270), .Z(n57381) );
  INV_X1 U8718 ( .I(n8444), .ZN(n30251) );
  NOR3_X1 U8719 ( .A1(n27719), .A2(n27718), .A3(n28507), .ZN(n27720) );
  INV_X1 U8723 ( .I(n30013), .ZN(n30763) );
  INV_X1 U8735 ( .I(n18060), .ZN(n28584) );
  CLKBUF_X2 U8737 ( .I(n30736), .Z(n59096) );
  NAND3_X1 U8739 ( .A1(n29888), .A2(n31259), .A3(n29886), .ZN(n5689) );
  INV_X1 U8762 ( .I(n30439), .ZN(n27306) );
  NAND2_X1 U8767 ( .A1(n15126), .A2(n30455), .ZN(n29426) );
  NAND2_X1 U8772 ( .A1(n29500), .A2(n10068), .ZN(n29501) );
  OAI21_X1 U8781 ( .A1(n30487), .A2(n5070), .B(n6609), .ZN(n30489) );
  NAND2_X1 U8784 ( .A1(n29579), .A2(n29580), .ZN(n19885) );
  NAND2_X1 U8795 ( .A1(n30148), .A2(n16279), .ZN(n30108) );
  NAND3_X1 U8797 ( .A1(n30487), .A2(n61162), .A3(n30478), .ZN(n26710) );
  OAI21_X1 U8808 ( .A1(n26112), .A2(n5285), .B(n59810), .ZN(n27727) );
  AND3_X1 U8820 ( .A1(n13030), .A2(n19721), .A3(n30745), .Z(n59087) );
  INV_X2 U8831 ( .I(n31105), .ZN(n10734) );
  NOR2_X1 U8835 ( .A1(n1552), .A2(n30120), .ZN(n60210) );
  OAI22_X1 U8837 ( .A1(n30294), .A2(n30293), .B1(n30295), .B2(n30296), .ZN(
        n30297) );
  NAND3_X1 U8855 ( .A1(n1853), .A2(n31160), .A3(n18573), .ZN(n25990) );
  NAND2_X1 U8860 ( .A1(n31147), .A2(n57789), .ZN(n30589) );
  NOR2_X1 U8862 ( .A1(n31049), .A2(n15333), .ZN(n31061) );
  AOI21_X1 U8865 ( .A1(n19841), .A2(n30001), .B(n31211), .ZN(n11965) );
  INV_X1 U8869 ( .I(n18248), .ZN(n61403) );
  NAND2_X1 U8882 ( .A1(n29441), .A2(n6041), .ZN(n29439) );
  NOR2_X1 U8883 ( .A1(n16110), .A2(n30082), .ZN(n21405) );
  NAND2_X1 U8884 ( .A1(n15135), .A2(n29206), .ZN(n7468) );
  INV_X1 U8893 ( .I(n27735), .ZN(n27071) );
  INV_X1 U8896 ( .I(n30264), .ZN(n30727) );
  AND3_X1 U8903 ( .A1(n25013), .A2(n4257), .A3(n61251), .Z(n30513) );
  INV_X1 U8914 ( .I(n13766), .ZN(n30549) );
  CLKBUF_X2 U8916 ( .I(n23053), .Z(n58409) );
  NAND3_X1 U8922 ( .A1(n14765), .A2(n29480), .A3(n12858), .ZN(n27728) );
  NAND3_X1 U8929 ( .A1(n9001), .A2(n8999), .A3(n8998), .ZN(n59351) );
  NOR2_X1 U8930 ( .A1(n30559), .A2(n60529), .ZN(n25029) );
  AOI21_X1 U8937 ( .A1(n30728), .A2(n23772), .B(n14389), .ZN(n14384) );
  CLKBUF_X2 U8949 ( .I(n30709), .Z(n23072) );
  NAND2_X1 U8956 ( .A1(n29514), .A2(n18736), .ZN(n28748) );
  NAND3_X1 U8960 ( .A1(n30546), .A2(n1277), .A3(n30549), .ZN(n1921) );
  NAND3_X1 U8964 ( .A1(n31184), .A2(n29568), .A3(n13444), .ZN(n809) );
  NOR2_X1 U8967 ( .A1(n29906), .A2(n29905), .ZN(n30864) );
  OAI21_X1 U8974 ( .A1(n16164), .A2(n18461), .B(n13417), .ZN(n61309) );
  INV_X1 U8995 ( .I(n19535), .ZN(n31206) );
  NAND2_X1 U9001 ( .A1(n60110), .A2(n60108), .ZN(n27733) );
  INV_X1 U9012 ( .I(n23794), .ZN(n26920) );
  NOR3_X1 U9025 ( .A1(n30592), .A2(n30591), .A3(n30590), .ZN(n30596) );
  OAI21_X1 U9029 ( .A1(n6179), .A2(n6180), .B(n6178), .ZN(n3607) );
  NAND3_X1 U9034 ( .A1(n24839), .A2(n7812), .A3(n28769), .ZN(n16738) );
  AOI22_X1 U9086 ( .A1(n57417), .A2(n30877), .B1(n1857), .B2(n6317), .ZN(
        n59594) );
  CLKBUF_X1 U9091 ( .I(n61732), .Z(n58531) );
  INV_X1 U9099 ( .I(n21094), .ZN(n16401) );
  CLKBUF_X2 U9112 ( .I(n3389), .Z(n3260) );
  CLKBUF_X2 U9122 ( .I(n9977), .Z(n61538) );
  INV_X2 U9125 ( .I(n31122), .ZN(n24283) );
  CLKBUF_X2 U9128 ( .I(n21321), .Z(n17182) );
  INV_X1 U9130 ( .I(n31706), .ZN(n61279) );
  INV_X1 U9140 ( .I(n3260), .ZN(n32747) );
  INV_X1 U9145 ( .I(n14847), .ZN(n31774) );
  INV_X1 U9169 ( .I(n32392), .ZN(n58781) );
  CLKBUF_X2 U9174 ( .I(n24672), .Z(n12559) );
  INV_X1 U9181 ( .I(n59773), .ZN(n14960) );
  INV_X1 U9191 ( .I(n31612), .ZN(n60264) );
  INV_X1 U9196 ( .I(n877), .ZN(n61129) );
  INV_X1 U9215 ( .I(n35667), .ZN(n35677) );
  NOR3_X1 U9228 ( .A1(n15756), .A2(n35031), .A3(n34632), .ZN(n9131) );
  INV_X1 U9235 ( .I(n32891), .ZN(n5733) );
  INV_X1 U9241 ( .I(n15288), .ZN(n57760) );
  AOI21_X1 U9265 ( .A1(n34159), .A2(n34158), .B(n34157), .ZN(n34160) );
  NAND2_X1 U9274 ( .A1(n20785), .A2(n35026), .ZN(n17896) );
  NAND2_X1 U9313 ( .A1(n34382), .A2(n34388), .ZN(n653) );
  NAND2_X1 U9327 ( .A1(n35827), .A2(n57169), .ZN(n60900) );
  OR2_X1 U9329 ( .A1(n34194), .A2(n34193), .Z(n20313) );
  OAI21_X1 U9341 ( .A1(n35679), .A2(n32765), .B(n33601), .ZN(n59711) );
  OAI21_X1 U9343 ( .A1(n34201), .A2(n17041), .B(n34194), .ZN(n17040) );
  NAND2_X1 U9354 ( .A1(n34219), .A2(n34305), .ZN(n22253) );
  NAND2_X1 U9356 ( .A1(n34754), .A2(n34755), .ZN(n60620) );
  NOR2_X1 U9363 ( .A1(n34535), .A2(n22419), .ZN(n34528) );
  AOI21_X1 U9371 ( .A1(n33), .A2(n62045), .B(n34658), .ZN(n33998) );
  INV_X1 U9376 ( .I(n35811), .ZN(n35815) );
  NAND2_X1 U9379 ( .A1(n33950), .A2(n60892), .ZN(n34125) );
  INV_X1 U9390 ( .I(n33300), .ZN(n33303) );
  AOI21_X1 U9417 ( .A1(n34126), .A2(n31354), .B(n33944), .ZN(n31355) );
  NAND2_X1 U9424 ( .A1(n34133), .A2(n34142), .ZN(n59482) );
  NAND2_X1 U9449 ( .A1(n61287), .A2(n34999), .ZN(n35008) );
  NAND2_X1 U9451 ( .A1(n33977), .A2(n33423), .ZN(n11763) );
  CLKBUF_X1 U9459 ( .I(n24006), .Z(n57732) );
  NAND3_X1 U9463 ( .A1(n13768), .A2(n35965), .A3(n35964), .ZN(n35141) );
  NAND2_X1 U9466 ( .A1(n34304), .A2(n34219), .ZN(n2388) );
  NOR2_X1 U9481 ( .A1(n57696), .A2(n57680), .ZN(n33367) );
  AOI21_X1 U9483 ( .A1(n22063), .A2(n16155), .B(n30896), .ZN(n21908) );
  AND2_X1 U9497 ( .A1(n8029), .A2(n34658), .Z(n14669) );
  OAI22_X1 U9498 ( .A1(n32864), .A2(n32789), .B1(n34125), .B2(n1809), .ZN(
        n32791) );
  INV_X2 U9521 ( .I(n3082), .ZN(n14247) );
  AOI21_X1 U9523 ( .A1(n23777), .A2(n31297), .B(n5123), .ZN(n16234) );
  AND2_X1 U9529 ( .A1(n11347), .A2(n34472), .Z(n57444) );
  CLKBUF_X1 U9556 ( .I(n1533), .Z(n59930) );
  AOI21_X1 U9558 ( .A1(n32871), .A2(n32872), .B(n60700), .ZN(n2535) );
  OAI21_X1 U9565 ( .A1(n34086), .A2(n34628), .B(n34624), .ZN(n33441) );
  NAND2_X1 U9595 ( .A1(n37043), .A2(n1793), .ZN(n58401) );
  NOR2_X1 U9600 ( .A1(n22169), .A2(n36422), .ZN(n57656) );
  NOR2_X1 U9623 ( .A1(n20455), .A2(n34630), .ZN(n60546) );
  INV_X1 U9676 ( .I(n10317), .ZN(n36492) );
  NAND2_X1 U9679 ( .A1(n34816), .A2(n22595), .ZN(n34811) );
  NAND2_X1 U9698 ( .A1(n33579), .A2(n35214), .ZN(n33580) );
  NAND2_X1 U9712 ( .A1(n35139), .A2(n21018), .ZN(n58900) );
  NOR2_X1 U9720 ( .A1(n57210), .A2(n652), .ZN(n35464) );
  NOR2_X1 U9740 ( .A1(n10596), .A2(n1779), .ZN(n35884) );
  NAND2_X1 U9754 ( .A1(n17243), .A2(n37269), .ZN(n37132) );
  OAI21_X1 U9755 ( .A1(n35996), .A2(n58401), .B(n58400), .ZN(n58399) );
  NAND2_X1 U9762 ( .A1(n60292), .A2(n60925), .ZN(n60291) );
  NOR2_X1 U9793 ( .A1(n12110), .A2(n36233), .ZN(n36487) );
  INV_X1 U9809 ( .I(n32813), .ZN(n58504) );
  NAND2_X1 U9811 ( .A1(n22317), .A2(n37363), .ZN(n18061) );
  NAND3_X1 U9813 ( .A1(n18313), .A2(n36413), .A3(n36412), .ZN(n14264) );
  NAND2_X1 U9814 ( .A1(n35983), .A2(n15720), .ZN(n10963) );
  NOR2_X1 U9850 ( .A1(n33122), .A2(n36384), .ZN(n59607) );
  NAND2_X1 U9852 ( .A1(n35979), .A2(n35983), .ZN(n25050) );
  CLKBUF_X8 U9860 ( .I(n35882), .Z(n1779) );
  NAND2_X1 U9869 ( .A1(n34942), .A2(n36212), .ZN(n36722) );
  OAI22_X1 U9871 ( .A1(n35113), .A2(n35112), .B1(n55), .B2(n36408), .ZN(n35114) );
  INV_X1 U9878 ( .I(n36979), .ZN(n37219) );
  INV_X1 U9895 ( .I(n37273), .ZN(n58257) );
  NAND2_X1 U9903 ( .A1(n58162), .A2(n21839), .ZN(n36872) );
  NAND2_X1 U9910 ( .A1(n23503), .A2(n35363), .ZN(n36185) );
  NAND2_X1 U9919 ( .A1(n22632), .A2(n2594), .ZN(n36590) );
  AOI21_X1 U9927 ( .A1(n34851), .A2(n34852), .B(n20309), .ZN(n4510) );
  NAND2_X1 U9944 ( .A1(n17191), .A2(n35574), .ZN(n17189) );
  OAI22_X1 U9953 ( .A1(n57617), .A2(n57616), .B1(n35124), .B2(n36188), .ZN(
        n35125) );
  NAND2_X1 U9965 ( .A1(n34486), .A2(n34485), .ZN(n24398) );
  NAND3_X1 U9974 ( .A1(n35171), .A2(n35896), .A3(n34491), .ZN(n17387) );
  INV_X1 U9992 ( .I(n38806), .ZN(n61105) );
  INV_X2 U9998 ( .I(n6889), .ZN(n39722) );
  CLKBUF_X4 U10001 ( .I(n38770), .Z(n24018) );
  CLKBUF_X2 U10007 ( .I(n12381), .Z(n60039) );
  CLKBUF_X1 U10013 ( .I(n7601), .Z(n16972) );
  INV_X1 U10020 ( .I(n37686), .ZN(n18428) );
  CLKBUF_X2 U10030 ( .I(n9255), .Z(n60489) );
  INV_X1 U10039 ( .I(n21918), .ZN(n3604) );
  INV_X1 U10041 ( .I(n24223), .ZN(n21462) );
  NOR2_X1 U10043 ( .A1(n60957), .A2(n25201), .ZN(n37510) );
  NOR2_X1 U10047 ( .A1(n19990), .A2(n19611), .ZN(n25650) );
  INV_X1 U10051 ( .I(n5728), .ZN(n61149) );
  INV_X1 U10053 ( .I(n14645), .ZN(n60151) );
  NAND2_X1 U10054 ( .A1(n62106), .A2(n971), .ZN(n18421) );
  CLKBUF_X1 U10062 ( .I(n39621), .Z(n25324) );
  NOR2_X1 U10077 ( .A1(n41031), .A2(n21736), .ZN(n40515) );
  NOR2_X1 U10080 ( .A1(n40595), .A2(n64459), .ZN(n39960) );
  CLKBUF_X2 U10090 ( .I(n6932), .Z(n58970) );
  NAND2_X1 U10091 ( .A1(n40274), .A2(n9802), .ZN(n21927) );
  NAND2_X1 U10110 ( .A1(n41017), .A2(n19458), .ZN(n19078) );
  NAND2_X1 U10113 ( .A1(n41240), .A2(n61950), .ZN(n40745) );
  INV_X1 U10116 ( .I(n41816), .ZN(n21206) );
  NAND2_X1 U10123 ( .A1(n60522), .A2(n37775), .ZN(n16357) );
  NOR2_X1 U10156 ( .A1(n40092), .A2(n40316), .ZN(n40131) );
  NOR2_X1 U10171 ( .A1(n36650), .A2(n36651), .ZN(n9184) );
  AND2_X1 U10180 ( .A1(n40939), .A2(n40256), .Z(n57382) );
  NAND2_X1 U10181 ( .A1(n40716), .A2(n41453), .ZN(n41451) );
  NAND2_X1 U10189 ( .A1(n41225), .A2(n12943), .ZN(n9795) );
  NAND2_X1 U10194 ( .A1(n6153), .A2(n40133), .ZN(n40135) );
  INV_X2 U10206 ( .I(n6467), .ZN(n12466) );
  CLKBUF_X2 U10207 ( .I(n18623), .Z(n58047) );
  NAND2_X1 U10208 ( .A1(n2247), .A2(n42266), .ZN(n42271) );
  NAND2_X1 U10216 ( .A1(n13384), .A2(n40364), .ZN(n172) );
  INV_X1 U10220 ( .I(n41066), .ZN(n25817) );
  NOR3_X1 U10221 ( .A1(n11994), .A2(n21207), .A3(n16497), .ZN(n42429) );
  NOR2_X1 U10231 ( .A1(n40204), .A2(n61712), .ZN(n40192) );
  NAND2_X1 U10237 ( .A1(n41890), .A2(n41889), .ZN(n41891) );
  CLKBUF_X2 U10246 ( .I(n25020), .Z(n60567) );
  OAI22_X1 U10258 ( .A1(n57303), .A2(n5709), .B1(n60764), .B2(n9711), .ZN(
        n5708) );
  NAND2_X1 U10271 ( .A1(n42785), .A2(n8538), .ZN(n42787) );
  NOR2_X1 U10273 ( .A1(n41294), .A2(n57545), .ZN(n58097) );
  INV_X1 U10276 ( .I(n12353), .ZN(n18016) );
  INV_X2 U10291 ( .I(n5980), .ZN(n42237) );
  NOR2_X1 U10294 ( .A1(n39948), .A2(n14099), .ZN(n58583) );
  OAI22_X1 U10295 ( .A1(n57773), .A2(n42242), .B1(n449), .B2(n21459), .ZN(
        n21958) );
  AOI22_X1 U10297 ( .A1(n42508), .A2(n42507), .B1(n42509), .B2(n22448), .ZN(
        n42512) );
  NAND2_X1 U10302 ( .A1(n42294), .A2(n9954), .ZN(n42296) );
  OR3_X1 U10308 ( .A1(n40128), .A2(n40092), .A3(n16118), .Z(n39890) );
  INV_X1 U10330 ( .I(n43306), .ZN(n43257) );
  NAND2_X1 U10337 ( .A1(n6262), .A2(n1399), .ZN(n57514) );
  AOI22_X1 U10344 ( .A1(n58097), .A2(n42529), .B1(n42524), .B2(n2586), .ZN(
        n12865) );
  AOI22_X1 U10352 ( .A1(n60219), .A2(n60218), .B1(n40992), .B2(n40991), .ZN(
        n19351) );
  CLKBUF_X2 U10369 ( .I(n43381), .Z(n57651) );
  AOI21_X1 U10383 ( .A1(n17478), .A2(n41062), .B(n41067), .ZN(n17477) );
  INV_X1 U10386 ( .I(n44841), .ZN(n33226) );
  NAND3_X1 U10393 ( .A1(n10652), .A2(n43015), .A3(n43012), .ZN(n10651) );
  NAND3_X1 U10394 ( .A1(n43712), .A2(n6005), .A3(n43992), .ZN(n13208) );
  NAND2_X1 U10407 ( .A1(n42641), .A2(n25210), .ZN(n43197) );
  NAND2_X1 U10416 ( .A1(n42968), .A2(n26020), .ZN(n42412) );
  NOR2_X1 U10430 ( .A1(n43958), .A2(n16890), .ZN(n17266) );
  NAND2_X1 U10431 ( .A1(n60471), .A2(n39829), .ZN(n60470) );
  OAI21_X1 U10432 ( .A1(n22168), .A2(n40410), .B(n40409), .ZN(n6876) );
  NAND2_X1 U10444 ( .A1(n1398), .A2(n8373), .ZN(n61119) );
  NAND2_X1 U10465 ( .A1(n43162), .A2(n43163), .ZN(n61594) );
  NAND2_X1 U10469 ( .A1(n11476), .A2(n22657), .ZN(n42012) );
  NAND2_X1 U10472 ( .A1(n41984), .A2(n41982), .ZN(n12925) );
  NAND2_X1 U10477 ( .A1(n42703), .A2(n2160), .ZN(n40172) );
  NAND2_X1 U10481 ( .A1(n22673), .A2(n8589), .ZN(n43847) );
  NOR2_X1 U10516 ( .A1(n24002), .A2(n41347), .ZN(n17744) );
  NAND2_X1 U10531 ( .A1(n12445), .A2(n12444), .ZN(n60608) );
  NAND3_X1 U10538 ( .A1(n59896), .A2(n3787), .A3(n3782), .ZN(n59149) );
  NOR4_X1 U10539 ( .A1(n42553), .A2(n42555), .A3(n42554), .A4(n20180), .ZN(
        n9563) );
  NOR2_X1 U10542 ( .A1(n43439), .A2(n65179), .ZN(n40016) );
  NOR2_X1 U10543 ( .A1(n42093), .A2(n42094), .ZN(n58222) );
  OAI21_X1 U10583 ( .A1(n42968), .A2(n42072), .B(n42417), .ZN(n13753) );
  NAND2_X1 U10644 ( .A1(n61595), .A2(n61594), .ZN(n61593) );
  NAND2_X1 U10662 ( .A1(n12355), .A2(n5364), .ZN(n41989) );
  NOR2_X1 U10672 ( .A1(n40172), .A2(n42697), .ZN(n41330) );
  NOR2_X1 U10691 ( .A1(n15695), .A2(n23488), .ZN(n43532) );
  OAI21_X1 U10694 ( .A1(n43177), .A2(n43185), .B(n61744), .ZN(n3025) );
  NAND2_X1 U10700 ( .A1(n16921), .A2(n57647), .ZN(n42763) );
  NAND4_X1 U10707 ( .A1(n59833), .A2(n6043), .A3(n42346), .A4(n42344), .ZN(
        n42351) );
  OAI21_X1 U10713 ( .A1(n43427), .A2(n43428), .B(n43426), .ZN(n43432) );
  AND3_X1 U10724 ( .A1(n8653), .A2(n8655), .A3(n8656), .Z(n58831) );
  CLKBUF_X2 U10730 ( .I(n19241), .Z(n57788) );
  OAI21_X1 U10761 ( .A1(n1398), .A2(n57177), .B(n43123), .ZN(n43125) );
  NOR2_X1 U10773 ( .A1(n40171), .A2(n41528), .ZN(n41977) );
  NAND2_X1 U10789 ( .A1(n2735), .A2(n1493), .ZN(n40882) );
  AOI21_X1 U10807 ( .A1(n22519), .A2(n41702), .B(n41706), .ZN(n24648) );
  NAND3_X1 U10809 ( .A1(n58343), .A2(n42392), .A3(n42394), .ZN(n60724) );
  NOR2_X1 U10810 ( .A1(n24130), .A2(n22030), .ZN(n60363) );
  CLKBUF_X2 U10871 ( .I(n24021), .Z(n61142) );
  INV_X1 U10873 ( .I(n46440), .ZN(n14882) );
  INV_X1 U10876 ( .I(n16599), .ZN(n17494) );
  INV_X1 U10887 ( .I(n44994), .ZN(n23270) );
  INV_X2 U10889 ( .I(n10449), .ZN(n13463) );
  CLKBUF_X2 U10910 ( .I(n60606), .Z(n59585) );
  INV_X1 U10919 ( .I(n15698), .ZN(n16557) );
  INV_X1 U10928 ( .I(n45862), .ZN(n58301) );
  INV_X1 U10931 ( .I(n59585), .ZN(n2479) );
  CLKBUF_X2 U10932 ( .I(n10241), .Z(n58750) );
  INV_X1 U10946 ( .I(n1011), .ZN(n58619) );
  INV_X1 U10974 ( .I(n48557), .ZN(n46765) );
  INV_X1 U10990 ( .I(n46906), .ZN(n45775) );
  NOR2_X1 U11000 ( .A1(n47115), .A2(n3686), .ZN(n46809) );
  NAND2_X1 U11007 ( .A1(n46905), .A2(n46906), .ZN(n179) );
  AND2_X1 U11013 ( .A1(n47231), .A2(n19715), .Z(n57298) );
  NOR2_X1 U11015 ( .A1(n59818), .A2(n59670), .ZN(n8271) );
  NAND2_X1 U11019 ( .A1(n23061), .A2(n7931), .ZN(n7930) );
  NOR2_X1 U11024 ( .A1(n47201), .A2(n48208), .ZN(n15295) );
  OAI21_X1 U11027 ( .A1(n48653), .A2(n48659), .B(n48654), .ZN(n48650) );
  AOI22_X1 U11032 ( .A1(n47834), .A2(n62952), .B1(n59695), .B2(n64944), .ZN(
        n2642) );
  CLKBUF_X2 U11033 ( .I(n45643), .Z(n59859) );
  INV_X1 U11053 ( .I(n23934), .ZN(n15162) );
  CLKBUF_X1 U11054 ( .I(n45724), .Z(n4569) );
  NOR2_X1 U11056 ( .A1(n64922), .A2(n12993), .ZN(n12992) );
  NAND2_X1 U11057 ( .A1(n47616), .A2(n47236), .ZN(n47238) );
  INV_X1 U11059 ( .I(n44194), .ZN(n44774) );
  NAND2_X1 U11060 ( .A1(n45673), .A2(n45674), .ZN(n60191) );
  INV_X1 U11061 ( .I(n45554), .ZN(n45976) );
  NAND2_X1 U11070 ( .A1(n4678), .A2(n58705), .ZN(n4262) );
  CLKBUF_X2 U11097 ( .I(n59695), .Z(n61543) );
  OAI22_X1 U11103 ( .A1(n6191), .A2(n8047), .B1(n47806), .B2(n23061), .ZN(n224) );
  NAND2_X1 U11105 ( .A1(n45953), .A2(n45951), .ZN(n19855) );
  NOR2_X1 U11115 ( .A1(n17951), .A2(n45432), .ZN(n47373) );
  NOR2_X1 U11135 ( .A1(n48176), .A2(n48584), .ZN(n48582) );
  AOI21_X1 U11139 ( .A1(n6957), .A2(n20162), .B(n17153), .ZN(n16702) );
  AND2_X1 U11142 ( .A1(n19039), .A2(n48654), .Z(n57243) );
  AOI21_X1 U11143 ( .A1(n47500), .A2(n9907), .B(n47503), .ZN(n12826) );
  NAND2_X1 U11145 ( .A1(n44872), .A2(n63734), .ZN(n58094) );
  INV_X1 U11156 ( .I(n46919), .ZN(n46925) );
  NAND2_X1 U11169 ( .A1(n47218), .A2(n20624), .ZN(n536) );
  NAND3_X1 U11171 ( .A1(n47544), .A2(n48614), .A3(n47174), .ZN(n22704) );
  INV_X2 U11176 ( .I(n45521), .ZN(n46979) );
  INV_X1 U11211 ( .I(n48155), .ZN(n22599) );
  AOI21_X1 U11214 ( .A1(n15566), .A2(n47255), .B(n60191), .ZN(n20787) );
  NAND2_X1 U11216 ( .A1(n24261), .A2(n61628), .ZN(n45945) );
  INV_X1 U11219 ( .I(n2223), .ZN(n47594) );
  AOI21_X1 U11220 ( .A1(n46075), .A2(n4262), .B(n4260), .ZN(n22206) );
  NOR2_X1 U11227 ( .A1(n57530), .A2(n57529), .ZN(n61680) );
  NAND2_X1 U11230 ( .A1(n47027), .A2(n47026), .ZN(n47032) );
  INV_X1 U11234 ( .I(n50268), .ZN(n45920) );
  INV_X1 U11236 ( .I(n48625), .ZN(n48620) );
  NAND3_X1 U11239 ( .A1(n17670), .A2(n13782), .A3(n64447), .ZN(n45903) );
  INV_X1 U11242 ( .I(n47801), .ZN(n47702) );
  INV_X1 U11245 ( .I(n14833), .ZN(n58414) );
  INV_X1 U11249 ( .I(n2786), .ZN(n12114) );
  NAND2_X1 U11255 ( .A1(n48198), .A2(n48197), .ZN(n58043) );
  NAND2_X1 U11260 ( .A1(n47376), .A2(n23718), .ZN(n25346) );
  NAND2_X1 U11267 ( .A1(n45541), .A2(n61017), .ZN(n61331) );
  AOI21_X1 U11290 ( .A1(n47509), .A2(n47508), .B(n57550), .ZN(n47522) );
  NAND2_X1 U11320 ( .A1(n50428), .A2(n23063), .ZN(n45466) );
  INV_X1 U11325 ( .I(n3472), .ZN(n2904) );
  INV_X1 U11328 ( .I(n47976), .ZN(n49775) );
  AOI22_X1 U11333 ( .A1(n46942), .A2(n18127), .B1(n46941), .B2(n60038), .ZN(
        n47981) );
  CLKBUF_X2 U11351 ( .I(n49493), .Z(n12701) );
  NAND2_X1 U11362 ( .A1(n48979), .A2(n62975), .ZN(n17514) );
  NOR2_X1 U11366 ( .A1(n60467), .A2(n50330), .ZN(n17901) );
  NOR2_X1 U11368 ( .A1(n45916), .A2(n50267), .ZN(n60066) );
  OAI21_X1 U11369 ( .A1(n44001), .A2(n47798), .B(n1657), .ZN(n44002) );
  NAND2_X1 U11371 ( .A1(n49610), .A2(n49319), .ZN(n49313) );
  NAND2_X1 U11376 ( .A1(n17335), .A2(n15724), .ZN(n49301) );
  OAI21_X1 U11380 ( .A1(n25555), .A2(n50398), .B(n50074), .ZN(n58123) );
  NAND2_X1 U11400 ( .A1(n3093), .A2(n3094), .ZN(n61209) );
  INV_X1 U11404 ( .I(n14617), .ZN(n50295) );
  INV_X1 U11409 ( .I(n7288), .ZN(n48791) );
  NOR2_X1 U11413 ( .A1(n12536), .A2(n8729), .ZN(n61210) );
  NAND2_X1 U11424 ( .A1(n50269), .A2(n50268), .ZN(n50270) );
  CLKBUF_X4 U11435 ( .I(n50045), .Z(n3335) );
  NOR2_X1 U11456 ( .A1(n48780), .A2(n49377), .ZN(n59639) );
  CLKBUF_X1 U11459 ( .I(n37713), .Z(n30564) );
  INV_X1 U11470 ( .I(n39210), .ZN(n58078) );
  INV_X1 U11486 ( .I(n52232), .ZN(n13830) );
  NOR2_X1 U11490 ( .A1(n50290), .A2(n50289), .ZN(n61392) );
  NAND2_X1 U11519 ( .A1(n5661), .A2(n48819), .ZN(n12840) );
  NAND2_X1 U11522 ( .A1(n58123), .A2(n59200), .ZN(n46725) );
  NAND2_X1 U11528 ( .A1(n50023), .A2(n47759), .ZN(n60695) );
  NOR2_X1 U11536 ( .A1(n50345), .A2(n21870), .ZN(n50351) );
  INV_X1 U11551 ( .I(n49476), .ZN(n48269) );
  NOR2_X1 U11552 ( .A1(n2810), .A2(n48067), .ZN(n46973) );
  NAND2_X1 U11560 ( .A1(n50295), .A2(n62035), .ZN(n61050) );
  INV_X1 U11569 ( .I(n56143), .ZN(n60828) );
  INV_X1 U11572 ( .I(n49257), .ZN(n3151) );
  NAND2_X1 U11575 ( .A1(n58844), .A2(n24802), .ZN(n14203) );
  NAND2_X1 U11580 ( .A1(n49847), .A2(n59101), .ZN(n59100) );
  NAND2_X1 U11582 ( .A1(n50048), .A2(n49572), .ZN(n22308) );
  NAND2_X1 U11601 ( .A1(n49421), .A2(n50397), .ZN(n59733) );
  CLKBUF_X2 U11614 ( .I(n49817), .Z(n721) );
  INV_X1 U11634 ( .I(n49798), .ZN(n58885) );
  OAI22_X1 U11640 ( .A1(n50364), .A2(n49133), .B1(n49201), .B2(n49132), .ZN(
        n49134) );
  NAND3_X1 U11641 ( .A1(n48853), .A2(n4724), .A3(n19175), .ZN(n48857) );
  OAI21_X1 U11670 ( .A1(n49365), .A2(n47642), .B(n49681), .ZN(n47645) );
  NOR2_X1 U11705 ( .A1(n61721), .A2(n19510), .ZN(n6214) );
  NAND3_X1 U11711 ( .A1(n49247), .A2(n49248), .A3(n61235), .ZN(n49252) );
  INV_X1 U11713 ( .I(n50611), .ZN(n50523) );
  OAI21_X1 U11731 ( .A1(n3032), .A2(n50383), .B(n50382), .ZN(n50384) );
  CLKBUF_X1 U11734 ( .I(n51940), .Z(n22614) );
  NAND2_X1 U11749 ( .A1(n49062), .A2(n49833), .ZN(n60732) );
  OAI21_X1 U11752 ( .A1(n3699), .A2(n47971), .B(n48825), .ZN(n3698) );
  NOR2_X1 U11754 ( .A1(n48018), .A2(n23612), .ZN(n49553) );
  INV_X2 U11769 ( .I(n1466), .ZN(n52538) );
  CLKBUF_X2 U11770 ( .I(n22153), .Z(n22152) );
  INV_X1 U11780 ( .I(n52601), .ZN(n58184) );
  INV_X1 U11794 ( .I(n51749), .ZN(n22141) );
  INV_X1 U11798 ( .I(n51036), .ZN(n51042) );
  INV_X1 U11801 ( .I(n51786), .ZN(n4350) );
  CLKBUF_X4 U11809 ( .I(n52445), .Z(n22795) );
  INV_X1 U11810 ( .I(n52541), .ZN(n1461) );
  INV_X1 U11816 ( .I(n58819), .ZN(n1462) );
  INV_X1 U11828 ( .I(n60934), .ZN(n59952) );
  CLKBUF_X2 U11829 ( .I(n51763), .Z(n61571) );
  CLKBUF_X2 U11839 ( .I(n25968), .Z(n5878) );
  INV_X1 U11841 ( .I(n24053), .ZN(n60395) );
  INV_X1 U11844 ( .I(n51737), .ZN(n58629) );
  INV_X1 U11849 ( .I(n51298), .ZN(n50167) );
  NAND2_X1 U11855 ( .A1(n15498), .A2(n59951), .ZN(n59950) );
  INV_X1 U11880 ( .I(n52349), .ZN(n59039) );
  CLKBUF_X2 U11891 ( .I(n12681), .Z(n60642) );
  OR2_X1 U11895 ( .A1(n53848), .A2(n64832), .Z(n57317) );
  CLKBUF_X1 U11899 ( .I(n1287), .Z(n58225) );
  INV_X1 U11906 ( .I(n54055), .ZN(n1599) );
  NAND2_X1 U11912 ( .A1(n56627), .A2(n63038), .ZN(n51453) );
  NOR2_X1 U11918 ( .A1(n1603), .A2(n55690), .ZN(n55694) );
  CLKBUF_X2 U11937 ( .I(n53847), .Z(n4473) );
  INV_X1 U11938 ( .I(n54062), .ZN(n16797) );
  CLKBUF_X2 U11955 ( .I(n11207), .Z(n59970) );
  NOR2_X1 U11990 ( .A1(n57390), .A2(n10237), .ZN(n60335) );
  CLKBUF_X2 U12012 ( .I(n8121), .Z(n22977) );
  NAND2_X1 U12043 ( .A1(n54105), .A2(n2959), .ZN(n49930) );
  INV_X1 U12052 ( .I(n57067), .ZN(n52255) );
  INV_X2 U12073 ( .I(n13312), .ZN(n15804) );
  NAND3_X1 U12082 ( .A1(n8062), .A2(n52945), .A3(n63194), .ZN(n8061) );
  NAND2_X1 U12086 ( .A1(n52901), .A2(n55245), .ZN(n55419) );
  AOI21_X1 U12095 ( .A1(n24647), .A2(n13920), .B(n56600), .ZN(n56981) );
  AOI21_X1 U12100 ( .A1(n53548), .A2(n51710), .B(n54105), .ZN(n51715) );
  CLKBUF_X2 U12122 ( .I(n54823), .Z(n61463) );
  NAND2_X1 U12129 ( .A1(n56252), .A2(n57203), .ZN(n57693) );
  INV_X1 U12132 ( .I(n52779), .ZN(n61559) );
  CLKBUF_X4 U12149 ( .I(n54323), .Z(n23736) );
  INV_X2 U12184 ( .I(n56414), .ZN(n9388) );
  INV_X1 U12186 ( .I(n56619), .ZN(n21069) );
  NOR2_X1 U12189 ( .A1(n60336), .A2(n60335), .ZN(n60334) );
  CLKBUF_X1 U12190 ( .I(n55906), .Z(n58655) );
  AOI21_X1 U12197 ( .A1(n21070), .A2(n56623), .B(n21069), .ZN(n58060) );
  INV_X2 U12200 ( .I(n54102), .ZN(n12917) );
  NAND3_X1 U12207 ( .A1(n55928), .A2(n60373), .A3(n57361), .ZN(n55930) );
  AOI21_X1 U12210 ( .A1(n54311), .A2(n54310), .B(n26154), .ZN(n26153) );
  AOI21_X1 U12211 ( .A1(n25461), .A2(n53606), .B(n25067), .ZN(n447) );
  OAI21_X1 U12222 ( .A1(n57185), .A2(n58418), .B(n55906), .ZN(n55919) );
  NOR2_X1 U12224 ( .A1(n53407), .A2(n54039), .ZN(n60042) );
  NAND2_X1 U12226 ( .A1(n53897), .A2(n53896), .ZN(n59929) );
  OAI21_X1 U12235 ( .A1(n56548), .A2(n56547), .B(n21643), .ZN(n56549) );
  INV_X1 U12248 ( .I(n52295), .ZN(n59609) );
  NOR2_X1 U12253 ( .A1(n25022), .A2(n14708), .ZN(n61567) );
  NAND2_X1 U12258 ( .A1(n56817), .A2(n56803), .ZN(n56747) );
  NAND2_X1 U12288 ( .A1(n55821), .A2(n20447), .ZN(n55772) );
  NAND2_X1 U12289 ( .A1(n60563), .A2(n60564), .ZN(n58796) );
  NAND2_X1 U12300 ( .A1(n14708), .A2(n56961), .ZN(n13693) );
  NAND2_X1 U12304 ( .A1(n55565), .A2(n55575), .ZN(n55586) );
  INV_X1 U12317 ( .I(n55135), .ZN(n26094) );
  NAND2_X1 U12318 ( .A1(n53690), .A2(n23935), .ZN(n53664) );
  NOR2_X1 U12319 ( .A1(n54162), .A2(n54192), .ZN(n54135) );
  OAI21_X1 U12330 ( .A1(n13693), .A2(n56964), .B(n6902), .ZN(n10218) );
  CLKBUF_X2 U12331 ( .I(n58811), .Z(n21) );
  INV_X1 U12346 ( .I(n55886), .ZN(n19077) );
  NAND3_X1 U12348 ( .A1(n12915), .A2(n25344), .A3(n23292), .ZN(n53994) );
  NOR2_X1 U12353 ( .A1(n55166), .A2(n55108), .ZN(n55112) );
  INV_X1 U12362 ( .I(n1919), .ZN(n57997) );
  AOI21_X1 U12369 ( .A1(n53694), .A2(n53650), .B(n53658), .ZN(n53651) );
  NAND2_X1 U12371 ( .A1(n23956), .A2(n19735), .ZN(n53264) );
  AOI22_X1 U12381 ( .A1(n54665), .A2(n54664), .B1(n54700), .B2(n22122), .ZN(
        n54674) );
  CLKBUF_X4 U12385 ( .I(Key[10]), .Z(n53174) );
  NOR2_X1 U12390 ( .A1(n56513), .A2(n56514), .ZN(n59779) );
  OAI21_X1 U12394 ( .A1(n3507), .A2(n53167), .B(n2820), .ZN(n59260) );
  NAND2_X1 U12398 ( .A1(n53647), .A2(n53648), .ZN(n10021) );
  CLKBUF_X4 U12404 ( .I(Key[28]), .Z(n23929) );
  AND2_X1 U12405 ( .A1(n56809), .A2(n56796), .Z(n57212) );
  AND3_X1 U12409 ( .A1(n13296), .A2(n46773), .A3(n48576), .Z(n57213) );
  OR2_X1 U12411 ( .A1(n29192), .A2(n59883), .Z(n57214) );
  AND4_X1 U12426 ( .A1(n28563), .A2(n29088), .A3(n30340), .A4(n13361), .Z(
        n57216) );
  AND2_X1 U12433 ( .A1(n19432), .A2(n19431), .Z(n57217) );
  XOR2_X1 U12438 ( .A1(n32324), .A2(n18434), .Z(n57218) );
  AND2_X1 U12442 ( .A1(n31845), .A2(n6125), .Z(n57220) );
  XNOR2_X1 U12448 ( .A1(n50926), .A2(n39685), .ZN(n57221) );
  OR2_X1 U12449 ( .A1(n54202), .A2(n54203), .Z(n57222) );
  XNOR2_X1 U12468 ( .A1(n43683), .A2(n52199), .ZN(n57223) );
  AND3_X1 U12472 ( .A1(n1324), .A2(n55910), .A3(n59792), .Z(n57225) );
  XNOR2_X1 U12473 ( .A1(n51548), .A2(n24132), .ZN(n57226) );
  XNOR2_X1 U12475 ( .A1(n44390), .A2(n31477), .ZN(n57227) );
  AND3_X1 U12487 ( .A1(n12310), .A2(n51713), .A3(n53879), .Z(n57228) );
  XNOR2_X1 U12488 ( .A1(n52162), .A2(n52161), .ZN(n57229) );
  XNOR2_X1 U12500 ( .A1(n46251), .A2(n43618), .ZN(n57230) );
  XNOR2_X1 U12501 ( .A1(n46666), .A2(n14806), .ZN(n57232) );
  AND2_X1 U12505 ( .A1(n5569), .A2(n58283), .Z(n57236) );
  XNOR2_X1 U12508 ( .A1(n37823), .A2(n37819), .ZN(n57237) );
  XNOR2_X1 U12510 ( .A1(n46215), .A2(n45884), .ZN(n57240) );
  AND2_X1 U12522 ( .A1(n54115), .A2(n54113), .Z(n57247) );
  XNOR2_X1 U12523 ( .A1(n1680), .A2(n62136), .ZN(n57250) );
  NAND2_X1 U12525 ( .A1(n41983), .A2(n40885), .ZN(n57251) );
  AND3_X1 U12533 ( .A1(n10170), .A2(n29549), .A3(n29548), .Z(n57253) );
  AND2_X1 U12535 ( .A1(n54111), .A2(n9124), .Z(n57254) );
  AND3_X1 U12542 ( .A1(n55089), .A2(n674), .A3(n15520), .Z(n57260) );
  AND2_X1 U12548 ( .A1(n21903), .A2(n60135), .Z(n57263) );
  AND2_X1 U12549 ( .A1(n55324), .A2(n55441), .Z(n57264) );
  AND2_X1 U12550 ( .A1(n36775), .A2(n20060), .Z(n57266) );
  AND2_X1 U12553 ( .A1(n34164), .A2(n34168), .Z(n57268) );
  XNOR2_X1 U12554 ( .A1(n52187), .A2(n52186), .ZN(n57269) );
  AND4_X1 U12557 ( .A1(n22934), .A2(n31269), .A3(n23269), .A4(n31271), .Z(
        n57271) );
  XNOR2_X1 U12559 ( .A1(n33238), .A2(n1314), .ZN(n57272) );
  AND2_X1 U12561 ( .A1(n33019), .A2(n35690), .Z(n57273) );
  XNOR2_X1 U12564 ( .A1(n1419), .A2(n7705), .ZN(n57275) );
  XNOR2_X1 U12566 ( .A1(n45044), .A2(n14251), .ZN(n57276) );
  OR2_X1 U12575 ( .A1(n60510), .A2(n17379), .Z(n57277) );
  AND2_X1 U12582 ( .A1(n34218), .A2(n32945), .Z(n57279) );
  AND3_X2 U12600 ( .A1(n43173), .A2(n61744), .A3(n61442), .Z(n57281) );
  XNOR2_X1 U12604 ( .A1(n18922), .A2(n31772), .ZN(n57285) );
  INV_X1 U12613 ( .I(n3117), .ZN(n2902) );
  AND3_X1 U12616 ( .A1(n54641), .A2(n17935), .A3(n20740), .Z(n57287) );
  NAND3_X1 U12623 ( .A1(n1477), .A2(n21639), .A3(n21638), .ZN(n57288) );
  AND3_X1 U12626 ( .A1(n49225), .A2(n22526), .A3(n49224), .Z(n57290) );
  AND2_X1 U12631 ( .A1(n2524), .A2(n55295), .Z(n57291) );
  XNOR2_X1 U12632 ( .A1(n24062), .A2(n60918), .ZN(n57292) );
  OR2_X1 U12637 ( .A1(n55298), .A2(n55685), .Z(n57293) );
  AND2_X1 U12647 ( .A1(n34383), .A2(n35279), .Z(n57294) );
  OR2_X1 U12651 ( .A1(n49929), .A2(n6130), .Z(n57297) );
  AND2_X1 U12655 ( .A1(n17267), .A2(n17266), .Z(n57299) );
  OR2_X2 U12662 ( .A1(n20209), .A2(n60368), .Z(n57300) );
  XNOR2_X1 U12669 ( .A1(n44523), .A2(n10370), .ZN(n57301) );
  NOR2_X1 U12674 ( .A1(n48847), .A2(n49525), .ZN(n57302) );
  INV_X1 U12681 ( .I(n59225), .ZN(n41102) );
  XNOR2_X1 U12698 ( .A1(n23120), .A2(n957), .ZN(n57311) );
  INV_X1 U12717 ( .I(n837), .ZN(n28066) );
  AND3_X2 U12719 ( .A1(n17387), .A2(n17385), .A3(n34494), .Z(n57313) );
  XNOR2_X1 U12721 ( .A1(n8449), .A2(n37547), .ZN(n57314) );
  CLKBUF_X2 U12726 ( .I(n61202), .Z(n60962) );
  OR2_X1 U12731 ( .A1(n12423), .A2(n26612), .Z(n57318) );
  NAND2_X1 U12732 ( .A1(n54073), .A2(n60794), .ZN(n57319) );
  AND4_X1 U12733 ( .A1(n61627), .A2(n1591), .A3(n58755), .A4(n59180), .Z(
        n57320) );
  XNOR2_X1 U12734 ( .A1(n15676), .A2(n1823), .ZN(n57321) );
  XNOR2_X1 U12736 ( .A1(n30604), .A2(n32475), .ZN(n57323) );
  XNOR2_X1 U12742 ( .A1(n32476), .A2(n32475), .ZN(n57324) );
  INV_X2 U12749 ( .I(n26823), .ZN(n27839) );
  XNOR2_X1 U12757 ( .A1(n22334), .A2(n14818), .ZN(n57326) );
  AND2_X2 U12761 ( .A1(n40320), .A2(n13984), .Z(n57327) );
  AND3_X1 U12763 ( .A1(n29009), .A2(n8584), .A3(n61007), .Z(n57329) );
  XNOR2_X1 U12768 ( .A1(n39776), .A2(n39775), .ZN(n57331) );
  XNOR2_X1 U12772 ( .A1(n52369), .A2(n52368), .ZN(n57336) );
  NAND2_X1 U12774 ( .A1(n34277), .A2(n61108), .ZN(n57338) );
  AND3_X1 U12779 ( .A1(n35936), .A2(n58220), .A3(n35517), .Z(n57339) );
  NOR2_X1 U12783 ( .A1(n40221), .A2(n1737), .ZN(n57340) );
  OR2_X2 U12800 ( .A1(n42084), .A2(n42404), .Z(n57341) );
  AND2_X1 U12819 ( .A1(n42282), .A2(n42281), .Z(n57345) );
  OR2_X1 U12824 ( .A1(n48434), .A2(n47947), .Z(n57346) );
  CLKBUF_X8 U12828 ( .I(n22898), .Z(n1708) );
  OR3_X1 U12832 ( .A1(n54200), .A2(n9968), .A3(n54205), .Z(n57348) );
  AND3_X1 U12857 ( .A1(n50431), .A2(n50429), .A3(n50430), .Z(n57349) );
  AND3_X1 U12858 ( .A1(n314), .A2(n11045), .A3(n11046), .Z(n57350) );
  XNOR2_X1 U12861 ( .A1(n52527), .A2(n52526), .ZN(n57351) );
  XNOR2_X1 U12864 ( .A1(n39753), .A2(n49122), .ZN(n57352) );
  INV_X1 U12894 ( .I(n15715), .ZN(n1441) );
  OR2_X1 U12896 ( .A1(n6635), .A2(n54848), .Z(n57354) );
  AND3_X1 U12901 ( .A1(n22172), .A2(n22171), .A3(n61959), .Z(n57355) );
  XNOR2_X1 U12923 ( .A1(n25608), .A2(n7070), .ZN(n57356) );
  AND2_X1 U12925 ( .A1(n48057), .A2(n49848), .Z(n57357) );
  CLKBUF_X4 U12934 ( .I(n26489), .Z(n19452) );
  CLKBUF_X1 U12936 ( .I(n31138), .Z(n7461) );
  XNOR2_X1 U12947 ( .A1(n31753), .A2(n29974), .ZN(n57358) );
  XNOR2_X1 U12949 ( .A1(n5630), .A2(n44220), .ZN(n57359) );
  XNOR2_X1 U12952 ( .A1(n14855), .A2(n44880), .ZN(n57360) );
  AND3_X2 U12953 ( .A1(n28241), .A2(n28065), .A3(n28066), .Z(n57363) );
  AND2_X1 U12959 ( .A1(n33634), .A2(n24093), .Z(n57364) );
  XNOR2_X1 U12963 ( .A1(n32199), .A2(n31651), .ZN(n57365) );
  AND2_X1 U12968 ( .A1(n376), .A2(n24374), .Z(n57366) );
  AND2_X1 U12970 ( .A1(n15761), .A2(n18629), .Z(n57367) );
  OR2_X1 U12978 ( .A1(n54277), .A2(n14354), .Z(n57370) );
  XNOR2_X1 U12980 ( .A1(n58341), .A2(n50773), .ZN(n57371) );
  NAND2_X1 U12987 ( .A1(n19208), .A2(n54069), .ZN(n57372) );
  XNOR2_X1 U12988 ( .A1(n46229), .A2(n46132), .ZN(n57373) );
  OR2_X2 U12991 ( .A1(n35658), .A2(n35646), .Z(n57375) );
  XNOR2_X1 U13001 ( .A1(n24018), .A2(n38260), .ZN(n57376) );
  AND2_X1 U13003 ( .A1(n60989), .A2(n60988), .Z(n57377) );
  XNOR2_X1 U13004 ( .A1(n21094), .A2(n16309), .ZN(n57378) );
  XOR2_X1 U13010 ( .A1(n51799), .A2(n14870), .Z(n57379) );
  XNOR2_X1 U13032 ( .A1(n42816), .A2(n42815), .ZN(n57380) );
  OR2_X2 U13035 ( .A1(n52393), .A2(n52389), .Z(n57383) );
  AND2_X2 U13040 ( .A1(n21343), .A2(n26143), .Z(n57390) );
  AND2_X1 U13045 ( .A1(n16689), .A2(n22072), .Z(n57393) );
  XNOR2_X1 U13052 ( .A1(n46204), .A2(n46203), .ZN(n57394) );
  AND3_X2 U13053 ( .A1(n28170), .A2(n19223), .A3(n28169), .Z(n57395) );
  INV_X1 U13063 ( .I(n11197), .ZN(n43373) );
  OR2_X1 U13065 ( .A1(n60043), .A2(n60042), .Z(n57396) );
  OR2_X1 U13131 ( .A1(n56264), .A2(n14324), .Z(n57401) );
  AND2_X1 U13133 ( .A1(n40938), .A2(n40939), .Z(n57402) );
  INV_X1 U13139 ( .I(n58369), .ZN(n39110) );
  XNOR2_X1 U13141 ( .A1(n12774), .A2(n21826), .ZN(n57403) );
  OR2_X2 U13145 ( .A1(n54949), .A2(n26095), .Z(n57404) );
  INV_X1 U13152 ( .I(n35314), .ZN(n35754) );
  INV_X1 U13161 ( .I(n35534), .ZN(n36090) );
  INV_X1 U13170 ( .I(n46326), .ZN(n57525) );
  INV_X1 U13199 ( .I(n25866), .ZN(n46835) );
  INV_X1 U13203 ( .I(n15551), .ZN(n33518) );
  OR2_X2 U13218 ( .A1(n23352), .A2(n14439), .Z(n57412) );
  AND2_X2 U13223 ( .A1(n14919), .A2(n24301), .Z(n57414) );
  AND2_X1 U13229 ( .A1(n20360), .A2(n34458), .Z(n57416) );
  INV_X1 U13238 ( .I(n24172), .ZN(n31142) );
  INV_X1 U13239 ( .I(n6276), .ZN(n59376) );
  XNOR2_X1 U13251 ( .A1(n38156), .A2(n48387), .ZN(n57420) );
  INV_X2 U13255 ( .I(n21064), .ZN(n22044) );
  OR2_X2 U13264 ( .A1(n33729), .A2(n3669), .Z(n57423) );
  AND2_X1 U13285 ( .A1(n3869), .A2(n3868), .Z(n57427) );
  CLKBUF_X8 U13286 ( .I(n21492), .Z(n22713) );
  INV_X1 U13287 ( .I(n60690), .ZN(n41883) );
  INV_X1 U13306 ( .I(n27626), .ZN(n9475) );
  INV_X1 U13312 ( .I(n35980), .ZN(n19354) );
  CLKBUF_X1 U13320 ( .I(n50406), .Z(n7494) );
  OR2_X1 U13322 ( .A1(n40872), .A2(n42394), .Z(n57431) );
  XNOR2_X1 U13323 ( .A1(n5712), .A2(n44604), .ZN(n57432) );
  INV_X1 U13324 ( .I(n52223), .ZN(n55628) );
  CLKBUF_X4 U13350 ( .I(n37681), .Z(n14228) );
  XNOR2_X1 U13352 ( .A1(n31327), .A2(n31326), .ZN(n57435) );
  INV_X2 U13372 ( .I(n9558), .ZN(n56585) );
  INV_X2 U13377 ( .I(n56585), .ZN(n56245) );
  AND2_X2 U13398 ( .A1(n19624), .A2(n31097), .Z(n57437) );
  XOR2_X1 U13399 ( .A1(n32666), .A2(n31154), .Z(n57438) );
  XNOR2_X1 U13401 ( .A1(n38332), .A2(n38331), .ZN(n57439) );
  XNOR2_X1 U13402 ( .A1(n24414), .A2(n31766), .ZN(n57440) );
  XNOR2_X1 U13414 ( .A1(n32645), .A2(n32646), .ZN(n57441) );
  OR2_X1 U13418 ( .A1(n30704), .A2(n23056), .Z(n57442) );
  INV_X1 U13431 ( .I(n23781), .ZN(n1430) );
  XNOR2_X1 U13445 ( .A1(n4339), .A2(n4340), .ZN(n57445) );
  AND2_X1 U13447 ( .A1(n8373), .A2(n65217), .Z(n57446) );
  XNOR2_X1 U13459 ( .A1(n38777), .A2(n4525), .ZN(n57448) );
  CLKBUF_X2 U13468 ( .I(n24378), .Z(n17400) );
  XOR2_X1 U13469 ( .A1(n37980), .A2(n37302), .Z(n57450) );
  INV_X1 U13475 ( .I(n25292), .ZN(n12409) );
  AND3_X1 U13484 ( .A1(n35352), .A2(n35548), .A3(n35964), .Z(n57453) );
  XNOR2_X1 U13492 ( .A1(n17889), .A2(n17888), .ZN(n57455) );
  AND2_X1 U13494 ( .A1(n46328), .A2(n10487), .Z(n57456) );
  CLKBUF_X1 U13502 ( .I(n34606), .Z(n20946) );
  CLKBUF_X4 U13505 ( .I(n46269), .Z(n3449) );
  XOR2_X1 U13525 ( .A1(n19803), .A2(n59895), .Z(n57458) );
  OR2_X1 U13526 ( .A1(n57837), .A2(n61511), .Z(n57459) );
  AND2_X1 U13533 ( .A1(n42260), .A2(n59271), .Z(n57461) );
  OR2_X2 U13549 ( .A1(n15215), .A2(n19770), .Z(n57462) );
  INV_X1 U13559 ( .I(n48130), .ZN(n24545) );
  AND2_X1 U13574 ( .A1(n45803), .A2(n11693), .Z(n57466) );
  CLKBUF_X4 U13577 ( .I(n48728), .Z(n6130) );
  INV_X1 U13587 ( .I(n22947), .ZN(n55262) );
  OR2_X2 U13596 ( .A1(n13485), .A2(n26143), .Z(n57470) );
  CLKBUF_X2 U13603 ( .I(n148), .Z(n10748) );
  CLKBUF_X2 U13625 ( .I(n51214), .Z(n19202) );
  AND2_X1 U13636 ( .A1(n52717), .A2(n52716), .Z(n57476) );
  BUF_X4 U13641 ( .I(n56644), .Z(n56731) );
  INV_X4 U13642 ( .I(n56731), .ZN(n56703) );
  INV_X1 U13685 ( .I(n52007), .ZN(n52131) );
  NOR3_X2 U13689 ( .A1(n15452), .A2(n15450), .A3(n61943), .ZN(n37107) );
  XOR2_X1 U13693 ( .A1(n18644), .A2(n57477), .Z(n57747) );
  XOR2_X1 U13697 ( .A1(n4265), .A2(n23422), .Z(n57477) );
  AOI22_X1 U13721 ( .A1(n27256), .A2(n1320), .B1(n8628), .B2(n597), .ZN(n26745) );
  XOR2_X1 U13735 ( .A1(n46526), .A2(n16050), .Z(n13545) );
  NAND2_X2 U13747 ( .A1(n1272), .A2(n984), .ZN(n14965) );
  INV_X2 U13750 ( .I(n57480), .ZN(n984) );
  NOR2_X2 U13751 ( .A1(n40595), .A2(n41078), .ZN(n57480) );
  XOR2_X1 U13762 ( .A1(n3402), .A2(n57379), .Z(n57481) );
  XOR2_X1 U13775 ( .A1(n3894), .A2(n57482), .Z(n60366) );
  XOR2_X1 U13776 ( .A1(n13069), .A2(n5898), .Z(n57482) );
  INV_X2 U13793 ( .I(n18951), .ZN(n59670) );
  NAND3_X2 U13794 ( .A1(n58354), .A2(n30866), .A3(n30867), .ZN(n33863) );
  XOR2_X1 U13796 ( .A1(n57486), .A2(n57485), .Z(n4038) );
  XOR2_X1 U13797 ( .A1(n25483), .A2(n531), .Z(n57485) );
  INV_X2 U13820 ( .I(n11340), .ZN(n23812) );
  AND2_X1 U13825 ( .A1(n44344), .A2(n44343), .Z(n57488) );
  XOR2_X1 U13833 ( .A1(n44307), .A2(n57292), .Z(n57489) );
  NOR2_X2 U13835 ( .A1(n10124), .A2(n26428), .ZN(n26429) );
  NOR3_X2 U13838 ( .A1(n14402), .A2(n14400), .A3(n48036), .ZN(n15473) );
  NOR2_X2 U13852 ( .A1(n16722), .A2(n16720), .ZN(n16719) );
  XOR2_X1 U13856 ( .A1(n10393), .A2(n46510), .Z(n57490) );
  NAND2_X1 U13874 ( .A1(n4019), .A2(n46089), .ZN(n4018) );
  INV_X1 U13880 ( .I(n58823), .ZN(n59637) );
  XOR2_X1 U13885 ( .A1(n12524), .A2(n11113), .Z(n10677) );
  NAND2_X2 U13891 ( .A1(n16645), .A2(n16644), .ZN(n14761) );
  BUF_X2 U13906 ( .I(n25188), .Z(n57492) );
  NAND2_X2 U13931 ( .A1(n57494), .A2(n2561), .ZN(n9337) );
  NAND2_X2 U13940 ( .A1(n21561), .A2(n57000), .ZN(n57495) );
  OAI21_X2 U13959 ( .A1(n22799), .A2(n21263), .B(n30197), .ZN(n57496) );
  OR2_X1 U13963 ( .A1(n9281), .A2(n30076), .Z(n7735) );
  OAI21_X2 U13978 ( .A1(n57497), .A2(n34988), .B(n34986), .ZN(n58790) );
  NOR2_X1 U13988 ( .A1(n58697), .A2(n63421), .ZN(n57497) );
  NAND4_X2 U13994 ( .A1(n57219), .A2(n20966), .A3(n29020), .A4(n57499), .ZN(
        n11360) );
  NAND2_X2 U14006 ( .A1(n42259), .A2(n42267), .ZN(n5319) );
  OAI22_X1 U14017 ( .A1(n8896), .A2(n49811), .B1(n8895), .B2(n4109), .ZN(
        n57501) );
  NAND2_X2 U14025 ( .A1(n57502), .A2(n27035), .ZN(n13174) );
  NOR2_X2 U14030 ( .A1(n58214), .A2(n58215), .ZN(n57502) );
  XOR2_X1 U14055 ( .A1(n25348), .A2(n12501), .Z(n45865) );
  XOR2_X1 U14063 ( .A1(n33292), .A2(n33293), .Z(n25891) );
  XOR2_X1 U14081 ( .A1(n32206), .A2(n23143), .Z(n33292) );
  XOR2_X1 U14082 ( .A1(n5245), .A2(n11446), .Z(n58838) );
  NOR3_X1 U14083 ( .A1(n6983), .A2(n6982), .A3(n4881), .ZN(n6981) );
  OR2_X2 U14100 ( .A1(n58823), .A2(n16657), .Z(n40571) );
  NOR2_X2 U14102 ( .A1(n35816), .A2(n10232), .ZN(n22797) );
  NAND2_X2 U14109 ( .A1(n24097), .A2(n15533), .ZN(n29254) );
  NOR2_X2 U14132 ( .A1(n54860), .A2(n54640), .ZN(n7148) );
  NAND2_X2 U14148 ( .A1(n34816), .A2(n35938), .ZN(n3767) );
  XOR2_X1 U14163 ( .A1(n21513), .A2(n12392), .Z(n57507) );
  NAND2_X1 U14196 ( .A1(n27741), .A2(n27740), .ZN(n60408) );
  AND2_X1 U14219 ( .A1(n18398), .A2(n62353), .Z(n43374) );
  AND2_X1 U14222 ( .A1(n4320), .A2(n33628), .Z(n33624) );
  OAI21_X1 U14243 ( .A1(n60103), .A2(n60102), .B(n55721), .ZN(n9867) );
  XOR2_X1 U14253 ( .A1(n57510), .A2(n21412), .Z(n20449) );
  XOR2_X1 U14326 ( .A1(n57517), .A2(n5810), .Z(n11102) );
  XOR2_X1 U14330 ( .A1(n5809), .A2(n45400), .Z(n57517) );
  OAI22_X1 U14344 ( .A1(n53881), .A2(n54015), .B1(n9613), .B2(n54349), .ZN(
        n53038) );
  AND2_X2 U14352 ( .A1(n2766), .A2(n47467), .Z(n47473) );
  NAND4_X2 U14355 ( .A1(n57519), .A2(n49336), .A3(n49334), .A4(n13788), .ZN(
        n51810) );
  AND2_X1 U14356 ( .A1(n10454), .A2(n49335), .Z(n57519) );
  NOR2_X2 U14374 ( .A1(n1419), .A2(n1792), .ZN(n36226) );
  NAND2_X1 U14403 ( .A1(n43250), .A2(n9440), .ZN(n57521) );
  INV_X1 U14417 ( .I(n760), .ZN(n57522) );
  NAND2_X1 U14425 ( .A1(n28972), .A2(n57679), .ZN(n28973) );
  XOR2_X1 U14440 ( .A1(n5520), .A2(n57523), .Z(n3776) );
  XOR2_X1 U14442 ( .A1(n2328), .A2(n2327), .Z(n57523) );
  OAI22_X1 U14467 ( .A1(n45450), .A2(n47730), .B1(n46731), .B2(n63647), .ZN(
        n43751) );
  INV_X2 U14471 ( .I(n47728), .ZN(n45450) );
  NAND2_X2 U14472 ( .A1(n46731), .A2(n47748), .ZN(n47728) );
  NAND2_X2 U14512 ( .A1(n61744), .A2(n43513), .ZN(n46331) );
  NAND2_X1 U14519 ( .A1(n15693), .A2(n49393), .ZN(n18950) );
  AOI21_X1 U14529 ( .A1(n37926), .A2(n6276), .B(n40470), .ZN(n60213) );
  NOR2_X2 U14531 ( .A1(n18538), .A2(n22295), .ZN(n33782) );
  NAND2_X2 U14533 ( .A1(n65160), .A2(n35130), .ZN(n22295) );
  NAND2_X1 U14536 ( .A1(n8800), .A2(n34747), .ZN(n34750) );
  NOR2_X2 U14543 ( .A1(n59275), .A2(n57456), .ZN(n46520) );
  NOR2_X2 U14544 ( .A1(n21467), .A2(n1310), .ZN(n59809) );
  INV_X2 U14578 ( .I(n55738), .ZN(n55473) );
  NAND2_X2 U14580 ( .A1(n23941), .A2(n22499), .ZN(n55738) );
  OR2_X1 U14583 ( .A1(n8336), .A2(n9281), .Z(n30075) );
  NAND3_X2 U14588 ( .A1(n35867), .A2(n35868), .A3(n35866), .ZN(n38433) );
  NAND3_X2 U14593 ( .A1(n24482), .A2(n53034), .A3(n53039), .ZN(n6743) );
  NAND3_X2 U14603 ( .A1(n5043), .A2(n11757), .A3(n11756), .ZN(n23495) );
  NAND2_X2 U14610 ( .A1(n42868), .A2(n16850), .ZN(n10827) );
  OAI21_X1 U14615 ( .A1(n28731), .A2(n29842), .B(n29845), .ZN(n28732) );
  NAND3_X2 U14643 ( .A1(n5208), .A2(n5209), .A3(n5210), .ZN(n14108) );
  NAND3_X1 U14647 ( .A1(n56780), .A2(n56779), .A3(n56806), .ZN(n56781) );
  NOR2_X2 U14652 ( .A1(n58753), .A2(n58754), .ZN(n8994) );
  NOR2_X1 U14655 ( .A1(n22900), .A2(n12692), .ZN(n57538) );
  NAND2_X1 U14658 ( .A1(n45648), .A2(n45645), .ZN(n58529) );
  NOR2_X2 U14681 ( .A1(n22505), .A2(n7760), .ZN(n28518) );
  BUF_X2 U14692 ( .I(n1209), .Z(n57543) );
  INV_X2 U14702 ( .I(n42527), .ZN(n57545) );
  XOR2_X1 U14705 ( .A1(n38222), .A2(n25914), .Z(n16795) );
  XOR2_X1 U14706 ( .A1(n16796), .A2(n15371), .Z(n38222) );
  OR2_X1 U14715 ( .A1(n57547), .A2(n26940), .Z(n10222) );
  NOR2_X1 U14716 ( .A1(n58708), .A2(n26937), .ZN(n57547) );
  OR3_X1 U14721 ( .A1(n28243), .A2(n27380), .A3(n28240), .Z(n57613) );
  NOR2_X1 U14729 ( .A1(n1865), .A2(n13174), .ZN(n29877) );
  NOR2_X1 U14739 ( .A1(n30285), .A2(n23772), .ZN(n29039) );
  OAI21_X1 U14750 ( .A1(n16485), .A2(n57549), .B(n16470), .ZN(n27722) );
  NOR2_X1 U14751 ( .A1(n27710), .A2(n27852), .ZN(n57549) );
  INV_X2 U14753 ( .I(n20139), .ZN(n46813) );
  XOR2_X1 U14755 ( .A1(n2948), .A2(n10700), .Z(n20139) );
  OAI22_X1 U14756 ( .A1(n47504), .A2(n1064), .B1(n47506), .B2(n47505), .ZN(
        n57550) );
  XOR2_X1 U14758 ( .A1(n24274), .A2(n16476), .Z(n38620) );
  NOR2_X2 U14778 ( .A1(n35898), .A2(n35886), .ZN(n13297) );
  NOR4_X2 U14807 ( .A1(n52695), .A2(n57555), .A3(n19732), .A4(n470), .ZN(
        n20485) );
  XOR2_X1 U14822 ( .A1(n24058), .A2(n1200), .Z(n8038) );
  INV_X2 U14843 ( .I(n24431), .ZN(n1569) );
  NAND2_X2 U14846 ( .A1(n7760), .A2(n9556), .ZN(n24431) );
  NAND2_X1 U14852 ( .A1(n2958), .A2(n9830), .ZN(n37190) );
  NAND2_X1 U14856 ( .A1(n40196), .A2(n19148), .ZN(n40189) );
  OR2_X2 U14865 ( .A1(n12287), .A2(n13799), .Z(n3057) );
  XOR2_X1 U14894 ( .A1(n19226), .A2(n46557), .Z(n21307) );
  AOI22_X2 U14909 ( .A1(n58398), .A2(n56987), .B1(n51446), .B2(n51445), .ZN(
        n51447) );
  XOR2_X1 U14929 ( .A1(n33264), .A2(n17920), .Z(n18167) );
  XOR2_X1 U14932 ( .A1(n57563), .A2(n16209), .Z(n24631) );
  AOI22_X2 U14967 ( .A1(n22211), .A2(n24647), .B1(n7835), .B2(n61405), .ZN(
        n56982) );
  INV_X2 U14970 ( .I(n53537), .ZN(n21982) );
  XOR2_X1 U14991 ( .A1(n57564), .A2(n55087), .Z(Plaintext[94]) );
  NAND3_X1 U14995 ( .A1(n60524), .A2(n55085), .A3(n55086), .ZN(n57564) );
  NAND2_X2 U15011 ( .A1(n55567), .A2(n55568), .ZN(n8949) );
  BUF_X2 U15012 ( .I(n54793), .Z(n24075) );
  AND2_X1 U15015 ( .A1(n842), .A2(n57566), .Z(n8088) );
  NAND2_X1 U15046 ( .A1(n3243), .A2(n2731), .ZN(n58759) );
  BUF_X2 U15055 ( .I(n50426), .Z(n57572) );
  NAND3_X2 U15056 ( .A1(n57350), .A2(n57958), .A3(n15670), .ZN(n42651) );
  NOR2_X1 U15091 ( .A1(n56052), .A2(n61865), .ZN(n56055) );
  INV_X2 U15112 ( .I(n57580), .ZN(n28542) );
  XNOR2_X1 U15117 ( .A1(Ciphertext[97]), .A2(Key[188]), .ZN(n57580) );
  NAND2_X2 U15122 ( .A1(n25191), .A2(n52444), .ZN(n9553) );
  NOR2_X2 U15123 ( .A1(n47453), .A2(n25193), .ZN(n52444) );
  OAI22_X2 U15125 ( .A1(n43093), .A2(n4659), .B1(n43092), .B2(n58874), .ZN(
        n14510) );
  NOR3_X2 U15134 ( .A1(n57582), .A2(n30963), .A3(n30964), .ZN(n25329) );
  AOI21_X1 U15160 ( .A1(n13766), .A2(n30537), .B(n58747), .ZN(n29980) );
  XOR2_X1 U15182 ( .A1(n59694), .A2(n57586), .Z(n44800) );
  INV_X2 U15185 ( .I(n42091), .ZN(n57586) );
  OAI22_X1 U15196 ( .A1(n27529), .A2(n23362), .B1(n27203), .B2(n20929), .ZN(
        n26352) );
  XOR2_X1 U15208 ( .A1(n57587), .A2(n23983), .Z(n18031) );
  XOR2_X1 U15209 ( .A1(n38314), .A2(n23493), .Z(n57587) );
  XOR2_X1 U15214 ( .A1(n32301), .A2(n31327), .Z(n18571) );
  NOR3_X2 U15215 ( .A1(n31376), .A2(n31378), .A3(n31377), .ZN(n32301) );
  NOR2_X2 U15228 ( .A1(n59429), .A2(n57589), .ZN(n1990) );
  BUF_X2 U15230 ( .I(n61261), .Z(n57590) );
  XOR2_X1 U15242 ( .A1(n24383), .A2(n2355), .Z(n39396) );
  NAND2_X2 U15250 ( .A1(n57593), .A2(n32827), .ZN(n20571) );
  NAND2_X1 U15266 ( .A1(n2004), .A2(n19078), .ZN(n59574) );
  XOR2_X1 U15272 ( .A1(n38159), .A2(n9896), .Z(n22561) );
  XOR2_X1 U15276 ( .A1(n33288), .A2(n33287), .Z(n59431) );
  XOR2_X1 U15293 ( .A1(n57595), .A2(n32353), .Z(n58238) );
  XOR2_X1 U15296 ( .A1(n32377), .A2(n24258), .Z(n57595) );
  AOI21_X1 U15299 ( .A1(n27653), .A2(n5268), .B(n59994), .ZN(n27654) );
  OAI21_X2 U15305 ( .A1(n29583), .A2(n64867), .B(n57596), .ZN(n29584) );
  NOR2_X2 U15309 ( .A1(n59330), .A2(n21814), .ZN(n57596) );
  NAND2_X1 U15315 ( .A1(n57597), .A2(n59703), .ZN(n8321) );
  NAND2_X1 U15317 ( .A1(n41678), .A2(n41677), .ZN(n57597) );
  XOR2_X1 U15320 ( .A1(n1819), .A2(n57598), .Z(n6590) );
  XOR2_X1 U15326 ( .A1(n14345), .A2(n31321), .Z(n4696) );
  NOR2_X2 U15332 ( .A1(n21305), .A2(n21304), .ZN(n48104) );
  AND2_X1 U15333 ( .A1(n22840), .A2(n57600), .Z(n918) );
  NAND2_X2 U15334 ( .A1(n24179), .A2(n43288), .ZN(n42423) );
  NAND2_X1 U15335 ( .A1(n24230), .A2(n24229), .ZN(n54158) );
  OR2_X1 U15340 ( .A1(n36226), .A2(n57171), .Z(n35599) );
  AOI22_X1 U15347 ( .A1(n29229), .A2(n29228), .B1(n57605), .B2(n29227), .ZN(
        n29230) );
  NAND3_X1 U15349 ( .A1(n29225), .A2(n30276), .A3(n30285), .ZN(n57605) );
  XOR2_X1 U15350 ( .A1(n19956), .A2(n57606), .Z(n58957) );
  NOR3_X2 U15397 ( .A1(n20947), .A2(n57611), .A3(n21151), .ZN(n24813) );
  NOR2_X1 U15398 ( .A1(n57613), .A2(n57612), .ZN(n57611) );
  XOR2_X1 U15411 ( .A1(n39638), .A2(n38913), .Z(n38919) );
  XOR2_X1 U15413 ( .A1(n11534), .A2(n38912), .Z(n39638) );
  NAND3_X2 U15415 ( .A1(n30483), .A2(n30493), .A3(n30484), .ZN(n15193) );
  OR2_X2 U15420 ( .A1(n61735), .A2(n59272), .Z(n34623) );
  AOI22_X2 U15444 ( .A1(n14043), .A2(n14044), .B1(n11059), .B2(n2148), .ZN(
        n17326) );
  AOI21_X1 U15500 ( .A1(n4907), .A2(n27415), .B(n27414), .ZN(n27418) );
  XOR2_X1 U15513 ( .A1(n31977), .A2(n25402), .Z(n32028) );
  XOR2_X1 U15527 ( .A1(n23070), .A2(n20234), .Z(n38649) );
  XOR2_X1 U15531 ( .A1(n21734), .A2(n38395), .Z(n57623) );
  OAI22_X2 U15532 ( .A1(n8853), .A2(n40190), .B1(n40189), .B2(n58599), .ZN(
        n57624) );
  INV_X2 U15537 ( .I(n36401), .ZN(n35361) );
  NAND3_X1 U15582 ( .A1(n36049), .A2(n36773), .A3(n36050), .ZN(n36051) );
  NAND2_X2 U15587 ( .A1(n11656), .A2(n12164), .ZN(n30048) );
  NOR2_X2 U15591 ( .A1(n37428), .A2(n23801), .ZN(n36916) );
  AND2_X1 U15601 ( .A1(n46103), .A2(n48653), .Z(n57626) );
  BUF_X2 U15622 ( .I(n732), .Z(n57628) );
  AOI22_X1 U15624 ( .A1(n29107), .A2(n29106), .B1(n2276), .B2(n10404), .ZN(
        n5484) );
  NAND2_X2 U15634 ( .A1(n5045), .A2(n57629), .ZN(n4198) );
  NAND3_X2 U15657 ( .A1(n48585), .A2(n48482), .A3(n178), .ZN(n48480) );
  NOR2_X2 U15666 ( .A1(n22184), .A2(n36123), .ZN(n57631) );
  XOR2_X1 U15676 ( .A1(n44734), .A2(n44732), .Z(n5576) );
  XOR2_X1 U15678 ( .A1(n12234), .A2(n12232), .Z(n44732) );
  OAI22_X1 U15689 ( .A1(n48995), .A2(n48994), .B1(n49318), .B2(n48996), .ZN(
        n24710) );
  NOR3_X2 U15691 ( .A1(n48699), .A2(n57640), .A3(n57639), .ZN(n49237) );
  NAND4_X2 U15700 ( .A1(n39945), .A2(n40833), .A3(n60693), .A4(n23420), .ZN(
        n39515) );
  NAND3_X1 U15708 ( .A1(n56238), .A2(n12468), .A3(n57239), .ZN(n56244) );
  NOR2_X1 U15722 ( .A1(n30188), .A2(n30189), .ZN(n58248) );
  NOR2_X1 U15730 ( .A1(n48783), .A2(n49545), .ZN(n48784) );
  AOI21_X2 U15733 ( .A1(n32429), .A2(n34775), .B(n64276), .ZN(n16679) );
  OR2_X1 U15758 ( .A1(n42756), .A2(n577), .Z(n57647) );
  OR2_X1 U15759 ( .A1(n26002), .A2(n57648), .Z(n59259) );
  XOR2_X1 U15770 ( .A1(n38213), .A2(n38205), .Z(n57649) );
  INV_X2 U15775 ( .I(n19569), .ZN(n1086) );
  NAND2_X2 U15777 ( .A1(n3271), .A2(n47518), .ZN(n19569) );
  OAI21_X2 U15783 ( .A1(n21178), .A2(n57195), .B(n58934), .ZN(n47194) );
  INV_X1 U15786 ( .I(n27256), .ZN(n57652) );
  XOR2_X1 U15801 ( .A1(n59465), .A2(n6357), .Z(n6157) );
  INV_X1 U15808 ( .I(n42451), .ZN(n41312) );
  AOI22_X1 U15820 ( .A1(n10481), .A2(n4918), .B1(n58262), .B2(n57655), .ZN(
        n3455) );
  NAND3_X2 U15825 ( .A1(n41318), .A2(n41319), .A3(n22016), .ZN(n61071) );
  NAND4_X2 U15828 ( .A1(n42296), .A2(n61930), .A3(n42298), .A4(n42295), .ZN(
        n42308) );
  NOR2_X1 U15829 ( .A1(n51714), .A2(n51715), .ZN(n12650) );
  NAND3_X2 U15830 ( .A1(n19682), .A2(n19686), .A3(n47355), .ZN(n22098) );
  XOR2_X1 U15832 ( .A1(n57657), .A2(n54289), .Z(Plaintext[65]) );
  NOR2_X2 U15860 ( .A1(n48625), .A2(n47541), .ZN(n48218) );
  XOR2_X1 U15883 ( .A1(n10595), .A2(n50993), .Z(n57660) );
  NAND3_X1 U15884 ( .A1(n40733), .A2(n39025), .A3(n20555), .ZN(n2090) );
  NAND2_X2 U15918 ( .A1(n57748), .A2(n57264), .ZN(n55385) );
  OR2_X2 U15964 ( .A1(n21899), .A2(n60937), .Z(n30832) );
  XOR2_X1 U15977 ( .A1(n22103), .A2(n21900), .Z(n60937) );
  XOR2_X1 U16010 ( .A1(n3214), .A2(n57664), .Z(n2407) );
  XOR2_X1 U16012 ( .A1(n22033), .A2(n22035), .Z(n57664) );
  XOR2_X1 U16037 ( .A1(n61947), .A2(n6458), .Z(n7432) );
  XOR2_X1 U16041 ( .A1(n37724), .A2(n8449), .Z(n6458) );
  XOR2_X1 U16065 ( .A1(n52006), .A2(n52005), .Z(n57665) );
  XOR2_X1 U16086 ( .A1(n37549), .A2(n14010), .Z(n11005) );
  INV_X2 U16099 ( .I(n18441), .ZN(n11016) );
  NAND2_X2 U16105 ( .A1(n60693), .A2(n41132), .ZN(n18441) );
  XOR2_X1 U16133 ( .A1(n32676), .A2(n57667), .Z(n26220) );
  XOR2_X1 U16139 ( .A1(n32675), .A2(n32674), .Z(n57667) );
  NAND2_X1 U16157 ( .A1(n57668), .A2(n17740), .ZN(n27824) );
  NAND3_X1 U16162 ( .A1(n17743), .A2(n28621), .A3(n20743), .ZN(n57668) );
  INV_X4 U16201 ( .I(n7979), .ZN(n60030) );
  XOR2_X1 U16204 ( .A1(n30835), .A2(n30834), .Z(n30837) );
  XOR2_X1 U16205 ( .A1(n51677), .A2(n61681), .Z(n25854) );
  OR2_X2 U16252 ( .A1(n60513), .A2(n60587), .Z(n60602) );
  OAI21_X2 U16315 ( .A1(n36041), .A2(n34819), .B(n35583), .ZN(n25242) );
  NAND2_X2 U16330 ( .A1(n52933), .A2(n22592), .ZN(n55480) );
  NAND2_X1 U16333 ( .A1(n57674), .A2(n57673), .ZN(n57672) );
  NAND2_X1 U16336 ( .A1(n55466), .A2(n55465), .ZN(n57674) );
  XOR2_X1 U16341 ( .A1(n55637), .A2(n55638), .Z(Plaintext[124]) );
  INV_X2 U16354 ( .I(n57678), .ZN(n29303) );
  OAI22_X1 U16366 ( .A1(n9039), .A2(n9169), .B1(n6033), .B2(n19435), .ZN(
        n57680) );
  NAND2_X2 U16367 ( .A1(n13931), .A2(n57681), .ZN(n50045) );
  AOI21_X2 U16372 ( .A1(n12618), .A2(n13178), .B(n13177), .ZN(n57681) );
  XOR2_X1 U16382 ( .A1(n57683), .A2(n60699), .Z(n13592) );
  XOR2_X1 U16387 ( .A1(n9010), .A2(n11801), .Z(n57683) );
  NAND2_X2 U16402 ( .A1(n10866), .A2(n16403), .ZN(n19570) );
  NAND2_X2 U16407 ( .A1(n5472), .A2(n1816), .ZN(n10866) );
  XOR2_X1 U16420 ( .A1(n11574), .A2(n17599), .Z(n17944) );
  XOR2_X1 U16425 ( .A1(n5435), .A2(n12022), .Z(n32099) );
  XOR2_X1 U16427 ( .A1(n14218), .A2(n57687), .Z(n58338) );
  XOR2_X1 U16442 ( .A1(n25402), .A2(n11663), .Z(n57687) );
  XOR2_X1 U16447 ( .A1(n11456), .A2(n57688), .Z(n12480) );
  XOR2_X1 U16448 ( .A1(n32285), .A2(n11455), .Z(n57688) );
  NAND2_X2 U16451 ( .A1(n57689), .A2(n59083), .ZN(n43979) );
  AOI22_X2 U16452 ( .A1(n33094), .A2(n8780), .B1(n33096), .B2(n33095), .ZN(
        n33108) );
  XOR2_X1 U16453 ( .A1(n58717), .A2(n57690), .Z(n15801) );
  XOR2_X1 U16457 ( .A1(n57984), .A2(n57324), .Z(n57690) );
  BUF_X2 U16464 ( .I(n56585), .Z(n57691) );
  NOR2_X2 U16465 ( .A1(n56261), .A2(n57692), .ZN(n56344) );
  NAND2_X1 U16467 ( .A1(n56251), .A2(n56250), .ZN(n57694) );
  NOR2_X2 U16469 ( .A1(n48546), .A2(n48544), .ZN(n47096) );
  XOR2_X1 U16473 ( .A1(n14608), .A2(n14607), .Z(n61132) );
  OAI21_X2 U16474 ( .A1(n57236), .A2(n57695), .B(n57235), .ZN(n60761) );
  XOR2_X1 U16493 ( .A1(n23674), .A2(n1466), .Z(n6140) );
  INV_X2 U16494 ( .I(n57697), .ZN(n25594) );
  XOR2_X1 U16495 ( .A1(n46224), .A2(n44594), .Z(n57697) );
  BUF_X4 U16497 ( .I(n26217), .Z(n60543) );
  INV_X2 U16528 ( .I(n54036), .ZN(n57700) );
  INV_X2 U16533 ( .I(n57701), .ZN(n17156) );
  NAND3_X2 U16565 ( .A1(n58572), .A2(n42361), .A3(n41614), .ZN(n4197) );
  XOR2_X1 U16568 ( .A1(n25845), .A2(n21260), .Z(n57704) );
  OR2_X2 U16572 ( .A1(n61354), .A2(n57901), .Z(n58514) );
  NAND2_X2 U16576 ( .A1(n15215), .A2(n3246), .ZN(n40729) );
  XOR2_X1 U16578 ( .A1(n3889), .A2(n57706), .Z(n54062) );
  XOR2_X1 U16581 ( .A1(n411), .A2(n51821), .Z(n57706) );
  OR2_X1 U16584 ( .A1(n14007), .A2(n49013), .Z(n5636) );
  OR2_X2 U16606 ( .A1(n16938), .A2(n25298), .Z(n3942) );
  XNOR2_X1 U16607 ( .A1(n49241), .A2(n49240), .ZN(n58661) );
  NOR2_X1 U16618 ( .A1(n576), .A2(n23626), .ZN(n34462) );
  XOR2_X1 U16636 ( .A1(n52530), .A2(n12509), .Z(n52156) );
  XOR2_X1 U16669 ( .A1(n46347), .A2(n44769), .Z(n57708) );
  XOR2_X1 U16684 ( .A1(n45111), .A2(n44990), .Z(n106) );
  NAND2_X2 U16715 ( .A1(n57709), .A2(n59184), .ZN(n11070) );
  NAND3_X2 U16716 ( .A1(n20569), .A2(n33396), .A3(n33395), .ZN(n33401) );
  AND2_X1 U16727 ( .A1(n22559), .A2(n19231), .Z(n9042) );
  XOR2_X1 U16745 ( .A1(n39589), .A2(n59023), .Z(n8209) );
  XOR2_X1 U16749 ( .A1(n25984), .A2(n21429), .Z(n39589) );
  NOR2_X2 U16752 ( .A1(n28886), .A2(n27508), .ZN(n29356) );
  OR2_X1 U16784 ( .A1(n22169), .A2(n59261), .Z(n36125) );
  XNOR2_X1 U16793 ( .A1(n19878), .A2(n32205), .ZN(n58137) );
  NAND2_X2 U16798 ( .A1(n23650), .A2(n5283), .ZN(n49619) );
  NOR2_X2 U16803 ( .A1(n21445), .A2(n62880), .ZN(n48151) );
  NOR2_X1 U16809 ( .A1(n5280), .A2(n5773), .ZN(n9564) );
  XOR2_X1 U16823 ( .A1(n38319), .A2(n38318), .Z(n38320) );
  NAND2_X2 U16849 ( .A1(n33570), .A2(n33096), .ZN(n33350) );
  XOR2_X1 U16875 ( .A1(n49962), .A2(n52187), .Z(n57714) );
  NAND2_X2 U16896 ( .A1(n58564), .A2(n7645), .ZN(n41997) );
  NAND4_X2 U16912 ( .A1(n63697), .A2(n36837), .A3(n26213), .A4(n36852), .ZN(
        n57716) );
  NOR2_X2 U16919 ( .A1(n21364), .A2(n54088), .ZN(n54589) );
  OR2_X1 U16923 ( .A1(n13669), .A2(n41412), .Z(n40742) );
  AND3_X1 U16924 ( .A1(n28345), .A2(n28344), .A3(n28343), .Z(n13056) );
  NOR2_X2 U16938 ( .A1(n2995), .A2(n43572), .ZN(n2898) );
  AND2_X1 U16945 ( .A1(n53374), .A2(n1448), .Z(n1179) );
  NAND2_X2 U16947 ( .A1(n12667), .A2(n53361), .ZN(n53374) );
  NAND2_X2 U16970 ( .A1(n6219), .A2(n6218), .ZN(n11556) );
  NOR2_X2 U16972 ( .A1(n37203), .A2(n57719), .ZN(n9201) );
  NAND2_X1 U16980 ( .A1(n55815), .A2(n55816), .ZN(n12432) );
  NAND2_X2 U16988 ( .A1(n57720), .A2(n55476), .ZN(n55724) );
  NOR3_X2 U17018 ( .A1(n57722), .A2(n30427), .A3(n57721), .ZN(n30434) );
  NOR2_X1 U17020 ( .A1(n30423), .A2(n60064), .ZN(n57722) );
  XOR2_X1 U17022 ( .A1(n23853), .A2(n9873), .Z(n17284) );
  OAI22_X1 U17033 ( .A1(n49016), .A2(n49017), .B1(n49018), .B2(n14007), .ZN(
        n57723) );
  BUF_X2 U17047 ( .I(n49226), .Z(n10030) );
  XOR2_X1 U17053 ( .A1(n51618), .A2(n21616), .Z(n51620) );
  INV_X2 U17083 ( .I(n24529), .ZN(n24063) );
  XOR2_X1 U17095 ( .A1(n57727), .A2(n5749), .Z(n32571) );
  XOR2_X1 U17100 ( .A1(n7948), .A2(n31849), .Z(n57727) );
  XOR2_X1 U17104 ( .A1(n1929), .A2(n8342), .Z(n8596) );
  AND2_X1 U17108 ( .A1(n58563), .A2(n34691), .Z(n7299) );
  INV_X2 U17109 ( .I(n2255), .ZN(n58164) );
  NAND2_X2 U17115 ( .A1(n1391), .A2(n5398), .ZN(n2255) );
  NAND3_X1 U17126 ( .A1(n41009), .A2(n58851), .A3(n23355), .ZN(n58340) );
  OAI22_X1 U17138 ( .A1(n3467), .A2(n21906), .B1(n1813), .B2(n60054), .ZN(
        n34688) );
  NAND2_X2 U17140 ( .A1(n2891), .A2(n25251), .ZN(n21906) );
  NOR2_X2 U17158 ( .A1(n54221), .A2(n23731), .ZN(n54225) );
  NAND2_X1 U17159 ( .A1(n33294), .A2(n22909), .ZN(n57729) );
  XOR2_X1 U17173 ( .A1(n24828), .A2(n57272), .Z(n57730) );
  INV_X2 U17180 ( .I(n24825), .ZN(n59546) );
  BUF_X4 U17215 ( .I(n59634), .Z(n59409) );
  NOR2_X2 U17235 ( .A1(n61047), .A2(n21529), .ZN(n41918) );
  NOR2_X2 U17280 ( .A1(n1256), .A2(n54259), .ZN(n54276) );
  NOR2_X2 U17295 ( .A1(n47415), .A2(n45267), .ZN(n47688) );
  OR2_X1 U17298 ( .A1(n35224), .A2(n35835), .Z(n35844) );
  NOR2_X2 U17319 ( .A1(n29716), .A2(n57746), .ZN(n31276) );
  NAND3_X2 U17320 ( .A1(n20401), .A2(n20088), .A3(n20089), .ZN(n57746) );
  NOR3_X2 U17328 ( .A1(n30861), .A2(n30859), .A3(n30860), .ZN(n58354) );
  XOR2_X1 U17332 ( .A1(n7533), .A2(n57747), .Z(n59763) );
  AND3_X1 U17334 ( .A1(n31273), .A2(n8182), .A3(n31268), .Z(n59735) );
  XOR2_X1 U17335 ( .A1(n38656), .A2(n38204), .Z(n38205) );
  XOR2_X1 U17336 ( .A1(n25326), .A2(n5555), .Z(n38656) );
  NOR3_X2 U17339 ( .A1(n61286), .A2(n55315), .A3(n55326), .ZN(n57748) );
  NAND2_X2 U17366 ( .A1(n21454), .A2(n11542), .ZN(n36443) );
  NOR2_X1 U17378 ( .A1(n57749), .A2(n14784), .ZN(n4870) );
  NOR2_X1 U17389 ( .A1(n14789), .A2(n12546), .ZN(n57749) );
  NAND3_X2 U17395 ( .A1(n26204), .A2(n57751), .A3(n26205), .ZN(n41549) );
  NAND2_X2 U17406 ( .A1(n14555), .A2(n3896), .ZN(n57752) );
  AND2_X1 U17438 ( .A1(n47339), .A2(n47338), .Z(n57754) );
  NOR2_X2 U17458 ( .A1(n1715), .A2(n6426), .ZN(n42650) );
  AND2_X2 U17473 ( .A1(n3482), .A2(n12049), .Z(n20860) );
  NAND2_X2 U17480 ( .A1(n19331), .A2(n18473), .ZN(n58307) );
  AOI22_X1 U17490 ( .A1(n3435), .A2(n65183), .B1(n65111), .B2(n27392), .ZN(
        n3434) );
  NAND2_X2 U17498 ( .A1(n14019), .A2(n28448), .ZN(n6273) );
  XOR2_X1 U17500 ( .A1(n44883), .A2(n44881), .Z(n57759) );
  XOR2_X1 U17524 ( .A1(n15289), .A2(n57760), .Z(n58294) );
  NAND2_X1 U17526 ( .A1(n23231), .A2(n12120), .ZN(n15286) );
  OR2_X1 U17527 ( .A1(n3510), .A2(n19329), .Z(n12203) );
  NOR2_X2 U17538 ( .A1(n48644), .A2(n26226), .ZN(n57762) );
  XOR2_X1 U17570 ( .A1(n52545), .A2(n4915), .Z(n12086) );
  XOR2_X1 U17582 ( .A1(n12088), .A2(n12087), .Z(n52545) );
  NAND3_X2 U17611 ( .A1(n58920), .A2(n50124), .A3(n11449), .ZN(n52616) );
  XOR2_X1 U17626 ( .A1(n43807), .A2(n44120), .Z(n45053) );
  OAI21_X1 U17637 ( .A1(n57766), .A2(n4176), .B(n47096), .ZN(n21821) );
  OAI21_X2 U17646 ( .A1(n1779), .A2(n35567), .B(n9721), .ZN(n35880) );
  NAND2_X2 U17649 ( .A1(n22632), .A2(n6682), .ZN(n34378) );
  NAND2_X2 U17653 ( .A1(n8305), .A2(n61198), .ZN(n43351) );
  AND2_X1 U17677 ( .A1(n28595), .A2(n29643), .Z(n28147) );
  XOR2_X1 U17678 ( .A1(n57775), .A2(n16274), .Z(n5119) );
  XOR2_X1 U17680 ( .A1(n51738), .A2(n58629), .Z(n57775) );
  XOR2_X1 U17681 ( .A1(n57776), .A2(n30959), .Z(n7417) );
  XOR2_X1 U17683 ( .A1(n27008), .A2(n27007), .Z(n57776) );
  OR2_X1 U17687 ( .A1(n62045), .A2(n2974), .Z(n8029) );
  XOR2_X1 U17691 ( .A1(n57777), .A2(n1129), .Z(n6641) );
  XOR2_X1 U17694 ( .A1(n58184), .A2(n52523), .Z(n57777) );
  NAND3_X1 U17696 ( .A1(n42003), .A2(n43011), .A3(n42004), .ZN(n57778) );
  INV_X2 U17744 ( .I(n20270), .ZN(n1519) );
  NAND3_X2 U17757 ( .A1(n61242), .A2(n61241), .A3(n45927), .ZN(n57780) );
  AOI21_X2 U17773 ( .A1(n10088), .A2(n45224), .B(n16597), .ZN(n16596) );
  BUF_X2 U17780 ( .I(n29661), .Z(n57781) );
  NOR2_X1 U17798 ( .A1(n57783), .A2(n57447), .ZN(n57782) );
  NOR2_X1 U17799 ( .A1(n41787), .A2(n41789), .ZN(n57783) );
  XOR2_X1 U17804 ( .A1(n57784), .A2(n18562), .Z(n7308) );
  XOR2_X1 U17810 ( .A1(n5878), .A2(n61606), .Z(n57784) );
  NAND2_X1 U17824 ( .A1(n59044), .A2(n59107), .ZN(n7355) );
  XOR2_X1 U17844 ( .A1(n60918), .A2(n57380), .Z(n831) );
  XOR2_X1 U17845 ( .A1(n57786), .A2(n21825), .Z(n21824) );
  XOR2_X1 U17846 ( .A1(n31965), .A2(n31964), .Z(n57786) );
  BUF_X2 U17859 ( .I(n19830), .Z(n57790) );
  INV_X2 U17863 ( .I(n57792), .ZN(n15763) );
  NAND2_X2 U17866 ( .A1(n7651), .A2(n22498), .ZN(n57792) );
  NOR2_X1 U17884 ( .A1(n10003), .A2(n43422), .ZN(n43424) );
  BUF_X2 U17907 ( .I(n23163), .Z(n19999) );
  NAND2_X2 U17963 ( .A1(n4547), .A2(n43572), .ZN(n42341) );
  XOR2_X1 U17974 ( .A1(n64269), .A2(n32305), .Z(n656) );
  OAI22_X2 U17995 ( .A1(n27388), .A2(n26272), .B1(n26271), .B2(n22095), .ZN(
        n26273) );
  NAND2_X2 U18006 ( .A1(n37206), .A2(n4388), .ZN(n37217) );
  NOR2_X2 U18007 ( .A1(n54860), .A2(n1373), .ZN(n7800) );
  NAND3_X1 U18028 ( .A1(n57799), .A2(n19523), .A3(n3738), .ZN(n24694) );
  NOR2_X1 U18033 ( .A1(n49922), .A2(n49921), .ZN(n57799) );
  NAND2_X1 U18063 ( .A1(n60943), .A2(n60942), .ZN(n37194) );
  XOR2_X1 U18080 ( .A1(n51990), .A2(n3842), .Z(n58947) );
  XOR2_X1 U18086 ( .A1(n19228), .A2(n51942), .Z(n3842) );
  NAND4_X2 U18088 ( .A1(n3360), .A2(n57802), .A3(n3357), .A4(n3468), .ZN(
        n16539) );
  AOI21_X2 U18091 ( .A1(n48243), .A2(n209), .B(n58548), .ZN(n57802) );
  NAND2_X1 U18099 ( .A1(n21272), .A2(n55594), .ZN(n55547) );
  XOR2_X1 U18101 ( .A1(n57803), .A2(n55516), .Z(Plaintext[114]) );
  NAND3_X1 U18115 ( .A1(n55515), .A2(n55513), .A3(n55514), .ZN(n57803) );
  NAND2_X1 U18131 ( .A1(n55504), .A2(n55590), .ZN(n55505) );
  NAND3_X2 U18159 ( .A1(n11224), .A2(n11222), .A3(n41551), .ZN(n41697) );
  XOR2_X1 U18163 ( .A1(n15081), .A2(n39258), .Z(n57809) );
  NOR2_X1 U18167 ( .A1(n38683), .A2(n38686), .ZN(n60272) );
  INV_X2 U18169 ( .I(n62535), .ZN(n57810) );
  AND2_X2 U18179 ( .A1(n7439), .A2(n6845), .Z(n41059) );
  XOR2_X1 U18186 ( .A1(n5676), .A2(n9157), .Z(n5607) );
  XOR2_X1 U18198 ( .A1(n58027), .A2(n45333), .Z(n42955) );
  XOR2_X1 U18207 ( .A1(n19759), .A2(n17284), .Z(n19066) );
  NOR3_X2 U18209 ( .A1(n57819), .A2(n14622), .A3(n5509), .ZN(n5510) );
  NOR2_X1 U18216 ( .A1(n40576), .A2(n40581), .ZN(n57819) );
  AND2_X1 U18219 ( .A1(n45546), .A2(n17793), .Z(n57821) );
  NAND2_X1 U18220 ( .A1(n1775), .A2(n948), .ZN(n11054) );
  AND2_X1 U18221 ( .A1(n24836), .A2(n28318), .Z(n28052) );
  XOR2_X1 U18222 ( .A1(n57822), .A2(n3431), .Z(n8782) );
  XOR2_X1 U18225 ( .A1(n18248), .A2(n9787), .Z(n57822) );
  XOR2_X1 U18233 ( .A1(Ciphertext[39]), .A2(Key[166]), .Z(n28317) );
  AOI22_X1 U18255 ( .A1(n57824), .A2(n23934), .B1(n47141), .B2(n47380), .ZN(
        n45433) );
  NAND2_X1 U18259 ( .A1(n45414), .A2(n1072), .ZN(n57824) );
  OR2_X1 U18272 ( .A1(n33391), .A2(n157), .Z(n32821) );
  NOR2_X2 U18285 ( .A1(n57826), .A2(n9584), .ZN(n30441) );
  NAND4_X2 U18287 ( .A1(n27267), .A2(n27265), .A3(n23000), .A4(n27266), .ZN(
        n57826) );
  INV_X2 U18290 ( .I(n50054), .ZN(n50142) );
  NAND2_X1 U18300 ( .A1(n57829), .A2(n57828), .ZN(n33415) );
  NAND2_X1 U18301 ( .A1(n33414), .A2(n57830), .ZN(n57829) );
  NOR2_X1 U18305 ( .A1(n43531), .A2(n15695), .ZN(n43493) );
  XOR2_X1 U18307 ( .A1(n13069), .A2(n18133), .Z(n7420) );
  AND2_X1 U18309 ( .A1(n19638), .A2(n42477), .Z(n40346) );
  OR2_X1 U18324 ( .A1(n17192), .A2(n35394), .Z(n57831) );
  NAND4_X2 U18470 ( .A1(n59488), .A2(n39033), .A3(n39032), .A4(n39034), .ZN(
        n39035) );
  NAND3_X1 U18492 ( .A1(n22657), .A2(n8676), .A3(n42993), .ZN(n43091) );
  NOR2_X1 U18511 ( .A1(n1444), .A2(n27976), .ZN(n3435) );
  XOR2_X1 U18522 ( .A1(n63011), .A2(n38710), .Z(n8500) );
  XOR2_X1 U18534 ( .A1(n3429), .A2(n64241), .Z(n38487) );
  XOR2_X1 U18548 ( .A1(n32099), .A2(n57842), .Z(n2260) );
  XOR2_X1 U18558 ( .A1(n33177), .A2(n23491), .Z(n57842) );
  NAND3_X2 U18589 ( .A1(n21165), .A2(n21167), .A3(n57846), .ZN(n21166) );
  NOR2_X2 U18660 ( .A1(n57851), .A2(n42723), .ZN(n58457) );
  NAND2_X2 U18665 ( .A1(n42721), .A2(n61891), .ZN(n57851) );
  NAND3_X2 U18672 ( .A1(n61231), .A2(n45686), .A3(n45687), .ZN(n48294) );
  INV_X1 U18693 ( .I(n741), .ZN(n57854) );
  AOI21_X1 U18706 ( .A1(n25046), .A2(n45504), .B(n6786), .ZN(n57856) );
  NOR3_X2 U18719 ( .A1(n11430), .A2(n57862), .A3(n57861), .ZN(n11429) );
  NAND2_X1 U18726 ( .A1(n30200), .A2(n30201), .ZN(n57861) );
  NAND2_X2 U18730 ( .A1(n34763), .A2(n15830), .ZN(n18440) );
  NOR2_X2 U18737 ( .A1(n34766), .A2(n34309), .ZN(n34763) );
  NAND2_X2 U18742 ( .A1(n2532), .A2(n57863), .ZN(n24357) );
  NOR3_X2 U18744 ( .A1(n61868), .A2(n21258), .A3(n2535), .ZN(n57863) );
  NAND3_X2 U18755 ( .A1(n17069), .A2(n57274), .A3(n57865), .ZN(n21187) );
  INV_X1 U18764 ( .I(n57866), .ZN(n57865) );
  OAI22_X1 U18772 ( .A1(n34314), .A2(n34315), .B1(n34313), .B2(n34312), .ZN(
        n57866) );
  XOR2_X1 U18779 ( .A1(n23957), .A2(n46118), .Z(n9010) );
  XOR2_X1 U18781 ( .A1(n44736), .A2(n58586), .Z(n46118) );
  NAND2_X2 U18804 ( .A1(n4415), .A2(n27196), .ZN(n57868) );
  NAND2_X2 U18816 ( .A1(n50343), .A2(n60099), .ZN(n11504) );
  XOR2_X1 U18818 ( .A1(n57869), .A2(n31294), .Z(n22732) );
  XOR2_X1 U18823 ( .A1(n46668), .A2(n13998), .Z(n13997) );
  NAND4_X1 U18827 ( .A1(n26366), .A2(n27580), .A3(n22541), .A4(n26660), .ZN(
        n26367) );
  OR2_X1 U18862 ( .A1(n25465), .A2(n26214), .Z(n12547) );
  XOR2_X1 U18888 ( .A1(n30717), .A2(n44797), .Z(n22472) );
  XOR2_X1 U18902 ( .A1(n37836), .A2(n52461), .Z(n44797) );
  XOR2_X1 U18903 ( .A1(n57870), .A2(n17402), .Z(n24547) );
  XOR2_X1 U18904 ( .A1(n30733), .A2(n19627), .Z(n57870) );
  XOR2_X1 U18910 ( .A1(n57871), .A2(n52154), .Z(n7612) );
  XOR2_X1 U18912 ( .A1(n1197), .A2(n52153), .Z(n57871) );
  OR2_X1 U18919 ( .A1(n24836), .A2(n57872), .Z(n26557) );
  NAND2_X1 U18925 ( .A1(n47603), .A2(n47819), .ZN(n45967) );
  OR2_X1 U18930 ( .A1(n16939), .A2(n33561), .Z(n18070) );
  XOR2_X1 U18934 ( .A1(n61955), .A2(n43764), .Z(n43906) );
  NOR2_X1 U18940 ( .A1(n45562), .A2(n59813), .ZN(n17563) );
  XOR2_X1 U18941 ( .A1(n32057), .A2(n33906), .Z(n22336) );
  NAND3_X2 U18943 ( .A1(n19178), .A2(n29742), .A3(n19179), .ZN(n32057) );
  NAND4_X2 U18958 ( .A1(n34409), .A2(n34410), .A3(n34407), .A4(n34408), .ZN(
        n57874) );
  INV_X2 U18970 ( .I(n29269), .ZN(n13731) );
  NAND2_X2 U18971 ( .A1(n13055), .A2(n13056), .ZN(n29269) );
  INV_X1 U18973 ( .I(n54272), .ZN(n21288) );
  NAND2_X2 U18975 ( .A1(n7784), .A2(n51709), .ZN(n54272) );
  XOR2_X1 U18976 ( .A1(n11205), .A2(n29580), .Z(n28430) );
  OAI21_X1 U18998 ( .A1(n48293), .A2(n1468), .B(n20458), .ZN(n57878) );
  NAND3_X2 U19043 ( .A1(n1381), .A2(n50398), .A3(n58840), .ZN(n49731) );
  OR2_X1 U19052 ( .A1(n18225), .A2(n49541), .Z(n57881) );
  XOR2_X1 U19065 ( .A1(n57882), .A2(n15056), .Z(n15055) );
  XOR2_X1 U19067 ( .A1(n15401), .A2(n46656), .Z(n57882) );
  XOR2_X1 U19070 ( .A1(n57883), .A2(n6512), .Z(n16945) );
  XOR2_X1 U19079 ( .A1(n52529), .A2(n5778), .Z(n57883) );
  XOR2_X1 U19092 ( .A1(n57885), .A2(n59228), .Z(n59296) );
  XOR2_X1 U19098 ( .A1(n60188), .A2(n46345), .Z(n57885) );
  OR2_X2 U19107 ( .A1(n19006), .A2(n9762), .Z(n32435) );
  XOR2_X1 U19168 ( .A1(n9876), .A2(n57888), .Z(n3375) );
  XOR2_X1 U19169 ( .A1(n7847), .A2(n37570), .Z(n57888) );
  NAND2_X2 U19172 ( .A1(n4263), .A2(n36404), .ZN(n36408) );
  NAND2_X2 U19176 ( .A1(n48063), .A2(n59808), .ZN(n47354) );
  XOR2_X1 U19202 ( .A1(n18098), .A2(n45400), .Z(n61102) );
  NAND2_X2 U19215 ( .A1(n22637), .A2(n61419), .ZN(n25676) );
  XOR2_X1 U19263 ( .A1(n1466), .A2(n50964), .Z(n25968) );
  NAND2_X2 U19270 ( .A1(n5580), .A2(n5579), .ZN(n50964) );
  XOR2_X1 U19283 ( .A1(n50997), .A2(n25005), .Z(n8123) );
  XOR2_X1 U19298 ( .A1(n7320), .A2(n8179), .Z(n50997) );
  AOI21_X1 U19335 ( .A1(n40612), .A2(n61308), .B(n59574), .ZN(n19296) );
  CLKBUF_X12 U19340 ( .I(n24918), .Z(n57894) );
  NAND2_X1 U19348 ( .A1(n57896), .A2(n4827), .ZN(n4826) );
  INV_X2 U19382 ( .I(n57735), .ZN(n48953) );
  NOR2_X2 U19400 ( .A1(n53036), .A2(n24415), .ZN(n25127) );
  NAND2_X1 U19402 ( .A1(n46086), .A2(n46085), .ZN(n4012) );
  XOR2_X1 U19418 ( .A1(n57900), .A2(n44499), .Z(n45726) );
  XOR2_X1 U19422 ( .A1(n44497), .A2(n7162), .Z(n57900) );
  OR2_X1 U19427 ( .A1(n55794), .A2(n55820), .Z(n11688) );
  NAND2_X2 U19429 ( .A1(n55821), .A2(n55812), .ZN(n55794) );
  NOR2_X2 U19460 ( .A1(n13842), .A2(n12897), .ZN(n7627) );
  NAND3_X2 U19461 ( .A1(n13845), .A2(n25181), .A3(n13843), .ZN(n13842) );
  OR2_X1 U19472 ( .A1(n55738), .A2(n55728), .Z(n52926) );
  AOI22_X2 U19477 ( .A1(n14241), .A2(n11410), .B1(n23949), .B2(n37866), .ZN(
        n14242) );
  INV_X2 U19487 ( .I(n51214), .ZN(n57908) );
  NAND3_X2 U19490 ( .A1(n57910), .A2(n57909), .A3(n41228), .ZN(n41242) );
  AND2_X1 U19505 ( .A1(n41226), .A2(n41225), .Z(n57909) );
  XOR2_X1 U19506 ( .A1(n57911), .A2(n52970), .Z(Plaintext[102]) );
  OAI22_X1 U19529 ( .A1(n57893), .A2(n23167), .B1(n44840), .B2(n47575), .ZN(
        n44858) );
  NOR2_X2 U19530 ( .A1(n47570), .A2(n47901), .ZN(n177) );
  INV_X2 U19549 ( .I(n57912), .ZN(n49331) );
  NOR2_X2 U19550 ( .A1(n49384), .A2(n15693), .ZN(n57912) );
  OR2_X2 U19552 ( .A1(n43733), .A2(n18104), .Z(n42843) );
  XOR2_X1 U19553 ( .A1(n1943), .A2(n61240), .Z(n5263) );
  NAND3_X1 U19570 ( .A1(n35024), .A2(n1803), .A3(n33520), .ZN(n61312) );
  NAND3_X1 U19578 ( .A1(n41369), .A2(n42677), .A3(n6706), .ZN(n4609) );
  XNOR2_X1 U19596 ( .A1(n46433), .A2(n24278), .ZN(n57918) );
  XOR2_X1 U19603 ( .A1(n57919), .A2(n23989), .Z(Plaintext[157]) );
  NAND2_X2 U19623 ( .A1(n57920), .A2(n12548), .ZN(n98) );
  NAND3_X2 U19631 ( .A1(n242), .A2(n60054), .A3(n34520), .ZN(n57920) );
  NAND4_X2 U19641 ( .A1(n50138), .A2(n50139), .A3(n49144), .A4(n60786), .ZN(
        n57921) );
  OR2_X2 U19644 ( .A1(n23936), .A2(n55135), .Z(n55166) );
  NOR2_X2 U19663 ( .A1(n10289), .A2(n57922), .ZN(n56451) );
  NOR2_X2 U19683 ( .A1(n58513), .A2(n55476), .ZN(n52932) );
  INV_X2 U19730 ( .I(n19768), .ZN(n46553) );
  XOR2_X1 U19731 ( .A1(n46213), .A2(n57926), .Z(n19768) );
  INV_X1 U19738 ( .I(n55349), .ZN(n57926) );
  AOI22_X2 U19741 ( .A1(n57927), .A2(n28341), .B1(n26054), .B2(n28352), .ZN(
        n4415) );
  INV_X2 U19758 ( .I(n26680), .ZN(n57927) );
  NAND2_X2 U19764 ( .A1(n7975), .A2(n5124), .ZN(n26680) );
  NOR2_X1 U19778 ( .A1(n57978), .A2(n18396), .ZN(n41100) );
  AND2_X1 U19785 ( .A1(n37168), .A2(n59362), .Z(n13890) );
  OR2_X1 U19818 ( .A1(n16601), .A2(n37529), .Z(n41001) );
  XOR2_X1 U19862 ( .A1(n57930), .A2(n23968), .Z(Plaintext[161]) );
  NAND4_X2 U19876 ( .A1(n56526), .A2(n56525), .A3(n59779), .A4(n59780), .ZN(
        n57930) );
  XOR2_X1 U19945 ( .A1(n61947), .A2(n13183), .Z(n57931) );
  INV_X4 U19946 ( .I(n15556), .ZN(n15557) );
  NOR2_X2 U19957 ( .A1(n57935), .A2(n41938), .ZN(n43549) );
  NOR2_X2 U19961 ( .A1(n60715), .A2(n60716), .ZN(n1466) );
  XOR2_X1 U19963 ( .A1(n57936), .A2(n43407), .Z(n43597) );
  XOR2_X1 U19965 ( .A1(n43406), .A2(n44920), .Z(n57936) );
  AOI21_X1 U19966 ( .A1(n61543), .A2(n62952), .B(n59697), .ZN(n59696) );
  OAI21_X1 U19967 ( .A1(n2915), .A2(n2914), .B(n59696), .ZN(n15596) );
  XOR2_X1 U19969 ( .A1(n43807), .A2(n43390), .Z(n43405) );
  NAND2_X2 U19970 ( .A1(n15007), .A2(n20942), .ZN(n58210) );
  OAI22_X1 U19972 ( .A1(n27369), .A2(n27010), .B1(n28225), .B2(n5627), .ZN(
        n27011) );
  INV_X4 U19973 ( .I(n13443), .ZN(n31189) );
  AND2_X1 U19983 ( .A1(n58179), .A2(n58178), .Z(n57938) );
  XOR2_X1 U19994 ( .A1(n52079), .A2(n51551), .Z(n51552) );
  NAND3_X2 U19997 ( .A1(n48762), .A2(n48761), .A3(n48763), .ZN(n52079) );
  AOI22_X1 U20003 ( .A1(n47026), .A2(n45529), .B1(n45528), .B2(n47035), .ZN(
        n45544) );
  NOR3_X2 U20009 ( .A1(n5865), .A2(n57941), .A3(n5864), .ZN(n12878) );
  NAND2_X1 U20014 ( .A1(n58900), .A2(n58898), .ZN(n35151) );
  OAI21_X1 U20015 ( .A1(n35949), .A2(n15171), .B(n36921), .ZN(n20611) );
  NAND2_X1 U20018 ( .A1(n23434), .A2(n43151), .ZN(n58180) );
  NOR2_X1 U20043 ( .A1(n34289), .A2(n17144), .ZN(n37437) );
  XOR2_X1 U20047 ( .A1(n38859), .A2(n3499), .Z(n39303) );
  INV_X2 U20050 ( .I(n57894), .ZN(n38859) );
  XOR2_X1 U20054 ( .A1(n38835), .A2(n39566), .Z(n24918) );
  NAND2_X2 U20055 ( .A1(n5196), .A2(n5198), .ZN(n5193) );
  NAND2_X1 U20056 ( .A1(n19326), .A2(n19325), .ZN(n57945) );
  INV_X1 U20060 ( .I(n56503), .ZN(n56485) );
  XOR2_X1 U20061 ( .A1(n44897), .A2(n42391), .Z(n11922) );
  OAI22_X2 U20064 ( .A1(n10798), .A2(n59048), .B1(n42389), .B2(n42390), .ZN(
        n44897) );
  NAND2_X2 U20068 ( .A1(n59407), .A2(n57947), .ZN(n37492) );
  NAND2_X2 U20071 ( .A1(n22587), .A2(n19322), .ZN(n36943) );
  XOR2_X1 U20085 ( .A1(n24458), .A2(n61100), .Z(n59305) );
  XNOR2_X1 U20087 ( .A1(n9752), .A2(n50876), .ZN(n59625) );
  NOR2_X1 U20089 ( .A1(n42177), .A2(n16545), .ZN(n59943) );
  OR2_X1 U20092 ( .A1(n57197), .A2(n40020), .Z(n18794) );
  NOR2_X2 U20097 ( .A1(n17293), .A2(n57951), .ZN(n6820) );
  NAND3_X2 U20100 ( .A1(n28737), .A2(n28738), .A3(n28739), .ZN(n57951) );
  NAND2_X2 U20118 ( .A1(n57953), .A2(n57952), .ZN(n28782) );
  INV_X1 U20119 ( .I(n22374), .ZN(n57952) );
  XOR2_X1 U20120 ( .A1(n50505), .A2(n52029), .Z(n38400) );
  XOR2_X1 U20121 ( .A1(n53344), .A2(n23754), .Z(n52029) );
  XOR2_X1 U20122 ( .A1(n26044), .A2(n39291), .Z(n6161) );
  XOR2_X1 U20123 ( .A1(n37821), .A2(n39769), .Z(n39291) );
  BUF_X2 U20124 ( .I(n1926), .Z(n57954) );
  XOR2_X1 U20136 ( .A1(n57956), .A2(n24248), .Z(n2578) );
  XOR2_X1 U20137 ( .A1(n39552), .A2(n19008), .Z(n57956) );
  XOR2_X1 U20138 ( .A1(n46396), .A2(n33832), .Z(n33833) );
  XOR2_X1 U20139 ( .A1(n50621), .A2(n56322), .Z(n46396) );
  NAND2_X2 U20154 ( .A1(n57957), .A2(n8533), .ZN(n6302) );
  NAND2_X2 U20163 ( .A1(n60726), .A2(n6411), .ZN(n48422) );
  NAND2_X1 U20164 ( .A1(n9692), .A2(n49014), .ZN(n15471) );
  NOR2_X2 U20167 ( .A1(n60021), .A2(n60602), .ZN(n982) );
  NAND2_X2 U20170 ( .A1(n57964), .A2(n57963), .ZN(n49375) );
  NOR2_X1 U20174 ( .A1(n47890), .A2(n47891), .ZN(n57964) );
  NAND2_X1 U20175 ( .A1(n42784), .A2(n42788), .ZN(n16262) );
  XOR2_X1 U20178 ( .A1(n57965), .A2(n61507), .Z(n12027) );
  XOR2_X1 U20183 ( .A1(n20272), .A2(n57966), .Z(n3231) );
  XOR2_X1 U20184 ( .A1(n38262), .A2(n57376), .Z(n57966) );
  AOI22_X2 U20194 ( .A1(n49531), .A2(n7358), .B1(n49530), .B2(n18769), .ZN(
        n60577) );
  XOR2_X1 U20195 ( .A1(n52207), .A2(n57113), .Z(n49189) );
  OR2_X1 U20199 ( .A1(n60969), .A2(n25746), .Z(n52763) );
  NAND3_X1 U20204 ( .A1(n36009), .A2(n19553), .A3(n61747), .ZN(n19552) );
  AOI21_X2 U20216 ( .A1(n2074), .A2(n2073), .B(n2072), .ZN(n24005) );
  OAI22_X2 U20217 ( .A1(n31285), .A2(n31284), .B1(n31287), .B2(n31286), .ZN(
        n31378) );
  NOR2_X2 U20222 ( .A1(n57970), .A2(n46904), .ZN(n16590) );
  NAND2_X2 U20228 ( .A1(n21453), .A2(n10237), .ZN(n52874) );
  INV_X2 U20237 ( .I(n61705), .ZN(n59158) );
  INV_X1 U20238 ( .I(n42651), .ZN(n57974) );
  INV_X2 U20252 ( .I(n1757), .ZN(n57975) );
  XOR2_X1 U20255 ( .A1(n20288), .A2(n39354), .Z(n57976) );
  NAND2_X2 U20274 ( .A1(n24081), .A2(n47748), .ZN(n18138) );
  NAND2_X2 U20276 ( .A1(n17133), .A2(n16657), .ZN(n57978) );
  NAND2_X2 U20284 ( .A1(n19294), .A2(n48685), .ZN(n17672) );
  NAND2_X2 U20285 ( .A1(n24325), .A2(n20094), .ZN(n23984) );
  NOR3_X2 U20299 ( .A1(n10550), .A2(n37400), .A3(n24041), .ZN(n36331) );
  BUF_X2 U20308 ( .I(n24103), .Z(n57984) );
  OAI21_X1 U20320 ( .A1(n13605), .A2(n42340), .B(n59746), .ZN(n57987) );
  NAND2_X2 U20336 ( .A1(n8688), .A2(n40570), .ZN(n59225) );
  XOR2_X1 U20340 ( .A1(n50906), .A2(n62455), .Z(n20169) );
  XOR2_X1 U20364 ( .A1(n13664), .A2(n57992), .Z(n26021) );
  XOR2_X1 U20367 ( .A1(n38468), .A2(n56949), .Z(n57992) );
  NOR2_X1 U20406 ( .A1(n54880), .A2(n54904), .ZN(n57996) );
  NOR2_X2 U20408 ( .A1(n58000), .A2(n57999), .ZN(n5013) );
  AND2_X1 U20415 ( .A1(n39992), .A2(n41378), .Z(n41123) );
  NAND2_X2 U20425 ( .A1(n4540), .A2(n53803), .ZN(n53774) );
  NOR2_X2 U20440 ( .A1(n47211), .A2(n48459), .ZN(n48126) );
  XOR2_X1 U20457 ( .A1(n49210), .A2(n49209), .Z(n51102) );
  XOR2_X1 U20458 ( .A1(n23690), .A2(n20403), .Z(n60840) );
  NAND3_X2 U20470 ( .A1(n25590), .A2(n20791), .A3(n35366), .ZN(n39346) );
  XOR2_X1 U20483 ( .A1(n39630), .A2(n17002), .Z(n58013) );
  XOR2_X1 U20484 ( .A1(n59679), .A2(n58378), .Z(n58014) );
  AOI21_X1 U20487 ( .A1(n664), .A2(n41306), .B(n41805), .ZN(n3493) );
  NAND2_X1 U20503 ( .A1(n17513), .A2(n45610), .ZN(n58016) );
  BUF_X2 U20521 ( .I(n5472), .Z(n58020) );
  NOR3_X2 U20522 ( .A1(n42844), .A2(n16232), .A3(n16607), .ZN(n10532) );
  OR2_X1 U20531 ( .A1(n23721), .A2(n49745), .Z(n60716) );
  NAND2_X2 U20533 ( .A1(n10983), .A2(n56268), .ZN(n56265) );
  NOR2_X2 U20545 ( .A1(n58022), .A2(n3583), .ZN(n14908) );
  NAND3_X2 U20546 ( .A1(n484), .A2(n3585), .A3(n37033), .ZN(n58022) );
  NAND2_X2 U20549 ( .A1(n59583), .A2(n41064), .ZN(n40845) );
  NAND3_X1 U20554 ( .A1(n27642), .A2(n27856), .A3(n23033), .ZN(n20050) );
  AOI22_X1 U20557 ( .A1(n19920), .A2(n27357), .B1(n19919), .B2(n29320), .ZN(
        n19918) );
  XOR2_X1 U20559 ( .A1(n38619), .A2(n58024), .Z(n5783) );
  XOR2_X1 U20562 ( .A1(n5785), .A2(n39768), .Z(n58024) );
  XOR2_X1 U20564 ( .A1(n58025), .A2(n19149), .Z(n9509) );
  XOR2_X1 U20566 ( .A1(n48753), .A2(n48752), .Z(n58025) );
  OR2_X1 U20569 ( .A1(n3582), .A2(n31539), .Z(n3581) );
  AND2_X2 U20570 ( .A1(n61735), .A2(n59272), .Z(n12539) );
  XOR2_X1 U20574 ( .A1(n58029), .A2(n39675), .Z(n25628) );
  XOR2_X1 U20578 ( .A1(n17845), .A2(n39587), .Z(n58029) );
  INV_X1 U20583 ( .I(n56264), .ZN(n1284) );
  AND2_X1 U20584 ( .A1(n56264), .A2(n15706), .Z(n5496) );
  OAI22_X2 U20590 ( .A1(n44559), .A2(n45505), .B1(n58705), .B2(n46950), .ZN(
        n58031) );
  NAND2_X1 U20592 ( .A1(n4334), .A2(n4335), .ZN(n4333) );
  NAND2_X1 U20596 ( .A1(n49968), .A2(n49969), .ZN(n49971) );
  OAI21_X2 U20607 ( .A1(n4187), .A2(n29168), .B(n18375), .ZN(n58215) );
  XOR2_X1 U20615 ( .A1(n39779), .A2(n61656), .Z(n58035) );
  OR2_X2 U20621 ( .A1(n21303), .A2(n48097), .Z(n47115) );
  NAND3_X2 U20624 ( .A1(n1832), .A2(n24869), .A3(n24868), .ZN(n5877) );
  XOR2_X1 U20628 ( .A1(n11828), .A2(n39728), .Z(n26146) );
  NAND2_X1 U20634 ( .A1(n59992), .A2(n48196), .ZN(n58042) );
  NOR2_X2 U20641 ( .A1(n2608), .A2(n50353), .ZN(n50366) );
  NAND2_X2 U20642 ( .A1(n9229), .A2(n23394), .ZN(n50353) );
  XOR2_X1 U20645 ( .A1(n59559), .A2(n58045), .Z(n21625) );
  XOR2_X1 U20647 ( .A1(n23827), .A2(n39257), .Z(n58045) );
  OR2_X2 U20668 ( .A1(n13418), .A2(n826), .Z(n48745) );
  NAND2_X2 U20675 ( .A1(n36838), .A2(n36851), .ZN(n60374) );
  NAND2_X1 U20708 ( .A1(n16524), .A2(n27833), .ZN(n26831) );
  INV_X2 U20723 ( .I(n18180), .ZN(n61647) );
  NAND2_X1 U20729 ( .A1(n22430), .A2(n25393), .ZN(n56300) );
  NOR2_X1 U20735 ( .A1(n23501), .A2(n3705), .ZN(n42519) );
  INV_X2 U20741 ( .I(n16912), .ZN(n3705) );
  XOR2_X1 U20742 ( .A1(n16795), .A2(n16251), .Z(n16912) );
  XNOR2_X1 U20743 ( .A1(n25316), .A2(n51010), .ZN(n58055) );
  NOR2_X1 U20751 ( .A1(n43549), .A2(n62535), .ZN(n43412) );
  XOR2_X1 U20752 ( .A1(n20874), .A2(n5603), .Z(n50114) );
  NAND2_X1 U20758 ( .A1(n47041), .A2(n6704), .ZN(n49487) );
  NAND3_X1 U20773 ( .A1(n16742), .A2(n46013), .A3(n12360), .ZN(n46020) );
  NOR2_X2 U20780 ( .A1(n16750), .A2(n22504), .ZN(n30339) );
  XOR2_X1 U20786 ( .A1(n58058), .A2(n8301), .Z(n3975) );
  XOR2_X1 U20787 ( .A1(n37867), .A2(n38716), .Z(n58058) );
  OAI21_X2 U20791 ( .A1(n22413), .A2(n65232), .B(n34131), .ZN(n33394) );
  NAND2_X2 U20794 ( .A1(n61598), .A2(n33390), .ZN(n34131) );
  XOR2_X1 U20800 ( .A1(n2911), .A2(n58061), .Z(n42819) );
  XOR2_X1 U20801 ( .A1(n25432), .A2(n831), .Z(n58061) );
  NAND2_X1 U20802 ( .A1(n23766), .A2(n61517), .ZN(n58062) );
  XOR2_X1 U20811 ( .A1(n58065), .A2(n20932), .Z(n37816) );
  XOR2_X1 U20815 ( .A1(n38181), .A2(n37814), .Z(n58065) );
  NAND3_X2 U20816 ( .A1(n31025), .A2(n31024), .A3(n31023), .ZN(n10478) );
  NOR2_X2 U20823 ( .A1(n11638), .A2(n29084), .ZN(n30620) );
  NAND3_X2 U20824 ( .A1(n16751), .A2(n28556), .A3(n28555), .ZN(n11638) );
  BUF_X4 U20825 ( .I(n53950), .Z(n54006) );
  NOR2_X2 U20833 ( .A1(n38926), .A2(n61094), .ZN(n22168) );
  NAND2_X2 U20841 ( .A1(n55820), .A2(n55812), .ZN(n55817) );
  OR2_X1 U20858 ( .A1(n36644), .A2(n37942), .Z(n58069) );
  XOR2_X1 U20874 ( .A1(n39482), .A2(n37347), .Z(n23204) );
  NAND2_X2 U20892 ( .A1(n35480), .A2(n23778), .ZN(n58073) );
  XOR2_X1 U20895 ( .A1(n58075), .A2(n14586), .Z(n38922) );
  BUF_X2 U20899 ( .I(n46112), .Z(n58077) );
  XOR2_X1 U20901 ( .A1(n31360), .A2(n58078), .Z(n50790) );
  XOR2_X1 U20903 ( .A1(n44925), .A2(n45371), .Z(n31360) );
  XOR2_X1 U20906 ( .A1(n58079), .A2(n38308), .Z(n16893) );
  XOR2_X1 U20907 ( .A1(n61468), .A2(n39237), .Z(n58079) );
  INV_X4 U20908 ( .I(n61700), .ZN(n32984) );
  NAND3_X1 U20917 ( .A1(n23006), .A2(n25495), .A3(n10077), .ZN(n25491) );
  BUF_X2 U20918 ( .I(n34822), .Z(n58080) );
  XOR2_X1 U20921 ( .A1(n18547), .A2(n19527), .Z(n24388) );
  OAI22_X1 U20928 ( .A1(n58082), .A2(n27467), .B1(n27466), .B2(n27465), .ZN(
        n27476) );
  AND2_X1 U20932 ( .A1(n60033), .A2(n27460), .Z(n58082) );
  NAND3_X1 U20933 ( .A1(n60754), .A2(n1298), .A3(n14605), .ZN(n42194) );
  NAND2_X2 U20939 ( .A1(n15824), .A2(n47307), .ZN(n45957) );
  XOR2_X1 U20957 ( .A1(n58085), .A2(n40458), .Z(n32226) );
  XOR2_X1 U20958 ( .A1(n45112), .A2(n39360), .Z(n58085) );
  NAND2_X2 U20959 ( .A1(n3705), .A2(n41289), .ZN(n59976) );
  XOR2_X1 U20964 ( .A1(n38330), .A2(n39733), .Z(n58910) );
  NAND2_X2 U20966 ( .A1(n6705), .A2(n8912), .ZN(n42824) );
  NAND3_X1 U20968 ( .A1(n58088), .A2(n54973), .A3(n54799), .ZN(n54805) );
  XOR2_X1 U20971 ( .A1(n14128), .A2(n52569), .Z(n16593) );
  NOR2_X1 U20972 ( .A1(n41323), .A2(n41788), .ZN(n41324) );
  NAND4_X2 U20974 ( .A1(n11344), .A2(n46796), .A3(n11342), .A4(n46797), .ZN(
        n9789) );
  INV_X2 U20977 ( .I(n58089), .ZN(n6330) );
  XOR2_X1 U20978 ( .A1(Key[112]), .A2(Ciphertext[141]), .Z(n58089) );
  OAI22_X1 U20983 ( .A1(n58090), .A2(n1583), .B1(n56902), .B2(n18111), .ZN(
        n52293) );
  NOR2_X1 U20987 ( .A1(n59736), .A2(n56926), .ZN(n58090) );
  NAND3_X2 U20995 ( .A1(n6613), .A2(n57341), .A3(n19490), .ZN(n58091) );
  OR2_X1 U21002 ( .A1(n10839), .A2(n53546), .Z(n10838) );
  XOR2_X1 U21003 ( .A1(n51764), .A2(n51154), .Z(n22360) );
  XOR2_X1 U21005 ( .A1(n7229), .A2(n52424), .Z(n51764) );
  NAND3_X1 U21027 ( .A1(n3032), .A2(n5282), .A3(n49721), .ZN(n58096) );
  XOR2_X1 U21028 ( .A1(n58098), .A2(n1039), .Z(n45265) );
  XOR2_X1 U21031 ( .A1(n45264), .A2(n45260), .Z(n58098) );
  XOR2_X1 U21048 ( .A1(n24095), .A2(n16401), .Z(n31851) );
  NAND2_X2 U21069 ( .A1(n10456), .A2(n49213), .ZN(n8963) );
  XOR2_X1 U21072 ( .A1(n9737), .A2(n25423), .Z(n41165) );
  XOR2_X1 U21086 ( .A1(n23464), .A2(n23927), .Z(n24223) );
  INV_X2 U21103 ( .I(n58103), .ZN(n2666) );
  XOR2_X1 U21105 ( .A1(n3310), .A2(n23343), .Z(n58103) );
  XOR2_X1 U21113 ( .A1(n53672), .A2(n53688), .Z(n53645) );
  NOR2_X1 U21147 ( .A1(n17615), .A2(n37067), .ZN(n21839) );
  NOR2_X2 U21150 ( .A1(n20106), .A2(n20101), .ZN(n17615) );
  OAI21_X2 U21164 ( .A1(n21215), .A2(n58107), .B(n59769), .ZN(n147) );
  AOI21_X2 U21166 ( .A1(n14980), .A2(n4097), .B(n34113), .ZN(n58107) );
  NAND3_X1 U21169 ( .A1(n8259), .A2(n19020), .A3(n19021), .ZN(n55615) );
  NAND2_X2 U21172 ( .A1(n40729), .A2(n40728), .ZN(n41205) );
  NOR2_X1 U21174 ( .A1(n58109), .A2(n21590), .ZN(n50740) );
  XOR2_X1 U21181 ( .A1(n58111), .A2(n32650), .Z(n58302) );
  XOR2_X1 U21185 ( .A1(n32638), .A2(n15464), .Z(n33289) );
  NOR2_X2 U21196 ( .A1(n62120), .A2(n56812), .ZN(n56815) );
  INV_X4 U21197 ( .I(n25112), .ZN(n30695) );
  NAND2_X2 U21200 ( .A1(n59334), .A2(n59335), .ZN(n25112) );
  NOR3_X2 U21202 ( .A1(n23545), .A2(n5033), .A3(n23546), .ZN(n58112) );
  XOR2_X1 U21204 ( .A1(n58113), .A2(n39501), .Z(n24834) );
  XOR2_X1 U21212 ( .A1(n51474), .A2(n27640), .Z(n50625) );
  NAND4_X2 U21214 ( .A1(n49707), .A2(n49704), .A3(n49706), .A4(n49705), .ZN(
        n51474) );
  OAI21_X1 U21215 ( .A1(n40569), .A2(n39958), .B(n25943), .ZN(n18419) );
  NAND3_X2 U21217 ( .A1(n60549), .A2(n20654), .A3(n7741), .ZN(n7738) );
  NAND3_X2 U21219 ( .A1(n58963), .A2(n49535), .A3(n49536), .ZN(n18733) );
  INV_X2 U21224 ( .I(n58115), .ZN(n24391) );
  XOR2_X1 U21225 ( .A1(Ciphertext[180]), .A2(Key[97]), .Z(n58115) );
  AOI21_X2 U21230 ( .A1(n49485), .A2(n15724), .B(n7745), .ZN(n49507) );
  AND2_X1 U21231 ( .A1(n34327), .A2(n34326), .Z(n58160) );
  NAND2_X1 U21236 ( .A1(n46968), .A2(n57430), .ZN(n58116) );
  XOR2_X1 U21238 ( .A1(n58117), .A2(n32654), .Z(n24434) );
  XOR2_X1 U21240 ( .A1(n31828), .A2(n32338), .Z(n58117) );
  OR3_X2 U21260 ( .A1(n58766), .A2(n7878), .A3(n18764), .Z(n18765) );
  NOR2_X1 U21263 ( .A1(n23200), .A2(n27476), .ZN(n61609) );
  XOR2_X1 U21291 ( .A1(n8208), .A2(n944), .Z(n14732) );
  NAND3_X1 U21292 ( .A1(n2240), .A2(n6790), .A3(n53301), .ZN(n53307) );
  NAND2_X2 U21295 ( .A1(n2698), .A2(n2014), .ZN(n2240) );
  AND2_X1 U21299 ( .A1(n49631), .A2(n64406), .Z(n48385) );
  XOR2_X1 U21301 ( .A1(n44948), .A2(n46573), .Z(n44586) );
  NAND2_X2 U21305 ( .A1(n36723), .A2(n35349), .ZN(n20161) );
  NAND2_X2 U21306 ( .A1(n35345), .A2(n36725), .ZN(n36723) );
  NAND2_X2 U21309 ( .A1(n3935), .A2(n33467), .ZN(n7932) );
  OR2_X1 U21314 ( .A1(n2380), .A2(n49407), .Z(n58122) );
  NOR2_X2 U21315 ( .A1(n33598), .A2(n24688), .ZN(n33299) );
  NAND3_X2 U21318 ( .A1(n58124), .A2(n47226), .A3(n44651), .ZN(n44655) );
  XOR2_X1 U21325 ( .A1(n58125), .A2(n24053), .Z(n12509) );
  NAND2_X2 U21330 ( .A1(n15171), .A2(n34927), .ZN(n24358) );
  OR3_X1 U21335 ( .A1(n35399), .A2(n36130), .A3(n36803), .Z(n36142) );
  NOR2_X2 U21352 ( .A1(n18162), .A2(n58129), .ZN(n19285) );
  NOR2_X2 U21355 ( .A1(n58130), .A2(n35892), .ZN(n13172) );
  OAI21_X2 U21358 ( .A1(n35897), .A2(n35881), .B(n35880), .ZN(n58130) );
  XOR2_X1 U21359 ( .A1(n60204), .A2(n58131), .Z(n15777) );
  NOR2_X1 U21374 ( .A1(n58132), .A2(n15842), .ZN(n23793) );
  AOI21_X1 U21375 ( .A1(n28489), .A2(n27834), .B(n27664), .ZN(n58132) );
  NAND2_X1 U21376 ( .A1(n47802), .A2(n47801), .ZN(n58133) );
  INV_X1 U21381 ( .I(n45306), .ZN(n58134) );
  XOR2_X1 U21393 ( .A1(n11440), .A2(n11439), .Z(n58135) );
  NAND3_X1 U21395 ( .A1(n2104), .A2(n55463), .A3(n55476), .ZN(n55284) );
  INV_X2 U21404 ( .I(n4324), .ZN(n7748) );
  NOR2_X2 U21413 ( .A1(n47356), .A2(n23156), .ZN(n58136) );
  NOR2_X1 U21414 ( .A1(n19457), .A2(n34783), .ZN(n33775) );
  XOR2_X1 U21420 ( .A1(n19879), .A2(n58137), .Z(n19876) );
  NAND3_X1 U21426 ( .A1(n56615), .A2(n56704), .A3(n56722), .ZN(n56649) );
  NOR2_X1 U21428 ( .A1(n6376), .A2(n6377), .ZN(n6375) );
  AOI22_X1 U21437 ( .A1(n49058), .A2(n49057), .B1(n19294), .B2(n49056), .ZN(
        n49059) );
  XOR2_X1 U21461 ( .A1(n51911), .A2(n23173), .Z(n51202) );
  AOI21_X1 U21483 ( .A1(n2514), .A2(n20708), .B(n49790), .ZN(n47948) );
  NAND2_X2 U21484 ( .A1(n23802), .A2(n15220), .ZN(n2514) );
  XOR2_X1 U21489 ( .A1(n58147), .A2(n18831), .Z(n38621) );
  AOI21_X2 U21503 ( .A1(n36079), .A2(n23842), .B(n59277), .ZN(n58148) );
  INV_X4 U21504 ( .I(n27085), .ZN(n31129) );
  NAND3_X2 U21505 ( .A1(n27084), .A2(n27082), .A3(n27083), .ZN(n27085) );
  INV_X2 U21523 ( .I(n58852), .ZN(n31147) );
  NAND3_X2 U21524 ( .A1(n27686), .A2(n27687), .A3(n27685), .ZN(n58852) );
  NAND2_X2 U21525 ( .A1(n50738), .A2(n52739), .ZN(n58151) );
  NAND2_X2 U21528 ( .A1(n50238), .A2(n19634), .ZN(n14266) );
  XOR2_X1 U21530 ( .A1(n50879), .A2(n58152), .Z(n6975) );
  XOR2_X1 U21539 ( .A1(n51509), .A2(n11488), .Z(n58152) );
  NAND2_X2 U21540 ( .A1(n34639), .A2(n35037), .ZN(n15466) );
  INV_X4 U21544 ( .I(n58153), .ZN(n61107) );
  NOR2_X2 U21547 ( .A1(n5060), .A2(n39010), .ZN(n58153) );
  NAND2_X1 U21561 ( .A1(n3448), .A2(n15858), .ZN(n58154) );
  XOR2_X1 U21565 ( .A1(n61061), .A2(n38468), .Z(n38262) );
  AND2_X1 U21574 ( .A1(n22498), .A2(n28542), .Z(n26756) );
  NAND3_X2 U21576 ( .A1(n8018), .A2(n23279), .A3(n43897), .ZN(n43144) );
  XOR2_X1 U21577 ( .A1(n49626), .A2(n58157), .Z(n20770) );
  NAND2_X1 U21581 ( .A1(n9533), .A2(n2037), .ZN(n59373) );
  NAND3_X2 U21586 ( .A1(n16526), .A2(n38346), .A3(n41248), .ZN(n7993) );
  NAND2_X1 U21599 ( .A1(n21593), .A2(n25110), .ZN(n58158) );
  NAND2_X1 U21611 ( .A1(n1452), .A2(n5614), .ZN(n3543) );
  INV_X2 U21614 ( .I(n3285), .ZN(n1452) );
  NAND2_X2 U21615 ( .A1(n2040), .A2(n53163), .ZN(n3285) );
  NOR3_X2 U21616 ( .A1(n58160), .A2(n18799), .A3(n34325), .ZN(n59407) );
  OR2_X1 U21624 ( .A1(n28187), .A2(n59604), .Z(n15305) );
  OR2_X1 U21626 ( .A1(n3123), .A2(n50306), .Z(n49661) );
  NAND4_X2 U21628 ( .A1(n58163), .A2(n40975), .A3(n40976), .A4(n40977), .ZN(
        n40979) );
  NAND2_X1 U21629 ( .A1(n40960), .A2(n40959), .ZN(n58163) );
  AOI21_X1 U21630 ( .A1(n58164), .A2(n6865), .B(n13854), .ZN(n5566) );
  OAI21_X2 U21631 ( .A1(n8396), .A2(n8395), .B(n54979), .ZN(n55011) );
  NOR2_X2 U21633 ( .A1(n9229), .A2(n23394), .ZN(n49471) );
  INV_X4 U21636 ( .I(n9228), .ZN(n9229) );
  AND2_X1 U21641 ( .A1(n12443), .A2(n31241), .Z(n12442) );
  NAND2_X2 U21649 ( .A1(n16766), .A2(n16765), .ZN(n50213) );
  NAND2_X2 U21657 ( .A1(n57073), .A2(n57079), .ZN(n57068) );
  NOR2_X2 U21668 ( .A1(n58168), .A2(n6024), .ZN(n28690) );
  AOI21_X2 U21673 ( .A1(n26277), .A2(n26276), .B(n28032), .ZN(n58168) );
  AND2_X1 U21678 ( .A1(n33603), .A2(n33602), .Z(n58169) );
  OAI21_X1 U21679 ( .A1(n17879), .A2(n29374), .B(n29373), .ZN(n58667) );
  NAND2_X2 U21698 ( .A1(n8320), .A2(n8322), .ZN(n25638) );
  NOR3_X2 U21707 ( .A1(n59176), .A2(n59177), .A3(n25266), .ZN(n24444) );
  NOR2_X2 U21742 ( .A1(n24091), .A2(n55671), .ZN(n13774) );
  OAI22_X1 U21754 ( .A1(n10988), .A2(n17500), .B1(n55612), .B2(n55611), .ZN(
        n21032) );
  NOR2_X2 U21765 ( .A1(n35153), .A2(n35154), .ZN(n36490) );
  NAND2_X2 U21767 ( .A1(n10829), .A2(n36232), .ZN(n35154) );
  XOR2_X1 U21769 ( .A1(n51130), .A2(n58176), .Z(n4112) );
  XOR2_X1 U21770 ( .A1(n51522), .A2(n52541), .Z(n58176) );
  NOR2_X1 U21783 ( .A1(n43150), .A2(n43167), .ZN(n58178) );
  NAND4_X2 U21784 ( .A1(n54832), .A2(n54829), .A3(n54830), .A4(n54831), .ZN(
        n2348) );
  NAND3_X1 U21797 ( .A1(n30759), .A2(n31215), .A3(n30760), .ZN(n17505) );
  NOR3_X2 U21798 ( .A1(n1218), .A2(n19929), .A3(n7426), .ZN(n31215) );
  NOR2_X2 U21801 ( .A1(n23405), .A2(n17128), .ZN(n5532) );
  AOI22_X1 U21820 ( .A1(n54297), .A2(n54296), .B1(n54294), .B2(n54295), .ZN(
        n54305) );
  INV_X2 U21823 ( .I(n19148), .ZN(n18612) );
  NAND4_X2 U21825 ( .A1(n23285), .A2(n54358), .A3(n54357), .A4(n54359), .ZN(
        n58213) );
  XOR2_X1 U21832 ( .A1(n58185), .A2(n46159), .Z(n46160) );
  XOR2_X1 U21838 ( .A1(n46156), .A2(n46157), .Z(n58185) );
  XOR2_X1 U21841 ( .A1(n31666), .A2(n59909), .Z(n31667) );
  XOR2_X1 U21844 ( .A1(n9787), .A2(n31668), .Z(n32394) );
  XOR2_X1 U21845 ( .A1(n22244), .A2(n55610), .Z(n31668) );
  NAND3_X1 U21855 ( .A1(n899), .A2(n4175), .A3(n36325), .ZN(n12451) );
  AOI21_X2 U21861 ( .A1(n58187), .A2(n57375), .B(n58186), .ZN(n20262) );
  NAND2_X2 U21864 ( .A1(n8040), .A2(n47510), .ZN(n47505) );
  NAND2_X2 U21865 ( .A1(n58189), .A2(n11287), .ZN(n8040) );
  INV_X2 U21869 ( .I(n46262), .ZN(n58189) );
  NAND2_X2 U21893 ( .A1(n12835), .A2(n44077), .ZN(n4287) );
  OAI22_X1 U21896 ( .A1(n40843), .A2(n41051), .B1(n39795), .B2(n62241), .ZN(
        n39796) );
  XOR2_X1 U21897 ( .A1(n23264), .A2(n58193), .Z(n44260) );
  XOR2_X1 U21904 ( .A1(n6677), .A2(n44258), .Z(n58193) );
  INV_X4 U21905 ( .I(n58522), .ZN(n15738) );
  NAND2_X2 U21918 ( .A1(n11243), .A2(n23348), .ZN(n11704) );
  XOR2_X1 U21920 ( .A1(n51808), .A2(n51190), .Z(n6965) );
  XOR2_X1 U21921 ( .A1(n23054), .A2(n62989), .Z(n51190) );
  INV_X4 U21922 ( .I(n14054), .ZN(n12652) );
  NAND2_X2 U21930 ( .A1(n7226), .A2(n11579), .ZN(n14054) );
  NAND2_X2 U21933 ( .A1(n18278), .A2(n11278), .ZN(n25306) );
  INV_X2 U21948 ( .I(n59398), .ZN(n19663) );
  NOR2_X2 U21952 ( .A1(n4685), .A2(n19373), .ZN(n18180) );
  XOR2_X1 U21958 ( .A1(n58201), .A2(n44518), .Z(n5766) );
  NOR3_X2 U21960 ( .A1(n15491), .A2(n15492), .A3(n15490), .ZN(n44518) );
  INV_X2 U21961 ( .I(n25621), .ZN(n61361) );
  NAND2_X2 U21962 ( .A1(n12786), .A2(n7228), .ZN(n25621) );
  XOR2_X1 U21965 ( .A1(n11236), .A2(n31630), .Z(n20143) );
  XOR2_X1 U21966 ( .A1(n33863), .A2(n32669), .Z(n11236) );
  XOR2_X1 U21972 ( .A1(n22101), .A2(n50318), .Z(n50783) );
  BUF_X2 U21978 ( .I(n37670), .Z(n58203) );
  XOR2_X1 U22000 ( .A1(n58207), .A2(n6331), .Z(n11373) );
  AND3_X1 U22010 ( .A1(n49982), .A2(n49981), .A3(n49983), .Z(n58208) );
  NOR2_X2 U22016 ( .A1(n28167), .A2(n58211), .ZN(n31097) );
  XOR2_X1 U22029 ( .A1(n58213), .A2(n54360), .Z(Plaintext[66]) );
  NOR2_X2 U22030 ( .A1(n19588), .A2(n31104), .ZN(n9787) );
  AOI21_X2 U22035 ( .A1(n4982), .A2(n31096), .B(n64484), .ZN(n19588) );
  NAND2_X2 U22047 ( .A1(n6369), .A2(n6370), .ZN(n26849) );
  NOR3_X2 U22056 ( .A1(n57210), .A2(n20147), .A3(n15720), .ZN(n58267) );
  NOR2_X2 U22062 ( .A1(n56719), .A2(n56722), .ZN(n7977) );
  INV_X2 U22064 ( .I(n56616), .ZN(n56722) );
  INV_X2 U22075 ( .I(n2928), .ZN(n1521) );
  OR2_X1 U22084 ( .A1(n6841), .A2(n16461), .Z(n12999) );
  OAI22_X1 U22085 ( .A1(n17862), .A2(n57123), .B1(n25147), .B2(n57108), .ZN(
        n57089) );
  INV_X2 U22091 ( .I(n21828), .ZN(n17862) );
  NOR2_X2 U22095 ( .A1(n21829), .A2(n21570), .ZN(n21828) );
  NAND2_X1 U22117 ( .A1(n24649), .A2(n21506), .ZN(n18659) );
  XOR2_X1 U22119 ( .A1(n39987), .A2(n38758), .Z(n21506) );
  NOR2_X2 U22124 ( .A1(n24352), .A2(n24353), .ZN(n57051) );
  NAND4_X2 U22125 ( .A1(n10733), .A2(n10731), .A3(n61913), .A4(n10732), .ZN(
        n31104) );
  BUF_X2 U22134 ( .I(n22503), .Z(n58220) );
  BUF_X4 U22136 ( .I(n15693), .Z(n61513) );
  NAND3_X2 U22139 ( .A1(n59141), .A2(n13109), .A3(n59140), .ZN(n19527) );
  NOR2_X2 U22141 ( .A1(n49459), .A2(n49739), .ZN(n19756) );
  XOR2_X1 U22150 ( .A1(n50990), .A2(n57371), .Z(n1111) );
  XOR2_X1 U22161 ( .A1(n30989), .A2(n58221), .Z(n30993) );
  XOR2_X1 U22164 ( .A1(n14866), .A2(n30990), .Z(n58221) );
  XOR2_X1 U22165 ( .A1(n246), .A2(n15876), .Z(n58348) );
  XOR2_X1 U22168 ( .A1(n51937), .A2(n52159), .Z(n15876) );
  XOR2_X1 U22169 ( .A1(n52157), .A2(n61137), .Z(n58357) );
  NOR3_X2 U22174 ( .A1(n13080), .A2(n58223), .A3(n58222), .ZN(n20796) );
  AOI21_X1 U22176 ( .A1(n55217), .A2(n55235), .B(n55208), .ZN(n55198) );
  NOR2_X2 U22177 ( .A1(n16943), .A2(n55231), .ZN(n55235) );
  NAND3_X2 U22179 ( .A1(n22753), .A2(n41752), .A3(n41753), .ZN(n44723) );
  NOR2_X2 U22189 ( .A1(n14428), .A2(n3251), .ZN(n55339) );
  NAND3_X2 U22191 ( .A1(n18383), .A2(n58227), .A3(n58226), .ZN(n24323) );
  NAND2_X1 U22206 ( .A1(n18381), .A2(n33823), .ZN(n58227) );
  XOR2_X1 U22219 ( .A1(n60107), .A2(n39756), .Z(n7216) );
  NAND3_X2 U22224 ( .A1(n17718), .A2(n17717), .A3(n58229), .ZN(n17715) );
  NAND3_X1 U22225 ( .A1(n29917), .A2(n29564), .A3(n29566), .ZN(n58229) );
  XOR2_X1 U22255 ( .A1(n13104), .A2(n52364), .Z(n52383) );
  NAND2_X2 U22261 ( .A1(n61816), .A2(n3227), .ZN(n39936) );
  AOI21_X1 U22264 ( .A1(n28703), .A2(n29007), .B(n24949), .ZN(n6085) );
  NAND2_X2 U22265 ( .A1(n2795), .A2(n30391), .ZN(n28703) );
  BUF_X2 U22266 ( .I(n1816), .Z(n58231) );
  OR3_X1 U22270 ( .A1(n5982), .A2(n27098), .A3(n26568), .Z(n26572) );
  NAND2_X2 U22273 ( .A1(n58233), .A2(n58232), .ZN(n2026) );
  XOR2_X1 U22274 ( .A1(n3420), .A2(n3421), .Z(n3419) );
  NOR2_X2 U22276 ( .A1(n59245), .A2(n58036), .ZN(n35015) );
  NAND2_X2 U22277 ( .A1(n22326), .A2(n25444), .ZN(n46907) );
  OAI21_X1 U22279 ( .A1(n27899), .A2(n27898), .B(n31187), .ZN(n58236) );
  OR2_X1 U22282 ( .A1(n58867), .A2(n44578), .Z(n2511) );
  BUF_X2 U22294 ( .I(n27789), .Z(n58237) );
  NAND2_X2 U22295 ( .A1(n21104), .A2(n36691), .ZN(n8039) );
  NAND2_X2 U22297 ( .A1(n11088), .A2(n16891), .ZN(n21104) );
  XOR2_X1 U22306 ( .A1(n32355), .A2(n58238), .Z(n3841) );
  XOR2_X1 U22323 ( .A1(n37657), .A2(n4779), .Z(n58240) );
  NAND2_X2 U22330 ( .A1(n58241), .A2(n17326), .ZN(n12502) );
  NAND2_X2 U22335 ( .A1(n10134), .A2(n32875), .ZN(n33433) );
  OR2_X1 U22339 ( .A1(n37091), .A2(n57686), .Z(n35079) );
  NOR2_X1 U22345 ( .A1(n4980), .A2(n4981), .ZN(n58575) );
  NAND2_X2 U22348 ( .A1(n57428), .A2(n43356), .ZN(n46166) );
  XNOR2_X1 U22349 ( .A1(n60832), .A2(n49127), .ZN(n58296) );
  NOR2_X1 U22351 ( .A1(n34542), .A2(n33723), .ZN(n58243) );
  XOR2_X1 U22353 ( .A1(n51057), .A2(n1462), .Z(n11191) );
  XOR2_X1 U22356 ( .A1(n51140), .A2(n51138), .Z(n51057) );
  NOR2_X2 U22358 ( .A1(n58244), .A2(n58033), .ZN(n45750) );
  XOR2_X1 U22359 ( .A1(n58245), .A2(n32493), .Z(n17324) );
  XOR2_X1 U22369 ( .A1(n32632), .A2(n33158), .Z(n58245) );
  NAND2_X2 U22374 ( .A1(n687), .A2(n2357), .ZN(n48885) );
  BUF_X4 U22379 ( .I(n27516), .Z(n30285) );
  AOI22_X2 U22383 ( .A1(n28081), .A2(n2120), .B1(n29826), .B2(n29278), .ZN(
        n58246) );
  XOR2_X1 U22384 ( .A1(n58247), .A2(n24051), .Z(Plaintext[87]) );
  AOI21_X1 U22386 ( .A1(n34554), .A2(n35020), .B(n34553), .ZN(n34561) );
  INV_X2 U22393 ( .I(n24246), .ZN(n39102) );
  XOR2_X1 U22394 ( .A1(n17312), .A2(n57450), .Z(n24246) );
  NAND2_X2 U22396 ( .A1(n11429), .A2(n58248), .ZN(n21944) );
  NOR3_X2 U22417 ( .A1(n18851), .A2(n5040), .A3(n58249), .ZN(n18852) );
  XOR2_X1 U22421 ( .A1(n44387), .A2(n45017), .Z(n60915) );
  XOR2_X1 U22423 ( .A1(n18957), .A2(n7698), .Z(n45017) );
  INV_X2 U22426 ( .I(n6425), .ZN(n44386) );
  OAI21_X2 U22434 ( .A1(n17580), .A2(n40627), .B(n17579), .ZN(n17578) );
  INV_X2 U22447 ( .I(n26088), .ZN(n58252) );
  XOR2_X1 U22457 ( .A1(n37761), .A2(n23199), .Z(n58254) );
  XOR2_X1 U22459 ( .A1(n60606), .A2(n12452), .Z(n16028) );
  XOR2_X1 U22460 ( .A1(n44549), .A2(n2960), .Z(n60606) );
  XOR2_X1 U22462 ( .A1(n58255), .A2(n32760), .Z(n33336) );
  XOR2_X1 U22468 ( .A1(n24255), .A2(n32758), .Z(n58255) );
  INV_X2 U22489 ( .I(n30033), .ZN(n25927) );
  NAND3_X2 U22490 ( .A1(n30029), .A2(n23315), .A3(n28989), .ZN(n30033) );
  NAND2_X2 U22501 ( .A1(n58232), .A2(n25517), .ZN(n6034) );
  XOR2_X1 U22502 ( .A1(n58259), .A2(n23999), .Z(Plaintext[101]) );
  NAND2_X1 U22504 ( .A1(n55174), .A2(n55173), .ZN(n58259) );
  OR2_X1 U22507 ( .A1(n11594), .A2(n58261), .Z(n59661) );
  XOR2_X1 U22508 ( .A1(n38531), .A2(n39260), .Z(n38465) );
  XOR2_X1 U22509 ( .A1(n38645), .A2(n29407), .Z(n38531) );
  NOR3_X1 U22516 ( .A1(n59588), .A2(n56023), .A3(n59587), .ZN(n56025) );
  NOR2_X2 U22521 ( .A1(n23785), .A2(n56708), .ZN(n56704) );
  XOR2_X1 U22524 ( .A1(n58265), .A2(n56714), .Z(Plaintext[166]) );
  NOR2_X1 U22525 ( .A1(n56605), .A2(n56606), .ZN(n56607) );
  NOR2_X2 U22526 ( .A1(n48953), .A2(n62700), .ZN(n49774) );
  NOR2_X1 U22530 ( .A1(n54543), .A2(n58896), .ZN(n54573) );
  BUF_X2 U22534 ( .I(n5481), .Z(n58269) );
  NAND2_X1 U22537 ( .A1(n60059), .A2(n34516), .ZN(n8398) );
  AND2_X2 U22540 ( .A1(n10737), .A2(n7814), .Z(n33004) );
  NAND2_X1 U22545 ( .A1(n7117), .A2(n54406), .ZN(n24004) );
  NOR3_X1 U22549 ( .A1(n40633), .A2(n6891), .A3(n39028), .ZN(n6890) );
  XOR2_X1 U22552 ( .A1(n13947), .A2(n2666), .Z(n15629) );
  NAND2_X2 U22553 ( .A1(n1611), .A2(n6737), .ZN(n11375) );
  NOR2_X2 U22558 ( .A1(n1432), .A2(n22745), .ZN(n30740) );
  XOR2_X1 U22559 ( .A1(n58272), .A2(n17729), .Z(n44064) );
  INV_X2 U22565 ( .I(n58275), .ZN(n12379) );
  XNOR2_X1 U22566 ( .A1(n15788), .A2(n51504), .ZN(n58275) );
  INV_X1 U22567 ( .I(n61549), .ZN(n24561) );
  XOR2_X1 U22573 ( .A1(n58279), .A2(n3139), .Z(n3136) );
  XOR2_X1 U22574 ( .A1(n3140), .A2(n61524), .Z(n58279) );
  NOR2_X1 U22584 ( .A1(n58280), .A2(n51441), .ZN(n59074) );
  NAND2_X1 U22586 ( .A1(n51439), .A2(n51440), .ZN(n58280) );
  OR3_X1 U22589 ( .A1(n555), .A2(n28151), .A3(n28596), .Z(n19625) );
  NAND2_X1 U22596 ( .A1(n6198), .A2(n39903), .ZN(n60985) );
  NAND2_X2 U22598 ( .A1(n35177), .A2(n35176), .ZN(n37555) );
  NOR2_X2 U22601 ( .A1(n19795), .A2(n19796), .ZN(n35173) );
  OAI21_X1 U22627 ( .A1(n49912), .A2(n3394), .B(n58282), .ZN(n49913) );
  OR2_X1 U22635 ( .A1(n49911), .A2(n13839), .Z(n58282) );
  XOR2_X1 U22636 ( .A1(n23534), .A2(n58284), .Z(n44328) );
  XOR2_X1 U22642 ( .A1(n59382), .A2(n44326), .Z(n58284) );
  XOR2_X1 U22669 ( .A1(n58286), .A2(n46528), .Z(n46561) );
  AND2_X1 U22671 ( .A1(n18608), .A2(n50117), .Z(n49891) );
  NAND2_X1 U22673 ( .A1(n41281), .A2(n41282), .ZN(n41283) );
  XOR2_X1 U22682 ( .A1(n8609), .A2(n58289), .Z(n5169) );
  XOR2_X1 U22687 ( .A1(n37562), .A2(n2905), .Z(n38232) );
  XOR2_X1 U22690 ( .A1(n21494), .A2(n38106), .Z(n37562) );
  NAND2_X2 U22699 ( .A1(n8096), .A2(n58290), .ZN(n50138) );
  XOR2_X1 U22702 ( .A1(n1753), .A2(n58293), .Z(n58292) );
  INV_X2 U22706 ( .I(n58294), .ZN(n15318) );
  XOR2_X1 U22719 ( .A1(n8220), .A2(n46637), .Z(n605) );
  NAND3_X1 U22732 ( .A1(n13033), .A2(n13031), .A3(n13032), .ZN(n61578) );
  NAND2_X1 U22735 ( .A1(n58298), .A2(n4323), .ZN(n1100) );
  NOR2_X2 U22736 ( .A1(n19681), .A2(n24788), .ZN(n4323) );
  NAND2_X1 U22745 ( .A1(n53836), .A2(n57317), .ZN(n53837) );
  NOR2_X1 U22746 ( .A1(n53847), .A2(n54072), .ZN(n53836) );
  XOR2_X1 U22755 ( .A1(n50681), .A2(n15459), .Z(n60312) );
  NAND2_X2 U22761 ( .A1(n57735), .A2(n49783), .ZN(n23141) );
  AOI21_X1 U22762 ( .A1(n9089), .A2(n54291), .B(n23122), .ZN(n54297) );
  XOR2_X1 U22788 ( .A1(n18114), .A2(n45402), .Z(n45861) );
  INV_X2 U22791 ( .I(n58302), .ZN(n6530) );
  XOR2_X1 U22793 ( .A1(n44029), .A2(n14461), .Z(n8901) );
  XOR2_X1 U22795 ( .A1(n44892), .A2(n43255), .Z(n44029) );
  NAND2_X1 U22798 ( .A1(n60814), .A2(n16043), .ZN(n60813) );
  NAND2_X2 U22805 ( .A1(n20800), .A2(n64534), .ZN(n34621) );
  NAND2_X2 U22816 ( .A1(n58304), .A2(n18670), .ZN(n15309) );
  INV_X2 U22825 ( .I(n8238), .ZN(n10291) );
  XOR2_X1 U22826 ( .A1(n8238), .A2(n19862), .Z(n19861) );
  AND2_X1 U22828 ( .A1(n63485), .A2(n20844), .Z(n12386) );
  XOR2_X1 U22844 ( .A1(n10927), .A2(n24757), .Z(n17060) );
  NAND2_X2 U22874 ( .A1(n34309), .A2(n23470), .ZN(n32436) );
  XOR2_X1 U22887 ( .A1(n54926), .A2(n63022), .Z(n6622) );
  NOR2_X2 U22890 ( .A1(n54904), .A2(n13671), .ZN(n54926) );
  AOI22_X2 U22895 ( .A1(n37009), .A2(n37011), .B1(n37008), .B2(n24840), .ZN(
        n37014) );
  NAND2_X1 U22896 ( .A1(n1452), .A2(n2037), .ZN(n58312) );
  AND3_X1 U22909 ( .A1(n57277), .A2(n48412), .A3(n12840), .Z(n59715) );
  XOR2_X1 U22922 ( .A1(n8162), .A2(n8161), .Z(n31868) );
  AOI22_X1 U22924 ( .A1(n13723), .A2(n4181), .B1(n4184), .B2(n21706), .ZN(
        n21593) );
  NOR2_X2 U22925 ( .A1(n24007), .A2(n58313), .ZN(n16686) );
  INV_X2 U22932 ( .I(n11475), .ZN(n58313) );
  XOR2_X1 U22937 ( .A1(n58316), .A2(n20446), .Z(n38587) );
  XOR2_X1 U22954 ( .A1(n12129), .A2(n12128), .Z(n58316) );
  INV_X4 U22957 ( .I(n61531), .ZN(n16631) );
  XOR2_X1 U22964 ( .A1(n10826), .A2(n52146), .Z(n22589) );
  NOR3_X2 U22978 ( .A1(n414), .A2(n20676), .A3(n58318), .ZN(n17829) );
  OR2_X1 U22982 ( .A1(n21215), .A2(n16098), .Z(n58318) );
  NOR2_X2 U22983 ( .A1(n24078), .A2(n19206), .ZN(n4571) );
  NAND3_X2 U22999 ( .A1(n59486), .A2(n59485), .A3(n33011), .ZN(n60014) );
  NAND2_X2 U23003 ( .A1(n30526), .A2(n30125), .ZN(n29766) );
  NOR2_X1 U23017 ( .A1(n61969), .A2(n59533), .ZN(n680) );
  NAND3_X2 U23023 ( .A1(n11926), .A2(n42378), .A3(n42379), .ZN(n10798) );
  XOR2_X1 U23038 ( .A1(n58320), .A2(n52348), .Z(n22792) );
  XOR2_X1 U23044 ( .A1(n23239), .A2(n44369), .Z(n41144) );
  OR2_X2 U23045 ( .A1(n54813), .A2(n5141), .Z(n54823) );
  XOR2_X1 U23047 ( .A1(n59209), .A2(n58321), .Z(n5231) );
  XOR2_X1 U23051 ( .A1(n31464), .A2(n31682), .Z(n58321) );
  AND2_X1 U23052 ( .A1(n40993), .A2(n40149), .Z(n59286) );
  NOR2_X2 U23062 ( .A1(n49411), .A2(n49410), .ZN(n47059) );
  XOR2_X1 U23070 ( .A1(n58323), .A2(n39341), .Z(n10778) );
  XOR2_X1 U23071 ( .A1(n10780), .A2(n39342), .Z(n58323) );
  XOR2_X1 U23096 ( .A1(n46550), .A2(n46582), .Z(n21309) );
  NOR2_X1 U23098 ( .A1(n58325), .A2(n21235), .ZN(n52254) );
  INV_X2 U23101 ( .I(n21079), .ZN(n58326) );
  NAND2_X2 U23103 ( .A1(n13567), .A2(n52857), .ZN(n14091) );
  NOR2_X2 U23105 ( .A1(n60590), .A2(n10228), .ZN(n58327) );
  NAND3_X2 U23109 ( .A1(n58328), .A2(n43032), .A3(n43031), .ZN(n43764) );
  NOR3_X1 U23113 ( .A1(n43176), .A2(n40777), .A3(n13678), .ZN(n58635) );
  XOR2_X1 U23119 ( .A1(n32620), .A2(n7773), .Z(n58330) );
  NAND2_X1 U23122 ( .A1(n60746), .A2(n26726), .ZN(n6554) );
  NAND2_X2 U23123 ( .A1(n42486), .A2(n42489), .ZN(n60971) );
  NAND2_X2 U23124 ( .A1(n58332), .A2(n2907), .ZN(n2548) );
  XOR2_X1 U23125 ( .A1(n10645), .A2(n365), .Z(n10650) );
  NAND2_X1 U23132 ( .A1(n57414), .A2(n55404), .ZN(n58333) );
  NAND3_X2 U23140 ( .A1(n54978), .A2(n24075), .A3(n197), .ZN(n55403) );
  NAND2_X2 U23141 ( .A1(n3478), .A2(n21159), .ZN(n61048) );
  NOR2_X2 U23145 ( .A1(n29416), .A2(n1925), .ZN(n1924) );
  XOR2_X1 U23154 ( .A1(n52415), .A2(n20512), .Z(n52417) );
  OR2_X2 U23155 ( .A1(n32461), .A2(n9289), .Z(n4326) );
  NAND3_X1 U23172 ( .A1(n13334), .A2(n13333), .A3(n54432), .ZN(n13332) );
  OR2_X2 U23175 ( .A1(n25333), .A2(n61731), .Z(n34116) );
  XOR2_X1 U23184 ( .A1(n2278), .A2(n14095), .Z(n59868) );
  NOR2_X2 U23186 ( .A1(n40713), .A2(n1516), .ZN(n58367) );
  NAND3_X1 U23195 ( .A1(n18712), .A2(n28269), .A3(n17918), .ZN(n13164) );
  NOR2_X1 U23200 ( .A1(n4373), .A2(n58346), .ZN(n15882) );
  NAND2_X1 U23204 ( .A1(n6894), .A2(n6895), .ZN(n58346) );
  NOR2_X2 U23207 ( .A1(n40100), .A2(n19990), .ZN(n40051) );
  NAND4_X1 U23211 ( .A1(n59700), .A2(n38018), .A3(n25921), .A4(n16962), .ZN(
        n25070) );
  XOR2_X1 U23219 ( .A1(n32238), .A2(n32721), .Z(n31800) );
  XOR2_X1 U23220 ( .A1(n23719), .A2(n56905), .Z(n32238) );
  NAND2_X2 U23227 ( .A1(n23834), .A2(n551), .ZN(n30467) );
  XOR2_X1 U23229 ( .A1(n14697), .A2(n58347), .Z(n17312) );
  XOR2_X1 U23230 ( .A1(n17711), .A2(n17710), .Z(n58347) );
  OR2_X1 U23231 ( .A1(n29456), .A2(n29452), .Z(n28099) );
  NOR2_X1 U23240 ( .A1(n17613), .A2(n45198), .ZN(n17612) );
  NAND2_X1 U23243 ( .A1(n3095), .A2(n57288), .ZN(n61208) );
  INV_X1 U23245 ( .I(n8581), .ZN(n59964) );
  XOR2_X1 U23253 ( .A1(n58355), .A2(n2929), .Z(n23604) );
  XOR2_X1 U23254 ( .A1(n2933), .A2(n61091), .Z(n58355) );
  XOR2_X1 U23260 ( .A1(n58357), .A2(n16508), .Z(n52159) );
  XOR2_X1 U23273 ( .A1(n26025), .A2(n24979), .Z(n26129) );
  XOR2_X1 U23274 ( .A1(n9150), .A2(n1678), .Z(n26025) );
  NOR2_X2 U23293 ( .A1(n50446), .A2(n47761), .ZN(n50235) );
  XOR2_X1 U23301 ( .A1(n52611), .A2(n52610), .Z(n9928) );
  AND3_X1 U23302 ( .A1(n40491), .A2(n40658), .A3(n1404), .Z(n10517) );
  NOR2_X2 U23305 ( .A1(n48560), .A2(n48564), .ZN(n11708) );
  INV_X2 U23308 ( .I(n17891), .ZN(n48560) );
  XOR2_X1 U23322 ( .A1(n51405), .A2(n4156), .Z(n52584) );
  NAND3_X2 U23327 ( .A1(n58365), .A2(n671), .A3(n54453), .ZN(n273) );
  NAND3_X1 U23330 ( .A1(n55023), .A2(n54855), .A3(n54328), .ZN(n58365) );
  NAND2_X2 U23333 ( .A1(n26192), .A2(n609), .ZN(n22514) );
  NAND2_X2 U23335 ( .A1(n58368), .A2(n49954), .ZN(n51628) );
  XOR2_X1 U23337 ( .A1(n59701), .A2(n57358), .Z(n16275) );
  INV_X1 U23347 ( .I(n281), .ZN(n58526) );
  AOI22_X1 U23357 ( .A1(n45509), .A2(n45508), .B1(n45507), .B2(n46075), .ZN(
        n47355) );
  NAND2_X2 U23359 ( .A1(n58371), .A2(n16850), .ZN(n41775) );
  NOR3_X2 U23361 ( .A1(n30282), .A2(n30283), .A3(n30281), .ZN(n58372) );
  OR2_X1 U23368 ( .A1(n30264), .A2(n23317), .Z(n30280) );
  OAI22_X1 U23377 ( .A1(n47581), .A2(n47275), .B1(n2223), .B2(n47579), .ZN(
        n11813) );
  INV_X2 U23379 ( .I(n52888), .ZN(n56987) );
  NAND2_X2 U23380 ( .A1(n52270), .A2(n13920), .ZN(n52888) );
  OR2_X1 U23391 ( .A1(n28676), .A2(n28675), .Z(n12639) );
  XOR2_X1 U23392 ( .A1(n39629), .A2(n20533), .Z(n58378) );
  NAND2_X1 U23393 ( .A1(n19317), .A2(n58379), .ZN(n610) );
  AOI22_X1 U23395 ( .A1(n53298), .A2(n23411), .B1(n16097), .B2(n53300), .ZN(
        n58379) );
  NOR2_X1 U23397 ( .A1(n44784), .A2(n44785), .ZN(n44786) );
  OAI21_X2 U23402 ( .A1(n58382), .A2(n57476), .B(n56206), .ZN(n52723) );
  NAND2_X2 U23410 ( .A1(n43890), .A2(n43242), .ZN(n42858) );
  XOR2_X1 U23415 ( .A1(n58385), .A2(n58384), .Z(n60305) );
  OR4_X1 U23432 ( .A1(n35472), .A2(n35986), .A3(n61180), .A4(n652), .Z(n34898)
         );
  NOR2_X2 U23437 ( .A1(n21409), .A2(n33993), .ZN(n58447) );
  INV_X2 U23438 ( .I(n25920), .ZN(n40100) );
  XOR2_X1 U23440 ( .A1(n17149), .A2(n758), .Z(n25920) );
  INV_X4 U23449 ( .I(n5346), .ZN(n25444) );
  OR2_X1 U23457 ( .A1(n42079), .A2(n42397), .Z(n996) );
  AOI22_X2 U23459 ( .A1(n47227), .A2(n3080), .B1(n59922), .B2(n58009), .ZN(
        n45691) );
  XOR2_X1 U23461 ( .A1(n58392), .A2(n10902), .Z(n45074) );
  INV_X2 U23466 ( .I(n48157), .ZN(n46788) );
  NAND2_X1 U23475 ( .A1(n40055), .A2(n12285), .ZN(n59700) );
  NOR3_X2 U23476 ( .A1(n58393), .A2(n51271), .A3(n51273), .ZN(n51461) );
  AOI21_X1 U23479 ( .A1(n51267), .A2(n51266), .B(n8367), .ZN(n58393) );
  NAND2_X2 U23487 ( .A1(n12848), .A2(n33624), .ZN(n18475) );
  OAI21_X1 U23488 ( .A1(n55902), .A2(n55901), .B(n58394), .ZN(n55904) );
  NAND2_X2 U23490 ( .A1(n58396), .A2(n5156), .ZN(n6744) );
  OAI21_X2 U23509 ( .A1(n52892), .A2(n56605), .B(n22967), .ZN(n58398) );
  NAND3_X2 U23510 ( .A1(n57322), .A2(n35108), .A3(n57263), .ZN(n15275) );
  INV_X2 U23517 ( .I(n44788), .ZN(n13550) );
  INV_X2 U23522 ( .I(n58404), .ZN(n5346) );
  NAND2_X1 U23527 ( .A1(n23980), .A2(n49785), .ZN(n20012) );
  BUF_X4 U23530 ( .I(n62606), .Z(n58975) );
  AND2_X1 U23535 ( .A1(n41769), .A2(n41770), .Z(n58406) );
  INV_X2 U23542 ( .I(n46070), .ZN(n45503) );
  NAND2_X2 U23545 ( .A1(n58313), .A2(n24782), .ZN(n46070) );
  NAND2_X2 U23557 ( .A1(n11477), .A2(n35021), .ZN(n20439) );
  BUF_X4 U23558 ( .I(n19225), .Z(n58710) );
  XOR2_X1 U23559 ( .A1(n58407), .A2(n888), .Z(n25844) );
  XOR2_X1 U23584 ( .A1(n32207), .A2(n13626), .Z(n26062) );
  BUF_X2 U23594 ( .I(n50195), .Z(n51358) );
  NAND2_X2 U23595 ( .A1(n9372), .A2(n7118), .ZN(n58743) );
  NAND3_X2 U23609 ( .A1(n55993), .A2(n55992), .A3(n55991), .ZN(n55994) );
  INV_X1 U23611 ( .I(n35399), .ZN(n36140) );
  NOR2_X2 U23612 ( .A1(n61579), .A2(n24351), .ZN(n35399) );
  NAND2_X1 U23614 ( .A1(n5488), .A2(n38672), .ZN(n38677) );
  NAND3_X1 U23615 ( .A1(n23562), .A2(n58417), .A3(n54862), .ZN(n22148) );
  NAND2_X2 U23616 ( .A1(n6580), .A2(n25758), .ZN(n54862) );
  AND2_X1 U23617 ( .A1(n54460), .A2(n24009), .Z(n58417) );
  NOR2_X1 U23618 ( .A1(n55915), .A2(n55905), .ZN(n58418) );
  XOR2_X1 U23624 ( .A1(n58419), .A2(n60561), .Z(n8733) );
  XOR2_X1 U23625 ( .A1(n46714), .A2(n46706), .Z(n58419) );
  BUF_X2 U23642 ( .I(n15789), .Z(n58420) );
  INV_X1 U23643 ( .I(n31143), .ZN(n58423) );
  XOR2_X1 U23660 ( .A1(n16431), .A2(n16428), .Z(n16757) );
  XOR2_X1 U23661 ( .A1(n58426), .A2(n3575), .Z(n3579) );
  XOR2_X1 U23663 ( .A1(n3578), .A2(n20456), .Z(n58426) );
  INV_X2 U23667 ( .I(n39692), .ZN(n58827) );
  INV_X2 U23670 ( .I(n58427), .ZN(n61659) );
  NOR2_X2 U23675 ( .A1(n13321), .A2(n13322), .ZN(n59018) );
  XOR2_X1 U23677 ( .A1(n58428), .A2(n11961), .Z(n38658) );
  XOR2_X1 U23678 ( .A1(n38656), .A2(n9660), .Z(n58428) );
  XOR2_X1 U23680 ( .A1(n61178), .A2(n58429), .Z(n20579) );
  XOR2_X1 U23684 ( .A1(n63024), .A2(n50927), .Z(n58429) );
  OR2_X1 U23685 ( .A1(n56982), .A2(n56980), .Z(n52276) );
  BUF_X2 U23690 ( .I(n23056), .Z(n58430) );
  NOR2_X2 U23693 ( .A1(n28495), .A2(n1571), .ZN(n26823) );
  NOR2_X2 U23694 ( .A1(n13838), .A2(n1293), .ZN(n12546) );
  XOR2_X1 U23696 ( .A1(n44747), .A2(n9477), .Z(n44045) );
  NAND3_X2 U23697 ( .A1(n1939), .A2(n1936), .A3(n1935), .ZN(n44747) );
  NAND2_X1 U23704 ( .A1(n58575), .A2(n32912), .ZN(n23572) );
  XOR2_X1 U23714 ( .A1(n58431), .A2(n56762), .Z(Plaintext[168]) );
  NAND3_X2 U23721 ( .A1(n14519), .A2(n48468), .A3(n47092), .ZN(n48123) );
  XOR2_X1 U23724 ( .A1(n8774), .A2(n58433), .Z(n58432) );
  INV_X1 U23725 ( .I(n9528), .ZN(n58433) );
  NOR2_X2 U23727 ( .A1(n11912), .A2(n22550), .ZN(n54966) );
  OAI21_X1 U23734 ( .A1(n40232), .A2(n21701), .B(n40231), .ZN(n40235) );
  NOR2_X2 U23738 ( .A1(n9593), .A2(n17775), .ZN(n13699) );
  XOR2_X1 U23741 ( .A1(n38911), .A2(n3950), .Z(n58437) );
  OAI21_X1 U23750 ( .A1(n47042), .A2(n65275), .B(n10333), .ZN(n47044) );
  NOR2_X2 U23760 ( .A1(n59282), .A2(n47501), .ZN(n10333) );
  XOR2_X1 U23766 ( .A1(n20446), .A2(n8629), .Z(n58442) );
  NOR2_X1 U23768 ( .A1(n18425), .A2(n18422), .ZN(n54571) );
  NAND2_X2 U23770 ( .A1(n15724), .A2(n19175), .ZN(n49491) );
  XOR2_X1 U23779 ( .A1(n58446), .A2(n3777), .Z(n5520) );
  NOR2_X1 U23793 ( .A1(n17809), .A2(n17808), .ZN(n59400) );
  NOR2_X2 U23810 ( .A1(n22498), .A2(n7651), .ZN(n28526) );
  NAND2_X1 U23815 ( .A1(n49631), .A2(n60520), .ZN(n49632) );
  NOR2_X2 U23816 ( .A1(n49929), .A2(n49923), .ZN(n60520) );
  NAND2_X2 U23818 ( .A1(n13671), .A2(n22486), .ZN(n22864) );
  NAND2_X1 U23824 ( .A1(n58449), .A2(n40674), .ZN(n22814) );
  NAND3_X1 U23825 ( .A1(n40665), .A2(n40663), .A3(n1404), .ZN(n58449) );
  NOR2_X2 U23828 ( .A1(n56725), .A2(n6954), .ZN(n56677) );
  NAND2_X1 U23844 ( .A1(n58451), .A2(n54861), .ZN(n5217) );
  NAND3_X1 U23850 ( .A1(n54859), .A2(n20740), .A3(n54858), .ZN(n58451) );
  BUF_X2 U23861 ( .I(n11005), .Z(n1248) );
  OR3_X2 U23862 ( .A1(n26565), .A2(n57872), .A3(n61317), .Z(n27020) );
  NOR2_X2 U23863 ( .A1(n7127), .A2(n1865), .ZN(n30029) );
  NAND3_X2 U23865 ( .A1(n41982), .A2(n22999), .A3(n64663), .ZN(n41615) );
  NOR2_X2 U23866 ( .A1(n40896), .A2(n40897), .ZN(n41987) );
  INV_X2 U23879 ( .I(n13054), .ZN(n58453) );
  XOR2_X1 U23886 ( .A1(n58456), .A2(n31734), .Z(n31743) );
  NOR2_X2 U23887 ( .A1(n4515), .A2(n20445), .ZN(n19507) );
  NOR2_X2 U23888 ( .A1(n34611), .A2(n34610), .ZN(n4628) );
  NOR2_X2 U23889 ( .A1(n34041), .A2(n33420), .ZN(n34611) );
  OR2_X2 U23895 ( .A1(n34035), .A2(n34606), .Z(n20443) );
  XOR2_X1 U23896 ( .A1(n9780), .A2(n19771), .Z(n19770) );
  AOI21_X2 U23911 ( .A1(n58655), .A2(n5175), .B(n58460), .ZN(n5173) );
  OAI21_X1 U23917 ( .A1(n56186), .A2(n1590), .B(n56176), .ZN(n56152) );
  NAND2_X1 U23919 ( .A1(n56174), .A2(n11716), .ZN(n56186) );
  XOR2_X1 U23923 ( .A1(n38870), .A2(n39466), .Z(n25885) );
  NAND2_X1 U23925 ( .A1(n56916), .A2(n56958), .ZN(n59736) );
  NOR2_X2 U23926 ( .A1(n6359), .A2(n8475), .ZN(n13054) );
  NAND2_X2 U23932 ( .A1(n5551), .A2(n52223), .ZN(n5553) );
  XOR2_X1 U23933 ( .A1(n58462), .A2(n32241), .Z(n61130) );
  OAI22_X1 U23939 ( .A1(n27917), .A2(n27918), .B1(n28786), .B2(n22164), .ZN(
        n27919) );
  XOR2_X1 U23945 ( .A1(n2748), .A2(n2540), .Z(n46272) );
  BUF_X2 U23946 ( .I(n23646), .Z(n58463) );
  NAND3_X2 U23959 ( .A1(n14501), .A2(n54446), .A3(n60751), .ZN(n54688) );
  INV_X2 U23961 ( .I(n58466), .ZN(n26539) );
  NAND2_X2 U23964 ( .A1(n15715), .A2(n58420), .ZN(n58466) );
  XOR2_X1 U23969 ( .A1(n6140), .A2(n1461), .Z(n52372) );
  XOR2_X1 U23975 ( .A1(n24276), .A2(n52354), .Z(n38943) );
  NOR2_X2 U23979 ( .A1(n3756), .A2(n1307), .ZN(n40064) );
  NOR2_X2 U23982 ( .A1(n34186), .A2(n34594), .ZN(n33966) );
  XOR2_X1 U23984 ( .A1(n14880), .A2(n50634), .Z(n2724) );
  NAND3_X2 U23989 ( .A1(n22985), .A2(n25551), .A3(n25550), .ZN(n14880) );
  NOR2_X2 U23997 ( .A1(n14333), .A2(n23796), .ZN(n59020) );
  XOR2_X1 U23998 ( .A1(n58470), .A2(n15430), .Z(n19049) );
  XOR2_X1 U23999 ( .A1(n51317), .A2(n50707), .Z(n58470) );
  NAND3_X2 U24009 ( .A1(n5611), .A2(n5610), .A3(n5609), .ZN(n17892) );
  BUF_X2 U24012 ( .I(n34993), .Z(n58472) );
  XOR2_X1 U24018 ( .A1(n19273), .A2(n38509), .Z(n58473) );
  XOR2_X1 U24028 ( .A1(n58474), .A2(n56827), .Z(Plaintext[174]) );
  INV_X1 U24033 ( .I(n10762), .ZN(n58475) );
  OAI21_X2 U24048 ( .A1(n18009), .A2(n18008), .B(n23526), .ZN(n56452) );
  OAI21_X2 U24049 ( .A1(n60639), .A2(n20501), .B(n36976), .ZN(n20502) );
  OAI21_X2 U24054 ( .A1(n15902), .A2(n58476), .B(n56660), .ZN(n17348) );
  NOR2_X2 U24055 ( .A1(n56372), .A2(n58477), .ZN(n58476) );
  INV_X2 U24057 ( .I(n56362), .ZN(n58477) );
  NAND2_X2 U24062 ( .A1(n7057), .A2(n17930), .ZN(n39922) );
  NAND2_X2 U24063 ( .A1(n57208), .A2(n10554), .ZN(n40061) );
  XOR2_X1 U24068 ( .A1(n38206), .A2(n23120), .Z(n58479) );
  OR2_X1 U24088 ( .A1(n50345), .A2(n50348), .Z(n59369) );
  AND2_X1 U24090 ( .A1(n29662), .A2(n29663), .Z(n28191) );
  OR2_X2 U24113 ( .A1(n52281), .A2(n59294), .Z(n56368) );
  AOI22_X1 U24122 ( .A1(n16824), .A2(n58484), .B1(n16823), .B2(n41053), .ZN(
        n20643) );
  XOR2_X1 U24129 ( .A1(n9018), .A2(Ciphertext[11]), .Z(n58485) );
  OR2_X1 U24131 ( .A1(n36483), .A2(n24028), .Z(n943) );
  AOI22_X1 U24139 ( .A1(n29257), .A2(n29256), .B1(n62414), .B2(n29255), .ZN(
        n29258) );
  NOR2_X2 U24144 ( .A1(n1556), .A2(n29779), .ZN(n29256) );
  XOR2_X1 U24145 ( .A1(n16835), .A2(n58488), .Z(n19006) );
  XOR2_X1 U24146 ( .A1(n31966), .A2(n16833), .Z(n58488) );
  XOR2_X1 U24149 ( .A1(n5694), .A2(n18091), .Z(n5693) );
  NAND2_X2 U24160 ( .A1(n58663), .A2(n56597), .ZN(n56689) );
  BUF_X2 U24168 ( .I(n23941), .Z(n58490) );
  NOR2_X2 U24173 ( .A1(n14561), .A2(n22570), .ZN(n46968) );
  NOR2_X2 U24177 ( .A1(n6987), .A2(n60560), .ZN(n60145) );
  XOR2_X1 U24184 ( .A1(n13286), .A2(n55139), .Z(n50581) );
  NAND2_X2 U24185 ( .A1(n23640), .A2(n50147), .ZN(n13286) );
  XOR2_X1 U24200 ( .A1(n63008), .A2(n20446), .Z(n38718) );
  OAI22_X1 U24220 ( .A1(n55167), .A2(n55166), .B1(n21389), .B2(n55168), .ZN(
        n55169) );
  XOR2_X1 U24224 ( .A1(n4281), .A2(n5818), .Z(n31913) );
  NOR2_X2 U24226 ( .A1(n273), .A2(n18246), .ZN(n60149) );
  NAND2_X2 U24232 ( .A1(n11704), .A2(n23890), .ZN(n39505) );
  AND2_X1 U24233 ( .A1(n6229), .A2(n15267), .Z(n58498) );
  NAND2_X2 U24249 ( .A1(n42338), .A2(n42724), .ZN(n42721) );
  INV_X2 U24252 ( .I(n58502), .ZN(n875) );
  NAND2_X2 U24254 ( .A1(n13163), .A2(n18306), .ZN(n58502) );
  NAND3_X2 U24261 ( .A1(n32811), .A2(n32810), .A3(n32812), .ZN(n58503) );
  NAND2_X2 U24262 ( .A1(n63012), .A2(n56084), .ZN(n56091) );
  XOR2_X1 U24263 ( .A1(n58505), .A2(n19723), .Z(n24548) );
  XOR2_X1 U24271 ( .A1(n11528), .A2(n31748), .Z(n58505) );
  NAND2_X2 U24276 ( .A1(n6928), .A2(n58506), .ZN(n18715) );
  NAND2_X1 U24289 ( .A1(n52938), .A2(n52937), .ZN(n58534) );
  NAND2_X1 U24301 ( .A1(n56546), .A2(n52706), .ZN(n58511) );
  NOR2_X2 U24302 ( .A1(n22870), .A2(n52701), .ZN(n56546) );
  XOR2_X1 U24315 ( .A1(n58517), .A2(n32594), .Z(n9991) );
  NAND3_X1 U24323 ( .A1(n46265), .A2(n46267), .A3(n47502), .ZN(n9934) );
  NOR2_X2 U24324 ( .A1(n2180), .A2(n55476), .ZN(n55478) );
  NOR2_X2 U24330 ( .A1(n24375), .A2(n24486), .ZN(n24405) );
  XOR2_X1 U24331 ( .A1(n52155), .A2(n59463), .Z(n18466) );
  NAND2_X2 U24332 ( .A1(n58519), .A2(n58518), .ZN(n37158) );
  INV_X2 U24342 ( .I(n25994), .ZN(n37212) );
  NOR3_X2 U24349 ( .A1(n28892), .A2(n28891), .A3(n28890), .ZN(n58522) );
  INV_X2 U24357 ( .I(n58524), .ZN(n32940) );
  XOR2_X1 U24362 ( .A1(n58525), .A2(n8795), .Z(n1048) );
  XOR2_X1 U24363 ( .A1(n46135), .A2(n57373), .Z(n58525) );
  XOR2_X1 U24366 ( .A1(n13778), .A2(n10793), .Z(n10792) );
  XOR2_X1 U24372 ( .A1(n24178), .A2(n61152), .Z(n6250) );
  NAND2_X2 U24380 ( .A1(n4783), .A2(n54951), .ZN(n54614) );
  NAND2_X1 U24384 ( .A1(n18722), .A2(n57261), .ZN(n18721) );
  NAND3_X2 U24386 ( .A1(n8163), .A2(n4240), .A3(n4238), .ZN(n13330) );
  INV_X2 U24388 ( .I(n40128), .ZN(n60860) );
  NAND2_X2 U24389 ( .A1(n19102), .A2(n42488), .ZN(n40128) );
  NAND2_X2 U24394 ( .A1(n42800), .A2(n42799), .ZN(n45041) );
  NAND2_X2 U24396 ( .A1(n59553), .A2(n9524), .ZN(n8997) );
  INV_X2 U24397 ( .I(n32940), .ZN(n36574) );
  NOR2_X2 U24400 ( .A1(n7891), .A2(n58535), .ZN(n23936) );
  NAND4_X2 U24402 ( .A1(n57383), .A2(n7896), .A3(n60921), .A4(n52397), .ZN(
        n58535) );
  XOR2_X1 U24413 ( .A1(n63005), .A2(n14373), .Z(n17231) );
  NOR3_X2 U24414 ( .A1(n58538), .A2(n6638), .A3(n42537), .ZN(n3005) );
  XOR2_X1 U24416 ( .A1(n37583), .A2(n6302), .Z(n37802) );
  NOR2_X1 U24422 ( .A1(n6842), .A2(n1341), .ZN(n58544) );
  NOR2_X2 U24429 ( .A1(n14312), .A2(n27508), .ZN(n26974) );
  XOR2_X1 U24433 ( .A1(n1198), .A2(n10745), .Z(n6756) );
  NAND2_X2 U24435 ( .A1(n28852), .A2(n28162), .ZN(n28157) );
  XOR2_X1 U24457 ( .A1(n7663), .A2(n58549), .Z(n32051) );
  XOR2_X1 U24459 ( .A1(n12123), .A2(n32049), .Z(n58549) );
  NAND2_X2 U24464 ( .A1(n17972), .A2(n29633), .ZN(n25014) );
  NAND2_X1 U24465 ( .A1(n19730), .A2(n19729), .ZN(n60257) );
  NAND2_X2 U24469 ( .A1(n17492), .A2(n34849), .ZN(n5073) );
  NOR2_X1 U24474 ( .A1(n30238), .A2(n29208), .ZN(n18238) );
  NAND3_X1 U24475 ( .A1(n59916), .A2(n35150), .A3(n35149), .ZN(n16639) );
  NOR2_X2 U24476 ( .A1(n4647), .A2(n49410), .ZN(n58550) );
  NOR4_X2 U24497 ( .A1(n5305), .A2(n5303), .A3(n5304), .A4(n11385), .ZN(n5045)
         );
  NOR2_X2 U24502 ( .A1(n43979), .A2(n1719), .ZN(n5571) );
  NAND3_X1 U24506 ( .A1(n15244), .A2(n55975), .A3(n55976), .ZN(n55977) );
  NOR2_X1 U24507 ( .A1(n58555), .A2(n7802), .ZN(n7803) );
  XOR2_X1 U24518 ( .A1(n61010), .A2(n46507), .Z(n46681) );
  NAND3_X2 U24519 ( .A1(n58637), .A2(n23454), .A3(n55459), .ZN(n25636) );
  NAND2_X2 U24520 ( .A1(n28989), .A2(n29726), .ZN(n29731) );
  OAI22_X1 U24529 ( .A1(n12248), .A2(n35287), .B1(n24983), .B2(n904), .ZN(
        n58562) );
  OAI21_X1 U24533 ( .A1(n34689), .A2(n34688), .B(n34687), .ZN(n58563) );
  NAND3_X2 U24542 ( .A1(n15886), .A2(n594), .A3(n20014), .ZN(n20892) );
  OAI21_X1 U24547 ( .A1(n58567), .A2(n55632), .B(n23520), .ZN(n23519) );
  NAND2_X1 U24548 ( .A1(n55626), .A2(n55628), .ZN(n58567) );
  OAI21_X1 U24554 ( .A1(n59947), .A2(n59946), .B(n59945), .ZN(n41777) );
  AOI21_X1 U24563 ( .A1(n42100), .A2(n41717), .B(n16139), .ZN(n3657) );
  BUF_X4 U24564 ( .I(n53462), .Z(n53493) );
  NOR2_X2 U24567 ( .A1(n54278), .A2(n58568), .ZN(n23756) );
  OR2_X2 U24575 ( .A1(n5271), .A2(n22739), .Z(n14306) );
  XOR2_X1 U24578 ( .A1(n20429), .A2(n5913), .Z(n50493) );
  XOR2_X1 U24582 ( .A1(n51522), .A2(n50204), .Z(n20429) );
  XOR2_X1 U24595 ( .A1(n44045), .A2(n12507), .Z(n44154) );
  OR2_X1 U24599 ( .A1(n55966), .A2(n23900), .Z(n24464) );
  XOR2_X1 U24601 ( .A1(n58570), .A2(n51616), .Z(n18444) );
  XOR2_X1 U24607 ( .A1(n51615), .A2(n18446), .Z(n58570) );
  XOR2_X1 U24608 ( .A1(n58571), .A2(n9244), .Z(n61236) );
  XOR2_X1 U24609 ( .A1(n9246), .A2(n14675), .Z(n58571) );
  NAND2_X2 U24611 ( .A1(n14165), .A2(n39007), .ZN(n41402) );
  XOR2_X1 U24620 ( .A1(n21826), .A2(n38968), .Z(n13060) );
  XOR2_X1 U24621 ( .A1(n22487), .A2(n17583), .Z(n38968) );
  NAND2_X1 U24632 ( .A1(n28583), .A2(n5267), .ZN(n5760) );
  NAND2_X2 U24635 ( .A1(n24504), .A2(n29472), .ZN(n28583) );
  NAND3_X1 U24636 ( .A1(n32956), .A2(n60960), .A3(n61748), .ZN(n32961) );
  AND2_X1 U24644 ( .A1(n14369), .A2(n48600), .Z(n60939) );
  NAND2_X1 U24648 ( .A1(n58577), .A2(n10138), .ZN(n10942) );
  OR3_X1 U24649 ( .A1(n34560), .A2(n20785), .A3(n17368), .Z(n58577) );
  NOR2_X2 U24658 ( .A1(n24571), .A2(n15545), .ZN(n33583) );
  NAND3_X2 U24661 ( .A1(n37140), .A2(n37141), .A3(n37139), .ZN(n21239) );
  AND2_X1 U24666 ( .A1(n28797), .A2(n17824), .Z(n9719) );
  XOR2_X1 U24667 ( .A1(n4871), .A2(n14626), .Z(n60854) );
  XOR2_X1 U24670 ( .A1(n44970), .A2(n25612), .Z(n14626) );
  OR2_X1 U24673 ( .A1(n2026), .A2(n23407), .Z(n44563) );
  NAND3_X1 U24676 ( .A1(n18143), .A2(n41749), .A3(n63212), .ZN(n41751) );
  NOR2_X2 U24677 ( .A1(n43447), .A2(n43438), .ZN(n18143) );
  NAND2_X2 U24678 ( .A1(n11769), .A2(n58581), .ZN(n14174) );
  NOR3_X2 U24681 ( .A1(n27434), .A2(n14176), .A3(n14177), .ZN(n58581) );
  XOR2_X1 U24682 ( .A1(n39756), .A2(n58582), .Z(n14508) );
  XOR2_X1 U24686 ( .A1(n39653), .A2(n58585), .Z(n39656) );
  XOR2_X1 U24688 ( .A1(n19008), .A2(n39652), .Z(n58585) );
  INV_X2 U24690 ( .I(n11034), .ZN(n11035) );
  XOR2_X1 U24695 ( .A1(n5676), .A2(n59866), .Z(n58586) );
  NOR2_X2 U24698 ( .A1(n50220), .A2(n50218), .ZN(n3303) );
  NAND3_X2 U24705 ( .A1(n3221), .A2(n3219), .A3(n48180), .ZN(n5204) );
  NAND2_X2 U24711 ( .A1(n24418), .A2(n6330), .ZN(n555) );
  NOR3_X2 U24713 ( .A1(n57434), .A2(n36805), .A3(n15946), .ZN(n58589) );
  NOR2_X2 U24726 ( .A1(n17715), .A2(n17713), .ZN(n24839) );
  NOR2_X1 U24728 ( .A1(n40280), .A2(n40281), .ZN(n40286) );
  INV_X1 U24740 ( .I(n58888), .ZN(n35383) );
  NAND2_X2 U24751 ( .A1(n36536), .A2(n60014), .ZN(n58888) );
  BUF_X4 U24752 ( .I(n23956), .Z(n518) );
  AOI22_X1 U24756 ( .A1(n54762), .A2(n54761), .B1(n54763), .B2(n54764), .ZN(
        n54773) );
  NAND3_X1 U24788 ( .A1(n50334), .A2(n60467), .A3(n21052), .ZN(n7527) );
  XOR2_X1 U24799 ( .A1(n31600), .A2(n58603), .Z(n6309) );
  XOR2_X1 U24810 ( .A1(n31599), .A2(n24008), .Z(n58603) );
  NOR2_X1 U24812 ( .A1(n29676), .A2(n29677), .ZN(n29678) );
  NAND2_X1 U24814 ( .A1(n54591), .A2(n54592), .ZN(n59506) );
  XOR2_X1 U24825 ( .A1(n58608), .A2(n5037), .Z(n14595) );
  XOR2_X1 U24828 ( .A1(n58609), .A2(n45860), .Z(n630) );
  XOR2_X1 U24832 ( .A1(n44338), .A2(n4732), .Z(n58609) );
  NOR2_X2 U24839 ( .A1(n2483), .A2(n35096), .ZN(n37048) );
  NAND3_X1 U24840 ( .A1(n58610), .A2(n26514), .A3(n3117), .ZN(n26516) );
  NAND2_X1 U24844 ( .A1(n11076), .A2(n28418), .ZN(n58610) );
  NAND4_X2 U24866 ( .A1(n12357), .A2(n35135), .A3(n58615), .A4(n35136), .ZN(
        n23922) );
  NOR2_X2 U24871 ( .A1(n59388), .A2(n58616), .ZN(n6230) );
  OR2_X1 U24875 ( .A1(n6084), .A2(n6085), .Z(n58616) );
  INV_X4 U24891 ( .I(n41132), .ZN(n1742) );
  XOR2_X1 U24898 ( .A1(n6145), .A2(n1751), .Z(n4928) );
  NAND2_X1 U24903 ( .A1(n17879), .A2(n27329), .ZN(n17878) );
  XOR2_X1 U24916 ( .A1(n46383), .A2(n46384), .Z(n58617) );
  XOR2_X1 U24921 ( .A1(n2881), .A2(n58619), .Z(n58618) );
  NOR2_X2 U24925 ( .A1(n60759), .A2(n24963), .ZN(n24962) );
  BUF_X2 U24932 ( .I(n14518), .Z(n58620) );
  BUF_X2 U24933 ( .I(n31242), .Z(n58621) );
  OR2_X1 U24935 ( .A1(n4097), .A2(n60808), .Z(n32789) );
  XNOR2_X1 U24949 ( .A1(n6722), .A2(n4901), .ZN(n58969) );
  NAND2_X2 U24955 ( .A1(n58624), .A2(n33417), .ZN(n31537) );
  AOI21_X2 U24957 ( .A1(n31528), .A2(n34615), .B(n18935), .ZN(n58624) );
  NAND2_X2 U24967 ( .A1(n55590), .A2(n55569), .ZN(n55596) );
  XOR2_X1 U24970 ( .A1(n57405), .A2(n58625), .Z(n3575) );
  XOR2_X1 U24973 ( .A1(n33154), .A2(n61883), .Z(n58625) );
  OR2_X2 U24985 ( .A1(n17536), .A2(n60822), .Z(n1704) );
  NAND2_X1 U24986 ( .A1(n54963), .A2(n61736), .ZN(n54975) );
  NOR2_X2 U24989 ( .A1(n54487), .A2(n11912), .ZN(n54963) );
  XOR2_X1 U25003 ( .A1(n38530), .A2(n23280), .Z(n37988) );
  AND2_X1 U25005 ( .A1(n25220), .A2(n54960), .Z(n59320) );
  OR2_X2 U25009 ( .A1(n16858), .A2(n29576), .Z(n2806) );
  AND2_X1 U25011 ( .A1(n6330), .A2(n21021), .Z(n29644) );
  XOR2_X1 U25012 ( .A1(n58628), .A2(n1677), .Z(n44020) );
  XOR2_X1 U25021 ( .A1(n44017), .A2(n44018), .Z(n58628) );
  INV_X4 U25024 ( .I(n31055), .ZN(n60111) );
  NOR2_X2 U25029 ( .A1(n60010), .A2(n29640), .ZN(n31155) );
  NAND3_X2 U25030 ( .A1(n41215), .A2(n61316), .A3(n38935), .ZN(n40769) );
  NAND2_X2 U25033 ( .A1(n6852), .A2(n20652), .ZN(n41215) );
  NAND2_X1 U25043 ( .A1(n29015), .A2(n9197), .ZN(n29018) );
  NAND2_X2 U25044 ( .A1(n1318), .A2(n23370), .ZN(n29015) );
  NOR2_X2 U25055 ( .A1(n26004), .A2(n59259), .ZN(n15209) );
  INV_X1 U25056 ( .I(n7797), .ZN(n34571) );
  NAND2_X2 U25063 ( .A1(n57166), .A2(n7797), .ZN(n11423) );
  NAND2_X2 U25064 ( .A1(n1428), .A2(n12480), .ZN(n7797) );
  INV_X2 U25068 ( .I(n40832), .ZN(n39945) );
  NAND2_X2 U25071 ( .A1(n24716), .A2(n58633), .ZN(n23600) );
  NOR4_X2 U25072 ( .A1(n24719), .A2(n24720), .A3(n2019), .A4(n36341), .ZN(
        n58633) );
  XOR2_X1 U25073 ( .A1(n51605), .A2(n58634), .Z(n25805) );
  XOR2_X1 U25074 ( .A1(n19847), .A2(n52335), .Z(n58634) );
  NAND2_X1 U25075 ( .A1(n12167), .A2(n63123), .ZN(n12166) );
  AND2_X1 U25081 ( .A1(n6317), .A2(n31270), .Z(n59760) );
  AND2_X1 U25082 ( .A1(n55458), .A2(n55457), .Z(n58637) );
  NOR2_X1 U25083 ( .A1(n41470), .A2(n64655), .ZN(n40765) );
  OR2_X1 U25096 ( .A1(n46984), .A2(n46983), .Z(n58639) );
  XNOR2_X1 U25098 ( .A1(n16935), .A2(n30922), .ZN(n59172) );
  XOR2_X1 U25099 ( .A1(n58640), .A2(n50166), .Z(n18702) );
  XOR2_X1 U25102 ( .A1(n10497), .A2(n50105), .Z(n58640) );
  XOR2_X1 U25103 ( .A1(n19407), .A2(n58531), .Z(n31871) );
  XOR2_X1 U25113 ( .A1(n33905), .A2(n18295), .Z(n19407) );
  XOR2_X1 U25119 ( .A1(n15401), .A2(n11074), .Z(n44549) );
  INV_X2 U25121 ( .I(n58641), .ZN(n26431) );
  XNOR2_X1 U25124 ( .A1(Key[24]), .A2(Ciphertext[101]), .ZN(n58641) );
  NAND3_X2 U25129 ( .A1(n59289), .A2(n41535), .A3(n41536), .ZN(n24450) );
  NAND2_X2 U25153 ( .A1(n24250), .A2(n58874), .ZN(n5104) );
  NAND4_X2 U25170 ( .A1(n12570), .A2(n12571), .A3(n25784), .A4(n35449), .ZN(
        n4903) );
  BUF_X2 U25179 ( .I(n19701), .Z(n58644) );
  INV_X2 U25182 ( .I(n42170), .ZN(n58646) );
  NOR2_X2 U25183 ( .A1(n41779), .A2(n4945), .ZN(n42170) );
  OR2_X1 U25189 ( .A1(n8400), .A2(n8402), .Z(n58647) );
  INV_X1 U25191 ( .I(n36141), .ZN(n60292) );
  BUF_X2 U25195 ( .I(n16766), .Z(n58648) );
  NAND2_X2 U25196 ( .A1(n22657), .A2(n61388), .ZN(n58874) );
  NAND3_X2 U25198 ( .A1(n58649), .A2(n48904), .A3(n49536), .ZN(n12220) );
  OAI21_X2 U25199 ( .A1(n16408), .A2(n49540), .B(n47917), .ZN(n58649) );
  NOR2_X2 U25204 ( .A1(n3055), .A2(n4734), .ZN(n58913) );
  BUF_X4 U25215 ( .I(n48586), .Z(n23542) );
  NOR3_X2 U25217 ( .A1(n13164), .A2(n4799), .A3(n13203), .ZN(n13204) );
  OAI21_X1 U25218 ( .A1(n4821), .A2(n4822), .B(n28258), .ZN(n18712) );
  NOR3_X2 U25220 ( .A1(n8740), .A2(n8739), .A3(n50315), .ZN(n8738) );
  XOR2_X1 U25225 ( .A1(n46611), .A2(n19994), .Z(n44856) );
  XOR2_X1 U25226 ( .A1(n604), .A2(n26046), .Z(n59679) );
  INV_X2 U25231 ( .I(n15808), .ZN(n58651) );
  NAND2_X2 U25246 ( .A1(n54189), .A2(n54197), .ZN(n54172) );
  NAND3_X2 U25252 ( .A1(n7060), .A2(n7059), .A3(n7061), .ZN(n15507) );
  NAND3_X1 U25253 ( .A1(n20045), .A2(n1615), .A3(n101), .ZN(n17028) );
  XOR2_X1 U25263 ( .A1(n38708), .A2(n38648), .Z(n39716) );
  NOR2_X2 U25264 ( .A1(n61267), .A2(n35540), .ZN(n38648) );
  NAND2_X2 U25266 ( .A1(n40670), .A2(n40663), .ZN(n10133) );
  INV_X1 U25267 ( .I(n48376), .ZN(n59956) );
  OR2_X1 U25271 ( .A1(n26665), .A2(n27573), .Z(n457) );
  OR2_X1 U25280 ( .A1(n15279), .A2(n15278), .Z(n14991) );
  XOR2_X1 U25282 ( .A1(n4453), .A2(n21101), .Z(n47290) );
  AOI21_X2 U25291 ( .A1(n58654), .A2(n27530), .B(n58653), .ZN(n17416) );
  NAND2_X2 U25296 ( .A1(n26053), .A2(n26595), .ZN(n58653) );
  NAND3_X2 U25298 ( .A1(n20974), .A2(n23698), .A3(n17915), .ZN(n39514) );
  BUF_X2 U25303 ( .I(n23646), .Z(n8194) );
  NAND3_X2 U25313 ( .A1(n60772), .A2(n49921), .A3(n24692), .ZN(n9240) );
  NAND2_X2 U25314 ( .A1(n25026), .A2(n3733), .ZN(n47875) );
  NAND2_X2 U25317 ( .A1(n47876), .A2(n7579), .ZN(n25026) );
  NAND3_X1 U25319 ( .A1(n55880), .A2(n60203), .A3(n19307), .ZN(n55845) );
  NOR2_X1 U25355 ( .A1(n6984), .A2(n37410), .ZN(n35922) );
  NOR2_X2 U25369 ( .A1(n14770), .A2(n14768), .ZN(n18599) );
  XOR2_X1 U25373 ( .A1(n17898), .A2(n64512), .Z(n58660) );
  XOR2_X1 U25380 ( .A1(n51102), .A2(n58661), .Z(n10749) );
  NAND2_X1 U25381 ( .A1(n37412), .A2(n37413), .ZN(n37414) );
  XOR2_X1 U25397 ( .A1(n10725), .A2(n10722), .Z(n51962) );
  NOR3_X2 U25414 ( .A1(n7277), .A2(n15981), .A3(n19521), .ZN(n58663) );
  NAND3_X2 U25420 ( .A1(n34654), .A2(n34663), .A3(n34656), .ZN(n58664) );
  AND2_X1 U25425 ( .A1(n61578), .A2(n30741), .Z(n59140) );
  NAND2_X1 U25426 ( .A1(n58665), .A2(n23097), .ZN(n56682) );
  OAI21_X1 U25427 ( .A1(n8616), .A2(n8617), .B(n56703), .ZN(n58665) );
  INV_X2 U25430 ( .I(n19379), .ZN(n3707) );
  NAND2_X2 U25431 ( .A1(n19489), .A2(n49923), .ZN(n19379) );
  NOR2_X1 U25432 ( .A1(n11388), .A2(n30488), .ZN(n60958) );
  INV_X4 U25438 ( .I(n36052), .ZN(n36775) );
  AOI22_X2 U25444 ( .A1(n38344), .A2(n7571), .B1(n15894), .B2(n37593), .ZN(
        n58669) );
  NAND3_X2 U25450 ( .A1(n40150), .A2(n18706), .A3(n58364), .ZN(n3466) );
  NAND2_X2 U25457 ( .A1(n60957), .A2(n60652), .ZN(n58672) );
  NAND3_X2 U25461 ( .A1(n58674), .A2(n6968), .A3(n23602), .ZN(n46165) );
  NOR2_X2 U25467 ( .A1(n12737), .A2(n33675), .ZN(n22942) );
  XOR2_X1 U25468 ( .A1(n46309), .A2(n46308), .Z(n46310) );
  XOR2_X1 U25487 ( .A1(n58745), .A2(n57438), .Z(n59064) );
  XOR2_X1 U25499 ( .A1(n1346), .A2(n24672), .Z(n32321) );
  XOR2_X1 U25508 ( .A1(n21944), .A2(n15816), .Z(n9288) );
  NOR2_X2 U25510 ( .A1(n10951), .A2(n27919), .ZN(n15816) );
  OAI21_X1 U25520 ( .A1(n1927), .A2(n16869), .B(n34073), .ZN(n33485) );
  XOR2_X1 U25527 ( .A1(n26090), .A2(n51362), .Z(n58916) );
  NOR3_X2 U25537 ( .A1(n58680), .A2(n11415), .A3(n12214), .ZN(n58691) );
  NOR2_X2 U25539 ( .A1(n49274), .A2(n4436), .ZN(n58680) );
  XOR2_X1 U25543 ( .A1(n23330), .A2(n24151), .Z(n37726) );
  OR2_X1 U25562 ( .A1(n35666), .A2(n35667), .Z(n58684) );
  NAND3_X2 U25572 ( .A1(n58685), .A2(n1015), .A3(n41585), .ZN(n41587) );
  NAND2_X1 U25574 ( .A1(n41582), .A2(n41581), .ZN(n58685) );
  INV_X4 U25576 ( .I(n33540), .ZN(n33539) );
  XOR2_X1 U25580 ( .A1(n50992), .A2(n58689), .Z(n50686) );
  XOR2_X1 U25581 ( .A1(n724), .A2(n49088), .Z(n58689) );
  XOR2_X1 U25582 ( .A1(n44912), .A2(n46446), .Z(n16599) );
  NAND3_X2 U25592 ( .A1(n32778), .A2(n32779), .A3(n32777), .ZN(n39391) );
  XOR2_X1 U25608 ( .A1(n5664), .A2(n5663), .Z(n5662) );
  XOR2_X1 U25612 ( .A1(n39293), .A2(n39292), .Z(n39305) );
  XOR2_X1 U25614 ( .A1(n18539), .A2(n18540), .Z(n39292) );
  NOR2_X2 U25618 ( .A1(n8589), .A2(n22084), .ZN(n11747) );
  NAND2_X2 U25631 ( .A1(n8028), .A2(n1398), .ZN(n41322) );
  AOI21_X1 U25632 ( .A1(n42852), .A2(n59412), .B(n42850), .ZN(n42853) );
  XOR2_X1 U25635 ( .A1(n2289), .A2(n60959), .Z(n17731) );
  AND2_X1 U25637 ( .A1(n21840), .A2(n25310), .Z(n5072) );
  XOR2_X1 U25661 ( .A1(n63030), .A2(n8148), .Z(n58694) );
  NAND4_X2 U25663 ( .A1(n34792), .A2(n34793), .A3(n35013), .A4(n35005), .ZN(
        n9768) );
  NAND2_X2 U25664 ( .A1(n34791), .A2(n33468), .ZN(n35005) );
  BUF_X4 U25673 ( .I(n54570), .Z(n18422) );
  NAND2_X2 U25677 ( .A1(n47244), .A2(n59059), .ZN(n45990) );
  XOR2_X1 U25679 ( .A1(n58695), .A2(n38908), .Z(n3713) );
  XOR2_X1 U25684 ( .A1(n24169), .A2(n14228), .Z(n58695) );
  BUF_X2 U25699 ( .I(n1192), .Z(n58696) );
  AND2_X2 U25701 ( .A1(n1388), .A2(n45766), .Z(n45762) );
  NAND2_X2 U25709 ( .A1(n26095), .A2(n2199), .ZN(n54943) );
  NAND2_X2 U25714 ( .A1(n9012), .A2(n2033), .ZN(n16869) );
  INV_X2 U25725 ( .I(n30895), .ZN(n58700) );
  XOR2_X1 U25730 ( .A1(n39646), .A2(n23853), .Z(n7853) );
  NAND2_X2 U25734 ( .A1(n7300), .A2(n7299), .ZN(n60140) );
  OR2_X1 U25735 ( .A1(n50286), .A2(n17957), .Z(n60375) );
  INV_X1 U25742 ( .I(n55385), .ZN(n21210) );
  NAND2_X1 U25745 ( .A1(n57184), .A2(n55385), .ZN(n61058) );
  NAND2_X1 U25750 ( .A1(n46764), .A2(n13348), .ZN(n13346) );
  AOI21_X1 U25757 ( .A1(n17028), .A2(n17027), .B(n1595), .ZN(n15508) );
  BUF_X2 U25759 ( .I(n55639), .Z(n58701) );
  XOR2_X1 U25777 ( .A1(n58703), .A2(n39233), .Z(n16536) );
  XOR2_X1 U25782 ( .A1(n25713), .A2(n39234), .Z(n58703) );
  XOR2_X1 U25804 ( .A1(n3164), .A2(n3165), .Z(n3163) );
  INV_X2 U25807 ( .I(n2026), .ZN(n58705) );
  AND2_X1 U25809 ( .A1(n27548), .A2(n26938), .Z(n58708) );
  AOI22_X2 U25810 ( .A1(n61820), .A2(n26965), .B1(n27214), .B2(n7437), .ZN(
        n25646) );
  NOR2_X2 U25815 ( .A1(n60162), .A2(n18402), .ZN(n13628) );
  NAND2_X2 U25817 ( .A1(n41614), .A2(n17223), .ZN(n20817) );
  XOR2_X1 U25829 ( .A1(n37624), .A2(n58827), .Z(n37792) );
  XOR2_X1 U25837 ( .A1(n50543), .A2(n15847), .Z(n10273) );
  XOR2_X1 U25841 ( .A1(n48703), .A2(n51959), .Z(n50543) );
  NAND3_X1 U25849 ( .A1(n9511), .A2(n4274), .A3(n22989), .ZN(n43034) );
  NOR3_X2 U25871 ( .A1(n35122), .A2(n36193), .A3(n36408), .ZN(n36192) );
  NOR2_X2 U25886 ( .A1(n5705), .A2(n21178), .ZN(n48237) );
  BUF_X2 U25890 ( .I(n1545), .Z(n58713) );
  XOR2_X1 U25901 ( .A1(n5755), .A2(n5754), .Z(n58715) );
  XOR2_X1 U25906 ( .A1(n33870), .A2(n58718), .Z(n58717) );
  INV_X2 U25911 ( .I(n54764), .ZN(n54726) );
  NOR2_X1 U25913 ( .A1(n52305), .A2(n52303), .ZN(n58720) );
  AND2_X1 U25928 ( .A1(n12798), .A2(n35852), .Z(n37444) );
  NAND2_X2 U25929 ( .A1(n16186), .A2(n18106), .ZN(n49676) );
  AND2_X1 U25938 ( .A1(n5193), .A2(n64176), .Z(n5195) );
  AND2_X1 U25955 ( .A1(n8941), .A2(n8944), .Z(n58729) );
  NAND3_X1 U25961 ( .A1(n6076), .A2(n17108), .A3(n60798), .ZN(n23808) );
  XOR2_X1 U25965 ( .A1(n50561), .A2(n58730), .Z(n50768) );
  XOR2_X1 U25972 ( .A1(n50560), .A2(n58731), .Z(n58730) );
  XOR2_X1 U25977 ( .A1(n58732), .A2(n15865), .Z(n33846) );
  NAND2_X2 U25984 ( .A1(n22444), .A2(n16491), .ZN(n29900) );
  BUF_X4 U25992 ( .I(n28933), .Z(n30680) );
  NOR3_X2 U25993 ( .A1(n42771), .A2(n58736), .A3(n4420), .ZN(n10153) );
  NAND2_X2 U25996 ( .A1(n18525), .A2(n24249), .ZN(n36163) );
  OR2_X1 U26007 ( .A1(n50074), .A2(n58840), .Z(n50402) );
  BUF_X2 U26016 ( .I(n14253), .Z(n58740) );
  XOR2_X1 U26027 ( .A1(n58744), .A2(n60968), .Z(n9358) );
  XOR2_X1 U26030 ( .A1(n11231), .A2(n2043), .Z(n58744) );
  XOR2_X1 U26033 ( .A1(n4867), .A2(n13278), .Z(n58745) );
  XOR2_X1 U26036 ( .A1(n2458), .A2(n11307), .Z(n2266) );
  XOR2_X1 U26052 ( .A1(n46268), .A2(n6904), .Z(n46381) );
  BUF_X2 U26053 ( .I(n15205), .Z(n58747) );
  NAND4_X1 U26067 ( .A1(n36898), .A2(n36533), .A3(n36538), .A4(n36385), .ZN(
        n58749) );
  XOR2_X1 U26068 ( .A1(n26029), .A2(n25192), .Z(n58751) );
  NAND2_X1 U26071 ( .A1(n20381), .A2(n53649), .ZN(n53652) );
  XOR2_X1 U26072 ( .A1(n11852), .A2(n11446), .Z(n10241) );
  NAND2_X1 U26074 ( .A1(n50394), .A2(n8994), .ZN(n20174) );
  NAND2_X1 U26080 ( .A1(n46457), .A2(n46458), .ZN(n58753) );
  INV_X1 U26081 ( .I(n46456), .ZN(n58754) );
  NAND2_X1 U26092 ( .A1(n35022), .A2(n58756), .ZN(n34552) );
  NOR2_X1 U26095 ( .A1(n2210), .A2(n902), .ZN(n58756) );
  INV_X4 U26097 ( .I(n59106), .ZN(n29794) );
  INV_X2 U26104 ( .I(n58757), .ZN(n31692) );
  XOR2_X1 U26108 ( .A1(n33898), .A2(n29818), .Z(n58757) );
  AOI22_X1 U26109 ( .A1(n10755), .A2(n29664), .B1(n29666), .B2(n29665), .ZN(
        n29679) );
  NAND2_X1 U26112 ( .A1(n4929), .A2(n52273), .ZN(n58789) );
  NOR2_X2 U26114 ( .A1(n58759), .A2(n2729), .ZN(n2727) );
  XOR2_X1 U26115 ( .A1(n58760), .A2(n45108), .Z(n22483) );
  XOR2_X1 U26116 ( .A1(n45107), .A2(n22340), .Z(n58760) );
  XOR2_X1 U26131 ( .A1(n58762), .A2(n45341), .Z(n61564) );
  AND2_X1 U26139 ( .A1(n23411), .A2(n9481), .Z(n9943) );
  NOR2_X2 U26143 ( .A1(n57211), .A2(n36139), .ZN(n36794) );
  NAND2_X2 U26146 ( .A1(n58764), .A2(n25980), .ZN(n22699) );
  NOR2_X2 U26168 ( .A1(n43513), .A2(n43504), .ZN(n43521) );
  NOR4_X2 U26172 ( .A1(n27635), .A2(n30396), .A3(n30392), .A4(n29511), .ZN(
        n59671) );
  XOR2_X1 U26181 ( .A1(n39565), .A2(n7851), .Z(n961) );
  OAI22_X1 U26182 ( .A1(n2287), .A2(n61496), .B1(n15148), .B2(n35743), .ZN(
        n35196) );
  NAND3_X2 U26200 ( .A1(n39056), .A2(n39055), .A3(n39860), .ZN(n39081) );
  NAND2_X2 U26204 ( .A1(n1336), .A2(n42968), .ZN(n43458) );
  NAND2_X2 U26209 ( .A1(n56659), .A2(n24259), .ZN(n18121) );
  NAND2_X1 U26223 ( .A1(n51403), .A2(n20634), .ZN(n58767) );
  NOR2_X2 U26236 ( .A1(n58770), .A2(n25818), .ZN(n50948) );
  NOR3_X2 U26245 ( .A1(n19674), .A2(n60180), .A3(n60179), .ZN(n19672) );
  NOR2_X2 U26248 ( .A1(n18608), .A2(n1224), .ZN(n50286) );
  NAND2_X2 U26252 ( .A1(n14196), .A2(n24351), .ZN(n36072) );
  NOR2_X1 U26269 ( .A1(n37962), .A2(n37048), .ZN(n37057) );
  NOR3_X2 U26275 ( .A1(n36605), .A2(n21915), .A3(n62672), .ZN(n37962) );
  NOR2_X2 U26292 ( .A1(n9281), .A2(n22903), .ZN(n27913) );
  AND2_X1 U26293 ( .A1(n53462), .A2(n9595), .Z(n53491) );
  XOR2_X1 U26301 ( .A1(n31859), .A2(n58775), .Z(n60234) );
  XOR2_X1 U26302 ( .A1(n30848), .A2(n26444), .Z(n31859) );
  XOR2_X1 U26307 ( .A1(n58776), .A2(n56309), .Z(Plaintext[151]) );
  NAND2_X2 U26308 ( .A1(n1256), .A2(n57202), .ZN(n54254) );
  OR2_X1 U26322 ( .A1(n6720), .A2(n29242), .Z(n30823) );
  NOR2_X2 U26323 ( .A1(n34247), .A2(n34727), .ZN(n34726) );
  NOR2_X2 U26332 ( .A1(n30809), .A2(n8521), .ZN(n30816) );
  INV_X2 U26336 ( .I(n56327), .ZN(n1580) );
  NAND2_X2 U26338 ( .A1(n23318), .A2(n12058), .ZN(n56327) );
  NAND4_X1 U26341 ( .A1(n41129), .A2(n13846), .A3(n41380), .A4(n41128), .ZN(
        n60822) );
  XOR2_X1 U26343 ( .A1(n20776), .A2(n58780), .Z(n22355) );
  XOR2_X1 U26361 ( .A1(n33207), .A2(n58781), .Z(n58780) );
  NOR2_X2 U26365 ( .A1(n1339), .A2(n32940), .ZN(n18850) );
  XOR2_X1 U26367 ( .A1(n46289), .A2(n46290), .Z(n58782) );
  XOR2_X1 U26378 ( .A1(n58783), .A2(n39759), .Z(n39642) );
  XOR2_X1 U26381 ( .A1(n39637), .A2(n39638), .Z(n58783) );
  OAI21_X2 U26389 ( .A1(n33018), .A2(n33019), .B(n11061), .ZN(n58785) );
  NOR2_X1 U26394 ( .A1(n3613), .A2(n56343), .ZN(n56340) );
  NOR2_X1 U26410 ( .A1(n55748), .A2(n55749), .ZN(n55755) );
  BUF_X4 U26412 ( .I(n49072), .Z(n11950) );
  XOR2_X1 U26429 ( .A1(n4616), .A2(n5181), .Z(n9396) );
  NOR2_X2 U26452 ( .A1(n59536), .A2(n46937), .ZN(n47982) );
  NAND3_X2 U26455 ( .A1(n59547), .A2(n10437), .A3(n47106), .ZN(n50229) );
  XOR2_X1 U26456 ( .A1(n46519), .A2(n46136), .Z(n6326) );
  NAND2_X2 U26470 ( .A1(n58790), .A2(n15254), .ZN(n36623) );
  NOR2_X2 U26471 ( .A1(n56958), .A2(n14708), .ZN(n56919) );
  NAND2_X2 U26474 ( .A1(n5017), .A2(n58791), .ZN(n49598) );
  NOR2_X1 U26475 ( .A1(n9449), .A2(n25033), .ZN(n58791) );
  OAI22_X1 U26486 ( .A1(n2020), .A2(n36336), .B1(n36335), .B2(n63593), .ZN(
        n2019) );
  AND2_X2 U26487 ( .A1(n48546), .A2(n48555), .Z(n48155) );
  OR2_X1 U26488 ( .A1(n55244), .A2(n54980), .Z(n19505) );
  NAND3_X1 U26499 ( .A1(n5949), .A2(n6297), .A3(n61107), .ZN(n13099) );
  NAND2_X2 U26502 ( .A1(n36170), .A2(n22169), .ZN(n12804) );
  NOR3_X2 U26503 ( .A1(n30465), .A2(n58793), .A3(n30466), .ZN(n30473) );
  NOR3_X1 U26506 ( .A1(n1532), .A2(n34069), .A3(n21008), .ZN(n58793) );
  NAND3_X2 U26507 ( .A1(n7993), .A2(n17094), .A3(n17093), .ZN(n58863) );
  BUF_X2 U26508 ( .I(n1743), .Z(n58794) );
  OAI21_X1 U26516 ( .A1(n58796), .A2(n58795), .B(n56731), .ZN(n23097) );
  NOR2_X1 U26524 ( .A1(n17532), .A2(n56707), .ZN(n58795) );
  INV_X2 U26552 ( .I(n40716), .ZN(n58798) );
  XOR2_X1 U26553 ( .A1(n59490), .A2(n51584), .Z(n12606) );
  XOR2_X1 U26556 ( .A1(n6959), .A2(n6960), .Z(n51584) );
  NAND2_X2 U26558 ( .A1(n4734), .A2(n50054), .ZN(n50059) );
  XOR2_X1 U26559 ( .A1(n22530), .A2(n58799), .Z(n52543) );
  XOR2_X1 U26560 ( .A1(n52539), .A2(n52540), .Z(n58799) );
  OAI21_X1 U26564 ( .A1(n36607), .A2(n35105), .B(n35104), .ZN(n60135) );
  NAND3_X2 U26571 ( .A1(n22394), .A2(n45438), .A3(n16658), .ZN(n58800) );
  XOR2_X1 U26572 ( .A1(n60206), .A2(n58801), .Z(n60423) );
  XOR2_X1 U26575 ( .A1(n58802), .A2(n25582), .Z(n58801) );
  NOR3_X2 U26577 ( .A1(n8751), .A2(n25955), .A3(n25954), .ZN(n8750) );
  XNOR2_X1 U26588 ( .A1(n45030), .A2(n46291), .ZN(n5214) );
  AOI22_X2 U26591 ( .A1(n41735), .A2(n41736), .B1(n41737), .B2(n42834), .ZN(
        n45030) );
  AOI21_X2 U26605 ( .A1(n18096), .A2(n23526), .B(n56830), .ZN(n18095) );
  NAND2_X1 U26616 ( .A1(n4985), .A2(n59320), .ZN(n55043) );
  NAND3_X2 U26617 ( .A1(n53097), .A2(n23212), .A3(n1281), .ZN(n53048) );
  NOR2_X2 U26627 ( .A1(n54960), .A2(n25220), .ZN(n55064) );
  NAND2_X2 U26633 ( .A1(n49649), .A2(n3123), .ZN(n50053) );
  INV_X4 U26634 ( .I(n1301), .ZN(n42361) );
  BUF_X4 U26638 ( .I(n24948), .Z(n59658) );
  AOI22_X1 U26640 ( .A1(n4046), .A2(n36718), .B1(n21468), .B2(n36719), .ZN(
        n19012) );
  NOR2_X2 U26646 ( .A1(n2403), .A2(n59071), .ZN(n48581) );
  AND2_X1 U26647 ( .A1(n50399), .A2(n58840), .Z(n1067) );
  BUF_X4 U26652 ( .I(n36955), .Z(n60694) );
  NOR2_X2 U26662 ( .A1(n25220), .A2(n9068), .ZN(n55057) );
  AOI21_X2 U26665 ( .A1(n40891), .A2(n40890), .B(n1301), .ZN(n42354) );
  NAND2_X2 U26667 ( .A1(n3055), .A2(n50142), .ZN(n50306) );
  INV_X2 U26669 ( .I(n27516), .ZN(n30271) );
  BUF_X4 U26681 ( .I(n56552), .Z(n56719) );
  AOI21_X1 U26684 ( .A1(n52702), .A2(n23095), .B(n1153), .ZN(n52703) );
  NAND4_X1 U26686 ( .A1(n56688), .A2(n56678), .A3(n56725), .A4(n20696), .ZN(
        n56679) );
  INV_X1 U26695 ( .I(n14761), .ZN(n15811) );
  NAND2_X1 U26703 ( .A1(n15281), .A2(n22544), .ZN(n15346) );
  NAND2_X1 U26711 ( .A1(n15281), .A2(n26095), .ZN(n54948) );
  INV_X1 U26721 ( .I(n51855), .ZN(n54314) );
  CLKBUF_X2 U26727 ( .I(n56687), .Z(n20696) );
  NOR2_X1 U26728 ( .A1(n56708), .A2(n56687), .ZN(n56674) );
  NAND2_X1 U26746 ( .A1(n53676), .A2(n53672), .ZN(n53667) );
  CLKBUF_X4 U26753 ( .I(n51628), .Z(n10101) );
  OAI21_X1 U26754 ( .A1(n64872), .A2(n56848), .B(n56861), .ZN(n17648) );
  OAI21_X1 U26757 ( .A1(n61123), .A2(n59970), .B(n54026), .ZN(n53884) );
  OAI21_X1 U26761 ( .A1(n60226), .A2(n16487), .B(n10425), .ZN(n21971) );
  AOI21_X1 U26769 ( .A1(n16713), .A2(n17928), .B(n43733), .ZN(n42124) );
  NOR2_X1 U26775 ( .A1(n16713), .A2(n43733), .ZN(n19047) );
  INV_X2 U26782 ( .I(n47748), .ZN(n24252) );
  NAND2_X1 U26793 ( .A1(n53781), .A2(n61415), .ZN(n61414) );
  INV_X1 U26803 ( .I(n2367), .ZN(n44118) );
  INV_X1 U26811 ( .I(n5219), .ZN(n48446) );
  AND2_X2 U26817 ( .A1(n5348), .A2(n59786), .Z(n10174) );
  INV_X1 U26819 ( .I(n15935), .ZN(n13426) );
  INV_X1 U26825 ( .I(n49499), .ZN(n9294) );
  AOI21_X1 U26839 ( .A1(n20671), .A2(n9292), .B(n9290), .ZN(n4626) );
  NOR2_X1 U26850 ( .A1(n11841), .A2(n59445), .ZN(n11654) );
  INV_X1 U26867 ( .I(n50964), .ZN(n59555) );
  NOR2_X1 U26877 ( .A1(n56248), .A2(n56245), .ZN(n61492) );
  CLKBUF_X4 U26881 ( .I(n4808), .Z(n2820) );
  NAND2_X1 U26882 ( .A1(n6431), .A2(n60313), .ZN(n152) );
  AOI22_X1 U26895 ( .A1(n56217), .A2(n56216), .B1(n64345), .B2(n56619), .ZN(
        n56218) );
  NAND2_X1 U26897 ( .A1(n7055), .A2(n13026), .ZN(n55425) );
  XOR2_X1 U26901 ( .A1(n5406), .A2(n5403), .Z(n58806) );
  INV_X4 U26908 ( .I(n15425), .ZN(n15615) );
  NAND3_X1 U26911 ( .A1(n53555), .A2(n53404), .A3(n54044), .ZN(n53405) );
  NAND2_X1 U26922 ( .A1(n21705), .A2(n1085), .ZN(n58883) );
  INV_X1 U26926 ( .I(n56587), .ZN(n24321) );
  AOI21_X1 U26928 ( .A1(n56587), .A2(n56245), .B(n55957), .ZN(n5020) );
  NAND2_X1 U26948 ( .A1(n21833), .A2(n49951), .ZN(n58917) );
  OAI21_X2 U26954 ( .A1(n8621), .A2(n2630), .B(n51213), .ZN(n2221) );
  NAND2_X1 U26961 ( .A1(n56673), .A2(n13249), .ZN(n60564) );
  NOR2_X1 U26963 ( .A1(n13249), .A2(n23785), .ZN(n17532) );
  CLKBUF_X2 U26966 ( .I(n56084), .Z(n60672) );
  OAI22_X1 U26980 ( .A1(n54322), .A2(n54321), .B1(n1368), .B2(n6211), .ZN(
        n6459) );
  NAND2_X1 U26981 ( .A1(n54472), .A2(n54594), .ZN(n6211) );
  INV_X1 U26988 ( .I(n17972), .ZN(n28836) );
  BUF_X1 U26989 ( .I(n20623), .Z(n10325) );
  INV_X2 U26996 ( .I(n109), .ZN(n10481) );
  CLKBUF_X2 U27021 ( .I(n51570), .Z(n6384) );
  CLKBUF_X4 U27025 ( .I(n21470), .Z(n15700) );
  OR2_X1 U27026 ( .A1(n61829), .A2(n11275), .Z(n11248) );
  XOR2_X1 U27029 ( .A1(n24733), .A2(n19268), .Z(n58807) );
  OAI21_X1 U27035 ( .A1(n42641), .A2(n20888), .B(n43184), .ZN(n43196) );
  NAND3_X1 U27036 ( .A1(n50221), .A2(n50216), .A3(n1262), .ZN(n49101) );
  NAND2_X1 U27042 ( .A1(n3618), .A2(n16850), .ZN(n42167) );
  OR2_X1 U27048 ( .A1(n49546), .A2(n49528), .Z(n47914) );
  AOI22_X1 U27053 ( .A1(n56864), .A2(n56865), .B1(n56866), .B2(n22667), .ZN(
        n60956) );
  AOI22_X1 U27054 ( .A1(n53994), .A2(n53993), .B1(n59662), .B2(n53991), .ZN(
        n5650) );
  AOI22_X1 U27055 ( .A1(n55897), .A2(n55870), .B1(n15716), .B2(n55847), .ZN(
        n59630) );
  AOI21_X1 U27069 ( .A1(n62886), .A2(n57070), .B(n57083), .ZN(n51470) );
  CLKBUF_X4 U27070 ( .I(n36245), .Z(n22431) );
  INV_X1 U27072 ( .I(n53455), .ZN(n60310) );
  NAND2_X1 U27073 ( .A1(n53586), .A2(n53455), .ZN(n9296) );
  AOI21_X1 U27076 ( .A1(n59232), .A2(n59231), .B(n1008), .ZN(n26036) );
  INV_X1 U27078 ( .I(n45766), .ZN(n6599) );
  NAND2_X1 U27080 ( .A1(n4283), .A2(n53294), .ZN(n53295) );
  NOR2_X2 U27081 ( .A1(n52963), .A2(n59256), .ZN(n58808) );
  NAND4_X1 U27086 ( .A1(n53259), .A2(n53260), .A3(n53268), .A4(n53261), .ZN(
        n58932) );
  OAI21_X1 U27103 ( .A1(n55696), .A2(n1285), .B(n18548), .ZN(n11023) );
  AND4_X1 U27109 ( .A1(n26145), .A2(n3364), .A3(n48659), .A4(n16616), .Z(
        n58809) );
  NOR2_X1 U27113 ( .A1(n9795), .A2(n59340), .ZN(n12947) );
  NAND2_X1 U27119 ( .A1(n4830), .A2(n60553), .ZN(n60552) );
  OAI21_X1 U27121 ( .A1(n53192), .A2(n53198), .B(n52752), .ZN(n52753) );
  NAND2_X1 U27126 ( .A1(n22720), .A2(n10198), .ZN(n17993) );
  NOR2_X1 U27131 ( .A1(n1541), .A2(n60175), .ZN(n905) );
  INV_X2 U27133 ( .I(n19803), .ZN(n20288) );
  INV_X2 U27134 ( .I(n23900), .ZN(n1260) );
  NOR2_X1 U27162 ( .A1(n65276), .A2(n49429), .ZN(n49431) );
  NAND2_X1 U27173 ( .A1(n6987), .A2(n22484), .ZN(n48229) );
  NOR2_X1 U27175 ( .A1(n6987), .A2(n8732), .ZN(n8749) );
  NOR2_X1 U27177 ( .A1(n59049), .A2(n54450), .ZN(n58810) );
  INV_X2 U27178 ( .I(n8147), .ZN(n52103) );
  CLKBUF_X4 U27182 ( .I(n51832), .Z(n10461) );
  INV_X1 U27183 ( .I(n7811), .ZN(n11284) );
  OAI21_X1 U27184 ( .A1(n54835), .A2(n58283), .B(n54843), .ZN(n60629) );
  NAND2_X1 U27197 ( .A1(n60075), .A2(n21493), .ZN(n11525) );
  INV_X1 U27200 ( .I(n19890), .ZN(n51823) );
  NAND4_X1 U27205 ( .A1(n56333), .A2(n56334), .A3(n56332), .A4(n56331), .ZN(
        n9763) );
  INV_X1 U27209 ( .I(n49790), .ZN(n46000) );
  AND2_X1 U27210 ( .A1(n55133), .A2(n55135), .Z(n58884) );
  NAND3_X1 U27211 ( .A1(n53365), .A2(n16778), .A3(n53369), .ZN(n53372) );
  NOR2_X1 U27240 ( .A1(n1259), .A2(n9514), .ZN(n53855) );
  CLKBUF_X4 U27242 ( .I(n50462), .Z(n61560) );
  NOR2_X1 U27254 ( .A1(n24117), .A2(n22343), .ZN(n52964) );
  INV_X1 U27257 ( .I(n52964), .ZN(n55217) );
  CLKBUF_X8 U27269 ( .I(n23585), .Z(n20124) );
  NAND2_X1 U27276 ( .A1(n55818), .A2(n22925), .ZN(n55781) );
  INV_X2 U27279 ( .I(n52122), .ZN(n55915) );
  NAND2_X1 U27281 ( .A1(n52122), .A2(n15454), .ZN(n55719) );
  BUF_X4 U27283 ( .I(n5194), .Z(n5172) );
  NAND2_X1 U27285 ( .A1(n54713), .A2(n54726), .ZN(n59094) );
  NAND3_X1 U27286 ( .A1(n54853), .A2(n54854), .A3(n54855), .ZN(n59030) );
  NAND3_X2 U27295 ( .A1(n19748), .A2(n59389), .A3(n19743), .ZN(n58814) );
  NAND4_X1 U27299 ( .A1(n26198), .A2(n53914), .A3(n58656), .A4(n53557), .ZN(
        n485) );
  NAND2_X1 U27314 ( .A1(n56100), .A2(n56108), .ZN(n9569) );
  INV_X2 U27318 ( .I(n13567), .ZN(n58815) );
  INV_X2 U27322 ( .I(n46455), .ZN(n48459) );
  NAND3_X1 U27325 ( .A1(n9099), .A2(n14520), .A3(n46455), .ZN(n46456) );
  OAI21_X1 U27327 ( .A1(n15005), .A2(n15006), .B(n3123), .ZN(n9499) );
  NAND2_X1 U27330 ( .A1(n22304), .A2(n40628), .ZN(n39025) );
  NAND2_X1 U27341 ( .A1(n23141), .A2(n22869), .ZN(n22022) );
  NOR2_X2 U27342 ( .A1(n1255), .A2(n56867), .ZN(n59273) );
  NAND2_X1 U27349 ( .A1(n60781), .A2(n60780), .ZN(n60779) );
  INV_X1 U27357 ( .I(n53181), .ZN(n52746) );
  NOR2_X2 U27359 ( .A1(n13440), .A2(n48676), .ZN(n49441) );
  NAND2_X1 U27362 ( .A1(n25989), .A2(n4257), .ZN(n31278) );
  NAND2_X1 U27371 ( .A1(n54714), .A2(n54768), .ZN(n59095) );
  INV_X1 U27374 ( .I(n31476), .ZN(n58876) );
  BUF_X2 U27375 ( .I(n23604), .Z(n2951) );
  INV_X1 U27377 ( .I(n23604), .ZN(n9160) );
  NAND2_X1 U27379 ( .A1(n47425), .A2(n57852), .ZN(n46755) );
  NAND2_X1 U27381 ( .A1(n47687), .A2(n47425), .ZN(n47413) );
  INV_X1 U27382 ( .I(n47425), .ZN(n47427) );
  NAND4_X1 U27383 ( .A1(n56792), .A2(n56791), .A3(n65064), .A4(n7209), .ZN(
        n56751) );
  XOR2_X1 U27387 ( .A1(n51628), .A2(n58818), .Z(n20675) );
  INV_X1 U27389 ( .I(n50646), .ZN(n58818) );
  INV_X1 U27390 ( .I(n51628), .ZN(n51404) );
  NAND2_X1 U27397 ( .A1(n49226), .A2(n5587), .ZN(n7328) );
  NAND2_X1 U27402 ( .A1(n60159), .A2(n23874), .ZN(n53365) );
  NOR2_X1 U27408 ( .A1(n7328), .A2(n16595), .ZN(n60718) );
  AND2_X2 U27423 ( .A1(n48676), .A2(n18502), .Z(n15124) );
  NOR2_X1 U27425 ( .A1(n5275), .A2(n1143), .ZN(n60762) );
  NOR2_X1 U27430 ( .A1(n54457), .A2(n58526), .ZN(n61551) );
  NOR2_X1 U27432 ( .A1(n54636), .A2(n54640), .ZN(n61552) );
  NAND3_X1 U27434 ( .A1(n54403), .A2(n54419), .A3(n54393), .ZN(n6559) );
  NAND2_X1 U27438 ( .A1(n2676), .A2(n54403), .ZN(n6558) );
  INV_X1 U27439 ( .I(n51510), .ZN(n60300) );
  NAND2_X1 U27441 ( .A1(n59928), .A2(n64307), .ZN(n59927) );
  OAI21_X1 U27442 ( .A1(n64307), .A2(n54596), .B(n22065), .ZN(n22064) );
  OAI21_X1 U27456 ( .A1(n56756), .A2(n56778), .B(n56790), .ZN(n5895) );
  OAI21_X1 U27457 ( .A1(n49891), .A2(n50122), .B(n47956), .ZN(n10112) );
  NAND2_X1 U27459 ( .A1(n63355), .A2(n29244), .ZN(n13338) );
  NAND3_X1 U27461 ( .A1(n58710), .A2(n29244), .A3(n63355), .ZN(n28945) );
  INV_X4 U27481 ( .I(n53950), .ZN(n54001) );
  BUF_X4 U27483 ( .I(n22084), .Z(n60583) );
  NAND2_X1 U27484 ( .A1(n22084), .A2(n43852), .ZN(n43842) );
  AOI22_X1 U27492 ( .A1(n56986), .A2(n13757), .B1(n56984), .B2(n56985), .ZN(
        n56996) );
  XOR2_X1 U27496 ( .A1(n9876), .A2(n7847), .Z(n58819) );
  INV_X1 U27505 ( .I(n8781), .ZN(n4008) );
  OAI22_X1 U27524 ( .A1(n56981), .A2(n7835), .B1(n56984), .B2(n52687), .ZN(
        n17543) );
  NAND2_X1 U27525 ( .A1(n30743), .A2(n30632), .ZN(n28683) );
  INV_X2 U27536 ( .I(n30632), .ZN(n24564) );
  BUF_X2 U27539 ( .I(n30632), .Z(n22745) );
  AND2_X2 U27553 ( .A1(n20139), .A2(n15728), .Z(n48102) );
  NAND3_X1 U27567 ( .A1(n43577), .A2(n43573), .A3(n42726), .ZN(n42342) );
  NOR2_X1 U27569 ( .A1(n43573), .A2(n64946), .ZN(n43578) );
  NAND2_X1 U27570 ( .A1(n43573), .A2(n5398), .ZN(n13605) );
  NAND2_X1 U27572 ( .A1(n7165), .A2(n41473), .ZN(n61526) );
  INV_X2 U27579 ( .I(n31077), .ZN(n29472) );
  BUF_X2 U27588 ( .I(n31077), .Z(n22411) );
  CLKBUF_X4 U27596 ( .I(n54758), .Z(n14848) );
  INV_X1 U27611 ( .I(n52507), .ZN(n60483) );
  NAND2_X1 U27612 ( .A1(n13389), .A2(n1270), .ZN(n42806) );
  AOI21_X1 U27628 ( .A1(n42900), .A2(n43147), .B(n13528), .ZN(n42568) );
  AND2_X2 U27638 ( .A1(n40096), .A2(n22050), .Z(n42070) );
  NOR2_X1 U27644 ( .A1(n57298), .A2(n9064), .ZN(n60313) );
  NAND3_X1 U27647 ( .A1(n138), .A2(n56919), .A3(n56936), .ZN(n59853) );
  NOR2_X1 U27650 ( .A1(n56659), .A2(n24259), .ZN(n59783) );
  AOI21_X1 U27653 ( .A1(n46905), .A2(n6599), .B(n62366), .ZN(n44778) );
  NAND2_X1 U27664 ( .A1(n2011), .A2(n2010), .ZN(n2009) );
  AOI22_X1 U27674 ( .A1(n6622), .A2(n18740), .B1(n54905), .B2(n6621), .ZN(
        n59226) );
  INV_X1 U27679 ( .I(n55017), .ZN(n14457) );
  CLKBUF_X2 U27685 ( .I(n54860), .Z(n10523) );
  INV_X1 U27686 ( .I(n54860), .ZN(n22900) );
  INV_X2 U27697 ( .I(n20996), .ZN(n9045) );
  INV_X1 U27704 ( .I(n56424), .ZN(n55980) );
  CLKBUF_X4 U27709 ( .I(n15306), .Z(n14316) );
  OAI21_X1 U27713 ( .A1(n56688), .A2(n2422), .B(n22024), .ZN(n11851) );
  INV_X4 U27715 ( .I(n56719), .ZN(n56725) );
  NAND3_X1 U27719 ( .A1(n53491), .A2(n23611), .A3(n53528), .ZN(n53529) );
  INV_X2 U27724 ( .I(n17775), .ZN(n35416) );
  NAND2_X1 U27730 ( .A1(n35943), .A2(n2607), .ZN(n3763) );
  INV_X1 U27731 ( .I(n35943), .ZN(n36914) );
  NOR2_X1 U27735 ( .A1(n47154), .A2(n48484), .ZN(n46469) );
  INV_X1 U27750 ( .I(n47154), .ZN(n48585) );
  INV_X1 U27752 ( .I(n12835), .ZN(n61032) );
  INV_X1 U27758 ( .I(n12835), .ZN(n24094) );
  INV_X1 U27765 ( .I(n46201), .ZN(n61591) );
  XOR2_X1 U27769 ( .A1(n61947), .A2(n13183), .Z(n58822) );
  CLKBUF_X12 U27781 ( .I(n7388), .Z(n58824) );
  NOR2_X2 U27787 ( .A1(n6743), .A2(n6742), .ZN(n58825) );
  BUF_X2 U27792 ( .I(n6744), .Z(n5155) );
  NAND3_X1 U27794 ( .A1(n658), .A2(n55962), .A3(n55964), .ZN(n58826) );
  NOR2_X1 U27813 ( .A1(n23750), .A2(n37006), .ZN(n37015) );
  NOR2_X1 U27826 ( .A1(n47696), .A2(n47798), .ZN(n45309) );
  CLKBUF_X4 U27827 ( .I(n26278), .Z(n28048) );
  NOR2_X1 U27829 ( .A1(n48233), .A2(n48232), .ZN(n60144) );
  AOI22_X1 U27836 ( .A1(n35402), .A2(n2885), .B1(n36790), .B2(n35401), .ZN(
        n35403) );
  XOR2_X1 U27844 ( .A1(n11285), .A2(n11283), .Z(n58830) );
  NAND2_X2 U27852 ( .A1(n36394), .A2(n36529), .ZN(n19206) );
  NAND2_X1 U27858 ( .A1(n7846), .A2(n14335), .ZN(n50212) );
  BUF_X2 U27861 ( .I(n43844), .Z(n22673) );
  AND3_X1 U27865 ( .A1(n50281), .A2(n50280), .A3(n50282), .Z(n58832) );
  INV_X1 U27868 ( .I(n48483), .ZN(n24185) );
  NAND2_X1 U27883 ( .A1(n59409), .A2(n41887), .ZN(n37828) );
  CLKBUF_X2 U27887 ( .I(n41887), .Z(n59803) );
  NAND2_X1 U27889 ( .A1(n14488), .A2(n50257), .ZN(n15793) );
  INV_X1 U27892 ( .I(n61350), .ZN(n33635) );
  BUF_X2 U27899 ( .I(n2674), .Z(n61350) );
  NAND2_X1 U27901 ( .A1(n49496), .A2(n49493), .ZN(n47041) );
  NAND2_X1 U27902 ( .A1(n43099), .A2(n42993), .ZN(n43094) );
  INV_X1 U27908 ( .I(n43099), .ZN(n7285) );
  XOR2_X1 U27922 ( .A1(n17584), .A2(n44434), .Z(n58835) );
  NAND3_X1 U27923 ( .A1(n63721), .A2(n42865), .A3(n6764), .ZN(n16546) );
  NAND2_X1 U27928 ( .A1(n59948), .A2(n6764), .ZN(n59947) );
  INV_X1 U27930 ( .I(n16582), .ZN(n58836) );
  INV_X1 U27931 ( .I(n58836), .ZN(n58837) );
  INV_X2 U27936 ( .I(n23230), .ZN(n9663) );
  INV_X1 U27942 ( .I(n44077), .ZN(n9157) );
  BUF_X2 U27943 ( .I(n26095), .Z(n22749) );
  XOR2_X1 U27948 ( .A1(n3279), .A2(n3277), .Z(n58839) );
  INV_X2 U27953 ( .I(n50395), .ZN(n4173) );
  CLKBUF_X1 U27972 ( .I(n25315), .Z(n25787) );
  NAND2_X1 U27983 ( .A1(n45715), .A2(n24578), .ZN(n12597) );
  NAND2_X1 U27984 ( .A1(n19375), .A2(n45715), .ZN(n44556) );
  CLKBUF_X4 U27990 ( .I(n24277), .Z(n8449) );
  AND4_X1 U27993 ( .A1(n35503), .A2(n35501), .A3(n18509), .A4(n35502), .Z(
        n58842) );
  AOI21_X1 U27998 ( .A1(n48529), .A2(n20878), .B(n57728), .ZN(n48112) );
  NAND3_X1 U27999 ( .A1(n21177), .A2(n20878), .A3(n46716), .ZN(n48528) );
  AND3_X2 U28001 ( .A1(n57728), .A2(n12100), .A3(n20878), .Z(n48120) );
  INV_X2 U28006 ( .I(n20878), .ZN(n6987) );
  INV_X2 U28008 ( .I(n62768), .ZN(n19137) );
  NAND3_X2 U28034 ( .A1(n45755), .A2(n45754), .A3(n58845), .ZN(n48069) );
  XOR2_X1 U28037 ( .A1(n39713), .A2(n39712), .Z(n39719) );
  XOR2_X1 U28045 ( .A1(n21331), .A2(n61569), .Z(n39713) );
  NAND3_X2 U28055 ( .A1(n59074), .A2(n51447), .A3(n51448), .ZN(n51449) );
  NOR2_X1 U28101 ( .A1(n21633), .A2(n27398), .ZN(n58855) );
  BUF_X4 U28115 ( .I(n36070), .Z(n61579) );
  XOR2_X1 U28123 ( .A1(n31597), .A2(n13475), .Z(n58858) );
  XOR2_X1 U28124 ( .A1(n31346), .A2(n31351), .Z(n58859) );
  NOR2_X2 U28126 ( .A1(n22782), .A2(n11557), .ZN(n11275) );
  NAND2_X2 U28128 ( .A1(n15204), .A2(n15203), .ZN(n22782) );
  NAND4_X2 U28146 ( .A1(n24994), .A2(n21584), .A3(n60022), .A4(n10849), .ZN(
        n36699) );
  NAND2_X1 U28153 ( .A1(n20045), .A2(n50932), .ZN(n20016) );
  AOI21_X2 U28164 ( .A1(n30768), .A2(n30790), .B(n58862), .ZN(n16603) );
  OAI22_X2 U28165 ( .A1(n29962), .A2(n29961), .B1(n29960), .B2(n30786), .ZN(
        n58862) );
  NAND2_X2 U28169 ( .A1(n17057), .A2(n3888), .ZN(n25080) );
  NAND4_X1 U28171 ( .A1(n37928), .A2(n37927), .A3(n40932), .A4(n40470), .ZN(
        n58864) );
  NAND2_X2 U28172 ( .A1(n65269), .A2(n7732), .ZN(n20842) );
  OAI21_X2 U28182 ( .A1(n14726), .A2(n31779), .B(n1420), .ZN(n7732) );
  AND2_X1 U28183 ( .A1(n11184), .A2(n6277), .Z(n61677) );
  NOR2_X2 U28184 ( .A1(n4347), .A2(n4346), .ZN(n58867) );
  NAND2_X1 U28188 ( .A1(n53781), .A2(n53794), .ZN(n58868) );
  NAND2_X1 U28226 ( .A1(n4139), .A2(n4140), .ZN(n4138) );
  XOR2_X1 U28231 ( .A1(n4343), .A2(n58878), .Z(n5094) );
  INV_X1 U28233 ( .I(n54776), .ZN(n58878) );
  NAND2_X1 U28247 ( .A1(n47100), .A2(n47101), .ZN(n58881) );
  AOI21_X1 U28248 ( .A1(n56602), .A2(n56601), .B(n13920), .ZN(n59404) );
  NOR2_X1 U28251 ( .A1(n40983), .A2(n40984), .ZN(n41000) );
  XNOR2_X1 U28253 ( .A1(n39491), .A2(n37563), .ZN(n3053) );
  OR2_X2 U28271 ( .A1(n28711), .A2(n30413), .Z(n30651) );
  XOR2_X1 U28274 ( .A1(n51017), .A2(n57351), .Z(n52529) );
  NOR3_X2 U28287 ( .A1(n49802), .A2(n58886), .A3(n58885), .ZN(n8292) );
  AND2_X1 U28292 ( .A1(n4043), .A2(n19163), .Z(n20096) );
  BUF_X4 U28320 ( .I(n35680), .Z(n59534) );
  OR3_X2 U28324 ( .A1(n3669), .A2(n34973), .A3(n7883), .Z(n34531) );
  NAND2_X2 U28333 ( .A1(n1639), .A2(n23247), .ZN(n19003) );
  NAND4_X2 U28346 ( .A1(n46853), .A2(n49726), .A3(n47934), .A4(n58892), .ZN(
        n49621) );
  XOR2_X1 U28356 ( .A1(n58895), .A2(n20081), .Z(n7884) );
  XOR2_X1 U28361 ( .A1(n20083), .A2(n20084), .Z(n58895) );
  OR2_X1 U28362 ( .A1(n54523), .A2(n18425), .Z(n54522) );
  NAND2_X1 U28391 ( .A1(n59125), .A2(n24093), .ZN(n33638) );
  NAND4_X2 U28401 ( .A1(n58897), .A2(n24680), .A3(n19096), .A4(n15165), .ZN(
        n11502) );
  NAND2_X1 U28403 ( .A1(n15170), .A2(n49733), .ZN(n58897) );
  NAND2_X1 U28422 ( .A1(n47984), .A2(n47232), .ZN(n6496) );
  NAND3_X2 U28432 ( .A1(n22724), .A2(n22942), .A3(n33367), .ZN(n36245) );
  NAND3_X1 U28434 ( .A1(n55147), .A2(n55148), .A3(n7890), .ZN(n55149) );
  XOR2_X1 U28442 ( .A1(n58904), .A2(n32736), .Z(n5747) );
  XOR2_X1 U28443 ( .A1(n31933), .A2(n23683), .Z(n58904) );
  XOR2_X1 U28445 ( .A1(n52206), .A2(n31931), .Z(n44351) );
  XOR2_X1 U28448 ( .A1(n61238), .A2(n50798), .Z(n52206) );
  XOR2_X1 U28452 ( .A1(n58905), .A2(n23886), .Z(Plaintext[51]) );
  XOR2_X1 U28461 ( .A1(n4901), .A2(n59496), .Z(n17112) );
  OR2_X1 U28464 ( .A1(n35324), .A2(n35787), .Z(n32136) );
  OAI21_X1 U28472 ( .A1(n53843), .A2(n53844), .B(n54065), .ZN(n58908) );
  XOR2_X1 U28474 ( .A1(n39385), .A2(n36322), .Z(n36323) );
  NAND2_X1 U28475 ( .A1(n37185), .A2(n24661), .ZN(n60942) );
  NAND2_X2 U28478 ( .A1(n35031), .A2(n15144), .ZN(n5927) );
  NAND2_X2 U28480 ( .A1(n59582), .A2(n25450), .ZN(n7693) );
  NAND2_X2 U28486 ( .A1(n1235), .A2(n36821), .ZN(n10550) );
  INV_X2 U28490 ( .I(n58910), .ZN(n25376) );
  XOR2_X1 U28492 ( .A1(n38987), .A2(n38979), .Z(n12611) );
  INV_X2 U28501 ( .I(n58913), .ZN(n50305) );
  NAND2_X2 U28502 ( .A1(n58914), .A2(n16358), .ZN(n37917) );
  XOR2_X1 U28506 ( .A1(n58916), .A2(n15881), .Z(n25288) );
  NAND2_X2 U28509 ( .A1(n2089), .A2(n9590), .ZN(n40631) );
  XOR2_X1 U28531 ( .A1(n19753), .A2(n25845), .Z(n58921) );
  XOR2_X1 U28532 ( .A1(n58922), .A2(n4558), .Z(n5023) );
  XOR2_X1 U28535 ( .A1(n5451), .A2(n61661), .Z(n58922) );
  XOR2_X1 U28536 ( .A1(n21022), .A2(n58923), .Z(n25823) );
  XOR2_X1 U28538 ( .A1(n45885), .A2(n57240), .Z(n58923) );
  NAND2_X1 U28541 ( .A1(n9289), .A2(n33005), .ZN(n59138) );
  NAND3_X2 U28565 ( .A1(n29464), .A2(n29466), .A3(n29465), .ZN(n10057) );
  XOR2_X1 U28589 ( .A1(n31600), .A2(n32035), .Z(n31673) );
  XOR2_X1 U28591 ( .A1(n58932), .A2(n53262), .Z(Plaintext[14]) );
  NOR2_X2 U28612 ( .A1(n19735), .A2(n23956), .ZN(n23411) );
  AOI22_X1 U28640 ( .A1(n53304), .A2(n59907), .B1(n53307), .B2(n53306), .ZN(
        n19317) );
  NOR2_X2 U28645 ( .A1(n46718), .A2(n58937), .ZN(n50395) );
  NAND3_X2 U28648 ( .A1(n18631), .A2(n18632), .A3(n18630), .ZN(n58937) );
  NAND2_X2 U28650 ( .A1(n16746), .A2(n58939), .ZN(n13884) );
  NAND2_X1 U28657 ( .A1(n36752), .A2(n36753), .ZN(n10493) );
  NAND3_X2 U28680 ( .A1(n40043), .A2(n40042), .A3(n40044), .ZN(n59165) );
  NAND2_X2 U28691 ( .A1(n33607), .A2(n36195), .ZN(n36109) );
  NOR2_X2 U28697 ( .A1(n55), .A2(n16968), .ZN(n33607) );
  NOR2_X2 U28705 ( .A1(n58941), .A2(n58940), .ZN(n59239) );
  INV_X2 U28707 ( .I(n4632), .ZN(n58941) );
  AOI22_X1 U28708 ( .A1(n53566), .A2(n21743), .B1(n53561), .B2(n53411), .ZN(
        n53412) );
  NOR3_X2 U28711 ( .A1(n22180), .A2(n12816), .A3(n13088), .ZN(n58943) );
  NOR2_X2 U28717 ( .A1(n15738), .A2(n10888), .ZN(n30759) );
  NOR2_X2 U28730 ( .A1(n29472), .A2(n30430), .ZN(n31073) );
  AOI21_X2 U28731 ( .A1(n27000), .A2(n24476), .B(n20771), .ZN(n31077) );
  NOR2_X2 U28744 ( .A1(n55680), .A2(n55456), .ZN(n55976) );
  XOR2_X1 U28745 ( .A1(n43425), .A2(n292), .Z(n18993) );
  BUF_X4 U28746 ( .I(n42894), .Z(n61237) );
  NAND4_X2 U28754 ( .A1(n6907), .A2(n35085), .A3(n6910), .A4(n6909), .ZN(
        n16025) );
  XOR2_X1 U28762 ( .A1(n58946), .A2(n60532), .Z(n12543) );
  XOR2_X1 U28764 ( .A1(n3665), .A2(n38818), .Z(n58946) );
  XOR2_X1 U28769 ( .A1(n11737), .A2(n52442), .Z(n11860) );
  XOR2_X1 U28773 ( .A1(n58947), .A2(n51989), .Z(n52007) );
  NAND4_X1 U28778 ( .A1(n56055), .A2(n56057), .A3(n56054), .A4(n56056), .ZN(
        n56079) );
  NOR2_X2 U28785 ( .A1(n3091), .A2(n48521), .ZN(n48503) );
  XOR2_X1 U28809 ( .A1(n31407), .A2(n21128), .Z(n30400) );
  NOR2_X2 U28821 ( .A1(n49451), .A2(n49842), .ZN(n48980) );
  NAND3_X2 U28851 ( .A1(n18080), .A2(n60674), .A3(n18078), .ZN(n51213) );
  NOR2_X2 U28854 ( .A1(n60209), .A2(n9229), .ZN(n50000) );
  NAND2_X2 U28856 ( .A1(n60209), .A2(n16336), .ZN(n7972) );
  NAND2_X2 U28867 ( .A1(n8211), .A2(n20391), .ZN(n31211) );
  AOI21_X2 U28869 ( .A1(n60767), .A2(n29645), .B(n28597), .ZN(n28599) );
  XOR2_X1 U28880 ( .A1(n8792), .A2(n2406), .Z(n59131) );
  NAND2_X2 U28894 ( .A1(n50006), .A2(n48228), .ZN(n50358) );
  OR2_X1 U28895 ( .A1(n18322), .A2(n21159), .Z(n29421) );
  XOR2_X1 U28907 ( .A1(n58954), .A2(n63031), .Z(n2361) );
  INV_X2 U28912 ( .I(n42822), .ZN(n42827) );
  BUF_X2 U28924 ( .I(n1362), .Z(n58955) );
  NOR2_X2 U28942 ( .A1(n22464), .A2(n47186), .ZN(n48239) );
  XOR2_X1 U28947 ( .A1(n5951), .A2(n58957), .Z(n5950) );
  NOR2_X2 U28951 ( .A1(n8790), .A2(n8679), .ZN(n8789) );
  NAND2_X1 U28952 ( .A1(n47318), .A2(n47319), .ZN(n58958) );
  NAND2_X1 U28954 ( .A1(n9731), .A2(n53351), .ZN(n53339) );
  NAND2_X2 U28963 ( .A1(n13659), .A2(n53873), .ZN(n13939) );
  INV_X4 U28973 ( .I(n58959), .ZN(n23215) );
  NOR2_X2 U28981 ( .A1(n2883), .A2(n7817), .ZN(n58959) );
  INV_X1 U28985 ( .I(n21751), .ZN(n34337) );
  OR2_X1 U28986 ( .A1(n21751), .A2(n25256), .Z(n10072) );
  NAND2_X2 U28987 ( .A1(n59057), .A2(n26059), .ZN(n36233) );
  INV_X2 U28989 ( .I(n24731), .ZN(n24733) );
  NOR2_X2 U29019 ( .A1(n23003), .A2(n42598), .ZN(n42606) );
  INV_X1 U29033 ( .I(n12379), .ZN(n14836) );
  XOR2_X1 U29047 ( .A1(n32585), .A2(n58962), .Z(n31490) );
  XOR2_X1 U29054 ( .A1(n31487), .A2(n45126), .Z(n58962) );
  NAND2_X2 U29063 ( .A1(n3597), .A2(n47670), .ZN(n47863) );
  XOR2_X1 U29068 ( .A1(n56097), .A2(n53477), .Z(n60692) );
  OAI22_X1 U29079 ( .A1(n36046), .A2(n7028), .B1(n36777), .B2(n17096), .ZN(
        n36047) );
  XOR2_X1 U29091 ( .A1(n14038), .A2(n2747), .Z(n13989) );
  INV_X1 U29094 ( .I(n45544), .ZN(n61332) );
  NAND2_X2 U29104 ( .A1(n11959), .A2(n38672), .ZN(n22304) );
  XOR2_X1 U29109 ( .A1(n58967), .A2(n18069), .Z(n5000) );
  XOR2_X1 U29114 ( .A1(n42591), .A2(n11317), .Z(n58967) );
  NAND3_X2 U29115 ( .A1(n27282), .A2(n1355), .A3(n22351), .ZN(n28560) );
  NOR2_X2 U29124 ( .A1(n44453), .A2(n44451), .ZN(n44457) );
  XOR2_X1 U29155 ( .A1(n7058), .A2(n31341), .Z(n31809) );
  NAND3_X2 U29157 ( .A1(n6820), .A2(n28740), .A3(n16085), .ZN(n31341) );
  NAND3_X1 U29158 ( .A1(n41511), .A2(n37924), .A3(n60213), .ZN(n37930) );
  NAND2_X2 U29166 ( .A1(n38021), .A2(n1410), .ZN(n40272) );
  XOR2_X1 U29195 ( .A1(n6057), .A2(n5824), .Z(n6055) );
  INV_X2 U29198 ( .I(n30620), .ZN(n30608) );
  NAND2_X1 U29203 ( .A1(n59268), .A2(n30620), .ZN(n29077) );
  XNOR2_X1 U29206 ( .A1(n39722), .A2(n37099), .ZN(n61160) );
  NAND2_X2 U29210 ( .A1(n8225), .A2(n25166), .ZN(n59695) );
  INV_X2 U29215 ( .I(n37374), .ZN(n1769) );
  NAND2_X2 U29216 ( .A1(n24634), .A2(n24635), .ZN(n37374) );
  XOR2_X1 U29217 ( .A1(n22979), .A2(n13831), .Z(n51136) );
  NAND2_X2 U29218 ( .A1(n36790), .A2(n36793), .ZN(n36813) );
  NAND2_X2 U29225 ( .A1(n50081), .A2(n50400), .ZN(n49425) );
  NAND2_X2 U29236 ( .A1(n13260), .A2(n49422), .ZN(n52446) );
  NOR2_X1 U29238 ( .A1(n11691), .A2(n57466), .ZN(n60278) );
  INV_X4 U29239 ( .I(n4437), .ZN(n15252) );
  NAND2_X2 U29241 ( .A1(n11854), .A2(n12189), .ZN(n4437) );
  AND2_X1 U29242 ( .A1(n58105), .A2(n57546), .Z(n35199) );
  NAND2_X1 U29244 ( .A1(n46732), .A2(n18590), .ZN(n46733) );
  NAND2_X2 U29250 ( .A1(n43726), .A2(n9046), .ZN(n18590) );
  NAND2_X1 U29256 ( .A1(n30285), .A2(n61734), .ZN(n29041) );
  NOR2_X2 U29262 ( .A1(n48082), .A2(n46770), .ZN(n48080) );
  NAND3_X1 U29272 ( .A1(n54810), .A2(n54809), .A3(n1146), .ZN(n58976) );
  BUF_X2 U29297 ( .I(n54802), .Z(n58978) );
  XOR2_X1 U29302 ( .A1(n17898), .A2(n46637), .Z(n46646) );
  NAND2_X1 U29337 ( .A1(n28914), .A2(n22262), .ZN(n59175) );
  NAND2_X1 U29339 ( .A1(n55066), .A2(n54960), .ZN(n55047) );
  OR3_X1 U29346 ( .A1(n40550), .A2(n21377), .A3(n9334), .Z(n41557) );
  NAND2_X2 U29354 ( .A1(n23763), .A2(n55400), .ZN(n54983) );
  NAND2_X2 U29356 ( .A1(n34734), .A2(n64812), .ZN(n34260) );
  AND2_X1 U29358 ( .A1(n34447), .A2(n1221), .Z(n34443) );
  NOR2_X2 U29385 ( .A1(n5024), .A2(n23266), .ZN(n6015) );
  NOR2_X2 U29386 ( .A1(n58984), .A2(n19064), .ZN(n18352) );
  XOR2_X1 U29387 ( .A1(n37793), .A2(n37792), .Z(n2850) );
  XOR2_X1 U29388 ( .A1(n38992), .A2(n18057), .Z(n37793) );
  NOR2_X1 U29391 ( .A1(n59473), .A2(n33332), .ZN(n58985) );
  AOI21_X2 U29405 ( .A1(n45627), .A2(n60893), .B(n58987), .ZN(n45628) );
  XOR2_X1 U29412 ( .A1(n32184), .A2(n32544), .Z(n12813) );
  OR2_X1 U29416 ( .A1(n1734), .A2(n41851), .Z(n59267) );
  NAND2_X1 U29427 ( .A1(n55644), .A2(n58463), .ZN(n52299) );
  NAND2_X2 U29432 ( .A1(n13038), .A2(n25857), .ZN(n49510) );
  NAND2_X1 U29434 ( .A1(n40025), .A2(n6932), .ZN(n40293) );
  AOI21_X1 U29442 ( .A1(n34866), .A2(n58990), .B(n34865), .ZN(n34868) );
  NAND3_X1 U29448 ( .A1(n20915), .A2(n37028), .A3(n37027), .ZN(n58990) );
  XOR2_X1 U29459 ( .A1(n30977), .A2(n11026), .Z(n31315) );
  NOR2_X2 U29461 ( .A1(n4620), .A2(n47486), .ZN(n4619) );
  XOR2_X1 U29480 ( .A1(n39270), .A2(n8204), .Z(n61494) );
  NAND2_X1 U29482 ( .A1(n28592), .A2(n28591), .ZN(n28600) );
  NOR2_X1 U29489 ( .A1(n58995), .A2(n11017), .ZN(n22027) );
  XOR2_X1 U29502 ( .A1(n10409), .A2(n24698), .Z(n31640) );
  NAND2_X1 U29523 ( .A1(n54054), .A2(n53407), .ZN(n58997) );
  AOI22_X1 U29524 ( .A1(n13149), .A2(n49884), .B1(n13148), .B2(n49883), .ZN(
        n13147) );
  BUF_X2 U29525 ( .I(n7517), .Z(n58998) );
  INV_X2 U29527 ( .I(n44388), .ZN(n60701) );
  XOR2_X1 U29536 ( .A1(n51243), .A2(n1140), .Z(n59000) );
  XNOR2_X1 U29555 ( .A1(n37581), .A2(n37875), .ZN(n15425) );
  NOR2_X2 U29565 ( .A1(n1716), .A2(n42585), .ZN(n8619) );
  NAND2_X2 U29585 ( .A1(n22123), .A2(n59006), .ZN(n54717) );
  XOR2_X1 U29603 ( .A1(n21244), .A2(n21243), .Z(n23505) );
  OR2_X1 U29612 ( .A1(n13525), .A2(n42239), .Z(n40559) );
  XOR2_X1 U29615 ( .A1(n52145), .A2(n61305), .Z(n10826) );
  XOR2_X1 U29622 ( .A1(n10476), .A2(n52559), .Z(n52145) );
  OAI21_X1 U29624 ( .A1(n18229), .A2(n54537), .B(n18422), .ZN(n54538) );
  NAND2_X2 U29626 ( .A1(n54565), .A2(n54561), .ZN(n18229) );
  NAND2_X2 U29628 ( .A1(n24501), .A2(n59012), .ZN(n50218) );
  NAND3_X1 U29634 ( .A1(n47172), .A2(n47173), .A3(n47171), .ZN(n59012) );
  AND2_X1 U29641 ( .A1(n10699), .A2(n34164), .Z(n60164) );
  NAND2_X2 U29646 ( .A1(n59056), .A2(n8012), .ZN(n47014) );
  INV_X2 U29657 ( .I(n59014), .ZN(n24420) );
  XOR2_X1 U29663 ( .A1(Ciphertext[93]), .A2(Key[160]), .Z(n59014) );
  NAND2_X1 U29664 ( .A1(n59491), .A2(n4250), .ZN(n1942) );
  INV_X2 U29669 ( .I(n59017), .ZN(n7175) );
  XNOR2_X1 U29671 ( .A1(n17378), .A2(n23998), .ZN(n59017) );
  BUF_X2 U29672 ( .I(n21493), .Z(n59019) );
  XOR2_X1 U29702 ( .A1(n38385), .A2(n38384), .Z(n59023) );
  XOR2_X1 U29703 ( .A1(n59024), .A2(n57314), .Z(n952) );
  XOR2_X1 U29711 ( .A1(n37550), .A2(n18428), .Z(n59024) );
  AOI22_X2 U29727 ( .A1(n1405), .A2(n1507), .B1(n59026), .B2(n58367), .ZN(
        n40717) );
  NAND2_X1 U29734 ( .A1(n59028), .A2(n48468), .ZN(n47207) );
  OR3_X1 U29744 ( .A1(n47204), .A2(n7186), .A3(n48460), .Z(n59028) );
  AND2_X2 U29746 ( .A1(n48612), .A2(n24519), .Z(n48626) );
  XOR2_X1 U29749 ( .A1(n37576), .A2(n37575), .Z(n19531) );
  XOR2_X1 U29750 ( .A1(n59029), .A2(n3600), .Z(n3602) );
  NOR2_X2 U29773 ( .A1(n52840), .A2(n52756), .ZN(n52836) );
  AND2_X1 U29780 ( .A1(n53604), .A2(n11997), .Z(n1160) );
  XOR2_X1 U29784 ( .A1(n59032), .A2(n60483), .Z(n60482) );
  NOR3_X2 U29786 ( .A1(n55068), .A2(n25220), .A3(n55096), .ZN(n55066) );
  NOR2_X2 U29787 ( .A1(n12725), .A2(n8337), .ZN(n45900) );
  XOR2_X1 U29800 ( .A1(n4031), .A2(n59188), .Z(n10784) );
  NOR2_X2 U29803 ( .A1(n23875), .A2(n41146), .ZN(n41155) );
  INV_X2 U29804 ( .I(n3685), .ZN(n41146) );
  XOR2_X1 U29807 ( .A1(n59036), .A2(n52562), .Z(n59905) );
  XOR2_X1 U29813 ( .A1(n2257), .A2(n52550), .Z(n59036) );
  NAND4_X2 U29819 ( .A1(n16520), .A2(n1083), .A3(n46109), .A4(n4448), .ZN(
        n16815) );
  XOR2_X1 U29827 ( .A1(n21598), .A2(n59039), .Z(n21597) );
  OR2_X2 U29829 ( .A1(n26000), .A2(n12003), .Z(n5713) );
  NAND2_X2 U29843 ( .A1(n20162), .A2(n48659), .ZN(n47000) );
  AND2_X2 U29858 ( .A1(n23505), .A2(n52476), .Z(n21268) );
  NAND3_X1 U29859 ( .A1(n8211), .A2(n30631), .A3(n59096), .ZN(n4764) );
  XOR2_X1 U29860 ( .A1(n59045), .A2(n46407), .Z(n24639) );
  NAND2_X2 U29869 ( .A1(n25617), .A2(n262), .ZN(n34129) );
  XOR2_X1 U29878 ( .A1(n22059), .A2(n22058), .Z(n59053) );
  NAND3_X2 U29911 ( .A1(n30864), .A2(n30865), .A3(n1353), .ZN(n11532) );
  BUF_X2 U29921 ( .I(n45992), .Z(n59059) );
  BUF_X2 U29943 ( .I(n15705), .Z(n59063) );
  INV_X2 U29944 ( .I(n59064), .ZN(n15144) );
  AOI21_X1 U29951 ( .A1(n1685), .A2(n42745), .B(n59065), .ZN(n6424) );
  BUF_X2 U29952 ( .I(n1335), .Z(n59067) );
  OAI21_X2 U29954 ( .A1(n6405), .A2(n31122), .B(n120), .ZN(n5247) );
  XOR2_X1 U29955 ( .A1(n59068), .A2(n59665), .Z(n7099) );
  XOR2_X1 U29956 ( .A1(n38206), .A2(n37072), .Z(n59068) );
  XOR2_X1 U29960 ( .A1(n31344), .A2(n33139), .Z(n25042) );
  NAND2_X2 U29961 ( .A1(n18337), .A2(n30563), .ZN(n31344) );
  NAND3_X2 U29963 ( .A1(n14495), .A2(n14478), .A3(n14497), .ZN(n14477) );
  XOR2_X1 U29964 ( .A1(n59069), .A2(n56976), .Z(Plaintext[185]) );
  BUF_X2 U29983 ( .I(n47156), .Z(n59071) );
  XOR2_X1 U30006 ( .A1(n12771), .A2(n46174), .Z(n59072) );
  NAND2_X2 U30026 ( .A1(n48126), .A2(n1479), .ZN(n8138) );
  XOR2_X1 U30029 ( .A1(n59075), .A2(n1976), .Z(n1973) );
  NAND2_X2 U30034 ( .A1(n36233), .A2(n32610), .ZN(n10317) );
  AOI21_X2 U30035 ( .A1(n1380), .A2(n48757), .B(n50426), .ZN(n14642) );
  NAND3_X2 U30037 ( .A1(n50281), .A2(n50280), .A3(n50282), .ZN(n51797) );
  NAND2_X2 U30044 ( .A1(n33540), .A2(n13942), .ZN(n59078) );
  OR2_X1 U30061 ( .A1(n54941), .A2(n59081), .Z(n59080) );
  INV_X2 U30066 ( .I(n26097), .ZN(n26095) );
  NOR2_X1 U30070 ( .A1(n30145), .A2(n19598), .ZN(n30709) );
  NAND3_X2 U30082 ( .A1(n26858), .A2(n26857), .A3(n26859), .ZN(n19598) );
  INV_X2 U30084 ( .I(n59082), .ZN(n61658) );
  OAI22_X1 U30086 ( .A1(n30137), .A2(n12871), .B1(n13531), .B2(n30136), .ZN(
        n30138) );
  NAND2_X1 U30089 ( .A1(n59248), .A2(n10711), .ZN(n59088) );
  OAI21_X1 U30091 ( .A1(n59090), .A2(n555), .B(n59089), .ZN(n28592) );
  NAND3_X1 U30095 ( .A1(n7150), .A2(n33507), .A3(n59091), .ZN(n10047) );
  NAND2_X1 U30097 ( .A1(n33497), .A2(n8431), .ZN(n59091) );
  NAND2_X2 U30107 ( .A1(n21468), .A2(n22528), .ZN(n4046) );
  NOR2_X2 U30112 ( .A1(n24558), .A2(n47266), .ZN(n46885) );
  NAND3_X2 U30114 ( .A1(n17538), .A2(n25256), .A3(n34268), .ZN(n8800) );
  NOR2_X1 U30121 ( .A1(n17666), .A2(n19554), .ZN(n17665) );
  NAND2_X2 U30123 ( .A1(n24933), .A2(n2795), .ZN(n22513) );
  XOR2_X1 U30130 ( .A1(n59097), .A2(n981), .Z(n6577) );
  XOR2_X1 U30132 ( .A1(n4854), .A2(n39189), .Z(n59097) );
  XOR2_X1 U30135 ( .A1(n59098), .A2(n36992), .Z(n9217) );
  XOR2_X1 U30136 ( .A1(n7573), .A2(n819), .Z(n59098) );
  AOI22_X2 U30156 ( .A1(n53193), .A2(n53192), .B1(n53190), .B2(n59649), .ZN(
        n53203) );
  NOR2_X2 U30159 ( .A1(n14773), .A2(n1518), .ZN(n59199) );
  NAND2_X2 U30160 ( .A1(n59103), .A2(n7500), .ZN(n17661) );
  NAND2_X1 U30165 ( .A1(n36372), .A2(n36558), .ZN(n20855) );
  NAND2_X2 U30166 ( .A1(n8356), .A2(n1339), .ZN(n36558) );
  NOR2_X1 U30178 ( .A1(n43210), .A2(n43212), .ZN(n59437) );
  AOI21_X2 U30181 ( .A1(n36572), .A2(n8356), .B(n25261), .ZN(n59105) );
  NAND2_X2 U30183 ( .A1(n10288), .A2(n14678), .ZN(n59106) );
  NAND2_X1 U30187 ( .A1(n45965), .A2(n45964), .ZN(n59107) );
  NAND2_X2 U30189 ( .A1(n19451), .A2(n11987), .ZN(n12300) );
  XOR2_X1 U30194 ( .A1(n59109), .A2(n24140), .Z(n9285) );
  XOR2_X1 U30196 ( .A1(n18854), .A2(n21133), .Z(n13755) );
  XOR2_X1 U30197 ( .A1(n59110), .A2(n21700), .Z(n51130) );
  OR2_X1 U30208 ( .A1(n4277), .A2(n9511), .Z(n4276) );
  NAND2_X2 U30214 ( .A1(n18482), .A2(n43701), .ZN(n9511) );
  AND2_X2 U30215 ( .A1(n3055), .A2(n15394), .Z(n49649) );
  XOR2_X1 U30216 ( .A1(n15704), .A2(n15309), .Z(n37863) );
  NOR2_X2 U30221 ( .A1(n59113), .A2(n3119), .ZN(n25794) );
  NAND3_X2 U30222 ( .A1(n49654), .A2(n22682), .A3(n49652), .ZN(n59113) );
  NOR2_X2 U30238 ( .A1(n26273), .A2(n26274), .ZN(n59115) );
  NOR2_X2 U30240 ( .A1(n54037), .A2(n23217), .ZN(n21919) );
  XOR2_X1 U30246 ( .A1(n10677), .A2(n10552), .Z(n9083) );
  NAND2_X2 U30248 ( .A1(n20275), .A2(n5961), .ZN(n59116) );
  XOR2_X1 U30249 ( .A1(n51163), .A2(n51164), .Z(n59572) );
  XOR2_X1 U30250 ( .A1(n51036), .A2(n50833), .Z(n51164) );
  AOI22_X1 U30253 ( .A1(n93), .A2(n15829), .B1(n28240), .B2(n28073), .ZN(
        n28074) );
  NOR2_X2 U30256 ( .A1(n12410), .A2(n12409), .ZN(n40980) );
  NAND2_X1 U30268 ( .A1(n59860), .A2(n59120), .ZN(n5336) );
  OAI21_X2 U30269 ( .A1(n51213), .A2(n2222), .B(n2221), .ZN(n10510) );
  NAND3_X2 U30274 ( .A1(n3854), .A2(n41520), .A3(n41521), .ZN(n301) );
  AOI21_X2 U30280 ( .A1(n59239), .A2(n59238), .B(n10341), .ZN(n60783) );
  INV_X1 U30283 ( .I(n59126), .ZN(n5042) );
  OAI21_X1 U30285 ( .A1(n59128), .A2(n59127), .B(n45672), .ZN(n59126) );
  NOR2_X1 U30292 ( .A1(n45673), .A2(n46885), .ZN(n59128) );
  NOR2_X1 U30296 ( .A1(n53732), .A2(n16489), .ZN(n53715) );
  INV_X4 U30297 ( .I(n36394), .ZN(n60196) );
  NOR3_X1 U30298 ( .A1(n60890), .A2(n26946), .A3(n28137), .ZN(n26950) );
  BUF_X2 U30300 ( .I(n30558), .Z(n59129) );
  NAND2_X2 U30307 ( .A1(n15346), .A2(n54616), .ZN(n54783) );
  XOR2_X1 U30310 ( .A1(n16095), .A2(n57336), .Z(n2486) );
  XOR2_X1 U30313 ( .A1(n22032), .A2(n6363), .Z(n16095) );
  XOR2_X1 U30320 ( .A1(n2407), .A2(n59131), .Z(n2409) );
  XOR2_X1 U30321 ( .A1(n31200), .A2(n31641), .Z(n33914) );
  INV_X1 U30322 ( .I(n59136), .ZN(n59135) );
  NAND2_X1 U30323 ( .A1(n35490), .A2(n25671), .ZN(n59136) );
  NAND2_X2 U30343 ( .A1(n31275), .A2(n31274), .ZN(n6321) );
  NAND2_X1 U30350 ( .A1(n14941), .A2(n29615), .ZN(n61618) );
  XOR2_X1 U30356 ( .A1(n10285), .A2(n5913), .Z(n9820) );
  XOR2_X1 U30379 ( .A1(n7862), .A2(n12890), .Z(n38923) );
  XOR2_X1 U30390 ( .A1(n45053), .A2(n45054), .Z(n45055) );
  AOI21_X1 U30397 ( .A1(n54576), .A2(n54577), .B(n54575), .ZN(n54578) );
  NOR2_X2 U30403 ( .A1(n26641), .A2(n20437), .ZN(n27594) );
  XOR2_X1 U30407 ( .A1(n3480), .A2(n24170), .Z(n19441) );
  NAND2_X2 U30409 ( .A1(n26172), .A2(n26171), .ZN(n24170) );
  NAND2_X2 U30411 ( .A1(n54035), .A2(n53905), .ZN(n54036) );
  OR2_X1 U30413 ( .A1(n60883), .A2(n33759), .Z(n34792) );
  AND3_X1 U30428 ( .A1(n42398), .A2(n42396), .A3(n42397), .Z(n18344) );
  NOR2_X1 U30429 ( .A1(n10125), .A2(n27668), .ZN(n27838) );
  NAND2_X1 U30430 ( .A1(n54043), .A2(n54044), .ZN(n60043) );
  NAND2_X1 U30435 ( .A1(n47287), .A2(n47286), .ZN(n3661) );
  NAND2_X1 U30438 ( .A1(n59146), .A2(n39970), .ZN(n39971) );
  NAND2_X1 U30439 ( .A1(n39968), .A2(n14132), .ZN(n59146) );
  NOR2_X2 U30455 ( .A1(n59150), .A2(n42630), .ZN(n41706) );
  NAND2_X2 U30462 ( .A1(n14263), .A2(n43090), .ZN(n44453) );
  XOR2_X1 U30469 ( .A1(n31809), .A2(n10229), .Z(n24911) );
  NAND2_X1 U30471 ( .A1(n29797), .A2(n9281), .ZN(n59151) );
  XOR2_X1 U30478 ( .A1(n50034), .A2(n50033), .Z(n50035) );
  NAND3_X1 U30480 ( .A1(n61174), .A2(n54585), .A3(n24489), .ZN(n7525) );
  NAND2_X2 U30481 ( .A1(n30695), .A2(n58999), .ZN(n31049) );
  NAND2_X2 U30482 ( .A1(n4619), .A2(n59153), .ZN(n4534) );
  XOR2_X1 U30488 ( .A1(n37581), .A2(n50494), .Z(n38203) );
  INV_X2 U30490 ( .I(n15246), .ZN(n59154) );
  XOR2_X1 U30498 ( .A1(n36685), .A2(n23493), .Z(n59663) );
  NAND3_X1 U30503 ( .A1(n59155), .A2(n7094), .A3(n42454), .ZN(n17185) );
  NAND4_X1 U30512 ( .A1(n59156), .A2(n42792), .A3(n43956), .A4(n59709), .ZN(
        n42797) );
  NOR3_X2 U30514 ( .A1(n56808), .A2(n56817), .A3(n56796), .ZN(n56790) );
  INV_X2 U30518 ( .I(n51461), .ZN(n56796) );
  NAND3_X1 U30526 ( .A1(n59157), .A2(n51264), .A3(n187), .ZN(n51267) );
  NAND2_X2 U30528 ( .A1(n7721), .A2(n59158), .ZN(n753) );
  XOR2_X1 U30530 ( .A1(n26181), .A2(n59159), .Z(n18458) );
  XOR2_X1 U30531 ( .A1(n46624), .A2(n46623), .Z(n59159) );
  NOR2_X2 U30533 ( .A1(n20555), .A2(n38691), .ZN(n41199) );
  NAND2_X1 U30544 ( .A1(n20730), .A2(n48892), .ZN(n48890) );
  NOR3_X1 U30545 ( .A1(n57248), .A2(n47251), .A3(n47255), .ZN(n16176) );
  NAND2_X2 U30565 ( .A1(n23738), .A2(n49006), .ZN(n48039) );
  NOR3_X2 U30566 ( .A1(n7433), .A2(n36491), .A3(n36490), .ZN(n36504) );
  NOR2_X2 U30574 ( .A1(n23658), .A2(n28716), .ZN(n30776) );
  XOR2_X1 U30576 ( .A1(n44466), .A2(n14313), .Z(n46252) );
  NAND2_X2 U30590 ( .A1(n59481), .A2(n18472), .ZN(n29744) );
  NOR2_X2 U30594 ( .A1(n61208), .A2(n61209), .ZN(n8727) );
  NOR2_X2 U30595 ( .A1(n59165), .A2(n40046), .ZN(n40096) );
  XOR2_X1 U30599 ( .A1(n3379), .A2(n3380), .Z(n59166) );
  NOR2_X1 U30603 ( .A1(n56572), .A2(n8367), .ZN(n15179) );
  BUF_X4 U30609 ( .I(n15727), .Z(n60162) );
  INV_X2 U30610 ( .I(n59168), .ZN(n14863) );
  XOR2_X1 U30614 ( .A1(n14864), .A2(n38335), .Z(n59168) );
  OAI22_X1 U30619 ( .A1(n15269), .A2(n17000), .B1(n29427), .B2(n29059), .ZN(
        n59169) );
  AOI21_X2 U30624 ( .A1(n42541), .A2(n61171), .B(n3980), .ZN(n3969) );
  NOR2_X2 U30627 ( .A1(n43039), .A2(n12965), .ZN(n3980) );
  XOR2_X1 U30629 ( .A1(n59173), .A2(n59172), .Z(n3735) );
  XOR2_X1 U30635 ( .A1(n13015), .A2(n24794), .Z(n59173) );
  NOR2_X2 U30643 ( .A1(n59175), .A2(n25506), .ZN(n31989) );
  NAND3_X2 U30659 ( .A1(n25265), .A2(n25264), .A3(n48119), .ZN(n59176) );
  NAND3_X2 U30660 ( .A1(n60681), .A2(n43576), .A3(n2690), .ZN(n2293) );
  NOR2_X2 U30663 ( .A1(n59983), .A2(n12226), .ZN(n12229) );
  OR2_X1 U30671 ( .A1(n61475), .A2(n22002), .Z(n43165) );
  NAND2_X1 U30679 ( .A1(n4641), .A2(n57168), .ZN(n35291) );
  NAND2_X2 U30683 ( .A1(n59181), .A2(n3857), .ZN(n36246) );
  NOR2_X2 U30687 ( .A1(n6581), .A2(n40987), .ZN(n59183) );
  NAND3_X2 U30689 ( .A1(n18042), .A2(n18041), .A3(n18043), .ZN(n43844) );
  NAND3_X2 U30692 ( .A1(n5873), .A2(n59924), .A3(n4798), .ZN(n36687) );
  XOR2_X1 U30709 ( .A1(n59186), .A2(n5240), .Z(n7096) );
  XOR2_X1 U30712 ( .A1(n16028), .A2(n18513), .Z(n59186) );
  NAND2_X1 U30716 ( .A1(n40711), .A2(n40710), .ZN(n59817) );
  XOR2_X1 U30727 ( .A1(n51302), .A2(n51301), .Z(n59188) );
  NAND2_X1 U30728 ( .A1(n47424), .A2(n47423), .ZN(n60399) );
  AND2_X2 U30753 ( .A1(n19716), .A2(n5348), .Z(n52281) );
  NAND2_X2 U30757 ( .A1(n212), .A2(n1226), .ZN(n4632) );
  NOR3_X2 U30763 ( .A1(n1970), .A2(n28471), .A3(n27810), .ZN(n28475) );
  XOR2_X1 U30777 ( .A1(n39696), .A2(n2770), .Z(n37059) );
  OAI21_X2 U30787 ( .A1(n5773), .A2(n20180), .B(n41715), .ZN(n42110) );
  AND2_X1 U30791 ( .A1(n35351), .A2(n59208), .Z(n15594) );
  NOR2_X2 U30797 ( .A1(n10236), .A2(n23596), .ZN(n28852) );
  XOR2_X1 U30802 ( .A1(n31463), .A2(n18595), .Z(n59209) );
  OR2_X2 U30807 ( .A1(n19695), .A2(n59210), .Z(n15982) );
  NAND4_X1 U30811 ( .A1(n19001), .A2(n30581), .A3(n61913), .A4(n31094), .ZN(
        n59210) );
  OAI21_X2 U30812 ( .A1(n59211), .A2(n4794), .B(n58369), .ZN(n22348) );
  INV_X1 U30815 ( .I(n19918), .ZN(n59335) );
  XOR2_X1 U30820 ( .A1(n59212), .A2(n15464), .Z(n30974) );
  XOR2_X1 U30821 ( .A1(n23424), .A2(n8329), .Z(n59212) );
  NOR2_X1 U30838 ( .A1(n30160), .A2(n30689), .ZN(n59214) );
  XOR2_X1 U30839 ( .A1(n59215), .A2(n4782), .Z(n40947) );
  XOR2_X1 U30843 ( .A1(n38131), .A2(n37386), .Z(n59215) );
  XOR2_X1 U30847 ( .A1(n7971), .A2(n12002), .Z(n43797) );
  NAND2_X1 U30856 ( .A1(n27437), .A2(n57306), .ZN(n27439) );
  NAND3_X2 U30876 ( .A1(n29708), .A2(n8087), .A3(n29707), .ZN(n29716) );
  NAND2_X2 U30877 ( .A1(n59728), .A2(n52681), .ZN(n56897) );
  OAI21_X2 U30894 ( .A1(n15745), .A2(n59650), .B(n59217), .ZN(n318) );
  NAND2_X2 U30895 ( .A1(n39936), .A2(n521), .ZN(n59217) );
  NOR2_X1 U30897 ( .A1(n30271), .A2(n61734), .ZN(n30277) );
  NAND2_X1 U30905 ( .A1(n59221), .A2(n61929), .ZN(n35091) );
  NAND2_X1 U30912 ( .A1(n7600), .A2(n23651), .ZN(n59221) );
  XOR2_X1 U30914 ( .A1(n44524), .A2(n59222), .Z(n44551) );
  NAND3_X1 U30932 ( .A1(n50219), .A2(n1262), .A3(n50220), .ZN(n47994) );
  AND2_X1 U30933 ( .A1(n59224), .A2(n41116), .Z(n5584) );
  AOI22_X1 U30937 ( .A1(n62106), .A2(n15139), .B1(n59637), .B2(n41113), .ZN(
        n59224) );
  NOR2_X2 U30945 ( .A1(n19278), .A2(n22503), .ZN(n35943) );
  NOR2_X2 U30946 ( .A1(n2387), .A2(n2389), .ZN(n19278) );
  NOR3_X1 U30947 ( .A1(n18398), .A2(n62353), .A3(n43376), .ZN(n3786) );
  NAND4_X2 U30948 ( .A1(n25706), .A2(n59226), .A3(n54869), .A4(n54868), .ZN(
        n107) );
  NAND2_X2 U30957 ( .A1(n22182), .A2(n41571), .ZN(n40453) );
  AOI21_X1 U30968 ( .A1(n15837), .A2(n50409), .B(n46729), .ZN(n59227) );
  OAI21_X1 U30986 ( .A1(n27286), .A2(n27413), .B(n21086), .ZN(n27288) );
  NOR3_X2 U30988 ( .A1(n8703), .A2(n15146), .A3(n29976), .ZN(n8702) );
  NOR2_X1 U30989 ( .A1(n17937), .A2(n1373), .ZN(n17936) );
  BUF_X2 U30995 ( .I(n15171), .Z(n59229) );
  OAI21_X1 U31006 ( .A1(n11893), .A2(n20611), .B(n36926), .ZN(n59230) );
  INV_X1 U31014 ( .I(n16713), .ZN(n59231) );
  XOR2_X1 U31021 ( .A1(n22535), .A2(n59233), .Z(n15002) );
  XOR2_X1 U31026 ( .A1(n39755), .A2(n57352), .Z(n59233) );
  XOR2_X1 U31055 ( .A1(n23345), .A2(n60610), .Z(n46453) );
  XOR2_X1 U31057 ( .A1(n62399), .A2(n39659), .Z(n60897) );
  NAND4_X2 U31060 ( .A1(n36349), .A2(n36347), .A3(n36615), .A4(n36348), .ZN(
        n59236) );
  NOR2_X2 U31064 ( .A1(n47670), .A2(n6730), .ZN(n17670) );
  NAND2_X2 U31066 ( .A1(n45905), .A2(n60417), .ZN(n45897) );
  AND2_X1 U31093 ( .A1(n33599), .A2(n11060), .Z(n59240) );
  XOR2_X1 U31113 ( .A1(n65274), .A2(n59241), .Z(n11614) );
  XOR2_X1 U31114 ( .A1(n15480), .A2(n22247), .Z(n59241) );
  XNOR2_X1 U31120 ( .A1(n6425), .A2(n44385), .ZN(n15705) );
  AOI21_X1 U31122 ( .A1(n49004), .A2(n49003), .B(n11639), .ZN(n13196) );
  NAND2_X2 U31130 ( .A1(n61717), .A2(n2571), .ZN(n45596) );
  NOR2_X1 U31143 ( .A1(n3168), .A2(n30361), .ZN(n3167) );
  NAND2_X2 U31154 ( .A1(n7041), .A2(n55164), .ZN(n21389) );
  NAND3_X2 U31155 ( .A1(n27732), .A2(n27731), .A3(n27733), .ZN(n20882) );
  NOR3_X1 U31156 ( .A1(n59244), .A2(n36876), .A3(n36878), .ZN(n36879) );
  XOR2_X1 U31161 ( .A1(n33161), .A2(n31796), .Z(n32369) );
  NOR2_X2 U31164 ( .A1(n20418), .A2(n37025), .ZN(n39276) );
  XOR2_X1 U31166 ( .A1(n46625), .A2(n46307), .Z(n43935) );
  XOR2_X1 U31169 ( .A1(n46162), .A2(n43909), .Z(n46625) );
  XOR2_X1 U31170 ( .A1(n32331), .A2(n32591), .Z(n14162) );
  NAND2_X2 U31173 ( .A1(n5483), .A2(n57209), .ZN(n35443) );
  NOR3_X2 U31182 ( .A1(n40986), .A2(n40997), .A3(n5362), .ZN(n40983) );
  XOR2_X1 U31183 ( .A1(n730), .A2(n31854), .Z(n13278) );
  XOR2_X1 U31185 ( .A1(n31336), .A2(n5247), .Z(n31854) );
  NAND3_X1 U31195 ( .A1(n59249), .A2(n49899), .A3(n14315), .ZN(n48336) );
  BUF_X2 U31220 ( .I(n14462), .Z(n59252) );
  NAND2_X1 U31229 ( .A1(n10150), .A2(n38693), .ZN(n24122) );
  NAND2_X1 U31230 ( .A1(n31112), .A2(n24199), .ZN(n14272) );
  BUF_X2 U31231 ( .I(n39094), .Z(n59255) );
  XOR2_X1 U31233 ( .A1(n59431), .A2(n33289), .Z(n61575) );
  AND2_X2 U31234 ( .A1(n23155), .A2(n15795), .Z(n42263) );
  NAND3_X2 U31242 ( .A1(n22752), .A2(n52961), .A3(n52962), .ZN(n59256) );
  NOR2_X2 U31250 ( .A1(n55644), .A2(n59610), .ZN(n52298) );
  NAND2_X1 U31252 ( .A1(n21052), .A2(n50345), .ZN(n21427) );
  OAI21_X2 U31253 ( .A1(n14435), .A2(n49858), .B(n50331), .ZN(n50345) );
  NAND3_X2 U31254 ( .A1(n60880), .A2(n59258), .A3(n59257), .ZN(n25942) );
  INV_X1 U31260 ( .I(n18413), .ZN(n59257) );
  NAND2_X1 U31262 ( .A1(n18414), .A2(n18416), .ZN(n59258) );
  NAND2_X1 U31271 ( .A1(n16406), .A2(n1382), .ZN(n61327) );
  NAND2_X2 U31272 ( .A1(n5615), .A2(n25525), .ZN(n22755) );
  NOR2_X1 U31276 ( .A1(n57004), .A2(n22114), .ZN(n52873) );
  NAND2_X2 U31285 ( .A1(n30547), .A2(n30441), .ZN(n30437) );
  NAND2_X1 U31294 ( .A1(n49532), .A2(n60592), .ZN(n60591) );
  XOR2_X1 U31299 ( .A1(n50512), .A2(n21342), .Z(n59262) );
  AND2_X1 U31308 ( .A1(n14412), .A2(n14411), .Z(n59918) );
  NAND2_X2 U31312 ( .A1(n32748), .A2(n15318), .ZN(n11060) );
  XOR2_X1 U31325 ( .A1(n8556), .A2(n24090), .Z(n11555) );
  XOR2_X1 U31326 ( .A1(n20545), .A2(n52077), .Z(n52078) );
  NOR2_X1 U31328 ( .A1(n59483), .A2(n59482), .ZN(n941) );
  NOR2_X2 U31331 ( .A1(n771), .A2(n11502), .ZN(n24679) );
  XOR2_X1 U31353 ( .A1(n59264), .A2(n13883), .Z(n45021) );
  XOR2_X1 U31355 ( .A1(n44723), .A2(n51029), .Z(n59264) );
  AOI22_X2 U31362 ( .A1(n59267), .A2(n59266), .B1(n1403), .B2(n16099), .ZN(
        n18693) );
  INV_X2 U31368 ( .I(n59270), .ZN(n3935) );
  XNOR2_X1 U31370 ( .A1(n5139), .A2(n11169), .ZN(n59272) );
  INV_X2 U31377 ( .I(n59273), .ZN(n56890) );
  NOR2_X2 U31388 ( .A1(n59569), .A2(n16773), .ZN(n7204) );
  OR2_X1 U31389 ( .A1(n46337), .A2(n59276), .Z(n59275) );
  XOR2_X1 U31392 ( .A1(n38866), .A2(n38806), .Z(n18545) );
  NAND3_X2 U31397 ( .A1(n34380), .A2(n34381), .A3(n18546), .ZN(n38866) );
  NAND2_X2 U31402 ( .A1(n1787), .A2(n36026), .ZN(n34828) );
  NAND2_X2 U31411 ( .A1(n36886), .A2(n37233), .ZN(n37240) );
  XOR2_X1 U31424 ( .A1(n31655), .A2(n57365), .Z(n8333) );
  XOR2_X1 U31428 ( .A1(n65041), .A2(n59622), .Z(n31655) );
  XOR2_X1 U31437 ( .A1(n8594), .A2(n31868), .Z(n8593) );
  INV_X1 U31442 ( .I(n59724), .ZN(n34311) );
  AND2_X1 U31478 ( .A1(n30510), .A2(n4387), .Z(n59287) );
  XOR2_X1 U31479 ( .A1(n61219), .A2(n10743), .Z(n4533) );
  NAND2_X1 U31481 ( .A1(n61720), .A2(n59523), .ZN(n47686) );
  NOR4_X2 U31489 ( .A1(n41530), .A2(n41529), .A3(n41527), .A4(n41528), .ZN(
        n59289) );
  NAND4_X2 U31490 ( .A1(n32961), .A2(n32959), .A3(n61299), .A4(n35005), .ZN(
        n60516) );
  XOR2_X1 U31492 ( .A1(n12253), .A2(n17447), .Z(n12919) );
  NAND2_X2 U31499 ( .A1(n17989), .A2(n29629), .ZN(n29291) );
  BUF_X2 U31523 ( .I(n11609), .Z(n59292) );
  AOI22_X1 U31537 ( .A1(n46003), .A2(n46002), .B1(n46001), .B2(n858), .ZN(
        n46010) );
  AOI21_X2 U31538 ( .A1(n59393), .A2(n64762), .B(n28442), .ZN(n28465) );
  XOR2_X1 U31547 ( .A1(n31123), .A2(n59521), .Z(n33849) );
  OR2_X1 U31549 ( .A1(n24862), .A2(n41069), .Z(n41076) );
  NAND2_X2 U31554 ( .A1(n20153), .A2(n59297), .ZN(n20308) );
  NOR4_X2 U31560 ( .A1(n20273), .A2(n30520), .A3(n20152), .A4(n20151), .ZN(
        n59297) );
  NAND2_X2 U31565 ( .A1(n13417), .A2(n8891), .ZN(n17084) );
  NOR2_X2 U31567 ( .A1(n59299), .A2(n6574), .ZN(n48729) );
  XOR2_X1 U31569 ( .A1(n59300), .A2(n21266), .Z(Plaintext[189]) );
  AOI21_X1 U31593 ( .A1(n59303), .A2(n57233), .B(n59302), .ZN(n59301) );
  NOR2_X1 U31606 ( .A1(n57138), .A2(n57233), .ZN(n59302) );
  INV_X1 U31609 ( .I(n57137), .ZN(n59303) );
  AOI21_X1 U31620 ( .A1(n61598), .A2(n10251), .B(n157), .ZN(n32694) );
  INV_X2 U31645 ( .I(n59307), .ZN(n892) );
  XOR2_X1 U31649 ( .A1(n2172), .A2(n2174), .Z(n59307) );
  NAND3_X2 U31650 ( .A1(n5076), .A2(n4973), .A3(n14420), .ZN(n33258) );
  NAND3_X1 U31667 ( .A1(n10025), .A2(n19756), .A3(n16595), .ZN(n59310) );
  NOR2_X2 U31677 ( .A1(n1205), .A2(n6314), .ZN(n2692) );
  XOR2_X1 U31679 ( .A1(n33159), .A2(n22652), .Z(n2863) );
  NAND2_X1 U31680 ( .A1(n57610), .A2(n49462), .ZN(n5396) );
  XOR2_X1 U31689 ( .A1(n45477), .A2(n45476), .Z(n59312) );
  INV_X4 U31720 ( .I(n60630), .ZN(n55270) );
  XOR2_X1 U31733 ( .A1(n53932), .A2(n6134), .Z(n21125) );
  NOR2_X1 U31735 ( .A1(n2851), .A2(n6168), .ZN(n53932) );
  NOR2_X2 U31744 ( .A1(n3082), .A2(n34018), .ZN(n20785) );
  AOI21_X2 U31747 ( .A1(n59322), .A2(n18328), .B(n37663), .ZN(n18327) );
  XOR2_X1 U31754 ( .A1(n32307), .A2(n59323), .Z(n638) );
  XOR2_X1 U31755 ( .A1(n10645), .A2(n14249), .Z(n59323) );
  XOR2_X1 U31759 ( .A1(n59324), .A2(n17656), .Z(n4065) );
  XOR2_X1 U31760 ( .A1(n61410), .A2(n25872), .Z(n59324) );
  NOR3_X2 U31761 ( .A1(n59326), .A2(n36893), .A3(n59325), .ZN(n5525) );
  NOR2_X2 U31765 ( .A1(n31767), .A2(n33995), .ZN(n23036) );
  NOR2_X2 U31775 ( .A1(n57210), .A2(n15720), .ZN(n36706) );
  NAND3_X2 U31786 ( .A1(n34416), .A2(n34418), .A3(n34417), .ZN(n59329) );
  NOR2_X2 U31788 ( .A1(n3684), .A2(n50419), .ZN(n59690) );
  NOR3_X1 U31790 ( .A1(n63890), .A2(n30293), .A3(n29580), .ZN(n59330) );
  NAND2_X2 U31792 ( .A1(n16626), .A2(n16627), .ZN(n20620) );
  AOI22_X1 U31795 ( .A1(n15763), .A2(n3211), .B1(n28526), .B2(n28525), .ZN(
        n24909) );
  OR2_X1 U31798 ( .A1(n53162), .A2(n3285), .Z(n3284) );
  XOR2_X1 U31803 ( .A1(n59331), .A2(n31403), .Z(n26050) );
  XOR2_X1 U31808 ( .A1(n31404), .A2(n31408), .Z(n59331) );
  XOR2_X1 U31817 ( .A1(n59332), .A2(n14666), .Z(n11050) );
  XOR2_X1 U31819 ( .A1(n32002), .A2(n23869), .Z(n59332) );
  OAI21_X1 U31820 ( .A1(n59081), .A2(n22749), .B(n14469), .ZN(n54781) );
  NOR2_X2 U31821 ( .A1(n17987), .A2(n59333), .ZN(n29028) );
  XOR2_X1 U31833 ( .A1(n8596), .A2(n44397), .Z(n45343) );
  NOR2_X2 U31842 ( .A1(n19911), .A2(n19914), .ZN(n59334) );
  NAND3_X2 U31843 ( .A1(n11543), .A2(n11544), .A3(n918), .ZN(n36453) );
  NAND4_X2 U31845 ( .A1(n10967), .A2(n10962), .A3(n10964), .A4(n34896), .ZN(
        n37873) );
  NAND2_X1 U31848 ( .A1(n25080), .A2(n53848), .ZN(n53843) );
  NOR2_X1 U31851 ( .A1(n59336), .A2(n15850), .ZN(n16816) );
  NAND3_X1 U31860 ( .A1(n1858), .A2(n15407), .A3(n25157), .ZN(n30158) );
  AND2_X1 U31863 ( .A1(n13802), .A2(n2640), .Z(n60239) );
  OAI22_X1 U31872 ( .A1(n38936), .A2(n38939), .B1(n13052), .B2(n59203), .ZN(
        n59340) );
  INV_X4 U31887 ( .I(n59342), .ZN(n34335) );
  NOR2_X2 U31888 ( .A1(n19868), .A2(n34268), .ZN(n59342) );
  NAND2_X2 U31891 ( .A1(n22580), .A2(n59343), .ZN(n59515) );
  AOI22_X2 U31893 ( .A1(n33442), .A2(n33447), .B1(n31296), .B2(n34014), .ZN(
        n59343) );
  NAND2_X1 U31903 ( .A1(n59344), .A2(n64400), .ZN(n7530) );
  NAND2_X1 U31904 ( .A1(n34129), .A2(n34128), .ZN(n59348) );
  NAND2_X2 U31919 ( .A1(n59354), .A2(n24970), .ZN(n23705) );
  NOR3_X2 U31921 ( .A1(n57214), .A2(n24969), .A3(n24968), .ZN(n59354) );
  XNOR2_X1 U31922 ( .A1(n46540), .A2(n46539), .ZN(n61128) );
  XOR2_X1 U31930 ( .A1(n1906), .A2(n1905), .Z(n4216) );
  NAND2_X1 U31936 ( .A1(n9569), .A2(n20876), .ZN(n56123) );
  NOR2_X2 U31938 ( .A1(n4534), .A2(n25729), .ZN(n13042) );
  INV_X2 U31940 ( .I(n6221), .ZN(n24195) );
  NAND3_X2 U31951 ( .A1(n3492), .A2(n3491), .A3(n41313), .ZN(n6221) );
  INV_X2 U31986 ( .I(n59358), .ZN(n54105) );
  NOR2_X2 U31991 ( .A1(n53545), .A2(n53876), .ZN(n59358) );
  OAI21_X2 U31995 ( .A1(n17288), .A2(n17289), .B(n59361), .ZN(n53755) );
  NOR3_X2 U32010 ( .A1(n60201), .A2(n49933), .A3(n60400), .ZN(n59361) );
  NOR2_X1 U32012 ( .A1(n909), .A2(n22427), .ZN(n36884) );
  NAND2_X2 U32017 ( .A1(n37454), .A2(n461), .ZN(n59362) );
  INV_X1 U32019 ( .I(n12752), .ZN(n13627) );
  XOR2_X1 U32023 ( .A1(n19352), .A2(n14697), .Z(n59363) );
  NAND2_X2 U32025 ( .A1(n20170), .A2(n20171), .ZN(n30632) );
  NAND2_X2 U32029 ( .A1(n41514), .A2(n41512), .ZN(n60268) );
  NOR2_X2 U32049 ( .A1(n57328), .A2(n59364), .ZN(n3393) );
  NAND3_X2 U32051 ( .A1(n59366), .A2(n59365), .A3(n28679), .ZN(n59364) );
  NAND2_X1 U32052 ( .A1(n59467), .A2(n33746), .ZN(n33748) );
  NAND2_X2 U32061 ( .A1(n23805), .A2(n10739), .ZN(n29660) );
  NAND3_X2 U32092 ( .A1(n32535), .A2(n32534), .A3(n32533), .ZN(n36493) );
  OR2_X1 U32094 ( .A1(n18374), .A2(n49568), .Z(n18372) );
  XOR2_X1 U32113 ( .A1(n10864), .A2(n31768), .Z(n59377) );
  AND2_X2 U32137 ( .A1(n21607), .A2(n6577), .Z(n7067) );
  XOR2_X1 U32138 ( .A1(n59378), .A2(n21142), .Z(n60094) );
  XOR2_X1 U32166 ( .A1(n19389), .A2(n46241), .Z(n59378) );
  INV_X2 U32168 ( .I(n26014), .ZN(n54960) );
  BUF_X2 U32179 ( .I(n36477), .Z(n59379) );
  NAND2_X2 U32191 ( .A1(n18301), .A2(n7534), .ZN(n2331) );
  NAND2_X1 U32192 ( .A1(n20414), .A2(n54098), .ZN(n59387) );
  AOI21_X2 U32197 ( .A1(n6089), .A2(n6087), .B(n29511), .ZN(n59388) );
  NOR2_X1 U32203 ( .A1(n48718), .A2(n49881), .ZN(n48719) );
  XOR2_X1 U32221 ( .A1(n59390), .A2(n61610), .Z(n31632) );
  XOR2_X1 U32231 ( .A1(n18336), .A2(n24258), .Z(n59390) );
  AND2_X1 U32240 ( .A1(n9567), .A2(n56106), .Z(n59588) );
  NAND3_X2 U32247 ( .A1(n14986), .A2(n14982), .A3(n59391), .ZN(n15280) );
  AND3_X1 U32249 ( .A1(n41477), .A2(n61519), .A3(n14985), .Z(n59391) );
  XOR2_X1 U32251 ( .A1(n24276), .A2(n38754), .Z(n59392) );
  NOR2_X2 U32258 ( .A1(n34973), .A2(n34530), .ZN(n476) );
  NAND3_X2 U32259 ( .A1(n30673), .A2(n60750), .A3(n60749), .ZN(n33872) );
  OAI22_X2 U32262 ( .A1(n28435), .A2(n10544), .B1(n28434), .B2(n28614), .ZN(
        n59393) );
  BUF_X2 U32265 ( .I(n42407), .Z(n59394) );
  XOR2_X1 U32282 ( .A1(n59395), .A2(n22883), .Z(n8219) );
  NAND2_X2 U32286 ( .A1(n21753), .A2(n21754), .ZN(n22883) );
  BUF_X2 U32287 ( .I(n36247), .Z(n59396) );
  XOR2_X1 U32290 ( .A1(n16449), .A2(n17241), .Z(n15406) );
  NOR2_X1 U32293 ( .A1(n59399), .A2(n59397), .ZN(n18909) );
  NAND3_X2 U32297 ( .A1(n59400), .A2(n17806), .A3(n17810), .ZN(n49486) );
  OAI22_X2 U32298 ( .A1(n3958), .A2(n17949), .B1(n42751), .B2(n61812), .ZN(
        n3957) );
  XOR2_X1 U32332 ( .A1(n5435), .A2(n50817), .Z(n59402) );
  NOR3_X2 U32339 ( .A1(n19685), .A2(n19683), .A3(n59403), .ZN(n19682) );
  NOR2_X2 U32367 ( .A1(n55175), .A2(n16937), .ZN(n55176) );
  OR2_X2 U32399 ( .A1(n25292), .A2(n4673), .Z(n40995) );
  AND2_X1 U32408 ( .A1(n1232), .A2(n61361), .Z(n53258) );
  NAND2_X2 U32409 ( .A1(n6628), .A2(n38548), .ZN(n38708) );
  XOR2_X1 U32410 ( .A1(n26202), .A2(n33171), .Z(n7377) );
  XOR2_X1 U32411 ( .A1(n13778), .A2(n61464), .Z(n59417) );
  AOI21_X2 U32415 ( .A1(n40187), .A2(n40186), .B(n40185), .ZN(n45357) );
  AND2_X1 U32416 ( .A1(n18099), .A2(n4660), .Z(n4176) );
  NAND4_X2 U32423 ( .A1(n5510), .A2(n5511), .A3(n5513), .A4(n5515), .ZN(n23132) );
  INV_X2 U32432 ( .I(n21792), .ZN(n59418) );
  NAND2_X1 U32438 ( .A1(n26258), .A2(n59420), .ZN(n2354) );
  NOR2_X2 U32448 ( .A1(n54337), .A2(n59421), .ZN(n54411) );
  OR2_X1 U32449 ( .A1(n10954), .A2(n12410), .Z(n10936) );
  NAND3_X1 U32455 ( .A1(n64080), .A2(n41537), .A3(n429), .ZN(n41541) );
  AOI21_X1 U32466 ( .A1(n8830), .A2(n60129), .B(n8829), .ZN(n59424) );
  NAND2_X2 U32470 ( .A1(n50383), .A2(n47925), .ZN(n49726) );
  NAND2_X2 U32475 ( .A1(n59409), .A2(n20598), .ZN(n41060) );
  NAND2_X2 U32478 ( .A1(n5282), .A2(n23707), .ZN(n14265) );
  NAND2_X1 U32489 ( .A1(n15007), .A2(n15091), .ZN(n59426) );
  NOR2_X2 U32492 ( .A1(n16447), .A2(n43415), .ZN(n11910) );
  NOR2_X2 U32500 ( .A1(n56631), .A2(n56627), .ZN(n56205) );
  NOR2_X1 U32514 ( .A1(n2329), .A2(n54901), .ZN(n54911) );
  NAND2_X1 U32515 ( .A1(n2904), .A2(n7622), .ZN(n49534) );
  XOR2_X1 U32516 ( .A1(n672), .A2(n22883), .Z(n18330) );
  XOR2_X1 U32522 ( .A1(n61546), .A2(n8866), .Z(n59634) );
  XOR2_X1 U32524 ( .A1(n32744), .A2(n32543), .Z(n30535) );
  XOR2_X1 U32536 ( .A1(n18709), .A2(n45057), .Z(n59428) );
  OR2_X1 U32543 ( .A1(n45968), .A2(n3510), .Z(n45960) );
  OAI22_X1 U32545 ( .A1(n55640), .A2(n5552), .B1(n55642), .B2(n55641), .ZN(
        n55647) );
  NOR2_X1 U32552 ( .A1(n25990), .A2(n31162), .ZN(n59429) );
  NAND3_X2 U32565 ( .A1(n6824), .A2(n6823), .A3(n6822), .ZN(n21314) );
  INV_X2 U32572 ( .I(n17620), .ZN(n21860) );
  NAND2_X2 U32578 ( .A1(n624), .A2(n17621), .ZN(n17620) );
  NOR2_X2 U32579 ( .A1(n17998), .A2(n17997), .ZN(n37292) );
  AND2_X2 U32580 ( .A1(n61893), .A2(n60630), .Z(n18737) );
  OR2_X1 U32590 ( .A1(n50406), .A2(n49732), .Z(n25555) );
  XOR2_X1 U32602 ( .A1(n52407), .A2(n7941), .Z(n59435) );
  NAND3_X1 U32614 ( .A1(n59437), .A2(n8290), .A3(n43741), .ZN(n24997) );
  NAND3_X1 U32630 ( .A1(n49905), .A2(n48739), .A3(n19243), .ZN(n24305) );
  AOI21_X1 U32631 ( .A1(n4940), .A2(n56017), .B(n59590), .ZN(n56028) );
  NOR2_X1 U32650 ( .A1(n36747), .A2(n36740), .ZN(n36753) );
  NOR2_X1 U32655 ( .A1(n33955), .A2(n32867), .ZN(n2533) );
  NAND3_X2 U32667 ( .A1(n20274), .A2(n17023), .A3(n59446), .ZN(n25811) );
  OR2_X1 U32670 ( .A1(n6892), .A2(n6599), .Z(n59447) );
  NOR3_X2 U32685 ( .A1(n59452), .A2(n15576), .A3(n59451), .ZN(n17717) );
  AOI22_X2 U32694 ( .A1(n40248), .A2(n37200), .B1(n65206), .B2(n39164), .ZN(
        n59453) );
  NAND2_X1 U32709 ( .A1(n56567), .A2(n56389), .ZN(n51253) );
  NOR2_X2 U32710 ( .A1(n28011), .A2(n59454), .ZN(n16382) );
  NAND3_X2 U32716 ( .A1(n41188), .A2(n40626), .A3(n16102), .ZN(n40623) );
  NAND2_X2 U32743 ( .A1(n21281), .A2(n27594), .ZN(n27073) );
  INV_X2 U32744 ( .I(n59460), .ZN(n1213) );
  INV_X2 U32751 ( .I(n49510), .ZN(n1374) );
  XOR2_X1 U32758 ( .A1(n51687), .A2(n65142), .Z(n51478) );
  NOR2_X2 U32760 ( .A1(n59514), .A2(n3320), .ZN(n8147) );
  NAND2_X2 U32763 ( .A1(n1330), .A2(n6588), .ZN(n11113) );
  XOR2_X1 U32770 ( .A1(n50722), .A2(n59464), .Z(n59463) );
  XOR2_X1 U32775 ( .A1(n59565), .A2(n31619), .Z(n59667) );
  NAND3_X2 U32780 ( .A1(n13011), .A2(n13009), .A3(n13012), .ZN(n13008) );
  XOR2_X1 U32790 ( .A1(n14720), .A2(n44807), .Z(n59465) );
  NAND2_X2 U32792 ( .A1(n16808), .A2(n22596), .ZN(n29805) );
  OAI21_X1 U32803 ( .A1(n24974), .A2(n2349), .B(n24973), .ZN(n10200) );
  NAND2_X1 U32805 ( .A1(n2063), .A2(n60604), .ZN(n59467) );
  BUF_X2 U32806 ( .I(n13799), .Z(n59468) );
  XOR2_X1 U32829 ( .A1(n32348), .A2(n33883), .Z(n61641) );
  XOR2_X1 U32831 ( .A1(n59469), .A2(n7238), .Z(n8368) );
  OAI21_X1 U32843 ( .A1(n16419), .A2(n28504), .B(n59470), .ZN(n7809) );
  NOR2_X1 U32844 ( .A1(n27847), .A2(n27846), .ZN(n59470) );
  OAI22_X1 U32845 ( .A1(n33328), .A2(n36588), .B1(n33329), .B2(n18061), .ZN(
        n59473) );
  XOR2_X1 U32847 ( .A1(n59474), .A2(n61807), .Z(n60867) );
  XOR2_X1 U32848 ( .A1(n59993), .A2(n5048), .Z(n59474) );
  XOR2_X1 U32850 ( .A1(n17102), .A2(n59475), .Z(n44637) );
  XOR2_X1 U32851 ( .A1(n1057), .A2(n44636), .Z(n59475) );
  BUF_X2 U32853 ( .I(n43874), .Z(n59476) );
  NOR2_X2 U32857 ( .A1(n125), .A2(n59477), .ZN(n24471) );
  NOR2_X2 U32886 ( .A1(n29339), .A2(n29340), .ZN(n29341) );
  NAND2_X2 U32889 ( .A1(n23504), .A2(n27507), .ZN(n29339) );
  NAND3_X2 U32893 ( .A1(n5851), .A2(n43206), .A3(n10937), .ZN(n60519) );
  XOR2_X1 U32916 ( .A1(n7420), .A2(n59487), .Z(n10393) );
  XOR2_X1 U32921 ( .A1(n14059), .A2(n57230), .Z(n59487) );
  NAND3_X2 U32928 ( .A1(n47950), .A2(n47951), .A3(n47952), .ZN(n26007) );
  NAND2_X1 U32931 ( .A1(n29942), .A2(n30409), .ZN(n29948) );
  NAND2_X2 U32935 ( .A1(n33701), .A2(n33561), .ZN(n33342) );
  NAND2_X1 U32937 ( .A1(n25023), .A2(n59492), .ZN(n4027) );
  OAI21_X1 U32940 ( .A1(n57007), .A2(n20484), .B(n57006), .ZN(n59492) );
  XOR2_X1 U32970 ( .A1(n24891), .A2(n15591), .Z(n59495) );
  XOR2_X1 U32974 ( .A1(n24598), .A2(n4761), .Z(n20386) );
  XOR2_X1 U32975 ( .A1(n3424), .A2(n9698), .Z(n59496) );
  NAND3_X2 U32988 ( .A1(n8922), .A2(n8921), .A3(n41238), .ZN(n59497) );
  NAND2_X2 U32991 ( .A1(n49732), .A2(n50398), .ZN(n50074) );
  INV_X2 U32997 ( .I(n46719), .ZN(n50398) );
  NAND2_X2 U33005 ( .A1(n46467), .A2(n59499), .ZN(n46719) );
  AND2_X1 U33009 ( .A1(n46466), .A2(n47540), .Z(n59499) );
  NOR2_X2 U33010 ( .A1(n45601), .A2(n60250), .ZN(n45604) );
  XOR2_X1 U33013 ( .A1(n1676), .A2(n46293), .Z(n59501) );
  OR2_X2 U33025 ( .A1(n25668), .A2(n26214), .Z(n8304) );
  NOR2_X2 U33041 ( .A1(n54727), .A2(n22385), .ZN(n54669) );
  AND2_X1 U33052 ( .A1(n57731), .A2(n6081), .Z(n59505) );
  NOR3_X2 U33057 ( .A1(n15690), .A2(n59507), .A3(n59506), .ZN(n54670) );
  XOR2_X1 U33059 ( .A1(n17438), .A2(n1670), .Z(n7178) );
  XOR2_X1 U33060 ( .A1(n59508), .A2(n51699), .Z(n59931) );
  NAND3_X2 U33064 ( .A1(n37948), .A2(n37323), .A3(n10556), .ZN(n38573) );
  NAND2_X2 U33076 ( .A1(n59842), .A2(n1421), .ZN(n34484) );
  NAND2_X2 U33078 ( .A1(n12523), .A2(n1275), .ZN(n39118) );
  NAND2_X1 U33084 ( .A1(n47219), .A2(n21641), .ZN(n11391) );
  NAND3_X1 U33096 ( .A1(n54116), .A2(n54117), .A3(n54194), .ZN(n54125) );
  XOR2_X1 U33101 ( .A1(n59510), .A2(n38870), .Z(n37526) );
  XOR2_X1 U33102 ( .A1(n37524), .A2(n22953), .Z(n59510) );
  NOR2_X2 U33103 ( .A1(n22606), .A2(n11727), .ZN(n41788) );
  NAND3_X2 U33106 ( .A1(n22074), .A2(n22078), .A3(n22073), .ZN(n35490) );
  NAND2_X1 U33117 ( .A1(n47223), .A2(n47224), .ZN(n59514) );
  NOR2_X2 U33122 ( .A1(n60908), .A2(n59515), .ZN(n21780) );
  XOR2_X1 U33123 ( .A1(n13569), .A2(n13568), .Z(n15046) );
  INV_X2 U33142 ( .I(n56224), .ZN(n18119) );
  NAND3_X2 U33144 ( .A1(n56277), .A2(n25411), .A3(n25410), .ZN(n56224) );
  BUF_X2 U33154 ( .I(n15725), .Z(n59521) );
  AOI21_X1 U33175 ( .A1(n15484), .A2(n52120), .B(n55905), .ZN(n7268) );
  NAND2_X2 U33177 ( .A1(n8479), .A2(n10341), .ZN(n40948) );
  OAI21_X2 U33181 ( .A1(n35681), .A2(n33299), .B(n33599), .ZN(n33311) );
  NOR2_X2 U33187 ( .A1(n1540), .A2(n63888), .ZN(n35681) );
  NAND2_X2 U33208 ( .A1(n8121), .A2(n63034), .ZN(n56269) );
  INV_X2 U33261 ( .I(n59533), .ZN(n55092) );
  NAND2_X2 U33263 ( .A1(n15520), .A2(n5051), .ZN(n59533) );
  XOR2_X1 U33272 ( .A1(n6322), .A2(n32719), .Z(n10649) );
  XOR2_X1 U33279 ( .A1(n30828), .A2(n54734), .Z(n32719) );
  AND2_X1 U33284 ( .A1(n55088), .A2(n59538), .Z(n2675) );
  XOR2_X1 U33288 ( .A1(n38063), .A2(n59576), .Z(n8600) );
  OR2_X2 U33290 ( .A1(n17978), .A2(n31261), .Z(n25013) );
  NOR2_X2 U33295 ( .A1(n16138), .A2(n23972), .ZN(n17978) );
  NAND2_X2 U33296 ( .A1(n58294), .A2(n15687), .ZN(n4231) );
  NOR3_X2 U33322 ( .A1(n9460), .A2(n60872), .A3(n7171), .ZN(n9457) );
  OR2_X1 U33338 ( .A1(n61167), .A2(n33647), .Z(n9760) );
  XOR2_X1 U33341 ( .A1(n59542), .A2(n57237), .Z(n970) );
  XOR2_X1 U33342 ( .A1(n2317), .A2(n2870), .Z(n59542) );
  XOR2_X1 U33348 ( .A1(n32744), .A2(n59544), .Z(n32745) );
  XOR2_X1 U33349 ( .A1(n32743), .A2(n45011), .Z(n59544) );
  INV_X2 U33351 ( .I(n22867), .ZN(n59545) );
  INV_X4 U33352 ( .I(n9337), .ZN(n16982) );
  NOR2_X2 U33353 ( .A1(n48148), .A2(n46753), .ZN(n4660) );
  INV_X2 U33354 ( .I(n59550), .ZN(n20344) );
  XOR2_X1 U33355 ( .A1(n20345), .A2(n24592), .Z(n59550) );
  XOR2_X1 U33357 ( .A1(n25455), .A2(n14981), .Z(n15869) );
  NAND3_X2 U33358 ( .A1(n10858), .A2(n29836), .A3(n29837), .ZN(n14981) );
  INV_X2 U33359 ( .I(n59551), .ZN(n17845) );
  XOR2_X1 U33364 ( .A1(n44594), .A2(n44592), .Z(n15480) );
  NOR2_X2 U33366 ( .A1(n41967), .A2(n41968), .ZN(n44594) );
  NAND2_X2 U33386 ( .A1(n25427), .A2(n22477), .ZN(n33374) );
  BUF_X2 U33387 ( .I(n41186), .Z(n59554) );
  NAND2_X1 U33416 ( .A1(n17467), .A2(n59560), .ZN(n41732) );
  NOR2_X1 U33419 ( .A1(n42676), .A2(n42672), .ZN(n59560) );
  OR2_X2 U33426 ( .A1(n11329), .A2(n20786), .Z(n491) );
  XOR2_X1 U33432 ( .A1(n10116), .A2(n24201), .Z(n13283) );
  NAND2_X2 U33451 ( .A1(n1622), .A2(n22350), .ZN(n11882) );
  NOR2_X2 U33460 ( .A1(n47963), .A2(n47962), .ZN(n22350) );
  NOR2_X2 U33463 ( .A1(n23888), .A2(n59563), .ZN(n23887) );
  NAND3_X2 U33473 ( .A1(n25044), .A2(n25043), .A3(n27833), .ZN(n59563) );
  NAND2_X2 U33489 ( .A1(n14904), .A2(n37034), .ZN(n22267) );
  XOR2_X1 U33497 ( .A1(n32229), .A2(n57445), .Z(n59565) );
  INV_X2 U33498 ( .I(n59566), .ZN(n4784) );
  XOR2_X1 U33500 ( .A1(Ciphertext[84]), .A2(Key[1]), .Z(n59566) );
  NAND3_X2 U33502 ( .A1(n60127), .A2(n51113), .A3(n52721), .ZN(n61222) );
  OR2_X2 U33510 ( .A1(n58830), .A2(n7487), .Z(n47510) );
  NOR2_X2 U33520 ( .A1(n57204), .A2(n1640), .ZN(n7113) );
  NAND3_X2 U33523 ( .A1(n216), .A2(n215), .A3(n59567), .ZN(n29232) );
  AND3_X1 U33531 ( .A1(n26453), .A2(n27225), .A3(n26448), .Z(n59567) );
  AOI21_X1 U33538 ( .A1(n30811), .A2(n6720), .B(n8521), .ZN(n30813) );
  OAI22_X1 U33540 ( .A1(n2418), .A2(n34937), .B1(n1766), .B2(n36719), .ZN(
        n34938) );
  XOR2_X1 U33553 ( .A1(n14857), .A2(n6872), .Z(n59568) );
  AND2_X1 U33561 ( .A1(n46565), .A2(n20624), .Z(n61205) );
  OAI21_X1 U33565 ( .A1(n32784), .A2(n32458), .B(n33612), .ZN(n16887) );
  NAND2_X2 U33570 ( .A1(n20996), .A2(n3112), .ZN(n2499) );
  OR2_X1 U33573 ( .A1(n45968), .A2(n19329), .Z(n13879) );
  XOR2_X1 U33583 ( .A1(n44169), .A2(n46234), .Z(n44354) );
  NAND2_X2 U33584 ( .A1(n23065), .A2(n15786), .ZN(n60054) );
  NAND2_X2 U33585 ( .A1(n23449), .A2(n37224), .ZN(n59570) );
  NOR3_X2 U33593 ( .A1(n11669), .A2(n11671), .A3(n11670), .ZN(n11088) );
  XOR2_X1 U33596 ( .A1(n32036), .A2(n59571), .Z(n5148) );
  XOR2_X1 U33598 ( .A1(n4901), .A2(n57326), .Z(n59571) );
  XOR2_X1 U33605 ( .A1(n19357), .A2(n59572), .Z(n60204) );
  XNOR2_X1 U33625 ( .A1(n6250), .A2(n32029), .ZN(n4917) );
  OAI22_X1 U33632 ( .A1(n40667), .A2(n5775), .B1(n40656), .B2(n40491), .ZN(
        n40493) );
  NOR2_X2 U33652 ( .A1(n6177), .A2(n10766), .ZN(n16885) );
  NAND3_X2 U33669 ( .A1(n57217), .A2(n21776), .A3(n30221), .ZN(n2378) );
  XOR2_X1 U33670 ( .A1(n32084), .A2(n33838), .Z(n16522) );
  XOR2_X1 U33673 ( .A1(n19993), .A2(n1826), .Z(n32084) );
  XOR2_X1 U33708 ( .A1(n37118), .A2(n1248), .Z(n20367) );
  XOR2_X1 U33739 ( .A1(n25062), .A2(n18987), .Z(n59581) );
  INV_X2 U33745 ( .I(n50361), .ZN(n26208) );
  NOR3_X2 U33758 ( .A1(n21468), .A2(n1310), .A3(n22528), .ZN(n36197) );
  AND2_X2 U33761 ( .A1(n35152), .A2(n12887), .Z(n36106) );
  AOI22_X2 U33768 ( .A1(n59586), .A2(n49203), .B1(n7972), .B2(n49202), .ZN(
        n60538) );
  AND2_X1 U33801 ( .A1(n30823), .A2(n30824), .Z(n59589) );
  OR2_X2 U33805 ( .A1(n11340), .A2(n35685), .Z(n4496) );
  OAI22_X1 U33806 ( .A1(n56015), .A2(n56047), .B1(n56024), .B2(n56014), .ZN(
        n59590) );
  NAND3_X2 U33829 ( .A1(n59594), .A2(n30881), .A3(n30882), .ZN(n32669) );
  NOR2_X2 U33835 ( .A1(n4577), .A2(n35698), .ZN(n23908) );
  NAND2_X1 U33857 ( .A1(n48382), .A2(n21875), .ZN(n59962) );
  BUF_X2 U33858 ( .I(n9655), .Z(n59599) );
  NAND3_X1 U33868 ( .A1(n26585), .A2(n23446), .A3(n30392), .ZN(n5866) );
  INV_X2 U33872 ( .I(n25134), .ZN(n22794) );
  NAND3_X2 U33880 ( .A1(n9128), .A2(n9129), .A3(n9134), .ZN(n59602) );
  NAND2_X2 U33883 ( .A1(n33445), .A2(n23014), .ZN(n35045) );
  INV_X2 U33885 ( .I(n54063), .ZN(n54318) );
  NAND2_X2 U33895 ( .A1(n14323), .A2(n25841), .ZN(n47696) );
  AND2_X1 U33897 ( .A1(n13126), .A2(n9806), .Z(n35937) );
  OAI21_X2 U33903 ( .A1(n13057), .A2(n13059), .B(n26156), .ZN(n56666) );
  NOR2_X2 U33914 ( .A1(n59603), .A2(n24457), .ZN(n37184) );
  AOI21_X2 U33917 ( .A1(n34335), .A2(n34263), .B(n20989), .ZN(n34264) );
  INV_X4 U33919 ( .I(n21470), .ZN(n59610) );
  NOR3_X1 U33924 ( .A1(n28648), .A2(n28640), .A3(n491), .ZN(n28185) );
  INV_X2 U33945 ( .I(n20786), .ZN(n59604) );
  AOI22_X1 U33955 ( .A1(n47475), .A2(n47476), .B1(n47473), .B2(n47474), .ZN(
        n47477) );
  NAND2_X2 U33958 ( .A1(n34268), .A2(n15041), .ZN(n23354) );
  NAND2_X2 U33967 ( .A1(n63582), .A2(n59607), .ZN(n36065) );
  INV_X2 U33976 ( .I(n19206), .ZN(n59608) );
  NAND2_X2 U33977 ( .A1(n63105), .A2(n5090), .ZN(n47080) );
  XOR2_X1 U33978 ( .A1(n3843), .A2(n32556), .Z(n15640) );
  XOR2_X1 U33985 ( .A1(n13742), .A2(n32186), .Z(n3843) );
  OAI21_X1 U33991 ( .A1(n36394), .A2(n36538), .B(n36053), .ZN(n60874) );
  NOR2_X2 U33995 ( .A1(n18459), .A2(n50229), .ZN(n59621) );
  OR2_X2 U34002 ( .A1(n20337), .A2(n36717), .Z(n36725) );
  NOR2_X2 U34006 ( .A1(n44), .A2(n35641), .ZN(n36986) );
  OR2_X1 U34007 ( .A1(n3246), .A2(n60567), .Z(n38691) );
  OAI22_X1 U34011 ( .A1(n17964), .A2(n22523), .B1(n41027), .B2(n38498), .ZN(
        n13311) );
  INV_X2 U34013 ( .I(n12384), .ZN(n41027) );
  NAND2_X2 U34017 ( .A1(n21057), .A2(n41034), .ZN(n12384) );
  XOR2_X1 U34030 ( .A1(n7935), .A2(n61857), .Z(n741) );
  BUF_X2 U34032 ( .I(n29915), .Z(n59613) );
  XOR2_X1 U34036 ( .A1(n59615), .A2(n40785), .Z(n44369) );
  XOR2_X1 U34037 ( .A1(n24055), .A2(n43941), .Z(n59615) );
  NAND2_X2 U34044 ( .A1(n41875), .A2(n14624), .ZN(n11895) );
  NOR2_X1 U34054 ( .A1(n5742), .A2(n30637), .ZN(n5741) );
  XOR2_X1 U34069 ( .A1(n44511), .A2(n60650), .Z(n44375) );
  NAND3_X2 U34087 ( .A1(n61411), .A2(n52982), .A3(n486), .ZN(n53816) );
  XOR2_X1 U34096 ( .A1(n59866), .A2(n43966), .Z(n59620) );
  BUF_X2 U34109 ( .I(n19654), .Z(n59622) );
  XOR2_X1 U34115 ( .A1(n32261), .A2(n32260), .Z(n32262) );
  NAND2_X2 U34156 ( .A1(n2247), .A2(n41900), .ZN(n42258) );
  OAI22_X1 U34194 ( .A1(n53351), .A2(n13667), .B1(n1450), .B2(n63931), .ZN(
        n53363) );
  XOR2_X1 U34212 ( .A1(n46347), .A2(n46346), .Z(n10628) );
  OR2_X2 U34224 ( .A1(n24873), .A2(n6698), .Z(n46959) );
  OAI21_X1 U34227 ( .A1(n4133), .A2(n4134), .B(n40569), .ZN(n4132) );
  NOR2_X2 U34242 ( .A1(n11666), .A2(n11667), .ZN(n16891) );
  NOR2_X2 U34244 ( .A1(n35755), .A2(n35318), .ZN(n31955) );
  NOR2_X1 U34249 ( .A1(n2100), .A2(n29998), .ZN(n60248) );
  OAI21_X2 U34252 ( .A1(n49731), .A2(n59200), .B(n50082), .ZN(n15170) );
  INV_X2 U34260 ( .I(n49433), .ZN(n59640) );
  XOR2_X1 U34263 ( .A1(n50385), .A2(n12986), .Z(n50184) );
  XOR2_X1 U34264 ( .A1(n49189), .A2(n12985), .Z(n50385) );
  NOR2_X2 U34267 ( .A1(n59642), .A2(n11728), .ZN(n14397) );
  NOR2_X2 U34281 ( .A1(n23328), .A2(n27171), .ZN(n21281) );
  XOR2_X1 U34286 ( .A1(n31499), .A2(n57440), .Z(n10911) );
  XOR2_X1 U34287 ( .A1(n31490), .A2(n807), .Z(n31499) );
  NAND2_X1 U34288 ( .A1(n47932), .A2(n5282), .ZN(n47933) );
  NAND2_X2 U34306 ( .A1(n20242), .A2(n22989), .ZN(n20243) );
  NAND3_X2 U34309 ( .A1(n50384), .A2(n59644), .A3(n9487), .ZN(n19349) );
  NAND2_X1 U34310 ( .A1(n50379), .A2(n50380), .ZN(n59644) );
  NOR2_X1 U34312 ( .A1(n17211), .A2(n51268), .ZN(n59646) );
  XOR2_X1 U34319 ( .A1(n38661), .A2(n20355), .Z(n13190) );
  XOR2_X1 U34325 ( .A1(n37709), .A2(n4691), .Z(n38661) );
  INV_X1 U34326 ( .I(n52846), .ZN(n59649) );
  NAND2_X2 U34327 ( .A1(n2018), .A2(n25067), .ZN(n52846) );
  BUF_X2 U34329 ( .I(n39935), .Z(n59650) );
  NOR2_X2 U34341 ( .A1(n3847), .A2(n14185), .ZN(n14370) );
  OR2_X1 U34351 ( .A1(n20845), .A2(n20846), .Z(n59660) );
  XOR2_X1 U34352 ( .A1(n3214), .A2(n59789), .Z(n4055) );
  XOR2_X1 U34355 ( .A1(n44892), .A2(n44891), .Z(n13959) );
  NAND2_X2 U34362 ( .A1(n4634), .A2(n56249), .ZN(n56587) );
  OAI22_X1 U34364 ( .A1(n56292), .A2(n56291), .B1(n56311), .B2(n24585), .ZN(
        n24584) );
  NAND2_X1 U34367 ( .A1(n56342), .A2(n1591), .ZN(n56291) );
  INV_X4 U34381 ( .I(n24332), .ZN(n617) );
  XOR2_X1 U34382 ( .A1(n59663), .A2(n33127), .Z(n33334) );
  NAND3_X1 U34383 ( .A1(n8129), .A2(n1639), .A3(n49317), .ZN(n47445) );
  NAND3_X2 U34394 ( .A1(n17194), .A2(n5383), .A3(n17196), .ZN(n39222) );
  AND2_X2 U34398 ( .A1(n8337), .A2(n6728), .Z(n637) );
  INV_X2 U34405 ( .I(n59667), .ZN(n9289) );
  CLKBUF_X8 U34406 ( .I(n21240), .Z(n61134) );
  OAI21_X1 U34407 ( .A1(n38198), .A2(n38199), .B(n1401), .ZN(n38201) );
  NAND2_X2 U34416 ( .A1(n1530), .A2(n12652), .ZN(n36627) );
  OAI22_X1 U34420 ( .A1(n35848), .A2(n2168), .B1(n35847), .B2(n21252), .ZN(
        n35849) );
  NOR2_X2 U34425 ( .A1(n35834), .A2(n25188), .ZN(n34392) );
  XOR2_X1 U34426 ( .A1(n59668), .A2(n62380), .Z(n38287) );
  XOR2_X1 U34430 ( .A1(n5555), .A2(n9956), .Z(n59668) );
  NAND3_X2 U34433 ( .A1(n29732), .A2(n29731), .A3(n61753), .ZN(n19852) );
  XOR2_X1 U34434 ( .A1(n38140), .A2(n59669), .Z(n9810) );
  XOR2_X1 U34441 ( .A1(n38139), .A2(n3625), .Z(n59669) );
  NAND2_X1 U34442 ( .A1(n48966), .A2(n59975), .ZN(n59974) );
  NOR2_X1 U34444 ( .A1(n59974), .A2(n48964), .ZN(n2645) );
  OAI21_X1 U34453 ( .A1(n12515), .A2(n33774), .B(n33766), .ZN(n12514) );
  NOR3_X2 U34465 ( .A1(n24851), .A2(n29505), .A3(n59671), .ZN(n7211) );
  XOR2_X1 U34472 ( .A1(n59673), .A2(n53328), .Z(Plaintext[20]) );
  INV_X1 U34474 ( .I(n36850), .ZN(n35494) );
  AOI22_X1 U34475 ( .A1(n6807), .A2(n19553), .B1(n36850), .B2(n60824), .ZN(
        n19607) );
  XOR2_X1 U34484 ( .A1(n33879), .A2(n32289), .Z(n14049) );
  NAND3_X2 U34487 ( .A1(n28976), .A2(n28975), .A3(n28974), .ZN(n33879) );
  NAND2_X1 U34495 ( .A1(n47954), .A2(n50285), .ZN(n47959) );
  XOR2_X1 U34498 ( .A1(n59675), .A2(n5595), .Z(n8540) );
  XOR2_X1 U34502 ( .A1(n3397), .A2(n3395), .Z(n59675) );
  NAND2_X1 U34503 ( .A1(n56191), .A2(n5172), .ZN(n56184) );
  XOR2_X1 U34521 ( .A1(n57836), .A2(n10898), .Z(n3396) );
  NAND3_X1 U34524 ( .A1(n53999), .A2(n6135), .A3(n7492), .ZN(n54003) );
  XOR2_X1 U34532 ( .A1(n32193), .A2(n32194), .Z(n59678) );
  NAND4_X2 U34537 ( .A1(n53893), .A2(n53891), .A3(n54592), .A4(n53892), .ZN(
        n53900) );
  NOR2_X1 U34539 ( .A1(n30680), .A2(n26740), .ZN(n14393) );
  NAND2_X2 U34548 ( .A1(n13489), .A2(n22029), .ZN(n8784) );
  NOR2_X2 U34554 ( .A1(n26912), .A2(n29690), .ZN(n20581) );
  AND2_X1 U34569 ( .A1(n41173), .A2(n41186), .Z(n39144) );
  NAND2_X2 U34571 ( .A1(n39147), .A2(n40666), .ZN(n41173) );
  NAND2_X2 U34576 ( .A1(n3761), .A2(n22745), .ZN(n31209) );
  XOR2_X1 U34591 ( .A1(n19066), .A2(n59689), .Z(n19065) );
  XOR2_X1 U34595 ( .A1(n19760), .A2(n22451), .Z(n59689) );
  XOR2_X1 U34599 ( .A1(Ciphertext[128]), .A2(Key[117]), .Z(n9995) );
  NOR3_X2 U34609 ( .A1(n21555), .A2(n21552), .A3(n59691), .ZN(n21551) );
  OAI22_X1 U34620 ( .A1(n46059), .A2(n45957), .B1(n46060), .B2(n47324), .ZN(
        n59691) );
  XOR2_X1 U34623 ( .A1(n8353), .A2(n19545), .Z(n59751) );
  INV_X2 U34625 ( .I(n43358), .ZN(n1685) );
  NAND2_X2 U34631 ( .A1(n6426), .A2(n21644), .ZN(n43358) );
  OAI21_X1 U34635 ( .A1(n40493), .A2(n40492), .B(n41172), .ZN(n59692) );
  NAND3_X1 U34651 ( .A1(n42239), .A2(n7728), .A3(n25247), .ZN(n41915) );
  NOR2_X1 U34652 ( .A1(n2066), .A2(n58601), .ZN(n28198) );
  NOR2_X2 U34671 ( .A1(n15595), .A2(n47873), .ZN(n7358) );
  XOR2_X1 U34675 ( .A1(n50736), .A2(n50844), .Z(n12704) );
  XOR2_X1 U34680 ( .A1(n63263), .A2(n24880), .Z(n50844) );
  NAND2_X2 U34694 ( .A1(n47266), .A2(n25004), .ZN(n46882) );
  NAND2_X1 U34704 ( .A1(n1233), .A2(n55015), .ZN(n55038) );
  XOR2_X1 U34715 ( .A1(n13662), .A2(n59705), .Z(n7608) );
  XOR2_X1 U34716 ( .A1(n8974), .A2(n59706), .Z(n59705) );
  XOR2_X1 U34733 ( .A1(n59708), .A2(n5924), .Z(n5923) );
  XOR2_X1 U34736 ( .A1(n22053), .A2(n10141), .Z(n59708) );
  NAND2_X2 U34745 ( .A1(n7836), .A2(n56599), .ZN(n7835) );
  NAND2_X1 U34753 ( .A1(n1), .A2(n2), .ZN(n10658) );
  XOR2_X1 U34759 ( .A1(n15308), .A2(n39231), .Z(n39261) );
  XOR2_X1 U34774 ( .A1(n22142), .A2(n2218), .Z(n46149) );
  AND3_X1 U34787 ( .A1(n12467), .A2(n16118), .A3(n6467), .Z(n12464) );
  BUF_X2 U34809 ( .I(n29586), .Z(n59710) );
  NOR3_X1 U34812 ( .A1(n43690), .A2(n43694), .A3(n41495), .ZN(n37916) );
  XOR2_X1 U34817 ( .A1(n32471), .A2(n19886), .Z(n33870) );
  XOR2_X1 U34822 ( .A1(n5973), .A2(n17078), .Z(n20355) );
  OAI21_X1 U34843 ( .A1(n54548), .A2(n54549), .B(n54547), .ZN(n54550) );
  NOR2_X2 U34850 ( .A1(n6244), .A2(n21334), .ZN(n48053) );
  NAND2_X2 U34855 ( .A1(n41970), .A2(n42693), .ZN(n9672) );
  OR2_X1 U34874 ( .A1(n39415), .A2(n36648), .Z(n40233) );
  NAND3_X2 U34889 ( .A1(n59715), .A2(n26103), .A3(n59714), .ZN(n50797) );
  XOR2_X1 U34890 ( .A1(n59716), .A2(n54676), .Z(Plaintext[78]) );
  NAND2_X1 U34894 ( .A1(n59719), .A2(n50364), .ZN(n59718) );
  NAND2_X1 U34906 ( .A1(n16711), .A2(n18598), .ZN(n59719) );
  XOR2_X1 U34922 ( .A1(n11147), .A2(n925), .Z(n59721) );
  NAND2_X2 U34925 ( .A1(n59722), .A2(n56237), .ZN(n14578) );
  XOR2_X1 U34938 ( .A1(n59723), .A2(n56950), .Z(Plaintext[184]) );
  NOR2_X1 U34943 ( .A1(n56947), .A2(n56948), .ZN(n59723) );
  NAND2_X1 U34948 ( .A1(n37236), .A2(n62992), .ZN(n37238) );
  NAND2_X2 U34974 ( .A1(n4780), .A2(n48711), .ZN(n49684) );
  NOR2_X2 U34999 ( .A1(n52861), .A2(n50601), .ZN(n57061) );
  NOR2_X1 U35003 ( .A1(n3175), .A2(n1808), .ZN(n3174) );
  INV_X2 U35027 ( .I(n40056), .ZN(n40274) );
  NAND2_X2 U35038 ( .A1(n1410), .A2(n8427), .ZN(n40056) );
  NAND2_X2 U35051 ( .A1(n10627), .A2(n18951), .ZN(n45618) );
  NOR2_X2 U35052 ( .A1(n5299), .A2(n45075), .ZN(n18951) );
  XOR2_X1 U35056 ( .A1(n51191), .A2(n59732), .Z(n7844) );
  XOR2_X1 U35064 ( .A1(n2153), .A2(n2603), .Z(n59732) );
  XOR2_X1 U35070 ( .A1(n39716), .A2(n38203), .Z(n39630) );
  NAND2_X2 U35075 ( .A1(n9782), .A2(n59734), .ZN(n31376) );
  NAND2_X2 U35081 ( .A1(n58811), .A2(n19085), .ZN(n53803) );
  NAND3_X1 U35109 ( .A1(n2047), .A2(n45792), .A3(n48071), .ZN(n17673) );
  INV_X1 U35122 ( .I(n4430), .ZN(n60276) );
  AND2_X1 U35128 ( .A1(n41870), .A2(n64986), .Z(n41867) );
  NAND2_X1 U35154 ( .A1(n51636), .A2(n51635), .ZN(n59741) );
  NAND2_X1 U35197 ( .A1(n15293), .A2(n17270), .ZN(n4485) );
  NOR2_X2 U35205 ( .A1(n48586), .A2(n24185), .ZN(n46176) );
  NOR3_X1 U35211 ( .A1(n55331), .A2(n61765), .A3(n59744), .ZN(n55334) );
  NAND2_X1 U35218 ( .A1(n55329), .A2(n55338), .ZN(n59744) );
  NAND2_X1 U35226 ( .A1(n46481), .A2(n19200), .ZN(n12766) );
  BUF_X2 U35242 ( .I(n1704), .Z(n59746) );
  XOR2_X1 U35258 ( .A1(n38285), .A2(n38284), .Z(n61009) );
  AOI22_X1 U35265 ( .A1(n13877), .A2(n40056), .B1(n40058), .B2(n40057), .ZN(
        n13875) );
  XOR2_X1 U35274 ( .A1(n59747), .A2(n79), .Z(n7313) );
  XOR2_X1 U35286 ( .A1(n16502), .A2(n7708), .Z(n59747) );
  XOR2_X1 U35293 ( .A1(n23481), .A2(n39481), .Z(n24213) );
  NAND3_X1 U35294 ( .A1(n43022), .A2(n42788), .A3(n42782), .ZN(n41662) );
  XOR2_X1 U35340 ( .A1(n44021), .A2(n9221), .Z(n59749) );
  NOR2_X2 U35350 ( .A1(n34349), .A2(n59750), .ZN(n21194) );
  NAND3_X2 U35354 ( .A1(n16819), .A2(n34731), .A3(n34730), .ZN(n59750) );
  AND3_X1 U35404 ( .A1(n35652), .A2(n6829), .A3(n22909), .Z(n61649) );
  XOR2_X1 U35425 ( .A1(n23915), .A2(n32414), .Z(n59776) );
  XOR2_X1 U35427 ( .A1(n32669), .A2(n53246), .Z(n32414) );
  XOR2_X1 U35440 ( .A1(n42819), .A2(n42909), .Z(n59758) );
  XOR2_X1 U35475 ( .A1(n4669), .A2(n59759), .Z(n8178) );
  XOR2_X1 U35476 ( .A1(n32421), .A2(n10535), .Z(n59759) );
  NAND3_X2 U35492 ( .A1(n17004), .A2(n48044), .A3(n48045), .ZN(n22741) );
  XOR2_X1 U35524 ( .A1(n37735), .A2(n37734), .Z(n12392) );
  XOR2_X1 U35525 ( .A1(n23280), .A2(n233), .Z(n37735) );
  NOR3_X1 U35527 ( .A1(n54006), .A2(n53927), .A3(n53926), .ZN(n53928) );
  NOR2_X2 U35546 ( .A1(n60768), .A2(n27040), .ZN(n27036) );
  XOR2_X1 U35568 ( .A1(n59763), .A2(n5913), .Z(n3889) );
  NOR2_X2 U35575 ( .A1(n23479), .A2(n29371), .ZN(n28813) );
  XOR2_X1 U35586 ( .A1(n31772), .A2(n881), .Z(n59765) );
  NOR2_X2 U35602 ( .A1(n13837), .A2(n55656), .ZN(n14324) );
  NAND2_X1 U35605 ( .A1(n50351), .A2(n60378), .ZN(n21352) );
  NAND3_X2 U35612 ( .A1(n48000), .A2(n47999), .A3(n48001), .ZN(n7847) );
  NAND2_X1 U35618 ( .A1(n61846), .A2(n49340), .ZN(n47223) );
  INV_X2 U35650 ( .I(n48656), .ZN(n17153) );
  NAND2_X2 U35656 ( .A1(n6957), .A2(n22283), .ZN(n48656) );
  NAND2_X2 U35669 ( .A1(n6977), .A2(n20894), .ZN(n2608) );
  NOR2_X2 U35694 ( .A1(n59772), .A2(n42015), .ZN(n6110) );
  NAND2_X2 U35700 ( .A1(n7400), .A2(n7401), .ZN(n59772) );
  NAND2_X2 U35714 ( .A1(n20060), .A2(n36775), .ZN(n36773) );
  NOR2_X1 U35725 ( .A1(n2593), .A2(n24366), .ZN(n14342) );
  NAND2_X2 U35726 ( .A1(n6102), .A2(n26131), .ZN(n6101) );
  XOR2_X1 U35740 ( .A1(n31481), .A2(n60555), .Z(n19) );
  OR2_X1 U35786 ( .A1(n30871), .A2(n6317), .Z(n30873) );
  XOR2_X1 U35848 ( .A1(n14087), .A2(n59781), .Z(n13689) );
  XOR2_X1 U35861 ( .A1(n44768), .A2(n57359), .Z(n59781) );
  XOR2_X1 U35890 ( .A1(n59782), .A2(n60514), .Z(n32255) );
  XOR2_X1 U35892 ( .A1(n32253), .A2(n15464), .Z(n59782) );
  OAI22_X1 U35895 ( .A1(n48801), .A2(n7485), .B1(n49710), .B2(n1469), .ZN(
        n2072) );
  NAND2_X2 U35910 ( .A1(n17860), .A2(n59783), .ZN(n56238) );
  AOI22_X1 U35921 ( .A1(n1596), .A2(n12468), .B1(n56362), .B2(n17860), .ZN(
        n56363) );
  NOR3_X2 U35926 ( .A1(n59785), .A2(n40466), .A3(n40941), .ZN(n163) );
  NOR2_X1 U35939 ( .A1(n40463), .A2(n40468), .ZN(n59785) );
  XOR2_X1 U35941 ( .A1(n46587), .A2(n46282), .Z(n7410) );
  NAND3_X2 U35955 ( .A1(n11880), .A2(n41786), .A3(n41785), .ZN(n46587) );
  AOI22_X1 U35990 ( .A1(n54413), .A2(n54423), .B1(n54412), .B2(n54414), .ZN(
        n54429) );
  XOR2_X1 U35992 ( .A1(n2367), .A2(n18920), .Z(n2911) );
  INV_X2 U35994 ( .I(n28135), .ZN(n28128) );
  NOR2_X2 U36015 ( .A1(n62263), .A2(n56430), .ZN(n55985) );
  NOR2_X1 U36023 ( .A1(n21357), .A2(n30303), .ZN(n30304) );
  NAND2_X2 U36031 ( .A1(n9865), .A2(n29575), .ZN(n30302) );
  NAND2_X2 U36037 ( .A1(n12741), .A2(n29609), .ZN(n28676) );
  NAND2_X2 U36053 ( .A1(n12635), .A2(n18881), .ZN(n30743) );
  NAND2_X2 U36093 ( .A1(n56451), .A2(n56452), .ZN(n15237) );
  XOR2_X1 U36128 ( .A1(n51127), .A2(n51186), .Z(n59789) );
  NAND3_X2 U36146 ( .A1(n11348), .A2(n11350), .A3(n34472), .ZN(n23294) );
  XOR2_X1 U36153 ( .A1(n31985), .A2(n24098), .Z(n31748) );
  XOR2_X1 U36179 ( .A1(n59794), .A2(n24355), .Z(Plaintext[39]) );
  NAND4_X2 U36184 ( .A1(n50826), .A2(n50823), .A3(n50824), .A4(n50825), .ZN(
        n59794) );
  NOR2_X2 U36202 ( .A1(n7448), .A2(n59795), .ZN(n5679) );
  XOR2_X1 U36231 ( .A1(n146), .A2(n59797), .Z(n10098) );
  INV_X1 U36233 ( .I(n19511), .ZN(n59797) );
  NAND2_X1 U36236 ( .A1(n17286), .A2(n25117), .ZN(n50818) );
  BUF_X4 U36253 ( .I(n49940), .Z(n61624) );
  XOR2_X1 U36267 ( .A1(n12716), .A2(n59799), .Z(n51699) );
  XOR2_X1 U36274 ( .A1(n14730), .A2(n51697), .Z(n59799) );
  NAND2_X1 U36286 ( .A1(n45010), .A2(n14417), .ZN(n59801) );
  XOR2_X1 U36289 ( .A1(n25432), .A2(n19926), .Z(n61347) );
  NAND2_X2 U36291 ( .A1(n24869), .A2(n24868), .ZN(n60525) );
  XOR2_X1 U36304 ( .A1(n13486), .A2(n2616), .Z(n2615) );
  XOR2_X1 U36354 ( .A1(n17869), .A2(n6571), .Z(n59804) );
  NAND2_X2 U36359 ( .A1(n26280), .A2(n28048), .ZN(n24836) );
  INV_X2 U36368 ( .I(n59805), .ZN(n7760) );
  XOR2_X1 U36376 ( .A1(Ciphertext[103]), .A2(Key[38]), .Z(n59805) );
  OR2_X2 U36396 ( .A1(n20953), .A2(n20739), .Z(n34634) );
  XOR2_X1 U36423 ( .A1(n9820), .A2(n60736), .Z(n21276) );
  AND2_X1 U36436 ( .A1(n25233), .A2(n50283), .Z(n49882) );
  AOI22_X1 U36449 ( .A1(n53929), .A2(n53930), .B1(n53928), .B2(n53946), .ZN(
        n53943) );
  NAND3_X2 U36450 ( .A1(n1861), .A2(n20606), .A3(n23918), .ZN(n29485) );
  NAND3_X2 U36457 ( .A1(n331), .A2(n18575), .A3(n12143), .ZN(n45115) );
  INV_X1 U36458 ( .I(n47611), .ZN(n59813) );
  NAND2_X1 U36509 ( .A1(n60046), .A2(n52992), .ZN(n52995) );
  NAND3_X2 U36540 ( .A1(n59817), .A2(n40717), .A3(n40718), .ZN(n42639) );
  XOR2_X1 U36546 ( .A1(n298), .A2(n38587), .Z(n18899) );
  XOR2_X1 U36553 ( .A1(n23674), .A2(n51651), .Z(n11255) );
  NAND2_X1 U36566 ( .A1(n30870), .A2(n31264), .ZN(n20069) );
  NOR2_X2 U36580 ( .A1(n4257), .A2(n6316), .ZN(n30870) );
  NAND2_X1 U36602 ( .A1(n59822), .A2(n59821), .ZN(n59820) );
  NAND2_X1 U36604 ( .A1(n45770), .A2(n23480), .ZN(n59822) );
  NOR2_X2 U36620 ( .A1(n59823), .A2(n2653), .ZN(n24869) );
  NOR2_X1 U36627 ( .A1(n42758), .A2(n42759), .ZN(n42762) );
  BUF_X2 U36637 ( .I(n57342), .Z(n59824) );
  INV_X4 U36649 ( .I(n24357), .ZN(n36926) );
  INV_X2 U36652 ( .I(n54316), .ZN(n20965) );
  OAI21_X1 U36657 ( .A1(n17768), .A2(n40605), .B(n16462), .ZN(n61597) );
  OAI22_X1 U36698 ( .A1(n26579), .A2(n26578), .B1(n28232), .B2(n21301), .ZN(
        n26582) );
  NAND2_X2 U36706 ( .A1(n21301), .A2(n26577), .ZN(n26579) );
  XOR2_X1 U36711 ( .A1(n59018), .A2(n38999), .Z(n59826) );
  XOR2_X1 U36731 ( .A1(n25804), .A2(n51211), .Z(n18186) );
  XOR2_X1 U36736 ( .A1(n50796), .A2(n61423), .Z(n51211) );
  XOR2_X1 U36753 ( .A1(n4876), .A2(n45346), .Z(n14748) );
  NAND2_X2 U36758 ( .A1(n47252), .A2(n63793), .ZN(n45674) );
  BUF_X2 U36762 ( .I(n56829), .Z(n59827) );
  XOR2_X1 U36773 ( .A1(n13441), .A2(n2777), .Z(n21452) );
  AOI21_X2 U36805 ( .A1(n14893), .A2(n8819), .B(n14892), .ZN(n14894) );
  INV_X2 U36812 ( .I(n15282), .ZN(n49540) );
  NAND2_X2 U36814 ( .A1(n49377), .A2(n49374), .ZN(n15282) );
  OAI21_X1 U36819 ( .A1(n8760), .A2(n36113), .B(n36115), .ZN(n8759) );
  XOR2_X1 U36823 ( .A1(n12428), .A2(n21923), .Z(n59829) );
  NAND2_X2 U36832 ( .A1(n48757), .A2(n50426), .ZN(n23992) );
  INV_X1 U36834 ( .I(n6438), .ZN(n39477) );
  NOR2_X2 U36835 ( .A1(n58808), .A2(n55223), .ZN(n18786) );
  OAI21_X1 U36853 ( .A1(n60501), .A2(n41004), .B(n41003), .ZN(n41012) );
  AND2_X1 U36859 ( .A1(n7809), .A2(n7808), .Z(n60807) );
  XOR2_X1 U36868 ( .A1(n12942), .A2(n51987), .Z(n59832) );
  NAND2_X2 U36913 ( .A1(n19868), .A2(n34268), .ZN(n21751) );
  XOR2_X1 U36919 ( .A1(n10635), .A2(n20742), .Z(n49210) );
  NAND2_X1 U36927 ( .A1(n59836), .A2(n59834), .ZN(n10137) );
  NOR2_X1 U36936 ( .A1(n59835), .A2(n22063), .ZN(n59834) );
  NAND2_X1 U36966 ( .A1(n34051), .A2(n21906), .ZN(n59835) );
  INV_X1 U36971 ( .I(n24084), .ZN(n59836) );
  NAND2_X1 U36996 ( .A1(n17333), .A2(n29373), .ZN(n27444) );
  NOR2_X1 U37014 ( .A1(n32784), .A2(n32457), .ZN(n60189) );
  NOR2_X2 U37021 ( .A1(n60426), .A2(n54001), .ZN(n53947) );
  NAND2_X2 U37032 ( .A1(n1782), .A2(n10829), .ZN(n19064) );
  XOR2_X1 U37056 ( .A1(n15447), .A2(n59843), .Z(n10090) );
  XOR2_X1 U37062 ( .A1(n52073), .A2(n52072), .Z(n59843) );
  INV_X2 U37067 ( .I(n59844), .ZN(n5115) );
  XOR2_X1 U37068 ( .A1(n18783), .A2(n18784), .Z(n59844) );
  XOR2_X1 U37076 ( .A1(n17944), .A2(n17943), .Z(n17942) );
  AND2_X2 U37081 ( .A1(n39502), .A2(n8576), .Z(n40570) );
  NAND3_X2 U37132 ( .A1(n59848), .A2(n19150), .A3(n47692), .ZN(n18976) );
  XOR2_X1 U37136 ( .A1(n45813), .A2(n45271), .Z(n59849) );
  NOR3_X2 U37171 ( .A1(n39897), .A2(n39898), .A3(n39896), .ZN(n39935) );
  INV_X1 U37186 ( .I(n5522), .ZN(n15701) );
  XOR2_X1 U37200 ( .A1(n37987), .A2(n39230), .Z(n5522) );
  NOR2_X2 U37201 ( .A1(n31041), .A2(n21176), .ZN(n30701) );
  NOR2_X2 U37209 ( .A1(n57873), .A2(n5261), .ZN(n42329) );
  NAND2_X2 U37228 ( .A1(n26853), .A2(n27345), .ZN(n19700) );
  NOR2_X2 U37235 ( .A1(n12325), .A2(n59862), .ZN(n49054) );
  NAND3_X2 U37247 ( .A1(n59949), .A2(n45739), .A3(n6507), .ZN(n59862) );
  XOR2_X1 U37253 ( .A1(n59863), .A2(n964), .Z(n2665) );
  NAND2_X2 U37275 ( .A1(n19598), .A2(n30145), .ZN(n31041) );
  XOR2_X1 U37276 ( .A1(n13060), .A2(n12436), .Z(n39383) );
  XOR2_X1 U37299 ( .A1(n4052), .A2(n39223), .Z(n12436) );
  OAI21_X2 U37350 ( .A1(n8484), .A2(n8485), .B(n8483), .ZN(n59867) );
  XOR2_X1 U37352 ( .A1(n59868), .A2(n14096), .Z(n52608) );
  AOI22_X1 U37365 ( .A1(n14212), .A2(n26863), .B1(n29702), .B2(n27813), .ZN(
        n26869) );
  NAND3_X2 U37381 ( .A1(n60461), .A2(n18533), .A3(n18532), .ZN(n18531) );
  XOR2_X1 U37383 ( .A1(n9477), .A2(n1573), .Z(n45057) );
  XOR2_X1 U37406 ( .A1(n33876), .A2(n59875), .Z(n12240) );
  XOR2_X1 U37410 ( .A1(n33874), .A2(n708), .Z(n59875) );
  XOR2_X1 U37415 ( .A1(n63016), .A2(n59876), .Z(n13211) );
  XOR2_X1 U37432 ( .A1(n16700), .A2(n4800), .Z(n59876) );
  XOR2_X1 U37435 ( .A1(n13975), .A2(n6133), .Z(n8983) );
  NOR2_X2 U37436 ( .A1(n23782), .A2(n35271), .ZN(n13975) );
  NOR2_X1 U37441 ( .A1(n435), .A2(n17904), .ZN(n2276) );
  XOR2_X1 U37448 ( .A1(n59877), .A2(n60713), .Z(n7306) );
  NOR2_X2 U37452 ( .A1(n17291), .A2(n59878), .ZN(n28717) );
  NAND2_X2 U37453 ( .A1(n2066), .A2(n2067), .ZN(n29662) );
  XOR2_X1 U37467 ( .A1(n59880), .A2(n54708), .Z(Plaintext[79]) );
  XOR2_X1 U37487 ( .A1(n59881), .A2(n52612), .Z(n14459) );
  XOR2_X1 U37500 ( .A1(n52339), .A2(n52338), .Z(n59881) );
  NOR3_X2 U37501 ( .A1(n19496), .A2(n19500), .A3(n7475), .ZN(n60315) );
  XOR2_X1 U37508 ( .A1(n44219), .A2(n44183), .Z(n26191) );
  NAND2_X2 U37525 ( .A1(n59884), .A2(n11108), .ZN(n49951) );
  AND3_X1 U37530 ( .A1(n22148), .A2(n62760), .A3(n54464), .Z(n61341) );
  NAND2_X2 U37541 ( .A1(n40258), .A2(n40934), .ZN(n6276) );
  NAND2_X1 U37549 ( .A1(n33699), .A2(n33560), .ZN(n32525) );
  XOR2_X1 U37560 ( .A1(n51808), .A2(n19079), .Z(n51809) );
  XOR2_X1 U37564 ( .A1(n64102), .A2(n6740), .Z(n19079) );
  XOR2_X1 U37571 ( .A1(n11056), .A2(n11373), .Z(n14023) );
  NAND2_X1 U37573 ( .A1(n18550), .A2(n59890), .ZN(n14691) );
  NAND2_X1 U37580 ( .A1(n19804), .A2(n63913), .ZN(n59890) );
  NOR2_X2 U37604 ( .A1(n24797), .A2(n16109), .ZN(n50271) );
  AOI21_X1 U37607 ( .A1(n45512), .A2(n59893), .B(n59892), .ZN(n16200) );
  OR2_X1 U37617 ( .A1(n45513), .A2(n46906), .Z(n59893) );
  XOR2_X1 U37621 ( .A1(n45129), .A2(n9249), .Z(n60065) );
  XOR2_X1 U37625 ( .A1(n31584), .A2(n31684), .Z(n26127) );
  NAND3_X2 U37628 ( .A1(n45158), .A2(n45159), .A3(n45157), .ZN(n45160) );
  XOR2_X1 U37630 ( .A1(n17365), .A2(n59894), .Z(n14466) );
  XOR2_X1 U37640 ( .A1(n24663), .A2(n24662), .Z(n59894) );
  NOR2_X2 U37646 ( .A1(n8495), .A2(n8496), .ZN(n19803) );
  NAND3_X2 U37672 ( .A1(n12001), .A2(n50100), .A3(n61612), .ZN(n50521) );
  XOR2_X1 U37674 ( .A1(n23096), .A2(n33139), .Z(n31815) );
  NAND2_X1 U37691 ( .A1(n59899), .A2(n50092), .ZN(n46833) );
  OAI21_X1 U37695 ( .A1(n23650), .A2(n61612), .B(n59900), .ZN(n59899) );
  NAND4_X1 U37702 ( .A1(n28207), .A2(n31114), .A3(n10102), .A4(n31118), .ZN(
        n19001) );
  XOR2_X1 U37703 ( .A1(n11322), .A2(n12716), .Z(n51163) );
  NOR4_X2 U37709 ( .A1(n17189), .A2(n5385), .A3(n32861), .A4(n32860), .ZN(
        n5384) );
  BUF_X2 U37727 ( .I(n29639), .Z(n59903) );
  XOR2_X1 U37730 ( .A1(n59904), .A2(n59905), .Z(n61067) );
  XOR2_X1 U37756 ( .A1(n22922), .A2(n9084), .Z(n52416) );
  NOR2_X2 U37759 ( .A1(n26089), .A2(n53001), .ZN(n6792) );
  NAND2_X1 U37787 ( .A1(n49721), .A2(n47932), .ZN(n21490) );
  NAND2_X2 U37817 ( .A1(n15386), .A2(n46850), .ZN(n49721) );
  XOR2_X1 U37822 ( .A1(n52602), .A2(n23841), .Z(n10477) );
  XOR2_X1 U37823 ( .A1(n6596), .A2(n6595), .Z(n52602) );
  BUF_X2 U37832 ( .I(n19863), .Z(n59909) );
  XOR2_X1 U37840 ( .A1(n59911), .A2(n60118), .Z(n7961) );
  XOR2_X1 U37842 ( .A1(n18468), .A2(n22975), .Z(n8159) );
  AOI21_X1 U37846 ( .A1(n57370), .A2(n59914), .B(n54282), .ZN(n54284) );
  NAND2_X2 U37848 ( .A1(n31216), .A2(n30312), .ZN(n10926) );
  INV_X2 U37850 ( .I(n59915), .ZN(n30312) );
  NOR2_X2 U37853 ( .A1(n19929), .A2(n1218), .ZN(n59915) );
  NAND2_X1 U37858 ( .A1(n35143), .A2(n35971), .ZN(n59916) );
  AND3_X1 U37894 ( .A1(n7697), .A2(n54459), .A3(n55024), .Z(n22150) );
  NAND2_X1 U37896 ( .A1(n60415), .A2(n34798), .ZN(n33469) );
  NAND2_X2 U37902 ( .A1(n5322), .A2(n61261), .ZN(n60415) );
  XOR2_X1 U37903 ( .A1(n20707), .A2(n59923), .Z(n2923) );
  XNOR2_X1 U37908 ( .A1(n17060), .A2(n51647), .ZN(n39) );
  NOR3_X2 U37922 ( .A1(n24541), .A2(n24540), .A3(n32221), .ZN(n24539) );
  AOI21_X2 U37931 ( .A1(n60518), .A2(n29179), .B(n59934), .ZN(n25940) );
  XOR2_X1 U37942 ( .A1(n8540), .A2(n38221), .Z(n41920) );
  XOR2_X1 U37943 ( .A1(n1239), .A2(n3527), .Z(n38221) );
  NOR2_X2 U37947 ( .A1(n1212), .A2(n11380), .ZN(n61191) );
  AOI21_X1 U37953 ( .A1(n47765), .A2(n3281), .B(n17446), .ZN(n8724) );
  INV_X1 U37966 ( .I(n6369), .ZN(n29635) );
  NAND2_X1 U37967 ( .A1(n59935), .A2(n6369), .ZN(n6514) );
  NAND2_X2 U37969 ( .A1(n26856), .A2(n24418), .ZN(n6369) );
  INV_X2 U37970 ( .I(n6513), .ZN(n59935) );
  XOR2_X1 U37975 ( .A1(n7009), .A2(n7008), .Z(n59936) );
  NOR2_X1 U37979 ( .A1(n37902), .A2(n40797), .ZN(n59937) );
  XOR2_X1 U37992 ( .A1(n25174), .A2(n59938), .Z(n6605) );
  NOR2_X1 U37998 ( .A1(n60134), .A2(n24808), .ZN(n24810) );
  NAND3_X1 U38001 ( .A1(n59939), .A2(n25767), .A3(n54528), .ZN(n19140) );
  INV_X4 U38007 ( .I(n12592), .ZN(n6581) );
  NAND3_X2 U38017 ( .A1(n21851), .A2(n8290), .A3(n62461), .ZN(n16713) );
  NAND2_X1 U38023 ( .A1(n43441), .A2(n9366), .ZN(n59940) );
  AND2_X2 U38026 ( .A1(n12702), .A2(n20770), .Z(n53455) );
  XOR2_X1 U38028 ( .A1(n59941), .A2(n58234), .Z(n9882) );
  XOR2_X1 U38031 ( .A1(n24919), .A2(n31440), .Z(n59941) );
  XOR2_X1 U38033 ( .A1(n10823), .A2(n22363), .Z(n15291) );
  AND2_X1 U38034 ( .A1(n53244), .A2(n53251), .Z(n6949) );
  AND2_X1 U38038 ( .A1(n34666), .A2(n64461), .Z(n34525) );
  NAND2_X2 U38051 ( .A1(n59942), .A2(n12577), .ZN(n25021) );
  NAND2_X1 U38052 ( .A1(n59943), .A2(n16546), .ZN(n16547) );
  XOR2_X1 U38062 ( .A1(n59944), .A2(n45033), .Z(n586) );
  OR2_X1 U38080 ( .A1(n43816), .A2(n41779), .Z(n59945) );
  XOR2_X1 U38083 ( .A1(n10017), .A2(n37556), .Z(n9400) );
  NAND2_X2 U38094 ( .A1(n28073), .A2(n59102), .ZN(n60020) );
  NAND2_X2 U38110 ( .A1(n28663), .A2(n28677), .ZN(n19787) );
  NOR2_X2 U38111 ( .A1(n28600), .A2(n19788), .ZN(n28663) );
  NAND2_X2 U38118 ( .A1(n59962), .A2(n9240), .ZN(n6365) );
  BUF_X2 U38129 ( .I(n1664), .Z(n59967) );
  AOI22_X1 U38133 ( .A1(n53778), .A2(n53829), .B1(n53776), .B2(n53777), .ZN(
        n53785) );
  OAI21_X1 U38155 ( .A1(n53030), .A2(n53031), .B(n54348), .ZN(n53032) );
  INV_X1 U38161 ( .I(n59968), .ZN(n11667) );
  INV_X2 U38166 ( .I(n59969), .ZN(n6726) );
  XOR2_X1 U38170 ( .A1(Ciphertext[174]), .A2(Key[55]), .Z(n59969) );
  NOR2_X2 U38173 ( .A1(n27223), .A2(n27222), .ZN(n18738) );
  NOR2_X2 U38178 ( .A1(n59972), .A2(n23058), .ZN(n30311) );
  OR2_X1 U38185 ( .A1(n28830), .A2(n28829), .Z(n59972) );
  XOR2_X1 U38188 ( .A1(n24416), .A2(n22053), .Z(n19299) );
  NOR2_X1 U38196 ( .A1(n28309), .A2(n27080), .ZN(n9364) );
  OR2_X1 U38199 ( .A1(n49272), .A2(n21367), .Z(n59975) );
  OR2_X2 U38205 ( .A1(n21856), .A2(n2409), .Z(n22029) );
  NOR2_X1 U38222 ( .A1(n31044), .A2(n31045), .ZN(n31048) );
  BUF_X4 U38223 ( .I(n30558), .Z(n60895) );
  NOR2_X2 U38224 ( .A1(n14906), .A2(n61555), .ZN(n60930) );
  NOR2_X1 U38229 ( .A1(n9858), .A2(n59979), .ZN(n545) );
  NOR2_X1 U38235 ( .A1(n42786), .A2(n42787), .ZN(n59979) );
  OAI21_X2 U38261 ( .A1(n47535), .A2(n48604), .B(n12225), .ZN(n59983) );
  NAND2_X2 U38267 ( .A1(n59987), .A2(n9834), .ZN(n30584) );
  INV_X4 U38277 ( .I(n59988), .ZN(n11413) );
  NAND2_X2 U38293 ( .A1(n5289), .A2(n26454), .ZN(n59989) );
  OR2_X1 U38299 ( .A1(n2761), .A2(n59468), .Z(n35128) );
  NAND2_X2 U38302 ( .A1(n18410), .A2(n18479), .ZN(n7331) );
  XOR2_X1 U38312 ( .A1(n2862), .A2(n2861), .Z(n59991) );
  NOR2_X1 U38313 ( .A1(n60226), .A2(n10969), .ZN(n1157) );
  OAI22_X1 U38315 ( .A1(n48212), .A2(n48194), .B1(n48193), .B2(n8842), .ZN(
        n59992) );
  NOR2_X2 U38322 ( .A1(n18240), .A2(n38023), .ZN(n205) );
  NOR2_X1 U38323 ( .A1(n4322), .A2(n22282), .ZN(n42656) );
  NAND2_X1 U38338 ( .A1(n55811), .A2(n24958), .ZN(n55815) );
  NAND2_X2 U38344 ( .A1(n55828), .A2(n55812), .ZN(n55811) );
  XOR2_X1 U38354 ( .A1(n31815), .A2(n31344), .Z(n60392) );
  OR2_X1 U38358 ( .A1(n7728), .A2(n42252), .Z(n42248) );
  NOR2_X2 U38360 ( .A1(n27304), .A2(n27303), .ZN(n27305) );
  XOR2_X1 U38362 ( .A1(n21891), .A2(n18518), .Z(n60559) );
  XOR2_X1 U38375 ( .A1(n8078), .A2(n1188), .Z(n21891) );
  NOR2_X1 U38377 ( .A1(n49544), .A2(n18821), .ZN(n18820) );
  OAI22_X1 U38378 ( .A1(n27651), .A2(n27650), .B1(n63330), .B2(n6273), .ZN(
        n59994) );
  XOR2_X1 U38389 ( .A1(n20403), .A2(n22296), .Z(n12102) );
  XOR2_X1 U38398 ( .A1(n60001), .A2(n32093), .Z(n22841) );
  XOR2_X1 U38399 ( .A1(n32315), .A2(n7390), .Z(n60001) );
  BUF_X2 U38401 ( .I(n148), .Z(n60002) );
  NOR2_X1 U38404 ( .A1(n6075), .A2(n53498), .ZN(n60798) );
  NAND2_X1 U38406 ( .A1(n34572), .A2(n34573), .ZN(n21610) );
  NAND2_X1 U38409 ( .A1(n14463), .A2(n32965), .ZN(n34572) );
  INV_X2 U38416 ( .I(n42845), .ZN(n60006) );
  NOR2_X2 U38422 ( .A1(n60006), .A2(n58210), .ZN(n1007) );
  NAND2_X2 U38427 ( .A1(n2059), .A2(n36422), .ZN(n36169) );
  NAND2_X1 U38431 ( .A1(n56519), .A2(n60008), .ZN(n56526) );
  OR2_X1 U38447 ( .A1(n56521), .A2(n56520), .Z(n60008) );
  XOR2_X1 U38452 ( .A1(n13936), .A2(n13937), .Z(n16755) );
  AND2_X1 U38472 ( .A1(n21203), .A2(n19712), .Z(n60011) );
  XOR2_X1 U38477 ( .A1(n60013), .A2(n60012), .Z(n23052) );
  XOR2_X1 U38478 ( .A1(n1548), .A2(n25190), .Z(n60012) );
  XOR2_X1 U38481 ( .A1(n23590), .A2(n22215), .Z(n60013) );
  XNOR2_X1 U38484 ( .A1(n18571), .A2(n21503), .ZN(n33837) );
  NAND2_X2 U38493 ( .A1(n1571), .A2(n26391), .ZN(n18006) );
  INV_X2 U38495 ( .I(n30177), .ZN(n30688) );
  NAND2_X2 U38497 ( .A1(n579), .A2(n30174), .ZN(n30177) );
  NOR2_X2 U38547 ( .A1(n7021), .A2(n53516), .ZN(n53527) );
  NOR2_X2 U38549 ( .A1(n60018), .A2(n17453), .ZN(n37563) );
  NAND2_X1 U38550 ( .A1(n9744), .A2(n32986), .ZN(n60018) );
  NAND2_X2 U38551 ( .A1(n48252), .A2(n7834), .ZN(n20624) );
  INV_X2 U38556 ( .I(n60019), .ZN(n28244) );
  XNOR2_X1 U38567 ( .A1(Ciphertext[49]), .A2(Key[44]), .ZN(n60019) );
  XOR2_X1 U38582 ( .A1(n44638), .A2(n44637), .Z(n22941) );
  NAND2_X2 U38583 ( .A1(n22391), .A2(n1482), .ZN(n18127) );
  XOR2_X1 U38584 ( .A1(n673), .A2(n44628), .Z(n44630) );
  BUF_X2 U38586 ( .I(n18205), .Z(n60022) );
  XOR2_X1 U38596 ( .A1(n31336), .A2(n3070), .Z(n3072) );
  NAND4_X1 U38597 ( .A1(n13798), .A2(n10971), .A3(n25924), .A4(n10824), .ZN(
        n42385) );
  NOR2_X2 U38604 ( .A1(n35691), .A2(n33600), .ZN(n60456) );
  INV_X1 U38625 ( .I(n41531), .ZN(n60026) );
  NAND2_X2 U38629 ( .A1(n56624), .A2(n21893), .ZN(n56214) );
  NAND3_X2 U38630 ( .A1(n46052), .A2(n44653), .A3(n44652), .ZN(n44654) );
  XOR2_X1 U38632 ( .A1(n7684), .A2(n44193), .Z(n46912) );
  NOR3_X2 U38636 ( .A1(n1417), .A2(n12863), .A3(n36742), .ZN(n36747) );
  NAND2_X2 U38637 ( .A1(n20755), .A2(n29452), .ZN(n29451) );
  OR2_X1 U38679 ( .A1(n41256), .A2(n60826), .Z(n41259) );
  OR2_X1 U38684 ( .A1(n29453), .A2(n29452), .Z(n60031) );
  INV_X2 U38694 ( .I(n60034), .ZN(n36029) );
  NOR3_X2 U38695 ( .A1(n60891), .A2(n21328), .A3(n61066), .ZN(n60034) );
  NAND2_X1 U38718 ( .A1(n18108), .A2(n55685), .ZN(n60045) );
  AOI22_X1 U38719 ( .A1(n52988), .A2(n54307), .B1(n52989), .B2(n52990), .ZN(
        n60046) );
  XOR2_X1 U38723 ( .A1(n63040), .A2(n3517), .Z(n1051) );
  XOR2_X1 U38730 ( .A1(n2126), .A2(n2125), .Z(n15739) );
  XOR2_X1 U38738 ( .A1(n3479), .A2(n38755), .Z(n60050) );
  NAND2_X2 U38749 ( .A1(n27236), .A2(n60055), .ZN(n29457) );
  NOR2_X1 U38755 ( .A1(n60058), .A2(n60056), .ZN(n60055) );
  NOR2_X1 U38758 ( .A1(n27226), .A2(n25786), .ZN(n60058) );
  NAND3_X1 U38783 ( .A1(n36067), .A2(n36069), .A3(n36068), .ZN(n36071) );
  NAND2_X1 U38829 ( .A1(n33434), .A2(n33433), .ZN(n10885) );
  NAND2_X2 U38842 ( .A1(n41717), .A2(n1269), .ZN(n42915) );
  XOR2_X1 U38843 ( .A1(n22848), .A2(n940), .Z(n4991) );
  NOR2_X2 U38852 ( .A1(n2994), .A2(n43573), .ZN(n42724) );
  NAND2_X2 U38862 ( .A1(n33945), .A2(n32795), .ZN(n34117) );
  NAND2_X2 U38864 ( .A1(n33948), .A2(n25972), .ZN(n33945) );
  NAND2_X2 U38876 ( .A1(n31074), .A2(n31077), .ZN(n23708) );
  XOR2_X1 U38878 ( .A1(n60065), .A2(n16195), .Z(n21067) );
  XOR2_X1 U38883 ( .A1(n44947), .A2(n2540), .Z(n45342) );
  NOR3_X2 U38887 ( .A1(n17578), .A2(n17575), .A3(n17574), .ZN(n43166) );
  NAND2_X2 U38892 ( .A1(n25333), .A2(n61731), .ZN(n32870) );
  NAND3_X2 U38895 ( .A1(n3393), .A2(n60070), .A3(n6107), .ZN(n5726) );
  INV_X1 U38898 ( .I(n60071), .ZN(n60070) );
  AOI22_X1 U38902 ( .A1(n11967), .A2(n14641), .B1(n28682), .B2(n59096), .ZN(
        n60071) );
  XOR2_X1 U38903 ( .A1(n4844), .A2(n60072), .Z(n50723) );
  XOR2_X1 U38909 ( .A1(n18466), .A2(n50997), .Z(n60072) );
  NAND2_X2 U38910 ( .A1(n3368), .A2(n2766), .ZN(n4380) );
  XOR2_X1 U38911 ( .A1(n60074), .A2(n60073), .Z(n2767) );
  XOR2_X1 U38912 ( .A1(n44021), .A2(n44020), .Z(n60074) );
  NAND2_X2 U38916 ( .A1(n25632), .A2(n61261), .ZN(n60960) );
  NOR2_X2 U38924 ( .A1(n60076), .A2(n60075), .ZN(n978) );
  INV_X1 U38931 ( .I(n27384), .ZN(n27385) );
  NAND2_X1 U38934 ( .A1(n28241), .A2(n27043), .ZN(n27384) );
  NAND2_X2 U38935 ( .A1(n49400), .A2(n60078), .ZN(n14034) );
  AOI22_X2 U38948 ( .A1(n49397), .A2(n49396), .B1(n49399), .B2(n49398), .ZN(
        n60078) );
  NAND2_X2 U38956 ( .A1(n25381), .A2(n60081), .ZN(n125) );
  NOR2_X2 U38957 ( .A1(n28578), .A2(n26231), .ZN(n60081) );
  NAND2_X2 U38963 ( .A1(n32528), .A2(n33561), .ZN(n33564) );
  NAND2_X1 U38964 ( .A1(n55431), .A2(n8969), .ZN(n8965) );
  NAND2_X1 U38965 ( .A1(n60082), .A2(n43375), .ZN(n3787) );
  NOR2_X1 U38966 ( .A1(n42756), .A2(n65228), .ZN(n60082) );
  NAND3_X1 U38968 ( .A1(n24578), .A2(n4086), .A3(n45718), .ZN(n44552) );
  NAND2_X2 U38974 ( .A1(n45716), .A2(n1666), .ZN(n24578) );
  XOR2_X1 U39004 ( .A1(n60086), .A2(n50884), .Z(n10501) );
  NAND3_X2 U39005 ( .A1(n14245), .A2(n16576), .A3(n16578), .ZN(n35030) );
  OR2_X1 U39007 ( .A1(n205), .A2(n39095), .Z(n40514) );
  XOR2_X1 U39011 ( .A1(n31977), .A2(n17092), .Z(n60087) );
  NAND2_X2 U39030 ( .A1(n19567), .A2(n19556), .ZN(n6351) );
  INV_X2 U39049 ( .I(n6607), .ZN(n1646) );
  NAND2_X2 U39056 ( .A1(n9972), .A2(n1648), .ZN(n6607) );
  XOR2_X1 U39062 ( .A1(n23426), .A2(n43909), .Z(n44829) );
  NAND2_X1 U39065 ( .A1(n60088), .A2(n1163), .ZN(n53271) );
  OAI21_X1 U39067 ( .A1(n9943), .A2(n53279), .B(n53296), .ZN(n60088) );
  XOR2_X1 U39086 ( .A1(n13152), .A2(n13151), .Z(n61072) );
  NOR2_X1 U39092 ( .A1(n3900), .A2(n3902), .ZN(n3899) );
  NOR2_X2 U39098 ( .A1(n5658), .A2(n56867), .ZN(n5585) );
  NAND2_X1 U39102 ( .A1(n55899), .A2(n55854), .ZN(n55851) );
  NOR2_X2 U39106 ( .A1(n17774), .A2(n55896), .ZN(n55899) );
  NOR2_X2 U39115 ( .A1(n61181), .A2(n60093), .ZN(n5017) );
  NAND2_X1 U39116 ( .A1(n52046), .A2(n57293), .ZN(n51965) );
  XOR2_X1 U39125 ( .A1(n52544), .A2(n60531), .Z(n19103) );
  XOR2_X1 U39126 ( .A1(n60094), .A2(n8932), .Z(n8931) );
  AOI22_X1 U39128 ( .A1(n29031), .A2(n29030), .B1(n13481), .B2(n29032), .ZN(
        n60095) );
  NAND2_X1 U39181 ( .A1(n50332), .A2(n50339), .ZN(n60099) );
  INV_X1 U39189 ( .I(n50769), .ZN(n8276) );
  NAND3_X2 U39192 ( .A1(n49120), .A2(n49121), .A3(n49119), .ZN(n50769) );
  NOR3_X1 U39194 ( .A1(n54422), .A2(n54421), .A3(n54420), .ZN(n60104) );
  XOR2_X1 U39198 ( .A1(n39224), .A2(n60106), .Z(n16372) );
  XOR2_X1 U39199 ( .A1(n38159), .A2(n5841), .Z(n60106) );
  XOR2_X1 U39203 ( .A1(n6322), .A2(n8952), .Z(n16502) );
  NAND2_X2 U39230 ( .A1(n18063), .A2(n54507), .ZN(n25172) );
  XOR2_X1 U39236 ( .A1(n60114), .A2(n4990), .Z(n146) );
  NAND2_X1 U39240 ( .A1(n61398), .A2(n41946), .ZN(n60116) );
  NOR2_X1 U39246 ( .A1(n4748), .A2(n60578), .ZN(n13860) );
  BUF_X4 U39253 ( .I(n36026), .Z(n60891) );
  NAND3_X1 U39256 ( .A1(n25488), .A2(n35536), .A3(n32979), .ZN(n17453) );
  XOR2_X1 U39267 ( .A1(n60119), .A2(n13635), .Z(n13383) );
  OAI22_X2 U39276 ( .A1(n17343), .A2(n17457), .B1(n28803), .B2(n28802), .ZN(
        n60121) );
  AND2_X1 U39277 ( .A1(n18678), .A2(n13141), .Z(n60122) );
  XOR2_X1 U39292 ( .A1(n3258), .A2(n60124), .Z(n3257) );
  INV_X2 U39303 ( .I(n60125), .ZN(n61503) );
  NAND3_X2 U39311 ( .A1(n25738), .A2(n25737), .A3(n7142), .ZN(n60125) );
  NAND2_X2 U39312 ( .A1(n19609), .A2(n19610), .ZN(n34603) );
  NAND2_X2 U39313 ( .A1(n60126), .A2(n15229), .ZN(n61087) );
  NAND2_X1 U39314 ( .A1(n19603), .A2(n19602), .ZN(n60126) );
  INV_X2 U39318 ( .I(n42686), .ZN(n1686) );
  NOR2_X2 U39348 ( .A1(n42499), .A2(n41850), .ZN(n11079) );
  XOR2_X1 U39353 ( .A1(n32649), .A2(n32648), .Z(n32650) );
  XOR2_X1 U39354 ( .A1(n31867), .A2(n14129), .Z(n32649) );
  AOI21_X2 U39377 ( .A1(n22627), .A2(n7964), .B(n60130), .ZN(n5855) );
  OAI22_X2 U39379 ( .A1(n12247), .A2(n5857), .B1(n24172), .B2(n24171), .ZN(
        n60130) );
  BUF_X2 U39392 ( .I(n64367), .Z(n60132) );
  NAND3_X1 U39395 ( .A1(n24807), .A2(n22990), .A3(n56177), .ZN(n60134) );
  NOR2_X2 U39416 ( .A1(n2005), .A2(n18129), .ZN(n30787) );
  INV_X2 U39426 ( .I(n21699), .ZN(n33643) );
  NAND2_X2 U39454 ( .A1(n30771), .A2(n30767), .ZN(n29743) );
  NAND4_X2 U39461 ( .A1(n8344), .A2(n8346), .A3(n34074), .A4(n34075), .ZN(
        n17202) );
  NAND2_X1 U39464 ( .A1(n22089), .A2(n43676), .ZN(n22088) );
  XOR2_X1 U39467 ( .A1(n46579), .A2(n46589), .Z(n24593) );
  AND3_X1 U39473 ( .A1(n34751), .A2(n34750), .A3(n34749), .Z(n60621) );
  NAND2_X2 U39475 ( .A1(n37050), .A2(n35990), .ZN(n37957) );
  XOR2_X1 U39476 ( .A1(n2876), .A2(n11318), .Z(n25754) );
  NAND2_X2 U39478 ( .A1(n6170), .A2(n39904), .ZN(n41806) );
  OAI21_X2 U39492 ( .A1(n60145), .A2(n60144), .B(n59616), .ZN(n14771) );
  AND2_X1 U39500 ( .A1(n30237), .A2(n26740), .Z(n4735) );
  INV_X4 U39508 ( .I(n60147), .ZN(n15805) );
  NAND3_X2 U39512 ( .A1(n10137), .A2(n21908), .A3(n21909), .ZN(n60147) );
  XOR2_X1 U39513 ( .A1(n6037), .A2(n44328), .Z(n60148) );
  INV_X1 U39515 ( .I(n36554), .ZN(n36563) );
  NAND2_X1 U39523 ( .A1(n23215), .A2(n36377), .ZN(n36554) );
  NOR2_X2 U39537 ( .A1(n9532), .A2(n48349), .ZN(n48894) );
  NAND2_X2 U39546 ( .A1(n60149), .A2(n6462), .ZN(n25510) );
  NOR2_X2 U39551 ( .A1(n56562), .A2(n56666), .ZN(n56687) );
  AND2_X2 U39555 ( .A1(n12810), .A2(n51557), .Z(n56234) );
  XNOR2_X1 U39564 ( .A1(n33862), .A2(n33034), .ZN(n24672) );
  XOR2_X1 U39567 ( .A1(n15153), .A2(n6544), .Z(n15186) );
  XOR2_X1 U39579 ( .A1(n7065), .A2(n60151), .Z(n972) );
  BUF_X2 U39580 ( .I(n1426), .Z(n60152) );
  AND2_X1 U39588 ( .A1(n27879), .A2(n27880), .Z(n60154) );
  XOR2_X1 U39597 ( .A1(n60156), .A2(n13545), .Z(n13544) );
  NOR2_X2 U39604 ( .A1(n48511), .A2(n48499), .ZN(n48506) );
  XOR2_X1 U39605 ( .A1(n60157), .A2(n1751), .Z(n12963) );
  AND2_X1 U39609 ( .A1(n60456), .A2(n4231), .Z(n12023) );
  INV_X4 U39615 ( .I(n60159), .ZN(n52762) );
  AND2_X2 U39616 ( .A1(n52760), .A2(n52761), .Z(n60159) );
  OR3_X1 U39620 ( .A1(n52845), .A2(n53602), .A3(n53605), .Z(n52757) );
  INV_X2 U39652 ( .I(n42102), .ZN(n42100) );
  XOR2_X1 U39676 ( .A1(n60941), .A2(n11233), .Z(n15201) );
  OR2_X1 U39681 ( .A1(n33126), .A2(n33125), .Z(n60161) );
  XOR2_X1 U39688 ( .A1(n33837), .A2(n32565), .Z(n32229) );
  XOR2_X1 U39689 ( .A1(n32206), .A2(n31654), .Z(n24279) );
  XOR2_X1 U39694 ( .A1(n14104), .A2(Key[79]), .Z(n28135) );
  NAND2_X2 U39697 ( .A1(n4547), .A2(n25328), .ZN(n25327) );
  XOR2_X1 U39703 ( .A1(n51960), .A2(n51959), .Z(n50660) );
  NOR2_X1 U39715 ( .A1(n11643), .A2(n34167), .ZN(n34170) );
  NAND2_X2 U39722 ( .A1(n15152), .A2(n24664), .ZN(n11643) );
  XOR2_X1 U39725 ( .A1(n33035), .A2(n30945), .Z(n25741) );
  NAND3_X2 U39726 ( .A1(n27428), .A2(n27427), .A3(n27426), .ZN(n30945) );
  INV_X1 U39730 ( .I(n60168), .ZN(n21715) );
  AOI21_X1 U39731 ( .A1(n5484), .A2(n873), .B(n14102), .ZN(n60168) );
  NAND3_X2 U39735 ( .A1(n30261), .A2(n30046), .A3(n2310), .ZN(n27423) );
  NAND2_X1 U39736 ( .A1(n33658), .A2(n60169), .ZN(n33668) );
  OAI21_X1 U39740 ( .A1(n33657), .A2(n33653), .B(n33652), .ZN(n60169) );
  NAND2_X2 U39751 ( .A1(n39102), .A2(n15101), .ZN(n19148) );
  OAI21_X1 U39754 ( .A1(n30744), .A2(n20172), .B(n13243), .ZN(n13030) );
  BUF_X2 U39761 ( .I(n27374), .Z(n60171) );
  XOR2_X1 U39790 ( .A1(n25641), .A2(n25642), .Z(n60174) );
  NAND2_X1 U39799 ( .A1(n5883), .A2(n5578), .ZN(n60715) );
  INV_X2 U39800 ( .I(n60176), .ZN(n12028) );
  NAND2_X1 U39807 ( .A1(n18592), .A2(n40622), .ZN(n16013) );
  NAND3_X2 U39825 ( .A1(n60554), .A2(n57268), .A3(n34658), .ZN(n25893) );
  AND3_X1 U39826 ( .A1(n30218), .A2(n2495), .A3(n21778), .Z(n60185) );
  NAND2_X1 U39828 ( .A1(n34798), .A2(n5322), .ZN(n12582) );
  XOR2_X1 U39830 ( .A1(n2975), .A2(n60186), .Z(n2974) );
  XOR2_X1 U39831 ( .A1(n32285), .A2(n13255), .Z(n60186) );
  BUF_X2 U39837 ( .I(n17872), .Z(n60187) );
  XOR2_X1 U39838 ( .A1(n15055), .A2(n15053), .Z(n60188) );
  NAND2_X1 U39840 ( .A1(n60189), .A2(n32459), .ZN(n7839) );
  NOR2_X2 U39842 ( .A1(n13981), .A2(n13980), .ZN(n13532) );
  NAND2_X2 U39844 ( .A1(n13533), .A2(n13534), .ZN(n13981) );
  XOR2_X1 U39854 ( .A1(n8074), .A2(n24388), .Z(n8306) );
  XOR2_X1 U39866 ( .A1(n60194), .A2(n38437), .Z(n11187) );
  OAI22_X1 U39872 ( .A1(n26424), .A2(n10239), .B1(n27851), .B2(n26834), .ZN(
        n26425) );
  NAND4_X2 U39880 ( .A1(n16799), .A2(n16887), .A3(n16888), .A4(n31660), .ZN(
        n16886) );
  OAI21_X1 U39881 ( .A1(n41030), .A2(n38496), .B(n60195), .ZN(n39093) );
  NAND2_X1 U39885 ( .A1(n41030), .A2(n39094), .ZN(n60195) );
  NAND3_X1 U39886 ( .A1(n53711), .A2(n53718), .A3(n21973), .ZN(n22021) );
  NOR2_X2 U39895 ( .A1(n57462), .A2(n64858), .ZN(n41193) );
  AOI21_X1 U39896 ( .A1(n28876), .A2(n4483), .B(n1875), .ZN(n4482) );
  NOR3_X2 U39899 ( .A1(n60198), .A2(n29289), .A3(n29288), .ZN(n12361) );
  NOR2_X1 U39900 ( .A1(n2957), .A2(n54119), .ZN(n54124) );
  NOR2_X1 U39902 ( .A1(n58806), .A2(n51606), .ZN(n13218) );
  NOR2_X2 U39915 ( .A1(n28875), .A2(n60199), .ZN(n30761) );
  NAND3_X2 U39923 ( .A1(n10918), .A2(n10920), .A3(n10917), .ZN(n60199) );
  NAND2_X2 U39927 ( .A1(n60200), .A2(n57192), .ZN(n11041) );
  NOR2_X1 U39942 ( .A1(n49930), .A2(n49931), .ZN(n60201) );
  OAI21_X1 U39956 ( .A1(n56592), .A2(n56593), .B(n56591), .ZN(n56594) );
  NAND2_X2 U39966 ( .A1(n21957), .A2(n56585), .ZN(n56591) );
  BUF_X2 U39971 ( .I(n51891), .Z(n60203) );
  INV_X1 U39996 ( .I(n11866), .ZN(n60319) );
  XOR2_X1 U40029 ( .A1(n688), .A2(n15960), .Z(n60206) );
  XOR2_X1 U40031 ( .A1(n46531), .A2(n50999), .Z(n31511) );
  XOR2_X1 U40040 ( .A1(n37883), .A2(n36734), .Z(n46531) );
  AND2_X1 U40055 ( .A1(n50215), .A2(n50220), .Z(n49344) );
  NOR2_X1 U40067 ( .A1(n49353), .A2(n49354), .ZN(n7341) );
  NOR2_X1 U40069 ( .A1(n49352), .A2(n49351), .ZN(n49353) );
  XOR2_X1 U40080 ( .A1(n60212), .A2(n54888), .Z(Plaintext[85]) );
  BUF_X2 U40083 ( .I(n30526), .Z(n60214) );
  NAND2_X2 U40089 ( .A1(n3364), .A2(n1667), .ZN(n60839) );
  NOR2_X2 U40098 ( .A1(n60216), .A2(n60215), .ZN(n6797) );
  NAND4_X2 U40099 ( .A1(n9870), .A2(n41136), .A3(n41135), .A4(n41137), .ZN(
        n60215) );
  INV_X2 U40106 ( .I(n53632), .ZN(n53692) );
  NAND3_X2 U40111 ( .A1(n11870), .A2(n11868), .A3(n53627), .ZN(n53632) );
  NAND3_X1 U40114 ( .A1(n52409), .A2(n14676), .A3(n48023), .ZN(n9207) );
  NAND2_X2 U40121 ( .A1(n25348), .A2(n16954), .ZN(n10077) );
  OR2_X1 U40126 ( .A1(n35532), .A2(n36567), .Z(n32981) );
  NAND4_X2 U40152 ( .A1(n35503), .A2(n35501), .A3(n18509), .A4(n35502), .ZN(
        n13322) );
  AND2_X1 U40170 ( .A1(n41232), .A2(n60132), .Z(n15342) );
  XOR2_X1 U40177 ( .A1(n32307), .A2(n32306), .Z(n13508) );
  XOR2_X1 U40185 ( .A1(n38967), .A2(n60220), .Z(n307) );
  XOR2_X1 U40192 ( .A1(n11474), .A2(n60221), .Z(n60220) );
  NAND3_X1 U40194 ( .A1(n60757), .A2(n14924), .A3(n60222), .ZN(n9833) );
  OAI22_X1 U40204 ( .A1(n28186), .A2(n28183), .B1(n28184), .B2(n28646), .ZN(
        n60222) );
  NAND4_X2 U40218 ( .A1(n3131), .A2(n20550), .A3(n3132), .A4(n3130), .ZN(
        n20548) );
  NAND3_X1 U40221 ( .A1(n60224), .A2(n48179), .A3(n48180), .ZN(n48182) );
  OAI21_X1 U40223 ( .A1(n8043), .A2(n46177), .B(n60687), .ZN(n60224) );
  OR2_X1 U40228 ( .A1(n38675), .A2(n40729), .Z(n41195) );
  NOR2_X2 U40255 ( .A1(n7705), .A2(n1531), .ZN(n7656) );
  INV_X4 U40257 ( .I(n36435), .ZN(n7705) );
  NAND2_X2 U40261 ( .A1(n52828), .A2(n25936), .ZN(n60225) );
  INV_X2 U40268 ( .I(n60226), .ZN(n1158) );
  NAND2_X2 U40269 ( .A1(n9160), .A2(n1459), .ZN(n60226) );
  XOR2_X1 U40270 ( .A1(n60228), .A2(n2935), .Z(n61091) );
  NAND2_X2 U40280 ( .A1(n14397), .A2(n21457), .ZN(n9885) );
  NAND3_X2 U40319 ( .A1(n20565), .A2(n45303), .A3(n20567), .ZN(n45304) );
  INV_X2 U40321 ( .I(n60233), .ZN(n45267) );
  XOR2_X1 U40337 ( .A1(n44524), .A2(n45265), .Z(n60233) );
  XOR2_X1 U40342 ( .A1(n23305), .A2(n7506), .Z(n44524) );
  NOR2_X2 U40345 ( .A1(n33662), .A2(n31701), .ZN(n262) );
  XOR2_X1 U40351 ( .A1(n60234), .A2(n13914), .Z(n30367) );
  NAND2_X2 U40372 ( .A1(n6989), .A2(n6990), .ZN(n18276) );
  NAND2_X1 U40380 ( .A1(n8669), .A2(n1528), .ZN(n35980) );
  NOR4_X2 U40382 ( .A1(n26934), .A2(n26931), .A3(n26933), .A4(n26932), .ZN(
        n27003) );
  NOR2_X1 U40385 ( .A1(n7464), .A2(n8826), .ZN(n7463) );
  NOR2_X2 U40394 ( .A1(n47712), .A2(n47713), .ZN(n49548) );
  NAND3_X1 U40407 ( .A1(n55958), .A2(n56591), .A3(n20737), .ZN(n60236) );
  NOR2_X2 U40420 ( .A1(n60237), .A2(n15115), .ZN(n30648) );
  XOR2_X1 U40433 ( .A1(n60238), .A2(n20554), .Z(n15292) );
  XOR2_X1 U40442 ( .A1(n25042), .A2(n32746), .Z(n60238) );
  INV_X2 U40447 ( .I(n4326), .ZN(n32782) );
  OR2_X1 U40448 ( .A1(n42040), .A2(n13678), .Z(n42037) );
  INV_X2 U40457 ( .I(n60241), .ZN(n25166) );
  NOR2_X2 U40460 ( .A1(n30583), .A2(n30584), .ZN(n24064) );
  AOI22_X1 U40464 ( .A1(n47561), .A2(n60242), .B1(n45216), .B2(n23361), .ZN(
        n45220) );
  NOR2_X1 U40469 ( .A1(n59119), .A2(n64944), .ZN(n60242) );
  NAND2_X2 U40471 ( .A1(n60243), .A2(n57341), .ZN(n18018) );
  XOR2_X1 U40489 ( .A1(n15398), .A2(n60251), .Z(n24579) );
  XOR2_X1 U40491 ( .A1(n6031), .A2(n44606), .Z(n60251) );
  OAI21_X1 U40498 ( .A1(n18085), .A2(n18086), .B(n17833), .ZN(n60252) );
  NOR2_X1 U40503 ( .A1(n20464), .A2(n28185), .ZN(n60757) );
  XOR2_X1 U40517 ( .A1(n46288), .A2(n23722), .Z(n3573) );
  NAND2_X2 U40522 ( .A1(n14658), .A2(n14657), .ZN(n46549) );
  NAND2_X2 U40545 ( .A1(n1334), .A2(n1495), .ZN(n43305) );
  NOR2_X2 U40552 ( .A1(n40020), .A2(n43444), .ZN(n43446) );
  INV_X4 U40553 ( .I(n25458), .ZN(n43444) );
  NAND2_X1 U40567 ( .A1(n56462), .A2(n56445), .ZN(n60256) );
  NAND2_X2 U40571 ( .A1(n60258), .A2(n34272), .ZN(n13126) );
  XOR2_X1 U40578 ( .A1(n50519), .A2(n13155), .Z(n349) );
  XOR2_X1 U40584 ( .A1(n10502), .A2(n48955), .Z(n50519) );
  XOR2_X1 U40589 ( .A1(n32357), .A2(n32504), .Z(n6484) );
  XOR2_X1 U40591 ( .A1(n5342), .A2(n3798), .Z(n32504) );
  XOR2_X1 U40600 ( .A1(n13286), .A2(n51601), .Z(n52030) );
  XOR2_X1 U40602 ( .A1(n60261), .A2(n3570), .Z(n24697) );
  NAND3_X2 U40606 ( .A1(n54971), .A2(n54970), .A3(n51779), .ZN(n54977) );
  NAND2_X2 U40608 ( .A1(n23766), .A2(n1528), .ZN(n20146) );
  BUF_X2 U40610 ( .I(n1318), .Z(n60262) );
  NOR2_X2 U40626 ( .A1(n28400), .A2(n3117), .ZN(n243) );
  XOR2_X1 U40629 ( .A1(n60267), .A2(n37632), .Z(n13581) );
  XOR2_X1 U40630 ( .A1(n63011), .A2(n61489), .Z(n60267) );
  NAND3_X2 U40632 ( .A1(n60467), .A2(n21870), .A3(n49972), .ZN(n50337) );
  NAND2_X2 U40638 ( .A1(n14624), .A2(n15934), .ZN(n41887) );
  OR2_X1 U40641 ( .A1(n30082), .A2(n60270), .Z(n30091) );
  NOR2_X1 U40642 ( .A1(n30084), .A2(n23111), .ZN(n60270) );
  NOR2_X2 U40645 ( .A1(n27915), .A2(n29015), .ZN(n30082) );
  XOR2_X1 U40662 ( .A1(n26202), .A2(n11050), .Z(n32486) );
  NOR2_X2 U40668 ( .A1(n40656), .A2(n40662), .ZN(n40484) );
  NAND2_X1 U40674 ( .A1(n56848), .A2(n56868), .ZN(n56820) );
  NOR2_X2 U40680 ( .A1(n21879), .A2(n56894), .ZN(n56868) );
  NOR3_X2 U40684 ( .A1(n60276), .A2(n11349), .A3(n60275), .ZN(n11348) );
  AOI21_X1 U40695 ( .A1(n4573), .A2(n1502), .B(n60951), .ZN(n22831) );
  NAND2_X2 U40696 ( .A1(n2541), .A2(n49681), .ZN(n60279) );
  NOR2_X2 U40708 ( .A1(n60280), .A2(n61314), .ZN(n17015) );
  XOR2_X1 U40713 ( .A1(n5685), .A2(n4278), .Z(n17201) );
  XOR2_X1 U40714 ( .A1(n2275), .A2(n60959), .Z(n20113) );
  XOR2_X1 U40733 ( .A1(n61927), .A2(n60282), .Z(n8882) );
  XOR2_X1 U40735 ( .A1(n8885), .A2(n8884), .Z(n60282) );
  INV_X2 U40736 ( .I(n60283), .ZN(n16938) );
  BUF_X2 U40737 ( .I(n27756), .Z(n60284) );
  XOR2_X1 U40743 ( .A1(n52154), .A2(n60287), .Z(n2264) );
  XOR2_X1 U40746 ( .A1(n51924), .A2(n51922), .Z(n60287) );
  INV_X1 U40749 ( .I(n60290), .ZN(n60289) );
  OAI21_X1 U40753 ( .A1(n36142), .A2(n60925), .B(n60291), .ZN(n60290) );
  XOR2_X1 U40769 ( .A1(n24048), .A2(n1756), .Z(n37966) );
  BUF_X4 U40784 ( .I(n44788), .Z(n49276) );
  NAND2_X1 U40787 ( .A1(n18185), .A2(n49284), .ZN(n18184) );
  AND2_X1 U40793 ( .A1(n28147), .A2(n27345), .Z(n61006) );
  XOR2_X1 U40803 ( .A1(n12122), .A2(n57378), .Z(n4369) );
  XOR2_X1 U40805 ( .A1(n21172), .A2(n11336), .Z(n12122) );
  BUF_X4 U40807 ( .I(n36595), .Z(n60297) );
  XOR2_X1 U40811 ( .A1(n52404), .A2(n60300), .Z(n2152) );
  NAND2_X2 U40812 ( .A1(n48359), .A2(n48358), .ZN(n52404) );
  NOR2_X1 U40813 ( .A1(n59203), .A2(n41211), .ZN(n41219) );
  NAND2_X1 U40820 ( .A1(n19124), .A2(n60301), .ZN(n356) );
  NOR2_X2 U40827 ( .A1(n1505), .A2(n6058), .ZN(n42302) );
  XOR2_X1 U40830 ( .A1(n17322), .A2(n14337), .Z(n60303) );
  INV_X2 U40855 ( .I(n60305), .ZN(n5377) );
  XOR2_X1 U40859 ( .A1(n39476), .A2(n3532), .Z(n3531) );
  OAI21_X1 U40871 ( .A1(n60306), .A2(n23068), .B(n28905), .ZN(n27761) );
  NOR2_X2 U40872 ( .A1(n28903), .A2(n1352), .ZN(n60306) );
  INV_X2 U40893 ( .I(n60309), .ZN(n17452) );
  AOI22_X1 U40895 ( .A1(n53051), .A2(n53050), .B1(n53052), .B2(n53053), .ZN(
        n53062) );
  OR2_X1 U40914 ( .A1(n47229), .A2(n9758), .Z(n44647) );
  NOR2_X2 U40917 ( .A1(n23643), .A2(n6747), .ZN(n47229) );
  XOR2_X1 U40920 ( .A1(n10749), .A2(n26107), .Z(n148) );
  XOR2_X1 U40922 ( .A1(n60314), .A2(n51528), .Z(n25997) );
  XOR2_X1 U40923 ( .A1(n18308), .A2(n9342), .Z(n60314) );
  NOR2_X2 U40928 ( .A1(n50369), .A2(n24134), .ZN(n49991) );
  NAND2_X2 U40934 ( .A1(n19493), .A2(n60315), .ZN(n19491) );
  XOR2_X1 U40939 ( .A1(n60316), .A2(n61149), .Z(n12380) );
  XOR2_X1 U40940 ( .A1(n5729), .A2(n12381), .Z(n60316) );
  AND2_X1 U40956 ( .A1(n54956), .A2(n54618), .Z(n19497) );
  NAND4_X2 U40957 ( .A1(n4690), .A2(n17487), .A3(n16058), .A4(n36038), .ZN(
        n20522) );
  NAND3_X1 U40979 ( .A1(n36549), .A2(n36384), .A3(n14763), .ZN(n60321) );
  OAI21_X2 U40980 ( .A1(n19550), .A2(n60767), .B(n60323), .ZN(n6407) );
  AOI21_X2 U40992 ( .A1(n19783), .A2(n29639), .B(n6408), .ZN(n60324) );
  AND2_X1 U40994 ( .A1(n36546), .A2(n60326), .Z(n60325) );
  AND2_X1 U40998 ( .A1(n36544), .A2(n36545), .Z(n60326) );
  BUF_X2 U40999 ( .I(n23955), .Z(n60327) );
  XOR2_X1 U41001 ( .A1(n60328), .A2(n586), .Z(n21241) );
  NAND3_X1 U41010 ( .A1(n43515), .A2(n43518), .A3(n43504), .ZN(n43180) );
  NOR2_X2 U41046 ( .A1(n1413), .A2(n21881), .ZN(n36866) );
  NOR2_X2 U41064 ( .A1(n3246), .A2(n3247), .ZN(n23492) );
  AOI21_X1 U41094 ( .A1(n14013), .A2(n14015), .B(n14018), .ZN(n14012) );
  NAND3_X1 U41095 ( .A1(n55604), .A2(n55619), .A3(n52295), .ZN(n52297) );
  OR2_X1 U41109 ( .A1(n50263), .A2(n4594), .Z(n48168) );
  XOR2_X1 U41122 ( .A1(n1094), .A2(n22305), .Z(n50559) );
  OR2_X1 U41129 ( .A1(n2608), .A2(n64562), .Z(n49128) );
  XOR2_X1 U41146 ( .A1(n21220), .A2(n60338), .Z(n21243) );
  XOR2_X1 U41150 ( .A1(n52550), .A2(n52456), .Z(n60338) );
  AOI21_X1 U41178 ( .A1(n42797), .A2(n42796), .B(n60862), .ZN(n42800) );
  NAND2_X2 U41185 ( .A1(n6059), .A2(n18511), .ZN(n22780) );
  NAND2_X1 U41196 ( .A1(n2562), .A2(n9852), .ZN(n34124) );
  NAND2_X1 U41198 ( .A1(n6758), .A2(n30277), .ZN(n60339) );
  XOR2_X1 U41199 ( .A1(n51391), .A2(n63021), .Z(n51397) );
  NOR2_X2 U41211 ( .A1(n36846), .A2(n36851), .ZN(n36841) );
  NOR2_X1 U41216 ( .A1(n47014), .A2(n60342), .ZN(n1084) );
  XOR2_X1 U41217 ( .A1(n51402), .A2(n60344), .Z(n52686) );
  XOR2_X1 U41224 ( .A1(n51400), .A2(n51399), .Z(n60344) );
  INV_X2 U41227 ( .I(n12028), .ZN(n16629) );
  NOR3_X1 U41239 ( .A1(n60858), .A2(n30638), .A3(n18691), .ZN(n30645) );
  XOR2_X1 U41246 ( .A1(n16969), .A2(n51919), .Z(n2265) );
  INV_X2 U41250 ( .I(n60345), .ZN(n863) );
  NAND3_X2 U41266 ( .A1(n57421), .A2(n21645), .A3(n60349), .ZN(n22939) );
  OAI22_X2 U41313 ( .A1(n25306), .A2(n40352), .B1(n61708), .B2(n6911), .ZN(
        n18869) );
  NOR2_X2 U41329 ( .A1(n23256), .A2(n64714), .ZN(n2455) );
  NAND3_X2 U41333 ( .A1(n28134), .A2(n28133), .A3(n28132), .ZN(n28143) );
  XOR2_X1 U41335 ( .A1(n2222), .A2(n56508), .Z(n52458) );
  XOR2_X1 U41355 ( .A1(n20554), .A2(n31442), .Z(n14961) );
  NOR2_X2 U41395 ( .A1(n56867), .A2(n56863), .ZN(n12454) );
  XOR2_X1 U41429 ( .A1(n13289), .A2(n13290), .Z(n10065) );
  XOR2_X1 U41445 ( .A1(n51478), .A2(n51593), .Z(n23273) );
  INV_X1 U41447 ( .I(n60362), .ZN(n60361) );
  AOI21_X1 U41450 ( .A1(n40601), .A2(n42156), .B(n42585), .ZN(n60362) );
  NOR3_X2 U41459 ( .A1(n5133), .A2(n34619), .A3(n896), .ZN(n60364) );
  XOR2_X1 U41460 ( .A1(n60365), .A2(n60366), .Z(n3890) );
  XOR2_X1 U41465 ( .A1(n60367), .A2(n10663), .Z(n6810) );
  XOR2_X1 U41472 ( .A1(n17907), .A2(n19656), .Z(n60367) );
  NOR3_X2 U41477 ( .A1(n22680), .A2(n22679), .A3(n15942), .ZN(n16655) );
  XOR2_X1 U41479 ( .A1(n51158), .A2(n4252), .Z(n50034) );
  NOR2_X2 U41482 ( .A1(n20209), .A2(n60368), .ZN(n10160) );
  NOR2_X2 U41485 ( .A1(n43779), .A2(n12091), .ZN(n60368) );
  NAND2_X2 U41500 ( .A1(n34149), .A2(n32846), .ZN(n6033) );
  XOR2_X1 U41501 ( .A1(n4289), .A2(n38090), .Z(n22515) );
  NOR2_X2 U41508 ( .A1(n14019), .A2(n28607), .ZN(n18213) );
  XOR2_X1 U41510 ( .A1(n60380), .A2(n33908), .Z(n33911) );
  XOR2_X1 U41511 ( .A1(n33909), .A2(n33907), .Z(n60380) );
  OAI21_X2 U41513 ( .A1(n5171), .A2(n43086), .B(n43085), .ZN(n14263) );
  NOR3_X2 U41514 ( .A1(n24981), .A2(n10203), .A3(n24250), .ZN(n5171) );
  XOR2_X1 U41515 ( .A1(n60381), .A2(n20409), .Z(n24447) );
  XOR2_X1 U41523 ( .A1(n32725), .A2(n32573), .Z(n60382) );
  XOR2_X1 U41539 ( .A1(n60383), .A2(n3113), .Z(n23114) );
  BUF_X2 U41549 ( .I(n5090), .Z(n60386) );
  NOR2_X2 U41565 ( .A1(n13144), .A2(n30408), .ZN(n30415) );
  NAND2_X1 U41574 ( .A1(n15397), .A2(n41904), .ZN(n60522) );
  NAND2_X2 U41581 ( .A1(n60393), .A2(n24422), .ZN(n56886) );
  XOR2_X1 U41591 ( .A1(n6566), .A2(n60395), .Z(n60394) );
  XOR2_X1 U41593 ( .A1(n33828), .A2(n33829), .Z(n33835) );
  NOR2_X1 U41597 ( .A1(n21972), .A2(n64076), .ZN(n60400) );
  OR2_X1 U41616 ( .A1(n32212), .A2(n22176), .Z(n60404) );
  XOR2_X1 U41618 ( .A1(n11442), .A2(n11488), .Z(n11487) );
  XOR2_X1 U41626 ( .A1(n52157), .A2(n25158), .Z(n11488) );
  INV_X2 U41627 ( .I(n60405), .ZN(n14038) );
  NAND3_X2 U41637 ( .A1(n60408), .A2(n61644), .A3(n60407), .ZN(n342) );
  XOR2_X1 U41638 ( .A1(n60409), .A2(n14793), .Z(n15429) );
  XOR2_X1 U41642 ( .A1(n6975), .A2(n14794), .Z(n60409) );
  AOI21_X2 U41644 ( .A1(n60411), .A2(n60410), .B(n59269), .ZN(n22547) );
  NAND2_X1 U41648 ( .A1(n16772), .A2(n57407), .ZN(n14326) );
  NAND2_X1 U41654 ( .A1(n14729), .A2(n30271), .ZN(n30719) );
  XOR2_X1 U41658 ( .A1(n19441), .A2(n9362), .Z(n37721) );
  INV_X2 U41664 ( .I(n3310), .ZN(n28796) );
  XOR2_X1 U41665 ( .A1(n3310), .A2(n12591), .Z(n32377) );
  NOR2_X2 U41666 ( .A1(n2668), .A2(n2667), .ZN(n3310) );
  BUF_X2 U41667 ( .I(n19005), .Z(n60416) );
  INV_X2 U41682 ( .I(n13836), .ZN(n60417) );
  NAND2_X2 U41685 ( .A1(n17967), .A2(n60417), .ZN(n47669) );
  INV_X2 U41694 ( .I(n60420), .ZN(n38338) );
  XNOR2_X1 U41699 ( .A1(n22060), .A2(n5039), .ZN(n60420) );
  NAND2_X2 U41700 ( .A1(n34459), .A2(n57416), .ZN(n38806) );
  NAND2_X2 U41730 ( .A1(n20559), .A2(n60425), .ZN(n53736) );
  INV_X1 U41751 ( .I(n45571), .ZN(n60429) );
  BUF_X2 U41753 ( .I(n37224), .Z(n60431) );
  XOR2_X1 U41757 ( .A1(n2998), .A2(n58831), .Z(n20044) );
  NOR3_X2 U41758 ( .A1(n24411), .A2(n10206), .A3(n15958), .ZN(n28677) );
  NOR2_X1 U41763 ( .A1(n6442), .A2(n54476), .ZN(n54477) );
  NAND2_X1 U41773 ( .A1(n11145), .A2(n60435), .ZN(n11920) );
  NAND2_X1 U41783 ( .A1(n56336), .A2(n61727), .ZN(n60435) );
  XOR2_X1 U41791 ( .A1(n37735), .A2(n8205), .Z(n8204) );
  XOR2_X1 U41798 ( .A1(n44154), .A2(n60350), .Z(n45320) );
  XOR2_X1 U41800 ( .A1(n19407), .A2(n62548), .Z(n32595) );
  NAND3_X2 U41811 ( .A1(n3814), .A2(n3813), .A3(n30454), .ZN(n29069) );
  NAND4_X2 U41818 ( .A1(n43756), .A2(n60444), .A3(n43753), .A4(n43754), .ZN(
        n44004) );
  AOI22_X1 U41819 ( .A1(n46737), .A2(n43749), .B1(n11821), .B2(n18980), .ZN(
        n60444) );
  NOR2_X1 U41835 ( .A1(n17799), .A2(n55225), .ZN(n2531) );
  INV_X2 U41839 ( .I(n12944), .ZN(n56403) );
  XOR2_X1 U41842 ( .A1(n12945), .A2(n19224), .Z(n12944) );
  AND2_X2 U41849 ( .A1(n24748), .A2(n3039), .Z(n2524) );
  XOR2_X1 U41867 ( .A1(n60717), .A2(n31795), .Z(n881) );
  XOR2_X1 U41871 ( .A1(n13457), .A2(n60449), .Z(n13456) );
  XOR2_X1 U41874 ( .A1(n39289), .A2(n39288), .Z(n60449) );
  NAND2_X2 U41888 ( .A1(n48648), .A2(n23416), .ZN(n48513) );
  NOR2_X2 U41893 ( .A1(n2548), .A2(n2546), .ZN(n60450) );
  NAND3_X2 U41900 ( .A1(n27995), .A2(n60451), .A3(n15898), .ZN(n15105) );
  AOI21_X2 U41903 ( .A1(n54686), .A2(n54650), .B(n54684), .ZN(n18463) );
  NAND2_X2 U41904 ( .A1(n54842), .A2(n54649), .ZN(n54684) );
  NAND2_X2 U41907 ( .A1(n34980), .A2(n23834), .ZN(n34069) );
  XOR2_X1 U41945 ( .A1(n60453), .A2(n2677), .Z(n10319) );
  AOI21_X1 U41948 ( .A1(n15359), .A2(n7541), .B(n22468), .ZN(n8643) );
  NAND2_X2 U41968 ( .A1(n8800), .A2(n22278), .ZN(n35300) );
  XOR2_X1 U41976 ( .A1(n60455), .A2(n11149), .Z(n23278) );
  XOR2_X1 U41979 ( .A1(n8416), .A2(n32037), .Z(n25388) );
  INV_X2 U41992 ( .I(n60459), .ZN(n12477) );
  XOR2_X1 U41995 ( .A1(Ciphertext[136]), .A2(Key[173]), .Z(n60459) );
  AND2_X1 U42028 ( .A1(n13144), .A2(n28711), .Z(n21678) );
  XOR2_X1 U42029 ( .A1(n44161), .A2(n44160), .Z(n7203) );
  AND2_X1 U42030 ( .A1(n36567), .A2(n23215), .Z(n3809) );
  INV_X1 U42032 ( .I(n29058), .ZN(n60508) );
  NAND2_X2 U42041 ( .A1(n15747), .A2(n52768), .ZN(n53572) );
  NOR2_X2 U42056 ( .A1(n1402), .A2(n15731), .ZN(n24477) );
  OR2_X1 U42076 ( .A1(n61563), .A2(n64063), .Z(n60465) );
  OR2_X1 U42091 ( .A1(n4115), .A2(n31841), .Z(n6124) );
  XOR2_X1 U42119 ( .A1(n60466), .A2(n24023), .Z(n61365) );
  NAND2_X2 U42124 ( .A1(n2442), .A2(n2436), .ZN(n24023) );
  XOR2_X1 U42125 ( .A1(n6092), .A2(n7998), .Z(n37876) );
  NOR2_X1 U42137 ( .A1(n56843), .A2(n56842), .ZN(n17654) );
  NAND3_X2 U42142 ( .A1(n56867), .A2(n56885), .A3(n56892), .ZN(n56842) );
  XOR2_X1 U42145 ( .A1(n11846), .A2(n11845), .Z(n13082) );
  XNOR2_X1 U42148 ( .A1(n3840), .A2(n3841), .ZN(n33467) );
  NAND2_X1 U42150 ( .A1(n28074), .A2(n28075), .ZN(n4602) );
  NAND2_X2 U42152 ( .A1(n36469), .A2(n36470), .ZN(n22254) );
  NOR3_X2 U42153 ( .A1(n60470), .A2(n26130), .A3(n60469), .ZN(n1020) );
  NAND2_X1 U42166 ( .A1(n39815), .A2(n39816), .ZN(n60469) );
  INV_X1 U42167 ( .I(n13016), .ZN(n21365) );
  XOR2_X1 U42168 ( .A1(n13016), .A2(n57323), .Z(n61441) );
  OR2_X1 U42171 ( .A1(n60413), .A2(n60960), .Z(n33463) );
  AOI21_X1 U42179 ( .A1(n21158), .A2(n28072), .B(n60473), .ZN(n15829) );
  NOR2_X2 U42186 ( .A1(n3376), .A2(n25213), .ZN(n61168) );
  XOR2_X1 U42188 ( .A1(n63024), .A2(n17085), .Z(n50036) );
  NOR2_X2 U42189 ( .A1(n16868), .A2(n17089), .ZN(n17085) );
  NAND2_X2 U42193 ( .A1(n8309), .A2(n8308), .ZN(n33010) );
  NOR2_X1 U42195 ( .A1(n53054), .A2(n53094), .ZN(n53113) );
  NOR2_X1 U42200 ( .A1(n20389), .A2(n30628), .ZN(n20388) );
  NAND4_X2 U42209 ( .A1(n25016), .A2(n60479), .A3(n25014), .A4(n23973), .ZN(
        n23972) );
  NAND2_X1 U42215 ( .A1(n60480), .A2(n21582), .ZN(n6950) );
  OAI21_X1 U42217 ( .A1(n25198), .A2(n6952), .B(n15434), .ZN(n60480) );
  XOR2_X1 U42232 ( .A1(n60482), .A2(n50658), .Z(n25948) );
  NOR2_X2 U42233 ( .A1(n19118), .A2(n6316), .ZN(n7596) );
  INV_X2 U42239 ( .I(n25855), .ZN(n48625) );
  NAND2_X1 U42246 ( .A1(n50254), .A2(n50342), .ZN(n13683) );
  XOR2_X1 U42247 ( .A1(n15560), .A2(n15561), .Z(n45237) );
  NOR2_X1 U42259 ( .A1(n261), .A2(n54984), .ZN(n60488) );
  XOR2_X1 U42262 ( .A1(n24653), .A2(n60490), .Z(n13538) );
  XOR2_X1 U42271 ( .A1(n21027), .A2(n12518), .Z(n60490) );
  XOR2_X1 U42273 ( .A1(n13552), .A2(n14081), .Z(n14080) );
  NAND4_X2 U42278 ( .A1(n38680), .A2(n60493), .A3(n2090), .A4(n40631), .ZN(
        n2087) );
  OR2_X1 U42290 ( .A1(n42916), .A2(n42914), .Z(n10617) );
  NAND3_X2 U42294 ( .A1(n53446), .A2(n13401), .A3(n60494), .ZN(n10027) );
  XOR2_X1 U42314 ( .A1(n60495), .A2(n53076), .Z(Plaintext[2]) );
  INV_X2 U42337 ( .I(n60496), .ZN(n1164) );
  NAND2_X2 U42339 ( .A1(n9338), .A2(n1232), .ZN(n60496) );
  XOR2_X1 U42351 ( .A1(n52322), .A2(n63031), .Z(n60497) );
  BUF_X2 U42362 ( .I(n38648), .Z(n60499) );
  INV_X2 U42370 ( .I(n42225), .ZN(n3090) );
  NAND2_X2 U42371 ( .A1(n24989), .A2(n28244), .ZN(n60505) );
  INV_X2 U42373 ( .I(n2023), .ZN(n31993) );
  XOR2_X1 U42381 ( .A1(n2023), .A2(n60500), .Z(n25364) );
  INV_X4 U42385 ( .I(n61503), .ZN(n25698) );
  OAI21_X1 U42388 ( .A1(n41002), .A2(n61308), .B(n41001), .ZN(n60501) );
  BUF_X2 U42391 ( .I(n24343), .Z(n60502) );
  NOR2_X2 U42395 ( .A1(n1787), .A2(n36026), .ZN(n34821) );
  NAND3_X2 U42398 ( .A1(n16549), .A2(n16548), .A3(n16550), .ZN(n12478) );
  AOI21_X1 U42399 ( .A1(n42482), .A2(n42481), .B(n18242), .ZN(n60503) );
  NOR3_X2 U42412 ( .A1(n60508), .A2(n883), .A3(n61391), .ZN(n2143) );
  INV_X1 U42429 ( .I(n60735), .ZN(n60734) );
  OR3_X1 U42436 ( .A1(n30391), .A2(n5242), .A3(n4037), .Z(n4063) );
  XOR2_X1 U42441 ( .A1(n18133), .A2(n44384), .Z(n60511) );
  INV_X2 U42446 ( .I(n60513), .ZN(n42225) );
  XNOR2_X1 U42456 ( .A1(n5783), .A2(n5780), .ZN(n60513) );
  NAND3_X2 U42462 ( .A1(n13671), .A2(n54904), .A3(n22486), .ZN(n61529) );
  XOR2_X1 U42469 ( .A1(n7388), .A2(n6336), .Z(n19703) );
  XOR2_X1 U42472 ( .A1(n46165), .A2(n43370), .Z(n44129) );
  NAND3_X1 U42473 ( .A1(n53450), .A2(n1605), .A3(n53587), .ZN(n53454) );
  NOR2_X2 U42477 ( .A1(n7021), .A2(n53462), .ZN(n53507) );
  XOR2_X1 U42496 ( .A1(n49804), .A2(n47947), .Z(n60515) );
  OR2_X1 U42505 ( .A1(n27276), .A2(n27277), .Z(n60518) );
  AOI21_X2 U42506 ( .A1(n60519), .A2(n41350), .B(n5849), .ZN(n5848) );
  NAND2_X1 U42517 ( .A1(n50424), .A2(n50425), .ZN(n50431) );
  NAND3_X1 U42521 ( .A1(n57201), .A2(n54727), .A3(n54769), .ZN(n7307) );
  NAND2_X2 U42544 ( .A1(n36477), .A2(n4893), .ZN(n36152) );
  NAND3_X2 U42551 ( .A1(n4361), .A2(n26572), .A3(n26571), .ZN(n60523) );
  NAND2_X2 U42557 ( .A1(n24451), .A2(n60526), .ZN(n51035) );
  NOR2_X2 U42571 ( .A1(n4322), .A2(n57974), .ZN(n42735) );
  NAND2_X1 U42574 ( .A1(n46177), .A2(n48176), .ZN(n60687) );
  AND2_X1 U42580 ( .A1(n5594), .A2(n24504), .Z(n60529) );
  XOR2_X1 U42591 ( .A1(n52371), .A2(n52064), .Z(n60531) );
  XOR2_X1 U42607 ( .A1(n60534), .A2(n769), .Z(n15544) );
  XOR2_X1 U42608 ( .A1(n6505), .A2(n33230), .Z(n60534) );
  NAND3_X1 U42641 ( .A1(n16635), .A2(n35544), .A3(n16634), .ZN(n16633) );
  NAND2_X2 U42662 ( .A1(n49207), .A2(n60538), .ZN(n17173) );
  NAND4_X2 U42664 ( .A1(n33707), .A2(n33708), .A3(n33705), .A4(n33706), .ZN(
        n33709) );
  OR2_X1 U42678 ( .A1(n19887), .A2(n21019), .Z(n26914) );
  NOR2_X2 U42680 ( .A1(n60542), .A2(n60540), .ZN(n26897) );
  NAND2_X2 U42682 ( .A1(n26074), .A2(n60541), .ZN(n60540) );
  INV_X2 U42683 ( .I(n27668), .ZN(n60541) );
  NAND3_X2 U42691 ( .A1(n60544), .A2(n19933), .A3(n44134), .ZN(n19932) );
  BUF_X2 U42693 ( .I(n27665), .Z(n60545) );
  XOR2_X1 U42700 ( .A1(n1548), .A2(n20212), .Z(n11169) );
  INV_X1 U42717 ( .I(n60550), .ZN(n52134) );
  OAI21_X1 U42721 ( .A1(n3567), .A2(n60552), .B(n60551), .ZN(n60550) );
  NAND2_X1 U42727 ( .A1(n14142), .A2(n62991), .ZN(n60551) );
  XOR2_X1 U42730 ( .A1(n4692), .A2(n5155), .Z(n60555) );
  BUF_X2 U42744 ( .I(n53477), .Z(n60556) );
  INV_X2 U42752 ( .I(n60557), .ZN(n45673) );
  OR3_X1 U42766 ( .A1(n12300), .A2(n5688), .A3(n463), .Z(n26708) );
  XOR2_X1 U42772 ( .A1(n14447), .A2(n19335), .Z(n60561) );
  NOR2_X2 U42785 ( .A1(n24402), .A2(n5070), .ZN(n5179) );
  XOR2_X1 U42788 ( .A1(n32734), .A2(n32068), .Z(n4056) );
  XOR2_X1 U42794 ( .A1(n31194), .A2(n31193), .Z(n32734) );
  NOR2_X2 U42807 ( .A1(n40728), .A2(n16102), .ZN(n61407) );
  OAI21_X2 U42811 ( .A1(n14723), .A2(n14722), .B(n31791), .ZN(n38591) );
  XOR2_X1 U42815 ( .A1(n24731), .A2(n45136), .Z(n60568) );
  XOR2_X1 U42818 ( .A1(n45813), .A2(n46609), .Z(n60570) );
  XOR2_X1 U42828 ( .A1(n60571), .A2(n10724), .Z(n10727) );
  XOR2_X1 U42832 ( .A1(n50851), .A2(n17941), .Z(n60571) );
  NAND3_X2 U42836 ( .A1(n50337), .A2(n21476), .A3(n21352), .ZN(n11503) );
  INV_X1 U42837 ( .I(n36699), .ZN(n623) );
  NAND2_X1 U42839 ( .A1(n1252), .A2(n39175), .ZN(n42004) );
  XOR2_X1 U42848 ( .A1(n60572), .A2(n45385), .Z(n10202) );
  NOR2_X2 U42852 ( .A1(n45412), .A2(n4090), .ZN(n47140) );
  NAND2_X2 U42857 ( .A1(n45437), .A2(n20902), .ZN(n4090) );
  NOR2_X1 U42862 ( .A1(n25107), .A2(n60573), .ZN(n12133) );
  NOR2_X2 U42865 ( .A1(n20025), .A2(n29727), .ZN(n29879) );
  OR2_X1 U42893 ( .A1(n20034), .A2(n29628), .Z(n28823) );
  NAND2_X1 U42894 ( .A1(n43577), .A2(n59746), .ZN(n41965) );
  XOR2_X1 U42923 ( .A1(n24178), .A2(n60580), .Z(n8463) );
  INV_X2 U42927 ( .I(n60581), .ZN(n38600) );
  XOR2_X1 U42930 ( .A1(n24480), .A2(n60582), .Z(n24479) );
  XOR2_X1 U42931 ( .A1(n50853), .A2(n50941), .Z(n60582) );
  NAND2_X2 U42933 ( .A1(n47208), .A2(n48460), .ZN(n3111) );
  XOR2_X1 U42939 ( .A1(n39750), .A2(n60584), .Z(n3437) );
  XOR2_X1 U42940 ( .A1(n3440), .A2(n37900), .Z(n60584) );
  OAI22_X1 U42941 ( .A1(n14139), .A2(n60585), .B1(n8489), .B2(n14141), .ZN(
        n24957) );
  NAND2_X1 U42943 ( .A1(n1600), .A2(n55975), .ZN(n60585) );
  XNOR2_X1 U42947 ( .A1(n13190), .A2(n16049), .ZN(n60587) );
  XOR2_X1 U42986 ( .A1(n51997), .A2(n9632), .Z(n50869) );
  AOI21_X2 U42990 ( .A1(n7333), .A2(n56209), .B(n22382), .ZN(n25411) );
  NOR3_X1 U42998 ( .A1(n61089), .A2(n49547), .A3(n24394), .ZN(n13631) );
  XOR2_X1 U42999 ( .A1(n38621), .A2(n60594), .Z(n8543) );
  XOR2_X1 U43002 ( .A1(n38623), .A2(n15957), .Z(n60594) );
  OAI21_X1 U43009 ( .A1(n60595), .A2(n17897), .B(n902), .ZN(n34031) );
  XOR2_X1 U43029 ( .A1(n39586), .A2(n37698), .Z(n5785) );
  XOR2_X1 U43030 ( .A1(n39670), .A2(n20667), .Z(n39586) );
  XOR2_X1 U43038 ( .A1(n2823), .A2(n37708), .Z(n37709) );
  NOR2_X2 U43039 ( .A1(n28128), .A2(n23578), .ZN(n28137) );
  NAND2_X1 U43041 ( .A1(n16335), .A2(n49989), .ZN(n16334) );
  XOR2_X1 U43075 ( .A1(n60599), .A2(n16843), .Z(n32529) );
  XOR2_X1 U43080 ( .A1(n4949), .A2(n32510), .Z(n60599) );
  NAND3_X2 U43096 ( .A1(n9817), .A2(n9816), .A3(n60600), .ZN(n23839) );
  OAI21_X2 U43097 ( .A1(n19801), .A2(n47140), .B(n47143), .ZN(n60600) );
  INV_X2 U43104 ( .I(n60602), .ZN(n976) );
  NAND2_X2 U43110 ( .A1(n12034), .A2(n1705), .ZN(n41496) );
  NOR2_X2 U43113 ( .A1(n40063), .A2(n42441), .ZN(n40314) );
  NOR2_X2 U43115 ( .A1(n48251), .A2(n48504), .ZN(n48494) );
  NAND2_X2 U43116 ( .A1(n7854), .A2(n48521), .ZN(n48251) );
  NOR3_X2 U43129 ( .A1(n5204), .A2(n1065), .A3(n48491), .ZN(n5203) );
  NOR2_X1 U43138 ( .A1(n29189), .A2(n27273), .ZN(n27277) );
  INV_X4 U43139 ( .I(n24298), .ZN(n1277) );
  NAND2_X2 U43150 ( .A1(n25940), .A2(n25939), .ZN(n24298) );
  NAND2_X2 U43159 ( .A1(n41924), .A2(n42252), .ZN(n37895) );
  XOR2_X1 U43163 ( .A1(n8620), .A2(n46434), .Z(n60610) );
  NAND2_X2 U43170 ( .A1(n40028), .A2(n23904), .ZN(n6153) );
  XOR2_X1 U43179 ( .A1(n26181), .A2(n44908), .Z(n20717) );
  XOR2_X1 U43196 ( .A1(n61352), .A2(n51097), .Z(n51104) );
  OR2_X1 U43198 ( .A1(n29417), .A2(n30437), .Z(n60615) );
  XOR2_X1 U43220 ( .A1(n65144), .A2(n60617), .Z(n27) );
  XOR2_X1 U43221 ( .A1(n44238), .A2(n43811), .Z(n60617) );
  NOR2_X1 U43226 ( .A1(n42607), .A2(n42594), .ZN(n37534) );
  NOR2_X1 U43230 ( .A1(n11505), .A2(n39985), .ZN(n39986) );
  NAND2_X2 U43232 ( .A1(n19539), .A2(n36233), .ZN(n36234) );
  NOR2_X2 U43234 ( .A1(n52477), .A2(n52476), .ZN(n21248) );
  NOR2_X2 U43252 ( .A1(n10379), .A2(n57393), .ZN(n61433) );
  INV_X1 U43257 ( .I(n60619), .ZN(n13094) );
  NAND2_X2 U43275 ( .A1(n14709), .A2(n60961), .ZN(n52287) );
  XOR2_X1 U43287 ( .A1(n13089), .A2(n4953), .Z(n31982) );
  NAND4_X1 U43294 ( .A1(n46862), .A2(n45713), .A3(n62571), .A4(n45714), .ZN(
        n45722) );
  NAND2_X2 U43296 ( .A1(n21829), .A2(n21570), .ZN(n9953) );
  OR3_X1 U43297 ( .A1(n47970), .A2(n19681), .A3(n19589), .Z(n19900) );
  XOR2_X1 U43306 ( .A1(n60624), .A2(n31962), .Z(n21825) );
  XOR2_X1 U43310 ( .A1(n21944), .A2(n33158), .Z(n60624) );
  OAI21_X2 U43315 ( .A1(n60105), .A2(n11571), .B(n6350), .ZN(n53183) );
  OR2_X1 U43319 ( .A1(n30429), .A2(n31083), .Z(n60625) );
  BUF_X2 U43321 ( .I(n1547), .Z(n60628) );
  AOI21_X2 U43322 ( .A1(n7555), .A2(n57231), .B(n60629), .ZN(n54874) );
  NOR2_X2 U43337 ( .A1(n52476), .A2(n21169), .ZN(n60630) );
  NAND2_X2 U43341 ( .A1(n7130), .A2(n30552), .ZN(n24503) );
  NOR2_X1 U43353 ( .A1(n45763), .A2(n60632), .ZN(n60631) );
  XOR2_X1 U43358 ( .A1(n20469), .A2(n32618), .Z(n60661) );
  NAND2_X2 U43359 ( .A1(n61939), .A2(n19587), .ZN(n20469) );
  XOR2_X1 U43360 ( .A1(n54708), .A2(n55191), .Z(n30602) );
  XOR2_X1 U43362 ( .A1(n3229), .A2(n60634), .Z(n20528) );
  XOR2_X1 U43367 ( .A1(n39660), .A2(n38263), .Z(n60634) );
  XOR2_X1 U43369 ( .A1(n9166), .A2(n60635), .Z(n26134) );
  XOR2_X1 U43381 ( .A1(n42625), .A2(n46239), .Z(n60635) );
  NAND3_X2 U43395 ( .A1(n36881), .A2(n36880), .A3(n36879), .ZN(n3480) );
  NAND3_X2 U43397 ( .A1(n26999), .A2(n26998), .A3(n26997), .ZN(n20771) );
  BUF_X4 U43425 ( .I(n21055), .Z(n4723) );
  INV_X2 U43434 ( .I(n36883), .ZN(n60639) );
  NOR2_X2 U43437 ( .A1(n7074), .A2(n12798), .ZN(n36883) );
  XOR2_X1 U43439 ( .A1(n1994), .A2(n14443), .Z(n1993) );
  AND3_X1 U43444 ( .A1(n38043), .A2(n38042), .A3(n40149), .Z(n7474) );
  NOR2_X2 U43445 ( .A1(n5129), .A2(n20653), .ZN(n55906) );
  OR2_X1 U43448 ( .A1(n30561), .A2(n30562), .Z(n25030) );
  INV_X2 U43464 ( .I(n60641), .ZN(n17632) );
  XOR2_X1 U43470 ( .A1(Ciphertext[151]), .A2(Key[182]), .Z(n60641) );
  AND2_X1 U43475 ( .A1(n60894), .A2(n57289), .Z(n60890) );
  NOR2_X1 U43484 ( .A1(n60643), .A2(n11876), .ZN(n10661) );
  NAND3_X1 U43485 ( .A1(n270), .A2(n24238), .A3(n31251), .ZN(n60643) );
  NAND4_X1 U43486 ( .A1(n56921), .A2(n52289), .A3(n52288), .A4(n56919), .ZN(
        n60644) );
  NAND2_X2 U43493 ( .A1(n56719), .A2(n56733), .ZN(n56707) );
  NOR2_X1 U43527 ( .A1(n45581), .A2(n45580), .ZN(n45582) );
  NOR2_X2 U43531 ( .A1(n42662), .A2(n21377), .ZN(n40547) );
  NAND2_X2 U43532 ( .A1(n48838), .A2(n48286), .ZN(n49516) );
  NOR2_X2 U43535 ( .A1(n3694), .A2(n15709), .ZN(n48838) );
  NAND2_X2 U43536 ( .A1(n12850), .A2(n60645), .ZN(n1064) );
  NOR2_X2 U43541 ( .A1(n21044), .A2(n47501), .ZN(n60645) );
  OR2_X2 U43546 ( .A1(n15524), .A2(n24697), .Z(n22468) );
  AOI22_X1 U43548 ( .A1(n45193), .A2(n18000), .B1(n45195), .B2(n17317), .ZN(
        n17316) );
  INV_X1 U43554 ( .I(n60502), .ZN(n19927) );
  XOR2_X1 U43557 ( .A1(n60649), .A2(n19713), .Z(n14187) );
  NAND2_X1 U43571 ( .A1(n42105), .A2(n42555), .ZN(n61194) );
  NAND3_X1 U43573 ( .A1(n20709), .A2(n25091), .A3(n49050), .ZN(n49051) );
  XOR2_X1 U43575 ( .A1(n44369), .A2(n44370), .Z(n60650) );
  NAND2_X2 U43580 ( .A1(n19701), .A2(n58273), .ZN(n8211) );
  XOR2_X1 U43593 ( .A1(n31913), .A2(n60654), .Z(n879) );
  XOR2_X1 U43594 ( .A1(n60655), .A2(n51832), .Z(n8143) );
  INV_X2 U43603 ( .I(n52424), .ZN(n60655) );
  NAND3_X2 U43604 ( .A1(n22488), .A2(n48724), .A3(n48723), .ZN(n51832) );
  XOR2_X1 U43639 ( .A1(n46408), .A2(n45821), .Z(n60656) );
  BUF_X4 U43642 ( .I(n3932), .Z(n61177) );
  OAI22_X2 U43652 ( .A1(n6137), .A2(n28031), .B1(n7775), .B2(n6215), .ZN(
        n28234) );
  AOI22_X1 U43674 ( .A1(n18145), .A2(n55006), .B1(n55310), .B2(n14927), .ZN(
        n21392) );
  NAND4_X2 U43684 ( .A1(n9700), .A2(n55071), .A3(n83), .A4(n55070), .ZN(n61602) );
  INV_X2 U43701 ( .I(n60662), .ZN(n815) );
  XOR2_X1 U43706 ( .A1(Ciphertext[133]), .A2(Key[56]), .Z(n60662) );
  NAND3_X1 U43711 ( .A1(n41899), .A2(n41901), .A3(n41900), .ZN(n41902) );
  NOR2_X1 U43713 ( .A1(n60663), .A2(n56721), .ZN(n56728) );
  AOI22_X1 U43717 ( .A1(n56718), .A2(n23785), .B1(n56731), .B2(n56719), .ZN(
        n60663) );
  INV_X2 U43718 ( .I(n9289), .ZN(n4880) );
  NOR3_X2 U43721 ( .A1(n6542), .A2(n6541), .A3(n35262), .ZN(n37397) );
  NAND3_X2 U43722 ( .A1(n40952), .A2(n23986), .A3(n40199), .ZN(n40207) );
  NOR2_X2 U43738 ( .A1(n1546), .A2(n16402), .ZN(n35316) );
  INV_X2 U43747 ( .I(n60668), .ZN(n61662) );
  XOR2_X1 U43750 ( .A1(n62646), .A2(n13313), .Z(n60668) );
  INV_X2 U43752 ( .I(n60670), .ZN(n3697) );
  XOR2_X1 U43768 ( .A1(Ciphertext[60]), .A2(Key[25]), .Z(n60670) );
  NAND2_X2 U43777 ( .A1(n5584), .A2(n5400), .ZN(n23017) );
  NAND2_X2 U43778 ( .A1(n63549), .A2(n19278), .ZN(n17144) );
  NAND2_X2 U43783 ( .A1(n54058), .A2(n54035), .ZN(n53557) );
  NAND2_X1 U43791 ( .A1(n18250), .A2(n10768), .ZN(n60674) );
  NAND2_X1 U43792 ( .A1(n17638), .A2(n60675), .ZN(Plaintext[47]) );
  NAND4_X1 U43795 ( .A1(n17637), .A2(n17055), .A3(n17644), .A4(n17056), .ZN(
        n60675) );
  OR2_X1 U43806 ( .A1(n30666), .A2(n60676), .Z(n6406) );
  OAI22_X1 U43807 ( .A1(n30313), .A2(n25052), .B1(n30314), .B2(n30758), .ZN(
        n60676) );
  XOR2_X1 U43814 ( .A1(n25524), .A2(n60677), .Z(n33005) );
  XOR2_X1 U43818 ( .A1(n33233), .A2(n31628), .Z(n60677) );
  XOR2_X1 U43826 ( .A1(n46228), .A2(n11878), .Z(n269) );
  NAND2_X2 U43830 ( .A1(n5525), .A2(n5523), .ZN(n39230) );
  XOR2_X1 U43842 ( .A1(n31412), .A2(n31413), .Z(n60682) );
  NOR2_X1 U43847 ( .A1(n16633), .A2(n60691), .ZN(n16637) );
  OR2_X1 U43849 ( .A1(n33989), .A2(n60684), .Z(n60683) );
  NAND2_X1 U43861 ( .A1(n10924), .A2(n30666), .ZN(n60750) );
  NAND2_X1 U43864 ( .A1(n22491), .A2(n60688), .ZN(n54715) );
  NAND3_X2 U43880 ( .A1(n12273), .A2(n12277), .A3(n16425), .ZN(n19225) );
  XOR2_X1 U43896 ( .A1(n60692), .A2(n27013), .Z(n28003) );
  XOR2_X1 U43909 ( .A1(n37864), .A2(n13634), .Z(n5640) );
  NAND3_X1 U43911 ( .A1(n8602), .A2(n2310), .A3(n2636), .ZN(n884) );
  NOR3_X2 U43939 ( .A1(n60762), .A2(n60761), .A3(n8744), .ZN(n1958) );
  XOR2_X1 U43943 ( .A1(n383), .A2(n9007), .Z(n60699) );
  NOR2_X1 U43946 ( .A1(n11836), .A2(n1414), .ZN(n61246) );
  XOR2_X1 U44019 ( .A1(n60702), .A2(n20948), .Z(n39730) );
  XOR2_X1 U44046 ( .A1(n38711), .A2(n39618), .Z(n60702) );
  XOR2_X1 U44078 ( .A1(n25364), .A2(n9698), .Z(n31442) );
  XOR2_X1 U44089 ( .A1(n60707), .A2(n1620), .Z(n25351) );
  XOR2_X1 U44114 ( .A1(n50531), .A2(n50532), .Z(n60707) );
  BUF_X2 U44139 ( .I(n20552), .Z(n60709) );
  XOR2_X1 U44192 ( .A1(n31902), .A2(n2612), .Z(n3578) );
  XOR2_X1 U44239 ( .A1(n21009), .A2(n38728), .Z(n60711) );
  XOR2_X1 U44326 ( .A1(n2637), .A2(n18711), .Z(n60713) );
  XOR2_X1 U44371 ( .A1(n60720), .A2(n25075), .Z(n18518) );
  XOR2_X1 U44373 ( .A1(n36505), .A2(n16346), .Z(n60720) );
  NAND2_X1 U44379 ( .A1(n1593), .A2(n55132), .ZN(n55163) );
  NAND2_X1 U44382 ( .A1(n25724), .A2(n60721), .ZN(n25725) );
  NAND2_X1 U44383 ( .A1(n55138), .A2(n55137), .ZN(n60721) );
  AOI21_X1 U44403 ( .A1(n52642), .A2(n60723), .B(n60722), .ZN(n26119) );
  NAND3_X1 U44408 ( .A1(n52640), .A2(n52639), .A3(n54849), .ZN(n60722) );
  OR2_X1 U44414 ( .A1(n52643), .A2(n54852), .Z(n60723) );
  NOR2_X2 U44454 ( .A1(n20461), .A2(n23532), .ZN(n21269) );
  NAND2_X2 U44455 ( .A1(n25001), .A2(n25003), .ZN(n23532) );
  NAND3_X2 U44466 ( .A1(n2236), .A2(n1061), .A3(n2235), .ZN(n44385) );
  NOR2_X2 U44468 ( .A1(n60728), .A2(n28380), .ZN(n27555) );
  XOR2_X1 U44484 ( .A1(n7627), .A2(n32398), .Z(n60731) );
  OAI21_X1 U44494 ( .A1(n49833), .A2(n11950), .B(n49069), .ZN(n60735) );
  XOR2_X1 U44574 ( .A1(n50923), .A2(n20578), .Z(n60736) );
  NAND3_X2 U44576 ( .A1(n10887), .A2(n28820), .A3(n60737), .ZN(n31221) );
  NOR2_X1 U44578 ( .A1(n17462), .A2(n28807), .ZN(n60737) );
  NOR2_X2 U44596 ( .A1(n29501), .A2(n3993), .ZN(n30398) );
  XOR2_X1 U44635 ( .A1(n46509), .A2(n46508), .Z(n60740) );
  AOI22_X1 U44650 ( .A1(n60741), .A2(n21690), .B1(n51876), .B2(n22315), .ZN(
        n51877) );
  INV_X1 U44656 ( .I(n60742), .ZN(n60741) );
  XOR2_X1 U44660 ( .A1(n21172), .A2(n4615), .Z(n60743) );
  XOR2_X1 U44678 ( .A1(n6106), .A2(n6105), .Z(n6115) );
  XOR2_X1 U44712 ( .A1(n60744), .A2(n18687), .Z(n51344) );
  AND3_X1 U44750 ( .A1(n48987), .A2(n48985), .A3(n48986), .Z(n61682) );
  NAND2_X2 U44753 ( .A1(n8734), .A2(n21293), .ZN(n37875) );
  NOR2_X2 U44756 ( .A1(n21691), .A2(n10100), .ZN(n8734) );
  OR2_X2 U44832 ( .A1(n815), .A2(n12477), .Z(n28176) );
  XOR2_X1 U44878 ( .A1(n52352), .A2(n26022), .Z(n22059) );
  XOR2_X1 U44912 ( .A1(n23016), .A2(n52465), .Z(n52352) );
  NAND2_X2 U44920 ( .A1(n24522), .A2(n2323), .ZN(n6867) );
  NAND2_X1 U44932 ( .A1(n25170), .A2(n54960), .ZN(n55031) );
  INV_X1 U44972 ( .I(n10922), .ZN(n60749) );
  NOR2_X1 U44984 ( .A1(n21440), .A2(n21441), .ZN(n21439) );
  XOR2_X1 U44987 ( .A1(n60752), .A2(n54716), .Z(Plaintext[80]) );
  NAND2_X1 U44989 ( .A1(n54656), .A2(n54657), .ZN(n54660) );
  NAND2_X1 U45017 ( .A1(n30544), .A2(n29977), .ZN(n3816) );
  NAND2_X1 U45056 ( .A1(n24779), .A2(n59139), .ZN(n60754) );
  XOR2_X1 U45078 ( .A1(n44184), .A2(n8108), .Z(n46161) );
  XOR2_X1 U45128 ( .A1(n7535), .A2(n6722), .Z(n60755) );
  XOR2_X1 U45157 ( .A1(n44129), .A2(n16599), .Z(n45844) );
  NOR3_X2 U45209 ( .A1(n35434), .A2(n35435), .A3(n14629), .ZN(n60759) );
  XOR2_X1 U45211 ( .A1(n32722), .A2(n20862), .Z(n32573) );
  OAI21_X2 U45212 ( .A1(n25635), .A2(n23794), .B(n61374), .ZN(n32722) );
  XOR2_X1 U45250 ( .A1(n5332), .A2(n60760), .Z(n60967) );
  BUF_X2 U45251 ( .I(n17922), .Z(n60763) );
  BUF_X2 U45272 ( .I(n7323), .Z(n60765) );
  NAND2_X1 U45277 ( .A1(n28147), .A2(n59935), .ZN(n60766) );
  XOR2_X1 U45305 ( .A1(n60776), .A2(n25599), .Z(n3568) );
  XOR2_X1 U45340 ( .A1(n44964), .A2(n46384), .Z(n60776) );
  XOR2_X1 U45354 ( .A1(n15149), .A2(n15047), .Z(n13574) );
  XOR2_X1 U45372 ( .A1(n19433), .A2(n5448), .Z(n60777) );
  XOR2_X1 U45396 ( .A1(n43935), .A2(n43934), .Z(n60778) );
  XOR2_X1 U45417 ( .A1(n32230), .A2(n4341), .Z(n4339) );
  INV_X4 U45485 ( .I(n56757), .ZN(n56808) );
  OR2_X2 U45547 ( .A1(n51353), .A2(n51352), .Z(n56757) );
  NAND3_X1 U45552 ( .A1(n17635), .A2(n9555), .A3(n51347), .ZN(n51349) );
  NAND2_X1 U45586 ( .A1(n52725), .A2(n56868), .ZN(n60780) );
  NAND2_X1 U45587 ( .A1(n21752), .A2(n30251), .ZN(n60782) );
  NOR2_X2 U45612 ( .A1(n60784), .A2(n60783), .ZN(n4873) );
  NOR2_X2 U45613 ( .A1(n40948), .A2(n40949), .ZN(n60784) );
  NOR2_X1 U45657 ( .A1(n15753), .A2(n617), .ZN(n49329) );
  XOR2_X1 U45688 ( .A1(n17518), .A2(n43766), .Z(n17517) );
  XOR2_X1 U45698 ( .A1(n44084), .A2(n45099), .Z(n43766) );
  NOR3_X2 U45704 ( .A1(n15094), .A2(n28248), .A3(n28253), .ZN(n30450) );
  XOR2_X1 U45716 ( .A1(n60788), .A2(n52735), .Z(Plaintext[177]) );
  NAND2_X1 U45717 ( .A1(n60789), .A2(n53159), .ZN(n22281) );
  NAND2_X2 U45753 ( .A1(n54754), .A2(n54728), .ZN(n54736) );
  NOR2_X2 U45758 ( .A1(n12468), .A2(n56659), .ZN(n56374) );
  NAND2_X2 U45774 ( .A1(n44082), .A2(n45373), .ZN(n8319) );
  NAND4_X1 U45777 ( .A1(n54236), .A2(n54234), .A3(n54235), .A4(n54237), .ZN(
        n54248) );
  XNOR2_X1 U45819 ( .A1(n44596), .A2(n44597), .ZN(n16196) );
  XOR2_X1 U45840 ( .A1(n15489), .A2(n60795), .Z(n31455) );
  XOR2_X1 U45859 ( .A1(n31450), .A2(n31449), .Z(n60795) );
  BUF_X2 U45881 ( .I(n56030), .Z(n60797) );
  NAND2_X2 U45921 ( .A1(n1484), .A2(n45724), .ZN(n4233) );
  NOR3_X2 U45958 ( .A1(n23159), .A2(n6473), .A3(n60804), .ZN(n60803) );
  INV_X2 U45960 ( .I(n16658), .ZN(n46822) );
  NAND2_X2 U46008 ( .A1(n47372), .A2(n15162), .ZN(n16658) );
  XOR2_X1 U46020 ( .A1(n31568), .A2(n26133), .Z(n31577) );
  NAND3_X2 U46047 ( .A1(n41040), .A2(n41038), .A3(n41039), .ZN(n41041) );
  NAND3_X2 U46049 ( .A1(n22010), .A2(n47285), .A3(n22008), .ZN(n60898) );
  AOI21_X2 U46060 ( .A1(n34343), .A2(n35295), .B(n60805), .ZN(n61501) );
  NAND2_X2 U46098 ( .A1(n56983), .A2(n56986), .ZN(n52682) );
  AND3_X1 U46109 ( .A1(n48330), .A2(n47787), .A3(n6027), .Z(n14843) );
  NAND2_X2 U46111 ( .A1(n7806), .A2(n60807), .ZN(n16491) );
  INV_X2 U46139 ( .I(n5029), .ZN(n4686) );
  NAND4_X2 U46156 ( .A1(n24603), .A2(n27779), .A3(n27778), .A4(n27777), .ZN(
        n23130) );
  NAND2_X1 U46157 ( .A1(n56218), .A2(n56219), .ZN(n56223) );
  BUF_X4 U46161 ( .I(n21945), .Z(n60808) );
  XOR2_X1 U46179 ( .A1(n38491), .A2(n57455), .Z(n3213) );
  NAND2_X2 U46222 ( .A1(n15759), .A2(n17452), .ZN(n48234) );
  BUF_X2 U46226 ( .I(n23873), .Z(n60809) );
  BUF_X2 U46228 ( .I(n40713), .Z(n60810) );
  INV_X1 U46376 ( .I(n6333), .ZN(n60814) );
  OAI22_X1 U46422 ( .A1(n10900), .A2(n35749), .B1(n35748), .B2(n15148), .ZN(
        n35752) );
  NOR2_X2 U46434 ( .A1(n11552), .A2(n47629), .ZN(n48711) );
  NOR2_X1 U46442 ( .A1(n40958), .A2(n60820), .ZN(n965) );
  NAND2_X2 U46454 ( .A1(n38600), .A2(n25139), .ZN(n40958) );
  INV_X2 U46466 ( .I(n60821), .ZN(n25742) );
  NAND2_X2 U46485 ( .A1(n3580), .A2(n8478), .ZN(n29118) );
  OAI21_X1 U46543 ( .A1(n36719), .A2(n34937), .B(n19012), .ZN(n60823) );
  NOR2_X2 U46549 ( .A1(n12933), .A2(n33916), .ZN(n35086) );
  NOR2_X2 U46586 ( .A1(n17615), .A2(n21104), .ZN(n13767) );
  XOR2_X1 U46601 ( .A1(n56762), .A2(n60828), .Z(n38388) );
  INV_X1 U46633 ( .I(n60829), .ZN(n17291) );
  OAI21_X1 U46634 ( .A1(n26408), .A2(n26409), .B(n21068), .ZN(n60829) );
  NOR2_X2 U46700 ( .A1(n2811), .A2(n60830), .ZN(n25598) );
  NOR3_X1 U46755 ( .A1(n36725), .A2(n1418), .A3(n59147), .ZN(n22494) );
  XNOR2_X1 U46768 ( .A1(n39660), .A2(n13686), .ZN(n61109) );
  NAND3_X1 U46805 ( .A1(n42438), .A2(n1981), .A3(n41820), .ZN(n41821) );
  XOR2_X1 U46860 ( .A1(n26100), .A2(n50414), .Z(n6210) );
  BUF_X2 U46861 ( .I(n35240), .Z(n60835) );
  NAND2_X1 U46903 ( .A1(n48244), .A2(n6957), .ZN(n60838) );
  XOR2_X1 U46904 ( .A1(n60840), .A2(n10553), .Z(n33232) );
  NOR2_X2 U46942 ( .A1(n377), .A2(n10673), .ZN(n826) );
  XOR2_X1 U47077 ( .A1(n4370), .A2(n60842), .Z(n4532) );
  XOR2_X1 U47090 ( .A1(n20229), .A2(n806), .Z(n60842) );
  NAND2_X2 U47140 ( .A1(n21495), .A2(n16666), .ZN(n15817) );
  NOR2_X2 U47158 ( .A1(n49948), .A2(n1209), .ZN(n376) );
  XOR2_X1 U47179 ( .A1(n60844), .A2(n32562), .Z(n1953) );
  XOR2_X1 U47184 ( .A1(n1955), .A2(n31682), .Z(n60844) );
  INV_X1 U47204 ( .I(n34306), .ZN(n34760) );
  NAND3_X1 U47340 ( .A1(n44710), .A2(n44711), .A3(n45784), .ZN(n60850) );
  BUF_X2 U47410 ( .I(n16342), .Z(n60855) );
  NOR2_X2 U47434 ( .A1(n61499), .A2(n16056), .ZN(n17236) );
  INV_X2 U47514 ( .I(n48338), .ZN(n49904) );
  NAND4_X2 U47527 ( .A1(n18320), .A2(n18318), .A3(n18324), .A4(n18319), .ZN(
        n48338) );
  NAND3_X2 U47529 ( .A1(n61326), .A2(n47915), .A3(n61327), .ZN(n60856) );
  BUF_X2 U47530 ( .I(n48764), .Z(n60857) );
  AND2_X1 U47531 ( .A1(n30639), .A2(n23901), .Z(n60858) );
  XOR2_X1 U47548 ( .A1(n50844), .A2(n50848), .Z(n60859) );
  NAND3_X1 U47549 ( .A1(n61859), .A2(n1708), .A3(n43601), .ZN(n1006) );
  NAND2_X2 U47565 ( .A1(n12677), .A2(n22228), .ZN(n17176) );
  NOR2_X1 U47594 ( .A1(n13828), .A2(n14030), .ZN(n60861) );
  NAND2_X2 U47612 ( .A1(n25118), .A2(n40928), .ZN(n20871) );
  NAND2_X2 U47628 ( .A1(n40481), .A2(n40255), .ZN(n40896) );
  XOR2_X1 U47630 ( .A1(n60863), .A2(n19341), .Z(n30999) );
  XOR2_X1 U47631 ( .A1(n30996), .A2(n15725), .Z(n60863) );
  XOR2_X1 U47673 ( .A1(n39196), .A2(n38699), .Z(n39707) );
  NAND2_X2 U47689 ( .A1(n55157), .A2(n55132), .ZN(n55148) );
  NOR2_X2 U47717 ( .A1(n2618), .A2(n1430), .ZN(n34277) );
  XOR2_X1 U47750 ( .A1(n2059), .A2(n35130), .Z(n7168) );
  NOR3_X2 U47813 ( .A1(n57468), .A2(n7666), .A3(n7408), .ZN(n60865) );
  NAND3_X2 U47825 ( .A1(n19024), .A2(n3308), .A3(n10175), .ZN(n33771) );
  NAND2_X2 U47842 ( .A1(n3425), .A2(n7513), .ZN(n46283) );
  XOR2_X1 U47850 ( .A1(n10713), .A2(n43856), .Z(n3038) );
  NAND4_X2 U47852 ( .A1(n60868), .A2(n34537), .A3(n34540), .A4(n34541), .ZN(
        n684) );
  NAND3_X1 U47859 ( .A1(n34533), .A2(n34532), .A3(n20895), .ZN(n60868) );
  NAND2_X2 U47860 ( .A1(n24100), .A2(n24101), .ZN(n46282) );
  XOR2_X1 U47914 ( .A1(n19395), .A2(n30906), .Z(n60869) );
  XOR2_X1 U47925 ( .A1(n4144), .A2(n4146), .Z(n61653) );
  XOR2_X1 U47926 ( .A1(n60870), .A2(n56933), .Z(Plaintext[183]) );
  NAND2_X2 U47943 ( .A1(n2852), .A2(n60871), .ZN(n53997) );
  NOR2_X2 U47948 ( .A1(n21755), .A2(n47036), .ZN(n11416) );
  INV_X2 U47975 ( .I(n60875), .ZN(n5147) );
  XOR2_X1 U47976 ( .A1(n13366), .A2(n5148), .Z(n60875) );
  XOR2_X1 U47984 ( .A1(n25331), .A2(n60876), .Z(n30998) );
  XOR2_X1 U47986 ( .A1(n31446), .A2(n20673), .Z(n60876) );
  INV_X2 U48006 ( .I(n1681), .ZN(n14059) );
  XOR2_X1 U48012 ( .A1(n60877), .A2(n45281), .Z(n1681) );
  NOR2_X2 U48058 ( .A1(n17410), .A2(n16631), .ZN(n60878) );
  OAI22_X1 U48059 ( .A1(n17687), .A2(n36777), .B1(n17685), .B2(n12031), .ZN(
        n11300) );
  AND2_X1 U48060 ( .A1(n18419), .A2(n18411), .Z(n60880) );
  BUF_X2 U48102 ( .I(n47843), .Z(n60881) );
  NAND2_X2 U48156 ( .A1(n21035), .A2(n21487), .ZN(n35820) );
  BUF_X4 U48157 ( .I(n15738), .Z(n61215) );
  XOR2_X1 U48230 ( .A1(n21984), .A2(n5165), .Z(n25483) );
  XOR2_X1 U48239 ( .A1(n14867), .A2(n32568), .Z(n60887) );
  XOR2_X1 U48244 ( .A1(n60888), .A2(n21369), .Z(n4057) );
  XOR2_X1 U48293 ( .A1(n60927), .A2(n5854), .Z(n4570) );
  NOR2_X2 U48305 ( .A1(n13983), .A2(n36959), .ZN(n5483) );
  BUF_X2 U48306 ( .I(n33948), .Z(n60892) );
  NOR2_X2 U48328 ( .A1(n60899), .A2(n10698), .ZN(n36052) );
  XOR2_X1 U48368 ( .A1(n3035), .A2(n45128), .Z(n60903) );
  XOR2_X1 U48372 ( .A1(n60904), .A2(n52499), .Z(n52475) );
  XOR2_X1 U48375 ( .A1(n1915), .A2(n52469), .Z(n60904) );
  OR2_X1 U48415 ( .A1(n35036), .A2(n31302), .Z(n60908) );
  NOR2_X2 U48416 ( .A1(n1868), .A2(n26084), .ZN(n31114) );
  NOR2_X2 U48418 ( .A1(n19080), .A2(n63006), .ZN(n53097) );
  AOI21_X2 U48420 ( .A1(n52848), .A2(n52846), .B(n50676), .ZN(n60909) );
  OR2_X1 U48433 ( .A1(n47030), .A2(n45536), .Z(n19326) );
  XOR2_X1 U48465 ( .A1(n24978), .A2(n9605), .Z(n60910) );
  NAND2_X2 U48467 ( .A1(n219), .A2(n60911), .ZN(n1196) );
  XOR2_X1 U48500 ( .A1(n60912), .A2(n52326), .Z(n55676) );
  XOR2_X1 U48503 ( .A1(n52028), .A2(n24470), .Z(n60912) );
  XOR2_X1 U48511 ( .A1(n61681), .A2(n60913), .Z(n52026) );
  XOR2_X1 U48512 ( .A1(n20780), .A2(n23670), .Z(n60913) );
  XOR2_X1 U48517 ( .A1(n50325), .A2(n17143), .Z(n60914) );
  XOR2_X1 U48535 ( .A1(n60915), .A2(n44397), .Z(n16994) );
  NOR3_X2 U48540 ( .A1(n7637), .A2(n60916), .A3(n777), .ZN(n8317) );
  OR2_X2 U48570 ( .A1(n47290), .A2(n14888), .Z(n2973) );
  XOR2_X1 U48580 ( .A1(n16369), .A2(n60919), .Z(n5836) );
  XOR2_X1 U48581 ( .A1(n39226), .A2(n39225), .Z(n60919) );
  XOR2_X1 U48606 ( .A1(n46409), .A2(n44625), .Z(n9497) );
  XOR2_X1 U48610 ( .A1(n2107), .A2(n2108), .Z(n60922) );
  NOR2_X2 U48618 ( .A1(n22814), .A2(n22813), .ZN(n61475) );
  NOR2_X1 U48636 ( .A1(n19281), .A2(n35399), .ZN(n60923) );
  NAND2_X2 U48639 ( .A1(n5250), .A2(n33540), .ZN(n33112) );
  BUF_X2 U48672 ( .I(n12479), .Z(n60926) );
  XOR2_X1 U48673 ( .A1(n39189), .A2(n57174), .Z(n60927) );
  BUF_X2 U48675 ( .I(n41007), .Z(n60928) );
  XOR2_X1 U48682 ( .A1(n3501), .A2(n20324), .Z(n4956) );
  XOR2_X1 U48695 ( .A1(n19551), .A2(n8374), .Z(n33031) );
  XOR2_X1 U48706 ( .A1(n60931), .A2(n129), .Z(n731) );
  INV_X2 U48719 ( .I(n7522), .ZN(n60931) );
  NAND3_X2 U48755 ( .A1(n4721), .A2(n43291), .A3(n60932), .ZN(n6565) );
  XOR2_X1 U48781 ( .A1(n31407), .A2(n26081), .Z(n5521) );
  XOR2_X1 U48801 ( .A1(n51677), .A2(n52559), .Z(n60) );
  INV_X2 U48827 ( .I(n33945), .ZN(n32864) );
  AND2_X1 U48870 ( .A1(n28772), .A2(n23317), .Z(n8357) );
  NAND2_X2 U48927 ( .A1(n58546), .A2(n14312), .ZN(n29351) );
  OAI21_X1 U48955 ( .A1(n56546), .A2(n51347), .B(n56386), .ZN(n51346) );
  NAND2_X2 U48956 ( .A1(n49465), .A2(n6313), .ZN(n5146) );
  NOR2_X2 U48983 ( .A1(n15587), .A2(n15586), .ZN(n16037) );
  NOR3_X2 U49065 ( .A1(n19338), .A2(n10222), .A3(n19339), .ZN(n25093) );
  NAND2_X1 U49066 ( .A1(n36396), .A2(n36538), .ZN(n60940) );
  XOR2_X1 U49072 ( .A1(n33060), .A2(n11383), .Z(n60941) );
  NAND2_X1 U49076 ( .A1(n60945), .A2(n6779), .ZN(n60943) );
  NAND2_X1 U49103 ( .A1(n16192), .A2(n17444), .ZN(n60945) );
  NOR3_X1 U49139 ( .A1(n25384), .A2(n60895), .A3(n31085), .ZN(n30555) );
  BUF_X2 U49153 ( .I(n36171), .Z(n60949) );
  INV_X2 U49218 ( .I(n22107), .ZN(n29993) );
  NAND2_X2 U49219 ( .A1(n17175), .A2(n17174), .ZN(n22107) );
  XOR2_X1 U49330 ( .A1(n9398), .A2(n60950), .Z(n22036) );
  XOR2_X1 U49331 ( .A1(n38916), .A2(n37656), .Z(n60950) );
  INV_X2 U49371 ( .I(n42867), .ZN(n60952) );
  NOR2_X2 U49386 ( .A1(n61039), .A2(n60955), .ZN(n41043) );
  NAND4_X2 U49409 ( .A1(n41025), .A2(n41026), .A3(n19173), .A4(n41024), .ZN(
        n60955) );
  NOR2_X2 U49481 ( .A1(n31469), .A2(n11643), .ZN(n34000) );
  NAND4_X2 U49482 ( .A1(n11601), .A2(n36629), .A3(n5528), .A4(n5527), .ZN(
        n37987) );
  XOR2_X1 U49483 ( .A1(n9430), .A2(n60963), .Z(n312) );
  XOR2_X1 U49485 ( .A1(n9432), .A2(n57285), .Z(n60963) );
  XOR2_X1 U49487 ( .A1(n52079), .A2(n60964), .Z(n26047) );
  INV_X2 U49488 ( .I(n14975), .ZN(n60964) );
  INV_X2 U49509 ( .I(n60967), .ZN(n52476) );
  XOR2_X1 U49517 ( .A1(n61927), .A2(n2612), .Z(n60968) );
  XOR2_X1 U49541 ( .A1(n18330), .A2(n3500), .Z(n20324) );
  XOR2_X1 U49546 ( .A1(n2278), .A2(n51164), .Z(n16744) );
  NOR2_X1 U49558 ( .A1(n39887), .A2(n20751), .ZN(n39888) );
  NAND2_X1 U49562 ( .A1(n42486), .A2(n40315), .ZN(n39887) );
  AND2_X2 U49630 ( .A1(n26110), .A2(n19065), .Z(n42200) );
  OR2_X1 U49658 ( .A1(n24210), .A2(n49803), .Z(n48432) );
  NAND3_X1 U49782 ( .A1(n55674), .A2(n17708), .A3(n4836), .ZN(n9267) );
  NAND3_X1 U49822 ( .A1(n34547), .A2(n60973), .A3(n476), .ZN(n7056) );
  NAND2_X1 U49941 ( .A1(n436), .A2(n127), .ZN(n60973) );
  BUF_X2 U49954 ( .I(n15245), .Z(n60974) );
  NAND2_X2 U49978 ( .A1(n9228), .A2(n60975), .ZN(n49476) );
  INV_X2 U49985 ( .I(n50359), .ZN(n60975) );
  NAND2_X2 U50075 ( .A1(n8914), .A2(n8915), .ZN(n8913) );
  NAND2_X2 U50157 ( .A1(n60977), .A2(n18323), .ZN(n15966) );
  NAND2_X2 U50168 ( .A1(n10389), .A2(n56567), .ZN(n55937) );
  NAND2_X2 U50179 ( .A1(n52126), .A2(n15454), .ZN(n55905) );
  XOR2_X1 U50188 ( .A1(n13885), .A2(n10825), .Z(n24650) );
  XOR2_X1 U50195 ( .A1(n60981), .A2(n12106), .Z(n35685) );
  XOR2_X1 U50199 ( .A1(n32726), .A2(n12103), .Z(n60981) );
  NAND2_X2 U50263 ( .A1(n57353), .A2(n56362), .ZN(n56237) );
  XOR2_X1 U50385 ( .A1(n44092), .A2(n22890), .Z(n44966) );
  NOR2_X1 U50386 ( .A1(n41651), .A2(n1702), .ZN(n60982) );
  INV_X2 U50476 ( .I(n29332), .ZN(n31255) );
  NAND2_X2 U50504 ( .A1(n52814), .A2(n57051), .ZN(n53445) );
  NAND2_X2 U50514 ( .A1(n436), .A2(n33509), .ZN(n33511) );
  XOR2_X1 U50515 ( .A1(n731), .A2(n32495), .Z(n8374) );
  AND2_X1 U50522 ( .A1(n47380), .A2(n23934), .Z(n17630) );
  XOR2_X1 U50524 ( .A1(n12559), .A2(n60987), .Z(n13914) );
  XOR2_X1 U50526 ( .A1(n31385), .A2(n30365), .Z(n60987) );
  NAND2_X1 U50533 ( .A1(n12365), .A2(n29281), .ZN(n60988) );
  NAND2_X1 U50541 ( .A1(n12366), .A2(n29626), .ZN(n60989) );
  NAND2_X2 U50565 ( .A1(n3650), .A2(n3647), .ZN(n22487) );
  NOR3_X2 U50570 ( .A1(n2298), .A2(n33528), .A3(n61642), .ZN(n3650) );
  INV_X2 U50598 ( .I(n60992), .ZN(n61681) );
  BUF_X2 U50604 ( .I(n22044), .Z(n60993) );
  XOR2_X1 U50605 ( .A1(n60994), .A2(n57232), .Z(n6808) );
  XOR2_X1 U50618 ( .A1(n14807), .A2(n11200), .Z(n60994) );
  XOR2_X1 U50642 ( .A1(n60996), .A2(n8866), .Z(n37725) );
  XOR2_X1 U50665 ( .A1(n7432), .A2(n22097), .Z(n60996) );
  XOR2_X1 U50668 ( .A1(n60997), .A2(n970), .Z(n2324) );
  XOR2_X1 U50672 ( .A1(n8516), .A2(n57403), .Z(n60997) );
  XOR2_X1 U50685 ( .A1(n60998), .A2(n37952), .Z(n43398) );
  XOR2_X1 U50690 ( .A1(n37758), .A2(n22458), .Z(n60998) );
  XOR2_X1 U50704 ( .A1(n25961), .A2(n60999), .Z(n7137) );
  NOR2_X2 U50705 ( .A1(n13315), .A2(n13314), .ZN(n25961) );
  NOR2_X2 U50777 ( .A1(n20842), .A2(n61001), .ZN(n35177) );
  NOR2_X1 U50779 ( .A1(n53578), .A2(n53577), .ZN(n53584) );
  NOR2_X1 U50789 ( .A1(n2744), .A2(n2745), .ZN(n11937) );
  XOR2_X1 U50844 ( .A1(n30994), .A2(n33226), .Z(n4615) );
  NAND3_X2 U50845 ( .A1(n30180), .A2(n17491), .A3(n17490), .ZN(n30994) );
  XOR2_X1 U50856 ( .A1(n31985), .A2(n17700), .Z(n12590) );
  OR2_X2 U50857 ( .A1(n3983), .A2(n3990), .Z(n17700) );
  INV_X1 U50860 ( .I(n19098), .ZN(n61285) );
  XOR2_X1 U50863 ( .A1(n9269), .A2(n61009), .Z(n38288) );
  BUF_X2 U50866 ( .I(n20950), .Z(n61010) );
  XOR2_X1 U50878 ( .A1(n39562), .A2(n24147), .Z(n61011) );
  XOR2_X1 U50885 ( .A1(n25479), .A2(n23232), .Z(n12930) );
  BUF_X2 U50886 ( .I(n14165), .Z(n61013) );
  NAND4_X2 U50888 ( .A1(n34181), .A2(n34183), .A3(n8095), .A4(n34182), .ZN(
        n34184) );
  NAND3_X1 U50892 ( .A1(n45537), .A2(n45784), .A3(n45783), .ZN(n61017) );
  AOI21_X1 U50936 ( .A1(n61018), .A2(n47037), .B(n13655), .ZN(n47039) );
  AND2_X1 U50974 ( .A1(n47034), .A2(n21755), .Z(n20298) );
  XOR2_X1 U50989 ( .A1(n65270), .A2(n39498), .Z(n39501) );
  XOR2_X1 U50990 ( .A1(n5376), .A2(n39299), .Z(n39498) );
  OAI22_X1 U50992 ( .A1(n47656), .A2(n10420), .B1(n47657), .B2(n14741), .ZN(
        n47662) );
  NAND4_X2 U50996 ( .A1(n61020), .A2(n33492), .A3(n33771), .A4(n34284), .ZN(
        n61306) );
  NAND2_X1 U50998 ( .A1(n33490), .A2(n34276), .ZN(n61020) );
  NAND2_X2 U51000 ( .A1(n4119), .A2(n4118), .ZN(n23874) );
  OR2_X1 U51004 ( .A1(n53363), .A2(n53364), .Z(n15361) );
  XOR2_X1 U51015 ( .A1(n45129), .A2(n61022), .Z(n4814) );
  XOR2_X1 U51016 ( .A1(n43887), .A2(n44805), .Z(n61022) );
  NAND2_X1 U51061 ( .A1(n56695), .A2(n56731), .ZN(n22025) );
  NAND3_X2 U51064 ( .A1(n52917), .A2(n52916), .A3(n61023), .ZN(n55216) );
  BUF_X2 U51065 ( .I(n47603), .Z(n61025) );
  XOR2_X1 U51068 ( .A1(n61026), .A2(n16106), .Z(n15223) );
  XOR2_X1 U51076 ( .A1(n61027), .A2(n9071), .Z(n11475) );
  XOR2_X1 U51082 ( .A1(n45024), .A2(n3417), .Z(n61027) );
  XOR2_X1 U51099 ( .A1(n20824), .A2(n46552), .Z(n3418) );
  XOR2_X1 U51109 ( .A1(n23905), .A2(n51016), .Z(n46552) );
  XOR2_X1 U51120 ( .A1(n61030), .A2(n22102), .Z(n13663) );
  XOR2_X1 U51131 ( .A1(n61032), .A2(n7365), .Z(n454) );
  XOR2_X1 U51141 ( .A1(n2937), .A2(n61033), .Z(n35329) );
  XOR2_X1 U51143 ( .A1(n2940), .A2(n2939), .Z(n61033) );
  BUF_X2 U51209 ( .I(n28025), .Z(n61035) );
  NOR2_X2 U51211 ( .A1(n17538), .A2(n25256), .ZN(n35295) );
  XOR2_X1 U51246 ( .A1(n31966), .A2(n21824), .Z(n61037) );
  XOR2_X1 U51270 ( .A1(n51738), .A2(n51600), .Z(n18641) );
  XOR2_X1 U51271 ( .A1(n25805), .A2(n51602), .Z(n51738) );
  XOR2_X1 U51291 ( .A1(n57586), .A2(n14253), .Z(n46145) );
  OR2_X1 U51312 ( .A1(n36485), .A2(n10829), .Z(n35554) );
  XOR2_X1 U51333 ( .A1(n61042), .A2(n61041), .Z(n399) );
  XOR2_X1 U51334 ( .A1(n14180), .A2(n25433), .Z(n61042) );
  AOI21_X1 U51390 ( .A1(n56504), .A2(n56517), .B(n15765), .ZN(n56505) );
  XOR2_X1 U51417 ( .A1(n39464), .A2(n10069), .Z(n16681) );
  INV_X2 U51426 ( .I(n61046), .ZN(n11767) );
  XOR2_X1 U51427 ( .A1(Ciphertext[189]), .A2(Key[64]), .Z(n61046) );
  INV_X4 U51433 ( .I(n5247), .ZN(n33848) );
  NOR2_X2 U51447 ( .A1(n64324), .A2(n20650), .ZN(n21527) );
  NOR2_X2 U51517 ( .A1(n28250), .A2(n27040), .ZN(n27386) );
  NAND2_X2 U51538 ( .A1(n28244), .A2(n26270), .ZN(n27040) );
  NOR2_X2 U51542 ( .A1(n14869), .A2(n20519), .ZN(n27229) );
  XOR2_X1 U51547 ( .A1(n2241), .A2(n46407), .Z(n362) );
  BUF_X2 U51648 ( .I(n28279), .Z(n61064) );
  BUF_X2 U51663 ( .I(n22807), .Z(n61065) );
  INV_X2 U51691 ( .I(n61067), .ZN(n24301) );
  NAND2_X1 U51732 ( .A1(n8784), .A2(n56538), .ZN(n14762) );
  AND2_X1 U51733 ( .A1(n35928), .A2(n35929), .Z(n25963) );
  OR2_X1 U51742 ( .A1(n9063), .A2(n43889), .Z(n22016) );
  XOR2_X1 U51752 ( .A1(n44838), .A2(n61072), .Z(n44839) );
  XOR2_X1 U51761 ( .A1(n61074), .A2(n20838), .Z(n16361) );
  XOR2_X1 U51775 ( .A1(n32383), .A2(n32056), .Z(n61074) );
  XOR2_X1 U51800 ( .A1(n61732), .A2(n22806), .Z(n31316) );
  XOR2_X1 U51804 ( .A1(n61075), .A2(n32757), .Z(n23735) );
  XOR2_X1 U51805 ( .A1(n20940), .A2(n32059), .Z(n61075) );
  XOR2_X1 U51893 ( .A1(n61077), .A2(n859), .Z(n25413) );
  XOR2_X1 U51894 ( .A1(n51731), .A2(n51027), .Z(n61077) );
  OR2_X1 U51897 ( .A1(n25233), .A2(n18606), .Z(n21189) );
  BUF_X2 U51912 ( .I(n34083), .Z(n61078) );
  NOR2_X2 U51939 ( .A1(n7426), .A2(n15738), .ZN(n8364) );
  OAI21_X1 U51940 ( .A1(n12616), .A2(n3348), .B(n61079), .ZN(n3352) );
  BUF_X2 U51962 ( .I(n22947), .Z(n61081) );
  NAND2_X2 U51963 ( .A1(n17285), .A2(n26777), .ZN(n27278) );
  NAND4_X2 U51970 ( .A1(n57253), .A2(n29555), .A3(n29554), .A4(n202), .ZN(
        n26038) );
  XOR2_X1 U51990 ( .A1(n12119), .A2(n3193), .Z(n61082) );
  NAND2_X1 U52044 ( .A1(n21268), .A2(n24870), .ZN(n54647) );
  XOR2_X1 U52070 ( .A1(n2858), .A2(n24780), .Z(n32496) );
  OAI21_X1 U52073 ( .A1(n61086), .A2(n1405), .B(n41456), .ZN(n14948) );
  NOR2_X1 U52075 ( .A1(n58798), .A2(n41455), .ZN(n61086) );
  XOR2_X1 U52109 ( .A1(n11636), .A2(n38307), .Z(n36638) );
  NAND3_X2 U52120 ( .A1(n35413), .A2(n35412), .A3(n35411), .ZN(n38307) );
  AOI21_X2 U52121 ( .A1(n34612), .A2(n34611), .B(n61087), .ZN(n15227) );
  BUF_X2 U52144 ( .I(n9329), .Z(n61090) );
  NOR3_X2 U52153 ( .A1(n45310), .A2(n45309), .A3(n47708), .ZN(n45313) );
  NAND2_X2 U52182 ( .A1(n1433), .A2(n4567), .ZN(n30803) );
  INV_X2 U52205 ( .I(n61095), .ZN(n61668) );
  NAND2_X2 U52219 ( .A1(n12468), .A2(n56659), .ZN(n61202) );
  NAND2_X2 U52222 ( .A1(n29241), .A2(n10820), .ZN(n29929) );
  NAND2_X2 U52225 ( .A1(n24091), .A2(n55677), .ZN(n55973) );
  OAI21_X2 U52262 ( .A1(n13588), .A2(n48184), .B(n58974), .ZN(n48583) );
  NOR2_X2 U52330 ( .A1(n48176), .A2(n10621), .ZN(n48184) );
  OAI22_X1 U52370 ( .A1(n34186), .A2(n24153), .B1(n64234), .B2(n59328), .ZN(
        n7865) );
  NAND2_X2 U52389 ( .A1(n16392), .A2(n16393), .ZN(n43464) );
  XOR2_X1 U52391 ( .A1(n51042), .A2(n24031), .Z(n7752) );
  XOR2_X1 U52429 ( .A1(n58891), .A2(n39380), .Z(n61099) );
  INV_X2 U52436 ( .I(n23116), .ZN(n12111) );
  XOR2_X1 U52439 ( .A1(n6251), .A2(n17271), .Z(n61100) );
  XOR2_X1 U52513 ( .A1(n61101), .A2(n18809), .Z(n21016) );
  XOR2_X1 U52517 ( .A1(n39545), .A2(n39544), .Z(n61101) );
  XOR2_X1 U52528 ( .A1(n61102), .A2(n11185), .Z(n2917) );
  XOR2_X1 U52531 ( .A1(n52197), .A2(n51611), .Z(n36632) );
  XOR2_X1 U52537 ( .A1(n52317), .A2(n56155), .Z(n51611) );
  NAND2_X1 U52540 ( .A1(n61081), .A2(n21248), .ZN(n15974) );
  NAND3_X1 U52557 ( .A1(n41408), .A2(n41405), .A3(n1303), .ZN(n61103) );
  XOR2_X1 U52564 ( .A1(n25376), .A2(n61104), .Z(n38987) );
  XOR2_X1 U52567 ( .A1(n39743), .A2(n61105), .Z(n61104) );
  XOR2_X1 U52611 ( .A1(n61106), .A2(n7132), .Z(n46591) );
  XOR2_X1 U52627 ( .A1(n19232), .A2(n10160), .Z(n61106) );
  OAI21_X1 U52632 ( .A1(n30819), .A2(n30820), .B(n30818), .ZN(n30824) );
  NOR2_X2 U52659 ( .A1(n61187), .A2(n29835), .ZN(n30818) );
  NAND2_X2 U52662 ( .A1(n27966), .A2(n2295), .ZN(n28279) );
  NAND3_X2 U52671 ( .A1(n59601), .A2(n39959), .A3(n40568), .ZN(n39485) );
  XOR2_X1 U52708 ( .A1(n61110), .A2(n23207), .Z(n26210) );
  XOR2_X1 U52722 ( .A1(n2458), .A2(n4349), .Z(n61110) );
  NAND2_X2 U52723 ( .A1(n26756), .A2(n26797), .ZN(n27880) );
  NAND2_X1 U52732 ( .A1(n34274), .A2(n34273), .ZN(n61111) );
  NAND2_X1 U52737 ( .A1(n27098), .A2(n10537), .ZN(n6863) );
  NOR2_X1 U52746 ( .A1(n17551), .A2(n34024), .ZN(n34032) );
  OR2_X1 U52796 ( .A1(n13980), .A2(n13981), .Z(n61112) );
  OR2_X1 U52805 ( .A1(n6679), .A2(n5629), .Z(n47057) );
  NOR2_X2 U52823 ( .A1(n10968), .A2(n54112), .ZN(n9136) );
  INV_X2 U52845 ( .I(n61116), .ZN(n25244) );
  XOR2_X1 U52857 ( .A1(n32185), .A2(n12811), .Z(n61117) );
  AND2_X1 U52863 ( .A1(n43450), .A2(n43444), .Z(n455) );
  NAND2_X2 U52927 ( .A1(n42732), .A2(n14920), .ZN(n61121) );
  BUF_X2 U52934 ( .I(n54017), .Z(n61123) );
  INV_X1 U52972 ( .I(n53763), .ZN(n61127) );
  XOR2_X1 U52986 ( .A1(n31926), .A2(n31925), .Z(n32237) );
  XOR2_X1 U53003 ( .A1(n32044), .A2(n22820), .Z(n31926) );
  XOR2_X1 U53032 ( .A1(n12769), .A2(n61128), .Z(n46545) );
  XOR2_X1 U53035 ( .A1(n7628), .A2(n61663), .Z(n12769) );
  XOR2_X1 U53038 ( .A1(n61130), .A2(n61129), .Z(n5622) );
  AOI21_X1 U53040 ( .A1(n30341), .A2(n30342), .B(n61131), .ZN(n15979) );
  XOR2_X1 U53042 ( .A1(n61132), .A2(n9557), .Z(n9558) );
  BUF_X2 U53043 ( .I(n21364), .Z(n61133) );
  NAND3_X1 U53048 ( .A1(n17549), .A2(n49815), .A3(n50441), .ZN(n47148) );
  XOR2_X1 U53053 ( .A1(n61135), .A2(n53464), .Z(Plaintext[24]) );
  NOR4_X2 U53054 ( .A1(n5965), .A2(n5968), .A3(n5966), .A4(n25739), .ZN(n61135) );
  OR2_X2 U53075 ( .A1(n15777), .A2(n56585), .Z(n56592) );
  NOR2_X2 U53118 ( .A1(n20832), .A2(n23588), .ZN(n47312) );
  AND3_X1 U53139 ( .A1(n25779), .A2(n47608), .A3(n47825), .Z(n61138) );
  NAND3_X2 U53140 ( .A1(n61140), .A2(n15612), .A3(n15613), .ZN(n36116) );
  XOR2_X1 U53151 ( .A1(n61143), .A2(n26158), .Z(n47323) );
  XOR2_X1 U53167 ( .A1(n39600), .A2(n10488), .Z(n39842) );
  XOR2_X1 U53198 ( .A1(n33880), .A2(n33883), .Z(n10904) );
  NOR2_X2 U53234 ( .A1(n4941), .A2(n29300), .ZN(n18739) );
  XOR2_X1 U53256 ( .A1(n9255), .A2(n9121), .Z(n39249) );
  NAND2_X2 U53281 ( .A1(n2618), .A2(n1815), .ZN(n3308) );
  XOR2_X1 U53292 ( .A1(n2615), .A2(n61145), .Z(n353) );
  XOR2_X1 U53322 ( .A1(n15512), .A2(n8111), .Z(n61145) );
  BUF_X2 U53326 ( .I(n3271), .Z(n61146) );
  NOR3_X2 U53347 ( .A1(n27480), .A2(n27546), .A3(n27537), .ZN(n27544) );
  XOR2_X1 U53377 ( .A1(n256), .A2(n9855), .Z(n44744) );
  NOR2_X2 U53404 ( .A1(n16852), .A2(n1410), .ZN(n18649) );
  XOR2_X1 U53473 ( .A1(n7601), .A2(n5730), .Z(n5729) );
  NAND2_X1 U53485 ( .A1(n19704), .A2(n48823), .ZN(n61151) );
  XOR2_X1 U53500 ( .A1(n61153), .A2(n31917), .Z(n31754) );
  XOR2_X1 U53504 ( .A1(n9055), .A2(n766), .Z(n61153) );
  XOR2_X1 U53509 ( .A1(n22975), .A2(n21170), .Z(n43796) );
  INV_X2 U53528 ( .I(n61156), .ZN(n1239) );
  NOR3_X2 U53534 ( .A1(n61158), .A2(n6732), .A3(n61157), .ZN(n22509) );
  INV_X1 U53538 ( .I(n24333), .ZN(n61158) );
  NOR2_X2 U53553 ( .A1(n27480), .A2(n27481), .ZN(n27550) );
  OR2_X1 U53580 ( .A1(n48927), .A2(n48366), .Z(n48767) );
  NAND2_X2 U53589 ( .A1(n1780), .A2(n37084), .ZN(n7662) );
  NOR2_X2 U53620 ( .A1(n5108), .A2(n5107), .ZN(n5105) );
  AOI21_X1 U53624 ( .A1(n7465), .A2(n14330), .B(n18244), .ZN(n61167) );
  INV_X2 U53625 ( .I(n61169), .ZN(n28553) );
  NOR2_X2 U53628 ( .A1(n7355), .A2(n10530), .ZN(n24210) );
  XOR2_X1 U53640 ( .A1(n61173), .A2(n10884), .Z(n7309) );
  XOR2_X1 U53642 ( .A1(n19348), .A2(n16246), .Z(n61173) );
  INV_X1 U53651 ( .I(n36899), .ZN(n23764) );
  XOR2_X1 U53662 ( .A1(n3038), .A2(n3037), .Z(n45128) );
  AND2_X1 U53794 ( .A1(n63261), .A2(n16336), .Z(n3462) );
  AND2_X1 U53801 ( .A1(n2350), .A2(n30211), .Z(n2349) );
  NAND2_X2 U53809 ( .A1(n3733), .A2(n45183), .ZN(n8475) );
  NAND2_X2 U53811 ( .A1(n6157), .A2(n1664), .ZN(n3733) );
  OR2_X1 U53812 ( .A1(n39074), .A2(n61183), .Z(n39076) );
  NAND2_X2 U53818 ( .A1(n30419), .A2(n30558), .ZN(n18060) );
  NAND4_X2 U53823 ( .A1(n48270), .A2(n61184), .A3(n49997), .A4(n4391), .ZN(
        n61576) );
  NAND2_X1 U53832 ( .A1(n42808), .A2(n43316), .ZN(n14988) );
  XOR2_X1 U53855 ( .A1(n3724), .A2(n6358), .Z(n6357) );
  XOR2_X1 U53865 ( .A1(n11185), .A2(n8899), .Z(n3724) );
  NOR3_X2 U53868 ( .A1(n54632), .A2(n54631), .A3(n54633), .ZN(n54667) );
  INV_X2 U53896 ( .I(n22557), .ZN(n24352) );
  XOR2_X1 U53903 ( .A1(n25497), .A2(n50762), .Z(n22557) );
  XOR2_X1 U53967 ( .A1(n51572), .A2(n50038), .Z(n5725) );
  NOR2_X1 U53999 ( .A1(n17204), .A2(n61193), .ZN(n53508) );
  NOR2_X2 U54004 ( .A1(n14537), .A2(n53518), .ZN(n17204) );
  INV_X1 U54006 ( .I(n56894), .ZN(n61221) );
  NOR2_X2 U54020 ( .A1(n9959), .A2(n17305), .ZN(n25939) );
  INV_X2 U54065 ( .I(n26077), .ZN(n61196) );
  NAND3_X1 U54109 ( .A1(n27001), .A2(n23708), .A3(n28582), .ZN(n5136) );
  XOR2_X1 U54121 ( .A1(n21488), .A2(n2763), .Z(n2762) );
  NAND2_X1 U54174 ( .A1(n48026), .A2(n49948), .ZN(n10740) );
  NOR3_X2 U54202 ( .A1(n26763), .A2(n27883), .A3(n26762), .ZN(n28780) );
  NAND2_X2 U54253 ( .A1(n61609), .A2(n188), .ZN(n27516) );
  OR2_X1 U54254 ( .A1(n35673), .A2(n57200), .Z(n4677) );
  NOR2_X2 U54318 ( .A1(n52866), .A2(n5536), .ZN(n53241) );
  OR2_X1 U54348 ( .A1(n25589), .A2(n61210), .Z(n50242) );
  NOR2_X2 U54360 ( .A1(n14266), .A2(n19144), .ZN(n25589) );
  NAND3_X2 U54366 ( .A1(n21634), .A2(n17925), .A3(n17926), .ZN(n51918) );
  NOR2_X2 U54453 ( .A1(n61221), .A2(n60708), .ZN(n56880) );
  NAND3_X2 U54464 ( .A1(n52776), .A2(n52774), .A3(n52775), .ZN(n52803) );
  XOR2_X1 U54498 ( .A1(n61226), .A2(n20191), .Z(n17486) );
  NOR2_X2 U54595 ( .A1(n52712), .A2(n627), .ZN(n56894) );
  AND2_X1 U54620 ( .A1(n45685), .A2(n47588), .Z(n61231) );
  XOR2_X1 U54626 ( .A1(n51017), .A2(n57229), .Z(n52164) );
  XOR2_X1 U54631 ( .A1(n24277), .A2(n5200), .Z(n38526) );
  BUF_X2 U54637 ( .I(n23348), .Z(n61233) );
  XOR2_X1 U54642 ( .A1(n61234), .A2(n49337), .Z(n25745) );
  XOR2_X1 U54678 ( .A1(n4112), .A2(n3690), .Z(n61234) );
  NOR2_X2 U54682 ( .A1(n61889), .A2(n2570), .ZN(n16162) );
  INV_X2 U54738 ( .I(n61236), .ZN(n9243) );
  NOR2_X1 U54765 ( .A1(n57299), .A2(n43304), .ZN(n61283) );
  XOR2_X1 U54778 ( .A1(n6717), .A2(n1947), .Z(n61240) );
  XOR2_X1 U54799 ( .A1(n2182), .A2(n61243), .Z(n55280) );
  XOR2_X1 U54801 ( .A1(n2167), .A2(n7612), .Z(n61243) );
  OAI22_X1 U54803 ( .A1(n61169), .A2(n29187), .B1(n16812), .B2(n28557), .ZN(
        n26409) );
  BUF_X2 U54837 ( .I(n14352), .Z(n61247) );
  OAI21_X1 U54851 ( .A1(n40400), .A2(n61250), .B(n4383), .ZN(n41417) );
  NOR2_X1 U54862 ( .A1(n41419), .A2(n58794), .ZN(n61250) );
  BUF_X2 U54869 ( .I(n31264), .Z(n61251) );
  XOR2_X1 U54918 ( .A1(n61252), .A2(n14348), .Z(n14612) );
  INV_X2 U54929 ( .I(n61253), .ZN(n1161) );
  NAND2_X2 U54930 ( .A1(n25675), .A2(n23611), .ZN(n61253) );
  NAND2_X1 U54966 ( .A1(n27393), .A2(n27395), .ZN(n61255) );
  XOR2_X1 U54978 ( .A1(n18702), .A2(n61257), .Z(n18701) );
  XOR2_X1 U54982 ( .A1(n20008), .A2(n50110), .Z(n61257) );
  NOR2_X1 U54986 ( .A1(n6598), .A2(n39424), .ZN(n39426) );
  NAND4_X2 U54988 ( .A1(n15039), .A2(n20971), .A3(n49677), .A4(n49675), .ZN(
        n61258) );
  NOR2_X2 U54993 ( .A1(n43839), .A2(n10990), .ZN(n43205) );
  XOR2_X1 U54999 ( .A1(n6326), .A2(n44609), .Z(n61263) );
  XOR2_X1 U55021 ( .A1(n31013), .A2(n2650), .Z(n61265) );
  NOR2_X1 U55072 ( .A1(n14936), .A2(n61618), .ZN(n61617) );
  XOR2_X1 U55073 ( .A1(n6322), .A2(n33827), .Z(n2131) );
  XOR2_X1 U55078 ( .A1(n15153), .A2(n59938), .Z(n33827) );
  NAND4_X2 U55116 ( .A1(n35535), .A2(n35537), .A3(n35536), .A4(n35538), .ZN(
        n61267) );
  NAND2_X2 U55145 ( .A1(n19873), .A2(n37440), .ZN(n39566) );
  INV_X4 U55164 ( .I(n19313), .ZN(n22503) );
  INV_X2 U55169 ( .I(n61270), .ZN(n740) );
  OR3_X1 U55171 ( .A1(n30579), .A2(n28207), .A3(n14921), .Z(n61272) );
  XOR2_X1 U55176 ( .A1(n18453), .A2(n18832), .Z(n6501) );
  NAND2_X2 U55178 ( .A1(n20555), .A2(n61407), .ZN(n38692) );
  AOI21_X2 U55183 ( .A1(n61685), .A2(n52883), .B(n17540), .ZN(n61277) );
  OAI21_X2 U55204 ( .A1(n46861), .A2(n10910), .B(n20426), .ZN(n61278) );
  XOR2_X1 U55208 ( .A1(n24047), .A2(n44944), .Z(n45602) );
  XOR2_X1 U55213 ( .A1(n21707), .A2(n61279), .Z(n14847) );
  XOR2_X1 U55238 ( .A1(n51406), .A2(n52584), .Z(n13922) );
  XOR2_X1 U55243 ( .A1(n50767), .A2(n7711), .Z(n51406) );
  NAND2_X1 U55244 ( .A1(n4021), .A2(n4020), .ZN(n4024) );
  NAND4_X2 U55248 ( .A1(n12680), .A2(n16015), .A3(n61281), .A4(n61280), .ZN(
        n14409) );
  NOR2_X2 U55256 ( .A1(n42485), .A2(n42493), .ZN(n61281) );
  NAND3_X2 U55277 ( .A1(n61284), .A2(n19100), .A3(n61283), .ZN(n46701) );
  OAI21_X1 U55297 ( .A1(n55371), .A2(n19973), .B(n61288), .ZN(n55376) );
  BUF_X2 U55300 ( .I(n9421), .Z(n61293) );
  XOR2_X1 U55304 ( .A1(n61294), .A2(n1835), .Z(n32348) );
  XOR2_X1 U55307 ( .A1(n23693), .A2(n32345), .Z(n61294) );
  NAND3_X1 U55327 ( .A1(n60415), .A2(n7932), .A3(n9648), .ZN(n20157) );
  XOR2_X1 U55353 ( .A1(n61295), .A2(n61418), .Z(n5028) );
  NOR2_X2 U55357 ( .A1(n2339), .A2(n2335), .ZN(n26131) );
  OAI21_X1 U55365 ( .A1(n61298), .A2(n61297), .B(n36569), .ZN(n20165) );
  NOR2_X1 U55389 ( .A1(n3809), .A2(n36563), .ZN(n61297) );
  NAND2_X2 U55398 ( .A1(n5054), .A2(n55099), .ZN(n55036) );
  XOR2_X1 U55421 ( .A1(n12815), .A2(n12814), .Z(n12811) );
  XOR2_X1 U55429 ( .A1(n25254), .A2(n9847), .Z(n61305) );
  NAND4_X2 U55486 ( .A1(n19295), .A2(n231), .A3(n19296), .A4(n40509), .ZN(
        n40511) );
  INV_X2 U55511 ( .I(n14306), .ZN(n61308) );
  NAND2_X2 U55540 ( .A1(n29188), .A2(n63007), .ZN(n2342) );
  NAND2_X2 U55541 ( .A1(n55286), .A2(n55474), .ZN(n55471) );
  NAND2_X2 U55545 ( .A1(n13128), .A2(n61310), .ZN(n19313) );
  AND2_X1 U55548 ( .A1(n13131), .A2(n13127), .Z(n61310) );
  NAND2_X2 U55568 ( .A1(n41831), .A2(n41293), .ZN(n42211) );
  AND2_X1 U55571 ( .A1(n48121), .A2(n48119), .Z(n61313) );
  OAI21_X1 U55575 ( .A1(n29531), .A2(n29532), .B(n29813), .ZN(n61315) );
  NAND2_X2 U55584 ( .A1(n47186), .A2(n19361), .ZN(n5705) );
  NAND2_X2 U55585 ( .A1(n1789), .A2(n34908), .ZN(n35435) );
  NOR2_X2 U55596 ( .A1(n35431), .A2(n22737), .ZN(n34908) );
  NAND4_X2 U55599 ( .A1(n42221), .A2(n42219), .A3(n42218), .A4(n42220), .ZN(
        n42222) );
  NAND2_X2 U55619 ( .A1(n40968), .A2(n40617), .ZN(n18827) );
  NAND2_X2 U55625 ( .A1(n5172), .A2(n56167), .ZN(n56158) );
  INV_X2 U55631 ( .I(n56190), .ZN(n56167) );
  OR2_X1 U55633 ( .A1(n30787), .A2(n29747), .Z(n29962) );
  XOR2_X1 U55639 ( .A1(n304), .A2(n61318), .Z(n18155) );
  XOR2_X1 U55640 ( .A1(n21369), .A2(n29410), .Z(n61318) );
  XOR2_X1 U55648 ( .A1(n45285), .A2(n16932), .Z(n61319) );
  NOR2_X1 U55671 ( .A1(n40998), .A2(n61005), .ZN(n40212) );
  BUF_X2 U55686 ( .I(n27568), .Z(n61320) );
  NOR2_X1 U55712 ( .A1(n63355), .A2(n9250), .ZN(n29250) );
  OAI21_X1 U55754 ( .A1(n61325), .A2(n61320), .B(n61324), .ZN(n26621) );
  AND2_X1 U55758 ( .A1(n8022), .A2(n26615), .Z(n61325) );
  NAND2_X2 U55763 ( .A1(n49432), .A2(n48907), .ZN(n61326) );
  INV_X4 U55781 ( .I(n5205), .ZN(n36955) );
  NAND3_X2 U55800 ( .A1(n35050), .A2(n35051), .A3(n35052), .ZN(n5205) );
  NAND2_X2 U55801 ( .A1(n54939), .A2(n52958), .ZN(n15281) );
  XOR2_X1 U55843 ( .A1(n24714), .A2(n24713), .Z(n51148) );
  NAND2_X2 U55914 ( .A1(n61334), .A2(n11672), .ZN(n22296) );
  NAND3_X2 U55933 ( .A1(n17162), .A2(n21501), .A3(n61337), .ZN(n24934) );
  OAI21_X1 U55935 ( .A1(n61761), .A2(n11353), .B(n61338), .ZN(n55110) );
  NOR2_X2 U55949 ( .A1(n31032), .A2(n31038), .ZN(n30141) );
  NAND2_X2 U55974 ( .A1(n26512), .A2(n26511), .ZN(n31556) );
  NAND2_X1 U56011 ( .A1(n33222), .A2(n33221), .ZN(n61349) );
  XOR2_X1 U56056 ( .A1(n51156), .A2(n51096), .Z(n61352) );
  INV_X2 U56072 ( .I(n61354), .ZN(n2670) );
  NAND4_X2 U56077 ( .A1(n23316), .A2(n48518), .A3(n48644), .A4(n48514), .ZN(
        n48630) );
  AND2_X1 U56088 ( .A1(n4784), .A2(n19196), .Z(n315) );
  NAND2_X1 U56090 ( .A1(n61356), .A2(n6706), .ZN(n7177) );
  NOR2_X2 U56120 ( .A1(n3888), .A2(n53845), .ZN(n53847) );
  NAND2_X2 U56136 ( .A1(n21059), .A2(n21878), .ZN(n34306) );
  XOR2_X1 U56143 ( .A1(n61360), .A2(n44585), .Z(n5027) );
  BUF_X2 U56169 ( .I(n7587), .Z(n61362) );
  NAND2_X1 U56170 ( .A1(n56428), .A2(n51899), .ZN(n51900) );
  XOR2_X1 U56223 ( .A1(n51812), .A2(n61364), .Z(n10352) );
  XOR2_X1 U56234 ( .A1(n50792), .A2(n50791), .Z(n61364) );
  INV_X2 U56264 ( .I(n61365), .ZN(n18490) );
  XOR2_X1 U56293 ( .A1(n3172), .A2(n1759), .Z(n5728) );
  NOR2_X1 U56299 ( .A1(n61366), .A2(n1848), .ZN(n21752) );
  NAND2_X1 U56303 ( .A1(n21626), .A2(n22014), .ZN(n61366) );
  NOR2_X2 U56325 ( .A1(n7062), .A2(n16174), .ZN(n23138) );
  BUF_X2 U56330 ( .I(n56441), .Z(n61368) );
  NAND2_X1 U56338 ( .A1(n5131), .A2(n47443), .ZN(n12455) );
  INV_X2 U56339 ( .I(n25150), .ZN(n51730) );
  AOI22_X1 U56350 ( .A1(n48997), .A2(n48998), .B1(n23656), .B2(n48999), .ZN(
        n24711) );
  BUF_X2 U56356 ( .I(n23928), .Z(n61372) );
  XOR2_X1 U56363 ( .A1(n51945), .A2(n61373), .Z(n50894) );
  XOR2_X1 U56380 ( .A1(n51229), .A2(n50889), .Z(n61373) );
  NOR2_X2 U56409 ( .A1(n15007), .A2(n18104), .ZN(n12694) );
  BUF_X2 U56423 ( .I(n31040), .Z(n61376) );
  BUF_X2 U56450 ( .I(Key[70]), .Z(n61380) );
  XOR2_X1 U56480 ( .A1(n25721), .A2(n10898), .Z(n3381) );
  BUF_X2 U56498 ( .I(n31074), .Z(n61382) );
  NAND3_X2 U56502 ( .A1(n61384), .A2(n29478), .A3(n29477), .ZN(n9166) );
  BUF_X4 U56522 ( .I(n56559), .Z(n23526) );
  XOR2_X1 U56533 ( .A1(n51616), .A2(n48725), .Z(n48753) );
  XOR2_X1 U56539 ( .A1(n10461), .A2(n55191), .Z(n51616) );
  NOR2_X1 U56541 ( .A1(n61389), .A2(n21785), .ZN(n21784) );
  NOR2_X1 U56552 ( .A1(n61750), .A2(n30360), .ZN(n61390) );
  NOR3_X1 U56556 ( .A1(n2846), .A2(n1842), .A3(n62670), .ZN(n61391) );
  NAND2_X2 U56567 ( .A1(n11642), .A2(n11640), .ZN(n49004) );
  OAI22_X2 U56571 ( .A1(n64080), .A2(n41543), .B1(n9211), .B2(n64724), .ZN(
        n61395) );
  NOR2_X1 U56574 ( .A1(n41940), .A2(n41941), .ZN(n61398) );
  NOR2_X2 U56584 ( .A1(n28244), .A2(n26270), .ZN(n28241) );
  NAND2_X1 U56586 ( .A1(n61399), .A2(n29109), .ZN(n2138) );
  NAND2_X1 U56588 ( .A1(n27372), .A2(n27371), .ZN(n61399) );
  XOR2_X1 U56595 ( .A1(n61400), .A2(n54517), .Z(Plaintext[72]) );
  XOR2_X1 U56596 ( .A1(n32706), .A2(n61401), .Z(n52366) );
  XOR2_X1 U56599 ( .A1(n38850), .A2(n31661), .Z(n32706) );
  XOR2_X1 U56618 ( .A1(n31667), .A2(n61403), .Z(n61402) );
  XOR2_X1 U56620 ( .A1(n12379), .A2(n2000), .Z(n1999) );
  XOR2_X1 U56633 ( .A1(n7082), .A2(n13553), .Z(n7439) );
  XOR2_X1 U56645 ( .A1(n1681), .A2(n44384), .Z(n12712) );
  XOR2_X1 U56646 ( .A1(n51662), .A2(n18485), .Z(n22056) );
  XOR2_X1 U56649 ( .A1(n61409), .A2(n33891), .Z(n30573) );
  XOR2_X1 U56651 ( .A1(n30571), .A2(n21531), .Z(n61409) );
  NAND2_X1 U56665 ( .A1(n61416), .A2(n61414), .ZN(n53044) );
  INV_X1 U56667 ( .I(n9161), .ZN(n61415) );
  NAND2_X1 U56683 ( .A1(n53017), .A2(n9161), .ZN(n61416) );
  XOR2_X1 U56684 ( .A1(n38779), .A2(n10703), .Z(n61418) );
  AND2_X1 U56686 ( .A1(n53413), .A2(n53412), .Z(n61419) );
  NOR2_X1 U56687 ( .A1(n16500), .A2(n52493), .ZN(n25720) );
  NOR2_X1 U56701 ( .A1(n6077), .A2(n6078), .ZN(n6076) );
  NOR2_X1 U56709 ( .A1(n14574), .A2(n46748), .ZN(n14573) );
  NOR2_X1 U56718 ( .A1(n25197), .A2(n61420), .ZN(n10119) );
  NOR2_X1 U56729 ( .A1(n6344), .A2(n25175), .ZN(n61420) );
  NOR2_X2 U56731 ( .A1(n23572), .A2(n32913), .ZN(n38835) );
  NAND2_X2 U56738 ( .A1(n13743), .A2(n54102), .ZN(n53545) );
  OR3_X1 U56746 ( .A1(n35952), .A2(n62041), .A3(n20020), .Z(n32910) );
  AOI21_X1 U56747 ( .A1(n55269), .A2(n55270), .B(n55268), .ZN(n55273) );
  OAI22_X1 U56758 ( .A1(n27230), .A2(n25090), .B1(n27231), .B2(n27543), .ZN(
        n27235) );
  XOR2_X1 U56760 ( .A1(n61424), .A2(n18362), .Z(n11539) );
  OAI21_X1 U56767 ( .A1(n11176), .A2(n11683), .B(n24404), .ZN(n11682) );
  BUF_X2 U56768 ( .I(n24000), .Z(n61426) );
  XOR2_X1 U56789 ( .A1(n51504), .A2(n7111), .Z(n5666) );
  NAND3_X2 U56790 ( .A1(n15467), .A2(n5657), .A3(n15473), .ZN(n7111) );
  NAND4_X2 U56791 ( .A1(n56276), .A2(n4746), .A3(n56275), .A4(n56274), .ZN(
        n56323) );
  NAND2_X1 U56793 ( .A1(n54086), .A2(n54085), .ZN(n21005) );
  NAND3_X1 U56795 ( .A1(n38354), .A2(n38355), .A3(n403), .ZN(n61429) );
  NAND2_X1 U56797 ( .A1(n22676), .A2(n51260), .ZN(n7190) );
  NAND2_X1 U56798 ( .A1(n3262), .A2(n14201), .ZN(n3261) );
  XOR2_X1 U56801 ( .A1(n9200), .A2(n42026), .Z(n42029) );
  NOR2_X2 U56802 ( .A1(n2036), .A2(n18468), .ZN(n5431) );
  INV_X2 U56803 ( .I(n61432), .ZN(n61697) );
  NAND2_X2 U56805 ( .A1(n13900), .A2(n61433), .ZN(n14934) );
  OAI22_X1 U56806 ( .A1(n57175), .A2(n61434), .B1(n12734), .B2(n12733), .ZN(
        n12731) );
  NAND2_X1 U56807 ( .A1(n59577), .A2(n61435), .ZN(n61434) );
  INV_X2 U56808 ( .I(n13756), .ZN(n61435) );
  XOR2_X1 U56809 ( .A1(n15155), .A2(n14867), .Z(n16439) );
  NAND2_X2 U56810 ( .A1(n16040), .A2(n16440), .ZN(n14867) );
  NOR2_X2 U56811 ( .A1(n22768), .A2(n28533), .ZN(n28540) );
  NAND2_X1 U56812 ( .A1(n28541), .A2(n22768), .ZN(n61439) );
  NAND2_X1 U56813 ( .A1(n28544), .A2(n28543), .ZN(n61440) );
  AND2_X1 U56814 ( .A1(n14915), .A2(n2699), .Z(n34862) );
  XOR2_X1 U56815 ( .A1(n31199), .A2(n61441), .Z(n3757) );
  OR2_X1 U56816 ( .A1(n56587), .A2(n56592), .Z(n10168) );
  XOR2_X1 U56818 ( .A1(n51140), .A2(n51139), .Z(n51199) );
  NOR2_X2 U56819 ( .A1(n23353), .A2(n16254), .ZN(n1528) );
  INV_X2 U56820 ( .I(n61444), .ZN(n6996) );
  XOR2_X1 U56821 ( .A1(n6998), .A2(n6997), .Z(n61444) );
  XOR2_X1 U56823 ( .A1(n46650), .A2(n57394), .Z(n61445) );
  XOR2_X1 U56824 ( .A1(n59395), .A2(n61446), .Z(n1035) );
  XOR2_X1 U56825 ( .A1(n12507), .A2(n45850), .Z(n61446) );
  XOR2_X1 U56826 ( .A1(n10645), .A2(n31774), .Z(n3274) );
  NOR4_X2 U56827 ( .A1(n45188), .A2(n45186), .A3(n45187), .A4(n45185), .ZN(
        n45189) );
  XOR2_X1 U56828 ( .A1(n49126), .A2(n26022), .Z(n6694) );
  BUF_X2 U56830 ( .I(n25657), .Z(n61449) );
  AOI22_X1 U56840 ( .A1(n57134), .A2(n57133), .B1(n57135), .B2(n25145), .ZN(
        n57140) );
  XOR2_X1 U56844 ( .A1(n44119), .A2(n44118), .Z(n46346) );
  XOR2_X1 U56845 ( .A1(n112), .A2(n24255), .Z(n24432) );
  XOR2_X1 U56846 ( .A1(n31764), .A2(n24225), .Z(n24254) );
  NAND4_X2 U56847 ( .A1(n19735), .A2(n53303), .A3(n4283), .A4(n9481), .ZN(
        n53251) );
  NOR2_X1 U56848 ( .A1(n18113), .A2(n26661), .ZN(n18112) );
  XOR2_X1 U56849 ( .A1(n61461), .A2(n39626), .Z(n3069) );
  XOR2_X1 U56850 ( .A1(n38648), .A2(n38283), .Z(n61461) );
  OR2_X1 U56853 ( .A1(n12378), .A2(n42608), .Z(n61465) );
  NAND2_X2 U56854 ( .A1(n42031), .A2(n42027), .ZN(n41794) );
  XOR2_X1 U56856 ( .A1(n32385), .A2(n32515), .Z(n23287) );
  XOR2_X1 U56857 ( .A1(n61467), .A2(n65268), .Z(n9971) );
  XOR2_X1 U56858 ( .A1(n12055), .A2(n13584), .Z(n61467) );
  XOR2_X1 U56859 ( .A1(n39259), .A2(n57223), .Z(n61468) );
  INV_X1 U56861 ( .I(n26346), .ZN(n61470) );
  AOI21_X1 U56864 ( .A1(n47375), .A2(n61474), .B(n61473), .ZN(n47383) );
  AND2_X1 U56865 ( .A1(n47373), .A2(n10475), .Z(n61473) );
  NAND2_X1 U56866 ( .A1(n47372), .A2(n47371), .ZN(n61474) );
  NOR2_X1 U56868 ( .A1(n48314), .A2(n19003), .ZN(n48310) );
  NOR3_X1 U56869 ( .A1(n14326), .A2(n61476), .A3(n25107), .ZN(n16771) );
  XOR2_X1 U56871 ( .A1(n32516), .A2(n32387), .Z(n25165) );
  XOR2_X1 U56872 ( .A1(n38716), .A2(n18809), .Z(n20412) );
  XOR2_X1 U56873 ( .A1(n61478), .A2(n37887), .Z(n22242) );
  NAND3_X1 U56875 ( .A1(n61479), .A2(n14051), .A3(n43039), .ZN(n41581) );
  NAND3_X1 U56876 ( .A1(n43043), .A2(n41584), .A3(n24405), .ZN(n61479) );
  XOR2_X1 U56877 ( .A1(n31421), .A2(n22237), .Z(n12977) );
  XOR2_X1 U56878 ( .A1(n19094), .A2(n19093), .Z(n31421) );
  XOR2_X1 U56882 ( .A1(n9109), .A2(n9108), .Z(n32620) );
  NAND2_X2 U56883 ( .A1(n64994), .A2(n27485), .ZN(n26936) );
  NOR3_X2 U56885 ( .A1(n689), .A2(n2123), .A3(n29114), .ZN(n29203) );
  NAND3_X2 U56886 ( .A1(n13795), .A2(n13790), .A3(n16008), .ZN(n54191) );
  NAND3_X1 U56887 ( .A1(n8089), .A2(n28433), .A3(n8088), .ZN(n7219) );
  OR3_X1 U56888 ( .A1(n5765), .A2(n5764), .A3(n5763), .Z(n219) );
  NOR2_X2 U56890 ( .A1(n36623), .A2(n13358), .ZN(n36960) );
  BUF_X2 U56892 ( .I(n26391), .Z(n61491) );
  NAND2_X2 U56894 ( .A1(n61749), .A2(n5147), .ZN(n33972) );
  XOR2_X1 U56895 ( .A1(n22015), .A2(n306), .Z(n11440) );
  NAND2_X2 U56899 ( .A1(n30708), .A2(n23072), .ZN(n30142) );
  NOR2_X2 U56900 ( .A1(n30702), .A2(n1315), .ZN(n30708) );
  NOR2_X2 U56901 ( .A1(n27808), .A2(n1970), .ZN(n11065) );
  NAND2_X2 U56902 ( .A1(n28625), .A2(n22648), .ZN(n27808) );
  XOR2_X1 U56904 ( .A1(n39758), .A2(n39441), .Z(n16983) );
  XOR2_X1 U56906 ( .A1(n20113), .A2(n46694), .Z(n2274) );
  AOI21_X2 U56907 ( .A1(n9720), .A2(n61501), .B(n61500), .ZN(n61499) );
  NAND2_X2 U56908 ( .A1(n6195), .A2(n39909), .ZN(n22084) );
  OR2_X1 U56909 ( .A1(n55088), .A2(n22362), .Z(n55077) );
  NAND2_X2 U56910 ( .A1(n11912), .A2(n22550), .ZN(n54807) );
  NOR2_X1 U56915 ( .A1(n6984), .A2(n8223), .ZN(n35913) );
  INV_X4 U56916 ( .I(n16491), .ZN(n1353) );
  OR2_X1 U56917 ( .A1(n1146), .A2(n24192), .Z(n54623) );
  NAND2_X2 U56919 ( .A1(n38612), .A2(n38611), .ZN(n23702) );
  BUF_X2 U56920 ( .I(n19418), .Z(n61506) );
  XOR2_X1 U56921 ( .A1(n50869), .A2(n61508), .Z(n61507) );
  NOR2_X1 U56923 ( .A1(n35983), .A2(n61180), .ZN(n61511) );
  OAI22_X1 U56924 ( .A1(n53420), .A2(n53421), .B1(n53422), .B2(n53862), .ZN(
        n53423) );
  NAND2_X2 U56925 ( .A1(n53018), .A2(n4480), .ZN(n53420) );
  NAND2_X1 U56926 ( .A1(n12157), .A2(n53159), .ZN(n53172) );
  OAI21_X1 U56927 ( .A1(n54960), .A2(n55094), .B(n61512), .ZN(n55105) );
  NOR2_X1 U56928 ( .A1(n23307), .A2(n680), .ZN(n61512) );
  NAND2_X2 U56931 ( .A1(n7273), .A2(n59681), .ZN(n33695) );
  NOR2_X2 U56934 ( .A1(n22444), .A2(n31189), .ZN(n27886) );
  NAND3_X2 U56935 ( .A1(n23624), .A2(n52823), .A3(n52824), .ZN(n52826) );
  NAND2_X2 U56938 ( .A1(n8348), .A2(n61520), .ZN(n7955) );
  NOR2_X2 U56939 ( .A1(n54874), .A2(n54871), .ZN(n61520) );
  XOR2_X1 U56940 ( .A1(n24343), .A2(n24342), .Z(n8165) );
  NAND2_X2 U56942 ( .A1(n42810), .A2(n7386), .ZN(n15278) );
  AOI22_X1 U56944 ( .A1(n1282), .A2(n9424), .B1(n55388), .B2(n23554), .ZN(
        n61521) );
  OR2_X1 U56951 ( .A1(n41472), .A2(n61526), .Z(n41477) );
  NAND2_X2 U56952 ( .A1(n40748), .A2(n40755), .ZN(n41472) );
  NAND2_X1 U56953 ( .A1(n21211), .A2(n21212), .ZN(n14584) );
  AOI22_X2 U56954 ( .A1(n42657), .A2(n42658), .B1(n8052), .B2(n8053), .ZN(
        n21211) );
  OR2_X1 U56955 ( .A1(n47161), .A2(n47160), .Z(n13526) );
  XOR2_X1 U56956 ( .A1(n12608), .A2(n44991), .Z(n44992) );
  OR3_X1 U56957 ( .A1(n45984), .A2(n47621), .A3(n61527), .Z(n47246) );
  BUF_X2 U56958 ( .I(n56990), .Z(n61528) );
  BUF_X2 U56960 ( .I(n19489), .Z(n61530) );
  NOR2_X1 U56961 ( .A1(n22506), .A2(n21428), .ZN(n23245) );
  INV_X1 U56962 ( .I(n30724), .ZN(n61534) );
  NAND2_X1 U56963 ( .A1(n61536), .A2(n30724), .ZN(n61535) );
  NAND2_X1 U56964 ( .A1(n64538), .A2(n29215), .ZN(n61536) );
  INV_X2 U56968 ( .I(n45229), .ZN(n6314) );
  XOR2_X1 U56970 ( .A1(n39272), .A2(n38744), .Z(n715) );
  XOR2_X1 U56971 ( .A1(n23175), .A2(n23962), .Z(n38744) );
  XOR2_X1 U56972 ( .A1(n61545), .A2(n886), .Z(n5745) );
  XOR2_X1 U56973 ( .A1(n33190), .A2(n5747), .Z(n61545) );
  BUF_X2 U56974 ( .I(n35318), .Z(n61547) );
  XOR2_X1 U56975 ( .A1(n61548), .A2(n31890), .Z(n31892) );
  XOR2_X1 U56976 ( .A1(n23096), .A2(n14818), .Z(n61548) );
  OAI21_X1 U56977 ( .A1(n30740), .A2(n31201), .B(n18872), .ZN(n61549) );
  BUF_X2 U56978 ( .I(n38126), .Z(n61550) );
  NAND2_X2 U56979 ( .A1(n5903), .A2(n34634), .ZN(n34639) );
  NOR4_X2 U56980 ( .A1(n22150), .A2(n61552), .A3(n19131), .A4(n61551), .ZN(
        n15097) );
  XOR2_X1 U56983 ( .A1(n52584), .A2(n52583), .Z(n15914) );
  NAND3_X2 U56985 ( .A1(n28053), .A2(n27141), .A3(n27142), .ZN(n28324) );
  NAND3_X2 U56986 ( .A1(n25287), .A2(n40606), .A3(n37533), .ZN(n61555) );
  NAND2_X1 U56987 ( .A1(n54573), .A2(n54574), .ZN(n61556) );
  NAND3_X1 U56988 ( .A1(n41925), .A2(n41926), .A3(n11316), .ZN(n61557) );
  NAND2_X1 U56991 ( .A1(n22885), .A2(n53616), .ZN(n61558) );
  OR2_X1 U56992 ( .A1(n12360), .A2(n47296), .Z(n45931) );
  INV_X2 U56993 ( .I(n19595), .ZN(n61563) );
  NOR2_X2 U56995 ( .A1(n48460), .A2(n20897), .ZN(n47209) );
  OAI21_X2 U57002 ( .A1(n3289), .A2(n8870), .B(n47085), .ZN(n3288) );
  NAND3_X1 U57004 ( .A1(n4008), .A2(n36548), .A3(n22454), .ZN(n61566) );
  XOR2_X1 U57005 ( .A1(n51975), .A2(n8144), .Z(n17704) );
  XOR2_X1 U57006 ( .A1(n17705), .A2(n50976), .Z(n51975) );
  NAND2_X2 U57007 ( .A1(n1990), .A2(n31169), .ZN(n33283) );
  XOR2_X1 U57008 ( .A1(n20470), .A2(n9922), .Z(n61569) );
  XOR2_X1 U57011 ( .A1(n23818), .A2(n24030), .Z(n61573) );
  NAND3_X2 U57013 ( .A1(n15513), .A2(n1032), .A3(n4096), .ZN(n43852) );
  XOR2_X1 U57014 ( .A1(n8868), .A2(n65058), .Z(n45860) );
  XOR2_X1 U57015 ( .A1(n33291), .A2(n61575), .Z(n33293) );
  NOR2_X2 U57016 ( .A1(n2078), .A2(n61576), .ZN(n9230) );
  NAND2_X1 U57018 ( .A1(n17837), .A2(n17753), .ZN(n17836) );
  XOR2_X1 U57019 ( .A1(n51932), .A2(n2604), .Z(n52058) );
  AND2_X1 U57020 ( .A1(n64145), .A2(n11977), .Z(n4718) );
  NAND2_X2 U57023 ( .A1(n8097), .A2(n10240), .ZN(n30341) );
  NOR2_X2 U57024 ( .A1(n28481), .A2(n61581), .ZN(n25669) );
  XOR2_X1 U57027 ( .A1(n61583), .A2(n18656), .Z(n11305) );
  XOR2_X1 U57028 ( .A1(n37980), .A2(n37986), .Z(n61583) );
  XOR2_X1 U57029 ( .A1(n50850), .A2(n24074), .Z(n51418) );
  XOR2_X1 U57030 ( .A1(n50938), .A2(n51671), .Z(n50850) );
  NAND2_X2 U57031 ( .A1(n21791), .A2(n41213), .ZN(n22525) );
  INV_X2 U57032 ( .I(n61584), .ZN(n14312) );
  XOR2_X1 U57033 ( .A1(Ciphertext[171]), .A2(Key[130]), .Z(n61584) );
  OR2_X2 U57034 ( .A1(n24889), .A2(n15789), .Z(n12423) );
  NOR2_X2 U57038 ( .A1(n36955), .A2(n36959), .ZN(n5900) );
  XOR2_X1 U57043 ( .A1(n17932), .A2(n17933), .Z(n19362) );
  AOI21_X2 U57045 ( .A1(n40908), .A2(n43014), .B(n41679), .ZN(n43021) );
  NOR2_X2 U57046 ( .A1(n41684), .A2(n41996), .ZN(n41679) );
  NAND2_X1 U57047 ( .A1(n2829), .A2(n2833), .ZN(n4842) );
  XOR2_X1 U57050 ( .A1(n61591), .A2(n5957), .Z(n61590) );
  XOR2_X1 U57051 ( .A1(n39653), .A2(n61592), .Z(n17448) );
  XOR2_X1 U57052 ( .A1(n24169), .A2(n12356), .Z(n61592) );
  NAND2_X1 U57053 ( .A1(n43164), .A2(n4789), .ZN(n61595) );
  NAND2_X2 U57054 ( .A1(n61596), .A2(n16466), .ZN(n40651) );
  NOR3_X2 U57055 ( .A1(n61597), .A2(n16465), .A3(n16464), .ZN(n61596) );
  NAND2_X2 U57058 ( .A1(n1233), .A2(n59538), .ZN(n55076) );
  XOR2_X1 U57060 ( .A1(n191), .A2(n44046), .Z(n850) );
  XOR2_X1 U57061 ( .A1(n61602), .A2(n4561), .Z(Plaintext[93]) );
  XOR2_X1 U57063 ( .A1(n8214), .A2(n22512), .Z(n61603) );
  XOR2_X1 U57064 ( .A1(n51318), .A2(n21757), .Z(n21756) );
  XOR2_X1 U57065 ( .A1(n51202), .A2(n51201), .Z(n51318) );
  NOR2_X1 U57066 ( .A1(n61605), .A2(n61604), .ZN(n56712) );
  NOR2_X1 U57067 ( .A1(n56738), .A2(n56736), .ZN(n61604) );
  NOR2_X1 U57068 ( .A1(n56707), .A2(n56708), .ZN(n61605) );
  INV_X2 U57069 ( .I(n7738), .ZN(n49498) );
  OR2_X1 U57071 ( .A1(n5389), .A2(n17866), .Z(n17865) );
  NAND4_X2 U57072 ( .A1(n34206), .A2(n34207), .A3(n36705), .A4(n14719), .ZN(
        n38510) );
  AOI21_X2 U57076 ( .A1(n33459), .A2(n22993), .B(n61608), .ZN(n24306) );
  OAI22_X2 U57077 ( .A1(n130), .A2(n34908), .B1(n36940), .B2(n34907), .ZN(
        n61608) );
  XOR2_X1 U57079 ( .A1(n57331), .A2(n61611), .Z(n61656) );
  XOR2_X1 U57080 ( .A1(n5363), .A2(n23019), .Z(n61611) );
  NAND3_X2 U57081 ( .A1(n18610), .A2(n15915), .A3(n61712), .ZN(n16914) );
  INV_X2 U57082 ( .I(n63261), .ZN(n18600) );
  NAND2_X2 U57085 ( .A1(n61617), .A2(n14940), .ZN(n31261) );
  NAND4_X2 U57086 ( .A1(n61619), .A2(n37938), .A3(n37936), .A4(n37937), .ZN(
        n38056) );
  INV_X2 U57087 ( .I(n8380), .ZN(n13925) );
  XOR2_X1 U57090 ( .A1(n39439), .A2(n16250), .Z(n11802) );
  XOR2_X1 U57092 ( .A1(n22146), .A2(n18838), .Z(n32564) );
  XOR2_X1 U57093 ( .A1(n32733), .A2(n23491), .Z(n32207) );
  BUF_X2 U57100 ( .I(n17411), .Z(n61622) );
  INV_X2 U57101 ( .I(n61623), .ZN(n2295) );
  XOR2_X1 U57102 ( .A1(Ciphertext[57]), .A2(Key[100]), .Z(n61623) );
  NOR3_X2 U57103 ( .A1(n10976), .A2(n10975), .A3(n61625), .ZN(n10973) );
  XOR2_X1 U57104 ( .A1(n15615), .A2(n39372), .Z(n15081) );
  BUF_X2 U57105 ( .I(n47902), .Z(n61628) );
  XOR2_X1 U57109 ( .A1(n14827), .A2(n14828), .Z(n4405) );
  XOR2_X1 U57110 ( .A1(n61632), .A2(n45035), .Z(n24689) );
  XOR2_X1 U57111 ( .A1(n61), .A2(n44848), .Z(n61632) );
  XOR2_X1 U57112 ( .A1(n61633), .A2(n33079), .Z(n57) );
  XOR2_X1 U57113 ( .A1(n33077), .A2(n33076), .Z(n61633) );
  XOR2_X1 U57114 ( .A1(n3184), .A2(n3185), .Z(n3183) );
  XOR2_X1 U57116 ( .A1(n31810), .A2(n31438), .Z(n61634) );
  NOR3_X2 U57120 ( .A1(n41247), .A2(n42684), .A3(n42829), .ZN(n45835) );
  XOR2_X1 U57122 ( .A1(n18054), .A2(n38990), .Z(n39696) );
  BUF_X2 U57124 ( .I(n41384), .Z(n61638) );
  XOR2_X1 U57128 ( .A1(n38622), .A2(n13705), .Z(n8542) );
  XOR2_X1 U57130 ( .A1(n61640), .A2(n31839), .Z(n6127) );
  XOR2_X1 U57131 ( .A1(n44274), .A2(n32636), .Z(n61640) );
  XOR2_X1 U57133 ( .A1(n32284), .A2(n61641), .Z(n7937) );
  NOR2_X1 U57134 ( .A1(n2301), .A2(n3651), .ZN(n61642) );
  NAND2_X2 U57135 ( .A1(n14451), .A2(n24420), .ZN(n19679) );
  INV_X1 U57136 ( .I(n2246), .ZN(n49527) );
  AND2_X2 U57137 ( .A1(n18004), .A2(n6589), .Z(n61643) );
  NAND3_X1 U57138 ( .A1(n58560), .A2(n23315), .A3(n25978), .ZN(n61644) );
  INV_X2 U57139 ( .I(n24571), .ZN(n35240) );
  XNOR2_X1 U57141 ( .A1(n12682), .A2(n31678), .ZN(n61646) );
  NAND2_X2 U57142 ( .A1(n24522), .A2(n2033), .ZN(n34989) );
  INV_X4 U57143 ( .I(n81), .ZN(n36070) );
  OR2_X1 U57144 ( .A1(n33763), .A2(n2721), .Z(n61648) );
  INV_X1 U57145 ( .I(n25571), .ZN(n35908) );
  OR2_X2 U57146 ( .A1(n15243), .A2(n62514), .Z(n25571) );
  XNOR2_X1 U57147 ( .A1(n38364), .A2(n37840), .ZN(n61650) );
  XNOR2_X1 U57148 ( .A1(n7713), .A2(n37706), .ZN(n61651) );
  NAND2_X2 U57150 ( .A1(n25008), .A2(n34471), .ZN(n38796) );
  XNOR2_X1 U57153 ( .A1(n38731), .A2(n21722), .ZN(n61654) );
  INV_X2 U57154 ( .I(n24976), .ZN(n38672) );
  INV_X1 U57156 ( .I(n41257), .ZN(n41256) );
  XNOR2_X1 U57157 ( .A1(n21016), .A2(n39547), .ZN(n61655) );
  INV_X2 U57158 ( .I(n9711), .ZN(n5775) );
  XOR2_X1 U57159 ( .A1(n63730), .A2(n38706), .Z(n61657) );
  INV_X2 U57160 ( .I(n24645), .ZN(n3566) );
  OR2_X2 U57161 ( .A1(n9872), .A2(n13383), .Z(n42450) );
  INV_X2 U57162 ( .I(n3178), .ZN(n25118) );
  NAND2_X2 U57165 ( .A1(n38272), .A2(n38271), .ZN(n43874) );
  AND3_X1 U57166 ( .A1(n21206), .A2(n19256), .A3(n16497), .Z(n61660) );
  INV_X4 U57167 ( .I(n19946), .ZN(n42324) );
  XNOR2_X1 U57168 ( .A1(n43906), .A2(n43008), .ZN(n61661) );
  XNOR2_X1 U57169 ( .A1(n22639), .A2(n46162), .ZN(n61663) );
  BUF_X4 U57172 ( .I(n42846), .Z(n15007) );
  XOR2_X1 U57174 ( .A1(n25695), .A2(n23073), .Z(n61665) );
  INV_X2 U57175 ( .I(n11595), .ZN(n23548) );
  XNOR2_X1 U57176 ( .A1(n25835), .A2(n25833), .ZN(n61666) );
  XOR2_X1 U57177 ( .A1(n16242), .A2(n6171), .Z(n61667) );
  XNOR2_X1 U57178 ( .A1(n63005), .A2(n46665), .ZN(n61669) );
  AND2_X1 U57179 ( .A1(n13801), .A2(n10891), .Z(n61670) );
  XNOR2_X1 U57180 ( .A1(n13853), .A2(n44336), .ZN(n61671) );
  XNOR2_X1 U57183 ( .A1(n5897), .A2(n12712), .ZN(n61672) );
  CLKBUF_X8 U57184 ( .I(n5945), .Z(n1205) );
  INV_X4 U57185 ( .I(n25598), .ZN(n2810) );
  INV_X1 U57186 ( .I(n376), .ZN(n48317) );
  INV_X2 U57187 ( .I(n50096), .ZN(n3031) );
  OR3_X1 U57188 ( .A1(n1633), .A2(n49287), .A3(n49283), .Z(n61674) );
  OR3_X1 U57189 ( .A1(n48082), .A2(n48076), .A3(n15823), .Z(n61675) );
  OR2_X1 U57190 ( .A1(n18565), .A2(n8380), .Z(n61676) );
  AND2_X1 U57191 ( .A1(n48332), .A2(n49910), .Z(n61678) );
  AND4_X1 U57192 ( .A1(n49725), .A2(n12580), .A3(n5282), .A4(n12579), .Z(
        n61679) );
  INV_X2 U57193 ( .I(n13944), .ZN(n6363) );
  INV_X4 U57194 ( .I(n25233), .ZN(n18608) );
  INV_X4 U57195 ( .I(n8228), .ZN(n51572) );
  NAND2_X2 U57196 ( .A1(n18084), .A2(n18083), .ZN(n2222) );
  INV_X2 U57198 ( .I(n56559), .ZN(n24696) );
  INV_X2 U57200 ( .I(n5119), .ZN(n22550) );
  AND3_X1 U57201 ( .A1(n54317), .A2(n1610), .A3(n22372), .Z(n61683) );
  INV_X2 U57202 ( .I(n25267), .ZN(n9161) );
  INV_X2 U57203 ( .I(n54110), .ZN(n53871) );
  OR3_X1 U57204 ( .A1(n18255), .A2(n4943), .A3(n25167), .Z(n61684) );
  AND3_X1 U57205 ( .A1(n56987), .A2(n52683), .A3(n61902), .Z(n61685) );
  AND3_X1 U57206 ( .A1(n53216), .A2(n53215), .A3(n1612), .Z(n61686) );
  AND2_X2 U57207 ( .A1(n14934), .A2(n21830), .Z(n61687) );
  INV_X4 U57210 ( .I(n53997), .ZN(n6168) );
  OR2_X2 U57212 ( .A1(n6873), .A2(n58843), .Z(n5227) );
  INV_X2 U57213 ( .I(n23646), .ZN(n5551) );
  AND2_X1 U57214 ( .A1(n19817), .A2(n14927), .Z(n61691) );
  AND2_X1 U57216 ( .A1(n62074), .A2(n22775), .Z(n61694) );
  AND3_X1 U57217 ( .A1(n54004), .A2(n54003), .A3(n54002), .Z(n61695) );
  AND3_X1 U57218 ( .A1(n53792), .A2(n53813), .A3(n53791), .Z(n61696) );
  NAND2_X2 U21061 ( .A1(n22042), .A2(n22533), .ZN(n20204) );
  INV_X2 U2837 ( .I(n11620), .ZN(n24698) );
  INV_X4 U16278 ( .I(n48103), .ZN(n13838) );
  BUF_X4 U36256 ( .I(n30196), .Z(n59798) );
  INV_X2 U12886 ( .I(n27139), .ZN(n57872) );
  NOR2_X2 U3020 ( .A1(n30085), .A2(n23370), .ZN(n30071) );
  NAND2_X2 U6129 ( .A1(n9392), .A2(n5070), .ZN(n28898) );
  INV_X2 U2122 ( .I(n38072), .ZN(n17817) );
  NOR2_X2 U23597 ( .A1(n22023), .A2(n61300), .ZN(n61299) );
  NAND2_X2 U7245 ( .A1(n48644), .A2(n26226), .ZN(n12993) );
  INV_X2 U2301 ( .I(n36538), .ZN(n36384) );
  INV_X4 U1162 ( .I(n826), .ZN(n49948) );
  NAND2_X2 U7367 ( .A1(n56150), .A2(n17606), .ZN(n56149) );
  NOR2_X2 U23849 ( .A1(n36821), .A2(n1235), .ZN(n36829) );
  NAND2_X2 U21137 ( .A1(n2790), .A2(n26347), .ZN(n28417) );
  INV_X2 U4394 ( .I(n42639), .ZN(n43504) );
  OAI22_X2 U2835 ( .A1(n3311), .A2(n28796), .B1(n3310), .B2(n58440), .ZN(
        n31063) );
  NAND3_X2 U35263 ( .A1(n1530), .A2(n60694), .A3(n1781), .ZN(n35053) );
  BUF_X2 U7674 ( .I(n41147), .Z(n60077) );
  INV_X2 U8265 ( .I(n11477), .ZN(n34559) );
  INV_X2 U4323 ( .I(n39066), .ZN(n25397) );
  INV_X2 U20491 ( .I(n6306), .ZN(n18809) );
  NOR2_X2 U5309 ( .A1(n26823), .A2(n26898), .ZN(n26903) );
  NOR2_X2 U3144 ( .A1(n1530), .A2(n36965), .ZN(n35450) );
  INV_X4 U8574 ( .I(n16766), .ZN(n1262) );
  AOI22_X2 U10074 ( .A1(n39018), .A2(n39017), .B1(n64493), .B2(n39016), .ZN(
        n8315) );
  OR2_X2 U206 ( .A1(n19980), .A2(n19981), .Z(n58828) );
  NOR2_X2 U3391 ( .A1(n16446), .A2(n16667), .ZN(n23039) );
  NAND2_X2 U9736 ( .A1(n26823), .A2(n63094), .ZN(n27833) );
  INV_X4 U15111 ( .I(n50576), .ZN(n22747) );
  INV_X2 U12885 ( .I(n10128), .ZN(n1491) );
  INV_X2 U1058 ( .I(n19558), .ZN(n48238) );
  INV_X2 U3085 ( .I(n31261), .ZN(n23269) );
  INV_X2 U34332 ( .I(n45386), .ZN(n16518) );
  INV_X2 U1213 ( .I(n24047), .ZN(n46025) );
  INV_X2 U484 ( .I(n54465), .ZN(n54088) );
  INV_X2 U215 ( .I(n56687), .ZN(n56733) );
  NAND2_X2 U65 ( .A1(n55074), .A2(n4087), .ZN(n55041) );
  OAI21_X2 U23216 ( .A1(n7260), .A2(n22875), .B(n57012), .ZN(n4396) );
  BUF_X4 U4361 ( .I(n900), .Z(n7883) );
  NAND2_X2 U50190 ( .A1(n59427), .A2(n39102), .ZN(n39103) );
  OAI21_X2 U19027 ( .A1(n30672), .A2(n30671), .B(n30670), .ZN(n30673) );
  INV_X2 U14954 ( .I(n38903), .ZN(n7256) );
  INV_X2 U3539 ( .I(n48930), .ZN(n44791) );
  BUF_X2 U16264 ( .I(n8794), .Z(n10621) );
  BUF_X2 U10403 ( .I(n32669), .Z(n8186) );
  INV_X2 U30887 ( .I(n10459), .ZN(n45889) );
  INV_X2 U8734 ( .I(n40400), .ZN(n41415) );
  BUF_X4 U44531 ( .I(Key[42]), .Z(n53772) );
  INV_X4 U27527 ( .I(n42681), .ZN(n42672) );
  AND2_X2 U2297 ( .A1(n4893), .A2(n2116), .Z(n798) );
  NAND2_X2 U4171 ( .A1(n15157), .A2(n838), .ZN(n14741) );
  INV_X2 U5368 ( .I(n18748), .ZN(n21985) );
  INV_X2 U43400 ( .I(n5193), .ZN(n56185) );
  INV_X2 U1595 ( .I(n15705), .ZN(n1214) );
  NOR2_X2 U2313 ( .A1(n321), .A2(n14556), .ZN(n40287) );
  OAI22_X2 U10817 ( .A1(n9294), .A2(n49505), .B1(n49503), .B2(n49504), .ZN(
        n9293) );
  INV_X4 U1675 ( .I(n7202), .ZN(n44480) );
  NOR2_X2 U1988 ( .A1(n16962), .A2(n4581), .ZN(n40329) );
  INV_X2 U28216 ( .I(n26060), .ZN(n51960) );
  INV_X4 U1615 ( .I(n42404), .ZN(n42076) );
  BUF_X4 U6696 ( .I(n34308), .Z(n23366) );
  NAND2_X2 U667 ( .A1(n3347), .A2(n20199), .ZN(n49580) );
  INV_X2 U213 ( .I(n56886), .ZN(n5658) );
  INV_X2 U8193 ( .I(n10187), .ZN(n4186) );
  BUF_X2 U17487 ( .I(n19904), .Z(n4995) );
  INV_X2 U1445 ( .I(n48586), .ZN(n23813) );
  INV_X2 U8829 ( .I(n36030), .ZN(n36041) );
  NAND3_X2 U14707 ( .A1(n59143), .A2(n18016), .A3(n18015), .ZN(n16854) );
  INV_X4 U34316 ( .I(n56541), .ZN(n14943) );
  NOR3_X2 U1047 ( .A1(n695), .A2(n48571), .A3(n45892), .ZN(n45894) );
  INV_X2 U9971 ( .I(n37761), .ZN(n38283) );
  INV_X2 U43893 ( .I(n3211), .ZN(n26794) );
  INV_X2 U47523 ( .I(n33618), .ZN(n32780) );
  NAND2_X2 U11615 ( .A1(n17183), .A2(n22284), .ZN(n33618) );
  NAND2_X2 U48544 ( .A1(n35569), .A2(n23626), .ZN(n35572) );
  NOR2_X2 U8957 ( .A1(n29585), .A2(n29083), .ZN(n30351) );
  INV_X4 U1700 ( .I(n12677), .ZN(n11986) );
  NOR3_X2 U40846 ( .A1(n60860), .A2(n60971), .A3(n40129), .ZN(n42493) );
  BUF_X4 U6949 ( .I(n44077), .Z(n23267) );
  INV_X2 U3582 ( .I(n33215), .ZN(n35712) );
  BUF_X4 U164 ( .I(n11789), .Z(n60092) );
  NAND2_X2 U4099 ( .A1(n10414), .A2(n19968), .ZN(n52048) );
  NAND2_X2 U41420 ( .A1(n42518), .A2(n41831), .ZN(n42527) );
  NAND2_X2 U4488 ( .A1(n53752), .A2(n25117), .ZN(n20605) );
  NAND4_X2 U3197 ( .A1(n28501), .A2(n28500), .A3(n28499), .A4(n28498), .ZN(
        n28502) );
  OAI21_X2 U14811 ( .A1(n24923), .A2(n49085), .B(n54353), .ZN(n22000) );
  BUF_X4 U17613 ( .I(n23619), .Z(n11751) );
  INV_X2 U30405 ( .I(n22444), .ZN(n29896) );
  NAND2_X2 U19980 ( .A1(n1920), .A2(n50434), .ZN(n50550) );
  INV_X4 U3466 ( .I(n34392), .ZN(n2168) );
  INV_X2 U30254 ( .I(n56962), .ZN(n56958) );
  OAI21_X2 U40470 ( .A1(n23992), .A2(n1380), .B(n25680), .ZN(n20563) );
  NAND2_X2 U4087 ( .A1(n51964), .A2(n55295), .ZN(n55496) );
  INV_X2 U6718 ( .I(n14108), .ZN(n3388) );
  INV_X4 U221 ( .I(n55594), .ZN(n55597) );
  INV_X2 U8465 ( .I(n55584), .ZN(n55566) );
  NOR2_X2 U10859 ( .A1(n16745), .A2(n9395), .ZN(n49406) );
  BUF_X2 U7915 ( .I(n55691), .Z(n23982) );
  INV_X2 U4960 ( .I(n16539), .ZN(n16336) );
  NAND3_X2 U43223 ( .A1(n22889), .A2(n53294), .A3(n4283), .ZN(n53267) );
  NAND2_X2 U4906 ( .A1(n48054), .A2(n21269), .ZN(n48046) );
  NAND2_X2 U367 ( .A1(n57063), .A2(n21235), .ZN(n52670) );
  BUF_X4 U1863 ( .I(n41082), .Z(n9790) );
  NAND2_X2 U35962 ( .A1(n43439), .A2(n43437), .ZN(n42373) );
  NOR2_X2 U2578 ( .A1(n20279), .A2(n24737), .ZN(n34082) );
  NOR3_X2 U28777 ( .A1(n43087), .A2(n8343), .A3(n4659), .ZN(n14262) );
  INV_X2 U13135 ( .I(n40288), .ZN(n1737) );
  NAND2_X2 U31695 ( .A1(n19591), .A2(n63485), .ZN(n19454) );
  INV_X2 U34015 ( .I(n17204), .ZN(n53480) );
  OR2_X2 U1712 ( .A1(n41997), .A2(n462), .Z(n43014) );
  OAI21_X2 U1018 ( .A1(n45665), .A2(n44484), .B(n16964), .ZN(n16965) );
  INV_X2 U10196 ( .I(n39829), .ZN(n13419) );
  NAND3_X2 U51159 ( .A1(n41685), .A2(n42314), .A3(n42001), .ZN(n41686) );
  INV_X2 U11866 ( .I(n53881), .ZN(n54027) );
  BUF_X2 U4837 ( .I(n25323), .Z(n23112) );
  NOR2_X2 U1122 ( .A1(n4526), .A2(n62795), .ZN(n49007) );
  NAND2_X2 U8725 ( .A1(n41859), .A2(n6016), .ZN(n2787) );
  NAND3_X2 U3738 ( .A1(n57442), .A2(n31041), .A3(n12871), .ZN(n30112) );
  INV_X2 U41777 ( .I(n56265), .ZN(n56273) );
  NAND2_X2 U3303 ( .A1(n2059), .A2(n13799), .ZN(n36173) );
  INV_X2 U4744 ( .I(n46570), .ZN(n1488) );
  INV_X2 U12893 ( .I(n43655), .ZN(n1692) );
  INV_X2 U2654 ( .I(n57534), .ZN(n38903) );
  NAND2_X2 U5890 ( .A1(n24069), .A2(n49901), .ZN(n49914) );
  NAND4_X2 U9088 ( .A1(n6355), .A2(n54534), .A3(n54535), .A4(n6354), .ZN(n6353) );
  NAND2_X2 U15664 ( .A1(n36127), .A2(n57631), .ZN(n25354) );
  NAND3_X2 U3652 ( .A1(n64067), .A2(n40832), .A3(n25180), .ZN(n39949) );
  INV_X2 U22140 ( .I(n5942), .ZN(n15722) );
  INV_X2 U11983 ( .I(n28651), .ZN(n28182) );
  BUF_X2 U4988 ( .I(n24811), .Z(n7127) );
  INV_X2 U4294 ( .I(n27229), .ZN(n27480) );
  NOR2_X2 U42688 ( .A1(n33763), .A2(n34798), .ZN(n34795) );
  BUF_X4 U30241 ( .I(n40662), .Z(n10022) );
  NAND2_X2 U1065 ( .A1(n687), .A2(n48678), .ZN(n48882) );
  NAND2_X2 U20803 ( .A1(n16937), .A2(n1587), .ZN(n55237) );
  AOI21_X2 U11858 ( .A1(n30374), .A2(n5768), .B(n30585), .ZN(n5857) );
  NOR2_X2 U29281 ( .A1(n9311), .A2(n17795), .ZN(n56478) );
  INV_X2 U398 ( .I(n5570), .ZN(n1456) );
  INV_X2 U31125 ( .I(n13799), .ZN(n36121) );
  NAND2_X2 U2479 ( .A1(n3306), .A2(n40939), .ZN(n3304) );
  INV_X2 U9152 ( .I(n52987), .ZN(n54493) );
  INV_X4 U9448 ( .I(n39102), .ZN(n40199) );
  NAND3_X2 U3655 ( .A1(n21405), .A2(n21404), .A3(n27912), .ZN(n10951) );
  NAND2_X2 U3242 ( .A1(n1355), .A2(n14503), .ZN(n28554) );
  INV_X4 U26993 ( .I(n52808), .ZN(n25604) );
  BUF_X2 U2158 ( .I(n23495), .Z(n10992) );
  NAND2_X2 U34027 ( .A1(n61729), .A2(n25241), .ZN(n30076) );
  NAND2_X2 U12337 ( .A1(n53781), .A2(n9161), .ZN(n53815) );
  NAND2_X2 U12264 ( .A1(n3895), .A2(n53811), .ZN(n53812) );
  NAND2_X2 U2591 ( .A1(n24799), .A2(n57590), .ZN(n34789) );
  BUF_X4 U3172 ( .I(n21838), .Z(n19255) );
  NAND2_X2 U3776 ( .A1(n27742), .A2(n25978), .ZN(n60407) );
  NOR2_X2 U44757 ( .A1(n29732), .A2(n58696), .ZN(n27742) );
  NAND3_X2 U774 ( .A1(n44409), .A2(n49006), .A3(n49013), .ZN(n49003) );
  OAI21_X2 U336 ( .A1(n13402), .A2(n53437), .B(n17003), .ZN(n60494) );
  INV_X2 U2648 ( .I(n14969), .ZN(n59926) );
  OAI21_X2 U3665 ( .A1(n29500), .A2(n22513), .B(n19186), .ZN(n2653) );
  NOR3_X2 U26250 ( .A1(n60923), .A2(n58772), .A3(n36798), .ZN(n36299) );
  NAND2_X2 U4739 ( .A1(n40613), .A2(n40971), .ZN(n39058) );
  INV_X2 U24471 ( .I(n2989), .ZN(n5099) );
  NAND2_X2 U4684 ( .A1(n30787), .A2(n29747), .ZN(n29954) );
  INV_X2 U40539 ( .I(n35296), .ZN(n34734) );
  NOR2_X2 U3994 ( .A1(n24373), .A2(n3617), .ZN(n29150) );
  OAI21_X2 U5205 ( .A1(n20179), .A2(n30788), .B(n30770), .ZN(n23658) );
  NAND2_X2 U12365 ( .A1(n12037), .A2(n48454), .ZN(n6679) );
  INV_X4 U12704 ( .I(n47472), .ZN(n44680) );
  INV_X4 U41834 ( .I(n59809), .ZN(n36729) );
  NOR2_X2 U9465 ( .A1(n37856), .A2(n37850), .ZN(n6489) );
  BUF_X4 U19922 ( .I(Key[157]), .Z(n23989) );
  AOI21_X1 U29607 ( .A1(n43608), .A2(n42590), .B(n8874), .ZN(n8873) );
  BUF_X4 U30048 ( .I(n35886), .Z(n10596) );
  BUF_X4 U39711 ( .I(n30828), .Z(n33840) );
  INV_X2 U42493 ( .I(n23443), .ZN(n52270) );
  NAND2_X2 U1223 ( .A1(n8842), .A2(n48668), .ZN(n19804) );
  INV_X2 U31267 ( .I(n25867), .ZN(n47682) );
  NOR2_X2 U15433 ( .A1(n49999), .A2(n59633), .ZN(n49202) );
  INV_X2 U18140 ( .I(n37035), .ZN(n2699) );
  NOR2_X2 U835 ( .A1(n48957), .A2(n12673), .ZN(n47058) );
  INV_X2 U31301 ( .I(n18976), .ZN(n25128) );
  NAND2_X2 U1460 ( .A1(n45768), .A2(n6082), .ZN(n46911) );
  NAND2_X2 U1963 ( .A1(n22999), .A2(n5368), .ZN(n41720) );
  NAND2_X2 U15438 ( .A1(n54028), .A2(n6737), .ZN(n54341) );
  NAND3_X2 U2526 ( .A1(n35320), .A2(n35321), .A3(n31955), .ZN(n11000) );
  NAND2_X2 U27618 ( .A1(n53969), .A2(n53950), .ZN(n54007) );
  AND2_X2 U1044 ( .A1(n15708), .A2(n48847), .Z(n57267) );
  AOI21_X2 U16541 ( .A1(n20591), .A2(n5972), .B(n20590), .ZN(n20592) );
  INV_X2 U21004 ( .I(n2694), .ZN(n51625) );
  INV_X2 U27347 ( .I(n42620), .ZN(n22710) );
  INV_X2 U1641 ( .I(n46234), .ZN(n46136) );
  NOR2_X2 U172 ( .A1(n25675), .A2(n23611), .ZN(n10862) );
  NAND3_X2 U26865 ( .A1(n54582), .A2(n58810), .A3(n54561), .ZN(n18424) );
  NAND2_X2 U3865 ( .A1(n17945), .A2(n61708), .ZN(n21036) );
  INV_X2 U3498 ( .I(n13081), .ZN(n57619) );
  NOR2_X2 U653 ( .A1(n15365), .A2(n15363), .ZN(n2646) );
  BUF_X4 U56652 ( .I(n57187), .Z(n61410) );
  OAI21_X2 U45391 ( .A1(n29904), .A2(n1353), .B(n24777), .ZN(n29569) );
  INV_X2 U468 ( .I(n53443), .ZN(n60475) );
  NAND2_X2 U5047 ( .A1(n8212), .A2(n21304), .ZN(n22426) );
  INV_X2 U15547 ( .I(n47343), .ZN(n47943) );
  INV_X2 U3136 ( .I(n29209), .ZN(n30677) );
  INV_X2 U965 ( .I(n48688), .ZN(n47921) );
  AOI21_X2 U21250 ( .A1(n1497), .A2(n541), .B(n60131), .ZN(n41733) );
  INV_X2 U1609 ( .I(n43380), .ZN(n42754) );
  BUF_X4 U4010 ( .I(n28067), .Z(n60768) );
  INV_X2 U12072 ( .I(n26347), .ZN(n28414) );
  AOI21_X2 U17957 ( .A1(n36954), .A2(n20505), .B(n36941), .ZN(n5043) );
  NAND2_X2 U2621 ( .A1(n277), .A2(n39847), .ZN(n7848) );
  BUF_X4 U25456 ( .I(n39491), .Z(n3429) );
  INV_X4 U17437 ( .I(n26182), .ZN(n22384) );
  AOI21_X1 U29822 ( .A1(n55289), .A2(n22592), .B(n59038), .ZN(n15311) );
  BUF_X4 U39440 ( .I(n55648), .Z(n19021) );
  NAND2_X2 U3412 ( .A1(n27135), .A2(n26092), .ZN(n28045) );
  NAND2_X1 U56984 ( .A1(n28326), .A2(n28324), .ZN(n14533) );
  BUF_X4 U10888 ( .I(n44507), .Z(n23534) );
  NAND2_X2 U5145 ( .A1(n7336), .A2(n1262), .ZN(n50222) );
  AOI22_X1 U31737 ( .A1(n33664), .A2(n7183), .B1(n10251), .B2(n22598), .ZN(
        n59321) );
  NAND2_X2 U41100 ( .A1(n61888), .A2(n30296), .ZN(n30301) );
  INV_X4 U39218 ( .I(n50123), .ZN(n18609) );
  INV_X2 U31676 ( .I(n61202), .ZN(n12469) );
  BUF_X4 U23196 ( .I(n42404), .Z(n58343) );
  BUF_X4 U10679 ( .I(n53118), .Z(n23212) );
  NAND2_X2 U37821 ( .A1(n22633), .A2(n21035), .ZN(n16347) );
  INV_X2 U20029 ( .I(n13638), .ZN(n13626) );
  OAI21_X1 U31516 ( .A1(n35902), .A2(n14138), .B(n15488), .ZN(n59291) );
  NAND2_X2 U6218 ( .A1(n32892), .A2(n17199), .ZN(n34193) );
  INV_X4 U1577 ( .I(n43634), .ZN(n5972) );
  NAND3_X2 U3338 ( .A1(n5160), .A2(n5162), .A3(n25350), .ZN(n61096) );
  INV_X2 U26639 ( .I(n5477), .ZN(n19053) );
  INV_X2 U2028 ( .I(n39158), .ZN(n37931) );
  BUF_X4 U125 ( .I(n55223), .Z(n17155) );
  NAND3_X2 U15834 ( .A1(n45079), .A2(n45078), .A3(n45077), .ZN(n45084) );
  NAND2_X2 U28513 ( .A1(n41972), .A2(n19928), .ZN(n8425) );
  INV_X8 U40678 ( .I(n43516), .ZN(n43513) );
  NOR2_X2 U15900 ( .A1(n45971), .A2(n17570), .ZN(n17569) );
  NAND2_X2 U10985 ( .A1(n46176), .A2(n8683), .ZN(n46483) );
  NAND2_X2 U55518 ( .A1(n53724), .A2(n25116), .ZN(n53718) );
  INV_X4 U20571 ( .I(n36851), .ZN(n4754) );
  NAND2_X2 U43919 ( .A1(n48275), .A2(n48832), .ZN(n48276) );
  INV_X4 U11556 ( .I(n15754), .ZN(n35971) );
  INV_X2 U1552 ( .I(n42082), .ZN(n38055) );
  CLKBUF_X4 U24228 ( .I(n52608), .Z(n54860) );
  BUF_X4 U13192 ( .I(Key[103]), .Z(n55191) );
  INV_X2 U43361 ( .I(n22794), .ZN(n56393) );
  NAND2_X2 U4983 ( .A1(n36959), .A2(n1786), .ZN(n159) );
  NAND2_X2 U47691 ( .A1(n14329), .A2(n63866), .ZN(n33532) );
  BUF_X4 U28399 ( .I(n43053), .Z(n8305) );
  INV_X2 U25800 ( .I(n6149), .ZN(n30392) );
  NAND3_X2 U8989 ( .A1(n28140), .A2(n23973), .A3(n28139), .ZN(n28141) );
  OR2_X2 U43478 ( .A1(n17632), .A2(n29282), .Z(n60894) );
  NAND2_X2 U38194 ( .A1(n61198), .A2(n11609), .ZN(n23151) );
  BUF_X4 U29594 ( .I(n49582), .Z(n19773) );
  NAND2_X2 U1086 ( .A1(n13120), .A2(n1640), .ZN(n1630) );
  NOR2_X2 U3722 ( .A1(n31277), .A2(n19118), .ZN(n30871) );
  INV_X4 U31653 ( .I(n11655), .ZN(n22214) );
  INV_X2 U1802 ( .I(n42622), .ZN(n1296) );
  INV_X2 U9742 ( .I(n64145), .ZN(n12589) );
  NAND2_X2 U10625 ( .A1(n60837), .A2(n60836), .ZN(n20591) );
  INV_X2 U25900 ( .I(n6250), .ZN(n6251) );
  INV_X2 U18678 ( .I(n31955), .ZN(n35758) );
  NOR2_X2 U19404 ( .A1(n26854), .A2(n23564), .ZN(n26858) );
  INV_X2 U6235 ( .I(n26849), .ZN(n26853) );
  BUF_X4 U3781 ( .I(n11987), .Z(n61162) );
  NAND3_X2 U884 ( .A1(n49804), .A2(n15220), .A3(n7271), .ZN(n47348) );
  NAND2_X2 U52521 ( .A1(n63501), .A2(n46033), .ZN(n45651) );
  NAND4_X2 U56635 ( .A1(n56680), .A2(n56679), .A3(n56711), .A4(n56699), .ZN(
        n56681) );
  AOI22_X2 U4215 ( .A1(n56677), .A2(n56676), .B1(n56722), .B2(n56730), .ZN(
        n56680) );
  NAND2_X2 U3550 ( .A1(n60633), .A2(n61196), .ZN(n34150) );
  NAND2_X2 U4937 ( .A1(n55131), .A2(n55148), .ZN(n55143) );
  NOR2_X2 U47682 ( .A1(n33564), .A2(n59681), .ZN(n33341) );
  INV_X2 U15142 ( .I(n13674), .ZN(n19888) );
  INV_X2 U20665 ( .I(n243), .ZN(n27087) );
  BUF_X4 U10311 ( .I(n39502), .Z(n40568) );
  INV_X2 U21851 ( .I(n3302), .ZN(n43268) );
  INV_X2 U3840 ( .I(n30810), .ZN(n61187) );
  NAND2_X2 U217 ( .A1(n8194), .A2(n59610), .ZN(n52295) );
  NAND3_X2 U4474 ( .A1(n54641), .A2(n54459), .A3(n55024), .ZN(n54331) );
  INV_X4 U993 ( .I(n61673), .ZN(n1261) );
  INV_X2 U23811 ( .I(n20177), .ZN(n14224) );
  INV_X2 U15549 ( .I(n49010), .ZN(n1626) );
  INV_X4 U10619 ( .I(n24420), .ZN(n29188) );
  INV_X1 U25171 ( .I(n19053), .ZN(n35046) );
  NOR2_X2 U10286 ( .A1(n40572), .A2(n4137), .ZN(n4136) );
  NOR2_X2 U38663 ( .A1(n1895), .A2(n22735), .ZN(n26613) );
  INV_X2 U15062 ( .I(n21343), .ZN(n1614) );
  NAND2_X2 U31532 ( .A1(n59658), .A2(n11106), .ZN(n11105) );
  BUF_X4 U5384 ( .I(n25994), .Z(n23357) );
  BUF_X2 U10158 ( .I(n35152), .Z(n18240) );
  INV_X1 U17425 ( .I(n51474), .ZN(n57753) );
  NAND3_X2 U4162 ( .A1(n50041), .A2(n49441), .A3(n50042), .ZN(n49572) );
  NAND2_X2 U9346 ( .A1(n12338), .A2(n34670), .ZN(n12548) );
  INV_X4 U5273 ( .I(n49582), .ZN(n13440) );
  OAI21_X2 U53390 ( .A1(n47899), .A2(n47895), .B(n47894), .ZN(n47910) );
  INV_X4 U5328 ( .I(n11039), .ZN(n14920) );
  NOR2_X2 U2355 ( .A1(n14282), .A2(n35432), .ZN(n14281) );
  NAND2_X2 U8810 ( .A1(n29002), .A2(n1840), .ZN(n19186) );
  INV_X2 U1063 ( .I(n47773), .ZN(n46866) );
  INV_X4 U28763 ( .I(n61734), .ZN(n29220) );
  NOR2_X2 U25733 ( .A1(n26213), .A2(n60140), .ZN(n36671) );
  NAND2_X2 U20582 ( .A1(n41064), .A2(n41054), .ZN(n19045) );
  NAND2_X2 U99 ( .A1(n55045), .A2(n25220), .ZN(n55065) );
  INV_X2 U144 ( .I(n55076), .ZN(n55045) );
  INV_X2 U1524 ( .I(n13385), .ZN(n43364) );
  INV_X2 U3340 ( .I(n28547), .ZN(n26777) );
  OAI21_X2 U741 ( .A1(n49732), .A2(n1381), .B(n25944), .ZN(n50077) );
  NOR2_X2 U15790 ( .A1(n820), .A2(n63532), .ZN(n27256) );
  INV_X2 U3544 ( .I(n60415), .ZN(n33468) );
  NAND2_X2 U14180 ( .A1(n27888), .A2(n27675), .ZN(n28653) );
  INV_X2 U39384 ( .I(n38529), .ZN(n40959) );
  BUF_X4 U151 ( .I(n21879), .Z(n22667) );
  INV_X2 U10463 ( .I(n29992), .ZN(n1553) );
  INV_X2 U43354 ( .I(n51112), .ZN(n56414) );
  OAI21_X2 U55147 ( .A1(n56216), .A2(n56214), .B(n56621), .ZN(n52713) );
  BUF_X4 U18156 ( .I(n34846), .Z(n38550) );
  NOR3_X2 U42178 ( .A1(n4099), .A2(n4104), .A3(n4102), .ZN(n22100) );
  INV_X4 U7811 ( .I(n8337), .ZN(n47407) );
  NAND3_X2 U27571 ( .A1(n2255), .A2(n6865), .A3(n43577), .ZN(n60681) );
  NAND2_X2 U1817 ( .A1(n43583), .A2(n2898), .ZN(n43576) );
  NAND2_X2 U1873 ( .A1(n20598), .A2(n41051), .ZN(n16823) );
  BUF_X4 U7643 ( .I(n19539), .Z(n10413) );
  NAND3_X1 U23181 ( .A1(n41012), .A2(n58340), .A3(n58339), .ZN(n61039) );
  NAND3_X2 U4028 ( .A1(n1502), .A2(n3619), .A3(n16850), .ZN(n42872) );
  INV_X2 U13528 ( .I(n33684), .ZN(n19922) );
  NAND2_X2 U18497 ( .A1(n32897), .A2(n24287), .ZN(n33684) );
  BUF_X4 U4936 ( .I(n46427), .Z(n21170) );
  NOR2_X2 U13232 ( .A1(n34889), .A2(n34890), .ZN(n14008) );
  INV_X2 U8588 ( .I(n27166), .ZN(n11053) );
  INV_X2 U8554 ( .I(n15477), .ZN(n2706) );
  NAND2_X2 U2372 ( .A1(n37400), .A2(n6540), .ZN(n36327) );
  NOR2_X2 U22802 ( .A1(n47972), .A2(n4271), .ZN(n46082) );
  NOR2_X2 U33108 ( .A1(n22710), .A2(n63983), .ZN(n42621) );
  INV_X2 U546 ( .I(n53241), .ZN(n1283) );
  AND2_X2 U20774 ( .A1(n23489), .A2(n8293), .Z(n8117) );
  BUF_X4 U30735 ( .I(n14505), .Z(n11501) );
  INV_X4 U26890 ( .I(n21623), .ZN(n19544) );
  NOR2_X2 U11642 ( .A1(n7098), .A2(n50336), .ZN(n49867) );
  NOR4_X2 U3194 ( .A1(n16790), .A2(n26704), .A3(n27542), .A4(n26703), .ZN(
        n16789) );
  INV_X4 U5158 ( .I(n56554), .ZN(n1596) );
  NAND3_X2 U11613 ( .A1(n34061), .A2(n34060), .A3(n34059), .ZN(n34062) );
  NAND3_X2 U8635 ( .A1(n12347), .A2(n27187), .A3(n12346), .ZN(n28104) );
  INV_X2 U3295 ( .I(n1443), .ZN(n27868) );
  NOR2_X2 U14834 ( .A1(n5328), .A2(n8119), .ZN(n4746) );
  NOR2_X2 U2772 ( .A1(n34136), .A2(n33389), .ZN(n25617) );
  INV_X2 U43916 ( .I(n24209), .ZN(n47947) );
  OR2_X2 U1101 ( .A1(n4428), .A2(n12100), .Z(n8732) );
  NAND3_X2 U2221 ( .A1(n58262), .A2(n109), .A3(n4918), .ZN(n42276) );
  AOI21_X1 U3659 ( .A1(n7428), .A2(n7427), .B(n53576), .ZN(n53585) );
  INV_X2 U9562 ( .I(n36234), .ZN(n32775) );
  NAND2_X2 U3687 ( .A1(n9701), .A2(n9702), .ZN(n11158) );
  NOR2_X2 U22513 ( .A1(n40591), .A2(n40850), .ZN(n14131) );
  INV_X2 U547 ( .I(n53612), .ZN(n53861) );
  INV_X4 U30326 ( .I(n40174), .ZN(n42694) );
  NOR2_X2 U10471 ( .A1(n30343), .A2(n22504), .ZN(n13360) );
  OAI21_X2 U40686 ( .A1(n27542), .A2(n22456), .B(n27470), .ZN(n27474) );
  NAND4_X2 U6500 ( .A1(n36445), .A2(n35590), .A3(n35589), .A4(n36436), .ZN(
        n4611) );
  OAI21_X2 U17511 ( .A1(n42725), .A2(n2255), .B(n5399), .ZN(n58375) );
  BUF_X4 U9782 ( .I(Key[48]), .Z(n24044) );
  NAND3_X2 U1396 ( .A1(n1387), .A2(n12647), .A3(n45183), .ZN(n47721) );
  INV_X2 U33253 ( .I(n36080), .ZN(n13403) );
  INV_X2 U4309 ( .I(n12930), .ZN(n21826) );
  NAND2_X2 U12724 ( .A1(n57300), .A2(n20208), .ZN(n13864) );
  NAND3_X2 U41636 ( .A1(n51270), .A2(n15966), .A3(n51269), .ZN(n51271) );
  NAND4_X2 U6594 ( .A1(n21816), .A2(n8890), .A3(n8664), .A4(n36687), .ZN(n614)
         );
  NAND2_X2 U10230 ( .A1(n3534), .A2(n6016), .ZN(n41853) );
  INV_X4 U7885 ( .I(n10472), .ZN(n49673) );
  NAND2_X2 U3548 ( .A1(n32924), .A2(n34356), .ZN(n34351) );
  OAI22_X2 U6632 ( .A1(n42654), .A2(n42652), .B1(n1490), .B2(n60846), .ZN(
        n42658) );
  NOR3_X2 U28836 ( .A1(n58949), .A2(n29854), .A3(n15860), .ZN(n3961) );
  NOR2_X2 U26098 ( .A1(n29515), .A2(n17413), .ZN(n29857) );
  NAND2_X2 U4508 ( .A1(n29516), .A2(n58424), .ZN(n29515) );
  INV_X4 U43404 ( .I(n53376), .ZN(n52756) );
  NOR2_X2 U2244 ( .A1(n62720), .A2(n5873), .ZN(n37389) );
  INV_X2 U46976 ( .I(n35297), .ZN(n35302) );
  NAND2_X2 U10052 ( .A1(n41188), .A2(n5488), .ZN(n40720) );
  NAND2_X2 U43477 ( .A1(n46753), .A2(n48148), .ZN(n46794) );
  NOR2_X2 U13742 ( .A1(n37292), .A2(n57479), .ZN(n6835) );
  BUF_X4 U2138 ( .I(n39709), .Z(n21348) );
  NOR2_X2 U42126 ( .A1(n32958), .A2(n21317), .ZN(n61300) );
  NOR2_X2 U48536 ( .A1(n36574), .A2(n24102), .ZN(n35528) );
  BUF_X4 U5340 ( .I(n40416), .Z(n61561) );
  NOR2_X2 U34525 ( .A1(n22669), .A2(n23292), .ZN(n53999) );
  NAND2_X2 U2923 ( .A1(n1776), .A2(n10498), .ZN(n36580) );
  NOR2_X2 U42648 ( .A1(n50407), .A2(n50394), .ZN(n49419) );
  NAND3_X2 U9617 ( .A1(n64797), .A2(n36329), .A3(n37400), .ZN(n36822) );
  INV_X2 U25869 ( .I(n6364), .ZN(n8553) );
  BUF_X4 U8282 ( .I(n30609), .Z(n22504) );
  BUF_X4 U17462 ( .I(n41160), .Z(n10452) );
  INV_X2 U27828 ( .I(n59634), .ZN(n41052) );
  INV_X2 U13128 ( .I(n47700), .ZN(n1385) );
  INV_X4 U42677 ( .I(n22550), .ZN(n54487) );
  INV_X2 U37655 ( .I(n34151), .ZN(n33685) );
  INV_X2 U1626 ( .I(n5358), .ZN(n14313) );
  INV_X2 U31329 ( .I(n61732), .ZN(n32587) );
  NAND2_X2 U3250 ( .A1(n29120), .A2(n22714), .ZN(n29129) );
  NAND2_X1 U4736 ( .A1(n26085), .A2(n65277), .ZN(n635) );
  INV_X2 U9594 ( .I(n17420), .ZN(n1312) );
  NOR2_X2 U5101 ( .A1(n9914), .A2(n42129), .ZN(n42125) );
  INV_X4 U4048 ( .I(n47884), .ZN(n12647) );
  INV_X2 U2419 ( .I(n40061), .ZN(n7057) );
  INV_X2 U40249 ( .I(n11608), .ZN(n43345) );
  INV_X2 U11521 ( .I(n63406), .ZN(n34930) );
  NOR3_X2 U42716 ( .A1(n46870), .A2(n46869), .A3(n46868), .ZN(n46880) );
  AOI21_X2 U17168 ( .A1(n38339), .A2(n39922), .B(n11436), .ZN(n25825) );
  NAND3_X2 U2510 ( .A1(n20815), .A2(n11000), .A3(n35256), .ZN(n6542) );
  NAND2_X2 U8143 ( .A1(n61535), .A2(n61533), .ZN(n29231) );
  OAI21_X2 U11730 ( .A1(n4640), .A2(n5876), .B(n20058), .ZN(n5875) );
  NAND2_X2 U19114 ( .A1(n30340), .A2(n20557), .ZN(n30628) );
  INV_X2 U2659 ( .I(n35316), .ZN(n10327) );
  BUF_X4 U13329 ( .I(n49794), .Z(n23802) );
  BUF_X4 U13444 ( .I(n34469), .Z(n4304) );
  NOR2_X2 U2314 ( .A1(n40487), .A2(n8026), .ZN(n41174) );
  NAND2_X2 U39691 ( .A1(n42127), .A2(n42662), .ZN(n42665) );
  NOR2_X2 U24329 ( .A1(n13074), .A2(n59309), .ZN(n42542) );
  NAND2_X2 U3796 ( .A1(n59760), .A2(n19118), .ZN(n31274) );
  NAND2_X2 U4085 ( .A1(n23879), .A2(n56796), .ZN(n56786) );
  INV_X2 U30529 ( .I(n10202), .ZN(n21495) );
  INV_X2 U3473 ( .I(n24990), .ZN(n3403) );
  NAND2_X2 U36369 ( .A1(n2168), .A2(n18218), .ZN(n19312) );
  INV_X2 U39791 ( .I(n61681), .ZN(n51931) );
  INV_X2 U10128 ( .I(n40998), .ZN(n6768) );
  NAND2_X2 U2337 ( .A1(n58672), .A2(n16601), .ZN(n41015) );
  INV_X4 U37974 ( .I(n57199), .ZN(n25201) );
  OAI21_X2 U11818 ( .A1(n759), .A2(n18872), .B(n31202), .ZN(n20538) );
  BUF_X2 U15703 ( .I(n18599), .Z(n9772) );
  AOI21_X2 U56227 ( .A1(n55618), .A2(n55651), .B(n55617), .ZN(n55621) );
  NAND2_X2 U15161 ( .A1(n4513), .A2(n50929), .ZN(n9208) );
  NOR2_X2 U9580 ( .A1(n60926), .A2(n63617), .ZN(n33756) );
  INV_X4 U4878 ( .I(n15692), .ZN(n15693) );
  NOR2_X2 U127 ( .A1(n53351), .A2(n53355), .ZN(n53332) );
  NAND2_X2 U27515 ( .A1(n15548), .A2(n39007), .ZN(n39050) );
  INV_X2 U30024 ( .I(n22349), .ZN(n14451) );
  NAND2_X2 U4487 ( .A1(n18724), .A2(n42985), .ZN(n43297) );
  OAI21_X2 U15338 ( .A1(n2321), .A2(n49324), .B(n49323), .ZN(n13788) );
  NAND2_X2 U4507 ( .A1(n17414), .A2(n29516), .ZN(n61270) );
  NAND2_X2 U30340 ( .A1(n14103), .A2(n26041), .ZN(n54055) );
  NAND2_X1 U5651 ( .A1(n13372), .A2(n53670), .ZN(n320) );
  INV_X2 U38393 ( .I(n25094), .ZN(n27233) );
  INV_X1 U39723 ( .I(n55416), .ZN(n55252) );
  NAND2_X2 U4164 ( .A1(n50041), .A2(n19773), .ZN(n12966) );
  NOR2_X2 U5304 ( .A1(n40629), .A2(n41193), .ZN(n17579) );
  NOR3_X2 U19481 ( .A1(n48891), .A2(n4580), .A3(n4579), .ZN(n9993) );
  NOR3_X1 U40778 ( .A1(n8099), .A2(n8098), .A3(n8101), .ZN(n16457) );
  AND2_X2 U27050 ( .A1(n35025), .A2(n33519), .Z(n23125) );
  INV_X2 U2091 ( .I(n65271), .ZN(n20277) );
  INV_X2 U1599 ( .I(n41583), .ZN(n1297) );
  BUF_X4 U32355 ( .I(n20893), .Z(n12312) );
  INV_X2 U1297 ( .I(n11417), .ZN(n8048) );
  BUF_X4 U9229 ( .I(n46719), .Z(n50394) );
  INV_X2 U4698 ( .I(n43924), .ZN(n13730) );
  AOI22_X2 U3527 ( .A1(n8405), .A2(n23743), .B1(n14361), .B2(n35821), .ZN(
        n34319) );
  NAND2_X2 U50897 ( .A1(n41881), .A2(n41065), .ZN(n40847) );
  INV_X2 U41686 ( .I(n55692), .ZN(n55302) );
  INV_X2 U5181 ( .I(n26163), .ZN(n20800) );
  INV_X2 U10177 ( .I(n39136), .ZN(n39130) );
  INV_X8 U1738 ( .I(n24361), .ZN(n43733) );
  NAND3_X2 U20094 ( .A1(n49330), .A2(n1375), .A3(n49394), .ZN(n11843) );
  NAND2_X2 U30654 ( .A1(n14314), .A2(n49908), .ZN(n44663) );
  NAND2_X2 U41480 ( .A1(n23191), .A2(n23942), .ZN(n26612) );
  NOR2_X2 U2976 ( .A1(n29516), .A2(n17412), .ZN(n29864) );
  NAND2_X2 U25803 ( .A1(n6152), .A2(n1825), .ZN(n6151) );
  NAND3_X2 U1036 ( .A1(n1383), .A2(n62413), .A3(n50215), .ZN(n18833) );
  OAI22_X2 U4253 ( .A1(n19560), .A2(n36557), .B1(n36559), .B2(n36558), .ZN(
        n36560) );
  INV_X2 U37745 ( .I(n38093), .ZN(n41293) );
  INV_X2 U19290 ( .I(n29099), .ZN(n18716) );
  OAI21_X2 U30492 ( .A1(n17724), .A2(n27118), .B(n17721), .ZN(n14220) );
  NAND2_X2 U9427 ( .A1(n41472), .A2(n41470), .ZN(n40412) );
  NOR4_X2 U55680 ( .A1(n10464), .A2(n54127), .A3(n54195), .A4(n15969), .ZN(
        n54133) );
  INV_X2 U14960 ( .I(n55293), .ZN(n24904) );
  BUF_X2 U11974 ( .I(n54465), .Z(n23897) );
  BUF_X2 U5911 ( .I(n20086), .Z(n61198) );
  NOR2_X2 U47542 ( .A1(n33566), .A2(n32809), .ZN(n32811) );
  INV_X2 U22437 ( .I(n54325), .ZN(n3769) );
  INV_X4 U26579 ( .I(n25482), .ZN(n47542) );
  NAND2_X2 U28736 ( .A1(n9437), .A2(n8639), .ZN(n25482) );
  AND2_X2 U11537 ( .A1(n36070), .A2(n25677), .Z(n14196) );
  INV_X2 U10740 ( .I(n43316), .ZN(n43317) );
  NAND2_X2 U32779 ( .A1(n55108), .A2(n11353), .ZN(n61338) );
  NAND2_X2 U4540 ( .A1(n7041), .A2(n55151), .ZN(n55108) );
  BUF_X2 U10757 ( .I(n55444), .Z(n23522) );
  NAND3_X1 U28170 ( .A1(n58864), .A2(n37930), .A3(n62157), .ZN(n61619) );
  INV_X2 U2802 ( .I(n33869), .ZN(n18596) );
  NAND2_X2 U4657 ( .A1(n34602), .A2(n21106), .ZN(n31023) );
  NAND2_X2 U12677 ( .A1(n47737), .A2(n47434), .ZN(n46745) );
  NAND2_X2 U21696 ( .A1(n61658), .A2(n3356), .ZN(n40990) );
  NOR2_X2 U1959 ( .A1(n40173), .A2(n1393), .ZN(n41531) );
  INV_X4 U54465 ( .I(n36246), .ZN(n61223) );
  NAND2_X2 U2502 ( .A1(n41810), .A2(n2459), .ZN(n38194) );
  NOR2_X2 U7186 ( .A1(n1685), .A2(n41695), .ZN(n8053) );
  NOR3_X2 U2700 ( .A1(n20792), .A2(n35855), .A3(n8295), .ZN(n5557) );
  NAND2_X2 U2424 ( .A1(n42486), .A2(n59851), .ZN(n40092) );
  NAND3_X2 U11283 ( .A1(n47599), .A2(n47598), .A3(n47597), .ZN(n47600) );
  NOR2_X2 U7036 ( .A1(n59958), .A2(n41688), .ZN(n8322) );
  NAND3_X2 U5832 ( .A1(n41686), .A2(n10651), .A3(n22469), .ZN(n59958) );
  NAND3_X2 U1699 ( .A1(n41565), .A2(n41566), .A3(n16204), .ZN(n41575) );
  INV_X2 U1479 ( .I(n2634), .ZN(n48488) );
  NOR2_X2 U3292 ( .A1(n25206), .A2(n58664), .ZN(n25205) );
  NAND2_X2 U4497 ( .A1(n13332), .A2(n13327), .ZN(n13331) );
  NAND3_X1 U50742 ( .A1(n40382), .A2(n22638), .A3(n40381), .ZN(n40383) );
  INV_X4 U20507 ( .I(n2867), .ZN(n41054) );
  INV_X4 U33767 ( .I(n29915), .ZN(n14202) );
  INV_X4 U16999 ( .I(n55474), .ZN(n57720) );
  INV_X4 U13701 ( .I(n35691), .ZN(n10682) );
  NOR2_X2 U5433 ( .A1(n63520), .A2(n15700), .ZN(n59108) );
  NAND2_X2 U12062 ( .A1(n28003), .A2(n27014), .ZN(n28219) );
  NOR2_X2 U5726 ( .A1(n59532), .A2(n1295), .ZN(n45971) );
  OAI21_X2 U4368 ( .A1(n24337), .A2(n24336), .B(n63001), .ZN(n3861) );
  BUF_X4 U16934 ( .I(n42916), .Z(n5773) );
  INV_X1 U24724 ( .I(n24839), .ZN(n58591) );
  NOR3_X1 U51317 ( .A1(n42291), .A2(n43995), .A3(n16880), .ZN(n42310) );
  NAND2_X2 U10222 ( .A1(n36110), .A2(n36412), .ZN(n36409) );
  INV_X2 U31488 ( .I(n13811), .ZN(n12382) );
  INV_X4 U6880 ( .I(n12312), .ZN(n25851) );
  INV_X4 U907 ( .I(n57204), .ZN(n45547) );
  NAND2_X2 U16787 ( .A1(n41507), .A2(n19004), .ZN(n10196) );
  NAND2_X2 U55301 ( .A1(n53033), .A2(n64608), .ZN(n53034) );
  NAND2_X2 U8962 ( .A1(n12125), .A2(n19118), .ZN(n31281) );
  INV_X4 U43455 ( .I(n3510), .ZN(n47605) );
  NAND2_X2 U6841 ( .A1(n20260), .A2(n35841), .ZN(n34409) );
  INV_X2 U13799 ( .I(n29002), .ZN(n30390) );
  NAND2_X2 U21091 ( .A1(n25459), .A2(n49014), .ZN(n3885) );
  NOR2_X2 U8846 ( .A1(n5082), .A2(n5086), .ZN(n32458) );
  NAND2_X2 U3589 ( .A1(n1811), .A2(n58105), .ZN(n32678) );
  NAND2_X2 U2726 ( .A1(n22633), .A2(n35816), .ZN(n35309) );
  INV_X2 U37732 ( .I(n42804), .ZN(n19428) );
  INV_X2 U23604 ( .I(n45972), .ZN(n8603) );
  AOI21_X2 U5582 ( .A1(n49359), .A2(n49358), .B(n14171), .ZN(n14170) );
  INV_X4 U34515 ( .I(n15245), .ZN(n23554) );
  BUF_X4 U13699 ( .I(n22477), .Z(n5250) );
  NAND2_X1 U28979 ( .A1(n8964), .A2(n55432), .ZN(n8966) );
  INV_X2 U78 ( .I(n11275), .ZN(n54391) );
  NAND2_X2 U9694 ( .A1(n36452), .A2(n15038), .ZN(n36445) );
  NAND2_X2 U10787 ( .A1(n4528), .A2(n5700), .ZN(n5698) );
  NOR2_X1 U25988 ( .A1(n337), .A2(n55424), .ZN(n58735) );
  OAI21_X2 U1293 ( .A1(n1328), .A2(n59406), .B(n45503), .ZN(n59383) );
  OAI22_X2 U13491 ( .A1(n12539), .A2(n9517), .B1(n61078), .B2(n4075), .ZN(
        n33439) );
  NAND2_X2 U5403 ( .A1(n2351), .A2(n64950), .ZN(n24712) );
  INV_X2 U33074 ( .I(n47729), .ZN(n46736) );
  NAND2_X2 U18676 ( .A1(n33622), .A2(n58998), .ZN(n17183) );
  INV_X2 U11148 ( .I(n42401), .ZN(n41694) );
  OAI21_X2 U340 ( .A1(n55260), .A2(n55259), .B(n55264), .ZN(n24530) );
  NAND2_X2 U15766 ( .A1(n25863), .A2(n45800), .ZN(n25862) );
  INV_X1 U9031 ( .I(n13704), .ZN(n5548) );
  INV_X4 U497 ( .I(n61893), .ZN(n12074) );
  BUF_X4 U23193 ( .I(n24180), .Z(n6052) );
  NOR2_X2 U37741 ( .A1(n63454), .A2(n15791), .ZN(n29512) );
  NOR2_X2 U8446 ( .A1(n35723), .A2(n23742), .ZN(n37218) );
  NAND3_X2 U3261 ( .A1(n27178), .A2(n21281), .A3(n24878), .ZN(n27608) );
  INV_X2 U232 ( .I(n22782), .ZN(n54403) );
  NAND3_X2 U4322 ( .A1(n59982), .A2(n25397), .A3(n59981), .ZN(n22154) );
  NOR2_X2 U7056 ( .A1(n61748), .A2(n14111), .ZN(n34997) );
  NOR2_X2 U2568 ( .A1(n1409), .A2(n41020), .ZN(n19458) );
  NOR3_X2 U715 ( .A1(n4018), .A2(n4014), .A3(n46091), .ZN(n4013) );
  BUF_X8 U4547 ( .I(n15152), .Z(n33) );
  OAI21_X2 U27516 ( .A1(n56604), .A2(n56982), .B(n59404), .ZN(n56614) );
  OAI21_X2 U11504 ( .A1(n36790), .A2(n61579), .B(n57211), .ZN(n4680) );
  NAND3_X2 U9234 ( .A1(n139), .A2(n1812), .A3(n33949), .ZN(n34120) );
  NOR2_X2 U27479 ( .A1(n56607), .A2(n56608), .ZN(n20781) );
  NAND2_X2 U4753 ( .A1(n13757), .A2(n56978), .ZN(n56604) );
  INV_X8 U7527 ( .I(n12521), .ZN(n37400) );
  INV_X1 U15082 ( .I(n18308), .ZN(n26090) );
  NOR2_X2 U795 ( .A1(n19773), .A2(n20428), .ZN(n50049) );
  INV_X2 U31510 ( .I(n33467), .ZN(n61261) );
  NOR2_X2 U875 ( .A1(n15550), .A2(n49940), .ZN(n50272) );
  NAND2_X2 U12355 ( .A1(n14713), .A2(n20477), .ZN(n56921) );
  AOI21_X2 U4291 ( .A1(n56787), .A2(n56788), .B(n56786), .ZN(n56807) );
  NOR2_X2 U1984 ( .A1(n41568), .A2(n24884), .ZN(n41704) );
  AOI21_X2 U53249 ( .A1(n47389), .A2(n47388), .B(n47387), .ZN(n47394) );
  NOR2_X2 U162 ( .A1(n15245), .A2(n55385), .ZN(n9424) );
  AOI21_X2 U23390 ( .A1(n43570), .A2(n1696), .B(n58375), .ZN(n60817) );
  NAND4_X2 U1814 ( .A1(n1397), .A2(n43573), .A3(n43572), .A4(n5398), .ZN(n5399) );
  NAND2_X2 U11311 ( .A1(n40395), .A2(n63119), .ZN(n41081) );
  NAND2_X2 U2401 ( .A1(n36423), .A2(n2056), .ZN(n21801) );
  INV_X2 U9203 ( .I(n48876), .ZN(n1375) );
  NAND2_X2 U896 ( .A1(n8604), .A2(n15753), .ZN(n48876) );
  INV_X2 U13584 ( .I(n54950), .ZN(n59081) );
  NAND2_X2 U25157 ( .A1(n49674), .A2(n5463), .ZN(n49372) );
  INV_X4 U27370 ( .I(n9185), .ZN(n23003) );
  AOI21_X2 U429 ( .A1(n55302), .A2(n2524), .B(n55300), .ZN(n52920) );
  NOR2_X2 U5131 ( .A1(n16995), .A2(n55237), .ZN(n55179) );
  BUF_X4 U41733 ( .I(n6168), .Z(n60426) );
  BUF_X4 U11039 ( .I(n57630), .Z(n2540) );
  INV_X2 U2128 ( .I(n37625), .ZN(n39743) );
  INV_X2 U1533 ( .I(n15044), .ZN(n43873) );
  NAND2_X2 U8283 ( .A1(n6206), .A2(n61496), .ZN(n35286) );
  INV_X2 U17447 ( .I(n38024), .ZN(n8484) );
  NOR2_X2 U45944 ( .A1(n30889), .A2(n30888), .ZN(n31239) );
  AND2_X2 U19327 ( .A1(n25349), .A2(n5933), .Z(n30889) );
  INV_X4 U20257 ( .I(n3233), .ZN(n22113) );
  BUF_X2 U6217 ( .I(n6041), .Z(n58765) );
  NAND2_X2 U29187 ( .A1(n20180), .A2(n42923), .ZN(n42917) );
  INV_X2 U2120 ( .I(n36370), .ZN(n39598) );
  INV_X2 U2039 ( .I(n15930), .ZN(n25570) );
  NAND2_X2 U10867 ( .A1(n1327), .A2(n12579), .ZN(n50375) );
  INV_X2 U27681 ( .I(n26210), .ZN(n54317) );
  NOR3_X2 U19814 ( .A1(n15811), .A2(n57009), .A3(n56388), .ZN(n17621) );
  OAI21_X2 U9334 ( .A1(n43131), .A2(n22606), .B(n57177), .ZN(n26227) );
  NOR2_X2 U35778 ( .A1(n35863), .A2(n35065), .ZN(n16663) );
  INV_X4 U9367 ( .I(n61134), .ZN(n11606) );
  NAND2_X2 U47524 ( .A1(n33622), .A2(n64838), .ZN(n32781) );
  NAND2_X2 U33297 ( .A1(n36553), .A2(n1339), .ZN(n36098) );
  NOR3_X2 U6715 ( .A1(n8548), .A2(n8547), .A3(n8546), .ZN(n8630) );
  NAND2_X2 U35956 ( .A1(n43699), .A2(n14214), .ZN(n16677) );
  OAI21_X2 U5909 ( .A1(n18741), .A2(n1272), .B(n41079), .ZN(n39970) );
  NAND2_X2 U36482 ( .A1(n35575), .A2(n36037), .ZN(n17488) );
  NOR2_X2 U43160 ( .A1(n24586), .A2(n23482), .ZN(n54016) );
  NAND2_X2 U23093 ( .A1(n54950), .A2(n54605), .ZN(n4319) );
  NOR4_X2 U736 ( .A1(n23421), .A2(n57723), .A3(n25501), .A4(n49021), .ZN(n7431) );
  NOR3_X2 U27692 ( .A1(n41072), .A2(n41073), .A3(n7618), .ZN(n40855) );
  BUF_X2 U41830 ( .I(n54546), .Z(n22572) );
  NAND2_X2 U854 ( .A1(n48717), .A2(n1224), .ZN(n49881) );
  INV_X2 U53240 ( .I(n19847), .ZN(n47351) );
  NAND2_X2 U52593 ( .A1(n45652), .A2(n46039), .ZN(n46865) );
  INV_X2 U41767 ( .I(n44518), .ZN(n46535) );
  NOR2_X2 U6125 ( .A1(n10550), .A2(n36332), .ZN(n11006) );
  NOR2_X2 U4122 ( .A1(n5324), .A2(n54424), .ZN(n54402) );
  NOR2_X2 U5014 ( .A1(n45486), .A2(n11183), .ZN(n45710) );
  INV_X2 U39863 ( .I(n38134), .ZN(n23501) );
  AOI21_X2 U3835 ( .A1(n36600), .A2(n36599), .B(n36598), .ZN(n36601) );
  NAND2_X2 U4925 ( .A1(n15784), .A2(n24405), .ZN(n8351) );
  INV_X2 U42156 ( .I(n56638), .ZN(n56206) );
  BUF_X4 U54528 ( .I(n56182), .Z(n61228) );
  NAND2_X2 U16758 ( .A1(n42017), .A2(n42931), .ZN(n3970) );
  NAND2_X2 U10758 ( .A1(n43495), .A2(n20100), .ZN(n6071) );
  NAND2_X2 U2494 ( .A1(n34549), .A2(n3721), .ZN(n3720) );
  BUF_X4 U4691 ( .I(n55582), .Z(n21272) );
  NAND2_X2 U38697 ( .A1(n12907), .A2(n16279), .ZN(n31042) );
  INV_X2 U310 ( .I(n57009), .ZN(n13902) );
  INV_X2 U23752 ( .I(n46872), .ZN(n47772) );
  AOI21_X2 U14111 ( .A1(n28190), .A2(n26913), .B(n27675), .ZN(n20099) );
  NOR3_X2 U53095 ( .A1(n46866), .A2(n46864), .A3(n64849), .ZN(n46869) );
  BUF_X4 U12483 ( .I(n10636), .Z(n19294) );
  NAND2_X2 U14605 ( .A1(n504), .A2(n16337), .ZN(n36945) );
  INV_X2 U10869 ( .I(n49687), .ZN(n16922) );
  NAND2_X2 U4862 ( .A1(n54440), .A2(n54815), .ZN(n54441) );
  NOR2_X1 U17875 ( .A1(n61341), .A2(n61340), .ZN(n57857) );
  NAND2_X2 U33522 ( .A1(n34614), .A2(n33420), .ZN(n34033) );
  NAND3_X2 U4918 ( .A1(n10624), .A2(n48572), .A3(n48081), .ZN(n13296) );
  AOI21_X2 U10608 ( .A1(n41767), .A2(n41766), .B(n43167), .ZN(n40687) );
  BUF_X4 U9606 ( .I(n32754), .Z(n13520) );
  INV_X2 U957 ( .I(n45160), .ZN(n48349) );
  NAND2_X2 U22870 ( .A1(n19102), .A2(n64077), .ZN(n42495) );
  INV_X2 U41151 ( .I(n21395), .ZN(n55312) );
  BUF_X4 U16925 ( .I(n18742), .Z(n8028) );
  INV_X2 U20722 ( .I(n9436), .ZN(n18856) );
  AOI22_X2 U35625 ( .A1(n52705), .A2(n56381), .B1(n15988), .B2(n17198), .ZN(
        n21324) );
  NOR2_X2 U1353 ( .A1(n6494), .A2(n9064), .ZN(n6493) );
  NAND3_X1 U12985 ( .A1(n7337), .A2(n16775), .A3(n41944), .ZN(n13198) );
  INV_X2 U7543 ( .I(n22092), .ZN(n15454) );
  NOR2_X2 U10784 ( .A1(n20741), .A2(n48844), .ZN(n18479) );
  NAND2_X1 U38715 ( .A1(n60037), .A2(n15846), .ZN(n16976) );
  NAND4_X1 U24328 ( .A1(n56975), .A2(n56972), .A3(n56973), .A4(n56974), .ZN(
        n59069) );
  INV_X4 U33966 ( .I(n14498), .ZN(n18724) );
  OAI21_X2 U30148 ( .A1(n1626), .A2(n63389), .B(n14401), .ZN(n14400) );
  NAND2_X2 U36632 ( .A1(n25305), .A2(n23399), .ZN(n42470) );
  NOR2_X2 U53437 ( .A1(n5463), .A2(n4780), .ZN(n48011) );
  NAND2_X2 U1121 ( .A1(n62424), .A2(n59698), .ZN(n3808) );
  INV_X4 U26325 ( .I(n7175), .ZN(n11279) );
  NAND2_X2 U19127 ( .A1(n50367), .A2(n60209), .ZN(n49129) );
  NAND3_X1 U3669 ( .A1(n25904), .A2(n10436), .A3(n25906), .ZN(n7375) );
  BUF_X4 U6017 ( .I(n7641), .Z(n60957) );
  NAND2_X2 U2701 ( .A1(n16736), .A2(n5472), .ZN(n8009) );
  INV_X2 U10351 ( .I(n13942), .ZN(n33627) );
  INV_X4 U33554 ( .I(n57686), .ZN(n37096) );
  INV_X2 U146 ( .I(n22343), .ZN(n55222) );
  NOR2_X2 U2350 ( .A1(n13768), .A2(n35964), .ZN(n35551) );
  NAND2_X2 U4049 ( .A1(n47884), .A2(n64548), .ZN(n47725) );
  INV_X2 U12097 ( .I(n28349), .ZN(n1447) );
  CLKBUF_X4 U9989 ( .I(n11074), .Z(n5712) );
  INV_X2 U6737 ( .I(n35876), .ZN(n37327) );
  INV_X2 U3304 ( .I(n24373), .ZN(n1444) );
  NAND2_X2 U2561 ( .A1(n33509), .A2(n7883), .ZN(n34544) );
  NOR2_X2 U9231 ( .A1(n9818), .A2(n21449), .ZN(n9817) );
  INV_X2 U12310 ( .I(n10464), .ZN(n54187) );
  NAND2_X2 U27414 ( .A1(n40703), .A2(n17831), .ZN(n41438) );
  NAND4_X2 U5417 ( .A1(n53975), .A2(n53974), .A3(n53977), .A4(n53976), .ZN(
        n58905) );
  INV_X4 U32618 ( .I(n25623), .ZN(n24147) );
  INV_X2 U7368 ( .I(n57115), .ZN(n57134) );
  OR2_X2 U17258 ( .A1(n14903), .A2(n24406), .Z(n27203) );
  NOR2_X1 U25151 ( .A1(n43871), .A2(n5800), .ZN(n6146) );
  NOR2_X2 U29268 ( .A1(n1310), .A2(n9304), .ZN(n36212) );
  BUF_X4 U13998 ( .I(n30748), .Z(n3761) );
  BUF_X4 U18154 ( .I(n36080), .Z(n18496) );
  INV_X2 U11811 ( .I(n29814), .ZN(n30482) );
  INV_X2 U28487 ( .I(n8389), .ZN(n9139) );
  NOR2_X2 U26857 ( .A1(n17467), .A2(n6705), .ZN(n42837) );
  NOR3_X2 U14455 ( .A1(n26168), .A2(n60621), .A3(n60620), .ZN(n22668) );
  OAI21_X2 U5522 ( .A1(n28721), .A2(n28722), .B(n28720), .ZN(n20551) );
  NAND2_X2 U29496 ( .A1(n15515), .A2(n15516), .ZN(n16894) );
  NOR2_X2 U2227 ( .A1(n20161), .A2(n35343), .ZN(n20160) );
  NAND2_X2 U35072 ( .A1(n18128), .A2(n30786), .ZN(n29551) );
  NAND2_X2 U2589 ( .A1(n34746), .A2(n8800), .ZN(n34751) );
  NAND2_X2 U7217 ( .A1(n42067), .A2(n1193), .ZN(n42964) );
  NAND3_X2 U10200 ( .A1(n24066), .A2(n1746), .A3(n2459), .ZN(n4227) );
  NOR2_X2 U5108 ( .A1(n18422), .A2(n54507), .ZN(n54574) );
  NAND3_X2 U48689 ( .A1(n36412), .A2(n21591), .A3(n36404), .ZN(n36117) );
  INV_X4 U7238 ( .I(n59629), .ZN(n47821) );
  NAND2_X2 U5224 ( .A1(n33961), .A2(n12539), .ZN(n25634) );
  NAND2_X2 U948 ( .A1(n21870), .A2(n50257), .ZN(n49937) );
  INV_X2 U30845 ( .I(n10079), .ZN(n23778) );
  BUF_X4 U6250 ( .I(n60417), .Z(n11627) );
  NOR2_X2 U19013 ( .A1(n29807), .A2(n29806), .ZN(n29809) );
  NOR2_X2 U15318 ( .A1(n22038), .A2(n9379), .ZN(n9387) );
  OAI22_X2 U1196 ( .A1(n58258), .A2(n47404), .B1(n8126), .B2(n70), .ZN(n58604)
         );
  AOI22_X2 U45766 ( .A1(n2825), .A2(n30460), .B1(n30459), .B2(n30458), .ZN(
        n30474) );
  BUF_X4 U18134 ( .I(n31910), .Z(n35876) );
  NOR2_X2 U7016 ( .A1(n29566), .A2(n60886), .ZN(n28957) );
  NOR3_X2 U2518 ( .A1(n12859), .A2(n34628), .A3(n61078), .ZN(n3582) );
  NOR3_X1 U9475 ( .A1(n13343), .A2(n33790), .A3(n13342), .ZN(n13344) );
  NOR2_X2 U837 ( .A1(n48678), .A2(n49701), .ZN(n24049) );
  BUF_X4 U13216 ( .I(n20667), .Z(n9896) );
  INV_X4 U30450 ( .I(n13976), .ZN(n31141) );
  BUF_X4 U31079 ( .I(n37648), .Z(n41132) );
  INV_X2 U4522 ( .I(n9953), .ZN(n15877) );
  NAND3_X2 U52229 ( .A1(n52807), .A2(n52808), .A3(n52806), .ZN(n53322) );
  NOR2_X2 U43492 ( .A1(n3335), .A2(n1637), .ZN(n49356) );
  NAND2_X2 U26353 ( .A1(n25246), .A2(n40090), .ZN(n6702) );
  INV_X2 U15132 ( .I(n8550), .ZN(n50761) );
  AND2_X2 U20057 ( .A1(n9049), .A2(n58527), .Z(n42484) );
  NAND2_X1 U31042 ( .A1(n39885), .A2(n40128), .ZN(n10569) );
  NOR2_X2 U12798 ( .A1(n57454), .A2(n24518), .ZN(n12043) );
  NOR2_X2 U1679 ( .A1(n8799), .A2(n42608), .ZN(n24518) );
  NAND2_X2 U40927 ( .A1(n47184), .A2(n47183), .ZN(n21033) );
  AOI22_X2 U39897 ( .A1(n47178), .A2(n47179), .B1(n48219), .B2(n47177), .ZN(
        n47184) );
  NAND2_X2 U16505 ( .A1(n1942), .A2(n43495), .ZN(n1940) );
  INV_X2 U1343 ( .I(n25244), .ZN(n18584) );
  OAI21_X1 U35683 ( .A1(n30012), .A2(n31220), .B(n1278), .ZN(n59770) );
  BUF_X4 U24152 ( .I(n25051), .Z(n59046) );
  OAI22_X2 U31165 ( .A1(n26635), .A2(n22234), .B1(n28381), .B2(n26551), .ZN(
        n26552) );
  NOR2_X2 U1744 ( .A1(n1296), .A2(n42099), .ZN(n58223) );
  NOR2_X2 U3247 ( .A1(n36926), .A2(n15171), .ZN(n11780) );
  NOR2_X2 U9966 ( .A1(n58064), .A2(n47604), .ZN(n43192) );
  NAND2_X2 U168 ( .A1(n16383), .A2(n55218), .ZN(n55226) );
  INV_X2 U11547 ( .I(n7380), .ZN(n36463) );
  NOR2_X2 U23550 ( .A1(n19127), .A2(n36489), .ZN(n7433) );
  NAND2_X2 U3809 ( .A1(n22799), .A2(n29736), .ZN(n11195) );
  INV_X2 U7911 ( .I(n56568), .ZN(n11119) );
  NAND2_X2 U26780 ( .A1(n22619), .A2(n22618), .ZN(n56128) );
  AOI21_X2 U51332 ( .A1(n42367), .A2(n43439), .B(n42366), .ZN(n42368) );
  OAI21_X2 U28270 ( .A1(n39945), .A2(n64450), .B(n23698), .ZN(n39946) );
  AND3_X2 U12590 ( .A1(n41064), .A2(n40841), .A3(n6855), .Z(n57280) );
  INV_X2 U32639 ( .I(n24672), .ZN(n31924) );
  INV_X2 U42115 ( .I(n42127), .ZN(n41559) );
  NOR2_X2 U31109 ( .A1(n29303), .A2(n29292), .ZN(n27219) );
  NOR2_X2 U11509 ( .A1(n35482), .A2(n37049), .ZN(n36607) );
  AOI21_X2 U35566 ( .A1(n49561), .A2(n49566), .B(n25128), .ZN(n48282) );
  OAI21_X2 U8971 ( .A1(n59561), .A2(n13335), .B(n9250), .ZN(n12562) );
  OAI21_X2 U36520 ( .A1(n1419), .A2(n60562), .B(n1792), .ZN(n36227) );
  INV_X2 U3010 ( .I(n30691), .ZN(n31054) );
  INV_X2 U10367 ( .I(n35666), .ZN(n1341) );
  INV_X4 U6000 ( .I(n2564), .ZN(n23969) );
  NOR2_X2 U41099 ( .A1(n21945), .A2(n34127), .ZN(n32869) );
  NAND2_X2 U873 ( .A1(n48688), .A2(n1474), .ZN(n48685) );
  NAND2_X2 U9551 ( .A1(n35706), .A2(n5999), .ZN(n328) );
  INV_X4 U32426 ( .I(n16543), .ZN(n50367) );
  NOR4_X2 U4218 ( .A1(n25765), .A2(n25762), .A3(n54580), .A4(n54524), .ZN(
        n59939) );
  NOR2_X2 U53397 ( .A1(n47919), .A2(n48688), .ZN(n49047) );
  AOI21_X2 U19454 ( .A1(n27566), .A2(n23039), .B(n15534), .ZN(n14651) );
  NAND2_X2 U712 ( .A1(n5703), .A2(n57821), .ZN(n57820) );
  NOR2_X2 U12467 ( .A1(n23612), .A2(n49166), .ZN(n18690) );
  INV_X4 U4065 ( .I(n43912), .ZN(n15695) );
  NAND2_X2 U2246 ( .A1(n16337), .A2(n59842), .ZN(n36947) );
  NAND2_X2 U6361 ( .A1(n13535), .A2(n12489), .ZN(n13980) );
  INV_X4 U45219 ( .I(n53805), .ZN(n29070) );
  NAND2_X2 U39054 ( .A1(n23503), .A2(n18313), .ZN(n36407) );
  NAND2_X2 U6052 ( .A1(n130), .A2(n34906), .ZN(n34911) );
  NOR2_X2 U31541 ( .A1(n39418), .A2(n40070), .ZN(n40166) );
  INV_X2 U11635 ( .I(n15649), .ZN(n6301) );
  NOR2_X2 U4985 ( .A1(n54575), .A2(n18229), .ZN(n54524) );
  AOI21_X2 U26060 ( .A1(n48423), .A2(n6411), .B(n49711), .ZN(n17134) );
  INV_X4 U2632 ( .I(n8304), .ZN(n12338) );
  INV_X4 U3872 ( .I(n25685), .ZN(n11243) );
  NAND3_X2 U9995 ( .A1(n4637), .A2(n42154), .A3(n7829), .ZN(n7828) );
  OAI21_X2 U28633 ( .A1(n64510), .A2(n8537), .B(n42786), .ZN(n42191) );
  NAND2_X2 U1833 ( .A1(n16962), .A2(n3505), .ZN(n40102) );
  NAND2_X2 U8005 ( .A1(n33016), .A2(n36545), .ZN(n33022) );
  OAI21_X2 U9382 ( .A1(n36543), .A2(n36541), .B(n36542), .ZN(n33016) );
  INV_X2 U4430 ( .I(n863), .ZN(n59282) );
  NAND2_X2 U32876 ( .A1(n34626), .A2(n12859), .ZN(n23117) );
  BUF_X4 U51687 ( .I(n18385), .Z(n61066) );
  NAND2_X2 U5008 ( .A1(n42140), .A2(n43254), .ZN(n42128) );
  INV_X1 U32442 ( .I(n1197), .ZN(n12419) );
  INV_X4 U26898 ( .I(n60969), .ZN(n53590) );
  INV_X4 U18712 ( .I(n34316), .ZN(n34324) );
  NOR2_X2 U42095 ( .A1(n60488), .A2(n11549), .ZN(n55014) );
  AOI21_X2 U17000 ( .A1(n13466), .A2(n23420), .B(n22027), .ZN(n13467) );
  OAI22_X2 U28258 ( .A1(n8619), .A2(n43341), .B1(n22446), .B2(n8185), .ZN(
        n42162) );
  INV_X2 U54500 ( .I(n56403), .ZN(n56250) );
  INV_X8 U11154 ( .I(n4547), .ZN(n1391) );
  AOI21_X2 U12805 ( .A1(n11361), .A2(n16377), .B(n19454), .ZN(n9503) );
  NAND3_X2 U17066 ( .A1(n39874), .A2(n39873), .A3(n39872), .ZN(n39875) );
  INV_X4 U57182 ( .I(n25231), .ZN(n48654) );
  NAND2_X2 U21392 ( .A1(n4659), .A2(n11476), .ZN(n42014) );
  INV_X2 U1059 ( .I(n46026), .ZN(n46871) );
  NAND2_X2 U36445 ( .A1(n36990), .A2(n37212), .ZN(n37208) );
  NAND2_X2 U41247 ( .A1(n21623), .A2(n49767), .ZN(n49772) );
  NAND2_X2 U2335 ( .A1(n10907), .A2(n461), .ZN(n13647) );
  NAND2_X2 U35315 ( .A1(n93), .A2(n28072), .ZN(n24817) );
  NAND3_X1 U16916 ( .A1(n54596), .A2(n54589), .A3(n64681), .ZN(n3664) );
  INV_X2 U1903 ( .I(n41805), .ZN(n1401) );
  NOR2_X2 U9741 ( .A1(n26568), .A2(n9661), .ZN(n16981) );
  NAND2_X2 U8360 ( .A1(n23488), .A2(n61743), .ZN(n43910) );
  NAND2_X2 U52583 ( .A1(n46016), .A2(n20666), .ZN(n47305) );
  INV_X1 U37681 ( .I(n38300), .ZN(n39437) );
  BUF_X2 U6161 ( .I(n26127), .Z(n60633) );
  NAND2_X2 U4643 ( .A1(n18252), .A2(n11153), .ZN(n49090) );
  NAND2_X2 U26826 ( .A1(n23030), .A2(n56775), .ZN(n56749) );
  INV_X2 U9291 ( .I(n7365), .ZN(n44956) );
  BUF_X2 U13205 ( .I(n14010), .Z(n4351) );
  NAND2_X2 U40361 ( .A1(n43564), .A2(n42620), .ZN(n43552) );
  INV_X2 U33960 ( .I(n25378), .ZN(n52541) );
  BUF_X4 U1320 ( .I(n11417), .Z(n25895) );
  OR2_X2 U43681 ( .A1(n18482), .A2(n43693), .Z(n4229) );
  OAI21_X2 U818 ( .A1(n58551), .A2(n58550), .B(n49412), .ZN(n5210) );
  NOR4_X2 U38496 ( .A1(n17612), .A2(n47808), .A3(n47702), .A4(n17611), .ZN(
        n17484) );
  NAND2_X2 U7595 ( .A1(n16823), .A2(n62357), .ZN(n58484) );
  AOI22_X2 U7144 ( .A1(n39116), .A2(n38046), .B1(n40946), .B2(n40110), .ZN(
        n7314) );
  NAND2_X2 U1668 ( .A1(n43897), .A2(n20183), .ZN(n43231) );
  INV_X2 U5699 ( .I(n49799), .ZN(n47346) );
  INV_X8 U10878 ( .I(n50427), .ZN(n1380) );
  NAND2_X2 U3935 ( .A1(n13191), .A2(n10309), .ZN(n28269) );
  NAND2_X2 U1972 ( .A1(n41496), .A2(n58693), .ZN(n12503) );
  NOR2_X2 U882 ( .A1(n49355), .A2(n50044), .ZN(n49359) );
  INV_X2 U36798 ( .I(n42067), .ZN(n42966) );
  INV_X2 U32020 ( .I(n56323), .ZN(n11841) );
  BUF_X4 U11563 ( .I(n23215), .Z(n19364) );
  NOR2_X2 U13643 ( .A1(n35777), .A2(n16736), .ZN(n33920) );
  NAND3_X2 U34701 ( .A1(n15477), .A2(n26626), .A3(n18751), .ZN(n27554) );
  INV_X4 U13160 ( .I(n1409), .ZN(n7641) );
  NOR2_X2 U42781 ( .A1(n48360), .A2(n16986), .ZN(n48927) );
  NOR2_X2 U2626 ( .A1(n34130), .A2(n22598), .ZN(n33657) );
  NAND3_X2 U22201 ( .A1(n48767), .A2(n48766), .A3(n49283), .ZN(n3594) );
  INV_X2 U33 ( .I(n55878), .ZN(n1585) );
  INV_X2 U3848 ( .I(n9281), .ZN(n3150) );
  INV_X8 U12956 ( .I(n20922), .ZN(n1500) );
  NAND2_X2 U54797 ( .A1(n54318), .A2(n22372), .ZN(n54499) );
  INV_X2 U4869 ( .I(n43361), .ZN(n60351) );
  BUF_X2 U5096 ( .I(n55884), .Z(n15717) );
  NAND2_X2 U40844 ( .A1(n55597), .A2(n55569), .ZN(n55573) );
  OAI21_X2 U26699 ( .A1(n54981), .A2(n52564), .B(n61065), .ZN(n7668) );
  BUF_X4 U17469 ( .I(n39095), .Z(n22786) );
  NAND2_X2 U914 ( .A1(n1377), .A2(n49882), .ZN(n50289) );
  INV_X4 U41940 ( .I(n57109), .ZN(n23538) );
  NAND2_X2 U9634 ( .A1(n14138), .A2(n22524), .ZN(n35907) );
  INV_X2 U11643 ( .I(n16403), .ZN(n35778) );
  INV_X2 U13201 ( .I(n38453), .ZN(n39736) );
  INV_X4 U29273 ( .I(n21489), .ZN(n9304) );
  NAND2_X2 U9637 ( .A1(n29933), .A2(n30812), .ZN(n29934) );
  INV_X2 U3859 ( .I(n29929), .ZN(n29933) );
  NOR2_X1 U37567 ( .A1(n59888), .A2(n59887), .ZN(n43663) );
  INV_X2 U26569 ( .I(n6888), .ZN(n24373) );
  OAI21_X2 U14840 ( .A1(n8058), .A2(n8057), .B(n55262), .ZN(n8056) );
  INV_X2 U38928 ( .I(n15731), .ZN(n60076) );
  NAND2_X2 U20796 ( .A1(n18294), .A2(n2524), .ZN(n55303) );
  NOR2_X2 U1787 ( .A1(n5512), .A2(n5514), .ZN(n5511) );
  AOI21_X2 U16645 ( .A1(n21664), .A2(n21666), .B(n15020), .ZN(n43276) );
  NAND2_X2 U7280 ( .A1(n2735), .A2(n19591), .ZN(n21664) );
  INV_X2 U29861 ( .I(n41186), .ZN(n40667) );
  NOR2_X2 U8684 ( .A1(n30027), .A2(n23315), .ZN(n27734) );
  INV_X2 U10609 ( .I(n65217), .ZN(n3729) );
  NAND3_X2 U3760 ( .A1(n27791), .A2(n7450), .A3(n10580), .ZN(n58386) );
  NAND3_X2 U20604 ( .A1(n4211), .A2(n27738), .A3(n2374), .ZN(n21795) );
  NOR2_X2 U684 ( .A1(n49266), .A2(n49267), .ZN(n7383) );
  OAI21_X2 U33542 ( .A1(n24099), .A2(n65062), .B(n24354), .ZN(n45367) );
  INV_X2 U39947 ( .I(n6789), .ZN(n53288) );
  INV_X2 U10023 ( .I(n7418), .ZN(n13458) );
  NAND2_X2 U4503 ( .A1(n53384), .A2(n25047), .ZN(n53605) );
  NAND2_X2 U3515 ( .A1(n35307), .A2(n22797), .ZN(n35811) );
  NAND2_X2 U3497 ( .A1(n34676), .A2(n1813), .ZN(n34522) );
  NAND2_X2 U32550 ( .A1(n43258), .A2(n43995), .ZN(n43712) );
  AOI21_X1 U7044 ( .A1(n42550), .A2(n42549), .B(n59309), .ZN(n10107) );
  INV_X2 U27726 ( .I(n12634), .ZN(n10229) );
  CLKBUF_X4 U5387 ( .I(n25994), .Z(n58250) );
  INV_X2 U784 ( .I(n48053), .ZN(n49071) );
  NOR2_X2 U679 ( .A1(n58722), .A2(n10244), .ZN(n58540) );
  INV_X8 U30355 ( .I(n6052), .ZN(n23577) );
  BUF_X4 U1763 ( .I(n42104), .Z(n1718) );
  NAND2_X2 U19262 ( .A1(n21486), .A2(n29819), .ZN(n30317) );
  INV_X1 U2435 ( .I(n10079), .ZN(n17407) );
  INV_X4 U33762 ( .I(n14630), .ZN(n22386) );
  NAND2_X2 U36296 ( .A1(n57015), .A2(n21569), .ZN(n57108) );
  OAI22_X2 U36098 ( .A1(n47821), .A2(n45569), .B1(n45570), .B2(n45969), .ZN(
        n17570) );
  NAND2_X2 U4406 ( .A1(n52487), .A2(n14927), .ZN(n15100) );
  INV_X2 U1281 ( .I(n20340), .ZN(n21820) );
  INV_X2 U14185 ( .I(n57412), .ZN(n10458) );
  INV_X2 U40418 ( .I(n22925), .ZN(n20447) );
  BUF_X2 U27352 ( .I(n12299), .Z(n11318) );
  NOR2_X1 U13243 ( .A1(n10966), .A2(n10965), .ZN(n10964) );
  INV_X2 U41468 ( .I(n22190), .ZN(n28072) );
  NAND2_X1 U8844 ( .A1(n9391), .A2(n34730), .ZN(n9390) );
  NAND2_X2 U29333 ( .A1(n21489), .A2(n24934), .ZN(n36719) );
  NOR2_X2 U50778 ( .A1(n40923), .A2(n7201), .ZN(n40936) );
  INV_X4 U17546 ( .I(n25377), .ZN(n37745) );
  INV_X4 U8081 ( .I(n28690), .ZN(n5631) );
  NAND2_X2 U36547 ( .A1(n27120), .A2(n22735), .ZN(n28360) );
  NAND2_X2 U8617 ( .A1(n9758), .A2(n6497), .ZN(n45734) );
  NAND2_X2 U1600 ( .A1(n43243), .A2(n1333), .ZN(n9063) );
  INV_X4 U29884 ( .I(n20897), .ZN(n14518) );
  NOR2_X2 U11645 ( .A1(n34626), .A2(n4075), .ZN(n4716) );
  NOR2_X2 U48248 ( .A1(n1422), .A2(n36070), .ZN(n36312) );
  AND2_X2 U3600 ( .A1(n15687), .A2(n15318), .Z(n22597) );
  INV_X2 U36275 ( .I(n55896), .ZN(n55855) );
  AOI21_X2 U783 ( .A1(n24135), .A2(n60209), .B(n49991), .ZN(n61184) );
  INV_X4 U34200 ( .I(n1316), .ZN(n30375) );
  AOI22_X2 U56486 ( .A1(n56273), .A2(n56272), .B1(n56271), .B2(n56270), .ZN(
        n56274) );
  NAND2_X2 U10380 ( .A1(n42140), .A2(n42666), .ZN(n42138) );
  AND2_X2 U38807 ( .A1(n10485), .A2(n36746), .Z(n23648) );
  NOR2_X2 U186 ( .A1(n55345), .A2(n15703), .ZN(n5087) );
  NAND4_X2 U2462 ( .A1(n35267), .A2(n35266), .A3(n35265), .A4(n35264), .ZN(
        n36332) );
  BUF_X4 U2085 ( .I(n42651), .Z(n11039) );
  BUF_X4 U19938 ( .I(Key[113]), .Z(n55395) );
  BUF_X4 U14307 ( .I(Key[186]), .Z(n57096) );
  NAND2_X2 U1987 ( .A1(n42427), .A2(n42432), .ZN(n42446) );
  BUF_X4 U6149 ( .I(n33568), .Z(n59681) );
  NOR2_X2 U52359 ( .A1(n45165), .A2(n48882), .ZN(n49764) );
  INV_X4 U1210 ( .I(n20912), .ZN(n18227) );
  NAND2_X2 U22696 ( .A1(n20156), .A2(n22114), .ZN(n53238) );
  NAND2_X2 U30950 ( .A1(n22201), .A2(n53860), .ZN(n15362) );
  INV_X4 U23083 ( .I(n58324), .ZN(n61673) );
  NOR2_X2 U35745 ( .A1(n22801), .A2(n461), .ZN(n20501) );
  NAND3_X2 U23365 ( .A1(n30475), .A2(n26707), .A3(n29816), .ZN(n29542) );
  NAND2_X2 U4993 ( .A1(n17350), .A2(n64283), .ZN(n33965) );
  NOR2_X2 U9566 ( .A1(n34080), .A2(n34628), .ZN(n17350) );
  INV_X4 U24040 ( .I(n5243), .ZN(n24949) );
  NAND2_X2 U3355 ( .A1(n58961), .A2(n16264), .ZN(n35830) );
  INV_X1 U1573 ( .I(n43478), .ZN(n18722) );
  NAND2_X2 U9563 ( .A1(n22559), .A2(n3856), .ZN(n11027) );
  INV_X2 U986 ( .I(n49676), .ZN(n49687) );
  NAND2_X2 U48609 ( .A1(n35827), .A2(n35826), .ZN(n35828) );
  INV_X4 U8025 ( .I(n41020), .ZN(n37529) );
  BUF_X2 U15186 ( .I(n52443), .Z(n19847) );
  AND2_X2 U7931 ( .A1(n24870), .A2(n8023), .Z(n22947) );
  NOR2_X2 U8894 ( .A1(n29783), .A2(n28938), .ZN(n29255) );
  NAND2_X2 U9009 ( .A1(n27622), .A2(n22643), .ZN(n27613) );
  INV_X4 U11523 ( .I(n65061), .ZN(n49089) );
  NOR2_X2 U3325 ( .A1(n27622), .A2(n63100), .ZN(n26669) );
  INV_X2 U2041 ( .I(n14732), .ZN(n40644) );
  NOR2_X2 U10953 ( .A1(n47844), .A2(n47828), .ZN(n47837) );
  NAND2_X2 U53527 ( .A1(n57949), .A2(n24332), .ZN(n49390) );
  INV_X2 U1804 ( .I(n8619), .ZN(n43606) );
  BUF_X2 U6460 ( .I(n15804), .Z(n60370) );
  NAND2_X1 U16642 ( .A1(n42164), .A2(n42163), .ZN(n21862) );
  NAND2_X2 U32498 ( .A1(n22169), .A2(n13799), .ZN(n21615) );
  INV_X4 U26340 ( .I(n64683), .ZN(n23407) );
  NOR2_X2 U9494 ( .A1(n37426), .A2(n2383), .ZN(n35517) );
  INV_X2 U57171 ( .I(n42846), .ZN(n43736) );
  INV_X2 U8186 ( .I(n15189), .ZN(n37686) );
  NAND2_X2 U20210 ( .A1(n39959), .A2(n18396), .ZN(n2081) );
  NOR3_X2 U4499 ( .A1(n53533), .A2(n23047), .A3(n13370), .ZN(n53391) );
  INV_X2 U37761 ( .I(n37549), .ZN(n38364) );
  INV_X2 U9043 ( .I(n11226), .ZN(n14229) );
  NOR2_X2 U48383 ( .A1(n1793), .A2(n37049), .ZN(n35103) );
  INV_X2 U13675 ( .I(n35252), .ZN(n35759) );
  INV_X4 U32004 ( .I(n43601), .ZN(n41624) );
  INV_X4 U8636 ( .I(n45768), .ZN(n1267) );
  INV_X2 U5162 ( .I(n47252), .ZN(n21793) );
  BUF_X2 U19877 ( .I(n27159), .Z(n20721) );
  BUF_X2 U853 ( .I(n687), .Z(n64) );
  AOI21_X2 U51096 ( .A1(n41526), .A2(n42698), .B(n42383), .ZN(n41527) );
  AOI22_X2 U51638 ( .A1(n43545), .A2(n43544), .B1(n43543), .B2(n43542), .ZN(
        n43546) );
  NAND2_X2 U51635 ( .A1(n43538), .A2(n43540), .ZN(n43544) );
  NAND2_X2 U21289 ( .A1(n18834), .A2(n2899), .ZN(n35706) );
  NOR2_X2 U11038 ( .A1(n45208), .A2(n45207), .ZN(n45571) );
  NAND3_X2 U28325 ( .A1(n8242), .A2(n36523), .A3(n36585), .ZN(n8239) );
  NOR2_X1 U41296 ( .A1(n21711), .A2(n21710), .ZN(n21709) );
  NAND2_X2 U9840 ( .A1(n9721), .A2(n35887), .ZN(n35900) );
  INV_X4 U30907 ( .I(n20743), .ZN(n28625) );
  NOR2_X2 U4486 ( .A1(n18724), .A2(n23557), .ZN(n43295) );
  INV_X2 U9474 ( .I(n36269), .ZN(n36347) );
  NOR2_X2 U42867 ( .A1(n28615), .A2(n28606), .ZN(n28436) );
  NOR3_X1 U43995 ( .A1(n26318), .A2(n26611), .A3(n26317), .ZN(n26332) );
  INV_X2 U38927 ( .I(n14819), .ZN(n60075) );
  NAND2_X2 U2439 ( .A1(n10126), .A2(n41183), .ZN(n40487) );
  NAND2_X2 U28048 ( .A1(n60028), .A2(n60030), .ZN(n7980) );
  NAND2_X2 U20434 ( .A1(n58004), .A2(n58669), .ZN(n13235) );
  INV_X1 U1298 ( .I(n16993), .ZN(n45532) );
  NAND4_X1 U30033 ( .A1(n60539), .A2(n49989), .A3(n18585), .A4(n60209), .ZN(
        n59076) );
  BUF_X4 U20580 ( .I(n17892), .Z(n2362) );
  NOR2_X2 U32600 ( .A1(n36852), .A2(n36846), .ZN(n36010) );
  INV_X1 U8028 ( .I(n25320), .ZN(n49318) );
  NAND3_X2 U20631 ( .A1(n22453), .A2(n58040), .A3(n58039), .ZN(n17796) );
  INV_X2 U5175 ( .I(n13963), .ZN(n13961) );
  NAND3_X2 U55992 ( .A1(n61348), .A2(n22777), .A3(n42042), .ZN(n42043) );
  NAND2_X2 U5319 ( .A1(n18138), .A2(n47729), .ZN(n15336) );
  NAND2_X2 U7248 ( .A1(n43410), .A2(n43624), .ZN(n60837) );
  INV_X1 U9337 ( .I(n12378), .ZN(n41545) );
  NAND2_X2 U8864 ( .A1(n34146), .A2(n59626), .ZN(n9169) );
  NAND3_X1 U32434 ( .A1(n12398), .A2(n56904), .A3(n12397), .ZN(n12396) );
  NAND2_X2 U2422 ( .A1(n26243), .A2(n7118), .ZN(n35346) );
  NOR3_X2 U8873 ( .A1(n31075), .A2(n31076), .A3(n61382), .ZN(n14423) );
  INV_X2 U12658 ( .I(n14473), .ZN(n11899) );
  OAI22_X1 U33303 ( .A1(n29859), .A2(n1838), .B1(n13517), .B2(n17413), .ZN(
        n29861) );
  INV_X2 U42538 ( .I(n1545), .ZN(n34952) );
  NOR3_X2 U27393 ( .A1(n7430), .A2(n25850), .A3(n7429), .ZN(n9493) );
  NAND3_X2 U5676 ( .A1(n60063), .A2(n22213), .A3(n25283), .ZN(n25282) );
  NOR2_X2 U13841 ( .A1(n2430), .A2(n16612), .ZN(n16611) );
  NOR2_X2 U12587 ( .A1(n47398), .A2(n47397), .ZN(n47855) );
  BUF_X4 U23695 ( .I(n43726), .Z(n47435) );
  BUF_X8 U4898 ( .I(n47873), .Z(n49377) );
  AND2_X2 U1590 ( .A1(n16850), .A2(n1502), .Z(n775) );
  NOR2_X2 U2381 ( .A1(n21536), .A2(n4541), .ZN(n6830) );
  BUF_X4 U27710 ( .I(n50035), .Z(n54035) );
  INV_X2 U7138 ( .I(n40132), .ZN(n14018) );
  INV_X4 U26254 ( .I(n10737), .ZN(n11359) );
  NAND2_X2 U273 ( .A1(n55948), .A2(n56409), .ZN(n55964) );
  OAI22_X2 U25080 ( .A1(n9451), .A2(n9452), .B1(n9453), .B2(n47359), .ZN(
        n60093) );
  INV_X2 U2131 ( .I(n37158), .ZN(n38382) );
  NOR2_X2 U2316 ( .A1(n6831), .A2(n37359), .ZN(n36758) );
  INV_X2 U27376 ( .I(n47725), .ZN(n47717) );
  NAND2_X2 U1165 ( .A1(n45762), .A2(n6290), .ZN(n45773) );
  OAI21_X2 U2495 ( .A1(n32463), .A2(n31658), .B(n31657), .ZN(n16888) );
  NAND3_X2 U49957 ( .A1(n41197), .A2(n41188), .A3(n61407), .ZN(n40734) );
  NOR2_X2 U8663 ( .A1(n57454), .A2(n23928), .ZN(n42024) );
  NAND4_X2 U28479 ( .A1(n38415), .A2(n38416), .A3(n10587), .A4(n39069), .ZN(
        n5302) );
  OAI21_X2 U1819 ( .A1(n39417), .A2(n7392), .B(n21074), .ZN(n6435) );
  AOI21_X2 U40595 ( .A1(n36653), .A2(n36654), .B(n20724), .ZN(n21074) );
  NAND2_X2 U2881 ( .A1(n37945), .A2(n1244), .ZN(n37091) );
  OAI21_X2 U11524 ( .A1(n7028), .A2(n20060), .B(n36777), .ZN(n35417) );
  BUF_X4 U5649 ( .I(n49384), .Z(n57949) );
  INV_X4 U1761 ( .I(n6601), .ZN(n20844) );
  NAND2_X2 U41228 ( .A1(n60601), .A2(n12028), .ZN(n9022) );
  NAND3_X2 U3127 ( .A1(n57847), .A2(n35150), .A3(n35138), .ZN(n5107) );
  NAND3_X2 U28978 ( .A1(n11844), .A2(n11843), .A3(n8963), .ZN(n11890) );
  INV_X4 U41136 ( .I(n22717), .ZN(n50304) );
  AOI21_X2 U11410 ( .A1(n35559), .A2(n35558), .B(n15940), .ZN(n16604) );
  INV_X4 U985 ( .I(n21071), .ZN(n49074) );
  BUF_X2 U10848 ( .I(n46122), .Z(n10255) );
  INV_X4 U7585 ( .I(n25826), .ZN(n35031) );
  NAND2_X2 U37159 ( .A1(n16543), .A2(n16336), .ZN(n16542) );
  INV_X2 U4896 ( .I(n47873), .ZN(n49542) );
  NOR2_X2 U37307 ( .A1(n54340), .A2(n62102), .ZN(n53885) );
  INV_X2 U2669 ( .I(n157), .ZN(n34128) );
  NAND3_X2 U10687 ( .A1(n4971), .A2(n3006), .A3(n3007), .ZN(n2999) );
  NAND2_X2 U11594 ( .A1(n3707), .A2(n64406), .ZN(n15826) );
  NAND3_X2 U27049 ( .A1(n12469), .A2(n56370), .A3(n56660), .ZN(n12720) );
  NAND2_X1 U10811 ( .A1(n14309), .A2(n14310), .ZN(n7154) );
  INV_X2 U40810 ( .I(n25403), .ZN(n25004) );
  NAND2_X2 U11861 ( .A1(n18871), .A2(n28663), .ZN(n18872) );
  INV_X2 U20954 ( .I(n24243), .ZN(n23928) );
  AOI21_X2 U3517 ( .A1(n37451), .A2(n12457), .B(n37455), .ZN(n12456) );
  INV_X2 U45540 ( .I(n31274), .ZN(n29921) );
  NAND2_X2 U2347 ( .A1(n14004), .A2(n63303), .ZN(n41514) );
  NAND2_X2 U10272 ( .A1(n36821), .A2(n16501), .ZN(n37408) );
  AOI21_X2 U26512 ( .A1(n7531), .A2(n22909), .B(n6829), .ZN(n35244) );
  NAND2_X2 U4973 ( .A1(n54307), .A2(n64832), .ZN(n54308) );
  NAND2_X2 U6532 ( .A1(n60376), .A2(n60375), .ZN(n17952) );
  NAND2_X2 U13907 ( .A1(n29207), .A2(n61383), .ZN(n28934) );
  OAI21_X2 U8493 ( .A1(n28596), .A2(n28595), .B(n19712), .ZN(n28597) );
  INV_X2 U19822 ( .I(n19619), .ZN(n26061) );
  INV_X4 U435 ( .I(n57470), .ZN(n1602) );
  INV_X2 U15859 ( .I(n48218), .ZN(n47546) );
  INV_X4 U34857 ( .I(n31097), .ZN(n26084) );
  NOR2_X2 U10555 ( .A1(n6083), .A2(n13192), .ZN(n13191) );
  BUF_X4 U44130 ( .I(n56886), .Z(n60708) );
  NOR2_X2 U53446 ( .A1(n48323), .A2(n5629), .ZN(n48449) );
  BUF_X4 U19941 ( .I(Key[174]), .Z(n56827) );
  INV_X4 U27030 ( .I(n25522), .ZN(n52768) );
  INV_X2 U32446 ( .I(n17156), .ZN(n34136) );
  INV_X1 U9734 ( .I(n14212), .ZN(n28477) );
  NAND3_X2 U3203 ( .A1(n2176), .A2(n28271), .A3(n62631), .ZN(n28024) );
  NOR2_X2 U38162 ( .A1(n22416), .A2(n24196), .ZN(n16920) );
  INV_X4 U1147 ( .I(n50378), .ZN(n5283) );
  NOR4_X2 U56547 ( .A1(n56460), .A2(n56459), .A3(n56457), .A4(n56458), .ZN(
        n56470) );
  NAND2_X2 U23167 ( .A1(n39070), .A2(n40643), .ZN(n11386) );
  NAND2_X2 U37035 ( .A1(n697), .A2(n48076), .ZN(n47119) );
  AOI21_X1 U36011 ( .A1(n17115), .A2(n20315), .B(n27925), .ZN(n17114) );
  NAND2_X2 U1368 ( .A1(n13296), .A2(n45888), .ZN(n10976) );
  NOR3_X2 U30019 ( .A1(n18286), .A2(n18285), .A3(n18288), .ZN(n18284) );
  INV_X2 U1451 ( .I(n47696), .ZN(n47800) );
  INV_X2 U9458 ( .I(n33404), .ZN(n32463) );
  NOR2_X2 U4224 ( .A1(n56703), .A2(n23785), .ZN(n56688) );
  NAND3_X2 U53309 ( .A1(n47589), .A2(n47588), .A3(n47587), .ZN(n47601) );
  INV_X4 U27488 ( .I(n22683), .ZN(n55231) );
  INV_X2 U12071 ( .I(n11375), .ZN(n54345) );
  NOR2_X2 U4005 ( .A1(n13688), .A2(n37543), .ZN(n44850) );
  INV_X4 U16184 ( .I(n9505), .ZN(n6523) );
  AOI22_X2 U15441 ( .A1(n34084), .A2(n11992), .B1(n4075), .B2(n33960), .ZN(
        n33962) );
  INV_X4 U600 ( .I(n59294), .ZN(n56370) );
  BUF_X4 U11192 ( .I(n10970), .Z(n1393) );
  NAND2_X2 U17009 ( .A1(n18713), .A2(n40155), .ZN(n3361) );
  INV_X4 U32069 ( .I(n43254), .ZN(n21376) );
  NAND2_X2 U4186 ( .A1(n56629), .A2(n51450), .ZN(n56623) );
  BUF_X4 U16887 ( .I(n62535), .Z(n16447) );
  NAND4_X2 U6282 ( .A1(n56308), .A2(n56305), .A3(n56307), .A4(n56306), .ZN(
        n58776) );
  NOR3_X2 U45571 ( .A1(n52733), .A2(n19181), .A3(n60779), .ZN(n60788) );
  NAND2_X2 U30925 ( .A1(n22463), .A2(n22462), .ZN(n24385) );
  OAI21_X2 U51305 ( .A1(n42217), .A2(n42216), .B(n42528), .ZN(n42218) );
  INV_X2 U3956 ( .I(n27880), .ZN(n26798) );
  INV_X4 U26631 ( .I(n8453), .ZN(n24188) );
  INV_X2 U10922 ( .I(n45730), .ZN(n45733) );
  NOR2_X2 U4120 ( .A1(n45734), .A2(n46944), .ZN(n45730) );
  INV_X1 U9041 ( .I(n29142), .ZN(n17489) );
  NOR2_X2 U13158 ( .A1(n8051), .A2(n16402), .ZN(n35314) );
  NOR2_X2 U43456 ( .A1(n60895), .A2(n31079), .ZN(n30562) );
  NAND2_X2 U49134 ( .A1(n37403), .A2(n37402), .ZN(n37415) );
  OAI21_X2 U4084 ( .A1(n56775), .A2(n56806), .B(n23879), .ZN(n56792) );
  NOR2_X2 U6092 ( .A1(n61088), .A2(n34266), .ZN(n60258) );
  BUF_X4 U8364 ( .I(n57738), .Z(n19000) );
  NOR2_X2 U904 ( .A1(n49074), .A2(n7990), .ZN(n48302) );
  BUF_X4 U38175 ( .I(n55216), .Z(n16943) );
  INV_X2 U541 ( .I(n53226), .ZN(n16427) );
  INV_X2 U2198 ( .I(n65150), .ZN(n59280) );
  INV_X2 U16273 ( .I(n45726), .ZN(n47774) );
  INV_X2 U8747 ( .I(n39118), .ZN(n41003) );
  NOR2_X2 U24162 ( .A1(n14712), .A2(n14711), .ZN(n14710) );
  NOR3_X2 U40789 ( .A1(n28425), .A2(n64867), .A3(n29580), .ZN(n28423) );
  OAI21_X2 U47562 ( .A1(n35388), .A2(n63484), .B(n4802), .ZN(n32856) );
  NOR2_X1 U55465 ( .A1(n54033), .A2(n53558), .ZN(n53559) );
  INV_X2 U214 ( .I(n18652), .ZN(n54198) );
  INV_X2 U1331 ( .I(n1039), .ZN(n25582) );
  AOI21_X2 U24186 ( .A1(n34625), .A2(n5135), .B(n5134), .ZN(n5133) );
  NOR2_X2 U11612 ( .A1(n64132), .A2(n4716), .ZN(n5135) );
  BUF_X2 U11739 ( .I(n11236), .Z(n26202) );
  INV_X2 U5243 ( .I(n1265), .ZN(n9152) );
  BUF_X4 U1069 ( .I(n49500), .Z(n6704) );
  BUF_X4 U26995 ( .I(n15731), .Z(n109) );
  AND2_X2 U5223 ( .A1(n25467), .A2(n13288), .Z(n53598) );
  INV_X2 U27551 ( .I(n29456), .ZN(n29458) );
  INV_X4 U34869 ( .I(n18875), .ZN(n22936) );
  NAND2_X2 U12354 ( .A1(n7747), .A2(n7746), .ZN(n7745) );
  NAND2_X2 U5132 ( .A1(n46973), .A2(n49057), .ZN(n48068) );
  NOR3_X2 U17714 ( .A1(n36283), .A2(n36282), .A3(n14172), .ZN(n36284) );
  NAND3_X2 U11998 ( .A1(n54436), .A2(n4783), .A3(n54605), .ZN(n54957) );
  AOI21_X2 U4210 ( .A1(n54204), .A2(n26008), .B(n14643), .ZN(n54127) );
  OR2_X2 U36817 ( .A1(n26097), .A2(n54615), .Z(n25792) );
  NAND2_X2 U1448 ( .A1(n47576), .A2(n1669), .ZN(n45590) );
  INV_X2 U21094 ( .I(n53009), .ZN(n53006) );
  NAND2_X2 U12151 ( .A1(n52488), .A2(n12696), .ZN(n55434) );
  INV_X2 U176 ( .I(n21389), .ZN(n9551) );
  BUF_X4 U5275 ( .I(n49779), .Z(n21550) );
  INV_X1 U10954 ( .I(n47810), .ZN(n12495) );
  NAND3_X2 U4933 ( .A1(n34128), .A2(n33390), .A3(n19538), .ZN(n34144) );
  NOR2_X2 U27587 ( .A1(n49465), .A2(n49459), .ZN(n49224) );
  INV_X2 U6416 ( .I(n43131), .ZN(n23541) );
  NOR2_X2 U10688 ( .A1(n42567), .A2(n41766), .ZN(n42889) );
  INV_X2 U5133 ( .I(n49057), .ZN(n2047) );
  AOI21_X2 U24948 ( .A1(n7537), .A2(n12768), .B(n5264), .ZN(n7536) );
  NOR2_X2 U1124 ( .A1(n49904), .A2(n49901), .ZN(n47075) );
  OR2_X2 U1449 ( .A1(n24216), .A2(n21518), .Z(n16244) );
  OAI21_X2 U26161 ( .A1(n64667), .A2(n35762), .B(n61547), .ZN(n18393) );
  INV_X2 U2490 ( .I(n37388), .ZN(n8520) );
  INV_X2 U1094 ( .I(n58313), .ZN(n46948) );
  NAND3_X2 U1697 ( .A1(n60725), .A2(n9031), .A3(n60724), .ZN(n8481) );
  NAND2_X2 U10317 ( .A1(n1795), .A2(n34661), .ZN(n7731) );
  NOR2_X2 U4930 ( .A1(n24405), .A2(n15784), .ZN(n6297) );
  NAND2_X2 U10032 ( .A1(n7031), .A2(n63747), .ZN(n7033) );
  INV_X4 U6388 ( .I(n40934), .ZN(n40257) );
  OAI21_X2 U17087 ( .A1(n41119), .A2(n11587), .B(n39993), .ZN(n11586) );
  INV_X2 U7531 ( .I(n48097), .ZN(n21304) );
  INV_X4 U29357 ( .I(n47669), .ZN(n11599) );
  INV_X2 U5323 ( .I(n36377), .ZN(n36566) );
  INV_X4 U34849 ( .I(n24646), .ZN(n56600) );
  BUF_X4 U10884 ( .I(n50218), .Z(n1383) );
  NOR2_X2 U53448 ( .A1(n48323), .A2(n49013), .ZN(n48040) );
  AOI21_X2 U32637 ( .A1(n15966), .A2(n56396), .B(n12555), .ZN(n12554) );
  NAND2_X2 U38688 ( .A1(n61472), .A2(n62760), .ZN(n54637) );
  BUF_X4 U16384 ( .I(n25961), .Z(n7202) );
  AOI22_X2 U10808 ( .A1(n44664), .A2(n48736), .B1(n44668), .B2(n60730), .ZN(
        n19743) );
  NAND2_X1 U33706 ( .A1(n55027), .A2(n55026), .ZN(n14101) );
  INV_X2 U2053 ( .I(n11664), .ZN(n1725) );
  INV_X2 U43331 ( .I(n25063), .ZN(n32516) );
  INV_X1 U3601 ( .I(n12768), .ZN(n33652) );
  INV_X2 U43431 ( .I(n48514), .ZN(n48504) );
  NAND2_X2 U11913 ( .A1(n22817), .A2(n10983), .ZN(n11177) );
  INV_X2 U24669 ( .I(n30213), .ZN(n30215) );
  BUF_X4 U8583 ( .I(n14019), .Z(n23487) );
  AOI21_X2 U6355 ( .A1(n55663), .A2(n55662), .B(n11682), .ZN(n58249) );
  CLKBUF_X12 U4449 ( .I(n20893), .Z(n10457) );
  INV_X4 U39015 ( .I(n15780), .ZN(n18247) );
  INV_X4 U9776 ( .I(n764), .ZN(n13704) );
  NOR2_X2 U30896 ( .A1(n13142), .A2(n16043), .ZN(n16149) );
  BUF_X2 U12102 ( .I(Key[119]), .Z(n55603) );
  NAND2_X1 U5697 ( .A1(n58095), .A2(n58094), .ZN(n45667) );
  OAI21_X2 U53354 ( .A1(n47739), .A2(n47738), .B(n47737), .ZN(n47740) );
  NAND2_X1 U23163 ( .A1(n35144), .A2(n4368), .ZN(n33717) );
  INV_X2 U19317 ( .I(n30754), .ZN(n30753) );
  BUF_X4 U474 ( .I(n15777), .Z(n21957) );
  NOR2_X2 U1330 ( .A1(n46976), .A2(n14875), .ZN(n45740) );
  INV_X4 U30835 ( .I(n4734), .ZN(n50296) );
  NOR2_X2 U1537 ( .A1(n47154), .A2(n2634), .ZN(n2633) );
  NOR2_X2 U9256 ( .A1(n46976), .A2(n11250), .ZN(n45519) );
  AOI21_X2 U14611 ( .A1(n20489), .A2(n20156), .B(n20487), .ZN(n20486) );
  NAND2_X2 U36505 ( .A1(n36331), .A2(n37404), .ZN(n22462) );
  NAND2_X2 U35868 ( .A1(n24556), .A2(n63394), .ZN(n16517) );
  OAI21_X1 U33139 ( .A1(n59516), .A2(n577), .B(n660), .ZN(n40456) );
  NOR2_X2 U51238 ( .A1(n42317), .A2(n5261), .ZN(n43010) );
  INV_X2 U1295 ( .I(n45074), .ZN(n47307) );
  NAND2_X1 U24119 ( .A1(n41991), .A2(n41990), .ZN(n14754) );
  AOI21_X2 U7324 ( .A1(n57014), .A2(n14756), .B(n21655), .ZN(n10379) );
  NAND2_X2 U31708 ( .A1(n1421), .A2(n36944), .ZN(n35433) );
  NOR2_X2 U23506 ( .A1(n18046), .A2(n12851), .ZN(n18042) );
  NOR2_X2 U44580 ( .A1(n29150), .A2(n22482), .ZN(n27260) );
  OAI21_X2 U5827 ( .A1(n5853), .A2(n10807), .B(n22112), .ZN(n60100) );
  OAI21_X1 U50564 ( .A1(n40094), .A2(n40129), .B(n42494), .ZN(n39885) );
  NAND2_X2 U38781 ( .A1(n50364), .A2(n59633), .ZN(n48228) );
  BUF_X4 U10366 ( .I(n18088), .Z(n9085) );
  INV_X1 U4969 ( .I(n33391), .ZN(n34143) );
  NOR2_X2 U7176 ( .A1(n42180), .A2(n42784), .ZN(n39087) );
  NOR2_X2 U1940 ( .A1(n38672), .A2(n5488), .ZN(n8536) );
  NOR4_X2 U54129 ( .A1(n50364), .A2(n50363), .A3(n50362), .A4(n23394), .ZN(
        n50365) );
  NAND2_X2 U3553 ( .A1(n60808), .A2(n3363), .ZN(n32872) );
  INV_X2 U12628 ( .I(n47325), .ZN(n46066) );
  OAI21_X2 U9725 ( .A1(n1308), .A2(n10061), .B(n3622), .ZN(n9598) );
  NAND2_X1 U18330 ( .A1(n4964), .A2(n25634), .ZN(n33440) );
  INV_X2 U9611 ( .I(n35429), .ZN(n14282) );
  NOR3_X1 U23717 ( .A1(n20235), .A2(n13229), .A3(n20285), .ZN(n8189) );
  NAND2_X2 U1224 ( .A1(n44065), .A2(n58174), .ZN(n46976) );
  NAND2_X2 U3008 ( .A1(n29773), .A2(n13943), .ZN(n29767) );
  NOR2_X1 U12035 ( .A1(n12856), .A2(n28517), .ZN(n27715) );
  INV_X2 U1715 ( .I(n20601), .ZN(n42896) );
  AOI21_X2 U12199 ( .A1(n55682), .A2(n55681), .B(n11805), .ZN(n24959) );
  NAND3_X2 U27306 ( .A1(n8362), .A2(n28888), .A3(n28889), .ZN(n28890) );
  NAND2_X2 U16476 ( .A1(n43038), .A2(n43035), .ZN(n22131) );
  NAND2_X1 U13523 ( .A1(n35794), .A2(n24956), .ZN(n34294) );
  NOR2_X2 U33603 ( .A1(n2674), .A2(n21592), .ZN(n33118) );
  NAND2_X2 U9839 ( .A1(n35159), .A2(n36487), .ZN(n35560) );
  NOR2_X2 U29724 ( .A1(n36238), .A2(n36483), .ZN(n35159) );
  BUF_X4 U22704 ( .I(n20625), .Z(n4030) );
  NAND2_X2 U4680 ( .A1(n36202), .A2(n9372), .ZN(n36207) );
  CLKBUF_X8 U40709 ( .I(n57126), .Z(n21570) );
  INV_X2 U51710 ( .I(n44004), .ZN(n49393) );
  OAI21_X2 U18964 ( .A1(n8269), .A2(n8268), .B(n8267), .ZN(n8266) );
  AOI21_X2 U38538 ( .A1(n17554), .A2(n17553), .B(n57023), .ZN(n21577) );
  AOI22_X2 U37268 ( .A1(n1601), .A2(n21706), .B1(n63339), .B2(n57030), .ZN(
        n17554) );
  NAND2_X2 U39373 ( .A1(n40720), .A2(n3245), .ZN(n60128) );
  INV_X2 U21787 ( .I(n3247), .ZN(n15215) );
  NAND2_X2 U27702 ( .A1(n62334), .A2(n1473), .ZN(n47932) );
  NAND2_X2 U9825 ( .A1(n4838), .A2(n19968), .ZN(n19977) );
  NAND2_X2 U51543 ( .A1(n43200), .A2(n43199), .ZN(n46337) );
  BUF_X4 U34794 ( .I(n15631), .Z(n15630) );
  BUF_X4 U8783 ( .I(n29456), .Z(n23224) );
  INV_X2 U8944 ( .I(n29000), .ZN(n28115) );
  NOR3_X2 U47867 ( .A1(n33752), .A2(n1545), .A3(n1345), .ZN(n34570) );
  INV_X2 U6303 ( .I(n517), .ZN(n2564) );
  BUF_X2 U18158 ( .I(n24864), .Z(n10110) );
  NOR3_X1 U25544 ( .A1(n58681), .A2(n60210), .A3(n27926), .ZN(n17524) );
  NAND2_X2 U8889 ( .A1(n21228), .A2(n21227), .ZN(n6152) );
  NAND2_X2 U7768 ( .A1(n59360), .A2(n35073), .ZN(n10211) );
  OAI21_X2 U9818 ( .A1(n35070), .A2(n36334), .B(n23648), .ZN(n59360) );
  NAND3_X2 U25951 ( .A1(n46803), .A2(n24428), .A3(n47082), .ZN(n58727) );
  NAND2_X2 U4201 ( .A1(n50096), .A2(n1473), .ZN(n47924) );
  NAND2_X2 U10232 ( .A1(n58307), .A2(n1515), .ZN(n16749) );
  NAND2_X2 U41254 ( .A1(n21622), .A2(n21621), .ZN(n49768) );
  INV_X2 U28090 ( .I(n16936), .ZN(n32638) );
  BUF_X4 U40969 ( .I(n57075), .Z(n21079) );
  NOR2_X2 U32317 ( .A1(n41350), .A2(n60583), .ZN(n43079) );
  NAND2_X2 U3170 ( .A1(n1785), .A2(n1339), .ZN(n35534) );
  NOR2_X2 U37230 ( .A1(n22788), .A2(n49172), .ZN(n49570) );
  NAND3_X2 U12951 ( .A1(n14950), .A2(n14948), .A3(n21349), .ZN(n8658) );
  BUF_X2 U102 ( .I(n53351), .Z(n60517) );
  AOI21_X2 U9263 ( .A1(n34178), .A2(n34161), .B(n34168), .ZN(n34162) );
  OAI22_X2 U4654 ( .A1(n45935), .A2(n45599), .B1(n46014), .B2(n47297), .ZN(
        n60250) );
  INV_X2 U48431 ( .I(n35204), .ZN(n35628) );
  NOR2_X2 U48430 ( .A1(n22428), .A2(n35203), .ZN(n35204) );
  AOI21_X2 U17025 ( .A1(n40769), .A2(n62272), .B(n40768), .ZN(n40775) );
  INV_X8 U24203 ( .I(n23215), .ZN(n25261) );
  BUF_X2 U17475 ( .I(n15616), .Z(n11264) );
  INV_X8 U42514 ( .I(n24949), .ZN(n29511) );
  INV_X2 U2145 ( .I(n16120), .ZN(n39690) );
  NAND2_X2 U21478 ( .A1(n28054), .A2(n23209), .ZN(n27136) );
  NAND2_X2 U39087 ( .A1(n1644), .A2(n48688), .ZN(n48071) );
  NOR2_X2 U28269 ( .A1(n18483), .A2(n1407), .ZN(n39510) );
  INV_X2 U1429 ( .I(n59818), .ZN(n46930) );
  NAND3_X2 U44511 ( .A1(n28325), .A2(n27144), .A3(n27143), .ZN(n27145) );
  INV_X4 U4121 ( .I(n1643), .ZN(n8251) );
  OR3_X2 U18401 ( .A1(n35341), .A2(n24934), .A3(n36202), .Z(n36728) );
  NOR2_X1 U17161 ( .A1(n18669), .A2(n40753), .ZN(n18665) );
  INV_X1 U15970 ( .I(n47655), .ZN(n47656) );
  NOR2_X2 U39130 ( .A1(n54646), .A2(n54645), .ZN(n54695) );
  INV_X2 U12243 ( .I(n55099), .ZN(n59538) );
  INV_X1 U14014 ( .I(n31051), .ZN(n30696) );
  OAI21_X2 U11687 ( .A1(n34069), .A2(n7534), .B(n33720), .ZN(n34990) );
  NAND2_X2 U53980 ( .A1(n9003), .A2(n56268), .ZN(n61192) );
  NAND2_X2 U37090 ( .A1(n47670), .A2(n7395), .ZN(n24894) );
  AOI22_X2 U4420 ( .A1(n48010), .A2(n5463), .B1(n49096), .B2(n48009), .ZN(
        n48016) );
  BUF_X4 U14304 ( .I(Key[148]), .Z(n51261) );
  BUF_X4 U19915 ( .I(Key[102]), .Z(n52970) );
  INV_X2 U8941 ( .I(n29063), .ZN(n17268) );
  NAND2_X2 U10557 ( .A1(n9908), .A2(n22044), .ZN(n26253) );
  NAND2_X2 U9210 ( .A1(n9225), .A2(n25128), .ZN(n22788) );
  NOR2_X2 U18692 ( .A1(n33719), .A2(n33720), .ZN(n34988) );
  INV_X2 U342 ( .I(n13800), .ZN(n52695) );
  INV_X8 U7194 ( .I(n42607), .ZN(n8799) );
  NOR2_X2 U53675 ( .A1(n1261), .A2(n48847), .ZN(n48848) );
  AOI22_X2 U2382 ( .A1(n8797), .A2(n36106), .B1(n41037), .B2(n57791), .ZN(
        n57846) );
  AOI22_X1 U36925 ( .A1(n43337), .A2(n41624), .B1(n43335), .B2(n22446), .ZN(
        n41631) );
  NAND2_X2 U35332 ( .A1(n21478), .A2(n28989), .ZN(n30030) );
  NOR3_X2 U6967 ( .A1(n61035), .A2(n18497), .A3(n28281), .ZN(n21601) );
  INV_X2 U12245 ( .I(n52672), .ZN(n52860) );
  NAND2_X2 U13424 ( .A1(n37404), .A2(n36831), .ZN(n11008) );
  NAND2_X2 U16441 ( .A1(n7449), .A2(n42752), .ZN(n7448) );
  NAND2_X2 U5685 ( .A1(n48151), .A2(n48548), .ZN(n46800) );
  INV_X4 U28824 ( .I(n17615), .ZN(n25396) );
  INV_X4 U871 ( .I(n23707), .ZN(n50373) );
  INV_X4 U22613 ( .I(n13174), .ZN(n28989) );
  NAND4_X1 U47560 ( .A1(n32852), .A2(n32851), .A3(n32850), .A4(n32849), .ZN(
        n32853) );
  NAND2_X1 U15308 ( .A1(n14033), .A2(n14032), .ZN(n14031) );
  NAND2_X2 U29985 ( .A1(n33362), .A2(n34155), .ZN(n34151) );
  NOR2_X2 U11892 ( .A1(n25013), .A2(n6316), .ZN(n31163) );
  INV_X2 U899 ( .I(n17523), .ZN(n1376) );
  OR2_X1 U4225 ( .A1(n15817), .A2(n10475), .Z(n1072) );
  NAND3_X2 U3186 ( .A1(n21632), .A2(n21631), .A3(n15976), .ZN(n21630) );
  INV_X2 U10269 ( .I(n34849), .ZN(n36781) );
  INV_X4 U8786 ( .I(n60878), .ZN(n2310) );
  NAND3_X2 U36393 ( .A1(n35670), .A2(n24006), .A3(n24286), .ZN(n35673) );
  INV_X4 U28503 ( .I(n35723), .ZN(n37210) );
  AOI21_X2 U7867 ( .A1(n59570), .A2(n37227), .B(n37225), .ZN(n37228) );
  INV_X2 U10901 ( .I(n44627), .ZN(n60877) );
  NOR3_X2 U31288 ( .A1(n15370), .A2(n59973), .A3(n20648), .ZN(n4042) );
  INV_X2 U48733 ( .I(n37211), .ZN(n36265) );
  BUF_X4 U27997 ( .I(n21205), .Z(n16765) );
  INV_X2 U1253 ( .I(n18361), .ZN(n1648) );
  NOR2_X2 U26978 ( .A1(n52548), .A2(n55418), .ZN(n54981) );
  INV_X2 U37673 ( .I(n48721), .ZN(n21822) );
  INV_X2 U5710 ( .I(n45751), .ZN(n59384) );
  NOR2_X1 U12162 ( .A1(n8325), .A2(n7989), .ZN(n7988) );
  BUF_X4 U2155 ( .I(n39737), .Z(n15644) );
  NAND2_X2 U55133 ( .A1(n52672), .A2(n52671), .ZN(n52676) );
  NAND2_X2 U37308 ( .A1(n56606), .A2(n24647), .ZN(n22967) );
  INV_X4 U39070 ( .I(n18333), .ZN(n23420) );
  NAND3_X2 U24618 ( .A1(n6583), .A2(n49713), .A3(n49714), .ZN(n49715) );
  NAND3_X1 U16540 ( .A1(n16474), .A2(n22844), .A3(n16472), .ZN(n40690) );
  BUF_X4 U42237 ( .I(Key[69]), .Z(n23093) );
  BUF_X4 U26725 ( .I(n54239), .Z(n1256) );
  INV_X2 U224 ( .I(n54032), .ZN(n54199) );
  NAND2_X2 U5192 ( .A1(n36493), .A2(n32691), .ZN(n36485) );
  NAND2_X2 U3512 ( .A1(n61647), .A2(n9329), .ZN(n35631) );
  INV_X4 U1259 ( .I(n44779), .ZN(n22326) );
  INV_X2 U39146 ( .I(n48422), .ZN(n46969) );
  NAND2_X2 U806 ( .A1(n20458), .A2(n49063), .ZN(n49062) );
  NAND2_X1 U23732 ( .A1(n60815), .A2(n60813), .ZN(n60812) );
  NAND2_X2 U10675 ( .A1(n9724), .A2(n41794), .ZN(n23623) );
  OAI21_X2 U6866 ( .A1(n11099), .A2(n16151), .B(n12057), .ZN(n40789) );
  NOR2_X2 U27509 ( .A1(n8781), .A2(n36898), .ZN(n35451) );
  NOR2_X2 U8445 ( .A1(n27494), .A2(n1575), .ZN(n26965) );
  AOI21_X2 U11213 ( .A1(n6659), .A2(n57488), .B(n57487), .ZN(n391) );
  NOR2_X2 U2334 ( .A1(n41257), .A2(n7728), .ZN(n12057) );
  NAND2_X2 U11002 ( .A1(n45503), .A2(n13258), .ZN(n44344) );
  INV_X2 U361 ( .I(n21643), .ZN(n21655) );
  BUF_X2 U5795 ( .I(n22283), .Z(n57677) );
  NOR3_X2 U23236 ( .A1(n59472), .A2(n1098), .A3(n59471), .ZN(n58349) );
  OAI21_X2 U9819 ( .A1(n22621), .A2(n22620), .B(n56229), .ZN(n22619) );
  INV_X2 U51282 ( .I(n42148), .ZN(n42154) );
  NOR2_X2 U9340 ( .A1(n23561), .A2(n42155), .ZN(n43602) );
  INV_X2 U11738 ( .I(n22336), .ZN(n25063) );
  NAND2_X2 U6578 ( .A1(n2692), .A2(n6203), .ZN(n5947) );
  INV_X2 U32417 ( .I(n63854), .ZN(n25368) );
  NOR2_X2 U7206 ( .A1(n42158), .A2(n42585), .ZN(n43610) );
  BUF_X4 U10309 ( .I(n9274), .Z(n1339) );
  NOR2_X2 U34860 ( .A1(n26052), .A2(n63430), .ZN(n37277) );
  OR2_X2 U41978 ( .A1(n38134), .A2(n26110), .Z(n42215) );
  INV_X2 U1326 ( .I(n46824), .ZN(n47378) );
  INV_X1 U18762 ( .I(n32308), .ZN(n13507) );
  BUF_X4 U7540 ( .I(n15713), .Z(n23157) );
  INV_X2 U2756 ( .I(n9971), .ZN(n13583) );
  OAI21_X1 U11587 ( .A1(n4164), .A2(n4163), .B(n4162), .ZN(n4165) );
  NOR3_X1 U23740 ( .A1(n34371), .A2(n34005), .A3(n34006), .ZN(n60388) );
  NAND2_X2 U13142 ( .A1(n41473), .A2(n40755), .ZN(n38765) );
  INV_X2 U11462 ( .I(n36211), .ZN(n1766) );
  INV_X2 U16855 ( .I(n8425), .ZN(n42689) );
  AOI21_X2 U48380 ( .A1(n35079), .A2(n35078), .B(n37311), .ZN(n35084) );
  NOR2_X2 U1704 ( .A1(n43980), .A2(n6007), .ZN(n43258) );
  INV_X2 U21536 ( .I(n8391), .ZN(n14969) );
  OR2_X2 U1377 ( .A1(n19160), .A2(n60935), .Z(n18099) );
  INV_X4 U42670 ( .I(n23416), .ZN(n48521) );
  AND3_X2 U32807 ( .A1(n48851), .A2(n48850), .A3(n1374), .Z(n12750) );
  NAND2_X2 U40748 ( .A1(n30333), .A2(n30408), .ZN(n30409) );
  OAI21_X1 U53093 ( .A1(n46860), .A2(n24578), .B(n46859), .ZN(n46861) );
  NAND2_X1 U56241 ( .A1(n55675), .A2(n58626), .ZN(n55683) );
  INV_X2 U29209 ( .I(n25594), .ZN(n45376) );
  NAND2_X2 U4807 ( .A1(n27958), .A2(n28270), .ZN(n28018) );
  NAND2_X2 U13234 ( .A1(n36347), .A2(n23449), .ZN(n35722) );
  NOR3_X2 U52541 ( .A1(n60510), .A2(n23156), .A3(n11058), .ZN(n45545) );
  NAND2_X1 U710 ( .A1(n19445), .A2(n58096), .ZN(n49618) );
  INV_X4 U13259 ( .I(n22044), .ZN(n18497) );
  OAI21_X2 U2874 ( .A1(n1783), .A2(n1243), .B(n37945), .ZN(n15442) );
  INV_X4 U15030 ( .I(n21877), .ZN(n52958) );
  NAND2_X1 U7759 ( .A1(n36643), .A2(n58069), .ZN(n36646) );
  NAND2_X2 U4636 ( .A1(n13627), .A2(n11781), .ZN(n11615) );
  NOR2_X2 U10440 ( .A1(n28981), .A2(n13817), .ZN(n29260) );
  NAND3_X2 U45189 ( .A1(n1317), .A2(n23734), .A3(n29576), .ZN(n28981) );
  INV_X4 U511 ( .I(n52768), .ZN(n21082) );
  NOR3_X2 U31507 ( .A1(n36560), .A2(n20166), .A3(n20167), .ZN(n61122) );
  BUF_X4 U11565 ( .I(n36768), .Z(n20060) );
  BUF_X4 U13430 ( .I(n35178), .Z(n10067) );
  NAND3_X2 U2846 ( .A1(n30434), .A2(n30433), .A3(n30432), .ZN(n31425) );
  AOI21_X1 U12880 ( .A1(n43077), .A2(n41350), .B(n22695), .ZN(n10991) );
  NAND2_X2 U37296 ( .A1(n25648), .A2(n54597), .ZN(n54084) );
  CLKBUF_X4 U5359 ( .I(n21856), .Z(n2408) );
  BUF_X4 U16292 ( .I(n45411), .Z(n23934) );
  NOR2_X1 U29499 ( .A1(n61127), .A2(n61126), .ZN(n12745) );
  NAND2_X2 U7362 ( .A1(n1577), .A2(n53738), .ZN(n53763) );
  INV_X2 U8799 ( .I(n35901), .ZN(n35896) );
  NAND2_X2 U36219 ( .A1(n48929), .A2(n48367), .ZN(n25562) );
  NAND3_X2 U15655 ( .A1(n5302), .A2(n59315), .A3(n59252), .ZN(n57629) );
  NAND2_X2 U19054 ( .A1(n14647), .A2(n23176), .ZN(n14852) );
  NAND2_X2 U39071 ( .A1(n18333), .A2(n23698), .ZN(n18338) );
  NAND2_X2 U6419 ( .A1(n54957), .A2(n54956), .ZN(n10032) );
  NAND4_X1 U27075 ( .A1(n22497), .A2(n55224), .A3(n17155), .A4(n55225), .ZN(
        n55227) );
  NAND2_X2 U10712 ( .A1(n51256), .A2(n50883), .ZN(n22621) );
  NOR2_X2 U53374 ( .A1(n47789), .A2(n47788), .ZN(n47790) );
  INV_X4 U31167 ( .I(n12497), .ZN(n15825) );
  INV_X4 U2804 ( .I(n31461), .ZN(n19886) );
  NOR3_X2 U44623 ( .A1(n19967), .A2(n58108), .A3(n29321), .ZN(n27355) );
  INV_X4 U4582 ( .I(n22142), .ZN(n2367) );
  OAI21_X2 U9171 ( .A1(n9232), .A2(n9234), .B(n18271), .ZN(n23342) );
  INV_X4 U30131 ( .I(n22701), .ZN(n33319) );
  NAND4_X2 U20307 ( .A1(n48370), .A2(n48372), .A3(n48371), .A4(n48373), .ZN(
        n51510) );
  NAND3_X2 U10018 ( .A1(n41656), .A2(n25327), .A3(n43581), .ZN(n23692) );
  NOR2_X2 U403 ( .A1(n64657), .A2(n20982), .ZN(n57006) );
  NOR2_X2 U36598 ( .A1(n28270), .A2(n61021), .ZN(n28277) );
  NAND3_X2 U35753 ( .A1(n34823), .A2(n36040), .A3(n61066), .ZN(n36038) );
  INV_X1 U11451 ( .I(n61728), .ZN(n13554) );
  AND2_X2 U12278 ( .A1(n54481), .A2(n51779), .Z(n16043) );
  NOR2_X2 U37272 ( .A1(n54340), .A2(n1611), .ZN(n54022) );
  INV_X2 U42827 ( .I(n40570), .ZN(n41106) );
  NOR2_X2 U10998 ( .A1(n47329), .A2(n7389), .ZN(n47315) );
  NOR2_X2 U37332 ( .A1(n55914), .A2(n55721), .ZN(n51884) );
  INV_X2 U15120 ( .I(n5167), .ZN(n21361) );
  OAI21_X2 U11403 ( .A1(n8816), .A2(n63742), .B(n3471), .ZN(n7338) );
  INV_X2 U1749 ( .I(n41966), .ZN(n43570) );
  NAND3_X2 U36577 ( .A1(n57792), .A2(n28541), .A3(n27871), .ZN(n27254) );
  BUF_X4 U3070 ( .I(n37034), .Z(n60659) );
  INV_X2 U26025 ( .I(n28933), .ZN(n1863) );
  NOR2_X2 U9251 ( .A1(n34957), .A2(n5529), .ZN(n12169) );
  AOI22_X1 U32738 ( .A1(n31466), .A2(n14107), .B1(n31468), .B2(n59458), .ZN(
        n31475) );
  NOR2_X2 U27150 ( .A1(n46910), .A2(n44774), .ZN(n46918) );
  INV_X2 U33105 ( .I(n35490), .ZN(n1773) );
  BUF_X4 U5664 ( .I(n36158), .Z(n324) );
  BUF_X8 U15675 ( .I(n16590), .Z(n14561) );
  OAI22_X2 U29562 ( .A1(n43606), .A2(n43605), .B1(n62299), .B2(n42160), .ZN(
        n42159) );
  INV_X4 U31297 ( .I(n22236), .ZN(n35272) );
  NOR2_X1 U36147 ( .A1(n59791), .A2(n21236), .ZN(n16453) );
  INV_X2 U13438 ( .I(n10811), .ZN(n42288) );
  INV_X1 U4735 ( .I(n10391), .ZN(n38942) );
  NAND3_X2 U7062 ( .A1(n34384), .A2(n18771), .A3(n35276), .ZN(n15450) );
  AND2_X2 U12000 ( .A1(n7975), .A2(n27533), .Z(n7974) );
  NAND2_X2 U2362 ( .A1(n6830), .A2(n22659), .ZN(n37117) );
  INV_X4 U6220 ( .I(n57620), .ZN(n30492) );
  INV_X4 U31365 ( .I(n30338), .ZN(n59268) );
  INV_X2 U3629 ( .I(n24388), .ZN(n33159) );
  BUF_X4 U5262 ( .I(n15746), .Z(n15728) );
  AOI22_X2 U11104 ( .A1(n46789), .A2(n46790), .B1(n46788), .B2(n47101), .ZN(
        n11344) );
  NOR2_X2 U30525 ( .A1(n24364), .A2(n48555), .ZN(n46790) );
  NAND2_X2 U1685 ( .A1(n15029), .A2(n15160), .ZN(n41583) );
  NAND2_X2 U485 ( .A1(n5008), .A2(n53009), .ZN(n7027) );
  INV_X1 U32239 ( .I(n36233), .ZN(n36232) );
  INV_X4 U56769 ( .I(n57433), .ZN(n57132) );
  NOR2_X2 U36357 ( .A1(n23947), .A2(n1547), .ZN(n34178) );
  NOR2_X2 U5955 ( .A1(n2979), .A2(n2982), .ZN(n409) );
  OAI21_X2 U5588 ( .A1(n2980), .A2(n49634), .B(n15826), .ZN(n2979) );
  NAND2_X2 U938 ( .A1(n3738), .A2(n24362), .ZN(n49634) );
  INV_X2 U1625 ( .I(n44155), .ZN(n60133) );
  BUF_X2 U3641 ( .I(n37987), .Z(n23280) );
  NAND2_X2 U39531 ( .A1(n157), .A2(n33663), .ZN(n32699) );
  NAND2_X2 U43659 ( .A1(n23030), .A2(n56809), .ZN(n56773) );
  NOR3_X1 U23772 ( .A1(n17472), .A2(n41207), .A3(n17471), .ZN(n17470) );
  NAND2_X2 U28988 ( .A1(n15020), .A2(n1493), .ZN(n8981) );
  BUF_X4 U6535 ( .I(n49732), .Z(n22764) );
  INV_X2 U24325 ( .I(n40090), .ZN(n9980) );
  INV_X4 U13309 ( .I(n60209), .ZN(n50364) );
  NOR2_X2 U35768 ( .A1(n36515), .A2(n37369), .ZN(n36600) );
  INV_X2 U41784 ( .I(n55020), .ZN(n54641) );
  INV_X4 U41322 ( .I(n56547), .ZN(n56530) );
  NAND3_X1 U20283 ( .A1(n10073), .A2(n12916), .A3(n42546), .ZN(n57979) );
  NOR2_X2 U1933 ( .A1(n42370), .A2(n43438), .ZN(n43428) );
  INV_X4 U20243 ( .I(n7580), .ZN(n30195) );
  NOR2_X2 U10733 ( .A1(n42759), .A2(n43380), .ZN(n43377) );
  BUF_X2 U13197 ( .I(n15275), .Z(n4667) );
  INV_X2 U41411 ( .I(n37818), .ZN(n39776) );
  NOR2_X1 U48136 ( .A1(n60882), .A2(n36709), .ZN(n35351) );
  INV_X4 U5298 ( .I(n11989), .ZN(n59647) );
  NOR2_X2 U13426 ( .A1(n36842), .A2(n36841), .ZN(n36843) );
  NAND2_X2 U20246 ( .A1(n30192), .A2(n364), .ZN(n30198) );
  INV_X4 U2556 ( .I(n33720), .ZN(n34513) );
  NAND3_X2 U25924 ( .A1(n34990), .A2(n63444), .A3(n58472), .ZN(n13898) );
  NOR2_X2 U48515 ( .A1(n35483), .A2(n35996), .ZN(n37958) );
  NAND2_X2 U2415 ( .A1(n60437), .A2(n12652), .ZN(n35444) );
  NAND2_X2 U27037 ( .A1(n19557), .A2(n19558), .ZN(n49863) );
  AOI21_X2 U37096 ( .A1(n22694), .A2(n826), .B(n49940), .ZN(n16867) );
  NAND2_X2 U48450 ( .A1(n35273), .A2(n20736), .ZN(n35274) );
  NOR2_X2 U36891 ( .A1(n43043), .A2(n12962), .ZN(n43044) );
  NOR3_X2 U2343 ( .A1(n59016), .A2(n23884), .A3(n59015), .ZN(n39074) );
  NOR2_X2 U4264 ( .A1(n39066), .A2(n25424), .ZN(n3636) );
  INV_X4 U2984 ( .I(n60111), .ZN(n17627) );
  OR2_X2 U37297 ( .A1(n64738), .A2(n54067), .Z(n54065) );
  INV_X2 U43480 ( .I(n8794), .ZN(n48584) );
  NOR2_X2 U6561 ( .A1(n60879), .A2(n61677), .ZN(n5580) );
  NAND2_X2 U1676 ( .A1(n7754), .A2(n43452), .ZN(n46495) );
  NOR2_X2 U7742 ( .A1(n36375), .A2(n58520), .ZN(n58519) );
  NAND2_X2 U24206 ( .A1(n47054), .A2(n10563), .ZN(n11642) );
  NAND2_X1 U1513 ( .A1(n42092), .A2(n43553), .ZN(n17064) );
  NOR2_X2 U12397 ( .A1(n1261), .A2(n48845), .ZN(n48004) );
  INV_X2 U34971 ( .I(n18891), .ZN(n24886) );
  INV_X4 U39237 ( .I(n25467), .ZN(n53384) );
  INV_X2 U596 ( .I(n51268), .ZN(n18195) );
  NAND2_X2 U2693 ( .A1(n1817), .A2(n6001), .ZN(n35747) );
  NAND2_X2 U2345 ( .A1(n22801), .A2(n37249), .ZN(n20951) );
  NOR2_X2 U11337 ( .A1(n58587), .A2(n2867), .ZN(n41884) );
  BUF_X4 U7680 ( .I(n2867), .Z(n2325) );
  INV_X2 U5905 ( .I(n33570), .ZN(n33097) );
  INV_X2 U17263 ( .I(n40207), .ZN(n10741) );
  INV_X2 U3050 ( .I(n36163), .ZN(n36514) );
  INV_X2 U28465 ( .I(n47411), .ZN(n47691) );
  INV_X2 U3235 ( .I(n28329), .ZN(n27025) );
  BUF_X4 U5053 ( .I(n23610), .Z(n1405) );
  INV_X2 U25540 ( .I(n52281), .ZN(n56372) );
  NOR2_X2 U6695 ( .A1(n61136), .A2(n23409), .ZN(n3739) );
  OAI22_X2 U31104 ( .A1(n16664), .A2(n35865), .B1(n16663), .B2(n35423), .ZN(
        n16662) );
  NAND2_X2 U3281 ( .A1(n8478), .A2(n1926), .ZN(n27410) );
  BUF_X4 U41787 ( .I(n36960), .Z(n60437) );
  AOI21_X1 U15785 ( .A1(n27258), .A2(n57652), .B(n29153), .ZN(n9584) );
  OAI21_X2 U12996 ( .A1(n19387), .A2(n60653), .B(n64377), .ZN(n10876) );
  NAND2_X2 U6507 ( .A1(n49622), .A2(n14122), .ZN(n52569) );
  NOR2_X2 U39664 ( .A1(n21577), .A2(n21727), .ZN(n19280) );
  BUF_X4 U27319 ( .I(n45373), .Z(n23668) );
  AOI21_X2 U8412 ( .A1(n4511), .A2(n402), .B(n5715), .ZN(n15402) );
  INV_X2 U35493 ( .I(n44523), .ZN(n23305) );
  INV_X2 U17426 ( .I(n41882), .ZN(n41881) );
  OR2_X2 U8875 ( .A1(n34627), .A2(n31508), .Z(n15819) );
  INV_X2 U27047 ( .I(n18590), .ZN(n47743) );
  BUF_X4 U41898 ( .I(n37351), .Z(n22659) );
  NOR2_X2 U6097 ( .A1(n2288), .A2(n59329), .ZN(n24506) );
  NOR2_X2 U3756 ( .A1(n29220), .A2(n9426), .ZN(n30723) );
  BUF_X4 U19908 ( .I(Key[178]), .Z(n56879) );
  INV_X1 U13436 ( .I(n23585), .ZN(n36288) );
  INV_X2 U25175 ( .I(n15247), .ZN(n24300) );
  INV_X2 U7311 ( .I(n1288), .ZN(n18435) );
  NOR2_X2 U12806 ( .A1(n14262), .A2(n14261), .ZN(n14260) );
  NAND2_X2 U6455 ( .A1(n60708), .A2(n56867), .ZN(n56895) );
  NOR2_X2 U25485 ( .A1(n41597), .A2(n5802), .ZN(n43871) );
  NAND2_X2 U11119 ( .A1(n15044), .A2(n43868), .ZN(n5802) );
  AND2_X1 U8235 ( .A1(n24815), .A2(n13174), .Z(n13087) );
  INV_X2 U17848 ( .I(n37019), .ZN(n35089) );
  NAND2_X2 U20798 ( .A1(n58059), .A2(n42947), .ZN(n11517) );
  NAND2_X2 U4911 ( .A1(n56499), .A2(n59444), .ZN(n56498) );
  INV_X4 U3666 ( .I(n24848), .ZN(n56436) );
  INV_X2 U14930 ( .I(n55296), .ZN(n4838) );
  NOR3_X1 U631 ( .A1(n15602), .A2(n15601), .A3(n61679), .ZN(n15599) );
  NAND2_X2 U50817 ( .A1(n42854), .A2(n40553), .ZN(n45823) );
  NAND2_X2 U7192 ( .A1(n6007), .A2(n5571), .ZN(n43977) );
  NOR3_X2 U41556 ( .A1(n5884), .A2(n5887), .A3(n5885), .ZN(n60387) );
  NAND2_X2 U9013 ( .A1(n22214), .A2(n29691), .ZN(n27887) );
  OAI21_X2 U1287 ( .A1(n22899), .A2(n16493), .B(n47502), .ZN(n57625) );
  INV_X2 U2127 ( .I(n38848), .ZN(n38411) );
  BUF_X4 U12931 ( .I(n462), .Z(n5261) );
  INV_X1 U1747 ( .I(n42113), .ZN(n60274) );
  INV_X2 U9084 ( .I(n25856), .ZN(n33150) );
  INV_X2 U37996 ( .I(n30994), .ZN(n59938) );
  NOR2_X2 U22620 ( .A1(n11659), .A2(n3939), .ZN(n34421) );
  NAND2_X2 U41653 ( .A1(n6498), .A2(n19938), .ZN(n42265) );
  BUF_X4 U5723 ( .I(n1293), .Z(n58018) );
  INV_X4 U1158 ( .I(n47610), .ZN(n1295) );
  CLKBUF_X4 U41772 ( .I(n3566), .Z(n22502) );
  NAND4_X2 U13618 ( .A1(n33973), .A2(n63116), .A3(n34589), .A4(n33972), .ZN(
        n9540) );
  INV_X2 U8014 ( .I(n33511), .ZN(n34545) );
  CLKBUF_X8 U5185 ( .I(n16460), .Z(n12521) );
  NAND2_X2 U3465 ( .A1(n34351), .A2(n57164), .ZN(n57734) );
  INV_X4 U3607 ( .I(n17671), .ZN(n17795) );
  NOR2_X2 U33456 ( .A1(n48080), .A2(n10250), .ZN(n48084) );
  INV_X4 U7607 ( .I(n26147), .ZN(n36777) );
  INV_X4 U31065 ( .I(n45897), .ZN(n47670) );
  INV_X4 U2043 ( .I(n42502), .ZN(n13169) );
  NAND2_X2 U999 ( .A1(n15021), .A2(n49918), .ZN(n48386) );
  OR2_X1 U19463 ( .A1(n248), .A2(n55727), .Z(n52393) );
  BUF_X2 U12115 ( .I(Key[5]), .Z(n53124) );
  BUF_X4 U8089 ( .I(n32870), .Z(n59769) );
  BUF_X4 U19943 ( .I(Key[149]), .Z(n56202) );
  BUF_X4 U13564 ( .I(n14328), .Z(n14251) );
  NAND2_X1 U36951 ( .A1(n29416), .A2(n29415), .ZN(n18160) );
  INV_X2 U20894 ( .I(n24908), .ZN(n32505) );
  NOR2_X1 U31729 ( .A1(n28894), .A2(n7426), .ZN(n30005) );
  NOR2_X1 U16948 ( .A1(n13600), .A2(n16469), .ZN(n13599) );
  INV_X4 U42214 ( .I(n30311), .ZN(n31224) );
  INV_X4 U22286 ( .I(n65274), .ZN(n8381) );
  INV_X4 U989 ( .I(n9225), .ZN(n49166) );
  NAND2_X2 U44846 ( .A1(n27913), .A2(n30084), .ZN(n28786) );
  INV_X4 U32267 ( .I(n17411), .ZN(n12164) );
  AOI21_X2 U41386 ( .A1(n260), .A2(n59633), .B(n64562), .ZN(n50362) );
  INV_X2 U9138 ( .I(n3127), .ZN(n8446) );
  OAI22_X2 U52917 ( .A1(n48462), .A2(n10626), .B1(n48460), .B2(n7186), .ZN(
        n46454) );
  INV_X2 U1096 ( .I(n15749), .ZN(n48462) );
  NOR2_X2 U11544 ( .A1(n20174), .A2(n50400), .ZN(n18142) );
  INV_X1 U10312 ( .I(n13493), .ZN(n60548) );
  INV_X2 U7840 ( .I(n6157), .ZN(n7579) );
  CLKBUF_X4 U5339 ( .I(n30895), .Z(n242) );
  AOI21_X1 U56040 ( .A1(n55159), .A2(n55158), .B(n55168), .ZN(n55160) );
  INV_X2 U8980 ( .I(n29795), .ZN(n30084) );
  AOI22_X2 U20920 ( .A1(n46175), .A2(n2634), .B1(n4655), .B2(n46483), .ZN(
        n13472) );
  OAI22_X2 U18931 ( .A1(n30091), .A2(n30090), .B1(n30089), .B2(n30088), .ZN(
        n15622) );
  INV_X2 U3921 ( .I(n48975), .ZN(n25474) );
  NAND2_X2 U1998 ( .A1(n1725), .A2(n8523), .ZN(n7951) );
  INV_X2 U14849 ( .I(n5604), .ZN(n2924) );
  NOR2_X1 U7382 ( .A1(n40564), .A2(n40565), .ZN(n57773) );
  INV_X1 U2025 ( .I(n25247), .ZN(n286) );
  NAND2_X2 U43746 ( .A1(n32941), .A2(n60667), .ZN(n34218) );
  INV_X2 U28185 ( .I(n49325), .ZN(n10456) );
  INV_X1 U1539 ( .I(n22283), .ZN(n1667) );
  NAND2_X1 U20022 ( .A1(n7568), .A2(n7569), .ZN(n58396) );
  BUF_X2 U7604 ( .I(n9806), .Z(n2383) );
  BUF_X4 U7702 ( .I(n9337), .Z(n2557) );
  NOR3_X2 U12377 ( .A1(n48369), .A2(n49280), .A3(n48368), .ZN(n48370) );
  OAI21_X2 U43246 ( .A1(n14884), .A2(n24473), .B(n56436), .ZN(n56437) );
  BUF_X4 U5024 ( .I(n35852), .Z(n37249) );
  INV_X2 U2665 ( .I(n3148), .ZN(n2346) );
  NAND2_X1 U257 ( .A1(n24013), .A2(n51872), .ZN(n54257) );
  INV_X2 U482 ( .I(n51860), .ZN(n51866) );
  OAI21_X2 U8001 ( .A1(n1537), .A2(n11423), .B(n34951), .ZN(n58195) );
  INV_X1 U4723 ( .I(n63007), .ZN(n24419) );
  NOR2_X2 U17040 ( .A1(n15342), .A2(n15341), .ZN(n8922) );
  NAND3_X2 U11313 ( .A1(n41197), .A2(n22304), .A3(n38674), .ZN(n41189) );
  CLKBUF_X4 U13804 ( .I(n51303), .Z(n56541) );
  INV_X4 U7068 ( .I(n19790), .ZN(n19789) );
  NAND2_X2 U7288 ( .A1(n16986), .A2(n19107), .ZN(n48771) );
  INV_X4 U4738 ( .I(n10526), .ZN(n17141) );
  INV_X2 U9106 ( .I(n23369), .ZN(n17092) );
  BUF_X4 U5822 ( .I(n45319), .Z(n22975) );
  NOR2_X2 U17175 ( .A1(n18745), .A2(n18744), .ZN(n18743) );
  NOR4_X2 U51436 ( .A1(n42976), .A2(n42807), .A3(n14605), .A4(n1298), .ZN(
        n42769) );
  INV_X2 U11884 ( .I(n17737), .ZN(n17738) );
  NOR2_X1 U1728 ( .A1(n42053), .A2(n15376), .ZN(n4551) );
  NAND2_X2 U912 ( .A1(n12579), .A2(n1473), .ZN(n50374) );
  NAND2_X2 U2971 ( .A1(n18048), .A2(n24028), .ZN(n58984) );
  INV_X2 U11885 ( .I(n28938), .ZN(n28937) );
  OAI22_X2 U44706 ( .A1(n19122), .A2(n27620), .B1(n27619), .B2(n430), .ZN(
        n27625) );
  NAND2_X2 U43127 ( .A1(n22936), .A2(n37319), .ZN(n35080) );
  NOR2_X2 U16676 ( .A1(n18822), .A2(n42057), .ZN(n4806) );
  NOR3_X1 U2877 ( .A1(n25031), .A2(n25029), .A3(n25030), .ZN(n18337) );
  INV_X2 U26722 ( .I(n54276), .ZN(n54221) );
  NOR2_X2 U16829 ( .A1(n42890), .A2(n23434), .ZN(n42891) );
  INV_X2 U71 ( .I(n55895), .ZN(n55871) );
  AOI21_X2 U4686 ( .A1(n11465), .A2(n59481), .B(n29747), .ZN(n28720) );
  NAND2_X2 U31870 ( .A1(n11619), .A2(n11618), .ZN(n35225) );
  NAND2_X2 U31871 ( .A1(n58048), .A2(n35713), .ZN(n11619) );
  BUF_X4 U15050 ( .I(n8122), .Z(n22817) );
  INV_X2 U1601 ( .I(n43325), .ZN(n42973) );
  INV_X4 U21877 ( .I(n24871), .ZN(n32972) );
  OAI21_X2 U17674 ( .A1(n14485), .A2(n13890), .B(n37245), .ZN(n13889) );
  INV_X4 U32682 ( .I(n51264), .ZN(n56564) );
  INV_X2 U17293 ( .I(n42522), .ZN(n14279) );
  INV_X2 U56668 ( .I(n56805), .ZN(n56813) );
  NAND2_X2 U27995 ( .A1(n14743), .A2(n63406), .ZN(n35501) );
  NAND3_X1 U14802 ( .A1(n58777), .A2(n41995), .A3(n63036), .ZN(n57553) );
  INV_X4 U11566 ( .I(n24228), .ZN(n36944) );
  AOI22_X2 U48549 ( .A1(n35581), .A2(n35580), .B1(n36027), .B2(n35579), .ZN(
        n35585) );
  INV_X1 U583 ( .I(n22332), .ZN(n52406) );
  INV_X4 U8828 ( .I(n9593), .ZN(n17096) );
  INV_X2 U9372 ( .I(n33966), .ZN(n23178) );
  NAND2_X2 U21603 ( .A1(n60116), .A2(n13198), .ZN(n59569) );
  INV_X2 U8757 ( .I(n3705), .ZN(n1273) );
  CLKBUF_X4 U5267 ( .I(n62530), .Z(n43626) );
  NOR2_X1 U12067 ( .A1(n1895), .A2(n1364), .ZN(n28366) );
  OAI21_X2 U16617 ( .A1(n57297), .A2(n60772), .B(n3707), .ZN(n11114) );
  OR2_X2 U13378 ( .A1(n37095), .A2(n57686), .Z(n37314) );
  NOR2_X1 U16305 ( .A1(n4562), .A2(n12036), .ZN(n58879) );
  INV_X2 U8740 ( .I(n42224), .ZN(n22289) );
  BUF_X2 U6082 ( .I(n36080), .Z(n58580) );
  INV_X2 U3599 ( .I(n15927), .ZN(n2617) );
  INV_X1 U9990 ( .I(n38729), .ZN(n37989) );
  AOI22_X2 U5673 ( .A1(n13472), .A2(n13527), .B1(n13526), .B2(n23301), .ZN(
        n24202) );
  NAND3_X2 U53199 ( .A1(n48135), .A2(n24545), .A3(n60390), .ZN(n47206) );
  OAI21_X2 U42555 ( .A1(n48583), .A2(n23018), .B(n61577), .ZN(n60697) );
  NOR2_X2 U14155 ( .A1(n27615), .A2(n27619), .ZN(n26603) );
  NAND2_X2 U7321 ( .A1(n13292), .A2(n53198), .ZN(n53607) );
  AOI21_X2 U1480 ( .A1(n43836), .A2(n43059), .B(n22677), .ZN(n43061) );
  NOR2_X2 U2822 ( .A1(n60441), .A2(n60440), .ZN(n13535) );
  NAND2_X2 U2404 ( .A1(n9593), .A2(n10717), .ZN(n12141) );
  INV_X4 U31158 ( .I(n24682), .ZN(n2403) );
  NAND3_X1 U14773 ( .A1(n56241), .A2(n56240), .A3(n23526), .ZN(n56242) );
  NOR2_X2 U890 ( .A1(n48717), .A2(n1384), .ZN(n49885) );
  INV_X2 U56518 ( .I(n56660), .ZN(n56367) );
  INV_X2 U26086 ( .I(n62530), .ZN(n43634) );
  BUF_X4 U28607 ( .I(n30810), .Z(n8521) );
  INV_X2 U3293 ( .I(n26912), .ZN(n29695) );
  CLKBUF_X4 U37804 ( .I(Key[153]), .Z(n56322) );
  BUF_X4 U9707 ( .I(n58852), .Z(n30374) );
  NAND3_X2 U11762 ( .A1(n6769), .A2(n29927), .A3(n10573), .ZN(n30534) );
  BUF_X2 U19872 ( .I(n27160), .Z(n23940) );
  OAI21_X2 U4234 ( .A1(n12468), .A2(n17860), .B(n12282), .ZN(n5889) );
  AOI22_X2 U29937 ( .A1(n46722), .A2(n21183), .B1(n46720), .B2(n46721), .ZN(
        n9837) );
  NOR2_X2 U8926 ( .A1(n15626), .A2(n21176), .ZN(n31033) );
  INV_X2 U38459 ( .I(n18747), .ZN(n27431) );
  AOI21_X2 U10963 ( .A1(n57677), .A2(n44770), .B(n3364), .ZN(n3367) );
  AOI21_X1 U25629 ( .A1(n16261), .A2(n22693), .B(n37916), .ZN(n58690) );
  INV_X1 U5015 ( .I(n21073), .ZN(n43922) );
  NAND4_X1 U5503 ( .A1(n54935), .A2(n54932), .A3(n54933), .A4(n54934), .ZN(
        n275) );
  NAND3_X2 U10381 ( .A1(n41125), .A2(n1731), .A3(n2193), .ZN(n41380) );
  AOI21_X2 U49019 ( .A1(n38552), .A2(n37138), .B(n37137), .ZN(n37139) );
  OAI21_X2 U49017 ( .A1(n22733), .A2(n63838), .B(n16027), .ZN(n37138) );
  AOI22_X2 U25482 ( .A1(n13683), .A2(n50259), .B1(n13024), .B2(n13682), .ZN(
        n15299) );
  INV_X1 U11497 ( .I(n20007), .ZN(n36976) );
  NOR2_X2 U2216 ( .A1(n34840), .A2(n34839), .ZN(n37495) );
  NAND2_X2 U11264 ( .A1(n5847), .A2(n23399), .ZN(n19592) );
  NAND2_X2 U33939 ( .A1(n63878), .A2(n62490), .ZN(n45757) );
  BUF_X8 U39661 ( .I(n37945), .Z(n19252) );
  BUF_X2 U5632 ( .I(n49948), .Z(n61170) );
  INV_X2 U32406 ( .I(n21006), .ZN(n21084) );
  NOR2_X2 U33088 ( .A1(n29727), .A2(n13176), .ZN(n13175) );
  NAND4_X1 U53808 ( .A1(n55353), .A2(n55351), .A3(n55352), .A4(n55354), .ZN(
        n55361) );
  NOR3_X1 U30028 ( .A1(n12473), .A2(n49348), .A3(n12472), .ZN(n61273) );
  OAI22_X2 U32878 ( .A1(n33962), .A2(n63305), .B1(n13698), .B2(n12859), .ZN(
        n13697) );
  NAND2_X2 U1795 ( .A1(n20276), .A2(n61743), .ZN(n43531) );
  INV_X4 U23477 ( .I(n50088), .ZN(n49720) );
  INV_X2 U10870 ( .I(n47932), .ZN(n49039) );
  INV_X4 U3139 ( .I(n30196), .ZN(n30183) );
  NAND2_X2 U4500 ( .A1(n10869), .A2(n23047), .ZN(n57636) );
  NOR3_X1 U789 ( .A1(n61248), .A2(n10346), .A3(n49689), .ZN(n217) );
  NOR2_X2 U1961 ( .A1(n64793), .A2(n62175), .ZN(n40633) );
  NAND2_X2 U13922 ( .A1(n6351), .A2(n53537), .ZN(n6350) );
  NAND3_X2 U11178 ( .A1(n45900), .A2(n11599), .A3(n70), .ZN(n47400) );
  NAND2_X2 U23920 ( .A1(n6041), .A2(n24000), .ZN(n29561) );
  INV_X4 U11345 ( .I(n41852), .ZN(n1403) );
  INV_X2 U4963 ( .I(n61388), .ZN(n41353) );
  INV_X4 U6861 ( .I(n33539), .ZN(n14329) );
  AOI21_X2 U13928 ( .A1(n13412), .A2(n13411), .B(n30862), .ZN(n31191) );
  INV_X2 U37734 ( .I(n22487), .ZN(n25840) );
  NAND3_X2 U26364 ( .A1(n11423), .A2(n63344), .A3(n63123), .ZN(n32964) );
  NAND2_X2 U8458 ( .A1(n35876), .A2(n37184), .ZN(n24660) );
  NOR2_X2 U23516 ( .A1(n13550), .A2(n48362), .ZN(n13549) );
  INV_X2 U15195 ( .I(n26007), .ZN(n1622) );
  NAND2_X1 U19171 ( .A1(n57890), .A2(n57889), .ZN(n59083) );
  NOR2_X2 U24899 ( .A1(n11125), .A2(n40162), .ZN(n40158) );
  BUF_X4 U3609 ( .I(n55947), .Z(n56084) );
  NAND2_X2 U13499 ( .A1(n34053), .A2(n34052), .ZN(n34064) );
  NAND3_X1 U14341 ( .A1(n13077), .A2(n13076), .A3(n7185), .ZN(n7184) );
  NOR2_X2 U10263 ( .A1(n39992), .A2(n10074), .ZN(n40004) );
  NAND2_X2 U21834 ( .A1(n19144), .A2(n17885), .ZN(n3281) );
  AOI22_X2 U10025 ( .A1(n16670), .A2(n43121), .B1(n26227), .B2(n3328), .ZN(
        n4865) );
  INV_X2 U48466 ( .I(n58743), .ZN(n35345) );
  INV_X4 U29334 ( .I(n9372), .ZN(n21489) );
  NOR2_X1 U52958 ( .A1(n61125), .A2(n61124), .ZN(n39702) );
  NAND3_X2 U2857 ( .A1(n17857), .A2(n17855), .A3(n17852), .ZN(n25332) );
  INV_X4 U9686 ( .I(n16279), .ZN(n1315) );
  INV_X4 U2609 ( .I(n34613), .ZN(n34042) );
  OAI22_X2 U18469 ( .A1(n34601), .A2(n22086), .B1(n34604), .B2(n19621), .ZN(
        n31515) );
  NAND3_X2 U26685 ( .A1(n34522), .A2(n7173), .A3(n58683), .ZN(n34053) );
  AOI21_X2 U20916 ( .A1(n50357), .A2(n50358), .B(n61436), .ZN(n50370) );
  OAI21_X2 U36294 ( .A1(n56418), .A2(n62846), .B(n56422), .ZN(n20001) );
  INV_X2 U7502 ( .I(n46096), .ZN(n48603) );
  INV_X2 U7490 ( .I(n29834), .ZN(n10820) );
  INV_X4 U43311 ( .I(n10232), .ZN(n34316) );
  NAND2_X2 U3565 ( .A1(n13081), .A2(n34771), .ZN(n60667) );
  NOR2_X2 U13318 ( .A1(n7284), .A2(n20007), .ZN(n37248) );
  NAND2_X1 U25568 ( .A1(n35117), .A2(n36403), .ZN(n35118) );
  INV_X2 U15704 ( .I(n50331), .ZN(n13684) );
  NAND2_X2 U1355 ( .A1(n15749), .A2(n10626), .ZN(n14519) );
  INV_X1 U21167 ( .I(n2814), .ZN(n7519) );
  BUF_X2 U6084 ( .I(n36740), .Z(n58769) );
  INV_X4 U38462 ( .I(n27621), .ZN(n26671) );
  NOR2_X2 U8687 ( .A1(n60583), .A2(n43845), .ZN(n43848) );
  BUF_X4 U2446 ( .I(n36246), .Z(n3856) );
  NAND3_X2 U7102 ( .A1(n36584), .A2(n798), .A3(n1790), .ZN(n11271) );
  NAND2_X2 U886 ( .A1(n6977), .A2(n50359), .ZN(n50369) );
  BUF_X4 U6706 ( .I(n50359), .Z(n59633) );
  BUF_X2 U4132 ( .I(n57122), .Z(n22516) );
  BUF_X4 U26654 ( .I(n18524), .Z(n6979) );
  AOI21_X2 U5602 ( .A1(n61541), .A2(n61540), .B(n50086), .ZN(n14041) );
  NAND2_X2 U15130 ( .A1(n8276), .A2(n4311), .ZN(n8275) );
  NAND2_X2 U52307 ( .A1(n23588), .A2(n20832), .ZN(n45619) );
  NAND2_X2 U55211 ( .A1(n58815), .A2(n60934), .ZN(n52849) );
  INV_X4 U3134 ( .I(n1192), .ZN(n21478) );
  BUF_X2 U13017 ( .I(n41432), .Z(n23406) );
  NAND2_X2 U7863 ( .A1(n18566), .A2(n60874), .ZN(n36056) );
  NAND3_X1 U8538 ( .A1(n47336), .A2(n15826), .A3(n47335), .ZN(n47337) );
  NOR3_X2 U2280 ( .A1(n35506), .A2(n4304), .A3(n34927), .ZN(n35954) );
  NAND3_X1 U55894 ( .A1(n54712), .A2(n19492), .A3(n54711), .ZN(n54714) );
  AND2_X2 U43779 ( .A1(n54667), .A2(n54666), .Z(n26015) );
  INV_X2 U1851 ( .I(n13673), .ZN(n42264) );
  OAI21_X1 U7530 ( .A1(n39503), .A2(n1732), .B(n2560), .ZN(n60069) );
  NAND3_X1 U23771 ( .A1(n35386), .A2(n35385), .A3(n36900), .ZN(n35395) );
  OAI22_X2 U53655 ( .A1(n18566), .A2(n19206), .B1(n35378), .B2(n36384), .ZN(
        n36899) );
  INV_X2 U6597 ( .I(n47858), .ZN(n47852) );
  NOR2_X2 U18447 ( .A1(n33578), .A2(n22850), .ZN(n33581) );
  OAI22_X2 U35022 ( .A1(n33577), .A2(n24286), .B1(n1341), .B2(n6979), .ZN(
        n22850) );
  AOI22_X2 U13384 ( .A1(n36345), .A2(n35072), .B1(n36749), .B2(n36343), .ZN(
        n35073) );
  INV_X1 U56946 ( .I(n63042), .ZN(n61523) );
  INV_X1 U55129 ( .I(n57072), .ZN(n57057) );
  INV_X4 U10174 ( .I(n39994), .ZN(n12158) );
  NAND2_X2 U10535 ( .A1(n13393), .A2(n42049), .ZN(n43429) );
  INV_X2 U1369 ( .I(n61960), .ZN(n1329) );
  OAI21_X2 U5399 ( .A1(n27216), .A2(n29304), .B(n27215), .ZN(n27223) );
  INV_X4 U4634 ( .I(n6727), .ZN(n25532) );
  OAI22_X1 U22454 ( .A1(n3781), .A2(n1254), .B1(n57090), .B2(n14778), .ZN(
        n57092) );
  OR2_X1 U29891 ( .A1(n57032), .A2(n60225), .Z(n2742) );
  NAND2_X2 U11996 ( .A1(n10324), .A2(n29304), .ZN(n24231) );
  INV_X2 U31034 ( .I(n30145), .ZN(n31039) );
  NAND2_X2 U8041 ( .A1(n22444), .A2(n57621), .ZN(n29904) );
  INV_X2 U41092 ( .I(n21303), .ZN(n48095) );
  NOR2_X2 U17876 ( .A1(n36500), .A2(n19641), .ZN(n36501) );
  AOI22_X2 U8677 ( .A1(n42125), .A2(n42128), .B1(n41784), .B2(n11881), .ZN(
        n11880) );
  OAI21_X1 U53669 ( .A1(n48831), .A2(n48830), .B(n48829), .ZN(n48836) );
  INV_X2 U51296 ( .I(n42185), .ZN(n42186) );
  OAI21_X2 U48703 ( .A1(n36327), .A2(n37404), .B(n17660), .ZN(n36159) );
  INV_X4 U42747 ( .I(n15753), .ZN(n49389) );
  AND2_X2 U26889 ( .A1(n20571), .A2(n36020), .Z(n34823) );
  BUF_X4 U13727 ( .I(n31701), .Z(n33654) );
  INV_X4 U2470 ( .I(n36443), .ZN(n1792) );
  BUF_X8 U12685 ( .I(n48135), .Z(n7186) );
  NAND2_X2 U6105 ( .A1(n34351), .A2(n32423), .ZN(n21456) );
  NAND2_X2 U23280 ( .A1(n47902), .A2(n47900), .ZN(n45595) );
  OAI21_X2 U688 ( .A1(n9696), .A2(n9695), .B(n1633), .ZN(n25064) );
  NOR2_X1 U33140 ( .A1(n59518), .A2(n59517), .ZN(n59516) );
  INV_X4 U32604 ( .I(n20514), .ZN(n47886) );
  AOI21_X2 U4213 ( .A1(n11510), .A2(n1930), .B(n28214), .ZN(n11509) );
  NOR2_X2 U38693 ( .A1(n60032), .A2(n57295), .ZN(n55185) );
  NOR2_X2 U45390 ( .A1(n1866), .A2(n17590), .ZN(n31173) );
  NAND2_X2 U34931 ( .A1(n1192), .A2(n29726), .ZN(n25470) );
  INV_X4 U1294 ( .I(n58018), .ZN(n24354) );
  AOI22_X2 U39491 ( .A1(n47596), .A2(n47595), .B1(n47594), .B2(n63338), .ZN(
        n47598) );
  NAND2_X2 U6756 ( .A1(n1080), .A2(n63953), .ZN(n44559) );
  NAND2_X2 U10055 ( .A1(n43220), .A2(n24981), .ZN(n43093) );
  INV_X4 U20275 ( .I(n57978), .ZN(n39959) );
  NAND2_X2 U38873 ( .A1(n18003), .A2(n58636), .ZN(n47633) );
  OAI21_X1 U6721 ( .A1(n45178), .A2(n57633), .B(n57632), .ZN(n45190) );
  INV_X2 U436 ( .I(n55270), .ZN(n55266) );
  NAND3_X2 U25459 ( .A1(n48396), .A2(n49465), .A3(n1205), .ZN(n48397) );
  INV_X1 U23358 ( .I(n41506), .ZN(n58371) );
  INV_X2 U3443 ( .I(n15790), .ZN(n11873) );
  NAND2_X2 U27079 ( .A1(n45532), .A2(n22905), .ZN(n45779) );
  NAND2_X2 U11821 ( .A1(n29205), .A2(n23349), .ZN(n30246) );
  NAND2_X2 U3499 ( .A1(n7534), .A2(n18300), .ZN(n34507) );
  NAND2_X2 U3323 ( .A1(n29297), .A2(n1575), .ZN(n26964) );
  BUF_X4 U57106 ( .I(n31085), .Z(n61629) );
  NAND3_X2 U24552 ( .A1(n47300), .A2(n18843), .A3(n15383), .ZN(n3662) );
  INV_X2 U11680 ( .I(n22597), .ZN(n15303) );
  NOR3_X1 U44736 ( .A1(n17652), .A2(n17650), .A3(n17651), .ZN(n17649) );
  INV_X12 U4506 ( .I(n29516), .ZN(n1838) );
  AND2_X2 U10333 ( .A1(n8217), .A2(n59134), .Z(n8365) );
  BUF_X4 U47442 ( .I(n32635), .Z(n35629) );
  NAND3_X2 U40025 ( .A1(n56478), .A2(n65216), .A3(n56510), .ZN(n19728) );
  NAND2_X2 U12198 ( .A1(n54958), .A2(n54957), .ZN(n20802) );
  NAND2_X2 U346 ( .A1(n14468), .A2(n4783), .ZN(n54958) );
  INV_X4 U3354 ( .I(n64445), .ZN(n27619) );
  INV_X4 U56937 ( .I(n32528), .ZN(n33701) );
  INV_X2 U9214 ( .I(n19489), .ZN(n1636) );
  NOR2_X2 U32003 ( .A1(n29568), .A2(n17590), .ZN(n29902) );
  NOR2_X2 U9900 ( .A1(n9041), .A2(n25125), .ZN(n34110) );
  BUF_X4 U13336 ( .I(n30024), .Z(n1192) );
  INV_X2 U1492 ( .I(n41588), .ZN(n1492) );
  INV_X2 U41789 ( .I(n60423), .ZN(n45991) );
  OAI22_X2 U2788 ( .A1(n13961), .A2(n17668), .B1(n13963), .B2(n13962), .ZN(
        n16434) );
  INV_X4 U1759 ( .I(n42355), .ZN(n1501) );
  NAND2_X2 U4236 ( .A1(n45988), .A2(n47622), .ZN(n45207) );
  NAND2_X1 U1440 ( .A1(n38060), .A2(n38059), .ZN(n13314) );
  NAND4_X2 U35032 ( .A1(n31419), .A2(n33433), .A3(n31418), .A4(n33435), .ZN(
        n31420) );
  NOR2_X2 U36661 ( .A1(n18752), .A2(n26633), .ZN(n26639) );
  NAND3_X2 U9615 ( .A1(n6538), .A2(n6535), .A3(n30686), .ZN(n32339) );
  NAND2_X2 U978 ( .A1(n62139), .A2(n48803), .ZN(n7288) );
  NOR2_X2 U48667 ( .A1(n36054), .A2(n36389), .ZN(n36055) );
  NAND2_X2 U40247 ( .A1(n20141), .A2(n9205), .ZN(n33611) );
  INV_X2 U40248 ( .I(n33004), .ZN(n20141) );
  INV_X1 U3827 ( .I(n10300), .ZN(n2777) );
  OAI21_X2 U4733 ( .A1(n17141), .A2(n34224), .B(n35806), .ZN(n17474) );
  INV_X2 U39217 ( .I(n579), .ZN(n60112) );
  INV_X2 U2489 ( .I(n19322), .ZN(n35427) );
  NOR2_X2 U20202 ( .A1(n8817), .A2(n7338), .ZN(n59925) );
  INV_X2 U53746 ( .I(n29254), .ZN(n61175) );
  NOR2_X1 U47883 ( .A1(n33501), .A2(n60579), .ZN(n33504) );
  NOR2_X2 U3132 ( .A1(n1316), .A2(n30588), .ZN(n29487) );
  NAND2_X2 U8357 ( .A1(n26883), .A2(n264), .ZN(n27696) );
  NOR2_X2 U5050 ( .A1(n45633), .A2(n3641), .ZN(n46022) );
  NAND2_X2 U1423 ( .A1(n46016), .A2(n46013), .ZN(n45633) );
  INV_X2 U492 ( .I(n56269), .ZN(n1370) );
  NAND2_X2 U12574 ( .A1(n48186), .A2(n46483), .ZN(n47152) );
  INV_X2 U28849 ( .I(n13538), .ZN(n8794) );
  BUF_X4 U31001 ( .I(n16764), .Z(n10525) );
  NAND2_X2 U40740 ( .A1(n49420), .A2(n50074), .ZN(n49421) );
  INV_X2 U5076 ( .I(n6001), .ZN(n21938) );
  OAI21_X2 U47677 ( .A1(n35217), .A2(n33083), .B(n35210), .ZN(n33086) );
  AOI21_X2 U27304 ( .A1(n54012), .A2(n54013), .B(n59872), .ZN(n54014) );
  NAND2_X2 U3381 ( .A1(n23352), .A2(n14439), .ZN(n11850) );
  AOI21_X2 U8958 ( .A1(n18236), .A2(n29206), .B(n22496), .ZN(n18235) );
  CLKBUF_X4 U8405 ( .I(n15739), .Z(n1238) );
  INV_X2 U9280 ( .I(n46794), .ZN(n48146) );
  BUF_X4 U1139 ( .I(n3658), .Z(n60772) );
  NAND2_X2 U683 ( .A1(n49646), .A2(n49644), .ZN(n11216) );
  OR2_X2 U2631 ( .A1(n38529), .A2(n40961), .Z(n39136) );
  INV_X4 U8952 ( .I(n16764), .ZN(n13810) );
  AOI21_X2 U32413 ( .A1(n42024), .A2(n42022), .B(n12378), .ZN(n42023) );
  INV_X4 U28341 ( .I(n892), .ZN(n35229) );
  OAI21_X1 U49657 ( .A1(n41806), .A2(n41306), .B(n40361), .ZN(n38198) );
  BUF_X4 U6253 ( .I(n49929), .Z(n502) );
  INV_X2 U2646 ( .I(n11373), .ZN(n37072) );
  INV_X4 U22001 ( .I(n15615), .ZN(n58207) );
  NOR2_X1 U19440 ( .A1(n27514), .A2(n27513), .ZN(n8670) );
  NAND3_X2 U2523 ( .A1(n35220), .A2(n23859), .A3(n7710), .ZN(n35707) );
  NAND2_X2 U7328 ( .A1(n52844), .A2(n53198), .ZN(n53386) );
  INV_X4 U33754 ( .I(n25162), .ZN(n49459) );
  NAND3_X1 U38922 ( .A1(n1537), .A2(n32298), .A3(n18077), .ZN(n32299) );
  NAND2_X2 U3001 ( .A1(n21532), .A2(n30216), .ZN(n30225) );
  CLKBUF_X4 U7757 ( .I(n23696), .Z(n2748) );
  NAND3_X2 U18645 ( .A1(n30830), .A2(n30831), .A3(n21910), .ZN(n21909) );
  NAND2_X2 U7029 ( .A1(n29220), .A2(n9426), .ZN(n30718) );
  NAND2_X1 U15216 ( .A1(n10855), .A2(n5600), .ZN(n5599) );
  INV_X2 U11036 ( .I(n44252), .ZN(n1390) );
  INV_X4 U7532 ( .I(n23904), .ZN(n40304) );
  NAND2_X1 U6911 ( .A1(n13197), .A2(n7431), .ZN(n52581) );
  INV_X4 U38424 ( .I(n15875), .ZN(n17860) );
  INV_X2 U5546 ( .I(n19146), .ZN(n1617) );
  NAND2_X2 U545 ( .A1(n5227), .A2(n1371), .ZN(n5226) );
  NOR2_X1 U103 ( .A1(n54213), .A2(n23731), .ZN(n54233) );
  NAND2_X2 U37825 ( .A1(n22461), .A2(n64967), .ZN(n35511) );
  BUF_X4 U9983 ( .I(n39365), .Z(n23790) );
  INV_X1 U18768 ( .I(n24012), .ZN(n4630) );
  NAND2_X2 U6064 ( .A1(n10165), .A2(n15794), .ZN(n10705) );
  AOI22_X2 U22756 ( .A1(n58303), .A2(n54493), .B1(n54068), .B2(n54307), .ZN(
        n52993) );
  INV_X2 U1405 ( .I(n45357), .ZN(n19864) );
  OAI21_X2 U38614 ( .A1(n60026), .A2(n40179), .B(n40177), .ZN(n40184) );
  INV_X2 U1706 ( .I(n9672), .ZN(n40173) );
  BUF_X4 U12342 ( .I(n11270), .Z(n11269) );
  NAND2_X2 U8802 ( .A1(n36384), .A2(n6440), .ZN(n36532) );
  NAND2_X2 U14521 ( .A1(n54508), .A2(n62629), .ZN(n54551) );
  INV_X2 U9159 ( .I(n25214), .ZN(n54802) );
  INV_X4 U19320 ( .I(n30736), .ZN(n13280) );
  NOR2_X1 U8139 ( .A1(n59088), .A2(n59087), .ZN(n59141) );
  INV_X1 U27399 ( .I(n53904), .ZN(n21124) );
  NOR2_X2 U2512 ( .A1(n38338), .A2(n42432), .ZN(n42438) );
  BUF_X2 U8769 ( .I(n25479), .Z(n17154) );
  NAND3_X2 U53530 ( .A1(n48340), .A2(n49909), .A3(n48339), .ZN(n48342) );
  INV_X2 U30883 ( .I(n10455), .ZN(n13811) );
  NAND3_X2 U21234 ( .A1(n2875), .A2(n4063), .A3(n26586), .ZN(n2874) );
  NAND3_X2 U31988 ( .A1(n11792), .A2(n37582), .A3(n58842), .ZN(n11790) );
  NAND3_X2 U56794 ( .A1(n38357), .A2(n61429), .A3(n7139), .ZN(n38358) );
  BUF_X4 U24975 ( .I(n55680), .Z(n58626) );
  BUF_X4 U4094 ( .I(n56812), .Z(n23879) );
  AOI21_X2 U11079 ( .A1(n41989), .A2(n41988), .B(n24569), .ZN(n24568) );
  NOR2_X2 U6964 ( .A1(n27380), .A2(n27381), .ZN(n26527) );
  NAND2_X1 U2851 ( .A1(n20695), .A2(n23154), .ZN(n22715) );
  INV_X2 U808 ( .I(n45547), .ZN(n11058) );
  INV_X2 U5056 ( .I(n21667), .ZN(n43289) );
  INV_X2 U12891 ( .I(n14905), .ZN(n41539) );
  INV_X1 U20973 ( .I(n6686), .ZN(n21346) );
  NAND4_X2 U15835 ( .A1(n54287), .A2(n54288), .A3(n21037), .A4(n26250), .ZN(
        n57657) );
  INV_X4 U1994 ( .I(n8523), .ZN(n20190) );
  NOR2_X2 U9627 ( .A1(n25671), .A2(n37034), .ZN(n14136) );
  NAND2_X2 U9515 ( .A1(n4263), .A2(n36193), .ZN(n36114) );
  OAI21_X2 U45546 ( .A1(n10821), .A2(n29937), .B(n29936), .ZN(n29938) );
  INV_X2 U12311 ( .I(n53213), .ZN(n52828) );
  INV_X2 U433 ( .I(n54802), .ZN(n54806) );
  NOR2_X2 U36333 ( .A1(n16489), .A2(n17286), .ZN(n17287) );
  INV_X2 U54590 ( .I(n56894), .ZN(n56881) );
  INV_X2 U9207 ( .I(n48957), .ZN(n49176) );
  AOI21_X2 U18450 ( .A1(n22253), .A2(n32941), .B(n57571), .ZN(n24514) );
  NAND2_X2 U8796 ( .A1(n13666), .A2(n37945), .ZN(n37022) );
  INV_X2 U9749 ( .I(n29155), .ZN(n27974) );
  INV_X2 U39350 ( .I(n25078), .ZN(n33573) );
  NOR2_X2 U2996 ( .A1(n30679), .A2(n13810), .ZN(n26781) );
  INV_X2 U12434 ( .I(n33573), .ZN(n35670) );
  NAND3_X2 U22069 ( .A1(n30667), .A2(n30760), .A3(n1278), .ZN(n30749) );
  INV_X2 U15108 ( .I(n52094), .ZN(n7743) );
  OR2_X2 U1923 ( .A1(n15252), .A2(n43319), .Z(n41483) );
  NOR2_X2 U16799 ( .A1(n5474), .A2(n57711), .ZN(n5473) );
  NAND4_X2 U52542 ( .A1(n7113), .A2(n23156), .A3(n19705), .A4(n47970), .ZN(
        n45546) );
  BUF_X4 U6073 ( .I(n36052), .Z(n10165) );
  NAND2_X2 U32059 ( .A1(n36775), .A2(n15794), .ZN(n36764) );
  NAND2_X2 U42050 ( .A1(n49910), .A2(n49904), .ZN(n49899) );
  INV_X2 U10494 ( .I(n20315), .ZN(n21559) );
  AOI21_X2 U10701 ( .A1(n56612), .A2(n56611), .B(n56610), .ZN(n56613) );
  INV_X4 U32180 ( .I(n13955), .ZN(n22505) );
  NAND2_X2 U4173 ( .A1(n55016), .A2(n7800), .ZN(n54457) );
  INV_X4 U31383 ( .I(n10909), .ZN(n21409) );
  OAI21_X1 U34257 ( .A1(n59640), .A2(n59639), .B(n48781), .ZN(n48787) );
  INV_X4 U9421 ( .I(n17866), .ZN(n5386) );
  NAND3_X2 U2698 ( .A1(n21146), .A2(n21147), .A3(n20131), .ZN(n20130) );
  INV_X4 U10183 ( .I(n40944), .ZN(n40203) );
  INV_X2 U8177 ( .I(n40947), .ZN(n40949) );
  INV_X2 U25771 ( .I(n48728), .ZN(n49918) );
  INV_X1 U21697 ( .I(n15616), .ZN(n40145) );
  AOI21_X2 U53687 ( .A1(n48879), .A2(n49215), .B(n48878), .ZN(n48880) );
  OAI21_X2 U53686 ( .A1(n48877), .A2(n48876), .B(n49322), .ZN(n48878) );
  INV_X4 U582 ( .I(n7800), .ZN(n7697) );
  NAND3_X2 U321 ( .A1(n61213), .A2(n55982), .A3(n24473), .ZN(n56428) );
  NAND2_X2 U13353 ( .A1(n35863), .A2(n9013), .ZN(n35421) );
  NAND2_X2 U3272 ( .A1(n4324), .A2(n26654), .ZN(n27180) );
  INV_X1 U35230 ( .I(n25333), .ZN(n32868) );
  NAND2_X2 U9729 ( .A1(n62942), .A2(n35497), .ZN(n60356) );
  INV_X2 U3363 ( .I(n12221), .ZN(n28342) );
  OAI22_X2 U16255 ( .A1(n12506), .A2(n63375), .B1(n35670), .B2(n18879), .ZN(
        n33083) );
  BUF_X2 U55713 ( .I(n13837), .Z(n61321) );
  NAND2_X2 U3400 ( .A1(n28128), .A2(n28127), .ZN(n29283) );
  OAI21_X2 U55289 ( .A1(n53451), .A2(n53572), .B(n53002), .ZN(n53003) );
  INV_X2 U2247 ( .I(n36921), .ZN(n1414) );
  NAND2_X2 U12621 ( .A1(n45639), .A2(n47292), .ZN(n45630) );
  NOR2_X2 U4419 ( .A1(n49096), .A2(n58645), .ZN(n49098) );
  NAND2_X2 U17670 ( .A1(n12451), .A2(n12450), .ZN(n14892) );
  CLKBUF_X4 U18575 ( .I(n33391), .Z(n22413) );
  INV_X2 U2385 ( .I(n35363), .ZN(n36402) );
  INV_X2 U2379 ( .I(n35898), .ZN(n35885) );
  BUF_X4 U13654 ( .I(n33763), .Z(n23761) );
  NAND2_X1 U189 ( .A1(n9068), .A2(n59538), .ZN(n55035) );
  INV_X2 U16920 ( .I(n42892), .ZN(n41767) );
  NOR2_X2 U38003 ( .A1(n61811), .A2(n16661), .ZN(n16660) );
  INV_X4 U43133 ( .I(n37351), .ZN(n37359) );
  NAND3_X2 U4125 ( .A1(n13925), .A2(n50042), .A3(n3335), .ZN(n50048) );
  NAND2_X2 U26902 ( .A1(n56045), .A2(n56107), .ZN(n56050) );
  NAND3_X2 U11243 ( .A1(n17577), .A2(n40638), .A3(n17576), .ZN(n17575) );
  BUF_X2 U37658 ( .I(n33810), .Z(n35755) );
  INV_X2 U3278 ( .I(n23039), .ZN(n26635) );
  NAND2_X2 U8316 ( .A1(n14361), .A2(n22797), .ZN(n24942) );
  NAND2_X2 U20327 ( .A1(n11719), .A2(n2267), .ZN(n30253) );
  NAND2_X2 U44201 ( .A1(n27109), .A2(n26626), .ZN(n26623) );
  NOR2_X2 U4966 ( .A1(n12411), .A2(n13603), .ZN(n2753) );
  NAND2_X2 U4938 ( .A1(n23692), .A2(n42721), .ZN(n12411) );
  BUF_X2 U6930 ( .I(n44994), .Z(n59218) );
  BUF_X4 U10186 ( .I(n4995), .Z(n8523) );
  OAI21_X1 U56369 ( .A1(n56003), .A2(n63699), .B(n56002), .ZN(n56004) );
  INV_X2 U17064 ( .I(n23406), .ZN(n19387) );
  OAI21_X1 U51833 ( .A1(n44070), .A2(n47471), .B(n44069), .ZN(n44076) );
  NOR2_X2 U7196 ( .A1(n43092), .A2(n11476), .ZN(n43227) );
  NAND3_X2 U52561 ( .A1(n47574), .A2(n47900), .A3(n47577), .ZN(n45586) );
  NAND2_X2 U9657 ( .A1(n22595), .A2(n34816), .ZN(n16354) );
  INV_X2 U5914 ( .I(n16493), .ZN(n12825) );
  NOR2_X2 U867 ( .A1(n50373), .A2(n5282), .ZN(n50098) );
  INV_X4 U39741 ( .I(n27665), .ZN(n28492) );
  BUF_X4 U20942 ( .I(Key[183]), .Z(n58084) );
  NOR2_X2 U18513 ( .A1(n33219), .A2(n33538), .ZN(n32604) );
  INV_X4 U34628 ( .I(n24293), .ZN(n34708) );
  INV_X2 U37516 ( .I(n52117), .ZN(n55437) );
  NAND2_X2 U17886 ( .A1(n36758), .A2(n37289), .ZN(n36291) );
  INV_X2 U486 ( .I(n55445), .ZN(n55006) );
  NAND2_X2 U7040 ( .A1(n20989), .A2(n34752), .ZN(n34740) );
  NAND3_X1 U11412 ( .A1(n36907), .A2(n36906), .A3(n36905), .ZN(n36919) );
  INV_X1 U45660 ( .I(n30184), .ZN(n30185) );
  NOR2_X2 U45761 ( .A1(n1860), .A2(n23478), .ZN(n30444) );
  INV_X4 U7517 ( .I(n24299), .ZN(n1860) );
  NAND3_X1 U23469 ( .A1(n10445), .A2(n24193), .A3(n54385), .ZN(n4622) );
  INV_X2 U8362 ( .I(n19000), .ZN(n43189) );
  BUF_X4 U12227 ( .I(n54813), .Z(n23849) );
  NAND2_X2 U23072 ( .A1(n59614), .A2(n10493), .ZN(n12941) );
  INV_X2 U629 ( .I(n60867), .ZN(n54102) );
  NAND4_X1 U34970 ( .A1(n18633), .A2(n8732), .A3(n47189), .A4(n48533), .ZN(
        n18632) );
  OR2_X1 U20495 ( .A1(n5582), .A2(n33928), .Z(n16782) );
  INV_X1 U4857 ( .I(n22601), .ZN(n32845) );
  NOR3_X2 U5398 ( .A1(n64684), .A2(n34578), .A3(n34579), .ZN(n34581) );
  NOR2_X2 U762 ( .A1(n49377), .A2(n58983), .ZN(n16406) );
  AND2_X2 U13429 ( .A1(n11348), .A2(n11350), .Z(n11347) );
  INV_X2 U18032 ( .I(n35430), .ZN(n5959) );
  INV_X2 U9689 ( .I(n58273), .ZN(n20172) );
  BUF_X2 U9777 ( .I(n22190), .Z(n28240) );
  NAND3_X1 U19002 ( .A1(n31058), .A2(n31056), .A3(n31057), .ZN(n14725) );
  NOR2_X2 U10277 ( .A1(n40958), .A2(n64040), .ZN(n39124) );
  NAND3_X2 U11758 ( .A1(n61755), .A2(n27792), .A3(n3794), .ZN(n7813) );
  AOI22_X1 U1367 ( .A1(n15567), .A2(n15568), .B1(n45670), .B2(n15566), .ZN(
        n59699) );
  INV_X4 U21931 ( .I(n16617), .ZN(n26145) );
  OAI21_X2 U16620 ( .A1(n41545), .A2(n42031), .B(n41539), .ZN(n9713) );
  NAND2_X2 U984 ( .A1(n7868), .A2(n19144), .ZN(n12536) );
  BUF_X2 U17464 ( .I(n41419), .Z(n20652) );
  INV_X1 U24872 ( .I(n5206), .ZN(n24947) );
  INV_X2 U32028 ( .I(n15758), .ZN(n11849) );
  INV_X2 U354 ( .I(n8597), .ZN(n56988) );
  NAND2_X1 U4237 ( .A1(n3734), .A2(n7588), .ZN(n11036) );
  NOR2_X1 U28453 ( .A1(n8367), .A2(n12553), .ZN(n12552) );
  BUF_X4 U2403 ( .I(n11413), .Z(n11272) );
  NOR2_X1 U6187 ( .A1(n60849), .A2(n63140), .ZN(n29756) );
  NOR2_X2 U53546 ( .A1(n15021), .A2(n10958), .ZN(n49921) );
  BUF_X4 U9170 ( .I(n10635), .Z(n11071) );
  NAND2_X2 U11995 ( .A1(n24980), .A2(n55695), .ZN(n19456) );
  NOR2_X2 U8954 ( .A1(n1432), .A2(n30736), .ZN(n25512) );
  NOR3_X2 U6713 ( .A1(n3444), .A2(n3443), .A3(n12657), .ZN(n13216) );
  NAND2_X2 U4290 ( .A1(n14019), .A2(n28607), .ZN(n27854) );
  AOI22_X1 U5420 ( .A1(n10835), .A2(n10834), .B1(n52312), .B2(n19120), .ZN(
        n57638) );
  INV_X4 U3351 ( .I(n15758), .ZN(n13672) );
  INV_X2 U52592 ( .I(n45651), .ZN(n45652) );
  OAI21_X2 U44510 ( .A1(n27140), .A2(n7438), .B(n27139), .ZN(n27144) );
  INV_X2 U9544 ( .I(n35822), .ZN(n34717) );
  AOI21_X2 U36125 ( .A1(n45451), .A2(n46737), .B(n46730), .ZN(n45454) );
  INV_X1 U2980 ( .I(n62999), .ZN(n29963) );
  BUF_X2 U32347 ( .I(n21751), .Z(n59676) );
  NOR3_X1 U7109 ( .A1(n36799), .A2(n19185), .A3(n36798), .ZN(n36816) );
  NAND2_X2 U7343 ( .A1(n53147), .A2(n20735), .ZN(n53162) );
  BUF_X2 U31524 ( .I(n476), .Z(n59293) );
  BUF_X4 U43870 ( .I(n50723), .Z(n53214) );
  NAND3_X2 U48137 ( .A1(n35822), .A2(n34232), .A3(n34324), .ZN(n34235) );
  CLKBUF_X8 U27637 ( .I(n15866), .Z(n1209) );
  BUF_X4 U45878 ( .I(Key[154]), .Z(n56335) );
  NAND2_X2 U7202 ( .A1(n60952), .A2(n775), .ZN(n41781) );
  BUF_X4 U6102 ( .I(n1225), .Z(n2330) );
  BUF_X4 U11898 ( .I(n23138), .Z(n1433) );
  INV_X2 U9817 ( .I(n24660), .ZN(n37334) );
  NOR3_X2 U23563 ( .A1(n46742), .A2(n46741), .A3(n46744), .ZN(n23106) );
  BUF_X2 U18882 ( .I(n32327), .Z(n23424) );
  INV_X4 U27589 ( .I(n54758), .ZN(n22385) );
  OAI21_X2 U48331 ( .A1(n7488), .A2(n35881), .B(n35901), .ZN(n34873) );
  NAND2_X1 U28308 ( .A1(n12522), .A2(n8223), .ZN(n35919) );
  INV_X2 U937 ( .I(n60726), .ZN(n1469) );
  OAI21_X2 U11256 ( .A1(n40635), .A2(n6890), .B(n40634), .ZN(n17577) );
  OAI21_X2 U44176 ( .A1(n26547), .A2(n26546), .B(n26627), .ZN(n26556) );
  BUF_X2 U14962 ( .I(n55445), .Z(n24454) );
  BUF_X2 U27683 ( .I(n22782), .Z(n15202) );
  OR2_X1 U26561 ( .A1(n9346), .A2(n23912), .Z(n9727) );
  INV_X4 U21168 ( .I(n22882), .ZN(n42502) );
  BUF_X2 U4127 ( .I(n8473), .Z(n8472) );
  NAND2_X2 U17850 ( .A1(n35421), .A2(n36750), .ZN(n10210) );
  NAND2_X2 U26495 ( .A1(n34507), .A2(n2322), .ZN(n34512) );
  NAND2_X2 U38330 ( .A1(n24641), .A2(n63593), .ZN(n36750) );
  NAND2_X2 U1669 ( .A1(n43327), .A2(n9663), .ZN(n41481) );
  INV_X1 U42609 ( .I(n42522), .ZN(n42209) );
  NAND3_X2 U33906 ( .A1(n28934), .A2(n28781), .A3(n18198), .ZN(n14391) );
  BUF_X2 U27031 ( .I(n46377), .Z(n10282) );
  NOR2_X1 U27012 ( .A1(n46102), .A2(n46101), .ZN(n48649) );
  NOR2_X2 U6844 ( .A1(n46101), .A2(n209), .ZN(n13506) );
  BUF_X2 U16308 ( .I(n16617), .Z(n3365) );
  NOR2_X1 U30681 ( .A1(n48649), .A2(n47489), .ZN(n13177) );
  NOR2_X2 U1901 ( .A1(n40025), .A2(n40229), .ZN(n40228) );
  OAI21_X2 U44873 ( .A1(n27993), .A2(n27992), .B(n27991), .ZN(n27994) );
  OAI21_X2 U12684 ( .A1(n57677), .A2(n44770), .B(n3365), .ZN(n3366) );
  NAND2_X2 U3372 ( .A1(n837), .A2(n22190), .ZN(n27381) );
  INV_X2 U37059 ( .I(n44064), .ZN(n45520) );
  BUF_X4 U10105 ( .I(n24631), .Z(n1226) );
  AOI22_X1 U29522 ( .A1(n45571), .A2(n45985), .B1(n9549), .B2(n22468), .ZN(
        n14412) );
  NAND3_X1 U1312 ( .A1(n9173), .A2(n25691), .A3(n1655), .ZN(n58140) );
  NOR2_X2 U30360 ( .A1(n14330), .A2(n12849), .ZN(n12848) );
  INV_X2 U26777 ( .I(n8237), .ZN(n17238) );
  INV_X4 U27838 ( .I(n8361), .ZN(n9792) );
  INV_X4 U25732 ( .I(n6168), .ZN(n6135) );
  INV_X2 U32932 ( .I(n53415), .ZN(n53625) );
  AOI21_X2 U16083 ( .A1(n47466), .A2(n8155), .B(n61738), .ZN(n8153) );
  NAND3_X2 U11203 ( .A1(n11298), .A2(n14962), .A3(n47512), .ZN(n11293) );
  OAI21_X2 U6761 ( .A1(n19568), .A2(n47045), .B(n47517), .ZN(n11298) );
  AOI21_X2 U38792 ( .A1(n29954), .A2(n21886), .B(n30786), .ZN(n29955) );
  BUF_X1 U13397 ( .I(n34524), .Z(n23065) );
  NAND2_X2 U41208 ( .A1(n27292), .A2(n62714), .ZN(n21511) );
  NAND2_X2 U358 ( .A1(n61560), .A2(n53859), .ZN(n53852) );
  NAND3_X2 U48139 ( .A1(n34319), .A2(n35304), .A3(n35811), .ZN(n34243) );
  NAND2_X2 U37333 ( .A1(n54350), .A2(n1611), .ZN(n24637) );
  INV_X2 U40535 ( .I(n21499), .ZN(n27292) );
  NOR2_X2 U1791 ( .A1(n11941), .A2(n23855), .ZN(n40299) );
  INV_X4 U829 ( .I(n49777), .ZN(n22869) );
  INV_X2 U17898 ( .I(n6329), .ZN(n36489) );
  OAI21_X2 U16653 ( .A1(n24715), .A2(n42633), .B(n61894), .ZN(n8934) );
  NAND2_X2 U27465 ( .A1(n7632), .A2(n62711), .ZN(n55200) );
  AOI21_X2 U36772 ( .A1(n25707), .A2(n30857), .B(n13412), .ZN(n30860) );
  INV_X1 U38258 ( .I(n17133), .ZN(n41112) );
  BUF_X4 U30916 ( .I(n23347), .Z(n10475) );
  AND2_X2 U32519 ( .A1(n30632), .A2(n20391), .Z(n30746) );
  NOR2_X2 U42121 ( .A1(n14848), .A2(n54727), .ZN(n54762) );
  NAND2_X2 U3155 ( .A1(n29586), .A2(n59268), .ZN(n29085) );
  INV_X2 U26648 ( .I(n2633), .ZN(n48186) );
  BUF_X4 U9837 ( .I(n12798), .Z(n24033) );
  INV_X8 U19349 ( .I(n29586), .ZN(n8097) );
  NAND3_X1 U45399 ( .A1(n65233), .A2(n59710), .A3(n10240), .ZN(n29587) );
  NAND2_X2 U1160 ( .A1(n1082), .A2(n209), .ZN(n48246) );
  NOR2_X2 U3302 ( .A1(n27930), .A2(n27298), .ZN(n29138) );
  NOR2_X1 U15724 ( .A1(n14694), .A2(n14693), .ZN(n14692) );
  NAND2_X2 U36495 ( .A1(n1779), .A2(n9721), .ZN(n34876) );
  NAND2_X2 U13532 ( .A1(n9028), .A2(n9030), .ZN(n19316) );
  NAND2_X2 U21776 ( .A1(n40631), .A2(n40639), .ZN(n17574) );
  NAND2_X2 U39149 ( .A1(n28684), .A2(n18476), .ZN(n28686) );
  OAI21_X2 U35816 ( .A1(n36490), .A2(n18048), .B(n18093), .ZN(n36241) );
  NAND2_X2 U7150 ( .A1(n40401), .A2(n40400), .ZN(n41423) );
  NAND3_X1 U13834 ( .A1(n40454), .A2(n40453), .A3(n1691), .ZN(n59518) );
  NOR2_X1 U30164 ( .A1(n40836), .A2(n40837), .ZN(n59103) );
  BUF_X2 U9788 ( .I(Key[173]), .Z(n56819) );
  INV_X2 U9063 ( .I(n28025), .ZN(n21154) );
  BUF_X2 U10397 ( .I(n32346), .Z(n23693) );
  BUF_X2 U4365 ( .I(n52719), .Z(n21066) );
  INV_X2 U11929 ( .I(n56629), .ZN(n56216) );
  INV_X2 U16874 ( .I(n43029), .ZN(n42777) );
  NAND2_X2 U5102 ( .A1(n15040), .A2(n1371), .ZN(n54447) );
  NAND3_X2 U45776 ( .A1(n30480), .A2(n30481), .A3(n19451), .ZN(n30484) );
  INV_X4 U3747 ( .I(n24078), .ZN(n36061) );
  BUF_X4 U35452 ( .I(n22939), .Z(n21644) );
  NOR2_X2 U23591 ( .A1(n58651), .A2(n30538), .ZN(n9186) );
  INV_X4 U9512 ( .I(n1786), .ZN(n1338) );
  NAND2_X2 U35481 ( .A1(n37772), .A2(n41894), .ZN(n16358) );
  NOR3_X2 U2570 ( .A1(n7534), .A2(n21008), .A3(n1424), .ZN(n34991) );
  NAND2_X2 U6520 ( .A1(n15545), .A2(n24571), .ZN(n34448) );
  OAI21_X2 U11050 ( .A1(n43061), .A2(n39937), .B(n22112), .ZN(n39944) );
  BUF_X4 U15595 ( .I(n50378), .Z(n5282) );
  NAND2_X2 U22365 ( .A1(n61052), .A2(n1208), .ZN(n21486) );
  NAND4_X2 U33998 ( .A1(n48313), .A2(n49309), .A3(n49597), .A4(n59084), .ZN(
        n9384) );
  NAND2_X2 U50107 ( .A1(n59203), .A2(n38932), .ZN(n40771) );
  INV_X2 U9863 ( .I(n64753), .ZN(n36454) );
  INV_X1 U17478 ( .I(n25214), .ZN(n58492) );
  NOR2_X2 U3679 ( .A1(n29952), .A2(n30647), .ZN(n59317) );
  BUF_X4 U27869 ( .I(n3376), .Z(n61509) );
  INV_X2 U9646 ( .I(n29884), .ZN(n30220) );
  NAND2_X2 U17828 ( .A1(n25152), .A2(n18215), .ZN(n12862) );
  NAND2_X2 U10264 ( .A1(n41185), .A2(n41184), .ZN(n41187) );
  AND2_X2 U5037 ( .A1(n14584), .A2(n64714), .Z(n2456) );
  NAND4_X1 U5471 ( .A1(n7444), .A2(n31257), .A3(n31258), .A4(n31256), .ZN(n270) );
  NOR2_X2 U4485 ( .A1(n18864), .A2(n18863), .ZN(n13786) );
  AOI21_X2 U15430 ( .A1(n10740), .A2(n48315), .B(n62244), .ZN(n18864) );
  NAND2_X2 U17355 ( .A1(n40573), .A2(n40571), .ZN(n15199) );
  INV_X2 U2048 ( .I(n3295), .ZN(n41082) );
  NAND4_X2 U56233 ( .A1(n55636), .A2(n55635), .A3(n55634), .A4(n55633), .ZN(
        n55637) );
  INV_X4 U41520 ( .I(n36178), .ZN(n36423) );
  INV_X2 U9930 ( .I(n48491), .ZN(n7911) );
  NAND2_X2 U1908 ( .A1(n43428), .A2(n42371), .ZN(n58059) );
  NAND2_X1 U26360 ( .A1(n6709), .A2(n30394), .ZN(n6708) );
  NAND2_X1 U30414 ( .A1(n6708), .A2(n59658), .ZN(n59685) );
  INV_X1 U26363 ( .I(n12480), .ZN(n12479) );
  AOI22_X2 U28191 ( .A1(n36307), .A2(n36306), .B1(n24351), .B2(n36305), .ZN(
        n58873) );
  OAI21_X2 U48754 ( .A1(n36304), .A2(n21605), .B(n60925), .ZN(n36306) );
  NAND2_X2 U2371 ( .A1(n37034), .A2(n25671), .ZN(n14915) );
  NAND3_X2 U265 ( .A1(n20018), .A2(n20017), .A3(n18750), .ZN(n594) );
  INV_X2 U1534 ( .I(n10827), .ZN(n43814) );
  NOR2_X2 U15727 ( .A1(n11293), .A2(n11292), .ZN(n11291) );
  NOR2_X2 U55302 ( .A1(n54015), .A2(n53035), .ZN(n54343) );
  BUF_X2 U14251 ( .I(n28230), .Z(n10537) );
  NOR2_X2 U11683 ( .A1(n47918), .A2(n3971), .ZN(n11184) );
  INV_X1 U50542 ( .I(n29281), .ZN(n60990) );
  BUF_X4 U5256 ( .I(Key[11]), .Z(n52232) );
  NOR2_X2 U4178 ( .A1(n22124), .A2(n54697), .ZN(n22123) );
  INV_X2 U27009 ( .I(n46918), .ZN(n44200) );
  INV_X2 U36470 ( .I(n34446), .ZN(n34442) );
  INV_X4 U3955 ( .I(n23217), .ZN(n14103) );
  INV_X8 U17994 ( .I(n37945), .ZN(n12050) );
  NAND2_X2 U3475 ( .A1(n7534), .A2(n57304), .ZN(n34073) );
  NAND3_X2 U6332 ( .A1(n53027), .A2(n53026), .A3(n59739), .ZN(n53029) );
  BUF_X4 U8453 ( .I(n36595), .Z(n22632) );
  BUF_X4 U18927 ( .I(n20308), .Z(n19388) );
  NAND3_X1 U44994 ( .A1(n28456), .A2(n28455), .A3(n28454), .ZN(n28457) );
  NAND2_X1 U18754 ( .A1(n537), .A2(n536), .ZN(n57864) );
  INV_X4 U2551 ( .I(n34165), .ZN(n14107) );
  NAND2_X2 U7080 ( .A1(n60659), .A2(n22524), .ZN(n8487) );
  BUF_X2 U19832 ( .I(n27859), .Z(n20872) );
  INV_X1 U10763 ( .I(n51632), .ZN(n54651) );
  INV_X2 U11488 ( .I(n59825), .ZN(n37018) );
  NOR3_X2 U5344 ( .A1(n317), .A2(n15177), .A3(n15605), .ZN(n7075) );
  NAND2_X2 U44896 ( .A1(n22556), .A2(n29988), .ZN(n28696) );
  NAND2_X2 U47869 ( .A1(n34513), .A2(n2033), .ZN(n33484) );
  INV_X4 U26504 ( .I(n21314), .ZN(n22556) );
  NAND2_X2 U4179 ( .A1(n58463), .A2(n21470), .ZN(n55641) );
  BUF_X4 U5198 ( .I(n37917), .Z(n4274) );
  INV_X2 U31636 ( .I(n18878), .ZN(n35666) );
  NAND2_X2 U9758 ( .A1(n29155), .A2(n6522), .ZN(n21589) );
  OAI21_X2 U10240 ( .A1(n15870), .A2(n35892), .B(n35568), .ZN(n13300) );
  NAND2_X2 U1696 ( .A1(n43225), .A2(n10203), .ZN(n43098) );
  NOR3_X2 U9470 ( .A1(n8680), .A2(n6122), .A3(n34883), .ZN(n6121) );
  BUF_X4 U14574 ( .I(n53729), .Z(n17286) );
  INV_X2 U32836 ( .I(n12799), .ZN(n50892) );
  BUF_X4 U11382 ( .I(n23600), .Z(n17583) );
  INV_X8 U9278 ( .I(n7854), .ZN(n48644) );
  INV_X2 U9321 ( .I(n1020), .ZN(n16649) );
  NAND2_X2 U10127 ( .A1(n6855), .A2(n41884), .ZN(n2895) );
  BUF_X4 U18911 ( .I(n31985), .Z(n23096) );
  BUF_X4 U28699 ( .I(n10205), .Z(n8602) );
  NOR3_X2 U27147 ( .A1(n57006), .A2(n1602), .A3(n6943), .ZN(n470) );
  NAND2_X2 U4377 ( .A1(n55696), .A2(n51961), .ZN(n17979) );
  NAND3_X1 U49480 ( .A1(n4276), .A2(n37915), .A3(n37914), .ZN(n37922) );
  OAI21_X2 U23593 ( .A1(n61557), .A2(n13094), .B(n42251), .ZN(n60901) );
  BUF_X4 U33792 ( .I(n16382), .Z(n14230) );
  NAND3_X1 U51929 ( .A1(n20281), .A2(n36749), .A3(n23648), .ZN(n20934) );
  INV_X2 U23349 ( .I(n7976), .ZN(n4457) );
  INV_X1 U5447 ( .I(n60851), .ZN(n58688) );
  INV_X1 U4561 ( .I(n41743), .ZN(n18770) );
  INV_X2 U3290 ( .I(n23191), .ZN(n26605) );
  INV_X4 U2624 ( .I(n14994), .ZN(n40755) );
  BUF_X4 U17476 ( .I(n61659), .Z(n23698) );
  BUF_X4 U14270 ( .I(n26459), .Z(n27621) );
  BUF_X4 U18839 ( .I(n17758), .Z(n5009) );
  NAND2_X1 U18288 ( .A1(n18896), .A2(n2390), .ZN(n2389) );
  NAND2_X2 U6587 ( .A1(n48027), .A2(n61170), .ZN(n58209) );
  INV_X2 U15554 ( .I(n48315), .ZN(n48027) );
  AOI22_X2 U18430 ( .A1(n34616), .A2(n34615), .B1(n34613), .B2(n34614), .ZN(
        n15229) );
  NOR2_X2 U11651 ( .A1(n2346), .A2(n34185), .ZN(n34190) );
  NOR2_X2 U3572 ( .A1(n52784), .A2(n23921), .ZN(n4119) );
  OAI22_X2 U55185 ( .A1(n52781), .A2(n52780), .B1(n4481), .B2(n53614), .ZN(
        n52784) );
  NAND2_X2 U55153 ( .A1(n23074), .A2(n64230), .ZN(n52729) );
  NOR3_X1 U6273 ( .A1(n17116), .A2(n17114), .A3(n30520), .ZN(n17525) );
  NAND2_X2 U124 ( .A1(n59610), .A2(n63520), .ZN(n52309) );
  INV_X2 U41598 ( .I(n55463), .ZN(n52933) );
  NOR2_X1 U1027 ( .A1(n46076), .A2(n44562), .ZN(n44567) );
  NAND3_X2 U13932 ( .A1(n1860), .A2(n11565), .A3(n1277), .ZN(n13572) );
  NAND3_X2 U5855 ( .A1(n10676), .A2(n20109), .A3(n10675), .ZN(n377) );
  OAI21_X2 U6365 ( .A1(n11023), .A2(n57291), .B(n55301), .ZN(n55305) );
  AOI21_X2 U8062 ( .A1(n39861), .A2(n42996), .B(n60472), .ZN(n4431) );
  NOR2_X2 U9359 ( .A1(n20922), .A2(n1499), .ZN(n41610) );
  AOI21_X2 U12889 ( .A1(n5364), .A2(n12355), .B(n62435), .ZN(n4409) );
  OAI21_X1 U11586 ( .A1(n34561), .A2(n10944), .B(n10942), .ZN(n34562) );
  INV_X4 U25311 ( .I(n49005), .ZN(n5629) );
  INV_X4 U30361 ( .I(n13655), .ZN(n22905) );
  INV_X4 U2725 ( .I(n16451), .ZN(n34784) );
  NAND2_X2 U2302 ( .A1(n37361), .A2(n20124), .ZN(n37289) );
  INV_X2 U28201 ( .I(n20517), .ZN(n46753) );
  OAI21_X2 U4184 ( .A1(n53067), .A2(n62412), .B(n53108), .ZN(n53106) );
  INV_X2 U10816 ( .I(n46493), .ZN(n2109) );
  INV_X1 U6616 ( .I(n63051), .ZN(n33948) );
  INV_X1 U6961 ( .I(n28040), .ZN(n28033) );
  NAND3_X1 U27024 ( .A1(n48229), .A2(n48231), .A3(n61715), .ZN(n14772) );
  INV_X2 U2601 ( .I(n22278), .ZN(n21464) );
  NAND4_X1 U41989 ( .A1(n25684), .A2(n25683), .A3(n55116), .A4(n25682), .ZN(
        n25681) );
  INV_X2 U3079 ( .I(n8336), .ZN(n22164) );
  NAND2_X2 U51106 ( .A1(n61894), .A2(n41564), .ZN(n41566) );
  OAI21_X2 U27526 ( .A1(n971), .A2(n23046), .B(n40571), .ZN(n40432) );
  INV_X2 U21558 ( .I(n42288), .ZN(n3078) );
  CLKBUF_X8 U13433 ( .I(n10717), .Z(n7028) );
  NAND2_X2 U30532 ( .A1(n26306), .A2(n26307), .ZN(n23580) );
  AOI22_X2 U36775 ( .A1(n16979), .A2(n30190), .B1(n30096), .B2(n22799), .ZN(
        n26306) );
  CLKBUF_X8 U14556 ( .I(n52287), .Z(n1583) );
  INV_X2 U15004 ( .I(n24749), .ZN(n1603) );
  OAI21_X1 U41558 ( .A1(n30274), .A2(n30275), .B(n30273), .ZN(n30282) );
  NAND3_X2 U2275 ( .A1(n36201), .A2(n36207), .A3(n1418), .ZN(n34941) );
  NOR2_X1 U13235 ( .A1(n14029), .A2(n8534), .ZN(n8533) );
  NAND4_X1 U42345 ( .A1(n45164), .A2(n48889), .A3(n45163), .A4(n45162), .ZN(
        n45170) );
  NAND3_X2 U52257 ( .A1(n46025), .A2(n46017), .A3(n20666), .ZN(n44943) );
  NOR2_X2 U28820 ( .A1(n48980), .A2(n48981), .ZN(n48987) );
  AOI21_X2 U53721 ( .A1(n48979), .A2(n48978), .B(n48977), .ZN(n48981) );
  AOI21_X2 U17393 ( .A1(n57750), .A2(n62213), .B(n62234), .ZN(n29159) );
  NOR2_X2 U319 ( .A1(n19068), .A2(n52845), .ZN(n25456) );
  BUF_X4 U2027 ( .I(n43845), .Z(n60052) );
  AND3_X1 U6887 ( .A1(n8759), .A2(n8761), .A3(n36120), .Z(n707) );
  INV_X1 U27598 ( .I(n49060), .ZN(n2697) );
  CLKBUF_X4 U42681 ( .I(n52189), .Z(n55474) );
  CLKBUF_X8 U9710 ( .I(n26429), .Z(n30786) );
  INV_X1 U2286 ( .I(n21915), .ZN(n15582) );
  INV_X2 U31573 ( .I(n46753), .ZN(n48545) );
  NAND2_X2 U11968 ( .A1(n17046), .A2(n21956), .ZN(n27967) );
  INV_X4 U26675 ( .I(n7376), .ZN(n30841) );
  BUF_X4 U20732 ( .I(n10079), .Z(n2483) );
  INV_X1 U37890 ( .I(n24733), .ZN(n46229) );
  NAND2_X1 U30964 ( .A1(n50413), .A2(n59227), .ZN(n50938) );
  NAND3_X2 U14828 ( .A1(n39168), .A2(n39166), .A3(n39167), .ZN(n39169) );
  INV_X4 U4287 ( .I(n40064), .ZN(n42433) );
  NAND2_X2 U22710 ( .A1(n4034), .A2(n32807), .ZN(n33690) );
  BUF_X2 U16389 ( .I(n23067), .Z(n5011) );
  OAI21_X1 U44669 ( .A1(n30727), .A2(n28773), .B(n29036), .ZN(n27515) );
  NOR3_X1 U5777 ( .A1(n2855), .A2(n39799), .A3(n2854), .ZN(n2853) );
  INV_X4 U2461 ( .I(n36955), .ZN(n13983) );
  INV_X1 U32490 ( .I(n59786), .ZN(n19716) );
  NAND2_X2 U11483 ( .A1(n36781), .A2(n19368), .ZN(n34362) );
  NOR2_X2 U56536 ( .A1(n20587), .A2(n21860), .ZN(n56523) );
  AOI21_X1 U36259 ( .A1(n53853), .A2(n18499), .B(n53852), .ZN(n53854) );
  INV_X2 U18741 ( .I(n35629), .ZN(n1811) );
  NOR2_X2 U32887 ( .A1(n49374), .A2(n58983), .ZN(n49532) );
  NAND4_X1 U18991 ( .A1(n2103), .A2(n29990), .A3(n29989), .A4(n61052), .ZN(
        n2102) );
  AOI21_X1 U55859 ( .A1(n61630), .A2(n25462), .B(n447), .ZN(n61330) );
  NOR2_X1 U19398 ( .A1(n27654), .A2(n5770), .ZN(n5769) );
  INV_X4 U32346 ( .I(n17240), .ZN(n31842) );
  INV_X4 U17535 ( .I(n57762), .ZN(n48254) );
  BUF_X2 U18760 ( .I(n32828), .Z(n10277) );
  INV_X1 U26655 ( .I(n33573), .ZN(n18549) );
  INV_X2 U24089 ( .I(n21938), .ZN(n6051) );
  INV_X2 U30122 ( .I(n12798), .ZN(n10907) );
  INV_X4 U31139 ( .I(n8986), .ZN(n21851) );
  OR2_X1 U10470 ( .A1(n16971), .A2(n3478), .Z(n29059) );
  NAND2_X2 U1485 ( .A1(n14518), .A2(n48460), .ZN(n47084) );
  INV_X2 U2733 ( .I(n35710), .ZN(n34404) );
  NAND2_X2 U33773 ( .A1(n29564), .A2(n14213), .ZN(n29912) );
  BUF_X4 U34067 ( .I(n36979), .Z(n59617) );
  OR2_X2 U19229 ( .A1(n30288), .A2(n23317), .Z(n30273) );
  NOR2_X2 U48898 ( .A1(n36781), .A2(n37268), .ZN(n36782) );
  NOR2_X2 U49472 ( .A1(n52283), .A2(n52284), .ZN(n60961) );
  NOR2_X2 U32679 ( .A1(n37454), .A2(n10907), .ZN(n36975) );
  BUF_X4 U10005 ( .I(n6604), .Z(n2823) );
  NOR2_X1 U36840 ( .A1(n28577), .A2(n30562), .ZN(n25381) );
  NAND2_X2 U2978 ( .A1(n24504), .A2(n30430), .ZN(n28574) );
  INV_X4 U488 ( .I(n52270), .ZN(n56978) );
  INV_X2 U8702 ( .I(n15280), .ZN(n1270) );
  NAND2_X2 U703 ( .A1(n9408), .A2(n49726), .ZN(n2502) );
  NOR2_X2 U10161 ( .A1(n42433), .A2(n62291), .ZN(n40310) );
  INV_X2 U9357 ( .I(n13493), .ZN(n43270) );
  NAND2_X2 U25410 ( .A1(n43476), .A2(n12312), .ZN(n42411) );
  INV_X4 U11538 ( .I(n10717), .ZN(n15794) );
  NAND3_X2 U39877 ( .A1(n19905), .A2(n16163), .A3(n56596), .ZN(n19446) );
  NAND2_X2 U22878 ( .A1(n1381), .A2(n4174), .ZN(n50410) );
  INV_X1 U24431 ( .I(n29343), .ZN(n58546) );
  INV_X2 U45778 ( .I(n30490), .ZN(n30491) );
  INV_X4 U11768 ( .I(n52530), .ZN(n1619) );
  INV_X2 U2761 ( .I(n62045), .ZN(n23947) );
  NOR2_X1 U4434 ( .A1(n53854), .A2(n53867), .ZN(n2852) );
  BUF_X4 U41916 ( .I(n33709), .Z(n35962) );
  OR2_X2 U416 ( .A1(n22105), .A2(n53615), .Z(n53421) );
  NAND2_X1 U29558 ( .A1(n707), .A2(n8764), .ZN(n37581) );
  BUF_X4 U9050 ( .I(n26375), .Z(n29154) );
  AOI21_X2 U53495 ( .A1(n48215), .A2(n48666), .B(n48214), .ZN(n48216) );
  NOR2_X2 U10939 ( .A1(n47196), .A2(n19804), .ZN(n46996) );
  INV_X2 U27278 ( .I(n45053), .ZN(n44907) );
  AOI21_X2 U19063 ( .A1(n13765), .A2(n28090), .B(n13571), .ZN(n8701) );
  INV_X2 U25981 ( .I(n18571), .ZN(n6322) );
  INV_X4 U2080 ( .I(n14863), .ZN(n42432) );
  NAND3_X1 U3765 ( .A1(n34373), .A2(n36161), .A3(n37373), .ZN(n34381) );
  NAND4_X1 U4104 ( .A1(n56470), .A2(n56469), .A3(n56468), .A4(n56467), .ZN(
        n57919) );
  NAND2_X2 U56543 ( .A1(n23920), .A2(n21859), .ZN(n56456) );
  NAND2_X1 U46704 ( .A1(n31731), .A2(n31728), .ZN(n31729) );
  INV_X2 U5241 ( .I(n3270), .ZN(n47518) );
  INV_X4 U12187 ( .I(n53677), .ZN(n53695) );
  BUF_X4 U5978 ( .I(n23472), .Z(n61417) );
  OAI21_X2 U53783 ( .A1(n6896), .A2(n49176), .B(n21367), .ZN(n49180) );
  INV_X8 U6499 ( .I(n49195), .ZN(n3694) );
  NOR2_X2 U15192 ( .A1(n49621), .A2(n49617), .ZN(n46856) );
  NAND3_X2 U12990 ( .A1(n3728), .A2(n3726), .A3(n3725), .ZN(n22972) );
  NOR2_X2 U4756 ( .A1(n11771), .A2(n11770), .ZN(n11769) );
  OAI22_X2 U19111 ( .A1(n25930), .A2(n48213), .B1(n48211), .B2(n48212), .ZN(
        n48214) );
  AOI21_X1 U17036 ( .A1(n6875), .A2(n41222), .B(n6874), .ZN(n6880) );
  NOR4_X1 U44835 ( .A1(n27886), .A2(n30854), .A3(n24556), .A4(n29905), .ZN(
        n27899) );
  INV_X4 U38914 ( .I(n18068), .ZN(n18333) );
  NAND2_X2 U15906 ( .A1(n47463), .A2(n45748), .ZN(n2812) );
  NAND2_X1 U36398 ( .A1(n33298), .A2(n35683), .ZN(n25101) );
  AOI22_X2 U18901 ( .A1(n3263), .A2(n16140), .B1(n27804), .B2(n3261), .ZN(
        n16440) );
  NOR3_X1 U15346 ( .A1(n7013), .A2(n2075), .A3(n5812), .ZN(n2071) );
  NAND3_X2 U4517 ( .A1(n54715), .A2(n59095), .A3(n59094), .ZN(n60752) );
  INV_X2 U32344 ( .I(n17873), .ZN(n17874) );
  INV_X2 U41306 ( .I(n25876), .ZN(n26023) );
  BUF_X4 U8267 ( .I(n16490), .Z(n1866) );
  BUF_X4 U4148 ( .I(n1133), .Z(n13920) );
  NOR2_X1 U15294 ( .A1(n7002), .A2(n49311), .ZN(n7001) );
  NAND2_X1 U14497 ( .A1(n63020), .A2(n2475), .ZN(n2474) );
  NAND2_X2 U2453 ( .A1(n14054), .A2(n7729), .ZN(n14331) );
  OAI22_X1 U50688 ( .A1(n40222), .A2(n40221), .B1(n40220), .B2(n9091), .ZN(
        n40227) );
  NAND2_X2 U6305 ( .A1(n59108), .A2(n55628), .ZN(n10988) );
  NOR2_X2 U8608 ( .A1(n16438), .A2(n47367), .ZN(n16437) );
  NAND2_X2 U24013 ( .A1(n19243), .A2(n49910), .ZN(n48340) );
  OR3_X2 U4175 ( .A1(n56792), .A2(n58688), .A3(n65064), .Z(n56800) );
  INV_X4 U5216 ( .I(n25348), .ZN(n46279) );
  NAND4_X1 U23792 ( .A1(n17360), .A2(n17359), .A3(n17363), .A4(n56826), .ZN(
        n58474) );
  NAND2_X2 U13635 ( .A1(n34583), .A2(n2346), .ZN(n33435) );
  BUF_X4 U42712 ( .I(n39324), .Z(n23752) );
  NAND2_X2 U17839 ( .A1(n35955), .A2(n15409), .ZN(n15411) );
  OAI21_X2 U34185 ( .A1(n35954), .A2(n14743), .B(n36923), .ZN(n15409) );
  NOR3_X1 U15599 ( .A1(n16414), .A2(n57626), .A3(n16413), .ZN(n16412) );
  INV_X1 U34390 ( .I(n15092), .ZN(n21955) );
  NAND4_X1 U6285 ( .A1(n53075), .A2(n53074), .A3(n53073), .A4(n53072), .ZN(
        n60495) );
  BUF_X4 U3108 ( .I(n37363), .Z(n60980) );
  BUF_X2 U2123 ( .I(n18545), .Z(n12669) );
  NAND2_X2 U7157 ( .A1(n42536), .A2(n42534), .ZN(n58538) );
  INV_X2 U5748 ( .I(n47535), .ZN(n60343) );
  NAND2_X2 U16542 ( .A1(n5104), .A2(n43097), .ZN(n5103) );
  INV_X1 U33135 ( .I(n26150), .ZN(n13245) );
  INV_X4 U1249 ( .I(n2344), .ZN(n47535) );
  NAND2_X2 U3219 ( .A1(n28030), .A2(n61177), .ZN(n6137) );
  NAND2_X2 U31715 ( .A1(n11386), .A2(n38406), .ZN(n59315) );
  AOI21_X2 U17715 ( .A1(n17947), .A2(n36200), .B(n9769), .ZN(n16682) );
  NAND3_X2 U35278 ( .A1(n10596), .A2(n1779), .A3(n35883), .ZN(n35568) );
  INV_X2 U11020 ( .I(n44861), .ZN(n1669) );
  NAND3_X2 U29040 ( .A1(n35828), .A2(n23556), .A3(n16919), .ZN(n58961) );
  AOI22_X2 U41817 ( .A1(n22552), .A2(n10226), .B1(n32143), .B2(n37333), .ZN(
        n32148) );
  OAI21_X1 U36110 ( .A1(n47856), .A2(n47855), .B(n70), .ZN(n47866) );
  NAND3_X1 U9113 ( .A1(n24866), .A2(n9867), .A3(n9866), .ZN(n24865) );
  INV_X4 U25470 ( .I(n33623), .ZN(n33644) );
  OAI21_X1 U4557 ( .A1(n6399), .A2(n6397), .B(n33537), .ZN(n12749) );
  NOR3_X1 U7018 ( .A1(n29278), .A2(n24896), .A3(n4103), .ZN(n4102) );
  NAND2_X1 U18347 ( .A1(n33381), .A2(n33379), .ZN(n3860) );
  INV_X1 U37023 ( .I(n44905), .ZN(n17729) );
  INV_X4 U22442 ( .I(n58205), .ZN(n3772) );
  NOR2_X2 U17724 ( .A1(n17911), .A2(n22968), .ZN(n4449) );
  CLKBUF_X8 U13206 ( .I(n20620), .Z(n11239) );
  INV_X1 U42537 ( .I(n23286), .ZN(n28004) );
  INV_X4 U12941 ( .I(n16982), .ZN(n8962) );
  INV_X2 U27811 ( .I(n7721), .ZN(n26113) );
  BUF_X2 U1523 ( .I(n20897), .Z(n60390) );
  BUF_X4 U4721 ( .I(n14335), .Z(n7824) );
  OAI21_X2 U1020 ( .A1(n48048), .A2(n20460), .B(n57574), .ZN(n48050) );
  NAND2_X2 U23458 ( .A1(n59647), .A2(n59646), .ZN(n59157) );
  OAI21_X2 U10132 ( .A1(n39117), .A2(n38421), .B(n41014), .ZN(n37533) );
  NAND3_X2 U11110 ( .A1(n41538), .A2(n41539), .A3(n61372), .ZN(n9724) );
  INV_X2 U13651 ( .I(n53161), .ZN(n53167) );
  NAND2_X2 U32855 ( .A1(n41027), .A2(n36106), .ZN(n39097) );
  NAND2_X1 U18217 ( .A1(n10119), .A2(n10118), .ZN(n22339) );
  INV_X2 U13450 ( .I(n37184), .ZN(n37335) );
  NAND3_X1 U15564 ( .A1(n32023), .A2(n20819), .A3(n16267), .ZN(n59603) );
  BUF_X4 U11342 ( .I(n1238), .Z(n23986) );
  OAI21_X2 U747 ( .A1(n5806), .A2(n24374), .B(n50267), .ZN(n5805) );
  NOR2_X1 U24485 ( .A1(n10355), .A2(n10354), .ZN(n13871) );
  NOR2_X1 U11733 ( .A1(n12414), .A2(n8461), .ZN(n8460) );
  INV_X2 U2722 ( .I(n65205), .ZN(n35321) );
  AOI21_X2 U15370 ( .A1(n48292), .A2(n21335), .B(n21333), .ZN(n23910) );
  INV_X2 U6331 ( .I(n63473), .ZN(n57201) );
  NAND2_X2 U900 ( .A1(n64764), .A2(n47073), .ZN(n60983) );
  NAND2_X2 U9560 ( .A1(n3691), .A2(n37224), .ZN(n3693) );
  NAND2_X1 U6607 ( .A1(n7782), .A2(n57465), .ZN(n7779) );
  INV_X2 U35752 ( .I(n37270), .ZN(n37491) );
  OR2_X2 U3298 ( .A1(n27366), .A2(n28221), .Z(n28002) );
  NAND3_X2 U10327 ( .A1(n5261), .A2(n43012), .A3(n42327), .ZN(n58777) );
  INV_X4 U3002 ( .I(n18306), .ZN(n20859) );
  OAI21_X2 U44496 ( .A1(n28007), .A2(n180), .B(n1893), .ZN(n27090) );
  NOR3_X2 U21585 ( .A1(n27728), .A2(n27729), .A3(n27730), .ZN(n27732) );
  NOR2_X2 U1950 ( .A1(n20397), .A2(n20396), .ZN(n20395) );
  NAND3_X1 U55562 ( .A1(n53832), .A2(n53831), .A3(n53830), .ZN(n53834) );
  INV_X8 U7175 ( .I(n12034), .ZN(n20242) );
  NOR3_X2 U37149 ( .A1(n44662), .A2(n19747), .A3(n48337), .ZN(n19746) );
  NAND3_X2 U669 ( .A1(n15467), .A2(n5657), .A3(n15473), .ZN(n58834) );
  BUF_X4 U39948 ( .I(n19059), .Z(n60202) );
  INV_X2 U17443 ( .I(n24931), .ZN(n39994) );
  INV_X2 U39572 ( .I(n40020), .ZN(n43433) );
  AOI22_X2 U6337 ( .A1(n4224), .A2(n53860), .B1(n4222), .B2(n53024), .ZN(
        n60425) );
  CLKBUF_X4 U15076 ( .I(n48060), .Z(n54025) );
  NOR2_X2 U14871 ( .A1(n1456), .A2(n61870), .ZN(n8057) );
  INV_X4 U3422 ( .I(n21087), .ZN(n21956) );
  NAND2_X1 U298 ( .A1(n20933), .A2(n54602), .ZN(n59507) );
  NAND2_X1 U15546 ( .A1(n6670), .A2(n54342), .ZN(n6674) );
  NAND3_X2 U5986 ( .A1(n2812), .A2(n45741), .A3(n45744), .ZN(n2811) );
  INV_X2 U9347 ( .I(n43898), .ZN(n7516) );
  NAND2_X2 U14770 ( .A1(n56575), .A2(n62769), .ZN(n57551) );
  INV_X2 U19282 ( .I(n29502), .ZN(n1840) );
  NAND2_X2 U9436 ( .A1(n7012), .A2(n7011), .ZN(n8201) );
  NOR2_X2 U54943 ( .A1(n61255), .A2(n27394), .ZN(n3710) );
  INV_X4 U3239 ( .I(n22726), .ZN(n27390) );
  NAND2_X2 U16810 ( .A1(n43120), .A2(n43270), .ZN(n41789) );
  NAND2_X2 U7289 ( .A1(n8962), .A2(n43124), .ZN(n43120) );
  BUF_X4 U11894 ( .I(n22106), .Z(n10629) );
  NOR2_X2 U22809 ( .A1(n2394), .A2(n2392), .ZN(n2400) );
  NOR2_X1 U681 ( .A1(n6898), .A2(n10070), .ZN(n4373) );
  NAND4_X2 U48908 ( .A1(n36813), .A2(n36812), .A3(n36811), .A4(n36810), .ZN(
        n36814) );
  INV_X2 U962 ( .I(n7358), .ZN(n49545) );
  NOR2_X1 U266 ( .A1(n19477), .A2(n53544), .ZN(n19476) );
  OAI22_X2 U15784 ( .A1(n10590), .A2(n47871), .B1(n12738), .B2(n43827), .ZN(
        n47872) );
  AOI21_X2 U8643 ( .A1(n43680), .A2(n22553), .B(n43681), .ZN(n25877) );
  NAND3_X2 U48705 ( .A1(n60980), .A2(n10087), .A3(n592), .ZN(n36167) );
  INV_X4 U11305 ( .I(n40804), .ZN(n41894) );
  INV_X4 U28620 ( .I(n28711), .ZN(n8522) );
  NAND2_X2 U14078 ( .A1(n27433), .A2(n26468), .ZN(n26602) );
  NAND2_X2 U43389 ( .A1(n17283), .A2(n60801), .ZN(n12822) );
  INV_X2 U17889 ( .I(n22116), .ZN(n35549) );
  NAND2_X2 U11432 ( .A1(n6612), .A2(n34888), .ZN(n34889) );
  OAI22_X2 U27606 ( .A1(n54009), .A2(n54010), .B1(n60426), .B2(n54007), .ZN(
        n59872) );
  OAI21_X1 U50715 ( .A1(n40297), .A2(n14014), .B(n40293), .ZN(n40302) );
  AND2_X1 U25192 ( .A1(n9596), .A2(n9597), .Z(n2187) );
  AOI21_X1 U1831 ( .A1(n40166), .A2(n11130), .B(n11128), .ZN(n11127) );
  AOI21_X1 U11100 ( .A1(n42029), .A2(n42028), .B(n42035), .ZN(n2709) );
  INV_X1 U27890 ( .I(n7834), .ZN(n48495) );
  INV_X4 U15027 ( .I(n53036), .ZN(n54026) );
  NAND2_X1 U54998 ( .A1(n52313), .A2(n52312), .ZN(n52314) );
  NAND3_X2 U28516 ( .A1(n61218), .A2(n16494), .A3(n50119), .ZN(n58920) );
  AND2_X2 U24412 ( .A1(n17661), .A2(n40839), .Z(n19358) );
  NOR2_X2 U328 ( .A1(n58784), .A2(n52222), .ZN(n8119) );
  AOI21_X1 U6711 ( .A1(n57705), .A2(n11903), .B(n11898), .ZN(n23565) );
  INV_X1 U13992 ( .I(n28711), .ZN(n3085) );
  NAND2_X2 U20300 ( .A1(n2149), .A2(n45935), .ZN(n45634) );
  BUF_X4 U15697 ( .I(n15595), .Z(n10422) );
  INV_X2 U2557 ( .I(n15819), .ZN(n1807) );
  BUF_X2 U3803 ( .I(n39306), .Z(n40028) );
  INV_X2 U42722 ( .I(n23301), .ZN(n48481) );
  INV_X2 U6758 ( .I(n3663), .ZN(n45966) );
  INV_X2 U20413 ( .I(n2225), .ZN(n26089) );
  NOR3_X2 U50741 ( .A1(n40378), .A2(n40377), .A3(n40376), .ZN(n40385) );
  BUF_X8 U5166 ( .I(n11359), .Z(n23127) );
  NAND2_X2 U16722 ( .A1(n43564), .A2(n11910), .ZN(n43422) );
  INV_X2 U22481 ( .I(n57603), .ZN(n47565) );
  INV_X2 U10725 ( .I(n64714), .ZN(n15355) );
  NAND2_X2 U11231 ( .A1(n3896), .A2(n40230), .ZN(n4642) );
  INV_X4 U6393 ( .I(n31804), .ZN(n19204) );
  INV_X1 U22399 ( .I(n7102), .ZN(n12918) );
  NAND2_X2 U2910 ( .A1(n37957), .A2(n15582), .ZN(n59117) );
  NAND2_X1 U14990 ( .A1(n23408), .A2(n58958), .ZN(n61136) );
  INV_X2 U17496 ( .I(n57173), .ZN(n3756) );
  NAND4_X2 U19511 ( .A1(n525), .A2(n524), .A3(n52969), .A4(n52968), .ZN(n57911) );
  NAND2_X1 U16819 ( .A1(n3126), .A2(n42359), .ZN(n23339) );
  BUF_X2 U7373 ( .I(n42016), .Z(n57557) );
  INV_X2 U1770 ( .I(n10945), .ZN(n42894) );
  NAND2_X2 U38454 ( .A1(n59522), .A2(n59328), .ZN(n33973) );
  NAND2_X2 U29571 ( .A1(n59910), .A2(n17096), .ZN(n16191) );
  OAI22_X2 U21654 ( .A1(n64234), .A2(n22333), .B1(n20607), .B2(n118), .ZN(
        n19253) );
  CLKBUF_X8 U8464 ( .I(n22997), .Z(n1253) );
  INV_X2 U23860 ( .I(n21624), .ZN(n24047) );
  INV_X1 U10764 ( .I(n53213), .ZN(n1372) );
  INV_X4 U1141 ( .I(n49768), .ZN(n49777) );
  INV_X1 U13167 ( .I(n57614), .ZN(n16921) );
  CLKBUF_X4 U14296 ( .I(Key[53]), .Z(n24061) );
  CLKBUF_X2 U9078 ( .I(Key[66]), .Z(n54360) );
  CLKBUF_X4 U14305 ( .I(Key[43]), .Z(n53787) );
  BUF_X2 U19904 ( .I(Key[117]), .Z(n24057) );
  BUF_X2 U12117 ( .I(Key[22]), .Z(n53359) );
  CLKBUF_X4 U44794 ( .I(Key[171]), .Z(n56784) );
  BUF_X2 U9083 ( .I(Key[180]), .Z(n56905) );
  CLKBUF_X4 U19940 ( .I(Key[168]), .Z(n51492) );
  CLKBUF_X4 U14317 ( .I(Key[156]), .Z(n24105) );
  BUF_X4 U10627 ( .I(n3385), .Z(n3117) );
  INV_X1 U43959 ( .I(n28317), .ZN(n26280) );
  CLKBUF_X2 U42289 ( .I(n28224), .Z(n23166) );
  INV_X2 U34084 ( .I(n27160), .ZN(n19522) );
  CLKBUF_X4 U41543 ( .I(n26293), .Z(n27114) );
  INV_X1 U1371 ( .I(n50494), .ZN(n1576) );
  CLKBUF_X4 U7981 ( .I(n26860), .Z(n28633) );
  BUF_X2 U19928 ( .I(n59130), .Z(n53102) );
  CLKBUF_X1 U24515 ( .I(n26826), .Z(n58559) );
  INV_X1 U1382 ( .I(n56905), .ZN(n18728) );
  CLKBUF_X2 U4816 ( .I(n61380), .Z(n54407) );
  CLKBUF_X4 U6779 ( .I(n6589), .Z(n3932) );
  CLKBUF_X4 U4895 ( .I(n24889), .Z(n15715) );
  INV_X2 U8544 ( .I(n16446), .ZN(n28379) );
  BUF_X2 U5798 ( .I(n26362), .Z(n27188) );
  CLKBUF_X2 U3976 ( .I(n24419), .Z(n61260) );
  CLKBUF_X2 U8491 ( .I(n27479), .Z(n23823) );
  CLKBUF_X4 U14264 ( .I(n26790), .Z(n28616) );
  CLKBUF_X4 U12080 ( .I(n28604), .Z(n23649) );
  INV_X2 U3349 ( .I(n27366), .ZN(n23716) );
  INV_X2 U28522 ( .I(n15093), .ZN(n21087) );
  CLKBUF_X2 U5457 ( .I(n27930), .Z(n266) );
  INV_X2 U10615 ( .I(n13079), .ZN(n1442) );
  BUF_X2 U9047 ( .I(n29972), .Z(n15735) );
  CLKBUF_X1 U19793 ( .I(n20508), .Z(n4617) );
  CLKBUF_X2 U4743 ( .I(n27380), .Z(n97) );
  INV_X2 U26509 ( .I(n22482), .ZN(n27976) );
  INV_X1 U14242 ( .I(n46398), .ZN(n1888) );
  INV_X2 U19767 ( .I(n24853), .ZN(n11110) );
  NAND2_X1 U21563 ( .A1(n27674), .A2(n20581), .ZN(n23937) );
  CLKBUF_X2 U56889 ( .I(n28327), .Z(n61484) );
  INV_X2 U37984 ( .I(n19679), .ZN(n28549) );
  CLKBUF_X2 U46910 ( .I(n29145), .Z(n60841) );
  CLKBUF_X4 U3971 ( .I(n243), .Z(n60265) );
  NOR2_X1 U12066 ( .A1(n28414), .A2(n1891), .ZN(n3254) );
  OR2_X1 U12974 ( .A1(n27522), .A2(n296), .Z(n57368) );
  INV_X1 U19618 ( .I(n28183), .ZN(n18824) );
  AND2_X1 U20560 ( .A1(n2342), .A2(n19679), .Z(n24967) );
  NAND2_X1 U44300 ( .A1(n26906), .A2(n28447), .ZN(n27860) );
  INV_X1 U14202 ( .I(n27592), .ZN(n28302) );
  OAI21_X1 U56517 ( .A1(n3409), .A2(n61387), .B(n29147), .ZN(n3407) );
  NAND2_X1 U14114 ( .A1(n27295), .A2(n26719), .ZN(n7024) );
  INV_X2 U3311 ( .I(n17047), .ZN(n18377) );
  NOR2_X1 U15401 ( .A1(n27386), .A2(n27042), .ZN(n57612) );
  NAND2_X1 U6231 ( .A1(n15358), .A2(n1884), .ZN(n26926) );
  AOI21_X1 U35361 ( .A1(n27120), .A2(n27121), .B(n1895), .ZN(n17722) );
  INV_X1 U11956 ( .I(n29698), .ZN(n3428) );
  NAND2_X1 U30324 ( .A1(n28618), .A2(n10084), .ZN(n28456) );
  OR3_X1 U37963 ( .A1(n26517), .A2(n61470), .A3(n60265), .Z(n26262) );
  NAND3_X1 U41243 ( .A1(n29156), .A2(n597), .A3(n65183), .ZN(n27259) );
  NOR2_X1 U11964 ( .A1(n29149), .A2(n65198), .ZN(n3828) );
  NAND2_X1 U8991 ( .A1(n24499), .A2(n21126), .ZN(n25732) );
  NAND2_X1 U40617 ( .A1(n26262), .A2(n26257), .ZN(n61144) );
  NAND3_X1 U11946 ( .A1(n4606), .A2(n19287), .A3(n28624), .ZN(n28468) );
  NOR2_X1 U3933 ( .A1(n26741), .A2(n9561), .ZN(n26747) );
  OAI21_X1 U57057 ( .A1(n60841), .A2(n26381), .B(n61599), .ZN(n15942) );
  INV_X1 U19615 ( .I(n16570), .ZN(n27539) );
  OAI21_X1 U44043 ( .A1(n27390), .A2(n27983), .B(n26377), .ZN(n26380) );
  NOR2_X1 U19449 ( .A1(n18263), .A2(n14152), .ZN(n14151) );
  NOR2_X1 U44620 ( .A1(n27351), .A2(n27350), .ZN(n27352) );
  NAND3_X1 U19476 ( .A1(n27317), .A2(n27316), .A3(n27315), .ZN(n27318) );
  NOR2_X1 U19451 ( .A1(n13377), .A2(n13374), .ZN(n13381) );
  NOR3_X1 U14057 ( .A1(n26838), .A2(n8888), .A3(n16516), .ZN(n19829) );
  NOR2_X1 U30710 ( .A1(n25453), .A2(n20760), .ZN(n25452) );
  NOR3_X1 U43243 ( .A1(n25732), .A2(n25733), .A3(n27385), .ZN(n25738) );
  NAND2_X1 U19586 ( .A1(n57915), .A2(n57249), .ZN(n57914) );
  CLKBUF_X4 U40131 ( .I(n30664), .Z(n19929) );
  BUF_X2 U14029 ( .I(n30730), .Z(n14729) );
  CLKBUF_X2 U38652 ( .I(n29457), .Z(n60028) );
  INV_X2 U33793 ( .I(n16382), .ZN(n23094) );
  CLKBUF_X1 U17858 ( .I(n13976), .Z(n57789) );
  AOI21_X1 U8624 ( .A1(n61054), .A2(n61053), .B(n61049), .ZN(n28020) );
  CLKBUF_X2 U37669 ( .I(n29726), .Z(n22748) );
  CLKBUF_X4 U19366 ( .I(n28948), .Z(n24097) );
  NAND2_X1 U19585 ( .A1(n18034), .A2(n57914), .ZN(n18033) );
  INV_X2 U3873 ( .I(n64169), .ZN(n57937) );
  CLKBUF_X4 U10498 ( .I(n17496), .Z(n8891) );
  CLKBUF_X2 U24522 ( .I(n29727), .Z(n58560) );
  CLKBUF_X4 U19378 ( .I(n64169), .Z(n24556) );
  CLKBUF_X4 U42497 ( .I(n29003), .Z(n23446) );
  CLKBUF_X2 U56730 ( .I(n20755), .Z(n61421) );
  INV_X2 U43302 ( .I(n24993), .ZN(n29773) );
  INV_X1 U13986 ( .I(n14334), .ZN(n30579) );
  BUF_X2 U8716 ( .I(n30338), .Z(n21029) );
  BUF_X1 U14893 ( .I(n29575), .Z(n57559) );
  NAND2_X2 U10493 ( .A1(n57789), .A2(n30588), .ZN(n31143) );
  INV_X1 U8945 ( .I(n29411), .ZN(n1859) );
  CLKBUF_X2 U38840 ( .I(n23708), .Z(n60064) );
  INV_X1 U10436 ( .I(n29050), .ZN(n30096) );
  INV_X2 U27820 ( .I(n12420), .ZN(n30078) );
  NOR2_X1 U32690 ( .A1(n14213), .A2(n31124), .ZN(n59452) );
  INV_X1 U45689 ( .I(n30277), .ZN(n30278) );
  NAND2_X1 U45192 ( .A1(n29729), .A2(n23315), .ZN(n28985) );
  NAND2_X1 U36070 ( .A1(n20364), .A2(n1351), .ZN(n30127) );
  NAND2_X1 U7011 ( .A1(n22893), .A2(n5631), .ZN(n28687) );
  OR2_X1 U15416 ( .A1(n5688), .A2(n61162), .Z(n9701) );
  INV_X1 U45575 ( .I(n29986), .ZN(n29987) );
  INV_X1 U45750 ( .I(n30422), .ZN(n30424) );
  NAND2_X1 U19021 ( .A1(n755), .A2(n27790), .ZN(n10580) );
  CLKBUF_X4 U51468 ( .I(n16961), .Z(n61052) );
  NAND3_X1 U45783 ( .A1(n30506), .A2(n30505), .A3(n30504), .ZN(n30507) );
  NAND3_X1 U35953 ( .A1(n30161), .A2(n30687), .A3(n30160), .ZN(n30162) );
  NAND2_X1 U38276 ( .A1(n30575), .A2(n59841), .ZN(n59987) );
  OAI22_X1 U17661 ( .A1(n57772), .A2(n57392), .B1(n29022), .B2(n29021), .ZN(
        n11864) );
  AOI21_X1 U18948 ( .A1(n5692), .A2(n12808), .B(n5691), .ZN(n5690) );
  NOR2_X1 U4713 ( .A1(n4736), .A2(n4735), .ZN(n13845) );
  AOI22_X1 U39630 ( .A1(n29013), .A2(n1554), .B1(n21251), .B2(n30071), .ZN(
        n20966) );
  NAND2_X1 U34547 ( .A1(n59685), .A2(n59684), .ZN(n59823) );
  OR3_X1 U14042 ( .A1(n29424), .A2(n29425), .A3(n19207), .Z(n58129) );
  AND2_X1 U27614 ( .A1(n7556), .A2(n30417), .Z(n22971) );
  NOR3_X1 U31912 ( .A1(n872), .A2(n9002), .A3(n59351), .ZN(n14475) );
  OAI21_X1 U53867 ( .A1(n30559), .A2(n30556), .B(n5136), .ZN(n4934) );
  NAND2_X1 U19019 ( .A1(n23080), .A2(n14109), .ZN(n6545) );
  AOI21_X1 U44584 ( .A1(n64694), .A2(n5653), .B(n29506), .ZN(n21414) );
  NAND2_X1 U23268 ( .A1(n6552), .A2(n30263), .ZN(n6551) );
  INV_X1 U18891 ( .I(n18120), .ZN(n4778) );
  INV_X1 U13752 ( .I(n22674), .ZN(n7568) );
  CLKBUF_X4 U11741 ( .I(n8109), .Z(n3523) );
  INV_X2 U39193 ( .I(n15155), .ZN(n24943) );
  INV_X2 U18845 ( .I(n7616), .ZN(n19993) );
  CLKBUF_X4 U18887 ( .I(n15816), .Z(n7522) );
  CLKBUF_X2 U18870 ( .I(n18434), .Z(n4795) );
  BUF_X2 U9612 ( .I(n32339), .Z(n23786) );
  INV_X1 U3633 ( .I(n33872), .ZN(n9374) );
  CLKBUF_X4 U3630 ( .I(n24730), .Z(n20573) );
  INV_X1 U10389 ( .I(n33048), .ZN(n13990) );
  INV_X2 U37739 ( .I(n7199), .ZN(n32338) );
  INV_X1 U13746 ( .I(n1313), .ZN(n13089) );
  INV_X1 U18829 ( .I(n32010), .ZN(n32059) );
  INV_X2 U33285 ( .I(n24943), .ZN(n13449) );
  INV_X2 U20956 ( .I(n2666), .ZN(n32544) );
  INV_X2 U11723 ( .I(n21509), .ZN(n1548) );
  INV_X1 U28652 ( .I(n32738), .ZN(n8558) );
  BUF_X2 U9375 ( .I(n24965), .Z(n10340) );
  CLKBUF_X4 U4493 ( .I(n32430), .Z(n34309) );
  BUF_X2 U6415 ( .I(n22316), .Z(n551) );
  CLKBUF_X4 U41878 ( .I(n31833), .Z(n35805) );
  CLKBUF_X2 U5366 ( .I(n33519), .Z(n24077) );
  CLKBUF_X4 U18743 ( .I(n31710), .Z(n34132) );
  CLKBUF_X2 U4860 ( .I(n889), .Z(n127) );
  CLKBUF_X2 U42834 ( .I(n33971), .Z(n23945) );
  CLKBUF_X4 U4853 ( .I(n32885), .Z(n15152) );
  CLKBUF_X2 U57056 ( .I(n33389), .Z(n61598) );
  CLKBUF_X4 U6151 ( .I(n23689), .Z(n60669) );
  CLKBUF_X4 U18728 ( .I(n33663), .Z(n22598) );
  CLKBUF_X4 U16778 ( .I(n34783), .Z(n57710) );
  BUF_X2 U27445 ( .I(n34585), .Z(n7453) );
  BUF_X2 U18720 ( .I(n14039), .Z(n22601) );
  INV_X2 U48145 ( .I(n35820), .ZN(n35813) );
  CLKBUF_X4 U18709 ( .I(n32512), .Z(n7359) );
  CLKBUF_X2 U52700 ( .I(n1815), .Z(n61108) );
  BUF_X2 U13421 ( .I(n35805), .Z(n61458) );
  INV_X1 U48163 ( .I(n34713), .ZN(n34321) );
  CLKBUF_X2 U10365 ( .I(n18884), .Z(n7183) );
  INV_X1 U18681 ( .I(n34150), .ZN(n33670) );
  INV_X2 U4992 ( .I(n23119), .ZN(n34626) );
  INV_X1 U11696 ( .I(n32454), .ZN(n32457) );
  INV_X2 U2713 ( .I(n34088), .ZN(n12039) );
  BUF_X2 U8073 ( .I(n35747), .Z(n60819) );
  INV_X2 U2547 ( .I(n33953), .ZN(n14980) );
  INV_X2 U18619 ( .I(n476), .ZN(n11247) );
  CLKBUF_X4 U11675 ( .I(n34972), .Z(n13818) );
  NOR2_X1 U9255 ( .A1(n7321), .A2(n23179), .ZN(n33824) );
  INV_X1 U18667 ( .I(n35309), .ZN(n3489) );
  INV_X1 U32877 ( .I(n34134), .ZN(n59483) );
  NAND2_X1 U13570 ( .A1(n14247), .A2(n2207), .ZN(n2206) );
  INV_X2 U28032 ( .I(n58702), .ZN(n34595) );
  NAND2_X1 U8058 ( .A1(n15085), .A2(n21008), .ZN(n2333) );
  CLKBUF_X1 U6132 ( .I(n33513), .Z(n58076) );
  INV_X2 U2616 ( .I(n11992), .ZN(n20279) );
  INV_X2 U9377 ( .I(n34201), .ZN(n19823) );
  INV_X2 U27045 ( .I(n15298), .ZN(n8780) );
  OR2_X1 U18480 ( .A1(n32976), .A2(n13352), .Z(n33766) );
  NAND2_X1 U47585 ( .A1(n32914), .A2(n7883), .ZN(n34526) );
  INV_X2 U13677 ( .I(n34661), .ZN(n1534) );
  CLKBUF_X4 U9369 ( .I(n17420), .Z(n59522) );
  NOR2_X1 U21777 ( .A1(n32700), .A2(n32699), .ZN(n33385) );
  NAND2_X1 U47822 ( .A1(n33354), .A2(n65052), .ZN(n33355) );
  NAND2_X1 U8255 ( .A1(n25625), .A2(n10358), .ZN(n33434) );
  INV_X1 U18500 ( .I(n33435), .ZN(n11396) );
  NAND2_X1 U11617 ( .A1(n60684), .A2(n10562), .ZN(n12877) );
  AOI21_X1 U37144 ( .A1(n33447), .A2(n34014), .B(n24296), .ZN(n24295) );
  OAI21_X1 U33408 ( .A1(n35196), .A2(n35702), .B(n60527), .ZN(n13610) );
  NAND2_X1 U22145 ( .A1(n33964), .A2(n3560), .ZN(n34090) );
  OR2_X1 U23290 ( .A1(n33350), .A2(n16939), .Z(n33105) );
  NAND3_X1 U8013 ( .A1(n22063), .A2(n34680), .A3(n34679), .ZN(n60059) );
  NAND2_X1 U15418 ( .A1(n34312), .A2(n57619), .ZN(n57618) );
  INV_X1 U46236 ( .I(n31298), .ZN(n31296) );
  INV_X2 U6732 ( .I(n61262), .ZN(n34796) );
  NAND3_X2 U3386 ( .A1(n19246), .A2(n11247), .A3(n34962), .ZN(n34537) );
  INV_X1 U11631 ( .I(n25634), .ZN(n34086) );
  NAND2_X1 U18319 ( .A1(n34135), .A2(n6923), .ZN(n6922) );
  OAI21_X1 U38163 ( .A1(n18393), .A2(n35319), .B(n16906), .ZN(n59968) );
  OAI21_X1 U43857 ( .A1(n60686), .A2(n19823), .B(n33989), .ZN(n60685) );
  NOR2_X1 U40206 ( .A1(n33955), .A2(n33954), .ZN(n20066) );
  OR2_X1 U13220 ( .A1(n21848), .A2(n35297), .Z(n57413) );
  NAND2_X1 U18311 ( .A1(n33424), .A2(n14285), .ZN(n21110) );
  NOR3_X1 U9554 ( .A1(n19823), .A2(n32890), .A3(n34200), .ZN(n2398) );
  OAI21_X1 U4922 ( .A1(n33692), .A2(n33691), .B(n10267), .ZN(n33708) );
  AOI22_X1 U47932 ( .A1(n63103), .A2(n33631), .B1(n33630), .B2(n33629), .ZN(
        n33633) );
  OAI21_X1 U18411 ( .A1(n61915), .A2(n34785), .B(n62373), .ZN(n18507) );
  NAND3_X1 U18329 ( .A1(n4537), .A2(n35004), .A3(n35003), .ZN(n35007) );
  NAND3_X1 U18351 ( .A1(n33355), .A2(n33356), .A3(n64100), .ZN(n33361) );
  NAND3_X1 U18432 ( .A1(n18947), .A2(n35661), .A3(n35649), .ZN(n18946) );
  AOI21_X1 U22350 ( .A1(n58243), .A2(n33728), .B(n33726), .ZN(n33735) );
  NAND2_X1 U56003 ( .A1(n61349), .A2(n33632), .ZN(n5254) );
  NOR2_X1 U6244 ( .A1(n13501), .A2(n32363), .ZN(n13500) );
  NAND3_X1 U30115 ( .A1(n20769), .A2(n33632), .A3(n33633), .ZN(n33648) );
  NAND2_X1 U34238 ( .A1(n35623), .A2(n8977), .ZN(n61359) );
  OR2_X1 U30027 ( .A1(n32142), .A2(n32140), .Z(n12302) );
  NAND2_X1 U52724 ( .A1(n61111), .A2(n34284), .ZN(n13129) );
  NOR2_X1 U18262 ( .A1(n21610), .A2(n14231), .ZN(n14084) );
  OAI22_X1 U9590 ( .A1(n34499), .A2(n34640), .B1(n34498), .B2(n61452), .ZN(
        n5130) );
  NOR2_X1 U18234 ( .A1(n9515), .A2(n2420), .ZN(n2419) );
  NOR2_X1 U18138 ( .A1(n5255), .A2(n5254), .ZN(n5253) );
  CLKBUF_X2 U30928 ( .I(n17202), .Z(n10485) );
  NAND2_X1 U18227 ( .A1(n16729), .A2(n16728), .ZN(n34453) );
  NOR2_X1 U30684 ( .A1(n3860), .A2(n59442), .ZN(n59181) );
  OAI21_X1 U18183 ( .A1(n32211), .A2(n26232), .B(n32210), .ZN(n32216) );
  CLKBUF_X4 U18113 ( .I(n36953), .Z(n22993) );
  INV_X1 U18170 ( .I(n36579), .ZN(n2116) );
  CLKBUF_X8 U5167 ( .I(n25677), .Z(n21605) );
  CLKBUF_X4 U9609 ( .I(n36233), .Z(n24028) );
  CLKBUF_X4 U7608 ( .I(n26147), .Z(n3622) );
  AND2_X1 U33029 ( .A1(n61940), .A2(n60562), .Z(n35165) );
  CLKBUF_X8 U6855 ( .I(n25611), .Z(n4541) );
  BUF_X2 U3177 ( .I(n15742), .Z(n61517) );
  CLKBUF_X4 U2474 ( .I(n21104), .Z(n5873) );
  BUF_X4 U18152 ( .I(n36030), .Z(n1787) );
  INV_X1 U34921 ( .I(n36943), .ZN(n34903) );
  CLKBUF_X4 U3183 ( .I(n36717), .Z(n20867) );
  INV_X2 U2436 ( .I(n19278), .ZN(n37426) );
  CLKBUF_X4 U2402 ( .I(n19278), .Z(n22595) );
  CLKBUF_X8 U8394 ( .I(n7693), .Z(n1235) );
  CLKBUF_X4 U4015 ( .I(n1422), .Z(n60925) );
  INV_X1 U4808 ( .I(n37136), .ZN(n17492) );
  INV_X1 U9921 ( .I(n34372), .ZN(n36161) );
  NAND2_X1 U18092 ( .A1(n36808), .A2(n36075), .ZN(n35397) );
  INV_X2 U25423 ( .I(n8039), .ZN(n5734) );
  INV_X1 U17823 ( .I(n37091), .ZN(n37017) );
  INV_X1 U31050 ( .I(n15442), .ZN(n36640) );
  AOI21_X1 U47815 ( .A1(n37365), .A2(n2594), .B(n37364), .ZN(n33329) );
  INV_X1 U48502 ( .I(n35444), .ZN(n35446) );
  AOI21_X1 U48702 ( .A1(n36153), .A2(n36152), .B(n36583), .ZN(n36156) );
  INV_X1 U48905 ( .I(n36804), .ZN(n36806) );
  NAND2_X1 U10223 ( .A1(n64423), .A2(n35174), .ZN(n35563) );
  OR2_X1 U9853 ( .A1(n34821), .A2(n34820), .Z(n16058) );
  INV_X1 U6063 ( .I(n35995), .ZN(n58074) );
  NOR3_X1 U13339 ( .A1(n36223), .A2(n36221), .A3(n57171), .ZN(n7644) );
  INV_X1 U17984 ( .I(n17851), .ZN(n2117) );
  INV_X1 U35729 ( .I(n36515), .ZN(n36518) );
  INV_X1 U17978 ( .I(n36001), .ZN(n31305) );
  OAI21_X1 U48066 ( .A1(n20251), .A2(n33931), .B(n35087), .ZN(n33932) );
  INV_X1 U17916 ( .I(n7245), .ZN(n7244) );
  AOI21_X1 U48763 ( .A1(n36340), .A2(n58769), .B(n36339), .ZN(n36341) );
  NAND2_X1 U13256 ( .A1(n36872), .A2(n35335), .ZN(n36694) );
  OAI21_X1 U10225 ( .A1(n35464), .A2(n20712), .B(n35463), .ZN(n35466) );
  OR2_X1 U27407 ( .A1(n35487), .A2(n35911), .Z(n7434) );
  AOI21_X1 U2262 ( .A1(n35418), .A2(n34007), .B(n34369), .ZN(n35420) );
  AOI21_X1 U32245 ( .A1(n34110), .A2(n12116), .B(n19231), .ZN(n24630) );
  OAI22_X1 U32957 ( .A1(n34096), .A2(n36584), .B1(n63247), .B2(n12967), .ZN(
        n25752) );
  AOI21_X1 U17792 ( .A1(n37047), .A2(n63469), .B(n37045), .ZN(n37058) );
  NAND2_X1 U29910 ( .A1(n59122), .A2(n37369), .ZN(n59058) );
  NAND2_X1 U7735 ( .A1(n24341), .A2(n34832), .ZN(n20521) );
  NAND2_X1 U17723 ( .A1(n36455), .A2(n36456), .ZN(n14398) );
  INV_X1 U17899 ( .I(n36705), .ZN(n12763) );
  NOR2_X1 U7772 ( .A1(n15082), .A2(n12358), .ZN(n12357) );
  INV_X1 U48940 ( .I(n37434), .ZN(n36917) );
  NAND2_X1 U15367 ( .A1(n11779), .A2(n11561), .ZN(n57607) );
  OAI22_X1 U13252 ( .A1(n37104), .A2(n37356), .B1(n6389), .B2(n2279), .ZN(
        n17912) );
  AND2_X2 U13237 ( .A1(n14895), .A2(n11304), .Z(n14891) );
  AOI22_X1 U17690 ( .A1(n15010), .A2(n15009), .B1(n20956), .B2(n7244), .ZN(
        n25688) );
  NAND3_X1 U17782 ( .A1(n14686), .A2(n36433), .A3(n14685), .ZN(n14684) );
  INV_X1 U7836 ( .I(n36822), .ZN(n35916) );
  NAND2_X1 U38986 ( .A1(n60085), .A2(n60084), .ZN(n61289) );
  NAND3_X1 U48740 ( .A1(n36957), .A2(n36274), .A3(n36273), .ZN(n36277) );
  NAND2_X1 U48742 ( .A1(n36277), .A2(n36276), .ZN(n36285) );
  NOR2_X1 U9929 ( .A1(n36682), .A2(n36681), .ZN(n36683) );
  NOR3_X1 U7734 ( .A1(n59037), .A2(n7821), .A3(n36556), .ZN(n4817) );
  NAND2_X1 U30452 ( .A1(n36458), .A2(n14398), .ZN(n59642) );
  NAND3_X1 U23602 ( .A1(n5152), .A2(n11466), .A3(n37965), .ZN(n58416) );
  NOR2_X1 U22817 ( .A1(n59337), .A2(n20680), .ZN(n58304) );
  OAI21_X1 U35288 ( .A1(n37020), .A2(n37021), .B(n20419), .ZN(n20418) );
  AOI21_X1 U40809 ( .A1(n33410), .A2(n33411), .B(n24629), .ZN(n24628) );
  OAI21_X1 U11436 ( .A1(n33527), .A2(n7933), .B(n2299), .ZN(n2298) );
  NAND2_X1 U10213 ( .A1(n19608), .A2(n19607), .ZN(n9579) );
  CLKBUF_X4 U3566 ( .I(n24151), .Z(n11142) );
  CLKBUF_X4 U17667 ( .I(n38535), .Z(n10017) );
  CLKBUF_X4 U17676 ( .I(n39769), .Z(n23019) );
  CLKBUF_X4 U13208 ( .I(n14798), .Z(n5555) );
  NAND2_X1 U4542 ( .A1(n36683), .A2(n30), .ZN(n24382) );
  INV_X1 U13211 ( .I(n23637), .ZN(n18354) );
  INV_X2 U29578 ( .I(n466), .ZN(n18831) );
  CLKBUF_X4 U2652 ( .I(n38856), .Z(n19303) );
  CLKBUF_X2 U17584 ( .I(n22277), .Z(n7713) );
  NOR2_X1 U50627 ( .A1(n24382), .A2(n24381), .ZN(n19184) );
  CLKBUF_X4 U4300 ( .I(n39254), .Z(n16594) );
  CLKBUF_X2 U11381 ( .I(n23949), .Z(n2334) );
  BUF_X2 U17579 ( .I(n39687), .Z(n22855) );
  BUF_X4 U17568 ( .I(n39346), .Z(n23927) );
  BUF_X2 U7720 ( .I(n39186), .Z(n61489) );
  CLKBUF_X2 U8209 ( .I(n39543), .Z(n23655) );
  CLKBUF_X4 U27640 ( .I(n11829), .Z(n7573) );
  CLKBUF_X4 U4445 ( .I(n38537), .Z(n233) );
  CLKBUF_X2 U17561 ( .I(n38729), .Z(n21009) );
  INV_X1 U10033 ( .I(n3479), .ZN(n21560) );
  NAND2_X1 U13183 ( .A1(n12267), .A2(n1763), .ZN(n7958) );
  CLKBUF_X2 U10069 ( .I(n25998), .Z(n58587) );
  CLKBUF_X4 U6014 ( .I(n36105), .Z(n41034) );
  BUF_X2 U8763 ( .I(n40961), .Z(n23787) );
  INV_X2 U22110 ( .I(n1239), .ZN(n8539) );
  CLKBUF_X2 U11358 ( .I(n39604), .Z(n40697) );
  BUF_X2 U25177 ( .I(n9606), .Z(n5488) );
  INV_X1 U2077 ( .I(n11188), .ZN(n22564) );
  INV_X2 U2473 ( .I(n15934), .ZN(n41875) );
  CLKBUF_X2 U17485 ( .I(n15930), .Z(n23319) );
  CLKBUF_X4 U26941 ( .I(n41474), .Z(n7165) );
  CLKBUF_X4 U7622 ( .I(n15934), .Z(n59583) );
  CLKBUF_X4 U17483 ( .I(n38922), .Z(n1743) );
  CLKBUF_X2 U37635 ( .I(n38924), .Z(n41212) );
  CLKBUF_X2 U34878 ( .I(n39317), .Z(n40026) );
  CLKBUF_X2 U10085 ( .I(n23720), .Z(n21057) );
  INV_X1 U30975 ( .I(n22564), .ZN(n39147) );
  INV_X2 U33824 ( .I(n42200), .ZN(n14280) );
  INV_X2 U38753 ( .I(n41162), .ZN(n41164) );
  CLKBUF_X4 U8750 ( .I(n38291), .Z(n40063) );
  CLKBUF_X2 U8751 ( .I(n38493), .Z(n40664) );
  CLKBUF_X4 U43587 ( .I(n40697), .Z(n60653) );
  CLKBUF_X4 U17463 ( .I(n42284), .Z(n21492) );
  INV_X1 U2067 ( .I(n20348), .ZN(n20339) );
  CLKBUF_X2 U6015 ( .I(n10044), .Z(n59531) );
  INV_X2 U13171 ( .I(n19638), .ZN(n19331) );
  BUF_X2 U4079 ( .I(n38336), .Z(n40308) );
  CLKBUF_X4 U1975 ( .I(n40850), .Z(n18741) );
  CLKBUF_X4 U3528 ( .I(n38600), .Z(n40968) );
  INV_X1 U10088 ( .I(n41445), .ZN(n25430) );
  INV_X2 U38165 ( .I(n18242), .ZN(n17945) );
  INV_X1 U28545 ( .I(n10669), .ZN(n60509) );
  BUF_X2 U1948 ( .I(n42508), .Z(n9954) );
  BUF_X2 U10304 ( .I(n36648), .Z(n2159) );
  INV_X2 U3586 ( .I(n41078), .ZN(n3345) );
  NOR2_X1 U51357 ( .A1(n42479), .A2(n42480), .ZN(n42478) );
  BUF_X2 U2567 ( .I(n22525), .Z(n61316) );
  AOI21_X1 U26776 ( .A1(n971), .A2(n40444), .B(n19343), .ZN(n40446) );
  INV_X2 U24458 ( .I(n42450), .ZN(n41810) );
  CLKBUF_X2 U12877 ( .I(n15503), .Z(n9725) );
  NOR2_X1 U30813 ( .A1(n40194), .A2(n59427), .ZN(n59211) );
  INV_X2 U2310 ( .I(n22168), .ZN(n66) );
  CLKBUF_X2 U33686 ( .I(n42226), .Z(n59577) );
  NAND2_X1 U50011 ( .A1(n38765), .A2(n38763), .ZN(n38764) );
  INV_X1 U11287 ( .I(n38765), .ZN(n40761) );
  BUF_X2 U10155 ( .I(n11765), .Z(n10593) );
  NAND2_X1 U29046 ( .A1(n21255), .A2(n59199), .ZN(n40236) );
  OAI21_X1 U29795 ( .A1(n40678), .A2(n40677), .B(n40676), .ZN(n59034) );
  INV_X1 U10076 ( .I(n40967), .ZN(n38543) );
  NAND2_X1 U17155 ( .A1(n40764), .A2(n58047), .ZN(n18667) );
  INV_X1 U8710 ( .I(n38420), .ZN(n40612) );
  OR2_X1 U13471 ( .A1(n25424), .A2(n10452), .Z(n57451) );
  INV_X1 U17146 ( .I(n40702), .ZN(n17831) );
  OAI21_X1 U41609 ( .A1(n10500), .A2(n5506), .B(n5505), .ZN(n60401) );
  OR3_X1 U23210 ( .A1(n42228), .A2(n22290), .A3(n41949), .Z(n17073) );
  INV_X2 U1910 ( .I(n18856), .ZN(n1303) );
  NOR2_X1 U8738 ( .A1(n61785), .A2(n64895), .ZN(n13034) );
  INV_X1 U1853 ( .I(n10500), .ZN(n41899) );
  INV_X2 U8103 ( .I(n61708), .ZN(n41844) );
  NAND2_X1 U36738 ( .A1(n16680), .A2(n10481), .ZN(n17981) );
  NAND2_X1 U32713 ( .A1(n59455), .A2(n17581), .ZN(n17580) );
  NAND2_X1 U29791 ( .A1(n40680), .A2(n59034), .ZN(n40682) );
  OAI21_X1 U51224 ( .A1(n41943), .A2(n20190), .B(n41942), .ZN(n41946) );
  CLKBUF_X2 U30673 ( .I(n40491), .Z(n59179) );
  INV_X2 U36989 ( .I(n60612), .ZN(n41924) );
  NAND2_X1 U50481 ( .A1(n40003), .A2(n61638), .ZN(n39699) );
  NAND2_X1 U17129 ( .A1(n6752), .A2(n6751), .ZN(n6582) );
  OAI21_X1 U12975 ( .A1(n15776), .A2(n42214), .B(n42213), .ZN(n42219) );
  NOR2_X1 U5942 ( .A1(n40165), .A2(n40158), .ZN(n61626) );
  NOR2_X1 U5938 ( .A1(n13724), .A2(n1403), .ZN(n59266) );
  INV_X1 U7474 ( .I(n38194), .ZN(n60123) );
  NAND2_X1 U13075 ( .A1(n15679), .A2(n15680), .ZN(n12101) );
  NOR2_X1 U10305 ( .A1(n42208), .A2(n20669), .ZN(n42221) );
  AND4_X2 U21638 ( .A1(n3135), .A2(n3134), .A3(n5395), .A4(n5391), .Z(n3133)
         );
  AOI22_X1 U17318 ( .A1(n40264), .A2(n40939), .B1(n40477), .B2(n3306), .ZN(
        n40265) );
  OAI21_X1 U50780 ( .A1(n60229), .A2(n40930), .B(n40468), .ZN(n40478) );
  NAND2_X1 U16960 ( .A1(n38846), .A2(n38845), .ZN(n20474) );
  NAND2_X1 U50645 ( .A1(n40244), .A2(n60113), .ZN(n40080) );
  NAND2_X1 U17131 ( .A1(n15427), .A2(n15426), .ZN(n15428) );
  NAND2_X1 U4369 ( .A1(n41172), .A2(n40487), .ZN(n701) );
  OAI21_X1 U3688 ( .A1(n15541), .A2(n15542), .B(n41813), .ZN(n1932) );
  AOI21_X1 U17276 ( .A1(n38479), .A2(n59179), .B(n5707), .ZN(n5706) );
  OAI21_X1 U52959 ( .A1(n39699), .A2(n39700), .B(n57257), .ZN(n61124) );
  NAND2_X1 U8699 ( .A1(n41842), .A2(n16643), .ZN(n41847) );
  NAND2_X1 U27401 ( .A1(n41903), .A2(n41902), .ZN(n41911) );
  AOI21_X1 U13031 ( .A1(n24950), .A2(n40642), .B(n22007), .ZN(n22006) );
  NAND2_X1 U13047 ( .A1(n41231), .A2(n41397), .ZN(n8919) );
  OAI21_X1 U20033 ( .A1(n40274), .A2(n16970), .B(n38020), .ZN(n59143) );
  NOR2_X1 U24651 ( .A1(n59855), .A2(n7188), .ZN(n58578) );
  AOI21_X1 U11246 ( .A1(n7681), .A2(n41308), .B(n61916), .ZN(n3495) );
  NOR3_X1 U25533 ( .A1(n17296), .A2(n16289), .A3(n17295), .ZN(n5869) );
  NOR2_X1 U16978 ( .A1(n13000), .A2(n12998), .ZN(n17029) );
  AOI21_X1 U24535 ( .A1(n39119), .A2(n25201), .B(n58565), .ZN(n58564) );
  CLKBUF_X4 U4950 ( .I(n24294), .Z(n2995) );
  NAND3_X1 U34634 ( .A1(n59692), .A2(n40497), .A3(n40495), .ZN(n40498) );
  NOR2_X1 U7390 ( .A1(n61292), .A2(n61290), .ZN(n16392) );
  NAND2_X1 U32801 ( .A1(n42238), .A2(n12730), .ZN(n43717) );
  CLKBUF_X4 U4900 ( .I(n42175), .Z(n3618) );
  INV_X4 U1734 ( .I(n42347), .ZN(n1502) );
  CLKBUF_X2 U34541 ( .I(n43549), .Z(n59682) );
  CLKBUF_X4 U10060 ( .I(n13493), .Z(n11727) );
  OAI21_X1 U10082 ( .A1(n8442), .A2(n8441), .B(n8439), .ZN(n13797) );
  NOR2_X1 U12960 ( .A1(n40822), .A2(n40821), .ZN(n40823) );
  CLKBUF_X1 U12943 ( .I(n19946), .Z(n4714) );
  CLKBUF_X4 U30827 ( .I(n42914), .Z(n10415) );
  CLKBUF_X4 U16967 ( .I(n44227), .Z(n22716) );
  INV_X1 U4020 ( .I(n43376), .ZN(n41571) );
  INV_X4 U53854 ( .I(n61739), .ZN(n61186) );
  CLKBUF_X2 U5906 ( .I(n43464), .Z(n58530) );
  CLKBUF_X4 U16834 ( .I(n20351), .Z(n23488) );
  BUF_X4 U5059 ( .I(n21667), .Z(n15020) );
  BUF_X4 U30054 ( .I(n42662), .Z(n9914) );
  NOR2_X1 U16573 ( .A1(n38685), .A2(n42922), .ZN(n42113) );
  INV_X1 U9303 ( .I(n14659), .ZN(n42805) );
  NOR2_X1 U16646 ( .A1(n9511), .A2(n16527), .ZN(n20235) );
  NOR2_X1 U35976 ( .A1(n43447), .A2(n43449), .ZN(n18796) );
  CLKBUF_X4 U39386 ( .I(n8911), .Z(n60131) );
  NAND2_X1 U51380 ( .A1(n42915), .A2(n42552), .ZN(n42556) );
  AOI21_X1 U12836 ( .A1(n43028), .A2(n43024), .B(n41665), .ZN(n10298) );
  NOR2_X1 U3455 ( .A1(n43633), .A2(n42098), .ZN(n17244) );
  NAND2_X1 U1974 ( .A1(n42776), .A2(n43024), .ZN(n58574) );
  CLKBUF_X2 U16757 ( .I(n46331), .Z(n10487) );
  NOR2_X1 U36994 ( .A1(n3652), .A2(n38686), .ZN(n23635) );
  NOR2_X1 U16657 ( .A1(n43959), .A2(n14408), .ZN(n14407) );
  NOR2_X1 U24852 ( .A1(n42113), .A2(n58613), .ZN(n58612) );
  INV_X1 U11101 ( .I(n43677), .ZN(n21519) );
  INV_X1 U50184 ( .I(n39086), .ZN(n40914) );
  AOI21_X1 U32264 ( .A1(n13547), .A2(n12154), .B(n42716), .ZN(n42723) );
  INV_X1 U7087 ( .I(n42419), .ZN(n43475) );
  INV_X1 U4899 ( .I(n42398), .ZN(n1688) );
  NAND2_X1 U16510 ( .A1(n42767), .A2(n42801), .ZN(n13123) );
  NAND2_X1 U56112 ( .A1(n42825), .A2(n42835), .ZN(n61356) );
  NAND2_X1 U5848 ( .A1(n58574), .A2(n42786), .ZN(n5906) );
  AOI21_X1 U16547 ( .A1(n24494), .A2(n41762), .B(n41765), .ZN(n23107) );
  NAND2_X1 U12902 ( .A1(n42667), .A2(n41560), .ZN(n22500) );
  NAND2_X1 U16529 ( .A1(n12972), .A2(n8171), .ZN(n24130) );
  AOI22_X1 U22563 ( .A1(n58274), .A2(n37919), .B1(n37920), .B2(n42018), .ZN(
        n37921) );
  INV_X1 U31967 ( .I(n59356), .ZN(n43363) );
  INV_X2 U25458 ( .I(n25327), .ZN(n42338) );
  OR2_X1 U7142 ( .A1(n42405), .A2(n42397), .Z(n60243) );
  NOR2_X1 U36922 ( .A1(n43451), .A2(n43450), .ZN(n25119) );
  INV_X1 U10527 ( .I(n41550), .ZN(n13453) );
  OAI21_X1 U16500 ( .A1(n6396), .A2(n5827), .B(n43352), .ZN(n5826) );
  INV_X1 U16739 ( .I(n19346), .ZN(n43311) );
  INV_X1 U12851 ( .I(n43271), .ZN(n3730) );
  AOI21_X1 U35488 ( .A1(n41710), .A2(n21934), .B(n21933), .ZN(n41712) );
  INV_X1 U36083 ( .I(n43237), .ZN(n43235) );
  NOR2_X1 U16641 ( .A1(n43363), .A2(n42732), .ZN(n42733) );
  NOR2_X1 U10568 ( .A1(n1193), .A2(n16480), .ZN(n42066) );
  NOR3_X1 U30618 ( .A1(n19939), .A2(n43609), .A3(n43610), .ZN(n10258) );
  INV_X1 U16612 ( .I(n13882), .ZN(n41637) );
  NAND2_X1 U1821 ( .A1(n43236), .A2(n43237), .ZN(n59672) );
  NAND2_X1 U7079 ( .A1(n5906), .A2(n57196), .ZN(n59767) );
  NAND2_X1 U36879 ( .A1(n41680), .A2(n41999), .ZN(n17859) );
  NAND2_X1 U12799 ( .A1(n14754), .A2(n42319), .ZN(n23427) );
  NAND3_X1 U25583 ( .A1(n43932), .A2(n43931), .A3(n43930), .ZN(n44912) );
  NAND3_X1 U21258 ( .A1(n19336), .A2(n9713), .A3(n2884), .ZN(n21681) );
  NAND2_X1 U36979 ( .A1(n42824), .A2(n41246), .ZN(n41247) );
  NOR2_X1 U51605 ( .A1(n43456), .A2(n43455), .ZN(n43482) );
  NOR3_X1 U24127 ( .A1(n25579), .A2(n25578), .A3(n57431), .ZN(n25576) );
  NAND4_X1 U5732 ( .A1(n42884), .A2(n42882), .A3(n42883), .A4(n42885), .ZN(
        n25009) );
  NAND2_X1 U12797 ( .A1(n9366), .A2(n24087), .ZN(n24085) );
  AOI21_X1 U26904 ( .A1(n41366), .A2(n41365), .B(n41364), .ZN(n41374) );
  NOR2_X1 U50861 ( .A1(n61285), .A2(n9247), .ZN(n61284) );
  NOR2_X1 U12764 ( .A1(n16341), .A2(n16340), .ZN(n16339) );
  CLKBUF_X4 U13545 ( .I(n46321), .Z(n3104) );
  NOR2_X1 U51486 ( .A1(n44234), .A2(n44232), .ZN(n42960) );
  CLKBUF_X4 U16433 ( .I(n22973), .Z(n7424) );
  NAND3_X1 U16438 ( .A1(n42996), .A2(n41358), .A3(n41357), .ZN(n41359) );
  NAND2_X1 U42964 ( .A1(n43389), .A2(n24129), .ZN(n46538) );
  CLKBUF_X2 U12740 ( .I(n45019), .Z(n23078) );
  CLKBUF_X4 U12730 ( .I(n17984), .Z(n17983) );
  INV_X2 U51754 ( .I(n65177), .ZN(n44608) );
  CLKBUF_X4 U1402 ( .I(n46283), .Z(n23687) );
  BUF_X2 U10885 ( .I(n44834), .Z(n58027) );
  INV_X2 U3623 ( .I(n14760), .ZN(n18331) );
  INV_X2 U37724 ( .I(n58027), .ZN(n45261) );
  CLKBUF_X4 U10882 ( .I(n14752), .Z(n12377) );
  CLKBUF_X4 U57170 ( .I(n46233), .Z(n11317) );
  INV_X2 U12727 ( .I(n22551), .ZN(n3339) );
  CLKBUF_X2 U12720 ( .I(n11555), .Z(n11554) );
  CLKBUF_X2 U6922 ( .I(n14055), .Z(n60350) );
  CLKBUF_X2 U7800 ( .I(n19483), .Z(n13746) );
  CLKBUF_X4 U26925 ( .I(n44064), .Z(n46985) );
  OR2_X2 U1444 ( .A1(n13298), .A2(n17891), .Z(n46771) );
  CLKBUF_X2 U5778 ( .I(n11150), .Z(n60979) );
  CLKBUF_X2 U9282 ( .I(n44670), .Z(n21044) );
  CLKBUF_X4 U29965 ( .I(n45218), .Z(n9860) );
  CLKBUF_X2 U7826 ( .I(n16993), .Z(n10428) );
  CLKBUF_X4 U29588 ( .I(n47748), .Z(n59008) );
  CLKBUF_X2 U6856 ( .I(n48564), .Z(n697) );
  INV_X2 U1271 ( .I(n25340), .ZN(n22736) );
  INV_X1 U1290 ( .I(n16783), .ZN(n48244) );
  BUF_X2 U6895 ( .I(n47541), .Z(n58675) );
  INV_X2 U26462 ( .I(n46959), .ZN(n46951) );
  BUF_X2 U16285 ( .I(n61714), .Z(n22391) );
  CLKBUF_X2 U42401 ( .I(n23588), .Z(n60504) );
  INV_X1 U53285 ( .I(n8012), .ZN(n48605) );
  CLKBUF_X2 U12705 ( .I(n16836), .Z(n23661) );
  INV_X2 U38838 ( .I(n17967), .ZN(n45905) );
  CLKBUF_X2 U47324 ( .I(n47127), .Z(n60848) );
  BUF_X2 U6896 ( .I(n47467), .Z(n58174) );
  CLKBUF_X4 U1425 ( .I(n61961), .Z(n59629) );
  INV_X2 U4399 ( .I(n6730), .ZN(n45901) );
  INV_X1 U5877 ( .I(n47020), .ZN(n20238) );
  CLKBUF_X4 U18271 ( .I(n26145), .Z(n20162) );
  NAND2_X1 U16144 ( .A1(n10624), .A2(n48561), .ZN(n46782) );
  INV_X2 U11049 ( .I(n47465), .ZN(n46977) );
  INV_X1 U53164 ( .I(n47096), .ZN(n47099) );
  NOR2_X1 U37362 ( .A1(n60398), .A2(n60358), .ZN(n47210) );
  INV_X2 U16214 ( .I(n46817), .ZN(n48096) );
  NOR2_X1 U1481 ( .A1(n13655), .A2(n61563), .ZN(n16074) );
  INV_X2 U11187 ( .I(n18127), .ZN(n22389) );
  INV_X1 U16078 ( .I(n47885), .ZN(n47714) );
  INV_X2 U23016 ( .I(n4678), .ZN(n46958) );
  NAND2_X1 U1195 ( .A1(n20238), .A2(n19595), .ZN(n47022) );
  CLKBUF_X2 U11202 ( .I(n4678), .Z(n60727) );
  NAND2_X1 U52577 ( .A1(n45953), .A2(n63700), .ZN(n45629) );
  AOI21_X1 U12603 ( .A1(n20574), .A2(n16012), .B(n21198), .ZN(n20576) );
  NAND2_X1 U1079 ( .A1(n46911), .A2(n44201), .ZN(n44204) );
  INV_X1 U29788 ( .I(n46022), .ZN(n46012) );
  NAND2_X1 U15881 ( .A1(n48486), .A2(n48485), .ZN(n8025) );
  CLKBUF_X2 U5698 ( .I(n22684), .Z(n61212) );
  NOR2_X1 U12576 ( .A1(n47702), .A2(n47701), .ZN(n47711) );
  NAND2_X1 U52138 ( .A1(n44683), .A2(n44682), .ZN(n44688) );
  OAI22_X1 U15052 ( .A1(n48498), .A2(n48497), .B1(n48496), .B2(n48648), .ZN(
        n57570) );
  NAND2_X1 U15910 ( .A1(n47906), .A2(n47571), .ZN(n4353) );
  INV_X1 U1125 ( .I(n45565), .ZN(n17572) );
  NAND2_X1 U22269 ( .A1(n1661), .A2(n47295), .ZN(n3640) );
  OAI22_X1 U52923 ( .A1(n46465), .A2(n46464), .B1(n46463), .B2(n46462), .ZN(
        n46467) );
  INV_X1 U52624 ( .I(n45710), .ZN(n45711) );
  OAI21_X1 U11212 ( .A1(n22011), .A2(n22012), .B(n45975), .ZN(n22010) );
  AOI22_X1 U52609 ( .A1(n45679), .A2(n45678), .B1(n47277), .B2(n45677), .ZN(
        n45687) );
  AND3_X1 U42055 ( .A1(n47313), .A2(n47312), .A3(n47311), .Z(n23409) );
  NAND2_X1 U11090 ( .A1(n22872), .A2(n45529), .ZN(n10375) );
  NAND2_X1 U53376 ( .A1(n47814), .A2(n1481), .ZN(n47815) );
  OAI21_X1 U36121 ( .A1(n22871), .A2(n22872), .B(n20938), .ZN(n18318) );
  NOR2_X1 U15738 ( .A1(n47021), .A2(n44576), .ZN(n18324) );
  INV_X1 U15993 ( .I(n45630), .ZN(n45632) );
  NAND3_X1 U21909 ( .A1(n44286), .A2(n44285), .A3(n57262), .ZN(n60308) );
  NOR2_X1 U12524 ( .A1(n22872), .A2(n45540), .ZN(n45541) );
  NOR2_X1 U12539 ( .A1(n12824), .A2(n45483), .ZN(n11294) );
  NAND2_X1 U12607 ( .A1(n47362), .A2(n8953), .ZN(n45182) );
  NOR2_X1 U5677 ( .A1(n47116), .A2(n48094), .ZN(n59471) );
  NAND2_X1 U43411 ( .A1(n60637), .A2(n45647), .ZN(n45606) );
  AOI21_X1 U51998 ( .A1(n44404), .A2(n44403), .B(n44402), .ZN(n44405) );
  INV_X1 U16150 ( .I(n47875), .ZN(n11907) );
  NAND2_X1 U1042 ( .A1(n17746), .A2(n23048), .ZN(n4095) );
  NOR2_X1 U15782 ( .A1(n44688), .A2(n44687), .ZN(n44689) );
  NOR2_X1 U29798 ( .A1(n14623), .A2(n1098), .ZN(n59035) );
  NOR2_X1 U53137 ( .A1(n61139), .A2(n61138), .ZN(n15781) );
  NAND2_X1 U15719 ( .A1(n16879), .A2(n17032), .ZN(n16878) );
  CLKBUF_X4 U6785 ( .I(n50422), .Z(n23063) );
  CLKBUF_X4 U34376 ( .I(n1110), .Z(n15021) );
  NAND2_X1 U28282 ( .A1(n58883), .A2(n45944), .ZN(n23104) );
  CLKBUF_X4 U26691 ( .I(n50054), .Z(n3054) );
  CLKBUF_X4 U42916 ( .I(n48338), .Z(n24069) );
  OAI21_X1 U52787 ( .A1(n47018), .A2(n48603), .B(n47525), .ZN(n46098) );
  CLKBUF_X2 U5639 ( .I(n49701), .Z(n22646) );
  CLKBUF_X1 U10874 ( .I(n11034), .Z(n10045) );
  CLKBUF_X4 U1035 ( .I(n5587), .Z(n4888) );
  INV_X2 U3493 ( .I(n50229), .ZN(n5258) );
  INV_X4 U30327 ( .I(n50346), .ZN(n21870) );
  CLKBUF_X4 U26303 ( .I(n49012), .Z(n6654) );
  CLKBUF_X4 U7886 ( .I(n10472), .Z(n4780) );
  INV_X1 U15611 ( .I(n47919), .ZN(n25967) );
  BUF_X2 U5595 ( .I(n49114), .Z(n59493) );
  CLKBUF_X4 U4465 ( .I(n48362), .Z(n22457) );
  INV_X1 U6645 ( .I(n10961), .ZN(n16197) );
  CLKBUF_X2 U5161 ( .I(n17379), .Z(n201) );
  CLKBUF_X4 U6659 ( .I(n49171), .Z(n58907) );
  INV_X1 U27404 ( .I(n7328), .ZN(n60648) );
  NAND2_X1 U25982 ( .A1(n6323), .A2(n1644), .ZN(n19714) );
  CLKBUF_X4 U5951 ( .I(n49637), .Z(n10958) );
  INV_X2 U27952 ( .I(n4173), .ZN(n58840) );
  INV_X1 U11421 ( .I(n48445), .ZN(n26069) );
  NOR2_X1 U8551 ( .A1(n63943), .A2(n19773), .ZN(n12616) );
  CLKBUF_X4 U1131 ( .I(n12646), .Z(n359) );
  NAND2_X1 U12417 ( .A1(n49138), .A2(n17200), .ZN(n49997) );
  INV_X1 U15533 ( .I(n49980), .ZN(n48167) );
  OR2_X2 U23524 ( .A1(n49500), .A2(n22780), .Z(n20363) );
  AOI21_X1 U53775 ( .A1(n22526), .A2(n3237), .B(n49153), .ZN(n49154) );
  INV_X1 U9205 ( .I(n22926), .ZN(n3032) );
  NAND2_X1 U41512 ( .A1(n22174), .A2(n49777), .ZN(n22173) );
  NAND2_X1 U15405 ( .A1(n50077), .A2(n15166), .ZN(n15165) );
  INV_X1 U9886 ( .I(n48690), .ZN(n49050) );
  OR2_X1 U756 ( .A1(n49731), .A2(n46728), .Z(n1095) );
  INV_X2 U1062 ( .I(n48745), .ZN(n50277) );
  OAI21_X1 U21835 ( .A1(n50241), .A2(n3281), .B(n50233), .ZN(n22198) );
  BUF_X2 U4766 ( .I(n48802), .Z(n59004) );
  CLKBUF_X4 U21906 ( .I(n9799), .Z(n3347) );
  OAI21_X1 U649 ( .A1(n47997), .A2(n47998), .B(n50221), .ZN(n47999) );
  INV_X1 U53434 ( .I(n48007), .ZN(n48008) );
  INV_X2 U30073 ( .I(n17818), .ZN(n9924) );
  AOI21_X1 U6686 ( .A1(n48168), .A2(n49972), .B(n48167), .ZN(n21466) );
  NOR2_X1 U3680 ( .A1(n9727), .A2(n48962), .ZN(n49270) );
  NAND2_X1 U5570 ( .A1(n60666), .A2(n18683), .ZN(n48851) );
  NAND2_X1 U30143 ( .A1(n59100), .A2(n14069), .ZN(n14067) );
  NAND2_X1 U5579 ( .A1(n58016), .A2(n17516), .ZN(n14068) );
  NOR2_X1 U15288 ( .A1(n15848), .A2(n25040), .ZN(n17707) );
  NOR2_X1 U15389 ( .A1(n49609), .A2(n64256), .ZN(n14127) );
  AOI22_X1 U53895 ( .A1(n49601), .A2(n49600), .B1(n49599), .B2(n23656), .ZN(
        n49603) );
  AOI21_X1 U53942 ( .A1(n49791), .A2(n49790), .B(n10015), .ZN(n49802) );
  AND3_X1 U10788 ( .A1(n49001), .A2(n24711), .A3(n24710), .Z(n25500) );
  NAND2_X1 U11650 ( .A1(n59310), .A2(n3241), .ZN(n3240) );
  NOR2_X1 U43920 ( .A1(n49157), .A2(n49156), .ZN(n49165) );
  NOR3_X1 U53886 ( .A1(n50047), .A2(n18565), .A3(n49580), .ZN(n49586) );
  OAI21_X1 U12366 ( .A1(n49192), .A2(n16484), .B(n18431), .ZN(n9234) );
  OAI21_X1 U11756 ( .A1(n12337), .A2(n49191), .B(n49516), .ZN(n12336) );
  NAND2_X1 U15198 ( .A1(n4012), .A2(n4011), .ZN(n4010) );
  OAI21_X1 U12375 ( .A1(n49409), .A2(n49408), .B(n2382), .ZN(n2381) );
  NAND2_X1 U28948 ( .A1(n8789), .A2(n65208), .ZN(n7782) );
  CLKBUF_X2 U42428 ( .I(n50796), .Z(n23344) );
  NAND2_X1 U31132 ( .A1(n12333), .A2(n49197), .ZN(n12332) );
  NOR2_X1 U15234 ( .A1(n47053), .A2(n47052), .ZN(n47056) );
  CLKBUF_X4 U15180 ( .I(n52424), .Z(n9635) );
  BUF_X2 U10779 ( .I(n9156), .Z(n9154) );
  CLKBUF_X2 U6523 ( .I(n8147), .Z(n3318) );
  INV_X2 U26038 ( .I(n22979), .ZN(n50792) );
  CLKBUF_X4 U13624 ( .I(n52409), .Z(n18645) );
  BUF_X4 U15148 ( .I(n50550), .Z(n52073) );
  INV_X1 U12324 ( .I(n23342), .ZN(n7340) );
  CLKBUF_X4 U6538 ( .I(n50797), .Z(n61423) );
  CLKBUF_X4 U25305 ( .I(n7111), .Z(n5626) );
  CLKBUF_X1 U15118 ( .I(n19189), .Z(n8180) );
  BUF_X2 U5560 ( .I(n23883), .Z(n61092) );
  INV_X1 U15081 ( .I(n52586), .ZN(n8615) );
  INV_X2 U501 ( .I(n51962), .ZN(n55299) );
  INV_X1 U15077 ( .I(n51722), .ZN(n6105) );
  CLKBUF_X4 U4644 ( .I(n52686), .Z(n24647) );
  CLKBUF_X2 U25333 ( .I(n54037), .Z(n58656) );
  CLKBUF_X4 U574 ( .I(n52381), .Z(n54605) );
  CLKBUF_X2 U634 ( .I(n51837), .Z(n54067) );
  CLKBUF_X2 U48825 ( .I(n57074), .Z(n60934) );
  INV_X2 U7920 ( .I(n57074), .ZN(n15498) );
  CLKBUF_X2 U42353 ( .I(n52862), .Z(n60498) );
  INV_X2 U40273 ( .I(n52952), .ZN(n52488) );
  CLKBUF_X2 U15002 ( .I(n55656), .Z(n23447) );
  INV_X2 U44162 ( .I(n60710), .ZN(n61693) );
  NAND2_X1 U55227 ( .A1(n56980), .A2(n52888), .ZN(n52889) );
  NOR2_X1 U8523 ( .A1(n52237), .A2(n1372), .ZN(n52737) );
  CLKBUF_X4 U528 ( .I(n25936), .Z(n15434) );
  INV_X1 U432 ( .I(n23248), .ZN(n53205) );
  INV_X2 U7900 ( .I(n53023), .ZN(n50462) );
  INV_X2 U22693 ( .I(n21453), .ZN(n57000) );
  CLKBUF_X1 U30738 ( .I(n55908), .Z(n59192) );
  INV_X2 U42946 ( .I(n55287), .ZN(n6531) );
  CLKBUF_X2 U5535 ( .I(n56269), .Z(n58050) );
  INV_X2 U426 ( .I(n12573), .ZN(n1601) );
  NAND2_X1 U14915 ( .A1(n53192), .A2(n64910), .ZN(n9963) );
  NAND2_X1 U27391 ( .A1(n53590), .A2(n23025), .ZN(n7427) );
  NAND2_X1 U35607 ( .A1(n56254), .A2(n56411), .ZN(n19908) );
  OR2_X1 U24846 ( .A1(n51884), .A2(n57225), .Z(n5175) );
  NOR2_X1 U12032 ( .A1(n5569), .A2(n16848), .ZN(n55263) );
  NAND2_X1 U12234 ( .A1(n53435), .A2(n57047), .ZN(n8448) );
  CLKBUF_X2 U5518 ( .I(n25080), .Z(n58303) );
  NAND2_X1 U55820 ( .A1(n54502), .A2(n59764), .ZN(n54503) );
  NAND3_X1 U37344 ( .A1(n54462), .A2(n17935), .A3(n54463), .ZN(n54464) );
  INV_X2 U3960 ( .I(n2997), .ZN(n2890) );
  NAND2_X1 U47292 ( .A1(n54801), .A2(n23122), .ZN(n60845) );
  NAND2_X1 U8502 ( .A1(n54100), .A2(n54446), .ZN(n13793) );
  NAND3_X1 U34980 ( .A1(n52046), .A2(n52045), .A3(n52920), .ZN(n19132) );
  NAND2_X1 U35187 ( .A1(n21643), .A2(n23334), .ZN(n52241) );
  AOI21_X1 U4586 ( .A1(n57401), .A2(n9003), .B(n5550), .ZN(n57641) );
  NAND2_X1 U335 ( .A1(n59812), .A2(n61371), .ZN(n58912) );
  NAND2_X1 U35649 ( .A1(n17138), .A2(n15909), .ZN(n54648) );
  NAND2_X1 U6383 ( .A1(n9003), .A2(n55924), .ZN(n60373) );
  NAND2_X1 U12174 ( .A1(n51712), .A2(n13940), .ZN(n53878) );
  NAND2_X1 U34877 ( .A1(n53392), .A2(n20630), .ZN(n53394) );
  NAND2_X1 U10702 ( .A1(n4864), .A2(n55970), .ZN(n9264) );
  OAI21_X1 U14671 ( .A1(n8447), .A2(n53434), .B(n8445), .ZN(n53447) );
  NAND2_X1 U4568 ( .A1(n56557), .A2(n56554), .ZN(n5330) );
  NAND2_X1 U48419 ( .A1(n53853), .A2(n53617), .ZN(n11869) );
  NAND3_X1 U17699 ( .A1(n52874), .A2(n10237), .A3(n52873), .ZN(n50547) );
  NAND2_X1 U14602 ( .A1(n20927), .A2(n20926), .ZN(n25089) );
  OAI21_X1 U30549 ( .A1(n52765), .A2(n53575), .B(n53589), .ZN(n10214) );
  INV_X1 U31035 ( .I(n22232), .ZN(n17054) );
  NAND2_X1 U29267 ( .A1(n58976), .A2(n54811), .ZN(n13142) );
  NOR2_X1 U39159 ( .A1(n17010), .A2(n60097), .ZN(n4117) );
  NAND2_X1 U14683 ( .A1(n24319), .A2(n24320), .ZN(n20588) );
  NAND2_X1 U5593 ( .A1(n7893), .A2(n7892), .ZN(n7891) );
  BUF_X4 U26874 ( .I(n2348), .Z(n2329) );
  NAND2_X1 U42874 ( .A1(n60574), .A2(n56663), .ZN(n56562) );
  NAND2_X1 U277 ( .A1(n57950), .A2(n50206), .ZN(n17261) );
  CLKBUF_X8 U203 ( .I(n56965), .Z(n14708) );
  CLKBUF_X8 U3642 ( .I(n52248), .Z(n1257) );
  CLKBUF_X4 U13327 ( .I(n52223), .Z(n55644) );
  INV_X1 U14503 ( .I(n56845), .ZN(n56844) );
  CLKBUF_X4 U23963 ( .I(n53518), .Z(n25789) );
  INV_X1 U37364 ( .I(n57120), .ZN(n57154) );
  CLKBUF_X2 U9803 ( .I(n25604), .Z(n7093) );
  INV_X1 U4057 ( .I(n53140), .ZN(n53128) );
  INV_X2 U133 ( .I(n63931), .ZN(n53320) );
  INV_X1 U35639 ( .I(n50830), .ZN(n20300) );
  OAI21_X1 U5821 ( .A1(n53048), .A2(n53109), .B(n53104), .ZN(n53049) );
  NAND2_X1 U5000 ( .A1(n8949), .A2(n15933), .ZN(n4874) );
  NOR2_X1 U14496 ( .A1(n52879), .A2(n53070), .ZN(n5620) );
  NAND3_X1 U55704 ( .A1(n54179), .A2(n10480), .A3(n54188), .ZN(n54157) );
  NAND2_X1 U7380 ( .A1(n53665), .A2(n53649), .ZN(n53670) );
  NOR2_X1 U3833 ( .A1(n53131), .A2(n12209), .ZN(n12208) );
  NOR2_X1 U4579 ( .A1(n20605), .A2(n1579), .ZN(n61126) );
  NAND3_X1 U55773 ( .A1(n54356), .A2(n54390), .A3(n54394), .ZN(n54357) );
  NAND2_X1 U10649 ( .A1(n13712), .A2(n54186), .ZN(n10318) );
  NAND2_X1 U56434 ( .A1(n56110), .A2(n9567), .ZN(n56111) );
  NAND2_X1 U14524 ( .A1(n15858), .A2(n9533), .ZN(n53159) );
  INV_X1 U14359 ( .I(n16828), .ZN(n16827) );
  NOR2_X1 U12378 ( .A1(n52304), .A2(n55617), .ZN(n58721) );
  NAND2_X1 U32529 ( .A1(n55230), .A2(n22815), .ZN(n55240) );
  NAND3_X1 U37455 ( .A1(n22859), .A2(n55791), .A3(n22858), .ZN(n23633) );
  NOR2_X1 U14383 ( .A1(n56970), .A2(n1257), .ZN(n12400) );
  BUF_X2 U9068 ( .I(Key[35]), .Z(n53705) );
  CLKBUF_X4 U14309 ( .I(Key[138]), .Z(n56008) );
  CLKBUF_X4 U19929 ( .I(Key[182]), .Z(n56915) );
  BUF_X2 U19860 ( .I(n26161), .Z(n11514) );
  CLKBUF_X2 U19878 ( .I(n26986), .Z(n23800) );
  BUF_X2 U44340 ( .I(n26866), .Z(n27822) );
  INV_X1 U37775 ( .I(n26866), .ZN(n28470) );
  INV_X1 U1 ( .I(n58084), .ZN(n56933) );
  CLKBUF_X2 U31406 ( .I(n16446), .Z(n59279) );
  BUF_X4 U5841 ( .I(n26264), .Z(n28067) );
  BUF_X2 U19823 ( .I(n24920), .Z(n9884) );
  CLKBUF_X2 U8585 ( .I(n26811), .Z(n58971) );
  BUF_X2 U19851 ( .I(n51977), .Z(n9722) );
  INV_X2 U19781 ( .I(n29709), .ZN(n29714) );
  AND2_X1 U33589 ( .A1(n28217), .A2(n3087), .Z(n13917) );
  CLKBUF_X2 U41358 ( .I(n27097), .Z(n60355) );
  CLKBUF_X2 U6267 ( .I(n34834), .Z(n59638) );
  BUF_X2 U9028 ( .I(n20734), .Z(n1891) );
  CLKBUF_X2 U12057 ( .I(n13763), .Z(n11605) );
  INV_X1 U14245 ( .I(n27121), .ZN(n21204) );
  BUF_X2 U19763 ( .I(n29312), .Z(n20665) );
  INV_X1 U43155 ( .I(n23487), .ZN(n28445) );
  CLKBUF_X4 U3389 ( .I(n28106), .Z(n23071) );
  BUF_X4 U9027 ( .I(n29628), .Z(n19290) );
  NAND2_X1 U45143 ( .A1(n28860), .A2(n20665), .ZN(n28861) );
  BUF_X1 U5324 ( .I(n32232), .Z(n238) );
  INV_X2 U22256 ( .I(n3626), .ZN(n28222) );
  NOR2_X1 U28604 ( .A1(n27615), .A2(n8518), .ZN(n14757) );
  AOI21_X1 U19508 ( .A1(n29369), .A2(n29368), .B(n17460), .ZN(n17882) );
  OAI21_X1 U44960 ( .A1(n28334), .A2(n28333), .B(n28332), .ZN(n28337) );
  AOI21_X1 U14062 ( .A1(n28218), .A2(n28219), .B(n24060), .ZN(n14152) );
  AOI21_X1 U26034 ( .A1(n28845), .A2(n27349), .B(n6382), .ZN(n27350) );
  NAND2_X1 U38471 ( .A1(n22442), .A2(n60011), .ZN(n60010) );
  NOR3_X1 U19425 ( .A1(n2113), .A2(n2111), .A3(n2110), .ZN(n8511) );
  OAI21_X1 U21102 ( .A1(n28413), .A2(n28412), .B(n58927), .ZN(n16860) );
  BUF_X4 U19368 ( .I(n30413), .Z(n11092) );
  CLKBUF_X4 U3145 ( .I(n29010), .Z(n23918) );
  CLKBUF_X2 U42886 ( .I(n29432), .Z(n60575) );
  BUF_X4 U11887 ( .I(n26650), .Z(n18736) );
  INV_X2 U20526 ( .I(n22181), .ZN(n17411) );
  CLKBUF_X4 U8976 ( .I(n29269), .Z(n15689) );
  INV_X1 U5088 ( .I(n12894), .ZN(n28942) );
  INV_X1 U8223 ( .I(n31049), .ZN(n31052) );
  INV_X1 U10439 ( .I(n18872), .ZN(n31204) );
  CLKBUF_X2 U54567 ( .I(n24123), .Z(n61229) );
  INV_X1 U44443 ( .I(n30551), .ZN(n30556) );
  OAI22_X1 U45207 ( .A1(n29037), .A2(n30724), .B1(n29036), .B2(n29224), .ZN(
        n29038) );
  NOR2_X1 U19149 ( .A1(n13444), .A2(n13447), .ZN(n27910) );
  INV_X1 U7567 ( .I(n30263), .ZN(n1348) );
  INV_X1 U19039 ( .I(n29936), .ZN(n30814) );
  INV_X2 U4672 ( .I(n9787), .ZN(n1835) );
  CLKBUF_X2 U11753 ( .I(n16759), .Z(n16758) );
  NOR3_X1 U5577 ( .A1(n19635), .A2(n29243), .A3(n15665), .ZN(n302) );
  BUF_X2 U11742 ( .I(n33889), .Z(n13181) );
  CLKBUF_X4 U2807 ( .I(n17617), .Z(n17668) );
  INV_X1 U18860 ( .I(n33178), .ZN(n2427) );
  BUF_X2 U6171 ( .I(n31438), .Z(n433) );
  CLKBUF_X2 U48360 ( .I(n20469), .Z(n60902) );
  CLKBUF_X2 U22275 ( .I(n9883), .Z(n58234) );
  BUF_X2 U26840 ( .I(n32420), .Z(n10535) );
  CLKBUF_X4 U8886 ( .I(n35002), .Z(n15588) );
  CLKBUF_X2 U6168 ( .I(n227), .Z(n59553) );
  CLKBUF_X2 U3469 ( .I(n11981), .Z(n2232) );
  BUF_X2 U13706 ( .I(n23834), .Z(n10091) );
  CLKBUF_X2 U18724 ( .I(n32295), .Z(n20660) );
  INV_X2 U34581 ( .I(n15318), .ZN(n35687) );
  INV_X2 U4303 ( .I(n15552), .ZN(n1543) );
  CLKBUF_X1 U9190 ( .I(n2989), .Z(n7272) );
  CLKBUF_X2 U42934 ( .I(n33628), .Z(n24093) );
  CLKBUF_X2 U6136 ( .I(n60883), .Z(n58036) );
  CLKBUF_X2 U19408 ( .I(n262), .Z(n57898) );
  INV_X2 U29328 ( .I(n9369), .ZN(n34353) );
  INV_X1 U18729 ( .I(n35785), .ZN(n34422) );
  CLKBUF_X2 U18615 ( .I(n32975), .Z(n7116) );
  CLKBUF_X2 U27691 ( .I(n6206), .Z(n60527) );
  CLKBUF_X4 U6072 ( .I(n6529), .Z(n445) );
  BUF_X2 U44579 ( .I(n34766), .Z(n60738) );
  NAND3_X1 U18504 ( .A1(n34134), .A2(n34142), .A3(n33660), .ZN(n33666) );
  NAND2_X1 U47593 ( .A1(n63249), .A2(n34356), .ZN(n32931) );
  INV_X1 U8054 ( .I(n34142), .ZN(n59399) );
  NAND2_X1 U18506 ( .A1(n34189), .A2(n17420), .ZN(n3122) );
  NAND2_X1 U36409 ( .A1(n33956), .A2(n33957), .ZN(n18451) );
  INV_X1 U26201 ( .I(n6526), .ZN(n35623) );
  NAND2_X1 U24117 ( .A1(n3670), .A2(n3668), .ZN(n58483) );
  NAND2_X1 U23536 ( .A1(n14147), .A2(n32360), .ZN(n13501) );
  NOR2_X1 U7984 ( .A1(n57273), .A2(n9717), .ZN(n26059) );
  AOI21_X1 U18178 ( .A1(n35323), .A2(n6520), .B(n35322), .ZN(n11669) );
  AOI21_X1 U35041 ( .A1(n34090), .A2(n34089), .B(n4075), .ZN(n34091) );
  NAND2_X1 U18346 ( .A1(n34176), .A2(n60628), .ZN(n34183) );
  AOI21_X1 U18149 ( .A1(n33223), .A2(n18475), .B(n20582), .ZN(n5255) );
  NAND2_X1 U32640 ( .A1(n33380), .A2(n33378), .ZN(n59442) );
  NOR2_X1 U21097 ( .A1(n58483), .A2(n9277), .ZN(n58102) );
  BUF_X4 U8227 ( .I(n36453), .Z(n1419) );
  CLKBUF_X4 U3670 ( .I(n35898), .Z(n23584) );
  NAND2_X1 U27011 ( .A1(n7730), .A2(n31721), .ZN(n16698) );
  BUF_X2 U27232 ( .I(n24357), .Z(n4151) );
  BUF_X2 U18004 ( .I(n37405), .Z(n17660) );
  BUF_X2 U9531 ( .I(n61703), .Z(n9633) );
  OAI22_X1 U33030 ( .A1(n61940), .A2(n15034), .B1(n7705), .B2(n23257), .ZN(
        n36223) );
  OAI21_X1 U13368 ( .A1(n36456), .A2(n1792), .B(n15034), .ZN(n20956) );
  NAND2_X1 U2231 ( .A1(n36676), .A2(n60374), .ZN(n17663) );
  CLKBUF_X4 U13443 ( .I(n60014), .Z(n6440) );
  INV_X1 U5012 ( .I(n35379), .ZN(n35382) );
  NAND2_X1 U13379 ( .A1(n35065), .A2(n35423), .ZN(n26016) );
  NAND2_X1 U17998 ( .A1(n65234), .A2(n12885), .ZN(n36339) );
  NOR2_X1 U38231 ( .A1(n17030), .A2(n63838), .ZN(n34838) );
  INV_X1 U18087 ( .I(n63838), .ZN(n36077) );
  NOR2_X1 U13392 ( .A1(n35423), .A2(n12885), .ZN(n35064) );
  NOR2_X1 U24858 ( .A1(n5185), .A2(n5900), .ZN(n35059) );
  NAND2_X1 U35787 ( .A1(n18076), .A2(n36275), .ZN(n23367) );
  NAND2_X1 U2205 ( .A1(n35563), .A2(n35562), .ZN(n13301) );
  NOR2_X1 U8787 ( .A1(n2279), .A2(n63817), .ZN(n15449) );
  NOR2_X1 U48504 ( .A1(n36389), .A2(n36385), .ZN(n35455) );
  INV_X1 U17953 ( .I(n37387), .ZN(n12236) );
  INV_X1 U17679 ( .I(n37396), .ZN(n6139) );
  NOR2_X1 U17966 ( .A1(n19777), .A2(n18677), .ZN(n60882) );
  NAND2_X1 U2762 ( .A1(n36267), .A2(n22301), .ZN(n59973) );
  AOI21_X1 U17830 ( .A1(n36496), .A2(n64093), .B(n34488), .ZN(n21673) );
  AOI21_X1 U28489 ( .A1(n34694), .A2(n63697), .B(n58909), .ZN(n34699) );
  NAND2_X1 U2695 ( .A1(n59058), .A2(n59123), .ZN(n33333) );
  NOR2_X1 U2821 ( .A1(n23367), .A2(n59657), .ZN(n13534) );
  INV_X2 U26796 ( .I(n37821), .ZN(n21494) );
  BUF_X2 U20857 ( .I(n23535), .Z(n2583) );
  CLKBUF_X2 U25937 ( .I(n14737), .Z(n58725) );
  BUF_X4 U6156 ( .I(n41383), .Z(n473) );
  CLKBUF_X2 U33812 ( .I(n23933), .Z(n59591) );
  CLKBUF_X4 U6392 ( .I(n39817), .Z(n41384) );
  BUF_X2 U41895 ( .I(n38811), .Z(n41453) );
  CLKBUF_X4 U17471 ( .I(n61705), .Z(n22759) );
  BUF_X2 U17472 ( .I(n1410), .Z(n4581) );
  BUF_X4 U17530 ( .I(n15963), .Z(n59601) );
  BUF_X1 U6010 ( .I(n17966), .Z(n58046) );
  CLKBUF_X2 U6024 ( .I(n38023), .Z(n57791) );
  CLKBUF_X2 U2089 ( .I(n20348), .Z(n11664) );
  CLKBUF_X1 U5218 ( .I(n40947), .Z(n212) );
  CLKBUF_X2 U11349 ( .I(n39007), .Z(n41397) );
  CLKBUF_X2 U13157 ( .I(n39904), .Z(n9808) );
  NAND2_X1 U36716 ( .A1(n17752), .A2(n42477), .ZN(n42466) );
  INV_X1 U35074 ( .I(n38939), .ZN(n41222) );
  NOR2_X1 U51221 ( .A1(n109), .A2(n8017), .ZN(n41929) );
  INV_X1 U27690 ( .I(n7618), .ZN(n40853) );
  OAI21_X1 U50517 ( .A1(n40591), .A2(n41073), .B(n14132), .ZN(n39783) );
  BUF_X2 U7616 ( .I(n41017), .Z(n58851) );
  CLKBUF_X2 U50712 ( .I(n40980), .Z(n61000) );
  NAND2_X1 U39249 ( .A1(n40754), .A2(n7165), .ZN(n18664) );
  BUF_X2 U39481 ( .I(n11664), .Z(n60143) );
  CLKBUF_X2 U40281 ( .I(n40469), .Z(n60229) );
  INV_X2 U39280 ( .I(n41289), .ZN(n18717) );
  INV_X2 U2071 ( .I(n39904), .ZN(n1733) );
  OAI21_X1 U25052 ( .A1(n23833), .A2(n5362), .B(n7257), .ZN(n5392) );
  INV_X1 U10107 ( .I(n40759), .ZN(n39806) );
  NOR3_X1 U50667 ( .A1(n11345), .A2(n25661), .A3(n2234), .ZN(n40165) );
  INV_X1 U17171 ( .I(n988), .ZN(n41274) );
  OAI21_X1 U27262 ( .A1(n40751), .A2(n40750), .B(n41470), .ZN(n10611) );
  NAND2_X1 U40882 ( .A1(n20991), .A2(n40643), .ZN(n40538) );
  NAND2_X1 U50646 ( .A1(n40074), .A2(n63952), .ZN(n40078) );
  INV_X1 U11265 ( .I(n41954), .ZN(n1727) );
  NAND2_X1 U17278 ( .A1(n40761), .A2(n40760), .ZN(n18668) );
  OAI21_X1 U23871 ( .A1(n41310), .A2(n41810), .B(n7094), .ZN(n4683) );
  OAI22_X1 U49553 ( .A1(n39418), .A2(n6576), .B1(n38031), .B2(n11126), .ZN(
        n38032) );
  NAND2_X1 U43272 ( .A1(n58599), .A2(n10341), .ZN(n40111) );
  AOI22_X1 U17065 ( .A1(n40240), .A2(n2159), .B1(n40242), .B2(n40241), .ZN(
        n40243) );
  NAND2_X1 U13072 ( .A1(n42516), .A2(n42517), .ZN(n12868) );
  NAND2_X1 U10165 ( .A1(n42450), .A2(n25606), .ZN(n41307) );
  BUF_X2 U7482 ( .I(n4968), .Z(n61159) );
  NAND2_X2 U7165 ( .A1(n8131), .A2(n40833), .ZN(n41137) );
  NAND2_X1 U10075 ( .A1(n40158), .A2(n9215), .ZN(n11124) );
  INV_X1 U17225 ( .I(n40221), .ZN(n40289) );
  INV_X1 U10081 ( .I(n16970), .ZN(n7696) );
  NAND2_X1 U9408 ( .A1(n40107), .A2(n64566), .ZN(n8440) );
  NAND2_X1 U17103 ( .A1(n10569), .A2(n22983), .ZN(n39898) );
  OAI21_X1 U10089 ( .A1(n41937), .A2(n41936), .B(n41935), .ZN(n41938) );
  INV_X1 U6579 ( .I(n41823), .ZN(n608) );
  OAI22_X1 U56837 ( .A1(n39830), .A2(n40434), .B1(n39831), .B2(n41113), .ZN(
        n61455) );
  NOR2_X1 U12929 ( .A1(n17294), .A2(n6223), .ZN(n5870) );
  NOR2_X1 U12969 ( .A1(n7356), .A2(n3495), .ZN(n3492) );
  CLKBUF_X4 U24960 ( .I(n23230), .Z(n13389) );
  BUF_X4 U5907 ( .I(n41614), .Z(n1499) );
  CLKBUF_X4 U1731 ( .I(n42636), .Z(n24884) );
  CLKBUF_X4 U16903 ( .I(n43656), .Z(n2824) );
  CLKBUF_X2 U35693 ( .I(n23877), .Z(n59771) );
  CLKBUF_X2 U1745 ( .I(n19537), .Z(n23350) );
  NAND3_X1 U4383 ( .A1(n40270), .A2(n21925), .A3(n21924), .ZN(n42356) );
  INV_X2 U13280 ( .I(n16850), .ZN(n4575) );
  AND2_X1 U12513 ( .A1(n41675), .A2(n4714), .Z(n57241) );
  CLKBUF_X2 U5915 ( .I(n41997), .Z(n60792) );
  NOR2_X1 U1648 ( .A1(n42865), .A2(n295), .ZN(n21336) );
  CLKBUF_X1 U47297 ( .I(n11039), .Z(n60846) );
  NAND2_X1 U51288 ( .A1(n42161), .A2(n8185), .ZN(n43611) );
  INV_X1 U3830 ( .I(n21935), .ZN(n43118) );
  BUF_X2 U16797 ( .I(n43289), .Z(n7349) );
  NAND2_X1 U36822 ( .A1(n43816), .A2(n42347), .ZN(n17706) );
  NOR2_X1 U1639 ( .A1(n24779), .A2(n12775), .ZN(n42980) );
  CLKBUF_X4 U23041 ( .I(n18482), .Z(n4275) );
  CLKBUF_X2 U25659 ( .I(n43695), .Z(n58693) );
  AOI21_X1 U50181 ( .A1(n41661), .A2(n17848), .B(n43028), .ZN(n39084) );
  INV_X2 U10059 ( .I(n42407), .ZN(n1396) );
  OAI22_X1 U22097 ( .A1(n20690), .A2(n43316), .B1(n43327), .B2(n59139), .ZN(
        n42767) );
  NOR2_X1 U16672 ( .A1(n42772), .A2(n20690), .ZN(n4420) );
  INV_X1 U16556 ( .I(n43697), .ZN(n37920) );
  NAND2_X1 U36054 ( .A1(n43690), .A2(n62326), .ZN(n16409) );
  INV_X1 U50915 ( .I(n40886), .ZN(n40887) );
  NAND2_X1 U51587 ( .A1(n43392), .A2(n43690), .ZN(n43394) );
  NAND3_X1 U10011 ( .A1(n43715), .A2(n10303), .A3(n10302), .ZN(n4519) );
  NOR2_X1 U16532 ( .A1(n43153), .A2(n13528), .ZN(n43172) );
  NAND2_X1 U4870 ( .A1(n43361), .A2(n14920), .ZN(n59066) );
  NAND2_X1 U16554 ( .A1(n43837), .A2(n59650), .ZN(n11748) );
  NOR2_X1 U51399 ( .A1(n65228), .A2(n42630), .ZN(n42631) );
  INV_X1 U8673 ( .I(n40899), .ZN(n6937) );
  NAND3_X2 U51289 ( .A1(n42162), .A2(n43336), .A3(n43611), .ZN(n42164) );
  NAND2_X1 U14582 ( .A1(n42941), .A2(n42943), .ZN(n9849) );
  AOI21_X1 U16397 ( .A1(n15234), .A2(n42555), .B(n15233), .ZN(n15232) );
  NOR2_X1 U5835 ( .A1(n57315), .A2(n58171), .ZN(n42887) );
  OAI22_X1 U51385 ( .A1(n42575), .A2(n42574), .B1(n42573), .B2(n42892), .ZN(
        n42576) );
  AOI21_X1 U6118 ( .A1(n43126), .A2(n43127), .B(n43125), .ZN(n43128) );
  INV_X1 U10801 ( .I(n43021), .ZN(n59686) );
  INV_X1 U7223 ( .I(n22802), .ZN(n58882) );
  OAI22_X1 U5839 ( .A1(n42013), .A2(n42012), .B1(n24981), .B2(n43091), .ZN(
        n42015) );
  NAND2_X1 U34574 ( .A1(n59686), .A2(n39173), .ZN(n1912) );
  NAND3_X1 U51612 ( .A1(n43474), .A2(n43473), .A3(n43472), .ZN(n43480) );
  INV_X2 U31889 ( .I(n60486), .ZN(n46251) );
  CLKBUF_X2 U8641 ( .I(n20208), .Z(n7132) );
  NAND3_X1 U50771 ( .A1(n40452), .A2(n40451), .A3(n40450), .ZN(n40457) );
  NAND2_X1 U1431 ( .A1(n10532), .A2(n26036), .ZN(n46292) );
  CLKBUF_X2 U16378 ( .I(n45041), .Z(n24062) );
  BUF_X2 U6931 ( .I(n22890), .Z(n59984) );
  CLKBUF_X2 U56841 ( .I(n22143), .Z(n61457) );
  INV_X1 U16334 ( .I(n11879), .ZN(n45356) );
  CLKBUF_X1 U5793 ( .I(n48546), .Z(n59160) );
  CLKBUF_X4 U23436 ( .I(n44861), .Z(n47900) );
  CLKBUF_X4 U37714 ( .I(n48097), .Z(n24099) );
  CLKBUF_X4 U12696 ( .I(n47819), .Z(n14630) );
  INV_X1 U30074 ( .I(n9926), .ZN(n16194) );
  CLKBUF_X2 U16291 ( .I(n48555), .Z(n22874) );
  INV_X1 U12708 ( .I(n21067), .ZN(n45140) );
  BUF_X2 U16298 ( .I(n48130), .Z(n22574) );
  BUF_X2 U16258 ( .I(n21231), .Z(n10626) );
  CLKBUF_X4 U41723 ( .I(n61668), .Z(n22436) );
  INV_X2 U29327 ( .I(n9368), .ZN(n48212) );
  INV_X2 U1315 ( .I(n48095), .ZN(n21305) );
  BUF_X2 U5782 ( .I(n47860), .Z(n10405) );
  INV_X2 U33469 ( .I(n1085), .ZN(n47578) );
  CLKBUF_X2 U12694 ( .I(n47314), .Z(n7389) );
  CLKBUF_X2 U41437 ( .I(n24545), .Z(n60358) );
  INV_X2 U12680 ( .I(n6933), .ZN(n3203) );
  OAI21_X1 U11084 ( .A1(n60386), .A2(n22574), .B(n7186), .ZN(n3105) );
  NOR3_X1 U10993 ( .A1(n1082), .A2(n48654), .A3(n46106), .ZN(n5717) );
  BUF_X2 U5729 ( .I(n48577), .Z(n59269) );
  NAND2_X1 U52551 ( .A1(n45964), .A2(n23894), .ZN(n45563) );
  INV_X1 U52813 ( .I(n48581), .ZN(n46175) );
  CLKBUF_X2 U5967 ( .I(n45591), .Z(n412) );
  INV_X1 U53578 ( .I(n48494), .ZN(n48498) );
  CLKBUF_X1 U5727 ( .I(n61717), .Z(n59959) );
  OAI22_X1 U15967 ( .A1(n47464), .A2(n47465), .B1(n47468), .B2(n4380), .ZN(
        n8156) );
  NAND2_X1 U1152 ( .A1(n45222), .A2(n23894), .ZN(n45565) );
  NAND2_X1 U16005 ( .A1(n12699), .A2(n12700), .ZN(n9642) );
  NAND2_X1 U16123 ( .A1(n46930), .A2(n47329), .ZN(n45622) );
  INV_X1 U16016 ( .I(n47813), .ZN(n47814) );
  OAI21_X1 U43415 ( .A1(n25476), .A2(n47292), .B(n47295), .ZN(n60637) );
  NOR2_X1 U38837 ( .A1(n9743), .A2(n9742), .ZN(n60063) );
  NOR2_X1 U12589 ( .A1(n47813), .A2(n12495), .ZN(n45310) );
  NAND3_X1 U52526 ( .A1(n60727), .A2(n45751), .A3(n15076), .ZN(n45500) );
  OAI22_X1 U53034 ( .A1(n47437), .A2(n46740), .B1(n46739), .B2(n46738), .ZN(
        n46741) );
  INV_X1 U52594 ( .I(n46865), .ZN(n45653) );
  OAI22_X1 U15920 ( .A1(n13446), .A2(n44485), .B1(n47261), .B2(n21793), .ZN(
        n13445) );
  AOI21_X1 U1179 ( .A1(n47805), .A2(n47804), .B(n57508), .ZN(n23266) );
  OAI21_X1 U23918 ( .A1(n47899), .A2(n47898), .B(n47897), .ZN(n47909) );
  NAND2_X1 U33514 ( .A1(n43831), .A2(n13782), .ZN(n23048) );
  NAND2_X1 U12534 ( .A1(n47027), .A2(n20725), .ZN(n47023) );
  INV_X1 U6819 ( .I(n44775), .ZN(n44199) );
  AOI21_X1 U33003 ( .A1(n45368), .A2(n46814), .B(n13053), .ZN(n15849) );
  CLKBUF_X4 U43443 ( .I(n44004), .Z(n49395) );
  NAND3_X1 U1051 ( .A1(n16877), .A2(n17033), .A3(n6607), .ZN(n16876) );
  NAND2_X1 U12555 ( .A1(n19652), .A2(n47139), .ZN(n14775) );
  OAI22_X1 U1260 ( .A1(n44281), .A2(n57625), .B1(n44283), .B2(n44282), .ZN(
        n44289) );
  OAI21_X1 U41856 ( .A1(n1646), .A2(n44204), .B(n44203), .ZN(n22603) );
  CLKBUF_X4 U7860 ( .I(n22805), .Z(n2878) );
  CLKBUF_X4 U39595 ( .I(n48852), .Z(n19175) );
  BUF_X2 U5638 ( .I(n17887), .Z(n60622) );
  CLKBUF_X4 U8575 ( .I(n20600), .Z(n23912) );
  CLKBUF_X4 U1033 ( .I(n16985), .Z(n16986) );
  CLKBUF_X4 U27138 ( .I(n23532), .Z(n6243) );
  CLKBUF_X2 U50891 ( .I(n47970), .Z(n61016) );
  BUF_X2 U1010 ( .I(n15386), .Z(n61612) );
  INV_X4 U24227 ( .I(n49063), .ZN(n11705) );
  CLKBUF_X4 U4880 ( .I(n15692), .Z(n8604) );
  INV_X1 U31196 ( .I(n22263), .ZN(n59249) );
  INV_X2 U6649 ( .I(n49684), .ZN(n17906) );
  INV_X1 U15647 ( .I(n49371), .ZN(n15039) );
  INV_X1 U12446 ( .I(n49600), .ZN(n48309) );
  NAND2_X1 U4810 ( .A1(n5517), .A2(n48332), .ZN(n47770) );
  NAND2_X1 U53742 ( .A1(n49039), .A2(n12580), .ZN(n49041) );
  OAI21_X1 U37220 ( .A1(n49099), .A2(n48709), .B(n49371), .ZN(n23028) );
  NAND2_X1 U15362 ( .A1(n19752), .A2(n48336), .ZN(n26120) );
  CLKBUF_X2 U23795 ( .I(n5743), .Z(n4647) );
  INV_X1 U11559 ( .I(n50428), .ZN(n50424) );
  INV_X1 U53435 ( .I(n49369), .ZN(n48010) );
  INV_X1 U52360 ( .I(n49764), .ZN(n45166) );
  NAND3_X1 U5912 ( .A1(n49066), .A2(n49067), .A3(n49068), .ZN(n393) );
  OAI21_X1 U23835 ( .A1(n406), .A2(n64170), .B(n49192), .ZN(n49193) );
  CLKBUF_X1 U10774 ( .I(n52079), .Z(n22790) );
  INV_X1 U37259 ( .I(n18479), .ZN(n18408) );
  CLKBUF_X2 U6541 ( .I(n50938), .Z(n58738) );
  BUF_X2 U11820 ( .I(n14975), .Z(n14974) );
  NOR2_X1 U32596 ( .A1(n15366), .A2(n48959), .ZN(n15365) );
  CLKBUF_X4 U617 ( .I(n52447), .Z(n22783) );
  CLKBUF_X2 U28747 ( .I(n50942), .Z(n58945) );
  CLKBUF_X4 U31069 ( .I(n51504), .Z(n10584) );
  CLKBUF_X4 U6551 ( .I(n51741), .Z(n20774) );
  CLKBUF_X2 U5564 ( .I(n51581), .Z(n59891) );
  INV_X2 U8529 ( .I(n51191), .ZN(n1288) );
  BUF_X2 U15049 ( .I(n20738), .Z(n10040) );
  INV_X2 U28089 ( .I(n24870), .ZN(n52479) );
  CLKBUF_X4 U6473 ( .I(n25519), .Z(n61443) );
  CLKBUF_X4 U607 ( .I(n1614), .Z(n61572) );
  INV_X2 U43692 ( .I(n25792), .ZN(n54436) );
  NAND2_X1 U38215 ( .A1(n833), .A2(n17003), .ZN(n52818) );
  INV_X2 U37774 ( .I(n61123), .ZN(n54023) );
  INV_X2 U10751 ( .I(n54599), .ZN(n1608) );
  INV_X1 U50166 ( .I(n55937), .ZN(n60977) );
  OR2_X1 U30053 ( .A1(n54942), .A2(n58994), .Z(n59079) );
  AND2_X1 U55923 ( .A1(n55250), .A2(n55401), .Z(n54791) );
  INV_X1 U12266 ( .I(n53436), .ZN(n53438) );
  NOR2_X1 U42476 ( .A1(n7027), .A2(n53586), .ZN(n53000) );
  OAI21_X1 U54958 ( .A1(n63339), .A2(n4181), .B(n57023), .ZN(n52233) );
  NOR3_X1 U7331 ( .A1(n1608), .A2(n54469), .A3(n54468), .ZN(n4895) );
  OAI21_X1 U9832 ( .A1(n55292), .A2(n9263), .B(n55974), .ZN(n4864) );
  NAND3_X1 U397 ( .A1(n53589), .A2(n533), .A3(n53587), .ZN(n2584) );
  NOR2_X1 U28943 ( .A1(n8904), .A2(n8903), .ZN(n8902) );
  NAND2_X1 U27153 ( .A1(n54648), .A2(n1613), .ZN(n54650) );
  NAND2_X1 U14731 ( .A1(n12729), .A2(n52239), .ZN(n14711) );
  AND3_X2 U10697 ( .A1(n55970), .A2(n55969), .A3(n1182), .Z(n55971) );
  NAND2_X1 U35596 ( .A1(n52767), .A2(n64521), .ZN(n16435) );
  NOR2_X1 U55650 ( .A1(n54316), .A2(n54066), .ZN(n54070) );
  NOR2_X1 U24484 ( .A1(n58553), .A2(n58552), .ZN(n7892) );
  NAND2_X1 U9827 ( .A1(n56557), .A2(n56556), .ZN(n56658) );
  NOR2_X1 U29997 ( .A1(n12833), .A2(n52842), .ZN(n12832) );
  OAI21_X1 U4158 ( .A1(n20965), .A2(n52986), .B(n54319), .ZN(n26151) );
  NOR2_X1 U20093 ( .A1(n17263), .A2(n17265), .ZN(n57950) );
  BUF_X2 U14579 ( .I(n56085), .Z(n24092) );
  CLKBUF_X8 U30336 ( .I(n55423), .Z(n55569) );
  CLKBUF_X2 U12340 ( .I(n63473), .Z(n23448) );
  CLKBUF_X4 U210 ( .I(n25621), .Z(n9338) );
  NOR2_X1 U27099 ( .A1(n24092), .A2(n56106), .ZN(n59587) );
  CLKBUF_X4 U39905 ( .I(n53677), .Z(n19475) );
  INV_X1 U14535 ( .I(n56158), .ZN(n15663) );
  AND3_X1 U40412 ( .A1(n56047), .A2(n63023), .A3(n61740), .Z(n56100) );
  CLKBUF_X1 U12284 ( .I(n53368), .Z(n60115) );
  INV_X2 U8469 ( .I(n61933), .ZN(n1579) );
  INV_X1 U55341 ( .I(n53165), .ZN(n53136) );
  NAND2_X1 U21761 ( .A1(n54892), .A2(n7680), .ZN(n54893) );
  NAND2_X1 U23774 ( .A1(n54584), .A2(n61556), .ZN(n58444) );
  INV_X1 U55725 ( .I(n54188), .ZN(n54190) );
  AOI21_X1 U54162 ( .A1(n1579), .A2(n50465), .B(n53759), .ZN(n50467) );
  NAND2_X1 U36519 ( .A1(n13492), .A2(n53815), .ZN(n7239) );
  NAND2_X1 U26894 ( .A1(n13512), .A2(n53313), .ZN(n61469) );
  NAND2_X2 U4088 ( .A1(n47274), .A2(n45551), .ZN(n47581) );
  INV_X2 U11235 ( .I(n40238), .ZN(n39419) );
  INV_X4 U19820 ( .I(n29641), .ZN(n20907) );
  INV_X2 U8315 ( .I(n28844), .ZN(n59090) );
  NAND2_X2 U3399 ( .A1(n29642), .A2(n28593), .ZN(n28844) );
  NAND3_X2 U20661 ( .A1(n2431), .A2(n45556), .A3(n45557), .ZN(n2434) );
  INV_X2 U18049 ( .I(n35602), .ZN(n17761) );
  INV_X4 U9968 ( .I(n47274), .ZN(n47281) );
  BUF_X2 U16364 ( .I(n45093), .Z(n23264) );
  BUF_X4 U12312 ( .I(n50111), .Z(n53915) );
  BUF_X4 U6121 ( .I(n37234), .Z(n461) );
  OAI22_X2 U34408 ( .A1(n8444), .A2(n30046), .B1(n25698), .B2(n30250), .ZN(
        n29052) );
  INV_X2 U6020 ( .I(n48554), .ZN(n48152) );
  INV_X4 U31822 ( .I(n1866), .ZN(n31187) );
  AOI22_X2 U8744 ( .A1(n29547), .A2(n18128), .B1(n29546), .B2(n20179), .ZN(
        n10170) );
  INV_X4 U19725 ( .I(n19223), .ZN(n28669) );
  INV_X2 U45036 ( .I(n28611), .ZN(n28612) );
  BUF_X2 U18750 ( .I(n32069), .Z(n21035) );
  OAI21_X2 U15292 ( .A1(n48687), .A2(n48686), .B(n48685), .ZN(n48695) );
  NOR2_X2 U12383 ( .A1(n48683), .A2(n48682), .ZN(n48687) );
  AOI22_X2 U55616 ( .A1(n53965), .A2(n53964), .B1(n53984), .B2(n54012), .ZN(
        n53977) );
  NAND2_X2 U19303 ( .A1(n4376), .A2(n2046), .ZN(n60879) );
  INV_X4 U13136 ( .I(n41859), .ZN(n1505) );
  NOR2_X2 U7219 ( .A1(n19792), .A2(n41658), .ZN(n2752) );
  OAI21_X2 U17923 ( .A1(n42717), .A2(n16135), .B(n41966), .ZN(n19792) );
  BUF_X4 U4106 ( .I(n12262), .Z(n244) );
  NOR2_X1 U12335 ( .A1(n46972), .A2(n46971), .ZN(n18474) );
  NOR2_X2 U50300 ( .A1(n40229), .A2(n15378), .ZN(n40288) );
  NOR3_X2 U7071 ( .A1(n77), .A2(n61547), .A3(n35755), .ZN(n33814) );
  NAND2_X1 U11589 ( .A1(n58116), .A2(n6583), .ZN(n46971) );
  INV_X2 U39839 ( .I(n40167), .ZN(n40069) );
  INV_X2 U48491 ( .I(n36842), .ZN(n35407) );
  NOR3_X2 U14051 ( .A1(n27940), .A2(n14257), .A3(n14256), .ZN(n23770) );
  NAND2_X2 U9768 ( .A1(n64614), .A2(n2902), .ZN(n8340) );
  BUF_X2 U8021 ( .I(n36638), .Z(n39646) );
  BUF_X2 U8490 ( .I(n14255), .Z(n1230) );
  INV_X2 U19389 ( .I(n11140), .ZN(n11139) );
  NOR2_X2 U11343 ( .A1(n10456), .A2(n49393), .ZN(n49332) );
  AOI22_X2 U45427 ( .A1(n29717), .A2(n31268), .B1(n31166), .B2(n31163), .ZN(
        n29720) );
  NAND3_X2 U22385 ( .A1(n54909), .A2(n23531), .A3(n54908), .ZN(n58247) );
  NAND2_X2 U2588 ( .A1(n13952), .A2(n16904), .ZN(n11666) );
  BUF_X4 U27277 ( .I(n51557), .Z(n56829) );
  BUF_X2 U666 ( .I(n51213), .Z(n22658) );
  NOR3_X1 U6100 ( .A1(n455), .A2(n40024), .A3(n40021), .ZN(n12147) );
  BUF_X4 U12707 ( .I(n45300), .Z(n47415) );
  BUF_X4 U15715 ( .I(n18976), .Z(n18918) );
  BUF_X4 U14623 ( .I(n56689), .Z(n20269) );
  INV_X2 U28753 ( .I(n10969), .ZN(n16487) );
  NOR2_X2 U753 ( .A1(n62593), .A2(n48768), .ZN(n9695) );
  INV_X4 U24624 ( .I(n9203), .ZN(n5903) );
  NOR4_X1 U51603 ( .A1(n43446), .A2(n43445), .A3(n43449), .A4(n43444), .ZN(
        n43451) );
  INV_X4 U16245 ( .I(n15757), .ZN(n48208) );
  NAND3_X2 U27409 ( .A1(n60252), .A2(n40704), .A3(n41438), .ZN(n40705) );
  OAI21_X2 U804 ( .A1(n18819), .A2(n18820), .B(n58983), .ZN(n58963) );
  INV_X4 U28721 ( .I(n10510), .ZN(n19228) );
  AOI21_X1 U20799 ( .A1(n40147), .A2(n1509), .B(n10542), .ZN(n2713) );
  NOR2_X1 U16482 ( .A1(n9503), .A2(n11363), .ZN(n19758) );
  INV_X2 U8791 ( .I(n36812), .ZN(n36307) );
  INV_X4 U16239 ( .I(n61668), .ZN(n47490) );
  NOR2_X1 U697 ( .A1(n45708), .A2(n58723), .ZN(n58541) );
  NOR2_X2 U24095 ( .A1(n47623), .A2(n45991), .ZN(n47245) );
  NOR2_X2 U26040 ( .A1(n38681), .A2(n6388), .ZN(n41716) );
  NAND2_X2 U25190 ( .A1(n10415), .A2(n4077), .ZN(n38681) );
  NAND3_X2 U32447 ( .A1(n14229), .A2(n28007), .A3(n28396), .ZN(n59420) );
  NOR2_X2 U35622 ( .A1(n19413), .A2(n19412), .ZN(n53419) );
  NOR2_X2 U37313 ( .A1(n53414), .A2(n61560), .ZN(n19413) );
  BUF_X4 U508 ( .I(n50601), .Z(n57070) );
  BUF_X4 U25564 ( .I(n6255), .Z(n5913) );
  NOR2_X2 U2467 ( .A1(n37394), .A2(n35934), .ZN(n36878) );
  INV_X4 U43069 ( .I(n41914), .ZN(n41258) );
  INV_X2 U13599 ( .I(n6205), .ZN(n24983) );
  NAND2_X2 U22250 ( .A1(n62975), .A2(n3596), .ZN(n48970) );
  AOI21_X2 U31072 ( .A1(n49433), .A2(n49374), .B(n49379), .ZN(n18226) );
  NAND3_X2 U27392 ( .A1(n53595), .A2(n53596), .A3(n53594), .ZN(n53597) );
  NAND3_X2 U11745 ( .A1(n49343), .A2(n50213), .A3(n50222), .ZN(n49105) );
  INV_X2 U39431 ( .I(n19004), .ZN(n42176) );
  INV_X2 U972 ( .I(n50213), .ZN(n18249) );
  AOI21_X2 U4681 ( .A1(n47244), .A2(n1069), .B(n22303), .ZN(n60430) );
  OAI21_X2 U50972 ( .A1(n23046), .A2(n25358), .B(n61710), .ZN(n41107) );
  INV_X2 U2358 ( .I(n36728), .ZN(n141) );
  NAND3_X2 U39294 ( .A1(n18750), .A2(n20653), .A3(n1324), .ZN(n55716) );
  INV_X2 U25989 ( .I(n6330), .ZN(n26856) );
  INV_X2 U10604 ( .I(n29154), .ZN(n9562) );
  INV_X1 U8385 ( .I(n22861), .ZN(n20929) );
  INV_X2 U6252 ( .I(n9548), .ZN(n9465) );
  CLKBUF_X2 U28581 ( .I(n24039), .Z(n58927) );
  BUF_X2 U19821 ( .I(n815), .Z(n4613) );
  BUF_X2 U9060 ( .I(n7322), .Z(n3617) );
  INV_X2 U40930 ( .I(n21265), .ZN(n28271) );
  BUF_X2 U8423 ( .I(n21265), .Z(n61021) );
  BUF_X2 U19852 ( .I(n26339), .Z(n28314) );
  NOR2_X1 U4635 ( .A1(n6727), .A2(n6726), .ZN(n57678) );
  INV_X2 U19863 ( .I(n23037), .ZN(n1893) );
  INV_X2 U20513 ( .I(n2295), .ZN(n23745) );
  INV_X1 U24126 ( .I(n58485), .ZN(n9017) );
  INV_X1 U38403 ( .I(n26986), .ZN(n27435) );
  INV_X1 U14285 ( .I(n26826), .ZN(n1571) );
  INV_X2 U12094 ( .I(n26431), .ZN(n28539) );
  INV_X1 U14262 ( .I(n27479), .ZN(n14603) );
  INV_X2 U29011 ( .I(n9017), .ZN(n27524) );
  AOI21_X1 U36612 ( .A1(n28400), .A2(n28004), .B(n26344), .ZN(n26346) );
  INV_X1 U22041 ( .I(n21955), .ZN(n3473) );
  BUF_X2 U14268 ( .I(n26192), .Z(n23596) );
  BUF_X2 U33373 ( .I(n22410), .Z(n59552) );
  CLKBUF_X2 U14187 ( .I(n11110), .Z(n4443) );
  INV_X2 U9039 ( .I(n7561), .ZN(n27690) );
  BUF_X2 U3420 ( .I(n29623), .Z(n23578) );
  INV_X2 U32786 ( .I(n27930), .ZN(n16654) );
  BUF_X2 U19853 ( .I(n29318), .Z(n23797) );
  INV_X2 U12075 ( .I(n23337), .ZN(n8889) );
  NOR2_X1 U3376 ( .A1(n10236), .A2(n29317), .ZN(n28853) );
  NAND2_X1 U42958 ( .A1(n27188), .A2(n28106), .ZN(n27573) );
  INV_X2 U23981 ( .I(n20519), .ZN(n26935) );
  INV_X2 U19892 ( .I(n27114), .ZN(n1895) );
  NAND2_X1 U42825 ( .A1(n29370), .A2(n29371), .ZN(n28812) );
  INV_X2 U33843 ( .I(n14312), .ZN(n28886) );
  NAND2_X1 U3383 ( .A1(n27171), .A2(n23328), .ZN(n27595) );
  AND2_X1 U6268 ( .A1(n24391), .A2(n23297), .Z(n20508) );
  INV_X1 U26404 ( .I(n25992), .ZN(n58792) );
  INV_X1 U7425 ( .I(n26414), .ZN(n28504) );
  INV_X1 U30581 ( .I(n13694), .ZN(n16446) );
  INV_X1 U43102 ( .I(n27709), .ZN(n27846) );
  CLKBUF_X2 U10612 ( .I(n27966), .Z(n9908) );
  NAND2_X1 U30723 ( .A1(n28271), .A2(n21946), .ZN(n28280) );
  INV_X2 U10554 ( .I(n28281), .ZN(n2176) );
  INV_X2 U43501 ( .I(n26670), .ZN(n27620) );
  BUF_X2 U8406 ( .I(n29310), .Z(n58108) );
  INV_X1 U19709 ( .I(n29325), .ZN(n20093) );
  NOR2_X1 U44637 ( .A1(n1444), .A2(n29153), .ZN(n27977) );
  NAND2_X1 U9010 ( .A1(n26527), .A2(n28241), .ZN(n24499) );
  NOR2_X1 U22830 ( .A1(n27962), .A2(n64374), .ZN(n27065) );
  NOR2_X1 U3322 ( .A1(n266), .A2(n23591), .ZN(n29147) );
  NAND2_X1 U5395 ( .A1(n26640), .A2(n26641), .ZN(n28301) );
  INV_X1 U3984 ( .I(n8528), .ZN(n7976) );
  NAND2_X1 U40544 ( .A1(n14604), .A2(n27483), .ZN(n27547) );
  NOR2_X1 U33590 ( .A1(n3580), .A2(n8478), .ZN(n28217) );
  INV_X2 U9016 ( .I(n26376), .ZN(n1320) );
  NOR2_X1 U3380 ( .A1(n21955), .A2(n15093), .ZN(n28216) );
  INV_X1 U35343 ( .I(n28808), .ZN(n17460) );
  NOR2_X1 U3310 ( .A1(n28414), .A2(n180), .ZN(n28405) );
  INV_X1 U26892 ( .I(n20716), .ZN(n7129) );
  INV_X1 U19602 ( .I(n65111), .ZN(n9561) );
  NAND2_X1 U32784 ( .A1(n29145), .A2(n16654), .ZN(n26714) );
  INV_X1 U3312 ( .I(n20473), .ZN(n27675) );
  INV_X1 U3297 ( .I(n28008), .ZN(n28418) );
  NOR2_X1 U44345 ( .A1(n28624), .A2(n28630), .ZN(n27821) );
  INV_X1 U9746 ( .I(n24921), .ZN(n17046) );
  INV_X2 U38257 ( .I(n29188), .ZN(n22351) );
  INV_X2 U19801 ( .I(n21774), .ZN(n14947) );
  INV_X1 U6414 ( .I(n28842), .ZN(n1358) );
  INV_X1 U3294 ( .I(n17522), .ZN(n28805) );
  INV_X1 U4875 ( .I(n22144), .ZN(n26968) );
  INV_X1 U50848 ( .I(n19566), .ZN(n61004) );
  INV_X1 U12076 ( .I(n22765), .ZN(n1570) );
  INV_X1 U42180 ( .I(n60505), .ZN(n60473) );
  NAND2_X1 U44352 ( .A1(n28632), .A2(n28630), .ZN(n27810) );
  INV_X2 U12053 ( .I(n20627), .ZN(n28622) );
  CLKBUF_X2 U8533 ( .I(n2342), .Z(n522) );
  NOR2_X1 U36607 ( .A1(n27136), .A2(n22408), .ZN(n28334) );
  INV_X1 U3271 ( .I(n28279), .ZN(n7558) );
  OAI22_X1 U8496 ( .A1(n28471), .A2(n63495), .B1(n28620), .B2(n28625), .ZN(
        n4606) );
  NOR2_X1 U8625 ( .A1(n27614), .A2(n23940), .ZN(n26468) );
  OAI22_X1 U56519 ( .A1(n29143), .A2(n29144), .B1(n60841), .B2(n18231), .ZN(
        n61387) );
  BUF_X2 U6144 ( .I(n10187), .Z(n6083) );
  INV_X1 U10584 ( .I(n28049), .ZN(n28320) );
  BUF_X2 U4003 ( .I(n27125), .Z(n61317) );
  INV_X1 U27965 ( .I(n17824), .ZN(n17879) );
  NAND2_X1 U8462 ( .A1(n28383), .A2(n23039), .ZN(n18753) );
  INV_X1 U8022 ( .I(n25993), .ZN(n22159) );
  INV_X1 U3233 ( .I(n26719), .ZN(n29132) );
  INV_X1 U22193 ( .I(n3591), .ZN(n28618) );
  INV_X1 U3273 ( .I(n28549), .ZN(n16812) );
  INV_X1 U28838 ( .I(n28012), .ZN(n8778) );
  CLKBUF_X4 U41886 ( .I(n27621), .Z(n22643) );
  NAND3_X1 U25943 ( .A1(n59935), .A2(n6382), .A3(n61004), .ZN(n6293) );
  INV_X1 U12056 ( .I(n22505), .ZN(n1568) );
  BUF_X4 U9040 ( .I(n27674), .Z(n1889) );
  NOR2_X1 U9753 ( .A1(n28034), .A2(n6215), .ZN(n27102) );
  NOR2_X1 U3276 ( .A1(n491), .A2(n22214), .ZN(n28183) );
  NOR2_X1 U31083 ( .A1(n10754), .A2(n28200), .ZN(n11374) );
  BUF_X2 U6140 ( .I(n25807), .Z(n469) );
  NAND2_X1 U23707 ( .A1(n26974), .A2(n58977), .ZN(n29358) );
  NOR2_X1 U29417 ( .A1(n27523), .A2(n9465), .ZN(n28352) );
  NOR2_X1 U3255 ( .A1(n27298), .A2(n29142), .ZN(n27928) );
  NAND2_X1 U3967 ( .A1(n28510), .A2(n28518), .ZN(n28506) );
  NAND2_X1 U22302 ( .A1(n27374), .A2(n23568), .ZN(n3904) );
  NOR2_X1 U14141 ( .A1(n13764), .A2(n27287), .ZN(n3793) );
  INV_X1 U39581 ( .I(n20714), .ZN(n28121) );
  NAND2_X1 U43985 ( .A1(n27120), .A2(n26533), .ZN(n26316) );
  INV_X2 U24628 ( .I(n4998), .ZN(n27532) );
  INV_X1 U14230 ( .I(n28350), .ZN(n26592) );
  NAND2_X1 U33534 ( .A1(n24734), .A2(n1894), .ZN(n27520) );
  INV_X2 U8486 ( .I(n27529), .ZN(n28341) );
  INV_X1 U3246 ( .I(n27936), .ZN(n28258) );
  NAND2_X1 U3962 ( .A1(n27274), .A2(n19328), .ZN(n29189) );
  INV_X1 U43309 ( .I(n23007), .ZN(n27560) );
  INV_X1 U3916 ( .I(n3087), .ZN(n1931) );
  NOR2_X1 U42313 ( .A1(n29616), .A2(n28176), .ZN(n28664) );
  INV_X1 U3301 ( .I(n27871), .ZN(n27875) );
  INV_X2 U28334 ( .I(n8437), .ZN(n8436) );
  INV_X1 U30580 ( .I(n26765), .ZN(n27877) );
  INV_X1 U8402 ( .I(n24836), .ZN(n28333) );
  NAND2_X1 U51295 ( .A1(n20930), .A2(n28884), .ZN(n28883) );
  INV_X1 U9049 ( .I(n28630), .ZN(n27812) );
  INV_X1 U39557 ( .I(n27328), .ZN(n28801) );
  NOR2_X1 U26820 ( .A1(n29353), .A2(n23496), .ZN(n29335) );
  INV_X1 U35857 ( .I(n27526), .ZN(n26054) );
  INV_X1 U25875 ( .I(n27047), .ZN(n6222) );
  AND2_X1 U3346 ( .A1(n23825), .A2(n28470), .Z(n29712) );
  INV_X1 U3279 ( .I(n18515), .ZN(n10625) );
  INV_X1 U8541 ( .I(n29351), .ZN(n27500) );
  INV_X1 U8450 ( .I(n10187), .ZN(n29162) );
  INV_X2 U3289 ( .I(n58977), .ZN(n29334) );
  NAND2_X1 U5448 ( .A1(n28471), .A2(n63495), .ZN(n28474) );
  NAND2_X1 U14161 ( .A1(n28007), .A2(n28401), .ZN(n3294) );
  NAND2_X1 U35320 ( .A1(n24499), .A2(n26528), .ZN(n25547) );
  NOR2_X1 U35833 ( .A1(n28176), .A2(n28175), .ZN(n26883) );
  INV_X1 U9008 ( .I(n26660), .ZN(n26661) );
  NAND2_X1 U8473 ( .A1(n28801), .A2(n19423), .ZN(n28815) );
  NOR2_X1 U44259 ( .A1(n1568), .A2(n23753), .ZN(n26733) );
  NAND2_X1 U34320 ( .A1(n28217), .A2(n14947), .ZN(n21805) );
  OAI21_X1 U44675 ( .A1(n27508), .A2(n7495), .B(n20930), .ZN(n27510) );
  AOI21_X1 U37924 ( .A1(n16523), .A2(n27483), .B(n27485), .ZN(n27466) );
  NOR2_X1 U45303 ( .A1(n29351), .A2(n29334), .ZN(n29336) );
  NAND2_X1 U17769 ( .A1(n29670), .A2(n19279), .ZN(n29667) );
  NOR2_X1 U8335 ( .A1(n57577), .A2(n57576), .ZN(n60537) );
  NOR3_X1 U8205 ( .A1(n7437), .A2(n5218), .A3(n29304), .ZN(n29300) );
  INV_X1 U37677 ( .I(n28620), .ZN(n28621) );
  NOR2_X1 U38575 ( .A1(n17619), .A2(n16278), .ZN(n27327) );
  NAND2_X1 U14206 ( .A1(n22234), .A2(n7886), .ZN(n20539) );
  INV_X1 U10550 ( .I(n28157), .ZN(n29308) );
  INV_X1 U45302 ( .I(n29333), .ZN(n29337) );
  NOR2_X1 U10567 ( .A1(n27976), .A2(n26742), .ZN(n27983) );
  NAND2_X1 U29705 ( .A1(n28808), .A2(n17824), .ZN(n26992) );
  NAND2_X1 U4293 ( .A1(n26706), .A2(n27229), .ZN(n16570) );
  NAND2_X1 U10548 ( .A1(n17047), .A2(n2662), .ZN(n27934) );
  NAND2_X1 U6972 ( .A1(n24001), .A2(n21132), .ZN(n28107) );
  NOR3_X1 U9021 ( .A1(n18006), .A2(n27655), .A3(n28483), .ZN(n28486) );
  NOR2_X1 U34446 ( .A1(n1565), .A2(n8436), .ZN(n27412) );
  NOR3_X1 U41444 ( .A1(n28137), .A2(n29286), .A3(n20034), .ZN(n29632) );
  NAND2_X1 U20008 ( .A1(n1880), .A2(n1931), .ZN(n3555) );
  NOR2_X1 U44149 ( .A1(n26979), .A2(n23504), .ZN(n29357) );
  NAND2_X1 U6697 ( .A1(n26680), .A2(n27523), .ZN(n28347) );
  INV_X1 U3204 ( .I(n10404), .ZN(n29111) );
  INV_X1 U33929 ( .I(n28127), .ZN(n29285) );
  INV_X1 U42685 ( .I(n28497), .ZN(n60542) );
  INV_X1 U12063 ( .I(n27568), .ZN(n1440) );
  NAND2_X1 U12021 ( .A1(n1359), .A2(n28260), .ZN(n29172) );
  INV_X1 U44140 ( .I(n26974), .ZN(n29350) );
  INV_X2 U3284 ( .I(n26626), .ZN(n28380) );
  INV_X1 U22579 ( .I(n3904), .ZN(n29108) );
  NOR3_X1 U3917 ( .A1(n14947), .A2(n8436), .A3(n10399), .ZN(n28214) );
  NAND2_X1 U19988 ( .A1(n1930), .A2(n57954), .ZN(n29131) );
  OAI22_X1 U21241 ( .A1(n28407), .A2(n9751), .B1(n11226), .B2(n2789), .ZN(
        n28413) );
  INV_X1 U11984 ( .I(n27614), .ZN(n22956) );
  AOI21_X1 U44294 ( .A1(n28451), .A2(n28453), .B(n28615), .ZN(n26788) );
  NAND2_X1 U34754 ( .A1(n26469), .A2(n26602), .ZN(n26472) );
  NOR2_X1 U44684 ( .A1(n27532), .A2(n27529), .ZN(n27531) );
  NAND4_X1 U43632 ( .A1(n29345), .A2(n25619), .A3(n7495), .A4(n62341), .ZN(
        n29346) );
  AOI22_X1 U45315 ( .A1(n29377), .A2(n29376), .B1(n29671), .B2(n57270), .ZN(
        n29390) );
  NAND2_X1 U41357 ( .A1(n21854), .A2(n28444), .ZN(n27861) );
  INV_X1 U14076 ( .I(n11065), .ZN(n20401) );
  AOI21_X1 U44180 ( .A1(n26550), .A2(n27109), .B(n26549), .ZN(n26553) );
  INV_X1 U31515 ( .I(n1970), .ZN(n28476) );
  OAI21_X1 U22494 ( .A1(n1320), .A2(n3823), .B(n3822), .ZN(n3821) );
  INV_X1 U3205 ( .I(n7437), .ZN(n14887) );
  AOI22_X1 U14038 ( .A1(n24232), .A2(n5290), .B1(n11875), .B2(n24231), .ZN(
        n11163) );
  NOR2_X1 U44037 ( .A1(n27572), .A2(n27579), .ZN(n26619) );
  OAI21_X1 U36679 ( .A1(n27565), .A2(n28380), .B(n20540), .ZN(n27566) );
  OAI22_X1 U14171 ( .A1(n10239), .A2(n28509), .B1(n24431), .B2(n8889), .ZN(
        n26415) );
  NOR2_X1 U44943 ( .A1(n93), .A2(n28235), .ZN(n28236) );
  NOR2_X1 U8527 ( .A1(n28471), .A2(n28624), .ZN(n26871) );
  INV_X1 U20004 ( .I(n1930), .ZN(n13657) );
  AOI22_X1 U44827 ( .A1(n27870), .A2(n28541), .B1(n27869), .B2(n28543), .ZN(
        n27873) );
  AOI22_X1 U32381 ( .A1(n26619), .A2(n12347), .B1(n26664), .B2(n27580), .ZN(
        n26368) );
  AOI22_X1 U3879 ( .A1(n28435), .A2(n28460), .B1(n26792), .B2(n28453), .ZN(
        n17528) );
  AOI22_X1 U19573 ( .A1(n28387), .A2(n7886), .B1(n64481), .B2(n28386), .ZN(
        n28390) );
  NAND3_X1 U40854 ( .A1(n27324), .A2(n27322), .A3(n27323), .ZN(n27335) );
  AOI22_X1 U19521 ( .A1(n14918), .A2(n13657), .B1(n29124), .B2(n13654), .ZN(
        n2544) );
  NOR2_X1 U35465 ( .A1(n26602), .A2(n22952), .ZN(n18759) );
  OAI22_X1 U37940 ( .A1(n17279), .A2(n17277), .B1(n27278), .B2(n60543), .ZN(
        n59934) );
  AOI21_X1 U11923 ( .A1(n27170), .A2(n9467), .B(n27176), .ZN(n9466) );
  AOI21_X1 U44178 ( .A1(n26548), .A2(n65037), .B(n27555), .ZN(n26555) );
  OAI21_X1 U39097 ( .A1(n18536), .A2(n27975), .B(n62234), .ZN(n60461) );
  NOR2_X1 U39803 ( .A1(n26639), .A2(n28378), .ZN(n20198) );
  NOR2_X1 U10576 ( .A1(n26805), .A2(n26794), .ZN(n27883) );
  NOR2_X1 U44488 ( .A1(n27176), .A2(n27075), .ZN(n27084) );
  OAI21_X1 U36614 ( .A1(n20628), .A2(n27809), .B(n28476), .ZN(n27819) );
  NOR2_X1 U38291 ( .A1(n59990), .A2(n59989), .ZN(n216) );
  INV_X1 U14106 ( .I(n28044), .ZN(n28047) );
  NOR3_X1 U6986 ( .A1(n26058), .A2(n26057), .A3(n26596), .ZN(n26056) );
  NAND2_X1 U8982 ( .A1(n28104), .A2(n27191), .ZN(n27192) );
  BUF_X4 U6716 ( .I(n19787), .Z(n19701) );
  NAND2_X1 U19386 ( .A1(n18937), .A2(n18936), .ZN(n26239) );
  CLKBUF_X2 U19344 ( .I(n30267), .Z(n22139) );
  NAND2_X1 U26434 ( .A1(n23772), .A2(n22139), .ZN(n29215) );
  INV_X2 U9713 ( .I(n21222), .ZN(n1318) );
  BUF_X2 U3874 ( .I(n22181), .Z(n17410) );
  CLKBUF_X1 U8278 ( .I(n26650), .Z(n58424) );
  BUF_X2 U5784 ( .I(n7580), .Z(n364) );
  BUF_X4 U8291 ( .I(n29028), .Z(n58999) );
  BUF_X2 U42063 ( .I(n28792), .Z(n22877) );
  INV_X2 U9719 ( .I(n16894), .ZN(n1319) );
  INV_X2 U3065 ( .I(n30183), .ZN(n21263) );
  INV_X2 U3160 ( .I(n25157), .ZN(n31059) );
  INV_X2 U3149 ( .I(n21512), .ZN(n30223) );
  INV_X2 U4915 ( .I(n13392), .ZN(n31098) );
  INV_X1 U3068 ( .I(n30347), .ZN(n30616) );
  INV_X1 U19362 ( .I(n25639), .ZN(n7026) );
  INV_X1 U11909 ( .I(n30722), .ZN(n1438) );
  INV_X1 U20382 ( .I(n29053), .ZN(n30252) );
  INV_X1 U33054 ( .I(n19059), .ZN(n30334) );
  BUF_X2 U14026 ( .I(n25349), .Z(n1561) );
  BUF_X2 U6214 ( .I(n16490), .Z(n57621) );
  CLKBUF_X2 U47561 ( .I(n28932), .Z(n61383) );
  INV_X1 U3135 ( .I(n30845), .ZN(n30216) );
  NAND3_X1 U38359 ( .A1(n27305), .A2(n25940), .A3(n25939), .ZN(n29411) );
  NOR2_X1 U2969 ( .A1(n30334), .A2(n23140), .ZN(n30332) );
  NOR2_X1 U4435 ( .A1(n30430), .A2(n31074), .ZN(n28571) );
  BUF_X2 U4565 ( .I(n30608), .Z(n40) );
  NAND3_X1 U26848 ( .A1(n31155), .A2(n31276), .A3(n31156), .ZN(n31267) );
  NOR2_X1 U3023 ( .A1(n30192), .A2(n2351), .ZN(n30184) );
  INV_X2 U24769 ( .I(n9411), .ZN(n9392) );
  NOR2_X1 U21114 ( .A1(n30441), .A2(n1253), .ZN(n19649) );
  NOR2_X1 U25232 ( .A1(n58651), .A2(n30547), .ZN(n27307) );
  NAND2_X1 U9667 ( .A1(n29241), .A2(n29835), .ZN(n29235) );
  INV_X2 U24279 ( .I(n18075), .ZN(n30124) );
  NAND3_X1 U3091 ( .A1(n29457), .A2(n18739), .A3(n18738), .ZN(n29846) );
  INV_X1 U19350 ( .I(n23140), .ZN(n8640) );
  INV_X2 U19381 ( .I(n21532), .ZN(n1869) );
  INV_X2 U37769 ( .I(n23705), .ZN(n22416) );
  NAND2_X1 U18499 ( .A1(n61531), .A2(n57537), .ZN(n30261) );
  BUF_X2 U8806 ( .I(n20809), .Z(n14399) );
  INV_X2 U33951 ( .I(n30781), .ZN(n30771) );
  INV_X2 U19293 ( .I(n24097), .ZN(n14063) );
  INV_X1 U6995 ( .I(n29860), .ZN(n12979) );
  INV_X2 U32905 ( .I(n31241), .ZN(n12893) );
  NOR2_X1 U44939 ( .A1(n10734), .A2(n26084), .ZN(n31115) );
  INV_X2 U32456 ( .I(n25349), .ZN(n23008) );
  INV_X2 U30236 ( .I(n31264), .ZN(n31279) );
  INV_X2 U27265 ( .I(n26438), .ZN(n29747) );
  INV_X2 U11908 ( .I(n23004), .ZN(n1437) );
  BUF_X2 U3131 ( .I(n29916), .Z(n9904) );
  NOR2_X1 U40115 ( .A1(n27516), .A2(n30267), .ZN(n30728) );
  INV_X2 U3064 ( .I(n29726), .ZN(n23315) );
  INV_X1 U3166 ( .I(n30609), .ZN(n29083) );
  NOR2_X1 U49155 ( .A1(n14230), .A2(n29993), .ZN(n29986) );
  INV_X2 U3129 ( .I(n10052), .ZN(n31277) );
  INV_X2 U9700 ( .I(n2005), .ZN(n2965) );
  INV_X1 U13950 ( .I(n31144), .ZN(n1843) );
  INV_X1 U3073 ( .I(n30267), .ZN(n30276) );
  INV_X1 U13989 ( .I(n22374), .ZN(n1862) );
  INV_X1 U31525 ( .I(n30413), .ZN(n30408) );
  INV_X1 U11888 ( .I(n29506), .ZN(n11106) );
  BUF_X2 U39760 ( .I(n23168), .Z(n60170) );
  NAND2_X1 U21868 ( .A1(n21222), .A2(n29801), .ZN(n30077) );
  INV_X1 U33433 ( .I(n1871), .ZN(n1556) );
  NAND3_X1 U19281 ( .A1(n30276), .A2(n9426), .A3(n23317), .ZN(n30279) );
  INV_X2 U3844 ( .I(n12112), .ZN(n57953) );
  BUF_X2 U6212 ( .I(n31254), .Z(n58395) );
  NAND2_X1 U24491 ( .A1(n19118), .A2(n31277), .ZN(n31262) );
  INV_X1 U4447 ( .I(n3993), .ZN(n6088) );
  INV_X2 U11823 ( .I(n1351), .ZN(n9618) );
  NAND2_X1 U8631 ( .A1(n29787), .A2(n14063), .ZN(n14062) );
  NOR3_X1 U15583 ( .A1(n30048), .A2(n2269), .A3(n30261), .ZN(n29055) );
  NAND3_X1 U20345 ( .A1(n22799), .A2(n30183), .A3(n2177), .ZN(n29045) );
  AOI21_X1 U31373 ( .A1(n1436), .A2(n1435), .B(n5933), .ZN(n30497) );
  OAI21_X1 U13958 ( .A1(n30396), .A2(n22742), .B(n4270), .ZN(n11104) );
  NOR3_X1 U44789 ( .A1(n14063), .A2(n58486), .A3(n29779), .ZN(n27788) );
  NAND2_X1 U11813 ( .A1(n2795), .A2(n29511), .ZN(n29503) );
  INV_X1 U3786 ( .I(n23269), .ZN(n59755) );
  INV_X1 U39552 ( .I(n30728), .ZN(n29036) );
  NAND2_X1 U38707 ( .A1(n26429), .A2(n1319), .ZN(n26441) );
  INV_X4 U7007 ( .I(n1253), .ZN(n30537) );
  NAND2_X1 U30345 ( .A1(n8182), .A2(n30870), .ZN(n31275) );
  NAND2_X1 U39767 ( .A1(n15727), .A2(n18306), .ZN(n18322) );
  NOR2_X1 U38388 ( .A1(n27763), .A2(n25527), .ZN(n60000) );
  INV_X2 U3036 ( .I(n30538), .ZN(n1434) );
  NOR2_X1 U36857 ( .A1(n29506), .A2(n10068), .ZN(n27634) );
  NAND2_X1 U3027 ( .A1(n23317), .A2(n29220), .ZN(n29224) );
  INV_X1 U5105 ( .I(n24987), .ZN(n13417) );
  INV_X1 U13987 ( .I(n20809), .ZN(n29453) );
  NOR2_X1 U24811 ( .A1(n31264), .A2(n6317), .ZN(n31271) );
  NAND2_X1 U2995 ( .A1(n31074), .A2(n30419), .ZN(n31079) );
  NAND2_X1 U3088 ( .A1(n5070), .A2(n24728), .ZN(n29813) );
  BUF_X2 U19310 ( .I(n24298), .Z(n16694) );
  NAND2_X1 U39289 ( .A1(n29862), .A2(n29860), .ZN(n29514) );
  BUF_X2 U42520 ( .I(n30547), .Z(n23478) );
  BUF_X2 U4537 ( .I(n30781), .Z(n21886) );
  NAND2_X1 U40309 ( .A1(n31255), .A2(n30891), .ZN(n29886) );
  INV_X1 U13840 ( .I(n28688), .ZN(n7594) );
  NOR2_X1 U42803 ( .A1(n31059), .A2(n31051), .ZN(n31053) );
  BUF_X2 U3787 ( .I(n2005), .Z(n59481) );
  NAND2_X1 U28143 ( .A1(n24949), .A2(n23502), .ZN(n6709) );
  NAND2_X1 U6103 ( .A1(n8097), .A2(n29083), .ZN(n29591) );
  NOR2_X1 U44790 ( .A1(n28943), .A2(n29779), .ZN(n27790) );
  INV_X1 U8697 ( .I(n22555), .ZN(n30618) );
  NAND2_X1 U34183 ( .A1(n23053), .A2(n30538), .ZN(n14739) );
  AOI21_X1 U5284 ( .A1(n12907), .A2(n23056), .B(n16279), .ZN(n31029) );
  INV_X4 U10489 ( .I(n30786), .ZN(n20179) );
  INV_X1 U25979 ( .I(n31270), .ZN(n25989) );
  NOR2_X1 U23739 ( .A1(n23955), .A2(n31098), .ZN(n31110) );
  INV_X1 U19239 ( .I(n13411), .ZN(n10140) );
  NOR2_X1 U9663 ( .A1(n58560), .A2(n23315), .ZN(n30025) );
  NOR2_X1 U4785 ( .A1(n22878), .A2(n5267), .ZN(n29474) );
  NOR2_X1 U44213 ( .A1(n64565), .A2(n29860), .ZN(n29855) );
  NAND2_X1 U3752 ( .A1(n11092), .A2(n23140), .ZN(n17903) );
  INV_X1 U39207 ( .I(n29397), .ZN(n30496) );
  INV_X1 U32686 ( .I(n29910), .ZN(n59451) );
  INV_X1 U37684 ( .I(n21832), .ZN(n29579) );
  INV_X1 U3083 ( .I(n26084), .ZN(n10427) );
  OR2_X1 U4514 ( .A1(n1866), .A2(n16491), .Z(n29568) );
  NAND2_X1 U2959 ( .A1(n9426), .A2(n1438), .ZN(n29221) );
  INV_X2 U2981 ( .I(n15738), .ZN(n1875) );
  NOR2_X1 U31372 ( .A1(n1436), .A2(n1435), .ZN(n30884) );
  CLKBUF_X2 U27358 ( .I(n1433), .Z(n58816) );
  NAND2_X1 U9661 ( .A1(n22496), .A2(n12112), .ZN(n15136) );
  CLKBUF_X2 U3863 ( .I(n19118), .Z(n327) );
  NAND2_X1 U28174 ( .A1(n8097), .A2(n59268), .ZN(n29594) );
  NAND2_X1 U28175 ( .A1(n8097), .A2(n30608), .ZN(n30342) );
  NAND2_X1 U10506 ( .A1(n15738), .A2(n30664), .ZN(n30013) );
  AOI21_X1 U38407 ( .A1(n30724), .A2(n14389), .B(n30275), .ZN(n17338) );
  INV_X1 U36862 ( .I(n30659), .ZN(n30330) );
  OAI21_X1 U19048 ( .A1(n2042), .A2(n58395), .B(n30496), .ZN(n30499) );
  NAND3_X1 U21708 ( .A1(n30654), .A2(n17903), .A3(n8770), .ZN(n30329) );
  NOR2_X1 U46221 ( .A1(n31267), .A2(n25013), .ZN(n31266) );
  OAI21_X1 U53759 ( .A1(n29778), .A2(n7943), .B(n61175), .ZN(n3794) );
  AOI21_X1 U8748 ( .A1(n25384), .A2(n31083), .B(n22411), .ZN(n31088) );
  NOR2_X1 U3098 ( .A1(n30343), .A2(n30614), .ZN(n29592) );
  NOR2_X1 U2990 ( .A1(n31098), .A2(n1868), .ZN(n28209) );
  NAND3_X1 U39965 ( .A1(n162), .A2(n58816), .A3(n10820), .ZN(n30811) );
  NAND2_X1 U3800 ( .A1(n16808), .A2(n30216), .ZN(n29195) );
  NAND2_X1 U8951 ( .A1(n27759), .A2(n1352), .ZN(n28905) );
  NAND2_X1 U3766 ( .A1(n11195), .A2(n29045), .ZN(n57558) );
  NAND2_X1 U19076 ( .A1(n23502), .A2(n6088), .ZN(n6087) );
  NOR2_X1 U18490 ( .A1(n24196), .A2(n30844), .ZN(n29194) );
  NAND2_X1 U8782 ( .A1(n30351), .A2(n30343), .ZN(n29088) );
  NAND2_X1 U21180 ( .A1(n60202), .A2(n63537), .ZN(n27990) );
  NAND2_X1 U8950 ( .A1(n13144), .A2(n23140), .ZN(n13145) );
  INV_X1 U19198 ( .I(n7774), .ZN(n29999) );
  INV_X2 U37742 ( .I(n29512), .ZN(n30954) );
  INV_X1 U37880 ( .I(n31092), .ZN(n19572) );
  NAND2_X1 U16345 ( .A1(n24777), .A2(n31187), .ZN(n57676) );
  NAND2_X1 U44158 ( .A1(n30799), .A2(n10820), .ZN(n30807) );
  NAND2_X1 U26984 ( .A1(n1838), .A2(n29099), .ZN(n29524) );
  NAND2_X1 U44850 ( .A1(n1351), .A2(n30124), .ZN(n27923) );
  NAND2_X1 U2931 ( .A1(n14230), .A2(n29988), .ZN(n30321) );
  NAND2_X1 U45625 ( .A1(n21176), .A2(n30702), .ZN(n31031) );
  OAI21_X1 U19023 ( .A1(n20009), .A2(n30285), .B(n8685), .ZN(n23064) );
  NAND4_X1 U45023 ( .A1(n61629), .A2(n28574), .A3(n25384), .A4(n60895), .ZN(
        n28575) );
  NAND2_X1 U8909 ( .A1(n29052), .A2(n61622), .ZN(n2843) );
  INV_X1 U22934 ( .I(n4210), .ZN(n30018) );
  AOI21_X1 U23980 ( .A1(n30280), .A2(n30279), .B(n30278), .ZN(n30281) );
  CLKBUF_X2 U10482 ( .I(n1863), .Z(n10431) );
  NAND2_X1 U19228 ( .A1(n60142), .A2(n30696), .ZN(n30160) );
  NAND3_X1 U21416 ( .A1(n30781), .A2(n26441), .A3(n2965), .ZN(n17281) );
  NAND2_X1 U11837 ( .A1(n13360), .A2(n30344), .ZN(n13361) );
  NAND2_X1 U4259 ( .A1(n18306), .A2(n16971), .ZN(n29422) );
  NOR2_X1 U34789 ( .A1(n3180), .A2(n16907), .ZN(n29505) );
  NAND2_X1 U45785 ( .A1(n19118), .A2(n6316), .ZN(n30509) );
  NAND2_X1 U42579 ( .A1(n29935), .A2(n8521), .ZN(n29936) );
  NOR2_X1 U45214 ( .A1(n60162), .A2(n21095), .ZN(n30362) );
  NOR2_X1 U7019 ( .A1(n12632), .A2(n29455), .ZN(n29842) );
  NOR2_X1 U37572 ( .A1(n31254), .A2(n31247), .ZN(n30890) );
  NOR2_X1 U45357 ( .A1(n24504), .A2(n61382), .ZN(n30422) );
  INV_X1 U5380 ( .I(n58931), .ZN(n30560) );
  INV_X1 U10452 ( .I(n30410), .ZN(n30641) );
  INV_X1 U14003 ( .I(n29787), .ZN(n14064) );
  INV_X1 U10488 ( .I(n30225), .ZN(n1350) );
  NOR2_X1 U36782 ( .A1(n28986), .A2(n21478), .ZN(n30020) );
  NOR2_X1 U2987 ( .A1(n30374), .A2(n5768), .ZN(n30593) );
  NOR2_X1 U4786 ( .A1(n5267), .A2(n18060), .ZN(n30551) );
  INV_X1 U3067 ( .I(n23708), .ZN(n1852) );
  NOR2_X1 U33908 ( .A1(n20809), .A2(n29452), .ZN(n29844) );
  NOR2_X1 U40832 ( .A1(n11987), .A2(n28899), .ZN(n30479) );
  NAND2_X1 U8839 ( .A1(n59046), .A2(n30752), .ZN(n31218) );
  INV_X1 U11832 ( .I(n28902), .ZN(n30478) );
  INV_X1 U2938 ( .I(n3052), .ZN(n28092) );
  INV_X1 U11862 ( .I(n29900), .ZN(n30854) );
  NAND3_X1 U45782 ( .A1(n31253), .A2(n5933), .A3(n58395), .ZN(n30504) );
  INV_X1 U45855 ( .I(n30654), .ZN(n30657) );
  NAND2_X1 U8758 ( .A1(n29987), .A2(n10345), .ZN(n29990) );
  NAND3_X1 U34854 ( .A1(n18867), .A2(n29824), .A3(n29988), .ZN(n30326) );
  NOR2_X1 U45084 ( .A1(n17413), .A2(n17414), .ZN(n29856) );
  OAI22_X1 U45467 ( .A1(n2636), .A2(n30054), .B1(n22014), .B2(n8602), .ZN(
        n29757) );
  NAND3_X1 U44906 ( .A1(n29844), .A2(n23224), .A3(n29842), .ZN(n28118) );
  NOR3_X1 U23442 ( .A1(n30391), .A2(n30396), .A3(n2795), .ZN(n4497) );
  NAND4_X1 U8947 ( .A1(n12112), .A2(n30680), .A3(n19461), .A4(n30239), .ZN(
        n14390) );
  NAND2_X1 U9633 ( .A1(n30890), .A2(n30883), .ZN(n31260) );
  AOI22_X1 U3520 ( .A1(n30578), .A2(n31114), .B1(n4993), .B2(n30577), .ZN(
        n19396) );
  NAND2_X1 U10424 ( .A1(n30685), .A2(n30239), .ZN(n29206) );
  NAND2_X1 U8915 ( .A1(n16147), .A2(n64894), .ZN(n3814) );
  AOI22_X1 U42684 ( .A1(n29091), .A2(n64940), .B1(n29090), .B2(n64565), .ZN(
        n29095) );
  NAND2_X1 U45119 ( .A1(n30680), .A2(n10525), .ZN(n28777) );
  NOR2_X1 U45261 ( .A1(n30225), .A2(n30841), .ZN(n29197) );
  NAND2_X1 U10423 ( .A1(n30759), .A2(n30750), .ZN(n30766) );
  INV_X1 U19151 ( .I(n17281), .ZN(n29552) );
  NOR2_X1 U33282 ( .A1(n17084), .A2(n30517), .ZN(n20151) );
  NAND2_X1 U38671 ( .A1(n31136), .A2(n8584), .ZN(n17792) );
  AOI21_X1 U9641 ( .A1(n30519), .A2(n30523), .B(n30518), .ZN(n20273) );
  NAND4_X1 U45857 ( .A1(n30659), .A2(n30658), .A3(n30657), .A4(n30656), .ZN(
        n30660) );
  AOI21_X1 U19020 ( .A1(n13119), .A2(n28938), .B(n58710), .ZN(n15531) );
  NAND3_X1 U23573 ( .A1(n31217), .A2(n30762), .A3(n31224), .ZN(n17506) );
  NAND2_X1 U39771 ( .A1(n30215), .A2(n16808), .ZN(n19431) );
  NAND2_X1 U34172 ( .A1(n24299), .A2(n58651), .ZN(n30541) );
  NOR2_X1 U38005 ( .A1(n29516), .A2(n30954), .ZN(n18763) );
  NOR2_X1 U13855 ( .A1(n27923), .A2(n29766), .ZN(n30520) );
  INV_X1 U17662 ( .I(n30141), .ZN(n57772) );
  NAND2_X1 U11878 ( .A1(n29905), .A2(n1353), .ZN(n27906) );
  NAND3_X1 U19195 ( .A1(n24777), .A2(n29900), .A3(n1431), .ZN(n13448) );
  INV_X1 U45893 ( .I(n30784), .ZN(n30791) );
  NOR2_X1 U39279 ( .A1(n28750), .A2(n18716), .ZN(n23159) );
  INV_X1 U5601 ( .I(n20364), .ZN(n1552) );
  NAND2_X1 U39179 ( .A1(n17590), .A2(n57937), .ZN(n27902) );
  INV_X1 U20117 ( .I(n28782), .ZN(n6038) );
  NOR2_X1 U25795 ( .A1(n3167), .A2(n13629), .ZN(n58704) );
  NAND3_X1 U22488 ( .A1(n29979), .A2(n29978), .A3(n8476), .ZN(n3818) );
  NAND3_X1 U10433 ( .A1(n30481), .A2(n61162), .A3(n30482), .ZN(n30483) );
  BUF_X2 U45520 ( .I(n63396), .Z(n55833) );
  NAND2_X1 U42582 ( .A1(n1852), .A2(n30430), .ZN(n30559) );
  NAND2_X1 U27797 ( .A1(n31127), .A2(n6041), .ZN(n31131) );
  NOR2_X1 U21700 ( .A1(n13145), .A2(n30409), .ZN(n30647) );
  BUF_X2 U19879 ( .I(n19171), .Z(n55379) );
  NAND3_X1 U35906 ( .A1(n30193), .A2(n30183), .A3(n5631), .ZN(n30200) );
  NAND2_X1 U13882 ( .A1(n28695), .A2(n16026), .ZN(n8424) );
  OR2_X1 U8938 ( .A1(n21176), .A2(n16279), .Z(n57392) );
  INV_X1 U21443 ( .I(n2996), .ZN(n29441) );
  INV_X1 U11790 ( .I(n30364), .ZN(n30456) );
  NAND3_X1 U13926 ( .A1(n29900), .A2(n1431), .A3(n29905), .ZN(n13447) );
  NOR3_X1 U45862 ( .A1(n18198), .A2(n10525), .A3(n30679), .ZN(n30675) );
  OAI21_X1 U23589 ( .A1(n13594), .A2(n16694), .B(n8476), .ZN(n13593) );
  NAND3_X1 U19032 ( .A1(n31260), .A2(n31252), .A3(n31259), .ZN(n11876) );
  NOR4_X1 U30836 ( .A1(n30062), .A2(n59214), .A3(n31061), .A4(n30061), .ZN(
        n30068) );
  INV_X1 U8983 ( .I(n6720), .ZN(n30822) );
  AOI21_X1 U54802 ( .A1(n30508), .A2(n30511), .B(n29921), .ZN(n29922) );
  NOR3_X1 U44842 ( .A1(n1431), .A2(n27907), .A3(n29896), .ZN(n27908) );
  OAI21_X1 U34174 ( .A1(n30540), .A2(n58651), .B(n23478), .ZN(n30543) );
  AOI22_X1 U5020 ( .A1(n31099), .A2(n65), .B1(n31101), .B2(n14276), .ZN(n10733) );
  NAND2_X1 U28450 ( .A1(n31217), .A2(n8364), .ZN(n25121) );
  AOI21_X1 U13957 ( .A1(n30319), .A2(n29820), .B(n29993), .ZN(n29273) );
  NAND4_X1 U38469 ( .A1(n10068), .A2(n30392), .A3(n30396), .A4(n24949), .ZN(
        n26586) );
  NAND4_X1 U45200 ( .A1(n29018), .A2(n64589), .A3(n29797), .A4(n29017), .ZN(
        n29020) );
  NOR2_X1 U5762 ( .A1(n25960), .A2(n14423), .ZN(n5076) );
  AOI21_X1 U9651 ( .A1(n28950), .A2(n28949), .B(n29244), .ZN(n14050) );
  INV_X1 U45939 ( .I(n30858), .ZN(n30859) );
  NAND2_X1 U35470 ( .A1(n29236), .A2(n18905), .ZN(n18904) );
  NAND3_X1 U8443 ( .A1(n20682), .A2(n29402), .A3(n29401), .ZN(n1989) );
  NAND2_X1 U25786 ( .A1(n58704), .A2(n3169), .ZN(n18637) );
  NOR2_X1 U26211 ( .A1(n30253), .A2(n61892), .ZN(n6547) );
  OAI21_X1 U2903 ( .A1(n5863), .A2(n5862), .B(n5861), .ZN(n28908) );
  NAND2_X1 U31727 ( .A1(n16971), .A2(n11425), .ZN(n28291) );
  NAND2_X1 U2871 ( .A1(n25185), .A2(n25183), .ZN(n12897) );
  NAND2_X1 U8745 ( .A1(n17631), .A2(n30749), .ZN(n30672) );
  NOR3_X1 U36852 ( .A1(n58502), .A2(n28291), .A3(n18402), .ZN(n28293) );
  AOI22_X1 U36957 ( .A1(n30325), .A2(n30324), .B1(n30323), .B2(n16026), .ZN(
        n30328) );
  AOI21_X1 U56503 ( .A1(n61386), .A2(n31083), .B(n61385), .ZN(n61384) );
  AOI21_X1 U19132 ( .A1(n27628), .A2(n27627), .B(n29255), .ZN(n12561) );
  NOR3_X1 U26149 ( .A1(n5425), .A2(n21657), .A3(n5421), .ZN(n58764) );
  NAND3_X1 U20328 ( .A1(n27425), .A2(n30047), .A3(n2267), .ZN(n27426) );
  NOR3_X1 U36952 ( .A1(n30081), .A2(n30080), .A3(n30079), .ZN(n30092) );
  NOR2_X1 U30616 ( .A1(n12060), .A2(n59169), .ZN(n6228) );
  NOR2_X1 U26231 ( .A1(n6584), .A2(n30397), .ZN(n30399) );
  CLKBUF_X2 U18916 ( .I(n30907), .Z(n18248) );
  INV_X1 U18917 ( .I(n33239), .ZN(n17546) );
  NOR2_X1 U28205 ( .A1(n21414), .A2(n16161), .ZN(n21228) );
  NAND2_X1 U8897 ( .A1(n28929), .A2(n20731), .ZN(n21885) );
  NOR4_X1 U2854 ( .A1(n12898), .A2(n14050), .A3(n13842), .A4(n12897), .ZN(
        n12896) );
  NAND2_X1 U8149 ( .A1(n21796), .A2(n21795), .ZN(n2373) );
  NOR4_X1 U39610 ( .A1(n29828), .A2(n29829), .A3(n29827), .A4(n29826), .ZN(
        n29830) );
  INV_X1 U13756 ( .I(n24869), .ZN(n4640) );
  INV_X1 U33703 ( .I(n19863), .ZN(n59933) );
  NAND2_X1 U5707 ( .A1(n19993), .A2(n7615), .ZN(n7617) );
  NAND2_X1 U3648 ( .A1(n58591), .A2(n31439), .ZN(n10013) );
  NAND3_X1 U2847 ( .A1(n25631), .A2(n23679), .A3(n25630), .ZN(n15732) );
  NAND4_X1 U18985 ( .A1(n31573), .A2(n31572), .A3(n31571), .A4(n31570), .ZN(
        n31576) );
  NAND2_X1 U20656 ( .A1(n24327), .A2(n5741), .ZN(n31863) );
  INV_X1 U3631 ( .I(n53764), .ZN(n1573) );
  NAND2_X1 U37689 ( .A1(n25027), .A2(n28897), .ZN(n33139) );
  INV_X1 U19056 ( .I(n20316), .ZN(n26845) );
  INV_X1 U28417 ( .I(n26038), .ZN(n26039) );
  INV_X1 U33869 ( .I(n30985), .ZN(n32382) );
  BUF_X2 U44349 ( .I(n8810), .Z(n60717) );
  BUF_X2 U3636 ( .I(n32324), .Z(n9283) );
  INV_X1 U11725 ( .I(n6544), .ZN(n7949) );
  BUF_X2 U2843 ( .I(n12414), .Z(n9055) );
  BUF_X2 U42686 ( .I(n32317), .Z(n23726) );
  BUF_X2 U5702 ( .I(n30921), .Z(n15464) );
  BUF_X2 U2845 ( .I(n15511), .Z(n15510) );
  INV_X2 U42210 ( .I(n31433), .ZN(n32617) );
  INV_X1 U2818 ( .I(n22674), .ZN(n23950) );
  INV_X1 U32996 ( .I(n839), .ZN(n13045) );
  INV_X1 U35428 ( .I(n31912), .ZN(n32181) );
  INV_X1 U38763 ( .I(n21503), .ZN(n31849) );
  INV_X1 U2850 ( .I(n31341), .ZN(n30897) );
  INV_X1 U18883 ( .I(n22476), .ZN(n1830) );
  BUF_X2 U3624 ( .I(n22296), .Z(n10553) );
  INV_X1 U10399 ( .I(n12414), .ZN(n31753) );
  CLKBUF_X1 U10392 ( .I(n24471), .Z(n19348) );
  INV_X1 U39687 ( .I(n1826), .ZN(n25203) );
  INV_X1 U26489 ( .I(n23152), .ZN(n8492) );
  BUF_X2 U2805 ( .I(n16958), .Z(n5436) );
  BUF_X2 U2820 ( .I(n32383), .Z(n23714) );
  INV_X1 U34862 ( .I(n33173), .ZN(n17616) );
  INV_X1 U6077 ( .I(n21172), .ZN(n33829) );
  INV_X1 U2812 ( .I(n32585), .ZN(n22769) );
  BUF_X2 U2806 ( .I(n31193), .Z(n25887) );
  BUF_X2 U32159 ( .I(n32733), .Z(n12022) );
  INV_X1 U20403 ( .I(n57405), .ZN(n13486) );
  INV_X1 U7033 ( .I(n5489), .ZN(n20617) );
  INV_X2 U25039 ( .I(n9883), .ZN(n5342) );
  INV_X1 U33155 ( .I(n14218), .ZN(n21586) );
  INV_X2 U9226 ( .I(n21586), .ZN(n1549) );
  INV_X1 U9165 ( .I(n30735), .ZN(n16952) );
  INV_X1 U3618 ( .I(n32207), .ZN(n18838) );
  INV_X1 U9183 ( .I(n18156), .ZN(n25843) );
  INV_X1 U18817 ( .I(n30400), .ZN(n1819) );
  INV_X1 U3884 ( .I(n6885), .ZN(n31749) );
  INV_X1 U56893 ( .I(n5147), .ZN(n34586) );
  INV_X2 U6438 ( .I(n33662), .ZN(n32695) );
  INV_X2 U28222 ( .I(n8146), .ZN(n34268) );
  INV_X2 U46985 ( .I(n32017), .ZN(n34752) );
  INV_X1 U9240 ( .I(n32497), .ZN(n15393) );
  INV_X1 U21431 ( .I(n2974), .ZN(n5412) );
  CLKBUF_X2 U9320 ( .I(n13487), .Z(n58048) );
  BUF_X2 U41880 ( .I(n34317), .Z(n22633) );
  INV_X2 U41576 ( .I(n13559), .ZN(n34798) );
  INV_X2 U2766 ( .I(n63586), .ZN(n1342) );
  INV_X2 U32535 ( .I(n1817), .ZN(n35748) );
  BUF_X2 U11703 ( .I(n15552), .Z(n2208) );
  INV_X2 U24734 ( .I(n4880), .ZN(n6304) );
  BUF_X2 U5802 ( .I(n33662), .Z(n10251) );
  INV_X2 U18747 ( .I(n34127), .ZN(n1812) );
  INV_X1 U18751 ( .I(n2271), .ZN(n2323) );
  INV_X1 U2743 ( .I(n32828), .ZN(n32834) );
  INV_X1 U42457 ( .I(n31905), .ZN(n25372) );
  INV_X1 U11719 ( .I(n24965), .ZN(n1427) );
  INV_X1 U2763 ( .I(n14080), .ZN(n1428) );
  INV_X1 U24596 ( .I(n33972), .ZN(n32875) );
  INV_X1 U8887 ( .I(n32409), .ZN(n34727) );
  INV_X1 U18748 ( .I(n61749), .ZN(n3148) );
  INV_X1 U5364 ( .I(n33519), .ZN(n34018) );
  OR2_X1 U25690 ( .A1(n13559), .A2(n13781), .Z(n60883) );
  INV_X2 U22107 ( .I(n11359), .ZN(n7517) );
  INV_X2 U11702 ( .I(n5082), .ZN(n33622) );
  NAND2_X1 U3871 ( .A1(n12582), .A2(n57590), .ZN(n34998) );
  INV_X1 U2773 ( .I(n35031), .ZN(n1814) );
  BUF_X4 U31049 ( .I(n18651), .Z(n61496) );
  NAND2_X1 U35222 ( .A1(n15740), .A2(n13583), .ZN(n35215) );
  CLKBUF_X2 U54842 ( .I(n2891), .Z(n61249) );
  NOR2_X1 U30171 ( .A1(n24093), .A2(n33540), .ZN(n33372) );
  NOR2_X1 U29116 ( .A1(n25657), .A2(n34632), .ZN(n35037) );
  INV_X2 U31386 ( .I(n24256), .ZN(n33993) );
  NOR2_X1 U7597 ( .A1(n35027), .A2(n1427), .ZN(n902) );
  INV_X2 U21244 ( .I(n19005), .ZN(n34761) );
  NAND2_X1 U29979 ( .A1(n15809), .A2(n23945), .ZN(n34594) );
  INV_X2 U7575 ( .I(n25657), .ZN(n9130) );
  INV_X1 U9285 ( .I(n23354), .ZN(n34747) );
  INV_X2 U7579 ( .I(n20865), .ZN(n35731) );
  INV_X1 U38327 ( .I(n60883), .ZN(n34791) );
  BUF_X2 U13423 ( .I(n32489), .Z(n33561) );
  CLKBUF_X2 U34518 ( .I(n2618), .Z(n61256) );
  INV_X1 U25112 ( .I(n5411), .ZN(n14703) );
  INV_X2 U22328 ( .I(n35738), .ZN(n35743) );
  INV_X1 U27316 ( .I(n6304), .ZN(n3549) );
  NOR2_X1 U21042 ( .A1(n33465), .A2(n2721), .ZN(n34787) );
  INV_X1 U4892 ( .I(n24083), .ZN(n34056) );
  CLKBUF_X2 U27510 ( .I(n32409), .Z(n34719) );
  INV_X1 U2687 ( .I(n15740), .ZN(n24614) );
  NOR2_X1 U2718 ( .A1(n35305), .A2(n16347), .ZN(n24488) );
  INV_X1 U38078 ( .I(n5322), .ZN(n61262) );
  INV_X1 U2689 ( .I(n16402), .ZN(n35764) );
  NAND2_X1 U2711 ( .A1(n64387), .A2(n16451), .ZN(n34275) );
  INV_X1 U4956 ( .I(n22316), .ZN(n34980) );
  NAND2_X1 U32390 ( .A1(n1545), .A2(n22185), .ZN(n12354) );
  INV_X1 U18696 ( .I(n2208), .ZN(n2207) );
  INV_X2 U5062 ( .I(n34973), .ZN(n25404) );
  INV_X1 U23623 ( .I(n4565), .ZN(n33098) );
  INV_X1 U11690 ( .I(n35750), .ZN(n12248) );
  INV_X1 U38126 ( .I(n16857), .ZN(n32512) );
  AND2_X1 U2729 ( .A1(n227), .A2(n9118), .Z(n33614) );
  INV_X1 U2630 ( .I(n10358), .ZN(n34587) );
  OAI21_X1 U2757 ( .A1(n25509), .A2(n5082), .B(n8997), .ZN(n5083) );
  INV_X2 U2696 ( .I(n34972), .ZN(n33730) );
  CLKBUF_X2 U18769 ( .I(n15740), .Z(n24006) );
  INV_X2 U18698 ( .I(n23470), .ZN(n34766) );
  INV_X1 U2612 ( .I(n15783), .ZN(n32795) );
  INV_X1 U2549 ( .I(n21252), .ZN(n35220) );
  NAND3_X1 U47938 ( .A1(n33651), .A2(n34137), .A3(n33650), .ZN(n33653) );
  INV_X2 U20636 ( .I(n34221), .ZN(n20736) );
  OAI22_X1 U38456 ( .A1(n34587), .A2(n34188), .B1(n23223), .B2(n59522), .ZN(
        n32878) );
  NAND2_X1 U22578 ( .A1(n35235), .A2(n7710), .ZN(n35708) );
  NOR2_X1 U26697 ( .A1(n32831), .A2(n17866), .ZN(n7017) );
  NAND2_X1 U47964 ( .A1(n63581), .A2(n34353), .ZN(n33738) );
  NAND2_X1 U16708 ( .A1(n18884), .A2(n33660), .ZN(n33396) );
  NAND2_X1 U18579 ( .A1(n35325), .A2(n11659), .ZN(n35326) );
  INV_X1 U38127 ( .I(n32512), .ZN(n33103) );
  NAND2_X1 U38761 ( .A1(n23127), .A2(n32782), .ZN(n22284) );
  INV_X1 U27695 ( .I(n6206), .ZN(n35287) );
  CLKBUF_X2 U6167 ( .I(n32846), .Z(n59626) );
  BUF_X2 U11674 ( .I(n9203), .Z(n4851) );
  NAND2_X1 U31162 ( .A1(n65119), .A2(n60960), .ZN(n59245) );
  NOR2_X1 U13600 ( .A1(n12248), .A2(n60175), .ZN(n35195) );
  INV_X1 U2604 ( .I(n15809), .ZN(n34589) );
  AOI21_X1 U36394 ( .A1(n34306), .A2(n60416), .B(n34309), .ZN(n34213) );
  CLKBUF_X1 U32558 ( .I(n34566), .Z(n59432) );
  BUF_X2 U11684 ( .I(n4189), .Z(n2322) );
  NOR2_X1 U2697 ( .A1(n9205), .A2(n1542), .ZN(n33408) );
  NOR2_X1 U2706 ( .A1(n31842), .A2(n35805), .ZN(n35803) );
  NAND2_X1 U22313 ( .A1(n7883), .A2(n34973), .ZN(n34971) );
  INV_X2 U34522 ( .I(n33763), .ZN(n24799) );
  NOR2_X1 U21780 ( .A1(n2617), .A2(n19894), .ZN(n25216) );
  NAND2_X1 U31756 ( .A1(n35743), .A2(n34415), .ZN(n1541) );
  NAND2_X1 U25552 ( .A1(n5903), .A2(n9130), .ZN(n31298) );
  NOR2_X1 U2623 ( .A1(n34309), .A2(n34761), .ZN(n34208) );
  INV_X1 U2618 ( .I(n14464), .ZN(n34948) );
  INV_X2 U11697 ( .I(n34956), .ZN(n1537) );
  NAND2_X1 U48162 ( .A1(n34316), .A2(n22633), .ZN(n34713) );
  NAND2_X1 U9243 ( .A1(n6979), .A2(n24006), .ZN(n18380) );
  INV_X1 U5130 ( .I(n32869), .ZN(n1809) );
  INV_X1 U9586 ( .I(n34185), .ZN(n34583) );
  BUF_X2 U6157 ( .I(n35031), .Z(n60984) );
  INV_X1 U32269 ( .I(n34958), .ZN(n22342) );
  NOR2_X1 U43495 ( .A1(n32892), .A2(n32834), .ZN(n34201) );
  INV_X1 U11709 ( .I(n33464), .ZN(n23645) );
  INV_X1 U2692 ( .I(n34708), .ZN(n35817) );
  INV_X1 U43855 ( .I(n34193), .ZN(n60684) );
  INV_X1 U34755 ( .I(n61196), .ZN(n33362) );
  INV_X1 U36380 ( .I(n33944), .ZN(n32862) );
  INV_X1 U4231 ( .I(n22797), .ZN(n18199) );
  INV_X1 U2660 ( .I(n34725), .ZN(n34246) );
  NOR2_X1 U4797 ( .A1(n34594), .A2(n23223), .ZN(n11403) );
  INV_X1 U8851 ( .I(n3325), .ZN(n33767) );
  INV_X2 U16816 ( .I(n32436), .ZN(n1804) );
  NOR2_X1 U34301 ( .A1(n34658), .A2(n5410), .ZN(n14913) );
  NAND2_X1 U21779 ( .A1(n18884), .A2(n262), .ZN(n32700) );
  INV_X1 U10372 ( .I(n25999), .ZN(n34643) );
  NOR2_X1 U34452 ( .A1(n15148), .A2(n10566), .ZN(n35701) );
  INV_X1 U3546 ( .I(n6033), .ZN(n33354) );
  NOR2_X1 U48076 ( .A1(n34080), .A2(n61078), .ZN(n33957) );
  INV_X1 U13682 ( .I(n35198), .ZN(n35619) );
  OAI21_X1 U42632 ( .A1(n23645), .A2(n23644), .B(n24799), .ZN(n32361) );
  NAND2_X1 U13540 ( .A1(n2899), .A2(n35735), .ZN(n4641) );
  NOR2_X1 U23571 ( .A1(n34535), .A2(n34971), .ZN(n32917) );
  NAND2_X1 U31094 ( .A1(n18394), .A2(n35315), .ZN(n11670) );
  INV_X1 U27607 ( .I(n34639), .ZN(n34647) );
  NAND2_X1 U33725 ( .A1(n65119), .A2(n23761), .ZN(n14147) );
  NAND2_X1 U47913 ( .A1(n35670), .A2(n17401), .ZN(n33577) );
  NOR2_X1 U38503 ( .A1(n35806), .A2(n10337), .ZN(n17498) );
  NAND2_X1 U21950 ( .A1(n57898), .A2(n65232), .ZN(n59397) );
  OAI21_X1 U16191 ( .A1(n23223), .A2(n20607), .B(n57669), .ZN(n15099) );
  NAND2_X1 U6139 ( .A1(n19663), .A2(n34132), .ZN(n59347) );
  NAND2_X1 U48559 ( .A1(n32684), .A2(n19373), .ZN(n35617) );
  NAND3_X1 U56406 ( .A1(n10448), .A2(n61458), .A3(n34385), .ZN(n35276) );
  NAND2_X1 U31881 ( .A1(n21751), .A2(n34335), .ZN(n34741) );
  NAND3_X1 U8277 ( .A1(n63103), .A2(n33624), .A3(n59125), .ZN(n33632) );
  NOR2_X1 U3574 ( .A1(n11247), .A2(n33509), .ZN(n33506) );
  NAND3_X1 U23483 ( .A1(n35300), .A2(n31976), .A3(n20105), .ZN(n59319) );
  NAND2_X1 U11646 ( .A1(n12338), .A2(n21906), .ZN(n3746) );
  NAND2_X1 U20321 ( .A1(n35799), .A2(n11182), .ZN(n34382) );
  NAND3_X1 U2559 ( .A1(n1804), .A2(n34305), .A3(n34306), .ZN(n32948) );
  NAND3_X1 U22053 ( .A1(n34138), .A2(n33390), .A3(n19663), .ZN(n34135) );
  NAND2_X1 U9281 ( .A1(n10750), .A2(n24737), .ZN(n33956) );
  NAND4_X1 U2576 ( .A1(n10448), .A2(n35802), .A3(n11182), .A4(n35799), .ZN(
        n34384) );
  CLKBUF_X2 U25557 ( .I(n60054), .Z(n58683) );
  NOR2_X1 U24043 ( .A1(n34415), .A2(n35738), .ZN(n35745) );
  BUF_X2 U13619 ( .I(n16403), .Z(n12184) );
  NOR2_X1 U24395 ( .A1(n8997), .A2(n4880), .ZN(n8308) );
  CLKBUF_X2 U2639 ( .I(n21938), .Z(n19265) );
  NOR2_X1 U47844 ( .A1(n10340), .A2(n35027), .ZN(n34020) );
  BUF_X2 U2640 ( .I(n15298), .Z(n11024) );
  NAND2_X1 U2529 ( .A1(n11064), .A2(n33993), .ZN(n33989) );
  INV_X1 U2560 ( .I(n60456), .ZN(n1808) );
  INV_X1 U18659 ( .I(n34670), .ZN(n17503) );
  NAND2_X1 U2637 ( .A1(n35802), .A2(n35799), .ZN(n35280) );
  NOR2_X1 U2555 ( .A1(n18878), .A2(n33820), .ZN(n35217) );
  INV_X1 U18658 ( .I(n35032), .ZN(n34631) );
  NOR2_X1 U39940 ( .A1(n34973), .A2(n7883), .ZN(n21041) );
  INV_X1 U13546 ( .I(n34033), .ZN(n33980) );
  INV_X1 U10338 ( .I(n17759), .ZN(n31609) );
  NOR2_X1 U11707 ( .A1(n34324), .A2(n34708), .ZN(n3488) );
  INV_X1 U9557 ( .I(n33542), .ZN(n35618) );
  INV_X1 U5830 ( .I(n34558), .ZN(n33520) );
  INV_X1 U5789 ( .I(n1813), .ZN(n34668) );
  NOR2_X1 U8857 ( .A1(n5085), .A2(n63085), .ZN(n33619) );
  INV_X2 U18683 ( .I(n10682), .ZN(n11061) );
  NAND2_X1 U3588 ( .A1(n11060), .A2(n4231), .ZN(n33598) );
  NAND2_X1 U6723 ( .A1(n34277), .A2(n33776), .ZN(n33494) );
  AND2_X1 U8051 ( .A1(n8405), .A2(n35303), .Z(n57337) );
  INV_X1 U7063 ( .I(n35662), .ZN(n35210) );
  INV_X1 U2651 ( .I(n35705), .ZN(n35749) );
  AND2_X1 U39295 ( .A1(n34614), .A2(n17922), .Z(n33977) );
  INV_X1 U13629 ( .I(n35038), .ZN(n33442) );
  INV_X1 U3541 ( .I(n5927), .ZN(n34014) );
  INV_X1 U25211 ( .I(n4496), .ZN(n33601) );
  NAND2_X1 U28585 ( .A1(n33), .A2(n34658), .ZN(n34001) );
  INV_X1 U3480 ( .I(n35765), .ZN(n7345) );
  INV_X1 U4409 ( .I(n15148), .ZN(n35740) );
  NAND2_X1 U2597 ( .A1(n35629), .A2(n33319), .ZN(n35625) );
  INV_X1 U18181 ( .I(n30467), .ZN(n18301) );
  INV_X1 U13678 ( .I(n8431), .ZN(n33499) );
  OR2_X1 U21829 ( .A1(n25465), .A2(n30895), .Z(n34676) );
  INV_X2 U2607 ( .I(n33560), .ZN(n33693) );
  INV_X1 U32139 ( .I(n13770), .ZN(n35312) );
  CLKBUF_X2 U8877 ( .I(n32528), .Z(n33345) );
  INV_X1 U36360 ( .I(n34335), .ZN(n34343) );
  INV_X1 U2614 ( .I(n35240), .ZN(n35643) );
  NAND2_X1 U2581 ( .A1(n35273), .A2(n10526), .ZN(n18771) );
  NAND2_X1 U21862 ( .A1(n3308), .A2(n62373), .ZN(n13470) );
  NAND2_X1 U3453 ( .A1(n11643), .A2(n5410), .ZN(n59458) );
  NAND2_X1 U2596 ( .A1(n21906), .A2(n3467), .ZN(n34057) );
  OAI21_X1 U48576 ( .A1(n35748), .A2(n35735), .B(n35731), .ZN(n35700) );
  AOI21_X1 U41315 ( .A1(n34262), .A2(n21751), .B(n34746), .ZN(n32221) );
  NOR2_X1 U47629 ( .A1(n33599), .A2(n33338), .ZN(n33015) );
  NOR2_X1 U38958 ( .A1(n33564), .A2(n16939), .ZN(n33094) );
  NAND2_X1 U18663 ( .A1(n5123), .A2(n35032), .ZN(n34503) );
  OAI21_X1 U11667 ( .A1(n34448), .A2(n34447), .B(n35247), .ZN(n35644) );
  INV_X1 U18599 ( .I(n8308), .ZN(n33006) );
  NOR2_X1 U2524 ( .A1(n35730), .A2(n63671), .ZN(n35704) );
  NAND3_X1 U24994 ( .A1(n10401), .A2(n5731), .A3(n5389), .ZN(n32835) );
  NOR2_X1 U10328 ( .A1(n34991), .A2(n34992), .ZN(n13899) );
  NOR2_X1 U40570 ( .A1(n60554), .A2(n14954), .ZN(n31466) );
  NAND2_X1 U13608 ( .A1(n12338), .A2(n34666), .ZN(n24543) );
  AOI21_X1 U9469 ( .A1(n34621), .A2(n12039), .B(n15819), .ZN(n34624) );
  NAND2_X1 U35026 ( .A1(n19253), .A2(n34187), .ZN(n19781) );
  INV_X1 U18457 ( .I(n35217), .ZN(n4169) );
  NAND2_X1 U22868 ( .A1(n1804), .A2(n15830), .ZN(n17426) );
  NAND4_X1 U14363 ( .A1(n34764), .A2(n23366), .A3(n64304), .A4(n64276), .ZN(
        n57600) );
  NAND2_X1 U48200 ( .A1(n63220), .A2(n77), .ZN(n34434) );
  OAI21_X1 U47681 ( .A1(n33701), .A2(n7359), .B(n33693), .ZN(n33691) );
  NAND3_X1 U9406 ( .A1(n17141), .A2(n897), .A3(n35799), .ZN(n35801) );
  NAND2_X1 U18437 ( .A1(n62190), .A2(n33644), .ZN(n6398) );
  NAND4_X1 U13557 ( .A1(n34282), .A2(n34281), .A3(n15927), .A4(n34280), .ZN(
        n34283) );
  NAND2_X1 U13463 ( .A1(n33773), .A2(n33771), .ZN(n22180) );
  NAND2_X1 U20414 ( .A1(n34647), .A2(n34646), .ZN(n58002) );
  NOR2_X1 U9548 ( .A1(n13892), .A2(n35011), .ZN(n35017) );
  NAND3_X1 U47918 ( .A1(n35656), .A2(n34447), .A3(n60835), .ZN(n33587) );
  INV_X1 U23289 ( .I(n33350), .ZN(n33566) );
  NAND2_X1 U2530 ( .A1(n25216), .A2(n62373), .ZN(n34284) );
  NAND2_X1 U47692 ( .A1(n33539), .A2(n33375), .ZN(n33119) );
  NOR2_X1 U22711 ( .A1(n33702), .A2(n4034), .ZN(n9796) );
  NAND2_X1 U2590 ( .A1(n26242), .A2(n35821), .ZN(n34710) );
  NOR2_X1 U47967 ( .A1(n33741), .A2(n33740), .ZN(n33750) );
  INV_X1 U11660 ( .I(n8217), .ZN(n8366) );
  NAND2_X1 U13633 ( .A1(n23774), .A2(n34646), .ZN(n34017) );
  OAI22_X1 U41764 ( .A1(n32437), .A2(n32436), .B1(n32438), .B2(n34759), .ZN(
        n24513) );
  OAI22_X1 U9559 ( .A1(n18089), .A2(n20137), .B1(n33619), .B2(n9085), .ZN(
        n34472) );
  AOI21_X1 U21517 ( .A1(n20736), .A2(n10448), .B(n35799), .ZN(n58150) );
  NAND3_X1 U47605 ( .A1(n33763), .A2(n9648), .A3(n5322), .ZN(n33462) );
  NOR2_X1 U7060 ( .A1(n1535), .A2(n3013), .ZN(n34176) );
  NOR3_X1 U7070 ( .A1(n12350), .A2(n21008), .A3(n33720), .ZN(n34065) );
  NAND2_X1 U11692 ( .A1(n34646), .A2(n34643), .ZN(n34504) );
  NOR2_X1 U4615 ( .A1(n32842), .A2(n17283), .ZN(n33674) );
  NOR2_X1 U18275 ( .A1(n6980), .A2(n6981), .ZN(n4160) );
  NOR3_X1 U42765 ( .A1(n2695), .A2(n25972), .A3(n4097), .ZN(n21215) );
  NAND2_X1 U36401 ( .A1(n10504), .A2(n77), .ZN(n33811) );
  NOR2_X1 U33216 ( .A1(n13352), .A2(n32972), .ZN(n34780) );
  NOR2_X1 U9482 ( .A1(n10267), .A2(n33342), .ZN(n33704) );
  NAND2_X1 U9567 ( .A1(n34084), .A2(n58421), .ZN(n34625) );
  NOR2_X1 U18366 ( .A1(n33894), .A2(n34413), .ZN(n33915) );
  NOR3_X1 U7058 ( .A1(n7047), .A2(n60765), .A3(n34168), .ZN(n34179) );
  NAND2_X1 U13467 ( .A1(n33618), .A2(n33617), .ZN(n11350) );
  NAND2_X1 U10332 ( .A1(n436), .A2(n13818), .ZN(n34547) );
  INV_X1 U8842 ( .I(n11064), .ZN(n34195) );
  INV_X1 U40162 ( .I(n35325), .ZN(n35783) );
  INV_X1 U2625 ( .I(n35307), .ZN(n35826) );
  NAND2_X1 U4737 ( .A1(n18488), .A2(n17141), .ZN(n34298) );
  NAND3_X1 U47517 ( .A1(n33599), .A2(n33304), .A3(n33017), .ZN(n32766) );
  INV_X1 U2548 ( .I(n21906), .ZN(n34518) );
  NAND4_X1 U38457 ( .A1(n61917), .A2(n58702), .A3(n25625), .A4(n59522), .ZN(
        n31419) );
  NOR3_X1 U42231 ( .A1(n35036), .A2(n35035), .A3(n35034), .ZN(n35052) );
  OAI21_X1 U13504 ( .A1(n15466), .A2(n61452), .B(n34502), .ZN(n18646) );
  OAI21_X1 U23029 ( .A1(n60434), .A2(n14269), .B(n4266), .ZN(n6399) );
  NAND3_X1 U36370 ( .A1(n35235), .A2(n57492), .A3(n35848), .ZN(n34399) );
  NAND2_X1 U13485 ( .A1(n22118), .A2(n1807), .ZN(n10757) );
  OAI21_X1 U6104 ( .A1(n33915), .A2(n58562), .B(n61496), .ZN(n12938) );
  NAND4_X1 U2545 ( .A1(n35740), .A2(n2287), .A3(n6051), .A4(n35739), .ZN(
        n35741) );
  NAND2_X1 U18338 ( .A1(n905), .A2(n2899), .ZN(n13651) );
  OAI21_X1 U7076 ( .A1(n11396), .A2(n33966), .B(n58702), .ZN(n11397) );
  NAND3_X1 U13566 ( .A1(n18301), .A2(n34512), .A3(n1424), .ZN(n12952) );
  INV_X1 U7997 ( .I(n33010), .ZN(n5065) );
  AOI22_X1 U34266 ( .A1(n33101), .A2(n63185), .B1(n33104), .B2(n63064), .ZN(
        n59641) );
  AOI21_X1 U3454 ( .A1(n33610), .A2(n32999), .B(n25509), .ZN(n25508) );
  NOR2_X1 U18409 ( .A1(n34988), .A2(n2764), .ZN(n3515) );
  AOI22_X1 U48443 ( .A1(n35244), .A2(n35243), .B1(n35242), .B2(n35655), .ZN(
        n35245) );
  NOR2_X1 U20359 ( .A1(n57991), .A2(n57990), .ZN(n3857) );
  NOR3_X1 U11567 ( .A1(n32865), .A2(n2533), .A3(n64407), .ZN(n2532) );
  NAND2_X1 U38002 ( .A1(n16660), .A2(n34057), .ZN(n34061) );
  NAND2_X1 U22997 ( .A1(n4249), .A2(n34434), .ZN(n12067) );
  INV_X1 U3521 ( .I(n18475), .ZN(n10104) );
  NAND2_X1 U17455 ( .A1(n34733), .A2(n57413), .ZN(n16056) );
  NAND2_X1 U18191 ( .A1(n33748), .A2(n33749), .ZN(n3049) );
  AOI21_X1 U35251 ( .A1(n15838), .A2(n19265), .B(n35701), .ZN(n35703) );
  INV_X1 U48571 ( .I(n35681), .ZN(n35682) );
  NAND2_X1 U30642 ( .A1(n32601), .A2(n14329), .ZN(n59174) );
  NAND2_X1 U47680 ( .A1(n33751), .A2(n33750), .ZN(n3050) );
  NAND3_X1 U39742 ( .A1(n35797), .A2(n35796), .A3(n35798), .ZN(n22586) );
  NOR3_X1 U33661 ( .A1(n35282), .A2(n21764), .A3(n21765), .ZN(n14024) );
  NAND3_X1 U13474 ( .A1(n23177), .A2(n23178), .A3(n9542), .ZN(n9538) );
  NAND2_X1 U20411 ( .A1(n58002), .A2(n58001), .ZN(n58000) );
  OAI21_X1 U13585 ( .A1(n33303), .A2(n33302), .B(n33301), .ZN(n33310) );
  NAND2_X1 U35254 ( .A1(n21456), .A2(n23914), .ZN(n21454) );
  NAND2_X1 U10313 ( .A1(n3995), .A2(n18281), .ZN(n3994) );
  NOR2_X1 U18320 ( .A1(n24513), .A2(n24514), .ZN(n11544) );
  NAND3_X1 U20617 ( .A1(n31906), .A2(n34764), .A3(n23366), .ZN(n34220) );
  OAI21_X1 U13588 ( .A1(n35642), .A2(n58598), .B(n15328), .ZN(n35246) );
  NAND3_X1 U27994 ( .A1(n33469), .A2(n23761), .A3(n560), .ZN(n33470) );
  NAND4_X1 U20616 ( .A1(n18895), .A2(n2388), .A3(n34303), .A4(n34220), .ZN(
        n2387) );
  NAND3_X1 U48243 ( .A1(n34547), .A2(n59293), .A3(n34546), .ZN(n34548) );
  NAND3_X1 U4781 ( .A1(n35761), .A2(n35314), .A3(n61532), .ZN(n35768) );
  AOI22_X1 U35012 ( .A1(n33084), .A2(n24317), .B1(n19789), .B2(n57200), .ZN(
        n33085) );
  AOI21_X1 U6098 ( .A1(n34261), .A2(n34262), .B(n34260), .ZN(n61088) );
  NAND2_X1 U3378 ( .A1(n57734), .A2(n34352), .ZN(n21191) );
  NOR2_X1 U13479 ( .A1(n15141), .A2(n18646), .ZN(n15140) );
  OAI21_X1 U9538 ( .A1(n13892), .A2(n33761), .B(n33760), .ZN(n13891) );
  NOR2_X1 U10319 ( .A1(n35703), .A2(n904), .ZN(n6000) );
  INV_X1 U3328 ( .I(n25893), .ZN(n60165) );
  NAND3_X1 U13568 ( .A1(n15998), .A2(n34055), .A3(n34054), .ZN(n34063) );
  OAI21_X1 U18232 ( .A1(n21807), .A2(n33758), .B(n58713), .ZN(n21806) );
  NOR2_X1 U13451 ( .A1(n19997), .A2(n19996), .ZN(n35790) );
  NOR2_X1 U3337 ( .A1(n5065), .A2(n33002), .ZN(n59485) );
  OAI21_X1 U9540 ( .A1(n19661), .A2(n35250), .B(n9027), .ZN(n9026) );
  NAND2_X1 U2506 ( .A1(n34329), .A2(n34427), .ZN(n16725) );
  INV_X2 U39780 ( .I(n60758), .ZN(n15754) );
  NAND3_X1 U40688 ( .A1(n32793), .A2(n21216), .A3(n32792), .ZN(n22622) );
  BUF_X2 U10292 ( .I(n36116), .Z(n16968) );
  NAND2_X1 U47525 ( .A1(n32780), .A2(n32781), .ZN(n32788) );
  INV_X2 U18025 ( .I(n6606), .ZN(n34478) );
  BUF_X2 U19986 ( .I(n19765), .Z(n57939) );
  INV_X4 U2475 ( .I(n36959), .ZN(n1527) );
  AOI21_X1 U18353 ( .A1(n7293), .A2(n33463), .B(n15575), .ZN(n7068) );
  NAND4_X1 U42475 ( .A1(n35792), .A2(n35791), .A3(n35789), .A4(n35790), .ZN(
        n35793) );
  NAND2_X1 U18355 ( .A1(n34536), .A2(n34548), .ZN(n3718) );
  CLKBUF_X2 U13435 ( .I(n2900), .Z(n4798) );
  INV_X2 U20611 ( .I(n9806), .ZN(n37424) );
  INV_X2 U3858 ( .I(n35341), .ZN(n7118) );
  INV_X1 U37816 ( .I(n16420), .ZN(n22587) );
  INV_X2 U2488 ( .I(n36410), .ZN(n36193) );
  INV_X1 U26907 ( .I(n37411), .ZN(n16501) );
  NOR2_X1 U35796 ( .A1(n20262), .A2(n20261), .ZN(n20252) );
  NOR2_X1 U11485 ( .A1(n36436), .A2(n36444), .ZN(n36219) );
  INV_X2 U9532 ( .I(n36717), .ZN(n1310) );
  NOR3_X1 U27996 ( .A1(n33475), .A2(n35015), .A3(n33474), .ZN(n36470) );
  INV_X4 U42409 ( .I(n34841), .ZN(n37268) );
  CLKBUF_X2 U18142 ( .I(n24365), .Z(n18525) );
  BUF_X2 U16410 ( .I(n33933), .Z(n57686) );
  CLKBUF_X2 U8299 ( .I(n17615), .Z(n8808) );
  INV_X4 U30647 ( .I(n23577), .ZN(n13768) );
  INV_X2 U2481 ( .I(n37358), .ZN(n37361) );
  BUF_X2 U5190 ( .I(n16886), .Z(n35883) );
  INV_X2 U32881 ( .I(n20280), .ZN(n12863) );
  INV_X2 U27101 ( .I(n34846), .ZN(n37269) );
  BUF_X2 U10289 ( .I(n17132), .Z(n8010) );
  INV_X1 U6376 ( .I(n21921), .ZN(n13734) );
  NAND2_X1 U9527 ( .A1(n19507), .A2(n20908), .ZN(n35910) );
  INV_X1 U23508 ( .I(n36768), .ZN(n59910) );
  AND2_X1 U27466 ( .A1(n36410), .A2(n36116), .Z(n35363) );
  INV_X1 U42898 ( .I(n20548), .ZN(n34927) );
  NAND2_X1 U38499 ( .A1(n37130), .A2(n34841), .ZN(n37136) );
  INV_X1 U9905 ( .I(n36818), .ZN(n35238) );
  INV_X4 U2378 ( .I(n57210), .ZN(n18677) );
  NOR2_X1 U36499 ( .A1(n21584), .A2(n652), .ZN(n19778) );
  INV_X2 U2398 ( .I(n9783), .ZN(n37364) );
  CLKBUF_X2 U17947 ( .I(n20531), .Z(n10086) );
  BUF_X2 U2414 ( .I(n36579), .Z(n10498) );
  NAND2_X1 U39138 ( .A1(n37376), .A2(n22317), .ZN(n36597) );
  NOR2_X1 U48523 ( .A1(n22503), .A2(n2383), .ZN(n36910) );
  INV_X2 U9528 ( .I(n37233), .ZN(n1309) );
  INV_X2 U31096 ( .I(n20571), .ZN(n35570) );
  BUF_X2 U15461 ( .I(n15045), .Z(n59261) );
  INV_X2 U5044 ( .I(n35994), .ZN(n21915) );
  NOR3_X1 U8341 ( .A1(n61223), .A2(n59396), .A3(n64263), .ZN(n36257) );
  CLKBUF_X2 U18189 ( .I(n36401), .Z(n10601) );
  BUF_X2 U13273 ( .I(n25788), .Z(n10849) );
  NAND2_X1 U33127 ( .A1(n36909), .A2(n13126), .ZN(n36908) );
  BUF_X2 U6079 ( .I(n23766), .Z(n61180) );
  NAND3_X1 U5627 ( .A1(n16337), .A2(n22993), .A3(n22737), .ZN(n35429) );
  BUF_X2 U42787 ( .I(n36435), .Z(n60562) );
  INV_X2 U2388 ( .I(n35178), .ZN(n12116) );
  NAND2_X1 U2412 ( .A1(n35876), .A2(n37181), .ZN(n37188) );
  INV_X1 U8313 ( .I(n37374), .ZN(n37369) );
  INV_X1 U13440 ( .I(n16337), .ZN(n1789) );
  INV_X1 U42453 ( .I(n33785), .ZN(n35130) );
  NAND2_X1 U19536 ( .A1(n3233), .A2(n36579), .ZN(n7380) );
  NAND2_X1 U38428 ( .A1(n20280), .A2(n20812), .ZN(n36340) );
  AND2_X1 U20567 ( .A1(n58026), .A2(n20908), .Z(n20431) );
  NAND2_X1 U23662 ( .A1(n10829), .A2(n24028), .ZN(n16268) );
  NAND2_X1 U9473 ( .A1(n36777), .A2(n7028), .ZN(n14952) );
  NOR2_X1 U2299 ( .A1(n36691), .A2(n1416), .ZN(n36870) );
  NAND2_X1 U9511 ( .A1(n18144), .A2(n36898), .ZN(n36386) );
  INV_X2 U25570 ( .I(n36195), .ZN(n36412) );
  INV_X2 U2471 ( .I(n6159), .ZN(n21536) );
  INV_X1 U3053 ( .I(n20146), .ZN(n35350) );
  NAND2_X1 U31379 ( .A1(n59910), .A2(n17775), .ZN(n12031) );
  INV_X1 U13432 ( .I(n35899), .ZN(n1788) );
  INV_X1 U2387 ( .I(n61703), .ZN(n36224) );
  INV_X1 U9588 ( .I(n26213), .ZN(n36013) );
  INV_X1 U9722 ( .I(n1417), .ZN(n12885) );
  NOR2_X1 U27783 ( .A1(n36818), .A2(n1235), .ZN(n37399) );
  NOR2_X1 U5379 ( .A1(n25994), .A2(n36979), .ZN(n36980) );
  NOR2_X1 U2340 ( .A1(n35353), .A2(n35974), .ZN(n35352) );
  INV_X2 U9792 ( .I(n22503), .ZN(n37435) );
  AND2_X1 U5189 ( .A1(n36444), .A2(n36435), .Z(n57171) );
  NAND2_X1 U5326 ( .A1(n32984), .A2(n36377), .ZN(n36572) );
  INV_X2 U34793 ( .I(n37363), .ZN(n36589) );
  NAND2_X1 U34641 ( .A1(n1781), .A2(n7729), .ZN(n19052) );
  OAI21_X1 U30012 ( .A1(n61180), .A2(n10849), .B(n19778), .ZN(n19777) );
  NOR2_X1 U9504 ( .A1(n2958), .A2(n37188), .ZN(n2942) );
  NAND3_X1 U4285 ( .A1(n35907), .A2(n64609), .A3(n14904), .ZN(n3585) );
  INV_X1 U37839 ( .I(n12031), .ZN(n36765) );
  NAND2_X1 U17778 ( .A1(n14763), .A2(n60196), .ZN(n35453) );
  NOR2_X1 U2917 ( .A1(n8041), .A2(n6918), .ZN(n35465) );
  NOR2_X1 U38204 ( .A1(n20060), .A2(n15794), .ZN(n16987) );
  NAND2_X1 U36511 ( .A1(n4541), .A2(n37359), .ZN(n18779) );
  NAND2_X1 U17784 ( .A1(n37409), .A2(n37408), .ZN(n5005) );
  INV_X1 U35271 ( .I(n35422), .ZN(n24641) );
  NAND2_X1 U9816 ( .A1(n59963), .A2(n35909), .ZN(n37033) );
  INV_X1 U13425 ( .I(n37326), .ZN(n37183) );
  NAND2_X1 U2425 ( .A1(n18313), .A2(n33607), .ZN(n36190) );
  INV_X1 U18047 ( .I(n34815), .ZN(n35944) );
  INV_X1 U13422 ( .I(n37133), .ZN(n34837) );
  INV_X1 U20875 ( .I(n15011), .ZN(n37375) );
  NAND3_X1 U7083 ( .A1(n57209), .A2(n36959), .A3(n1786), .ZN(n36966) );
  INV_X1 U2359 ( .I(n11077), .ZN(n37371) );
  BUF_X4 U18122 ( .I(n36898), .Z(n7103) );
  CLKBUF_X2 U28063 ( .I(n3149), .Z(n58853) );
  CLKBUF_X2 U7929 ( .I(n22737), .Z(n59842) );
  CLKBUF_X2 U54170 ( .I(n36851), .Z(n61207) );
  NAND2_X1 U30496 ( .A1(n37376), .A2(n1769), .ZN(n34372) );
  CLKBUF_X2 U29984 ( .I(n37454), .Z(n9869) );
  NAND2_X1 U27108 ( .A1(n38551), .A2(n7269), .ZN(n36786) );
  NAND2_X1 U2341 ( .A1(n9593), .A2(n59910), .ZN(n36774) );
  NAND2_X1 U11515 ( .A1(n13983), .A2(n59852), .ZN(n36620) );
  NOR2_X1 U24983 ( .A1(n36852), .A2(n36847), .ZN(n36672) );
  NOR2_X1 U5279 ( .A1(n35454), .A2(n60196), .ZN(n36534) );
  NAND2_X1 U28449 ( .A1(n36494), .A2(n36232), .ZN(n8363) );
  NAND2_X1 U28206 ( .A1(n58876), .A2(n14904), .ZN(n34859) );
  NOR2_X1 U2390 ( .A1(n1779), .A2(n1788), .ZN(n34875) );
  NAND2_X1 U11480 ( .A1(n36875), .A2(n21881), .ZN(n5872) );
  NOR2_X1 U9493 ( .A1(n35357), .A2(n13768), .ZN(n35976) );
  NOR2_X1 U25823 ( .A1(n5936), .A2(n9456), .ZN(n14629) );
  NOR2_X1 U33756 ( .A1(n14189), .A2(n17364), .ZN(n36343) );
  NAND3_X1 U32799 ( .A1(n22559), .A2(n1415), .A3(n35178), .ZN(n36244) );
  INV_X1 U30417 ( .I(n60374), .ZN(n36009) );
  INV_X2 U24763 ( .I(n35353), .ZN(n35543) );
  INV_X1 U35269 ( .I(n21591), .ZN(n16851) );
  INV_X2 U9535 ( .I(n22559), .ZN(n1311) );
  NAND2_X1 U2325 ( .A1(n34914), .A2(n1789), .ZN(n36938) );
  INV_X1 U8452 ( .I(n22632), .ZN(n37365) );
  INV_X1 U34233 ( .I(n35398), .ZN(n36309) );
  INV_X1 U31477 ( .I(n11020), .ZN(n20712) );
  AND2_X1 U33826 ( .A1(n36952), .A2(n22993), .Z(n35432) );
  INV_X1 U33125 ( .I(n36908), .ZN(n37420) );
  NAND2_X1 U11510 ( .A1(n10165), .A2(n35416), .ZN(n36049) );
  NAND2_X1 U2384 ( .A1(n22528), .A2(n21467), .ZN(n35608) );
  INV_X1 U20539 ( .I(n17892), .ZN(n36477) );
  NOR2_X1 U36451 ( .A1(n23146), .A2(n26213), .ZN(n36848) );
  AND2_X1 U17928 ( .A1(n36517), .A2(n9783), .Z(n36511) );
  NAND2_X1 U2389 ( .A1(n35096), .A2(n15805), .ZN(n35483) );
  INV_X1 U37699 ( .I(n20251), .ZN(n23651) );
  INV_X2 U31559 ( .I(n7598), .ZN(n35903) );
  INV_X1 U17996 ( .I(n34852), .ZN(n34365) );
  AND2_X1 U7591 ( .A1(n1235), .A2(n37397), .Z(n899) );
  NOR2_X1 U36486 ( .A1(n22524), .A2(n37030), .ZN(n34860) );
  NAND2_X1 U4078 ( .A1(n20060), .A2(n36777), .ZN(n34368) );
  NOR2_X1 U3101 ( .A1(n21605), .A2(n1422), .ZN(n21606) );
  NAND2_X1 U2290 ( .A1(n36483), .A2(n36494), .ZN(n35153) );
  INV_X1 U11477 ( .I(n36725), .ZN(n35344) );
  INV_X1 U7092 ( .I(n23742), .ZN(n37222) );
  INV_X1 U2311 ( .I(n22737), .ZN(n36889) );
  NAND2_X1 U28525 ( .A1(n1781), .A2(n8438), .ZN(n35449) );
  NOR2_X1 U23796 ( .A1(n11413), .A2(n2362), .ZN(n36462) );
  NOR2_X1 U34232 ( .A1(n36304), .A2(n36803), .ZN(n14810) );
  INV_X4 U21529 ( .I(n57211), .ZN(n36796) );
  INV_X1 U2291 ( .I(n36579), .ZN(n36472) );
  NOR2_X1 U35788 ( .A1(n22461), .A2(n22503), .ZN(n37423) );
  OR2_X1 U7625 ( .A1(n38551), .A2(n57860), .Z(n16027) );
  INV_X2 U33179 ( .I(n36022), .ZN(n36040) );
  INV_X1 U20896 ( .I(n2607), .ZN(n36915) );
  AOI21_X1 U48464 ( .A1(n35340), .A2(n35346), .B(n35344), .ZN(n35343) );
  INV_X1 U2326 ( .I(n17030), .ZN(n37276) );
  NAND2_X1 U49067 ( .A1(n37225), .A2(n3691), .ZN(n37207) );
  NAND2_X1 U5278 ( .A1(n36534), .A2(n20530), .ZN(n4005) );
  NOR2_X1 U17722 ( .A1(n36922), .A2(n11563), .ZN(n11562) );
  NAND2_X1 U2861 ( .A1(n1524), .A2(n36755), .ZN(n60831) );
  OAI21_X1 U13404 ( .A1(n36803), .A2(n61579), .B(n21606), .ZN(n36067) );
  INV_X1 U35264 ( .I(n36188), .ZN(n36118) );
  NAND2_X1 U22430 ( .A1(n35937), .A2(n37435), .ZN(n3766) );
  NAND3_X1 U23203 ( .A1(n37204), .A2(n37205), .A3(n37225), .ZN(n4388) );
  NOR2_X1 U17918 ( .A1(n35944), .A2(n22503), .ZN(n35941) );
  NAND2_X1 U18068 ( .A1(n22559), .A2(n61223), .ZN(n33414) );
  NAND2_X1 U57119 ( .A1(n35543), .A2(n35548), .ZN(n61636) );
  INV_X1 U13369 ( .I(n34368), .ZN(n36050) );
  NOR2_X1 U41797 ( .A1(n35440), .A2(n12652), .ZN(n60441) );
  NOR2_X1 U48381 ( .A1(n35081), .A2(n35080), .ZN(n37098) );
  NOR3_X1 U28122 ( .A1(n8041), .A2(n35979), .A3(n652), .ZN(n10966) );
  AOI21_X1 U9579 ( .A1(n3561), .A2(n36921), .B(n20020), .ZN(n26125) );
  NAND2_X1 U26518 ( .A1(n37112), .A2(n6831), .ZN(n17997) );
  INV_X1 U48897 ( .I(n36780), .ZN(n36783) );
  INV_X1 U17834 ( .I(n19699), .ZN(n6049) );
  INV_X1 U48668 ( .I(n36395), .ZN(n36059) );
  NOR2_X1 U35284 ( .A1(n38551), .A2(n38550), .ZN(n36076) );
  INV_X1 U13406 ( .I(n36310), .ZN(n36801) );
  NAND2_X1 U18133 ( .A1(n35962), .A2(n15754), .ZN(n34475) );
  INV_X1 U13315 ( .I(n7802), .ZN(n14726) );
  INV_X1 U13416 ( .I(n36020), .ZN(n36021) );
  NOR2_X1 U7089 ( .A1(n1243), .A2(n13666), .ZN(n2512) );
  INV_X1 U47896 ( .I(n34100), .ZN(n33522) );
  INV_X1 U23765 ( .I(n37350), .ZN(n4636) );
  OAI21_X1 U20335 ( .A1(n36209), .A2(n36210), .B(n1418), .ZN(n57988) );
  BUF_X2 U42071 ( .I(n22113), .Z(n60462) );
  NAND3_X1 U17719 ( .A1(n5872), .A2(n12236), .A3(n5871), .ZN(n12235) );
  NAND2_X1 U17849 ( .A1(n35549), .A2(n35550), .ZN(n7350) );
  NAND2_X1 U2266 ( .A1(n14904), .A2(n21010), .ZN(n35485) );
  NAND2_X1 U2257 ( .A1(n36309), .A2(n14810), .ZN(n36133) );
  NAND2_X1 U11430 ( .A1(n37341), .A2(n64620), .ZN(n35878) );
  NOR2_X1 U3006 ( .A1(n9041), .A2(n10067), .ZN(n11030) );
  NAND2_X1 U36404 ( .A1(n14196), .A2(n10110), .ZN(n36804) );
  NAND2_X1 U5013 ( .A1(n18144), .A2(n60196), .ZN(n35379) );
  NAND2_X1 U10247 ( .A1(n1788), .A2(n35887), .ZN(n34872) );
  NAND2_X1 U17925 ( .A1(n36864), .A2(n1413), .ZN(n37069) );
  NOR2_X1 U9509 ( .A1(n36580), .A2(n36471), .ZN(n36480) );
  NAND2_X1 U9815 ( .A1(n36875), .A2(n8520), .ZN(n3471) );
  NAND2_X1 U2249 ( .A1(n37424), .A2(n8177), .ZN(n36904) );
  INV_X1 U53581 ( .I(n7662), .ZN(n61165) );
  NOR2_X1 U32747 ( .A1(n34822), .A2(n36040), .ZN(n34827) );
  NOR2_X1 U24679 ( .A1(n36304), .A2(n10110), .ZN(n12393) );
  BUF_X2 U29072 ( .I(n35876), .Z(n61574) );
  BUF_X2 U24523 ( .I(n37181), .Z(n58561) );
  NOR2_X1 U2315 ( .A1(n36169), .A2(n3057), .ZN(n36431) );
  NAND2_X1 U7078 ( .A1(n4541), .A2(n19573), .ZN(n37113) );
  NAND2_X1 U20181 ( .A1(n36423), .A2(n2059), .ZN(n21802) );
  INV_X1 U11500 ( .I(n37393), .ZN(n37065) );
  NOR2_X1 U21058 ( .A1(n37335), .A2(n37328), .ZN(n37324) );
  NAND2_X1 U2957 ( .A1(n57686), .A2(n22936), .ZN(n16380) );
  NAND3_X1 U8461 ( .A1(n61747), .A2(n36850), .A3(n61207), .ZN(n8299) );
  NOR2_X1 U31239 ( .A1(n21058), .A2(n10413), .ZN(n35552) );
  INV_X1 U2899 ( .I(n59362), .ZN(n909) );
  NAND2_X1 U33090 ( .A1(n24118), .A2(n10596), .ZN(n35894) );
  NOR2_X1 U39288 ( .A1(n6918), .A2(n57210), .ZN(n24994) );
  OR2_X1 U22284 ( .A1(n18583), .A2(n23357), .Z(n36348) );
  NAND2_X1 U2268 ( .A1(n18583), .A2(n37210), .ZN(n7759) );
  INV_X1 U2264 ( .I(n36773), .ZN(n1308) );
  INV_X1 U2320 ( .I(n25125), .ZN(n25584) );
  NAND2_X1 U9491 ( .A1(n35972), .A2(n35543), .ZN(n35150) );
  NOR2_X1 U7086 ( .A1(n1415), .A2(n22559), .ZN(n35181) );
  NOR2_X1 U2306 ( .A1(n10067), .A2(n3856), .ZN(n948) );
  AND2_X1 U2890 ( .A1(n1793), .A2(n37049), .Z(n57391) );
  NOR2_X1 U40618 ( .A1(n34914), .A2(n9456), .ZN(n23739) );
  NOR2_X1 U2214 ( .A1(n36796), .A2(n21605), .ZN(n36809) );
  NOR2_X1 U10248 ( .A1(n37096), .A2(n37945), .ZN(n36639) );
  OR2_X1 U2895 ( .A1(n37358), .A2(n4541), .Z(n37111) );
  OAI21_X1 U13376 ( .A1(n9013), .A2(n17720), .B(n35863), .ZN(n18215) );
  NAND2_X1 U9520 ( .A1(n36584), .A2(n1217), .ZN(n12352) );
  NAND2_X1 U35762 ( .A1(n31308), .A2(n35996), .ZN(n19334) );
  NAND2_X1 U34388 ( .A1(n36170), .A2(n59261), .ZN(n35369) );
  INV_X1 U17911 ( .I(n36973), .ZN(n37237) );
  NAND2_X1 U13428 ( .A1(n64405), .A2(n36574), .ZN(n36374) );
  NOR3_X1 U17725 ( .A1(n25056), .A2(n3171), .A3(n36612), .ZN(n25055) );
  NAND3_X1 U11448 ( .A1(n11081), .A2(n36464), .A3(n36583), .ZN(n36468) );
  NOR2_X1 U32181 ( .A1(n12050), .A2(n1244), .ZN(n33931) );
  OAI21_X1 U18015 ( .A1(n2460), .A2(n63593), .B(n12885), .ZN(n35859) );
  NOR2_X1 U22477 ( .A1(n37132), .A2(n37133), .ZN(n37272) );
  INV_X1 U13241 ( .I(n22853), .ZN(n13206) );
  NOR2_X1 U7888 ( .A1(n10317), .A2(n36485), .ZN(n19038) );
  OAI21_X1 U13305 ( .A1(n25585), .A2(n25584), .B(n9041), .ZN(n10506) );
  OAI21_X1 U32327 ( .A1(n59468), .A2(n36427), .B(n12288), .ZN(n36429) );
  NAND2_X1 U8794 ( .A1(n899), .A2(n37400), .ZN(n36819) );
  AOI22_X1 U31430 ( .A1(n35988), .A2(n35987), .B1(n22895), .B2(n36708), .ZN(
        n10967) );
  NOR2_X1 U13373 ( .A1(n1420), .A2(n24118), .ZN(n35565) );
  INV_X1 U13308 ( .I(n19064), .ZN(n35559) );
  NOR2_X1 U2848 ( .A1(n21605), .A2(n36308), .ZN(n36311) );
  NOR2_X1 U49068 ( .A1(n37208), .A2(n37207), .ZN(n37216) );
  INV_X1 U17738 ( .I(n36407), .ZN(n17395) );
  NAND2_X1 U17697 ( .A1(n35263), .A2(n19666), .ZN(n35270) );
  NOR2_X1 U37991 ( .A1(n36301), .A2(n63848), .ZN(n36798) );
  INV_X1 U33436 ( .I(n37943), .ZN(n35087) );
  NOR2_X1 U18119 ( .A1(n37050), .A2(n37049), .ZN(n24775) );
  NOR2_X1 U41801 ( .A1(n37208), .A2(n18583), .ZN(n22531) );
  NAND2_X1 U57003 ( .A1(n61566), .A2(n36551), .ZN(n4001) );
  NAND2_X1 U43094 ( .A1(n19368), .A2(n38550), .ZN(n36084) );
  INV_X1 U13370 ( .I(n35576), .ZN(n17168) );
  NOR2_X1 U35709 ( .A1(n26213), .A2(n61207), .ZN(n18151) );
  OAI21_X1 U11440 ( .A1(n37361), .A2(n4541), .B(n1524), .ZN(n6389) );
  INV_X1 U13289 ( .I(n3649), .ZN(n36466) );
  NAND2_X1 U5184 ( .A1(n36348), .A2(n59617), .ZN(n57542) );
  NAND2_X1 U55685 ( .A1(n21694), .A2(n21693), .ZN(n10100) );
  AOI21_X1 U3814 ( .A1(n36915), .A2(n36916), .B(n36914), .ZN(n37434) );
  NAND2_X1 U41093 ( .A1(n4005), .A2(n4006), .ZN(n60337) );
  NOR3_X1 U2284 ( .A1(n37113), .A2(n1524), .A3(n21536), .ZN(n19677) );
  NAND3_X1 U56981 ( .A1(n61553), .A2(n21769), .A3(n21768), .ZN(n4769) );
  NAND3_X1 U2245 ( .A1(n1311), .A2(n36262), .A3(n63897), .ZN(n12834) );
  NOR2_X1 U22070 ( .A1(n1787), .A2(n21329), .ZN(n35582) );
  NOR2_X1 U26274 ( .A1(n36787), .A2(n22733), .ZN(n37475) );
  NAND2_X1 U7831 ( .A1(n35466), .A2(n35467), .ZN(n60770) );
  NOR2_X1 U13277 ( .A1(n35557), .A2(n36489), .ZN(n19482) );
  NAND2_X1 U2240 ( .A1(n22528), .A2(n9304), .ZN(n35607) );
  INV_X1 U3496 ( .I(n10550), .ZN(n36834) );
  NOR2_X1 U40279 ( .A1(n36663), .A2(n36669), .ZN(n20203) );
  INV_X1 U46509 ( .I(n34863), .ZN(n37031) );
  NAND3_X1 U9867 ( .A1(n36040), .A2(n60891), .A3(n36021), .ZN(n34460) );
  NOR2_X1 U9937 ( .A1(n61770), .A2(n36259), .ZN(n17960) );
  NOR2_X1 U20540 ( .A1(n60462), .A2(n2362), .ZN(n33526) );
  OR2_X1 U11467 ( .A1(n34872), .A2(n7802), .Z(n35170) );
  INV_X1 U17712 ( .I(n37252), .ZN(n18209) );
  NAND2_X1 U48545 ( .A1(n35571), .A2(n576), .ZN(n36019) );
  INV_X1 U18057 ( .I(n34828), .ZN(n35569) );
  AOI21_X1 U35290 ( .A1(n36109), .A2(n36402), .B(n33606), .ZN(n17392) );
  NAND3_X1 U22244 ( .A1(n3620), .A2(n36771), .A3(n35414), .ZN(n35415) );
  NAND2_X1 U17802 ( .A1(n12050), .A2(n2512), .ZN(n37315) );
  NOR2_X1 U28557 ( .A1(n60891), .A2(n8474), .ZN(n35579) );
  INV_X1 U36526 ( .I(n35863), .ZN(n36337) );
  NAND4_X1 U2212 ( .A1(n37477), .A2(n61890), .A3(n37476), .A4(n38544), .ZN(
        n37478) );
  NAND2_X1 U35743 ( .A1(n34908), .A2(n9456), .ZN(n33458) );
  NAND2_X1 U17709 ( .A1(n10506), .A2(n35606), .ZN(n8532) );
  OAI22_X1 U34034 ( .A1(n36744), .A2(n36745), .B1(n36747), .B2(n62617), .ZN(
        n59614) );
  NAND2_X1 U2672 ( .A1(n35170), .A2(n35171), .ZN(n61001) );
  AOI21_X1 U22714 ( .A1(n19560), .A2(n36558), .B(n4035), .ZN(n36375) );
  NAND3_X1 U13210 ( .A1(n13206), .A2(n37415), .A3(n6139), .ZN(n4268) );
  OAI21_X1 U32371 ( .A1(n18812), .A2(n18811), .B(n36959), .ZN(n12341) );
  AOI21_X1 U7783 ( .A1(n60636), .A2(n11337), .B(n17960), .ZN(n14009) );
  NAND3_X1 U16025 ( .A1(n37223), .A2(n37230), .A3(n3171), .ZN(n37232) );
  INV_X1 U7101 ( .I(n13078), .ZN(n1765) );
  AOI21_X1 U17716 ( .A1(n4914), .A2(n63817), .B(n37350), .ZN(n16564) );
  NAND2_X1 U2209 ( .A1(n36124), .A2(n36175), .ZN(n3047) );
  OAI21_X1 U35761 ( .A1(n19334), .A2(n22578), .B(n15582), .ZN(n31309) );
  NOR2_X1 U11407 ( .A1(n19482), .A2(n21131), .ZN(n16606) );
  NAND3_X1 U11466 ( .A1(n931), .A2(n36583), .A3(n12351), .ZN(n2096) );
  AOI21_X1 U48939 ( .A1(n36913), .A2(n36912), .B(n36911), .ZN(n36918) );
  NOR2_X1 U35792 ( .A1(n36780), .A2(n17243), .ZN(n36088) );
  NAND2_X1 U17659 ( .A1(n36065), .A2(n36066), .ZN(n24437) );
  OAI21_X1 U49073 ( .A1(n37230), .A2(n37229), .B(n37228), .ZN(n37231) );
  NAND2_X1 U13360 ( .A1(n36843), .A2(n62920), .ZN(n16455) );
  NOR2_X1 U26973 ( .A1(n20502), .A2(n37443), .ZN(n37453) );
  NOR2_X1 U8780 ( .A1(n36478), .A2(n59379), .ZN(n2095) );
  AOI21_X1 U41091 ( .A1(n20530), .A2(n36537), .B(n60337), .ZN(n4003) );
  INV_X1 U8789 ( .I(n36551), .ZN(n35381) );
  NOR2_X1 U48210 ( .A1(n34463), .A2(n63484), .ZN(n34464) );
  NOR2_X1 U13307 ( .A1(n36616), .A2(n23449), .ZN(n15370) );
  OAI21_X1 U2717 ( .A1(n34462), .A2(n35388), .B(n34821), .ZN(n37616) );
  NAND3_X1 U48750 ( .A1(n36292), .A2(n36291), .A3(n36290), .ZN(n36295) );
  INV_X1 U48833 ( .I(n36585), .ZN(n36594) );
  INV_X1 U17902 ( .I(n37322), .ZN(n37016) );
  INV_X1 U57095 ( .I(n17409), .ZN(n24961) );
  AOI22_X1 U48623 ( .A1(n35864), .A2(n35863), .B1(n35862), .B2(n35861), .ZN(
        n35867) );
  AOI21_X1 U26799 ( .A1(n5287), .A2(n36842), .B(n36014), .ZN(n58909) );
  NAND3_X1 U11383 ( .A1(n23976), .A2(n38702), .A3(n23977), .ZN(n12809) );
  AOI22_X1 U23785 ( .A1(n36607), .A2(n36606), .B1(n36604), .B2(n36605), .ZN(
        n7856) );
  AOI22_X1 U48070 ( .A1(n37023), .A2(n37016), .B1(n37018), .B2(n33935), .ZN(
        n33940) );
  NAND4_X1 U8379 ( .A1(n18150), .A2(n18148), .A3(n18147), .A4(n8299), .ZN(
        n18146) );
  NAND3_X1 U17908 ( .A1(n35368), .A2(n35905), .A3(n35909), .ZN(n7858) );
  NAND3_X1 U35789 ( .A1(n37240), .A2(n37162), .A3(n461), .ZN(n37171) );
  OAI21_X1 U13230 ( .A1(n57453), .A2(n5088), .B(n22116), .ZN(n11321) );
  AOI21_X1 U13242 ( .A1(n36045), .A2(n10165), .B(n11300), .ZN(n11299) );
  AOI22_X1 U11464 ( .A1(n36608), .A2(n61831), .B1(n2483), .B2(n57391), .ZN(
        n7855) );
  NOR3_X1 U11386 ( .A1(n26170), .A2(n34940), .A3(n34938), .ZN(n26171) );
  NAND3_X1 U41238 ( .A1(n36294), .A2(n36297), .A3(n36295), .ZN(n21579) );
  AOI21_X1 U6398 ( .A1(n36025), .A2(n36024), .B(n17166), .ZN(n36036) );
  AOI21_X1 U17791 ( .A1(n34366), .A2(n35414), .B(n34370), .ZN(n17923) );
  NAND2_X1 U20162 ( .A1(n57962), .A2(n57960), .ZN(n37601) );
  INV_X2 U54632 ( .I(n13532), .ZN(n5200) );
  BUF_X2 U9985 ( .I(n6441), .Z(n4947) );
  AOI21_X1 U13226 ( .A1(n37125), .A2(n37493), .B(n20402), .ZN(n13856) );
  INV_X1 U13189 ( .I(n38994), .ZN(n8392) );
  OAI21_X1 U2178 ( .A1(n3648), .A2(n33524), .B(n60462), .ZN(n3647) );
  NAND4_X1 U28733 ( .A1(n25212), .A2(n8637), .A3(n34292), .A4(n8636), .ZN(
        n38004) );
  INV_X2 U2170 ( .I(n703), .ZN(n10898) );
  CLKBUF_X2 U2168 ( .I(n38972), .Z(n23429) );
  INV_X1 U2141 ( .I(n5266), .ZN(n22) );
  AOI21_X1 U4889 ( .A1(n11600), .A2(n12341), .B(n23495), .ZN(n9122) );
  NOR2_X1 U24865 ( .A1(n5200), .A2(n38367), .ZN(n13505) );
  NAND3_X1 U34136 ( .A1(n18059), .A2(n36417), .A3(n14687), .ZN(n39687) );
  BUF_X2 U9986 ( .I(n39310), .Z(n7370) );
  NAND2_X1 U33211 ( .A1(n13344), .A2(n18613), .ZN(n20667) );
  NAND2_X1 U2157 ( .A1(n25342), .A2(n37042), .ZN(n38871) );
  NAND2_X1 U20965 ( .A1(n34699), .A2(n34698), .ZN(n38330) );
  BUF_X2 U51577 ( .I(n2928), .Z(n61061) );
  BUF_X2 U31816 ( .I(n13975), .Z(n11534) );
  BUF_X2 U3825 ( .I(n39714), .Z(n24058) );
  INV_X1 U2164 ( .I(n25130), .ZN(n24435) );
  INV_X2 U6873 ( .I(n37555), .ZN(n38530) );
  INV_X1 U8030 ( .I(n61489), .ZN(n26063) );
  INV_X1 U2147 ( .I(n11828), .ZN(n38578) );
  INV_X1 U11372 ( .I(n24342), .ZN(n39314) );
  INV_X1 U7998 ( .I(n22048), .ZN(n38916) );
  NAND3_X1 U32660 ( .A1(n18700), .A2(n22081), .A3(n63000), .ZN(n12577) );
  INV_X2 U7110 ( .I(n59018), .ZN(n39253) );
  INV_X1 U9457 ( .I(n4667), .ZN(n38909) );
  INV_X1 U49292 ( .I(n59250), .ZN(n38084) );
  BUF_X2 U13464 ( .I(n38745), .Z(n25995) );
  BUF_X2 U2135 ( .I(n23232), .Z(n21098) );
  BUF_X2 U11378 ( .I(n22988), .Z(n9398) );
  BUF_X2 U2149 ( .I(n39222), .Z(n23493) );
  BUF_X2 U17618 ( .I(n38063), .Z(n38645) );
  INV_X1 U25234 ( .I(n63133), .ZN(n18579) );
  BUF_X2 U4329 ( .I(n39592), .Z(n23573) );
  INV_X1 U2144 ( .I(n24536), .ZN(n39710) );
  INV_X1 U2132 ( .I(n38106), .ZN(n24189) );
  INV_X1 U2167 ( .I(n19410), .ZN(n39544) );
  INV_X1 U20412 ( .I(n26044), .ZN(n39385) );
  INV_X1 U2125 ( .I(n38377), .ZN(n39284) );
  INV_X1 U29680 ( .I(n1411), .ZN(n9667) );
  INV_X1 U17585 ( .I(n5244), .ZN(n1756) );
  INV_X1 U34929 ( .I(n23927), .ZN(n25965) );
  INV_X2 U49754 ( .I(n11239), .ZN(n38360) );
  BUF_X2 U3782 ( .I(n39385), .Z(n4563) );
  BUF_X2 U43440 ( .I(n37699), .Z(n39582) );
  NAND2_X1 U4840 ( .A1(n14259), .A2(n18699), .ZN(n18698) );
  BUF_X2 U22303 ( .I(n8353), .Z(n3665) );
  INV_X1 U2126 ( .I(n19687), .ZN(n39238) );
  BUF_X4 U22065 ( .I(n3715), .Z(n3499) );
  NAND2_X1 U10193 ( .A1(n18698), .A2(n22080), .ZN(n39629) );
  BUF_X2 U13509 ( .I(n20048), .Z(n19990) );
  INV_X1 U13179 ( .I(n21607), .ZN(n1518) );
  INV_X1 U29428 ( .I(n24890), .ZN(n40662) );
  INV_X1 U33659 ( .I(n37173), .ZN(n37198) );
  INV_X1 U4080 ( .I(n38336), .ZN(n42441) );
  CLKBUF_X2 U34824 ( .I(n24991), .Z(n61047) );
  INV_X2 U2072 ( .I(n41213), .ZN(n1739) );
  INV_X1 U17474 ( .I(n8576), .ZN(n20856) );
  INV_X2 U32549 ( .I(n24990), .ZN(n21529) );
  INV_X2 U5596 ( .I(n39011), .ZN(n41401) );
  INV_X1 U2605 ( .I(n58527), .ZN(n9143) );
  INV_X2 U10176 ( .I(n41856), .ZN(n42507) );
  INV_X1 U32955 ( .I(n59495), .ZN(n15590) );
  INV_X1 U4392 ( .I(n36649), .ZN(n9215) );
  INV_X1 U40640 ( .I(n39306), .ZN(n40132) );
  INV_X1 U17488 ( .I(n61659), .ZN(n1745) );
  INV_X2 U26866 ( .I(n38026), .ZN(n39418) );
  INV_X2 U42876 ( .I(n38480), .ZN(n40656) );
  INV_X1 U25254 ( .I(n24644), .ZN(n11677) );
  INV_X2 U2064 ( .I(n40070), .ZN(n2234) );
  INV_X1 U9443 ( .I(n11264), .ZN(n6625) );
  INV_X2 U2098 ( .I(n40970), .ZN(n40963) );
  CLKBUF_X2 U30391 ( .I(n41078), .Z(n23484) );
  BUF_X2 U32517 ( .I(n41019), .Z(n12523) );
  INV_X2 U10163 ( .I(n40695), .ZN(n41435) );
  CLKBUF_X2 U17467 ( .I(n38134), .Z(n9875) );
  CLKBUF_X2 U37396 ( .I(n60077), .Z(n59871) );
  NOR2_X1 U26002 ( .A1(n22617), .A2(n1747), .ZN(n40519) );
  BUF_X2 U43184 ( .I(n41469), .Z(n24649) );
  CLKBUF_X2 U7671 ( .I(n40962), .Z(n61333) );
  INV_X2 U42653 ( .I(n41105), .ZN(n40443) );
  CLKBUF_X2 U14634 ( .I(n40100), .Z(n57536) );
  INV_X1 U32554 ( .I(n23348), .ZN(n39509) );
  INV_X2 U23877 ( .I(n42484), .ZN(n25246) );
  INV_X1 U2097 ( .I(n39842), .ZN(n41433) );
  NOR2_X1 U41359 ( .A1(n39241), .A2(n25258), .ZN(n42465) );
  INV_X1 U2082 ( .I(n12382), .ZN(n25229) );
  INV_X1 U2044 ( .I(n23875), .ZN(n20994) );
  INV_X2 U6929 ( .I(n14462), .ZN(n7012) );
  INV_X1 U13174 ( .I(n9872), .ZN(n21920) );
  INV_X1 U2046 ( .I(n40961), .ZN(n40613) );
  INV_X1 U43462 ( .I(n42504), .ZN(n41270) );
  INV_X1 U26838 ( .I(n42285), .ZN(n21493) );
  INV_X1 U2051 ( .I(n38811), .ZN(n1516) );
  INV_X2 U21508 ( .I(n41874), .ZN(n41051) );
  INV_X1 U41553 ( .I(n40962), .ZN(n25137) );
  INV_X1 U2038 ( .I(n23634), .ZN(n40650) );
  NAND2_X1 U5332 ( .A1(n25131), .A2(n40416), .ZN(n10883) );
  NAND3_X1 U3968 ( .A1(n9875), .A2(n18717), .A3(n1274), .ZN(n42517) );
  INV_X1 U13126 ( .I(n40939), .ZN(n40250) );
  NOR2_X1 U7158 ( .A1(n10883), .A2(n40748), .ZN(n40760) );
  NOR2_X1 U36567 ( .A1(n41470), .A2(n40755), .ZN(n18658) );
  INV_X1 U7148 ( .I(n21920), .ZN(n1746) );
  NAND2_X1 U2018 ( .A1(n42477), .A2(n25258), .ZN(n39242) );
  NAND2_X1 U34471 ( .A1(n61477), .A2(n41914), .ZN(n40794) );
  INV_X2 U27198 ( .I(n60075), .ZN(n8017) );
  CLKBUF_X2 U10135 ( .I(n42285), .Z(n16680) );
  NOR2_X1 U1996 ( .A1(n41469), .A2(n40755), .ZN(n40413) );
  BUF_X2 U42791 ( .I(n41162), .Z(n23884) );
  INV_X2 U13169 ( .I(n40315), .ZN(n13984) );
  NAND2_X1 U20581 ( .A1(n59409), .A2(n41054), .ZN(n41066) );
  INV_X1 U9441 ( .I(n7257), .ZN(n40154) );
  INV_X1 U10268 ( .I(n41109), .ZN(n25356) );
  INV_X2 U1990 ( .I(n11279), .ZN(n42480) );
  INV_X1 U1997 ( .I(n41858), .ZN(n22609) );
  INV_X2 U39152 ( .I(n42477), .ZN(n25666) );
  INV_X1 U33226 ( .I(n13357), .ZN(n40708) );
  INV_X2 U20451 ( .I(n40577), .ZN(n2247) );
  INV_X2 U41050 ( .I(n23492), .ZN(n3245) );
  INV_X1 U11268 ( .I(n10041), .ZN(n1730) );
  NAND2_X1 U11303 ( .A1(n22786), .A2(n18241), .ZN(n41039) );
  NOR2_X1 U8743 ( .A1(n40963), .A2(n40959), .ZN(n40614) );
  BUF_X2 U7681 ( .I(n37197), .Z(n40470) );
  INV_X2 U47606 ( .I(n20871), .ZN(n3306) );
  INV_X1 U9387 ( .I(n18278), .ZN(n25305) );
  INV_X2 U43454 ( .I(n40218), .ZN(n40229) );
  INV_X1 U5755 ( .I(n1238), .ZN(n15558) );
  INV_X1 U30540 ( .I(n22809), .ZN(n39164) );
  INV_X1 U6496 ( .I(n12410), .ZN(n10542) );
  INV_X1 U23737 ( .I(n6576), .ZN(n58435) );
  NAND2_X1 U2009 ( .A1(n40970), .A2(n25137), .ZN(n39123) );
  INV_X1 U10209 ( .I(n40962), .ZN(n38607) );
  INV_X1 U5117 ( .I(n40959), .ZN(n60820) );
  INV_X8 U34302 ( .I(n14317), .ZN(n42452) );
  NOR2_X1 U2468 ( .A1(n5319), .A2(n23145), .ZN(n6498) );
  INV_X1 U1829 ( .I(n40025), .ZN(n11941) );
  NAND2_X1 U10072 ( .A1(n41261), .A2(n11316), .ZN(n11099) );
  NOR2_X1 U50858 ( .A1(n63510), .A2(n40721), .ZN(n40724) );
  INV_X1 U17326 ( .I(n2800), .ZN(n11080) );
  NOR2_X1 U28706 ( .A1(n40944), .A2(n40943), .ZN(n58940) );
  NOR2_X1 U12993 ( .A1(n1721), .A2(n2233), .ZN(n40168) );
  BUF_X2 U2434 ( .I(n42259), .Z(n59271) );
  NOR2_X1 U28875 ( .A1(n8812), .A2(n22289), .ZN(n41941) );
  NAND2_X1 U34722 ( .A1(n9725), .A2(n3756), .ZN(n15541) );
  NOR2_X1 U25666 ( .A1(n6016), .A2(n41858), .ZN(n41279) );
  INV_X1 U49297 ( .I(n40557), .ZN(n40826) );
  INV_X1 U17270 ( .I(n40424), .ZN(n39818) );
  INV_X1 U10190 ( .I(n23933), .ZN(n1748) );
  INV_X1 U20271 ( .I(n2124), .ZN(n40951) );
  INV_X1 U17466 ( .I(n23477), .ZN(n14014) );
  NAND2_X1 U50614 ( .A1(n64655), .A2(n41470), .ZN(n39985) );
  NAND2_X1 U13086 ( .A1(n1304), .A2(n17915), .ZN(n13465) );
  NAND2_X1 U10140 ( .A1(n64067), .A2(n60091), .ZN(n40825) );
  NAND2_X1 U23672 ( .A1(n40104), .A2(n40274), .ZN(n37996) );
  BUF_X2 U3608 ( .I(n40218), .Z(n23855) );
  NAND2_X1 U43569 ( .A1(n23046), .A2(n64183), .ZN(n39836) );
  NOR2_X1 U1951 ( .A1(n40924), .A2(n40923), .ZN(n37934) );
  NOR2_X1 U1811 ( .A1(n7618), .A2(n63914), .ZN(n40858) );
  NAND2_X1 U29007 ( .A1(n38049), .A2(n9015), .ZN(n40204) );
  CLKBUF_X2 U29625 ( .I(n42477), .Z(n9627) );
  NAND2_X1 U22249 ( .A1(n41405), .A2(n41400), .ZN(n13669) );
  NAND2_X1 U8095 ( .A1(n40604), .A2(n14306), .ZN(n40609) );
  INV_X2 U2087 ( .I(n23752), .ZN(n23833) );
  INV_X2 U17449 ( .I(n23420), .ZN(n7501) );
  NAND2_X1 U1931 ( .A1(n24633), .A2(n5837), .ZN(n42474) );
  NAND2_X1 U1929 ( .A1(n57615), .A2(n10173), .ZN(n13049) );
  NOR2_X1 U25525 ( .A1(n42477), .A2(n25258), .ZN(n5847) );
  INV_X2 U1913 ( .I(n40713), .ZN(n41149) );
  INV_X1 U34105 ( .I(n20856), .ZN(n18396) );
  NAND2_X1 U50343 ( .A1(n23298), .A2(n9802), .ZN(n40328) );
  NAND3_X1 U5007 ( .A1(n59409), .A2(n59583), .A3(n41874), .ZN(n41888) );
  NAND2_X1 U49063 ( .A1(n40939), .A2(n40464), .ZN(n40933) );
  INV_X1 U8230 ( .I(n9143), .ZN(n42488) );
  INV_X1 U20313 ( .I(n4918), .ZN(n19982) );
  INV_X1 U20098 ( .I(n40603), .ZN(n17450) );
  INV_X1 U50589 ( .I(n41851), .ZN(n42498) );
  OR2_X1 U1845 ( .A1(n20277), .A2(n42299), .Z(n988) );
  INV_X1 U42417 ( .I(n39095), .ZN(n41030) );
  NOR2_X1 U50204 ( .A1(n40523), .A2(n23787), .ZN(n40532) );
  INV_X1 U41561 ( .I(n825), .ZN(n40946) );
  INV_X1 U17397 ( .I(n6932), .ZN(n9091) );
  INV_X1 U28750 ( .I(n40708), .ZN(n41460) );
  INV_X1 U1943 ( .I(n5774), .ZN(n40491) );
  INV_X1 U11282 ( .I(n23472), .ZN(n2193) );
  INV_X1 U2592 ( .I(n40196), .ZN(n19277) );
  INV_X1 U36639 ( .I(n41177), .ZN(n40654) );
  INV_X1 U43215 ( .I(n41017), .ZN(n24743) );
  INV_X1 U43128 ( .I(n3246), .ZN(n40628) );
  NOR2_X1 U1971 ( .A1(n40025), .A2(n40028), .ZN(n20807) );
  NOR2_X1 U19223 ( .A1(n5319), .A2(n40577), .ZN(n12416) );
  NAND2_X1 U28423 ( .A1(n40944), .A2(n22593), .ZN(n39111) );
  INV_X1 U8731 ( .I(n21529), .ZN(n42239) );
  NAND2_X1 U33444 ( .A1(n37773), .A2(n42259), .ZN(n13673) );
  NAND2_X1 U49248 ( .A1(n8017), .A2(n16680), .ZN(n37590) );
  INV_X1 U28200 ( .I(n8117), .ZN(n8303) );
  NOR2_X1 U8733 ( .A1(n42452), .A2(n9808), .ZN(n41310) );
  INV_X1 U10117 ( .I(n8812), .ZN(n42236) );
  OAI21_X1 U35887 ( .A1(n40732), .A2(n57462), .B(n3245), .ZN(n40722) );
  NOR2_X1 U17398 ( .A1(n63119), .A2(n40591), .ZN(n14656) );
  NAND2_X1 U50747 ( .A1(n40854), .A2(n1272), .ZN(n40395) );
  INV_X1 U6402 ( .I(n41432), .ZN(n39845) );
  NAND2_X1 U9434 ( .A1(n1273), .A2(n42215), .ZN(n41833) );
  NAND2_X1 U41400 ( .A1(n21960), .A2(n38604), .ZN(n39127) );
  AOI21_X1 U51348 ( .A1(n42453), .A2(n664), .B(n42452), .ZN(n42454) );
  NOR2_X1 U9394 ( .A1(n40500), .A2(n24743), .ZN(n3611) );
  NAND3_X1 U1838 ( .A1(n40039), .A2(n22943), .A3(n25258), .ZN(n40355) );
  OAI21_X1 U50478 ( .A1(n39999), .A2(n41122), .B(n39992), .ZN(n39697) );
  NAND2_X1 U11317 ( .A1(n40732), .A2(n23492), .ZN(n41206) );
  NOR3_X1 U50753 ( .A1(n40750), .A2(n24649), .A3(n61561), .ZN(n40420) );
  NAND2_X1 U2304 ( .A1(n42433), .A2(n42427), .ZN(n19256) );
  INV_X1 U50898 ( .I(n40855), .ZN(n40860) );
  NOR2_X1 U50304 ( .A1(n23752), .A2(n61986), .ZN(n39325) );
  INV_X1 U10210 ( .I(n39099), .ZN(n41029) );
  NAND4_X1 U24631 ( .A1(n39506), .A2(n11704), .A3(n23890), .A4(n64450), .ZN(
        n3728) );
  NOR2_X1 U1859 ( .A1(n42269), .A2(n59271), .ZN(n41097) );
  NAND2_X1 U21556 ( .A1(n978), .A2(n3078), .ZN(n42279) );
  CLKBUF_X2 U13100 ( .I(n24477), .Z(n7571) );
  NAND2_X1 U13022 ( .A1(n12416), .A2(n42263), .ZN(n20287) );
  AOI21_X1 U1862 ( .A1(n1725), .A2(n8523), .B(n22289), .ZN(n42234) );
  NAND2_X1 U26547 ( .A1(n25816), .A2(n61008), .ZN(n15890) );
  NAND2_X1 U1938 ( .A1(n41234), .A2(n41237), .ZN(n41231) );
  NAND2_X1 U7137 ( .A1(n12975), .A2(n62134), .ZN(n40814) );
  NAND2_X1 U49249 ( .A1(n109), .A2(n37590), .ZN(n40813) );
  NOR2_X1 U1930 ( .A1(n41164), .A2(n23634), .ZN(n40542) );
  NOR2_X1 U1856 ( .A1(n40470), .A2(n40938), .ZN(n40477) );
  NAND2_X1 U2307 ( .A1(n41400), .A2(n41234), .ZN(n41399) );
  INV_X1 U2023 ( .I(n40602), .ZN(n1728) );
  NOR2_X1 U17277 ( .A1(n1505), .A2(n38264), .ZN(n42304) );
  INV_X1 U1875 ( .I(n13909), .ZN(n41172) );
  INV_X1 U33138 ( .I(n205), .ZN(n17964) );
  NAND2_X1 U7134 ( .A1(n6058), .A2(n41858), .ZN(n42293) );
  INV_X1 U2374 ( .I(n41405), .ZN(n58081) );
  NOR2_X1 U21902 ( .A1(n41077), .A2(n64224), .ZN(n40390) );
  INV_X1 U13085 ( .I(n7094), .ZN(n6200) );
  INV_X1 U9431 ( .I(n41414), .ZN(n40405) );
  INV_X1 U10168 ( .I(n41220), .ZN(n40403) );
  INV_X1 U17367 ( .I(n8688), .ZN(n19343) );
  NOR2_X1 U9438 ( .A1(n40804), .A2(n23145), .ZN(n40582) );
  INV_X1 U10235 ( .I(n7907), .ZN(n41083) );
  NOR2_X1 U8459 ( .A1(n4171), .A2(n40315), .ZN(n40087) );
  NOR2_X1 U7146 ( .A1(n40092), .A2(n25246), .ZN(n40319) );
  AND2_X1 U57022 ( .A1(n41105), .A2(n59601), .Z(n40444) );
  INV_X1 U1850 ( .I(n40267), .ZN(n40103) );
  INV_X1 U1841 ( .I(n9393), .ZN(n40670) );
  INV_X1 U17399 ( .I(n14131), .ZN(n2760) );
  NAND2_X1 U42795 ( .A1(n61950), .A2(n41234), .ZN(n39052) );
  INV_X1 U26921 ( .I(n60132), .ZN(n17063) );
  OR2_X1 U40866 ( .A1(n41162), .A2(n23634), .Z(n41168) );
  INV_X1 U2441 ( .I(n10452), .ZN(n59015) );
  INV_X1 U49655 ( .I(n753), .ZN(n40363) );
  INV_X1 U40335 ( .I(n1274), .ZN(n42199) );
  NOR2_X1 U50600 ( .A1(n41082), .A2(n40854), .ZN(n39973) );
  INV_X1 U4801 ( .I(n40472), .ZN(n40935) );
  NOR2_X1 U11296 ( .A1(n3245), .A2(n41197), .ZN(n40636) );
  NOR2_X1 U1896 ( .A1(n42453), .A2(n25606), .ZN(n42447) );
  NOR3_X1 U21117 ( .A1(n41924), .A2(n64768), .A3(n41256), .ZN(n40565) );
  NAND3_X1 U50765 ( .A1(n41113), .A2(n61984), .A3(n18418), .ZN(n40435) );
  NAND2_X1 U43187 ( .A1(n40223), .A2(n40306), .ZN(n24667) );
  NAND3_X1 U13099 ( .A1(n3245), .A2(n61407), .A3(n41197), .ZN(n40638) );
  NAND2_X1 U7129 ( .A1(n22738), .A2(n1728), .ZN(n40502) );
  NAND2_X1 U10097 ( .A1(n40249), .A2(n40248), .ZN(n37938) );
  NAND2_X1 U36727 ( .A1(n8942), .A2(n14512), .ZN(n39809) );
  INV_X1 U9396 ( .I(n6200), .ZN(n1399) );
  NAND2_X1 U11288 ( .A1(n40405), .A2(n41220), .ZN(n41424) );
  NOR2_X1 U32076 ( .A1(n25816), .A2(n11895), .ZN(n25815) );
  NAND2_X1 U10073 ( .A1(n40038), .A2(n5847), .ZN(n40043) );
  NAND2_X1 U10288 ( .A1(n41853), .A2(n41849), .ZN(n16099) );
  NOR2_X1 U23729 ( .A1(n40378), .A2(n39601), .ZN(n39603) );
  OAI21_X1 U7159 ( .A1(n11122), .A2(n11132), .B(n39414), .ZN(n11131) );
  INV_X1 U55600 ( .I(n18827), .ZN(n40615) );
  INV_X1 U1852 ( .I(n41402), .ZN(n41239) );
  OAI22_X1 U13049 ( .A1(n40299), .A2(n40298), .B1(n61994), .B2(n40297), .ZN(
        n11940) );
  OR2_X1 U7699 ( .A1(n41079), .A2(n2693), .Z(n983) );
  NAND2_X1 U2339 ( .A1(n60123), .A2(n40363), .ZN(n41313) );
  NOR2_X1 U13088 ( .A1(n40437), .A2(n39957), .ZN(n40569) );
  NAND2_X1 U5936 ( .A1(n17357), .A2(n58305), .ZN(n17356) );
  NAND2_X1 U50038 ( .A1(n59871), .A2(n41453), .ZN(n41145) );
  NAND2_X1 U20272 ( .A1(n18612), .A2(n2124), .ZN(n40190) );
  NAND2_X1 U43428 ( .A1(n39124), .A2(n39060), .ZN(n40975) );
  OR2_X1 U30808 ( .A1(n1304), .A2(n39950), .Z(n10395) );
  NOR2_X1 U9414 ( .A1(n22079), .A2(n64895), .ZN(n5642) );
  NOR2_X1 U11257 ( .A1(n39048), .A2(n40737), .ZN(n41241) );
  INV_X1 U10261 ( .I(n41918), .ZN(n42247) );
  INV_X1 U1848 ( .I(n41035), .ZN(n20726) );
  OR2_X1 U17272 ( .A1(n40275), .A2(n40107), .Z(n40333) );
  INV_X1 U9425 ( .I(n41166), .ZN(n1729) );
  AOI21_X1 U2265 ( .A1(n41145), .A2(n58996), .B(n41460), .ZN(n41463) );
  NAND3_X1 U11237 ( .A1(n41442), .A2(n41449), .A3(n40381), .ZN(n8243) );
  INV_X1 U50172 ( .I(n40527), .ZN(n39062) );
  NAND2_X1 U37934 ( .A1(n16189), .A2(n16526), .ZN(n41932) );
  AOI22_X1 U45268 ( .A1(n40659), .A2(n40656), .B1(n41186), .B2(n41182), .ZN(
        n60764) );
  OAI21_X1 U13006 ( .A1(n41241), .A2(n41240), .B(n23780), .ZN(n8915) );
  AOI22_X1 U29184 ( .A1(n39092), .A2(n9189), .B1(n38499), .B2(n64147), .ZN(
        n21716) );
  OAI21_X1 U7156 ( .A1(n42302), .A2(n42301), .B(n42300), .ZN(n42307) );
  AOI21_X1 U2181 ( .A1(n4259), .A2(n39505), .B(n40556), .ZN(n59322) );
  OAI21_X1 U33865 ( .A1(n41804), .A2(n41812), .B(n41811), .ZN(n14344) );
  NAND2_X1 U51320 ( .A1(n42304), .A2(n1403), .ZN(n42305) );
  NAND2_X1 U17411 ( .A1(n20726), .A2(n22617), .ZN(n9314) );
  NOR2_X1 U27870 ( .A1(n40439), .A2(n18418), .ZN(n39831) );
  NAND2_X1 U49793 ( .A1(n1729), .A2(n41161), .ZN(n38415) );
  NAND2_X1 U1801 ( .A1(n16842), .A2(n19277), .ZN(n15918) );
  NAND2_X1 U43549 ( .A1(n25397), .A2(n40542), .ZN(n38416) );
  NAND2_X1 U2113 ( .A1(n37598), .A2(n57844), .ZN(n17352) );
  INV_X1 U50969 ( .I(n41081), .ZN(n41087) );
  OAI21_X1 U35085 ( .A1(n39320), .A2(n39321), .B(n61994), .ZN(n25626) );
  AOI21_X1 U41410 ( .A1(n39426), .A2(n39425), .B(n40054), .ZN(n21966) );
  AOI22_X1 U50834 ( .A1(n41880), .A2(n41879), .B1(n24791), .B2(n59803), .ZN(
        n41893) );
  OAI22_X1 U50056 ( .A1(n40707), .A2(n38843), .B1(n1507), .B2(n41149), .ZN(
        n41457) );
  OAI21_X1 U20365 ( .A1(n39827), .A2(n2193), .B(n6103), .ZN(n39828) );
  AOI21_X1 U37347 ( .A1(n38025), .A2(n8486), .B(n59867), .ZN(n13305) );
  NAND2_X1 U8724 ( .A1(n1729), .A2(n3636), .ZN(n40543) );
  NAND3_X1 U17149 ( .A1(n13395), .A2(n41137), .A3(n13465), .ZN(n13466) );
  OAI21_X1 U10217 ( .A1(n61159), .A2(n40465), .B(n40925), .ZN(n40466) );
  AOI22_X1 U8706 ( .A1(n3490), .A2(n1399), .B1(n3493), .B2(n61838), .ZN(n3491)
         );
  NOR3_X1 U4067 ( .A1(n61707), .A2(n8201), .A3(n23634), .ZN(n5304) );
  NAND2_X1 U22271 ( .A1(n25227), .A2(n3642), .ZN(n5303) );
  OAI21_X1 U50794 ( .A1(n41013), .A2(n40508), .B(n41003), .ZN(n40509) );
  NAND3_X1 U50568 ( .A1(n39895), .A2(n40127), .A3(n42483), .ZN(n39896) );
  AOI21_X1 U35988 ( .A1(n39070), .A2(n39071), .B(n24766), .ZN(n24765) );
  NAND2_X1 U2088 ( .A1(n25865), .A2(n3466), .ZN(n40151) );
  NAND2_X1 U17107 ( .A1(n21716), .A2(n13133), .ZN(n13132) );
  NAND2_X1 U6294 ( .A1(n11588), .A2(n11586), .ZN(n19210) );
  OAI22_X1 U23892 ( .A1(n41076), .A2(n41075), .B1(n41074), .B2(n41073), .ZN(
        n41090) );
  NAND3_X1 U50744 ( .A1(n40389), .A2(n41073), .A3(n40388), .ZN(n40392) );
  NOR2_X1 U17037 ( .A1(n39952), .A2(n11015), .ZN(n15380) );
  AOI21_X1 U31450 ( .A1(n59286), .A2(n40148), .B(n59285), .ZN(n60774) );
  OAI21_X1 U10461 ( .A1(n24272), .A2(n39981), .B(n24271), .ZN(n39816) );
  NOR3_X1 U50782 ( .A1(n40935), .A2(n40474), .A3(n62157), .ZN(n40475) );
  NOR2_X1 U40174 ( .A1(n41847), .A2(n41846), .ZN(n43486) );
  NAND2_X1 U30426 ( .A1(n40266), .A2(n40265), .ZN(n40897) );
  INV_X2 U56577 ( .I(n13823), .ZN(n23877) );
  AOI22_X1 U50783 ( .A1(n40478), .A2(n40477), .B1(n40476), .B2(n40475), .ZN(
        n40479) );
  NAND3_X1 U1765 ( .A1(n38839), .A2(n38840), .A3(n39021), .ZN(n20863) );
  NAND2_X1 U20721 ( .A1(n14288), .A2(n14286), .ZN(n39860) );
  NOR2_X1 U12930 ( .A1(n5796), .A2(n5795), .ZN(n5794) );
  BUF_X4 U7298 ( .I(n15557), .Z(n57873) );
  NAND2_X1 U16998 ( .A1(n41187), .A2(n59554), .ZN(n41229) );
  NOR2_X1 U10524 ( .A1(n65262), .A2(n1717), .ZN(n43185) );
  INV_X2 U21009 ( .I(n15539), .ZN(n23557) );
  INV_X2 U27497 ( .I(n43281), .ZN(n24179) );
  INV_X2 U12914 ( .I(n63485), .ZN(n1493) );
  INV_X2 U1657 ( .I(n20942), .ZN(n18104) );
  INV_X2 U57164 ( .I(n19248), .ZN(n19241) );
  NAND2_X1 U1760 ( .A1(n21055), .A2(n13306), .ZN(n19517) );
  INV_X2 U27091 ( .I(n23877), .ZN(n42600) );
  BUF_X4 U3563 ( .I(n43166), .Z(n4789) );
  BUF_X4 U56898 ( .I(n23017), .Z(n5398) );
  INV_X4 U30398 ( .I(n43733), .ZN(n42118) );
  NAND3_X1 U12860 ( .A1(n25928), .A2(n24360), .A3(n18104), .ZN(n42842) );
  BUF_X4 U17024 ( .I(n40015), .Z(n43438) );
  CLKBUF_X2 U41555 ( .I(n42986), .Z(n22228) );
  NAND2_X1 U1709 ( .A1(n42324), .A2(n15557), .ZN(n5262) );
  BUF_X2 U16807 ( .I(n63485), .Z(n10111) );
  BUF_X2 U16904 ( .I(n15539), .Z(n12864) );
  INV_X2 U24509 ( .I(n43572), .ZN(n43569) );
  INV_X2 U5917 ( .I(n25942), .ZN(n57197) );
  INV_X2 U42880 ( .I(n41987), .ZN(n41980) );
  INV_X2 U51023 ( .I(n43241), .ZN(n43657) );
  INV_X2 U7195 ( .I(n1494), .ZN(n42750) );
  INV_X2 U48182 ( .I(n41997), .ZN(n42327) );
  INV_X1 U1579 ( .I(n21644), .ZN(n42732) );
  INV_X2 U29186 ( .I(n9190), .ZN(n42554) );
  NAND2_X1 U5063 ( .A1(n21667), .A2(n6601), .ZN(n21950) );
  NAND2_X1 U10438 ( .A1(n20602), .A2(n43161), .ZN(n42564) );
  INV_X2 U1726 ( .I(n23003), .ZN(n42608) );
  NAND2_X1 U4453 ( .A1(n20601), .A2(n11179), .ZN(n43157) );
  INV_X2 U21218 ( .I(n1225), .ZN(n43130) );
  BUF_X8 U3710 ( .I(n23132), .Z(n11229) );
  INV_X8 U21637 ( .I(n3133), .ZN(n42355) );
  INV_X2 U33072 ( .I(n43319), .ZN(n42807) );
  INV_X1 U32601 ( .I(n41242), .ZN(n42835) );
  NAND2_X1 U1574 ( .A1(n1715), .A2(n41695), .ZN(n42739) );
  NAND3_X1 U8664 ( .A1(n63666), .A2(n42784), .A3(n42785), .ZN(n9634) );
  INV_X1 U9366 ( .I(n43874), .ZN(n1709) );
  INV_X1 U10078 ( .I(n42784), .ZN(n42781) );
  BUF_X2 U5118 ( .I(n43693), .Z(n22989) );
  NOR3_X1 U30179 ( .A1(n20942), .A2(n41635), .A3(n41634), .ZN(n42120) );
  NOR2_X1 U9338 ( .A1(n8537), .A2(n42180), .ZN(n42775) );
  BUF_X4 U4000 ( .I(n8289), .Z(n8290) );
  BUF_X4 U41770 ( .I(n40482), .Z(n42140) );
  NAND2_X1 U3794 ( .A1(n16447), .A2(n43415), .ZN(n43416) );
  NOR2_X1 U4182 ( .A1(n20888), .A2(n43504), .ZN(n42642) );
  BUF_X2 U5931 ( .I(n43468), .Z(n57198) );
  CLKBUF_X2 U1741 ( .I(n17950), .Z(n7451) );
  BUF_X2 U47097 ( .I(n5787), .Z(n60843) );
  NAND2_X1 U6539 ( .A1(n16447), .A2(n43679), .ZN(n42097) );
  INV_X2 U1769 ( .I(n15557), .ZN(n23184) );
  NOR2_X1 U33846 ( .A1(n8538), .A2(n39081), .ZN(n43029) );
  INV_X2 U37728 ( .I(n42668), .ZN(n42670) );
  NAND3_X1 U43368 ( .A1(n1301), .A2(n40898), .A3(n25169), .ZN(n41719) );
  BUF_X2 U2021 ( .I(n18724), .Z(n16890) );
  INV_X1 U32145 ( .I(n20700), .ZN(n43741) );
  AND2_X1 U2005 ( .A1(n5125), .A2(n13823), .Z(n41796) );
  NAND2_X1 U9328 ( .A1(n63485), .A2(n39427), .ZN(n42422) );
  NAND2_X1 U1688 ( .A1(n15540), .A2(n12864), .ZN(n43953) );
  NAND2_X1 U4962 ( .A1(n61388), .A2(n43099), .ZN(n43102) );
  INV_X1 U36904 ( .I(n42858), .ZN(n20338) );
  NAND2_X1 U1691 ( .A1(n26020), .A2(n43460), .ZN(n43476) );
  NAND2_X1 U43723 ( .A1(n24884), .A2(n41568), .ZN(n43375) );
  INV_X4 U50963 ( .I(n41046), .ZN(n42871) );
  INV_X4 U41678 ( .I(n57197), .ZN(n43437) );
  NAND2_X1 U1677 ( .A1(n43845), .A2(n57591), .ZN(n39938) );
  NOR2_X1 U1729 ( .A1(n40866), .A2(n20942), .ZN(n43734) );
  NOR2_X1 U28518 ( .A1(n42080), .A2(n19793), .ZN(n16148) );
  NAND2_X1 U35209 ( .A1(n10457), .A2(n26020), .ZN(n42419) );
  NAND2_X1 U1693 ( .A1(n1717), .A2(n20888), .ZN(n43183) );
  INV_X1 U31451 ( .I(n11747), .ZN(n43836) );
  NAND2_X1 U24665 ( .A1(n64536), .A2(n41789), .ZN(n372) );
  AOI21_X1 U51280 ( .A1(n42139), .A2(n43254), .B(n42666), .ZN(n42142) );
  NAND2_X1 U2036 ( .A1(n42410), .A2(n58343), .ZN(n59737) );
  OAI21_X1 U10341 ( .A1(n2160), .A2(n42694), .B(n19928), .ZN(n42696) );
  NOR2_X1 U51081 ( .A1(n43700), .A2(n62346), .ZN(n41489) );
  BUF_X2 U7253 ( .I(n8247), .Z(n60866) );
  NAND2_X1 U24045 ( .A1(n43734), .A2(n8290), .ZN(n17928) );
  NOR2_X1 U55997 ( .A1(n3026), .A2(n43183), .ZN(n43177) );
  AOI21_X1 U43813 ( .A1(n42670), .A2(n43254), .B(n42140), .ZN(n42141) );
  NOR2_X1 U1703 ( .A1(n42357), .A2(n1500), .ZN(n41612) );
  NAND3_X1 U51129 ( .A1(n11229), .A2(n23561), .A3(n41624), .ZN(n41628) );
  NOR2_X1 U36986 ( .A1(n8799), .A2(n429), .ZN(n37539) );
  NAND2_X1 U32906 ( .A1(n3674), .A2(n1714), .ZN(n12965) );
  NAND2_X1 U6336 ( .A1(n43449), .A2(n43439), .ZN(n40017) );
  NAND2_X1 U1551 ( .A1(n42607), .A2(n42605), .ZN(n8798) );
  INV_X1 U51044 ( .I(n41554), .ZN(n41339) );
  OAI21_X1 U10582 ( .A1(n8468), .A2(n8469), .B(n43288), .ZN(n60932) );
  NAND2_X1 U43490 ( .A1(n41353), .A2(n43225), .ZN(n42013) );
  NAND2_X1 U38279 ( .A1(n43457), .A2(n62686), .ZN(n42414) );
  NAND2_X1 U33550 ( .A1(n43582), .A2(n43569), .ZN(n13854) );
  BUF_X4 U5018 ( .I(n42826), .Z(n6705) );
  OAI21_X1 U16535 ( .A1(n42025), .A2(n42031), .B(n42023), .ZN(n2708) );
  NAND3_X1 U32574 ( .A1(n60952), .A2(n41779), .A3(n42871), .ZN(n42169) );
  NOR2_X1 U1521 ( .A1(n43444), .A2(n43438), .ZN(n42372) );
  NOR2_X1 U33112 ( .A1(n1495), .A2(n43980), .ZN(n43975) );
  CLKBUF_X2 U34764 ( .I(n12677), .Z(n59709) );
  NOR2_X1 U16564 ( .A1(n4197), .A2(n20922), .ZN(n42352) );
  NOR2_X1 U9355 ( .A1(n23700), .A2(n2735), .ZN(n41711) );
  NAND2_X1 U12816 ( .A1(n42782), .A2(n9792), .ZN(n42184) );
  NAND2_X1 U26096 ( .A1(n4575), .A2(n295), .ZN(n42876) );
  NOR2_X1 U6081 ( .A1(n1716), .A2(n22898), .ZN(n43612) );
  NOR2_X1 U1642 ( .A1(n43288), .A2(n23700), .ZN(n43116) );
  BUF_X2 U5908 ( .I(n11197), .Z(n11198) );
  INV_X2 U34476 ( .I(n18398), .ZN(n22182) );
  NAND2_X1 U1667 ( .A1(n42605), .A2(n9200), .ZN(n42594) );
  INV_X2 U6030 ( .I(n2824), .ZN(n23279) );
  NOR2_X1 U32123 ( .A1(n14496), .A2(n12864), .ZN(n24191) );
  INV_X1 U12937 ( .I(n42916), .ZN(n42555) );
  BUF_X2 U16973 ( .I(n14620), .Z(n22446) );
  NOR2_X1 U1531 ( .A1(n1706), .A2(n6007), .ZN(n43984) );
  INV_X2 U32612 ( .I(n1708), .ZN(n43341) );
  BUF_X2 U1724 ( .I(n14955), .Z(n14605) );
  INV_X1 U12900 ( .I(n42397), .ZN(n1695) );
  INV_X1 U25602 ( .I(n1714), .ZN(n43042) );
  NAND2_X1 U49484 ( .A1(n20242), .A2(n1705), .ZN(n41490) );
  NAND2_X1 U30602 ( .A1(n11039), .A2(n1335), .ZN(n59356) );
  INV_X1 U1917 ( .I(n42922), .ZN(n1698) );
  NAND2_X1 U33568 ( .A1(n43733), .A2(n15007), .ZN(n13882) );
  NOR2_X1 U1532 ( .A1(n5939), .A2(n41970), .ZN(n41522) );
  INV_X1 U26039 ( .I(n6388), .ZN(n42910) );
  INV_X1 U1607 ( .I(n8912), .ZN(n18858) );
  BUF_X2 U6375 ( .I(n2879), .Z(n541) );
  INV_X1 U3484 ( .I(n42676), .ZN(n1497) );
  NAND2_X1 U27435 ( .A1(n21667), .A2(n43288), .ZN(n21935) );
  INV_X1 U28354 ( .I(n42008), .ZN(n42998) );
  INV_X2 U22852 ( .I(n42140), .ZN(n42667) );
  NAND2_X1 U7744 ( .A1(n4077), .A2(n4198), .ZN(n42553) );
  NAND2_X1 U43021 ( .A1(n19928), .A2(n42387), .ZN(n42377) );
  NOR2_X1 U33881 ( .A1(n41779), .A2(n42865), .ZN(n42866) );
  NOR2_X1 U1578 ( .A1(n12677), .A2(n23557), .ZN(n43303) );
  NAND2_X1 U28375 ( .A1(n19358), .A2(n8290), .ZN(n14405) );
  INV_X2 U5089 ( .I(n43444), .ZN(n43447) );
  OAI21_X1 U11147 ( .A1(n42076), .A2(n42082), .B(n42075), .ZN(n42077) );
  OAI21_X1 U10446 ( .A1(n17755), .A2(n63455), .B(n43297), .ZN(n10275) );
  NAND2_X1 U1849 ( .A1(n61344), .A2(n42788), .ZN(n24762) );
  OAI22_X1 U25889 ( .A1(n16705), .A2(n43339), .B1(n12972), .B2(n8185), .ZN(
        n21549) );
  NOR2_X1 U4195 ( .A1(n41558), .A2(n41784), .ZN(n42137) );
  NAND3_X1 U27909 ( .A1(n43284), .A2(n43292), .A3(n43285), .ZN(n24275) );
  OAI21_X1 U5996 ( .A1(n42607), .A2(n42600), .B(n42599), .ZN(n42602) );
  NAND3_X1 U7191 ( .A1(n9162), .A2(n4282), .A3(n43714), .ZN(n13207) );
  OAI22_X1 U51083 ( .A1(n43395), .A2(n41491), .B1(n43391), .B2(n14214), .ZN(
        n41492) );
  NAND2_X1 U1893 ( .A1(n41604), .A2(n5773), .ZN(n59439) );
  NAND4_X1 U27396 ( .A1(n9504), .A2(n4789), .A3(n43155), .A4(n20601), .ZN(
        n14700) );
  INV_X1 U3568 ( .I(n43170), .ZN(n18822) );
  AOI21_X1 U11130 ( .A1(n9377), .A2(n42768), .B(n60432), .ZN(n42771) );
  INV_X1 U22280 ( .I(n3653), .ZN(n8213) );
  NOR2_X1 U1827 ( .A1(n3606), .A2(n43326), .ZN(n58736) );
  NOR3_X1 U13168 ( .A1(n65228), .A2(n43381), .A3(n11198), .ZN(n57614) );
  INV_X1 U1557 ( .I(n43365), .ZN(n1490) );
  AOI21_X1 U10009 ( .A1(n9032), .A2(n1695), .B(n14506), .ZN(n41708) );
  OR2_X1 U45687 ( .A1(n1714), .A2(n15784), .Z(n43041) );
  NOR2_X1 U29224 ( .A1(n43300), .A2(n43299), .ZN(n43955) );
  NAND2_X1 U43093 ( .A1(n43703), .A2(n12034), .ZN(n43036) );
  NAND2_X1 U56852 ( .A1(n41794), .A2(n61465), .ZN(n9214) );
  INV_X1 U12873 ( .I(n41567), .ZN(n1691) );
  NAND2_X1 U6482 ( .A1(n42697), .A2(n42703), .ZN(n42701) );
  NOR2_X1 U50462 ( .A1(n42118), .A2(n14405), .ZN(n43214) );
  INV_X2 U34650 ( .I(n43699), .ZN(n43690) );
  NAND2_X1 U51265 ( .A1(n43624), .A2(n43626), .ZN(n42092) );
  INV_X2 U1654 ( .I(n41350), .ZN(n22112) );
  NAND2_X1 U10027 ( .A1(n6297), .A2(n1297), .ZN(n42927) );
  BUF_X2 U1911 ( .I(n43383), .Z(n577) );
  BUF_X2 U10726 ( .I(n43679), .Z(n22553) );
  NAND2_X1 U7180 ( .A1(n42998), .A2(n11476), .ZN(n41354) );
  NAND2_X1 U1633 ( .A1(n16527), .A2(n4275), .ZN(n43392) );
  NAND2_X1 U11093 ( .A1(n23485), .A2(n60583), .ZN(n43202) );
  NAND3_X1 U38983 ( .A1(n23838), .A2(n41550), .A3(n1491), .ZN(n41547) );
  NAND2_X1 U1627 ( .A1(n8911), .A2(n42681), .ZN(n42836) );
  NAND2_X1 U11184 ( .A1(n19702), .A2(n43079), .ZN(n43843) );
  NAND2_X1 U1542 ( .A1(n43290), .A2(n23700), .ZN(n16377) );
  NAND2_X1 U1619 ( .A1(n5261), .A2(n57873), .ZN(n42332) );
  NOR2_X1 U50710 ( .A1(n22999), .A2(n1499), .ZN(n42362) );
  NAND2_X1 U10727 ( .A1(n4659), .A2(n1020), .ZN(n42996) );
  INV_X1 U25791 ( .I(n6144), .ZN(n43352) );
  NAND2_X1 U1518 ( .A1(n1708), .A2(n61859), .ZN(n43607) );
  NAND2_X1 U1614 ( .A1(n8912), .A2(n541), .ZN(n20784) );
  NOR2_X1 U10499 ( .A1(n65217), .A2(n63529), .ZN(n7620) );
  NAND2_X1 U39659 ( .A1(n6388), .A2(n10415), .ZN(n42102) );
  NAND2_X1 U12853 ( .A1(n12760), .A2(n43341), .ZN(n42156) );
  INV_X1 U9352 ( .I(n14051), .ZN(n42931) );
  INV_X1 U1927 ( .I(n43027), .ZN(n57196) );
  NAND2_X1 U1529 ( .A1(n8028), .A2(n8962), .ZN(n6926) );
  INV_X2 U1680 ( .I(n5939), .ZN(n42383) );
  NAND2_X1 U1620 ( .A1(n12962), .A2(n1714), .ZN(n42926) );
  NOR2_X1 U21056 ( .A1(n43286), .A2(n2735), .ZN(n43117) );
  NAND2_X1 U10736 ( .A1(n42672), .A2(n42676), .ZN(n42839) );
  NOR2_X1 U51101 ( .A1(n5126), .A2(n42608), .ZN(n42601) );
  NOR2_X1 U37977 ( .A1(n43736), .A2(n8290), .ZN(n43738) );
  NAND2_X1 U10021 ( .A1(n22989), .A2(n12034), .ZN(n43697) );
  NOR2_X1 U35473 ( .A1(n5939), .A2(n2160), .ZN(n42687) );
  NAND2_X1 U1585 ( .A1(n43513), .A2(n1717), .ZN(n43511) );
  INV_X1 U35431 ( .I(n42962), .ZN(n42971) );
  OR2_X1 U12540 ( .A1(n42784), .A2(n8361), .Z(n57256) );
  INV_X1 U51127 ( .I(n42589), .ZN(n41626) );
  INV_X1 U9351 ( .I(n43612), .ZN(n43336) );
  INV_X1 U4989 ( .I(n42650), .ZN(n42654) );
  INV_X1 U9360 ( .I(n43094), .ZN(n43220) );
  INV_X1 U1666 ( .I(n1392), .ZN(n12073) );
  NAND3_X1 U1909 ( .A1(n8028), .A2(n43270), .A3(n1398), .ZN(n25556) );
  NAND2_X1 U5983 ( .A1(n12760), .A2(n8619), .ZN(n8171) );
  NOR2_X1 U4119 ( .A1(n63036), .A2(n57873), .ZN(n40908) );
  NAND2_X1 U8012 ( .A1(n42019), .A2(n12034), .ZN(n43696) );
  AOI22_X1 U1790 ( .A1(n42338), .A2(n43581), .B1(n2994), .B2(n5398), .ZN(
        n41964) );
  OAI21_X1 U23115 ( .A1(n43273), .A2(n8028), .B(n43272), .ZN(n4332) );
  NAND2_X1 U9316 ( .A1(n3606), .A2(n2496), .ZN(n8654) );
  OAI21_X1 U4292 ( .A1(n41694), .A2(n12073), .B(n11817), .ZN(n12140) );
  NOR3_X1 U16828 ( .A1(n6685), .A2(n43736), .A3(n15089), .ZN(n15090) );
  NOR2_X1 U28632 ( .A1(n43023), .A2(n8537), .ZN(n20852) );
  OAI21_X1 U41280 ( .A1(n42648), .A2(n42655), .B(n60351), .ZN(n8052) );
  AOI21_X1 U50810 ( .A1(n41559), .A2(n21376), .B(n42848), .ZN(n40546) );
  NOR2_X1 U16839 ( .A1(n43029), .A2(n43022), .ZN(n20853) );
  NOR2_X1 U36992 ( .A1(n42097), .A2(n43548), .ZN(n17246) );
  OAI21_X1 U12884 ( .A1(n57177), .A2(n2557), .B(n65217), .ZN(n10848) );
  NAND3_X1 U7177 ( .A1(n42314), .A2(n42324), .A3(n42328), .ZN(n42323) );
  NAND3_X1 U22952 ( .A1(n43036), .A2(n18363), .A3(n63386), .ZN(n43038) );
  NAND2_X1 U36898 ( .A1(n61744), .A2(n25210), .ZN(n19397) );
  NAND3_X1 U11138 ( .A1(n43868), .A2(n43351), .A3(n43350), .ZN(n6396) );
  AOI21_X1 U21884 ( .A1(n42777), .A2(n9792), .B(n57196), .ZN(n58192) );
  AOI21_X1 U21634 ( .A1(n9043), .A2(n4197), .B(n3126), .ZN(n5367) );
  NAND2_X1 U12822 ( .A1(n41986), .A2(n41611), .ZN(n5365) );
  NAND3_X1 U1558 ( .A1(n1500), .A2(n41980), .A3(n1499), .ZN(n41983) );
  INV_X1 U36934 ( .I(n42724), .ZN(n42725) );
  INV_X1 U12815 ( .I(n26227), .ZN(n8786) );
  OAI21_X1 U11071 ( .A1(n43719), .A2(n43718), .B(n64156), .ZN(n13670) );
  AOI22_X1 U1560 ( .A1(n42166), .A2(n41779), .B1(n41509), .B2(n42871), .ZN(
        n41521) );
  NAND2_X1 U29611 ( .A1(n61859), .A2(n11229), .ZN(n43608) );
  NOR2_X1 U9365 ( .A1(n43043), .A2(n1714), .ZN(n42545) );
  NOR2_X1 U25873 ( .A1(n16850), .A2(n42878), .ZN(n42345) );
  NOR2_X1 U25636 ( .A1(n43559), .A2(n5972), .ZN(n20590) );
  NAND2_X1 U1564 ( .A1(n43391), .A2(n7282), .ZN(n43692) );
  NAND2_X1 U22160 ( .A1(n43521), .A2(n43518), .ZN(n42042) );
  NAND2_X1 U51116 ( .A1(n5773), .A2(n9191), .ZN(n42557) );
  BUF_X2 U38951 ( .I(n11179), .Z(n60079) );
  AOI21_X1 U10793 ( .A1(n1395), .A2(n65181), .B(n42151), .ZN(n41243) );
  INV_X1 U1495 ( .I(n43345), .ZN(n403) );
  NAND2_X1 U8686 ( .A1(n43079), .A2(n10990), .ZN(n15502) );
  NAND3_X1 U9348 ( .A1(n43270), .A2(n2330), .A3(n1398), .ZN(n15219) );
  NAND2_X1 U51744 ( .A1(n60583), .A2(n60052), .ZN(n43846) );
  INV_X1 U37886 ( .I(n42756), .ZN(n42753) );
  AOI21_X1 U11109 ( .A1(n42184), .A2(n42781), .B(n43023), .ZN(n42187) );
  NAND2_X1 U1884 ( .A1(n42338), .A2(n59746), .ZN(n59416) );
  NAND3_X1 U41337 ( .A1(n42564), .A2(n20602), .A3(n42892), .ZN(n16474) );
  OAI22_X1 U11076 ( .A1(n41966), .A2(n43572), .B1(n42716), .B2(n5340), .ZN(
        n5339) );
  NAND4_X1 U9308 ( .A1(n43253), .A2(n43252), .A3(n43251), .A4(n64105), .ZN(
        n2010) );
  NAND2_X1 U39432 ( .A1(n19004), .A2(n43814), .ZN(n42349) );
  AOI21_X1 U51520 ( .A1(n43097), .A2(n64651), .B(n43096), .ZN(n43101) );
  OAI22_X1 U26295 ( .A1(n43210), .A2(n1702), .B1(n21851), .B2(n43733), .ZN(
        n18021) );
  NOR3_X1 U16718 ( .A1(n43434), .A2(n58850), .A3(n18407), .ZN(n15856) );
  NOR4_X1 U4071 ( .A1(n43118), .A2(n43116), .A3(n20844), .A4(n40882), .ZN(
        n16387) );
  AOI22_X1 U27886 ( .A1(n42147), .A2(n42149), .B1(n42152), .B2(n42827), .ZN(
        n7830) );
  NAND2_X1 U30752 ( .A1(n15119), .A2(n16569), .ZN(n10354) );
  NAND3_X1 U5231 ( .A1(n5773), .A2(n42919), .A3(n1718), .ZN(n15494) );
  NOR2_X1 U9310 ( .A1(n43219), .A2(n43225), .ZN(n43223) );
  NAND2_X1 U12747 ( .A1(n4531), .A2(n42185), .ZN(n4530) );
  NAND2_X1 U16651 ( .A1(n41596), .A2(n43350), .ZN(n7449) );
  AOI21_X1 U21882 ( .A1(n58192), .A2(n58191), .B(n777), .ZN(n22538) );
  AOI21_X1 U51506 ( .A1(n43040), .A2(n43039), .B(n62546), .ZN(n43049) );
  NAND2_X1 U50593 ( .A1(n43061), .A2(n39941), .ZN(n39942) );
  NAND3_X1 U24133 ( .A1(n1005), .A2(n18995), .A3(n1006), .ZN(n12761) );
  NAND3_X1 U19014 ( .A1(n14305), .A2(n60079), .A3(n43150), .ZN(n42571) );
  AOI21_X1 U11062 ( .A1(n65147), .A2(n43344), .B(n43054), .ZN(n5825) );
  OAI21_X1 U11081 ( .A1(n42058), .A2(n42896), .B(n4806), .ZN(n42061) );
  AOI21_X1 U11128 ( .A1(n43256), .A2(n44226), .B(n43992), .ZN(n20321) );
  NAND3_X1 U26133 ( .A1(n43977), .A2(n43710), .A3(n23314), .ZN(n21136) );
  NOR2_X1 U10674 ( .A1(n59650), .A2(n43068), .ZN(n43854) );
  NAND3_X1 U9314 ( .A1(n8654), .A2(n42196), .A3(n61739), .ZN(n8653) );
  OAI21_X1 U27619 ( .A1(n21140), .A2(n42310), .B(n42309), .ZN(n21139) );
  OAI21_X1 U23110 ( .A1(n20852), .A2(n20853), .B(n9792), .ZN(n58328) );
  NOR2_X1 U16544 ( .A1(n8192), .A2(n8191), .ZN(n8190) );
  NAND2_X1 U16705 ( .A1(n40546), .A2(n22500), .ZN(n41785) );
  NAND2_X1 U9293 ( .A1(n13202), .A2(n13200), .ZN(n43681) );
  NAND2_X1 U11095 ( .A1(n7033), .A2(n7032), .ZN(n39014) );
  INV_X1 U8642 ( .I(n20208), .ZN(n13866) );
  AOI22_X1 U20461 ( .A1(n41965), .A2(n2255), .B1(n41966), .B2(n2898), .ZN(
        n41967) );
  OAI21_X1 U31412 ( .A1(n42892), .A2(n60079), .B(n14305), .ZN(n42056) );
  NAND3_X1 U50187 ( .A1(n39089), .A2(n42185), .A3(n39088), .ZN(n39090) );
  INV_X1 U16531 ( .I(n42975), .ZN(n7819) );
  INV_X2 U37740 ( .I(n25638), .ZN(n44082) );
  OAI21_X1 U32651 ( .A1(n43510), .A2(n57281), .B(n1717), .ZN(n42046) );
  AOI21_X1 U16472 ( .A1(n42063), .A2(n42062), .B(n1940), .ZN(n1939) );
  NAND2_X1 U30707 ( .A1(n13866), .A2(n10160), .ZN(n13865) );
  NAND3_X1 U1491 ( .A1(n42055), .A2(n24895), .A3(n42056), .ZN(n9479) );
  NOR3_X1 U30798 ( .A1(n41344), .A2(n41343), .A3(n41342), .ZN(n41345) );
  NOR2_X1 U16524 ( .A1(n17398), .A2(n24623), .ZN(n17397) );
  NOR2_X1 U12789 ( .A1(n25537), .A2(n42997), .ZN(n7404) );
  NOR2_X1 U16530 ( .A1(n17559), .A2(n43509), .ZN(n43526) );
  INV_X2 U1428 ( .I(n20371), .ZN(n46558) );
  NAND2_X1 U47957 ( .A1(n21211), .A2(n21212), .ZN(n23256) );
  NOR3_X1 U25516 ( .A1(n16244), .A2(n21517), .A3(n20371), .ZN(n5839) );
  NAND3_X1 U22398 ( .A1(n42569), .A2(n42903), .A3(n42568), .ZN(n42577) );
  INV_X1 U24393 ( .I(n45041), .ZN(n15277) );
  AOI21_X1 U1435 ( .A1(n42680), .A2(n42679), .B(n42678), .ZN(n44541) );
  BUF_X2 U6076 ( .I(n20347), .Z(n10449) );
  INV_X1 U20772 ( .I(n44578), .ZN(n44957) );
  INV_X1 U10920 ( .I(n44592), .ZN(n46216) );
  INV_X1 U27761 ( .I(n7679), .ZN(n45045) );
  BUF_X2 U16426 ( .I(n46432), .Z(n24055) );
  NAND3_X1 U1398 ( .A1(n43820), .A2(n43819), .A3(n43818), .ZN(n44911) );
  BUF_X2 U1391 ( .I(n46701), .Z(n22212) );
  BUF_X2 U1397 ( .I(n13884), .Z(n13883) );
  BUF_X2 U12743 ( .I(n46213), .Z(n19226) );
  BUF_X2 U1390 ( .I(n12478), .Z(n12507) );
  CLKBUF_X2 U7023 ( .I(n9242), .Z(n61498) );
  CLKBUF_X2 U1401 ( .I(n25809), .Z(n14253) );
  BUF_X2 U1392 ( .I(n46493), .Z(n23953) );
  NAND2_X1 U33495 ( .A1(n15119), .A2(n16569), .ZN(n24090) );
  BUF_X2 U4551 ( .I(n46150), .Z(n23818) );
  BUF_X2 U10835 ( .I(n9477), .Z(n6872) );
  BUF_X2 U7994 ( .I(n18468), .Z(n14760) );
  BUF_X2 U6981 ( .I(n44723), .Z(n10536) );
  INV_X1 U1653 ( .I(n58127), .ZN(n5358) );
  INV_X1 U25312 ( .I(n46353), .ZN(n46507) );
  INV_X1 U37012 ( .I(n46433), .ZN(n46162) );
  INV_X1 U5245 ( .I(n44422), .ZN(n45325) );
  INV_X1 U1388 ( .I(n45246), .ZN(n45875) );
  INV_X2 U1364 ( .I(n59984), .ZN(n45136) );
  INV_X1 U9298 ( .I(n10278), .ZN(n46298) );
  INV_X1 U10866 ( .I(n5180), .ZN(n24401) );
  BUF_X2 U9982 ( .I(n45357), .Z(n23893) );
  BUF_X2 U11064 ( .I(n45326), .Z(n23426) );
  INV_X1 U12904 ( .I(n11852), .ZN(n15773) );
  INV_X1 U1383 ( .I(n13261), .ZN(n13313) );
  INV_X1 U16400 ( .I(n23987), .ZN(n1680) );
  BUF_X2 U11042 ( .I(n46691), .Z(n23618) );
  INV_X1 U31484 ( .I(n12872), .ZN(n46319) );
  BUF_X2 U43600 ( .I(n43774), .Z(n25530) );
  INV_X1 U13886 ( .I(n10678), .ZN(n12524) );
  INV_X1 U27874 ( .I(n8042), .ZN(n12265) );
  INV_X1 U32046 ( .I(n11858), .ZN(n43807) );
  INV_X1 U1359 ( .I(n46690), .ZN(n44223) );
  INV_X1 U51654 ( .I(n44478), .ZN(n45811) );
  INV_X1 U22629 ( .I(n7971), .ZN(n3941) );
  INV_X1 U1594 ( .I(n24992), .ZN(n673) );
  INV_X1 U10902 ( .I(n14900), .ZN(n15810) );
  INV_X1 U34091 ( .I(n15773), .ZN(n59619) );
  INV_X1 U1361 ( .I(n13313), .ZN(n46680) );
  INV_X1 U1570 ( .I(n57918), .ZN(n45047) );
  INV_X1 U4251 ( .I(n10098), .ZN(n17907) );
  INV_X1 U4470 ( .I(n14901), .ZN(n15734) );
  INV_X1 U1635 ( .I(n45401), .ZN(n46137) );
  INV_X1 U1336 ( .I(n43425), .ZN(n21316) );
  INV_X1 U16323 ( .I(n46210), .ZN(n12518) );
  INV_X1 U1592 ( .I(n8220), .ZN(n16932) );
  INV_X1 U9976 ( .I(n7506), .ZN(n44920) );
  INV_X4 U23256 ( .I(n4413), .ZN(n15697) );
  INV_X1 U43564 ( .I(n44944), .ZN(n25429) );
  INV_X2 U30573 ( .I(n24615), .ZN(n14323) );
  INV_X1 U31548 ( .I(n59296), .ZN(n24850) );
  INV_X1 U22262 ( .I(n47290), .ZN(n23186) );
  INV_X1 U34290 ( .I(n14888), .ZN(n47270) );
  INV_X1 U1296 ( .I(n46148), .ZN(n8683) );
  INV_X1 U1226 ( .I(n45551), .ZN(n47593) );
  INV_X8 U7805 ( .I(n9243), .ZN(n15757) );
  INV_X8 U30192 ( .I(n11443), .ZN(n13655) );
  INV_X8 U9279 ( .I(n10863), .ZN(n1294) );
  BUF_X2 U12699 ( .I(n1203), .Z(n22703) );
  INV_X1 U4819 ( .I(n15824), .ZN(n45076) );
  INV_X2 U6805 ( .I(n25896), .ZN(n23180) );
  NOR2_X1 U42754 ( .A1(n47252), .A2(n16020), .ZN(n60557) );
  INV_X1 U52069 ( .I(n44551), .ZN(n45718) );
  INV_X1 U3503 ( .I(n47617), .ZN(n45985) );
  CLKBUF_X2 U11045 ( .I(n10863), .Z(n195) );
  INV_X2 U38433 ( .I(n17452), .ZN(n48533) );
  NAND2_X1 U26021 ( .A1(n47717), .A2(n14473), .ZN(n6359) );
  INV_X2 U25116 ( .I(n63926), .ZN(n47530) );
  BUF_X2 U1507 ( .I(n20996), .Z(n60398) );
  INV_X2 U7823 ( .I(n23969), .ZN(n47575) );
  NAND2_X1 U52354 ( .A1(n23186), .A2(n22908), .ZN(n47280) );
  INV_X1 U1285 ( .I(n21090), .ZN(n1482) );
  NOR2_X1 U52035 ( .A1(n25004), .A2(n46897), .ZN(n44868) );
  INV_X2 U5049 ( .I(n3641), .ZN(n47295) );
  INV_X2 U12678 ( .I(n6934), .ZN(n20832) );
  INV_X1 U32917 ( .I(n45300), .ZN(n47683) );
  INV_X2 U11204 ( .I(n47407), .ZN(n47853) );
  INV_X1 U16193 ( .I(n47581), .ZN(n45978) );
  INV_X1 U17287 ( .I(n23666), .ZN(n57740) );
  INV_X1 U16284 ( .I(n45140), .ZN(n47275) );
  INV_X1 U12695 ( .I(n47501), .ZN(n1480) );
  INV_X1 U28127 ( .I(n47156), .ZN(n48484) );
  INV_X1 U43489 ( .I(n45576), .ZN(n47615) );
  INV_X1 U43325 ( .I(n44944), .ZN(n46017) );
  INV_X1 U1275 ( .I(n45905), .ZN(n1266) );
  INV_X1 U41011 ( .I(n22772), .ZN(n47592) );
  INV_X1 U25953 ( .I(n25444), .ZN(n44781) );
  INV_X2 U8157 ( .I(n2403), .ZN(n48588) );
  NAND2_X1 U52831 ( .A1(n16533), .A2(n48208), .ZN(n47196) );
  INV_X2 U39583 ( .I(n19160), .ZN(n26032) );
  NAND2_X1 U12664 ( .A1(n48588), .A2(n23542), .ZN(n8200) );
  NAND2_X1 U10973 ( .A1(n47825), .A2(n45964), .ZN(n59532) );
  INV_X1 U28790 ( .I(n47843), .ZN(n8692) );
  BUF_X2 U42218 ( .I(n47799), .Z(n23061) );
  NAND3_X1 U10967 ( .A1(n47827), .A2(n61025), .A3(n22386), .ZN(n45570) );
  BUF_X2 U4050 ( .I(n47884), .Z(n10225) );
  INV_X2 U9969 ( .I(n64548), .ZN(n47882) );
  INV_X1 U1191 ( .I(n12360), .ZN(n45935) );
  INV_X2 U9262 ( .I(n2973), .ZN(n47596) );
  NOR2_X1 U1163 ( .A1(n1064), .A2(n12825), .ZN(n12824) );
  BUF_X2 U5779 ( .I(n8225), .Z(n57603) );
  NAND3_X1 U7258 ( .A1(n46024), .A2(n12360), .A3(n46017), .ZN(n45647) );
  NAND2_X1 U11034 ( .A1(n2403), .A2(n59071), .ZN(n46468) );
  NOR2_X1 U1465 ( .A1(n47328), .A2(n5299), .ZN(n59818) );
  BUF_X2 U16257 ( .I(n16020), .Z(n47255) );
  NAND2_X1 U40860 ( .A1(n2564), .A2(n23167), .ZN(n45594) );
  NOR2_X1 U33487 ( .A1(n47505), .A2(n19569), .ZN(n47045) );
  INV_X2 U1306 ( .I(n16798), .ZN(n8842) );
  INV_X2 U11014 ( .I(n47881), .ZN(n1387) );
  NAND2_X1 U1232 ( .A1(n61714), .A2(n21090), .ZN(n46944) );
  NOR2_X1 U28466 ( .A1(n23666), .A2(n47421), .ZN(n47411) );
  INV_X1 U21364 ( .I(n2944), .ZN(n7799) );
  INV_X2 U6637 ( .I(n45498), .ZN(n1080) );
  INV_X1 U1443 ( .I(n1267), .ZN(n59892) );
  INV_X1 U28872 ( .I(n65074), .ZN(n45225) );
  INV_X2 U16296 ( .I(n47518), .ZN(n47502) );
  NOR2_X1 U27185 ( .A1(n57740), .A2(n45267), .ZN(n47414) );
  INV_X1 U10976 ( .I(n47084), .ZN(n1479) );
  INV_X1 U34089 ( .I(n47826), .ZN(n45566) );
  INV_X1 U16194 ( .I(n3942), .ZN(n25066) );
  NAND3_X1 U1228 ( .A1(n48518), .A2(n48511), .A3(n23416), .ZN(n48632) );
  NAND2_X1 U1230 ( .A1(n47472), .A2(n9256), .ZN(n8152) );
  INV_X1 U1321 ( .I(n21755), .ZN(n47035) );
  INV_X1 U28051 ( .I(n45682), .ZN(n45979) );
  INV_X2 U26184 ( .I(n48095), .ZN(n16950) );
  NAND2_X1 U42553 ( .A1(n46039), .A2(n46033), .ZN(n45486) );
  INV_X1 U21685 ( .I(n6497), .ZN(n19715) );
  INV_X2 U8623 ( .I(n59523), .ZN(n1263) );
  INV_X1 U34285 ( .I(n25689), .ZN(n48487) );
  INV_X1 U1483 ( .I(n47245), .ZN(n22303) );
  INV_X1 U16183 ( .I(n25702), .ZN(n47282) );
  NAND2_X1 U40400 ( .A1(n1666), .A2(n1484), .ZN(n46027) );
  INV_X1 U4998 ( .I(n24558), .ZN(n21976) );
  INV_X1 U11011 ( .I(n47579), .ZN(n47288) );
  INV_X1 U1243 ( .I(n47197), .ZN(n18787) );
  INV_X1 U43200 ( .I(n47244), .ZN(n47621) );
  BUF_X8 U41624 ( .I(n46382), .Z(n48460) );
  INV_X1 U52701 ( .I(n47119), .ZN(n45887) );
  INV_X2 U1256 ( .I(n46106), .ZN(n48659) );
  NAND2_X1 U33837 ( .A1(n45716), .A2(n46033), .ZN(n14300) );
  INV_X2 U1432 ( .I(n48135), .ZN(n48472) );
  INV_X2 U4523 ( .I(n47851), .ZN(n24893) );
  INV_X2 U23444 ( .I(n48460), .ZN(n48134) );
  INV_X2 U27989 ( .I(n7931), .ZN(n47386) );
  NOR2_X1 U1314 ( .A1(n47880), .A2(n14473), .ZN(n14472) );
  INV_X1 U38045 ( .I(n48199), .ZN(n16718) );
  NAND2_X1 U22496 ( .A1(n1080), .A2(n6034), .ZN(n60347) );
  NAND3_X1 U37137 ( .A1(n48665), .A2(n48208), .A3(n23661), .ZN(n18551) );
  NOR2_X1 U16186 ( .A1(n8692), .A2(n9860), .ZN(n8691) );
  BUF_X2 U20455 ( .I(n9758), .Z(n58009) );
  OAI21_X1 U53206 ( .A1(n12993), .A2(n7335), .B(n48254), .ZN(n47219) );
  NOR2_X1 U33621 ( .A1(n45961), .A2(n10088), .ZN(n45561) );
  NAND2_X1 U21427 ( .A1(n47282), .A2(n2973), .ZN(n45684) );
  BUF_X2 U34578 ( .I(n46919), .Z(n59687) );
  AOI21_X1 U12645 ( .A1(n14121), .A2(n47717), .B(n47886), .ZN(n9452) );
  NOR2_X1 U39200 ( .A1(n20031), .A2(n18590), .ZN(n46730) );
  NAND3_X1 U16138 ( .A1(n45673), .A2(n45674), .A3(n47262), .ZN(n45675) );
  INV_X2 U16090 ( .I(n21177), .ZN(n48529) );
  NAND3_X1 U52702 ( .A1(n45887), .A2(n23617), .A3(n24113), .ZN(n45888) );
  NAND2_X1 U37060 ( .A1(n18570), .A2(n16533), .ZN(n46997) );
  NAND2_X1 U7236 ( .A1(n1652), .A2(n3510), .ZN(n8582) );
  CLKBUF_X2 U5733 ( .I(n2026), .Z(n58033) );
  INV_X1 U31332 ( .I(n16974), .ZN(n45784) );
  AOI21_X1 U8296 ( .A1(n6497), .A2(n10193), .B(n46943), .ZN(n47984) );
  INV_X1 U10975 ( .I(n47839), .ZN(n47559) );
  INV_X1 U25108 ( .I(n8047), .ZN(n18766) );
  INV_X2 U33763 ( .I(n45964), .ZN(n47820) );
  NAND2_X1 U53222 ( .A1(n47302), .A2(n47301), .ZN(n47303) );
  INV_X2 U31566 ( .I(n11183), .ZN(n46863) );
  INV_X1 U1144 ( .I(n47432), .ZN(n47437) );
  CLKBUF_X2 U5715 ( .I(n2403), .Z(n58974) );
  CLKBUF_X2 U25079 ( .I(n20514), .Z(n58636) );
  NAND2_X1 U51658 ( .A1(n47886), .A2(n43596), .ZN(n47366) );
  NAND2_X1 U9963 ( .A1(n47542), .A2(n25481), .ZN(n25480) );
  BUF_X2 U10999 ( .I(n9140), .Z(n3340) );
  NAND2_X1 U4400 ( .A1(n3597), .A2(n6730), .ZN(n47864) );
  NOR2_X1 U52844 ( .A1(n48205), .A2(n48209), .ZN(n46995) );
  NAND2_X1 U31960 ( .A1(n47180), .A2(n25481), .ZN(n48619) );
  NAND2_X1 U12644 ( .A1(n14120), .A2(n47726), .ZN(n47365) );
  NAND2_X1 U37025 ( .A1(n6957), .A2(n46106), .ZN(n48652) );
  INV_X2 U1095 ( .I(n47262), .ZN(n45672) );
  INV_X2 U42624 ( .I(n47208), .ZN(n48136) );
  NAND2_X1 U42356 ( .A1(n47186), .A2(n19921), .ZN(n48540) );
  NAND2_X1 U30834 ( .A1(n45566), .A2(n23894), .ZN(n43191) );
  NAND3_X1 U24610 ( .A1(n22326), .A2(n46914), .A3(n25444), .ZN(n44194) );
  NAND2_X1 U1117 ( .A1(n43192), .A2(n3510), .ZN(n47823) );
  CLKBUF_X2 U5788 ( .I(n25866), .Z(n57852) );
  NAND2_X1 U1170 ( .A1(n3365), .A2(n44770), .ZN(n47481) );
  INV_X1 U1399 ( .I(n6081), .ZN(n59821) );
  INV_X2 U10980 ( .I(n637), .ZN(n47857) );
  INV_X1 U47941 ( .I(n46911), .ZN(n5225) );
  NAND2_X1 U53474 ( .A1(n48503), .A2(n48511), .ZN(n48261) );
  INV_X1 U32494 ( .I(n45436), .ZN(n47144) );
  INV_X1 U1149 ( .I(n64250), .ZN(n47232) );
  NOR2_X1 U31078 ( .A1(n59419), .A2(n47255), .ZN(n45670) );
  INV_X1 U16093 ( .I(n63913), .ZN(n47202) );
  INV_X1 U17286 ( .I(n47688), .ZN(n1649) );
  NAND2_X1 U52300 ( .A1(n46927), .A2(n5299), .ZN(n47325) );
  NOR2_X1 U28611 ( .A1(n9730), .A2(n47263), .ZN(n45663) );
  NOR2_X1 U11055 ( .A1(n4086), .A2(n47774), .ZN(n46858) );
  INV_X1 U1237 ( .I(n45482), .ZN(n1647) );
  INV_X1 U11175 ( .I(n22255), .ZN(n48236) );
  INV_X1 U20347 ( .I(n2179), .ZN(n47806) );
  INV_X1 U1182 ( .I(n13356), .ZN(n47574) );
  INV_X1 U16014 ( .I(n45594), .ZN(n47906) );
  INV_X1 U1143 ( .I(n15421), .ZN(n18980) );
  NAND2_X1 U52641 ( .A1(n46950), .A2(n1328), .ZN(n45758) );
  INV_X1 U16173 ( .I(n10397), .ZN(n47690) );
  INV_X1 U32341 ( .I(n23606), .ZN(n59406) );
  INV_X1 U1142 ( .I(n46943), .ZN(n47228) );
  INV_X1 U1135 ( .I(n26032), .ZN(n48543) );
  INV_X1 U26678 ( .I(n46013), .ZN(n47299) );
  INV_X1 U5640 ( .I(n18100), .ZN(n48145) );
  INV_X1 U7829 ( .I(n17128), .ZN(n5554) );
  INV_X2 U21390 ( .I(n46813), .ZN(n12698) );
  OAI21_X1 U8603 ( .A1(n16950), .A2(n15728), .B(n6805), .ZN(n47112) );
  NAND2_X1 U4920 ( .A1(n10624), .A2(n23617), .ZN(n45891) );
  NOR2_X1 U9268 ( .A1(n2973), .A2(n47579), .ZN(n47272) );
  NAND3_X1 U24817 ( .A1(n15076), .A2(n45503), .A3(n59406), .ZN(n59652) );
  NAND2_X1 U24598 ( .A1(n5705), .A2(n21178), .ZN(n58934) );
  OAI21_X1 U26194 ( .A1(n11813), .A2(n47273), .B(n6523), .ZN(n47287) );
  OAI22_X1 U29841 ( .A1(n47000), .A2(n17153), .B1(n48652), .B2(n48654), .ZN(
        n46107) );
  NAND2_X1 U53253 ( .A1(n1266), .A2(n7395), .ZN(n47397) );
  OAI21_X1 U16061 ( .A1(n45487), .A2(n13566), .B(n46858), .ZN(n45488) );
  NAND2_X1 U35172 ( .A1(n48530), .A2(n17905), .ZN(n18118) );
  INV_X1 U3721 ( .I(n47864), .ZN(n43831) );
  NAND2_X1 U53243 ( .A1(n47368), .A2(n47367), .ZN(n47369) );
  NOR2_X1 U1128 ( .A1(n47494), .A2(n16493), .ZN(n13072) );
  NOR2_X1 U37045 ( .A1(n47325), .A2(n45619), .ZN(n45958) );
  NOR2_X1 U21502 ( .A1(n48644), .A2(n48511), .ZN(n48512) );
  NAND3_X1 U15952 ( .A1(n45901), .A2(n13782), .A3(n3597), .ZN(n45902) );
  NOR2_X1 U16001 ( .A1(n47823), .A2(n47820), .ZN(n2315) );
  NAND2_X1 U12618 ( .A1(n5934), .A2(n47255), .ZN(n45665) );
  NAND3_X1 U1299 ( .A1(n16162), .A2(n47906), .A3(n47576), .ZN(n45942) );
  NAND2_X1 U8598 ( .A1(n47272), .A2(n45978), .ZN(n47588) );
  NAND2_X1 U22632 ( .A1(n45785), .A2(n3942), .ZN(n47025) );
  NAND2_X1 U33961 ( .A1(n14472), .A2(n47886), .ZN(n47877) );
  INV_X2 U30577 ( .I(n48552), .ZN(n21445) );
  NAND2_X1 U9266 ( .A1(n47494), .A2(n65275), .ZN(n11808) );
  NOR2_X1 U12620 ( .A1(n45672), .A2(n63734), .ZN(n44485) );
  NOR2_X1 U1354 ( .A1(n7050), .A2(n62748), .ZN(n45223) );
  NAND2_X1 U53588 ( .A1(n48642), .A2(n48518), .ZN(n48520) );
  NAND2_X1 U23751 ( .A1(n47772), .A2(n11183), .ZN(n20425) );
  OAI21_X1 U12627 ( .A1(n62755), .A2(n3686), .B(n65062), .ZN(n12699) );
  OAI21_X1 U1427 ( .A1(n17572), .A2(n45567), .B(n45566), .ZN(n17571) );
  NAND2_X1 U53247 ( .A1(n47386), .A2(n47803), .ZN(n47388) );
  CLKBUF_X2 U12682 ( .I(n46959), .Z(n6786) );
  NAND2_X1 U10955 ( .A1(n44284), .A2(n65275), .ZN(n44674) );
  NOR2_X1 U7842 ( .A1(n46919), .A2(n2944), .ZN(n2786) );
  AOI21_X1 U53200 ( .A1(n48460), .A2(n14520), .B(n47206), .ZN(n48124) );
  NOR2_X1 U1159 ( .A1(n22255), .A2(n47186), .ZN(n47190) );
  NAND2_X1 U22299 ( .A1(n12203), .A2(n3663), .ZN(n47817) );
  NAND2_X1 U1127 ( .A1(n48203), .A2(n12482), .ZN(n7436) );
  INV_X2 U32493 ( .I(n15825), .ZN(n47382) );
  NAND2_X1 U5318 ( .A1(n20031), .A2(n18138), .ZN(n47431) );
  NAND3_X1 U1357 ( .A1(n24113), .A2(n57398), .A3(n48561), .ZN(n48576) );
  INV_X1 U10960 ( .I(n47489), .ZN(n13759) );
  INV_X2 U28804 ( .I(n8732), .ZN(n49862) );
  CLKBUF_X2 U33210 ( .I(n47415), .Z(n59528) );
  INV_X1 U52601 ( .I(n46028), .ZN(n46864) );
  OR2_X1 U1099 ( .A1(n12546), .A2(n21304), .Z(n48094) );
  INV_X1 U43419 ( .I(n22700), .ZN(n46739) );
  AND2_X1 U31163 ( .A1(n15728), .A2(n46813), .Z(n12700) );
  NAND2_X1 U52500 ( .A1(n47737), .A2(n47437), .ZN(n45452) );
  NAND2_X1 U5724 ( .A1(n25895), .A2(n7931), .ZN(n47802) );
  INV_X1 U1078 ( .I(n19200), .ZN(n23018) );
  NOR2_X1 U9269 ( .A1(n16950), .A2(n23099), .ZN(n46758) );
  INV_X1 U16182 ( .I(n838), .ZN(n47845) );
  INV_X1 U22792 ( .I(n4090), .ZN(n5246) );
  INV_X1 U12683 ( .I(n46016), .ZN(n4214) );
  INV_X1 U5028 ( .I(n24578), .ZN(n46875) );
  NAND2_X1 U37064 ( .A1(n48511), .A2(n48521), .ZN(n48636) );
  NAND2_X1 U15969 ( .A1(n20140), .A2(n46817), .ZN(n13053) );
  OAI22_X1 U28119 ( .A1(n1064), .A2(n8040), .B1(n47494), .B2(n12850), .ZN(
        n44283) );
  OAI21_X1 U25703 ( .A1(n58244), .A2(n57839), .B(n45504), .ZN(n6651) );
  NAND3_X1 U7232 ( .A1(n21102), .A2(n47368), .A3(n45807), .ZN(n22394) );
  OAI21_X1 U12577 ( .A1(n58889), .A2(n47691), .B(n46840), .ZN(n14268) );
  NAND3_X1 U9948 ( .A1(n47190), .A2(n22464), .A3(n17905), .ZN(n48119) );
  AOI21_X1 U5580 ( .A1(n45762), .A2(n57731), .B(n1646), .ZN(n6281) );
  NAND3_X1 U53761 ( .A1(n48262), .A2(n48260), .A3(n48261), .ZN(n61176) );
  NAND3_X1 U12573 ( .A1(n10405), .A2(n59216), .A3(n45901), .ZN(n9726) );
  AOI22_X1 U11266 ( .A1(n47633), .A2(n47885), .B1(n47886), .B2(n47875), .ZN(
        n47640) );
  AOI21_X1 U1049 ( .A1(n13566), .A2(n45486), .B(n12597), .ZN(n16093) );
  OAI21_X1 U53251 ( .A1(n47391), .A2(n47390), .B(n47803), .ZN(n47393) );
  AOI22_X1 U22741 ( .A1(n44654), .A2(n47228), .B1(n22389), .B2(n44655), .ZN(
        n58299) );
  OAI21_X1 U12624 ( .A1(n1328), .A2(n63878), .B(n46959), .ZN(n46960) );
  OAI21_X1 U41392 ( .A1(n21954), .A2(n49862), .B(n20878), .ZN(n47135) );
  INV_X1 U6787 ( .I(n62220), .ZN(n57205) );
  NAND2_X1 U16211 ( .A1(n3340), .A2(n571), .ZN(n48608) );
  AOI21_X1 U12543 ( .A1(n8156), .A2(n64969), .B(n8153), .ZN(n47478) );
  NAND2_X1 U22570 ( .A1(n5721), .A2(n22389), .ZN(n59949) );
  NAND3_X1 U52562 ( .A1(n45588), .A2(n45587), .A3(n45586), .ZN(n45589) );
  INV_X1 U53271 ( .I(n47463), .ZN(n47479) );
  OAI22_X1 U15907 ( .A1(n5466), .A2(n11928), .B1(n47845), .B2(n5464), .ZN(
        n11927) );
  NAND2_X1 U33370 ( .A1(n13566), .A2(n20426), .ZN(n46867) );
  NOR2_X1 U34596 ( .A1(n15336), .A2(n46739), .ZN(n46744) );
  NOR2_X1 U1043 ( .A1(n45506), .A2(n46958), .ZN(n46074) );
  NOR2_X1 U21937 ( .A1(n46977), .A2(n4380), .ZN(n46984) );
  OR2_X1 U5617 ( .A1(n25691), .A2(n47464), .Z(n9170) );
  AOI21_X1 U1077 ( .A1(n47857), .A2(n70), .B(n11599), .ZN(n47399) );
  OR2_X1 U1282 ( .A1(n3716), .A2(n45619), .Z(n46062) );
  INV_X1 U29839 ( .I(n63710), .ZN(n11699) );
  NAND2_X1 U26191 ( .A1(n6523), .A2(n61967), .ZN(n16509) );
  AOI21_X1 U4238 ( .A1(n15295), .A2(n18757), .B(n46995), .ZN(n17005) );
  OAI21_X1 U10911 ( .A1(n49863), .A2(n49860), .B(n49862), .ZN(n48115) );
  OAI22_X1 U25479 ( .A1(n18047), .A2(n47900), .B1(n47568), .B2(n47896), .ZN(
        n2610) );
  AOI21_X1 U33371 ( .A1(n13566), .A2(n64654), .B(n4086), .ZN(n44557) );
  NAND4_X1 U7254 ( .A1(n47863), .A2(n43827), .A3(n43828), .A4(n24893), .ZN(
        n4093) );
  AOI22_X1 U26814 ( .A1(n44197), .A2(n44196), .B1(n46916), .B2(n44195), .ZN(
        n44198) );
  NAND4_X1 U4009 ( .A1(n323), .A2(n48144), .A3(n48157), .A4(n48553), .ZN(
        n46797) );
  OAI21_X1 U1052 ( .A1(n61863), .A2(n11343), .B(n47101), .ZN(n11342) );
  NAND3_X1 U15744 ( .A1(n47024), .A2(n10572), .A3(n47023), .ZN(n10571) );
  NAND2_X1 U43499 ( .A1(n47837), .A2(n45550), .ZN(n25283) );
  NAND2_X1 U6736 ( .A1(n47408), .A2(n70), .ZN(n58258) );
  NAND2_X1 U52660 ( .A1(n47426), .A2(n47418), .ZN(n45799) );
  OAI21_X1 U37091 ( .A1(n42618), .A2(n11929), .B(n47828), .ZN(n22213) );
  AOI22_X1 U9925 ( .A1(n47046), .A2(n22899), .B1(n61014), .B2(n47047), .ZN(
        n17806) );
  NAND2_X1 U52579 ( .A1(n46062), .A2(n45620), .ZN(n45627) );
  NOR2_X1 U16056 ( .A1(n47027), .A2(n45780), .ZN(n45790) );
  AOI22_X1 U1266 ( .A1(n48515), .A2(n20624), .B1(n48517), .B2(n48516), .ZN(
        n48524) );
  AOI21_X1 U12571 ( .A1(n46717), .A2(n15903), .B(n48238), .ZN(n18631) );
  OAI21_X1 U23689 ( .A1(n46960), .A2(n46961), .B(n58033), .ZN(n46962) );
  AOI21_X1 U6752 ( .A1(n57544), .A2(n65095), .B(n45937), .ZN(n45939) );
  NAND2_X1 U25176 ( .A1(n13802), .A2(n16183), .ZN(n20019) );
  NOR2_X1 U24348 ( .A1(n58521), .A2(n24430), .ZN(n21290) );
  NAND3_X1 U16092 ( .A1(n45733), .A2(n45737), .A3(n58445), .ZN(n12325) );
  NOR2_X1 U8582 ( .A1(n13970), .A2(n1295), .ZN(n13969) );
  NAND2_X1 U52071 ( .A1(n44553), .A2(n44552), .ZN(n47776) );
  NOR2_X1 U52438 ( .A1(n47386), .A2(n45308), .ZN(n47708) );
  NAND2_X1 U10899 ( .A1(n44000), .A2(n45203), .ZN(n15265) );
  INV_X2 U11487 ( .I(n23514), .ZN(n3596) );
  NAND2_X1 U52926 ( .A1(n47175), .A2(n47542), .ZN(n47540) );
  AND4_X1 U1008 ( .A1(n46078), .A2(n47259), .A3(n47261), .A4(n44486), .Z(
        n44487) );
  NAND4_X1 U53289 ( .A1(n47540), .A2(n48616), .A3(n48629), .A4(n47539), .ZN(
        n47553) );
  AOI21_X1 U55863 ( .A1(n19774), .A2(n20624), .B(n48635), .ZN(n17079) );
  AOI22_X1 U1235 ( .A1(n58639), .A2(n9299), .B1(n46981), .B2(n46980), .ZN(
        n7741) );
  OAI21_X1 U15827 ( .A1(n13041), .A2(n17805), .B(n13040), .ZN(n13039) );
  NAND2_X1 U10881 ( .A1(n2610), .A2(n47578), .ZN(n2609) );
  NAND2_X1 U8050 ( .A1(n18590), .A2(n64096), .ZN(n11821) );
  OAI21_X1 U1054 ( .A1(n48597), .A2(n48596), .B(n48595), .ZN(n14371) );
  NOR2_X1 U1183 ( .A1(n61205), .A2(n61204), .ZN(n61203) );
  NAND4_X1 U1019 ( .A1(n19988), .A2(n45518), .A3(n19987), .A4(n10184), .ZN(
        n45526) );
  NAND3_X1 U35570 ( .A1(n25864), .A2(n25861), .A3(n45799), .ZN(n25860) );
  BUF_X4 U6693 ( .I(n48414), .Z(n57204) );
  NAND3_X1 U22796 ( .A1(n4093), .A2(n4092), .A3(n4091), .ZN(n17629) );
  NOR2_X1 U42711 ( .A1(n60825), .A2(n57399), .ZN(n60549) );
  INV_X2 U8178 ( .I(n12988), .ZN(n50346) );
  INV_X2 U26621 ( .I(n49226), .ZN(n49465) );
  INV_X1 U21998 ( .I(n61716), .ZN(n58206) );
  INV_X1 U32135 ( .I(n16815), .ZN(n12003) );
  INV_X2 U20226 ( .I(n5587), .ZN(n6313) );
  BUF_X8 U42420 ( .I(n47480), .Z(n48847) );
  AOI21_X1 U8587 ( .A1(n14371), .A2(n48601), .B(n14366), .ZN(n14365) );
  INV_X2 U31622 ( .I(n47646), .ZN(n18252) );
  NAND2_X1 U15497 ( .A1(n3771), .A2(n16379), .ZN(n7454) );
  BUF_X2 U5141 ( .I(n7846), .Z(n7336) );
  CLKBUF_X2 U1173 ( .I(n49486), .Z(n15724) );
  BUF_X4 U1113 ( .I(n58297), .Z(n57735) );
  BUF_X2 U12495 ( .I(n23514), .Z(n2433) );
  BUF_X4 U42701 ( .I(n48322), .Z(n23738) );
  NAND2_X1 U969 ( .A1(n47970), .A2(n57204), .ZN(n47964) );
  NAND2_X1 U23151 ( .A1(n47093), .A2(n47094), .ZN(n47108) );
  BUF_X4 U29909 ( .I(n45662), .Z(n49063) );
  INV_X2 U4183 ( .I(n26000), .ZN(n9346) );
  INV_X1 U38518 ( .I(n49486), .ZN(n17334) );
  INV_X1 U22667 ( .I(n49053), .ZN(n47920) );
  INV_X1 U10863 ( .I(n49500), .ZN(n9594) );
  INV_X2 U13567 ( .I(n16963), .ZN(n48341) );
  INV_X4 U855 ( .I(n1209), .ZN(n15550) );
  INV_X2 U964 ( .I(n47347), .ZN(n24209) );
  AOI21_X1 U20725 ( .A1(n2477), .A2(n49842), .B(n16379), .ZN(n21526) );
  INV_X1 U12456 ( .I(n6341), .ZN(n17126) );
  NAND2_X1 U38030 ( .A1(n59633), .A2(n9772), .ZN(n49998) );
  NOR2_X1 U4062 ( .A1(n14931), .A2(n16765), .ZN(n339) );
  BUF_X4 U9890 ( .I(n6654), .Z(n10563) );
  BUF_X2 U35567 ( .I(n50236), .Z(n17885) );
  NAND2_X1 U25967 ( .A1(n49459), .A2(n6314), .ZN(n49150) );
  INV_X2 U15740 ( .I(n49803), .ZN(n1642) );
  INV_X2 U43623 ( .I(n49783), .ZN(n47977) );
  BUF_X2 U5425 ( .I(n50360), .Z(n260) );
  INV_X2 U971 ( .I(n49792), .ZN(n49114) );
  NAND2_X1 U42663 ( .A1(n24134), .A2(n50004), .ZN(n50354) );
  INV_X2 U13321 ( .I(n50406), .ZN(n25944) );
  INV_X2 U950 ( .I(n6243), .ZN(n23238) );
  INV_X2 U12504 ( .I(n15741), .ZN(n1471) );
  INV_X2 U10886 ( .I(n50283), .ZN(n1384) );
  INV_X2 U4463 ( .I(n48362), .ZN(n49283) );
  INV_X2 U15729 ( .I(n48411), .ZN(n1640) );
  CLKBUF_X2 U5691 ( .I(n22962), .Z(n2357) );
  INV_X2 U31047 ( .I(n15386), .ZN(n50093) );
  INV_X2 U990 ( .I(n12646), .ZN(n15753) );
  INV_X1 U15709 ( .I(n12003), .ZN(n10874) );
  INV_X2 U22884 ( .I(n49732), .ZN(n4174) );
  NAND2_X1 U11445 ( .A1(n50142), .A2(n22717), .ZN(n49655) );
  NOR2_X1 U30225 ( .A1(n7738), .A2(n15724), .ZN(n48391) );
  INV_X2 U26073 ( .I(n8994), .ZN(n50407) );
  INV_X1 U951 ( .I(n18502), .ZN(n20428) );
  INV_X2 U21760 ( .I(n9164), .ZN(n49411) );
  NAND2_X1 U1108 ( .A1(n21870), .A2(n50340), .ZN(n57995) );
  INV_X2 U5280 ( .I(n5498), .ZN(n49677) );
  INV_X1 U955 ( .I(n15595), .ZN(n49374) );
  INV_X1 U983 ( .I(n23247), .ZN(n1638) );
  INV_X1 U1114 ( .I(n21205), .ZN(n50221) );
  NAND2_X1 U8074 ( .A1(n1205), .A2(n16595), .ZN(n8887) );
  NAND2_X1 U881 ( .A1(n57204), .A2(n23156), .ZN(n48419) );
  INV_X1 U32553 ( .I(n49493), .ZN(n17335) );
  INV_X1 U4321 ( .I(n64416), .ZN(n1291) );
  INV_X2 U10851 ( .I(n49842), .ZN(n49452) );
  INV_X1 U7545 ( .I(n2810), .ZN(n49055) );
  INV_X2 U963 ( .I(n49929), .ZN(n24692) );
  INV_X1 U7242 ( .I(n49630), .ZN(n3738) );
  BUF_X8 U15710 ( .I(n48527), .Z(n3055) );
  NOR2_X1 U4163 ( .A1(n13440), .A2(n50041), .ZN(n3338) );
  NAND2_X1 U9908 ( .A1(n19756), .A2(n57610), .ZN(n49743) );
  INV_X8 U5274 ( .I(n11153), .ZN(n58645) );
  BUF_X8 U1112 ( .I(n49990), .Z(n60209) );
  INV_X1 U12420 ( .I(n48999), .ZN(n49609) );
  NAND2_X1 U53439 ( .A1(n18975), .A2(n58907), .ZN(n48021) );
  NAND3_X1 U35519 ( .A1(n50092), .A2(n50093), .A3(n50374), .ZN(n22038) );
  NOR2_X1 U15614 ( .A1(n12701), .A2(n9177), .ZN(n49494) );
  NOR2_X1 U42019 ( .A1(n49702), .A2(n48349), .ZN(n45161) );
  INV_X1 U8557 ( .I(n45171), .ZN(n2157) );
  AOI21_X1 U32064 ( .A1(n50123), .A2(n1384), .B(n1224), .ZN(n14833) );
  AOI21_X1 U33964 ( .A1(n49377), .A2(n58983), .B(n49538), .ZN(n49378) );
  NOR2_X1 U6404 ( .A1(n49075), .A2(n49074), .ZN(n48301) );
  INV_X1 U55565 ( .I(n13988), .ZN(n61311) );
  NOR2_X1 U25123 ( .A1(n49089), .A2(n49674), .ZN(n5428) );
  CLKBUF_X2 U6743 ( .I(n50283), .Z(n60487) );
  NOR2_X1 U37174 ( .A1(n13038), .A2(n48847), .ZN(n49520) );
  INV_X1 U30564 ( .I(n48039), .ZN(n48448) );
  BUF_X2 U9899 ( .I(n64416), .Z(n7098) );
  OAI21_X1 U25185 ( .A1(n5517), .A2(n13839), .B(n58037), .ZN(n47789) );
  NOR2_X1 U12457 ( .A1(n48377), .A2(n20055), .ZN(n49453) );
  NAND2_X1 U935 ( .A1(n49908), .A2(n14315), .ZN(n6028) );
  INV_X2 U885 ( .I(n50340), .ZN(n49868) );
  NOR2_X1 U880 ( .A1(n49283), .A2(n49276), .ZN(n48917) );
  CLKBUF_X2 U15602 ( .I(n49792), .Z(n20708) );
  BUF_X2 U12478 ( .I(n18502), .Z(n1637) );
  NAND3_X1 U831 ( .A1(n1468), .A2(n7990), .A3(n49063), .ZN(n49073) );
  INV_X2 U57197 ( .I(n49384), .ZN(n49323) );
  INV_X2 U10883 ( .I(n49538), .ZN(n1382) );
  NAND2_X1 U21665 ( .A1(n23063), .A2(n78), .ZN(n49255) );
  NAND2_X1 U842 ( .A1(n8129), .A2(n49318), .ZN(n49597) );
  NOR2_X1 U5920 ( .A1(n24821), .A2(n3694), .ZN(n49515) );
  NAND2_X1 U952 ( .A1(n1468), .A2(n7990), .ZN(n20460) );
  NOR2_X1 U26936 ( .A1(n16963), .A2(n14315), .ZN(n48737) );
  NOR2_X1 U29920 ( .A1(n23156), .A2(n1640), .ZN(n48825) );
  NAND2_X1 U24717 ( .A1(n62795), .A2(n4526), .ZN(n48030) );
  NAND2_X1 U825 ( .A1(n49114), .A2(n49803), .ZN(n49115) );
  NAND2_X1 U34385 ( .A1(n49673), .A2(n47646), .ZN(n49371) );
  CLKBUF_X2 U24157 ( .I(n20004), .Z(n58856) );
  INV_X2 U33345 ( .I(n50220), .ZN(n50216) );
  INV_X1 U8565 ( .I(n49937), .ZN(n50262) );
  OAI21_X1 U10868 ( .A1(n3031), .A2(n23707), .B(n49720), .ZN(n50094) );
  NAND2_X1 U41828 ( .A1(n44004), .A2(n359), .ZN(n43757) );
  NAND2_X1 U924 ( .A1(n18252), .A2(n4780), .ZN(n49686) );
  NAND2_X1 U32912 ( .A1(n1471), .A2(n50283), .ZN(n50287) );
  NAND2_X1 U25897 ( .A1(n20458), .A2(n65135), .ZN(n6244) );
  INV_X1 U43851 ( .I(n49065), .ZN(n48299) );
  NAND2_X1 U37526 ( .A1(n1956), .A2(n49940), .ZN(n13118) );
  INV_X1 U15763 ( .I(n49701), .ZN(n49757) );
  OR2_X1 U23633 ( .A1(n8044), .A2(n57204), .Z(n48413) );
  OR2_X1 U21582 ( .A1(n25233), .A2(n50283), .Z(n48721) );
  NAND2_X1 U4648 ( .A1(n61624), .A2(n15550), .ZN(n49947) );
  INV_X1 U5226 ( .I(n49462), .ZN(n49221) );
  AND2_X1 U5641 ( .A1(n49701), .A2(n22819), .Z(n15737) );
  OR2_X1 U55509 ( .A1(n15741), .A2(n23533), .Z(n22867) );
  OR2_X1 U5624 ( .A1(n23247), .A2(n25320), .Z(n10941) );
  INV_X1 U10831 ( .I(n15436), .ZN(n50060) );
  INV_X1 U11678 ( .I(n57473), .ZN(n49096) );
  NAND2_X1 U3924 ( .A1(n49063), .A2(n49076), .ZN(n21334) );
  NOR2_X1 U4202 ( .A1(n48678), .A2(n49702), .ZN(n49697) );
  CLKBUF_X2 U37864 ( .I(n7952), .Z(n60397) );
  INV_X1 U10860 ( .I(n49986), .ZN(n49989) );
  INV_X1 U25062 ( .I(n49319), .ZN(n49602) );
  INV_X1 U10857 ( .I(n9177), .ZN(n19042) );
  NOR2_X1 U6199 ( .A1(n49019), .A2(n9853), .ZN(n12037) );
  NOR2_X1 U53396 ( .A1(n61741), .A2(n49529), .ZN(n47916) );
  INV_X1 U15521 ( .I(n49597), .ZN(n49601) );
  NOR2_X1 U12395 ( .A1(n49634), .A2(n1629), .ZN(n7243) );
  NAND3_X1 U40514 ( .A1(n6341), .A2(n58206), .A3(n16379), .ZN(n48972) );
  NAND2_X1 U12419 ( .A1(n57949), .A2(n1376), .ZN(n49385) );
  INV_X1 U6307 ( .I(n48859), .ZN(n9354) );
  NOR3_X1 U27550 ( .A1(n48434), .A2(n7271), .A3(n47941), .ZN(n49112) );
  NOR2_X1 U9222 ( .A1(n25944), .A2(n58840), .ZN(n46727) );
  NAND3_X1 U27308 ( .A1(n49283), .A2(n49287), .A3(n49276), .ZN(n48360) );
  NAND2_X1 U36182 ( .A1(n9177), .A2(n6704), .ZN(n48855) );
  NAND2_X1 U31073 ( .A1(n49377), .A2(n49543), .ZN(n18817) );
  INV_X1 U11557 ( .I(n18833), .ZN(n57884) );
  NAND2_X1 U52543 ( .A1(n57204), .A2(n7115), .ZN(n48416) );
  INV_X1 U4516 ( .I(n19003), .ZN(n11170) );
  INV_X1 U24339 ( .I(n48046), .ZN(n48051) );
  NAND2_X1 U7269 ( .A1(n48366), .A2(n57425), .ZN(n9306) );
  NAND2_X1 U11316 ( .A1(n21870), .A2(n49868), .ZN(n21479) );
  NAND2_X1 U1105 ( .A1(n1382), .A2(n10422), .ZN(n18821) );
  INV_X1 U41566 ( .I(n50342), .ZN(n49969) );
  NAND2_X1 U5104 ( .A1(n48269), .A2(n24135), .ZN(n49130) );
  NAND2_X1 U53405 ( .A1(n63605), .A2(n1642), .ZN(n48441) );
  NAND2_X1 U26719 ( .A1(n19634), .A2(n7868), .ZN(n50239) );
  NAND2_X1 U994 ( .A1(n50304), .A2(n1643), .ZN(n58290) );
  NAND2_X1 U819 ( .A1(n58856), .A2(n8790), .ZN(n49408) );
  NOR2_X1 U42434 ( .A1(n50093), .A2(n12580), .ZN(n47925) );
  NAND3_X1 U4476 ( .A1(n49694), .A2(n24049), .A3(n22157), .ZN(n49705) );
  NAND2_X1 U8555 ( .A1(n49276), .A2(n16862), .ZN(n48367) );
  BUF_X2 U23912 ( .I(n50309), .Z(n4699) );
  NOR2_X1 U987 ( .A1(n50420), .A2(n23063), .ZN(n49245) );
  CLKBUF_X2 U5626 ( .I(n24073), .Z(n58306) );
  NAND2_X1 U922 ( .A1(n18975), .A2(n49166), .ZN(n49560) );
  NOR2_X1 U836 ( .A1(n5282), .A2(n23707), .ZN(n49038) );
  NAND2_X1 U4064 ( .A1(n50060), .A2(n3055), .ZN(n49142) );
  NOR2_X1 U3598 ( .A1(n50333), .A2(n50340), .ZN(n49972) );
  NAND2_X1 U32102 ( .A1(n10422), .A2(n49529), .ZN(n49428) );
  NAND2_X1 U53956 ( .A1(n3055), .A2(n50309), .ZN(n14617) );
  NOR2_X1 U31989 ( .A1(n11794), .A2(n23912), .ZN(n49260) );
  NAND2_X1 U33962 ( .A1(n58983), .A2(n49538), .ZN(n48907) );
  NAND2_X1 U39319 ( .A1(n10422), .A2(n49538), .ZN(n48906) );
  NOR2_X1 U51801 ( .A1(n61513), .A2(n49395), .ZN(n49391) );
  NAND2_X1 U32992 ( .A1(n21226), .A2(n50346), .ZN(n50259) );
  NAND2_X1 U37173 ( .A1(n24069), .A2(n49908), .ZN(n49909) );
  NAND2_X1 U33503 ( .A1(n15709), .A2(n13038), .ZN(n13819) );
  CLKBUF_X2 U4949 ( .I(n19544), .Z(n149) );
  NOR2_X1 U722 ( .A1(n64135), .A2(n61742), .ZN(n48431) );
  NOR2_X1 U7295 ( .A1(n49606), .A2(n49315), .ZN(n49000) );
  NOR2_X1 U11599 ( .A1(n60428), .A2(n1383), .ZN(n49340) );
  INV_X1 U37109 ( .I(n24049), .ZN(n48893) );
  INV_X1 U15548 ( .I(n13549), .ZN(n49278) );
  INV_X1 U1015 ( .I(n49602), .ZN(n59084) );
  NAND2_X1 U9912 ( .A1(n1473), .A2(n3031), .ZN(n22926) );
  INV_X1 U39808 ( .I(n49376), .ZN(n49533) );
  INV_X1 U24809 ( .I(n20055), .ZN(n49846) );
  NAND2_X1 U839 ( .A1(n18882), .A2(n19634), .ZN(n8729) );
  BUF_X2 U34347 ( .I(n19681), .Z(n60510) );
  INV_X1 U50836 ( .I(n5713), .ZN(n6896) );
  NOR2_X1 U7271 ( .A1(n49908), .A2(n13839), .ZN(n48330) );
  NAND2_X1 U10832 ( .A1(n858), .A2(n49109), .ZN(n49111) );
  NAND2_X1 U671 ( .A1(n4734), .A2(n22717), .ZN(n50294) );
  INV_X1 U3914 ( .I(n49007), .ZN(n47054) );
  INV_X1 U15610 ( .I(n49025), .ZN(n50083) );
  INV_X1 U954 ( .I(n23141), .ZN(n4017) );
  NAND2_X1 U7285 ( .A1(n1205), .A2(n49459), .ZN(n10831) );
  NOR2_X1 U17625 ( .A1(n4526), .A2(n23738), .ZN(n44409) );
  INV_X1 U792 ( .I(n7113), .ZN(n48063) );
  INV_X1 U12437 ( .I(n20363), .ZN(n48863) );
  INV_X1 U26934 ( .I(n14315), .ZN(n19243) );
  NAND2_X1 U12452 ( .A1(n9177), .A2(n12701), .ZN(n49296) );
  NOR2_X1 U24001 ( .A1(n48768), .A2(n48366), .ZN(n49284) );
  NAND2_X1 U1021 ( .A1(n58443), .A2(n9177), .ZN(n16730) );
  NAND2_X1 U21571 ( .A1(n9177), .A2(n65245), .ZN(n49504) );
  NAND2_X1 U23244 ( .A1(n7868), .A2(n22264), .ZN(n17446) );
  NAND2_X1 U31302 ( .A1(n49166), .A2(n18918), .ZN(n48280) );
  NAND2_X1 U41858 ( .A1(n50044), .A2(n20199), .ZN(n49581) );
  NAND3_X1 U849 ( .A1(n14265), .A2(n49722), .A3(n49721), .ZN(n49724) );
  NOR2_X1 U15471 ( .A1(n49452), .A2(n6341), .ZN(n20013) );
  OAI21_X1 U54001 ( .A1(n21052), .A2(n13684), .B(n50340), .ZN(n49976) );
  NOR2_X1 U4787 ( .A1(n48454), .A2(n11641), .ZN(n11640) );
  NAND2_X1 U37180 ( .A1(n502), .A2(n61530), .ZN(n47334) );
  NOR2_X1 U39850 ( .A1(n47456), .A2(n63876), .ZN(n47457) );
  INV_X1 U53394 ( .I(n49430), .ZN(n47912) );
  NAND3_X1 U35526 ( .A1(n50288), .A2(n50287), .A3(n21092), .ZN(n17955) );
  AOI21_X1 U10806 ( .A1(n49282), .A2(n14005), .B(n1633), .ZN(n12214) );
  AOI22_X1 U5687 ( .A1(n47955), .A2(n48716), .B1(n49885), .B2(n18607), .ZN(
        n47958) );
  NAND2_X1 U6651 ( .A1(n50083), .A2(n50082), .ZN(n61541) );
  NOR2_X1 U27605 ( .A1(n48956), .A2(n47058), .ZN(n15366) );
  NAND3_X1 U7281 ( .A1(n2542), .A2(n49365), .A3(n1089), .ZN(n2541) );
  NAND2_X1 U15499 ( .A1(n1380), .A2(n49253), .ZN(n19832) );
  NOR2_X1 U36209 ( .A1(n21127), .A2(n24393), .ZN(n48281) );
  AOI21_X1 U699 ( .A1(n49142), .A2(n50058), .B(n4699), .ZN(n49149) );
  NOR2_X1 U13740 ( .A1(n3394), .A2(n61678), .ZN(n10855) );
  NOR2_X1 U51795 ( .A1(n49393), .A2(n4815), .ZN(n44003) );
  NOR2_X1 U4905 ( .A1(n18814), .A2(n49543), .ZN(n18813) );
  NAND2_X1 U26574 ( .A1(n46261), .A2(n21367), .ZN(n6898) );
  NOR2_X1 U10854 ( .A1(n64006), .A2(n49674), .ZN(n47647) );
  OAI21_X1 U22880 ( .A1(n49023), .A2(n50394), .B(n4174), .ZN(n24681) );
  NOR2_X1 U21243 ( .A1(n48757), .A2(n2878), .ZN(n50430) );
  NAND2_X1 U52509 ( .A1(n49243), .A2(n50427), .ZN(n45459) );
  INV_X1 U11415 ( .I(n44009), .ZN(n2321) );
  INV_X1 U12445 ( .I(n60520), .ZN(n48381) );
  NAND2_X1 U37117 ( .A1(n48380), .A2(n696), .ZN(n20664) );
  NOR3_X1 U8561 ( .A1(n12580), .A2(n61355), .A3(n50093), .ZN(n12624) );
  NOR2_X1 U35542 ( .A1(n59084), .A2(n25032), .ZN(n49312) );
  NOR2_X1 U43323 ( .A1(n62054), .A2(n49767), .ZN(n25048) );
  NOR2_X1 U22879 ( .A1(n50082), .A2(n4174), .ZN(n8992) );
  NAND3_X1 U29290 ( .A1(n7289), .A2(n9052), .A3(n7288), .ZN(n49709) );
  NAND2_X1 U29280 ( .A1(n18609), .A2(n60487), .ZN(n19775) );
  NAND2_X1 U33769 ( .A1(n25103), .A2(n49201), .ZN(n59586) );
  NOR2_X1 U874 ( .A1(n49547), .A2(n48280), .ZN(n49168) );
  NAND2_X1 U38725 ( .A1(n57397), .A2(n1224), .ZN(n50292) );
  NOR2_X1 U41439 ( .A1(n50095), .A2(n17818), .ZN(n50522) );
  NOR2_X1 U25354 ( .A1(n25018), .A2(n23156), .ZN(n5661) );
  NAND3_X1 U53537 ( .A1(n58306), .A2(n15737), .A3(n64), .ZN(n48355) );
  NOR2_X1 U28084 ( .A1(n1469), .A2(n16590), .ZN(n48423) );
  NOR2_X1 U37860 ( .A1(n49428), .A2(n49377), .ZN(n16408) );
  NOR2_X1 U696 ( .A1(n50353), .A2(n6977), .ZN(n49135) );
  NAND2_X1 U53781 ( .A1(n24394), .A2(n49170), .ZN(n49559) );
  NAND2_X1 U34363 ( .A1(n8129), .A2(n25032), .ZN(n49314) );
  INV_X1 U24172 ( .I(n46968), .ZN(n48799) );
  NAND2_X1 U37092 ( .A1(n63664), .A2(n14561), .ZN(n47990) );
  NOR2_X1 U5069 ( .A1(n23992), .A2(n63876), .ZN(n47458) );
  NAND2_X1 U53748 ( .A1(n49832), .A2(n49065), .ZN(n49066) );
  OAI21_X1 U11512 ( .A1(n49313), .A2(n49314), .B(n11172), .ZN(n9442) );
  OAI21_X1 U54369 ( .A1(n61759), .A2(n50117), .B(n18607), .ZN(n61218) );
  NAND3_X1 U35907 ( .A1(n10915), .A2(n14561), .A3(n18469), .ZN(n49710) );
  AOI21_X1 U6511 ( .A1(n4212), .A2(n49648), .B(n50312), .ZN(n49653) );
  NOR2_X1 U37955 ( .A1(n16571), .A2(n49541), .ZN(n18816) );
  NAND2_X1 U14612 ( .A1(n48355), .A2(n48889), .ZN(n48356) );
  NOR2_X1 U22387 ( .A1(n60428), .A2(n64751), .ZN(n47998) );
  NOR2_X1 U6554 ( .A1(n57193), .A2(n17955), .ZN(n60376) );
  AOI21_X1 U52367 ( .A1(n45175), .A2(n48354), .B(n45174), .ZN(n45176) );
  NOR2_X1 U11604 ( .A1(n11867), .A2(n48691), .ZN(n57666) );
  AOI21_X1 U10805 ( .A1(n49849), .A2(n49848), .B(n49847), .ZN(n49853) );
  INV_X1 U53666 ( .I(n48809), .ZN(n48813) );
  NAND2_X1 U10856 ( .A1(n49682), .A2(n49090), .ZN(n48707) );
  NOR2_X1 U6525 ( .A1(n2381), .A2(n58122), .ZN(n5209) );
  OAI21_X1 U53708 ( .A1(n25065), .A2(n48933), .B(n48932), .ZN(n48934) );
  NAND3_X1 U32056 ( .A1(n21351), .A2(n7527), .A3(n59369), .ZN(n4425) );
  NAND2_X1 U11776 ( .A1(n5426), .A2(n2629), .ZN(n18083) );
  NOR2_X1 U45296 ( .A1(n5805), .A2(n57366), .ZN(n8377) );
  NOR2_X1 U21945 ( .A1(n15990), .A2(n58198), .ZN(n14042) );
  NAND2_X1 U30693 ( .A1(n24394), .A2(n18975), .ZN(n49167) );
  NOR2_X1 U53715 ( .A1(n20055), .A2(n48970), .ZN(n49854) );
  NOR2_X1 U52126 ( .A1(n63923), .A2(n49910), .ZN(n48736) );
  INV_X1 U27603 ( .I(n11108), .ZN(n14254) );
  INV_X1 U730 ( .I(n4908), .ZN(n48683) );
  INV_X1 U9916 ( .I(n43757), .ZN(n49215) );
  AND2_X1 U12470 ( .A1(n15832), .A2(n63186), .Z(n19752) );
  OAI22_X1 U40358 ( .A1(n48855), .A2(n49301), .B1(n48698), .B2(n20363), .ZN(
        n48699) );
  AOI21_X1 U19958 ( .A1(n2956), .A2(n10637), .B(n49431), .ZN(n11003) );
  NAND4_X1 U7302 ( .A1(n46725), .A2(n50400), .A3(n63238), .A4(n49420), .ZN(
        n46726) );
  NAND2_X1 U10791 ( .A1(n49853), .A2(n49852), .ZN(n49855) );
  NOR3_X1 U31092 ( .A1(n16233), .A2(n50448), .A3(n19618), .ZN(n17926) );
  NOR2_X1 U43588 ( .A1(n1626), .A2(n10563), .ZN(n25501) );
  OAI21_X1 U848 ( .A1(n62593), .A2(n48769), .B(n48923), .ZN(n48773) );
  NAND3_X1 U15236 ( .A1(n48348), .A2(n48811), .A3(n48347), .ZN(n2073) );
  OAI21_X1 U31076 ( .A1(n61741), .A2(n48911), .B(n48910), .ZN(n48912) );
  NOR2_X1 U717 ( .A1(n13363), .A2(n1115), .ZN(n59965) );
  NAND4_X1 U51453 ( .A1(n61050), .A2(n50298), .A3(n8251), .A4(n50300), .ZN(
        n50316) );
  NAND3_X1 U707 ( .A1(n8502), .A2(n48677), .A3(n62192), .ZN(n59184) );
  NOR3_X1 U645 ( .A1(n50051), .A2(n50052), .A3(n16917), .ZN(n16916) );
  NAND3_X1 U662 ( .A1(n12675), .A2(n47060), .A3(n12674), .ZN(n9156) );
  NOR2_X1 U751 ( .A1(n57349), .A2(n60083), .ZN(n1920) );
  NOR2_X1 U15261 ( .A1(n48399), .A2(n8579), .ZN(n8578) );
  NOR2_X1 U9172 ( .A1(n5637), .A2(n5635), .ZN(n5657) );
  NOR3_X1 U680 ( .A1(n11867), .A2(n19294), .A3(n48071), .ZN(n50755) );
  NAND2_X1 U6574 ( .A1(n47348), .A2(n57346), .ZN(n45999) );
  AND2_X1 U623 ( .A1(n49920), .A2(n1629), .Z(n24336) );
  NOR3_X1 U10814 ( .A1(n15348), .A2(n49168), .A3(n49169), .ZN(n10315) );
  INV_X1 U15205 ( .I(n50752), .ZN(n50758) );
  INV_X1 U639 ( .I(n52445), .ZN(n25191) );
  NOR2_X1 U11608 ( .A1(n48772), .A2(n48773), .ZN(n3593) );
  NOR2_X1 U642 ( .A1(n50755), .A2(n46974), .ZN(n50751) );
  INV_X2 U24147 ( .I(n8075), .ZN(n8076) );
  INV_X1 U8019 ( .I(n50648), .ZN(n12942) );
  INV_X1 U28158 ( .I(n8076), .ZN(n8077) );
  NAND3_X1 U15176 ( .A1(n50758), .A2(n50757), .A3(n50756), .ZN(n50759) );
  CLKBUF_X2 U10780 ( .I(n18103), .Z(n2603) );
  INV_X2 U33032 ( .I(n24803), .ZN(n51788) );
  INV_X1 U610 ( .I(n24005), .ZN(n1464) );
  BUF_X2 U598 ( .I(n23571), .Z(n20302) );
  INV_X1 U5356 ( .I(n52107), .ZN(n5167) );
  INV_X1 U613 ( .I(n25394), .ZN(n51298) );
  BUF_X2 U15141 ( .I(n51691), .Z(n4470) );
  INV_X1 U7312 ( .I(n51986), .ZN(n24776) );
  BUF_X2 U577 ( .I(n51748), .Z(n23022) );
  BUF_X2 U38201 ( .I(n23792), .Z(n16984) );
  BUF_X2 U7877 ( .I(n52404), .Z(n24053) );
  BUF_X2 U41163 ( .I(n24079), .Z(n21425) );
  INV_X1 U589 ( .I(n14372), .ZN(n23758) );
  CLKBUF_X2 U657 ( .I(n52177), .Z(n23016) );
  INV_X1 U20334 ( .I(n7246), .ZN(n15873) );
  INV_X1 U567 ( .I(n5878), .ZN(n22577) );
  BUF_X4 U4458 ( .I(n50716), .Z(n52530) );
  INV_X1 U54432 ( .I(n52335), .ZN(n51048) );
  INV_X1 U36220 ( .I(n22845), .ZN(n25814) );
  INV_X1 U15107 ( .I(n20512), .ZN(n12283) );
  BUF_X2 U668 ( .I(n51081), .Z(n7459) );
  INV_X1 U5803 ( .I(n21100), .ZN(n23674) );
  INV_X1 U27714 ( .I(n8143), .ZN(n15719) );
  INV_X1 U7310 ( .I(n16593), .ZN(n19029) );
  INV_X1 U37310 ( .I(n7711), .ZN(n18260) );
  INV_X1 U11830 ( .I(n19224), .ZN(n11650) );
  INV_X1 U31235 ( .I(n10727), .ZN(n23197) );
  INV_X1 U11864 ( .I(n19810), .ZN(n52114) );
  INV_X1 U31781 ( .I(n11487), .ZN(n51807) );
  INV_X1 U15095 ( .I(n62574), .ZN(n11955) );
  INV_X1 U30680 ( .I(n17441), .ZN(n52585) );
  INV_X1 U56922 ( .I(n5349), .ZN(n61508) );
  INV_X1 U32564 ( .I(n23197), .ZN(n17940) );
  BUF_X2 U553 ( .I(n50151), .Z(n53917) );
  INV_X2 U28086 ( .I(n8023), .ZN(n55261) );
  BUF_X2 U12308 ( .I(n51333), .Z(n56544) );
  INV_X2 U641 ( .I(n8121), .ZN(n24944) );
  BUF_X2 U5536 ( .I(n53917), .Z(n60049) );
  INV_X2 U4352 ( .I(n53845), .ZN(n17057) );
  INV_X1 U10765 ( .I(n14977), .ZN(n14978) );
  CLKBUF_X2 U26818 ( .I(n25047), .Z(n13292) );
  BUF_X2 U15020 ( .I(n12605), .Z(n56567) );
  INV_X2 U7938 ( .I(n19556), .ZN(n20349) );
  BUF_X2 U14997 ( .I(n25213), .Z(n10441) );
  CLKBUF_X2 U4307 ( .I(n14977), .Z(n14307) );
  INV_X1 U19430 ( .I(n57901), .ZN(n22499) );
  INV_X2 U30751 ( .I(n23157), .ZN(n52837) );
  BUF_X2 U27064 ( .I(n12027), .Z(n1237) );
  INV_X1 U10759 ( .I(n24352), .ZN(n57039) );
  INV_X2 U42627 ( .I(n55286), .ZN(n55476) );
  INV_X1 U37831 ( .I(n17251), .ZN(n19555) );
  INV_X1 U40235 ( .I(n25252), .ZN(n56249) );
  INV_X1 U22372 ( .I(n52861), .ZN(n21669) );
  INV_X1 U9162 ( .I(n25803), .ZN(n1287) );
  INV_X1 U626 ( .I(n57073), .ZN(n59951) );
  INV_X2 U23344 ( .I(n26095), .ZN(n54951) );
  CLKBUF_X2 U10753 ( .I(n25168), .Z(n10183) );
  INV_X2 U41379 ( .I(n21919), .ZN(n54057) );
  INV_X1 U54480 ( .I(n20737), .ZN(n51162) );
  INV_X1 U27221 ( .I(n53381), .ZN(n50674) );
  CLKBUF_X2 U415 ( .I(n54072), .Z(n61371) );
  NAND2_X1 U25340 ( .A1(n16427), .A2(n60002), .ZN(n52996) );
  NOR2_X1 U19998 ( .A1(n55476), .A2(n55727), .ZN(n55279) );
  BUF_X2 U23398 ( .I(n9388), .Z(n58380) );
  INV_X1 U27214 ( .I(n55443), .ZN(n7973) );
  NOR2_X1 U504 ( .A1(n13921), .A2(n52270), .ZN(n56985) );
  NAND2_X1 U430 ( .A1(n54072), .A2(n53848), .ZN(n52986) );
  CLKBUF_X2 U24124 ( .I(n54939), .Z(n4783) );
  INV_X2 U42185 ( .I(n56627), .ZN(n56635) );
  NAND2_X1 U6921 ( .A1(n23164), .A2(n26041), .ZN(n52975) );
  BUF_X2 U55271 ( .I(n55286), .Z(n61282) );
  INV_X2 U56948 ( .I(n58218), .ZN(n53444) );
  CLKBUF_X2 U12302 ( .I(n53214), .Z(n4658) );
  INV_X1 U20860 ( .I(n25746), .ZN(n53576) );
  INV_X2 U5282 ( .I(n58283), .ZN(n55265) );
  NOR2_X1 U522 ( .A1(n53915), .A2(n23217), .ZN(n53407) );
  INV_X2 U4209 ( .I(n18109), .ZN(n18294) );
  INV_X1 U34464 ( .I(n15804), .ZN(n24404) );
  INV_X1 U41088 ( .I(n54492), .ZN(n21296) );
  INV_X1 U31248 ( .I(n10748), .ZN(n53001) );
  AND2_X1 U624 ( .A1(n54292), .A2(n13184), .Z(n51779) );
  OR2_X1 U7478 ( .A1(n3673), .A2(n54323), .Z(n818) );
  INV_X1 U23605 ( .I(n2199), .ZN(n54949) );
  INV_X1 U31839 ( .I(n19567), .ZN(n23857) );
  INV_X1 U33173 ( .I(n25047), .ZN(n25067) );
  INV_X1 U4219 ( .I(n57048), .ZN(n17003) );
  INV_X1 U4893 ( .I(n18247), .ZN(n54858) );
  INV_X1 U417 ( .I(n24455), .ZN(n14142) );
  BUF_X2 U10752 ( .I(n53232), .Z(n20156) );
  INV_X1 U15018 ( .I(n52866), .ZN(n57004) );
  INV_X2 U490 ( .I(n22029), .ZN(n56381) );
  INV_X1 U34858 ( .I(n54323), .ZN(n54074) );
  INV_X8 U30303 ( .I(n24259), .ZN(n12468) );
  INV_X2 U11951 ( .I(n56417), .ZN(n56217) );
  NOR2_X1 U471 ( .A1(n6531), .A2(n55469), .ZN(n55726) );
  NOR2_X1 U55649 ( .A1(n54065), .A2(n7532), .ZN(n54066) );
  NOR2_X1 U34342 ( .A1(n56403), .A2(n14978), .ZN(n55952) );
  INV_X2 U54066 ( .I(n54035), .ZN(n54052) );
  NAND2_X1 U6474 ( .A1(n7973), .A2(n23275), .ZN(n52492) );
  NAND2_X1 U33273 ( .A1(n52819), .A2(n53444), .ZN(n52815) );
  INV_X1 U14890 ( .I(n18750), .ZN(n52125) );
  NOR2_X1 U56579 ( .A1(n56545), .A2(n57013), .ZN(n56529) );
  NAND2_X1 U56756 ( .A1(n57068), .A2(n21079), .ZN(n57069) );
  NAND2_X1 U54362 ( .A1(n64808), .A2(n56436), .ZN(n50882) );
  NOR2_X1 U9141 ( .A1(n51162), .A2(n56404), .ZN(n56595) );
  INV_X1 U483 ( .I(n1325), .ZN(n20921) );
  NAND2_X1 U33759 ( .A1(n23873), .A2(n56659), .ZN(n56239) );
  INV_X1 U31837 ( .I(n11571), .ZN(n53397) );
  NOR2_X1 U15723 ( .A1(n14226), .A2(n5907), .ZN(n52487) );
  BUF_X4 U42535 ( .I(n51632), .Z(n54659) );
  NAND2_X1 U21774 ( .A1(n24669), .A2(n56381), .ZN(n137) );
  INV_X1 U8522 ( .I(n56370), .ZN(n52282) );
  NAND3_X1 U55115 ( .A1(n14457), .A2(n54860), .A3(n54640), .ZN(n54460) );
  NOR2_X1 U40687 ( .A1(n22775), .A2(n54067), .ZN(n53835) );
  NOR2_X1 U37288 ( .A1(n53848), .A2(n54072), .ZN(n54502) );
  NOR2_X1 U55018 ( .A1(n52958), .A2(n54938), .ZN(n54431) );
  NAND2_X1 U28530 ( .A1(n52825), .A2(n7095), .ZN(n53435) );
  BUF_X2 U5283 ( .I(n54314), .Z(n60794) );
  NAND3_X1 U31480 ( .A1(n24749), .A2(n55486), .A3(n10362), .ZN(n18548) );
  NOR2_X1 U29591 ( .A1(n58218), .A2(n12574), .ZN(n53437) );
  NAND2_X1 U447 ( .A1(n1616), .A2(n64808), .ZN(n56430) );
  INV_X1 U420 ( .I(n13920), .ZN(n52687) );
  INV_X2 U439 ( .I(n22114), .ZN(n23110) );
  NOR2_X1 U33307 ( .A1(n23701), .A2(n53226), .ZN(n53586) );
  INV_X2 U7470 ( .I(n61443), .ZN(n54598) );
  INV_X1 U8514 ( .I(n57013), .ZN(n16644) );
  INV_X1 U521 ( .I(n55908), .ZN(n52124) );
  NOR2_X1 U3926 ( .A1(n56268), .A2(n61321), .ZN(n55922) );
  INV_X1 U25474 ( .I(n22544), .ZN(n5777) );
  INV_X1 U437 ( .I(n56397), .ZN(n56563) );
  INV_X1 U5496 ( .I(n56250), .ZN(n57203) );
  BUF_X2 U440 ( .I(n52044), .Z(n55695) );
  INV_X2 U487 ( .I(n61168), .ZN(n1146) );
  INV_X1 U477 ( .I(n15040), .ZN(n14358) );
  INV_X1 U21203 ( .I(n11938), .ZN(n15929) );
  NAND2_X1 U25392 ( .A1(n54057), .A2(n53907), .ZN(n54045) );
  INV_X1 U40259 ( .I(n60225), .ZN(n57031) );
  INV_X1 U32706 ( .I(n53535), .ZN(n53540) );
  INV_X2 U29002 ( .I(n15706), .ZN(n9003) );
  INV_X1 U479 ( .I(n59020), .ZN(n1612) );
  INV_X1 U37492 ( .I(n25167), .ZN(n56573) );
  INV_X1 U496 ( .I(n2959), .ZN(n13815) );
  INV_X1 U55401 ( .I(n53379), .ZN(n53602) );
  INV_X2 U19399 ( .I(n25127), .ZN(n54340) );
  INV_X1 U9845 ( .I(n53539), .ZN(n1455) );
  INV_X1 U5392 ( .I(n57051), .ZN(n53440) );
  AND2_X1 U38677 ( .A1(n25936), .A2(n53213), .Z(n57025) );
  NAND2_X1 U28020 ( .A1(n54652), .A2(n62768), .ZN(n54653) );
  CLKBUF_X2 U4865 ( .I(n54815), .Z(n60751) );
  NAND2_X1 U33886 ( .A1(n53848), .A2(n54314), .ZN(n54063) );
  INV_X1 U8525 ( .I(n53622), .ZN(n1259) );
  INV_X1 U23673 ( .I(n18597), .ZN(n24553) );
  OAI21_X1 U55643 ( .A1(n54047), .A2(n54046), .B(n54054), .ZN(n54050) );
  NAND3_X1 U37287 ( .A1(n56372), .A2(n56371), .A3(n23526), .ZN(n56373) );
  NAND3_X1 U8397 ( .A1(n55024), .A2(n7800), .A3(n20740), .ZN(n54453) );
  NAND3_X1 U27223 ( .A1(n53381), .A2(n52837), .A3(n52756), .ZN(n53608) );
  NOR2_X1 U37278 ( .A1(n53427), .A2(n53860), .ZN(n18520) );
  NAND2_X1 U8505 ( .A1(n53614), .A2(n53613), .ZN(n53853) );
  NAND2_X1 U32657 ( .A1(n12574), .A2(n17003), .ZN(n50803) );
  NAND3_X1 U4336 ( .A1(n56206), .A2(n56205), .A3(n56619), .ZN(n51113) );
  NAND2_X1 U32575 ( .A1(n56554), .A2(n24696), .ZN(n21844) );
  INV_X1 U14845 ( .I(n54341), .ZN(n54342) );
  NAND2_X1 U14950 ( .A1(n64850), .A2(n64808), .ZN(n56228) );
  NOR2_X1 U6537 ( .A1(n56408), .A2(n57691), .ZN(n56257) );
  INV_X1 U10693 ( .I(n52048), .ZN(n9912) );
  NAND3_X1 U3963 ( .A1(n23563), .A2(n58225), .A3(n52819), .ZN(n20765) );
  INV_X1 U7323 ( .I(n56993), .ZN(n52883) );
  NAND2_X1 U424 ( .A1(n57700), .A2(n57699), .ZN(n54044) );
  NOR2_X1 U401 ( .A1(n56214), .A2(n23165), .ZN(n56636) );
  OAI21_X1 U55986 ( .A1(n55310), .A2(n55000), .B(n54999), .ZN(n55004) );
  NAND3_X1 U27220 ( .A1(n52845), .A2(n52844), .A3(n53381), .ZN(n53609) );
  NOR2_X1 U53899 ( .A1(n52768), .A2(n60002), .ZN(n53223) );
  NAND2_X1 U25472 ( .A1(n5777), .A2(n1139), .ZN(n13329) );
  NAND2_X1 U40628 ( .A1(n23736), .A2(n54594), .ZN(n53894) );
  NAND2_X1 U360 ( .A1(n58283), .A2(n19167), .ZN(n54843) );
  NOR2_X1 U366 ( .A1(n54597), .A2(n53890), .ZN(n54590) );
  NOR2_X1 U21660 ( .A1(n57073), .A2(n52861), .ZN(n52854) );
  NAND3_X1 U56870 ( .A1(n1601), .A2(n15304), .A3(n52235), .ZN(n12729) );
  NAND2_X1 U8513 ( .A1(n53006), .A2(n5008), .ZN(n53578) );
  INV_X2 U40961 ( .I(n57068), .ZN(n52863) );
  INV_X1 U29009 ( .I(n52890), .ZN(n56605) );
  NAND2_X1 U20091 ( .A1(n53445), .A2(n52815), .ZN(n9253) );
  NAND2_X1 U43817 ( .A1(n53587), .A2(n23476), .ZN(n52767) );
  INV_X1 U14806 ( .I(n57025), .ZN(n57023) );
  INV_X1 U5792 ( .I(n52477), .ZN(n5279) );
  INV_X1 U394 ( .I(n25080), .ZN(n24510) );
  INV_X1 U21368 ( .I(n1158), .ZN(n53548) );
  NOR2_X1 U42004 ( .A1(n55982), .A2(n1616), .ZN(n22804) );
  NAND2_X1 U12208 ( .A1(n54589), .A2(n54596), .ZN(n15249) );
  INV_X1 U347 ( .I(n16948), .ZN(n54990) );
  INV_X1 U43832 ( .I(n56436), .ZN(n56434) );
  NAND2_X1 U21296 ( .A1(n61405), .A2(n61528), .ZN(n56601) );
  NAND2_X1 U376 ( .A1(n54431), .A2(n1139), .ZN(n54956) );
  AOI21_X1 U341 ( .A1(n16801), .A2(n53220), .B(n57024), .ZN(n25109) );
  NAND3_X1 U56139 ( .A1(n55463), .A2(n58490), .A3(n55476), .ZN(n55733) );
  OAI21_X1 U35615 ( .A1(n24510), .A2(n1610), .B(n60794), .ZN(n26154) );
  AOI21_X1 U6746 ( .A1(n54024), .A2(n54023), .B(n15945), .ZN(n21931) );
  NOR2_X1 U6458 ( .A1(n52846), .A2(n53386), .ZN(n52842) );
  NOR3_X1 U30550 ( .A1(n53409), .A2(n53551), .A3(n53408), .ZN(n53413) );
  NAND2_X1 U26821 ( .A1(n15935), .A2(n50205), .ZN(n17265) );
  NAND2_X1 U25541 ( .A1(n23873), .A2(n56359), .ZN(n13575) );
  NAND2_X1 U56528 ( .A1(n56420), .A2(n56417), .ZN(n56418) );
  AOI22_X1 U8184 ( .A1(n54611), .A2(n54434), .B1(n54955), .B2(n4783), .ZN(
        n8163) );
  NOR2_X1 U31767 ( .A1(n59052), .A2(n1607), .ZN(n13794) );
  NOR2_X1 U326 ( .A1(n58175), .A2(n56532), .ZN(n1153) );
  OAI21_X1 U333 ( .A1(n54016), .A2(n53038), .B(n53037), .ZN(n53039) );
  NOR2_X1 U42037 ( .A1(n53572), .A2(n23476), .ZN(n53575) );
  NAND2_X1 U4974 ( .A1(n53837), .A2(n54307), .ZN(n57742) );
  INV_X1 U4620 ( .I(n3077), .ZN(n54592) );
  OAI22_X1 U6223 ( .A1(n54655), .A2(n14501), .B1(n54654), .B2(n5711), .ZN(
        n54697) );
  NAND4_X1 U55150 ( .A1(n52720), .A2(n56632), .A3(n1286), .A4(n56627), .ZN(
        n56220) );
  NAND3_X1 U14943 ( .A1(n56415), .A2(n56632), .A3(n61914), .ZN(n56421) );
  OAI21_X1 U54965 ( .A1(n63743), .A2(n52253), .B(n52672), .ZN(n52659) );
  NAND2_X1 U400 ( .A1(n52264), .A2(n64657), .ZN(n20488) );
  NOR2_X1 U351 ( .A1(n53238), .A2(n1602), .ZN(n57007) );
  NAND2_X1 U365 ( .A1(n14943), .A2(n56547), .ZN(n52708) );
  NAND2_X1 U40731 ( .A1(n56991), .A2(n61528), .ZN(n52893) );
  INV_X1 U312 ( .I(n52222), .ZN(n56271) );
  INV_X1 U14661 ( .I(n57056), .ZN(n53446) );
  NAND3_X1 U306 ( .A1(n55666), .A2(n55665), .A3(n56271), .ZN(n56275) );
  AOI21_X1 U12219 ( .A1(n20488), .A2(n57008), .B(n57004), .ZN(n20487) );
  NAND3_X1 U54704 ( .A1(n54824), .A2(n60751), .A3(n5711), .ZN(n51637) );
  OAI21_X1 U14870 ( .A1(n22210), .A2(n1368), .B(n54588), .ZN(n53891) );
  NAND2_X1 U9829 ( .A1(n51257), .A2(n56432), .ZN(n22620) );
  AOI21_X1 U40171 ( .A1(n56419), .A2(n56420), .B(n56421), .ZN(n20003) );
  NAND2_X1 U26835 ( .A1(n53878), .A2(n13661), .ZN(n13660) );
  INV_X1 U43926 ( .I(n56630), .ZN(n56209) );
  NAND3_X1 U54644 ( .A1(n52860), .A2(n59952), .A3(n51465), .ZN(n51468) );
  AOI21_X1 U44450 ( .A1(n54638), .A2(n54639), .B(n57287), .ZN(n1171) );
  NAND3_X1 U6169 ( .A1(n56236), .A2(n56235), .A3(n56243), .ZN(n18023) );
  NOR2_X1 U296 ( .A1(n25109), .A2(n58151), .ZN(n12134) );
  NOR2_X1 U293 ( .A1(n52841), .A2(n60909), .ZN(n19083) );
  NAND2_X1 U279 ( .A1(n13328), .A2(n13329), .ZN(n54435) );
  NAND2_X1 U4022 ( .A1(n61463), .A2(n59052), .ZN(n54819) );
  NAND3_X1 U42336 ( .A1(n61920), .A2(n61516), .A3(n52863), .ZN(n51469) );
  OAI21_X1 U55932 ( .A1(n60751), .A2(n54814), .B(n62768), .ZN(n54816) );
  AOI21_X1 U34401 ( .A1(n17258), .A2(n15059), .B(n17257), .ZN(n17256) );
  NAND2_X1 U26423 ( .A1(n53040), .A2(n10527), .ZN(n6742) );
  NOR2_X1 U10698 ( .A1(n54435), .A2(n64989), .ZN(n7475) );
  OAI21_X1 U30598 ( .A1(n53910), .A2(n1141), .B(n10245), .ZN(n53923) );
  OAI21_X1 U26216 ( .A1(n58768), .A2(n58767), .B(n51435), .ZN(n51448) );
  NAND2_X1 U25819 ( .A1(n10214), .A2(n52766), .ZN(n52804) );
  BUF_X2 U14581 ( .I(n53632), .Z(n53699) );
  BUF_X4 U26842 ( .I(n59445), .Z(n59180) );
  NAND2_X1 U54887 ( .A1(n52040), .A2(n52039), .ZN(n55868) );
  INV_X2 U8482 ( .I(n7020), .ZN(n9595) );
  NAND2_X1 U247 ( .A1(n55156), .A2(n55157), .ZN(n52645) );
  INV_X2 U28004 ( .I(n23603), .ZN(n25299) );
  INV_X1 U48928 ( .I(n13939), .ZN(n6061) );
  BUF_X4 U42023 ( .I(n55015), .Z(n55089) );
  BUF_X2 U4541 ( .I(n55151), .Z(n10310) );
  INV_X2 U26704 ( .I(n9595), .ZN(n7021) );
  NAND2_X1 U43449 ( .A1(n14643), .A2(n54197), .ZN(n54188) );
  CLKBUF_X2 U231 ( .I(n55892), .Z(n13858) );
  INV_X2 U12926 ( .I(n20625), .ZN(n21569) );
  BUF_X2 U14586 ( .I(n54507), .Z(n54565) );
  INV_X1 U7969 ( .I(n53163), .ZN(n25484) );
  NAND2_X1 U29053 ( .A1(n1591), .A2(n59180), .ZN(n11144) );
  INV_X1 U57219 ( .I(n55892), .ZN(n55854) );
  INV_X2 U230 ( .I(n53672), .ZN(n53690) );
  INV_X1 U4380 ( .I(n52878), .ZN(n53094) );
  INV_X2 U37870 ( .I(n53740), .ZN(n53726) );
  INV_X1 U4692 ( .I(n55582), .ZN(n21273) );
  INV_X1 U126 ( .I(n53688), .ZN(n53691) );
  INV_X2 U34246 ( .I(n56084), .ZN(n56104) );
  INV_X2 U43292 ( .I(n63013), .ZN(n56108) );
  NAND2_X1 U29408 ( .A1(n16943), .A2(n17155), .ZN(n55175) );
  INV_X1 U14606 ( .I(n55151), .ZN(n55165) );
  INV_X2 U195 ( .I(n17795), .ZN(n1366) );
  INV_X4 U180 ( .I(n55089), .ZN(n55068) );
  INV_X1 U25747 ( .I(n54362), .ZN(n54393) );
  NOR2_X1 U21738 ( .A1(n23554), .A2(n24063), .ZN(n55350) );
  NAND2_X1 U56994 ( .A1(n56092), .A2(n63013), .ZN(n56080) );
  INV_X2 U7954 ( .I(n23212), .ZN(n4033) );
  NOR2_X1 U18953 ( .A1(n53355), .A2(n52808), .ZN(n53312) );
  INV_X1 U9110 ( .I(n12111), .ZN(n7182) );
  NAND2_X1 U31410 ( .A1(n3307), .A2(n58463), .ZN(n8222) );
  NOR2_X1 U5930 ( .A1(n6168), .A2(n6134), .ZN(n25344) );
  BUF_X2 U201 ( .I(n13939), .Z(n12915) );
  NAND2_X1 U54956 ( .A1(n55628), .A2(n19021), .ZN(n52301) );
  NAND2_X1 U188 ( .A1(n4030), .A2(n25147), .ZN(n57144) );
  NAND2_X1 U7376 ( .A1(n22401), .A2(n1367), .ZN(n54379) );
  NAND2_X1 U9810 ( .A1(n11716), .A2(n19161), .ZN(n8985) );
  INV_X4 U36352 ( .I(n54196), .ZN(n54192) );
  BUF_X2 U23326 ( .I(n54409), .Z(n271) );
  NOR2_X1 U39910 ( .A1(n53672), .A2(n53695), .ZN(n53694) );
  NOR2_X1 U38950 ( .A1(n15703), .A2(n14428), .ZN(n55384) );
  INV_X2 U14572 ( .I(n17155), .ZN(n1587) );
  NOR2_X1 U4128 ( .A1(n22516), .A2(n57124), .ZN(n57136) );
  INV_X2 U27639 ( .I(n23030), .ZN(n56806) );
  INV_X1 U6567 ( .I(n9102), .ZN(n55056) );
  INV_X1 U43466 ( .I(n54669), .ZN(n54723) );
  NOR2_X1 U3819 ( .A1(n12111), .A2(n15415), .ZN(n15858) );
  NAND2_X1 U42052 ( .A1(n55828), .A2(n24958), .ZN(n55796) );
  INV_X1 U38709 ( .I(n55224), .ZN(n60037) );
  INV_X2 U141 ( .I(n1232), .ZN(n53303) );
  NAND2_X1 U12256 ( .A1(n56502), .A2(n21860), .ZN(n56499) );
  OR2_X1 U8114 ( .A1(n53014), .A2(n19085), .Z(n53813) );
  NAND2_X1 U3911 ( .A1(n18859), .A2(n2984), .ZN(n54204) );
  NOR2_X1 U3654 ( .A1(n53692), .A2(n53676), .ZN(n53673) );
  INV_X1 U139 ( .I(n11556), .ZN(n54390) );
  OR2_X1 U6146 ( .A1(n18582), .A2(n56935), .Z(n9035) );
  CLKBUF_X1 U187 ( .I(n17795), .Z(n59444) );
  CLKBUF_X2 U14599 ( .I(n56757), .Z(n7209) );
  NAND2_X1 U22705 ( .A1(n57015), .A2(n4030), .ZN(n57123) );
  INV_X1 U159 ( .I(n12923), .ZN(n16778) );
  NAND2_X1 U23648 ( .A1(n56106), .A2(n56104), .ZN(n56099) );
  NAND2_X1 U220 ( .A1(n53265), .A2(n1232), .ZN(n53305) );
  NOR2_X1 U39442 ( .A1(n55627), .A2(n19021), .ZN(n55650) );
  NAND2_X1 U55832 ( .A1(n18422), .A2(n22572), .ZN(n54567) );
  NAND2_X1 U4086 ( .A1(n23879), .A2(n56808), .ZN(n58687) );
  NAND2_X1 U4459 ( .A1(n17012), .A2(n53351), .ZN(n53366) );
  INV_X1 U56262 ( .I(n24958), .ZN(n55752) );
  INV_X1 U29548 ( .I(n56047), .ZN(n9568) );
  BUF_X8 U42413 ( .I(n56144), .Z(n56191) );
  NAND2_X1 U36323 ( .A1(n54582), .A2(n54561), .ZN(n54508) );
  INV_X1 U36312 ( .I(n53097), .ZN(n53100) );
  NOR2_X1 U56913 ( .A1(n56080), .A2(n56081), .ZN(n56102) );
  NAND2_X1 U9805 ( .A1(n56502), .A2(n59444), .ZN(n56517) );
  NAND2_X1 U14421 ( .A1(n22667), .A2(n23074), .ZN(n2371) );
  NOR2_X1 U37372 ( .A1(n56906), .A2(n14708), .ZN(n56970) );
  NOR2_X1 U28497 ( .A1(n9067), .A2(n25220), .ZN(n8411) );
  INV_X2 U23928 ( .I(n5553), .ZN(n55651) );
  NAND2_X1 U56545 ( .A1(n61964), .A2(n17795), .ZN(n56455) );
  NAND2_X1 U12180 ( .A1(n518), .A2(n62199), .ZN(n53269) );
  NAND2_X1 U96 ( .A1(n61760), .A2(n57156), .ZN(n3937) );
  AOI21_X1 U8467 ( .A1(n54192), .A2(n2984), .B(n18859), .ZN(n13716) );
  NAND2_X1 U38747 ( .A1(n55893), .A2(n22681), .ZN(n19034) );
  NAND2_X1 U56681 ( .A1(n65064), .A2(n23879), .ZN(n56776) );
  INV_X1 U7357 ( .I(n61687), .ZN(n1254) );
  NAND2_X1 U42763 ( .A1(n56837), .A2(n56885), .ZN(n56872) );
  NAND2_X1 U56742 ( .A1(n14708), .A2(n25022), .ZN(n56966) );
  NAND2_X1 U81 ( .A1(n56104), .A2(n56107), .ZN(n56009) );
  INV_X1 U14498 ( .I(n17500), .ZN(n14549) );
  NAND2_X1 U105 ( .A1(n5195), .A2(n56196), .ZN(n56177) );
  NAND2_X1 U7358 ( .A1(n14643), .A2(n54196), .ZN(n54201) );
  NOR2_X1 U56781 ( .A1(n21570), .A2(n57125), .ZN(n57157) );
  NAND2_X1 U25344 ( .A1(n56881), .A2(n5658), .ZN(n56856) );
  NAND2_X1 U56374 ( .A1(n56108), .A2(n9567), .ZN(n56018) );
  NAND2_X1 U53526 ( .A1(n53325), .A2(n53324), .ZN(n53361) );
  NOR3_X1 U30117 ( .A1(n23212), .A2(n23243), .A3(n53108), .ZN(n53066) );
  NAND2_X1 U5075 ( .A1(n5122), .A2(n55846), .ZN(n55897) );
  NOR2_X1 U4093 ( .A1(n56791), .A2(n23879), .ZN(n56778) );
  NAND2_X1 U28441 ( .A1(n10310), .A2(n55170), .ZN(n55147) );
  NAND2_X1 U4077 ( .A1(n54741), .A2(n22122), .ZN(n54718) );
  NOR2_X1 U94 ( .A1(n57156), .A2(n21829), .ZN(n57148) );
  NAND2_X1 U60 ( .A1(n55590), .A2(n55597), .ZN(n55584) );
  NAND2_X1 U30076 ( .A1(n1593), .A2(n11353), .ZN(n55119) );
  BUF_X2 U92 ( .I(n15237), .Z(n15238) );
  NOR2_X1 U87 ( .A1(n55089), .A2(n9067), .ZN(n11548) );
  BUF_X2 U9797 ( .I(n63039), .Z(n24032) );
  INV_X1 U42888 ( .I(n55625), .ZN(n52300) );
  INV_X1 U85 ( .I(n56952), .ZN(n56940) );
  INV_X1 U161 ( .I(n55339), .ZN(n55342) );
  NAND2_X1 U27156 ( .A1(n51878), .A2(n63873), .ZN(n54243) );
  NAND2_X1 U83 ( .A1(n55829), .A2(n55760), .ZN(n55816) );
  NAND2_X1 U42143 ( .A1(n23302), .A2(n4030), .ZN(n57116) );
  NOR2_X1 U56553 ( .A1(n20587), .A2(n21859), .ZN(n56473) );
  AND2_X1 U42438 ( .A1(n56886), .A2(n56894), .Z(n56861) );
  OR2_X1 U7970 ( .A1(n53166), .A2(n53130), .Z(n1177) );
  INV_X1 U57 ( .I(n54898), .ZN(n54914) );
  NAND2_X1 U72 ( .A1(n15703), .A2(n14428), .ZN(n55381) );
  AND2_X1 U4780 ( .A1(n22486), .A2(n2329), .Z(n17959) );
  INV_X1 U20981 ( .I(n54392), .ZN(n2676) );
  NAND2_X1 U35236 ( .A1(n22667), .A2(n56892), .ZN(n56893) );
  NAND2_X1 U28098 ( .A1(n1593), .A2(n7890), .ZN(n55140) );
  NAND2_X1 U4208 ( .A1(n26008), .A2(n54198), .ZN(n54162) );
  NOR2_X1 U32894 ( .A1(n17893), .A2(n56510), .ZN(n56496) );
  AOI21_X1 U55382 ( .A1(n53320), .A2(n9731), .B(n53351), .ZN(n53314) );
  NAND2_X1 U12349 ( .A1(n19845), .A2(n55654), .ZN(n58468) );
  AOI22_X1 U14913 ( .A1(n53293), .A2(n53303), .B1(n53294), .B2(n53302), .ZN(
        n14267) );
  NAND3_X1 U8425 ( .A1(n56815), .A2(n56791), .A3(n65064), .ZN(n56759) );
  NAND2_X1 U10653 ( .A1(n2619), .A2(n53690), .ZN(n53647) );
  NAND3_X1 U55699 ( .A1(n10480), .A2(n26008), .A3(n25299), .ZN(n54148) );
  NAND2_X1 U55543 ( .A1(n53812), .A2(n53794), .ZN(n53778) );
  INV_X1 U32435 ( .I(n56902), .ZN(n12397) );
  NOR2_X1 U4045 ( .A1(n55197), .A2(n17155), .ZN(n55204) );
  NAND3_X1 U5436 ( .A1(n55864), .A2(n55895), .A3(n60092), .ZN(n55850) );
  INV_X1 U4026 ( .I(n52231), .ZN(n53143) );
  INV_X1 U55687 ( .I(n54144), .ZN(n54134) );
  NAND2_X1 U27565 ( .A1(n52797), .A2(n52798), .ZN(n9937) );
  OAI21_X1 U4205 ( .A1(n24146), .A2(n58813), .B(n55219), .ZN(n55230) );
  NAND2_X1 U26747 ( .A1(n53795), .A2(n53794), .ZN(n53821) );
  AOI21_X1 U39104 ( .A1(n25764), .A2(n25763), .B(n18424), .ZN(n25762) );
  NAND4_X1 U25200 ( .A1(n53371), .A2(n53372), .A3(n53373), .A4(n53370), .ZN(
        n19838) );
  NAND2_X1 U62 ( .A1(n53249), .A2(n53248), .ZN(n60180) );
  NOR2_X1 U56045 ( .A1(n55218), .A2(n63193), .ZN(n55234) );
  NOR2_X1 U22131 ( .A1(n7181), .A2(n53160), .ZN(n52230) );
  INV_X1 U30 ( .I(n56157), .ZN(n56188) );
  NOR3_X1 U38798 ( .A1(n17893), .A2(n19827), .A3(n56456), .ZN(n56460) );
  OAI21_X1 U56671 ( .A1(n56813), .A2(n56775), .B(n65064), .ZN(n56763) );
  NAND4_X1 U27181 ( .A1(n53744), .A2(n53763), .A3(n53742), .A4(n53743), .ZN(
        n53745) );
  AOI21_X1 U4211 ( .A1(n57133), .A2(n57115), .B(n57110), .ZN(n57111) );
  AOI21_X1 U20405 ( .A1(n57998), .A2(n57997), .B(n57996), .ZN(n54869) );
  NAND4_X1 U36322 ( .A1(n22021), .A2(n53721), .A3(n53707), .A4(n53708), .ZN(
        n19110) );
  NOR2_X1 U6292 ( .A1(n58468), .A2(n55647), .ZN(n16574) );
  NOR2_X1 U27566 ( .A1(n9937), .A2(n22581), .ZN(n52813) );
  NAND4_X1 U9 ( .A1(n54885), .A2(n54887), .A3(n54886), .A4(n54884), .ZN(n60212) );
  NAND2_X1 U10 ( .A1(n5895), .A2(n51567), .ZN(n5894) );
  NAND2_X1 U11 ( .A1(n62913), .A2(n55030), .ZN(n8406) );
  OAI21_X1 U12 ( .A1(n10318), .A2(n13710), .B(n18859), .ZN(n13709) );
  OAI22_X1 U17 ( .A1(n18290), .A2(n23129), .B1(n15864), .B2(n61293), .ZN(n63)
         );
  AOI22_X1 U21 ( .A1(n62288), .A2(n8259), .B1(n52307), .B2(n55651), .ZN(n52315) );
  NAND2_X1 U31 ( .A1(n62756), .A2(n64646), .ZN(n51567) );
  INV_X1 U35 ( .I(n54214), .ZN(n64780) );
  NAND4_X1 U36 ( .A1(n53741), .A2(n7240), .A3(n25011), .A4(n16489), .ZN(n53742) );
  OAI21_X1 U38 ( .A1(n56071), .A2(n56117), .B(n13960), .ZN(n55997) );
  OR2_X1 U40 ( .A1(n58896), .A2(n54542), .Z(n54575) );
  AND2_X1 U46 ( .A1(n23785), .A2(n56697), .Z(n61766) );
  INV_X1 U51 ( .I(n54709), .ZN(n54755) );
  NOR2_X1 U53 ( .A1(n3525), .A2(n53147), .ZN(n53135) );
  INV_X1 U56 ( .I(n65007), .ZN(n15969) );
  NOR2_X1 U59 ( .A1(n23682), .A2(n56895), .ZN(n56870) );
  NAND2_X1 U63 ( .A1(n25115), .A2(n25011), .ZN(n53759) );
  NOR2_X1 U64 ( .A1(n7138), .A2(n54403), .ZN(n54366) );
  BUF_X2 U67 ( .I(n54196), .Z(n10480) );
  OAI21_X1 U69 ( .A1(n19475), .A2(n53672), .B(n53688), .ZN(n20615) );
  NAND2_X1 U73 ( .A1(n53800), .A2(n13503), .ZN(n13492) );
  NAND2_X1 U74 ( .A1(n53731), .A2(n53732), .ZN(n53720) );
  NAND2_X1 U77 ( .A1(n12915), .A2(n6135), .ZN(n58817) );
  AOI21_X1 U79 ( .A1(n56808), .A2(n56796), .B(n56791), .ZN(n62596) );
  NAND2_X1 U80 ( .A1(n56775), .A2(n56808), .ZN(n51473) );
  NOR2_X1 U88 ( .A1(n58687), .A2(n56749), .ZN(n64646) );
  OR2_X1 U95 ( .A1(n56196), .A2(n11716), .Z(n61873) );
  AOI21_X1 U98 ( .A1(n53265), .A2(n23956), .B(n9338), .ZN(n25545) );
  NAND2_X1 U101 ( .A1(n54424), .A2(n7138), .ZN(n54410) );
  AOI21_X1 U106 ( .A1(n53354), .A2(n9731), .B(n53369), .ZN(n52796) );
  AOI21_X1 U107 ( .A1(n54170), .A2(n26008), .B(n54189), .ZN(n57568) );
  INV_X1 U109 ( .I(n56103), .ZN(n56013) );
  INV_X1 U114 ( .I(n55641), .ZN(n55611) );
  NOR2_X1 U115 ( .A1(n56892), .A2(n21879), .ZN(n56837) );
  NAND2_X1 U118 ( .A1(n54403), .A2(n20985), .ZN(n54363) );
  NOR2_X1 U120 ( .A1(n63931), .A2(n17012), .ZN(n53325) );
  INV_X1 U121 ( .I(n53755), .ZN(n53731) );
  AND2_X1 U122 ( .A1(n21569), .A2(n23538), .Z(n61760) );
  NAND2_X1 U131 ( .A1(n9655), .A2(n14708), .ZN(n8722) );
  INV_X1 U132 ( .I(n25859), .ZN(n53675) );
  INV_X1 U136 ( .I(n26135), .ZN(n9533) );
  NOR2_X1 U137 ( .A1(n4030), .A2(n21570), .ZN(n14776) );
  AND2_X1 U140 ( .A1(n53736), .A2(n53740), .Z(n53756) );
  INV_X1 U145 ( .I(n53969), .ZN(n53926) );
  NAND2_X1 U147 ( .A1(n60426), .A2(n54012), .ZN(n53902) );
  NOR2_X1 U148 ( .A1(n54768), .A2(n22385), .ZN(n54754) );
  CLKBUF_X2 U150 ( .I(n1281), .Z(n63767) );
  BUF_X2 U155 ( .I(n53736), .Z(n25115) );
  NAND2_X1 U156 ( .A1(n23453), .A2(n18422), .ZN(n14552) );
  AND2_X1 U157 ( .A1(n55132), .A2(n55170), .Z(n61761) );
  NAND2_X1 U165 ( .A1(n20985), .A2(n5324), .ZN(n54368) );
  NAND2_X1 U166 ( .A1(n16943), .A2(n22683), .ZN(n55228) );
  NAND2_X1 U169 ( .A1(n55643), .A2(n62550), .ZN(n62549) );
  NAND2_X1 U171 ( .A1(n54006), .A2(n54012), .ZN(n54009) );
  NAND2_X1 U174 ( .A1(n62579), .A2(n62578), .ZN(n62577) );
  AND2_X1 U178 ( .A1(n64897), .A2(n17180), .Z(n63006) );
  INV_X1 U179 ( .I(n58825), .ZN(n53817) );
  BUF_X2 U181 ( .I(n53901), .Z(n22669) );
  CLKBUF_X2 U183 ( .I(n22755), .Z(n5614) );
  NAND2_X1 U192 ( .A1(n17795), .A2(n23163), .ZN(n56454) );
  INV_X1 U194 ( .I(n8194), .ZN(n62550) );
  INV_X2 U196 ( .I(n10507), .ZN(n56892) );
  NAND2_X1 U198 ( .A1(n57146), .A2(n57109), .ZN(n64585) );
  INV_X8 U202 ( .I(n63591), .ZN(n56106) );
  BUF_X4 U205 ( .I(n52216), .Z(n55627) );
  INV_X2 U207 ( .I(n55164), .ZN(n55157) );
  INV_X1 U222 ( .I(n57146), .ZN(n57122) );
  NOR2_X1 U227 ( .A1(n61817), .A2(n65117), .ZN(n15951) );
  NAND2_X1 U233 ( .A1(n56998), .A2(n15924), .ZN(n62339) );
  NOR2_X1 U236 ( .A1(n62178), .A2(n61840), .ZN(n62599) );
  AND2_X1 U239 ( .A1(n54783), .A2(n54958), .Z(n61723) );
  NOR2_X1 U240 ( .A1(n64730), .A2(n64729), .ZN(n13230) );
  NAND2_X1 U242 ( .A1(n20239), .A2(n60236), .ZN(n64543) );
  NAND3_X1 U243 ( .A1(n51776), .A2(n54977), .A3(n51780), .ZN(n63122) );
  NOR2_X1 U244 ( .A1(n56263), .A2(n55932), .ZN(n55933) );
  NAND2_X1 U245 ( .A1(n64842), .A2(n64841), .ZN(n64840) );
  AOI21_X1 U246 ( .A1(n52662), .A2(n63781), .B(n52661), .ZN(n63884) );
  NAND2_X1 U249 ( .A1(n64038), .A2(n64037), .ZN(n5053) );
  AOI22_X1 U253 ( .A1(n6944), .A2(n56566), .B1(n56565), .B2(n56564), .ZN(
        n63648) );
  NAND4_X1 U255 ( .A1(n54352), .A2(n6676), .A3(n54351), .A4(n54353), .ZN(n6675) );
  NAND2_X1 U258 ( .A1(n2890), .A2(n20383), .ZN(n53879) );
  AOI21_X1 U260 ( .A1(n55272), .A2(n55273), .B(n64479), .ZN(n24527) );
  OAI21_X1 U261 ( .A1(n63138), .A2(n63137), .B(n12469), .ZN(n57924) );
  NOR2_X1 U262 ( .A1(n62960), .A2(n55258), .ZN(n14429) );
  NAND2_X1 U263 ( .A1(n57038), .A2(n8446), .ZN(n64836) );
  AOI21_X1 U270 ( .A1(n24637), .A2(n20610), .B(n24636), .ZN(n64820) );
  NAND2_X1 U271 ( .A1(n22588), .A2(n55739), .ZN(n62558) );
  NAND3_X1 U272 ( .A1(n61693), .A2(n22114), .A3(n20982), .ZN(n64078) );
  NAND2_X1 U278 ( .A1(n62329), .A2(n62328), .ZN(n62327) );
  INV_X1 U282 ( .I(n53614), .ZN(n62513) );
  NAND2_X1 U284 ( .A1(n53609), .A2(n52843), .ZN(n63268) );
  NOR2_X1 U285 ( .A1(n57083), .A2(n52863), .ZN(n52252) );
  BUF_X2 U287 ( .I(n54597), .Z(n64307) );
  INV_X1 U288 ( .I(n54437), .ZN(n6311) );
  INV_X1 U289 ( .I(n54945), .ZN(n64879) );
  AND2_X1 U290 ( .A1(n2104), .A2(n61282), .Z(n61769) );
  INV_X2 U294 ( .I(n23025), .ZN(n64521) );
  NAND2_X1 U295 ( .A1(n62343), .A2(n22884), .ZN(n53426) );
  NAND3_X1 U297 ( .A1(n59764), .A2(n25080), .A3(n54502), .ZN(n54500) );
  NAND3_X1 U299 ( .A1(n6792), .A2(n53590), .A3(n53009), .ZN(n9765) );
  CLKBUF_X1 U301 ( .I(n5140), .Z(n62648) );
  NOR2_X1 U320 ( .A1(n62682), .A2(n53621), .ZN(n53856) );
  NOR2_X1 U322 ( .A1(n62868), .A2(n18750), .ZN(n57185) );
  NOR2_X1 U325 ( .A1(n13920), .A2(n61528), .ZN(n56992) );
  NAND2_X1 U329 ( .A1(n19187), .A2(n55277), .ZN(n64479) );
  INV_X1 U338 ( .I(n15281), .ZN(n14469) );
  INV_X1 U343 ( .I(n57002), .ZN(n52264) );
  NOR2_X1 U352 ( .A1(n6531), .A2(n55470), .ZN(n52931) );
  NOR2_X1 U353 ( .A1(n56365), .A2(n17860), .ZN(n63137) );
  NOR2_X1 U355 ( .A1(n11375), .A2(n61123), .ZN(n62900) );
  NOR2_X1 U357 ( .A1(n10425), .A2(n54102), .ZN(n20383) );
  NAND2_X1 U359 ( .A1(n61405), .A2(n64031), .ZN(n64030) );
  NAND3_X1 U362 ( .A1(n1612), .A2(n57031), .A3(n4181), .ZN(n50738) );
  AOI21_X1 U363 ( .A1(n56417), .A2(n23165), .B(n63038), .ZN(n63360) );
  INV_X1 U368 ( .I(n56631), .ZN(n1286) );
  INV_X1 U373 ( .I(n15434), .ZN(n4184) );
  BUF_X2 U375 ( .I(n56539), .Z(n22229) );
  BUF_X2 U377 ( .I(n60710), .Z(n64657) );
  BUF_X2 U381 ( .I(n53214), .Z(n4181) );
  INV_X1 U384 ( .I(n52975), .ZN(n717) );
  CLKBUF_X2 U388 ( .I(n54501), .Z(n59764) );
  CLKBUF_X2 U393 ( .I(n18247), .Z(n62760) );
  CLKBUF_X2 U399 ( .I(n53376), .Z(n23974) );
  CLKBUF_X2 U404 ( .I(n54025), .Z(n23482) );
  INV_X1 U405 ( .I(n23784), .ZN(n62330) );
  NAND2_X1 U407 ( .A1(n58490), .A2(n55739), .ZN(n55465) );
  NAND3_X1 U413 ( .A1(n21028), .A2(n53444), .A3(n53443), .ZN(n62370) );
  NOR2_X1 U419 ( .A1(n14468), .A2(n15281), .ZN(n14467) );
  NAND2_X1 U422 ( .A1(n18291), .A2(n8203), .ZN(n52046) );
  BUF_X4 U431 ( .I(n51633), .Z(n54814) );
  INV_X1 U442 ( .I(n52786), .ZN(n57047) );
  CLKBUF_X2 U443 ( .I(n2951), .Z(n59831) );
  BUF_X2 U444 ( .I(n24352), .Z(n7095) );
  CLKBUF_X2 U445 ( .I(n19556), .Z(n23047) );
  AND2_X1 U448 ( .A1(n55275), .A2(n19167), .Z(n55267) );
  BUF_X2 U450 ( .I(n56414), .Z(n23165) );
  NOR2_X1 U451 ( .A1(n9160), .A2(n1459), .ZN(n2959) );
  CLKBUF_X2 U452 ( .I(n6095), .Z(n22760) );
  BUF_X2 U453 ( .I(n63555), .Z(n61736) );
  CLKBUF_X2 U455 ( .I(n54492), .Z(n7532) );
  CLKBUF_X2 U456 ( .I(n1326), .Z(n10113) );
  BUF_X2 U457 ( .I(n53023), .Z(n61147) );
  NAND3_X1 U461 ( .A1(n52837), .A2(n53198), .A3(n13292), .ZN(n59009) );
  INV_X2 U466 ( .I(n54025), .ZN(n54347) );
  INV_X8 U469 ( .I(n56539), .ZN(n24669) );
  INV_X2 U472 ( .I(n53383), .ZN(n52840) );
  INV_X1 U480 ( .I(n12605), .ZN(n55934) );
  BUF_X2 U481 ( .I(n52211), .Z(n55470) );
  NAND2_X1 U489 ( .A1(n52977), .A2(n14446), .ZN(n54039) );
  INV_X1 U493 ( .I(n13485), .ZN(n21343) );
  INV_X2 U503 ( .I(n53905), .ZN(n54058) );
  INV_X1 U507 ( .I(n63705), .ZN(n24748) );
  CLKBUF_X1 U510 ( .I(n4031), .Z(n63035) );
  INV_X1 U512 ( .I(n246), .ZN(n2406) );
  BUF_X2 U513 ( .I(n52505), .Z(n724) );
  BUF_X2 U515 ( .I(n24368), .Z(n2801) );
  CLKBUF_X4 U517 ( .I(n51572), .Z(n62574) );
  CLKBUF_X2 U525 ( .I(n6596), .Z(n22373) );
  INV_X1 U532 ( .I(n52629), .ZN(n1621) );
  INV_X1 U535 ( .I(n2604), .ZN(n51374) );
  INV_X1 U537 ( .I(n4894), .ZN(n26087) );
  BUF_X2 U542 ( .I(n52192), .Z(n52420) );
  BUF_X4 U543 ( .I(n52334), .Z(n24076) );
  BUF_X2 U548 ( .I(n11742), .Z(n11741) );
  BUF_X2 U550 ( .I(n52587), .Z(n10335) );
  BUF_X2 U557 ( .I(n6298), .Z(n6004) );
  BUF_X2 U562 ( .I(n16389), .Z(n59854) );
  INV_X1 U563 ( .I(n65279), .ZN(n20021) );
  INV_X1 U565 ( .I(n62183), .ZN(n25618) );
  BUF_X2 U568 ( .I(n25970), .Z(n61178) );
  BUF_X2 U569 ( .I(n17127), .Z(n6336) );
  NAND2_X1 U573 ( .A1(n62553), .A2(n58390), .ZN(n12800) );
  NOR2_X1 U578 ( .A1(n45999), .A2(n45998), .ZN(n46011) );
  NAND3_X1 U579 ( .A1(n61774), .A2(n58271), .A3(n49857), .ZN(n57310) );
  NAND2_X1 U586 ( .A1(n64478), .A2(n9069), .ZN(n60966) );
  OR2_X1 U590 ( .A1(n696), .A2(n49452), .Z(n61774) );
  INV_X1 U591 ( .I(n2630), .ZN(n18084) );
  NAND2_X1 U595 ( .A1(n47914), .A2(n47913), .ZN(n13490) );
  AOI22_X1 U597 ( .A1(n22173), .A2(n57355), .B1(n4302), .B2(n47975), .ZN(n4301) );
  OAI21_X1 U599 ( .A1(n48797), .A2(n48796), .B(n48795), .ZN(n62811) );
  NAND2_X1 U601 ( .A1(n62561), .A2(n62086), .ZN(n63291) );
  OAI22_X1 U604 ( .A1(n1117), .A2(n9442), .B1(n49316), .B2(n9443), .ZN(n62563)
         );
  NAND2_X1 U605 ( .A1(n14211), .A2(n62274), .ZN(n14210) );
  NAND2_X1 U609 ( .A1(n62915), .A2(n17693), .ZN(n6366) );
  NOR2_X1 U612 ( .A1(n64288), .A2(n49492), .ZN(n19437) );
  NOR2_X1 U615 ( .A1(n49308), .A2(n49608), .ZN(n11820) );
  NOR2_X1 U616 ( .A1(n64161), .A2(n64162), .ZN(n64539) );
  AOI21_X1 U619 ( .A1(n1067), .A2(n62255), .B(n8992), .ZN(n63192) );
  NAND2_X1 U621 ( .A1(n59718), .A2(n59717), .ZN(n63197) );
  AOI22_X1 U625 ( .A1(n59640), .A2(n49432), .B1(n48909), .B2(n48908), .ZN(
        n48910) );
  NAND2_X1 U627 ( .A1(n49524), .A2(n24821), .ZN(n14211) );
  OAI21_X1 U635 ( .A1(n46261), .A2(n63802), .B(n46370), .ZN(n10577) );
  NAND3_X1 U638 ( .A1(n49678), .A2(n61258), .A3(n49679), .ZN(n7147) );
  NOR2_X1 U640 ( .A1(n50342), .A2(n60467), .ZN(n58676) );
  OAI22_X1 U644 ( .A1(n3044), .A2(n62946), .B1(n50058), .B2(n50304), .ZN(n3043) );
  NAND4_X1 U647 ( .A1(n11114), .A2(n48381), .A3(n49634), .A4(n48386), .ZN(
        n62915) );
  AOI21_X1 U651 ( .A1(n49299), .A2(n49298), .B(n64326), .ZN(n49306) );
  NAND3_X1 U654 ( .A1(n47354), .A2(n5661), .A3(n61016), .ZN(n5703) );
  INV_X1 U655 ( .I(n49377), .ZN(n64561) );
  NAND3_X1 U656 ( .A1(n63959), .A2(n45923), .A3(n63958), .ZN(n61241) );
  NAND3_X1 U658 ( .A1(n23156), .A2(n25018), .A3(n1640), .ZN(n48418) );
  INV_X1 U660 ( .I(n6323), .ZN(n11867) );
  NOR2_X1 U664 ( .A1(n61742), .A2(n6411), .ZN(n10915) );
  OR2_X1 U670 ( .A1(n20311), .A2(n13440), .Z(n61776) );
  AND2_X1 U674 ( .A1(n48295), .A2(n48299), .Z(n61773) );
  NOR2_X1 U675 ( .A1(n64303), .A2(n48305), .ZN(n61972) );
  NAND3_X1 U677 ( .A1(n3703), .A2(n61150), .A3(n61151), .ZN(n3702) );
  NAND3_X1 U682 ( .A1(n50342), .A2(n50341), .A3(n50340), .ZN(n50343) );
  NAND4_X1 U689 ( .A1(n12475), .A2(n8355), .A3(n5188), .A4(n25081), .ZN(n5187)
         );
  OAI22_X1 U698 ( .A1(n16193), .A2(n49089), .B1(n48012), .B2(n48011), .ZN(
        n64529) );
  NAND2_X1 U700 ( .A1(n25783), .A2(n49490), .ZN(n64288) );
  NOR2_X1 U701 ( .A1(n48823), .A2(n739), .ZN(n5701) );
  NAND2_X1 U702 ( .A1(n48950), .A2(n57735), .ZN(n22171) );
  NOR2_X1 U706 ( .A1(n49411), .A2(n8789), .ZN(n58551) );
  NAND2_X1 U708 ( .A1(n49266), .A2(n46369), .ZN(n63802) );
  OAI21_X1 U709 ( .A1(n64669), .A2(n64668), .B(n49391), .ZN(n49400) );
  NAND2_X1 U713 ( .A1(n24694), .A2(n16030), .ZN(n62807) );
  NOR2_X1 U718 ( .A1(n49619), .A2(n49039), .ZN(n21491) );
  NAND2_X1 U720 ( .A1(n2889), .A2(n49383), .ZN(n7758) );
  INV_X1 U721 ( .I(n49504), .ZN(n64336) );
  NOR2_X1 U724 ( .A1(n11623), .A2(n13118), .ZN(n48319) );
  NAND2_X1 U726 ( .A1(n2514), .A2(n7146), .ZN(n62007) );
  NOR2_X1 U728 ( .A1(n64990), .A2(n24069), .ZN(n63358) );
  NOR2_X1 U731 ( .A1(n24643), .A2(n49705), .ZN(n64161) );
  NOR2_X1 U732 ( .A1(n49947), .A2(n61170), .ZN(n63958) );
  OAI22_X1 U734 ( .A1(n49296), .A2(n20363), .B1(n9354), .B2(n49301), .ZN(
        n64326) );
  NOR2_X1 U735 ( .A1(n63369), .A2(n50421), .ZN(n63368) );
  INV_X1 U738 ( .I(n17886), .ZN(n50441) );
  NAND2_X1 U739 ( .A1(n65135), .A2(n49074), .ZN(n47449) );
  NOR2_X1 U742 ( .A1(n8380), .A2(n50044), .ZN(n49440) );
  OR2_X1 U744 ( .A1(n1631), .A2(n48701), .Z(n49490) );
  NAND2_X1 U745 ( .A1(n50367), .A2(n3462), .ZN(n62499) );
  NOR2_X1 U748 ( .A1(n16985), .A2(n49281), .ZN(n11458) );
  NAND3_X1 U749 ( .A1(n60360), .A2(n22264), .A3(n23299), .ZN(n14353) );
  NAND2_X1 U750 ( .A1(n60648), .A2(n16595), .ZN(n49460) );
  NAND3_X1 U754 ( .A1(n11467), .A2(n60726), .A3(n47989), .ZN(n7485) );
  NAND2_X1 U755 ( .A1(n1377), .A2(n64404), .ZN(n50285) );
  NOR2_X1 U761 ( .A1(n64935), .A2(n64936), .ZN(n24643) );
  CLKBUF_X1 U763 ( .I(n9772), .Z(n63202) );
  NAND2_X1 U765 ( .A1(n16411), .A2(n22457), .ZN(n49275) );
  INV_X1 U767 ( .I(n47977), .ZN(n12845) );
  NOR2_X1 U770 ( .A1(n49763), .A2(n49764), .ZN(n64862) );
  NOR2_X1 U773 ( .A1(n61742), .A2(n48803), .ZN(n48346) );
  NAND2_X1 U777 ( .A1(n16595), .A2(n45231), .ZN(n64661) );
  NOR2_X1 U778 ( .A1(n49390), .A2(n49389), .ZN(n64669) );
  INV_X1 U785 ( .I(n49942), .ZN(n63959) );
  NAND3_X1 U790 ( .A1(n11950), .A2(n7990), .A3(n49063), .ZN(n48295) );
  NAND2_X1 U793 ( .A1(n15319), .A2(n18975), .ZN(n49567) );
  NAND2_X1 U796 ( .A1(n50123), .A2(n1224), .ZN(n63621) );
  BUF_X2 U798 ( .I(n5498), .Z(n5463) );
  NAND2_X1 U800 ( .A1(n49674), .A2(n11153), .ZN(n49093) );
  OR2_X1 U803 ( .A1(n61673), .A2(n49195), .Z(n61833) );
  NOR2_X1 U811 ( .A1(n6411), .A2(n48790), .ZN(n48798) );
  NAND2_X1 U817 ( .A1(n22694), .A2(n1209), .ZN(n48026) );
  NAND2_X1 U827 ( .A1(n26000), .A2(n20600), .ZN(n5743) );
  NAND2_X1 U830 ( .A1(n62653), .A2(n49319), .ZN(n49608) );
  NOR2_X1 U832 ( .A1(n15386), .A2(n5283), .ZN(n47935) );
  INV_X1 U834 ( .I(n60726), .ZN(n62905) );
  NAND2_X1 U844 ( .A1(n49676), .A2(n5498), .ZN(n49682) );
  BUF_X2 U850 ( .I(n49277), .Z(n16411) );
  CLKBUF_X2 U851 ( .I(n19646), .Z(n63605) );
  INV_X1 U856 ( .I(n2433), .ZN(n62927) );
  NAND2_X1 U862 ( .A1(n4724), .A2(n17335), .ZN(n49495) );
  NAND2_X1 U863 ( .A1(n49844), .A2(n49452), .ZN(n64206) );
  CLKBUF_X2 U865 ( .I(n49286), .Z(n64488) );
  AND2_X1 U866 ( .A1(n3658), .A2(n49637), .Z(n61867) );
  BUF_X2 U868 ( .I(n49053), .Z(n3971) );
  INV_X1 U869 ( .I(n48847), .ZN(n62744) );
  BUF_X2 U877 ( .I(n46367), .Z(n49410) );
  NAND2_X1 U879 ( .A1(n61070), .A2(n58205), .ZN(n49450) );
  NAND2_X1 U883 ( .A1(n48341), .A2(n49908), .ZN(n48734) );
  BUF_X2 U891 ( .I(n2736), .Z(n78) );
  NOR2_X1 U892 ( .A1(n62653), .A2(n49319), .ZN(n10761) );
  NOR2_X1 U905 ( .A1(n502), .A2(n49641), .ZN(n47796) );
  BUF_X4 U908 ( .I(n9229), .Z(n64562) );
  INV_X2 U909 ( .I(n9346), .ZN(n8790) );
  INV_X1 U911 ( .I(n46850), .ZN(n1327) );
  INV_X2 U918 ( .I(n11037), .ZN(n8044) );
  BUF_X2 U919 ( .I(n25320), .Z(n1639) );
  CLKBUF_X2 U921 ( .I(n49923), .Z(n19523) );
  NAND2_X1 U927 ( .A1(n15424), .A2(n63602), .ZN(n63865) );
  NOR3_X1 U928 ( .A1(n45440), .A2(n58800), .A3(n45439), .ZN(n62659) );
  NOR2_X1 U930 ( .A1(n21620), .A2(n46056), .ZN(n63145) );
  NAND3_X1 U940 ( .A1(n22602), .A2(n44208), .A3(n22603), .ZN(n63059) );
  NAND3_X1 U946 ( .A1(n48671), .A2(n48670), .A3(n48669), .ZN(n62238) );
  OAI21_X1 U949 ( .A1(n20970), .A2(n47752), .B(n62114), .ZN(n18982) );
  NAND2_X1 U953 ( .A1(n59505), .A2(n46918), .ZN(n63829) );
  AOI22_X1 U959 ( .A1(n64293), .A2(n48581), .B1(n12767), .B2(n12766), .ZN(
        n58068) );
  AOI21_X1 U966 ( .A1(n47855), .A2(n47399), .B(n63363), .ZN(n47403) );
  OR2_X1 U974 ( .A1(n48603), .A2(n61422), .Z(n61722) );
  AND2_X1 U975 ( .A1(n47187), .A2(n46716), .Z(n61876) );
  NOR2_X1 U976 ( .A1(n6651), .A2(n6662), .ZN(n63401) );
  OAI21_X1 U977 ( .A1(n62484), .A2(n61966), .B(n47513), .ZN(n47521) );
  NOR3_X1 U981 ( .A1(n20861), .A2(n16093), .A3(n19229), .ZN(n64711) );
  NOR2_X1 U982 ( .A1(n62131), .A2(n62130), .ZN(n5482) );
  NAND2_X1 U995 ( .A1(n46822), .A2(n46746), .ZN(n63418) );
  OAI21_X1 U997 ( .A1(n64313), .A2(n61862), .B(n59528), .ZN(n25863) );
  NAND2_X1 U1000 ( .A1(n48079), .A2(n48078), .ZN(n48092) );
  NOR3_X1 U1007 ( .A1(n63585), .A2(n6788), .A3(n63584), .ZN(n44566) );
  NOR2_X1 U1009 ( .A1(n23361), .A2(n2640), .ZN(n25281) );
  NAND2_X1 U1012 ( .A1(n19931), .A2(n20307), .ZN(n65215) );
  AOI21_X1 U1014 ( .A1(n46015), .A2(n1661), .B(n46014), .ZN(n61974) );
  OAI21_X1 U1016 ( .A1(n13472), .A2(n5202), .B(n23018), .ZN(n63452) );
  NAND2_X1 U1017 ( .A1(n12700), .A2(n46817), .ZN(n10450) );
  INV_X1 U1022 ( .I(n10910), .ZN(n64123) );
  NAND2_X1 U1024 ( .A1(n47512), .A2(n47511), .ZN(n62484) );
  NOR2_X1 U1025 ( .A1(n47568), .A2(n45948), .ZN(n65012) );
  OAI21_X1 U1026 ( .A1(n45602), .A2(n20666), .B(n344), .ZN(n46023) );
  NAND2_X1 U1030 ( .A1(n48258), .A2(n62824), .ZN(n62823) );
  NAND2_X1 U1034 ( .A1(n62181), .A2(n62180), .ZN(n19683) );
  NAND2_X1 U1037 ( .A1(n63706), .A2(n47529), .ZN(n19931) );
  INV_X1 U1038 ( .I(n48626), .ZN(n64913) );
  NAND2_X1 U1041 ( .A1(n13348), .A2(n48085), .ZN(n62121) );
  NAND2_X1 U1045 ( .A1(n24114), .A2(n47828), .ZN(n65024) );
  NOR3_X1 U1050 ( .A1(n64441), .A2(n64440), .A3(n45730), .ZN(n44657) );
  NAND2_X1 U1060 ( .A1(n48552), .A2(n57973), .ZN(n48150) );
  NAND2_X1 U1061 ( .A1(n48096), .A2(n45805), .ZN(n23925) );
  NOR2_X1 U1071 ( .A1(n16375), .A2(n47559), .ZN(n62021) );
  NAND2_X1 U1072 ( .A1(n1080), .A2(n46948), .ZN(n63309) );
  NAND2_X1 U1075 ( .A1(n47161), .A2(n48481), .ZN(n46472) );
  NOR2_X1 U1076 ( .A1(n48506), .A2(n12968), .ZN(n63135) );
  AOI22_X1 U1082 ( .A1(n46474), .A2(n46475), .B1(n46473), .B2(n2403), .ZN(
        n63523) );
  NOR2_X1 U1083 ( .A1(n64960), .A2(n6786), .ZN(n63584) );
  OAI22_X1 U1088 ( .A1(n48096), .A2(n45804), .B1(n11692), .B2(n11087), .ZN(
        n11691) );
  NOR3_X1 U1097 ( .A1(n47752), .A2(n18590), .A3(n47744), .ZN(n46742) );
  NAND4_X1 U1100 ( .A1(n7161), .A2(n46863), .A3(n46028), .A4(n46027), .ZN(
        n64296) );
  AOI22_X1 U1102 ( .A1(n47369), .A2(n47370), .B1(n21451), .B2(n65161), .ZN(
        n47375) );
  INV_X1 U1107 ( .I(n48234), .ZN(n57728) );
  NAND2_X1 U1109 ( .A1(n60727), .A2(n7191), .ZN(n62181) );
  INV_X1 U1111 ( .I(n2743), .ZN(n63710) );
  NAND2_X1 U1123 ( .A1(n64683), .A2(n14448), .ZN(n46949) );
  NAND3_X1 U1126 ( .A1(n46951), .A2(n23113), .A3(n16686), .ZN(n45495) );
  NAND4_X1 U1136 ( .A1(n24354), .A2(n23850), .A3(n21304), .A4(n16950), .ZN(
        n48098) );
  INV_X1 U1138 ( .I(n23361), .ZN(n1658) );
  NAND2_X1 U1140 ( .A1(n61719), .A2(n8138), .ZN(n58991) );
  NOR2_X1 U1145 ( .A1(n5771), .A2(n25148), .ZN(n63837) );
  OAI21_X1 U1151 ( .A1(n10979), .A2(n61675), .B(n48575), .ZN(n61625) );
  NAND2_X1 U1153 ( .A1(n47168), .A2(n48626), .ZN(n64597) );
  NOR2_X1 U1154 ( .A1(n61967), .A2(n9505), .ZN(n45679) );
  NAND3_X1 U1156 ( .A1(n48561), .A2(n48085), .A3(n63871), .ZN(n48086) );
  AOI21_X1 U1161 ( .A1(n48506), .A2(n57762), .B(n61861), .ZN(n62824) );
  NAND3_X1 U1164 ( .A1(n44401), .A2(n20938), .A3(n21755), .ZN(n44399) );
  INV_X1 U1172 ( .I(n18099), .ZN(n48153) );
  NAND3_X1 U1178 ( .A1(n47233), .A2(n47232), .A3(n60038), .ZN(n64466) );
  OAI21_X1 U1180 ( .A1(n45550), .A2(n5554), .B(n5145), .ZN(n16373) );
  NOR2_X1 U1185 ( .A1(n8012), .A2(n24820), .ZN(n44692) );
  INV_X1 U1186 ( .I(n57731), .ZN(n64386) );
  NAND3_X1 U1188 ( .A1(n2664), .A2(n9758), .A3(n64899), .ZN(n46936) );
  CLKBUF_X2 U1189 ( .I(n48095), .Z(n62755) );
  AND2_X1 U1190 ( .A1(n47851), .A2(n25007), .Z(n13782) );
  INV_X1 U1192 ( .I(n47834), .ZN(n45550) );
  NAND2_X1 U1199 ( .A1(n45536), .A2(n19595), .ZN(n45783) );
  OR2_X1 U1202 ( .A1(n1386), .A2(n46753), .Z(n48149) );
  AND2_X1 U1204 ( .A1(n22508), .A2(n25896), .Z(n61756) );
  AND2_X1 U1205 ( .A1(n25702), .A2(n45551), .Z(n61967) );
  NAND2_X1 U1208 ( .A1(n46882), .A2(n6148), .ZN(n5934) );
  OR2_X1 U1219 ( .A1(n47080), .A2(n14521), .Z(n61719) );
  NOR2_X1 U1220 ( .A1(n57670), .A2(n1294), .ZN(n44401) );
  INV_X1 U1229 ( .I(n17905), .ZN(n15276) );
  NAND2_X1 U1238 ( .A1(n61718), .A2(n48191), .ZN(n48203) );
  CLKBUF_X2 U1239 ( .I(n48252), .Z(n64922) );
  NAND3_X1 U1240 ( .A1(n47535), .A2(n47529), .A3(n22684), .ZN(n48602) );
  INV_X1 U1247 ( .I(n63144), .ZN(n46052) );
  BUF_X4 U1250 ( .I(n46874), .Z(n20426) );
  OR2_X1 U1261 ( .A1(n63017), .A2(n10364), .Z(n16628) );
  INV_X1 U1262 ( .I(n23894), .ZN(n45961) );
  AND2_X1 U1264 ( .A1(n24615), .A2(n25841), .Z(n47810) );
  OR2_X1 U1267 ( .A1(n45551), .A2(n47274), .Z(n2223) );
  INV_X1 U1277 ( .I(n2955), .ZN(n62633) );
  NAND2_X1 U1280 ( .A1(n15697), .A2(n18196), .ZN(n64250) );
  INV_X1 U1289 ( .I(n48205), .ZN(n48191) );
  CLKBUF_X1 U1301 ( .I(n48644), .Z(n64791) );
  NAND2_X1 U1303 ( .A1(n1085), .A2(n47572), .ZN(n45592) );
  INV_X2 U1305 ( .I(n14521), .ZN(n15749) );
  INV_X1 U1308 ( .I(n48642), .ZN(n62046) );
  INV_X1 U1322 ( .I(n10193), .ZN(n2664) );
  NAND2_X1 U1323 ( .A1(n16533), .A2(n15757), .ZN(n48193) );
  AOI21_X1 U1324 ( .A1(n64347), .A2(n22386), .B(n19329), .ZN(n32) );
  NAND3_X1 U1327 ( .A1(n21793), .A2(n47250), .A3(n60753), .ZN(n47254) );
  INV_X1 U1332 ( .I(n47580), .ZN(n45683) );
  INV_X1 U1333 ( .I(n44705), .ZN(n62110) );
  CLKBUF_X2 U1337 ( .I(n16020), .Z(n63793) );
  INV_X2 U1338 ( .I(n43750), .ZN(n47434) );
  INV_X1 U1347 ( .I(n46244), .ZN(n48668) );
  INV_X1 U1350 ( .I(n1652), .ZN(n47818) );
  INV_X2 U1351 ( .I(n64347), .ZN(n23894) );
  BUF_X2 U1356 ( .I(n46148), .Z(n8758) );
  BUF_X2 U1358 ( .I(n15871), .Z(n60753) );
  CLKBUF_X2 U1372 ( .I(n6157), .Z(n57637) );
  CLKBUF_X2 U1374 ( .I(n47749), .Z(n24081) );
  INV_X2 U1379 ( .I(n2024), .ZN(n58233) );
  BUF_X8 U1394 ( .I(n8525), .Z(n3510) );
  BUF_X4 U1400 ( .I(n47491), .Z(n16533) );
  INV_X1 U1403 ( .I(n10447), .ZN(n19680) );
  INV_X1 U1404 ( .I(n11339), .ZN(n62926) );
  CLKBUF_X2 U1411 ( .I(n45401), .Z(n61490) );
  INV_X1 U1420 ( .I(n14935), .ZN(n61220) );
  CLKBUF_X2 U1421 ( .I(n18624), .Z(n7034) );
  BUF_X2 U1422 ( .I(n44549), .Z(n24112) );
  INV_X1 U1424 ( .I(n46319), .ZN(n1672) );
  INV_X1 U1426 ( .I(n45021), .ZN(n65250) );
  INV_X2 U1430 ( .I(n8598), .ZN(n64837) );
  INV_X1 U1433 ( .I(n63027), .ZN(n61988) );
  INV_X1 U1434 ( .I(n1198), .ZN(n58212) );
  CLKBUF_X2 U1436 ( .I(n45030), .Z(n23210) );
  BUF_X2 U1437 ( .I(n44156), .Z(n46650) );
  CLKBUF_X2 U1439 ( .I(n22396), .Z(n64373) );
  BUF_X2 U1442 ( .I(n59382), .Z(n24521) );
  INV_X1 U1446 ( .I(n6678), .ZN(n5093) );
  INV_X1 U1450 ( .I(n20758), .ZN(n44169) );
  NAND2_X1 U1454 ( .A1(n63005), .A2(n14373), .ZN(n13868) );
  NOR2_X1 U1456 ( .A1(n59443), .A2(n14857), .ZN(n14856) );
  BUF_X2 U1457 ( .I(n6136), .Z(n3208) );
  NAND2_X1 U1459 ( .A1(n10258), .A2(n13108), .ZN(n22973) );
  BUF_X2 U1461 ( .I(n21940), .Z(n10619) );
  CLKBUF_X2 U1462 ( .I(n6678), .Z(n6677) );
  BUF_X2 U1463 ( .I(n44735), .Z(n59866) );
  NOR2_X1 U1471 ( .A1(n5327), .A2(n5326), .ZN(n62622) );
  NAND2_X1 U1473 ( .A1(n7819), .A2(n42974), .ZN(n14628) );
  NOR2_X1 U1475 ( .A1(n18297), .A2(n18299), .ZN(n62738) );
  NAND3_X1 U1477 ( .A1(n43560), .A2(n43558), .A3(n43559), .ZN(n63989) );
  NOR2_X1 U1484 ( .A1(n4551), .A2(n18405), .ZN(n62466) );
  NOR2_X1 U1490 ( .A1(n40687), .A2(n40688), .ZN(n40689) );
  OAI21_X1 U1498 ( .A1(n64380), .A2(n64379), .B(n64378), .ZN(n15279) );
  OAI21_X1 U1504 ( .A1(n15119), .A2(n18342), .B(n13873), .ZN(n13872) );
  INV_X1 U1512 ( .I(n10339), .ZN(n63872) );
  OAI21_X1 U1515 ( .A1(n8934), .A2(n57614), .B(n8937), .ZN(n8933) );
  NAND2_X1 U1522 ( .A1(n58965), .A2(n63380), .ZN(n15374) );
  NOR2_X1 U1530 ( .A1(n5930), .A2(n8349), .ZN(n62374) );
  NAND2_X1 U1535 ( .A1(n62847), .A2(n42861), .ZN(n65000) );
  NOR2_X1 U1541 ( .A1(n60230), .A2(n24764), .ZN(n24760) );
  NAND3_X1 U1545 ( .A1(n62269), .A2(n25757), .A3(n9822), .ZN(n8323) );
  OAI21_X1 U1546 ( .A1(n63479), .A2(n63478), .B(n4228), .ZN(n64588) );
  NOR2_X1 U1548 ( .A1(n42187), .A2(n42186), .ZN(n64127) );
  OAI21_X1 U1549 ( .A1(n64893), .A2(n64892), .B(n21851), .ZN(n24136) );
  OAI21_X1 U1550 ( .A1(n12137), .A2(n64226), .B(n42399), .ZN(n12135) );
  AOI21_X1 U1555 ( .A1(n10848), .A2(n14846), .B(n62567), .ZN(n7794) );
  OAI21_X1 U1556 ( .A1(n8786), .A2(n8785), .B(n63270), .ZN(n7795) );
  AOI22_X1 U1561 ( .A1(n42368), .A2(n24996), .B1(n16260), .B2(n42053), .ZN(
        n63068) );
  AOI22_X1 U1563 ( .A1(n42920), .A2(n42921), .B1(n13159), .B2(n42924), .ZN(
        n64569) );
  NOR2_X1 U1565 ( .A1(n6865), .A2(n43577), .ZN(n16201) );
  NAND4_X1 U1566 ( .A1(n43491), .A2(n43492), .A3(n43925), .A4(n43531), .ZN(
        n6070) );
  NAND4_X1 U1571 ( .A1(n42190), .A2(n42191), .A3(n57256), .A4(n42189), .ZN(
        n63104) );
  AOI21_X1 U1575 ( .A1(n8343), .A2(n43220), .B(n63095), .ZN(n2464) );
  AOI22_X1 U1584 ( .A1(n42975), .A2(n42804), .B1(n42805), .B2(n42980), .ZN(
        n42810) );
  INV_X1 U1597 ( .I(n18342), .ZN(n10355) );
  NOR2_X1 U1598 ( .A1(n58343), .A2(n42082), .ZN(n62239) );
  INV_X1 U1602 ( .I(n41321), .ZN(n62567) );
  OR2_X1 U1604 ( .A1(n43517), .A2(n25210), .Z(n61786) );
  NAND2_X1 U1605 ( .A1(n12932), .A2(n61171), .ZN(n1015) );
  NOR2_X1 U1610 ( .A1(n7877), .A2(n40453), .ZN(n42764) );
  NAND2_X1 U1612 ( .A1(n43327), .A2(n43325), .ZN(n41482) );
  NOR2_X1 U1616 ( .A1(n61397), .A2(n61395), .ZN(n9209) );
  NAND2_X1 U1624 ( .A1(n42542), .A2(n1297), .ZN(n12916) );
  NOR3_X1 U1628 ( .A1(n43129), .A2(n43130), .A3(n8962), .ZN(n43269) );
  OAI21_X1 U1629 ( .A1(n64333), .A2(n64332), .B(n64510), .ZN(n62269) );
  OR2_X1 U1630 ( .A1(n42717), .A2(n2994), .Z(n61891) );
  NAND2_X1 U1631 ( .A1(n25851), .A2(n62961), .ZN(n5719) );
  INV_X1 U1636 ( .I(n18363), .ZN(n63478) );
  NOR3_X1 U1643 ( .A1(n12043), .A2(n62391), .A3(n61976), .ZN(n12042) );
  OAI21_X1 U1644 ( .A1(n42181), .A2(n42788), .B(n64510), .ZN(n58191) );
  AOI21_X1 U1646 ( .A1(n11361), .A2(n24575), .B(n63482), .ZN(n3001) );
  NOR2_X1 U1647 ( .A1(n65129), .A2(n42067), .ZN(n62438) );
  NOR3_X1 U1649 ( .A1(n43454), .A2(n13750), .A3(n58530), .ZN(n42073) );
  NOR3_X1 U1655 ( .A1(n65181), .A2(n42827), .A3(n6705), .ZN(n64865) );
  NAND3_X1 U1656 ( .A1(n64323), .A2(n23279), .A3(n43655), .ZN(n62847) );
  AOI22_X1 U1660 ( .A1(n63276), .A2(n42604), .B1(n42602), .B2(n42601), .ZN(
        n42611) );
  NOR2_X1 U1663 ( .A1(n41726), .A2(n42353), .ZN(n23899) );
  NAND2_X1 U1672 ( .A1(n43275), .A2(n41711), .ZN(n62203) );
  NOR3_X1 U1673 ( .A1(n775), .A2(n42871), .A3(n63721), .ZN(n41505) );
  OAI21_X1 U1683 ( .A1(n1698), .A2(n42923), .B(n64363), .ZN(n13159) );
  NAND2_X1 U1686 ( .A1(n8213), .A2(n42917), .ZN(n42920) );
  NAND3_X1 U1689 ( .A1(n43338), .A2(n43337), .A3(n43341), .ZN(n18995) );
  NAND2_X1 U1690 ( .A1(n42940), .A2(n65179), .ZN(n42941) );
  OAI21_X1 U1692 ( .A1(n42860), .A2(n1692), .B(n42858), .ZN(n64104) );
  NAND2_X1 U1694 ( .A1(n64629), .A2(n61976), .ZN(n23622) );
  AOI22_X1 U1708 ( .A1(n20400), .A2(n42331), .B1(n42330), .B2(n42329), .ZN(
        n62367) );
  NOR2_X1 U1711 ( .A1(n57178), .A2(n24360), .ZN(n64892) );
  OAI22_X1 U1718 ( .A1(n6268), .A2(n42076), .B1(n58402), .B2(n42082), .ZN(
        n64226) );
  INV_X2 U1722 ( .I(n9792), .ZN(n64510) );
  AND2_X1 U1732 ( .A1(n41666), .A2(n42788), .Z(n777) );
  INV_X1 U1733 ( .I(n16659), .ZN(n63482) );
  INV_X1 U1737 ( .I(n19490), .ZN(n42078) );
  NOR2_X1 U1750 ( .A1(n42140), .A2(n42662), .ZN(n42669) );
  NAND2_X1 U1751 ( .A1(n25851), .A2(n13751), .ZN(n43454) );
  NOR2_X1 U1755 ( .A1(n59650), .A2(n23730), .ZN(n19487) );
  OR2_X1 U1762 ( .A1(n24386), .A2(n41549), .Z(n11223) );
  NAND2_X1 U1767 ( .A1(n62391), .A2(n8798), .ZN(n63276) );
  NAND2_X1 U1772 ( .A1(n42365), .A2(n40016), .ZN(n9366) );
  NOR2_X1 U1774 ( .A1(n41775), .A2(n1502), .ZN(n42343) );
  INV_X1 U1776 ( .I(n15031), .ZN(n23188) );
  NOR2_X1 U1778 ( .A1(n61951), .A2(n43897), .ZN(n43234) );
  NOR2_X1 U1781 ( .A1(n63091), .A2(n57177), .ZN(n43271) );
  NOR2_X1 U1782 ( .A1(n18019), .A2(n18020), .ZN(n15118) );
  CLKBUF_X2 U1784 ( .I(n1495), .Z(n64156) );
  OR2_X1 U1785 ( .A1(n62314), .A2(n1270), .Z(n41484) );
  INV_X1 U1786 ( .I(n62072), .ZN(n60836) );
  NOR2_X1 U1796 ( .A1(n42777), .A2(n42188), .ZN(n64333) );
  NAND3_X1 U1800 ( .A1(n43199), .A2(n13677), .A3(n13679), .ZN(n42643) );
  BUF_X2 U1806 ( .I(n42606), .Z(n61976) );
  NAND2_X1 U1807 ( .A1(n59309), .A2(n61107), .ZN(n12955) );
  AOI21_X1 U1810 ( .A1(n42976), .A2(n43327), .B(n63970), .ZN(n62332) );
  NAND2_X1 U1813 ( .A1(n42128), .A2(n42127), .ZN(n62388) );
  NOR2_X1 U1825 ( .A1(n43444), .A2(n58850), .ZN(n62467) );
  NOR2_X1 U1832 ( .A1(n42405), .A2(n42079), .ZN(n40872) );
  NOR2_X1 U1835 ( .A1(n60866), .A2(n61794), .ZN(n40023) );
  NAND2_X1 U1840 ( .A1(n1225), .A2(n43270), .ZN(n62899) );
  OAI22_X1 U1842 ( .A1(n42595), .A2(n42606), .B1(n59771), .B2(n42594), .ZN(
        n42596) );
  INV_X1 U1857 ( .I(n43023), .ZN(n64332) );
  NOR2_X1 U1861 ( .A1(n11229), .A2(n43601), .ZN(n2068) );
  OR2_X1 U1867 ( .A1(n24405), .A2(n15160), .Z(n43039) );
  OR2_X1 U1868 ( .A1(n13393), .A2(n42049), .Z(n43445) );
  INV_X1 U1871 ( .I(n6005), .ZN(n43714) );
  INV_X2 U1876 ( .I(n64363), .ZN(n9191) );
  NAND2_X1 U1878 ( .A1(n4437), .A2(n43319), .ZN(n15031) );
  NAND2_X1 U1879 ( .A1(n2557), .A2(n60548), .ZN(n25440) );
  NOR2_X1 U1882 ( .A1(n4198), .A2(n4077), .ZN(n41717) );
  NAND2_X1 U1885 ( .A1(n1501), .A2(n1301), .ZN(n4313) );
  BUF_X2 U1886 ( .I(n8361), .Z(n61344) );
  NAND2_X1 U1888 ( .A1(n43444), .A2(n65179), .ZN(n41744) );
  NOR2_X1 U1889 ( .A1(n43161), .A2(n61237), .ZN(n42566) );
  NAND2_X1 U1892 ( .A1(n12386), .A2(n2735), .ZN(n16659) );
  CLKBUF_X2 U1897 ( .I(n16447), .Z(n63983) );
  INV_X1 U1898 ( .I(n43299), .ZN(n63778) );
  NAND2_X1 U1914 ( .A1(n41665), .A2(n63666), .ZN(n57283) );
  AND2_X1 U1915 ( .A1(n43242), .A2(n24195), .Z(n8018) );
  NAND2_X1 U1920 ( .A1(n57198), .A2(n43460), .ZN(n62963) );
  NOR2_X1 U1926 ( .A1(n1008), .A2(n63437), .ZN(n63341) );
  AOI22_X1 U1928 ( .A1(n43167), .A2(n43168), .B1(n43169), .B2(n43170), .ZN(
        n64302) );
  INV_X1 U1932 ( .I(n13751), .ZN(n62962) );
  INV_X2 U1936 ( .I(n40015), .ZN(n43449) );
  BUF_X2 U1941 ( .I(n12312), .Z(n62686) );
  NOR2_X1 U1945 ( .A1(n5126), .A2(n42598), .ZN(n37535) );
  INV_X1 U1952 ( .I(n41963), .ZN(n41656) );
  NAND2_X1 U1954 ( .A1(n8361), .A2(n42784), .ZN(n43024) );
  INV_X2 U1956 ( .I(n43242), .ZN(n43898) );
  NOR2_X1 U1962 ( .A1(n59425), .A2(n59426), .ZN(n1008) );
  INV_X2 U1964 ( .I(n43852), .ZN(n10990) );
  BUF_X1 U1965 ( .I(n4198), .Z(n4199) );
  NOR2_X1 U1981 ( .A1(n59263), .A2(n25534), .ZN(n42074) );
  INV_X2 U1982 ( .I(n15029), .ZN(n61745) );
  NAND2_X1 U1985 ( .A1(n57810), .A2(n16710), .ZN(n43677) );
  INV_X1 U1999 ( .I(n64292), .ZN(n43184) );
  BUF_X2 U2000 ( .I(n40776), .Z(n43517) );
  INV_X2 U2010 ( .I(n43693), .ZN(n1705) );
  INV_X2 U2022 ( .I(n43382), .ZN(n25412) );
  OR2_X1 U2029 ( .A1(n20276), .A2(n61164), .Z(n57255) );
  INV_X2 U2035 ( .I(n8361), .ZN(n63666) );
  NAND2_X1 U2037 ( .A1(n64391), .A2(n19241), .ZN(n42084) );
  INV_X1 U2045 ( .I(n41538), .ZN(n57454) );
  NAND3_X1 U2055 ( .A1(n64709), .A2(n41400), .A3(n39049), .ZN(n39056) );
  NAND2_X1 U2060 ( .A1(n8660), .A2(n12567), .ZN(n8659) );
  NOR2_X1 U2061 ( .A1(n63312), .A2(n60985), .ZN(n6195) );
  OAI22_X1 U2062 ( .A1(n40072), .A2(n1721), .B1(n59199), .B2(n40163), .ZN(
        n40244) );
  AOI21_X1 U2068 ( .A1(n3060), .A2(n3061), .B(n10201), .ZN(n3059) );
  NOR2_X1 U2069 ( .A1(n62719), .A2(n17076), .ZN(n63703) );
  NOR2_X1 U2070 ( .A1(n64580), .A2(n64581), .ZN(n64579) );
  NAND2_X1 U2081 ( .A1(n63349), .A2(n3612), .ZN(n231) );
  NOR2_X1 U2083 ( .A1(n40402), .A2(n4383), .ZN(n998) );
  AOI21_X1 U2086 ( .A1(n61952), .A2(n42433), .B(n17930), .ZN(n39926) );
  OAI22_X1 U2092 ( .A1(n41422), .A2(n41414), .B1(n64364), .B2(n38935), .ZN(
        n41418) );
  AND2_X1 U2095 ( .A1(n6791), .A2(n40645), .Z(n61707) );
  NAND2_X1 U2096 ( .A1(n39069), .A2(n39068), .ZN(n24766) );
  NOR2_X1 U2115 ( .A1(n4607), .A2(n65056), .ZN(n4468) );
  NAND3_X1 U2118 ( .A1(n23971), .A2(n39822), .A3(n39823), .ZN(n39824) );
  NOR2_X1 U2136 ( .A1(n42471), .A2(n63101), .ZN(n60349) );
  NAND2_X1 U2139 ( .A1(n17073), .A2(n41955), .ZN(n62719) );
  NOR2_X1 U2143 ( .A1(n41459), .A2(n63464), .ZN(n63463) );
  AND2_X1 U2163 ( .A1(n41825), .A2(n42428), .Z(n61952) );
  NAND2_X1 U2176 ( .A1(n18869), .A2(n64914), .ZN(n62969) );
  AOI21_X1 U2177 ( .A1(n57415), .A2(n40820), .B(n7995), .ZN(n63940) );
  AOI21_X1 U2183 ( .A1(n41205), .A2(n40731), .B(n62144), .ZN(n22894) );
  OAI22_X1 U2185 ( .A1(n62009), .A2(n62008), .B1(n1737), .B2(n40224), .ZN(
        n39916) );
  INV_X1 U2186 ( .I(n41190), .ZN(n22329) );
  AOI21_X1 U2187 ( .A1(n41809), .A2(n64359), .B(n6259), .ZN(n57515) );
  AOI22_X1 U2189 ( .A1(n62071), .A2(n40967), .B1(n39130), .B2(n40619), .ZN(
        n39063) );
  NAND2_X1 U2196 ( .A1(n19438), .A2(n39408), .ZN(n64675) );
  AOI21_X1 U2199 ( .A1(n6236), .A2(n39809), .B(n39808), .ZN(n20983) );
  OAI22_X1 U2200 ( .A1(n1723), .A2(n40379), .B1(n40380), .B2(n41447), .ZN(
        n19575) );
  OAI22_X1 U2201 ( .A1(n40203), .A2(n40199), .B1(n40108), .B2(n59427), .ZN(
        n62819) );
  NAND2_X1 U2207 ( .A1(n39028), .A2(n60567), .ZN(n41190) );
  OR2_X1 U2211 ( .A1(n41918), .A2(n21459), .Z(n23741) );
  INV_X1 U2219 ( .I(n62018), .ZN(n10479) );
  NAND2_X1 U2223 ( .A1(n39982), .A2(n10683), .ZN(n6236) );
  NAND2_X1 U2224 ( .A1(n61233), .A2(n20879), .ZN(n4259) );
  NAND3_X1 U2229 ( .A1(n41258), .A2(n40563), .A3(n42252), .ZN(n41262) );
  NOR2_X1 U2232 ( .A1(n40682), .A2(n25776), .ZN(n63676) );
  NOR2_X1 U2236 ( .A1(n40985), .A2(n40986), .ZN(n62232) );
  INV_X1 U2239 ( .I(n63119), .ZN(n63093) );
  NOR2_X1 U2242 ( .A1(n40986), .A2(n58364), .ZN(n64066) );
  OAI22_X1 U2243 ( .A1(n64672), .A2(n62123), .B1(n64390), .B2(n11704), .ZN(
        n62168) );
  NAND2_X1 U2259 ( .A1(n62191), .A2(n40734), .ZN(n62144) );
  NAND2_X1 U2260 ( .A1(n64475), .A2(n40857), .ZN(n63806) );
  OAI21_X1 U2263 ( .A1(n41948), .A2(n982), .B(n41947), .ZN(n41955) );
  NAND2_X1 U2273 ( .A1(n41882), .A2(n11895), .ZN(n63236) );
  NOR2_X1 U2274 ( .A1(n40523), .A2(n38607), .ZN(n62071) );
  NAND2_X1 U2276 ( .A1(n62107), .A2(n41376), .ZN(n40002) );
  NAND2_X1 U2279 ( .A1(n42265), .A2(n20287), .ZN(n64396) );
  NAND2_X1 U2282 ( .A1(n39862), .A2(n6852), .ZN(n41225) );
  OAI22_X1 U2283 ( .A1(n22607), .A2(n41278), .B1(n42294), .B2(n42293), .ZN(
        n65246) );
  OAI22_X1 U2288 ( .A1(n64672), .A2(n18483), .B1(n18338), .B2(n18441), .ZN(
        n62169) );
  OAI22_X1 U2289 ( .A1(n41472), .A2(n40747), .B1(n40414), .B2(n64308), .ZN(
        n39984) );
  NOR2_X1 U2292 ( .A1(n42453), .A2(n59674), .ZN(n42458) );
  INV_X1 U2293 ( .I(n41850), .ZN(n1734) );
  NAND2_X1 U2303 ( .A1(n8812), .A2(n6305), .ZN(n42228) );
  NAND2_X1 U2308 ( .A1(n41401), .A2(n11472), .ZN(n41230) );
  NAND2_X1 U2317 ( .A1(n18856), .A2(n21471), .ZN(n39048) );
  BUF_X2 U2318 ( .I(n59583), .Z(n62241) );
  CLKBUF_X2 U2324 ( .I(n14343), .Z(n64359) );
  OR2_X1 U2330 ( .A1(n14317), .A2(n21920), .Z(n61916) );
  INV_X1 U2331 ( .I(n11895), .ZN(n62785) );
  NAND2_X1 U2338 ( .A1(n42236), .A2(n63435), .ZN(n41803) );
  NAND2_X1 U2348 ( .A1(n1405), .A2(n63464), .ZN(n5673) );
  INV_X1 U2353 ( .I(n39021), .ZN(n40683) );
  NAND2_X1 U2356 ( .A1(n41199), .A2(n64793), .ZN(n62191) );
  NOR2_X1 U2361 ( .A1(n12895), .A2(n38939), .ZN(n39862) );
  NAND2_X1 U2367 ( .A1(n41397), .A2(n41400), .ZN(n63937) );
  NAND2_X1 U2375 ( .A1(n40304), .A2(n14016), .ZN(n62856) );
  NOR2_X1 U2376 ( .A1(n5362), .A2(n10542), .ZN(n37060) );
  INV_X1 U2377 ( .I(n40438), .ZN(n40437) );
  INV_X1 U2383 ( .I(n40472), .ZN(n63801) );
  INV_X1 U2395 ( .I(n41446), .ZN(n39846) );
  OR2_X1 U2396 ( .A1(n40200), .A2(n19148), .Z(n61712) );
  AND2_X1 U2399 ( .A1(n22289), .A2(n38273), .Z(n41944) );
  NAND2_X1 U2400 ( .A1(n60143), .A2(n42230), .ZN(n41942) );
  NAND2_X1 U2406 ( .A1(n41455), .A2(n23610), .ZN(n39021) );
  NAND2_X1 U2420 ( .A1(n1725), .A2(n976), .ZN(n42231) );
  INV_X1 U2421 ( .I(n21471), .ZN(n41237) );
  CLKBUF_X2 U2423 ( .I(n21529), .Z(n64895) );
  NOR2_X1 U2426 ( .A1(n14863), .A2(n38338), .ZN(n62018) );
  NOR2_X1 U2427 ( .A1(n40987), .A2(n23752), .ZN(n58264) );
  INV_X1 U2428 ( .I(n40068), .ZN(n20724) );
  INV_X1 U2438 ( .I(n40220), .ZN(n14558) );
  NOR2_X1 U2440 ( .A1(n42251), .A2(n42240), .ZN(n62204) );
  NOR2_X1 U2443 ( .A1(n64040), .A2(n39136), .ZN(n20397) );
  NAND2_X1 U2447 ( .A1(n40039), .A2(n42480), .ZN(n62023) );
  NOR3_X1 U2451 ( .A1(n42240), .A2(n286), .A3(n41258), .ZN(n24856) );
  INV_X1 U2454 ( .I(n39786), .ZN(n40854) );
  OR2_X1 U2456 ( .A1(n38600), .A2(n38516), .Z(n40956) );
  CLKBUF_X4 U2458 ( .I(n40063), .Z(n62291) );
  OR2_X1 U2459 ( .A1(n41444), .A2(n8260), .Z(n40379) );
  OR2_X1 U2464 ( .A1(n8260), .A2(n62416), .Z(n41428) );
  INV_X1 U2465 ( .I(n64655), .ZN(n59961) );
  NAND2_X1 U2466 ( .A1(n23875), .A2(n3685), .ZN(n3667) );
  INV_X2 U2483 ( .I(n62580), .ZN(n40196) );
  BUF_X2 U2484 ( .I(n38672), .Z(n64793) );
  BUF_X2 U2485 ( .I(n41210), .Z(n59203) );
  NAND2_X1 U2486 ( .A1(n41429), .A2(n39847), .ZN(n40702) );
  BUF_X2 U2491 ( .I(n42224), .Z(n22290) );
  CLKBUF_X2 U2492 ( .I(n40387), .Z(n63914) );
  CLKBUF_X2 U2496 ( .I(n4171), .Z(n64077) );
  CLKBUF_X2 U2497 ( .I(n42267), .Z(n9716) );
  CLKBUF_X2 U2500 ( .I(n41213), .Z(n10173) );
  NAND2_X1 U2501 ( .A1(n39987), .A2(n40755), .ZN(n40750) );
  NOR2_X1 U2508 ( .A1(n40272), .A2(n25229), .ZN(n16970) );
  NAND2_X1 U2509 ( .A1(n40571), .A2(n59601), .ZN(n63203) );
  NAND2_X1 U2511 ( .A1(n39987), .A2(n40749), .ZN(n40754) );
  BUF_X2 U2521 ( .I(n1409), .Z(n1512) );
  INV_X1 U2528 ( .I(n1226), .ZN(n64085) );
  INV_X1 U2531 ( .I(n37059), .ZN(n10954) );
  CLKBUF_X2 U2538 ( .I(n41132), .Z(n60091) );
  INV_X2 U2542 ( .I(n64172), .ZN(n971) );
  BUF_X2 U2554 ( .I(n23489), .Z(n1402) );
  BUF_X2 U2562 ( .I(n40193), .Z(n59427) );
  INV_X2 U2566 ( .I(n59601), .ZN(n64183) );
  INV_X1 U2571 ( .I(n40928), .ZN(n12082) );
  INV_X1 U2573 ( .I(n62105), .ZN(n16511) );
  INV_X1 U2577 ( .I(n23277), .ZN(n63426) );
  BUF_X2 U2579 ( .I(n39566), .Z(n15711) );
  INV_X1 U2586 ( .I(n63008), .ZN(n19145) );
  BUF_X2 U2593 ( .I(n14969), .Z(n63768) );
  INV_X1 U2599 ( .I(n11005), .ZN(n3172) );
  INV_X1 U2600 ( .I(n7857), .ZN(n13809) );
  NOR2_X1 U2608 ( .A1(n5108), .A2(n5107), .ZN(n63011) );
  AND2_X1 U2610 ( .A1(n38367), .A2(n61112), .Z(n61851) );
  INV_X1 U2622 ( .I(n39737), .ZN(n60616) );
  OAI21_X1 U2636 ( .A1(n62733), .A2(n61801), .B(n32148), .ZN(n32157) );
  AOI22_X1 U2653 ( .A1(n62471), .A2(n36729), .B1(n59809), .B2(n36730), .ZN(
        n25915) );
  NAND3_X1 U2656 ( .A1(n3011), .A2(n62939), .A3(n3010), .ZN(n61998) );
  NOR2_X1 U2658 ( .A1(n8531), .A2(n8532), .ZN(n57957) );
  AOI22_X1 U2663 ( .A1(n63161), .A2(n36086), .B1(n36088), .B2(n36087), .ZN(
        n36089) );
  NOR2_X1 U2664 ( .A1(n4268), .A2(n63381), .ZN(n4269) );
  NAND3_X1 U2674 ( .A1(n32145), .A2(n58561), .A3(n32144), .ZN(n62733) );
  INV_X1 U2676 ( .I(n9375), .ZN(n63046) );
  NAND2_X1 U2677 ( .A1(n64876), .A2(n36482), .ZN(n3313) );
  OAI21_X1 U2684 ( .A1(n18206), .A2(n18207), .B(n38912), .ZN(n20158) );
  OAI22_X1 U2685 ( .A1(n35573), .A2(n35574), .B1(n35572), .B2(n36019), .ZN(
        n65259) );
  NAND2_X1 U2686 ( .A1(n36729), .A2(n58743), .ZN(n17947) );
  NAND2_X1 U2702 ( .A1(n37313), .A2(n37314), .ZN(n63115) );
  NOR2_X1 U2705 ( .A1(n64476), .A2(n21695), .ZN(n21293) );
  NAND2_X1 U2708 ( .A1(n35128), .A2(n63083), .ZN(n58615) );
  NOR2_X1 U2709 ( .A1(n64619), .A2(n63348), .ZN(n5460) );
  NAND3_X1 U2716 ( .A1(n63399), .A2(n6612), .A3(n63398), .ZN(n8531) );
  NAND4_X1 U2724 ( .A1(n36984), .A2(n36982), .A3(n36983), .A4(n36981), .ZN(
        n64005) );
  OAI22_X1 U2735 ( .A1(n36468), .A2(n36467), .B1(n36466), .B2(n7933), .ZN(
        n64876) );
  NAND3_X1 U2736 ( .A1(n63595), .A2(n37086), .A3(n11754), .ZN(n62690) );
  AOI21_X1 U2737 ( .A1(n36084), .A2(n37125), .B(n36083), .ZN(n63161) );
  NAND2_X1 U2742 ( .A1(n19252), .A2(n35080), .ZN(n63762) );
  OR2_X1 U2753 ( .A1(n7656), .A2(n36442), .Z(n7655) );
  NAND2_X1 U2758 ( .A1(n17168), .A2(n21329), .ZN(n35574) );
  NAND2_X1 U2764 ( .A1(n63990), .A2(n5073), .ZN(n59277) );
  AOI21_X1 U2765 ( .A1(n17664), .A2(n17665), .B(n62162), .ZN(n36017) );
  NOR2_X1 U2768 ( .A1(n6632), .A2(n36779), .ZN(n62704) );
  NOR2_X1 U2769 ( .A1(n11143), .A2(n36583), .ZN(n62575) );
  NOR3_X1 U2770 ( .A1(n26194), .A2(n64103), .A3(n36490), .ZN(n64114) );
  NOR3_X1 U2781 ( .A1(n61784), .A2(n35576), .A3(n60891), .ZN(n17166) );
  NOR2_X1 U2782 ( .A1(n63900), .A2(n63899), .ZN(n4450) );
  NAND3_X1 U2786 ( .A1(n57848), .A2(n8816), .A3(n61631), .ZN(n63511) );
  NAND3_X1 U2791 ( .A1(n36866), .A2(n59924), .A3(n8808), .ZN(n8890) );
  NAND2_X1 U2795 ( .A1(n35996), .A2(n35997), .ZN(n35999) );
  NAND2_X1 U2823 ( .A1(n37409), .A2(n1771), .ZN(n22463) );
  AOI21_X1 U2826 ( .A1(n36312), .A2(n36313), .B(n64684), .ZN(n23320) );
  NAND2_X1 U2832 ( .A1(n62592), .A2(n64093), .ZN(n440) );
  NAND3_X1 U2833 ( .A1(n38544), .A2(n6630), .A3(n37477), .ZN(n6629) );
  NAND2_X1 U2834 ( .A1(n13459), .A2(n6138), .ZN(n63381) );
  OAI21_X1 U2840 ( .A1(n33782), .A2(n3057), .B(n33781), .ZN(n33784) );
  NAND2_X1 U2844 ( .A1(n34877), .A2(n7802), .ZN(n62333) );
  NAND2_X1 U2849 ( .A1(n60770), .A2(n60771), .ZN(n62984) );
  NAND2_X1 U2855 ( .A1(n17444), .A2(n24660), .ZN(n63644) );
  NOR2_X1 U2862 ( .A1(n35996), .A2(n31303), .ZN(n62782) );
  INV_X1 U2867 ( .I(n36292), .ZN(n63820) );
  NOR2_X1 U2875 ( .A1(n36963), .A2(n1786), .ZN(n18811) );
  NAND2_X1 U2879 ( .A1(n63049), .A2(n57988), .ZN(n62649) );
  NOR2_X1 U2880 ( .A1(n20007), .A2(n63395), .ZN(n37247) );
  OAI21_X1 U2883 ( .A1(n37083), .A2(n23651), .B(n37096), .ZN(n63595) );
  NOR2_X1 U2885 ( .A1(n62246), .A2(n62245), .ZN(n57434) );
  AOI22_X1 U2886 ( .A1(n37449), .A2(n37448), .B1(n37447), .B2(n37446), .ZN(
        n63207) );
  AOI21_X1 U2887 ( .A1(n58285), .A2(n58933), .B(n36159), .ZN(n14893) );
  NAND2_X1 U2888 ( .A1(n35089), .A2(n37322), .ZN(n63665) );
  NAND2_X1 U2889 ( .A1(n61856), .A2(n36776), .ZN(n62500) );
  AOI21_X1 U2893 ( .A1(n35054), .A2(n35444), .B(n64011), .ZN(n13533) );
  NAND2_X1 U2896 ( .A1(n25225), .A2(n22559), .ZN(n63398) );
  NAND3_X1 U2898 ( .A1(n64798), .A2(n2220), .A3(n4636), .ZN(n11312) );
  NOR2_X1 U2900 ( .A1(n37112), .A2(n6831), .ZN(n63899) );
  OAI21_X1 U2905 ( .A1(n34817), .A2(n18427), .B(n22595), .ZN(n19689) );
  AOI21_X1 U2906 ( .A1(n13769), .A2(n35971), .B(n61636), .ZN(n64476) );
  NAND2_X1 U2911 ( .A1(n63845), .A2(n36606), .ZN(n37965) );
  NAND3_X1 U2915 ( .A1(n19552), .A2(n17663), .A3(n8299), .ZN(n62162) );
  NOR2_X1 U2918 ( .A1(n23778), .A2(n36001), .ZN(n62783) );
  OAI22_X1 U2925 ( .A1(n64164), .A2(n37214), .B1(n37212), .B2(n37211), .ZN(n29) );
  NAND2_X1 U2935 ( .A1(n36154), .A2(n3218), .ZN(n3907) );
  NAND2_X1 U2937 ( .A1(n25584), .A2(n19231), .ZN(n34105) );
  INV_X1 U2941 ( .I(n17144), .ZN(n37422) );
  NOR2_X1 U2947 ( .A1(n35946), .A2(n34816), .ZN(n62654) );
  OAI21_X1 U2949 ( .A1(n36550), .A2(n36538), .B(n62151), .ZN(n36066) );
  NAND2_X1 U2963 ( .A1(n36945), .A2(n36944), .ZN(n36949) );
  NAND2_X1 U2964 ( .A1(n3620), .A2(n17096), .ZN(n24427) );
  NOR2_X1 U2966 ( .A1(n36109), .A2(n9984), .ZN(n36112) );
  NOR2_X1 U2982 ( .A1(n35871), .A2(n4834), .ZN(n64619) );
  NAND2_X1 U2988 ( .A1(n61747), .A2(n7092), .ZN(n64905) );
  NOR2_X1 U2989 ( .A1(n1782), .A2(n36494), .ZN(n9513) );
  NAND3_X1 U3000 ( .A1(n14093), .A2(n8356), .A3(n1785), .ZN(n36576) );
  INV_X1 U3004 ( .I(n20501), .ZN(n63395) );
  CLKBUF_X2 U3016 ( .I(n34914), .Z(n64101) );
  OR2_X1 U3017 ( .A1(n36971), .A2(n35852), .Z(n61937) );
  NAND2_X1 U3032 ( .A1(n10086), .A2(n7103), .ZN(n36535) );
  INV_X1 U3039 ( .I(n16426), .ZN(n19666) );
  NAND2_X1 U3043 ( .A1(n36313), .A2(n3864), .ZN(n62245) );
  BUF_X2 U3048 ( .I(n36846), .Z(n62942) );
  NOR2_X1 U3051 ( .A1(n20712), .A2(n35979), .ZN(n18207) );
  NAND2_X1 U3052 ( .A1(n37428), .A2(n23801), .ZN(n37419) );
  NAND2_X1 U3055 ( .A1(n2002), .A2(n36775), .ZN(n34854) );
  NAND3_X1 U3059 ( .A1(n35068), .A2(n58769), .A3(n1417), .ZN(n36751) );
  NAND3_X1 U3061 ( .A1(n37395), .A2(n37394), .A3(n16910), .ZN(n22853) );
  NOR3_X1 U3062 ( .A1(n36063), .A2(n36062), .A3(n36898), .ZN(n62151) );
  NOR2_X1 U3075 ( .A1(n35991), .A2(n35997), .ZN(n63845) );
  NOR2_X1 U3086 ( .A1(n36010), .A2(n36841), .ZN(n63771) );
  NOR2_X1 U3087 ( .A1(n36728), .A2(n21489), .ZN(n63910) );
  NOR2_X1 U3094 ( .A1(n35470), .A2(n15720), .ZN(n64524) );
  OAI21_X1 U3095 ( .A1(n37352), .A2(n6831), .B(n22659), .ZN(n64798) );
  NAND3_X1 U3104 ( .A1(n36841), .A2(n23146), .A3(n61747), .ZN(n63402) );
  NOR2_X1 U3109 ( .A1(n16054), .A2(n57830), .ZN(n25585) );
  NOR3_X1 U3110 ( .A1(n35608), .A2(n36719), .A3(n36724), .ZN(n16059) );
  NOR3_X1 U3111 ( .A1(n23626), .A2(n34819), .A3(n36041), .ZN(n57592) );
  NAND2_X1 U3112 ( .A1(n36041), .A2(n35570), .ZN(n21328) );
  INV_X2 U3114 ( .I(n61747), .ZN(n63697) );
  AND2_X1 U3121 ( .A1(n35723), .A2(n61935), .Z(n37204) );
  NOR2_X1 U3123 ( .A1(n36304), .A2(n57211), .ZN(n36800) );
  CLKBUF_X2 U3124 ( .I(n1339), .Z(n64181) );
  CLKBUF_X2 U3133 ( .I(n22936), .Z(n4745) );
  NAND2_X1 U3140 ( .A1(n25964), .A2(n21921), .ZN(n37068) );
  NAND2_X1 U3143 ( .A1(n5900), .A2(n35447), .ZN(n36275) );
  NOR2_X1 U3154 ( .A1(n17144), .A2(n8177), .ZN(n16445) );
  NOR2_X1 U3158 ( .A1(n36224), .A2(n35591), .ZN(n35595) );
  NOR2_X1 U3159 ( .A1(n59988), .A2(n17892), .ZN(n11414) );
  NOR2_X1 U3167 ( .A1(n37035), .A2(n58876), .ZN(n35491) );
  NAND2_X1 U3169 ( .A1(n10717), .A2(n36775), .ZN(n34369) );
  NAND2_X1 U3171 ( .A1(n35551), .A2(n65178), .ZN(n258) );
  NOR3_X1 U3175 ( .A1(n36163), .A2(n22632), .A3(n37374), .ZN(n24366) );
  AOI21_X1 U3181 ( .A1(n34921), .A2(n4151), .B(n24198), .ZN(n7682) );
  INV_X4 U3192 ( .I(n22461), .ZN(n34816) );
  NAND2_X1 U3198 ( .A1(n36898), .A2(n36394), .ZN(n36389) );
  CLKBUF_X2 U3206 ( .I(n13126), .Z(n23801) );
  NAND2_X1 U3211 ( .A1(n35965), .A2(n35962), .ZN(n8608) );
  INV_X1 U3214 ( .I(n37400), .ZN(n58285) );
  NAND3_X1 U3224 ( .A1(n57209), .A2(n7729), .A3(n1527), .ZN(n7230) );
  INV_X1 U3225 ( .I(n25677), .ZN(n36075) );
  BUF_X2 U3229 ( .I(n37374), .Z(n2594) );
  BUF_X2 U3236 ( .I(n36838), .Z(n23146) );
  NOR2_X1 U3241 ( .A1(n34926), .A2(n24609), .ZN(n34921) );
  NAND2_X1 U3243 ( .A1(n35974), .A2(n6606), .ZN(n35142) );
  BUF_X2 U3244 ( .I(n20908), .Z(n64609) );
  INV_X1 U3249 ( .I(n36529), .ZN(n20531) );
  NAND2_X1 U3257 ( .A1(n60437), .A2(n1527), .ZN(n36964) );
  INV_X2 U3268 ( .I(n35140), .ZN(n35974) );
  BUF_X2 U3270 ( .I(n34078), .Z(n14189) );
  INV_X2 U3275 ( .I(n36953), .ZN(n35431) );
  BUF_X2 U3280 ( .I(n36691), .Z(n62720) );
  BUF_X4 U3309 ( .I(n12521), .Z(n6984) );
  NAND2_X1 U3317 ( .A1(n12239), .A2(n33495), .ZN(n63984) );
  AOI21_X1 U3324 ( .A1(n24544), .A2(n34522), .B(n20520), .ZN(n14194) );
  AOI21_X1 U3334 ( .A1(n63077), .A2(n5996), .B(n35704), .ZN(n5995) );
  NAND2_X1 U3350 ( .A1(n31541), .A2(n31534), .ZN(n63815) );
  NAND2_X1 U3359 ( .A1(n64112), .A2(n32938), .ZN(n64468) );
  NOR2_X1 U3361 ( .A1(n64381), .A2(n33429), .ZN(n16338) );
  NOR2_X1 U3375 ( .A1(n21322), .A2(n64407), .ZN(n32793) );
  AOI21_X1 U3405 ( .A1(n33460), .A2(n23761), .B(n64371), .ZN(n7293) );
  AOI21_X1 U3417 ( .A1(n17427), .A2(n64304), .B(n64314), .ZN(n31909) );
  AOI21_X1 U3421 ( .A1(n32832), .A2(n61896), .B(n63488), .ZN(n32840) );
  INV_X1 U3426 ( .I(n34656), .ZN(n13251) );
  AOI21_X1 U3441 ( .A1(n33531), .A2(n57364), .B(n16096), .ZN(n15620) );
  AOI21_X1 U3450 ( .A1(n35670), .A2(n58684), .B(n24286), .ZN(n62140) );
  NOR2_X1 U3451 ( .A1(n62692), .A2(n58544), .ZN(n63387) );
  OAI21_X1 U3458 ( .A1(n34513), .A2(n2476), .B(n24874), .ZN(n5610) );
  OAI21_X1 U3463 ( .A1(n17502), .A2(n64356), .B(n34517), .ZN(n9461) );
  NAND2_X1 U3464 ( .A1(n33997), .A2(n61841), .ZN(n7730) );
  OR2_X1 U3471 ( .A1(n19924), .A2(n17759), .Z(n61899) );
  OAI21_X1 U3474 ( .A1(n61701), .A2(n63669), .B(n20835), .ZN(n25350) );
  NOR2_X1 U3481 ( .A1(n59237), .A2(n32296), .ZN(n64016) );
  NAND3_X1 U3486 ( .A1(n8431), .A2(n34962), .A3(n476), .ZN(n34540) );
  NAND3_X1 U3495 ( .A1(n35635), .A2(n8365), .A3(n57546), .ZN(n63893) );
  NOR4_X1 U3500 ( .A1(n61982), .A2(n61818), .A3(n4701), .A4(n62078), .ZN(n414)
         );
  AND2_X1 U3501 ( .A1(n9085), .A2(n6620), .Z(n61842) );
  NAND3_X1 U3507 ( .A1(n33531), .A2(n7043), .A3(n7042), .ZN(n33535) );
  NAND2_X1 U3508 ( .A1(n19781), .A2(n10852), .ZN(n63446) );
  NOR2_X1 U3509 ( .A1(n62566), .A2(n63062), .ZN(n62692) );
  INV_X1 U3510 ( .I(n35250), .ZN(n58187) );
  NOR2_X1 U3513 ( .A1(n62158), .A2(n2386), .ZN(n2384) );
  NOR2_X1 U3514 ( .A1(n891), .A2(n33214), .ZN(n63862) );
  INV_X1 U3516 ( .I(n3432), .ZN(n64112) );
  AOI22_X1 U3522 ( .A1(n33015), .A2(n33014), .B1(n33013), .B2(n33599), .ZN(
        n36545) );
  OAI21_X1 U3523 ( .A1(n62440), .A2(n33341), .B(n33563), .ZN(n33092) );
  NAND3_X1 U3524 ( .A1(n62016), .A2(n33691), .A3(n33089), .ZN(n62287) );
  NOR2_X1 U3537 ( .A1(n57200), .A2(n12506), .ZN(n62351) );
  NOR2_X1 U3538 ( .A1(n34045), .A2(n34042), .ZN(n21113) );
  NOR2_X1 U3540 ( .A1(n18440), .A2(n32944), .ZN(n64782) );
  AOI21_X1 U3551 ( .A1(n34625), .A2(n12859), .B(n64677), .ZN(n16257) );
  NAND2_X1 U3558 ( .A1(n33997), .A2(n1535), .ZN(n62947) );
  NOR3_X1 U3560 ( .A1(n34034), .A2(n34033), .A3(n34602), .ZN(n63494) );
  NOR2_X1 U3573 ( .A1(n33385), .A2(n33384), .ZN(n33387) );
  INV_X1 U3577 ( .I(n19095), .ZN(n11038) );
  NOR2_X1 U3581 ( .A1(n35673), .A2(n62322), .ZN(n62352) );
  NAND3_X1 U3585 ( .A1(n35826), .A2(n34707), .A3(n35821), .ZN(n63048) );
  AOI21_X1 U3594 ( .A1(n24295), .A2(n34017), .B(n34632), .ZN(n20992) );
  NOR2_X1 U3596 ( .A1(n33567), .A2(n33566), .ZN(n61140) );
  OAI21_X1 U3597 ( .A1(n22118), .A2(n11281), .B(n18451), .ZN(n64300) );
  NAND2_X1 U3602 ( .A1(n33965), .A2(n34090), .ZN(n63754) );
  NAND2_X1 U3604 ( .A1(n60819), .A2(n904), .ZN(n63078) );
  NAND3_X1 U3610 ( .A1(n35715), .A2(n59824), .A3(n35841), .ZN(n34408) );
  INV_X1 U3611 ( .I(n33462), .ZN(n64371) );
  NAND3_X1 U3612 ( .A1(n61312), .A2(n14792), .A3(n34023), .ZN(n64381) );
  AOI22_X1 U3613 ( .A1(n34660), .A2(n14107), .B1(n1535), .B2(n34661), .ZN(
        n34662) );
  NAND4_X1 U3614 ( .A1(n35642), .A2(n35644), .A3(n35643), .A4(n22909), .ZN(
        n18944) );
  AND2_X1 U3616 ( .A1(n33960), .A2(n6721), .Z(n34619) );
  AND2_X1 U3619 ( .A1(n11992), .A2(n6721), .Z(n22118) );
  NAND2_X1 U3621 ( .A1(n7731), .A2(n34001), .ZN(n33997) );
  OAI21_X1 U3634 ( .A1(n34983), .A2(n10091), .B(n63443), .ZN(n15254) );
  INV_X2 U3638 ( .I(n7359), .ZN(n63064) );
  NOR2_X1 U3639 ( .A1(n35847), .A2(n34395), .ZN(n64473) );
  NAND2_X1 U3640 ( .A1(n35273), .A2(n11182), .ZN(n63132) );
  AOI21_X1 U3643 ( .A1(n31356), .A2(n34679), .B(n63861), .ZN(n64329) );
  INV_X1 U3644 ( .I(n35211), .ZN(n62566) );
  NAND2_X1 U3645 ( .A1(n59769), .A2(n32795), .ZN(n62078) );
  NAND3_X1 U3647 ( .A1(n17538), .A2(n64812), .A3(n20989), .ZN(n34344) );
  NAND2_X1 U3650 ( .A1(n35210), .A2(n57732), .ZN(n63062) );
  AOI22_X1 U3657 ( .A1(n6360), .A2(n1807), .B1(n11992), .B2(n64283), .ZN(
        n11281) );
  NOR2_X1 U3658 ( .A1(n34587), .A2(n20607), .ZN(n63669) );
  OAI22_X1 U3660 ( .A1(n19790), .A2(n35674), .B1(n57200), .B2(n7321), .ZN(
        n18379) );
  NOR2_X1 U3663 ( .A1(n34733), .A2(n34748), .ZN(n34739) );
  AOI22_X1 U3671 ( .A1(n35740), .A2(n60819), .B1(n61702), .B2(n35705), .ZN(
        n35285) );
  NOR2_X1 U3672 ( .A1(n23746), .A2(n34613), .ZN(n33978) );
  NAND2_X1 U3673 ( .A1(n24286), .A2(n17401), .ZN(n25563) );
  NAND2_X1 U3674 ( .A1(n33597), .A2(n35679), .ZN(n35683) );
  NAND2_X1 U3675 ( .A1(n18488), .A2(n34221), .ZN(n34293) );
  NAND3_X1 U3678 ( .A1(n5386), .A2(n11064), .A3(n18390), .ZN(n19805) );
  NOR2_X1 U3681 ( .A1(n33738), .A2(n34248), .ZN(n34349) );
  NAND2_X1 U3683 ( .A1(n21938), .A2(n35743), .ZN(n35730) );
  NAND2_X1 U3684 ( .A1(n64883), .A2(n20356), .ZN(n35839) );
  NAND2_X1 U3690 ( .A1(n1804), .A2(n23366), .ZN(n63843) );
  NAND3_X1 U3691 ( .A1(n32946), .A2(n60738), .A3(n65194), .ZN(n32429) );
  NAND2_X1 U3692 ( .A1(n13770), .A2(n60669), .ZN(n34441) );
  NOR2_X1 U3693 ( .A1(n35333), .A2(n33925), .ZN(n63254) );
  OAI21_X1 U3698 ( .A1(n34228), .A2(n17141), .B(n35273), .ZN(n63557) );
  NAND2_X1 U3699 ( .A1(n60413), .A2(n32951), .ZN(n63928) );
  INV_X1 U3703 ( .I(n34163), .ZN(n63579) );
  NAND2_X1 U3705 ( .A1(n35701), .A2(n63072), .ZN(n63827) );
  INV_X1 U3711 ( .I(n63581), .ZN(n32933) );
  NOR2_X1 U3712 ( .A1(n34957), .A2(n57166), .ZN(n12170) );
  INV_X1 U3718 ( .I(n65052), .ZN(n32897) );
  INV_X1 U3720 ( .I(n34784), .ZN(n34779) );
  INV_X1 U3727 ( .I(n34167), .ZN(n1795) );
  NAND2_X1 U3728 ( .A1(n22419), .A2(n13818), .ZN(n34969) );
  INV_X1 U3731 ( .I(n23743), .ZN(n35303) );
  AND2_X1 U3736 ( .A1(n34189), .A2(n2346), .Z(n61701) );
  BUF_X2 U3739 ( .I(n26163), .Z(n4075) );
  NOR2_X1 U3741 ( .A1(n34350), .A2(n23914), .ZN(n34721) );
  INV_X2 U3742 ( .I(n61522), .ZN(n33570) );
  NAND2_X1 U3745 ( .A1(n5409), .A2(n34658), .ZN(n34163) );
  CLKBUF_X2 U3750 ( .I(n59398), .Z(n65232) );
  NAND2_X1 U3751 ( .A1(n34972), .A2(n25404), .ZN(n33725) );
  INV_X1 U3753 ( .I(n20785), .ZN(n64706) );
  INV_X1 U3754 ( .I(n34353), .ZN(n63250) );
  NAND2_X1 U3757 ( .A1(n34588), .A2(n57165), .ZN(n57669) );
  NOR2_X1 U3759 ( .A1(n2064), .A2(n34727), .ZN(n6579) );
  OAI22_X1 U3761 ( .A1(n21938), .A2(n35731), .B1(n61702), .B2(n15148), .ZN(
        n59874) );
  INV_X1 U3764 ( .I(n35027), .ZN(n64708) );
  INV_X1 U3767 ( .I(n34358), .ZN(n63249) );
  INV_X1 U3772 ( .I(n24153), .ZN(n34189) );
  BUF_X2 U3783 ( .I(n34588), .Z(n23223) );
  BUF_X2 U3788 ( .I(n34961), .Z(n60579) );
  BUF_X2 U3790 ( .I(n32748), .Z(n33338) );
  NOR2_X1 U3791 ( .A1(n15184), .A2(n23914), .ZN(n60604) );
  BUF_X2 U3792 ( .I(n23470), .Z(n21388) );
  BUF_X2 U3797 ( .I(n24181), .Z(n10401) );
  BUF_X2 U3802 ( .I(n15809), .Z(n20835) );
  CLKBUF_X2 U3805 ( .I(n23410), .Z(n19512) );
  BUF_X2 U3807 ( .I(n32461), .Z(n65256) );
  CLKBUF_X4 U3813 ( .I(n13583), .Z(n63375) );
  BUF_X2 U3818 ( .I(n15588), .Z(n61748) );
  CLKBUF_X2 U3821 ( .I(n34209), .Z(n65194) );
  CLKBUF_X2 U3824 ( .I(n32425), .Z(n493) );
  BUF_X2 U3828 ( .I(n30944), .Z(n34961) );
  INV_X2 U3831 ( .I(n32846), .ZN(n61197) );
  INV_X1 U3837 ( .I(n1343), .ZN(n57342) );
  INV_X1 U3838 ( .I(n59936), .ZN(n7007) );
  INV_X1 U3841 ( .I(n63428), .ZN(n10232) );
  CLKBUF_X2 U3843 ( .I(n31456), .Z(n64360) );
  INV_X1 U3847 ( .I(n32369), .ZN(n62762) );
  CLKBUF_X2 U3849 ( .I(n32368), .Z(n496) );
  INV_X1 U3850 ( .I(n32321), .ZN(n32003) );
  INV_X1 U3853 ( .I(n16953), .ZN(n62548) );
  BUF_X2 U3854 ( .I(n30735), .Z(n32592) );
  INV_X1 U3855 ( .I(n33840), .ZN(n17035) );
  INV_X1 U3860 ( .I(n31322), .ZN(n32121) );
  CLKBUF_X2 U3861 ( .I(n32615), .Z(n33153) );
  INV_X1 U3862 ( .I(n16625), .ZN(n62147) );
  BUF_X2 U3869 ( .I(n15869), .Z(n61732) );
  INV_X1 U3875 ( .I(n25455), .ZN(n33248) );
  INV_X1 U3877 ( .I(n32001), .ZN(n1314) );
  INV_X2 U3878 ( .I(n2130), .ZN(n23152) );
  CLKBUF_X2 U3881 ( .I(n8074), .Z(n15844) );
  INV_X1 U3883 ( .I(n62354), .ZN(n823) );
  BUF_X2 U3885 ( .I(n24594), .Z(n10409) );
  AOI21_X1 U3890 ( .A1(n30129), .A2(n30128), .B(n64617), .ZN(n22353) );
  AOI21_X1 U3900 ( .A1(n27239), .A2(n63431), .B(n14668), .ZN(n14667) );
  AOI21_X1 U3902 ( .A1(n29252), .A2(n62414), .B(n61882), .ZN(n13083) );
  INV_X1 U3904 ( .I(n30833), .ZN(n61346) );
  NAND2_X1 U3909 ( .A1(n29928), .A2(n30534), .ZN(n29940) );
  NOR2_X1 U3910 ( .A1(n27903), .A2(n27904), .ZN(n20777) );
  AND2_X1 U3912 ( .A1(n25881), .A2(n29778), .Z(n61882) );
  OAI22_X1 U3913 ( .A1(n61912), .A2(n30751), .B1(n30310), .B2(n30309), .ZN(
        n30316) );
  NAND2_X1 U3919 ( .A1(n64907), .A2(n64906), .ZN(n10178) );
  NAND2_X1 U3923 ( .A1(n30234), .A2(n29212), .ZN(n29213) );
  OAI22_X1 U3925 ( .A1(n30127), .A2(n1551), .B1(n17084), .B2(n30126), .ZN(
        n64617) );
  OAI21_X1 U3930 ( .A1(n29832), .A2(n162), .B(n62793), .ZN(n10858) );
  OAI21_X1 U3942 ( .A1(n28117), .A2(n29844), .B(n29448), .ZN(n63431) );
  NOR2_X1 U3945 ( .A1(n30540), .A2(n58409), .ZN(n30435) );
  NAND2_X1 U3946 ( .A1(n30523), .A2(n22877), .ZN(n29768) );
  NOR2_X1 U3947 ( .A1(n19191), .A2(n19192), .ZN(n19190) );
  NAND2_X1 U3948 ( .A1(n7466), .A2(n63166), .ZN(n63165) );
  NAND2_X1 U3954 ( .A1(n31170), .A2(n64064), .ZN(n57589) );
  NAND2_X1 U3979 ( .A1(n61839), .A2(n63504), .ZN(n15665) );
  NAND3_X1 U3985 ( .A1(n9340), .A2(n28791), .A3(n28789), .ZN(n2667) );
  NAND2_X1 U3986 ( .A1(n62588), .A2(n62585), .ZN(n63362) );
  INV_X1 U3991 ( .I(n12632), .ZN(n65120) );
  NOR2_X1 U3995 ( .A1(n29740), .A2(n16979), .ZN(n63939) );
  NAND2_X1 U3996 ( .A1(n17792), .A2(n17791), .ZN(n63097) );
  AOI21_X1 U4006 ( .A1(n30804), .A2(n29929), .B(n30799), .ZN(n62793) );
  NOR3_X1 U4008 ( .A1(n30862), .A2(n57937), .A3(n24777), .ZN(n27904) );
  NAND2_X1 U4013 ( .A1(n29858), .A2(n29863), .ZN(n64917) );
  NAND3_X1 U4021 ( .A1(n29950), .A2(n27972), .A3(n63592), .ZN(n60451) );
  AND2_X1 U4027 ( .A1(n29516), .A2(n64565), .Z(n61825) );
  OAI22_X1 U4032 ( .A1(n61827), .A2(n18736), .B1(n29102), .B2(n28748), .ZN(
        n64699) );
  NAND3_X1 U4033 ( .A1(n29564), .A2(n28952), .A3(n14202), .ZN(n64907) );
  OAI21_X1 U4035 ( .A1(n30784), .A2(n29552), .B(n1319), .ZN(n29555) );
  OAI21_X1 U4037 ( .A1(n30194), .A2(n30193), .B(n2351), .ZN(n62968) );
  NOR2_X1 U4038 ( .A1(n29019), .A2(n64962), .ZN(n16082) );
  OAI21_X1 U4040 ( .A1(n23224), .A2(n29460), .B(n14399), .ZN(n20808) );
  AND2_X1 U4041 ( .A1(n30254), .A2(n2269), .Z(n61892) );
  NOR2_X1 U4043 ( .A1(n1351), .A2(n22877), .ZN(n27924) );
  OR2_X1 U4044 ( .A1(n18581), .A2(n59046), .Z(n61912) );
  INV_X1 U4046 ( .I(n30084), .ZN(n64962) );
  NOR2_X1 U4051 ( .A1(n30030), .A2(n27739), .ZN(n29876) );
  NOR2_X1 U4055 ( .A1(n29559), .A2(n29560), .ZN(n64911) );
  NAND2_X1 U4056 ( .A1(n21588), .A2(n6912), .ZN(n63646) );
  OR2_X1 U4060 ( .A1(n29242), .A2(n61187), .Z(n61839) );
  NOR2_X1 U4061 ( .A1(n30642), .A2(n30641), .ZN(n62953) );
  OAI21_X1 U4063 ( .A1(n30610), .A2(n61783), .B(n61897), .ZN(n15926) );
  NAND4_X1 U4066 ( .A1(n65032), .A2(n3761), .A3(n30747), .A4(n14217), .ZN(
        n59248) );
  NAND2_X1 U4068 ( .A1(n31081), .A2(n24504), .ZN(n63333) );
  OAI22_X1 U4070 ( .A1(n30522), .A2(n20315), .B1(n30524), .B2(n64057), .ZN(
        n64084) );
  NAND4_X1 U4074 ( .A1(n30654), .A2(n3901), .A3(n29949), .A4(n62285), .ZN(
        n28714) );
  NAND2_X1 U4090 ( .A1(n31218), .A2(n30754), .ZN(n64236) );
  AOI22_X1 U4092 ( .A1(n13412), .A2(n61777), .B1(n31174), .B2(n1431), .ZN(
        n24155) );
  NAND3_X1 U4109 ( .A1(n29516), .A2(n17413), .A3(n29512), .ZN(n29093) );
  NOR2_X1 U4111 ( .A1(n27743), .A2(n28989), .ZN(n29882) );
  INV_X1 U4114 ( .I(n24556), .ZN(n63256) );
  NOR2_X1 U4115 ( .A1(n23056), .A2(n16279), .ZN(n30135) );
  NOR2_X1 U4123 ( .A1(n28696), .A2(n29993), .ZN(n30000) );
  BUF_X2 U4126 ( .I(n30602), .Z(n61737) );
  AOI21_X1 U4134 ( .A1(n57733), .A2(n63259), .B(n63237), .ZN(n64538) );
  OR2_X1 U4138 ( .A1(n40), .A2(n22504), .Z(n61783) );
  OR2_X1 U4140 ( .A1(n29077), .A2(n30348), .Z(n61752) );
  INV_X1 U4142 ( .I(n9392), .ZN(n62103) );
  INV_X1 U4149 ( .I(n18581), .ZN(n64238) );
  NOR2_X1 U4150 ( .A1(n24949), .A2(n29502), .ZN(n65138) );
  NAND2_X1 U4153 ( .A1(n62670), .A2(n62669), .ZN(n30053) );
  NAND2_X1 U4157 ( .A1(n29942), .A2(n30333), .ZN(n6912) );
  NAND3_X1 U4159 ( .A1(n327), .A2(n31155), .A3(n31156), .ZN(n31160) );
  NOR3_X1 U4160 ( .A1(n8522), .A2(n11092), .A3(n30333), .ZN(n28712) );
  NAND2_X1 U4165 ( .A1(n14276), .A2(n10102), .ZN(n30574) );
  INV_X1 U4166 ( .I(n5768), .ZN(n63159) );
  OR2_X1 U4172 ( .A1(n13174), .A2(n24811), .Z(n61753) );
  INV_X2 U4176 ( .I(n7405), .ZN(n29460) );
  NAND2_X1 U4177 ( .A1(n1253), .A2(n30538), .ZN(n29981) );
  NOR2_X1 U4180 ( .A1(n16382), .A2(n22556), .ZN(n23237) );
  NOR2_X1 U4181 ( .A1(n8522), .A2(n23901), .ZN(n30640) );
  CLKBUF_X2 U4188 ( .I(n21532), .Z(n63691) );
  NAND2_X1 U4191 ( .A1(n5768), .A2(n29010), .ZN(n31145) );
  INV_X1 U4196 ( .I(n30953), .ZN(n64940) );
  INV_X1 U4197 ( .I(n31141), .ZN(n63158) );
  BUF_X2 U4200 ( .I(n14174), .Z(n9426) );
  CLKBUF_X2 U4203 ( .I(n30292), .Z(n23734) );
  BUF_X2 U4212 ( .I(n29834), .Z(n11830) );
  BUF_X2 U4214 ( .I(n19059), .Z(n13144) );
  CLKBUF_X2 U4221 ( .I(n1871), .Z(n58486) );
  INV_X1 U4222 ( .I(n62437), .ZN(n30264) );
  BUF_X2 U4226 ( .I(n27591), .Z(n60293) );
  BUF_X2 U4227 ( .I(n58606), .Z(n61733) );
  INV_X1 U4228 ( .I(n64950), .ZN(n22893) );
  BUF_X2 U4233 ( .I(n30722), .Z(n23772) );
  NAND2_X1 U4239 ( .A1(n12347), .A2(n18938), .ZN(n18936) );
  NAND2_X1 U4247 ( .A1(n28236), .A2(n64622), .ZN(n64621) );
  NAND2_X1 U4255 ( .A1(n63053), .A2(n2907), .ZN(n13806) );
  OAI21_X1 U4266 ( .A1(n8822), .A2(n8824), .B(n28514), .ZN(n8893) );
  NOR3_X1 U4268 ( .A1(n64959), .A2(n8338), .A3(n28005), .ZN(n9014) );
  NAND3_X1 U4270 ( .A1(n63299), .A2(n26288), .A3(n26287), .ZN(n63298) );
  NOR2_X1 U4271 ( .A1(n62271), .A2(n62270), .ZN(n15992) );
  INV_X1 U4275 ( .I(n29689), .ZN(n64929) );
  OAI21_X1 U4276 ( .A1(n28380), .A2(n469), .B(n64942), .ZN(n20898) );
  OAI21_X1 U4286 ( .A1(n28441), .A2(n28440), .B(n64572), .ZN(n28442) );
  AOI22_X1 U4288 ( .A1(n26343), .A2(n2789), .B1(n28406), .B2(n1893), .ZN(
        n26515) );
  INV_X1 U4289 ( .I(n29158), .ZN(n27975) );
  OAI21_X1 U4295 ( .A1(n62532), .A2(n11513), .B(n29124), .ZN(n62156) );
  AOI21_X1 U4296 ( .A1(n28550), .A2(n28551), .B(n29192), .ZN(n28555) );
  NAND3_X1 U4297 ( .A1(n63714), .A2(n17046), .A3(n63713), .ZN(n13562) );
  INV_X1 U4301 ( .I(n26469), .ZN(n27434) );
  AND2_X1 U4304 ( .A1(n64145), .A2(n13483), .Z(n13482) );
  NAND2_X1 U4305 ( .A1(n469), .A2(n27560), .ZN(n26551) );
  NOR2_X1 U4306 ( .A1(n5117), .A2(n27532), .ZN(n26678) );
  NOR2_X1 U4308 ( .A1(n8389), .A2(n28886), .ZN(n64810) );
  BUF_X2 U4311 ( .I(n15414), .Z(n17619) );
  BUF_X1 U4312 ( .I(n65111), .Z(n63532) );
  INV_X1 U4314 ( .I(n27390), .ZN(n62099) );
  OAI21_X1 U4315 ( .A1(n26330), .A2(n26539), .B(n26606), .ZN(n26319) );
  NAND3_X1 U4316 ( .A1(n27121), .A2(n26613), .A3(n10946), .ZN(n14135) );
  NOR2_X1 U4318 ( .A1(n5206), .A2(n26969), .ZN(n26689) );
  INV_X2 U4319 ( .I(n14947), .ZN(n63714) );
  INV_X1 U4324 ( .I(n27559), .ZN(n28376) );
  INV_X2 U4325 ( .I(n2971), .ZN(n27980) );
  CLKBUF_X2 U4328 ( .I(n28616), .Z(n63330) );
  CLKBUF_X2 U4331 ( .I(n28495), .Z(n10125) );
  AND2_X1 U4332 ( .A1(n64445), .A2(n11850), .Z(n61921) );
  NAND2_X1 U4333 ( .A1(n20473), .A2(n22214), .ZN(n18826) );
  BUF_X2 U4335 ( .I(n27823), .Z(n20743) );
  INV_X1 U4337 ( .I(n15092), .ZN(n62155) );
  OAI22_X2 U4339 ( .A1(n56968), .A2(n9035), .B1(n56967), .B2(n56966), .ZN(
        n65163) );
  BUF_X2 U4341 ( .I(n34233), .Z(n64458) );
  AOI21_X2 U4344 ( .A1(n54133), .A2(n54132), .B(n62651), .ZN(n54141) );
  NOR2_X2 U4348 ( .A1(n20374), .A2(n18704), .ZN(n20396) );
  NAND2_X2 U4350 ( .A1(n47623), .A2(n45991), .ZN(n47617) );
  NAND3_X2 U4366 ( .A1(n48253), .A2(n64922), .A3(n48165), .ZN(n200) );
  BUF_X4 U4375 ( .I(n53597), .Z(n53700) );
  INV_X4 U4376 ( .I(n58572), .ZN(n5368) );
  NAND3_X1 U4379 ( .A1(n15199), .A2(n61984), .A3(n40444), .ZN(n15198) );
  OAI21_X1 U4381 ( .A1(n15198), .A2(n16925), .B(n985), .ZN(n64682) );
  OAI21_X2 U4385 ( .A1(n41112), .A2(n15139), .B(n971), .ZN(n40573) );
  NAND2_X2 U4386 ( .A1(n57070), .A2(n13567), .ZN(n62225) );
  NAND2_X2 U4388 ( .A1(n54189), .A2(n54207), .ZN(n54144) );
  NAND2_X2 U4390 ( .A1(n23125), .A2(n34026), .ZN(n17895) );
  NOR2_X1 U4391 ( .A1(n61144), .A2(n2354), .ZN(n2352) );
  BUF_X8 U4393 ( .I(n61728), .Z(n1474) );
  INV_X2 U4395 ( .I(n57083), .ZN(n63781) );
  BUF_X4 U4396 ( .I(n52604), .Z(n24040) );
  NAND2_X2 U4398 ( .A1(n30341), .A2(n29083), .ZN(n28565) );
  NAND2_X1 U4403 ( .A1(n4676), .A2(n4677), .ZN(n63409) );
  BUF_X4 U4410 ( .I(n56600), .Z(n61405) );
  NOR2_X1 U4412 ( .A1(n16929), .A2(n64682), .ZN(n18399) );
  NAND3_X2 U4413 ( .A1(n58043), .A2(n58042), .A3(n48202), .ZN(n62029) );
  NAND3_X2 U4414 ( .A1(n34552), .A2(n34551), .A3(n17895), .ZN(n34563) );
  NAND2_X2 U4416 ( .A1(n16673), .A2(n16672), .ZN(n63719) );
  NOR3_X2 U4417 ( .A1(n28291), .A2(n17268), .A3(n58448), .ZN(n28295) );
  INV_X2 U4421 ( .I(n14871), .ZN(n64718) );
  AND2_X2 U4422 ( .A1(n40776), .A2(n43516), .Z(n43515) );
  INV_X2 U4424 ( .I(n50215), .ZN(n13537) );
  BUF_X4 U4425 ( .I(n36951), .Z(n5936) );
  NOR2_X2 U4431 ( .A1(n29148), .A2(n6888), .ZN(n64506) );
  NAND2_X2 U4437 ( .A1(n60962), .A2(n57353), .ZN(n64086) );
  BUF_X4 U4439 ( .I(n53755), .Z(n16489) );
  NAND2_X2 U4441 ( .A1(n22516), .A2(n57143), .ZN(n57102) );
  NOR3_X1 U4444 ( .A1(n48378), .A2(n48980), .A3(n49453), .ZN(n62079) );
  INV_X2 U4448 ( .I(n24529), .ZN(n3250) );
  NOR2_X2 U4450 ( .A1(n56616), .A2(n56689), .ZN(n13249) );
  NOR3_X2 U4452 ( .A1(n54198), .A2(n54187), .A3(n25299), .ZN(n13710) );
  NOR2_X2 U4460 ( .A1(n45787), .A2(n20299), .ZN(n47027) );
  BUF_X4 U4462 ( .I(n22573), .Z(n12153) );
  NAND2_X2 U4469 ( .A1(n24696), .A2(n15875), .ZN(n56364) );
  BUF_X2 U4479 ( .I(n9378), .Z(n63667) );
  NOR3_X2 U4480 ( .A1(n8198), .A2(n47159), .A3(n47158), .ZN(n63765) );
  NOR2_X2 U4489 ( .A1(n60786), .A2(n50303), .ZN(n48580) );
  NAND3_X2 U4492 ( .A1(n53601), .A2(n53602), .A3(n2001), .ZN(n53604) );
  NAND2_X2 U4502 ( .A1(n23316), .A2(n48518), .ZN(n48519) );
  INV_X2 U4504 ( .I(n7596), .ZN(n20491) );
  NAND3_X2 U4510 ( .A1(n23028), .A2(n48710), .A3(n49091), .ZN(n48715) );
  NAND2_X2 U4511 ( .A1(n1282), .A2(n14360), .ZN(n55352) );
  NAND2_X2 U4518 ( .A1(n54276), .A2(n51878), .ZN(n13263) );
  NAND2_X2 U4519 ( .A1(n8818), .A2(n1200), .ZN(n6019) );
  NAND3_X2 U4524 ( .A1(n52477), .A2(n54997), .A3(n24870), .ZN(n55269) );
  BUF_X4 U4526 ( .I(n54062), .Z(n3888) );
  BUF_X4 U4530 ( .I(n14522), .Z(n12112) );
  OAI21_X1 U4531 ( .A1(n2417), .A2(n28688), .B(n2416), .ZN(n65049) );
  NAND3_X2 U4532 ( .A1(n30738), .A2(n20172), .A3(n31208), .ZN(n13031) );
  INV_X2 U4536 ( .I(n37285), .ZN(n59576) );
  NOR2_X2 U4539 ( .A1(n28381), .A2(n13704), .ZN(n26633) );
  INV_X2 U4543 ( .I(n35842), .ZN(n64884) );
  NAND2_X1 U4544 ( .A1(n35458), .A2(n62198), .ZN(n63896) );
  AOI21_X2 U4545 ( .A1(n56280), .A2(n51262), .B(n56574), .ZN(n51273) );
  INV_X2 U4548 ( .I(n28494), .ZN(n27830) );
  BUF_X4 U4549 ( .I(n5349), .Z(n411) );
  NOR2_X2 U4550 ( .A1(n11425), .A2(n23168), .ZN(n28707) );
  NAND2_X2 U4553 ( .A1(n4035), .A2(n22785), .ZN(n36559) );
  OAI21_X2 U4554 ( .A1(n1860), .A2(n1277), .B(n9186), .ZN(n18397) );
  AND2_X2 U4558 ( .A1(n60583), .A2(n10990), .Z(n61816) );
  NAND2_X2 U4559 ( .A1(n6779), .A2(n32076), .ZN(n37187) );
  NAND2_X2 U4560 ( .A1(n56530), .A2(n56541), .ZN(n51347) );
  NOR3_X2 U4566 ( .A1(n13614), .A2(n24374), .A3(n48318), .ZN(n48024) );
  INV_X2 U4572 ( .I(n2842), .ZN(n6885) );
  BUF_X4 U4574 ( .I(n64950), .Z(n22799) );
  INV_X8 U4575 ( .I(n15252), .ZN(n1298) );
  AOI21_X2 U4581 ( .A1(n47254), .A2(n47253), .B(n47263), .ZN(n63373) );
  BUF_X2 U4583 ( .I(n38931), .Z(n40408) );
  INV_X2 U4584 ( .I(n6577), .ZN(n13166) );
  NOR3_X2 U4585 ( .A1(n30738), .A2(n14217), .A3(n31201), .ZN(n30742) );
  BUF_X4 U4588 ( .I(n28448), .Z(n22312) );
  BUF_X4 U4591 ( .I(n35723), .Z(n23449) );
  INV_X4 U4592 ( .I(n41444), .ZN(n39847) );
  INV_X2 U4598 ( .I(n16503), .ZN(n1282) );
  CLKBUF_X2 U4599 ( .I(n54862), .Z(n671) );
  NAND2_X1 U4604 ( .A1(n3939), .A2(n35775), .ZN(n35785) );
  INV_X2 U4607 ( .I(n35775), .ZN(n1544) );
  INV_X2 U4608 ( .I(n2641), .ZN(n2640) );
  NAND2_X1 U4609 ( .A1(n2640), .A2(n24114), .ZN(n2644) );
  NAND4_X1 U4612 ( .A1(n52657), .A2(n52658), .A3(n52656), .A4(n52655), .ZN(
        n20766) );
  INV_X2 U4619 ( .I(n4723), .ZN(n42399) );
  NOR2_X1 U4629 ( .A1(n1396), .A2(n4723), .ZN(n42410) );
  NAND3_X1 U4630 ( .A1(n1688), .A2(n41693), .A3(n4723), .ZN(n6613) );
  NAND2_X1 U4631 ( .A1(n4723), .A2(n42404), .ZN(n42079) );
  CLKBUF_X4 U4632 ( .I(n2950), .Z(n2876) );
  NAND2_X1 U4633 ( .A1(n55148), .A2(n7983), .ZN(n55136) );
  NOR2_X1 U4639 ( .A1(n53852), .A2(n53622), .ZN(n53025) );
  CLKBUF_X4 U4641 ( .I(n9550), .Z(n62699) );
  NOR3_X1 U4642 ( .A1(n1593), .A2(n9550), .A3(n55156), .ZN(n7983) );
  INV_X2 U4650 ( .I(n1334), .ZN(n9162) );
  AOI22_X1 U4651 ( .A1(n1334), .A2(n43309), .B1(n24071), .B2(n62462), .ZN(
        n21140) );
  NOR2_X1 U4653 ( .A1(n54560), .A2(n22217), .ZN(n54577) );
  BUF_X2 U4655 ( .I(n47290), .Z(n22549) );
  NOR2_X1 U4662 ( .A1(n23407), .A2(n14448), .ZN(n15076) );
  NAND2_X1 U4663 ( .A1(n62247), .A2(n23407), .ZN(n62180) );
  NAND4_X1 U4665 ( .A1(n17224), .A2(n47990), .A3(n59004), .A4(n22570), .ZN(
        n17088) );
  NOR2_X1 U4668 ( .A1(n20930), .A2(n29356), .ZN(n27504) );
  NAND3_X1 U4669 ( .A1(n61169), .A2(n26217), .A3(n29175), .ZN(n64388) );
  OAI21_X1 U4670 ( .A1(n29016), .A2(n25241), .B(n1318), .ZN(n21251) );
  INV_X1 U4671 ( .I(n38234), .ZN(n42503) );
  INV_X1 U4682 ( .I(n54087), .ZN(n54595) );
  INV_X1 U4683 ( .I(n53427), .ZN(n53416) );
  NAND3_X1 U4689 ( .A1(n53321), .A2(n16778), .A3(n9731), .ZN(n52797) );
  NOR2_X1 U4693 ( .A1(n54726), .A2(n54759), .ZN(n54737) );
  NAND2_X1 U4695 ( .A1(n47371), .A2(n23934), .ZN(n45412) );
  NOR2_X1 U4696 ( .A1(n64334), .A2(n64442), .ZN(n63160) );
  AOI21_X1 U4697 ( .A1(n61192), .A2(n55658), .B(n24404), .ZN(n64442) );
  NAND2_X1 U4703 ( .A1(n9346), .A2(n7086), .ZN(n49264) );
  NAND2_X1 U4704 ( .A1(n49068), .A2(n49073), .ZN(n58723) );
  NAND2_X1 U4706 ( .A1(n47452), .A2(n49068), .ZN(n47453) );
  NOR2_X1 U4711 ( .A1(n2820), .A2(n23856), .ZN(n58109) );
  NOR2_X1 U4712 ( .A1(n65196), .A2(n47736), .ZN(n47738) );
  NAND2_X1 U4716 ( .A1(n56635), .A2(n21066), .ZN(n56422) );
  INV_X1 U4718 ( .I(n55906), .ZN(n59806) );
  NAND3_X1 U4725 ( .A1(n16776), .A2(n53366), .A3(n53361), .ZN(n62020) );
  INV_X1 U4730 ( .I(n45990), .ZN(n47625) );
  NOR2_X1 U4731 ( .A1(n45990), .A2(n60979), .ZN(n45206) );
  OR3_X2 U4745 ( .A1(n45990), .A2(n62739), .A3(n61601), .Z(n47628) );
  BUF_X2 U4748 ( .I(n20349), .Z(n58763) );
  AOI21_X1 U4752 ( .A1(n608), .A2(n1517), .B(n40062), .ZN(n22051) );
  NAND2_X1 U4754 ( .A1(n1932), .A2(n41814), .ZN(n41824) );
  INV_X1 U4758 ( .I(n21279), .ZN(n22772) );
  CLKBUF_X2 U4761 ( .I(n54950), .Z(n58994) );
  CLKBUF_X2 U4764 ( .I(n46292), .Z(n10043) );
  INV_X1 U4765 ( .I(n12454), .ZN(n56850) );
  NOR2_X1 U4767 ( .A1(n15930), .A2(n21679), .ZN(n21171) );
  NAND2_X1 U4768 ( .A1(n22122), .A2(n62577), .ZN(n54740) );
  AND2_X1 U4772 ( .A1(n56531), .A2(n56546), .Z(n61871) );
  INV_X1 U4773 ( .I(n50305), .ZN(n8096) );
  NAND3_X1 U4775 ( .A1(n54192), .A2(n54198), .A3(n2984), .ZN(n54186) );
  NAND2_X1 U4776 ( .A1(n7977), .A2(n56716), .ZN(n62390) );
  NAND2_X1 U4777 ( .A1(n57720), .A2(n58514), .ZN(n58513) );
  INV_X2 U4778 ( .I(n58514), .ZN(n55469) );
  NOR2_X1 U4779 ( .A1(n14577), .A2(n11803), .ZN(n14576) );
  NAND3_X1 U4789 ( .A1(n39846), .A2(n64773), .A3(n40374), .ZN(n39602) );
  NAND3_X1 U4792 ( .A1(n53521), .A2(n62095), .A3(n62094), .ZN(n17098) );
  NOR3_X1 U4795 ( .A1(n7298), .A2(n57893), .A3(n412), .ZN(n44863) );
  CLKBUF_X1 U4796 ( .I(n177), .Z(n57893) );
  NAND2_X1 U4799 ( .A1(n13549), .A2(n57194), .ZN(n14005) );
  NOR2_X1 U4800 ( .A1(n56364), .A2(n60809), .ZN(n63138) );
  INV_X2 U4814 ( .I(n23538), .ZN(n25147) );
  NAND2_X1 U4817 ( .A1(n57124), .A2(n23538), .ZN(n57125) );
  NOR2_X1 U4820 ( .A1(n22764), .A2(n8995), .ZN(n62255) );
  BUF_X1 U4826 ( .I(n22764), .Z(n59021) );
  NAND2_X1 U4828 ( .A1(n57414), .A2(n55244), .ZN(n54792) );
  INV_X1 U4831 ( .I(n53480), .ZN(n53515) );
  NAND3_X1 U4832 ( .A1(n7866), .A2(n50441), .A3(n19144), .ZN(n50233) );
  NAND2_X1 U4833 ( .A1(n55829), .A2(n14890), .ZN(n62957) );
  INV_X2 U4834 ( .I(n16342), .ZN(n14890) );
  OR2_X1 U4836 ( .A1(n55709), .A2(n61368), .Z(n61817) );
  INV_X1 U4838 ( .I(n55153), .ZN(n55159) );
  NAND2_X1 U4839 ( .A1(n45991), .A2(n59802), .ZN(n47239) );
  OAI21_X1 U4842 ( .A1(n8324), .A2(n8323), .B(n25638), .ZN(n8318) );
  INV_X1 U4844 ( .I(n6790), .ZN(n53279) );
  BUF_X4 U4848 ( .I(n50399), .Z(n1381) );
  NAND2_X1 U4849 ( .A1(n50406), .A2(n50399), .ZN(n49729) );
  NOR2_X1 U4858 ( .A1(n53688), .A2(n19475), .ZN(n53665) );
  OAI22_X1 U4863 ( .A1(n22747), .A2(n14966), .B1(n50576), .B2(n52323), .ZN(
        n7614) );
  INV_X2 U4873 ( .I(n39517), .ZN(n23890) );
  BUF_X2 U4879 ( .I(n39517), .Z(n64672) );
  NOR2_X1 U4881 ( .A1(n56049), .A2(n56050), .ZN(n56089) );
  NAND2_X1 U4882 ( .A1(n55412), .A2(n55416), .ZN(n54790) );
  NAND2_X1 U4884 ( .A1(n4646), .A2(n48602), .ZN(n352) );
  NOR2_X1 U4888 ( .A1(n3086), .A2(n23140), .ZN(n29942) );
  INV_X1 U4891 ( .I(n15713), .ZN(n60200) );
  CLKBUF_X2 U4901 ( .I(n45614), .Z(n62975) );
  NOR2_X1 U4903 ( .A1(n56856), .A2(n56850), .ZN(n56873) );
  CLKBUF_X4 U4904 ( .I(n15785), .Z(n15713) );
  NOR2_X1 U4908 ( .A1(n56256), .A2(n56586), .ZN(n56411) );
  NOR2_X1 U4909 ( .A1(n63767), .A2(n63006), .ZN(n53092) );
  NAND2_X1 U4914 ( .A1(n58154), .A2(n1177), .ZN(n3545) );
  NAND4_X1 U4919 ( .A1(n780), .A2(n1177), .A3(n59260), .A4(n53137), .ZN(n53139) );
  NAND2_X1 U4924 ( .A1(n55092), .A2(n55056), .ZN(n55084) );
  NAND2_X1 U4927 ( .A1(n57694), .A2(n57693), .ZN(n57692) );
  NAND2_X1 U4928 ( .A1(n54531), .A2(n54572), .ZN(n54540) );
  INV_X1 U4929 ( .I(n51548), .ZN(n49209) );
  NAND2_X1 U4934 ( .A1(n39835), .A2(n39485), .ZN(n4951) );
  NAND4_X1 U4940 ( .A1(n39837), .A2(n39835), .A3(n25358), .A4(n39836), .ZN(
        n39838) );
  NAND2_X1 U4941 ( .A1(n39486), .A2(n25356), .ZN(n39835) );
  NAND3_X1 U4944 ( .A1(n28610), .A2(n28452), .A3(n63330), .ZN(n28455) );
  NOR2_X1 U4946 ( .A1(n28610), .A2(n28609), .ZN(n13010) );
  BUF_X2 U4947 ( .I(n50780), .Z(n17597) );
  NAND2_X1 U4948 ( .A1(n15606), .A2(n61719), .ZN(n58521) );
  NAND3_X1 U4952 ( .A1(n3111), .A2(n48466), .A3(n48464), .ZN(n15606) );
  BUF_X2 U4953 ( .I(n25253), .Z(n61070) );
  NAND2_X1 U4954 ( .A1(n58206), .A2(n25253), .ZN(n48059) );
  NAND2_X1 U4955 ( .A1(n56048), .A2(n9567), .ZN(n56014) );
  CLKBUF_X4 U4959 ( .I(n22083), .Z(n6216) );
  NAND2_X1 U4964 ( .A1(n1146), .A2(n54966), .ZN(n54968) );
  NAND3_X1 U4965 ( .A1(n54626), .A2(n1146), .A3(n23122), .ZN(n54627) );
  NOR4_X1 U4968 ( .A1(n9003), .A2(n11521), .A3(n60370), .A4(n55659), .ZN(
        n64334) );
  INV_X1 U4972 ( .I(n50236), .ZN(n17887) );
  NOR2_X1 U4975 ( .A1(n5129), .A2(n1324), .ZN(n55911) );
  OR2_X1 U4976 ( .A1(n5194), .A2(n56190), .Z(n56168) );
  NAND3_X1 U4978 ( .A1(n15132), .A2(n56433), .A3(n56434), .ZN(n56440) );
  BUF_X2 U4981 ( .I(n20548), .Z(n3129) );
  CLKBUF_X2 U4984 ( .I(n3129), .Z(n3128) );
  CLKBUF_X4 U4987 ( .I(n53163), .Z(n23856) );
  INV_X1 U4990 ( .I(n55619), .ZN(n55632) );
  OR2_X1 U4991 ( .A1(n13693), .A2(n9655), .Z(n56929) );
  BUF_X2 U4999 ( .I(n35019), .Z(n36965) );
  NOR2_X1 U5001 ( .A1(n1578), .A2(n59599), .ZN(n382) );
  INV_X1 U5005 ( .I(n14484), .ZN(n1578) );
  INV_X1 U5006 ( .I(n56824), .ZN(n56874) );
  OAI22_X1 U5010 ( .A1(n52732), .A2(n52731), .B1(n52730), .B2(n56824), .ZN(
        n52733) );
  NAND2_X1 U5011 ( .A1(n23682), .A2(n5585), .ZN(n56824) );
  NAND2_X1 U5016 ( .A1(n4541), .A2(n6159), .ZN(n37354) );
  CLKBUF_X2 U5017 ( .I(n6159), .Z(n59011) );
  INV_X1 U5019 ( .I(n23485), .ZN(n43837) );
  AOI21_X1 U5021 ( .A1(n56003), .A2(n55999), .B(n55998), .ZN(n56006) );
  INV_X1 U5023 ( .I(n56082), .ZN(n56003) );
  OAI21_X1 U5025 ( .A1(n54172), .A2(n54198), .B(n54192), .ZN(n54117) );
  INV_X1 U5029 ( .I(n3606), .ZN(n42195) );
  INV_X1 U5030 ( .I(n43549), .ZN(n20372) );
  NOR2_X1 U5042 ( .A1(n62530), .A2(n43549), .ZN(n16710) );
  INV_X1 U5043 ( .I(n25320), .ZN(n65057) );
  AOI21_X1 U5046 ( .A1(n47263), .A2(n21793), .B(n47262), .ZN(n47264) );
  INV_X1 U5052 ( .I(n53054), .ZN(n53111) );
  NOR3_X1 U5054 ( .A1(n53054), .A2(n52896), .A3(n63767), .ZN(n53116) );
  OAI21_X1 U5055 ( .A1(n53054), .A2(n23243), .B(n53080), .ZN(n23290) );
  INV_X1 U5058 ( .I(n50141), .ZN(n50297) );
  NAND3_X1 U5068 ( .A1(n50141), .A2(n9646), .A3(n1643), .ZN(n50313) );
  NAND2_X1 U5070 ( .A1(n61311), .A2(n1209), .ZN(n1121) );
  NOR2_X1 U5078 ( .A1(n43343), .A2(n61134), .ZN(n41592) );
  NAND2_X1 U5082 ( .A1(n40146), .A2(n6625), .ZN(n40993) );
  INV_X2 U5083 ( .I(n40146), .ZN(n40986) );
  AOI21_X1 U5085 ( .A1(n55477), .A2(n55478), .B(n55741), .ZN(n62605) );
  NOR3_X1 U5086 ( .A1(n55476), .A2(n55475), .A3(n22592), .ZN(n55741) );
  NOR2_X1 U5087 ( .A1(n20549), .A2(n34176), .ZN(n3131) );
  CLKBUF_X4 U5091 ( .I(n14731), .Z(n14730) );
  NAND2_X1 U5092 ( .A1(n23595), .A2(n53079), .ZN(n53081) );
  OAI22_X1 U5094 ( .A1(n57062), .A2(n13567), .B1(n57068), .B2(n21079), .ZN(
        n57064) );
  INV_X1 U5095 ( .I(n53513), .ZN(n14021) );
  NOR3_X1 U5097 ( .A1(n16779), .A2(n16777), .A3(n62020), .ZN(n59673) );
  NAND2_X1 U5098 ( .A1(n58380), .A2(n56214), .ZN(n63361) );
  NAND2_X1 U5099 ( .A1(n53410), .A2(n54055), .ZN(n53411) );
  INV_X1 U5100 ( .I(n52465), .ZN(n58731) );
  NAND2_X1 U5109 ( .A1(n36075), .A2(n36304), .ZN(n36793) );
  AOI21_X1 U5112 ( .A1(n52123), .A2(n55719), .B(n59806), .ZN(n9974) );
  AOI22_X1 U5119 ( .A1(n21028), .A2(n52786), .B1(n53444), .B2(n52814), .ZN(
        n64028) );
  NOR3_X1 U5120 ( .A1(n9825), .A2(n44792), .A3(n9824), .ZN(n25561) );
  NAND2_X1 U5121 ( .A1(n56962), .A2(n1583), .ZN(n56906) );
  INV_X2 U5122 ( .I(n14424), .ZN(n51790) );
  BUF_X2 U5136 ( .I(n55738), .Z(n22588) );
  NAND2_X1 U5137 ( .A1(n11556), .A2(n54409), .ZN(n54362) );
  BUF_X2 U5138 ( .I(n11556), .Z(n4688) );
  NAND2_X1 U5142 ( .A1(n25253), .A2(n5481), .ZN(n2477) );
  INV_X2 U5146 ( .I(n56344), .ZN(n56342) );
  NAND2_X1 U5147 ( .A1(n55644), .A2(n55631), .ZN(n55642) );
  OAI21_X1 U5148 ( .A1(n64227), .A2(n56631), .B(n63359), .ZN(n56130) );
  OAI21_X1 U5160 ( .A1(n56631), .A2(n21893), .B(n56417), .ZN(n52716) );
  NAND2_X1 U5164 ( .A1(n23165), .A2(n56631), .ZN(n56415) );
  BUF_X2 U5165 ( .I(n56631), .Z(n58846) );
  NAND2_X1 U5168 ( .A1(n61693), .A2(n57470), .ZN(n19658) );
  NOR2_X1 U5169 ( .A1(n53006), .A2(n53455), .ZN(n52771) );
  NAND2_X1 U5180 ( .A1(n22684), .A2(n9152), .ZN(n48599) );
  NOR2_X1 U5182 ( .A1(n9152), .A2(n5771), .ZN(n47005) );
  NAND2_X1 U5183 ( .A1(n55146), .A2(n55145), .ZN(n55154) );
  NAND2_X1 U5187 ( .A1(n14333), .A2(n23796), .ZN(n17555) );
  AOI21_X1 U5188 ( .A1(n56885), .A2(n64230), .B(n62800), .ZN(n52730) );
  NAND2_X1 U5193 ( .A1(n10862), .A2(n53519), .ZN(n53521) );
  NOR2_X1 U5194 ( .A1(n63948), .A2(n974), .ZN(n60329) );
  CLKBUF_X2 U5197 ( .I(n12615), .Z(n64896) );
  NAND2_X1 U5201 ( .A1(n22842), .A2(n46367), .ZN(n48957) );
  CLKBUF_X4 U5206 ( .I(n55746), .Z(n55821) );
  NOR3_X1 U5214 ( .A1(n52230), .A2(n58146), .A3(n52231), .ZN(n50816) );
  NOR2_X1 U5220 ( .A1(n57002), .A2(n23110), .ZN(n53239) );
  NAND4_X1 U5221 ( .A1(n56712), .A2(n56713), .A3(n56711), .A4(n56710), .ZN(
        n58265) );
  INV_X1 U5222 ( .I(n53737), .ZN(n1577) );
  NAND3_X1 U5227 ( .A1(n56407), .A2(n14307), .A3(n22473), .ZN(n56581) );
  NAND2_X1 U5230 ( .A1(n41980), .A2(n58572), .ZN(n42359) );
  BUF_X2 U5236 ( .I(n58572), .Z(n62435) );
  NAND2_X1 U5238 ( .A1(n20922), .A2(n58572), .ZN(n5075) );
  CLKBUF_X2 U5240 ( .I(n3172), .Z(n62399) );
  NOR2_X1 U5242 ( .A1(n9136), .A2(n23704), .ZN(n13601) );
  NOR2_X1 U5244 ( .A1(n53557), .A2(n53916), .ZN(n53566) );
  INV_X1 U5247 ( .I(n53557), .ZN(n53403) );
  NAND3_X1 U5248 ( .A1(n63228), .A2(n41206), .A3(n40733), .ZN(n63948) );
  NAND2_X1 U5250 ( .A1(n39029), .A2(n38677), .ZN(n40733) );
  CLKBUF_X2 U5251 ( .I(n30648), .Z(n63537) );
  CLKBUF_X4 U5254 ( .I(n30648), .Z(n3086) );
  NAND3_X1 U5255 ( .A1(n6947), .A2(n6949), .A3(n6946), .ZN(n62171) );
  NOR3_X1 U5259 ( .A1(n64483), .A2(n62293), .A3(n64482), .ZN(n6947) );
  NAND2_X1 U5260 ( .A1(n1366), .A2(n61964), .ZN(n645) );
  BUF_X2 U5264 ( .I(n22794), .Z(n10389) );
  NOR2_X1 U5265 ( .A1(n61529), .A2(n63020), .ZN(n54920) );
  NOR2_X1 U5270 ( .A1(n56731), .A2(n56722), .ZN(n56718) );
  CLKBUF_X4 U5271 ( .I(n56897), .Z(n23074) );
  NAND2_X1 U5272 ( .A1(n56225), .A2(n15132), .ZN(n55713) );
  NAND4_X1 U5276 ( .A1(n54674), .A2(n54675), .A3(n18564), .A4(n54673), .ZN(
        n59716) );
  OAI21_X1 U5277 ( .A1(n15706), .A2(n5550), .B(n56266), .ZN(n5328) );
  CLKBUF_X4 U5287 ( .I(n55280), .Z(n2180) );
  INV_X1 U5291 ( .I(n3741), .ZN(n51308) );
  CLKBUF_X2 U5292 ( .I(n3741), .Z(n59787) );
  INV_X2 U5293 ( .I(n47435), .ZN(n47746) );
  BUF_X2 U5297 ( .I(n47435), .Z(n63647) );
  CLKBUF_X2 U5303 ( .I(n25997), .Z(n64750) );
  AND2_X1 U5308 ( .A1(n53130), .A2(n53167), .Z(n53158) );
  NAND2_X1 U5311 ( .A1(n53167), .A2(n7182), .ZN(n7181) );
  NAND3_X1 U5313 ( .A1(n53167), .A2(n23856), .A3(n12111), .ZN(n12156) );
  CLKBUF_X2 U5314 ( .I(n22092), .Z(n15632) );
  NAND2_X1 U5321 ( .A1(n59695), .A2(n8691), .ZN(n47659) );
  CLKBUF_X4 U5325 ( .I(n23505), .Z(n21169) );
  OAI21_X1 U5330 ( .A1(n21983), .A2(n21982), .B(n53539), .ZN(n15059) );
  NOR2_X1 U5331 ( .A1(n53184), .A2(n1457), .ZN(n21983) );
  NOR2_X1 U5333 ( .A1(n61961), .A2(n61025), .ZN(n45222) );
  NAND2_X1 U5335 ( .A1(n54489), .A2(n21030), .ZN(n64491) );
  NOR2_X1 U5341 ( .A1(n53700), .A2(n53667), .ZN(n53697) );
  OAI22_X1 U5342 ( .A1(n4323), .A2(n47964), .B1(n48416), .B2(n12595), .ZN(
        n7692) );
  NAND3_X1 U5349 ( .A1(n56217), .A2(n60129), .A3(n56205), .ZN(n56213) );
  NAND2_X1 U5353 ( .A1(n21073), .A2(n43924), .ZN(n43490) );
  BUF_X2 U5361 ( .I(n43924), .Z(n20276) );
  INV_X1 U5371 ( .I(n44156), .ZN(n4049) );
  CLKBUF_X4 U5373 ( .I(n20547), .Z(n10869) );
  NAND2_X1 U5377 ( .A1(n20547), .A2(n19567), .ZN(n53184) );
  INV_X1 U5382 ( .I(n23116), .ZN(n2040) );
  NOR2_X1 U5385 ( .A1(n24421), .A2(n20657), .ZN(n60393) );
  INV_X1 U5390 ( .I(n53301), .ZN(n53293) );
  AOI21_X1 U5391 ( .A1(n53306), .A2(n53301), .B(n6790), .ZN(n62293) );
  NOR3_X1 U5393 ( .A1(n61228), .A2(n23258), .A3(n56168), .ZN(n56148) );
  INV_X1 U5394 ( .I(n3734), .ZN(n50209) );
  BUF_X2 U5396 ( .I(n3734), .Z(n60428) );
  NAND2_X1 U5404 ( .A1(n23411), .A2(n53303), .ZN(n53247) );
  NAND4_X1 U5405 ( .A1(n7654), .A2(n13328), .A3(n54436), .A4(n13329), .ZN(
        n13327) );
  CLKBUF_X4 U5406 ( .I(n56190), .Z(n11716) );
  INV_X1 U5407 ( .I(n17211), .ZN(n51263) );
  NAND3_X1 U5409 ( .A1(n54380), .A2(n54424), .A3(n1367), .ZN(n54397) );
  CLKBUF_X1 U5413 ( .I(n1519), .Z(n63032) );
  CLKBUF_X2 U5418 ( .I(n5382), .Z(n5317) );
  NAND2_X1 U5419 ( .A1(n53081), .A2(n19080), .ZN(n23289) );
  NAND2_X1 U5422 ( .A1(n63006), .A2(n19080), .ZN(n53082) );
  NOR2_X1 U5423 ( .A1(n43175), .A2(n43506), .ZN(n20495) );
  CLKBUF_X2 U5424 ( .I(n59538), .Z(n62822) );
  NAND2_X1 U5426 ( .A1(n56963), .A2(n19708), .ZN(n19707) );
  NAND2_X1 U5428 ( .A1(n54997), .A2(n11237), .ZN(n18790) );
  CLKBUF_X2 U5430 ( .I(n15252), .Z(n60432) );
  OR2_X1 U5431 ( .A1(n15252), .A2(n61739), .Z(n61858) );
  NOR2_X1 U5434 ( .A1(n47127), .A2(n48560), .ZN(n48567) );
  NAND2_X1 U5435 ( .A1(n53240), .A2(n53239), .ZN(n63987) );
  NOR2_X1 U5440 ( .A1(n19658), .A2(n57004), .ZN(n53240) );
  CLKBUF_X1 U5444 ( .I(n11528), .Z(n20072) );
  NAND3_X1 U5445 ( .A1(n18130), .A2(n12407), .A3(n62347), .ZN(n62592) );
  NOR2_X1 U5449 ( .A1(n17054), .A2(n17053), .ZN(n63562) );
  AND2_X1 U5450 ( .A1(n26200), .A2(n58526), .Z(n54451) );
  NAND4_X1 U5454 ( .A1(n54515), .A2(n23229), .A3(n678), .A4(n677), .ZN(n61400)
         );
  NAND4_X1 U5455 ( .A1(n50305), .A2(n50306), .A3(n50304), .A4(n50303), .ZN(
        n63803) );
  CLKBUF_X2 U5458 ( .I(n6853), .Z(n4383) );
  NAND2_X1 U5461 ( .A1(n4724), .A2(n47041), .ZN(n48393) );
  AOI21_X1 U5465 ( .A1(n50820), .A2(n50821), .B(n62539), .ZN(n50826) );
  CLKBUF_X2 U5467 ( .I(n18145), .Z(n16500) );
  NOR2_X1 U5474 ( .A1(n54526), .A2(n54576), .ZN(n54562) );
  NAND2_X1 U5480 ( .A1(n49277), .A2(n57194), .ZN(n48930) );
  NOR2_X1 U5488 ( .A1(n53145), .A2(n53147), .ZN(n64776) );
  INV_X1 U5489 ( .I(n21130), .ZN(n59250) );
  NAND2_X1 U5498 ( .A1(n63020), .A2(n14635), .ZN(n54880) );
  NAND2_X1 U5504 ( .A1(n52698), .A2(n13800), .ZN(n24421) );
  OAI22_X1 U5509 ( .A1(n23241), .A2(n36423), .B1(n6883), .B2(n12804), .ZN(
        n58988) );
  NAND3_X1 U5510 ( .A1(n36425), .A2(n36432), .A3(n12804), .ZN(n14683) );
  AOI22_X1 U5512 ( .A1(n36125), .A2(n12804), .B1(n36423), .B2(n59468), .ZN(
        n63083) );
  NOR2_X1 U5513 ( .A1(n23650), .A2(n12580), .ZN(n50090) );
  OAI21_X1 U5528 ( .A1(n50098), .A2(n50097), .B(n23650), .ZN(n12001) );
  NAND2_X1 U5531 ( .A1(n15386), .A2(n23650), .ZN(n24583) );
  NOR2_X1 U5532 ( .A1(n23650), .A2(n12579), .ZN(n50099) );
  NAND2_X1 U5538 ( .A1(n12692), .A2(n7148), .ZN(n54855) );
  INV_X1 U5543 ( .I(n19904), .ZN(n41950) );
  INV_X2 U5544 ( .I(n14624), .ZN(n41064) );
  CLKBUF_X4 U5545 ( .I(n14624), .Z(n20598) );
  NAND2_X1 U5549 ( .A1(n65150), .A2(n6305), .ZN(n7337) );
  CLKBUF_X2 U5552 ( .I(n1603), .Z(n64019) );
  INV_X1 U5554 ( .I(n1603), .ZN(n1285) );
  NAND2_X1 U5557 ( .A1(n20965), .A2(n61371), .ZN(n17051) );
  AOI21_X1 U5563 ( .A1(n10237), .A2(n1325), .B(n23836), .ZN(n5684) );
  BUF_X2 U5567 ( .I(n13286), .Z(n13285) );
  OAI21_X1 U5573 ( .A1(n43513), .A2(n61744), .B(n43511), .ZN(n43514) );
  NAND2_X1 U5576 ( .A1(n65262), .A2(n43513), .ZN(n3026) );
  NAND2_X1 U5581 ( .A1(n47302), .A2(n1078), .ZN(n25476) );
  OAI22_X1 U5589 ( .A1(n45936), .A2(n46016), .B1(n1078), .B2(n45935), .ZN(
        n57544) );
  CLKBUF_X2 U5591 ( .I(n8260), .Z(n1219) );
  NAND3_X1 U5592 ( .A1(n51858), .A2(n51859), .A3(n54499), .ZN(n17053) );
  OAI22_X1 U5594 ( .A1(n43506), .A2(n61744), .B1(n43189), .B2(n42045), .ZN(
        n43510) );
  AOI22_X1 U5597 ( .A1(n53242), .A2(n57000), .B1(n6608), .B2(n1602), .ZN(
        n52698) );
  CLKBUF_X4 U5598 ( .I(n17620), .Z(n9311) );
  NOR2_X1 U5603 ( .A1(n57483), .A2(n25475), .ZN(n64616) );
  NAND3_X1 U5604 ( .A1(n12175), .A2(n34882), .A3(n35878), .ZN(n57483) );
  NAND2_X1 U5605 ( .A1(n47529), .A2(n5235), .ZN(n48604) );
  CLKBUF_X1 U5606 ( .I(n5235), .Z(n64118) );
  NAND2_X1 U5611 ( .A1(n5235), .A2(n8666), .ZN(n46095) );
  INV_X2 U5620 ( .I(n5235), .ZN(n47018) );
  OAI22_X1 U5622 ( .A1(n50421), .A2(n50427), .B1(n50426), .B2(n50420), .ZN(
        n50423) );
  INV_X2 U5633 ( .I(n48614), .ZN(n48624) );
  OAI22_X1 U5642 ( .A1(n47546), .A2(n48614), .B1(n47545), .B2(n47180), .ZN(
        n47548) );
  NOR2_X1 U5646 ( .A1(n1501), .A2(n7595), .ZN(n41984) );
  AOI22_X1 U5647 ( .A1(n53183), .A2(n50477), .B1(n50476), .B2(n53185), .ZN(
        n50485) );
  NAND2_X1 U5648 ( .A1(n19973), .A2(n11726), .ZN(n61288) );
  NAND2_X1 U5654 ( .A1(n47028), .A2(n195), .ZN(n44704) );
  NAND3_X1 U5658 ( .A1(n47028), .A2(n195), .A3(n20299), .ZN(n47037) );
  NAND4_X1 U5660 ( .A1(n54707), .A2(n54705), .A3(n54706), .A4(n19383), .ZN(
        n59880) );
  NAND4_X1 U5666 ( .A1(n41936), .A2(n42275), .A3(n59019), .A4(n42281), .ZN(
        n57844) );
  OAI21_X1 U5669 ( .A1(n41934), .A2(n978), .B(n42281), .ZN(n37597) );
  INV_X1 U5670 ( .I(n46941), .ZN(n47227) );
  OAI21_X1 U5674 ( .A1(n63670), .A2(n46941), .B(n46936), .ZN(n63634) );
  NAND3_X1 U5679 ( .A1(n45731), .A2(n46941), .A3(n47231), .ZN(n58445) );
  NAND2_X1 U5680 ( .A1(n45161), .A2(n24073), .ZN(n48889) );
  NAND2_X1 U5681 ( .A1(n24073), .A2(n19302), .ZN(n48898) );
  NAND2_X1 U5682 ( .A1(n24073), .A2(n22646), .ZN(n45165) );
  NOR2_X1 U5686 ( .A1(n24073), .A2(n48894), .ZN(n64936) );
  INV_X1 U5694 ( .I(n25970), .ZN(n15322) );
  INV_X1 U5695 ( .I(n45715), .ZN(n46038) );
  OAI21_X1 U5701 ( .A1(n13703), .A2(n49758), .B(n49757), .ZN(n24566) );
  OAI21_X1 U5703 ( .A1(n13703), .A2(n48887), .B(n48886), .ZN(n48901) );
  AOI22_X1 U5704 ( .A1(n48884), .A2(n48885), .B1(n48882), .B2(n9863), .ZN(
        n13703) );
  NAND3_X1 U5706 ( .A1(n48599), .A2(n2344), .A3(n20091), .ZN(n14369) );
  NOR2_X1 U5709 ( .A1(n24820), .A2(n2344), .ZN(n62220) );
  NAND3_X1 U5711 ( .A1(n20529), .A2(n48443), .A3(n48442), .ZN(n25529) );
  INV_X2 U5714 ( .I(n22835), .ZN(n33925) );
  NAND3_X1 U5717 ( .A1(n35325), .A2(n22835), .A3(n35770), .ZN(n33927) );
  NOR2_X1 U5718 ( .A1(n22835), .A2(n1544), .ZN(n12150) );
  AOI21_X1 U5719 ( .A1(n29251), .A2(n58237), .B(n29246), .ZN(n27628) );
  INV_X1 U5722 ( .I(n47831), .ZN(n57532) );
  NOR2_X1 U5728 ( .A1(n1658), .A2(n47831), .ZN(n62022) );
  NAND3_X1 U5730 ( .A1(n15091), .A2(n24361), .A3(n60948), .ZN(n23819) );
  NOR2_X1 U5731 ( .A1(n47316), .A2(n47310), .ZN(n62003) );
  NOR2_X1 U5736 ( .A1(n1070), .A2(n57731), .ZN(n44773) );
  INV_X1 U5737 ( .I(n1070), .ZN(n18477) );
  NOR3_X1 U5739 ( .A1(n12845), .A2(n48947), .A3(n49780), .ZN(n12844) );
  NOR2_X1 U5741 ( .A1(n50275), .A2(n13614), .ZN(n65072) );
  NOR2_X1 U5747 ( .A1(n20138), .A2(n13614), .ZN(n49942) );
  AOI21_X1 U5749 ( .A1(n63266), .A2(n20138), .B(n13614), .ZN(n63054) );
  NAND3_X1 U5750 ( .A1(n56507), .A2(n56506), .A3(n25704), .ZN(n25703) );
  INV_X2 U5752 ( .I(n12563), .ZN(n44826) );
  INV_X1 U5753 ( .I(n50339), .ZN(n50341) );
  NOR2_X1 U5754 ( .A1(n13988), .A2(n11624), .ZN(n21835) );
  INV_X1 U5756 ( .I(n25676), .ZN(n14537) );
  AOI21_X1 U5759 ( .A1(n15969), .A2(n54189), .B(n25299), .ZN(n54116) );
  AOI21_X1 U5760 ( .A1(n54189), .A2(n25299), .B(n54192), .ZN(n54130) );
  NOR2_X1 U5761 ( .A1(n22891), .A2(n25393), .ZN(n56318) );
  OAI21_X1 U5766 ( .A1(n12176), .A2(n2942), .B(n5807), .ZN(n12175) );
  OAI22_X1 U5768 ( .A1(n28965), .A2(n29905), .B1(n16517), .B2(n1866), .ZN(
        n28966) );
  INV_X1 U5769 ( .I(n7860), .ZN(n17863) );
  NAND2_X1 U5771 ( .A1(n18688), .A2(n47420), .ZN(n45800) );
  NAND2_X1 U5773 ( .A1(n11628), .A2(n13391), .ZN(n18688) );
  NAND2_X1 U5774 ( .A1(n19867), .A2(n15319), .ZN(n49555) );
  NAND3_X1 U5775 ( .A1(n22571), .A2(n24394), .A3(n19867), .ZN(n49550) );
  AOI22_X1 U5780 ( .A1(n40615), .A2(n64571), .B1(n19015), .B2(n39057), .ZN(
        n59593) );
  INV_X1 U5783 ( .I(n50019), .ZN(n49810) );
  INV_X1 U5787 ( .I(n55973), .ZN(n1600) );
  NAND2_X1 U5796 ( .A1(n17708), .A2(n55973), .ZN(n55968) );
  NAND3_X1 U5797 ( .A1(n55294), .A2(n4830), .A3(n55973), .ZN(n55970) );
  OR2_X1 U5799 ( .A1(n3966), .A2(n3962), .Z(n26246) );
  CLKBUF_X4 U5806 ( .I(n56516), .Z(n20587) );
  CLKBUF_X2 U5807 ( .I(n56516), .Z(n62421) );
  NAND2_X1 U5810 ( .A1(n56412), .A2(n14978), .ZN(n51888) );
  BUF_X2 U5811 ( .I(n56249), .Z(n22473) );
  NOR2_X1 U5812 ( .A1(n23538), .A2(n57146), .ZN(n57120) );
  NAND2_X1 U5813 ( .A1(n47801), .A2(n47802), .ZN(n18735) );
  BUF_X1 U5818 ( .I(n21894), .Z(n60946) );
  NOR2_X1 U5819 ( .A1(n56593), .A2(n56245), .ZN(n55957) );
  NAND2_X1 U5820 ( .A1(n16815), .A2(n49177), .ZN(n49265) );
  AND2_X1 U5823 ( .A1(n55218), .A2(n55233), .Z(n61768) );
  OAI21_X1 U5828 ( .A1(n61725), .A2(n54590), .B(n54595), .ZN(n53893) );
  AOI21_X1 U5834 ( .A1(n49256), .A2(n45458), .B(n45457), .ZN(n45461) );
  NAND2_X1 U5842 ( .A1(n20708), .A2(n23802), .ZN(n62006) );
  NAND2_X1 U5846 ( .A1(n46882), .A2(n47255), .ZN(n47248) );
  NAND2_X1 U5852 ( .A1(n46882), .A2(n16212), .ZN(n46078) );
  NAND3_X1 U5853 ( .A1(n12111), .A2(n2037), .A3(n53165), .ZN(n2712) );
  OAI21_X1 U5856 ( .A1(n2037), .A2(n23856), .B(n5614), .ZN(n50814) );
  NAND2_X1 U5857 ( .A1(n61012), .A2(n51886), .ZN(n9976) );
  NAND3_X1 U5868 ( .A1(n42110), .A2(n10415), .A3(n64363), .ZN(n38682) );
  BUF_X2 U5870 ( .I(n52278), .Z(n56962) );
  NOR2_X1 U5874 ( .A1(n35354), .A2(n6606), .ZN(n13745) );
  INV_X1 U5878 ( .I(n35354), .ZN(n1770) );
  OAI21_X1 U5881 ( .A1(n35964), .A2(n35543), .B(n35354), .ZN(n5088) );
  INV_X1 U5883 ( .I(n31989), .ZN(n1834) );
  NOR3_X1 U5886 ( .A1(n8259), .A2(n10381), .A3(n8194), .ZN(n52296) );
  OAI22_X1 U5887 ( .A1(n32886), .A2(n1535), .B1(n5410), .B2(n7047), .ZN(n20549) );
  NOR2_X1 U5888 ( .A1(n49598), .A2(n47444), .ZN(n49600) );
  NAND3_X1 U5889 ( .A1(n20045), .A2(n1615), .A3(n1595), .ZN(n61012) );
  NAND2_X1 U5891 ( .A1(n43003), .A2(n42994), .ZN(n43224) );
  NAND2_X1 U5894 ( .A1(n2179), .A2(n8047), .ZN(n47801) );
  NAND2_X1 U5895 ( .A1(n25527), .A2(n24728), .ZN(n30487) );
  NAND2_X1 U5897 ( .A1(n9392), .A2(n24728), .ZN(n29538) );
  NOR2_X1 U5898 ( .A1(n463), .A2(n24728), .ZN(n18917) );
  INV_X1 U5903 ( .I(n10364), .ZN(n15775) );
  INV_X2 U5904 ( .I(n46497), .ZN(n8021) );
  NAND2_X1 U5910 ( .A1(n9418), .A2(n9898), .ZN(n61620) );
  NAND2_X1 U5913 ( .A1(n61716), .A2(n3654), .ZN(n48058) );
  CLKBUF_X2 U5921 ( .I(n53823), .Z(n4540) );
  NAND2_X1 U5928 ( .A1(n56539), .A2(n22870), .ZN(n21732) );
  NAND2_X1 U5935 ( .A1(n21314), .A2(n28060), .ZN(n23397) );
  INV_X1 U5937 ( .I(n15726), .ZN(n62658) );
  OAI21_X1 U5939 ( .A1(n37942), .A2(n59825), .B(n33932), .ZN(n36645) );
  OAI21_X1 U5940 ( .A1(n59825), .A2(n37319), .B(n16380), .ZN(n37020) );
  AOI21_X1 U5941 ( .A1(n47921), .A2(n1474), .B(n61525), .ZN(n4624) );
  INV_X1 U5945 ( .I(n50425), .ZN(n10063) );
  NAND2_X1 U5947 ( .A1(n62921), .A2(n21701), .ZN(n11123) );
  INV_X2 U5956 ( .I(n35021), .ZN(n34553) );
  INV_X1 U5957 ( .I(n40213), .ZN(n1509) );
  BUF_X2 U5960 ( .I(n40213), .Z(n58364) );
  NAND2_X1 U5961 ( .A1(n64267), .A2(n48081), .ZN(n64880) );
  INV_X2 U5975 ( .I(n64267), .ZN(n48572) );
  NOR2_X1 U5976 ( .A1(n46771), .A2(n64267), .ZN(n48571) );
  NOR2_X1 U5989 ( .A1(n1237), .A2(n56436), .ZN(n51902) );
  NOR2_X1 U5991 ( .A1(n25404), .A2(n60579), .ZN(n32921) );
  NOR2_X1 U5993 ( .A1(n60579), .A2(n33730), .ZN(n33496) );
  NOR2_X1 U5995 ( .A1(n56455), .A2(n26162), .ZN(n56458) );
  CLKBUF_X2 U5997 ( .I(n44948), .Z(n63941) );
  NAND4_X1 U6003 ( .A1(n14568), .A2(n17319), .A3(n46823), .A4(n14567), .ZN(
        n14566) );
  INV_X1 U6006 ( .I(n46823), .ZN(n12268) );
  CLKBUF_X2 U6011 ( .I(n14773), .Z(n60113) );
  NAND3_X1 U6012 ( .A1(n30869), .A2(n30508), .A3(n31272), .ZN(n64982) );
  NOR2_X1 U6016 ( .A1(n64183), .A2(n41105), .ZN(n40438) );
  NAND3_X1 U6027 ( .A1(n11808), .A2(n10333), .A3(n61014), .ZN(n11807) );
  NOR2_X1 U6037 ( .A1(n65262), .A2(n64462), .ZN(n63594) );
  BUF_X4 U6045 ( .I(n64462), .Z(n61744) );
  INV_X2 U6047 ( .I(n6153), .ZN(n40291) );
  NOR2_X1 U6054 ( .A1(n6153), .A2(n14016), .ZN(n40223) );
  OAI22_X1 U6057 ( .A1(n1737), .A2(n39319), .B1(n64613), .B2(n6153), .ZN(
        n39321) );
  NAND2_X1 U6058 ( .A1(n17619), .A2(n28813), .ZN(n28814) );
  OAI21_X1 U6065 ( .A1(n45794), .A2(n10397), .B(n63465), .ZN(n13391) );
  CLKBUF_X2 U6070 ( .I(n10397), .Z(n58889) );
  NOR2_X1 U6074 ( .A1(n24668), .A2(n56541), .ZN(n56531) );
  INV_X1 U6078 ( .I(n46907), .ZN(n45764) );
  NAND2_X1 U6085 ( .A1(n46907), .A2(n18361), .ZN(n45513) );
  NAND3_X1 U6090 ( .A1(n56105), .A2(n9567), .A3(n56104), .ZN(n56113) );
  AOI22_X1 U6093 ( .A1(n55997), .A2(n55996), .B1(n56105), .B2(n55995), .ZN(
        n56007) );
  OAI21_X1 U6099 ( .A1(n56105), .A2(n56103), .B(n56102), .ZN(n56114) );
  NOR2_X1 U6101 ( .A1(n34350), .A2(n32922), .ZN(n32934) );
  NOR2_X1 U6106 ( .A1(n21502), .A2(n17409), .ZN(n12171) );
  NAND2_X1 U6107 ( .A1(n48155), .A2(n18099), .ZN(n47098) );
  NAND2_X1 U6108 ( .A1(n13558), .A2(n2350), .ZN(n2495) );
  NAND2_X1 U6120 ( .A1(n30841), .A2(n13558), .ZN(n16863) );
  NAND2_X1 U6122 ( .A1(n61928), .A2(n13558), .ZN(n8458) );
  INV_X2 U6123 ( .I(n49375), .ZN(n58983) );
  CLKBUF_X4 U6124 ( .I(n49375), .Z(n61741) );
  INV_X1 U6126 ( .I(n12299), .ZN(n14128) );
  NAND3_X1 U6134 ( .A1(n48722), .A2(n57182), .A3(n48721), .ZN(n48723) );
  AOI21_X1 U6135 ( .A1(n3303), .A2(n50213), .B(n50212), .ZN(n10768) );
  NAND2_X1 U6142 ( .A1(n20374), .A2(n40523), .ZN(n17971) );
  NOR2_X1 U6143 ( .A1(n39129), .A2(n20374), .ZN(n40527) );
  NAND2_X1 U6148 ( .A1(n17673), .A2(n63627), .ZN(n17677) );
  NOR2_X1 U6150 ( .A1(n54000), .A2(n53998), .ZN(n53927) );
  NAND2_X1 U6152 ( .A1(n54000), .A2(n6168), .ZN(n53983) );
  CLKBUF_X4 U6170 ( .I(n54000), .Z(n23292) );
  INV_X1 U6173 ( .I(n34359), .ZN(n32922) );
  CLKBUF_X2 U6180 ( .I(n34359), .Z(n23281) );
  NAND2_X1 U6193 ( .A1(n13940), .A2(n16487), .ZN(n16748) );
  INV_X1 U6213 ( .I(n16487), .ZN(n1453) );
  CLKBUF_X4 U6221 ( .I(n1484), .Z(n63501) );
  INV_X2 U6222 ( .I(n1484), .ZN(n45716) );
  CLKBUF_X4 U6227 ( .I(n44550), .Z(n1484) );
  BUF_X2 U6234 ( .I(n15708), .Z(n15709) );
  NOR2_X1 U6247 ( .A1(n47480), .A2(n15708), .ZN(n65005) );
  INV_X2 U6258 ( .I(n15708), .ZN(n62606) );
  NAND3_X1 U6260 ( .A1(n15032), .A2(n43328), .A3(n15033), .ZN(n62974) );
  INV_X1 U6261 ( .I(n43328), .ZN(n41486) );
  NAND2_X1 U6265 ( .A1(n12576), .A2(n42978), .ZN(n43328) );
  INV_X1 U6266 ( .I(n45191), .ZN(n1483) );
  NOR2_X1 U6274 ( .A1(n517), .A2(n45191), .ZN(n63874) );
  INV_X1 U6279 ( .I(n47470), .ZN(n2828) );
  NAND2_X1 U6283 ( .A1(n47470), .A2(n44065), .ZN(n44067) );
  NOR2_X1 U6284 ( .A1(n50045), .A2(n50041), .ZN(n49360) );
  NOR2_X1 U6288 ( .A1(n7373), .A2(n7374), .ZN(n5680) );
  NAND3_X1 U6289 ( .A1(n17818), .A2(n49721), .A3(n3031), .ZN(n62630) );
  NAND2_X1 U6290 ( .A1(n10507), .A2(n56891), .ZN(n56845) );
  AOI21_X1 U6293 ( .A1(n40990), .A2(n5362), .B(n62681), .ZN(n5393) );
  OAI21_X1 U6300 ( .A1(n49502), .A2(n49495), .B(n48391), .ZN(n47049) );
  NAND3_X1 U6306 ( .A1(n48064), .A2(n19681), .A3(n7115), .ZN(n17793) );
  NAND2_X1 U6310 ( .A1(n19681), .A2(n7113), .ZN(n8433) );
  AOI21_X1 U6312 ( .A1(n19681), .A2(n12595), .B(n48416), .ZN(n5699) );
  NOR2_X1 U6315 ( .A1(n19681), .A2(n23156), .ZN(n18625) );
  NAND2_X1 U6319 ( .A1(n55619), .A2(n62549), .ZN(n55613) );
  INV_X1 U6320 ( .I(n28800), .ZN(n27441) );
  BUF_X2 U6321 ( .I(n28800), .Z(n23773) );
  NAND2_X1 U6322 ( .A1(n64708), .A2(n34025), .ZN(n64707) );
  NOR2_X1 U6328 ( .A1(n34025), .A2(n15552), .ZN(n15551) );
  NAND3_X1 U6329 ( .A1(n36309), .A2(n2885), .A3(n36139), .ZN(n36135) );
  NAND2_X1 U6330 ( .A1(n23702), .A2(n9190), .ZN(n41715) );
  NAND2_X1 U6335 ( .A1(n42104), .A2(n23702), .ZN(n42922) );
  NAND2_X1 U6339 ( .A1(n23702), .A2(n4199), .ZN(n41713) );
  NOR2_X1 U6340 ( .A1(n4198), .A2(n23702), .ZN(n3653) );
  INV_X1 U6342 ( .I(n56812), .ZN(n56809) );
  NOR2_X1 U6343 ( .A1(n56574), .A2(n56397), .ZN(n56571) );
  INV_X1 U6346 ( .I(n56574), .ZN(n56398) );
  OAI22_X1 U6351 ( .A1(n56574), .A2(n56573), .B1(n56572), .B2(n59647), .ZN(
        n56575) );
  NOR2_X1 U6353 ( .A1(n49308), .A2(n17874), .ZN(n48999) );
  NAND2_X1 U6358 ( .A1(n17874), .A2(n49317), .ZN(n49307) );
  INV_X2 U6359 ( .I(n17874), .ZN(n11172) );
  AOI22_X1 U6360 ( .A1(n8392), .A2(n23070), .B1(n8818), .B2(n1200), .ZN(n64244) );
  OAI22_X1 U6367 ( .A1(n9505), .A2(n47580), .B1(n47281), .B2(n2973), .ZN(
        n45154) );
  NOR2_X1 U6369 ( .A1(n47579), .A2(n47580), .ZN(n47586) );
  NAND2_X1 U6377 ( .A1(n47272), .A2(n47580), .ZN(n63230) );
  NOR2_X1 U6378 ( .A1(n47580), .A2(n23186), .ZN(n47283) );
  NOR2_X1 U6382 ( .A1(n47582), .A2(n47580), .ZN(n47273) );
  NAND3_X1 U6385 ( .A1(n57195), .A2(n48236), .A3(n48234), .ZN(n14990) );
  CLKBUF_X2 U6390 ( .I(n38769), .Z(n39658) );
  INV_X2 U6391 ( .I(n49850), .ZN(n25253) );
  BUF_X2 U6394 ( .I(n49850), .Z(n22756) );
  NOR2_X1 U6395 ( .A1(n19882), .A2(n42540), .ZN(n42925) );
  NOR2_X1 U6407 ( .A1(n42540), .A2(n3674), .ZN(n42541) );
  NOR2_X1 U6408 ( .A1(n59824), .A2(n8957), .ZN(n62598) );
  NOR2_X1 U6409 ( .A1(n17304), .A2(n8957), .ZN(n35222) );
  NOR2_X1 U6413 ( .A1(n8957), .A2(n35833), .ZN(n64472) );
  INV_X1 U6421 ( .I(n8957), .ZN(n35715) );
  NOR2_X1 U6423 ( .A1(n64884), .A2(n8957), .ZN(n64883) );
  INV_X2 U6424 ( .I(n23936), .ZN(n55156) );
  BUF_X2 U6427 ( .I(n23936), .Z(n7890) );
  CLKBUF_X2 U6428 ( .I(n20899), .Z(n4651) );
  INV_X1 U6432 ( .I(n20899), .ZN(n33146) );
  INV_X1 U6441 ( .I(n20899), .ZN(n60528) );
  INV_X1 U6444 ( .I(n60826), .ZN(n4635) );
  NOR2_X1 U6445 ( .A1(n42240), .A2(n60826), .ZN(n41264) );
  CLKBUF_X2 U6451 ( .I(n14857), .Z(n14855) );
  NAND2_X1 U6459 ( .A1(n57070), .A2(n52858), .ZN(n50602) );
  NAND2_X1 U6461 ( .A1(n60498), .A2(n52858), .ZN(n52256) );
  BUF_X2 U6464 ( .I(n52858), .Z(n61516) );
  INV_X1 U6465 ( .I(n26359), .ZN(n27574) );
  BUF_X2 U6468 ( .I(n26359), .Z(n27582) );
  OAI21_X1 U6469 ( .A1(n19456), .A2(n19455), .B(n19971), .ZN(n19978) );
  AOI21_X1 U6472 ( .A1(n62724), .A2(n7146), .B(n7271), .ZN(n48442) );
  BUF_X2 U6488 ( .I(n48440), .Z(n62724) );
  INV_X1 U6489 ( .I(n38159), .ZN(n39221) );
  INV_X1 U6492 ( .I(n50230), .ZN(n17929) );
  NAND2_X1 U6498 ( .A1(n17887), .A2(n50230), .ZN(n17886) );
  BUF_X2 U6502 ( .I(n50230), .Z(n22264) );
  BUF_X2 U6503 ( .I(n22780), .Z(n4724) );
  NOR2_X1 U6506 ( .A1(n22780), .A2(n49493), .ZN(n59838) );
  NAND2_X1 U6509 ( .A1(n22780), .A2(n7738), .ZN(n49488) );
  CLKBUF_X2 U6512 ( .I(n44045), .Z(n25629) );
  CLKBUF_X4 U6513 ( .I(n57738), .Z(n65262) );
  INV_X1 U6515 ( .I(n18136), .ZN(n35024) );
  NOR2_X1 U6519 ( .A1(n36529), .A2(n36536), .ZN(n63262) );
  BUF_X4 U6521 ( .I(n36529), .Z(n18144) );
  INV_X2 U6522 ( .I(n33893), .ZN(n35735) );
  OR2_X2 U6524 ( .A1(n6686), .A2(n33116), .Z(n59125) );
  OR2_X2 U6529 ( .A1(n12480), .A2(n14080), .Z(n18077) );
  AND2_X2 U6531 ( .A1(n15807), .A2(n6530), .Z(n61699) );
  INV_X2 U6533 ( .I(n33374), .ZN(n63103) );
  AND3_X2 U6543 ( .A1(n58102), .A2(n9278), .A3(n9279), .Z(n61700) );
  INV_X8 U6546 ( .I(n7729), .ZN(n1530) );
  OR2_X2 U6547 ( .A1(n6001), .A2(n1817), .Z(n61702) );
  INV_X1 U6549 ( .I(n18130), .ZN(n18093) );
  AND2_X2 U6552 ( .A1(n13500), .A2(n63331), .Z(n61703) );
  INV_X2 U6553 ( .I(n36853), .ZN(n36847) );
  INV_X2 U6555 ( .I(n15171), .ZN(n35506) );
  AND2_X2 U6556 ( .A1(n37363), .A2(n18525), .Z(n61704) );
  INV_X4 U6558 ( .I(n22431), .ZN(n57830) );
  CLKBUF_X4 U6559 ( .I(n1528), .Z(n652) );
  NAND2_X2 U6562 ( .A1(n22936), .A2(n37090), .ZN(n59825) );
  XOR2_X1 U6563 ( .A1(n59363), .A2(n38183), .Z(n61705) );
  OR2_X1 U6569 ( .A1(n15558), .A2(n22593), .Z(n61706) );
  BUF_X4 U6573 ( .I(n23364), .Z(n17848) );
  INV_X4 U6575 ( .I(n17848), .ZN(n41665) );
  OR2_X2 U6576 ( .A1(n8368), .A2(n13462), .Z(n7237) );
  AND2_X2 U6577 ( .A1(n6689), .A2(n7175), .Z(n61708) );
  INV_X1 U6585 ( .I(n19102), .ZN(n23654) );
  INV_X2 U6593 ( .I(n41363), .ZN(n1395) );
  AND2_X1 U6611 ( .A1(n42892), .A2(n20602), .Z(n61709) );
  OR2_X2 U6613 ( .A1(n41105), .A2(n59601), .Z(n61710) );
  INV_X1 U6619 ( .I(n42019), .ZN(n43694) );
  BUF_X4 U6639 ( .I(n37913), .Z(n42019) );
  OR2_X2 U6640 ( .A1(n41242), .A2(n42681), .Z(n42151) );
  OR3_X2 U6641 ( .A1(n8215), .A2(n57557), .A3(n63747), .Z(n61711) );
  INV_X4 U6647 ( .I(n13825), .ZN(n42031) );
  INV_X4 U6660 ( .I(n62106), .ZN(n18418) );
  NOR2_X2 U6664 ( .A1(n39065), .A2(n39064), .ZN(n8538) );
  INV_X4 U6665 ( .I(n14955), .ZN(n43327) );
  INV_X4 U6667 ( .I(n46549), .ZN(n46288) );
  AND2_X1 U6676 ( .A1(n62945), .A2(n43705), .Z(n61713) );
  XOR2_X1 U6677 ( .A1(n22941), .A2(n44642), .Z(n61714) );
  INV_X2 U6678 ( .I(n16686), .ZN(n58244) );
  INV_X1 U6680 ( .I(n10624), .ZN(n10981) );
  CLKBUF_X4 U6681 ( .I(n48161), .Z(n23416) );
  INV_X1 U6683 ( .I(n18608), .ZN(n48720) );
  AND2_X1 U6684 ( .A1(n46716), .A2(n48234), .Z(n61715) );
  AND2_X2 U6685 ( .A1(n62924), .A2(n45582), .Z(n61716) );
  INV_X4 U6688 ( .I(n687), .ZN(n22157) );
  INV_X2 U6689 ( .I(n49694), .ZN(n64935) );
  OR2_X2 U6692 ( .A1(n44802), .A2(n47901), .Z(n61717) );
  NOR2_X2 U6701 ( .A1(n59967), .A2(n47874), .ZN(n47634) );
  AND2_X1 U6707 ( .A1(n18570), .A2(n48194), .Z(n61718) );
  INV_X4 U6712 ( .I(n24429), .ZN(n15386) );
  INV_X2 U6714 ( .I(n24519), .ZN(n8639) );
  INV_X2 U6717 ( .I(n59086), .ZN(n63106) );
  INV_X1 U6719 ( .I(n48944), .ZN(n50042) );
  INV_X2 U6720 ( .I(n48177), .ZN(n1659) );
  AND2_X2 U6722 ( .A1(n47421), .A2(n23666), .Z(n61720) );
  CLKBUF_X12 U6730 ( .I(n48742), .Z(n11623) );
  BUF_X4 U6733 ( .I(n44558), .Z(n14314) );
  INV_X2 U6734 ( .I(n44558), .ZN(n13839) );
  AND3_X1 U6738 ( .A1(n61867), .A2(n6130), .A3(n19379), .Z(n61721) );
  BUF_X2 U6739 ( .I(n17251), .Z(n23784) );
  INV_X2 U6742 ( .I(n54983), .ZN(n65010) );
  INV_X4 U6745 ( .I(n12702), .ZN(n15747) );
  INV_X2 U6748 ( .I(n55648), .ZN(n55631) );
  AND2_X1 U6751 ( .A1(n56359), .A2(n56554), .Z(n61724) );
  INV_X1 U6754 ( .I(n62074), .ZN(n54498) );
  AND2_X2 U6765 ( .A1(n25519), .A2(n54323), .Z(n61725) );
  CLKBUF_X8 U6769 ( .I(n19974), .Z(n15703) );
  OR2_X1 U6771 ( .A1(n55225), .A2(n16978), .Z(n61726) );
  INV_X2 U6772 ( .I(n26143), .ZN(n1325) );
  INV_X2 U6776 ( .I(n22755), .ZN(n11578) );
  INV_X4 U6782 ( .I(n138), .ZN(n25987) );
  BUF_X4 U6783 ( .I(n18582), .Z(n138) );
  AND2_X2 U6784 ( .A1(n25393), .A2(n56344), .Z(n61727) );
  CLKBUF_X4 U6794 ( .I(n53146), .Z(n20735) );
  BUF_X2 U6796 ( .I(n41444), .Z(n357) );
  NAND2_X1 U6797 ( .A1(n1219), .A2(n41444), .ZN(n40691) );
  NOR2_X2 U6800 ( .A1(n64785), .A2(n61970), .ZN(n64625) );
  NOR2_X2 U6801 ( .A1(n11871), .A2(n53857), .ZN(n53619) );
  OAI22_X2 U6806 ( .A1(n53427), .A2(n62186), .B1(n9514), .B2(n65282), .ZN(
        n11871) );
  INV_X1 U6809 ( .I(n1663), .ZN(n61527) );
  NAND2_X1 U6812 ( .A1(n6991), .A2(n52687), .ZN(n56977) );
  INV_X2 U6814 ( .I(n6991), .ZN(n56991) );
  NOR2_X1 U6815 ( .A1(n56978), .A2(n6991), .ZN(n52685) );
  NAND2_X1 U6818 ( .A1(n13960), .A2(n56103), .ZN(n56069) );
  AND2_X2 U6822 ( .A1(n43327), .A2(n15031), .Z(n16258) );
  OR2_X2 U6828 ( .A1(n14605), .A2(n15031), .Z(n15033) );
  AOI22_X1 U6831 ( .A1(n55478), .A2(n52396), .B1(n55473), .B2(n55739), .ZN(
        n60921) );
  NAND4_X1 U6837 ( .A1(n55478), .A2(n55473), .A3(n22592), .A4(n55727), .ZN(
        n52213) );
  INV_X2 U6839 ( .I(n63589), .ZN(n2177) );
  OAI21_X1 U6848 ( .A1(n30192), .A2(n30195), .B(n63589), .ZN(n62153) );
  NOR2_X1 U6849 ( .A1(n57810), .A2(n5971), .ZN(n43410) );
  INV_X1 U6852 ( .I(n5971), .ZN(n64324) );
  BUF_X4 U6858 ( .I(n25517), .Z(n2024) );
  CLKBUF_X12 U6859 ( .I(n27499), .Z(n23822) );
  NAND2_X1 U6864 ( .A1(n4226), .A2(n53428), .ZN(n62682) );
  INV_X1 U6867 ( .I(n23036), .ZN(n34200) );
  NAND2_X1 U6868 ( .A1(n23036), .A2(n34201), .ZN(n10930) );
  NOR2_X1 U6874 ( .A1(n23036), .A2(n25731), .ZN(n25730) );
  INV_X2 U6876 ( .I(n24924), .ZN(n36404) );
  NAND2_X1 U6877 ( .A1(n21591), .A2(n24924), .ZN(n36188) );
  BUF_X2 U6878 ( .I(n24924), .Z(n22474) );
  NAND2_X1 U6882 ( .A1(n35605), .A2(n11049), .ZN(n36252) );
  INV_X1 U6892 ( .I(n50254), .ZN(n22506) );
  NAND2_X1 U6897 ( .A1(n50254), .A2(n7098), .ZN(n49968) );
  NOR3_X1 U6898 ( .A1(n49310), .A2(n7005), .A3(n49614), .ZN(n7004) );
  INV_X1 U6901 ( .I(n18482), .ZN(n43695) );
  CLKBUF_X8 U6902 ( .I(n49054), .Z(n61728) );
  NOR2_X1 U6903 ( .A1(n63162), .A2(n24624), .ZN(n62737) );
  INV_X1 U6906 ( .I(n47749), .ZN(n46731) );
  NOR2_X1 U6909 ( .A1(n6170), .A2(n26113), .ZN(n64898) );
  OAI21_X1 U6918 ( .A1(n60690), .A2(n58771), .B(n2325), .ZN(n18029) );
  NAND3_X1 U6920 ( .A1(n35599), .A2(n35598), .A3(n36442), .ZN(n25355) );
  NOR2_X1 U6927 ( .A1(n23257), .A2(n36442), .ZN(n36449) );
  OAI22_X1 U6928 ( .A1(n23610), .A2(n1516), .B1(n41455), .B2(n58996), .ZN(
        n39018) );
  NAND2_X1 U6935 ( .A1(n23610), .A2(n13737), .ZN(n40680) );
  INV_X1 U6936 ( .I(n47491), .ZN(n16836) );
  NAND2_X1 U6938 ( .A1(n17630), .A2(n47372), .ZN(n46823) );
  NAND2_X1 U6942 ( .A1(n41173), .A2(n8026), .ZN(n59408) );
  NAND2_X1 U6946 ( .A1(n41173), .A2(n11787), .ZN(n40489) );
  NOR2_X1 U6955 ( .A1(n47347), .A2(n49109), .ZN(n49789) );
  INV_X1 U6956 ( .I(n23489), .ZN(n37592) );
  NOR2_X1 U6975 ( .A1(n58975), .A2(n25857), .ZN(n48840) );
  AND2_X2 U6985 ( .A1(n6808), .A2(n6810), .Z(n6809) );
  INV_X2 U6991 ( .I(n14091), .ZN(n57060) );
  NOR2_X1 U6997 ( .A1(n14091), .A2(n58326), .ZN(n58325) );
  OR2_X1 U7001 ( .A1(n14091), .A2(n25437), .Z(n61907) );
  OR3_X2 U7008 ( .A1(n33486), .A2(n16869), .A3(n18300), .Z(n9757) );
  NAND2_X1 U7012 ( .A1(n16869), .A2(n18300), .ZN(n58697) );
  CLKBUF_X12 U7020 ( .I(n22652), .Z(n59355) );
  AOI21_X2 U7021 ( .A1(n43423), .A2(n22087), .B(n60474), .ZN(n6020) );
  INV_X1 U7031 ( .I(n5140), .ZN(n6312) );
  NAND2_X1 U7041 ( .A1(n24097), .A2(n1871), .ZN(n29248) );
  NAND2_X1 U7061 ( .A1(n60293), .A2(n1871), .ZN(n29245) );
  NOR2_X1 U7066 ( .A1(n41549), .A2(n22939), .ZN(n10128) );
  INV_X1 U7072 ( .I(n41549), .ZN(n42655) );
  CLKBUF_X12 U7073 ( .I(n23114), .Z(n3112) );
  BUF_X4 U7081 ( .I(n14547), .Z(n61729) );
  CLKBUF_X12 U7096 ( .I(n56894), .Z(n23682) );
  NAND2_X1 U7100 ( .A1(n30722), .A2(n14174), .ZN(n30265) );
  INV_X1 U7105 ( .I(n14174), .ZN(n14389) );
  NOR2_X1 U7107 ( .A1(n30722), .A2(n14174), .ZN(n62437) );
  NAND2_X1 U7112 ( .A1(n14174), .A2(n30267), .ZN(n30288) );
  CLKBUF_X12 U7115 ( .I(n61164), .Z(n43917) );
  NAND2_X1 U7117 ( .A1(n6791), .A2(n23634), .ZN(n40643) );
  NAND3_X1 U7121 ( .A1(n40541), .A2(n6791), .A3(n41163), .ZN(n3642) );
  INV_X1 U7122 ( .I(n6791), .ZN(n39072) );
  NAND2_X1 U7126 ( .A1(n22380), .A2(n6791), .ZN(n59981) );
  AOI22_X1 U7132 ( .A1(n35453), .A2(n36393), .B1(n35451), .B2(n35452), .ZN(
        n62198) );
  CLKBUF_X12 U7133 ( .I(n5266), .Z(n5244) );
  INV_X4 U7135 ( .I(n24509), .ZN(n1610) );
  NOR2_X1 U7145 ( .A1(n47920), .A2(n10636), .ZN(n4908) );
  NAND2_X1 U7155 ( .A1(n47920), .A2(n10636), .ZN(n47923) );
  INV_X2 U7162 ( .I(n37411), .ZN(n36831) );
  BUF_X2 U7166 ( .I(n37411), .Z(n24041) );
  INV_X1 U7187 ( .I(n23552), .ZN(n64478) );
  BUF_X2 U7189 ( .I(n23552), .Z(n9044) );
  NAND2_X1 U7201 ( .A1(n14372), .A2(n23552), .ZN(n5078) );
  CLKBUF_X2 U7205 ( .I(n52868), .Z(n61730) );
  AND2_X2 U7207 ( .A1(n46176), .A2(n10621), .Z(n13588) );
  INV_X2 U7211 ( .I(n46176), .ZN(n48587) );
  INV_X2 U7212 ( .I(n16528), .ZN(n16527) );
  BUF_X2 U7216 ( .I(n16528), .Z(n14214) );
  CLKBUF_X12 U7221 ( .I(n16528), .Z(n7282) );
  BUF_X2 U7222 ( .I(n62507), .Z(n61731) );
  NAND2_X1 U7231 ( .A1(n10660), .A2(n33597), .ZN(n1) );
  INV_X2 U7234 ( .I(n33597), .ZN(n1540) );
  NOR2_X1 U7239 ( .A1(n33597), .A2(n11060), .ZN(n3175) );
  NOR2_X1 U7243 ( .A1(n7596), .A2(n59754), .ZN(n59753) );
  NAND2_X1 U7246 ( .A1(n24370), .A2(n37090), .ZN(n37095) );
  INV_X2 U7249 ( .I(n37090), .ZN(n37085) );
  INV_X1 U7250 ( .I(n40200), .ZN(n23932) );
  NOR2_X1 U7252 ( .A1(n40200), .A2(n22593), .ZN(n4794) );
  NAND4_X1 U7262 ( .A1(n40196), .A2(n40200), .A3(n40199), .A4(n40203), .ZN(
        n40197) );
  NOR2_X1 U7268 ( .A1(n61187), .A2(n30808), .ZN(n30531) );
  NAND2_X1 U7274 ( .A1(n61187), .A2(n10821), .ZN(n30801) );
  INV_X1 U7276 ( .I(n48676), .ZN(n9799) );
  CLKBUF_X4 U7282 ( .I(n11884), .Z(n5676) );
  NAND2_X1 U7286 ( .A1(n6273), .A2(n10544), .ZN(n27857) );
  NOR2_X1 U7287 ( .A1(n10085), .A2(n6273), .ZN(n10084) );
  INV_X1 U7294 ( .I(n6273), .ZN(n28451) );
  OR2_X2 U7304 ( .A1(n7489), .A2(n62155), .Z(n21774) );
  NOR2_X1 U7307 ( .A1(n64712), .A2(n57390), .ZN(n62516) );
  INV_X1 U7314 ( .I(n64712), .ZN(n6608) );
  CLKBUF_X4 U7327 ( .I(n33255), .Z(n35247) );
  INV_X1 U7334 ( .I(n33255), .ZN(n35241) );
  INV_X2 U7335 ( .I(n53736), .ZN(n53732) );
  NAND2_X1 U7338 ( .A1(n53736), .A2(n14845), .ZN(n53737) );
  NOR2_X1 U7339 ( .A1(n53736), .A2(n53740), .ZN(n22200) );
  CLKBUF_X12 U7344 ( .I(n51474), .Z(n23670) );
  CLKBUF_X4 U7345 ( .I(n58606), .Z(n61734) );
  CLKBUF_X12 U7346 ( .I(n23368), .Z(n61735) );
  NOR2_X1 U7349 ( .A1(n6116), .A2(n6115), .ZN(n63555) );
  NOR3_X1 U7350 ( .A1(n18806), .A2(n4389), .A3(n18808), .ZN(n60377) );
  NAND2_X1 U7352 ( .A1(n53144), .A2(n53143), .ZN(n65106) );
  NAND2_X1 U7355 ( .A1(n5087), .A2(n55364), .ZN(n14359) );
  AOI21_X1 U7359 ( .A1(n56486), .A2(n56512), .B(n56454), .ZN(n56459) );
  CLKBUF_X2 U7364 ( .I(n55882), .Z(n63830) );
  CLKBUF_X2 U7370 ( .I(n53305), .Z(n59907) );
  BUF_X2 U7374 ( .I(n56189), .Z(n19853) );
  CLKBUF_X1 U7378 ( .I(n56953), .Z(n63420) );
  BUF_X2 U7379 ( .I(n54560), .Z(n62629) );
  CLKBUF_X1 U7387 ( .I(n10507), .Z(n62800) );
  CLKBUF_X2 U7399 ( .I(n5194), .Z(n64176) );
  CLKBUF_X2 U7400 ( .I(n54727), .Z(n65124) );
  CLKBUF_X2 U7409 ( .I(n52648), .Z(n7041) );
  NAND2_X1 U7411 ( .A1(n62327), .A2(n53540), .ZN(n52749) );
  CLKBUF_X4 U7412 ( .I(n54670), .Z(n54727) );
  NAND2_X1 U7415 ( .A1(n52751), .A2(n52846), .ZN(n62161) );
  NOR3_X1 U7421 ( .A1(n7785), .A2(n65204), .A3(n7791), .ZN(n7784) );
  OAI21_X1 U7435 ( .A1(n14539), .A2(n63775), .B(n24404), .ZN(n6666) );
  AOI21_X1 U7436 ( .A1(n54500), .A2(n54499), .B(n54498), .ZN(n23139) );
  NAND2_X1 U7444 ( .A1(n53416), .A2(n53616), .ZN(n62047) );
  NAND2_X1 U7445 ( .A1(n61787), .A2(n11989), .ZN(n51270) );
  INV_X2 U7449 ( .I(n9136), .ZN(n9137) );
  NAND2_X1 U7469 ( .A1(n53178), .A2(n6351), .ZN(n53392) );
  NAND2_X1 U7480 ( .A1(n52955), .A2(n52954), .ZN(n62178) );
  NAND2_X1 U7481 ( .A1(n2466), .A2(n2468), .ZN(n8904) );
  OAI22_X1 U7483 ( .A1(n64345), .A2(n21893), .B1(n59449), .B2(n63038), .ZN(
        n64339) );
  CLKBUF_X2 U7485 ( .I(n56401), .Z(n64719) );
  CLKBUF_X1 U7491 ( .I(n6351), .Z(n63126) );
  NOR2_X1 U7495 ( .A1(n57404), .A2(n14469), .ZN(n10033) );
  NAND2_X1 U7497 ( .A1(n15820), .A2(n23360), .ZN(n51887) );
  CLKBUF_X1 U7511 ( .I(n52665), .Z(n62434) );
  INV_X2 U7518 ( .I(n21028), .ZN(n833) );
  BUF_X4 U7520 ( .I(n65281), .Z(n56229) );
  CLKBUF_X2 U7521 ( .I(n54634), .Z(n4504) );
  CLKBUF_X2 U7522 ( .I(n50683), .Z(n62818) );
  BUF_X2 U7528 ( .I(n19859), .Z(n17598) );
  OAI21_X1 U7535 ( .A1(n46849), .A2(n49618), .B(n50373), .ZN(n63136) );
  CLKBUF_X2 U7541 ( .I(n52030), .Z(n64825) );
  BUF_X4 U7542 ( .I(n5272), .Z(n4156) );
  CLKBUF_X2 U7544 ( .I(n18734), .Z(n63343) );
  AOI21_X1 U7552 ( .A1(n8432), .A2(n48418), .B(n59808), .ZN(n15879) );
  INV_X1 U7555 ( .I(n49709), .ZN(n48797) );
  NAND2_X1 U7569 ( .A1(n62088), .A2(n62087), .ZN(n62086) );
  NAND2_X1 U7570 ( .A1(n50433), .A2(n50435), .ZN(n60083) );
  NOR2_X1 U7588 ( .A1(n9322), .A2(n63493), .ZN(n63656) );
  NAND2_X1 U7589 ( .A1(n20664), .A2(n20661), .ZN(n62597) );
  NOR2_X1 U7602 ( .A1(n63082), .A2(n21892), .ZN(n13260) );
  OAI21_X1 U7605 ( .A1(n64726), .A2(n64725), .B(n48834), .ZN(n18481) );
  AOI21_X1 U7611 ( .A1(n49665), .A2(n49664), .B(n63787), .ZN(n3119) );
  NAND2_X1 U7612 ( .A1(n49661), .A2(n49662), .ZN(n63787) );
  BUF_X4 U7613 ( .I(n61673), .Z(n406) );
  INV_X1 U7624 ( .I(n50002), .ZN(n64722) );
  INV_X1 U7627 ( .I(n1376), .ZN(n64668) );
  NAND2_X1 U7628 ( .A1(n62506), .A2(n62505), .ZN(n64726) );
  OAI21_X1 U7632 ( .A1(n18158), .A2(n49145), .B(n3123), .ZN(n63915) );
  INV_X1 U7634 ( .I(n49256), .ZN(n64004) );
  AOI22_X1 U7644 ( .A1(n48771), .A2(n48774), .B1(n64488), .B2(n22457), .ZN(
        n5602) );
  NOR2_X1 U7646 ( .A1(n49576), .A2(n62033), .ZN(n62088) );
  NOR2_X1 U7649 ( .A1(n49255), .A2(n2754), .ZN(n64003) );
  AOI21_X1 U7658 ( .A1(n24821), .A2(n62744), .B(n13819), .ZN(n3846) );
  NAND2_X1 U7660 ( .A1(n16157), .A2(n49560), .ZN(n62506) );
  AND2_X1 U7663 ( .A1(n6243), .A2(n49063), .Z(n61805) );
  INV_X1 U7672 ( .I(n49551), .ZN(n49174) );
  CLKBUF_X2 U7682 ( .I(n21737), .Z(n63724) );
  AND2_X1 U7684 ( .A1(n21092), .A2(n1471), .Z(n61759) );
  INV_X1 U7685 ( .I(n48058), .ZN(n49851) );
  CLKBUF_X2 U7688 ( .I(n49729), .Z(n63238) );
  CLKBUF_X2 U7691 ( .I(n13550), .Z(n62200) );
  CLKBUF_X1 U7696 ( .I(n7328), .Z(n62358) );
  OR2_X1 U7700 ( .A1(n22819), .A2(n45160), .Z(n45171) );
  CLKBUF_X2 U7707 ( .I(n1292), .Z(n63725) );
  CLKBUF_X1 U7709 ( .I(n60726), .Z(n62139) );
  BUF_X2 U7713 ( .I(n49904), .Z(n63923) );
  CLKBUF_X2 U7716 ( .I(n22819), .Z(n19302) );
  CLKBUF_X1 U7721 ( .I(n50041), .Z(n62033) );
  INV_X2 U7723 ( .I(n46367), .ZN(n20004) );
  NAND2_X1 U7726 ( .A1(n64280), .A2(n64278), .ZN(n46904) );
  NAND2_X1 U7729 ( .A1(n47875), .A2(n47874), .ZN(n63572) );
  NOR2_X1 U7733 ( .A1(n16036), .A2(n64851), .ZN(n20544) );
  NOR3_X1 U7736 ( .A1(n48568), .A2(n48569), .A3(n48570), .ZN(n63796) );
  NAND2_X1 U7737 ( .A1(n17034), .A2(n6081), .ZN(n63107) );
  INV_X1 U7740 ( .I(n48094), .ZN(n62290) );
  NAND2_X1 U7743 ( .A1(n45592), .A2(n61860), .ZN(n62215) );
  NAND2_X1 U7745 ( .A1(n62789), .A2(n48150), .ZN(n48158) );
  AOI21_X1 U7746 ( .A1(n63652), .A2(n48558), .B(n47122), .ZN(n62307) );
  AOI21_X1 U7752 ( .A1(n10624), .A2(n62709), .B(n61819), .ZN(n62708) );
  AND2_X1 U7754 ( .A1(n1647), .A2(n47510), .Z(n61966) );
  NOR2_X1 U7756 ( .A1(n44563), .A2(n9986), .ZN(n63585) );
  INV_X1 U7763 ( .I(n48542), .ZN(n62789) );
  NAND2_X1 U7765 ( .A1(n4781), .A2(n22700), .ZN(n62522) );
  NOR2_X1 U7766 ( .A1(n47115), .A2(n62633), .ZN(n62632) );
  CLKBUF_X2 U7770 ( .I(n45900), .Z(n64447) );
  AOI21_X1 U7776 ( .A1(n15757), .A2(n48664), .B(n61963), .ZN(n12484) );
  OAI21_X1 U7778 ( .A1(n60504), .A2(n10627), .B(n2944), .ZN(n22647) );
  INV_X2 U7784 ( .I(n47469), .ZN(n61738) );
  CLKBUF_X2 U7787 ( .I(n15817), .Z(n65161) );
  CLKBUF_X4 U7788 ( .I(n45889), .Z(n48085) );
  CLKBUF_X2 U7794 ( .I(n47266), .Z(n65145) );
  OR2_X1 U7802 ( .A1(n48668), .A2(n16628), .Z(n61963) );
  CLKBUF_X2 U7817 ( .I(n47617), .Z(n64470) );
  CLKBUF_X1 U7818 ( .I(n48560), .Z(n63871) );
  CLKBUF_X2 U7835 ( .I(n58313), .Z(n63953) );
  CLKBUF_X2 U7839 ( .I(n47518), .Z(n61980) );
  BUF_X2 U7844 ( .I(n46039), .Z(n64888) );
  BUF_X2 U7851 ( .I(n15823), .Z(n64859) );
  CLKBUF_X2 U7856 ( .I(n45425), .Z(n14824) );
  BUF_X1 U7864 ( .I(n5358), .Z(n60959) );
  NAND2_X1 U7872 ( .A1(n62951), .A2(n17735), .ZN(n62950) );
  INV_X1 U7874 ( .I(n24450), .ZN(n62411) );
  NAND2_X1 U7876 ( .A1(n64787), .A2(n40870), .ZN(n44242) );
  CLKBUF_X1 U7887 ( .I(n46165), .Z(n63448) );
  INV_X1 U7890 ( .I(n22212), .ZN(n63613) );
  INV_X1 U7891 ( .I(n6588), .ZN(n63058) );
  NOR2_X1 U7893 ( .A1(n40456), .A2(n40457), .ZN(n46253) );
  CLKBUF_X2 U7894 ( .I(n62529), .Z(n62518) );
  NAND2_X1 U7897 ( .A1(n19420), .A2(n42046), .ZN(n59443) );
  CLKBUF_X2 U7899 ( .I(n60486), .Z(n62477) );
  NAND2_X1 U7901 ( .A1(n43089), .A2(n43096), .ZN(n62376) );
  NAND2_X1 U7902 ( .A1(n43235), .A2(n20183), .ZN(n65002) );
  NOR2_X1 U7904 ( .A1(n40447), .A2(n42764), .ZN(n40452) );
  NAND2_X1 U7919 ( .A1(n14363), .A2(n65084), .ZN(n43779) );
  NOR2_X1 U7921 ( .A1(n60272), .A2(n23635), .ZN(n63739) );
  NAND2_X1 U7922 ( .A1(n1690), .A2(n1332), .ZN(n15445) );
  NAND3_X1 U7924 ( .A1(n61956), .A2(n6338), .A3(n61751), .ZN(n15234) );
  INV_X1 U7930 ( .I(n41788), .ZN(n64536) );
  NOR2_X2 U7935 ( .A1(n42979), .A2(n42980), .ZN(n62313) );
  NAND2_X1 U7942 ( .A1(n64531), .A2(n64530), .ZN(n1053) );
  NAND2_X1 U7947 ( .A1(n21519), .A2(n62072), .ZN(n64284) );
  NOR2_X1 U7952 ( .A1(n39080), .A2(n57256), .ZN(n63651) );
  AOI22_X1 U7953 ( .A1(n42855), .A2(n63818), .B1(n20183), .B2(n43242), .ZN(
        n42856) );
  NAND2_X1 U7956 ( .A1(n43272), .A2(n11727), .ZN(n64535) );
  INV_X1 U7958 ( .I(n13284), .ZN(n64048) );
  NAND2_X1 U7959 ( .A1(n62963), .A2(n62962), .ZN(n62961) );
  INV_X1 U7965 ( .I(n41706), .ZN(n40431) );
  CLKBUF_X2 U7967 ( .I(n42593), .Z(n64080) );
  NAND2_X1 U7977 ( .A1(n43011), .A2(n43012), .ZN(n43013) );
  CLKBUF_X2 U7985 ( .I(n4229), .Z(n63386) );
  CLKBUF_X2 U7986 ( .I(n43890), .Z(n63818) );
  CLKBUF_X1 U7989 ( .I(n10128), .Z(n62237) );
  INV_X1 U7993 ( .I(n43123), .ZN(n63206) );
  INV_X1 U8000 ( .I(n22898), .ZN(n63945) );
  CLKBUF_X4 U8002 ( .I(n22881), .Z(n20526) );
  CLKBUF_X2 U8007 ( .I(n61237), .Z(n64653) );
  CLKBUF_X2 U8016 ( .I(n42554), .Z(n63392) );
  BUF_X4 U8018 ( .I(n4198), .Z(n64363) );
  BUF_X1 U8024 ( .I(n1705), .Z(n62346) );
  BUF_X4 U8027 ( .I(n40174), .Z(n42703) );
  CLKBUF_X8 U8031 ( .I(n17623), .Z(n61739) );
  NOR2_X1 U8035 ( .A1(n41283), .A2(n65246), .ZN(n41285) );
  OAI21_X1 U8039 ( .A1(n64896), .A2(n63807), .B(n63806), .ZN(n63805) );
  NOR2_X1 U8045 ( .A1(n64774), .A2(n12190), .ZN(n12189) );
  NAND2_X1 U8061 ( .A1(n40434), .A2(n40433), .ZN(n19274) );
  NAND2_X1 U8064 ( .A1(n40860), .A2(n15073), .ZN(n64504) );
  NOR2_X1 U8068 ( .A1(n991), .A2(n64821), .ZN(n15797) );
  NOR2_X1 U8071 ( .A1(n14343), .A2(n63919), .ZN(n3490) );
  OAI21_X1 U8072 ( .A1(n63952), .A2(n62666), .B(n2159), .ZN(n21284) );
  AOI21_X1 U8077 ( .A1(n39818), .A2(n39648), .B(n41122), .ZN(n64249) );
  NAND2_X1 U8080 ( .A1(n41380), .A2(n62228), .ZN(n13000) );
  OAI21_X1 U8083 ( .A1(n62543), .A2(n12194), .B(n41438), .ZN(n64774) );
  NAND2_X1 U8084 ( .A1(n20074), .A2(n14278), .ZN(n64821) );
  NAND2_X1 U8092 ( .A1(n18668), .A2(n18667), .ZN(n64062) );
  NOR2_X1 U8094 ( .A1(n63867), .A2(n41893), .ZN(n63531) );
  NOR2_X1 U8097 ( .A1(n42251), .A2(n41914), .ZN(n63265) );
  BUF_X2 U8098 ( .I(n20879), .Z(n64067) );
  CLKBUF_X1 U8099 ( .I(n5775), .Z(n63174) );
  NAND2_X1 U8102 ( .A1(n40680), .A2(n58798), .ZN(n58797) );
  OAI22_X1 U8106 ( .A1(n60947), .A2(n42215), .B1(n42211), .B2(n1274), .ZN(
        n42214) );
  NOR2_X1 U8107 ( .A1(n41415), .A2(n41220), .ZN(n63467) );
  OR2_X1 U8109 ( .A1(n41397), .A2(n23108), .Z(n15584) );
  CLKBUF_X2 U8115 ( .I(n12895), .Z(n62272) );
  CLKBUF_X2 U8118 ( .I(n24066), .Z(n63795) );
  CLKBUF_X2 U8123 ( .I(n37592), .Z(n62134) );
  OR2_X1 U8127 ( .A1(n40602), .A2(n40605), .Z(n38420) );
  CLKBUF_X2 U8128 ( .I(n40308), .Z(n65128) );
  CLKBUF_X1 U8129 ( .I(n20925), .Z(n65021) );
  CLKBUF_X2 U8133 ( .I(n41052), .Z(n222) );
  BUF_X1 U8140 ( .I(n41875), .Z(n62357) );
  CLKBUF_X1 U8144 ( .I(n1274), .Z(n63233) );
  CLKBUF_X2 U8145 ( .I(n40749), .Z(n62611) );
  CLKBUF_X2 U8147 ( .I(n6748), .Z(n62681) );
  BUF_X2 U8156 ( .I(n39786), .Z(n40592) );
  AND2_X2 U8161 ( .A1(n64698), .A2(n62922), .Z(n63952) );
  CLKBUF_X2 U8164 ( .I(n41059), .Z(n61008) );
  INV_X1 U8167 ( .I(n37886), .ZN(n63882) );
  CLKBUF_X2 U8169 ( .I(n14242), .Z(n9376) );
  NOR2_X1 U8171 ( .A1(n5105), .A2(n1765), .ZN(n12267) );
  CLKBUF_X2 U8173 ( .I(n38742), .Z(n64786) );
  INV_X1 U8174 ( .I(n13928), .ZN(n1763) );
  NAND2_X1 U8188 ( .A1(n21692), .A2(n7350), .ZN(n21691) );
  NOR2_X1 U8189 ( .A1(n63771), .A2(n36671), .ZN(n63770) );
  NOR2_X1 U8190 ( .A1(n36187), .A2(n36186), .ZN(n13078) );
  NAND4_X1 U8196 ( .A1(n37431), .A2(n37429), .A3(n37432), .A4(n37430), .ZN(
        n63810) );
  NOR3_X1 U8197 ( .A1(n61919), .A2(n35500), .A3(n60356), .ZN(n64988) );
  AOI22_X1 U8198 ( .A1(n34875), .A2(n62333), .B1(n35883), .B2(n64198), .ZN(
        n17385) );
  INV_X1 U8203 ( .I(n37008), .ZN(n63645) );
  NAND2_X1 U8204 ( .A1(n37422), .A2(n37423), .ZN(n37431) );
  NAND2_X1 U8211 ( .A1(n36373), .A2(n36374), .ZN(n64425) );
  AOI21_X1 U8212 ( .A1(n19699), .A2(n35546), .B(n15070), .ZN(n62948) );
  AOI22_X1 U8220 ( .A1(n36949), .A2(n36950), .B1(n36947), .B2(n36948), .ZN(
        n11757) );
  NAND2_X1 U8224 ( .A1(n37327), .A2(n37328), .ZN(n65140) );
  INV_X1 U8234 ( .I(n33716), .ZN(n65178) );
  AOI21_X1 U8236 ( .A1(n35433), .A2(n36945), .B(n23944), .ZN(n63088) );
  AND3_X1 U8238 ( .A1(n63638), .A2(n36639), .A3(n37085), .Z(n61887) );
  AOI21_X1 U8241 ( .A1(n36456), .A2(n61940), .B(n15034), .ZN(n7245) );
  BUF_X1 U8243 ( .I(n35396), .Z(n63848) );
  OR2_X1 U8257 ( .A1(n23626), .A2(n36021), .Z(n61784) );
  BUF_X2 U8259 ( .I(n7208), .Z(n62920) );
  AND2_X1 U8262 ( .A1(n7208), .A2(n4754), .Z(n61919) );
  CLKBUF_X4 U8263 ( .I(n6682), .Z(n4969) );
  BUF_X4 U8268 ( .I(n24228), .Z(n9456) );
  OR2_X1 U8272 ( .A1(n36115), .A2(n35363), .Z(n61936) );
  OAI21_X1 U8275 ( .A1(n61701), .A2(n32878), .B(n34187), .ZN(n62447) );
  INV_X1 U8280 ( .I(n35839), .ZN(n64626) );
  AOI21_X1 U8288 ( .A1(n34192), .A2(n15099), .B(n63553), .ZN(n10853) );
  NAND3_X1 U8293 ( .A1(n35719), .A2(n35718), .A3(n35717), .ZN(n61996) );
  NAND2_X1 U8294 ( .A1(n34283), .A2(n34285), .ZN(n63996) );
  NOR2_X1 U8300 ( .A1(n63494), .A2(n34037), .ZN(n34050) );
  OAI21_X1 U8302 ( .A1(n35751), .A2(n35752), .B(n35750), .ZN(n62460) );
  NAND2_X1 U8312 ( .A1(n35730), .A2(n10608), .ZN(n35733) );
  NAND2_X1 U8317 ( .A1(n7017), .A2(n60684), .ZN(n64748) );
  NAND2_X1 U8318 ( .A1(n63103), .A2(n33537), .ZN(n63625) );
  NOR2_X1 U8330 ( .A1(n23223), .A2(n2346), .ZN(n34590) );
  CLKBUF_X1 U8333 ( .I(n20865), .Z(n63329) );
  NAND2_X1 U8338 ( .A1(n33489), .A2(n63319), .ZN(n63318) );
  BUF_X2 U8339 ( .I(n33534), .Z(n60434) );
  CLKBUF_X2 U8340 ( .I(n33780), .Z(n10175) );
  OR2_X1 U8345 ( .A1(n18878), .A2(n6914), .Z(n61934) );
  CLKBUF_X2 U8347 ( .I(n24737), .Z(n63305) );
  CLKBUF_X2 U8350 ( .I(n14464), .Z(n64958) );
  CLKBUF_X2 U8354 ( .I(n60883), .Z(n64158) );
  BUF_X2 U8363 ( .I(n4405), .Z(n62045) );
  INV_X4 U8371 ( .I(n9601), .ZN(n64603) );
  BUF_X2 U8383 ( .I(n35629), .Z(n7342) );
  CLKBUF_X1 U8393 ( .I(n12586), .Z(n32545) );
  CLKBUF_X2 U8395 ( .I(n30401), .Z(n65197) );
  NAND3_X1 U8398 ( .A1(n29761), .A2(n29760), .A3(n62747), .ZN(n62746) );
  NAND3_X1 U8399 ( .A1(n62695), .A2(n29598), .A3(n29597), .ZN(n16759) );
  OAI22_X1 U8404 ( .A1(n13629), .A2(n61390), .B1(n30362), .B2(n29431), .ZN(
        n62036) );
  NAND2_X1 U8407 ( .A1(n29928), .A2(n29936), .ZN(n63447) );
  OAI21_X1 U8410 ( .A1(n18101), .A2(n18102), .B(n58052), .ZN(n62721) );
  OAI21_X1 U8418 ( .A1(n64238), .A2(n59046), .B(n30755), .ZN(n64237) );
  NAND2_X1 U8432 ( .A1(n30479), .A2(n30478), .ZN(n65190) );
  NOR2_X1 U8436 ( .A1(n8458), .A2(n7040), .ZN(n63689) );
  NAND3_X1 U8447 ( .A1(n61849), .A2(n9654), .A3(n1435), .ZN(n30505) );
  INV_X2 U8448 ( .I(n25707), .ZN(n1431) );
  AND2_X1 U8449 ( .A1(n29904), .A2(n63394), .Z(n61777) );
  BUF_X4 U8454 ( .I(n31189), .Z(n24777) );
  NOR2_X1 U8456 ( .A1(n24556), .A2(n63394), .ZN(n62479) );
  BUF_X2 U8460 ( .I(n31098), .Z(n64128) );
  CLKBUF_X1 U8468 ( .I(n63355), .Z(n63272) );
  CLKBUF_X1 U8478 ( .I(n64169), .Z(n62053) );
  CLKBUF_X2 U8479 ( .I(n23094), .Z(n64154) );
  AOI22_X1 U8497 ( .A1(n2176), .A2(n27061), .B1(n60993), .B2(n61021), .ZN(
        n27062) );
  CLKBUF_X1 U8504 ( .I(n18213), .Z(n65039) );
  CLKBUF_X1 U8510 ( .I(n37691), .Z(n64355) );
  NAND2_X1 U8517 ( .A1(n23822), .A2(n19452), .ZN(n63797) );
  CLKBUF_X2 U8519 ( .I(n28534), .Z(n7354) );
  NAND2_X1 U8537 ( .A1(n22721), .A2(n27665), .ZN(n62271) );
  CLKBUF_X2 U8547 ( .I(n26824), .Z(n63094) );
  CLKBUF_X2 U8553 ( .I(n29171), .Z(n62005) );
  CLKBUF_X2 U8559 ( .I(Key[131]), .Z(n63396) );
  AOI21_X1 U8560 ( .A1(n12322), .A2(n12320), .B(n63457), .ZN(n12318) );
  NAND3_X1 U8566 ( .A1(n22280), .A2(n22279), .A3(n50816), .ZN(n64560) );
  NAND3_X1 U8568 ( .A1(n60377), .A2(n65169), .A3(n18803), .ZN(n63282) );
  NAND3_X1 U8571 ( .A1(n64365), .A2(n56493), .A3(n56494), .ZN(n19177) );
  NAND3_X1 U8573 ( .A1(n59599), .A2(n56943), .A3(n64845), .ZN(n56944) );
  NOR2_X1 U8579 ( .A1(n64656), .A2(n53132), .ZN(n12210) );
  NAND3_X1 U8580 ( .A1(n64743), .A2(n23088), .A3(n55195), .ZN(n23087) );
  NAND2_X1 U8586 ( .A1(n4645), .A2(n4644), .ZN(n53153) );
  NAND4_X1 U8594 ( .A1(n54167), .A2(n54166), .A3(n54165), .A4(n57222), .ZN(
        n54169) );
  NAND3_X1 U8596 ( .A1(n56964), .A2(n56908), .A3(n14708), .ZN(n56904) );
  NOR2_X1 U8604 ( .A1(n54235), .A2(n19884), .ZN(n21286) );
  NOR3_X1 U8605 ( .A1(n19376), .A2(n58444), .A3(n57334), .ZN(n61174) );
  AOI22_X1 U8613 ( .A1(n55181), .A2(n55210), .B1(n55182), .B2(n55234), .ZN(
        n63711) );
  NOR2_X1 U8626 ( .A1(n2372), .A2(n2371), .ZN(n17652) );
  NAND2_X1 U8628 ( .A1(n53167), .A2(n52231), .ZN(n59372) );
  NAND2_X1 U8634 ( .A1(n54769), .A2(n54669), .ZN(n57967) );
  INV_X1 U8644 ( .I(n64872), .ZN(n56838) );
  AOI21_X1 U8646 ( .A1(n21210), .A2(n14428), .B(n64598), .ZN(n4559) );
  CLKBUF_X4 U8648 ( .I(n18652), .Z(n14643) );
  INV_X1 U8652 ( .I(n56667), .ZN(n63858) );
  BUF_X2 U8655 ( .I(n62578), .Z(n61057) );
  INV_X1 U8674 ( .I(n18786), .ZN(n63822) );
  CLKBUF_X2 U8676 ( .I(n56886), .Z(n1255) );
  CLKBUF_X2 U8678 ( .I(n54272), .Z(n23731) );
  CLKBUF_X4 U8682 ( .I(n56522), .Z(n23920) );
  BUF_X4 U8690 ( .I(n53483), .Z(n23611) );
  NAND2_X1 U8692 ( .A1(n13902), .A2(n17455), .ZN(n13901) );
  NAND2_X1 U8694 ( .A1(n56281), .A2(n10389), .ZN(n64652) );
  AOI22_X1 U8696 ( .A1(n63580), .A2(n57002), .B1(n53239), .B2(n50548), .ZN(
        n5615) );
  NOR2_X1 U8698 ( .A1(n62077), .A2(n62076), .ZN(n62075) );
  NAND2_X1 U8703 ( .A1(n62161), .A2(n25894), .ZN(n61630) );
  NAND2_X1 U8707 ( .A1(n14376), .A2(n14374), .ZN(n2925) );
  BUF_X4 U8714 ( .I(n56107), .Z(n61740) );
  BUF_X4 U8722 ( .I(n56717), .Z(n23785) );
  BUF_X2 U8726 ( .I(n55868), .Z(n22681) );
  OAI22_X1 U8727 ( .A1(n61931), .A2(n61871), .B1(n52246), .B2(n52245), .ZN(
        n63786) );
  NOR2_X1 U8741 ( .A1(n53395), .A2(n22708), .ZN(n62076) );
  INV_X1 U8754 ( .I(n56130), .ZN(n63550) );
  NAND2_X1 U8759 ( .A1(n64741), .A2(n64740), .ZN(n62723) );
  NOR3_X1 U8766 ( .A1(n25718), .A2(n52119), .A3(n25719), .ZN(n62840) );
  NAND2_X1 U8771 ( .A1(n53454), .A2(n63481), .ZN(n53459) );
  NOR2_X1 U8773 ( .A1(n59387), .A2(n64739), .ZN(n13795) );
  NOR2_X1 U8775 ( .A1(n60814), .A2(n54619), .ZN(n21837) );
  INV_X1 U8777 ( .I(n53392), .ZN(n53179) );
  NOR3_X1 U8778 ( .A1(n53855), .A2(n53857), .A3(n53856), .ZN(n62211) );
  AND3_X1 U8785 ( .A1(n57057), .A2(n57058), .A3(n57067), .Z(n61767) );
  OAI21_X1 U8800 ( .A1(n57029), .A2(n1152), .B(n64586), .ZN(n21573) );
  NAND2_X1 U8805 ( .A1(n57007), .A2(n6608), .ZN(n63988) );
  NAND2_X1 U8807 ( .A1(n53872), .A2(n13601), .ZN(n64991) );
  AOI21_X1 U8809 ( .A1(n54309), .A2(n54308), .B(n60794), .ZN(n64596) );
  AOI21_X1 U8812 ( .A1(n64342), .A2(n52667), .B(n62434), .ZN(n52680) );
  NOR2_X1 U8817 ( .A1(n63126), .A2(n53534), .ZN(n62741) );
  AND2_X1 U8818 ( .A1(n52708), .A2(n21330), .Z(n61931) );
  OAI21_X1 U8819 ( .A1(n56997), .A2(n61572), .B(n23110), .ZN(n20200) );
  INV_X1 U8822 ( .I(n4078), .ZN(n52772) );
  NOR2_X1 U8824 ( .A1(n16620), .A2(n51901), .ZN(n64453) );
  NOR3_X1 U8830 ( .A1(n14325), .A2(n51895), .A3(n62752), .ZN(n60578) );
  NAND2_X1 U8836 ( .A1(n55263), .A2(n55264), .ZN(n62979) );
  NAND2_X1 U8840 ( .A1(n56212), .A2(n56213), .ZN(n22382) );
  NAND2_X1 U8847 ( .A1(n24526), .A2(n55276), .ZN(n62980) );
  NOR2_X1 U8848 ( .A1(n16384), .A2(n12695), .ZN(n64740) );
  INV_X1 U8849 ( .I(n56580), .ZN(n64189) );
  NAND2_X1 U8853 ( .A1(n1605), .A2(n53589), .ZN(n52769) );
  NAND2_X1 U8856 ( .A1(n63361), .A2(n63360), .ZN(n63359) );
  NAND2_X1 U8859 ( .A1(n64339), .A2(n51110), .ZN(n60127) );
  CLKBUF_X2 U8867 ( .I(n54346), .Z(n64608) );
  CLKBUF_X2 U8871 ( .I(n52668), .Z(n63743) );
  NAND3_X1 U8879 ( .A1(n55953), .A2(n55952), .A3(n55951), .ZN(n64190) );
  CLKBUF_X2 U8880 ( .I(n53871), .Z(n63679) );
  NOR2_X1 U8890 ( .A1(n53440), .A2(n23248), .ZN(n64772) );
  NAND2_X1 U8900 ( .A1(n56977), .A2(n64030), .ZN(n56979) );
  CLKBUF_X2 U8902 ( .I(n5277), .Z(n64255) );
  INV_X1 U8904 ( .I(n24404), .ZN(n62752) );
  NOR2_X1 U8905 ( .A1(n56256), .A2(n23952), .ZN(n56590) );
  OR2_X1 U8907 ( .A1(n15281), .A2(n54949), .Z(n23309) );
  BUF_X4 U8908 ( .I(n55474), .Z(n22592) );
  CLKBUF_X2 U8912 ( .I(n20737), .Z(n65175) );
  CLKBUF_X2 U8918 ( .I(n54594), .Z(n64129) );
  CLKBUF_X2 U8920 ( .I(n56215), .Z(n64345) );
  CLKBUF_X2 U8923 ( .I(n16797), .Z(n64832) );
  CLKBUF_X2 U8925 ( .I(n14178), .Z(n62186) );
  BUF_X4 U8934 ( .I(n51344), .Z(n56539) );
  BUF_X4 U8936 ( .I(n52091), .Z(n55440) );
  BUF_X2 U8942 ( .I(n51962), .Z(n55690) );
  CLKBUF_X1 U8953 ( .I(n25149), .Z(n63002) );
  INV_X1 U8955 ( .I(n52146), .ZN(n62475) );
  CLKBUF_X2 U8961 ( .I(n52458), .Z(n64454) );
  CLKBUF_X2 U8963 ( .I(n25618), .Z(n63690) );
  OAI21_X1 U8966 ( .A1(n48002), .A2(n12330), .B(n15709), .ZN(n62876) );
  INV_X1 U8968 ( .I(n24079), .ZN(n63424) );
  BUF_X2 U8972 ( .I(n24005), .Z(n9854) );
  NAND2_X1 U8973 ( .A1(n13923), .A2(n62531), .ZN(n8713) );
  NAND2_X1 U8987 ( .A1(n47460), .A2(n58980), .ZN(n20211) );
  BUF_X4 U8993 ( .I(n51804), .Z(n3741) );
  NOR2_X1 U9004 ( .A1(n63760), .A2(n49765), .ZN(n8675) );
  NAND2_X1 U9006 ( .A1(n63737), .A2(n20935), .ZN(n14975) );
  NAND2_X1 U9011 ( .A1(n18432), .A2(n9233), .ZN(n9232) );
  AOI22_X1 U9020 ( .A1(n393), .A2(n62861), .B1(n60732), .B2(n60734), .ZN(
        n49084) );
  OAI21_X1 U9023 ( .A1(n49042), .A2(n49041), .B(n62630), .ZN(n49045) );
  NOR2_X1 U9030 ( .A1(n12557), .A2(n49268), .ZN(n65030) );
  NAND2_X1 U9045 ( .A1(n25541), .A2(n49952), .ZN(n63061) );
  OAI21_X1 U9046 ( .A1(n13319), .A2(n64170), .B(n13316), .ZN(n64533) );
  NAND2_X1 U9058 ( .A1(n49574), .A2(n49573), .ZN(n62561) );
  NAND3_X1 U9065 ( .A1(n49924), .A2(n60772), .A3(n61808), .ZN(n47336) );
  AOI21_X1 U9085 ( .A1(n61773), .A2(n57878), .B(n63073), .ZN(n62302) );
  NAND2_X1 U9087 ( .A1(n45166), .A2(n49755), .ZN(n64143) );
  NOR3_X1 U9097 ( .A1(n49608), .A2(n63852), .A3(n64256), .ZN(n7002) );
  NAND2_X1 U9098 ( .A1(n64862), .A2(n49766), .ZN(n63760) );
  AOI22_X1 U9104 ( .A1(n47991), .A2(n17086), .B1(n16047), .B2(n63664), .ZN(
        n64803) );
  NAND2_X1 U9114 ( .A1(n23245), .A2(n50255), .ZN(n63180) );
  NAND2_X1 U9120 ( .A1(n50260), .A2(n50259), .ZN(n63182) );
  NAND2_X1 U9134 ( .A1(n64004), .A2(n64003), .ZN(n64002) );
  INV_X1 U9137 ( .I(n63621), .ZN(n57265) );
  NAND2_X1 U9142 ( .A1(n63915), .A2(n49147), .ZN(n22930) );
  NAND2_X1 U9143 ( .A1(n5602), .A2(n24906), .ZN(n63868) );
  INV_X1 U9147 ( .I(n49477), .ZN(n64723) );
  NAND2_X1 U9149 ( .A1(n48333), .A2(n62174), .ZN(n62173) );
  NAND2_X1 U9158 ( .A1(n64206), .A2(n57474), .ZN(n58204) );
  INV_X1 U9160 ( .I(n48298), .ZN(n63073) );
  INV_X1 U9175 ( .I(n49613), .ZN(n64926) );
  INV_X1 U9178 ( .I(n14353), .ZN(n61488) );
  NAND3_X1 U9179 ( .A1(n47785), .A2(n49914), .A3(n48734), .ZN(n47786) );
  NOR2_X1 U9184 ( .A1(n44795), .A2(n44794), .ZN(n62618) );
  NAND2_X1 U9187 ( .A1(n48059), .A2(n62927), .ZN(n59101) );
  OR2_X1 U9188 ( .A1(n20460), .A2(n49077), .Z(n64053) );
  NAND2_X1 U9192 ( .A1(n49499), .A2(n6704), .ZN(n64545) );
  INV_X1 U9212 ( .I(n49772), .ZN(n64108) );
  INV_X1 U9217 ( .I(n50053), .ZN(n62610) );
  INV_X2 U9224 ( .I(n49598), .ZN(n49308) );
  CLKBUF_X2 U9227 ( .I(n16963), .Z(n63186) );
  CLKBUF_X1 U9232 ( .I(n50257), .Z(n62538) );
  CLKBUF_X4 U9233 ( .I(n49076), .Z(n1468) );
  CLKBUF_X4 U9237 ( .I(n23532), .Z(n65135) );
  INV_X2 U9238 ( .I(n49277), .ZN(n49286) );
  BUF_X4 U9245 ( .I(n44569), .Z(n49908) );
  NOR2_X1 U9246 ( .A1(n16876), .A2(n16878), .ZN(n63108) );
  NOR2_X1 U9249 ( .A1(n63831), .A2(n49918), .ZN(n63610) );
  NOR2_X1 U9253 ( .A1(n17770), .A2(n12698), .ZN(n64196) );
  NAND2_X2 U9254 ( .A1(n21622), .A2(n21621), .ZN(n62700) );
  NOR2_X1 U9260 ( .A1(n61211), .A2(n60939), .ZN(n62496) );
  NAND2_X1 U9277 ( .A1(n3598), .A2(n64220), .ZN(n64219) );
  AOI21_X1 U9286 ( .A1(n57344), .A2(n23676), .B(n57333), .ZN(n64765) );
  CLKBUF_X8 U9287 ( .I(n48428), .Z(n61742) );
  NAND2_X1 U9292 ( .A1(n6288), .A2(n6285), .ZN(n6284) );
  CLKBUF_X2 U9295 ( .I(n18364), .Z(n64135) );
  NAND3_X1 U9300 ( .A1(n47005), .A2(n47006), .A3(n47004), .ZN(n47008) );
  NAND2_X1 U9307 ( .A1(n17206), .A2(n63057), .ZN(n57970) );
  NAND2_X1 U9317 ( .A1(n63572), .A2(n63571), .ZN(n57963) );
  AOI22_X1 U9318 ( .A1(n62215), .A2(n45594), .B1(n47904), .B2(n59959), .ZN(
        n57654) );
  INV_X1 U9319 ( .I(n62307), .ZN(n13350) );
  NAND2_X1 U9322 ( .A1(n6432), .A2(n46055), .ZN(n65103) );
  NAND2_X1 U9323 ( .A1(n47005), .A2(n61815), .ZN(n57344) );
  NAND2_X1 U9324 ( .A1(n62165), .A2(n64997), .ZN(n21978) );
  NAND2_X1 U9326 ( .A1(n14366), .A2(n47016), .ZN(n62082) );
  NAND3_X1 U9330 ( .A1(n61212), .A2(n47529), .A3(n8820), .ZN(n47007) );
  NAND2_X1 U9333 ( .A1(n46081), .A2(n46080), .ZN(n64997) );
  NAND2_X1 U9335 ( .A1(n62300), .A2(n48662), .ZN(n1083) );
  NAND2_X1 U9336 ( .A1(n45552), .A2(n63338), .ZN(n63824) );
  OAI21_X1 U9339 ( .A1(n47118), .A2(n10329), .B(n10328), .ZN(n47131) );
  NOR2_X1 U9349 ( .A1(n47892), .A2(n47634), .ZN(n63571) );
  AOI21_X1 U9350 ( .A1(n47437), .A2(n47436), .B(n62570), .ZN(n5373) );
  NAND2_X1 U9358 ( .A1(n45910), .A2(n45911), .ZN(n62523) );
  INV_X1 U9364 ( .I(n46037), .ZN(n64168) );
  NAND2_X1 U9368 ( .A1(n47025), .A2(n44570), .ZN(n22871) );
  NAND2_X1 U9380 ( .A1(n8603), .A2(n45222), .ZN(n64330) );
  NOR2_X1 U9381 ( .A1(n46104), .A2(n62301), .ZN(n62300) );
  NAND2_X1 U9388 ( .A1(n62632), .A2(n23850), .ZN(n57463) );
  AND3_X1 U9393 ( .A1(n64779), .A2(n48552), .A3(n59160), .Z(n61764) );
  AOI21_X1 U9395 ( .A1(n9175), .A2(n9176), .B(n61738), .ZN(n57399) );
  NAND2_X1 U9397 ( .A1(n64576), .A2(n47439), .ZN(n62570) );
  NOR2_X1 U9398 ( .A1(n44705), .A2(n18321), .ZN(n63171) );
  CLKBUF_X2 U9400 ( .I(n45972), .Z(n62748) );
  OAI21_X1 U9401 ( .A1(n61527), .A2(n47236), .B(n1069), .ZN(n8651) );
  AND2_X1 U9402 ( .A1(n4660), .A2(n26032), .Z(n61863) );
  NOR2_X1 U9403 ( .A1(n44647), .A2(n46944), .ZN(n64441) );
  BUF_X2 U9409 ( .I(n47312), .Z(n63700) );
  CLKBUF_X2 U9422 ( .I(n64250), .Z(n63670) );
  INV_X1 U9426 ( .I(n18127), .ZN(n64800) );
  NOR2_X1 U9435 ( .A1(n2743), .A2(n65062), .ZN(n63403) );
  NAND2_X1 U9437 ( .A1(n48474), .A2(n48475), .ZN(n63916) );
  INV_X1 U9446 ( .I(n44860), .ZN(n64584) );
  BUF_X1 U9447 ( .I(n16742), .Z(n61582) );
  INV_X2 U9450 ( .I(n61191), .ZN(n48252) );
  CLKBUF_X2 U9454 ( .I(n47465), .Z(n64061) );
  AND3_X1 U9464 ( .A1(n48080), .A2(n48085), .A3(n24113), .Z(n61819) );
  INV_X1 U9468 ( .I(n62230), .ZN(n63232) );
  BUF_X2 U9472 ( .I(n22852), .Z(n59922) );
  AND2_X1 U9477 ( .A1(n23263), .A2(n7335), .Z(n61861) );
  AND2_X1 U9480 ( .A1(n45908), .A2(n46731), .Z(n4781) );
  INV_X1 U9488 ( .I(n48162), .ZN(n48163) );
  AND2_X1 U9495 ( .A1(n6730), .A2(n24893), .Z(n61830) );
  CLKBUF_X2 U9496 ( .I(n62978), .Z(n62366) );
  CLKBUF_X2 U9500 ( .I(n46927), .Z(n63294) );
  CLKBUF_X2 U9505 ( .I(n45746), .Z(n63098) );
  CLKBUF_X2 U9510 ( .I(n1486), .Z(n64096) );
  AND2_X1 U9517 ( .A1(n9860), .A2(n47830), .Z(n61885) );
  BUF_X4 U9522 ( .I(n47868), .Z(n70) );
  CLKBUF_X2 U9525 ( .I(n23759), .Z(n64654) );
  BUF_X2 U9530 ( .I(n47367), .Z(n62501) );
  CLKBUF_X2 U9533 ( .I(n25702), .Z(n63338) );
  CLKBUF_X2 U9536 ( .I(n47680), .Z(n63465) );
  CLKBUF_X2 U9537 ( .I(n14448), .Z(n62490) );
  CLKBUF_X2 U9542 ( .I(n20091), .Z(n62115) );
  BUF_X2 U9543 ( .I(n22772), .Z(n548) );
  CLKBUF_X2 U9547 ( .I(n47181), .Z(n65059) );
  CLKBUF_X2 U9549 ( .I(n47034), .Z(n64063) );
  CLKBUF_X2 U9552 ( .I(n47830), .Z(n62952) );
  BUF_X2 U9553 ( .I(n23405), .Z(n64944) );
  CLKBUF_X4 U9561 ( .I(n46912), .Z(n23480) );
  INV_X1 U9575 ( .I(n21027), .ZN(n63308) );
  BUF_X2 U9578 ( .I(n23089), .Z(n22199) );
  INV_X1 U9587 ( .I(n45117), .ZN(n65003) );
  CLKBUF_X2 U9591 ( .I(n65273), .Z(n62646) );
  CLKBUF_X1 U9613 ( .I(n9628), .Z(n64512) );
  BUF_X2 U9619 ( .I(n4686), .Z(n20919) );
  CLKBUF_X2 U9620 ( .I(n46688), .Z(n64258) );
  CLKBUF_X2 U9628 ( .I(n46187), .Z(n65144) );
  CLKBUF_X2 U9642 ( .I(n46538), .Z(n64971) );
  NOR2_X1 U9645 ( .A1(n9941), .A2(n16547), .ZN(n16555) );
  NOR2_X1 U9648 ( .A1(n65122), .A2(n19047), .ZN(n1010) );
  NOR2_X1 U9650 ( .A1(n6971), .A2(n62137), .ZN(n58674) );
  NAND2_X1 U9662 ( .A1(n63341), .A2(n15658), .ZN(n65122) );
  NOR2_X1 U9682 ( .A1(n64886), .A2(n18576), .ZN(n63283) );
  CLKBUF_X2 U9690 ( .I(n44912), .Z(n65022) );
  NOR2_X1 U9699 ( .A1(n43329), .A2(n62974), .ZN(n14658) );
  NOR2_X1 U9703 ( .A1(n64688), .A2(n19718), .ZN(n19717) );
  AOI21_X1 U9704 ( .A1(n42615), .A2(n8788), .B(n63206), .ZN(n63222) );
  OAI22_X1 U9709 ( .A1(n59767), .A2(n63651), .B1(n39083), .B2(n39084), .ZN(
        n14060) );
  NOR2_X1 U9716 ( .A1(n4519), .A2(n20293), .ZN(n21753) );
  OAI21_X1 U9723 ( .A1(n42844), .A2(n1008), .B(n7435), .ZN(n62879) );
  NOR2_X1 U9724 ( .A1(n62971), .A2(n62970), .ZN(n5326) );
  NAND2_X1 U9730 ( .A1(n62058), .A2(n42424), .ZN(n3009) );
  BUF_X1 U9731 ( .I(n43100), .Z(n62297) );
  NOR2_X1 U9743 ( .A1(n41758), .A2(n42065), .ZN(n62439) );
  NAND2_X1 U9752 ( .A1(n62537), .A2(n62536), .ZN(n43676) );
  NOR2_X1 U9783 ( .A1(n43994), .A2(n17428), .ZN(n18460) );
  NOR2_X1 U9790 ( .A1(n43396), .A2(n43690), .ZN(n63479) );
  NAND2_X1 U9800 ( .A1(n64536), .A2(n64535), .ZN(n57447) );
  NOR2_X1 U9801 ( .A1(n42352), .A2(n42353), .ZN(n6162) );
  NAND2_X1 U9808 ( .A1(n63466), .A2(n14700), .ZN(n14699) );
  INV_X1 U9820 ( .I(n12972), .ZN(n43614) );
  OAI21_X1 U9821 ( .A1(n1938), .A2(n12091), .B(n63397), .ZN(n1936) );
  NAND2_X1 U9822 ( .A1(n43611), .A2(n12972), .ZN(n12971) );
  NOR2_X1 U9823 ( .A1(n12642), .A2(n19843), .ZN(n62971) );
  NOR2_X1 U9826 ( .A1(n65086), .A2(n65085), .ZN(n65084) );
  NOR2_X1 U9830 ( .A1(n64048), .A2(n42044), .ZN(n41764) );
  NAND2_X1 U9833 ( .A1(n63778), .A2(n63777), .ZN(n59156) );
  AOI21_X1 U9836 ( .A1(n2580), .A2(n42614), .B(n42613), .ZN(n63270) );
  INV_X1 U9838 ( .I(n43391), .ZN(n16997) );
  NAND2_X1 U9844 ( .A1(n42702), .A2(n42701), .ZN(n62303) );
  NAND2_X1 U9856 ( .A1(n18958), .A2(n43023), .ZN(n42779) );
  INV_X1 U9859 ( .I(n43631), .ZN(n62537) );
  NAND2_X1 U9864 ( .A1(n42100), .A2(n63506), .ZN(n5315) );
  BUF_X2 U9873 ( .I(n20942), .Z(n62461) );
  INV_X1 U9874 ( .I(n24576), .ZN(n64530) );
  INV_X1 U9876 ( .I(n43842), .ZN(n63792) );
  AND2_X1 U9881 ( .A1(n42915), .A2(n38613), .Z(n61956) );
  NAND2_X1 U9884 ( .A1(n42110), .A2(n42111), .ZN(n64792) );
  INV_X1 U9891 ( .I(n42188), .ZN(n1689) );
  NAND2_X2 U9892 ( .A1(n15020), .A2(n20844), .ZN(n16378) );
  CLKBUF_X2 U9893 ( .I(n2121), .Z(n64724) );
  NAND2_X1 U9894 ( .A1(n57255), .A2(n279), .ZN(n65086) );
  NAND2_X1 U9897 ( .A1(n16258), .A2(n61858), .ZN(n63774) );
  AOI21_X1 U9907 ( .A1(n65217), .A2(n43122), .B(n43268), .ZN(n43126) );
  CLKBUF_X2 U9911 ( .I(n23557), .Z(n63455) );
  OR2_X1 U9913 ( .A1(n3653), .A2(n41604), .Z(n3652) );
  NOR2_X1 U9914 ( .A1(n42585), .A2(n63945), .ZN(n63944) );
  BUF_X2 U9915 ( .I(n43852), .Z(n60706) );
  CLKBUF_X2 U9918 ( .I(n22716), .Z(n62462) );
  INV_X1 U9920 ( .I(n38684), .ZN(n42912) );
  BUF_X1 U9923 ( .I(n25534), .Z(n64492) );
  NOR2_X1 U9934 ( .A1(n63965), .A2(n64992), .ZN(n61973) );
  INV_X2 U9939 ( .I(n42049), .ZN(n43448) );
  NOR2_X1 U9940 ( .A1(n15340), .A2(n64253), .ZN(n8921) );
  INV_X1 U9943 ( .I(n63805), .ZN(n20584) );
  AOI21_X1 U9949 ( .A1(n1979), .A2(n1982), .B(n62423), .ZN(n62436) );
  BUF_X4 U9951 ( .I(n63372), .Z(n61743) );
  NOR2_X1 U9954 ( .A1(n64486), .A2(n64485), .ZN(n1032) );
  NAND2_X1 U9957 ( .A1(n38048), .A2(n62427), .ZN(n62426) );
  NAND2_X1 U9959 ( .A1(n62956), .A2(n62955), .ZN(n58565) );
  NAND2_X1 U9961 ( .A1(n58051), .A2(n9998), .ZN(n65154) );
  NAND2_X1 U9964 ( .A1(n39928), .A2(n64487), .ZN(n64486) );
  AOI22_X1 U9972 ( .A1(n40252), .A2(n40251), .B1(n40253), .B2(n40254), .ZN(
        n40255) );
  NAND2_X1 U9977 ( .A1(n39411), .A2(n39410), .ZN(n64852) );
  INV_X1 U9981 ( .I(n64249), .ZN(n64248) );
  NAND2_X1 U9988 ( .A1(n13137), .A2(n13135), .ZN(n64902) );
  NOR2_X1 U9993 ( .A1(n6582), .A2(n37060), .ZN(n64023) );
  AOI21_X1 U9996 ( .A1(n41413), .A2(n41412), .B(n63839), .ZN(n13265) );
  OAI21_X1 U9997 ( .A1(n62185), .A2(n61435), .B(n41954), .ZN(n8403) );
  NAND3_X1 U9999 ( .A1(n40439), .A2(n40438), .A3(n59591), .ZN(n64184) );
  NAND2_X1 U10000 ( .A1(n37719), .A2(n42234), .ZN(n41953) );
  NAND2_X1 U10002 ( .A1(n22359), .A2(n22357), .ZN(n62233) );
  NAND2_X1 U10012 ( .A1(n12868), .A2(n19962), .ZN(n58051) );
  OAI21_X1 U10015 ( .A1(n40245), .A2(n40244), .B(n40243), .ZN(n40246) );
  NAND2_X1 U10016 ( .A1(n40812), .A2(n42276), .ZN(n65116) );
  AOI22_X1 U10022 ( .A1(n61707), .A2(n40541), .B1(n17213), .B2(n40542), .ZN(
        n3868) );
  NAND2_X1 U10026 ( .A1(n58797), .A2(n60810), .ZN(n62827) );
  INV_X1 U10028 ( .I(n41307), .ZN(n63919) );
  NAND2_X1 U10029 ( .A1(n39930), .A2(n39929), .ZN(n64485) );
  NAND2_X1 U10031 ( .A1(n62870), .A2(n39806), .ZN(n39814) );
  AOI22_X1 U10038 ( .A1(n63467), .A2(n41222), .B1(n41223), .B2(n41224), .ZN(
        n41226) );
  NAND3_X1 U10042 ( .A1(n62857), .A2(n20807), .A3(n62856), .ZN(n22357) );
  NAND2_X1 U10056 ( .A1(n12191), .A2(n12192), .ZN(n12190) );
  NAND2_X1 U10057 ( .A1(n39421), .A2(n9215), .ZN(n62666) );
  NOR2_X1 U10058 ( .A1(n40794), .A2(n40797), .ZN(n62205) );
  AND3_X1 U10064 ( .A1(n19726), .A2(n64675), .A3(n40087), .Z(n61792) );
  NAND2_X1 U10066 ( .A1(n62368), .A2(n42261), .ZN(n41098) );
  INV_X1 U10070 ( .I(n42268), .ZN(n62482) );
  NOR2_X1 U10099 ( .A1(n41091), .A2(n22502), .ZN(n62524) );
  OAI21_X1 U10101 ( .A1(n63204), .A2(n63203), .B(n40443), .ZN(n25357) );
  AOI21_X1 U10103 ( .A1(n12345), .A2(n11895), .B(n12344), .ZN(n12343) );
  INV_X1 U10104 ( .I(n42231), .ZN(n62185) );
  NAND2_X1 U10106 ( .A1(n39678), .A2(n41122), .ZN(n64247) );
  NAND2_X1 U10108 ( .A1(n41892), .A2(n41891), .ZN(n63867) );
  NAND2_X1 U10114 ( .A1(n62018), .A2(n65128), .ZN(n64487) );
  NAND2_X1 U10118 ( .A1(n40854), .A2(n64224), .ZN(n24863) );
  NAND2_X1 U10121 ( .A1(n64831), .A2(n64830), .ZN(n59856) );
  NAND2_X1 U10122 ( .A1(n5775), .A2(n11787), .ZN(n39145) );
  NOR2_X1 U10129 ( .A1(n40420), .A2(n40760), .ZN(n63756) );
  BUF_X1 U10133 ( .I(n10500), .Z(n65202) );
  NAND2_X1 U10138 ( .A1(n41476), .A2(n40413), .ZN(n62870) );
  NAND2_X1 U10145 ( .A1(n40853), .A2(n40854), .ZN(n63092) );
  NAND2_X1 U10153 ( .A1(n40300), .A2(n40296), .ZN(n62008) );
  INV_X1 U10162 ( .I(n39912), .ZN(n62009) );
  OR2_X1 U10164 ( .A1(n2895), .A2(n19466), .Z(n61780) );
  BUF_X2 U10170 ( .I(n4632), .Z(n58599) );
  OR2_X1 U10175 ( .A1(n40603), .A2(n37532), .Z(n61800) );
  AOI21_X1 U10179 ( .A1(n40750), .A2(n62565), .B(n24649), .ZN(n39988) );
  CLKBUF_X2 U10191 ( .I(n3345), .Z(n64224) );
  AOI21_X1 U10192 ( .A1(n37827), .A2(n64590), .B(n19045), .ZN(n12344) );
  INV_X1 U10197 ( .I(n62474), .ZN(n5506) );
  NAND2_X1 U10201 ( .A1(n40792), .A2(n40791), .ZN(n63264) );
  CLKBUF_X4 U10218 ( .I(n41447), .Z(n64773) );
  INV_X2 U10219 ( .I(n9396), .ZN(n64367) );
  INV_X2 U10224 ( .I(n40987), .ZN(n40147) );
  NOR2_X1 U10226 ( .A1(n41877), .A2(n222), .ZN(n64590) );
  NOR2_X1 U10228 ( .A1(n40763), .A2(n41470), .ZN(n40764) );
  NOR2_X1 U10236 ( .A1(n40417), .A2(n24982), .ZN(n64830) );
  INV_X1 U10241 ( .I(n9091), .ZN(n62857) );
  CLKBUF_X2 U10243 ( .I(n40716), .Z(n64493) );
  CLKBUF_X4 U10256 ( .I(n38516), .Z(n40617) );
  CLKBUF_X2 U10259 ( .I(n3705), .Z(n65199) );
  CLKBUF_X2 U10260 ( .I(n40923), .Z(n63303) );
  CLKBUF_X2 U10274 ( .I(n3246), .Z(n62175) );
  CLKBUF_X2 U10279 ( .I(n61094), .Z(n64826) );
  NAND2_X1 U10282 ( .A1(n40470), .A2(n40258), .ZN(n63800) );
  INV_X2 U10285 ( .I(n63952), .ZN(n11345) );
  CLKBUF_X2 U10300 ( .I(n42504), .Z(n23744) );
  INV_X4 U10301 ( .I(n22759), .ZN(n61746) );
  BUF_X2 U10310 ( .I(n39842), .Z(n22832) );
  BUF_X2 U10323 ( .I(n41874), .Z(n64592) );
  BUF_X2 U10335 ( .I(n37059), .Z(n40996) );
  CLKBUF_X2 U10339 ( .I(n40842), .Z(n64732) );
  CLKBUF_X2 U10340 ( .I(n25021), .Z(n63730) );
  INV_X1 U10342 ( .I(n18578), .ZN(n18580) );
  CLKBUF_X1 U10345 ( .I(n22561), .Z(n62027) );
  BUF_X2 U10353 ( .I(n12253), .Z(n3244) );
  INV_X1 U10358 ( .I(n38537), .ZN(n58281) );
  CLKBUF_X4 U10361 ( .I(n24677), .Z(n64640) );
  BUF_X2 U10362 ( .I(n39578), .Z(n25914) );
  CLKBUF_X2 U10363 ( .I(n9885), .Z(n62966) );
  CLKBUF_X2 U10371 ( .I(n18831), .Z(n65046) );
  CLKBUF_X2 U10377 ( .I(n6045), .Z(n65210) );
  NAND2_X1 U10378 ( .A1(n6138), .A2(n6139), .ZN(n13460) );
  CLKBUF_X2 U10382 ( .I(n38330), .Z(n62864) );
  CLKBUF_X2 U10385 ( .I(n23637), .Z(n62502) );
  NOR2_X1 U10395 ( .A1(n614), .A2(n36690), .ZN(n21942) );
  INV_X1 U10401 ( .I(n11600), .ZN(n62266) );
  AOI21_X1 U10406 ( .A1(n35407), .A2(n23146), .B(n63770), .ZN(n35412) );
  BUF_X4 U10410 ( .I(n39644), .Z(n23330) );
  NOR2_X1 U10413 ( .A1(n63810), .A2(n19874), .ZN(n19873) );
  NAND2_X1 U10414 ( .A1(n23387), .A2(n13929), .ZN(n13928) );
  NOR2_X1 U10419 ( .A1(n64058), .A2(n7723), .ZN(n7722) );
  NAND2_X1 U10426 ( .A1(n23495), .A2(n12341), .ZN(n62267) );
  NOR2_X1 U10427 ( .A1(n11777), .A2(n57607), .ZN(n64742) );
  NAND2_X1 U10428 ( .A1(n11558), .A2(n7483), .ZN(n62223) );
  NAND2_X1 U10443 ( .A1(n36480), .A2(n36584), .ZN(n63982) );
  NAND2_X1 U10447 ( .A1(n35726), .A2(n35725), .ZN(n64074) );
  NOR2_X1 U10453 ( .A1(n64020), .A2(n37248), .ZN(n61652) );
  AOI21_X1 U10456 ( .A1(n64988), .A2(n7967), .B(n7966), .ZN(n9580) );
  AOI21_X1 U10457 ( .A1(n36261), .A2(n9042), .B(n9041), .ZN(n10671) );
  NAND2_X1 U10462 ( .A1(n14618), .A2(n8549), .ZN(n8548) );
  NAND2_X1 U10468 ( .A1(n34483), .A2(n63088), .ZN(n25983) );
  NAND3_X1 U10478 ( .A1(n36667), .A2(n20203), .A3(n36666), .ZN(n65121) );
  INV_X1 U10484 ( .I(n7643), .ZN(n36458) );
  INV_X1 U10487 ( .I(n62948), .ZN(n21692) );
  NOR2_X1 U10495 ( .A1(n63645), .A2(n63644), .ZN(n32154) );
  INV_X1 U10496 ( .I(n9513), .ZN(n36229) );
  AOI22_X1 U10503 ( .A1(n61782), .A2(n37375), .B1(n36596), .B2(n36514), .ZN(
        n58938) );
  NAND2_X1 U10507 ( .A1(n15442), .A2(n37018), .ZN(n35077) );
  OAI21_X1 U10508 ( .A1(n61855), .A2(n19252), .B(n63762), .ZN(n33941) );
  NAND2_X1 U10510 ( .A1(n37105), .A2(n2220), .ZN(n63191) );
  NAND2_X1 U10513 ( .A1(n35950), .A2(n3128), .ZN(n35951) );
  NAND2_X1 U10514 ( .A1(n63456), .A2(n61937), .ZN(n64020) );
  INV_X1 U10520 ( .I(n11081), .ZN(n62576) );
  NAND2_X1 U10525 ( .A1(n36077), .A2(n36076), .ZN(n63990) );
  OAI22_X1 U10526 ( .A1(n35939), .A2(n37419), .B1(n35941), .B2(n35940), .ZN(
        n35942) );
  INV_X1 U10537 ( .I(n11721), .ZN(n9273) );
  INV_X2 U10545 ( .I(n36588), .ZN(n36512) );
  AND3_X1 U10547 ( .A1(n37085), .A2(n37940), .A3(n37096), .Z(n61855) );
  NOR2_X1 U10552 ( .A1(n35061), .A2(n64429), .ZN(n64428) );
  NOR2_X1 U10563 ( .A1(n57573), .A2(n36904), .ZN(n62655) );
  NAND2_X1 U10572 ( .A1(n61919), .A2(n63697), .ZN(n63696) );
  INV_X2 U10577 ( .I(n36610), .ZN(n36987) );
  NOR2_X1 U10580 ( .A1(n37064), .A2(n8520), .ZN(n62148) );
  AOI22_X1 U10586 ( .A1(n35595), .A2(n64753), .B1(n36227), .B2(n36225), .ZN(
        n35600) );
  NAND2_X1 U10593 ( .A1(n36219), .A2(n1531), .ZN(n62092) );
  OR2_X1 U10597 ( .A1(n33716), .A2(n35974), .Z(n4368) );
  NOR2_X1 U10620 ( .A1(n36118), .A2(n35363), .ZN(n35113) );
  CLKBUF_X2 U10623 ( .I(n37328), .Z(n62734) );
  CLKBUF_X4 U10643 ( .I(n37492), .Z(n63430) );
  INV_X1 U10648 ( .I(n15940), .ZN(n62347) );
  NAND2_X1 U10656 ( .A1(n35491), .A2(n14904), .ZN(n35492) );
  INV_X1 U10667 ( .I(n65036), .ZN(n57278) );
  INV_X1 U10669 ( .I(n36308), .ZN(n36789) );
  CLKBUF_X2 U10670 ( .I(n7380), .Z(n63247) );
  NOR2_X1 U10681 ( .A1(n61936), .A2(n35121), .ZN(n57617) );
  INV_X1 U10682 ( .I(n3076), .ZN(n62858) );
  CLKBUF_X2 U10686 ( .I(n7118), .Z(n64679) );
  CLKBUF_X2 U10695 ( .I(n36853), .Z(n7208) );
  CLKBUF_X2 U10699 ( .I(n15805), .Z(n62672) );
  CLKBUF_X4 U10709 ( .I(n34695), .Z(n36846) );
  BUF_X2 U10710 ( .I(n36494), .Z(n64093) );
  INV_X2 U10719 ( .I(n35852), .ZN(n61438) );
  CLKBUF_X4 U10721 ( .I(n35427), .Z(n504) );
  BUF_X4 U10734 ( .I(n36986), .Z(n18583) );
  CLKBUF_X2 U10744 ( .I(n37036), .Z(n62514) );
  NOR2_X1 U10747 ( .A1(n31525), .A2(n63815), .ZN(n22074) );
  NAND2_X1 U10750 ( .A1(n62317), .A2(n34653), .ZN(n25206) );
  AOI21_X1 U10754 ( .A1(n35837), .A2(n33210), .B(n64626), .ZN(n64885) );
  INV_X1 U10770 ( .I(n62342), .ZN(n25308) );
  BUF_X8 U10771 ( .I(n60140), .Z(n61747) );
  INV_X1 U10772 ( .I(n62447), .ZN(n62446) );
  NOR2_X1 U10775 ( .A1(n13129), .A2(n63996), .ZN(n13128) );
  NOR2_X1 U10781 ( .A1(n61852), .A2(n61996), .ZN(n61995) );
  NAND2_X1 U10782 ( .A1(n63285), .A2(n33687), .ZN(n6053) );
  OAI22_X1 U10785 ( .A1(n35733), .A2(n35734), .B1(n904), .B2(n35732), .ZN(
        n62342) );
  NAND2_X1 U10790 ( .A1(n13469), .A2(n2510), .ZN(n63986) );
  INV_X1 U10795 ( .I(n64676), .ZN(n59815) );
  AOI21_X1 U10812 ( .A1(n32358), .A2(n34795), .B(n61823), .ZN(n63331) );
  INV_X1 U10813 ( .I(n62460), .ZN(n19275) );
  NOR2_X1 U10815 ( .A1(n62878), .A2(n12237), .ZN(n3224) );
  NOR2_X1 U10818 ( .A1(n33407), .A2(n33619), .ZN(n64153) );
  INV_X1 U10836 ( .I(n35700), .ZN(n63079) );
  NAND3_X1 U10837 ( .A1(n32696), .A2(n32697), .A3(n61854), .ZN(n59298) );
  OAI21_X1 U10838 ( .A1(n20607), .A2(n34596), .B(n7969), .ZN(n65167) );
  OAI21_X1 U10842 ( .A1(n19922), .A2(n33686), .B(n33685), .ZN(n63285) );
  NAND2_X1 U10844 ( .A1(n32953), .A2(n64933), .ZN(n64932) );
  AOI22_X1 U10845 ( .A1(n35234), .A2(n35235), .B1(n35233), .B2(n35842), .ZN(
        n35236) );
  NOR2_X1 U10850 ( .A1(n12849), .A2(n63625), .ZN(n15642) );
  NAND2_X1 U10853 ( .A1(n14045), .A2(n14046), .ZN(n62878) );
  NOR2_X1 U10858 ( .A1(n33978), .A2(n64618), .ZN(n19337) );
  NAND2_X1 U10861 ( .A1(n3560), .A2(n1807), .ZN(n9910) );
  AOI21_X1 U10877 ( .A1(n1803), .A2(n64707), .B(n64706), .ZN(n35029) );
  NOR2_X1 U10879 ( .A1(n18680), .A2(n18679), .ZN(n65134) );
  INV_X1 U10891 ( .I(n35202), .ZN(n62697) );
  NAND2_X1 U10893 ( .A1(n17425), .A2(n34305), .ZN(n63844) );
  AOI21_X1 U10894 ( .A1(n19780), .A2(n23223), .B(n62967), .ZN(n60318) );
  AOI21_X1 U10895 ( .A1(n64604), .A2(n64603), .B(n58421), .ZN(n2079) );
  NAND2_X1 U10897 ( .A1(n63318), .A2(n63317), .ZN(n32973) );
  CLKBUF_X4 U10903 ( .I(n60970), .Z(n64304) );
  BUF_X4 U10904 ( .I(n7661), .Z(n62373) );
  INV_X1 U10906 ( .I(n25563), .ZN(n9677) );
  CLKBUF_X2 U10907 ( .I(n15551), .Z(n64954) );
  NAND2_X1 U10912 ( .A1(n25175), .A2(n1810), .ZN(n64677) );
  INV_X1 U10913 ( .I(n35837), .ZN(n62698) );
  INV_X1 U10914 ( .I(n9766), .ZN(n64933) );
  INV_X1 U10923 ( .I(n34687), .ZN(n63861) );
  NOR2_X1 U10924 ( .A1(n31724), .A2(n19119), .ZN(n61982) );
  CLKBUF_X2 U10925 ( .I(n61249), .Z(n64358) );
  CLKBUF_X1 U10930 ( .I(n33098), .Z(n61483) );
  CLKBUF_X2 U10943 ( .I(n60633), .Z(n64100) );
  BUF_X2 U10948 ( .I(n33431), .Z(n34025) );
  BUF_X2 U10952 ( .I(n31840), .Z(n35806) );
  BUF_X2 U10957 ( .I(n31026), .Z(n33420) );
  BUF_X2 U10959 ( .I(n33453), .Z(n9687) );
  CLKBUF_X4 U10964 ( .I(n14872), .Z(n61749) );
  INV_X1 U10965 ( .I(n24548), .ZN(n64418) );
  INV_X1 U10969 ( .I(n26142), .ZN(n26141) );
  CLKBUF_X2 U10971 ( .I(n25106), .Z(n63892) );
  BUF_X2 U10972 ( .I(n26062), .Z(n23143) );
  BUF_X2 U10978 ( .I(n32495), .Z(n61497) );
  CLKBUF_X2 U10987 ( .I(n60259), .Z(n64035) );
  INV_X1 U10997 ( .I(n31431), .ZN(n63114) );
  NOR2_X1 U11001 ( .A1(n5296), .A2(n63447), .ZN(n5294) );
  CLKBUF_X2 U11005 ( .I(n32663), .Z(n65171) );
  NAND3_X1 U11006 ( .A1(n62721), .A2(n13945), .A3(n61309), .ZN(n14672) );
  CLKBUF_X2 U11012 ( .I(n33203), .Z(n63099) );
  NOR2_X1 U11016 ( .A1(n25036), .A2(n15926), .ZN(n25035) );
  NAND2_X1 U11017 ( .A1(n58408), .A2(n62036), .ZN(n18162) );
  NOR2_X1 U11028 ( .A1(n4482), .A2(n63513), .ZN(n25027) );
  NAND2_X1 U11030 ( .A1(n30791), .A2(n16647), .ZN(n16646) );
  AOI21_X1 U11035 ( .A1(n63535), .A2(n59202), .B(n61781), .ZN(n8093) );
  INV_X1 U11044 ( .I(n65049), .ZN(n58929) );
  AOI21_X1 U11046 ( .A1(n57733), .A2(n30729), .B(n61941), .ZN(n19628) );
  OR3_X1 U11048 ( .A1(n58388), .A2(n63450), .A3(n29242), .Z(n28755) );
  INV_X1 U11067 ( .I(n30838), .ZN(n17857) );
  INV_X1 U11068 ( .I(n62725), .ZN(n31285) );
  NOR3_X1 U11073 ( .A1(n65139), .A2(n65138), .A3(n29505), .ZN(n29507) );
  NOR2_X1 U11077 ( .A1(n30172), .A2(n62552), .ZN(n30180) );
  INV_X1 U11078 ( .I(n29757), .ZN(n62747) );
  INV_X1 U11082 ( .I(n63646), .ZN(n15898) );
  NOR2_X1 U11086 ( .A1(n64237), .A2(n64236), .ZN(n15883) );
  NAND2_X1 U11096 ( .A1(n63334), .A2(n63333), .ZN(n61386) );
  NAND3_X1 U11099 ( .A1(n28714), .A2(n28713), .A3(n6912), .ZN(n62773) );
  INV_X1 U11112 ( .I(n62806), .ZN(n62767) );
  NAND2_X1 U11114 ( .A1(n3723), .A2(n23237), .ZN(n8753) );
  INV_X1 U11118 ( .I(n64282), .ZN(n7878) );
  NAND2_X1 U11121 ( .A1(n28699), .A2(n3706), .ZN(n62509) );
  INV_X1 U11123 ( .I(n61229), .ZN(n63450) );
  NAND3_X1 U11125 ( .A1(n30594), .A2(n18810), .A3(n23918), .ZN(n14765) );
  AND2_X1 U11126 ( .A1(n30731), .A2(n14729), .Z(n61941) );
  NOR2_X1 U11127 ( .A1(n29789), .A2(n63304), .ZN(n29790) );
  INV_X1 U11132 ( .I(n31282), .ZN(n64998) );
  OR3_X1 U11141 ( .A1(n30262), .A2(n30261), .A3(n17410), .Z(n61904) );
  INV_X1 U11146 ( .I(n25526), .ZN(n62104) );
  AOI21_X1 U11149 ( .A1(n14944), .A2(n21263), .B(n62153), .ZN(n29051) );
  NAND2_X1 U11150 ( .A1(n3901), .A2(n63497), .ZN(n3900) );
  NOR2_X1 U11151 ( .A1(n22014), .A2(n1848), .ZN(n62669) );
  INV_X1 U11152 ( .I(n29949), .ZN(n27972) );
  OAI21_X1 U11155 ( .A1(n27788), .A2(n7947), .B(n7946), .ZN(n682) );
  INV_X1 U11160 ( .I(n22156), .ZN(n63259) );
  INV_X1 U11161 ( .I(n29235), .ZN(n65096) );
  INV_X1 U11162 ( .I(n30429), .ZN(n63334) );
  NAND2_X1 U11167 ( .A1(n28957), .A2(n3267), .ZN(n64906) );
  BUF_X1 U11168 ( .I(n29844), .Z(n63315) );
  INV_X1 U11180 ( .I(n30521), .ZN(n30522) );
  INV_X2 U11181 ( .I(n58448), .ZN(n61750) );
  INV_X1 U11185 ( .I(n22596), .ZN(n64229) );
  CLKBUF_X2 U11189 ( .I(n31105), .Z(n10102) );
  NOR2_X1 U11195 ( .A1(n26471), .A2(n26472), .ZN(n61985) );
  NOR2_X1 U11198 ( .A1(n27211), .A2(n27199), .ZN(n63241) );
  AOI21_X1 U11200 ( .A1(n5471), .A2(n29138), .B(n62284), .ZN(n5469) );
  NOR2_X1 U11201 ( .A1(n63512), .A2(n7807), .ZN(n7806) );
  NOR2_X1 U11207 ( .A1(n26406), .A2(n25159), .ZN(n65029) );
  NOR2_X1 U11209 ( .A1(n57395), .A2(n62895), .ZN(n11702) );
  AND2_X1 U11210 ( .A1(n14757), .A2(n22956), .Z(n61898) );
  NAND2_X1 U11218 ( .A1(n27291), .A2(n6519), .ZN(n62642) );
  NOR2_X1 U11221 ( .A1(n8777), .A2(n8778), .ZN(n27964) );
  AOI21_X1 U11224 ( .A1(n28190), .A2(n28189), .B(n64929), .ZN(n14922) );
  OAI21_X1 U11225 ( .A1(n26423), .A2(n7772), .B(n7771), .ZN(n63512) );
  NOR3_X1 U11226 ( .A1(n6773), .A2(n6774), .A3(n26457), .ZN(n6772) );
  INV_X1 U11228 ( .I(n7109), .ZN(n64942) );
  NOR2_X1 U11238 ( .A1(n61875), .A2(n27592), .ZN(n16088) );
  NAND2_X1 U11240 ( .A1(n64388), .A2(n91), .ZN(n61239) );
  INV_X1 U11250 ( .I(n7438), .ZN(n63302) );
  CLKBUF_X2 U11251 ( .I(n22514), .Z(n64451) );
  CLKBUF_X2 U11258 ( .I(n27821), .Z(n63525) );
  OR2_X1 U11262 ( .A1(n22648), .A2(n28620), .Z(n61771) );
  INV_X1 U11270 ( .I(n29123), .ZN(n63713) );
  CLKBUF_X2 U11271 ( .I(n38699), .Z(n63603) );
  CLKBUF_X2 U11281 ( .I(n25202), .Z(n62714) );
  CLKBUF_X2 U11298 ( .I(n29353), .Z(n62341) );
  CLKBUF_X2 U11302 ( .I(n28470), .Z(n63495) );
  INV_X1 U11306 ( .I(Ciphertext[130]), .ZN(n64857) );
  INV_X1 U11310 ( .I(n26936), .ZN(n26705) );
  INV_X1 U11319 ( .I(n19287), .ZN(n62715) );
  OAI21_X1 U11322 ( .A1(n26958), .A2(n7538), .B(n29303), .ZN(n6616) );
  NOR2_X1 U11323 ( .A1(n28034), .A2(n28033), .ZN(n28038) );
  INV_X1 U11324 ( .I(n26720), .ZN(n24941) );
  NAND2_X1 U11330 ( .A1(n27520), .A2(n27203), .ZN(n22857) );
  NOR2_X1 U11332 ( .A1(n27876), .A2(n7651), .ZN(n26797) );
  INV_X1 U11336 ( .I(n27386), .ZN(n21126) );
  OAI21_X1 U11340 ( .A1(n27560), .A2(n28383), .B(n7886), .ZN(n26628) );
  INV_X2 U11344 ( .I(n6345), .ZN(n28843) );
  NOR2_X1 U11348 ( .A1(n469), .A2(n28379), .ZN(n27562) );
  NAND2_X1 U11356 ( .A1(n60265), .A2(n63932), .ZN(n7220) );
  INV_X2 U11364 ( .I(n26536), .ZN(n27120) );
  NOR2_X1 U11367 ( .A1(n28008), .A2(n2790), .ZN(n22397) );
  NOR2_X1 U11370 ( .A1(n12707), .A2(n23591), .ZN(n27927) );
  OAI21_X1 U11377 ( .A1(n29147), .A2(n21511), .B(n18377), .ZN(n3413) );
  NOR2_X1 U11379 ( .A1(n2176), .A2(n27065), .ZN(n21949) );
  BUF_X2 U11388 ( .I(n24921), .Z(n10399) );
  INV_X1 U11393 ( .I(n24419), .ZN(n27274) );
  NOR2_X1 U11397 ( .A1(n22115), .A2(n26536), .ZN(n26614) );
  NAND2_X1 U11401 ( .A1(n1930), .A2(n1880), .ZN(n15207) );
  NOR2_X1 U11405 ( .A1(n26074), .A2(n27664), .ZN(n27829) );
  NOR2_X1 U11411 ( .A1(n61260), .A2(n28547), .ZN(n28550) );
  NAND2_X1 U11414 ( .A1(n13702), .A2(n28383), .ZN(n60728) );
  NAND2_X1 U11418 ( .A1(n28814), .A2(n28815), .ZN(n28817) );
  NOR2_X1 U11419 ( .A1(n27620), .A2(n27614), .ZN(n26461) );
  INV_X2 U11420 ( .I(n22234), .ZN(n20540) );
  AND2_X1 U11422 ( .A1(n29302), .A2(n5259), .Z(n61798) );
  NAND2_X1 U11425 ( .A1(n8302), .A2(n27849), .ZN(n7771) );
  AOI21_X1 U11431 ( .A1(n28622), .A2(n23540), .B(n26864), .ZN(n26865) );
  NAND2_X1 U11434 ( .A1(n60171), .A2(n2276), .ZN(n27370) );
  CLKBUF_X2 U11438 ( .I(n29119), .Z(n24080) );
  INV_X1 U11442 ( .I(n29150), .ZN(n1886) );
  NOR2_X1 U11447 ( .A1(n29334), .A2(n29338), .ZN(n28885) );
  OAI21_X1 U11449 ( .A1(n3828), .A2(n3827), .B(n9561), .ZN(n63727) );
  NOR2_X1 U11452 ( .A1(n59552), .A2(n63883), .ZN(n27491) );
  NAND2_X1 U11457 ( .A1(n26968), .A2(n856), .ZN(n19857) );
  OAI21_X1 U11458 ( .A1(n26739), .A2(n15648), .B(n26835), .ZN(n26420) );
  NAND2_X1 U11460 ( .A1(n26379), .A2(n26380), .ZN(n2008) );
  INV_X1 U11461 ( .I(n27203), .ZN(n28348) );
  AOI21_X1 U11463 ( .A1(n3294), .A2(n3293), .B(n11226), .ZN(n26520) );
  AOI22_X1 U11469 ( .A1(n28835), .A2(n28834), .B1(n29629), .B2(n28833), .ZN(
        n28841) );
  NAND2_X1 U11479 ( .A1(n26283), .A2(n7438), .ZN(n63299) );
  INV_X1 U11489 ( .I(n26500), .ZN(n27587) );
  CLKBUF_X1 U11491 ( .I(n64943), .Z(n63150) );
  BUF_X2 U11494 ( .I(n28223), .Z(n19170) );
  NAND3_X1 U11496 ( .A1(n28245), .A2(n27037), .A3(n60473), .ZN(n26528) );
  NAND2_X1 U11502 ( .A1(n3253), .A2(n64056), .ZN(n59454) );
  AOI21_X1 U11508 ( .A1(n27969), .A2(n27968), .B(n63722), .ZN(n15111) );
  NAND3_X1 U11513 ( .A1(n28278), .A2(n28279), .A3(n61021), .ZN(n28026) );
  OAI21_X1 U11514 ( .A1(n29361), .A2(n64810), .B(n10828), .ZN(n4885) );
  NOR2_X1 U11526 ( .A1(n31255), .A2(n31254), .ZN(n31257) );
  AOI21_X1 U11527 ( .A1(n24967), .A2(n27278), .B(n60543), .ZN(n24969) );
  AOI21_X1 U11529 ( .A1(n4457), .A2(n26376), .B(n62099), .ZN(n27394) );
  NAND2_X1 U11533 ( .A1(n29310), .A2(n10236), .ZN(n27450) );
  INV_X1 U11535 ( .I(n29304), .ZN(n27213) );
  NOR3_X1 U11540 ( .A1(n27296), .A2(n27295), .A3(n27928), .ZN(n27302) );
  INV_X1 U11542 ( .I(n3932), .ZN(n9685) );
  NAND3_X1 U11550 ( .A1(n28468), .A2(n28467), .A3(n8087), .ZN(n61581) );
  CLKBUF_X2 U11555 ( .I(n31261), .Z(n12125) );
  NOR2_X1 U11561 ( .A1(n30608), .A2(n30347), .ZN(n6271) );
  NOR2_X1 U11562 ( .A1(n27603), .A2(n28314), .ZN(n27077) );
  AOI21_X1 U11564 ( .A1(n60543), .A2(n28560), .B(n28559), .ZN(n29084) );
  NOR3_X1 U11568 ( .A1(n28176), .A2(n12741), .A3(n4715), .ZN(n6303) );
  NOR3_X1 U11573 ( .A1(n4188), .A2(n30183), .A3(n10629), .ZN(n30187) );
  NOR2_X1 U11576 ( .A1(n30223), .A2(n1869), .ZN(n24975) );
  INV_X1 U11581 ( .I(n31267), .ZN(n31273) );
  CLKBUF_X4 U11583 ( .I(n1445), .Z(n5153) );
  AOI21_X1 U11584 ( .A1(n28220), .A2(n5415), .B(n5414), .ZN(n14148) );
  INV_X1 U11588 ( .I(n28952), .ZN(n14200) );
  NAND2_X1 U11596 ( .A1(n29813), .A2(n19451), .ZN(n26707) );
  NOR2_X1 U11602 ( .A1(n58395), .A2(n29397), .ZN(n31238) );
  CLKBUF_X4 U11603 ( .I(n15791), .Z(n17412) );
  NOR2_X1 U11609 ( .A1(n3086), .A2(n11092), .ZN(n30655) );
  CLKBUF_X1 U11611 ( .I(n30523), .Z(n58052) );
  NOR2_X1 U11622 ( .A1(n16961), .A2(n23397), .ZN(n60665) );
  NAND2_X1 U11633 ( .A1(n30348), .A2(n21029), .ZN(n30345) );
  NAND3_X1 U11636 ( .A1(n28117), .A2(n1867), .A3(n29848), .ZN(n14745) );
  NAND2_X1 U11637 ( .A1(n5631), .A2(n30197), .ZN(n29050) );
  NAND2_X1 U11658 ( .A1(n62588), .A2(n22893), .ZN(n62587) );
  NOR2_X1 U11669 ( .A1(n23705), .A2(n30844), .ZN(n2350) );
  NAND2_X1 U11671 ( .A1(n4210), .A2(n25898), .ZN(n5423) );
  INV_X1 U11676 ( .I(n13628), .ZN(n29427) );
  INV_X1 U11679 ( .I(n31119), .ZN(n11701) );
  CLKBUF_X4 U11685 ( .I(n28426), .Z(n30296) );
  NOR2_X1 U11693 ( .A1(n17508), .A2(n6680), .ZN(n14525) );
  AOI21_X1 U11698 ( .A1(n29592), .A2(n28917), .B(n40), .ZN(n63535) );
  NAND3_X1 U11701 ( .A1(n29394), .A2(n29393), .A3(n20683), .ZN(n20682) );
  NAND2_X1 U11704 ( .A1(n29986), .A2(n30322), .ZN(n28699) );
  NAND3_X1 U11708 ( .A1(n29860), .A2(n18736), .A3(n17412), .ZN(n21134) );
  NAND2_X1 U11715 ( .A1(n28754), .A2(n11830), .ZN(n30825) );
  OAI21_X1 U11720 ( .A1(n28712), .A2(n30655), .B(n30410), .ZN(n28713) );
  NAND2_X1 U11722 ( .A1(n27905), .A2(n64169), .ZN(n29901) );
  AOI21_X1 U11724 ( .A1(n24503), .A2(n24502), .B(n30430), .ZN(n25960) );
  NAND2_X1 U11726 ( .A1(n30816), .A2(n11830), .ZN(n63504) );
  CLKBUF_X4 U11728 ( .I(n26438), .Z(n30767) );
  CLKBUF_X4 U11743 ( .I(n28060), .Z(n30319) );
  NAND3_X1 U11744 ( .A1(n30339), .A2(n30616), .A3(n8097), .ZN(n30340) );
  NAND2_X1 U11747 ( .A1(n15147), .A2(n28093), .ZN(n15146) );
  NAND2_X1 U11748 ( .A1(n58829), .A2(n2572), .ZN(n3908) );
  NAND2_X1 U11750 ( .A1(n22164), .A2(n29015), .ZN(n17794) );
  INV_X1 U11759 ( .I(n4188), .ZN(n30190) );
  NAND2_X1 U11764 ( .A1(n62968), .A2(n11195), .ZN(n57862) );
  NOR2_X1 U11771 ( .A1(n22311), .A2(n30144), .ZN(n30155) );
  CLKBUF_X2 U11772 ( .I(n31215), .Z(n62892) );
  CLKBUF_X1 U11785 ( .I(n23111), .Z(n7423) );
  NOR2_X1 U11786 ( .A1(n31127), .A2(n29442), .ZN(n29911) );
  NAND2_X1 U11787 ( .A1(n7405), .A2(n20809), .ZN(n63417) );
  NAND2_X1 U11803 ( .A1(n29881), .A2(n27746), .ZN(n63251) );
  OR2_X1 U11807 ( .A1(n29490), .A2(n31092), .Z(n61913) );
  CLKBUF_X4 U11827 ( .I(n7405), .Z(n12632) );
  NAND2_X1 U11843 ( .A1(n28755), .A2(n30825), .ZN(n6469) );
  NOR2_X1 U11846 ( .A1(n31571), .A2(n29901), .ZN(n58366) );
  OAI21_X1 U11852 ( .A1(n30540), .A2(n30541), .B(n58747), .ZN(n57526) );
  AOI21_X1 U11867 ( .A1(n12300), .A2(n463), .B(n5688), .ZN(n57941) );
  OAI21_X1 U11871 ( .A1(n27423), .A2(n27422), .B(n30050), .ZN(n27428) );
  NAND2_X1 U11872 ( .A1(n21703), .A2(n21704), .ZN(n63217) );
  NOR2_X1 U11873 ( .A1(n11965), .A2(n11968), .ZN(n6107) );
  CLKBUF_X2 U11893 ( .I(n7058), .Z(n61462) );
  OAI22_X1 U11903 ( .A1(n18635), .A2(n61750), .B1(n30364), .B2(n30363), .ZN(
        n18634) );
  AND3_X1 U11911 ( .A1(n30226), .A2(n1350), .A3(n30843), .Z(n872) );
  OAI22_X1 U11922 ( .A1(n30078), .A2(n30077), .B1(n58630), .B2(n30076), .ZN(
        n30079) );
  NOR2_X1 U11934 ( .A1(n11032), .A2(n30098), .ZN(n62081) );
  CLKBUF_X2 U11936 ( .I(n17624), .Z(n62323) );
  INV_X1 U11942 ( .I(n1213), .ZN(n4441) );
  OAI21_X1 U11945 ( .A1(n29589), .A2(n29590), .B(n22504), .ZN(n62695) );
  CLKBUF_X1 U11952 ( .I(n31912), .Z(n19220) );
  AOI21_X1 U11959 ( .A1(n28702), .A2(n28701), .B(n62509), .ZN(n3390) );
  NOR2_X1 U11967 ( .A1(n19636), .A2(n25279), .ZN(n62937) );
  NAND2_X1 U11976 ( .A1(n7253), .A2(n9787), .ZN(n19587) );
  CLKBUF_X4 U11978 ( .I(n32289), .Z(n22390) );
  NOR2_X1 U11985 ( .A1(n19088), .A2(n62254), .ZN(n19178) );
  BUF_X2 U12015 ( .I(n32541), .Z(n22781) );
  NAND3_X1 U12017 ( .A1(n21228), .A2(n21227), .A3(n16037), .ZN(n6150) );
  INV_X1 U12044 ( .I(n32292), .ZN(n24790) );
  CLKBUF_X4 U12046 ( .I(n32483), .Z(n20862) );
  INV_X1 U12051 ( .I(n57218), .ZN(n15840) );
  CLKBUF_X2 U12054 ( .I(n18204), .Z(n63213) );
  INV_X1 U12089 ( .I(n24698), .ZN(n63759) );
  INV_X2 U12124 ( .I(n11930), .ZN(n32068) );
  INV_X1 U12126 ( .I(n32247), .ZN(n32637) );
  INV_X1 U12130 ( .I(n21321), .ZN(n21332) );
  INV_X1 U12135 ( .I(n58099), .ZN(n32228) );
  CLKBUF_X4 U12138 ( .I(n23706), .Z(n61610) );
  INV_X1 U12152 ( .I(n25741), .ZN(n1346) );
  CLKBUF_X2 U12156 ( .I(n8463), .Z(n59539) );
  INV_X1 U12159 ( .I(n33897), .ZN(n64431) );
  INV_X1 U12161 ( .I(n31687), .ZN(n63496) );
  INV_X1 U12167 ( .I(n31654), .ZN(n32106) );
  INV_X1 U12170 ( .I(n32332), .ZN(n22188) );
  NAND2_X1 U12175 ( .A1(n127), .A2(n7883), .ZN(n33500) );
  INV_X1 U12177 ( .I(n33729), .ZN(n32914) );
  AOI21_X1 U12183 ( .A1(n15551), .A2(n10340), .B(n35027), .ZN(n4938) );
  NAND2_X1 U12192 ( .A1(n34783), .A2(n61028), .ZN(n63317) );
  BUF_X2 U12195 ( .I(n21522), .Z(n21509) );
  NAND2_X1 U12201 ( .A1(n10448), .A2(n7272), .ZN(n10822) );
  AOI21_X1 U12202 ( .A1(n32889), .A2(n17866), .B(n34194), .ZN(n2402) );
  NAND2_X1 U12205 ( .A1(n57423), .A2(n21041), .ZN(n3668) );
  INV_X1 U12206 ( .I(n32271), .ZN(n63631) );
  NAND2_X1 U12212 ( .A1(n23127), .A2(n4880), .ZN(n64254) );
  INV_X1 U12220 ( .I(n35215), .ZN(n62470) );
  NOR2_X1 U12225 ( .A1(n60628), .A2(n34168), .ZN(n62583) );
  NAND2_X1 U12231 ( .A1(n65052), .A2(n23351), .ZN(n63668) );
  INV_X1 U12232 ( .I(n11981), .ZN(n24054) );
  NAND2_X1 U12241 ( .A1(n65119), .A2(n61262), .ZN(n4537) );
  INV_X1 U12244 ( .I(n60604), .ZN(n33747) );
  INV_X2 U12254 ( .I(n35224), .ZN(n35847) );
  NAND2_X1 U12255 ( .A1(n9843), .A2(n34446), .ZN(n4911) );
  NOR2_X1 U12270 ( .A1(n6925), .A2(n157), .ZN(n33664) );
  INV_X1 U12271 ( .I(n33987), .ZN(n60686) );
  INV_X1 U12273 ( .I(n21863), .ZN(n60805) );
  INV_X1 U12274 ( .I(n30934), .ZN(n33207) );
  OAI21_X1 U12275 ( .A1(n34190), .A2(n1312), .B(n34189), .ZN(n34191) );
  NOR2_X1 U12277 ( .A1(n33345), .A2(n7359), .ZN(n33348) );
  NOR2_X1 U12280 ( .A1(n1535), .A2(n11643), .ZN(n14615) );
  OAI21_X1 U12290 ( .A1(n64276), .A2(n23366), .B(n13081), .ZN(n34314) );
  INV_X2 U12293 ( .I(n13781), .ZN(n33763) );
  AOI21_X1 U12294 ( .A1(n34595), .A2(n3148), .B(n34594), .ZN(n7969) );
  NAND2_X1 U12297 ( .A1(n35675), .A2(n35674), .ZN(n4676) );
  NAND3_X1 U12298 ( .A1(n4075), .A2(n33963), .A3(n12039), .ZN(n4964) );
  INV_X2 U12299 ( .I(n33390), .ZN(n6925) );
  NAND2_X1 U12301 ( .A1(n33300), .A2(n4496), .ZN(n36543) );
  INV_X1 U12314 ( .I(n34733), .ZN(n34745) );
  NOR2_X1 U12315 ( .A1(n22342), .A2(n58713), .ZN(n11709) );
  CLKBUF_X4 U12316 ( .I(n34973), .Z(n22419) );
  INV_X1 U12320 ( .I(n34676), .ZN(n33455) );
  NAND2_X1 U12321 ( .A1(n18379), .A2(n24286), .ZN(n58226) );
  NAND3_X1 U12322 ( .A1(n35750), .A2(n63329), .A3(n61702), .ZN(n34418) );
  NAND2_X1 U12334 ( .A1(n32872), .A2(n139), .ZN(n33955) );
  INV_X1 U12338 ( .I(n34129), .ZN(n34140) );
  NAND2_X1 U12339 ( .A1(n34427), .A2(n10769), .ZN(n35324) );
  CLKBUF_X2 U12357 ( .I(n34958), .Z(n63123) );
  NAND2_X1 U12360 ( .A1(n8009), .A2(n3939), .ZN(n34333) );
  OAI21_X1 U12361 ( .A1(n33824), .A2(n33823), .B(n24286), .ZN(n33825) );
  CLKBUF_X4 U12363 ( .I(n35709), .Z(n23859) );
  NAND2_X1 U12364 ( .A1(n63557), .A2(n34384), .ZN(n62158) );
  OR2_X1 U12379 ( .A1(n35222), .A2(n35713), .Z(n64465) );
  NAND2_X1 U12386 ( .A1(n32993), .A2(n445), .ZN(n20182) );
  OAI21_X1 U12387 ( .A1(n14615), .A2(n14613), .B(n34658), .ZN(n62317) );
  NAND2_X1 U12391 ( .A1(n63844), .A2(n63843), .ZN(n17071) );
  INV_X1 U12393 ( .I(n35753), .ZN(n35761) );
  AND2_X1 U12410 ( .A1(n32359), .A2(n23645), .Z(n61823) );
  NOR3_X1 U12414 ( .A1(n5927), .A2(n35032), .A3(n5477), .ZN(n35035) );
  NAND3_X1 U12416 ( .A1(n34545), .A2(n34544), .A3(n34546), .ZN(n34549) );
  NAND2_X1 U12421 ( .A1(n34995), .A2(n30463), .ZN(n30462) );
  AOI22_X1 U12425 ( .A1(n32974), .A2(n33767), .B1(n57710), .B2(n34779), .ZN(
        n2507) );
  NAND2_X1 U12427 ( .A1(n20124), .A2(n22659), .ZN(n22823) );
  CLKBUF_X2 U12428 ( .I(n1427), .Z(n65189) );
  NAND2_X1 U12432 ( .A1(n33372), .A2(n59125), .ZN(n18244) );
  AND3_X1 U12441 ( .A1(n34307), .A2(n34217), .A3(n23567), .Z(n908) );
  AOI21_X1 U12444 ( .A1(n35846), .A2(n1343), .B(n35849), .ZN(n23160) );
  INV_X1 U12447 ( .I(n2695), .ZN(n21218) );
  INV_X2 U12451 ( .I(n33338), .ZN(n33596) );
  OAI22_X1 U12461 ( .A1(n34685), .A2(n33451), .B1(n34675), .B2(n34677), .ZN(
        n64356) );
  INV_X1 U12464 ( .I(n59769), .ZN(n31731) );
  CLKBUF_X4 U12474 ( .I(n35329), .Z(n10769) );
  INV_X1 U12476 ( .I(n35322), .ZN(n31956) );
  NOR2_X1 U12481 ( .A1(n33610), .A2(n64838), .ZN(n33617) );
  NAND3_X1 U12491 ( .A1(n61811), .A2(n7173), .A3(n2968), .ZN(n34060) );
  AOI21_X1 U12492 ( .A1(n60700), .A2(n59769), .B(n34113), .ZN(n32790) );
  NAND2_X1 U12496 ( .A1(n35004), .A2(n35003), .ZN(n34799) );
  NAND3_X1 U12502 ( .A1(n34260), .A2(n34340), .A3(n32004), .ZN(n32023) );
  NAND3_X1 U12503 ( .A1(n35642), .A2(n35660), .A3(n35643), .ZN(n33796) );
  OAI22_X1 U12509 ( .A1(n8366), .A2(n20182), .B1(n33550), .B2(n35611), .ZN(
        n32996) );
  INV_X1 U12511 ( .I(n34275), .ZN(n10016) );
  NAND2_X1 U12512 ( .A1(n26052), .A2(n18496), .ZN(n5740) );
  INV_X1 U12519 ( .I(n35721), .ZN(n62661) );
  INV_X1 U12520 ( .I(n7321), .ZN(n35214) );
  AOI21_X1 U12521 ( .A1(n30462), .A2(n12350), .B(n30461), .ZN(n30466) );
  NOR2_X1 U12529 ( .A1(n1779), .A2(n35881), .ZN(n58555) );
  AOI21_X1 U12532 ( .A1(n35021), .A2(n1538), .B(n16580), .ZN(n14811) );
  INV_X1 U12536 ( .I(n35946), .ZN(n16444) );
  INV_X1 U12541 ( .I(n33675), .ZN(n12820) );
  OAI21_X1 U12544 ( .A1(n1310), .A2(n64679), .B(n59147), .ZN(n36209) );
  NAND2_X1 U12545 ( .A1(n59319), .A2(n20102), .ZN(n20101) );
  NAND2_X1 U12563 ( .A1(n64934), .A2(n64932), .ZN(n64931) );
  NOR2_X1 U12565 ( .A1(n22503), .A2(n8177), .ZN(n35938) );
  INV_X1 U12567 ( .I(n20020), .ZN(n62340) );
  NOR3_X1 U12594 ( .A1(n22632), .A2(n2594), .A3(n9783), .ZN(n36509) );
  NAND2_X1 U12598 ( .A1(n17615), .A2(n25964), .ZN(n8132) );
  AOI21_X1 U12601 ( .A1(n35567), .A2(n1788), .B(n1779), .ZN(n31779) );
  NAND2_X1 U12605 ( .A1(n35274), .A2(n35275), .ZN(n21766) );
  NAND3_X1 U12606 ( .A1(n1338), .A2(n36956), .A3(n13557), .ZN(n35055) );
  NAND2_X1 U12609 ( .A1(n36174), .A2(n12804), .ZN(n14618) );
  NAND2_X1 U12611 ( .A1(n37447), .A2(n37455), .ZN(n63456) );
  NAND2_X1 U12614 ( .A1(n36379), .A2(n3809), .ZN(n64179) );
  AOI22_X1 U12650 ( .A1(n33417), .A2(n21113), .B1(n33425), .B2(n33978), .ZN(
        n21112) );
  NAND2_X1 U12653 ( .A1(n36740), .A2(n12863), .ZN(n36743) );
  NOR2_X1 U12663 ( .A1(n37369), .A2(n37363), .ZN(n36508) );
  AOI21_X1 U12668 ( .A1(n59348), .A2(n59346), .B(n6922), .ZN(n60167) );
  OAI21_X1 U12671 ( .A1(n35422), .A2(n14189), .B(n65234), .ZN(n35061) );
  NAND2_X1 U12676 ( .A1(n22785), .A2(n64181), .ZN(n23677) );
  CLKBUF_X2 U12679 ( .I(n36533), .Z(n65075) );
  INV_X1 U12688 ( .I(n34877), .ZN(n34490) );
  CLKBUF_X4 U12691 ( .I(n23742), .Z(n3691) );
  INV_X1 U12697 ( .I(n37335), .ZN(n24661) );
  NAND2_X1 U12710 ( .A1(n26213), .A2(n36851), .ZN(n36673) );
  NAND3_X1 U12711 ( .A1(n37085), .A2(n37084), .A3(n12050), .ZN(n35078) );
  NOR3_X1 U12714 ( .A1(n9869), .A2(n37161), .A3(n37455), .ZN(n20792) );
  INV_X1 U12715 ( .I(n36841), .ZN(n36014) );
  NAND2_X1 U12735 ( .A1(n10110), .A2(n36794), .ZN(n36131) );
  INV_X1 U12739 ( .I(n37227), .ZN(n36264) );
  OAI21_X1 U12744 ( .A1(n36511), .A2(n37363), .B(n36512), .ZN(n59122) );
  NAND2_X1 U12745 ( .A1(n37446), .A2(n62992), .ZN(n37457) );
  NAND2_X1 U12750 ( .A1(n19252), .A2(n37085), .ZN(n37086) );
  INV_X1 U12752 ( .I(n34460), .ZN(n10271) );
  INV_X1 U12756 ( .I(n18857), .ZN(n35993) );
  NAND2_X1 U12765 ( .A1(n36961), .A2(n60437), .ZN(n60085) );
  INV_X2 U12769 ( .I(n4893), .ZN(n36471) );
  NOR2_X1 U12770 ( .A1(n8010), .A2(n37328), .ZN(n37011) );
  INV_X2 U12781 ( .I(n26052), .ZN(n7270) );
  NAND2_X1 U12782 ( .A1(n36800), .A2(n36808), .ZN(n36792) );
  NAND2_X1 U12788 ( .A1(n36483), .A2(n1525), .ZN(n19616) );
  NOR2_X1 U12790 ( .A1(n14904), .A2(n37030), .ZN(n35486) );
  NAND2_X1 U12803 ( .A1(n3128), .A2(n35508), .ZN(n35952) );
  NOR2_X1 U12807 ( .A1(n35985), .A2(n36706), .ZN(n35988) );
  INV_X1 U12810 ( .I(n35561), .ZN(n34874) );
  OAI21_X1 U12812 ( .A1(n35986), .A2(n35985), .B(n19354), .ZN(n3010) );
  AOI22_X1 U12814 ( .A1(n36708), .A2(n36707), .B1(n12763), .B2(n36706), .ZN(
        n36712) );
  NOR2_X1 U12831 ( .A1(n10317), .A2(n10413), .ZN(n36496) );
  INV_X1 U12833 ( .I(n21673), .ZN(n62636) );
  OAI21_X1 U12839 ( .A1(n37211), .A2(n59617), .B(n18583), .ZN(n36983) );
  AOI21_X1 U12846 ( .A1(n60831), .A2(n37111), .B(n36756), .ZN(n57479) );
  OAI21_X1 U12847 ( .A1(n3460), .A2(n37225), .B(n37222), .ZN(n36349) );
  NOR2_X1 U12848 ( .A1(n13321), .A2(n13322), .ZN(n62764) );
  AOI22_X1 U12852 ( .A1(n35094), .A2(n21904), .B1(n36606), .B2(n2483), .ZN(
        n21903) );
  NAND2_X1 U12859 ( .A1(n65121), .A2(n62942), .ZN(n30) );
  AOI22_X1 U12867 ( .A1(n36289), .A2(n36291), .B1(n36754), .B2(n15449), .ZN(
        n63661) );
  NOR2_X1 U12869 ( .A1(n63191), .A2(n61803), .ZN(n36297) );
  INV_X1 U12876 ( .I(n13767), .ZN(n37394) );
  OAI21_X1 U12887 ( .A1(n16988), .A2(n16987), .B(n35416), .ZN(n61553) );
  INV_X1 U12895 ( .I(n14010), .ZN(n60647) );
  NAND2_X1 U12903 ( .A1(n36943), .A2(n34914), .ZN(n35425) );
  INV_X1 U12907 ( .I(n23739), .ZN(n36892) );
  AOI21_X1 U12912 ( .A1(n37942), .A2(n37319), .B(n19252), .ZN(n2242) );
  NAND2_X1 U12919 ( .A1(n34864), .A2(n25663), .ZN(n57599) );
  OAI22_X1 U12920 ( .A1(n32859), .A2(n58080), .B1(n35573), .B2(n36031), .ZN(
        n32861) );
  OAI21_X1 U12928 ( .A1(n12116), .A2(n12834), .B(n24625), .ZN(n24624) );
  CLKBUF_X1 U12932 ( .I(n39618), .Z(n9931) );
  OAI22_X1 U12933 ( .A1(n7644), .A2(n7643), .B1(n36225), .B2(n36224), .ZN(
        n5459) );
  AOI22_X1 U12940 ( .A1(n17394), .A2(n17395), .B1(n17396), .B2(n16181), .ZN(
        n62415) );
  INV_X1 U12964 ( .I(n63661), .ZN(n2294) );
  AOI21_X1 U12967 ( .A1(n57541), .A2(n57542), .B(n61945), .ZN(n913) );
  NAND2_X1 U12971 ( .A1(n14397), .A2(n21457), .ZN(n6782) );
  CLKBUF_X2 U12977 ( .I(n25690), .Z(n61450) );
  CLKBUF_X2 U12989 ( .I(n21921), .Z(n59924) );
  CLKBUF_X4 U12998 ( .I(n39728), .Z(n23898) );
  NOR2_X1 U13016 ( .A1(n62267), .A2(n62266), .ZN(n62265) );
  OAI21_X1 U13033 ( .A1(n36922), .A2(n19763), .B(n24358), .ZN(n9495) );
  INV_X2 U13036 ( .I(n37582), .ZN(n39626) );
  INV_X1 U13038 ( .I(n35977), .ZN(n5110) );
  NOR2_X1 U13044 ( .A1(n34868), .A2(n57599), .ZN(n8494) );
  CLKBUF_X1 U13062 ( .I(n37875), .Z(n59882) );
  INV_X1 U13064 ( .I(n39690), .ZN(n39274) );
  CLKBUF_X4 U13080 ( .I(n39345), .Z(n15704) );
  CLKBUF_X4 U13105 ( .I(n39689), .Z(n22485) );
  INV_X1 U13106 ( .I(n38286), .ZN(n7998) );
  INV_X1 U13107 ( .I(n38659), .ZN(n38120) );
  INV_X1 U13119 ( .I(n21508), .ZN(n62070) );
  INV_X1 U13121 ( .I(n39385), .ZN(n12293) );
  CLKBUF_X2 U13130 ( .I(n58177), .Z(n62852) );
  INV_X1 U13140 ( .I(n39312), .ZN(n64612) );
  INV_X2 U13147 ( .I(n13548), .ZN(n13705) );
  AOI21_X1 U13153 ( .A1(n41453), .A2(n1507), .B(n40713), .ZN(n40676) );
  INV_X1 U13154 ( .I(n16511), .ZN(n14697) );
  INV_X1 U13156 ( .I(n37580), .ZN(n62324) );
  INV_X1 U13162 ( .I(n60039), .ZN(n64306) );
  INV_X1 U13165 ( .I(n42263), .ZN(n41091) );
  CLKBUF_X2 U13166 ( .I(n19687), .Z(n62923) );
  INV_X2 U13172 ( .I(n23962), .ZN(n4691) );
  NOR2_X1 U13173 ( .A1(n20598), .A2(n41051), .ZN(n61232) );
  CLKBUF_X2 U13175 ( .I(n22321), .Z(n60062) );
  CLKBUF_X2 U13181 ( .I(n795), .Z(n60532) );
  NAND2_X1 U13182 ( .A1(n22593), .A2(n15558), .ZN(n40194) );
  NAND2_X1 U13184 ( .A1(n41906), .A2(n37773), .ZN(n37774) );
  INV_X1 U13186 ( .I(n42273), .ZN(n63476) );
  INV_X1 U13187 ( .I(n38466), .ZN(n9474) );
  INV_X1 U13190 ( .I(n61494), .ZN(n65040) );
  NAND2_X1 U13193 ( .A1(n61233), .A2(n60091), .ZN(n59664) );
  NOR2_X1 U13194 ( .A1(n40104), .A2(n20047), .ZN(n38020) );
  NOR2_X1 U13196 ( .A1(n10341), .A2(n40949), .ZN(n25104) );
  NAND2_X1 U13198 ( .A1(n36648), .A2(n2234), .ZN(n2233) );
  INV_X1 U13202 ( .I(n11460), .ZN(n22653) );
  CLKBUF_X1 U13217 ( .I(n38758), .Z(n62565) );
  INV_X1 U13224 ( .I(n16980), .ZN(n63204) );
  NOR2_X1 U13227 ( .A1(n40577), .A2(n42259), .ZN(n62474) );
  INV_X1 U13245 ( .I(n42281), .ZN(n41933) );
  NAND2_X1 U13248 ( .A1(n11459), .A2(n41400), .ZN(n41403) );
  NAND3_X1 U13249 ( .A1(n59664), .A2(n1730), .A3(n23420), .ZN(n40831) );
  NAND2_X1 U13253 ( .A1(n64571), .A2(n38607), .ZN(n18592) );
  NAND2_X1 U13260 ( .A1(n40623), .A2(n40726), .ZN(n59455) );
  NAND2_X1 U13261 ( .A1(n40231), .A2(n11123), .ZN(n11122) );
  CLKBUF_X2 U13262 ( .I(n11278), .Z(n11244) );
  NAND2_X1 U13263 ( .A1(n41006), .A2(n40607), .ZN(n40611) );
  NAND2_X1 U13268 ( .A1(n22809), .A2(n40924), .ZN(n40263) );
  NAND2_X1 U13269 ( .A1(n41799), .A2(n8404), .ZN(n63540) );
  NAND2_X1 U13270 ( .A1(n42458), .A2(n42448), .ZN(n5816) );
  INV_X2 U13281 ( .I(n59199), .ZN(n40162) );
  INV_X1 U13288 ( .I(n40294), .ZN(n14016) );
  INV_X1 U13290 ( .I(n40729), .ZN(n39029) );
  CLKBUF_X4 U13292 ( .I(n990), .Z(n1741) );
  AOI21_X1 U13294 ( .A1(n37596), .A2(n37597), .B(n59019), .ZN(n17353) );
  NAND2_X1 U13295 ( .A1(n41009), .A2(n58851), .ZN(n62956) );
  OAI21_X1 U13296 ( .A1(n8797), .A2(n39091), .B(n40519), .ZN(n25566) );
  OAI22_X1 U13297 ( .A1(n40712), .A2(n20994), .B1(n25777), .B2(n63464), .ZN(
        n7629) );
  INV_X2 U13298 ( .I(n40755), .ZN(n10683) );
  NAND2_X1 U13299 ( .A1(n10669), .A2(n40578), .ZN(n42260) );
  INV_X1 U13313 ( .I(n7237), .ZN(n1304) );
  CLKBUF_X2 U13316 ( .I(n41153), .Z(n64366) );
  AOI21_X1 U13326 ( .A1(n40831), .A2(n40830), .B(n64450), .ZN(n40836) );
  NAND2_X1 U13330 ( .A1(n12999), .A2(n41381), .ZN(n12998) );
  NAND3_X1 U13332 ( .A1(n40502), .A2(n40611), .A3(n40501), .ZN(n40503) );
  NOR2_X1 U13338 ( .A1(n63540), .A2(n63541), .ZN(n63539) );
  AOI21_X1 U13340 ( .A1(n38033), .A2(n40162), .B(n38032), .ZN(n25074) );
  NAND2_X1 U13343 ( .A1(n37996), .A2(n40099), .ZN(n40049) );
  AOI22_X1 U13347 ( .A1(n40502), .A2(n38420), .B1(n39118), .B2(n3612), .ZN(
        n57711) );
  NOR3_X1 U13349 ( .A1(n41454), .A2(n40712), .A3(n1516), .ZN(n8662) );
  NAND2_X1 U13351 ( .A1(n41178), .A2(n23616), .ZN(n39038) );
  OAI21_X1 U13357 ( .A1(n40683), .A2(n7629), .B(n58367), .ZN(n8314) );
  OAI21_X1 U13365 ( .A1(n57925), .A2(n41230), .B(n41231), .ZN(n39856) );
  NOR2_X1 U13366 ( .A1(n24863), .A2(n7618), .ZN(n24862) );
  NOR2_X1 U13367 ( .A1(n42292), .A2(n22609), .ZN(n42510) );
  NAND2_X1 U13389 ( .A1(n42252), .A2(n1744), .ZN(n41261) );
  INV_X1 U13391 ( .I(n16497), .ZN(n42431) );
  AOI22_X1 U13395 ( .A1(n40147), .A2(n6581), .B1(n40217), .B2(n39325), .ZN(
        n39327) );
  NAND2_X1 U13396 ( .A1(n41934), .A2(n59019), .ZN(n42290) );
  INV_X1 U13400 ( .I(n41642), .ZN(n63654) );
  NAND2_X1 U13408 ( .A1(n63756), .A2(n59856), .ZN(n59855) );
  CLKBUF_X1 U13415 ( .I(n21055), .Z(n59263) );
  NOR2_X1 U13417 ( .A1(n41258), .A2(n42240), .ZN(n41916) );
  OAI21_X1 U13419 ( .A1(n41949), .A2(n41947), .B(n41799), .ZN(n6223) );
  AOI21_X1 U13437 ( .A1(n9091), .A2(n39914), .B(n40139), .ZN(n39915) );
  AOI21_X1 U13442 ( .A1(n59976), .A2(n42211), .B(n42523), .ZN(n41836) );
  NOR2_X1 U13448 ( .A1(n39127), .A2(n18827), .ZN(n40522) );
  NAND3_X1 U13454 ( .A1(n40269), .A2(n18649), .A3(n40268), .ZN(n40270) );
  NAND2_X1 U13456 ( .A1(n21527), .A2(n16447), .ZN(n16448) );
  INV_X1 U13458 ( .I(n63036), .ZN(n10652) );
  INV_X1 U13461 ( .I(n20374), .ZN(n39060) );
  NAND2_X1 U13462 ( .A1(n62819), .A2(n40110), .ZN(n40115) );
  NOR3_X1 U13476 ( .A1(n20249), .A2(n42493), .A3(n40130), .ZN(n20248) );
  AOI21_X1 U13478 ( .A1(n40820), .A2(n40819), .B(n42277), .ZN(n40821) );
  NAND2_X1 U13481 ( .A1(n1333), .A2(n43657), .ZN(n2587) );
  NOR2_X1 U13489 ( .A1(n61660), .A2(n15671), .ZN(n57958) );
  OAI21_X1 U13495 ( .A1(n41442), .A2(n10877), .B(n10876), .ZN(n10875) );
  NAND2_X1 U13497 ( .A1(n64248), .A2(n64247), .ZN(n39703) );
  NAND2_X1 U13501 ( .A1(n43516), .A2(n61442), .ZN(n43181) );
  NAND2_X1 U13507 ( .A1(n17371), .A2(n42781), .ZN(n63977) );
  NAND2_X1 U13510 ( .A1(n64972), .A2(n41267), .ZN(n63921) );
  NAND2_X1 U13511 ( .A1(n42352), .A2(n42355), .ZN(n41616) );
  INV_X1 U13512 ( .I(n43318), .ZN(n14119) );
  NOR3_X1 U13514 ( .A1(n40525), .A2(n40527), .A3(n40526), .ZN(n40535) );
  NOR2_X1 U13516 ( .A1(n11986), .A2(n1503), .ZN(n43300) );
  NAND2_X1 U13519 ( .A1(n19975), .A2(n4274), .ZN(n4924) );
  NOR2_X1 U13524 ( .A1(n42631), .A2(n22186), .ZN(n8940) );
  INV_X1 U13527 ( .I(n37917), .ZN(n43698) );
  AOI22_X1 U13535 ( .A1(n40972), .A2(n6508), .B1(n40974), .B2(n40973), .ZN(
        n40976) );
  NOR2_X1 U13538 ( .A1(n3003), .A2(n1712), .ZN(n62058) );
  INV_X1 U13539 ( .I(n11635), .ZN(n43891) );
  INV_X1 U13554 ( .I(n16710), .ZN(n43414) );
  NOR2_X1 U13556 ( .A1(n43573), .A2(n4547), .ZN(n41657) );
  OAI21_X1 U13558 ( .A1(n43573), .A2(n25328), .B(n1391), .ZN(n42719) );
  INV_X1 U13576 ( .I(n42776), .ZN(n62624) );
  NOR2_X1 U13581 ( .A1(n61344), .A2(n8538), .ZN(n40912) );
  NAND2_X1 U13591 ( .A1(n19000), .A2(n43504), .ZN(n42641) );
  CLKBUF_X1 U13597 ( .I(n43156), .Z(n64251) );
  INV_X1 U13602 ( .I(n42698), .ZN(n42700) );
  INV_X1 U13613 ( .I(n42423), .ZN(n1712) );
  OAI22_X1 U13617 ( .A1(n42169), .A2(n16850), .B1(n42172), .B2(n58646), .ZN(
        n9941) );
  NOR2_X1 U13622 ( .A1(n15214), .A2(n43155), .ZN(n42890) );
  NAND2_X1 U13630 ( .A1(n42399), .A2(n42076), .ZN(n14506) );
  OAI21_X1 U13632 ( .A1(n42338), .A2(n43573), .B(n59746), .ZN(n41140) );
  NOR2_X1 U13637 ( .A1(n43917), .A2(n43922), .ZN(n65085) );
  OAI21_X1 U13645 ( .A1(n42621), .A2(n43415), .B(n62072), .ZN(n13202) );
  NAND2_X1 U13650 ( .A1(n43170), .A2(n15214), .ZN(n42562) );
  NOR2_X1 U13653 ( .A1(n14119), .A2(n1298), .ZN(n42198) );
  NAND2_X1 U13655 ( .A1(n5075), .A2(n15283), .ZN(n42360) );
  AOI21_X1 U13659 ( .A1(n8415), .A2(n63386), .B(n4924), .ZN(n14043) );
  OAI21_X1 U13660 ( .A1(n42018), .A2(n20284), .B(n16527), .ZN(n57932) );
  INV_X1 U13664 ( .I(n41496), .ZN(n43691) );
  NAND3_X1 U13668 ( .A1(n42316), .A2(n57873), .A3(n57241), .ZN(n42322) );
  NAND3_X1 U13676 ( .A1(n62510), .A2(n42947), .A3(n58678), .ZN(n18576) );
  NAND3_X1 U13681 ( .A1(n1908), .A2(n41773), .A3(n16850), .ZN(n42346) );
  NAND2_X1 U13686 ( .A1(n21644), .A2(n14920), .ZN(n42648) );
  BUF_X4 U13702 ( .I(n41549), .Z(n1715) );
  INV_X2 U13704 ( .I(n64462), .ZN(n43518) );
  NAND2_X1 U13705 ( .A1(n25851), .A2(n43464), .ZN(n16480) );
  INV_X2 U13707 ( .I(n42554), .ZN(n42923) );
  NAND2_X1 U13708 ( .A1(n43445), .A2(n43429), .ZN(n43426) );
  AOI21_X1 U13710 ( .A1(n43187), .A2(n64292), .B(n1017), .ZN(n20468) );
  INV_X1 U13718 ( .I(n41969), .ZN(n42380) );
  OAI22_X1 U13719 ( .A1(n41367), .A2(n17501), .B1(n42149), .B2(n41368), .ZN(
        n41372) );
  NOR2_X1 U13722 ( .A1(n42110), .A2(n41607), .ZN(n63506) );
  NAND3_X1 U13730 ( .A1(n64302), .A2(n62765), .A3(n24895), .ZN(n57682) );
  INV_X1 U13737 ( .I(n43992), .ZN(n43994) );
  NAND2_X1 U13738 ( .A1(n57410), .A2(n43327), .ZN(n14659) );
  NOR2_X1 U13739 ( .A1(n57256), .A2(n42188), .ZN(n1012) );
  AOI22_X1 U13743 ( .A1(n43219), .A2(n41353), .B1(n62297), .B2(n24250), .ZN(
        n41358) );
  NOR2_X1 U13745 ( .A1(n42137), .A2(n25235), .ZN(n63224) );
  OAI22_X1 U13758 ( .A1(n11748), .A2(n43842), .B1(n11746), .B2(n23485), .ZN(
        n62365) );
  INV_X1 U13760 ( .I(n20784), .ZN(n63752) );
  AOI22_X1 U13769 ( .A1(n42901), .A2(n60079), .B1(n42566), .B2(n64251), .ZN(
        n42060) );
  NOR2_X1 U13773 ( .A1(n60706), .A2(n41350), .ZN(n43078) );
  CLKBUF_X4 U13778 ( .I(n43778), .Z(n12089) );
  INV_X1 U13782 ( .I(n3208), .ZN(n44898) );
  INV_X1 U13783 ( .I(n21326), .ZN(n41560) );
  NOR2_X1 U13784 ( .A1(n42661), .A2(n64105), .ZN(n9440) );
  NAND2_X1 U13785 ( .A1(n40886), .A2(n41980), .ZN(n40885) );
  NAND3_X1 U13787 ( .A1(n58882), .A2(n58693), .A3(n43691), .ZN(n43037) );
  OAI22_X1 U13788 ( .A1(n42556), .A2(n9565), .B1(n9564), .B2(n9563), .ZN(
        n12424) );
  NAND2_X1 U13801 ( .A1(n39880), .A2(n62297), .ZN(n62375) );
  OAI21_X1 U13803 ( .A1(n24086), .A2(n40019), .B(n24085), .ZN(n12145) );
  AOI21_X1 U13807 ( .A1(n7215), .A2(n41331), .B(n20244), .ZN(n64688) );
  OAI21_X1 U13808 ( .A1(n43344), .A2(n43873), .B(n43343), .ZN(n43348) );
  AOI21_X1 U13811 ( .A1(n43362), .A2(n62237), .B(n43361), .ZN(n43368) );
  NAND2_X1 U13814 ( .A1(n57241), .A2(n5261), .ZN(n41990) );
  AOI21_X1 U13819 ( .A1(n61786), .A2(n43518), .B(n62194), .ZN(n62193) );
  NOR2_X1 U13823 ( .A1(n12916), .A2(n43041), .ZN(n43048) );
  NOR2_X1 U13828 ( .A1(n13630), .A2(n13882), .ZN(n15659) );
  AOI21_X1 U13831 ( .A1(n16201), .A2(n16740), .B(n16739), .ZN(n24732) );
  OAI22_X1 U13836 ( .A1(n4149), .A2(n3628), .B1(n42137), .B2(n42667), .ZN(
        n63226) );
  NAND2_X1 U13845 ( .A1(n63280), .A2(n43055), .ZN(n59795) );
  NOR2_X1 U13853 ( .A1(n57682), .A2(n57938), .ZN(n58944) );
  NOR3_X1 U13854 ( .A1(n12677), .A2(n16911), .A3(n22228), .ZN(n43949) );
  NOR2_X1 U13860 ( .A1(n63225), .A2(n63224), .ZN(n26234) );
  NAND3_X1 U13864 ( .A1(n41363), .A2(n42672), .A3(n63752), .ZN(n4637) );
  INV_X1 U13866 ( .I(n43909), .ZN(n62951) );
  CLKBUF_X2 U13871 ( .I(n23256), .Z(n64610) );
  NAND2_X1 U13873 ( .A1(n58690), .A2(n37922), .ZN(n18554) );
  NOR2_X1 U13875 ( .A1(n1502), .A2(n4945), .ZN(n43817) );
  AOI21_X1 U13876 ( .A1(n43355), .A2(n43354), .B(n61813), .ZN(n57428) );
  INV_X1 U13877 ( .I(n4264), .ZN(n62146) );
  INV_X1 U13881 ( .I(n39014), .ZN(n43051) );
  INV_X1 U13883 ( .I(n45281), .ZN(n24686) );
  AOI21_X1 U13888 ( .A1(n43004), .A2(n43003), .B(n43002), .ZN(n43005) );
  INV_X1 U13894 ( .I(n46321), .ZN(n59395) );
  AOI21_X1 U13895 ( .A1(n43871), .A2(n23151), .B(n41595), .ZN(n5681) );
  CLKBUF_X4 U13901 ( .I(n24450), .Z(n24449) );
  INV_X1 U13903 ( .I(n23365), .ZN(n63633) );
  INV_X1 U13908 ( .I(n46428), .ZN(n12002) );
  CLKBUF_X4 U13910 ( .I(n46495), .Z(n23440) );
  NOR2_X1 U13911 ( .A1(n39172), .A2(n62398), .ZN(n1913) );
  BUF_X2 U13917 ( .I(n44385), .Z(n23006) );
  CLKBUF_X4 U13921 ( .I(n14880), .Z(n2722) );
  INV_X2 U13933 ( .I(n16700), .ZN(n44731) );
  INV_X2 U13938 ( .I(n25629), .ZN(n58964) );
  INV_X1 U13947 ( .I(n44938), .ZN(n45032) );
  INV_X2 U13948 ( .I(n17919), .ZN(n21580) );
  INV_X1 U13951 ( .I(n44744), .ZN(n63869) );
  CLKBUF_X2 U13954 ( .I(n18709), .Z(n21895) );
  INV_X1 U13970 ( .I(n65058), .ZN(n18069) );
  INV_X1 U13972 ( .I(n15074), .ZN(n5408) );
  NAND3_X1 U13982 ( .A1(n43820), .A2(n43819), .A3(n41049), .ZN(n43370) );
  INV_X1 U13983 ( .I(n62065), .ZN(n17982) );
  INV_X1 U13990 ( .I(n18726), .ZN(n63325) );
  INV_X2 U14000 ( .I(n14513), .ZN(n7698) );
  INV_X1 U14001 ( .I(n8813), .ZN(n63642) );
  CLKBUF_X4 U14019 ( .I(n46430), .Z(n22551) );
  NAND2_X1 U14020 ( .A1(n63404), .A2(n17464), .ZN(n57426) );
  INV_X1 U14023 ( .I(n61672), .ZN(n60365) );
  INV_X1 U14024 ( .I(n46528), .ZN(n60124) );
  NAND2_X1 U14028 ( .A1(n25492), .A2(n25491), .ZN(n46186) );
  CLKBUF_X2 U14032 ( .I(n58310), .Z(n57785) );
  INV_X1 U14033 ( .I(n19947), .ZN(n7880) );
  NAND2_X1 U14034 ( .A1(n48514), .A2(n48521), .ZN(n48645) );
  NAND2_X1 U14035 ( .A1(n13413), .A2(n2955), .ZN(n11689) );
  CLKBUF_X1 U14036 ( .I(n1212), .Z(n7335) );
  NOR2_X1 U14037 ( .A1(n47488), .A2(n20162), .ZN(n62301) );
  NAND2_X1 U14040 ( .A1(n45768), .A2(n10512), .ZN(n44780) );
  NAND2_X1 U14041 ( .A1(n47883), .A2(n47880), .ZN(n63841) );
  INV_X2 U14043 ( .I(n11380), .ZN(n48499) );
  NOR2_X1 U14044 ( .A1(n47881), .A2(n45183), .ZN(n47362) );
  NAND2_X1 U14058 ( .A1(n1388), .A2(n1070), .ZN(n45770) );
  NOR2_X1 U14059 ( .A1(n12698), .A2(n47115), .ZN(n45803) );
  NOR2_X1 U14067 ( .A1(n47414), .A2(n61720), .ZN(n15555) );
  INV_X1 U14072 ( .I(n46095), .ZN(n44135) );
  NAND2_X1 U14087 ( .A1(n3510), .A2(n14630), .ZN(n64790) );
  NAND2_X1 U14090 ( .A1(n46941), .A2(n18127), .ZN(n24339) );
  NOR2_X1 U14094 ( .A1(n22326), .A2(n45765), .ZN(n44660) );
  NOR2_X1 U14096 ( .A1(n59670), .A2(n45955), .ZN(n62004) );
  NAND2_X1 U14097 ( .A1(n58018), .A2(n63232), .ZN(n63231) );
  NOR2_X1 U14103 ( .A1(n15359), .A2(n22468), .ZN(n7296) );
  NAND3_X1 U14115 ( .A1(n65196), .A2(n46733), .A3(n18980), .ZN(n64544) );
  NOR2_X1 U14117 ( .A1(n48153), .A2(n46794), .ZN(n11343) );
  INV_X2 U14123 ( .I(n47623), .ZN(n22239) );
  AOI21_X1 U14129 ( .A1(n63547), .A2(n48549), .B(n24364), .ZN(n48551) );
  CLKBUF_X4 U14136 ( .I(n16930), .Z(n65074) );
  INV_X1 U14160 ( .I(n64654), .ZN(n63500) );
  NAND3_X1 U14173 ( .A1(n44067), .A2(n44066), .A3(n46978), .ZN(n24022) );
  INV_X1 U14174 ( .I(n15817), .ZN(n47381) );
  INV_X1 U14190 ( .I(n47370), .ZN(n46821) );
  NAND2_X1 U14192 ( .A1(n47503), .A2(n1647), .ZN(n46267) );
  NAND3_X1 U14197 ( .A1(n44135), .A2(n44133), .A3(n7104), .ZN(n20307) );
  AOI21_X1 U14198 ( .A1(n8199), .A2(n48479), .B(n64634), .ZN(n8198) );
  CLKBUF_X2 U14208 ( .I(n57740), .Z(n63686) );
  NOR2_X1 U14223 ( .A1(n11929), .A2(n47560), .ZN(n5466) );
  NAND2_X1 U14228 ( .A1(n21246), .A2(n20832), .ZN(n21245) );
  INV_X1 U14229 ( .I(n45203), .ZN(n1481) );
  INV_X1 U14234 ( .I(n64406), .ZN(n48383) );
  AOI22_X1 U14237 ( .A1(n64969), .A2(n44681), .B1(n46985), .B2(n44065), .ZN(
        n44682) );
  INV_X2 U14252 ( .I(n5145), .ZN(n59698) );
  INV_X1 U14255 ( .I(n17670), .ZN(n47667) );
  CLKBUF_X4 U14257 ( .I(n47291), .Z(n20666) );
  NAND3_X1 U14261 ( .A1(n9772), .A2(n23394), .A3(n6977), .ZN(n16712) );
  NOR2_X1 U14263 ( .A1(n18477), .A2(n45775), .ZN(n45763) );
  INV_X1 U14265 ( .I(n6148), .ZN(n47263) );
  NOR2_X1 U14274 ( .A1(n58675), .A2(n47542), .ZN(n64912) );
  NAND3_X1 U14275 ( .A1(n17670), .A2(n13782), .A3(n47407), .ZN(n17746) );
  AOI21_X1 U14279 ( .A1(n11906), .A2(n11907), .B(n11897), .ZN(n57705) );
  AOI22_X1 U14283 ( .A1(n47596), .A2(n47593), .B1(n47592), .B2(n45683), .ZN(
        n45556) );
  AOI21_X1 U14291 ( .A1(n47239), .A2(n45204), .B(n61968), .ZN(n63804) );
  CLKBUF_X1 U14298 ( .I(n8012), .Z(n61993) );
  NAND2_X1 U14308 ( .A1(n46999), .A2(n7504), .ZN(n63087) );
  NAND2_X1 U14321 ( .A1(n22239), .A2(n7541), .ZN(n45204) );
  OAI21_X1 U14322 ( .A1(n46867), .A2(n46866), .B(n46865), .ZN(n46868) );
  AOI21_X1 U14324 ( .A1(n45986), .A2(n45987), .B(n47236), .ZN(n64851) );
  NOR2_X1 U14325 ( .A1(n45590), .A2(n45591), .ZN(n47904) );
  CLKBUF_X2 U14327 ( .I(n48148), .Z(n60138) );
  AOI21_X1 U14331 ( .A1(n47364), .A2(n58636), .B(n47718), .ZN(n45181) );
  NAND2_X1 U14338 ( .A1(n23416), .A2(n1212), .ZN(n48162) );
  INV_X1 U14339 ( .I(n47400), .ZN(n25749) );
  NAND2_X1 U14343 ( .A1(n45710), .A2(n46026), .ZN(n45654) );
  CLKBUF_X2 U14346 ( .I(n47470), .Z(n64969) );
  NOR2_X1 U14348 ( .A1(n47229), .A2(n46049), .ZN(n6495) );
  NAND3_X1 U14351 ( .A1(n14769), .A2(n48240), .A3(n14990), .ZN(n14768) );
  INV_X1 U14354 ( .I(n9299), .ZN(n47471) );
  INV_X1 U14368 ( .I(n21246), .ZN(n46061) );
  NAND2_X1 U14369 ( .A1(n11810), .A2(n47493), .ZN(n14962) );
  CLKBUF_X1 U14372 ( .I(n20340), .Z(n64231) );
  OAI21_X1 U14382 ( .A1(n18735), .A2(n2901), .B(n47803), .ZN(n57508) );
  AOI21_X1 U14384 ( .A1(n25812), .A2(n48341), .B(n14315), .ZN(n47785) );
  NAND2_X1 U14385 ( .A1(n44698), .A2(n44705), .ZN(n47030) );
  NOR2_X1 U14389 ( .A1(n1078), .A2(n3641), .ZN(n45640) );
  NAND2_X1 U14391 ( .A1(n46893), .A2(n47250), .ZN(n47249) );
  NOR2_X1 U14392 ( .A1(n44646), .A2(n63670), .ZN(n64440) );
  OR2_X1 U14395 ( .A1(n61624), .A2(n13614), .Z(n61821) );
  NAND4_X1 U14396 ( .A1(n43599), .A2(n47366), .A3(n47359), .A4(n43598), .ZN(
        n43600) );
  OAI21_X1 U14399 ( .A1(n16276), .A2(n17315), .B(n61628), .ZN(n63439) );
  OAI21_X1 U14400 ( .A1(n61993), .A2(n48604), .B(n48602), .ZN(n61211) );
  NAND2_X1 U14419 ( .A1(n49014), .A2(n49006), .ZN(n48038) );
  OAI21_X1 U14424 ( .A1(n63804), .A2(n47618), .B(n14414), .ZN(n58450) );
  NOR2_X1 U14435 ( .A1(n18047), .A2(n64584), .ZN(n64583) );
  AND3_X1 U14437 ( .A1(n7104), .A2(n47016), .A3(n47018), .Z(n61910) );
  CLKBUF_X4 U14439 ( .I(n43597), .Z(n47874) );
  NAND2_X1 U14444 ( .A1(n46889), .A2(n64281), .ZN(n64280) );
  NAND2_X1 U14450 ( .A1(n47596), .A2(n548), .ZN(n45982) );
  OAI21_X1 U14456 ( .A1(n10155), .A2(n8749), .B(n60946), .ZN(n8748) );
  NAND3_X1 U14458 ( .A1(n47866), .A2(n24096), .A3(n47865), .ZN(n4629) );
  CLKBUF_X2 U14459 ( .I(n1386), .Z(n64766) );
  NOR2_X1 U14463 ( .A1(n47877), .A2(n45183), .ZN(n45187) );
  AOI21_X1 U14470 ( .A1(n8582), .A2(n45565), .B(n10088), .ZN(n16597) );
  NAND2_X1 U14478 ( .A1(n25749), .A2(n24893), .ZN(n64220) );
  NAND3_X1 U14481 ( .A1(n46950), .A2(n6034), .A3(n46948), .ZN(n46075) );
  NAND3_X1 U14484 ( .A1(n59652), .A2(n45495), .A3(n59651), .ZN(n59403) );
  NAND2_X1 U14506 ( .A1(n46012), .A2(n45636), .ZN(n62613) );
  NAND3_X1 U14511 ( .A1(n12114), .A2(n45617), .A3(n45618), .ZN(n46064) );
  NAND2_X1 U14515 ( .A1(n25032), .A2(n65057), .ZN(n49593) );
  INV_X1 U14520 ( .I(n23500), .ZN(n9367) );
  INV_X1 U14522 ( .I(n50272), .ZN(n50269) );
  OAI21_X1 U14523 ( .A1(n63423), .A2(n47096), .B(n21820), .ZN(n21817) );
  NAND2_X1 U14534 ( .A1(n6130), .A2(n49923), .ZN(n10961) );
  NOR2_X1 U14537 ( .A1(n10422), .A2(n49538), .ZN(n48779) );
  OAI21_X1 U14542 ( .A1(n45788), .A2(n20938), .B(n19595), .ZN(n63139) );
  AOI21_X1 U14545 ( .A1(n45663), .A2(n44483), .B(n47251), .ZN(n16964) );
  NAND2_X1 U14547 ( .A1(n61821), .A2(n64759), .ZN(n15569) );
  NAND2_X1 U14552 ( .A1(n1209), .A2(n13614), .ZN(n11624) );
  INV_X1 U14553 ( .I(n49281), .ZN(n49287) );
  NOR2_X1 U14555 ( .A1(n11705), .A2(n49074), .ZN(n48048) );
  INV_X1 U14557 ( .I(n46004), .ZN(n49788) );
  NOR2_X1 U14559 ( .A1(n47935), .A2(n1473), .ZN(n59900) );
  AOI21_X1 U14562 ( .A1(n152), .A2(n64899), .B(n65103), .ZN(n1093) );
  CLKBUF_X1 U14564 ( .I(n64631), .Z(n63785) );
  OAI21_X1 U14567 ( .A1(n47095), .A2(n10117), .B(n64766), .ZN(n47106) );
  INV_X1 U14568 ( .I(n47075), .ZN(n60756) );
  NAND2_X1 U14569 ( .A1(n23707), .A2(n3030), .ZN(n49723) );
  NAND2_X1 U14571 ( .A1(n48859), .A2(n12701), .ZN(n48392) );
  NAND2_X1 U14573 ( .A1(n48454), .A2(n49013), .ZN(n7014) );
  OAI21_X1 U14576 ( .A1(n18433), .A2(n49526), .B(n61833), .ZN(n18432) );
  NOR2_X1 U14584 ( .A1(n57735), .A2(n21550), .ZN(n22174) );
  NAND3_X1 U14587 ( .A1(n47912), .A2(n49377), .A3(n3472), .ZN(n47915) );
  INV_X1 U14590 ( .I(n49762), .ZN(n49759) );
  OAI22_X1 U14592 ( .A1(n49264), .A2(n16745), .B1(n49265), .B2(n12558), .ZN(
        n12557) );
  INV_X1 U14594 ( .I(n49512), .ZN(n48286) );
  NAND2_X1 U14597 ( .A1(n49478), .A2(n64722), .ZN(n64721) );
  NAND4_X1 U14598 ( .A1(n17523), .A2(n57949), .A3(n8604), .A4(n49395), .ZN(
        n47062) );
  NOR2_X1 U14601 ( .A1(n48318), .A2(n13614), .ZN(n10716) );
  CLKBUF_X2 U14607 ( .I(n15319), .Z(n61089) );
  OAI21_X1 U14608 ( .A1(n11950), .A2(n49063), .B(n8298), .ZN(n48300) );
  AOI21_X1 U14613 ( .A1(n49077), .A2(n49063), .B(n48299), .ZN(n48049) );
  CLKBUF_X1 U14618 ( .I(n1224), .Z(n58861) );
  CLKBUF_X1 U14619 ( .I(n13925), .Z(n62192) );
  NAND2_X1 U14620 ( .A1(n49003), .A2(n47051), .ZN(n47053) );
  OAI21_X1 U14621 ( .A1(n50428), .A2(n63876), .B(n57572), .ZN(n50429) );
  NAND3_X1 U14624 ( .A1(n50425), .A2(n60853), .A3(n49249), .ZN(n7194) );
  NAND2_X1 U14625 ( .A1(n18142), .A2(n1381), .ZN(n19096) );
  NAND2_X1 U14626 ( .A1(n48963), .A2(n49411), .ZN(n49179) );
  NAND2_X1 U14631 ( .A1(n23707), .A2(n15386), .ZN(n49722) );
  NAND2_X1 U14635 ( .A1(n50214), .A2(n1383), .ZN(n12475) );
  NOR2_X1 U14636 ( .A1(n49000), .A2(n48310), .ZN(n9383) );
  CLKBUF_X2 U14640 ( .I(n49019), .Z(n63389) );
  CLKBUF_X2 U14641 ( .I(n49512), .Z(n64170) );
  NOR2_X1 U14645 ( .A1(n61089), .A2(n42), .ZN(n48831) );
  NOR2_X1 U14646 ( .A1(n50288), .A2(n48720), .ZN(n50121) );
  NAND2_X1 U14651 ( .A1(n48375), .A2(n49856), .ZN(n59957) );
  NAND3_X1 U14653 ( .A1(n49813), .A2(n50441), .A3(n50437), .ZN(n8898) );
  NOR2_X1 U14654 ( .A1(n64564), .A2(n17122), .ZN(n58053) );
  NAND3_X1 U14656 ( .A1(n49437), .A2(n8380), .A3(n49436), .ZN(n19851) );
  NAND2_X1 U14659 ( .A1(n20594), .A2(n22847), .ZN(n19481) );
  NAND2_X1 U14663 ( .A1(n19043), .A2(n9177), .ZN(n7747) );
  NAND2_X1 U14664 ( .A1(n49603), .A2(n49602), .ZN(n59085) );
  AOI22_X1 U14666 ( .A1(n47457), .A2(n49254), .B1(n50428), .B2(n50430), .ZN(
        n47460) );
  NAND3_X1 U14667 ( .A1(n60696), .A2(n50233), .A3(n60695), .ZN(n8728) );
  NOR2_X1 U14670 ( .A1(n23612), .A2(n49170), .ZN(n49175) );
  INV_X1 U14674 ( .I(n50289), .ZN(n57193) );
  NAND2_X1 U14675 ( .A1(n25830), .A2(n381), .ZN(n59828) );
  OAI21_X1 U14676 ( .A1(n22869), .A2(n49772), .B(n21550), .ZN(n48410) );
  NAND2_X1 U14678 ( .A1(n61612), .A2(n5282), .ZN(n50379) );
  NOR2_X1 U14684 ( .A1(n9321), .A2(n48280), .ZN(n63655) );
  CLKBUF_X4 U14685 ( .I(n20763), .Z(n60786) );
  NAND2_X1 U14689 ( .A1(n57204), .A2(n25018), .ZN(n48412) );
  NOR2_X1 U14691 ( .A1(n50421), .A2(n2755), .ZN(n49257) );
  CLKBUF_X2 U14696 ( .I(n22042), .Z(n60853) );
  NAND2_X1 U14698 ( .A1(n48965), .A2(n49179), .ZN(n15363) );
  OAI21_X1 U14703 ( .A1(n60464), .A2(n57224), .B(n59733), .ZN(n63082) );
  OAI21_X1 U14704 ( .A1(n48843), .A2(n48842), .B(n48841), .ZN(n48844) );
  OAI21_X1 U14708 ( .A1(n1643), .A2(n3055), .B(n50297), .ZN(n50136) );
  INV_X1 U14709 ( .I(n50549), .ZN(n11288) );
  CLKBUF_X2 U14717 ( .I(n49561), .Z(n63493) );
  NAND2_X1 U14718 ( .A1(n61866), .A2(n63110), .ZN(n64162) );
  CLKBUF_X4 U14719 ( .I(n50695), .Z(n52537) );
  NAND2_X1 U14724 ( .A1(n13317), .A2(n48847), .ZN(n13316) );
  CLKBUF_X4 U14726 ( .I(n23342), .Z(n9231) );
  OAI21_X1 U14727 ( .A1(n50020), .A2(n50021), .B(n7868), .ZN(n63737) );
  NAND2_X1 U14730 ( .A1(n25605), .A2(n63518), .ZN(n2501) );
  CLKBUF_X1 U14734 ( .I(n1205), .Z(n59966) );
  OAI21_X1 U14736 ( .A1(n50075), .A2(n59021), .B(n50400), .ZN(n19262) );
  NAND3_X1 U14746 ( .A1(n14042), .A2(n50087), .A3(n14041), .ZN(n15669) );
  NOR2_X1 U14749 ( .A1(n20211), .A2(n16177), .ZN(n25200) );
  CLKBUF_X2 U14761 ( .I(n7847), .Z(n58989) );
  INV_X1 U14769 ( .I(n52370), .ZN(n64094) );
  CLKBUF_X4 U14780 ( .I(n7331), .Z(n65143) );
  NAND2_X1 U14783 ( .A1(n52568), .A2(n51033), .ZN(n60911) );
  INV_X1 U14791 ( .I(n14299), .ZN(n11914) );
  AOI21_X1 U14793 ( .A1(n23372), .A2(n50234), .B(n22198), .ZN(n17925) );
  CLKBUF_X2 U14795 ( .I(n24640), .Z(n6597) );
  INV_X1 U14796 ( .I(n11071), .ZN(n7232) );
  INV_X1 U14800 ( .I(n2167), .ZN(n52148) );
  CLKBUF_X2 U14801 ( .I(n50648), .Z(n23149) );
  INV_X1 U14805 ( .I(n51701), .ZN(n21545) );
  CLKBUF_X2 U14808 ( .I(n50717), .Z(n23678) );
  INV_X1 U14810 ( .I(n51528), .ZN(n64259) );
  INV_X1 U14817 ( .I(n50371), .ZN(n62208) );
  INV_X1 U14833 ( .I(n57070), .ZN(n62885) );
  INV_X1 U14837 ( .I(n52523), .ZN(n62527) );
  NAND2_X1 U14841 ( .A1(n61725), .A2(n54594), .ZN(n25648) );
  NAND2_X1 U14842 ( .A1(n23736), .A2(n21364), .ZN(n54466) );
  NAND2_X1 U14853 ( .A1(n54493), .A2(n4473), .ZN(n52989) );
  INV_X1 U14854 ( .I(n54996), .ZN(n16848) );
  NAND2_X1 U14855 ( .A1(n15718), .A2(n57025), .ZN(n4183) );
  AOI21_X1 U14857 ( .A1(n23919), .A2(n55721), .B(n1324), .ZN(n55424) );
  NOR2_X1 U14860 ( .A1(n62886), .A2(n62885), .ZN(n62884) );
  INV_X1 U14868 ( .I(n54966), .ZN(n54291) );
  NAND2_X1 U14872 ( .A1(n52996), .A2(n53009), .ZN(n2585) );
  INV_X1 U14883 ( .I(n8513), .ZN(n55278) );
  NAND2_X1 U14888 ( .A1(n8203), .A2(n59040), .ZN(n55498) );
  INV_X1 U14889 ( .I(n54054), .ZN(n53402) );
  NAND2_X1 U14897 ( .A1(n21982), .A2(n23784), .ZN(n62328) );
  INV_X1 U14901 ( .I(n53876), .ZN(n51711) );
  NAND2_X1 U14903 ( .A1(n64813), .A2(n22807), .ZN(n55414) );
  NOR2_X1 U14904 ( .A1(n54858), .A2(n17935), .ZN(n55023) );
  INV_X1 U14910 ( .I(n52858), .ZN(n57062) );
  INV_X1 U14924 ( .I(n56978), .ZN(n64031) );
  NAND3_X1 U14925 ( .A1(n57060), .A2(n21079), .A3(n57061), .ZN(n57066) );
  NAND3_X1 U14926 ( .A1(n14307), .A2(n56586), .A3(n4634), .ZN(n56402) );
  INV_X1 U14931 ( .I(n51716), .ZN(n53016) );
  INV_X2 U14941 ( .I(n54807), .ZN(n54971) );
  INV_X1 U14942 ( .I(n54028), .ZN(n51865) );
  CLKBUF_X2 U14945 ( .I(n22114), .Z(n62515) );
  NAND2_X1 U14946 ( .A1(n2585), .A2(n53455), .ZN(n4078) );
  INV_X1 U14952 ( .I(n54107), .ZN(n51712) );
  CLKBUF_X4 U14959 ( .I(n13774), .Z(n3567) );
  AND2_X1 U14965 ( .A1(n55684), .A2(n18294), .Z(n52047) );
  NAND2_X1 U14968 ( .A1(n54451), .A2(n55016), .ZN(n54636) );
  NAND3_X1 U14971 ( .A1(n53589), .A2(n53590), .A3(n16427), .ZN(n53591) );
  INV_X1 U14973 ( .I(n53240), .ZN(n4020) );
  NAND2_X1 U14976 ( .A1(n52721), .A2(n56220), .ZN(n58382) );
  INV_X1 U14977 ( .I(n56592), .ZN(n64187) );
  BUF_X1 U14981 ( .I(n6737), .Z(n4835) );
  NAND2_X1 U14982 ( .A1(n56424), .A2(n56433), .ZN(n55703) );
  CLKBUF_X1 U14983 ( .I(n54107), .Z(n64076) );
  NOR2_X1 U14985 ( .A1(n52949), .A2(n24454), .ZN(n52950) );
  NOR2_X1 U14988 ( .A1(n55415), .A2(n54983), .ZN(n55413) );
  NAND2_X1 U14989 ( .A1(n57239), .A2(n56370), .ZN(n56375) );
  CLKBUF_X2 U14993 ( .I(n52861), .Z(n507) );
  CLKBUF_X1 U14994 ( .I(n55293), .Z(n60181) );
  INV_X1 U14998 ( .I(n55676), .ZN(n55668) );
  NOR2_X1 U14999 ( .A1(n55413), .A2(n55412), .ZN(n55421) );
  OAI22_X1 U15000 ( .A1(n24511), .A2(n24510), .B1(n54307), .B2(n25080), .ZN(
        n22232) );
  NOR2_X1 U15005 ( .A1(n53871), .A2(n54102), .ZN(n53877) );
  CLKBUF_X1 U15007 ( .I(n54325), .Z(n64681) );
  NAND3_X1 U15008 ( .A1(n62886), .A2(n57073), .A3(n52671), .ZN(n21225) );
  CLKBUF_X2 U15010 ( .I(n57048), .Z(n23563) );
  NAND3_X1 U15014 ( .A1(n57636), .A2(n50480), .A3(n53539), .ZN(n62085) );
  OAI21_X1 U15019 ( .A1(n64189), .A2(n64190), .B(n56592), .ZN(n64188) );
  INV_X1 U15022 ( .I(n52696), .ZN(n53242) );
  INV_X1 U15024 ( .I(n52893), .ZN(n58768) );
  AOI21_X1 U15025 ( .A1(n24454), .A2(n52492), .B(n14224), .ZN(n52119) );
  OAI21_X1 U15028 ( .A1(n53452), .A2(n21082), .B(n53451), .ZN(n63481) );
  INV_X1 U15029 ( .I(n13423), .ZN(n62077) );
  NAND2_X1 U15032 ( .A1(n52844), .A2(n52837), .ZN(n53603) );
  NOR2_X1 U15034 ( .A1(n53572), .A2(n533), .ZN(n64522) );
  OAI21_X1 U15035 ( .A1(n52659), .A2(n57063), .B(n21079), .ZN(n65188) );
  NAND3_X1 U15038 ( .A1(n53590), .A2(n53001), .A3(n16427), .ZN(n53002) );
  NAND2_X1 U15040 ( .A1(n54818), .A2(n6312), .ZN(n54692) );
  CLKBUF_X1 U15041 ( .I(n818), .Z(n59530) );
  NAND2_X1 U15043 ( .A1(n52792), .A2(n64028), .ZN(n17010) );
  NAND2_X1 U15044 ( .A1(n22804), .A2(n62263), .ZN(n15949) );
  AND3_X1 U15045 ( .A1(n26096), .A2(n54430), .A3(n54952), .Z(n869) );
  CLKBUF_X2 U15047 ( .I(n53241), .Z(n64424) );
  OAI21_X1 U15048 ( .A1(n57316), .A2(n58912), .B(n62074), .ZN(n22718) );
  NAND2_X1 U15053 ( .A1(n52220), .A2(n52219), .ZN(n63775) );
  NAND2_X1 U15058 ( .A1(n64733), .A2(n56399), .ZN(n12549) );
  NOR2_X1 U15059 ( .A1(n55441), .A2(n55440), .ZN(n711) );
  OAI21_X1 U15060 ( .A1(n22760), .A2(n57538), .B(n55024), .ZN(n54863) );
  CLKBUF_X1 U15065 ( .I(n52825), .Z(n64666) );
  NOR2_X1 U15066 ( .A1(n16080), .A2(n17543), .ZN(n17542) );
  NAND2_X1 U15072 ( .A1(n55253), .A2(n55254), .ZN(n62960) );
  OAI21_X1 U15073 ( .A1(n54020), .A2(n19402), .B(n19400), .ZN(n54031) );
  AOI21_X1 U15075 ( .A1(n52490), .A2(n20175), .B(n52491), .ZN(n52495) );
  NOR2_X1 U15080 ( .A1(n24729), .A2(n24696), .ZN(n56830) );
  CLKBUF_X4 U15086 ( .I(n54110), .Z(n23704) );
  OAI21_X1 U15089 ( .A1(n56558), .A2(n56658), .B(n59461), .ZN(n60574) );
  AOI21_X1 U15090 ( .A1(n53394), .A2(n53393), .B(n62741), .ZN(n13424) );
  NAND2_X1 U15104 ( .A1(n53400), .A2(n54049), .ZN(n53555) );
  AOI22_X1 U15105 ( .A1(n60334), .A2(n52874), .B1(n1602), .B2(n53239), .ZN(
        n59003) );
  NAND2_X1 U15113 ( .A1(n65188), .A2(n65187), .ZN(n52681) );
  NAND2_X1 U15116 ( .A1(n51963), .A2(n55684), .ZN(n17834) );
  OAI21_X1 U15119 ( .A1(n4895), .A2(n22064), .B(n59530), .ZN(n9650) );
  INV_X1 U15127 ( .I(n25172), .ZN(n54583) );
  NOR2_X1 U15129 ( .A1(n26151), .A2(n26155), .ZN(n15204) );
  NOR2_X1 U15131 ( .A1(n13792), .A2(n57367), .ZN(n13790) );
  NAND2_X1 U15133 ( .A1(n63858), .A2(n20696), .ZN(n56645) );
  NOR2_X1 U15135 ( .A1(n10507), .A2(n21879), .ZN(n64872) );
  INV_X1 U15136 ( .I(n56868), .ZN(n64246) );
  OAI21_X1 U15137 ( .A1(n56350), .A2(n56342), .B(n56349), .ZN(n11145) );
  INV_X1 U15139 ( .I(n54577), .ZN(n25764) );
  NAND2_X1 U15140 ( .A1(n53322), .A2(n53355), .ZN(n53362) );
  NAND3_X1 U15150 ( .A1(n1281), .A2(n22980), .A3(n19080), .ZN(n53067) );
  NAND2_X1 U15155 ( .A1(n22933), .A2(n21403), .ZN(n55822) );
  NAND3_X1 U15156 ( .A1(n53507), .A2(n53501), .A3(n25789), .ZN(n60796) );
  NAND4_X1 U15158 ( .A1(n23920), .A2(n21859), .A3(n17795), .A4(n21860), .ZN(
        n56463) );
  AOI21_X1 U15165 ( .A1(n55384), .A2(n60974), .B(n8261), .ZN(n24670) );
  CLKBUF_X2 U15166 ( .I(n23538), .Z(n58277) );
  CLKBUF_X4 U15167 ( .I(n57015), .Z(n63784) );
  INV_X1 U15169 ( .I(n53526), .ZN(n1581) );
  NAND2_X1 U15170 ( .A1(n16976), .A2(n55177), .ZN(n55180) );
  INV_X1 U15173 ( .I(n56867), .ZN(n56848) );
  NAND3_X1 U15174 ( .A1(n54402), .A2(n7138), .A3(n271), .ZN(n54387) );
  INV_X1 U15179 ( .I(n56189), .ZN(n1590) );
  INV_X1 U15181 ( .I(n53296), .ZN(n13239) );
  AOI21_X1 U15183 ( .A1(n53775), .A2(n53826), .B(n53774), .ZN(n53829) );
  AOI21_X1 U15187 ( .A1(n61057), .A2(n54742), .B(n54740), .ZN(n54661) );
  NOR2_X1 U15191 ( .A1(n23274), .A2(n53082), .ZN(n53093) );
  NAND2_X1 U15193 ( .A1(n13858), .A2(n60203), .ZN(n55891) );
  AOI21_X1 U15200 ( .A1(n15700), .A2(n8259), .B(n55642), .ZN(n8258) );
  NOR2_X1 U15202 ( .A1(n19492), .A2(n57967), .ZN(n54700) );
  OAI21_X1 U15203 ( .A1(n53311), .A2(n53310), .B(n53321), .ZN(n16828) );
  AOI21_X1 U15204 ( .A1(n56952), .A2(n63420), .B(n6902), .ZN(n56956) );
  CLKBUF_X2 U15207 ( .I(n53265), .Z(n62199) );
  OAI22_X1 U15223 ( .A1(n53127), .A2(n53167), .B1(n25484), .B2(n53128), .ZN(
        n53131) );
  NAND2_X1 U15225 ( .A1(n54727), .A2(n54767), .ZN(n54750) );
  INV_X1 U15226 ( .I(n56870), .ZN(n52728) );
  INV_X1 U15231 ( .I(n56350), .ZN(n56330) );
  NAND2_X1 U15232 ( .A1(n53335), .A2(n53369), .ZN(n214) );
  CLKBUF_X2 U15233 ( .I(n23074), .Z(n64833) );
  AOI21_X1 U15235 ( .A1(n1254), .A2(n14619), .B(n57132), .ZN(n4389) );
  CLKBUF_X4 U15238 ( .I(n59374), .Z(n23030) );
  NAND2_X1 U15239 ( .A1(n56108), .A2(n56092), .ZN(n56024) );
  CLKBUF_X2 U15241 ( .I(n54259), .Z(n22545) );
  NAND2_X1 U15248 ( .A1(n54380), .A2(n22401), .ZN(n54415) );
  NOR3_X1 U15251 ( .A1(n54187), .A2(n10480), .A3(n54170), .ZN(n54174) );
  INV_X1 U15253 ( .I(n56842), .ZN(n56888) );
  NAND2_X1 U15256 ( .A1(n53527), .A2(n53528), .ZN(n62094) );
  CLKBUF_X1 U15262 ( .I(n56104), .Z(n63699) );
  INV_X1 U15265 ( .I(n53305), .ZN(n53275) );
  CLKBUF_X4 U15267 ( .I(n55164), .Z(n11353) );
  AOI22_X1 U15269 ( .A1(n53055), .A2(n53114), .B1(n53111), .B2(n63006), .ZN(
        n53061) );
  CLKBUF_X4 U15273 ( .I(Key[15]), .Z(n53272) );
  OAI21_X1 U15279 ( .A1(n56874), .A2(n56870), .B(n64833), .ZN(n17359) );
  NAND3_X1 U15284 ( .A1(n56704), .A2(n56722), .A3(n56731), .ZN(n56711) );
  CLKBUF_X4 U15285 ( .I(Key[107]), .Z(n55242) );
  CLKBUF_X4 U15289 ( .I(Key[71]), .Z(n23455) );
  CLKBUF_X2 U15301 ( .I(n13306), .Z(n19793) );
  NAND2_X1 U15312 ( .A1(n38684), .A2(n20180), .ZN(n61751) );
  CLKBUF_X4 U15314 ( .I(n25772), .Z(n18300) );
  CLKBUF_X2 U15319 ( .I(n18401), .Z(n18402) );
  INV_X2 U15323 ( .I(n18401), .ZN(n21159) );
  INV_X1 U15324 ( .I(n30193), .ZN(n1846) );
  XNOR2_X1 U15325 ( .A1(n50028), .A2(n50027), .ZN(n61754) );
  OR3_X2 U15327 ( .A1(n14062), .A2(n1556), .A3(n29779), .Z(n61755) );
  OR2_X1 U15329 ( .A1(n41895), .A2(n2247), .Z(n61757) );
  AND2_X1 U15336 ( .A1(n59957), .A2(n59956), .Z(n61758) );
  OR3_X2 U15337 ( .A1(n49221), .A2(n16595), .A3(n6314), .Z(n61762) );
  OR2_X1 U15339 ( .A1(n19973), .A2(n24063), .Z(n61763) );
  AND3_X1 U15341 ( .A1(n24063), .A2(n9065), .A3(n61293), .Z(n61765) );
  OR2_X2 U15344 ( .A1(n22431), .A2(n3856), .Z(n61770) );
  OR2_X1 U15345 ( .A1(n51462), .A2(n52854), .Z(n61772) );
  XNOR2_X1 U15351 ( .A1(n20228), .A2(n62324), .ZN(n61775) );
  OR2_X1 U15359 ( .A1(n43191), .A2(n64330), .Z(n61778) );
  AND2_X1 U15360 ( .A1(n48101), .A2(n62290), .Z(n61779) );
  AND2_X1 U15364 ( .A1(n28562), .A2(n40), .Z(n61781) );
  AND2_X1 U15371 ( .A1(n37363), .A2(n4969), .Z(n61782) );
  OR2_X2 U15380 ( .A1(n25247), .A2(n20552), .Z(n61785) );
  AND2_X2 U15385 ( .A1(n56564), .A2(n56282), .Z(n61787) );
  OR2_X1 U15392 ( .A1(n15206), .A2(n15211), .Z(n61788) );
  AND2_X1 U15394 ( .A1(n559), .A2(n35799), .Z(n61789) );
  XNOR2_X1 U15395 ( .A1(n6363), .A2(n51727), .ZN(n61790) );
  XNOR2_X1 U15396 ( .A1(n62487), .A2(n61949), .ZN(n61791) );
  AND2_X1 U15400 ( .A1(n35665), .A2(n57732), .Z(n61793) );
  OR2_X2 U15404 ( .A1(n43437), .A2(n43449), .Z(n61794) );
  AND2_X2 U15407 ( .A1(n21409), .A2(n24256), .Z(n61795) );
  AND2_X1 U15414 ( .A1(n2325), .A2(n41877), .Z(n61796) );
  AND2_X1 U15431 ( .A1(n51185), .A2(n56586), .Z(n61797) );
  AND2_X1 U15439 ( .A1(n21218), .A2(n21311), .Z(n61799) );
  CLKBUF_X2 U15443 ( .I(n49548), .Z(n22571) );
  AND3_X2 U15457 ( .A1(n32149), .A2(n5807), .A3(n61574), .Z(n61801) );
  XNOR2_X1 U15458 ( .A1(n61099), .A2(n8234), .ZN(n61802) );
  AND2_X1 U15459 ( .A1(n37352), .A2(n36287), .Z(n61803) );
  AND2_X1 U15464 ( .A1(n16749), .A2(n40349), .Z(n61804) );
  OR2_X1 U15465 ( .A1(n6243), .A2(n63200), .Z(n61806) );
  XNOR2_X1 U15468 ( .A1(n10896), .A2(n51548), .ZN(n61807) );
  AND2_X1 U15470 ( .A1(n60520), .A2(n49918), .Z(n61808) );
  OR3_X1 U15474 ( .A1(n12859), .A2(n34626), .A3(n20279), .Z(n61809) );
  OR2_X1 U15476 ( .A1(n35764), .A2(n21096), .Z(n61810) );
  AND2_X2 U15477 ( .A1(n60054), .A2(n30895), .Z(n61811) );
  AND2_X2 U15479 ( .A1(n8305), .A2(n7950), .Z(n61812) );
  AND2_X1 U15482 ( .A1(n43353), .A2(n23151), .Z(n61813) );
  OR3_X1 U15484 ( .A1(n49606), .A2(n49605), .A3(n19003), .Z(n61814) );
  NOR2_X1 U15485 ( .A1(n7318), .A2(n48594), .ZN(n61815) );
  AND3_X1 U15486 ( .A1(n34120), .A2(n31722), .A3(n33944), .Z(n61818) );
  AND2_X2 U15487 ( .A1(n29306), .A2(n29295), .Z(n61820) );
  AND2_X1 U15488 ( .A1(n55347), .A2(n55362), .Z(n61822) );
  AND2_X1 U15494 ( .A1(n37068), .A2(n4798), .Z(n61824) );
  AND2_X1 U15495 ( .A1(n40925), .A2(n40924), .Z(n61826) );
  AND2_X1 U15504 ( .A1(n29516), .A2(n29856), .Z(n61827) );
  NOR2_X1 U15509 ( .A1(n52123), .A2(n55908), .ZN(n61828) );
  OR2_X2 U15530 ( .A1(n5323), .A2(n22782), .Z(n61829) );
  OR2_X2 U15535 ( .A1(n35994), .A2(n35096), .Z(n61831) );
  OR2_X2 U15536 ( .A1(n36764), .A2(n3622), .Z(n61832) );
  XNOR2_X1 U15542 ( .A1(n16202), .A2(n16196), .ZN(n61834) );
  AND2_X1 U15544 ( .A1(n63610), .A2(n6575), .Z(n61835) );
  AND2_X1 U15545 ( .A1(n56397), .A2(n64295), .Z(n61836) );
  XOR2_X1 U15552 ( .A1(n22195), .A2(n33041), .Z(n61837) );
  CLKBUF_X4 U15558 ( .I(Key[109]), .Z(n55340) );
  OR2_X1 U15563 ( .A1(n42451), .A2(n7094), .Z(n61838) );
  AND2_X1 U15571 ( .A1(n24454), .A2(n62763), .Z(n61840) );
  AND2_X1 U15578 ( .A1(n1535), .A2(n14669), .Z(n61841) );
  XNOR2_X1 U15581 ( .A1(n21009), .A2(n37180), .ZN(n61843) );
  INV_X1 U15586 ( .I(n15795), .ZN(n25837) );
  CLKBUF_X2 U15588 ( .I(n15795), .Z(n23145) );
  AND2_X1 U15594 ( .A1(n29040), .A2(n29039), .Z(n61844) );
  AND2_X1 U15598 ( .A1(n45672), .A2(n47256), .Z(n61845) );
  AND2_X2 U15603 ( .A1(n50215), .A2(n16765), .Z(n61846) );
  CLKBUF_X4 U15605 ( .I(n56616), .Z(n56697) );
  OR2_X1 U15609 ( .A1(n40933), .A2(n63303), .Z(n61847) );
  CLKBUF_X4 U15612 ( .I(n30979), .Z(n34613) );
  AND3_X1 U15617 ( .A1(n41417), .A2(n41418), .A3(n66), .Z(n61848) );
  AND2_X1 U15618 ( .A1(n31241), .A2(n31254), .Z(n61849) );
  OR3_X2 U15619 ( .A1(n1743), .A2(n38932), .A3(n10173), .Z(n61850) );
  AND3_X1 U15620 ( .A1(n35715), .A2(n35714), .A3(n35833), .Z(n61852) );
  OR2_X1 U15626 ( .A1(n15635), .A2(n502), .Z(n61853) );
  OR2_X1 U15629 ( .A1(n33391), .A2(n18884), .Z(n61854) );
  INV_X1 U15649 ( .I(n19621), .ZN(n64618) );
  OR2_X1 U15656 ( .A1(n34009), .A2(n59910), .Z(n61856) );
  INV_X1 U15660 ( .I(n33431), .ZN(n35026) );
  XNOR2_X1 U15661 ( .A1(n63213), .A2(n9108), .ZN(n61857) );
  AND2_X2 U15662 ( .A1(n1716), .A2(n42585), .Z(n61859) );
  CLKBUF_X4 U15669 ( .I(n36202), .Z(n2418) );
  OR2_X1 U15671 ( .A1(n47575), .A2(n47576), .Z(n61860) );
  AND2_X1 U15680 ( .A1(n58889), .A2(n47418), .Z(n61862) );
  AND2_X1 U15683 ( .A1(n19365), .A2(n42996), .Z(n61864) );
  AND2_X1 U15684 ( .A1(n56069), .A2(n56090), .Z(n61865) );
  OR2_X1 U15685 ( .A1(n45167), .A2(n49757), .Z(n61866) );
  AND2_X1 U15686 ( .A1(n60245), .A2(n63609), .Z(n61868) );
  OR2_X1 U15687 ( .A1(n42925), .A2(n42541), .Z(n61869) );
  AND2_X2 U15688 ( .A1(n19167), .A2(n54997), .Z(n61870) );
  CLKBUF_X4 U15701 ( .I(Key[115]), .Z(n55534) );
  OR2_X1 U15702 ( .A1(n138), .A2(n56961), .Z(n61872) );
  XNOR2_X1 U15705 ( .A1(n45105), .A2(n31595), .ZN(n61874) );
  NAND2_X1 U15706 ( .A1(n28301), .A2(n23636), .ZN(n61875) );
  CLKBUF_X4 U15707 ( .I(n20586), .Z(n8185) );
  OR2_X1 U15713 ( .A1(n64562), .A2(n9772), .Z(n61877) );
  AND2_X1 U15716 ( .A1(n1315), .A2(n31039), .Z(n61878) );
  AND2_X1 U15717 ( .A1(n36175), .A2(n36122), .Z(n61879) );
  AND2_X1 U15720 ( .A1(n38682), .A2(n60274), .Z(n61880) );
  OR2_X1 U15721 ( .A1(n34597), .A2(n62967), .Z(n61881) );
  XNOR2_X1 U15725 ( .A1(n5009), .A2(n22390), .ZN(n61883) );
  OR3_X1 U15726 ( .A1(n29593), .A2(n29076), .A3(n59268), .Z(n61884) );
  AND2_X1 U15739 ( .A1(n28034), .A2(n10537), .Z(n61886) );
  AND2_X2 U15742 ( .A1(n9865), .A2(n1562), .Z(n61888) );
  AND2_X1 U15743 ( .A1(n47572), .A2(n47900), .Z(n61889) );
  OR2_X2 U15745 ( .A1(n37126), .A2(n37125), .Z(n61890) );
  INV_X1 U15747 ( .I(n54300), .ZN(n63569) );
  OR2_X2 U15748 ( .A1(n24870), .A2(n8023), .Z(n61893) );
  INV_X1 U15749 ( .I(n43199), .ZN(n43509) );
  CLKBUF_X2 U15752 ( .I(n56599), .Z(n19151) );
  OR2_X2 U15753 ( .A1(n41702), .A2(n41568), .Z(n61894) );
  OR2_X2 U15754 ( .A1(n55416), .A2(n24075), .Z(n61895) );
  NAND2_X1 U15755 ( .A1(n61388), .A2(n11476), .ZN(n43222) );
  INV_X1 U15756 ( .I(n43222), .ZN(n63095) );
  INV_X1 U15757 ( .I(n48929), .ZN(n25065) );
  AND2_X2 U15760 ( .A1(n21409), .A2(n33993), .Z(n61896) );
  NAND3_X1 U15761 ( .A1(n29964), .A2(n30782), .A3(n30786), .ZN(n30777) );
  INV_X1 U15765 ( .I(n30777), .ZN(n62202) );
  OR2_X2 U15767 ( .A1(n29079), .A2(n22504), .Z(n61897) );
  INV_X1 U15769 ( .I(n34598), .ZN(n62967) );
  AND2_X2 U15771 ( .A1(n21512), .A2(n24196), .Z(n61900) );
  AND2_X1 U15772 ( .A1(n20013), .A2(n45611), .Z(n61901) );
  OR2_X2 U15773 ( .A1(n56599), .A2(n15536), .Z(n61902) );
  OR2_X1 U15776 ( .A1(n30262), .A2(n2310), .Z(n61903) );
  AND2_X1 U15778 ( .A1(n8770), .A2(n29943), .Z(n61905) );
  INV_X1 U15779 ( .I(n54790), .ZN(n63708) );
  INV_X2 U15781 ( .I(n64869), .ZN(n57398) );
  INV_X1 U15791 ( .I(n62656), .ZN(n41981) );
  NAND2_X1 U15794 ( .A1(n58572), .A2(n42355), .ZN(n62656) );
  AND2_X1 U15796 ( .A1(n41823), .A2(n41821), .Z(n61906) );
  AND2_X1 U15802 ( .A1(n7047), .A2(n34003), .Z(n61908) );
  INV_X1 U15804 ( .I(n64291), .ZN(n42026) );
  OR2_X2 U15809 ( .A1(n47851), .A2(n12725), .Z(n61909) );
  XNOR2_X1 U15810 ( .A1(n11970), .A2(n50633), .ZN(n61911) );
  INV_X1 U15814 ( .I(n62247), .ZN(n9986) );
  OR2_X2 U15815 ( .A1(n56414), .A2(n25413), .Z(n61914) );
  AND2_X1 U15816 ( .A1(n18508), .A2(n34786), .Z(n61915) );
  CLKBUF_X4 U15818 ( .I(n36220), .Z(n15034) );
  OR2_X1 U15819 ( .A1(n10358), .A2(n15809), .Z(n61917) );
  XNOR2_X1 U15822 ( .A1(Ciphertext[8]), .A2(Key[45]), .ZN(n61918) );
  OR2_X2 U15836 ( .A1(n52668), .A2(n52665), .Z(n61920) );
  AND2_X1 U15838 ( .A1(n45740), .A2(n19305), .Z(n61922) );
  AND4_X1 U15840 ( .A1(n16506), .A2(n16505), .A3(n35228), .A4(n16507), .Z(
        n61923) );
  NAND2_X1 U15841 ( .A1(n40472), .A2(n4968), .ZN(n61924) );
  INV_X1 U15843 ( .I(n16631), .ZN(n16630) );
  AND2_X2 U15845 ( .A1(n16489), .A2(n22200), .Z(n61925) );
  INV_X2 U15852 ( .I(n55474), .ZN(n55472) );
  XNOR2_X1 U15856 ( .A1(n8492), .A2(n31522), .ZN(n61926) );
  XNOR2_X1 U15861 ( .A1(n16821), .A2(n33261), .ZN(n61927) );
  AND2_X2 U15868 ( .A1(n24196), .A2(n8470), .Z(n61928) );
  CLKBUF_X1 U15869 ( .I(n29148), .Z(n65198) );
  OR2_X1 U15873 ( .A1(n7662), .A2(n37310), .Z(n61929) );
  CLKBUF_X1 U15874 ( .I(n15726), .Z(n8652) );
  INV_X2 U15875 ( .I(n31189), .ZN(n13444) );
  OR3_X2 U15877 ( .A1(n39933), .A2(n41854), .A3(n41280), .Z(n61930) );
  INV_X2 U15879 ( .I(n40842), .ZN(n41877) );
  XOR2_X1 U15882 ( .A1(n15377), .A2(n20386), .Z(n61932) );
  OR2_X2 U15885 ( .A1(n53755), .A2(n53728), .Z(n61933) );
  INV_X1 U15886 ( .I(n40661), .ZN(n1404) );
  OR3_X2 U15888 ( .A1(n18943), .A2(n18946), .A3(n61649), .Z(n61935) );
  XNOR2_X1 U15889 ( .A1(n31395), .A2(n31394), .ZN(n61938) );
  OR2_X1 U15893 ( .A1(n19289), .A2(n7253), .Z(n61939) );
  AND2_X2 U15902 ( .A1(n36453), .A2(n36443), .Z(n61940) );
  NAND2_X1 U15905 ( .A1(n30288), .A2(n23772), .ZN(n61942) );
  AND2_X1 U15909 ( .A1(n34383), .A2(n11182), .Z(n61943) );
  OR2_X2 U15915 ( .A1(n59013), .A2(n57509), .Z(n61944) );
  NOR2_X1 U15919 ( .A1(n13656), .A2(n3460), .ZN(n61945) );
  CLKBUF_X4 U15926 ( .I(n37583), .Z(n39625) );
  XNOR2_X1 U15928 ( .A1(n32668), .A2(n31739), .ZN(n61946) );
  INV_X1 U15934 ( .I(n31026), .ZN(n19610) );
  INV_X1 U15935 ( .I(n43429), .ZN(n63212) );
  CLKBUF_X4 U15940 ( .I(n19010), .Z(n57199) );
  XOR2_X1 U15951 ( .A1(n15189), .A2(n16423), .Z(n61947) );
  BUF_X2 U15957 ( .I(n16423), .Z(n16346) );
  AND3_X2 U15960 ( .A1(n33532), .A2(n33118), .A3(n14330), .Z(n61948) );
  CLKBUF_X2 U15980 ( .I(n37755), .Z(n40578) );
  CLKBUF_X2 U15986 ( .I(n64387), .Z(n61028) );
  INV_X1 U15989 ( .I(n64387), .ZN(n63319) );
  OR2_X2 U15994 ( .A1(n15411), .A2(n6337), .Z(n61949) );
  CLKBUF_X4 U15996 ( .I(n35710), .Z(n24089) );
  INV_X1 U16000 ( .I(n25020), .ZN(n40728) );
  INV_X1 U16007 ( .I(n36671), .ZN(n36664) );
  CLKBUF_X4 U16013 ( .I(n40947), .Z(n22593) );
  OR2_X2 U16015 ( .A1(n64367), .A2(n11460), .Z(n61950) );
  INV_X2 U16017 ( .I(n57925), .ZN(n41412) );
  AND2_X2 U16018 ( .A1(n43657), .A2(n43242), .Z(n61951) );
  XNOR2_X1 U16030 ( .A1(n39291), .A2(n33529), .ZN(n61953) );
  AND3_X1 U16036 ( .A1(n41542), .A2(n426), .A3(n57179), .Z(n61954) );
  INV_X1 U16050 ( .I(n47868), .ZN(n47674) );
  OR2_X2 U16051 ( .A1(n64125), .A2(n9643), .Z(n61955) );
  XOR2_X1 U16057 ( .A1(n61665), .A2(n20694), .Z(n61957) );
  XNOR2_X1 U16062 ( .A1(n40554), .A2(n45823), .ZN(n61958) );
  OR2_X1 U16063 ( .A1(n49768), .A2(n49783), .Z(n61959) );
  XNOR2_X1 U16064 ( .A1(n46495), .A2(n43453), .ZN(n61960) );
  AND2_X2 U16072 ( .A1(n65074), .A2(n18357), .Z(n61961) );
  BUF_X2 U16079 ( .I(n53161), .Z(n2037) );
  AND2_X1 U16082 ( .A1(n36399), .A2(n36398), .Z(n61962) );
  CLKBUF_X1 U16088 ( .I(n44779), .Z(n10512) );
  CLKBUF_X4 U16094 ( .I(n1487), .Z(n63926) );
  INV_X2 U16097 ( .I(n3400), .ZN(n24509) );
  INV_X2 U16106 ( .I(n1237), .ZN(n14884) );
  AND2_X2 U16112 ( .A1(n23163), .A2(n56522), .Z(n61964) );
  CLKBUF_X2 U16113 ( .I(n23533), .Z(n21092) );
  XNOR2_X1 U16124 ( .A1(n13257), .A2(n57276), .ZN(n61965) );
  INV_X1 U16128 ( .I(n56600), .ZN(n56984) );
  INV_X1 U16129 ( .I(n6704), .ZN(n64335) );
  NAND2_X1 U16136 ( .A1(n15020), .A2(n63485), .ZN(n18228) );
  NOR2_X1 U16137 ( .A1(n47622), .A2(n60423), .ZN(n61968) );
  INV_X2 U16140 ( .I(n48294), .ZN(n20461) );
  CLKBUF_X2 U16147 ( .I(n48294), .Z(n7990) );
  CLKBUF_X4 U16153 ( .I(n51918), .Z(n17336) );
  OR2_X1 U16164 ( .A1(n9102), .A2(n1233), .Z(n61969) );
  AND3_X1 U16167 ( .A1(n54965), .A2(n54970), .A3(n54973), .Z(n61970) );
  AND2_X2 U16187 ( .A1(n56817), .A2(n51461), .Z(n61971) );
  BUF_X1 U16196 ( .I(n10823), .Z(n6722) );
  INV_X1 U16203 ( .I(n10823), .ZN(n64340) );
  NAND2_X2 U16207 ( .A1(n59858), .A2(n61730), .ZN(n6943) );
  NOR2_X1 U16231 ( .A1(n53233), .A2(n53232), .ZN(n52868) );
  AOI22_X2 U16237 ( .A1(n33130), .A2(n6842), .B1(n6979), .B2(n35675), .ZN(
        n33087) );
  NOR2_X2 U16241 ( .A1(n12506), .A2(n17401), .ZN(n35675) );
  NAND2_X2 U16242 ( .A1(n62855), .A2(n61972), .ZN(n59731) );
  NAND2_X2 U16247 ( .A1(n61973), .A2(n18399), .ZN(n43382) );
  NAND2_X2 U16250 ( .A1(n56401), .A2(n20737), .ZN(n56579) );
  NOR2_X2 U16251 ( .A1(n14307), .A2(n56403), .ZN(n56401) );
  NOR3_X2 U16259 ( .A1(n61974), .A2(n24214), .A3(n46022), .ZN(n21621) );
  NOR3_X2 U16260 ( .A1(n12750), .A2(n12751), .A3(n64533), .ZN(n18410) );
  XOR2_X1 U16269 ( .A1(n61603), .A2(n17733), .Z(n64501) );
  INV_X1 U16270 ( .I(n56225), .ZN(n12026) );
  NAND2_X2 U16271 ( .A1(n1237), .A2(n12028), .ZN(n56225) );
  NAND3_X2 U16274 ( .A1(n12843), .A2(n12841), .A3(n26101), .ZN(n4234) );
  XOR2_X1 U16281 ( .A1(n37873), .A2(n10351), .Z(n9967) );
  NOR2_X2 U16283 ( .A1(n61975), .A2(n28393), .ZN(n28426) );
  NAND4_X2 U16286 ( .A1(n28390), .A2(n28391), .A3(n63150), .A4(n28388), .ZN(
        n61975) );
  NAND2_X1 U16287 ( .A1(n61977), .A2(n4024), .ZN(n65132) );
  NOR2_X1 U16289 ( .A1(n4023), .A2(n52869), .ZN(n61977) );
  NAND2_X2 U16290 ( .A1(n62155), .A2(n7489), .ZN(n3087) );
  NOR2_X2 U16294 ( .A1(n59185), .A2(n16840), .ZN(n26000) );
  NAND2_X2 U16299 ( .A1(n61978), .A2(n10853), .ZN(n25788) );
  NOR2_X2 U16301 ( .A1(n63446), .A2(n60318), .ZN(n61978) );
  INV_X8 U16309 ( .I(n11395), .ZN(n29516) );
  NAND2_X2 U16310 ( .A1(n64664), .A2(n20195), .ZN(n11395) );
  NOR2_X2 U16314 ( .A1(n22547), .A2(n61979), .ZN(n22546) );
  AOI21_X2 U16316 ( .A1(n64880), .A2(n64881), .B(n11708), .ZN(n61979) );
  BUF_X2 U16337 ( .I(n44578), .Z(n22650) );
  XOR2_X1 U16340 ( .A1(n36298), .A2(n19314), .Z(n26044) );
  NAND3_X2 U16344 ( .A1(n58985), .A2(n33333), .A3(n18071), .ZN(n36298) );
  NOR2_X2 U16348 ( .A1(n49676), .A2(n5498), .ZN(n65253) );
  NAND2_X2 U16350 ( .A1(n58716), .A2(n18107), .ZN(n5498) );
  XOR2_X1 U16352 ( .A1(n43425), .A2(n1488), .Z(n44947) );
  NAND2_X2 U16355 ( .A1(n2749), .A2(n62177), .ZN(n43425) );
  AND2_X1 U16357 ( .A1(n5674), .A2(n5673), .Z(n63675) );
  XOR2_X1 U16360 ( .A1(n12608), .A2(n44478), .Z(n13261) );
  NAND2_X2 U16363 ( .A1(n12901), .A2(n13262), .ZN(n12608) );
  INV_X2 U16373 ( .I(n42826), .ZN(n6706) );
  NAND2_X2 U16375 ( .A1(n6707), .A2(n41229), .ZN(n42826) );
  NOR2_X2 U16376 ( .A1(n57557), .A2(n12961), .ZN(n64517) );
  NOR2_X2 U16377 ( .A1(n61981), .A2(n40227), .ZN(n40890) );
  NAND4_X2 U16385 ( .A1(n24667), .A2(n40226), .A3(n40225), .A4(n40293), .ZN(
        n61981) );
  NAND2_X1 U16388 ( .A1(n3599), .A2(n3614), .ZN(n64218) );
  NAND2_X2 U16390 ( .A1(n63440), .A2(n25823), .ZN(n64267) );
  XOR2_X1 U16391 ( .A1(n14372), .A2(n20621), .Z(n58954) );
  NAND2_X2 U16392 ( .A1(n193), .A2(n49587), .ZN(n20621) );
  INV_X1 U16394 ( .I(n47535), .ZN(n64121) );
  XOR2_X1 U16395 ( .A1(n44145), .A2(n8164), .Z(n45876) );
  XOR2_X1 U16399 ( .A1(n36298), .A2(n55876), .Z(n36685) );
  NAND2_X1 U16401 ( .A1(n56814), .A2(n58688), .ZN(n51568) );
  NAND2_X2 U16411 ( .A1(n25773), .A2(n49428), .ZN(n2956) );
  NAND3_X2 U16415 ( .A1(n49543), .A2(n61741), .A3(n7358), .ZN(n25773) );
  NAND3_X1 U16416 ( .A1(n8217), .A2(n58105), .A3(n33542), .ZN(n35202) );
  NOR2_X2 U16419 ( .A1(n6529), .A2(n15807), .ZN(n58105) );
  XOR2_X1 U16422 ( .A1(n61983), .A2(n63149), .Z(n63153) );
  XOR2_X1 U16423 ( .A1(n51289), .A2(n2801), .Z(n61983) );
  NOR2_X2 U16424 ( .A1(n21550), .A2(n48952), .ZN(n49776) );
  INV_X4 U16428 ( .I(n15243), .ZN(n22524) );
  AOI21_X2 U16430 ( .A1(n7598), .A2(n15243), .B(n64609), .ZN(n35906) );
  NOR2_X2 U16435 ( .A1(n21179), .A2(n14290), .ZN(n15243) );
  BUF_X2 U16436 ( .I(n48076), .Z(n64036) );
  INV_X2 U16439 ( .I(n61984), .ZN(n39957) );
  NAND2_X2 U16440 ( .A1(n8576), .A2(n5115), .ZN(n61984) );
  BUF_X2 U16445 ( .I(n56803), .Z(n60851) );
  NAND2_X2 U16449 ( .A1(n25412), .A2(n62353), .ZN(n65228) );
  NAND3_X1 U16454 ( .A1(n47833), .A2(n62424), .A3(n60881), .ZN(n57529) );
  NAND3_X2 U16459 ( .A1(n26473), .A2(n26475), .A3(n61985), .ZN(n30810) );
  BUF_X8 U16460 ( .I(n40994), .Z(n61986) );
  NAND3_X1 U16462 ( .A1(n42360), .A2(n63828), .A3(n1694), .ZN(n41985) );
  XOR2_X1 U16466 ( .A1(n61987), .A2(n57441), .Z(n58111) );
  XOR2_X1 U16478 ( .A1(n33289), .A2(n62694), .Z(n61987) );
  INV_X2 U16481 ( .I(n6324), .ZN(n45129) );
  XOR2_X1 U16483 ( .A1(n61988), .A2(n63279), .Z(n6324) );
  XOR2_X1 U16484 ( .A1(n38487), .A2(n61989), .Z(n37418) );
  XOR2_X1 U16491 ( .A1(n20684), .A2(n22487), .Z(n61989) );
  NOR2_X2 U16492 ( .A1(n23313), .A2(n23812), .ZN(n33597) );
  NAND2_X1 U16496 ( .A1(n54537), .A2(n18422), .ZN(n54525) );
  INV_X4 U16499 ( .I(n49910), .ZN(n25812) );
  XOR2_X1 U16501 ( .A1(n57481), .A2(n26211), .Z(n3400) );
  AOI22_X2 U16502 ( .A1(n55799), .A2(n61990), .B1(n55800), .B2(n55797), .ZN(
        n55808) );
  NOR2_X1 U16503 ( .A1(n55795), .A2(n55794), .ZN(n61990) );
  NAND3_X2 U16506 ( .A1(n16343), .A2(n61991), .A3(n16344), .ZN(n16342) );
  NAND2_X1 U16508 ( .A1(n55711), .A2(n55712), .ZN(n61991) );
  XOR2_X1 U16512 ( .A1(n33889), .A2(n60259), .Z(n5417) );
  NAND2_X2 U16514 ( .A1(n58498), .A2(n6228), .ZN(n33889) );
  NAND2_X2 U16517 ( .A1(n41158), .A2(n1306), .ZN(n6791) );
  NAND2_X2 U16519 ( .A1(n20897), .A2(n48460), .ZN(n14521) );
  AND2_X1 U16523 ( .A1(n3652), .A2(n25962), .Z(n65100) );
  NAND2_X1 U16527 ( .A1(n52940), .A2(n62280), .ZN(n59043) );
  NAND3_X2 U16538 ( .A1(n5246), .A2(n47367), .A3(n16486), .ZN(n17319) );
  NAND3_X2 U16545 ( .A1(n48676), .A2(n12829), .A3(n57467), .ZN(n8380) );
  NAND3_X2 U16546 ( .A1(n14370), .A2(n14365), .A3(n62496), .ZN(n48676) );
  XOR2_X1 U16555 ( .A1(n50879), .A2(n52530), .Z(n9038) );
  XOR2_X1 U16558 ( .A1(n16641), .A2(n51017), .Z(n50879) );
  NAND2_X2 U16566 ( .A1(n7668), .A2(n60865), .ZN(n55164) );
  NOR3_X2 U16567 ( .A1(n62407), .A2(n48470), .A3(n48469), .ZN(n5917) );
  BUF_X2 U16570 ( .I(n26671), .Z(n61992) );
  AOI22_X1 U16571 ( .A1(n22956), .A2(n27433), .B1(n22810), .B2(n64445), .ZN(
        n26668) );
  XOR2_X1 U16579 ( .A1(n62987), .A2(n7343), .Z(n6643) );
  XOR2_X1 U16580 ( .A1(n22678), .A2(n52207), .Z(n62987) );
  BUF_X2 U16582 ( .I(n40296), .Z(n61994) );
  NAND2_X2 U16589 ( .A1(n61995), .A2(n62661), .ZN(n63683) );
  NAND3_X2 U16592 ( .A1(n64778), .A2(n50803), .A3(n20765), .ZN(n50807) );
  XOR2_X1 U16594 ( .A1(n61997), .A2(n46381), .Z(n46382) );
  XOR2_X1 U16597 ( .A1(n13938), .A2(n9463), .Z(n61997) );
  NAND3_X1 U16601 ( .A1(n50046), .A2(n48942), .A3(n13925), .ZN(n62531) );
  NOR3_X2 U16604 ( .A1(n34899), .A2(n64312), .A3(n61998), .ZN(n37549) );
  XOR2_X1 U16608 ( .A1(n46392), .A2(n46283), .Z(n13173) );
  NAND3_X2 U16609 ( .A1(n43064), .A2(n43063), .A3(n43062), .ZN(n46392) );
  NOR3_X1 U16619 ( .A1(n60122), .A2(n23036), .A3(n34196), .ZN(n10933) );
  XOR2_X1 U16621 ( .A1(n6117), .A2(n64092), .Z(n6116) );
  XOR2_X1 U16623 ( .A1(n32327), .A2(n26038), .Z(n7352) );
  NAND3_X2 U16625 ( .A1(n30662), .A2(n26040), .A3(n22998), .ZN(n32327) );
  XOR2_X1 U16629 ( .A1(n62000), .A2(n45024), .Z(n60328) );
  XOR2_X1 U16631 ( .A1(n3416), .A2(n1677), .Z(n45024) );
  XOR2_X1 U16635 ( .A1(n4243), .A2(n61999), .Z(n2970) );
  XOR2_X1 U16640 ( .A1(n4244), .A2(n38306), .Z(n61999) );
  NAND2_X1 U16643 ( .A1(n55930), .A2(n10185), .ZN(n63694) );
  XOR2_X1 U16647 ( .A1(n45022), .A2(n65250), .Z(n62000) );
  NOR2_X2 U16650 ( .A1(n56084), .A2(n63023), .ZN(n56117) );
  XOR2_X1 U16652 ( .A1(n2183), .A2(n2185), .Z(n2182) );
  BUF_X2 U16656 ( .I(n43439), .Z(n62001) );
  NAND2_X2 U16663 ( .A1(n45959), .A2(n62002), .ZN(n63692) );
  NOR2_X2 U16666 ( .A1(n62004), .A2(n62003), .ZN(n62002) );
  XOR2_X1 U16667 ( .A1(n50992), .A2(n50991), .Z(n64513) );
  AOI21_X2 U16673 ( .A1(n62007), .A2(n62006), .B(n49799), .ZN(n58886) );
  INV_X4 U16686 ( .I(n57184), .ZN(n15245) );
  OR2_X2 U16688 ( .A1(n9265), .A2(n9264), .Z(n57184) );
  OAI21_X2 U16690 ( .A1(n10947), .A2(n47405), .B(n47852), .ZN(n47409) );
  AND2_X2 U16693 ( .A1(n13479), .A2(n4487), .Z(n6932) );
  NAND2_X2 U16696 ( .A1(n36226), .A2(n7656), .ZN(n64713) );
  NAND3_X2 U16697 ( .A1(n58534), .A2(n23101), .A3(n57383), .ZN(n63909) );
  NAND3_X2 U16702 ( .A1(n1024), .A2(n8657), .A3(n42194), .ZN(n8656) );
  OR2_X2 U16706 ( .A1(n15280), .A2(n4437), .Z(n43326) );
  NAND2_X2 U16713 ( .A1(n2754), .A2(n22805), .ZN(n50421) );
  BUF_X2 U16714 ( .I(n21915), .Z(n62010) );
  OAI21_X2 U16720 ( .A1(n24002), .A2(n10990), .B(n41350), .ZN(n43080) );
  NAND3_X1 U16725 ( .A1(n48776), .A2(n48914), .A3(n57425), .ZN(n48372) );
  XOR2_X1 U16728 ( .A1(n14588), .A2(n7602), .Z(n2576) );
  NAND2_X2 U16731 ( .A1(n5150), .A2(n25326), .ZN(n5149) );
  NAND2_X1 U16736 ( .A1(n53619), .A2(n53618), .ZN(n11870) );
  NOR2_X2 U16737 ( .A1(n23104), .A2(n62011), .ZN(n49107) );
  NAND3_X2 U16766 ( .A1(n45943), .A2(n45942), .A3(n45945), .ZN(n62011) );
  NAND2_X2 U16769 ( .A1(n64053), .A2(n49071), .ZN(n58722) );
  NAND2_X1 U16770 ( .A1(n4559), .A2(n55358), .ZN(n55359) );
  OAI21_X1 U16773 ( .A1(n62067), .A2(n62068), .B(n47577), .ZN(n2538) );
  XOR2_X1 U16774 ( .A1(n31902), .A2(n31982), .Z(n65195) );
  XOR2_X1 U16776 ( .A1(n62012), .A2(n17226), .Z(n10357) );
  XOR2_X1 U16779 ( .A1(n17230), .A2(n45862), .Z(n62012) );
  BUF_X4 U16789 ( .I(n24117), .Z(n16937) );
  XOR2_X1 U16790 ( .A1(n62013), .A2(n19079), .Z(n6739) );
  XOR2_X1 U16792 ( .A1(n6738), .A2(n50952), .Z(n62013) );
  XOR2_X1 U16795 ( .A1(n62014), .A2(n54143), .Z(Plaintext[55]) );
  NAND4_X2 U16796 ( .A1(n54141), .A2(n54138), .A3(n54139), .A4(n54140), .ZN(
        n62014) );
  NOR2_X2 U16804 ( .A1(n62015), .A2(n9962), .ZN(n23956) );
  NAND2_X1 U16811 ( .A1(n62448), .A2(n25903), .ZN(n62015) );
  OAI21_X2 U16812 ( .A1(n43277), .A2(n43276), .B(n24179), .ZN(n4721) );
  NAND3_X2 U16824 ( .A1(n11131), .A2(n11124), .A3(n11127), .ZN(n63695) );
  OR2_X1 U16841 ( .A1(n16957), .A2(n61522), .Z(n62016) );
  AOI21_X2 U16844 ( .A1(n30653), .A2(n62285), .B(n62017), .ZN(n30661) );
  INV_X2 U16846 ( .I(n3849), .ZN(n62017) );
  NAND2_X2 U16853 ( .A1(n30332), .A2(n8522), .ZN(n3849) );
  AND2_X1 U16857 ( .A1(n60940), .A2(n35384), .Z(n62281) );
  OAI21_X2 U16863 ( .A1(n53180), .A2(n53179), .B(n53539), .ZN(n20352) );
  NAND2_X2 U16865 ( .A1(n63128), .A2(n15935), .ZN(n53180) );
  XOR2_X1 U16868 ( .A1(n2722), .A2(n46305), .Z(n44120) );
  INV_X2 U16869 ( .I(n62019), .ZN(n6934) );
  XOR2_X1 U16870 ( .A1(n17158), .A2(n17157), .Z(n62019) );
  NOR2_X2 U16873 ( .A1(n23025), .A2(n60002), .ZN(n53589) );
  NOR3_X2 U16878 ( .A1(n15983), .A2(n62022), .A3(n62021), .ZN(n7035) );
  NAND3_X2 U16882 ( .A1(n43295), .A2(n43947), .A3(n15540), .ZN(n43951) );
  NAND2_X2 U16883 ( .A1(n42470), .A2(n62023), .ZN(n17750) );
  XNOR2_X1 U16888 ( .A1(n22535), .A2(n19821), .ZN(n62875) );
  NAND4_X2 U16889 ( .A1(n57111), .A2(n57112), .A3(n19195), .A4(n62024), .ZN(
        n62044) );
  AOI22_X2 U16895 ( .A1(n63356), .A2(n57116), .B1(n57132), .B2(n57104), .ZN(
        n62024) );
  XOR2_X1 U16901 ( .A1(n24037), .A2(n8767), .Z(n44162) );
  NAND2_X2 U16902 ( .A1(n11516), .A2(n63068), .ZN(n24037) );
  AND2_X1 U16907 ( .A1(n42016), .A2(n61745), .Z(n7031) );
  NAND2_X2 U16908 ( .A1(n7120), .A2(n62025), .ZN(n9224) );
  NAND3_X2 U16909 ( .A1(n64254), .A2(n9085), .A3(n33614), .ZN(n62025) );
  BUF_X2 U16910 ( .I(n6606), .Z(n62026) );
  NAND2_X2 U16911 ( .A1(n63803), .A2(n50314), .ZN(n8739) );
  NAND3_X1 U16914 ( .A1(n62104), .A2(n28902), .A3(n62103), .ZN(n27757) );
  NOR2_X2 U16917 ( .A1(n21532), .A2(n30216), .ZN(n13558) );
  NAND2_X1 U16932 ( .A1(n62028), .A2(n10193), .ZN(n45739) );
  NAND2_X2 U16940 ( .A1(n12249), .A2(n6747), .ZN(n10193) );
  INV_X2 U16943 ( .I(n45734), .ZN(n62028) );
  OR2_X1 U16949 ( .A1(n9286), .A2(n61236), .Z(n48205) );
  OAI21_X2 U16950 ( .A1(n42592), .A2(n42593), .B(n2884), .ZN(n42597) );
  NAND2_X2 U16951 ( .A1(n41796), .A2(n37535), .ZN(n2884) );
  XOR2_X1 U16952 ( .A1(n50037), .A2(n52414), .Z(n51722) );
  XOR2_X1 U16953 ( .A1(n52066), .A2(n58824), .Z(n50037) );
  NAND2_X1 U16955 ( .A1(n62390), .A2(n56672), .ZN(n8616) );
  NOR2_X2 U16957 ( .A1(n63619), .A2(n62029), .ZN(n9228) );
  XOR2_X1 U16958 ( .A1(n13544), .A2(n62030), .Z(n58286) );
  XOR2_X1 U16959 ( .A1(n21895), .A2(n46630), .Z(n62030) );
  NAND3_X2 U16963 ( .A1(n28298), .A2(n28296), .A3(n28297), .ZN(n5312) );
  NAND2_X2 U16964 ( .A1(n62032), .A2(n62031), .ZN(n37428) );
  NAND3_X2 U16968 ( .A1(n34244), .A2(n34242), .A3(n34243), .ZN(n62031) );
  AOI21_X2 U16977 ( .A1(n34236), .A2(n1801), .B(n62691), .ZN(n62032) );
  XOR2_X1 U16982 ( .A1(n8774), .A2(n8264), .Z(n3609) );
  NAND2_X2 U16983 ( .A1(n21252), .A2(n1343), .ZN(n35848) );
  NAND2_X2 U16993 ( .A1(n35229), .A2(n13487), .ZN(n21252) );
  XOR2_X1 U16996 ( .A1(n59306), .A2(n31809), .Z(n5798) );
  INV_X1 U17001 ( .I(n24405), .ZN(n62043) );
  INV_X2 U17002 ( .I(n41837), .ZN(n60947) );
  NOR2_X2 U17003 ( .A1(n41293), .A2(n41831), .ZN(n41837) );
  NAND2_X2 U17004 ( .A1(n55339), .A2(n15936), .ZN(n55373) );
  INV_X2 U17013 ( .I(n62034), .ZN(n15936) );
  NAND2_X2 U17015 ( .A1(n15245), .A2(n55385), .ZN(n62034) );
  BUF_X2 U17026 ( .I(n22717), .Z(n62035) );
  NAND2_X2 U17038 ( .A1(n11950), .A2(n11705), .ZN(n49832) );
  NOR2_X2 U17042 ( .A1(n35852), .A2(n37441), .ZN(n22427) );
  NOR2_X2 U17049 ( .A1(n2002), .A2(n10717), .ZN(n3620) );
  NAND2_X1 U17050 ( .A1(n36386), .A2(n58749), .ZN(n65244) );
  OAI21_X1 U17057 ( .A1(n40894), .A2(n40895), .B(n42362), .ZN(n40901) );
  AND2_X1 U17060 ( .A1(n17177), .A2(n52865), .Z(n64897) );
  OR2_X2 U17062 ( .A1(n11153), .A2(n5498), .Z(n49365) );
  XOR2_X1 U17063 ( .A1(n40922), .A2(n62873), .Z(n41142) );
  INV_X2 U17068 ( .I(n25686), .ZN(n62873) );
  XOR2_X1 U17069 ( .A1(n10278), .A2(n44238), .Z(n25686) );
  XOR2_X1 U17072 ( .A1(n62037), .A2(n38081), .Z(n38093) );
  XOR2_X1 U17074 ( .A1(n59977), .A2(n38402), .Z(n62037) );
  XOR2_X1 U17075 ( .A1(n8599), .A2(n16700), .Z(n8609) );
  XOR2_X1 U17076 ( .A1(n38080), .A2(n38079), .Z(n13225) );
  XOR2_X1 U17077 ( .A1(n37678), .A2(n24435), .Z(n38080) );
  NOR2_X2 U17078 ( .A1(n34466), .A2(n37615), .ZN(n22949) );
  NAND2_X2 U17085 ( .A1(n37616), .A2(n37620), .ZN(n37615) );
  INV_X2 U17086 ( .I(n32833), .ZN(n33992) );
  NAND2_X2 U17088 ( .A1(n18277), .A2(n33995), .ZN(n32833) );
  NOR2_X2 U17090 ( .A1(n5550), .A2(n55926), .ZN(n55920) );
  NAND2_X2 U17096 ( .A1(n24944), .A2(n8122), .ZN(n5550) );
  NAND2_X2 U17101 ( .A1(n57637), .A2(n47876), .ZN(n47880) );
  NOR2_X2 U17114 ( .A1(n44011), .A2(n62038), .ZN(n44013) );
  NAND4_X2 U17118 ( .A1(n44008), .A2(n44007), .A3(n44006), .A4(n44009), .ZN(
        n62038) );
  OAI21_X2 U17121 ( .A1(n62039), .A2(n9438), .B(n17962), .ZN(n44892) );
  NOR2_X1 U17122 ( .A1(n57521), .A2(n57522), .ZN(n62039) );
  NAND3_X1 U17128 ( .A1(n62040), .A2(n9189), .A3(n40514), .ZN(n63620) );
  NAND2_X1 U17132 ( .A1(n40513), .A2(n40512), .ZN(n62040) );
  AOI21_X1 U17135 ( .A1(n19955), .A2(n42548), .B(n19954), .ZN(n42550) );
  BUF_X2 U17139 ( .I(n4151), .Z(n62041) );
  NAND3_X1 U17143 ( .A1(n9266), .A2(n9267), .A3(n62042), .ZN(n9265) );
  NAND2_X1 U17147 ( .A1(n55291), .A2(n60181), .ZN(n62042) );
  OR2_X1 U17150 ( .A1(n25874), .A2(n42267), .Z(n40805) );
  XOR2_X1 U17151 ( .A1(n33174), .A2(n32467), .Z(n8667) );
  NAND2_X2 U17152 ( .A1(n29231), .A2(n29230), .ZN(n33174) );
  INV_X2 U17156 ( .I(n23283), .ZN(n14648) );
  XOR2_X1 U17157 ( .A1(n24279), .A2(n64607), .Z(n30977) );
  NAND4_X1 U17160 ( .A1(n53942), .A2(n53943), .A3(n53944), .A4(n53941), .ZN(
        n62060) );
  INV_X2 U17163 ( .I(n15160), .ZN(n42016) );
  NAND2_X1 U17165 ( .A1(n62043), .A2(n15160), .ZN(n42540) );
  NAND3_X2 U17166 ( .A1(n15899), .A2(n14800), .A3(n14801), .ZN(n15160) );
  XOR2_X1 U17167 ( .A1(n4871), .A2(n46147), .Z(n7882) );
  XOR2_X1 U17169 ( .A1(n45852), .A2(n43797), .Z(n46147) );
  XOR2_X1 U17172 ( .A1(n62044), .A2(n57113), .Z(Plaintext[187]) );
  AND2_X2 U17179 ( .A1(n17967), .A2(n13836), .Z(n6730) );
  NAND2_X2 U17182 ( .A1(n20971), .A2(n48007), .ZN(n49681) );
  NOR2_X2 U17186 ( .A1(n57864), .A2(n62488), .ZN(n11390) );
  NAND2_X2 U17189 ( .A1(n14934), .A2(n25147), .ZN(n57233) );
  NAND2_X2 U17198 ( .A1(n48845), .A2(n61673), .ZN(n47554) );
  NOR2_X2 U17201 ( .A1(n13688), .A2(n2691), .ZN(n24508) );
  NAND2_X2 U17202 ( .A1(n64752), .A2(n22318), .ZN(n13688) );
  AND2_X1 U17216 ( .A1(n7834), .A2(n62046), .Z(n21641) );
  NOR2_X2 U17221 ( .A1(n62047), .A2(n53426), .ZN(n53867) );
  NAND4_X2 U17226 ( .A1(n19301), .A2(n19280), .A3(n21574), .A4(n21573), .ZN(
        n57126) );
  NOR2_X2 U17229 ( .A1(n34184), .A2(n62048), .ZN(n34203) );
  NAND4_X2 U17233 ( .A1(n34174), .A2(n34175), .A3(n25893), .A4(n34173), .ZN(
        n62048) );
  XOR2_X1 U17238 ( .A1(n31912), .A2(n30550), .Z(n6940) );
  AOI21_X2 U17239 ( .A1(n25293), .A2(n28715), .B(n62773), .ZN(n31912) );
  XOR2_X1 U17242 ( .A1(n24516), .A2(n10628), .Z(n25855) );
  XOR2_X1 U17248 ( .A1(n6456), .A2(n6454), .Z(n227) );
  XOR2_X1 U17256 ( .A1(n31641), .A2(n32342), .Z(n32271) );
  XOR2_X1 U17265 ( .A1(n32011), .A2(n22336), .Z(n32342) );
  INV_X1 U17267 ( .I(n26210), .ZN(n64738) );
  XOR2_X1 U17282 ( .A1(n38907), .A2(n39551), .Z(n24277) );
  NAND4_X2 U17289 ( .A1(n22404), .A2(n37232), .A3(n20646), .A4(n37231), .ZN(
        n38907) );
  NOR2_X2 U17291 ( .A1(n28710), .A2(n62049), .ZN(n25293) );
  NAND2_X2 U17296 ( .A1(n61905), .A2(n62050), .ZN(n62049) );
  NAND2_X2 U17300 ( .A1(n30658), .A2(n30415), .ZN(n62050) );
  NAND3_X2 U17306 ( .A1(n19748), .A2(n59389), .A3(n19743), .ZN(n15788) );
  AOI21_X2 U17308 ( .A1(n19750), .A2(n19752), .B(n59116), .ZN(n19748) );
  NAND2_X2 U17310 ( .A1(n10909), .A2(n17867), .ZN(n17866) );
  XOR2_X1 U17311 ( .A1(n4265), .A2(n50964), .Z(n59110) );
  NOR2_X2 U17313 ( .A1(n20603), .A2(n9504), .ZN(n43153) );
  INV_X1 U17329 ( .I(n12329), .ZN(n62221) );
  XOR2_X1 U17333 ( .A1(n62207), .A2(n18331), .Z(n44104) );
  XOR2_X1 U17345 ( .A1(n39766), .A2(n25409), .Z(n7265) );
  XOR2_X1 U17350 ( .A1(n37988), .A2(n37989), .Z(n39766) );
  NAND2_X1 U17354 ( .A1(n55955), .A2(n64187), .ZN(n64186) );
  NAND2_X1 U17356 ( .A1(n64188), .A2(n64186), .ZN(n658) );
  NOR2_X2 U17358 ( .A1(n40295), .A2(n40218), .ZN(n40029) );
  NAND2_X2 U17359 ( .A1(n62051), .A2(n30336), .ZN(n30833) );
  NAND2_X2 U17362 ( .A1(n19420), .A2(n42046), .ZN(n59694) );
  NOR3_X2 U17368 ( .A1(n19421), .A2(n22880), .A3(n42043), .ZN(n19420) );
  NAND2_X2 U17400 ( .A1(n15890), .A2(n40864), .ZN(n4607) );
  NAND2_X2 U17405 ( .A1(n25816), .A2(n41876), .ZN(n40864) );
  INV_X4 U17413 ( .I(n62784), .ZN(n26657) );
  XOR2_X1 U17417 ( .A1(n10363), .A2(n31804), .Z(n32045) );
  XOR2_X1 U17419 ( .A1(n61346), .A2(n31556), .Z(n10363) );
  OR2_X1 U17420 ( .A1(n30337), .A2(n30416), .Z(n62051) );
  XOR2_X1 U17429 ( .A1(n62052), .A2(n45261), .Z(n44450) );
  XOR2_X1 U17436 ( .A1(n44448), .A2(n44910), .Z(n62052) );
  XOR2_X1 U17439 ( .A1(n44991), .A2(n23067), .Z(n14328) );
  AOI21_X2 U17442 ( .A1(n41697), .A2(n40373), .B(n3905), .ZN(n44991) );
  XOR2_X1 U17448 ( .A1(n38188), .A2(n22048), .Z(n22047) );
  NAND3_X2 U17451 ( .A1(n36918), .A2(n36919), .A3(n36917), .ZN(n38188) );
  BUF_X2 U17457 ( .I(n57735), .Z(n62054) );
  NAND3_X2 U17460 ( .A1(n62055), .A2(n35824), .A3(n35823), .ZN(n61076) );
  OAI21_X2 U17468 ( .A1(n35815), .A2(n57337), .B(n35813), .ZN(n62055) );
  XOR2_X1 U17470 ( .A1(n52067), .A2(n18494), .Z(n17252) );
  XOR2_X1 U17477 ( .A1(n18493), .A2(n24787), .Z(n52067) );
  OR2_X1 U17481 ( .A1(n21400), .A2(n40839), .Z(n43735) );
  NOR3_X2 U17484 ( .A1(n13599), .A2(n13660), .A3(n62056), .ZN(n13659) );
  NAND4_X2 U17486 ( .A1(n10008), .A2(n53879), .A3(n64991), .A4(n53880), .ZN(
        n62056) );
  NAND3_X2 U17489 ( .A1(n42251), .A2(n41918), .A3(n61477), .ZN(n40786) );
  NAND3_X2 U17494 ( .A1(n62057), .A2(n26604), .A3(n12033), .ZN(n18758) );
  OAI21_X2 U17497 ( .A1(n26603), .A2(n26669), .B(n19122), .ZN(n62057) );
  OAI21_X1 U17499 ( .A1(n1610), .A2(n54310), .B(n54071), .ZN(n53849) );
  NAND3_X2 U17501 ( .A1(n64885), .A2(n61923), .A3(n63862), .ZN(n36595) );
  NAND3_X1 U17502 ( .A1(n47527), .A2(n47526), .A3(n47525), .ZN(n62219) );
  NAND2_X2 U17504 ( .A1(n60343), .A2(n64122), .ZN(n47527) );
  NOR2_X2 U17513 ( .A1(n49528), .A2(n63785), .ZN(n49531) );
  XOR2_X1 U17514 ( .A1(n3232), .A2(n46681), .Z(n45269) );
  XOR2_X1 U17515 ( .A1(n25244), .A2(n19926), .Z(n3232) );
  NOR2_X2 U17517 ( .A1(n27621), .A2(n27611), .ZN(n64445) );
  NAND3_X2 U17522 ( .A1(n20796), .A2(n63117), .A3(n62059), .ZN(n62529) );
  OAI21_X2 U17531 ( .A1(n17064), .A2(n42621), .B(n62997), .ZN(n62059) );
  NAND2_X2 U17532 ( .A1(n43438), .A2(n43437), .ZN(n41743) );
  XOR2_X1 U17539 ( .A1(n39307), .A2(n14228), .Z(n39357) );
  XOR2_X1 U17540 ( .A1(n62060), .A2(n53945), .Z(Plaintext[49]) );
  AOI21_X2 U17558 ( .A1(n29092), .A2(n28750), .B(n6475), .ZN(n6474) );
  NOR3_X2 U17559 ( .A1(n43048), .A2(n43049), .A3(n62061), .ZN(n43050) );
  OAI22_X2 U17562 ( .A1(n43044), .A2(n43045), .B1(n12962), .B2(n14051), .ZN(
        n62061) );
  NOR2_X2 U17563 ( .A1(n22726), .A2(n27980), .ZN(n27985) );
  NOR2_X2 U17564 ( .A1(n11590), .A2(n23472), .ZN(n6841) );
  NOR2_X2 U17581 ( .A1(n41120), .A2(n26182), .ZN(n23472) );
  NOR2_X2 U17588 ( .A1(n23112), .A2(n22384), .ZN(n11590) );
  XOR2_X1 U17590 ( .A1(n44820), .A2(n44731), .Z(n8462) );
  XOR2_X1 U17596 ( .A1(n8598), .A2(n8599), .Z(n44820) );
  NOR3_X2 U17597 ( .A1(n61954), .A2(n59998), .A3(n62062), .ZN(n2236) );
  NAND2_X2 U17598 ( .A1(n5044), .A2(n12717), .ZN(n62062) );
  XOR2_X1 U17599 ( .A1(n62063), .A2(n63941), .Z(n44821) );
  XOR2_X1 U17606 ( .A1(n23006), .A2(n23440), .Z(n62063) );
  INV_X2 U17608 ( .I(n62064), .ZN(n57452) );
  NOR2_X2 U17610 ( .A1(n18617), .A2(n20130), .ZN(n62064) );
  NAND2_X2 U17612 ( .A1(n20132), .A2(n20136), .ZN(n18617) );
  XOR2_X1 U17614 ( .A1(n62066), .A2(n62065), .Z(n4398) );
  INV_X2 U17615 ( .I(n4674), .ZN(n62065) );
  XOR2_X1 U17622 ( .A1(n46162), .A2(n46197), .Z(n62066) );
  XOR2_X1 U17624 ( .A1(n14967), .A2(n8179), .Z(n46093) );
  NOR2_X1 U17628 ( .A1(n13356), .A2(n47576), .ZN(n62067) );
  NOR2_X2 U17632 ( .A1(n47578), .A2(n47575), .ZN(n62068) );
  XOR2_X1 U17634 ( .A1(n17975), .A2(n62069), .Z(n63780) );
  XOR2_X1 U17635 ( .A1(n39578), .A2(n62070), .Z(n62069) );
  NAND3_X1 U17638 ( .A1(n65149), .A2(n53849), .A3(n61371), .ZN(n24265) );
  NAND2_X2 U17639 ( .A1(n35723), .A2(n23742), .ZN(n37211) );
  NAND2_X2 U17643 ( .A1(n62949), .A2(n35678), .ZN(n35723) );
  XOR2_X1 U17645 ( .A1(n15788), .A2(n51783), .Z(n64507) );
  NOR2_X2 U17648 ( .A1(n65199), .A2(n18717), .ZN(n42213) );
  NOR2_X2 U17654 ( .A1(n42095), .A2(n5971), .ZN(n62072) );
  AND2_X1 U17655 ( .A1(n22726), .A2(n8528), .Z(n8626) );
  NAND2_X2 U17663 ( .A1(n21720), .A2(n3617), .ZN(n22726) );
  XOR2_X1 U17666 ( .A1(n11539), .A2(n11538), .Z(n13205) );
  XOR2_X1 U17671 ( .A1(n44338), .A2(n15698), .Z(n61424) );
  NAND3_X2 U17682 ( .A1(n41016), .A2(n41014), .A3(n41015), .ZN(n41025) );
  NAND2_X2 U17686 ( .A1(n15117), .A2(n15118), .ZN(n18342) );
  INV_X2 U17688 ( .I(n53678), .ZN(n53658) );
  NAND2_X2 U17710 ( .A1(n53695), .A2(n62073), .ZN(n53678) );
  INV_X1 U17711 ( .I(n24244), .ZN(n62073) );
  NOR2_X2 U17720 ( .A1(n54317), .A2(n24509), .ZN(n62074) );
  NAND3_X2 U17721 ( .A1(n62075), .A2(n13424), .A3(n13425), .ZN(n53518) );
  XOR2_X1 U17726 ( .A1(n16960), .A2(n10095), .Z(n62089) );
  XOR2_X1 U17730 ( .A1(n5458), .A2(n23637), .Z(n63008) );
  NOR2_X2 U17732 ( .A1(n5461), .A2(n4839), .ZN(n5458) );
  NOR2_X2 U17733 ( .A1(n10629), .A2(n64950), .ZN(n30193) );
  NAND2_X2 U17735 ( .A1(n14796), .A2(n59115), .ZN(n64950) );
  OAI22_X2 U17737 ( .A1(n59255), .A2(n41035), .B1(n1400), .B2(n40517), .ZN(
        n8797) );
  INV_X2 U17742 ( .I(n21171), .ZN(n40517) );
  NAND3_X2 U17746 ( .A1(n62597), .A2(n61758), .A3(n62079), .ZN(n19806) );
  NOR2_X1 U17751 ( .A1(n62081), .A2(n62080), .ZN(n15624) );
  NOR2_X1 U17752 ( .A1(n30200), .A2(n2351), .ZN(n62080) );
  AOI22_X1 U17756 ( .A1(n34544), .A2(n34528), .B1(n34527), .B2(n22419), .ZN(
        n34543) );
  OAI21_X1 U17760 ( .A1(n27091), .A2(n27092), .B(n27090), .ZN(n27093) );
  XOR2_X1 U17761 ( .A1(n4354), .A2(n2567), .Z(n416) );
  BUF_X4 U17765 ( .I(n5055), .Z(n4526) );
  NOR2_X1 U17766 ( .A1(n60069), .A2(n63972), .ZN(n57494) );
  NAND2_X2 U17768 ( .A1(n921), .A2(n34755), .ZN(n24541) );
  NAND2_X2 U17785 ( .A1(n62401), .A2(n34753), .ZN(n921) );
  NAND3_X2 U17787 ( .A1(n12230), .A2(n12229), .A3(n62082), .ZN(n59185) );
  BUF_X2 U17790 ( .I(n15715), .Z(n62083) );
  BUF_X2 U17794 ( .I(n5626), .Z(n62084) );
  NAND2_X1 U17796 ( .A1(n44135), .A2(n64352), .ZN(n60544) );
  NAND2_X2 U17797 ( .A1(n50482), .A2(n62085), .ZN(n62242) );
  INV_X2 U17809 ( .I(n50039), .ZN(n62087) );
  NAND2_X2 U17811 ( .A1(n1487), .A2(n63043), .ZN(n2344) );
  XOR2_X1 U17816 ( .A1(n62089), .A2(n57704), .Z(n10870) );
  NAND2_X2 U17822 ( .A1(n57205), .A2(n61722), .ZN(n3847) );
  NOR2_X1 U17827 ( .A1(n57570), .A2(n48501), .ZN(n48526) );
  NOR2_X2 U17832 ( .A1(n1714), .A2(n61107), .ZN(n62546) );
  BUF_X2 U17837 ( .I(n19434), .Z(n62090) );
  XOR2_X1 U17838 ( .A1(n50178), .A2(n18891), .Z(n50179) );
  XOR2_X1 U17841 ( .A1(n13285), .A2(n51335), .Z(n50177) );
  XOR2_X1 U17847 ( .A1(n62091), .A2(n22212), .Z(n44362) );
  XOR2_X1 U17851 ( .A1(n13463), .A2(n55546), .Z(n62091) );
  OR2_X1 U17854 ( .A1(n2794), .A2(n30398), .Z(n64693) );
  NAND2_X2 U17871 ( .A1(n64713), .A2(n62092), .ZN(n7643) );
  XOR2_X1 U17872 ( .A1(n62093), .A2(n12379), .Z(n60228) );
  XOR2_X1 U17874 ( .A1(n2876), .A2(n22845), .Z(n62093) );
  XOR2_X1 U17882 ( .A1(n64117), .A2(n24731), .Z(n43877) );
  XOR2_X1 U17887 ( .A1(n1523), .A2(n6441), .Z(n8391) );
  NOR2_X2 U17896 ( .A1(n62984), .A2(n62983), .ZN(n1523) );
  NAND2_X1 U17901 ( .A1(n1161), .A2(n53526), .ZN(n62095) );
  XOR2_X1 U17904 ( .A1(n9011), .A2(n62096), .Z(n16747) );
  XOR2_X1 U17913 ( .A1(n14058), .A2(n6385), .Z(n62096) );
  NAND2_X2 U17919 ( .A1(n6247), .A2(n45715), .ZN(n46862) );
  NOR2_X2 U17920 ( .A1(n4086), .A2(n23759), .ZN(n45715) );
  OAI22_X2 U17926 ( .A1(n46987), .A2(n46978), .B1(n45747), .B2(n4380), .ZN(
        n47463) );
  XOR2_X1 U17930 ( .A1(n44680), .A2(n9256), .Z(n45747) );
  NAND3_X2 U17935 ( .A1(n62097), .A2(n41262), .A3(n23741), .ZN(n3064) );
  OAI21_X2 U17937 ( .A1(n41264), .A2(n61477), .B(n41263), .ZN(n62097) );
  NOR2_X2 U17940 ( .A1(n11243), .A2(n23348), .ZN(n39517) );
  NOR3_X2 U17942 ( .A1(n63855), .A2(n25055), .A3(n5561), .ZN(n5560) );
  NAND2_X2 U17943 ( .A1(n35655), .A2(n6829), .ZN(n35642) );
  NOR2_X2 U17946 ( .A1(n62098), .A2(n39956), .ZN(n42049) );
  NAND3_X2 U17950 ( .A1(n8244), .A2(n39955), .A3(n8243), .ZN(n62098) );
  AND2_X1 U17954 ( .A1(n43898), .A2(n2824), .Z(n43654) );
  NAND3_X1 U17956 ( .A1(n62843), .A2(n1148), .A3(n54081), .ZN(n54086) );
  NOR2_X1 U17958 ( .A1(n16076), .A2(n63239), .ZN(n63148) );
  NAND2_X2 U17960 ( .A1(n42130), .A2(n42129), .ZN(n42132) );
  XOR2_X1 U17969 ( .A1(n14730), .A2(n52568), .Z(n52436) );
  XOR2_X1 U17980 ( .A1(n17336), .A2(n58814), .Z(n14356) );
  XOR2_X1 U17981 ( .A1(n62100), .A2(n58841), .Z(n9180) );
  XOR2_X1 U17983 ( .A1(n60682), .A2(n31414), .Z(n62100) );
  XOR2_X1 U17985 ( .A1(n46577), .A2(n62101), .Z(n20516) );
  XOR2_X1 U17992 ( .A1(n11852), .A2(n1488), .Z(n62101) );
  NOR2_X2 U18002 ( .A1(n11513), .A2(n29122), .ZN(n13564) );
  XOR2_X1 U18014 ( .A1(n51080), .A2(n50519), .Z(n11208) );
  XOR2_X1 U18039 ( .A1(n51749), .A2(n51148), .Z(n51080) );
  AND2_X1 U18042 ( .A1(n41446), .A2(n41433), .Z(n39609) );
  XOR2_X1 U18048 ( .A1(n45325), .A2(n44897), .Z(n44607) );
  BUF_X2 U18053 ( .I(n51870), .Z(n62102) );
  INV_X2 U18056 ( .I(n6015), .ZN(n64631) );
  OAI22_X1 U18059 ( .A1(n17131), .A2(n39052), .B1(n39051), .B2(n13669), .ZN(
        n17130) );
  AND2_X2 U18061 ( .A1(n58205), .A2(n61716), .Z(n3646) );
  XOR2_X1 U18062 ( .A1(n5487), .A2(n62315), .Z(n14180) );
  XOR2_X1 U18065 ( .A1(n20021), .A2(n6300), .Z(n5487) );
  XOR2_X1 U18066 ( .A1(n19687), .A2(n15755), .Z(n62105) );
  NOR2_X2 U18069 ( .A1(n25356), .A2(n18418), .ZN(n40434) );
  NOR2_X2 U18071 ( .A1(n23933), .A2(n58823), .ZN(n62106) );
  NAND3_X2 U18072 ( .A1(n37858), .A2(n6489), .A3(n6490), .ZN(n22452) );
  INV_X1 U18076 ( .I(n40012), .ZN(n62510) );
  NOR2_X2 U18078 ( .A1(n41743), .A2(n42944), .ZN(n43450) );
  INV_X2 U18082 ( .I(n39998), .ZN(n62107) );
  XOR2_X1 U18085 ( .A1(n43425), .A2(n62108), .Z(n65078) );
  XOR2_X1 U18095 ( .A1(n44948), .A2(n24449), .Z(n62108) );
  NOR3_X1 U18097 ( .A1(n44407), .A2(n15469), .A3(n15472), .ZN(n65211) );
  NAND3_X2 U18111 ( .A1(n31610), .A2(n62109), .A3(n61899), .ZN(n19795) );
  NOR2_X2 U18116 ( .A1(n19922), .A2(n19464), .ZN(n62109) );
  BUF_X4 U18117 ( .I(n30480), .Z(n62647) );
  NOR2_X2 U18120 ( .A1(n62110), .A2(n44577), .ZN(n22872) );
  NOR2_X2 U18121 ( .A1(n10428), .A2(n1294), .ZN(n44705) );
  NAND2_X1 U18124 ( .A1(n64639), .A2(n61315), .ZN(n60280) );
  OAI21_X1 U18125 ( .A1(n62111), .A2(n1031), .B(n59067), .ZN(n6423) );
  NOR2_X1 U18127 ( .A1(n6901), .A2(n41548), .ZN(n62111) );
  NOR2_X2 U18129 ( .A1(n24069), .A2(n49910), .ZN(n47787) );
  NOR2_X2 U18130 ( .A1(n65249), .A2(n19631), .ZN(n19630) );
  INV_X2 U18132 ( .I(n4860), .ZN(n7079) );
  NAND2_X2 U18135 ( .A1(n17015), .A2(n4824), .ZN(n4860) );
  AOI21_X2 U18139 ( .A1(n13382), .A2(n27187), .B(n62112), .ZN(n7297) );
  OAI22_X2 U18141 ( .A1(n27580), .A2(n26656), .B1(n26657), .B2(n26658), .ZN(
        n62112) );
  XOR2_X1 U18143 ( .A1(n15087), .A2(n33146), .Z(n62472) );
  INV_X4 U18145 ( .I(n62216), .ZN(n10448) );
  XOR2_X1 U18146 ( .A1(n15003), .A2(n38757), .Z(n39756) );
  XOR2_X1 U18147 ( .A1(n62113), .A2(n54208), .Z(Plaintext[59]) );
  NAND4_X2 U18148 ( .A1(n13706), .A2(n13713), .A3(n57348), .A4(n13709), .ZN(
        n62113) );
  XOR2_X1 U18155 ( .A1(n18887), .A2(n45319), .Z(n10678) );
  NAND3_X2 U18157 ( .A1(n8193), .A2(n8188), .A3(n8190), .ZN(n18887) );
  NAND3_X2 U18160 ( .A1(n54001), .A2(n53992), .A3(n6168), .ZN(n53903) );
  INV_X1 U18161 ( .I(n62529), .ZN(n62442) );
  OAI21_X2 U18164 ( .A1(n15919), .A2(n18590), .B(n18589), .ZN(n62114) );
  NOR3_X2 U18171 ( .A1(n57979), .A2(n10107), .A3(n61869), .ZN(n44893) );
  NOR2_X1 U18173 ( .A1(n62116), .A2(n13716), .ZN(n64799) );
  NAND2_X1 U18180 ( .A1(n54190), .A2(n54189), .ZN(n62116) );
  XOR2_X1 U18182 ( .A1(n62117), .A2(n57096), .Z(Plaintext[186]) );
  NAND3_X1 U18184 ( .A1(n57094), .A2(n57095), .A3(n57093), .ZN(n62117) );
  XOR2_X1 U18185 ( .A1(n62118), .A2(n51809), .Z(n62545) );
  XOR2_X1 U18190 ( .A1(n51806), .A2(n63687), .Z(n62118) );
  XOR2_X1 U18193 ( .A1(n62183), .A2(n62119), .Z(n51805) );
  INV_X2 U18194 ( .I(n51508), .ZN(n62119) );
  NOR2_X2 U18196 ( .A1(n3387), .A2(n3386), .ZN(n62183) );
  BUF_X2 U18197 ( .I(n59374), .Z(n62120) );
  AOI22_X2 U18199 ( .A1(n62121), .A2(n48084), .B1(n48081), .B2(n23617), .ZN(
        n48091) );
  AOI21_X2 U18201 ( .A1(n21296), .A2(n21135), .B(n53848), .ZN(n54071) );
  NOR2_X1 U18202 ( .A1(n20857), .A2(n64433), .ZN(n63169) );
  XOR2_X1 U18203 ( .A1(n13664), .A2(n38911), .Z(n12980) );
  XOR2_X1 U18204 ( .A1(n15487), .A2(n52559), .Z(n21219) );
  XOR2_X1 U18205 ( .A1(n23696), .A2(n11884), .Z(n46570) );
  NAND3_X2 U18206 ( .A1(n2752), .A2(n62677), .A3(n2753), .ZN(n23696) );
  NAND2_X2 U18208 ( .A1(n62122), .A2(n62197), .ZN(n24436) );
  OAI21_X2 U18211 ( .A1(n36056), .A2(n36055), .B(n10086), .ZN(n62122) );
  NAND2_X2 U18218 ( .A1(n62345), .A2(n33592), .ZN(n24926) );
  BUF_X2 U18229 ( .I(n39950), .Z(n62123) );
  XOR2_X1 U18235 ( .A1(n51741), .A2(n57753), .Z(n26185) );
  NOR2_X2 U18240 ( .A1(n47337), .A2(n57754), .ZN(n51741) );
  INV_X2 U18241 ( .I(n62124), .ZN(n62689) );
  XOR2_X1 U18248 ( .A1(n60311), .A2(n6500), .Z(n62124) );
  NAND3_X2 U18250 ( .A1(n53011), .A2(n53012), .A3(n53013), .ZN(n58811) );
  NOR2_X2 U18251 ( .A1(n53230), .A2(n53010), .ZN(n53011) );
  NOR2_X1 U18252 ( .A1(n36331), .A2(n35914), .ZN(n63598) );
  NAND2_X2 U18254 ( .A1(n53587), .A2(n58300), .ZN(n16708) );
  XOR2_X1 U18256 ( .A1(n21034), .A2(n63213), .Z(n65219) );
  XOR2_X1 U18263 ( .A1(n62850), .A2(n31004), .Z(n21034) );
  XOR2_X1 U18269 ( .A1(n8030), .A2(n24891), .Z(n24890) );
  NAND2_X2 U18270 ( .A1(n58128), .A2(n62125), .ZN(n9482) );
  NOR3_X2 U18280 ( .A1(n11435), .A2(n9812), .A3(n11434), .ZN(n62125) );
  XOR2_X1 U18281 ( .A1(n62126), .A2(n20580), .Z(n63895) );
  XOR2_X1 U18282 ( .A1(n18954), .A2(n18955), .Z(n62126) );
  XOR2_X1 U18293 ( .A1(n62127), .A2(n14871), .Z(n14872) );
  XOR2_X1 U18294 ( .A1(n11956), .A2(n7961), .Z(n62127) );
  XOR2_X1 U18295 ( .A1(n32737), .A2(n59274), .Z(n12019) );
  XOR2_X1 U18296 ( .A1(n13638), .A2(n31456), .Z(n59274) );
  XOR2_X1 U18297 ( .A1(n52177), .A2(n23371), .Z(n63659) );
  NAND3_X2 U18306 ( .A1(n61682), .A2(n48990), .A3(n2647), .ZN(n52177) );
  NAND2_X2 U18316 ( .A1(n9860), .A2(n47843), .ZN(n2641) );
  BUF_X2 U18318 ( .I(n23745), .Z(n62128) );
  XOR2_X1 U18321 ( .A1(n62129), .A2(n22821), .Z(Plaintext[13]) );
  NAND4_X2 U18326 ( .A1(n19672), .A2(n63981), .A3(n19676), .A4(n63980), .ZN(
        n62129) );
  NOR2_X2 U18328 ( .A1(n2644), .A2(n2642), .ZN(n62130) );
  OR2_X1 U18336 ( .A1(n17135), .A2(n17137), .Z(n62131) );
  XOR2_X1 U18349 ( .A1(n62132), .A2(n41144), .Z(n11519) );
  XOR2_X1 U18350 ( .A1(n41142), .A2(n45052), .Z(n62132) );
  NAND2_X1 U18361 ( .A1(n40904), .A2(n40905), .ZN(n64761) );
  AOI21_X1 U18364 ( .A1(n6790), .A2(n25545), .B(n19594), .ZN(n53250) );
  INV_X1 U18365 ( .I(n33825), .ZN(n62464) );
  NAND3_X2 U18371 ( .A1(n4115), .A2(n62268), .A3(n35806), .ZN(n13406) );
  NAND3_X2 U18375 ( .A1(n61789), .A2(n63132), .A3(n34386), .ZN(n4115) );
  XOR2_X1 U18377 ( .A1(n20882), .A2(n10599), .Z(n21025) );
  NAND2_X2 U18379 ( .A1(n62133), .A2(n23427), .ZN(n43261) );
  NOR2_X2 U18380 ( .A1(n63728), .A2(n64570), .ZN(n62133) );
  NAND3_X1 U18387 ( .A1(n12163), .A2(n63140), .A3(n29924), .ZN(n4889) );
  NAND2_X2 U18388 ( .A1(n39153), .A2(n62135), .ZN(n63736) );
  AOI22_X2 U18391 ( .A1(n39143), .A2(n9444), .B1(n41177), .B2(n39144), .ZN(
        n62135) );
  BUF_X2 U18395 ( .I(n2036), .Z(n62136) );
  OAI21_X1 U18400 ( .A1(n64374), .A2(n28271), .B(n62128), .ZN(n27401) );
  AOI21_X1 U18402 ( .A1(n42717), .A2(n42726), .B(n2255), .ZN(n62137) );
  XOR2_X1 U18403 ( .A1(n50549), .A2(n51081), .Z(n51987) );
  NAND3_X2 U18408 ( .A1(n48816), .A2(n62201), .A3(n62811), .ZN(n50549) );
  XOR2_X1 U18413 ( .A1(n44422), .A2(n12178), .Z(n12179) );
  NAND3_X2 U18422 ( .A1(n22538), .A2(n64127), .A3(n63104), .ZN(n44422) );
  NOR3_X2 U18424 ( .A1(n16914), .A2(n62138), .A3(n15482), .ZN(n10751) );
  AOI21_X1 U18425 ( .A1(n37416), .A2(n3109), .B(n40203), .ZN(n62138) );
  NOR3_X2 U18427 ( .A1(n62854), .A2(n62140), .A3(n22402), .ZN(n35678) );
  XOR2_X1 U18431 ( .A1(n20512), .A2(n22350), .Z(n6994) );
  AND2_X1 U18435 ( .A1(n30254), .A2(n16631), .Z(n29057) );
  XOR2_X1 U18439 ( .A1(n63271), .A2(n62141), .Z(n6181) );
  XOR2_X1 U18441 ( .A1(n39630), .A2(n37876), .Z(n62141) );
  OR2_X2 U18448 ( .A1(n25078), .A2(n15740), .Z(n7321) );
  XOR2_X1 U18452 ( .A1(n14755), .A2(n38286), .Z(n39482) );
  XOR2_X1 U18453 ( .A1(n38573), .A2(n20470), .Z(n38286) );
  XOR2_X1 U18454 ( .A1(n19), .A2(n25973), .Z(n62507) );
  NOR2_X2 U18455 ( .A1(n42596), .A2(n42597), .ZN(n42612) );
  NOR2_X2 U18458 ( .A1(n24188), .A2(n8452), .ZN(n38026) );
  NAND2_X2 U18460 ( .A1(n62142), .A2(n24612), .ZN(n43069) );
  NOR2_X2 U18462 ( .A1(n24611), .A2(n65073), .ZN(n62142) );
  NAND2_X2 U18465 ( .A1(n53625), .A2(n53622), .ZN(n53614) );
  NAND2_X2 U18467 ( .A1(n6129), .A2(n22105), .ZN(n53622) );
  NOR2_X2 U18494 ( .A1(n62143), .A2(n48159), .ZN(n50257) );
  NAND3_X2 U18495 ( .A1(n48158), .A2(n48156), .A3(n23076), .ZN(n62143) );
  NAND2_X1 U18498 ( .A1(n15357), .A2(n16030), .ZN(n14311) );
  OAI22_X2 U18515 ( .A1(n62170), .A2(n24089), .B1(n34404), .B2(n62598), .ZN(
        n33809) );
  XOR2_X1 U18516 ( .A1(n10447), .A2(n62145), .Z(n12754) );
  XOR2_X1 U18524 ( .A1(n8620), .A2(n62146), .Z(n62145) );
  OR2_X1 U18526 ( .A1(n13438), .A2(n63321), .Z(n16783) );
  XOR2_X1 U18529 ( .A1(n1749), .A2(n37647), .Z(n5911) );
  XOR2_X1 U18541 ( .A1(n1752), .A2(n6026), .Z(n37647) );
  XOR2_X1 U18543 ( .A1(n11733), .A2(n62147), .Z(n58099) );
  NOR3_X1 U18546 ( .A1(n62148), .A2(n25964), .A3(n37065), .ZN(n8817) );
  NAND2_X2 U18552 ( .A1(n17556), .A2(n62149), .ZN(n57738) );
  NOR3_X2 U18555 ( .A1(n18662), .A2(n18665), .A3(n63590), .ZN(n62149) );
  NAND2_X2 U18560 ( .A1(n25167), .A2(n56389), .ZN(n56396) );
  NOR2_X2 U18563 ( .A1(n22794), .A2(n18335), .ZN(n56389) );
  XOR2_X1 U18566 ( .A1(n16892), .A2(n16535), .Z(n26067) );
  NAND3_X1 U18571 ( .A1(n35024), .A2(n23125), .A3(n11477), .ZN(n34023) );
  NAND2_X2 U18577 ( .A1(n1543), .A2(n34025), .ZN(n11477) );
  OAI22_X2 U18578 ( .A1(n57684), .A2(n26749), .B1(n26750), .B2(n62213), .ZN(
        n65076) );
  XOR2_X1 U18582 ( .A1(n25660), .A2(n19511), .Z(n9739) );
  XOR2_X1 U18584 ( .A1(n11595), .A2(n44747), .Z(n25660) );
  XOR2_X1 U18588 ( .A1(n22066), .A2(n32228), .Z(n31950) );
  NAND2_X1 U18591 ( .A1(n60906), .A2(n7302), .ZN(n62177) );
  XOR2_X1 U18598 ( .A1(n50766), .A2(n23991), .Z(n50767) );
  NAND2_X2 U18600 ( .A1(n61565), .A2(n58499), .ZN(n23991) );
  INV_X2 U18602 ( .I(n32999), .ZN(n8309) );
  NAND2_X2 U18603 ( .A1(n18088), .A2(n65256), .ZN(n32999) );
  AND2_X2 U18608 ( .A1(n59912), .A2(n36394), .Z(n36550) );
  NAND3_X2 U18613 ( .A1(n14392), .A2(n14390), .A3(n14391), .ZN(n58481) );
  NOR2_X2 U18614 ( .A1(n13235), .A2(n62150), .ZN(n13234) );
  NAND3_X2 U18622 ( .A1(n37595), .A2(n37594), .A3(n18358), .ZN(n62150) );
  NOR2_X2 U18626 ( .A1(n22972), .A2(n63258), .ZN(n39522) );
  INV_X1 U18634 ( .I(n1866), .ZN(n62152) );
  AND2_X1 U18646 ( .A1(n16517), .A2(n62152), .Z(n29898) );
  INV_X1 U18648 ( .I(n38051), .ZN(n62427) );
  NOR2_X2 U18651 ( .A1(n62154), .A2(n39951), .ZN(n11731) );
  NOR2_X1 U18655 ( .A1(n39953), .A2(n7259), .ZN(n62154) );
  NAND3_X2 U18656 ( .A1(n11509), .A2(n62156), .A3(n22119), .ZN(n22121) );
  XOR2_X1 U18669 ( .A1(n4546), .A2(n22890), .Z(n1198) );
  NAND2_X2 U18671 ( .A1(n42351), .A2(n42350), .ZN(n22890) );
  BUF_X2 U18684 ( .I(n40924), .Z(n62157) );
  XOR2_X1 U18685 ( .A1(n62159), .A2(n51589), .Z(n61537) );
  XOR2_X1 U18687 ( .A1(n51592), .A2(n51591), .Z(n62159) );
  OAI21_X2 U18695 ( .A1(n44864), .A2(n17366), .B(n62160), .ZN(n44865) );
  NOR2_X2 U18697 ( .A1(n44862), .A2(n44863), .ZN(n62160) );
  XOR2_X1 U18700 ( .A1(n62163), .A2(n65270), .Z(n63314) );
  XOR2_X1 U18702 ( .A1(n58467), .A2(n21508), .Z(n62163) );
  XOR2_X1 U18708 ( .A1(n14424), .A2(n14425), .Z(n18639) );
  NAND2_X2 U18710 ( .A1(n892), .A2(n2614), .ZN(n1343) );
  NAND3_X2 U18714 ( .A1(n62690), .A2(n11753), .A3(n62164), .ZN(n23619) );
  OAI21_X1 U18716 ( .A1(n37093), .A2(n37094), .B(n37092), .ZN(n62164) );
  NAND2_X2 U18718 ( .A1(n1252), .A2(n23184), .ZN(n43011) );
  NAND2_X1 U18721 ( .A1(n62463), .A2(n62464), .ZN(n63388) );
  NAND2_X2 U18727 ( .A1(n43016), .A2(n40903), .ZN(n41999) );
  NOR2_X2 U18731 ( .A1(n1252), .A2(n23425), .ZN(n43016) );
  NAND2_X1 U18732 ( .A1(n46079), .A2(n21980), .ZN(n62165) );
  NAND2_X2 U18733 ( .A1(n6197), .A2(n62184), .ZN(n63312) );
  NAND4_X1 U18736 ( .A1(n53063), .A2(n53062), .A3(n53061), .A4(n53060), .ZN(
        n62459) );
  XOR2_X1 U18738 ( .A1(n62166), .A2(n65280), .Z(n16814) );
  XOR2_X1 U18740 ( .A1(n50559), .A2(n50558), .Z(n62166) );
  XOR2_X1 U18746 ( .A1(n62167), .A2(n44607), .Z(n22053) );
  XOR2_X1 U18749 ( .A1(n21141), .A2(n57892), .Z(n62167) );
  XOR2_X1 U18752 ( .A1(n16747), .A2(n1124), .Z(n11993) );
  XOR2_X1 U18753 ( .A1(n4311), .A2(n52073), .Z(n50557) );
  NOR2_X2 U18763 ( .A1(n26065), .A2(n24215), .ZN(n4311) );
  AOI22_X2 U18784 ( .A1(n39520), .A2(n62169), .B1(n40557), .B2(n62168), .ZN(
        n39521) );
  INV_X1 U18785 ( .I(n35717), .ZN(n62170) );
  XOR2_X1 U18788 ( .A1(n62171), .A2(n53246), .Z(Plaintext[12]) );
  INV_X2 U18791 ( .I(n45504), .ZN(n46076) );
  NAND2_X2 U18792 ( .A1(n16686), .A2(n45498), .ZN(n45504) );
  XOR2_X1 U18799 ( .A1(n7608), .A2(n62172), .Z(n7607) );
  XOR2_X1 U18803 ( .A1(n19146), .A2(n17272), .Z(n62172) );
  OAI21_X2 U18806 ( .A1(n62173), .A2(n26120), .B(n61115), .ZN(n51030) );
  AND2_X1 U18807 ( .A1(n48334), .A2(n48739), .Z(n62174) );
  NAND2_X2 U18811 ( .A1(n7580), .A2(n21014), .ZN(n63589) );
  NAND2_X2 U18819 ( .A1(n7715), .A2(n63885), .ZN(n7580) );
  XOR2_X1 U18826 ( .A1(n46395), .A2(n64552), .Z(n61252) );
  INV_X2 U18830 ( .I(n20255), .ZN(n20250) );
  NAND2_X2 U18831 ( .A1(n20258), .A2(n62176), .ZN(n20255) );
  AND2_X1 U18838 ( .A1(n20257), .A2(n20256), .Z(n62176) );
  BUF_X2 U18844 ( .I(n49908), .Z(n64990) );
  OR2_X1 U18847 ( .A1(n54106), .A2(n53549), .Z(n10842) );
  INV_X2 U18848 ( .I(n12697), .ZN(n11442) );
  NAND2_X2 U18851 ( .A1(n62252), .A2(n63178), .ZN(n12697) );
  XOR2_X1 U18855 ( .A1(n25643), .A2(n38910), .Z(n38769) );
  XOR2_X1 U18856 ( .A1(n38469), .A2(n39310), .Z(n38910) );
  XOR2_X1 U18857 ( .A1(n21130), .A2(n37670), .Z(n5266) );
  AOI21_X2 U18878 ( .A1(n13301), .A2(n13302), .B(n13300), .ZN(n37670) );
  NAND2_X1 U18884 ( .A1(n65167), .A2(n61881), .ZN(n34599) );
  INV_X2 U18885 ( .I(n62179), .ZN(n8576) );
  XNOR2_X1 U18895 ( .A1(n972), .A2(n2219), .ZN(n62179) );
  AOI21_X2 U18908 ( .A1(n35885), .A2(n35567), .B(n10596), .ZN(n35892) );
  NAND3_X1 U18909 ( .A1(n58808), .A2(n1967), .A3(n22343), .ZN(n7632) );
  NAND2_X2 U18918 ( .A1(n2352), .A2(n7584), .ZN(n21014) );
  NAND2_X2 U18928 ( .A1(n9170), .A2(n58140), .ZN(n60825) );
  NAND3_X2 U18932 ( .A1(n41809), .A2(n1401), .A3(n753), .ZN(n62184) );
  NAND2_X2 U18935 ( .A1(n1221), .A2(n33797), .ZN(n6829) );
  NAND3_X2 U18939 ( .A1(n34442), .A2(n33798), .A3(n35656), .ZN(n62844) );
  NAND3_X2 U18949 ( .A1(n59690), .A2(n3680), .A3(n3677), .ZN(n23054) );
  NAND3_X2 U18955 ( .A1(n62772), .A2(n4160), .A3(n4161), .ZN(n4166) );
  NOR2_X2 U18957 ( .A1(n1221), .A2(n33797), .ZN(n59005) );
  NAND3_X1 U18959 ( .A1(n5049), .A2(n55312), .A3(n15100), .ZN(n25717) );
  NOR2_X2 U18962 ( .A1(n61096), .A2(n31420), .ZN(n37035) );
  NOR3_X2 U18966 ( .A1(n761), .A2(n27633), .A3(n27632), .ZN(n27638) );
  AOI22_X2 U18969 ( .A1(n47142), .A2(n46746), .B1(n62634), .B2(n45435), .ZN(
        n45440) );
  AOI21_X2 U18977 ( .A1(n47372), .A2(n21451), .B(n62634), .ZN(n46746) );
  NAND2_X2 U18978 ( .A1(n26583), .A2(n4491), .ZN(n6149) );
  NOR2_X2 U18984 ( .A1(n23938), .A2(n26582), .ZN(n26583) );
  NAND2_X1 U18986 ( .A1(n35646), .A2(n62188), .ZN(n62187) );
  NAND3_X2 U18988 ( .A1(n41351), .A2(n4522), .A3(n41352), .ZN(n46620) );
  NAND2_X1 U18989 ( .A1(n62189), .A2(n62187), .ZN(n16728) );
  INV_X1 U18990 ( .I(n6829), .ZN(n62188) );
  NAND2_X1 U18992 ( .A1(n34446), .A2(n6829), .ZN(n62189) );
  NAND2_X2 U18993 ( .A1(n35655), .A2(n33583), .ZN(n34446) );
  NAND3_X1 U18994 ( .A1(n37355), .A2(n18123), .A3(n18779), .ZN(n63120) );
  XOR2_X1 U18995 ( .A1(n50780), .A2(n50716), .Z(n51119) );
  XOR2_X1 U18996 ( .A1(n19806), .A2(n14108), .Z(n50780) );
  XOR2_X1 U18997 ( .A1(n44806), .A2(n2960), .Z(n17586) );
  XOR2_X1 U19000 ( .A1(n24733), .A2(n63763), .Z(n44806) );
  NAND3_X2 U19005 ( .A1(n23099), .A2(n21304), .A3(n16950), .ZN(n11087) );
  BUF_X2 U19007 ( .I(n21699), .Z(n62190) );
  AOI21_X2 U19008 ( .A1(n43523), .A2(n62418), .B(n62193), .ZN(n62382) );
  OAI21_X1 U19010 ( .A1(n43518), .A2(n25210), .B(n43521), .ZN(n62194) );
  AND2_X2 U19015 ( .A1(n13418), .A2(n826), .Z(n11108) );
  XOR2_X1 U19022 ( .A1(n61037), .A2(n8796), .Z(n34342) );
  XOR2_X1 U19024 ( .A1(n19551), .A2(n21823), .Z(n8796) );
  XOR2_X1 U19025 ( .A1(n62646), .A2(n2367), .Z(n45366) );
  NAND2_X2 U19031 ( .A1(n43586), .A2(n9209), .ZN(n44442) );
  NOR2_X2 U19044 ( .A1(n9214), .A2(n41795), .ZN(n43586) );
  INV_X2 U19046 ( .I(n6133), .ZN(n37812) );
  NAND2_X2 U19050 ( .A1(n6132), .A2(n6131), .ZN(n6133) );
  NOR2_X2 U19053 ( .A1(n17761), .A2(n35182), .ZN(n36261) );
  XOR2_X1 U19074 ( .A1(n38952), .A2(n19418), .Z(n38643) );
  XOR2_X1 U19080 ( .A1(n63412), .A2(n48946), .Z(n8716) );
  NAND3_X2 U19088 ( .A1(n8713), .A2(n8715), .A3(n8714), .ZN(n48946) );
  XOR2_X1 U19090 ( .A1(n17252), .A2(n62195), .Z(n17251) );
  XOR2_X1 U19093 ( .A1(n18491), .A2(n23032), .Z(n62195) );
  NOR3_X2 U19099 ( .A1(n12924), .A2(n15550), .A3(n15549), .ZN(n18863) );
  NAND4_X1 U19101 ( .A1(n53654), .A2(n10021), .A3(n22707), .A4(n53653), .ZN(
        n64289) );
  NOR2_X1 U19113 ( .A1(n12042), .A2(n37538), .ZN(n64752) );
  NAND3_X2 U19117 ( .A1(n29823), .A2(n30322), .A3(n29820), .ZN(n3706) );
  NOR2_X2 U19118 ( .A1(n29988), .A2(n1208), .ZN(n29823) );
  AOI21_X2 U19122 ( .A1(n16182), .A2(n61888), .B(n62196), .ZN(n16608) );
  NOR2_X1 U19123 ( .A1(n16610), .A2(n29267), .ZN(n62196) );
  XOR2_X1 U19126 ( .A1(n1818), .A2(n64026), .Z(n13964) );
  OR2_X1 U19129 ( .A1(n19885), .A2(n13731), .Z(n29264) );
  NOR2_X2 U19143 ( .A1(n22428), .A2(n35629), .ZN(n33548) );
  NAND2_X2 U19145 ( .A1(n59912), .A2(n36538), .ZN(n24078) );
  NAND2_X2 U19146 ( .A1(n32998), .A2(n32997), .ZN(n36538) );
  AOI22_X2 U19157 ( .A1(n36058), .A2(n36059), .B1(n36061), .B2(n36060), .ZN(
        n62197) );
  NAND3_X2 U19163 ( .A1(n41185), .A2(n40485), .A3(n40486), .ZN(n40499) );
  NAND2_X2 U19174 ( .A1(n7402), .A2(n41177), .ZN(n41185) );
  XOR2_X1 U19175 ( .A1(n51910), .A2(n1462), .Z(n51317) );
  XOR2_X1 U19187 ( .A1(n25378), .A2(n21100), .Z(n51910) );
  OR2_X1 U19203 ( .A1(n8026), .A2(n9711), .Z(n64602) );
  INV_X2 U19205 ( .I(n46947), .ZN(n63663) );
  NAND2_X2 U19208 ( .A1(n6411), .A2(n18464), .ZN(n46947) );
  OAI21_X2 U19217 ( .A1(n48814), .A2(n48813), .B(n48812), .ZN(n62201) );
  XOR2_X1 U19218 ( .A1(n60382), .A2(n12662), .Z(n24108) );
  NOR3_X2 U19224 ( .A1(n62202), .A2(n26440), .A3(n30784), .ZN(n61334) );
  BUF_X4 U19225 ( .I(n33276), .Z(n1221) );
  NOR2_X2 U19232 ( .A1(n21282), .A2(n63695), .ZN(n21667) );
  NAND3_X2 U19243 ( .A1(n40883), .A2(n62203), .A3(n18228), .ZN(n18297) );
  XOR2_X1 U19244 ( .A1(n3333), .A2(n52172), .Z(n51140) );
  NAND2_X2 U19245 ( .A1(n16816), .A2(n16916), .ZN(n3333) );
  NOR2_X2 U19254 ( .A1(n62205), .A2(n62204), .ZN(n40799) );
  AND2_X1 U19273 ( .A1(n21400), .A2(n40839), .Z(n20700) );
  NOR2_X2 U19278 ( .A1(n37329), .A2(n35876), .ZN(n37182) );
  INV_X2 U19279 ( .I(n9830), .ZN(n37329) );
  NAND2_X2 U19280 ( .A1(n57220), .A2(n6124), .ZN(n9830) );
  NAND2_X2 U19308 ( .A1(n31841), .A2(n62206), .ZN(n34295) );
  NOR3_X2 U19315 ( .A1(n897), .A2(n17498), .A3(n35803), .ZN(n62206) );
  XOR2_X1 U19323 ( .A1(n45426), .A2(n44177), .Z(n43826) );
  XOR2_X1 U19324 ( .A1(n11857), .A2(n17982), .Z(n44177) );
  XOR2_X1 U19332 ( .A1(n6255), .A2(n21088), .Z(n64891) );
  XOR2_X1 U19333 ( .A1(n21100), .A2(n59555), .Z(n21088) );
  NAND2_X2 U19342 ( .A1(n48612), .A2(n8639), .ZN(n62308) );
  XOR2_X1 U19346 ( .A1(n20230), .A2(n55889), .Z(n62207) );
  XOR2_X1 U19356 ( .A1(n62209), .A2(n62208), .Z(n61041) );
  XOR2_X1 U19357 ( .A1(n22577), .A2(n50326), .Z(n62209) );
  BUF_X4 U19367 ( .I(n56817), .Z(n65064) );
  XOR2_X1 U19369 ( .A1(n62210), .A2(n5890), .Z(Plaintext[169]) );
  NOR4_X2 U19372 ( .A1(n5894), .A2(n5892), .A3(n5893), .A4(n5896), .ZN(n62210)
         );
  XOR2_X1 U19373 ( .A1(n32744), .A2(n60466), .Z(n62799) );
  NOR2_X2 U19374 ( .A1(n63218), .A2(n63217), .ZN(n60466) );
  AND2_X1 U19376 ( .A1(n53865), .A2(n62211), .Z(n60871) );
  XOR2_X1 U19387 ( .A1(n62212), .A2(n58145), .Z(n7559) );
  XOR2_X1 U19388 ( .A1(n59720), .A2(n19145), .Z(n62212) );
  NAND3_X1 U19391 ( .A1(n28270), .A2(n62663), .A3(n23876), .ZN(n27063) );
  NAND2_X2 U19393 ( .A1(n23745), .A2(n27966), .ZN(n62663) );
  OAI21_X1 U19395 ( .A1(n16014), .A2(n28697), .B(n23395), .ZN(n62556) );
  NOR2_X1 U19397 ( .A1(n5936), .A2(n36946), .ZN(n36948) );
  NAND2_X2 U19405 ( .A1(n16337), .A2(n35431), .ZN(n36946) );
  BUF_X2 U19406 ( .I(n29158), .Z(n62213) );
  NOR2_X2 U19410 ( .A1(n28020), .A2(n62214), .ZN(n28080) );
  NAND3_X2 U19411 ( .A1(n28016), .A2(n28017), .A3(n28015), .ZN(n62214) );
  NAND2_X2 U19415 ( .A1(n12003), .A2(n26000), .ZN(n9164) );
  XOR2_X1 U19420 ( .A1(n7559), .A2(n59575), .Z(n20348) );
  XNOR2_X1 U19428 ( .A1(n31480), .A2(n31481), .ZN(n62919) );
  XOR2_X1 U19432 ( .A1(n33132), .A2(n60392), .Z(n31481) );
  XOR2_X1 U19433 ( .A1(n19060), .A2(n13705), .Z(n64194) );
  AOI21_X2 U19439 ( .A1(n54471), .A2(n54599), .B(n64129), .ZN(n64665) );
  OAI22_X1 U19442 ( .A1(n11006), .A2(n6984), .B1(n11007), .B2(n36825), .ZN(
        n64015) );
  NAND2_X1 U19444 ( .A1(n18714), .A2(n62930), .ZN(n3362) );
  NAND2_X2 U19447 ( .A1(n22236), .A2(n17240), .ZN(n62216) );
  XOR2_X1 U19448 ( .A1(n7058), .A2(n30550), .Z(n31911) );
  NAND3_X2 U19455 ( .A1(n63462), .A2(n6818), .A3(n6817), .ZN(n7058) );
  NAND2_X1 U19456 ( .A1(n30187), .A2(n22799), .ZN(n62586) );
  INV_X2 U19458 ( .I(n62217), .ZN(n53537) );
  AND2_X1 U19459 ( .A1(n10870), .A2(n10868), .Z(n62217) );
  INV_X2 U19464 ( .I(n41163), .ZN(n25424) );
  NAND2_X1 U19465 ( .A1(n20925), .A2(n41163), .ZN(n38418) );
  NOR2_X2 U19466 ( .A1(n14732), .A2(n41165), .ZN(n41163) );
  XOR2_X1 U19468 ( .A1(n4074), .A2(n4073), .Z(n7510) );
  NOR3_X2 U19469 ( .A1(n20254), .A2(n20261), .A3(n20262), .ZN(n18875) );
  NOR3_X2 U19473 ( .A1(n62221), .A2(n62218), .A3(n12327), .ZN(n58324) );
  NOR2_X1 U19474 ( .A1(n62220), .A2(n62219), .ZN(n62218) );
  NAND4_X2 U19485 ( .A1(n5316), .A2(n5315), .A3(n41598), .A4(n41599), .ZN(
        n65226) );
  NOR2_X2 U19489 ( .A1(n9205), .A2(n4880), .ZN(n32784) );
  XOR2_X1 U19497 ( .A1(n14999), .A2(n62615), .Z(n24390) );
  XOR2_X1 U19514 ( .A1(n62222), .A2(n45377), .Z(n46581) );
  XOR2_X1 U19564 ( .A1(n8381), .A2(n44084), .Z(n62222) );
  NAND3_X2 U19583 ( .A1(n1922), .A2(n1924), .A3(n1921), .ZN(n33239) );
  NAND3_X2 U19592 ( .A1(n40847), .A2(n19045), .A3(n40846), .ZN(n41642) );
  NOR3_X2 U19595 ( .A1(n60983), .A2(n19107), .A3(n4436), .ZN(n62619) );
  NAND4_X1 U19619 ( .A1(n32907), .A2(n62223), .A3(n36921), .A4(n32908), .ZN(
        n32912) );
  NAND2_X2 U19633 ( .A1(n62224), .A2(n49893), .ZN(n58770) );
  NAND2_X1 U19640 ( .A1(n13147), .A2(n49895), .ZN(n62224) );
  NOR2_X1 U19649 ( .A1(n60982), .A2(n43214), .ZN(n13522) );
  XOR2_X1 U19668 ( .A1(n2998), .A2(n9242), .Z(n6636) );
  NAND2_X2 U19670 ( .A1(n3005), .A2(n3004), .ZN(n9242) );
  NAND2_X2 U19702 ( .A1(n25535), .A2(n25781), .ZN(n52568) );
  NOR2_X2 U19712 ( .A1(n52674), .A2(n62225), .ZN(n57083) );
  XOR2_X1 U19720 ( .A1(n62226), .A2(n22166), .Z(n59559) );
  XOR2_X1 U19726 ( .A1(n62383), .A2(n38903), .Z(n62226) );
  INV_X2 U19766 ( .I(n54944), .ZN(n54616) );
  NAND2_X2 U19768 ( .A1(n54778), .A2(n54605), .ZN(n54944) );
  OR2_X1 U19780 ( .A1(n61094), .A2(n41220), .Z(n40404) );
  NAND3_X2 U19783 ( .A1(n13350), .A2(n22546), .A3(n57213), .ZN(n62541) );
  XOR2_X1 U19794 ( .A1(n18888), .A2(n63716), .Z(n47491) );
  NAND2_X2 U19795 ( .A1(n62227), .A2(n17484), .ZN(n5587) );
  NOR3_X2 U19798 ( .A1(n6187), .A2(n224), .A3(n223), .ZN(n62227) );
  XOR2_X1 U19799 ( .A1(Ciphertext[80]), .A2(Key[165]), .Z(n6888) );
  XOR2_X1 U19802 ( .A1(n51918), .A2(n10584), .Z(n51590) );
  NAND4_X2 U19806 ( .A1(n45790), .A2(n20184), .A3(n63139), .A4(n20185), .ZN(
        n48074) );
  XOR2_X1 U19810 ( .A1(n1835), .A2(n61152), .Z(n12374) );
  NAND2_X2 U19824 ( .A1(n5294), .A2(n30533), .ZN(n61152) );
  NOR2_X2 U19825 ( .A1(n62446), .A2(n62445), .ZN(n58128) );
  AOI22_X2 U19856 ( .A1(n13002), .A2(n41379), .B1(n41377), .B2(n41378), .ZN(
        n62228) );
  NOR2_X2 U19925 ( .A1(n61739), .A2(n9663), .ZN(n43325) );
  NOR2_X1 U19931 ( .A1(n15171), .A2(n24609), .ZN(n14743) );
  NAND2_X2 U19933 ( .A1(n17525), .A2(n17524), .ZN(n31327) );
  NAND3_X2 U19942 ( .A1(n18363), .A2(n43692), .A3(n43691), .ZN(n62945) );
  NAND3_X1 U19944 ( .A1(n27924), .A2(n30523), .A3(n8891), .ZN(n17115) );
  XOR2_X1 U19948 ( .A1(n38708), .A2(n24536), .Z(n37801) );
  NAND2_X2 U19950 ( .A1(n57569), .A2(n12809), .ZN(n24536) );
  NAND2_X1 U19952 ( .A1(n60319), .A2(n42824), .ZN(n21173) );
  NAND3_X2 U19954 ( .A1(n25355), .A2(n35600), .A3(n62229), .ZN(n38702) );
  NAND2_X1 U19956 ( .A1(n35594), .A2(n4611), .ZN(n62229) );
  NOR2_X2 U19959 ( .A1(n26391), .A2(n26826), .ZN(n27837) );
  BUF_X2 U19962 ( .I(n24099), .Z(n62230) );
  XOR2_X1 U19968 ( .A1(n39709), .A2(n15631), .Z(n6832) );
  NAND2_X2 U19971 ( .A1(n58942), .A2(n6836), .ZN(n15631) );
  BUF_X2 U19976 ( .I(n29773), .Z(n62231) );
  XOR2_X1 U19981 ( .A1(n3479), .A2(n62399), .Z(n39660) );
  INV_X2 U19982 ( .I(n36587), .ZN(n36596) );
  NAND2_X2 U19987 ( .A1(n22632), .A2(n9783), .ZN(n36587) );
  XOR2_X1 U19993 ( .A1(n8901), .A2(n61490), .Z(n14720) );
  AND2_X2 U20001 ( .A1(n39011), .A2(n15590), .Z(n41405) );
  NAND2_X1 U20005 ( .A1(n15343), .A2(n41411), .ZN(n64253) );
  XOR2_X1 U20006 ( .A1(n50195), .A2(n6298), .Z(n12462) );
  NAND3_X2 U20007 ( .A1(n12216), .A2(n58691), .A3(n12215), .ZN(n50195) );
  XOR2_X1 U20011 ( .A1(n31851), .A2(n58099), .Z(n16833) );
  NOR3_X2 U20012 ( .A1(n40989), .A2(n62232), .A3(n59183), .ZN(n40999) );
  OAI21_X2 U20019 ( .A1(n21380), .A2(n57279), .B(n16133), .ZN(n2883) );
  NOR2_X2 U20027 ( .A1(n13506), .A2(n47489), .ZN(n46103) );
  XOR2_X1 U20028 ( .A1(Ciphertext[111]), .A2(Key[94]), .Z(n26826) );
  NAND2_X1 U20034 ( .A1(n32879), .A2(n32880), .ZN(n62445) );
  XOR2_X1 U20042 ( .A1(n9917), .A2(n38457), .Z(n13906) );
  XOR2_X1 U20044 ( .A1(n25995), .A2(n38870), .Z(n38457) );
  XOR2_X1 U20046 ( .A1(n60897), .A2(n5729), .Z(n13410) );
  NOR2_X2 U20051 ( .A1(n40033), .A2(n62233), .ZN(n43460) );
  BUF_X2 U20059 ( .I(n29156), .Z(n62234) );
  AOI22_X2 U20062 ( .A1(n5719), .A2(n5720), .B1(n42964), .B2(n42068), .ZN(
        n5718) );
  OAI21_X2 U20063 ( .A1(n8377), .A2(n61624), .B(n62235), .ZN(n24330) );
  OAI21_X2 U20072 ( .A1(n11678), .A2(n11108), .B(n61624), .ZN(n62235) );
  NAND2_X2 U20073 ( .A1(n60826), .A2(n61477), .ZN(n11316) );
  NOR2_X2 U20080 ( .A1(n3403), .A2(n1744), .ZN(n60826) );
  XOR2_X1 U20082 ( .A1(n45876), .A2(n45376), .Z(n15075) );
  XOR2_X1 U20083 ( .A1(n62236), .A2(n52232), .Z(Plaintext[11]) );
  NAND3_X1 U20086 ( .A1(n3544), .A2(n3540), .A3(n53126), .ZN(n62236) );
  NAND3_X2 U20095 ( .A1(n62238), .A2(n13397), .A3(n13396), .ZN(n18502) );
  XOR2_X1 U20101 ( .A1(n24213), .A2(n57809), .Z(n22068) );
  OR3_X1 U20108 ( .A1(n40217), .A2(n58264), .A3(n40146), .Z(n38041) );
  NOR3_X2 U20109 ( .A1(n3806), .A2(n62240), .A3(n62239), .ZN(n60725) );
  NOR2_X1 U20112 ( .A1(n64240), .A2(n64239), .ZN(n62240) );
  NAND2_X1 U20115 ( .A1(n62461), .A2(n8986), .ZN(n59425) );
  NAND2_X2 U20125 ( .A1(n18027), .A2(n18029), .ZN(n8986) );
  AOI22_X1 U20128 ( .A1(n28916), .A2(n28917), .B1(n28915), .B2(n30623), .ZN(
        n22262) );
  NOR2_X2 U20129 ( .A1(n30343), .A2(n29083), .ZN(n30623) );
  AOI21_X2 U20140 ( .A1(n53178), .A2(n62243), .B(n62242), .ZN(n50484) );
  OR2_X1 U20144 ( .A1(n50478), .A2(n53540), .Z(n62243) );
  INV_X2 U20145 ( .I(n3979), .ZN(n49770) );
  NAND2_X2 U20146 ( .A1(n57735), .A2(n4271), .ZN(n3979) );
  INV_X1 U20147 ( .I(n21724), .ZN(n1331) );
  NAND3_X2 U20148 ( .A1(n3657), .A2(n41718), .A3(n65100), .ZN(n21724) );
  INV_X1 U20149 ( .I(n32829), .ZN(n5731) );
  NAND2_X1 U20151 ( .A1(n7007), .A2(n32829), .ZN(n7016) );
  XOR2_X1 U20152 ( .A1(n58968), .A2(n4592), .Z(n32829) );
  INV_X2 U20155 ( .I(n11570), .ZN(n38367) );
  NAND2_X2 U20156 ( .A1(n4743), .A2(n11983), .ZN(n11570) );
  BUF_X2 U20157 ( .I(n1379), .Z(n62244) );
  XOR2_X1 U20158 ( .A1(n8342), .A2(n5094), .Z(n46577) );
  XOR2_X1 U20159 ( .A1(n46674), .A2(n5093), .Z(n8342) );
  NAND3_X1 U20160 ( .A1(n48154), .A2(n48155), .A3(n46798), .ZN(n46639) );
  INV_X2 U20161 ( .I(n36800), .ZN(n62246) );
  NOR2_X2 U20169 ( .A1(n24782), .A2(n11475), .ZN(n62247) );
  BUF_X2 U20176 ( .I(n39935), .Z(n43839) );
  XOR2_X1 U20182 ( .A1(n38512), .A2(n38123), .Z(n38992) );
  BUF_X2 U20185 ( .I(n23222), .Z(n12716) );
  NAND3_X2 U20186 ( .A1(n28465), .A2(n28463), .A3(n28464), .ZN(n28546) );
  XOR2_X1 U20189 ( .A1(n4876), .A2(n6416), .Z(n6415) );
  BUF_X2 U20197 ( .I(n18252), .Z(n62248) );
  NAND2_X2 U20203 ( .A1(n63794), .A2(n64116), .ZN(n21830) );
  NAND2_X2 U20205 ( .A1(n64494), .A2(n11760), .ZN(n11771) );
  NAND4_X1 U20206 ( .A1(n56114), .A2(n56113), .A3(n56112), .A4(n56111), .ZN(
        n56122) );
  INV_X4 U20207 ( .I(n62249), .ZN(n10717) );
  AND2_X2 U20208 ( .A1(n7030), .A2(n62429), .Z(n62249) );
  AOI21_X2 U20213 ( .A1(n28387), .A2(n27111), .B(n62250), .ZN(n27112) );
  OAI22_X2 U20215 ( .A1(n28380), .A2(n59279), .B1(n27109), .B2(n469), .ZN(
        n62250) );
  CLKBUF_X2 U20218 ( .I(n57146), .Z(n23302) );
  XOR2_X1 U20227 ( .A1(n62251), .A2(n55624), .Z(Plaintext[123]) );
  NAND4_X2 U20230 ( .A1(n55623), .A2(n55622), .A3(n55620), .A4(n55621), .ZN(
        n62251) );
  XOR2_X1 U20231 ( .A1(n52636), .A2(n12094), .Z(n12093) );
  INV_X1 U20233 ( .I(n18870), .ZN(n52636) );
  XOR2_X1 U20234 ( .A1(n51810), .A2(n10292), .Z(n18870) );
  OR2_X1 U20235 ( .A1(n23054), .A2(n18715), .Z(n62252) );
  NAND3_X1 U20236 ( .A1(n53723), .A2(n53721), .A3(n62253), .ZN(n53747) );
  NAND3_X1 U20240 ( .A1(n53719), .A2(n53720), .A3(n17286), .ZN(n62253) );
  AOI21_X1 U20244 ( .A1(n29737), .A2(n19087), .B(n4188), .ZN(n62254) );
  NOR3_X2 U20247 ( .A1(n8212), .A2(n47115), .A3(n23099), .ZN(n1098) );
  NOR2_X2 U20248 ( .A1(n62256), .A2(n14642), .ZN(n3684) );
  INV_X2 U20259 ( .I(n63368), .ZN(n62256) );
  XOR2_X1 U20261 ( .A1(n4650), .A2(n62257), .Z(n20535) );
  XOR2_X1 U20262 ( .A1(n32516), .A2(n33896), .Z(n62257) );
  XOR2_X1 U20263 ( .A1(n39261), .A2(n25624), .Z(n39348) );
  AND3_X1 U20264 ( .A1(n8348), .A2(n54872), .A3(n54873), .Z(n6511) );
  XOR2_X1 U20273 ( .A1(n62258), .A2(n51996), .Z(n59109) );
  XOR2_X1 U20279 ( .A1(n58787), .A2(n13755), .Z(n62258) );
  XOR2_X1 U20282 ( .A1(n52546), .A2(n52545), .Z(n52547) );
  NOR3_X2 U20288 ( .A1(n62259), .A2(n62365), .A3(n43849), .ZN(n62419) );
  NOR2_X1 U20289 ( .A1(n43841), .A2(n43842), .ZN(n62259) );
  NAND2_X1 U20290 ( .A1(n47685), .A2(n64704), .ZN(n59848) );
  BUF_X4 U20293 ( .I(n23839), .Z(n60360) );
  NOR3_X1 U20294 ( .A1(n62260), .A2(n21442), .A3(n21433), .ZN(n59300) );
  NAND2_X1 U20296 ( .A1(n21436), .A2(n21439), .ZN(n62260) );
  NAND2_X2 U20297 ( .A1(n61733), .A2(n23317), .ZN(n30286) );
  NAND2_X2 U20298 ( .A1(n8671), .A2(n8670), .ZN(n58606) );
  BUF_X2 U20301 ( .I(n1237), .Z(n62261) );
  AND2_X1 U20302 ( .A1(n33689), .A2(n63042), .Z(n33095) );
  XOR2_X1 U20306 ( .A1(n24342), .A2(n24343), .Z(n20270) );
  NAND2_X2 U20314 ( .A1(n63269), .A2(n4003), .ZN(n24342) );
  XOR2_X1 U20316 ( .A1(n7860), .A2(n24537), .Z(n8226) );
  XOR2_X1 U20325 ( .A1(n63684), .A2(n63685), .Z(n12062) );
  INV_X2 U20331 ( .I(n35212), .ZN(n62322) );
  NAND2_X2 U20333 ( .A1(n18879), .A2(n13583), .ZN(n35212) );
  NAND2_X2 U20338 ( .A1(n62262), .A2(n2609), .ZN(n11153) );
  NOR3_X2 U20343 ( .A1(n60348), .A2(n1071), .A3(n4352), .ZN(n62262) );
  INV_X2 U20349 ( .I(n64850), .ZN(n62263) );
  BUF_X2 U20353 ( .I(n1393), .Z(n62264) );
  NOR2_X2 U20354 ( .A1(n9122), .A2(n62265), .ZN(n13548) );
  OR2_X2 U20355 ( .A1(n21205), .A2(n17016), .Z(n2262) );
  NOR3_X2 U20357 ( .A1(n47195), .A2(n7672), .A3(n63994), .ZN(n21205) );
  NAND3_X2 U20358 ( .A1(n34298), .A2(n58150), .A3(n34300), .ZN(n62268) );
  NOR3_X2 U20360 ( .A1(n372), .A2(n1690), .A3(n57446), .ZN(n8756) );
  NOR2_X2 U20363 ( .A1(n57782), .A2(n8756), .ZN(n15478) );
  NAND3_X2 U20369 ( .A1(n47527), .A2(n47526), .A3(n64118), .ZN(n19933) );
  NOR2_X2 U20372 ( .A1(n49014), .A2(n48322), .ZN(n48454) );
  XOR2_X1 U20373 ( .A1(n5334), .A2(n8064), .Z(n5333) );
  NAND2_X2 U20374 ( .A1(n8319), .A2(n8318), .ZN(n8598) );
  XOR2_X1 U20376 ( .A1(n63559), .A2(n2391), .Z(n20707) );
  XOR2_X1 U20377 ( .A1(n6885), .A2(n60087), .Z(n2391) );
  AND2_X2 U20378 ( .A1(n64367), .A2(n11460), .Z(n57925) );
  BUF_X4 U20379 ( .I(n48404), .Z(n51863) );
  NAND2_X2 U20381 ( .A1(n4275), .A2(n1705), .ZN(n43391) );
  INV_X2 U20385 ( .I(n18006), .ZN(n62270) );
  OR2_X2 U20387 ( .A1(n37363), .A2(n9783), .Z(n34377) );
  AOI21_X2 U20388 ( .A1(n1655), .A2(n2826), .B(n61922), .ZN(n64171) );
  XOR2_X1 U20389 ( .A1(n38527), .A2(n3015), .Z(n62394) );
  XOR2_X1 U20393 ( .A1(n19311), .A2(n62273), .Z(n38527) );
  INV_X2 U20395 ( .I(n16346), .ZN(n62273) );
  NAND3_X1 U20399 ( .A1(n49514), .A2(n49515), .A3(n49513), .ZN(n62274) );
  NAND3_X1 U20400 ( .A1(n27142), .A2(n27141), .A3(n28049), .ZN(n27143) );
  INV_X2 U20401 ( .I(n62275), .ZN(n48213) );
  NOR2_X2 U20404 ( .A1(n16798), .A2(n9243), .ZN(n62275) );
  NOR2_X1 U20407 ( .A1(n62279), .A2(n20642), .ZN(n64430) );
  XOR2_X1 U20409 ( .A1(n58437), .A2(n62276), .Z(n58075) );
  XOR2_X1 U20410 ( .A1(n16558), .A2(n3713), .Z(n62276) );
  OAI21_X1 U20416 ( .A1(n34936), .A2(n35607), .B(n34935), .ZN(n62679) );
  NOR2_X1 U20418 ( .A1(n59149), .A2(n62277), .ZN(n41574) );
  NAND2_X1 U20419 ( .A1(n64660), .A2(n41570), .ZN(n62277) );
  NOR2_X2 U20420 ( .A1(n19212), .A2(n24844), .ZN(n62353) );
  XOR2_X1 U20421 ( .A1(n62278), .A2(n45375), .Z(n7635) );
  XOR2_X1 U20422 ( .A1(n58838), .A2(n16242), .Z(n62278) );
  NAND2_X1 U20423 ( .A1(n49052), .A2(n49051), .ZN(n62279) );
  AOI21_X2 U20426 ( .A1(n20425), .A2(n45723), .B(n63500), .ZN(n63499) );
  OAI21_X1 U20427 ( .A1(n20750), .A2(n55730), .B(n20749), .ZN(n62280) );
  NAND3_X2 U20435 ( .A1(n61962), .A2(n12387), .A3(n62281), .ZN(n39737) );
  XOR2_X1 U20437 ( .A1(n3232), .A2(n6253), .Z(n44905) );
  XOR2_X1 U20438 ( .A1(n13964), .A2(n15801), .Z(n16857) );
  AND2_X2 U20439 ( .A1(n16857), .A2(n4565), .Z(n33560) );
  AOI21_X1 U20441 ( .A1(n62282), .A2(n41655), .B(n57987), .ZN(n13603) );
  NOR2_X1 U20442 ( .A1(n43573), .A2(n42340), .ZN(n62282) );
  NAND2_X2 U20445 ( .A1(n50370), .A2(n62283), .ZN(n25970) );
  NOR3_X2 U20447 ( .A1(n3464), .A2(n50365), .A3(n50366), .ZN(n62283) );
  INV_X2 U20449 ( .I(n27962), .ZN(n28012) );
  NAND2_X2 U20450 ( .A1(n21946), .A2(n21265), .ZN(n27962) );
  NAND2_X1 U20453 ( .A1(n17250), .A2(n17249), .ZN(n62284) );
  BUF_X2 U20456 ( .I(n23140), .Z(n62285) );
  NOR2_X2 U20459 ( .A1(n64175), .A2(n37539), .ZN(n41795) );
  NOR2_X2 U20460 ( .A1(n61828), .A2(n62286), .ZN(n7059) );
  NAND2_X2 U20462 ( .A1(n52127), .A2(n19309), .ZN(n62286) );
  NOR2_X1 U20464 ( .A1(n8642), .A2(n8770), .ZN(n62766) );
  NAND2_X2 U20466 ( .A1(n53428), .A2(n50462), .ZN(n53427) );
  NAND4_X2 U20467 ( .A1(n8254), .A2(n57638), .A3(n10081), .A4(n8257), .ZN(
        n64204) );
  NAND2_X2 U20471 ( .A1(n41887), .A2(n6855), .ZN(n40840) );
  XOR2_X1 U20472 ( .A1(n46690), .A2(n44851), .Z(n16909) );
  NAND2_X2 U20474 ( .A1(n16339), .A2(n2853), .ZN(n46690) );
  XOR2_X1 U20478 ( .A1(n5607), .A2(n64157), .Z(n44143) );
  NAND2_X2 U20481 ( .A1(n63531), .A2(n64956), .ZN(n62535) );
  NAND3_X2 U20482 ( .A1(n62287), .A2(n33092), .A3(n3994), .ZN(n33109) );
  XOR2_X1 U20494 ( .A1(n25809), .A2(n62442), .Z(n2961) );
  NAND3_X2 U20496 ( .A1(n58457), .A2(n60817), .A3(n42720), .ZN(n25809) );
  NAND2_X2 U20497 ( .A1(n55654), .A2(n63382), .ZN(n62288) );
  NOR2_X2 U20498 ( .A1(n1603), .A2(n55486), .ZN(n19971) );
  XOR2_X1 U20499 ( .A1(n62289), .A2(n60502), .Z(n19311) );
  XOR2_X1 U20502 ( .A1(n14228), .A2(n189), .Z(n62289) );
  OAI21_X2 U20505 ( .A1(n35976), .A2(n35975), .B(n35974), .ZN(n57847) );
  INV_X2 U20506 ( .I(n462), .ZN(n62389) );
  XOR2_X1 U20510 ( .A1(n6889), .A2(n39721), .Z(n64642) );
  AOI22_X1 U20512 ( .A1(n29899), .A2(n29906), .B1(n31187), .B2(n29903), .ZN(
        n11530) );
  NOR2_X2 U20514 ( .A1(n8212), .A2(n12698), .ZN(n48101) );
  OAI21_X2 U20515 ( .A1(n62797), .A2(n7501), .B(n17915), .ZN(n3726) );
  OAI22_X1 U20517 ( .A1(n62479), .A2(n31189), .B1(n31177), .B2(n31182), .ZN(
        n25586) );
  NAND3_X2 U20518 ( .A1(n36035), .A2(n36036), .A3(n36044), .ZN(n39728) );
  NOR3_X2 U20519 ( .A1(n58504), .A2(n58503), .A3(n32815), .ZN(n36022) );
  XOR2_X1 U20520 ( .A1(n62292), .A2(n37634), .Z(n8387) );
  XOR2_X1 U20525 ( .A1(n37628), .A2(n8665), .Z(n62292) );
  XOR2_X1 U20527 ( .A1(n3099), .A2(n60854), .Z(n5265) );
  NAND2_X1 U20528 ( .A1(n62441), .A2(n63063), .ZN(n33353) );
  NAND3_X1 U20530 ( .A1(n32903), .A2(n22613), .A3(n32902), .ZN(n63323) );
  NAND2_X2 U20536 ( .A1(n62294), .A2(n20541), .ZN(n64735) );
  OAI21_X2 U20537 ( .A1(n55003), .A2(n55004), .B(n55442), .ZN(n62294) );
  NAND2_X2 U20538 ( .A1(n23439), .A2(n50065), .ZN(n52172) );
  INV_X2 U20542 ( .I(n62295), .ZN(n19973) );
  NOR2_X2 U20544 ( .A1(n62993), .A2(n55385), .ZN(n62295) );
  XOR2_X1 U20552 ( .A1(n62296), .A2(n56849), .Z(Plaintext[175]) );
  NAND4_X2 U20555 ( .A1(n17649), .A2(n64152), .A3(n17646), .A4(n17645), .ZN(
        n62296) );
  XOR2_X1 U20556 ( .A1(n16529), .A2(n5458), .Z(n37867) );
  NOR2_X2 U20565 ( .A1(n61914), .A2(n56417), .ZN(n56637) );
  NAND2_X2 U20572 ( .A1(n22273), .A2(n61921), .ZN(n26469) );
  INV_X2 U20573 ( .I(n62298), .ZN(n51112) );
  XNOR2_X1 U20579 ( .A1(n51068), .A2(n64091), .ZN(n62298) );
  NOR2_X1 U20586 ( .A1(n61693), .A2(n64712), .ZN(n53237) );
  NAND2_X2 U20587 ( .A1(n5536), .A2(n25649), .ZN(n64712) );
  NAND3_X1 U20588 ( .A1(n53536), .A2(n53534), .A3(n53535), .ZN(n7481) );
  BUF_X2 U20591 ( .I(n1716), .Z(n62299) );
  XOR2_X1 U20593 ( .A1(n8381), .A2(n44084), .Z(n25982) );
  NOR2_X2 U20594 ( .A1(n59731), .A2(n62302), .ZN(n23126) );
  NAND2_X2 U20595 ( .A1(n2160), .A2(n42694), .ZN(n42698) );
  NOR2_X2 U20598 ( .A1(n57592), .A2(n36034), .ZN(n17487) );
  NOR2_X2 U20601 ( .A1(n35576), .A2(n34822), .ZN(n36034) );
  NOR2_X2 U20603 ( .A1(n20521), .A2(n20522), .ZN(n24343) );
  NOR2_X2 U20606 ( .A1(n11806), .A2(n9740), .ZN(n11795) );
  XOR2_X1 U20608 ( .A1(n3269), .A2(n45357), .Z(n3268) );
  INV_X2 U20610 ( .I(n14846), .ZN(n1690) );
  NAND2_X2 U20613 ( .A1(n2330), .A2(n63205), .ZN(n14846) );
  NOR3_X2 U20618 ( .A1(n25361), .A2(n45640), .A3(n24597), .ZN(n25360) );
  NAND4_X2 U20620 ( .A1(n42708), .A2(n42705), .A3(n62304), .A4(n62303), .ZN(
        n22554) );
  AOI21_X2 U20622 ( .A1(n42700), .A2(n42699), .B(n62305), .ZN(n62304) );
  INV_X2 U20623 ( .I(n42707), .ZN(n62305) );
  XOR2_X1 U20625 ( .A1(n45844), .A2(n4264), .Z(n46543) );
  XOR2_X1 U20632 ( .A1(n25209), .A2(n24992), .Z(n4264) );
  OR2_X2 U20633 ( .A1(n61531), .A2(n29053), .Z(n2636) );
  NOR2_X2 U20638 ( .A1(n15947), .A2(n62306), .ZN(n22398) );
  NAND3_X2 U20646 ( .A1(n52921), .A2(n19903), .A3(n19902), .ZN(n62306) );
  NOR2_X1 U20648 ( .A1(n59557), .A2(n12486), .ZN(n61225) );
  NOR2_X2 U20649 ( .A1(n20055), .A2(n58205), .ZN(n49856) );
  NOR2_X2 U20651 ( .A1(n55214), .A2(n55200), .ZN(n59041) );
  XOR2_X1 U20652 ( .A1(n2779), .A2(n2782), .Z(n25569) );
  XOR2_X1 U20653 ( .A1(n1904), .A2(n14086), .Z(n64197) );
  XOR2_X1 U20666 ( .A1(n11011), .A2(n20772), .Z(n1904) );
  NAND2_X2 U20667 ( .A1(n39815), .A2(n39816), .ZN(n61388) );
  NOR3_X2 U20669 ( .A1(n20983), .A2(n39814), .A3(n24270), .ZN(n39815) );
  NAND2_X1 U20671 ( .A1(n56503), .A2(n10286), .ZN(n56504) );
  NAND2_X2 U20673 ( .A1(n23920), .A2(n20587), .ZN(n56503) );
  NAND3_X2 U20678 ( .A1(n2346), .A2(n10358), .A3(n59328), .ZN(n33437) );
  NAND2_X2 U20680 ( .A1(n3981), .A2(n23908), .ZN(n25994) );
  XOR2_X1 U20683 ( .A1(n10823), .A2(n6744), .Z(n5154) );
  XOR2_X1 U20684 ( .A1(n62309), .A2(n24105), .Z(Plaintext[156]) );
  NAND4_X2 U20686 ( .A1(n56448), .A2(n60257), .A3(n64855), .A4(n60256), .ZN(
        n62309) );
  NAND3_X2 U20688 ( .A1(n26069), .A2(n48323), .A3(n10563), .ZN(n48450) );
  XOR2_X1 U20691 ( .A1(n62310), .A2(n6965), .Z(n63766) );
  XOR2_X1 U20692 ( .A1(n51189), .A2(n1619), .Z(n62310) );
  XOR2_X1 U20698 ( .A1(n62311), .A2(n37527), .Z(n14864) );
  XOR2_X1 U20704 ( .A1(n14382), .A2(n57439), .Z(n62311) );
  XOR2_X1 U20705 ( .A1(n13689), .A2(n62312), .Z(n3270) );
  XOR2_X1 U20707 ( .A1(n45815), .A2(n44222), .Z(n62312) );
  BUF_X4 U20712 ( .I(n10064), .Z(n9608) );
  NAND2_X2 U20713 ( .A1(n43327), .A2(n61186), .ZN(n43316) );
  NAND2_X2 U20714 ( .A1(n62313), .A2(n42982), .ZN(n14627) );
  BUF_X2 U20715 ( .I(n14955), .Z(n62314) );
  NAND2_X1 U20716 ( .A1(n36844), .A2(n36847), .ZN(n16456) );
  AND2_X1 U20717 ( .A1(n41872), .A2(n42528), .Z(n63930) );
  NAND2_X2 U20731 ( .A1(n2646), .A2(n2645), .ZN(n23371) );
  NAND2_X2 U20733 ( .A1(n24557), .A2(n27865), .ZN(n64169) );
  XOR2_X1 U20738 ( .A1(n21289), .A2(n38119), .Z(n16796) );
  XOR2_X1 U20744 ( .A1(n10647), .A2(n10650), .Z(n62381) );
  NAND4_X2 U20749 ( .A1(n21684), .A2(n21683), .A3(n47268), .A4(n47269), .ZN(
        n48728) );
  INV_X1 U20755 ( .I(n6509), .ZN(n63168) );
  NOR3_X1 U20756 ( .A1(n63129), .A2(n30269), .A3(n30268), .ZN(n30283) );
  XOR2_X1 U20763 ( .A1(n51572), .A2(n50616), .Z(n62315) );
  NAND2_X2 U20764 ( .A1(n58372), .A2(n23211), .ZN(n7616) );
  NOR2_X1 U20765 ( .A1(n7154), .A2(n14311), .ZN(n64643) );
  XOR2_X1 U20770 ( .A1(n63768), .A2(n6438), .Z(n14970) );
  XOR2_X1 U20778 ( .A1(n59154), .A2(n38203), .Z(n6438) );
  XOR2_X1 U20781 ( .A1(n8782), .A2(n24908), .Z(n32556) );
  OAI22_X1 U20782 ( .A1(n34894), .A2(n35981), .B1(n34893), .B2(n35463), .ZN(
        n64312) );
  NAND3_X2 U20784 ( .A1(n35986), .A2(n60022), .A3(n20147), .ZN(n35463) );
  NAND3_X2 U20785 ( .A1(n64873), .A2(n6422), .A3(n6424), .ZN(n6425) );
  OAI22_X2 U20790 ( .A1(n34163), .A2(n34164), .B1(n34162), .B2(n34165), .ZN(
        n24036) );
  NOR2_X1 U20804 ( .A1(n32528), .A2(n4565), .ZN(n33689) );
  NAND2_X2 U20805 ( .A1(n12271), .A2(n62316), .ZN(n44388) );
  NOR4_X2 U20806 ( .A1(n41486), .A2(n41487), .A3(n41488), .A4(n42770), .ZN(
        n62316) );
  OAI21_X2 U20808 ( .A1(n62318), .A2(n4332), .B(n63205), .ZN(n4331) );
  NOR2_X2 U20810 ( .A1(n23541), .A2(n22606), .ZN(n62318) );
  XNOR2_X1 U20813 ( .A1(n12685), .A2(n63436), .ZN(n14827) );
  XOR2_X1 U20818 ( .A1(n6941), .A2(n64340), .Z(n12685) );
  INV_X2 U20821 ( .I(n62319), .ZN(n14994) );
  XNOR2_X1 U20826 ( .A1(n14997), .A2(n60714), .ZN(n62319) );
  XOR2_X1 U20839 ( .A1(n37174), .A2(n12879), .Z(n9019) );
  NAND2_X2 U20843 ( .A1(n5072), .A2(n62320), .ZN(n5163) );
  NOR3_X2 U20844 ( .A1(n5164), .A2(n5069), .A3(n61798), .ZN(n62320) );
  AOI22_X1 U20846 ( .A1(n62500), .A2(n35414), .B1(n35420), .B2(n34011), .ZN(
        n62450) );
  XOR2_X1 U20848 ( .A1(n44162), .A2(n578), .Z(n8237) );
  NAND2_X1 U20850 ( .A1(n52053), .A2(n9386), .ZN(n9382) );
  NAND4_X2 U20851 ( .A1(n9383), .A2(n9380), .A3(n9385), .A4(n9384), .ZN(n52053) );
  INV_X2 U20852 ( .I(n47429), .ZN(n62321) );
  OR2_X1 U20853 ( .A1(n10397), .A2(n62321), .Z(n47423) );
  XOR2_X1 U20854 ( .A1(n45290), .A2(n45291), .Z(n62403) );
  XOR2_X1 U20855 ( .A1(n10613), .A2(n25949), .Z(n25947) );
  AOI22_X1 U20856 ( .A1(n42133), .A2(n62388), .B1(n42132), .B2(n42131), .ZN(
        n42135) );
  AND3_X1 U20859 ( .A1(n24997), .A2(n11537), .A3(n11536), .Z(n61664) );
  NAND2_X2 U20861 ( .A1(n16863), .A2(n2495), .ZN(n30838) );
  NAND2_X2 U20862 ( .A1(n287), .A2(n1741), .ZN(n42240) );
  NAND2_X1 U20863 ( .A1(n35518), .A2(n35519), .ZN(n10096) );
  AND2_X2 U20865 ( .A1(n8470), .A2(n64192), .Z(n7376) );
  XOR2_X1 U20867 ( .A1(n8294), .A2(n18579), .Z(n20228) );
  NAND2_X2 U20871 ( .A1(n3302), .A2(n18742), .ZN(n43272) );
  NAND2_X2 U20872 ( .A1(n18743), .A2(n18746), .ZN(n3302) );
  XOR2_X1 U20873 ( .A1(n6181), .A2(n61775), .Z(n23489) );
  NAND2_X2 U20878 ( .A1(n15110), .A2(n1930), .ZN(n15109) );
  NAND2_X2 U20879 ( .A1(n21774), .A2(n3087), .ZN(n1930) );
  XOR2_X1 U20881 ( .A1(n9463), .A2(n20580), .Z(n8417) );
  XOR2_X1 U20891 ( .A1(n8418), .A2(n13359), .Z(n9463) );
  INV_X4 U20893 ( .I(n22050), .ZN(n26020) );
  NAND2_X2 U20904 ( .A1(n62436), .A2(n22051), .ZN(n22050) );
  OAI22_X1 U20909 ( .A1(n54806), .A2(n7518), .B1(n1146), .B2(n54300), .ZN(
        n64690) );
  NAND2_X1 U20915 ( .A1(n61824), .A2(n62325), .ZN(n57848) );
  XOR2_X1 U20919 ( .A1(n16885), .A2(n25964), .Z(n62325) );
  BUF_X2 U20927 ( .I(n16527), .Z(n62326) );
  AOI21_X2 U20929 ( .A1(n62330), .A2(n1457), .B(n10869), .ZN(n62329) );
  INV_X2 U20930 ( .I(n62331), .ZN(n57173) );
  XNOR2_X1 U20931 ( .A1(n2970), .A2(n58292), .ZN(n62331) );
  AOI22_X2 U20934 ( .A1(n17675), .A2(n1628), .B1(n4624), .B2(n63712), .ZN(
        n63627) );
  OR2_X1 U20935 ( .A1(n3302), .A2(n13493), .Z(n43273) );
  OR2_X1 U20947 ( .A1(n56981), .A2(n56980), .Z(n64113) );
  BUF_X4 U20948 ( .I(n17173), .Z(n17171) );
  NOR3_X2 U20950 ( .A1(n42769), .A2(n62332), .A3(n42770), .ZN(n10152) );
  OAI21_X1 U20952 ( .A1(n12905), .A2(n42930), .B(n12904), .ZN(n12903) );
  AND2_X1 U20967 ( .A1(n42117), .A2(n15007), .Z(n62432) );
  NAND2_X1 U20969 ( .A1(n15026), .A2(n18925), .ZN(n54278) );
  NAND2_X2 U20970 ( .A1(n54542), .A2(n22217), .ZN(n54568) );
  NOR2_X2 U20980 ( .A1(n59049), .A2(n54450), .ZN(n54542) );
  NOR2_X1 U20985 ( .A1(n3708), .A2(n15023), .ZN(n54827) );
  NAND2_X2 U20994 ( .A1(n15040), .A2(n2489), .ZN(n3708) );
  BUF_X2 U20996 ( .I(n24429), .Z(n62334) );
  OAI22_X2 U20997 ( .A1(n39048), .A2(n39047), .B1(n39050), .B2(n57925), .ZN(
        n19992) );
  NOR3_X1 U20998 ( .A1(n54443), .A2(n1371), .A3(n54823), .ZN(n54445) );
  AND2_X1 U21006 ( .A1(n11460), .A2(n9396), .Z(n9436) );
  XOR2_X1 U21007 ( .A1(n2061), .A2(n2060), .Z(n62455) );
  XOR2_X1 U21010 ( .A1(n5403), .A2(n5406), .Z(n54689) );
  XOR2_X1 U21020 ( .A1(n5405), .A2(n5404), .Z(n5403) );
  INV_X2 U21023 ( .I(n39081), .ZN(n42786) );
  AOI21_X2 U21029 ( .A1(n35874), .A2(n35873), .B(n62335), .ZN(n16531) );
  AOI21_X2 U21032 ( .A1(n5442), .A2(n61574), .B(n37007), .ZN(n62335) );
  XOR2_X1 U21033 ( .A1(n62337), .A2(n62336), .Z(n59786) );
  XOR2_X1 U21039 ( .A1(n51807), .A2(n51507), .Z(n62336) );
  XOR2_X1 U21040 ( .A1(n62377), .A2(n16006), .Z(n62337) );
  AND2_X1 U21043 ( .A1(n14178), .A2(n399), .Z(n53415) );
  NAND3_X2 U21046 ( .A1(n46863), .A2(n46027), .A3(n46028), .ZN(n45723) );
  NAND3_X1 U21047 ( .A1(n48976), .A2(n48975), .A3(n49850), .ZN(n48374) );
  NOR2_X2 U21049 ( .A1(n45589), .A2(n25637), .ZN(n49850) );
  NAND2_X1 U21051 ( .A1(n41999), .A2(n41998), .ZN(n64570) );
  XOR2_X1 U21052 ( .A1(n62338), .A2(n53124), .Z(Plaintext[5]) );
  NAND4_X1 U21059 ( .A1(n53121), .A2(n53123), .A3(n53120), .A4(n53122), .ZN(
        n62338) );
  AOI21_X2 U21063 ( .A1(n4029), .A2(n62339), .B(n4027), .ZN(n20625) );
  XOR2_X1 U21068 ( .A1(n7601), .A2(n64640), .Z(n38911) );
  INV_X4 U21070 ( .I(n12502), .ZN(n25348) );
  NOR2_X1 U21074 ( .A1(n59229), .A2(n62340), .ZN(n2793) );
  NAND2_X2 U21076 ( .A1(n57939), .A2(n4304), .ZN(n20020) );
  XOR2_X1 U21077 ( .A1(n46305), .A2(n42984), .Z(n44994) );
  NOR2_X2 U21078 ( .A1(n21682), .A2(n21681), .ZN(n42984) );
  NOR2_X2 U21079 ( .A1(n50043), .A2(n3348), .ZN(n49358) );
  XOR2_X1 U21084 ( .A1(n51119), .A2(n5778), .Z(n2487) );
  AOI21_X2 U21085 ( .A1(n3472), .A2(n23575), .B(n64225), .ZN(n58506) );
  NAND2_X2 U21087 ( .A1(n7303), .A2(n22885), .ZN(n62343) );
  NAND2_X2 U21088 ( .A1(n2021), .A2(n62344), .ZN(n2023) );
  AND3_X1 U21090 ( .A1(n12160), .A2(n29925), .A3(n14109), .Z(n62344) );
  XOR2_X1 U21101 ( .A1(n14969), .A2(n39716), .Z(n38446) );
  AND2_X1 U21109 ( .A1(n14863), .A2(n57173), .Z(n41816) );
  NOR2_X1 U21110 ( .A1(n44700), .A2(n45779), .ZN(n63172) );
  OAI21_X1 U21115 ( .A1(n63172), .A2(n63171), .B(n61166), .ZN(n19325) );
  NAND2_X2 U21118 ( .A1(n23484), .A2(n40387), .ZN(n63119) );
  XOR2_X1 U21119 ( .A1(n51804), .A2(n23571), .Z(n51509) );
  NAND2_X2 U21127 ( .A1(n3920), .A2(n3917), .ZN(n23571) );
  OR2_X1 U21129 ( .A1(n63047), .A2(n62896), .Z(n62693) );
  NOR3_X2 U21130 ( .A1(n7563), .A2(n33588), .A3(n7562), .ZN(n62345) );
  BUF_X4 U21131 ( .I(n33110), .Z(n36898) );
  AOI22_X2 U21132 ( .A1(n36520), .A2(n2594), .B1(n36589), .B2(n37375), .ZN(
        n62473) );
  NAND3_X2 U21133 ( .A1(n27112), .A2(n25800), .A3(n25801), .ZN(n28959) );
  NAND3_X2 U21135 ( .A1(n52821), .A2(n53439), .A3(n53436), .ZN(n23624) );
  INV_X2 U21136 ( .I(n14255), .ZN(n22234) );
  NAND2_X1 U21140 ( .A1(n764), .A2(n27559), .ZN(n14255) );
  XOR2_X1 U21143 ( .A1(n2583), .A2(n23898), .Z(n37628) );
  NAND2_X2 U21144 ( .A1(n62348), .A2(n61713), .ZN(n15401) );
  NOR3_X2 U21151 ( .A1(n60609), .A2(n43704), .A3(n60608), .ZN(n62348) );
  XOR2_X1 U21153 ( .A1(n32354), .A2(n62349), .Z(n30904) );
  XOR2_X1 U21154 ( .A1(n30901), .A2(n9977), .Z(n62349) );
  INV_X1 U21155 ( .I(n31873), .ZN(n62356) );
  NAND3_X1 U21158 ( .A1(n53087), .A2(n53089), .A3(n53088), .ZN(n63901) );
  NOR2_X2 U21165 ( .A1(n13395), .A2(n8394), .ZN(n7259) );
  NOR2_X2 U21170 ( .A1(n65110), .A2(n40829), .ZN(n13395) );
  NOR2_X1 U21173 ( .A1(n14484), .A2(n56958), .ZN(n7565) );
  NAND2_X2 U21176 ( .A1(n138), .A2(n3021), .ZN(n14484) );
  XNOR2_X1 U21178 ( .A1(n12957), .A2(n51940), .ZN(n63918) );
  NAND2_X2 U21179 ( .A1(n25951), .A2(n57921), .ZN(n12957) );
  XOR2_X1 U21182 ( .A1(n1676), .A2(n5214), .Z(n4900) );
  XOR2_X1 U21186 ( .A1(n5911), .A2(n62350), .Z(n37648) );
  XOR2_X1 U21187 ( .A1(n39757), .A2(n11013), .Z(n62350) );
  INV_X4 U21190 ( .I(n13393), .ZN(n42944) );
  XOR2_X1 U21191 ( .A1(n25111), .A2(n17624), .Z(n6765) );
  NAND2_X2 U21193 ( .A1(n7546), .A2(n17625), .ZN(n17624) );
  INV_X4 U21195 ( .I(n24370), .ZN(n37945) );
  NAND3_X2 U21198 ( .A1(n63387), .A2(n63388), .A3(n24371), .ZN(n24370) );
  INV_X2 U21201 ( .I(n15271), .ZN(n23168) );
  NAND3_X2 U21205 ( .A1(n60450), .A2(n2544), .A3(n13623), .ZN(n15271) );
  OAI21_X2 U21206 ( .A1(n62352), .A2(n62351), .B(n33081), .ZN(n33088) );
  XOR2_X1 U21207 ( .A1(n62356), .A2(n62354), .Z(n24154) );
  NAND2_X2 U21208 ( .A1(n62355), .A2(n24156), .ZN(n62354) );
  AND2_X1 U21210 ( .A1(n24155), .A2(n11816), .Z(n62355) );
  XOR2_X1 U21211 ( .A1(n15722), .A2(n60394), .Z(n51731) );
  XOR2_X1 U21216 ( .A1(n45373), .A2(n57630), .Z(n12234) );
  INV_X2 U21221 ( .I(n44569), .ZN(n21406) );
  NOR2_X1 U21233 ( .A1(n40202), .A2(n40201), .ZN(n11494) );
  NAND2_X2 U21235 ( .A1(n60843), .A2(n7451), .ZN(n43343) );
  NOR2_X2 U21255 ( .A1(n62359), .A2(n5792), .ZN(n5791) );
  NAND2_X2 U21256 ( .A1(n5790), .A2(n17077), .ZN(n62359) );
  NOR2_X1 U21257 ( .A1(n58727), .A2(n58728), .ZN(n64508) );
  XOR2_X1 U21259 ( .A1(n44377), .A2(n8214), .Z(n24798) );
  XOR2_X1 U21261 ( .A1(n12153), .A2(n54249), .Z(n44377) );
  OR2_X1 U21264 ( .A1(n37233), .A2(n12798), .Z(n36973) );
  XOR2_X1 U21266 ( .A1(n9255), .A2(n38080), .Z(n59720) );
  NAND2_X1 U21270 ( .A1(n37829), .A2(n18892), .ZN(n62362) );
  NOR2_X2 U21274 ( .A1(n9789), .A2(n62360), .ZN(n50096) );
  NAND4_X2 U21275 ( .A1(n46800), .A2(n46802), .A3(n46801), .A4(n46799), .ZN(
        n62360) );
  XOR2_X1 U21277 ( .A1(n51481), .A2(n51482), .Z(n51677) );
  NAND3_X2 U21278 ( .A1(n21602), .A2(n46975), .A3(n50751), .ZN(n51481) );
  NAND3_X2 U21279 ( .A1(n23357), .A2(n61935), .A3(n37210), .ZN(n64164) );
  XOR2_X1 U21281 ( .A1(n62361), .A2(n24067), .Z(Plaintext[19]) );
  NAND3_X2 U21284 ( .A1(n52813), .A2(n52812), .A3(n52811), .ZN(n62361) );
  AND2_X2 U21287 ( .A1(n8854), .A2(n25803), .Z(n21028) );
  XOR2_X1 U21288 ( .A1(n648), .A2(n8629), .Z(n61156) );
  NAND2_X2 U21290 ( .A1(n7958), .A2(n7957), .ZN(n8629) );
  XOR2_X1 U21298 ( .A1(n52415), .A2(n50616), .Z(n3184) );
  XOR2_X1 U21302 ( .A1(n6004), .A2(n52538), .Z(n52415) );
  INV_X1 U21304 ( .I(n64531), .ZN(n43108) );
  NAND2_X2 U21307 ( .A1(n31767), .A2(n18390), .ZN(n18678) );
  AOI21_X1 U21308 ( .A1(n56925), .A2(n14484), .B(n21370), .ZN(n21514) );
  AOI21_X1 U21312 ( .A1(n37825), .A2(n40848), .B(n62362), .ZN(n754) );
  XOR2_X1 U21313 ( .A1(n5098), .A2(n62363), .Z(n62603) );
  XOR2_X1 U21321 ( .A1(n11508), .A2(n8354), .Z(n62363) );
  NOR2_X2 U21323 ( .A1(n57194), .A2(n16985), .ZN(n4436) );
  INV_X2 U21324 ( .I(n18887), .ZN(n20230) );
  NOR2_X2 U21326 ( .A1(n62364), .A2(n14510), .ZN(n44456) );
  NAND2_X2 U21331 ( .A1(n4657), .A2(n2197), .ZN(n62364) );
  XOR2_X1 U21332 ( .A1(n14605), .A2(n61739), .Z(n1024) );
  NOR2_X2 U21339 ( .A1(n42968), .A2(n1336), .ZN(n43462) );
  INV_X4 U21343 ( .I(n43460), .ZN(n1336) );
  XOR2_X1 U21344 ( .A1(n3118), .A2(n2361), .Z(n2933) );
  NAND3_X2 U21345 ( .A1(n39140), .A2(n20393), .A3(n20392), .ZN(n462) );
  NAND3_X2 U21347 ( .A1(n8656), .A2(n8653), .A3(n8655), .ZN(n12178) );
  NAND3_X2 U21348 ( .A1(n42336), .A2(n62367), .A3(n42334), .ZN(n42337) );
  NOR2_X2 U21351 ( .A1(n42259), .A2(n42267), .ZN(n42261) );
  INV_X1 U21365 ( .I(n41898), .ZN(n62368) );
  XOR2_X1 U21366 ( .A1(n62369), .A2(n61807), .Z(n24284) );
  XOR2_X1 U21367 ( .A1(n18187), .A2(n10575), .Z(n62369) );
  AND2_X1 U21371 ( .A1(n36401), .A2(n36116), .Z(n36115) );
  NAND2_X2 U21372 ( .A1(n62370), .A2(n53445), .ZN(n57056) );
  XOR2_X1 U21373 ( .A1(n51617), .A2(n26047), .Z(n18189) );
  XOR2_X1 U21386 ( .A1(n9416), .A2(n51209), .Z(n51617) );
  XOR2_X1 U21387 ( .A1(n62371), .A2(n17737), .Z(n12585) );
  XOR2_X1 U21388 ( .A1(n50802), .A2(n12257), .Z(n62371) );
  NAND2_X2 U21389 ( .A1(n57757), .A2(n57758), .ZN(n57569) );
  XOR2_X1 U21394 ( .A1(n46231), .A2(n63872), .Z(n2574) );
  NAND3_X2 U21406 ( .A1(n7795), .A2(n63222), .A3(n7794), .ZN(n46231) );
  NAND2_X2 U21407 ( .A1(n62372), .A2(n57710), .ZN(n32210) );
  OAI21_X2 U21408 ( .A1(n7660), .A2(n32208), .B(n3308), .ZN(n62372) );
  NAND2_X2 U21409 ( .A1(n34161), .A2(n23947), .ZN(n34167) );
  AOI22_X1 U21410 ( .A1(n52860), .A2(n52859), .B1(n13567), .B2(n61516), .ZN(
        n17177) );
  NAND3_X2 U21412 ( .A1(n28726), .A2(n20551), .A3(n30776), .ZN(n30550) );
  INV_X2 U21417 ( .I(n19802), .ZN(n47141) );
  NAND2_X2 U21421 ( .A1(n16457), .A2(n61358), .ZN(n39310) );
  NAND3_X2 U21422 ( .A1(n13102), .A2(n62374), .A3(n7033), .ZN(n5928) );
  NAND2_X1 U21423 ( .A1(n39178), .A2(n39179), .ZN(n62398) );
  NOR2_X1 U21429 ( .A1(n13971), .A2(n45561), .ZN(n13970) );
  NAND4_X2 U21432 ( .A1(n63378), .A2(n39883), .A3(n62376), .A4(n62375), .ZN(
        n22143) );
  XOR2_X1 U21433 ( .A1(n59758), .A2(n8104), .Z(n8103) );
  XNOR2_X1 U21435 ( .A1(n13695), .A2(n18555), .ZN(n63905) );
  NAND3_X2 U21436 ( .A1(n63108), .A2(n63107), .A3(n63829), .ZN(n6410) );
  NOR2_X2 U21438 ( .A1(n10211), .A2(n10210), .ZN(n11983) );
  XOR2_X1 U21439 ( .A1(n24594), .A2(n11360), .Z(n24730) );
  AOI21_X2 U21441 ( .A1(n28091), .A2(n13573), .B(n1277), .ZN(n8703) );
  XOR2_X1 U21447 ( .A1(n62590), .A2(n19711), .Z(n62377) );
  XOR2_X1 U21448 ( .A1(n6731), .A2(n10802), .Z(n65019) );
  NAND3_X2 U21449 ( .A1(n10706), .A2(n18990), .A3(n10803), .ZN(n10802) );
  NOR3_X2 U21450 ( .A1(n43233), .A2(n43234), .A3(n11635), .ZN(n62433) );
  AND2_X2 U21451 ( .A1(n59786), .A2(n64635), .Z(n59294) );
  INV_X1 U21452 ( .I(n14315), .ZN(n63357) );
  XOR2_X1 U21453 ( .A1(n62378), .A2(n45400), .Z(n17438) );
  XOR2_X1 U21454 ( .A1(n244), .A2(n53064), .Z(n62378) );
  XOR2_X1 U21455 ( .A1(n62379), .A2(n14588), .Z(n13221) );
  XOR2_X1 U21459 ( .A1(n19803), .A2(n15664), .Z(n62379) );
  NOR2_X2 U21462 ( .A1(n40797), .A2(n41914), .ZN(n41263) );
  BUF_X2 U21463 ( .I(n16594), .Z(n62380) );
  INV_X2 U21468 ( .I(n25058), .ZN(n36612) );
  NAND2_X2 U21475 ( .A1(n58250), .A2(n59617), .ZN(n25058) );
  XOR2_X1 U21476 ( .A1(n62381), .A2(n11341), .Z(n11340) );
  NAND3_X2 U21480 ( .A1(n43526), .A2(n43525), .A3(n62382), .ZN(n46150) );
  XOR2_X1 U21481 ( .A1(n38891), .A2(n38890), .Z(n62383) );
  NOR2_X1 U21482 ( .A1(n11031), .A2(n7254), .ZN(n8083) );
  INV_X2 U21486 ( .I(n60793), .ZN(n32528) );
  INV_X2 U21487 ( .I(n62384), .ZN(n63185) );
  NAND2_X1 U21492 ( .A1(n60793), .A2(n61523), .ZN(n62384) );
  XOR2_X1 U21493 ( .A1(n60303), .A2(n60302), .Z(n60793) );
  NAND3_X2 U21495 ( .A1(n48316), .A2(n49939), .A3(n48315), .ZN(n11678) );
  NOR2_X1 U21497 ( .A1(n56466), .A2(n62385), .ZN(n56448) );
  AND2_X1 U21498 ( .A1(n56523), .A2(n23920), .Z(n62385) );
  XOR2_X1 U21500 ( .A1(n11858), .A2(n62386), .Z(n11857) );
  XOR2_X1 U21506 ( .A1(n2723), .A2(n2724), .Z(n62386) );
  NAND2_X1 U21507 ( .A1(n57173), .A2(n59168), .ZN(n42428) );
  NAND2_X2 U21509 ( .A1(n61716), .A2(n5481), .ZN(n20055) );
  NAND3_X2 U21510 ( .A1(n5482), .A2(n20019), .A3(n7035), .ZN(n5481) );
  NAND2_X2 U21511 ( .A1(n19666), .A2(n62387), .ZN(n8819) );
  NOR2_X2 U21512 ( .A1(n35918), .A2(n8509), .ZN(n62387) );
  INV_X2 U21513 ( .I(n42325), .ZN(n20400) );
  NAND2_X2 U21515 ( .A1(n62389), .A2(n57873), .ZN(n42325) );
  NAND4_X1 U21516 ( .A1(n52292), .A2(n52291), .A3(n52293), .A4(n60644), .ZN(
        n62568) );
  NOR2_X2 U21527 ( .A1(n44406), .A2(n44405), .ZN(n23581) );
  OR2_X1 U21531 ( .A1(n22835), .A2(n8009), .Z(n35782) );
  INV_X2 U21534 ( .I(n41540), .ZN(n62391) );
  XOR2_X1 U21535 ( .A1(n62392), .A2(n54153), .Z(Plaintext[56]) );
  NAND3_X1 U21537 ( .A1(n54152), .A2(n54151), .A3(n54193), .ZN(n62392) );
  NAND2_X2 U21541 ( .A1(n47142), .A2(n19802), .ZN(n19801) );
  XOR2_X1 U21543 ( .A1(n17025), .A2(n16522), .Z(n16521) );
  XOR2_X1 U21548 ( .A1(n51179), .A2(n51400), .Z(n4811) );
  XOR2_X1 U21549 ( .A1(n14609), .A2(n3318), .Z(n51179) );
  XOR2_X1 U21551 ( .A1(n14356), .A2(n51692), .Z(n59508) );
  NAND2_X1 U21554 ( .A1(n35091), .A2(n37940), .ZN(n6909) );
  NAND2_X2 U21562 ( .A1(n48543), .A2(n62393), .ZN(n48157) );
  NOR3_X1 U21564 ( .A1(n48148), .A2(n20517), .A3(n18100), .ZN(n62393) );
  NAND3_X1 U21566 ( .A1(n6236), .A2(n41466), .A3(n39809), .ZN(n14800) );
  XOR2_X1 U21567 ( .A1(n62395), .A2(n62394), .Z(n40928) );
  XOR2_X1 U21568 ( .A1(n65239), .A2(n59284), .Z(n62395) );
  NAND3_X1 U21570 ( .A1(n8083), .A2(n8084), .A3(n8085), .ZN(n65093) );
  INV_X2 U21572 ( .I(n62396), .ZN(n24571) );
  XNOR2_X1 U21580 ( .A1(n18873), .A2(n57730), .ZN(n62396) );
  NAND2_X2 U21587 ( .A1(n64537), .A2(n27519), .ZN(n33862) );
  XOR2_X1 U21588 ( .A1(n24686), .A2(n46688), .Z(n62562) );
  NAND2_X1 U21593 ( .A1(n36619), .A2(n36616), .ZN(n59337) );
  XOR2_X1 U21597 ( .A1(n8673), .A2(n7850), .Z(n8418) );
  XOR2_X1 U21601 ( .A1(n3750), .A2(n10939), .Z(n7850) );
  NOR4_X2 U21602 ( .A1(n40286), .A2(n5541), .A3(n4648), .A4(n4649), .ZN(n57252) );
  NAND2_X2 U21605 ( .A1(n15336), .A2(n18590), .ZN(n18589) );
  NAND2_X2 U21606 ( .A1(n56407), .A2(n4634), .ZN(n56580) );
  XOR2_X1 U21609 ( .A1(n62400), .A2(n59581), .Z(n47749) );
  XOR2_X1 U21617 ( .A1(n64402), .A2(n14935), .Z(n62400) );
  NOR2_X2 U21622 ( .A1(n41446), .A2(n41445), .ZN(n40378) );
  NAND2_X2 U21625 ( .A1(n1219), .A2(n39847), .ZN(n41446) );
  BUF_X4 U21640 ( .I(n56000), .Z(n56047) );
  INV_X2 U21643 ( .I(n34736), .ZN(n62401) );
  NAND3_X2 U21644 ( .A1(n3970), .A2(n3969), .A3(n61711), .ZN(n3966) );
  NOR3_X1 U21645 ( .A1(n27964), .A2(n62402), .A3(n26255), .ZN(n7715) );
  NOR2_X1 U21647 ( .A1(n26252), .A2(n28275), .ZN(n62402) );
  NAND2_X2 U21648 ( .A1(n49166), .A2(n25128), .ZN(n49551) );
  XOR2_X1 U21652 ( .A1(n62403), .A2(n18695), .Z(n10721) );
  OAI22_X1 U21653 ( .A1(n23077), .A2(n59205), .B1(n1649), .B2(n21200), .ZN(
        n64704) );
  NOR2_X1 U21655 ( .A1(n62404), .A2(n57001), .ZN(n57555) );
  NAND2_X2 U21658 ( .A1(n22114), .A2(n23836), .ZN(n57001) );
  NAND2_X1 U21662 ( .A1(n64712), .A2(n57470), .ZN(n62404) );
  XOR2_X1 U21663 ( .A1(n50576), .A2(n52323), .Z(n11322) );
  NAND2_X2 U21664 ( .A1(n25549), .A2(n10486), .ZN(n52323) );
  BUF_X2 U21669 ( .I(n4174), .Z(n62405) );
  BUF_X2 U21670 ( .I(n21087), .Z(n62406) );
  AOI21_X2 U21674 ( .A1(n1075), .A2(n48461), .B(n14611), .ZN(n62407) );
  NOR2_X2 U21675 ( .A1(n43077), .A2(n22673), .ZN(n43850) );
  INV_X2 U21688 ( .I(n62408), .ZN(n43077) );
  NAND2_X2 U21693 ( .A1(n43845), .A2(n39935), .ZN(n62408) );
  XOR2_X1 U21695 ( .A1(n62183), .A2(n3388), .Z(n61030) );
  NOR2_X2 U21699 ( .A1(n35962), .A2(n23577), .ZN(n15071) );
  NAND2_X2 U21702 ( .A1(n62409), .A2(n13493), .ZN(n57177) );
  INV_X2 U21703 ( .I(n18742), .ZN(n62409) );
  NAND2_X2 U21709 ( .A1(n39522), .A2(n39521), .ZN(n18742) );
  NAND3_X2 U21712 ( .A1(n62410), .A2(n24681), .A3(n6804), .ZN(n49728) );
  NAND2_X2 U21713 ( .A1(n46729), .A2(n46727), .ZN(n62410) );
  XOR2_X1 U21715 ( .A1(n58573), .A2(n1329), .Z(n64351) );
  XOR2_X1 U21716 ( .A1(n62411), .A2(n23162), .Z(n64343) );
  NAND2_X2 U21718 ( .A1(n64770), .A2(n17397), .ZN(n23162) );
  BUF_X2 U21719 ( .I(n53078), .Z(n62412) );
  NAND2_X2 U21724 ( .A1(n57184), .A2(n19974), .ZN(n62993) );
  NOR2_X2 U21725 ( .A1(n19980), .A2(n19981), .ZN(n19974) );
  XOR2_X1 U21730 ( .A1(n49727), .A2(n18870), .Z(n6386) );
  XOR2_X1 U21731 ( .A1(n50695), .A2(n22741), .Z(n49727) );
  BUF_X2 U21733 ( .I(n16765), .Z(n62413) );
  XOR2_X1 U21734 ( .A1(n15500), .A2(n5522), .Z(n39564) );
  INV_X2 U21743 ( .I(n13808), .ZN(n15500) );
  XOR2_X1 U21744 ( .A1(n39343), .A2(n7857), .Z(n13808) );
  BUF_X2 U21750 ( .I(n1556), .Z(n62414) );
  XOR2_X1 U21758 ( .A1(n31293), .A2(n15153), .Z(n2862) );
  XOR2_X1 U21759 ( .A1(n33828), .A2(n30828), .Z(n31293) );
  NAND3_X2 U21773 ( .A1(n17391), .A2(n17389), .A3(n62415), .ZN(n18072) );
  BUF_X2 U21775 ( .I(n961), .Z(n62416) );
  INV_X1 U21785 ( .I(n35646), .ZN(n62417) );
  AND2_X1 U21788 ( .A1(n6829), .A2(n62417), .Z(n7563) );
  NAND2_X1 U21789 ( .A1(n17799), .A2(n58808), .ZN(n52966) );
  NOR2_X2 U21790 ( .A1(n62602), .A2(n59041), .ZN(n55190) );
  NOR2_X1 U21792 ( .A1(n53592), .A2(n53593), .ZN(n53594) );
  NOR3_X2 U21794 ( .A1(n51906), .A2(n51907), .A3(n1138), .ZN(n63229) );
  AOI22_X1 U21804 ( .A1(n53700), .A2(n53690), .B1(n53691), .B2(n53692), .ZN(
        n53693) );
  XOR2_X1 U21805 ( .A1(n13678), .A2(n65262), .Z(n62418) );
  NAND2_X2 U21806 ( .A1(n62416), .A2(n41435), .ZN(n41440) );
  AOI21_X1 U21809 ( .A1(n55231), .A2(n7200), .B(n52965), .ZN(n58119) );
  BUF_X2 U21816 ( .I(n35685), .Z(n23313) );
  NAND3_X1 U21817 ( .A1(n42498), .A2(n41274), .A3(n2787), .ZN(n39934) );
  NOR2_X2 U21819 ( .A1(n4171), .A2(n19438), .ZN(n40320) );
  NAND2_X2 U21821 ( .A1(n63933), .A2(n11041), .ZN(n11999) );
  XOR2_X1 U21824 ( .A1(n8042), .A2(n44269), .Z(n7810) );
  NAND3_X2 U21826 ( .A1(n11749), .A2(n62419), .A3(n11156), .ZN(n44098) );
  NOR2_X1 U21827 ( .A1(n64583), .A2(n44859), .ZN(n44866) );
  NAND2_X1 U21828 ( .A1(n45637), .A2(n45638), .ZN(n62614) );
  NOR2_X1 U21839 ( .A1(n62614), .A2(n62613), .ZN(n62612) );
  NOR2_X2 U21840 ( .A1(n13408), .A2(n62420), .ZN(n331) );
  OR2_X1 U21843 ( .A1(n7366), .A2(n42066), .Z(n62420) );
  NAND2_X1 U21847 ( .A1(n56487), .A2(n56488), .ZN(n64365) );
  OR2_X1 U21859 ( .A1(n12521), .A2(n6540), .Z(n63957) );
  XOR2_X1 U21866 ( .A1(n51158), .A2(n62422), .Z(n24314) );
  XOR2_X1 U21867 ( .A1(n51156), .A2(n51155), .Z(n62422) );
  INV_X1 U21870 ( .I(n13888), .ZN(n62423) );
  AOI21_X1 U21872 ( .A1(n52739), .A2(n57018), .B(n57024), .ZN(n62444) );
  NAND3_X2 U21883 ( .A1(n42414), .A2(n15122), .A3(n42416), .ZN(n62860) );
  AOI22_X1 U21886 ( .A1(n1179), .A2(n15361), .B1(n1448), .B2(n19838), .ZN(
        n62443) );
  BUF_X2 U21888 ( .I(n47834), .Z(n62424) );
  XOR2_X1 U21889 ( .A1(n39223), .A2(n37821), .Z(n38314) );
  NAND2_X1 U21890 ( .A1(n24330), .A2(n48320), .ZN(n64955) );
  NOR2_X2 U21894 ( .A1(n62426), .A2(n62425), .ZN(n19248) );
  NAND2_X2 U21899 ( .A1(n7314), .A2(n38047), .ZN(n62425) );
  XOR2_X1 U21900 ( .A1(n50686), .A2(n62428), .Z(n2225) );
  XOR2_X1 U21901 ( .A1(n2230), .A2(n58296), .Z(n62428) );
  XOR2_X1 U21908 ( .A1(n1464), .A2(n6502), .Z(n63277) );
  XOR2_X1 U21910 ( .A1(n7843), .A2(n7844), .Z(n52408) );
  XOR2_X1 U21911 ( .A1(n44896), .A2(n64010), .Z(n62644) );
  XOR2_X1 U21914 ( .A1(n4068), .A2(n43781), .Z(n44896) );
  NOR2_X1 U21915 ( .A1(n20312), .A2(n33996), .ZN(n62429) );
  AOI22_X1 U21916 ( .A1(n11030), .A2(n57830), .B1(n10067), .B2(n11029), .ZN(
        n8084) );
  NAND3_X2 U21919 ( .A1(n1010), .A2(n62431), .A3(n62430), .ZN(n43453) );
  NOR3_X2 U21938 ( .A1(n23810), .A2(n23809), .A3(n15659), .ZN(n62430) );
  NOR2_X2 U21949 ( .A1(n62432), .A2(n15657), .ZN(n62431) );
  XOR2_X1 U21951 ( .A1(n52458), .A2(n13622), .Z(n64523) );
  XOR2_X1 U21954 ( .A1(n26044), .A2(n24274), .Z(n1910) );
  OAI21_X2 U21956 ( .A1(n62433), .A2(n43240), .B(n59672), .ZN(n43249) );
  OR2_X1 U21957 ( .A1(n14977), .A2(n12944), .Z(n56256) );
  XOR2_X1 U21959 ( .A1(n16202), .A2(n44941), .Z(n12921) );
  XOR2_X1 U21963 ( .A1(n45108), .A2(n24068), .Z(n16202) );
  NOR3_X2 U21964 ( .A1(n62439), .A2(n41759), .A3(n62438), .ZN(n58939) );
  INV_X2 U21967 ( .I(n20230), .ZN(n20232) );
  NOR2_X1 U21968 ( .A1(n33702), .A2(n33695), .ZN(n62440) );
  OR4_X1 U21971 ( .A1(n11038), .A2(n33698), .A3(n33704), .A4(n63064), .Z(
        n62441) );
  NOR2_X2 U21973 ( .A1(n57075), .A2(n57074), .ZN(n52858) );
  NOR2_X2 U21974 ( .A1(n63790), .A2(n51472), .ZN(n59374) );
  NOR2_X1 U21976 ( .A1(n45170), .A2(n64143), .ZN(n64540) );
  NAND2_X2 U21977 ( .A1(n43898), .A2(n3696), .ZN(n43243) );
  OAI21_X1 U21979 ( .A1(n65157), .A2(n19836), .B(n62443), .ZN(Plaintext[23])
         );
  AOI21_X1 U21980 ( .A1(n19833), .A2(n16769), .B(n62444), .ZN(n16768) );
  OAI21_X1 U21982 ( .A1(n53237), .A2(n20341), .B(n62517), .ZN(n62448) );
  NAND3_X2 U21983 ( .A1(n55305), .A2(n19978), .A3(n19977), .ZN(n19981) );
  XOR2_X1 U21985 ( .A1(n62449), .A2(n39307), .Z(n64025) );
  XOR2_X1 U21987 ( .A1(n4105), .A2(n11239), .Z(n62449) );
  AND2_X2 U21988 ( .A1(n24749), .A2(n63705), .Z(n8203) );
  AND2_X2 U21991 ( .A1(n60388), .A2(n62450), .Z(n21238) );
  CLKBUF_X8 U21993 ( .I(n50427), .Z(n63876) );
  XOR2_X1 U21997 ( .A1(n46499), .A2(n46498), .Z(n46509) );
  XOR2_X1 U22007 ( .A1(n12607), .A2(n23553), .Z(n46499) );
  NOR2_X2 U22011 ( .A1(n18023), .A2(n62451), .ZN(n56341) );
  NAND3_X2 U22013 ( .A1(n56242), .A2(n56244), .A3(n56237), .ZN(n62451) );
  NAND2_X2 U22014 ( .A1(n17452), .A2(n9770), .ZN(n17905) );
  AND2_X2 U22015 ( .A1(n42288), .A2(n42285), .Z(n12975) );
  NAND3_X1 U22018 ( .A1(n16443), .A2(n3766), .A3(n63131), .ZN(n35520) );
  NAND2_X2 U22019 ( .A1(n62452), .A2(n61944), .ZN(n63118) );
  NOR2_X2 U22021 ( .A1(n16652), .A2(n16653), .ZN(n62452) );
  NOR2_X2 U22022 ( .A1(n53160), .A2(n25484), .ZN(n52231) );
  NAND2_X2 U22024 ( .A1(n62480), .A2(n16453), .ZN(n4808) );
  NOR2_X2 U22025 ( .A1(n10381), .A2(n55642), .ZN(n55617) );
  NOR2_X2 U22034 ( .A1(n18209), .A2(n37247), .ZN(n60533) );
  NOR2_X2 U22040 ( .A1(n37943), .A2(n12050), .ZN(n37019) );
  NAND3_X2 U22045 ( .A1(n20040), .A2(n5718), .A3(n62456), .ZN(n26248) );
  NOR3_X2 U22046 ( .A1(n20037), .A2(n20039), .A3(n42073), .ZN(n62456) );
  XOR2_X1 U22051 ( .A1(n6294), .A2(n62457), .Z(n12127) );
  XOR2_X1 U22059 ( .A1(n6296), .A2(n15916), .Z(n62457) );
  INV_X1 U22060 ( .I(n63372), .ZN(n43916) );
  NAND4_X2 U22068 ( .A1(n57515), .A2(n14344), .A3(n57514), .A4(n41808), .ZN(
        n63372) );
  NOR3_X2 U22080 ( .A1(n61375), .A2(n50004), .A3(n64562), .ZN(n63244) );
  NAND2_X2 U22081 ( .A1(n60209), .A2(n50360), .ZN(n61375) );
  NAND3_X1 U22082 ( .A1(n28069), .A2(n28070), .A3(n28068), .ZN(n28075) );
  NOR2_X2 U22083 ( .A1(n17186), .A2(n62458), .ZN(n2130) );
  NAND3_X2 U22098 ( .A1(n28087), .A2(n58246), .A3(n28088), .ZN(n62458) );
  XOR2_X1 U22099 ( .A1(n62459), .A2(n53064), .Z(Plaintext[1]) );
  XOR2_X1 U22102 ( .A1(n38377), .A2(n7589), .Z(n9767) );
  NAND3_X2 U22103 ( .A1(n34807), .A2(n16682), .A3(n34808), .ZN(n38377) );
  NOR2_X2 U22104 ( .A1(n6551), .A2(n63391), .ZN(n6549) );
  AND2_X2 U22105 ( .A1(n9243), .A2(n63017), .Z(n9368) );
  NOR3_X2 U22106 ( .A1(n52826), .A2(n13422), .A3(n23507), .ZN(n13421) );
  NAND2_X1 U22108 ( .A1(n6881), .A2(n33826), .ZN(n62463) );
  AND2_X1 U22111 ( .A1(n28034), .A2(n9661), .Z(n27057) );
  XOR2_X1 U22112 ( .A1(n31454), .A2(n31452), .Z(n33042) );
  XOR2_X1 U22113 ( .A1(n59546), .A2(n11236), .Z(n31454) );
  XOR2_X1 U22115 ( .A1(n13233), .A2(n64775), .Z(n8854) );
  NAND2_X2 U22123 ( .A1(n8851), .A2(n53443), .ZN(n53439) );
  XOR2_X1 U22126 ( .A1(n30291), .A2(n2494), .Z(n12954) );
  OAI21_X1 U22127 ( .A1(n30185), .A2(n62587), .B(n62586), .ZN(n30188) );
  OAI21_X1 U22128 ( .A1(n47414), .A2(n47425), .B(n59528), .ZN(n23996) );
  XOR2_X1 U22132 ( .A1(n62465), .A2(n53714), .Z(Plaintext[36]) );
  NOR2_X1 U22135 ( .A1(n19110), .A2(n22017), .ZN(n62465) );
  NAND2_X2 U22144 ( .A1(n62621), .A2(n62466), .ZN(n14857) );
  NOR3_X2 U22146 ( .A1(n62467), .A2(n42366), .A3(n25806), .ZN(n42053) );
  AOI22_X2 U22147 ( .A1(n58353), .A2(n58352), .B1(n58031), .B2(n44560), .ZN(
        n44568) );
  XOR2_X1 U22159 ( .A1(n50194), .A2(n49898), .Z(n25257) );
  XOR2_X1 U22162 ( .A1(n8472), .A2(n63010), .Z(n50194) );
  NAND2_X2 U22163 ( .A1(n36716), .A2(n20867), .ZN(n36724) );
  AND2_X2 U22170 ( .A1(n60075), .A2(n10811), .Z(n4918) );
  NOR2_X1 U22178 ( .A1(n64731), .A2(n61767), .ZN(n63794) );
  XOR2_X1 U22184 ( .A1(n64995), .A2(n62468), .Z(n25333) );
  XOR2_X1 U22185 ( .A1(n58858), .A2(n1549), .Z(n62468) );
  NAND2_X2 U22188 ( .A1(n29794), .A2(n21222), .ZN(n9281) );
  NAND2_X2 U22190 ( .A1(n21223), .A2(n9014), .ZN(n21222) );
  BUF_X2 U22200 ( .I(n17589), .Z(n62469) );
  AND2_X1 U22203 ( .A1(n33573), .A2(n62470), .Z(n19791) );
  NOR2_X1 U22208 ( .A1(n40396), .A2(n41081), .ZN(n64925) );
  OAI22_X2 U22210 ( .A1(n36726), .A2(n58743), .B1(n36727), .B2(n36728), .ZN(
        n62471) );
  XOR2_X1 U22213 ( .A1(n62472), .A2(n31486), .Z(n31597) );
  XOR2_X1 U22214 ( .A1(n16439), .A2(n32230), .Z(n10583) );
  NAND3_X2 U22215 ( .A1(n36522), .A2(n37368), .A3(n62473), .ZN(n57764) );
  XOR2_X1 U22220 ( .A1(n64839), .A2(n45845), .Z(n9729) );
  XOR2_X1 U22221 ( .A1(n64266), .A2(n12265), .Z(n45845) );
  NAND2_X1 U22222 ( .A1(n63371), .A2(n20287), .ZN(n62640) );
  XOR2_X1 U22226 ( .A1(n26206), .A2(n11234), .Z(n60311) );
  XOR2_X1 U22227 ( .A1(n62607), .A2(n2457), .Z(n11234) );
  NAND2_X2 U22233 ( .A1(n61726), .A2(n55176), .ZN(n55214) );
  NAND2_X2 U22241 ( .A1(n6524), .A2(n703), .ZN(n11227) );
  NOR2_X2 U22243 ( .A1(n24596), .A2(n25445), .ZN(n6524) );
  OAI22_X2 U22247 ( .A1(n49020), .A2(n48323), .B1(n48031), .B2(n48030), .ZN(
        n65080) );
  XOR2_X1 U22258 ( .A1(n62476), .A2(n62475), .Z(n63705) );
  XOR2_X1 U22272 ( .A1(n10996), .A2(n21220), .Z(n62476) );
  INV_X2 U22278 ( .I(n27907), .ZN(n31174) );
  NAND2_X2 U22283 ( .A1(n62053), .A2(n31189), .ZN(n27907) );
  NOR2_X2 U22287 ( .A1(n33807), .A2(n35712), .ZN(n7710) );
  NAND2_X2 U22288 ( .A1(n4808), .A2(n53146), .ZN(n53160) );
  AND2_X1 U22289 ( .A1(n17170), .A2(n51469), .Z(n62480) );
  NAND3_X1 U22291 ( .A1(n61579), .A2(n36803), .A3(n10110), .ZN(n36068) );
  NAND2_X1 U22293 ( .A1(n14887), .A2(n27214), .ZN(n27215) );
  NAND2_X2 U22300 ( .A1(n3082), .A2(n34018), .ZN(n34558) );
  NAND3_X2 U22308 ( .A1(n61757), .A2(n62481), .A3(n63626), .ZN(n63405) );
  NOR2_X2 U22309 ( .A1(n62524), .A2(n62482), .ZN(n62481) );
  NAND3_X2 U22312 ( .A1(n22779), .A2(n49140), .A3(n49141), .ZN(n51940) );
  XOR2_X1 U22314 ( .A1(n16624), .A2(n62483), .Z(n64382) );
  XOR2_X1 U22315 ( .A1(n15297), .A2(n4256), .Z(n62483) );
  NAND3_X2 U22320 ( .A1(n48216), .A2(n62758), .A3(n48203), .ZN(n63619) );
  NOR2_X2 U22321 ( .A1(n15278), .A2(n15279), .ZN(n60486) );
  NOR2_X1 U22322 ( .A1(n63183), .A2(n63182), .ZN(n63181) );
  INV_X2 U22324 ( .I(n10939), .ZN(n46573) );
  OAI21_X2 U22326 ( .A1(n48152), .A2(n64779), .B(n48151), .ZN(n48156) );
  NAND2_X2 U22327 ( .A1(n60416), .A2(n59724), .ZN(n34764) );
  NAND2_X2 U22329 ( .A1(n34209), .A2(n21059), .ZN(n59724) );
  NAND2_X2 U22333 ( .A1(n46040), .A2(n46026), .ZN(n46859) );
  INV_X2 U22334 ( .I(n45725), .ZN(n46040) );
  NAND2_X2 U22340 ( .A1(n63501), .A2(n45718), .ZN(n45725) );
  NOR2_X2 U22342 ( .A1(n4328), .A2(n43271), .ZN(n4327) );
  NAND2_X2 U22347 ( .A1(n12244), .A2(n62485), .ZN(n13493) );
  AND3_X1 U22352 ( .A1(n39603), .A2(n39602), .A3(n40694), .Z(n62485) );
  INV_X2 U22357 ( .I(n38702), .ZN(n57757) );
  XOR2_X1 U22366 ( .A1(n23162), .A2(n44957), .Z(n58455) );
  AND2_X1 U22368 ( .A1(n61742), .A2(n18364), .Z(n48425) );
  NOR2_X2 U22370 ( .A1(n65259), .A2(n62486), .ZN(n37761) );
  NAND3_X2 U22376 ( .A1(n62917), .A2(n35585), .A3(n35584), .ZN(n62486) );
  NOR2_X1 U22380 ( .A1(n27866), .A2(n63252), .ZN(n24557) );
  BUF_X2 U22404 ( .I(n2583), .Z(n62487) );
  NAND2_X1 U22414 ( .A1(n200), .A2(n11391), .ZN(n62488) );
  BUF_X4 U22420 ( .I(n22657), .Z(n8343) );
  XOR2_X1 U22427 ( .A1(n22142), .A2(n1681), .Z(n11011) );
  XOR2_X1 U22431 ( .A1(n22143), .A2(n4111), .Z(n2217) );
  XOR2_X1 U22432 ( .A1(n2213), .A2(n11307), .Z(n64134) );
  XOR2_X1 U22433 ( .A1(n51939), .A2(n62489), .Z(n55691) );
  XOR2_X1 U22441 ( .A1(n52059), .A2(n52156), .Z(n62489) );
  NAND2_X2 U22445 ( .A1(n13258), .A2(n23407), .ZN(n57234) );
  INV_X1 U22449 ( .I(n39987), .ZN(n24982) );
  OR2_X1 U22450 ( .A1(n39987), .A2(n14994), .Z(n40756) );
  BUF_X2 U22451 ( .I(n5536), .Z(n59858) );
  XOR2_X1 U22458 ( .A1(n62491), .A2(n52358), .Z(n52362) );
  XOR2_X1 U22461 ( .A1(n9506), .A2(n52357), .Z(n62491) );
  NAND3_X2 U22464 ( .A1(n62492), .A2(n57717), .A3(n17477), .ZN(n24294) );
  NAND2_X1 U22465 ( .A1(n41057), .A2(n41056), .ZN(n62492) );
  NOR3_X2 U22466 ( .A1(n19641), .A2(n62493), .A3(n36237), .ZN(n60492) );
  NOR2_X2 U22473 ( .A1(n7831), .A2(n10317), .ZN(n62493) );
  NOR3_X2 U22474 ( .A1(n14210), .A2(n14206), .A3(n62494), .ZN(n25394) );
  NAND4_X2 U22479 ( .A1(n14203), .A2(n11615), .A3(n49516), .A4(n49522), .ZN(
        n62494) );
  XOR2_X1 U22485 ( .A1(n15844), .A2(n11797), .Z(n64217) );
  XOR2_X1 U22486 ( .A1(n11742), .A2(n52447), .Z(n60992) );
  NAND2_X2 U22487 ( .A1(n49469), .A2(n49470), .ZN(n52447) );
  BUF_X2 U22492 ( .I(n30343), .Z(n62495) );
  AOI21_X2 U22493 ( .A1(n20311), .A2(n63943), .B(n50043), .ZN(n49574) );
  XOR2_X1 U22499 ( .A1(n1390), .A2(n5676), .Z(n10538) );
  NAND2_X1 U22506 ( .A1(n34531), .A2(n8431), .ZN(n34533) );
  NAND2_X2 U22510 ( .A1(n33729), .A2(n34961), .ZN(n8431) );
  XOR2_X1 U22511 ( .A1(n17657), .A2(n26206), .Z(n17766) );
  XOR2_X1 U22515 ( .A1(n63538), .A2(n38220), .Z(n17657) );
  NAND2_X2 U22518 ( .A1(n50220), .A2(n7824), .ZN(n50211) );
  INV_X2 U22519 ( .I(n62497), .ZN(n24682) );
  XNOR2_X1 U22522 ( .A1(n2404), .A2(n46610), .ZN(n62497) );
  NOR3_X1 U22527 ( .A1(n62498), .A2(n55230), .A3(n61768), .ZN(n55221) );
  NAND3_X1 U22528 ( .A1(n55215), .A2(n55214), .A3(n55212), .ZN(n62498) );
  NAND2_X1 U22533 ( .A1(n63856), .A2(n59001), .ZN(n12271) );
  XOR2_X1 U22535 ( .A1(n52346), .A2(n52345), .Z(n58320) );
  NOR2_X2 U22539 ( .A1(n52963), .A2(n59256), .ZN(n16978) );
  XOR2_X1 U22543 ( .A1(n12269), .A2(n8673), .Z(n16242) );
  XOR2_X1 U22544 ( .A1(n60701), .A2(n45093), .Z(n12269) );
  NAND3_X2 U22546 ( .A1(n58453), .A2(n47365), .A3(n9454), .ZN(n61181) );
  NAND2_X2 U22547 ( .A1(n8880), .A2(n33296), .ZN(n15012) );
  OR2_X2 U22548 ( .A1(n592), .A2(n6682), .Z(n11077) );
  NAND2_X1 U22551 ( .A1(n20762), .A2(n28756), .ZN(n63453) );
  OAI22_X1 U22555 ( .A1(n40551), .A2(n42665), .B1(n42849), .B2(n42139), .ZN(
        n42850) );
  INV_X2 U22556 ( .I(n10939), .ZN(n60906) );
  NAND2_X2 U22560 ( .A1(n14428), .A2(n15245), .ZN(n55345) );
  XOR2_X1 U22561 ( .A1(n60118), .A2(n20573), .Z(n2978) );
  NAND2_X2 U22564 ( .A1(n62499), .A2(n467), .ZN(n3464) );
  NAND3_X2 U22569 ( .A1(n48108), .A2(n22464), .A3(n23331), .ZN(n19558) );
  INV_X2 U22571 ( .I(n3149), .ZN(n35985) );
  INV_X4 U22572 ( .I(n25788), .ZN(n15720) );
  OAI22_X1 U22576 ( .A1(n33990), .A2(n33989), .B1(n33991), .B2(n33992), .ZN(
        n33996) );
  XOR2_X1 U22582 ( .A1(n25828), .A2(n51691), .Z(n7885) );
  NOR2_X2 U22588 ( .A1(n57780), .A2(n59828), .ZN(n25828) );
  NOR2_X2 U22597 ( .A1(n20311), .A2(n49581), .ZN(n14171) );
  XOR2_X1 U22600 ( .A1(n19606), .A2(n25690), .Z(n21331) );
  NOR2_X2 U22603 ( .A1(n9580), .A2(n9579), .ZN(n19606) );
  OAI21_X1 U22604 ( .A1(n2697), .A2(n49047), .B(n49046), .ZN(n49052) );
  OR2_X1 U22605 ( .A1(n53427), .A2(n53625), .Z(n53418) );
  XOR2_X1 U22610 ( .A1(n5919), .A2(n38889), .Z(n38931) );
  XOR2_X1 U22617 ( .A1(n44317), .A2(n60511), .Z(n44531) );
  OR2_X1 U22621 ( .A1(n10717), .A2(n9536), .Z(n34009) );
  NOR2_X2 U22634 ( .A1(n18599), .A2(n26208), .ZN(n63261) );
  XNOR2_X1 U22637 ( .A1(n44734), .A2(n16700), .ZN(n62688) );
  XOR2_X1 U22643 ( .A1(n44757), .A2(n61573), .Z(n17815) );
  NOR3_X2 U22644 ( .A1(n6545), .A2(n6547), .A3(n6546), .ZN(n6548) );
  OR2_X1 U22645 ( .A1(n26648), .A2(n26647), .Z(n17415) );
  NAND3_X2 U22646 ( .A1(n12147), .A2(n12145), .A3(n63283), .ZN(n22573) );
  XOR2_X1 U22653 ( .A1(n6003), .A2(n64718), .Z(n4560) );
  NAND2_X2 U22661 ( .A1(n26671), .A2(n27611), .ZN(n27614) );
  XOR2_X1 U22662 ( .A1(n51080), .A2(n62503), .Z(n51084) );
  XOR2_X1 U22664 ( .A1(n51078), .A2(n51077), .Z(n62503) );
  INV_X2 U22665 ( .I(n13458), .ZN(n63030) );
  NOR2_X1 U22666 ( .A1(n62504), .A2(n56761), .ZN(n58431) );
  NAND4_X1 U22670 ( .A1(n56751), .A2(n56753), .A3(n56754), .A4(n56752), .ZN(
        n62504) );
  OR2_X1 U22672 ( .A1(n41743), .A2(n58678), .Z(n58965) );
  XOR2_X1 U22674 ( .A1(n10662), .A2(n5101), .Z(n3290) );
  XOR2_X1 U22675 ( .A1(n7034), .A2(n9025), .Z(n10662) );
  OR2_X1 U22676 ( .A1(n13460), .A2(n22853), .Z(n8150) );
  AND2_X2 U22677 ( .A1(n20438), .A2(n60851), .Z(n62756) );
  XNOR2_X1 U22680 ( .A1(n45269), .A2(n59849), .ZN(n45282) );
  NOR2_X2 U22684 ( .A1(n29516), .A2(n29523), .ZN(n29520) );
  INV_X2 U22685 ( .I(n49172), .ZN(n62505) );
  AND2_X1 U22689 ( .A1(n12539), .A2(n64603), .Z(n34081) );
  XOR2_X1 U22692 ( .A1(n18709), .A2(n17919), .Z(n2897) );
  XOR2_X1 U22697 ( .A1(n23587), .A2(n20754), .Z(n18709) );
  NOR2_X2 U22700 ( .A1(n5612), .A2(n62508), .ZN(n5611) );
  OAI21_X2 U22701 ( .A1(n2332), .A2(n3790), .B(n2331), .ZN(n62508) );
  NOR2_X2 U22707 ( .A1(n62511), .A2(n1348), .ZN(n2144) );
  NAND2_X2 U22708 ( .A1(n2843), .A2(n61903), .ZN(n62511) );
  NOR2_X2 U22715 ( .A1(n62512), .A2(n61908), .ZN(n31472) );
  NOR2_X2 U22720 ( .A1(n62582), .A2(n1535), .ZN(n62512) );
  INV_X2 U22722 ( .I(n37027), .ZN(n35911) );
  NAND2_X2 U22729 ( .A1(n2699), .A2(n22524), .ZN(n37027) );
  NAND3_X2 U22730 ( .A1(n64589), .A2(n29014), .A3(n29798), .ZN(n30074) );
  XOR2_X1 U22733 ( .A1(n15840), .A2(n8590), .Z(n32107) );
  OAI22_X2 U22734 ( .A1(n40691), .A2(n39845), .B1(n7848), .B2(n40380), .ZN(
        n40382) );
  NAND2_X2 U22737 ( .A1(n25976), .A2(n41433), .ZN(n40380) );
  NAND3_X1 U22738 ( .A1(n53785), .A2(n53786), .A3(n53784), .ZN(n64807) );
  OAI22_X1 U22739 ( .A1(n62513), .A2(n53428), .B1(n1259), .B2(n61147), .ZN(
        n4222) );
  INV_X2 U22748 ( .I(n19589), .ZN(n47356) );
  NAND3_X2 U22749 ( .A1(n19897), .A2(n48061), .A3(n19896), .ZN(n19976) );
  NAND2_X2 U22750 ( .A1(n62517), .A2(n62516), .ZN(n13800) );
  INV_X2 U22751 ( .I(n57001), .ZN(n62517) );
  XOR2_X1 U22752 ( .A1(n38367), .A2(n39315), .Z(n12253) );
  NOR3_X2 U22753 ( .A1(n49195), .A2(n61673), .A3(n62606), .ZN(n13317) );
  XOR2_X1 U22754 ( .A1(n62519), .A2(n13219), .Z(n11256) );
  XOR2_X1 U22760 ( .A1(n65227), .A2(n3244), .Z(n62519) );
  NAND2_X2 U22763 ( .A1(n19681), .A2(n45547), .ZN(n48823) );
  NOR2_X2 U22765 ( .A1(n64712), .A2(n22114), .ZN(n21561) );
  XOR2_X1 U22766 ( .A1(n62520), .A2(n7699), .Z(n7136) );
  XOR2_X1 U22768 ( .A1(n46178), .A2(n5969), .Z(n62520) );
  XOR2_X1 U22773 ( .A1(n59931), .A2(n51700), .Z(n15262) );
  INV_X2 U22776 ( .I(n5971), .ZN(n62997) );
  XOR2_X1 U22777 ( .A1(n62521), .A2(n9269), .Z(n38206) );
  XOR2_X1 U22785 ( .A1(n6092), .A2(n38142), .Z(n62521) );
  XOR2_X1 U22789 ( .A1(n51828), .A2(n17172), .Z(n25099) );
  NAND3_X2 U22800 ( .A1(n62523), .A2(n45914), .A3(n62522), .ZN(n24797) );
  INV_X2 U22803 ( .I(n41287), .ZN(n43890) );
  NAND3_X2 U22804 ( .A1(n41285), .A2(n987), .A3(n41286), .ZN(n41287) );
  XOR2_X1 U22810 ( .A1(n17171), .A2(n52192), .Z(n52193) );
  OAI21_X1 U22818 ( .A1(n61769), .A2(n64637), .B(n7894), .ZN(n7893) );
  INV_X2 U22819 ( .I(n62525), .ZN(n41859) );
  NOR2_X2 U22822 ( .A1(n41856), .A2(n22882), .ZN(n62525) );
  XOR2_X1 U22823 ( .A1(n52510), .A2(n62526), .Z(n54793) );
  XOR2_X1 U22827 ( .A1(n62527), .A2(n52524), .Z(n62526) );
  XOR2_X1 U22829 ( .A1(n4751), .A2(n57490), .Z(n10053) );
  XOR2_X1 U22833 ( .A1(n12092), .A2(n12095), .Z(n18774) );
  INV_X2 U22834 ( .I(n18489), .ZN(n35794) );
  NAND2_X2 U22835 ( .A1(n18488), .A2(n18489), .ZN(n34386) );
  NOR2_X2 U22845 ( .A1(n5604), .A2(n2989), .ZN(n18489) );
  NOR2_X1 U22846 ( .A1(n62528), .A2(n29038), .ZN(n7546) );
  NAND2_X1 U22847 ( .A1(n7548), .A2(n60339), .ZN(n62528) );
  OR2_X1 U22850 ( .A1(n63163), .A2(n10526), .Z(n20706) );
  XOR2_X1 U22853 ( .A1(n63879), .A2(n4209), .Z(n14999) );
  XOR2_X1 U22855 ( .A1(n13246), .A2(n13245), .Z(n4209) );
  NAND2_X2 U22861 ( .A1(n7204), .A2(n63703), .ZN(n62530) );
  NAND2_X2 U22862 ( .A1(n25987), .A2(n56957), .ZN(n56963) );
  NAND2_X2 U22863 ( .A1(n56880), .A2(n56867), .ZN(n2372) );
  XOR2_X1 U22872 ( .A1(n13643), .A2(n13640), .Z(n53233) );
  XOR2_X1 U22876 ( .A1(n14731), .A2(n25394), .Z(n1189) );
  NOR3_X2 U22877 ( .A1(n52288), .A2(n9655), .A3(n14708), .ZN(n56902) );
  NAND2_X2 U22883 ( .A1(n138), .A2(n1257), .ZN(n52288) );
  OAI22_X1 U22886 ( .A1(n63714), .A2(n29118), .B1(n3087), .B2(n8613), .ZN(
        n62532) );
  XOR2_X1 U22888 ( .A1(n7199), .A2(n32663), .Z(n25935) );
  NOR2_X2 U22889 ( .A1(n62746), .A2(n29756), .ZN(n7199) );
  XOR2_X1 U22892 ( .A1(n62533), .A2(n1818), .Z(n13214) );
  XOR2_X1 U22894 ( .A1(n63306), .A2(n32405), .Z(n62533) );
  NAND2_X2 U22900 ( .A1(n21678), .A2(n18691), .ZN(n21588) );
  NOR2_X2 U22901 ( .A1(n3086), .A2(n23901), .ZN(n18691) );
  XOR2_X1 U22903 ( .A1(n31599), .A2(n5726), .Z(n3389) );
  NAND2_X2 U22906 ( .A1(n62556), .A2(n3390), .ZN(n31599) );
  INV_X2 U22907 ( .I(n54015), .ZN(n51864) );
  NAND2_X2 U22910 ( .A1(n54017), .A2(n53036), .ZN(n54015) );
  NAND4_X2 U22915 ( .A1(n48526), .A2(n588), .A3(n48524), .A4(n62534), .ZN(
        n48527) );
  AOI22_X2 U22916 ( .A1(n48510), .A2(n21641), .B1(n63135), .B2(n48508), .ZN(
        n62534) );
  XOR2_X1 U22920 ( .A1(n38321), .A2(n50878), .Z(n37824) );
  XOR2_X1 U22921 ( .A1(n19184), .A2(n39579), .Z(n38321) );
  NAND3_X1 U22926 ( .A1(n17991), .A2(n17992), .A3(n27321), .ZN(n59333) );
  NOR2_X1 U22933 ( .A1(n42622), .A2(n42620), .ZN(n62536) );
  XOR2_X1 U22936 ( .A1(n62722), .A2(n64692), .Z(n24415) );
  NOR3_X1 U22938 ( .A1(n57839), .A2(n57234), .A3(n9986), .ZN(n44562) );
  NAND3_X2 U22947 ( .A1(n53011), .A2(n53012), .A3(n53013), .ZN(n53014) );
  NAND4_X1 U22949 ( .A1(n49905), .A2(n14315), .A3(n14314), .A4(n47787), .ZN(
        n5600) );
  NAND3_X2 U22953 ( .A1(n5189), .A2(n64207), .A3(n5187), .ZN(n23552) );
  OR3_X1 U22956 ( .A1(n40424), .A2(n40421), .A3(n61417), .Z(n39823) );
  NOR2_X2 U22959 ( .A1(n8324), .A2(n8323), .ZN(n45373) );
  NAND3_X2 U22966 ( .A1(n8317), .A2(n41668), .A3(n41669), .ZN(n8324) );
  NAND2_X2 U22967 ( .A1(n50338), .A2(n60467), .ZN(n21476) );
  NOR2_X2 U22969 ( .A1(n57995), .A2(n21052), .ZN(n50338) );
  NAND2_X2 U22975 ( .A1(n6205), .A2(n6206), .ZN(n2899) );
  NAND2_X2 U22979 ( .A1(n6001), .A2(n35748), .ZN(n6205) );
  NAND2_X1 U22985 ( .A1(n21982), .A2(n18487), .ZN(n53177) );
  NAND2_X2 U22986 ( .A1(n61165), .A2(n22935), .ZN(n37313) );
  OAI22_X1 U23005 ( .A1(n50818), .A2(n53717), .B1(n53706), .B2(n53751), .ZN(
        n62539) );
  XOR2_X1 U23007 ( .A1(n6596), .A2(n62540), .Z(n10579) );
  XOR2_X1 U23009 ( .A1(n22747), .A2(n50167), .Z(n62540) );
  NAND3_X1 U23013 ( .A1(n63864), .A2(n49037), .A3(n12625), .ZN(n62553) );
  INV_X1 U23015 ( .I(n65089), .ZN(n24644) );
  OR2_X1 U23020 ( .A1(n65089), .A2(n62689), .Z(n10669) );
  NAND3_X2 U23021 ( .A1(n21822), .A2(n59545), .A3(n18607), .ZN(n50293) );
  NAND2_X2 U23022 ( .A1(n48559), .A2(n47121), .ZN(n47128) );
  NOR2_X2 U23024 ( .A1(n62541), .A2(n12803), .ZN(n25233) );
  XOR2_X1 U23030 ( .A1(n6780), .A2(n24468), .Z(n39439) );
  OAI22_X2 U23037 ( .A1(n62966), .A2(n61061), .B1(n1521), .B2(n6781), .ZN(
        n6780) );
  XNOR2_X1 U23042 ( .A1(n32057), .A2(n31322), .ZN(n30715) );
  AOI21_X2 U23053 ( .A1(n29752), .A2(n29753), .B(n29751), .ZN(n31322) );
  XOR2_X1 U23055 ( .A1(n62542), .A2(n18890), .Z(n18889) );
  XOR2_X1 U23069 ( .A1(n46206), .A2(n61445), .Z(n62542) );
  INV_X2 U23073 ( .I(n30658), .ZN(n30416) );
  NAND2_X2 U23074 ( .A1(n63537), .A2(n28711), .ZN(n30658) );
  XOR2_X1 U23075 ( .A1(n6216), .A2(n21686), .Z(n21685) );
  NOR3_X2 U23076 ( .A1(n37217), .A2(n37216), .A3(n29), .ZN(n22404) );
  NOR2_X2 U23079 ( .A1(n41443), .A2(n41442), .ZN(n62543) );
  OR2_X1 U23080 ( .A1(n1341), .A2(n25563), .Z(n35669) );
  NOR2_X2 U23085 ( .A1(n41483), .A2(n43318), .ZN(n42770) );
  INV_X2 U23090 ( .I(n62544), .ZN(n57187) );
  XNOR2_X1 U23097 ( .A1(n44893), .A2(n22396), .ZN(n62544) );
  NOR2_X2 U23099 ( .A1(n25988), .A2(n18582), .ZN(n20477) );
  INV_X2 U23104 ( .I(n56935), .ZN(n25988) );
  NAND3_X2 U23114 ( .A1(n52261), .A2(n52259), .A3(n64119), .ZN(n56935) );
  XOR2_X1 U23117 ( .A1(n1684), .A2(n23587), .Z(n4521) );
  XOR2_X1 U23120 ( .A1(n62545), .A2(n17061), .Z(n3887) );
  XOR2_X1 U23121 ( .A1(n31336), .A2(n21986), .Z(n33866) );
  NAND2_X2 U23138 ( .A1(n17545), .A2(n17544), .ZN(n31336) );
  NAND4_X2 U23139 ( .A1(n16574), .A2(n16573), .A3(n55646), .A4(n55653), .ZN(
        n62557) );
  NAND3_X2 U23142 ( .A1(n61880), .A2(n63739), .A3(n15232), .ZN(n44478) );
  INV_X2 U23146 ( .I(n25323), .ZN(n41120) );
  XOR2_X1 U23147 ( .A1(n58014), .A2(n58013), .Z(n25323) );
  AND2_X1 U23148 ( .A1(n41985), .A2(n41986), .Z(n58434) );
  NAND3_X2 U23149 ( .A1(n5369), .A2(n1694), .A3(n41980), .ZN(n41986) );
  NAND2_X1 U23150 ( .A1(n23054), .A2(n18715), .ZN(n63178) );
  NAND3_X2 U23161 ( .A1(n56248), .A2(n16160), .A3(n20737), .ZN(n56596) );
  BUF_X4 U23162 ( .I(n8287), .Z(n2754) );
  INV_X2 U23164 ( .I(n62547), .ZN(n25068) );
  NAND3_X2 U23165 ( .A1(n25074), .A2(n25073), .A3(n38034), .ZN(n62547) );
  NAND3_X1 U23169 ( .A1(n45367), .A2(n23099), .A3(n2955), .ZN(n63709) );
  NAND4_X1 U23171 ( .A1(n52488), .A2(n55006), .A3(n55440), .A4(n55438), .ZN(
        n52118) );
  XOR2_X1 U23174 ( .A1(n32011), .A2(n62548), .Z(n31200) );
  NAND2_X1 U23176 ( .A1(n63769), .A2(n64223), .ZN(n18019) );
  XOR2_X1 U23177 ( .A1(n57187), .A2(n10139), .Z(n5273) );
  NAND4_X1 U23178 ( .A1(n19031), .A2(n19035), .A3(n55839), .A4(n55838), .ZN(
        n65136) );
  NAND4_X2 U23179 ( .A1(n58720), .A2(n58721), .A3(n52314), .A4(n52315), .ZN(
        n65130) );
  XOR2_X1 U23185 ( .A1(n11261), .A2(n18156), .Z(n15589) );
  XOR2_X1 U23187 ( .A1(n4057), .A2(n4056), .Z(n11261) );
  NAND2_X2 U23190 ( .A1(n62551), .A2(n52389), .ZN(n57993) );
  NAND3_X2 U23191 ( .A1(n55480), .A2(n52210), .A3(n22588), .ZN(n62551) );
  NAND2_X2 U23197 ( .A1(n14964), .A2(n19190), .ZN(n63337) );
  NAND2_X1 U23198 ( .A1(n4437), .A2(n15280), .ZN(n57410) );
  OAI21_X1 U23199 ( .A1(n30169), .A2(n30170), .B(n30168), .ZN(n62552) );
  NOR2_X2 U23202 ( .A1(n61107), .A2(n15784), .ZN(n41584) );
  OR2_X2 U23205 ( .A1(n38697), .A2(n38696), .Z(n15784) );
  NAND3_X1 U23206 ( .A1(n58388), .A2(n10821), .A3(n30804), .ZN(n28753) );
  NAND2_X2 U23208 ( .A1(n8521), .A2(n10820), .ZN(n58388) );
  NAND2_X1 U23209 ( .A1(n42805), .A2(n42802), .ZN(n64378) );
  NAND2_X1 U23212 ( .A1(n62555), .A2(n62554), .ZN(n52313) );
  NAND2_X1 U23213 ( .A1(n52310), .A2(n55631), .ZN(n62554) );
  NAND2_X1 U23215 ( .A1(n52311), .A2(n19021), .ZN(n62555) );
  NAND3_X1 U23222 ( .A1(n55742), .A2(n55744), .A3(n62558), .ZN(n64409) );
  XOR2_X1 U23223 ( .A1(n64269), .A2(n31290), .Z(n63860) );
  INV_X2 U23225 ( .I(n20059), .ZN(n64269) );
  XOR2_X1 U23226 ( .A1(n60743), .A2(n9288), .Z(n20059) );
  NOR2_X2 U23228 ( .A1(n9514), .A2(n53625), .ZN(n52781) );
  INV_X2 U23233 ( .I(n13489), .ZN(n17635) );
  NAND2_X2 U23242 ( .A1(n2408), .A2(n56540), .ZN(n13489) );
  NAND2_X2 U23250 ( .A1(n59271), .A2(n41900), .ZN(n41895) );
  NOR2_X2 U23251 ( .A1(n25874), .A2(n23145), .ZN(n41900) );
  XOR2_X1 U23255 ( .A1(n62557), .A2(n55655), .Z(Plaintext[125]) );
  NOR2_X2 U23257 ( .A1(n8259), .A2(n55644), .ZN(n55640) );
  NAND2_X1 U23259 ( .A1(n65203), .A2(n62535), .ZN(n43417) );
  NAND2_X2 U23261 ( .A1(n58475), .A2(n62559), .ZN(n59845) );
  AND2_X1 U23262 ( .A1(n60399), .A2(n24706), .Z(n62559) );
  XOR2_X1 U23264 ( .A1(n62560), .A2(n9709), .Z(n10719) );
  XOR2_X1 U23265 ( .A1(n10721), .A2(n15476), .Z(n62560) );
  XOR2_X1 U23266 ( .A1(n2960), .A2(n46343), .Z(n256) );
  NAND2_X2 U23270 ( .A1(n22653), .A2(n64367), .ZN(n21471) );
  INV_X2 U23272 ( .I(n6305), .ZN(n60021) );
  NAND2_X2 U23278 ( .A1(n20339), .A2(n41950), .ZN(n6305) );
  NAND2_X1 U23279 ( .A1(n55297), .A2(n55684), .ZN(n24745) );
  XOR2_X1 U23281 ( .A1(n62562), .A2(n3208), .Z(n46611) );
  NOR2_X2 U23284 ( .A1(n60009), .A2(n18075), .ZN(n30521) );
  XOR2_X1 U23285 ( .A1(n39249), .A2(n39247), .Z(n5098) );
  NAND3_X2 U23286 ( .A1(n62563), .A2(n7004), .A3(n7001), .ZN(n9084) );
  NOR2_X2 U23287 ( .A1(n62564), .A2(n3921), .ZN(n3920) );
  OAI21_X2 U23294 ( .A1(n3923), .A2(n49048), .B(n48068), .ZN(n62564) );
  NAND2_X2 U23295 ( .A1(n52932), .A2(n55463), .ZN(n55734) );
  NAND2_X2 U23300 ( .A1(n61934), .A2(n63342), .ZN(n35211) );
  AOI22_X1 U23310 ( .A1(n27412), .A2(n26732), .B1(n28212), .B2(n29125), .ZN(
        n60301) );
  XOR2_X1 U23317 ( .A1(n62568), .A2(n52294), .Z(Plaintext[181]) );
  BUF_X2 U23318 ( .I(n5712), .Z(n62569) );
  BUF_X2 U23319 ( .I(n46033), .Z(n62571) );
  NOR2_X2 U23320 ( .A1(n21087), .A2(n3473), .ZN(n29128) );
  XOR2_X1 U23321 ( .A1(n4894), .A2(n51404), .Z(n51405) );
  XOR2_X1 U23323 ( .A1(n2694), .A2(n12800), .Z(n4894) );
  NAND4_X2 U23324 ( .A1(n53804), .A2(n53801), .A3(n53803), .A4(n53802), .ZN(
        n63969) );
  XOR2_X1 U23329 ( .A1(n62572), .A2(n25307), .Z(n21939) );
  XOR2_X1 U23331 ( .A1(n22661), .A2(n21937), .Z(n62572) );
  XOR2_X1 U23338 ( .A1(n62573), .A2(n20406), .Z(n60381) );
  XOR2_X1 U23339 ( .A1(n38718), .A2(n63201), .Z(n62573) );
  XOR2_X1 U23346 ( .A1(n46529), .A2(n46166), .Z(n14427) );
  NAND3_X2 U23353 ( .A1(n22767), .A2(n7530), .A3(n43369), .ZN(n46529) );
  NOR3_X2 U23354 ( .A1(n932), .A2(n62576), .A3(n62575), .ZN(n2717) );
  XOR2_X1 U23360 ( .A1(n19501), .A2(n19503), .Z(n19419) );
  NAND2_X2 U23363 ( .A1(n2995), .A2(n43572), .ZN(n42717) );
  XOR2_X1 U23364 ( .A1(n26023), .A2(n33053), .Z(n64949) );
  NAND2_X2 U23366 ( .A1(n35212), .A2(n18878), .ZN(n63342) );
  AND3_X1 U23367 ( .A1(n30227), .A2(n30228), .A3(n8458), .Z(n822) );
  INV_X2 U23369 ( .I(n63473), .ZN(n62578) );
  INV_X2 U23370 ( .I(n54727), .ZN(n62579) );
  XOR2_X1 U23375 ( .A1(n5224), .A2(n5222), .Z(n65213) );
  NAND2_X2 U23376 ( .A1(n35650), .A2(n19316), .ZN(n35250) );
  NOR2_X2 U23378 ( .A1(n40193), .A2(n1238), .ZN(n62580) );
  XOR2_X1 U23381 ( .A1(n37681), .A2(n14738), .Z(n25643) );
  NAND2_X2 U23382 ( .A1(n63575), .A2(n61122), .ZN(n14738) );
  XOR2_X1 U23384 ( .A1(n52505), .A2(n51621), .Z(n62798) );
  INV_X2 U23385 ( .I(n24714), .ZN(n52505) );
  XOR2_X1 U23386 ( .A1(n23582), .A2(n52581), .Z(n24714) );
  NOR3_X2 U23387 ( .A1(n13563), .A2(n63069), .A3(n62581), .ZN(n19363) );
  NAND4_X2 U23388 ( .A1(n13561), .A2(n13562), .A3(n15025), .A4(n12085), .ZN(
        n62581) );
  XOR2_X1 U23389 ( .A1(n4178), .A2(n6098), .Z(n60935) );
  XOR2_X1 U23396 ( .A1(n43878), .A2(n22108), .Z(n2821) );
  NOR2_X2 U23399 ( .A1(n42337), .A2(n63442), .ZN(n43878) );
  NOR2_X2 U23400 ( .A1(n45764), .A2(n62366), .ZN(n46910) );
  NAND2_X2 U23403 ( .A1(n6082), .A2(n6617), .ZN(n62978) );
  NAND2_X2 U23405 ( .A1(n54651), .A2(n51633), .ZN(n62768) );
  NAND2_X2 U23409 ( .A1(n14107), .A2(n62583), .ZN(n62582) );
  NAND2_X2 U23411 ( .A1(n53383), .A2(n52756), .ZN(n50676) );
  XOR2_X1 U23414 ( .A1(n46578), .A2(n4080), .Z(n4079) );
  XOR2_X1 U23419 ( .A1(n1051), .A2(n84), .Z(n46578) );
  NAND3_X1 U23421 ( .A1(n45722), .A2(n45721), .A3(n20426), .ZN(n45728) );
  XOR2_X1 U23428 ( .A1(n4549), .A2(n6848), .Z(n6845) );
  INV_X2 U23430 ( .I(n56880), .ZN(n56840) );
  NAND2_X2 U23435 ( .A1(n35675), .A2(n6915), .ZN(n62772) );
  NOR2_X2 U23439 ( .A1(n27826), .A2(n62584), .ZN(n13443) );
  OR2_X1 U23447 ( .A1(n27825), .A2(n27824), .Z(n62584) );
  NAND2_X2 U23448 ( .A1(n7812), .A2(n28769), .ZN(n31439) );
  NOR2_X2 U23451 ( .A1(n7813), .A2(n28768), .ZN(n7812) );
  XOR2_X1 U23452 ( .A1(n24471), .A2(n13045), .Z(n31431) );
  BUF_X2 U23453 ( .I(n30192), .Z(n62585) );
  NAND3_X2 U23454 ( .A1(n24618), .A2(n22969), .A3(n15996), .ZN(n57146) );
  XOR2_X1 U23455 ( .A1(n7658), .A2(n32162), .Z(n7657) );
  INV_X2 U23462 ( .I(n22796), .ZN(n62588) );
  NAND2_X2 U23470 ( .A1(n10636), .A2(n61728), .ZN(n63712) );
  XOR2_X1 U23471 ( .A1(n14597), .A2(n15372), .Z(n14596) );
  BUF_X2 U23472 ( .I(n52617), .Z(n62589) );
  XOR2_X1 U23474 ( .A1(n51511), .A2(n52165), .Z(n62590) );
  XOR2_X1 U23481 ( .A1(n46521), .A2(n43261), .Z(n14752) );
  INV_X2 U23482 ( .I(n46885), .ZN(n46900) );
  XOR2_X1 U23484 ( .A1(n49126), .A2(n51941), .Z(n60832) );
  XOR2_X1 U23489 ( .A1(n11288), .A2(n50949), .Z(n49126) );
  NAND2_X1 U23491 ( .A1(n4491), .A2(n26583), .ZN(n58829) );
  NOR3_X2 U23492 ( .A1(n60523), .A2(n26576), .A3(n26575), .ZN(n4491) );
  OAI21_X2 U23495 ( .A1(n61886), .A2(n26570), .B(n26569), .ZN(n4361) );
  NAND2_X2 U23497 ( .A1(n62591), .A2(n44677), .ZN(n44793) );
  NOR2_X2 U23498 ( .A1(n19258), .A2(n44675), .ZN(n62591) );
  BUF_X2 U23501 ( .I(n64764), .Z(n62593) );
  BUF_X2 U23502 ( .I(n863), .Z(n9331) );
  XOR2_X1 U23505 ( .A1(n62594), .A2(n22521), .Z(n51386) );
  XOR2_X1 U23511 ( .A1(n22478), .A2(n51384), .Z(n62594) );
  NOR2_X1 U23512 ( .A1(n12479), .A2(n22185), .ZN(n57332) );
  XOR2_X1 U23514 ( .A1(n62595), .A2(n55191), .Z(Plaintext[103]) );
  NAND4_X2 U23515 ( .A1(n55190), .A2(n55189), .A3(n63711), .A4(n55187), .ZN(
        n62595) );
  BUF_X4 U23518 ( .I(n56540), .Z(n22870) );
  INV_X2 U23519 ( .I(n39117), .ZN(n41016) );
  NOR2_X2 U23521 ( .A1(n40500), .A2(n57199), .ZN(n39117) );
  AOI21_X1 U23525 ( .A1(n49847), .A2(n48983), .B(n6340), .ZN(n48986) );
  NOR2_X2 U23526 ( .A1(n58205), .A2(n49843), .ZN(n49847) );
  NAND2_X2 U23531 ( .A1(n63379), .A2(n60384), .ZN(n23863) );
  NAND4_X1 U23532 ( .A1(n60811), .A2(n56749), .A3(n56773), .A4(n62596), .ZN(
        n56753) );
  INV_X2 U23534 ( .I(n60833), .ZN(n53580) );
  NAND2_X2 U23537 ( .A1(n60002), .A2(n26089), .ZN(n60833) );
  NOR2_X2 U23538 ( .A1(n37334), .A2(n37339), .ZN(n63348) );
  INV_X1 U23539 ( .I(n62775), .ZN(n32438) );
  OR2_X1 U23540 ( .A1(n62775), .A2(n19005), .Z(n31906) );
  NAND2_X2 U23541 ( .A1(n62723), .A2(n62599), .ZN(n22343) );
  XOR2_X1 U23549 ( .A1(n52155), .A2(n2801), .Z(n2185) );
  NAND3_X1 U23551 ( .A1(n58205), .A2(n2433), .A3(n58269), .ZN(n48380) );
  BUF_X2 U23566 ( .I(n64946), .Z(n62600) );
  NAND2_X2 U23567 ( .A1(n60297), .A2(n22317), .ZN(n36588) );
  XOR2_X1 U23569 ( .A1(n4894), .A2(n52465), .Z(n51749) );
  NOR2_X1 U23572 ( .A1(n58880), .A2(n49045), .ZN(n58390) );
  NAND2_X1 U23574 ( .A1(n19274), .A2(n62601), .ZN(n63965) );
  NAND3_X1 U23576 ( .A1(n40432), .A2(n61984), .A3(n64183), .ZN(n62601) );
  INV_X1 U23578 ( .I(n52751), .ZN(n12440) );
  NAND3_X2 U23580 ( .A1(n59724), .A2(n60970), .A3(n34761), .ZN(n32941) );
  NOR2_X1 U23582 ( .A1(n61244), .A2(n13814), .ZN(n7889) );
  NAND3_X2 U23583 ( .A1(n57186), .A2(n55205), .A3(n55219), .ZN(n62602) );
  NAND2_X2 U23585 ( .A1(n40697), .A2(n22832), .ZN(n11855) );
  XOR2_X1 U23586 ( .A1(n62603), .A2(n64412), .Z(n39317) );
  INV_X4 U23590 ( .I(n21960), .ZN(n64040) );
  NAND3_X2 U23598 ( .A1(n41427), .A2(n41437), .A3(n64773), .ZN(n40694) );
  OR2_X1 U23599 ( .A1(n6033), .A2(n12412), .Z(n32901) );
  NOR3_X2 U23606 ( .A1(n59937), .A2(n37904), .A3(n62604), .ZN(n37911) );
  OAI22_X1 U23607 ( .A1(n42247), .A2(n40791), .B1(n42251), .B2(n60709), .ZN(
        n62604) );
  NAND3_X2 U23622 ( .A1(n55483), .A2(n55481), .A3(n62605), .ZN(n55484) );
  NOR2_X2 U23628 ( .A1(n5115), .A2(n8576), .ZN(n64172) );
  NOR2_X2 U23629 ( .A1(n35511), .A2(n17144), .ZN(n35947) );
  XOR2_X1 U23632 ( .A1(n105), .A2(n46668), .Z(n13441) );
  XOR2_X1 U23640 ( .A1(n39581), .A2(n2355), .Z(n39583) );
  XOR2_X1 U23646 ( .A1(n14242), .A2(n62639), .Z(n62607) );
  XOR2_X1 U23647 ( .A1(n62608), .A2(n43823), .Z(n43825) );
  XOR2_X1 U23649 ( .A1(n43821), .A2(n45263), .Z(n62608) );
  NAND2_X1 U23652 ( .A1(n18370), .A2(n35310), .ZN(n65105) );
  NOR2_X1 U23656 ( .A1(n65105), .A2(n60452), .ZN(n8754) );
  NOR2_X2 U23659 ( .A1(n57939), .A2(n4304), .ZN(n63406) );
  NOR3_X2 U23664 ( .A1(n3043), .A2(n62610), .A3(n62609), .ZN(n23439) );
  NAND2_X2 U23666 ( .A1(n3046), .A2(n50057), .ZN(n62609) );
  NAND2_X2 U23671 ( .A1(n64047), .A2(n62612), .ZN(n49072) );
  XOR2_X1 U23674 ( .A1(n20169), .A2(n50244), .Z(n62615) );
  BUF_X2 U23686 ( .I(n52172), .Z(n62616) );
  NOR2_X2 U23687 ( .A1(n49832), .A2(n62861), .ZN(n64887) );
  BUF_X2 U23688 ( .I(n20720), .Z(n62617) );
  NOR4_X2 U23691 ( .A1(n25559), .A2(n62619), .A3(n25562), .A4(n62618), .ZN(
        n25558) );
  XOR2_X1 U23698 ( .A1(n39345), .A2(n24257), .Z(n37301) );
  XOR2_X1 U23700 ( .A1(n2345), .A2(n305), .Z(n63043) );
  XOR2_X1 U23703 ( .A1(n8596), .A2(n45375), .Z(n305) );
  NAND2_X2 U23708 ( .A1(n49283), .A2(n57194), .ZN(n64764) );
  BUF_X2 U23710 ( .I(n8538), .Z(n62620) );
  NOR3_X2 U23713 ( .A1(n15374), .A2(n18406), .A3(n15856), .ZN(n62621) );
  NOR2_X1 U23715 ( .A1(n2444), .A2(n2443), .ZN(n2442) );
  NAND2_X2 U23716 ( .A1(n62622), .A2(n6068), .ZN(n14513) );
  NAND2_X2 U23720 ( .A1(n62623), .A2(n26720), .ZN(n6913) );
  XOR2_X1 U23726 ( .A1(Key[118]), .A2(Ciphertext[87]), .Z(n19196) );
  INV_X2 U23728 ( .I(n4784), .ZN(n62623) );
  NAND2_X2 U23733 ( .A1(n35674), .A2(n35667), .ZN(n6842) );
  NAND2_X2 U23735 ( .A1(n13583), .A2(n18524), .ZN(n35667) );
  NAND4_X2 U23742 ( .A1(n5443), .A2(n5445), .A3(n56818), .A4(n64209), .ZN(
        n64018) );
  AND2_X1 U23743 ( .A1(n43029), .A2(n62624), .Z(n42778) );
  XOR2_X1 U23744 ( .A1(n62625), .A2(n60556), .Z(Plaintext[25]) );
  NAND4_X2 U23745 ( .A1(n53476), .A2(n4963), .A3(n53474), .A4(n53475), .ZN(
        n62625) );
  XOR2_X1 U23755 ( .A1(n8238), .A2(n20620), .Z(n4919) );
  NOR3_X2 U23757 ( .A1(n57764), .A2(n8239), .A3(n8241), .ZN(n8238) );
  XOR2_X1 U23762 ( .A1(n62626), .A2(n44976), .Z(n44977) );
  XOR2_X1 U23763 ( .A1(n45058), .A2(n44974), .Z(n62626) );
  NOR2_X1 U23773 ( .A1(n37956), .A2(n37047), .ZN(n5152) );
  INV_X2 U23775 ( .I(n6237), .ZN(n39987) );
  XOR2_X1 U23776 ( .A1(n62627), .A2(n21531), .Z(n15444) );
  XOR2_X1 U23777 ( .A1(n33065), .A2(n23343), .Z(n62627) );
  NOR2_X1 U23778 ( .A1(n50340), .A2(n64416), .ZN(n60378) );
  AOI21_X2 U23780 ( .A1(n59497), .A2(n62628), .B(n8913), .ZN(n9427) );
  NAND2_X1 U23783 ( .A1(n8917), .A2(n8918), .ZN(n62628) );
  NOR2_X2 U23786 ( .A1(n63873), .A2(n57202), .ZN(n54235) );
  NAND2_X1 U23787 ( .A1(n64088), .A2(n54963), .ZN(n63961) );
  XOR2_X1 U23791 ( .A1(n2472), .A2(n64320), .Z(n63429) );
  XOR2_X1 U23794 ( .A1(n52065), .A2(n65279), .Z(n64177) );
  XOR2_X1 U23798 ( .A1(n63681), .A2(n6004), .Z(n52065) );
  NAND3_X1 U23799 ( .A1(n54972), .A2(n54970), .A3(n54971), .ZN(n63486) );
  XOR2_X1 U23800 ( .A1(n31590), .A2(n19048), .Z(n32011) );
  BUF_X2 U23801 ( .I(n7452), .Z(n62631) );
  BUF_X2 U23805 ( .I(n45436), .Z(n62634) );
  XOR2_X1 U23806 ( .A1(n13104), .A2(n51288), .Z(n52700) );
  XOR2_X1 U23807 ( .A1(n26086), .A2(n51274), .Z(n13104) );
  NAND2_X2 U23808 ( .A1(n56757), .A2(n56803), .ZN(n56805) );
  NOR2_X2 U23814 ( .A1(n56804), .A2(n56805), .ZN(n5444) );
  NAND2_X2 U23817 ( .A1(n56815), .A2(n56775), .ZN(n56804) );
  XOR2_X1 U23819 ( .A1(n25743), .A2(n39407), .Z(n60821) );
  XOR2_X1 U23820 ( .A1(n38991), .A2(n18054), .Z(n39407) );
  XOR2_X1 U23821 ( .A1(n45320), .A2(n62635), .Z(n3099) );
  XOR2_X1 U23822 ( .A1(n13841), .A2(n6803), .Z(n62635) );
  NOR3_X2 U23826 ( .A1(n62636), .A2(n21672), .A3(n21671), .ZN(n10284) );
  INV_X2 U23833 ( .I(n62637), .ZN(n15875) );
  NOR2_X2 U23834 ( .A1(n5348), .A2(n59786), .ZN(n62637) );
  NAND3_X1 U23838 ( .A1(n21490), .A2(n47933), .A3(n50375), .ZN(n62891) );
  NAND2_X2 U23839 ( .A1(n4689), .A2(n43839), .ZN(n43203) );
  XOR2_X1 U23840 ( .A1(n1904), .A2(n2241), .Z(n2740) );
  AOI22_X1 U23841 ( .A1(n62638), .A2(n30841), .B1(n29805), .B2(n7376), .ZN(
        n2437) );
  NAND2_X1 U23842 ( .A1(n10371), .A2(n30214), .ZN(n62638) );
  NOR2_X1 U23845 ( .A1(n14205), .A2(n65005), .ZN(n58844) );
  NAND2_X2 U23848 ( .A1(n16808), .A2(n23055), .ZN(n30226) );
  XOR2_X1 U23851 ( .A1(n466), .A2(n23790), .Z(n62639) );
  NOR2_X2 U23852 ( .A1(n62640), .A2(n15944), .ZN(n63379) );
  OAI21_X2 U23854 ( .A1(n5444), .A2(n56807), .B(n61688), .ZN(n5443) );
  NAND3_X2 U23856 ( .A1(n62642), .A2(n27293), .A3(n62641), .ZN(n27304) );
  NAND2_X1 U23857 ( .A1(n27933), .A2(n29144), .ZN(n62641) );
  OAI21_X2 U23867 ( .A1(n61830), .A2(n62643), .B(n64447), .ZN(n43834) );
  NAND2_X2 U23868 ( .A1(n24894), .A2(n70), .ZN(n62643) );
  XOR2_X1 U23869 ( .A1(n62644), .A2(n4065), .Z(n12426) );
  AND2_X2 U23872 ( .A1(n65089), .A2(n62689), .Z(n40577) );
  NAND3_X1 U23876 ( .A1(n62645), .A2(n49642), .A3(n19172), .ZN(n14309) );
  NAND2_X1 U23878 ( .A1(n48383), .A2(n19523), .ZN(n62645) );
  XOR2_X1 U23882 ( .A1(n59063), .A2(n44464), .Z(n62821) );
  NOR3_X2 U23884 ( .A1(n20029), .A2(n29876), .A3(n29882), .ZN(n58309) );
  XOR2_X1 U23885 ( .A1(n36685), .A2(n39290), .Z(n5376) );
  XOR2_X1 U23891 ( .A1(n39776), .A2(n39579), .Z(n39290) );
  AND2_X2 U23893 ( .A1(n1238), .A2(n2665), .Z(n10341) );
  NOR2_X2 U23894 ( .A1(n62649), .A2(n14243), .ZN(n9375) );
  NOR3_X1 U23898 ( .A1(n5082), .A2(n8997), .A3(n32457), .ZN(n18568) );
  XOR2_X1 U23899 ( .A1(n12177), .A2(n62650), .Z(n6906) );
  XOR2_X1 U23900 ( .A1(n6458), .A2(n18169), .Z(n62650) );
  XOR2_X1 U23903 ( .A1(n19861), .A2(n11239), .Z(n39227) );
  NAND2_X2 U23906 ( .A1(n41720), .A2(n41612), .ZN(n41726) );
  NOR3_X1 U23910 ( .A1(n57568), .A2(n54130), .A3(n54131), .ZN(n62651) );
  OR2_X1 U23914 ( .A1(n3394), .A2(n6030), .Z(n57409) );
  NAND2_X2 U23915 ( .A1(n25500), .A2(n59661), .ZN(n23582) );
  XOR2_X1 U23927 ( .A1(n62652), .A2(n18190), .Z(n10860) );
  XOR2_X1 U23929 ( .A1(n63141), .A2(n11675), .Z(n62652) );
  XOR2_X1 U23931 ( .A1(n8306), .A2(n31702), .Z(n32720) );
  XOR2_X1 U23934 ( .A1(n16581), .A2(n16582), .Z(n31702) );
  NAND3_X2 U23935 ( .A1(n12455), .A2(n5373), .A3(n8130), .ZN(n49319) );
  INV_X1 U23936 ( .I(n17873), .ZN(n62653) );
  NAND3_X2 U23940 ( .A1(n41621), .A2(n41622), .A3(n41620), .ZN(n44578) );
  XOR2_X1 U23941 ( .A1(n2978), .A2(n59539), .Z(n64420) );
  NOR2_X2 U23942 ( .A1(n43701), .A2(n37917), .ZN(n43699) );
  NOR3_X2 U23944 ( .A1(n35947), .A2(n62655), .A3(n62654), .ZN(n8173) );
  NAND2_X2 U23948 ( .A1(n16958), .A2(n19654), .ZN(n64444) );
  NAND2_X2 U23951 ( .A1(n22100), .A2(n22099), .ZN(n16958) );
  INV_X1 U23952 ( .I(n34258), .ZN(n62908) );
  AOI21_X1 U23953 ( .A1(n34255), .A2(n34356), .B(n62908), .ZN(n62907) );
  XOR2_X1 U23954 ( .A1(n24640), .A2(n23222), .Z(n51592) );
  NAND2_X2 U23956 ( .A1(n40890), .A2(n40891), .ZN(n17223) );
  NAND2_X2 U23957 ( .A1(n18144), .A2(n20530), .ZN(n36395) );
  OAI21_X2 U23958 ( .A1(n62657), .A2(n65265), .B(n9801), .ZN(n24570) );
  NAND2_X1 U23962 ( .A1(n12927), .A2(n42359), .ZN(n62657) );
  XOR2_X1 U23966 ( .A1(n38501), .A2(n38500), .Z(n39273) );
  XOR2_X1 U23967 ( .A1(n39406), .A2(n13458), .Z(n38501) );
  XOR2_X1 U23968 ( .A1(n2130), .A2(n62658), .Z(n32493) );
  AND2_X2 U23970 ( .A1(n21064), .A2(n28025), .Z(n7452) );
  XOR2_X1 U23971 ( .A1(Ciphertext[58]), .A2(Key[11]), .Z(n28025) );
  NAND2_X1 U23973 ( .A1(n35603), .A2(n36262), .ZN(n63399) );
  NOR2_X1 U23976 ( .A1(n63689), .A2(n29199), .ZN(n14303) );
  XOR2_X1 U23977 ( .A1(n2950), .A2(n58814), .Z(n51591) );
  NAND3_X2 U23983 ( .A1(n24608), .A2(n24607), .A3(n45469), .ZN(n2950) );
  OR3_X1 U23987 ( .A1(n56630), .A2(n56629), .A3(n56631), .Z(n51452) );
  NAND2_X2 U23993 ( .A1(n62659), .A2(n62705), .ZN(n45442) );
  OAI21_X1 U23994 ( .A1(n11863), .A2(n61376), .B(n62660), .ZN(n64148) );
  INV_X1 U23995 ( .I(n30151), .ZN(n62660) );
  BUF_X4 U23996 ( .I(n30148), .Z(n21176) );
  AND2_X1 U24002 ( .A1(n56813), .A2(n23879), .Z(n62771) );
  INV_X2 U24003 ( .I(n8287), .ZN(n22042) );
  BUF_X2 U24006 ( .I(n25794), .Z(n22521) );
  CLKBUF_X4 U24016 ( .I(n33721), .Z(n65160) );
  NAND2_X2 U24022 ( .A1(n10205), .A2(n11656), .ZN(n30250) );
  AND2_X1 U24026 ( .A1(n47101), .A2(n18099), .Z(n23795) );
  NAND2_X2 U24027 ( .A1(n51463), .A2(n57060), .ZN(n64550) );
  OAI21_X2 U24029 ( .A1(n61772), .A2(n57060), .B(n64550), .ZN(n51472) );
  AND3_X1 U24030 ( .A1(n36608), .A2(n62010), .A3(n35103), .Z(n63761) );
  NAND2_X2 U24035 ( .A1(n53493), .A2(n53506), .ZN(n53513) );
  NAND2_X2 U24039 ( .A1(n62662), .A2(n58053), .ZN(n17127) );
  NOR2_X1 U24041 ( .A1(n57357), .A2(n58204), .ZN(n62662) );
  BUF_X2 U24044 ( .I(n4226), .Z(n62664) );
  NAND2_X2 U24046 ( .A1(n57621), .A2(n16491), .ZN(n25707) );
  XOR2_X1 U24053 ( .A1(n62665), .A2(n3875), .Z(n2309) );
  XOR2_X1 U24058 ( .A1(n64658), .A2(n45096), .Z(n62665) );
  NAND3_X2 U24059 ( .A1(n50808), .A2(n62779), .A3(n64666), .ZN(n64767) );
  NAND3_X2 U24064 ( .A1(n62667), .A2(n54959), .A3(n60530), .ZN(n26014) );
  NAND3_X2 U24066 ( .A1(n59080), .A2(n64879), .A3(n59079), .ZN(n62667) );
  NAND2_X1 U24069 ( .A1(n54522), .A2(n63155), .ZN(n63154) );
  XOR2_X1 U24073 ( .A1(n62668), .A2(n56784), .Z(Plaintext[171]) );
  NAND3_X1 U24076 ( .A1(n56783), .A2(n56782), .A3(n56781), .ZN(n62668) );
  NAND2_X1 U24079 ( .A1(n2333), .A2(n58472), .ZN(n2332) );
  AOI22_X2 U24080 ( .A1(n10788), .A2(n10789), .B1(n16263), .B2(n36149), .ZN(
        n64368) );
  NAND2_X2 U24082 ( .A1(n17018), .A2(n2323), .ZN(n4189) );
  INV_X2 U24085 ( .I(n8602), .ZN(n62670) );
  XOR2_X1 U24086 ( .A1(n21321), .A2(n30897), .Z(n12173) );
  XOR2_X1 U24093 ( .A1(n2023), .A2(n58440), .Z(n21321) );
  NOR2_X1 U24097 ( .A1(n26173), .A2(n62679), .ZN(n26172) );
  XOR2_X1 U24104 ( .A1(n62671), .A2(n6722), .Z(n23760) );
  XOR2_X1 U24106 ( .A1(n61538), .A2(n29908), .Z(n62671) );
  AOI21_X1 U24107 ( .A1(n18519), .A2(n18523), .B(n7303), .ZN(n20560) );
  NOR2_X1 U24108 ( .A1(n28619), .A2(n61771), .ZN(n28638) );
  NAND2_X2 U24110 ( .A1(n14212), .A2(n63525), .ZN(n28619) );
  NOR2_X1 U24114 ( .A1(n20391), .A2(n30748), .ZN(n30002) );
  NOR2_X2 U24118 ( .A1(n37050), .A2(n31306), .ZN(n35480) );
  NOR2_X2 U24120 ( .A1(n25312), .A2(n21564), .ZN(n51482) );
  NAND2_X1 U24121 ( .A1(n59820), .A2(n45772), .ZN(n6285) );
  NAND4_X2 U24132 ( .A1(n36504), .A2(n62673), .A3(n36503), .A4(n36501), .ZN(
        n39551) );
  AOI22_X2 U24134 ( .A1(n36499), .A2(n36498), .B1(n36497), .B2(n36496), .ZN(
        n62673) );
  XOR2_X1 U24138 ( .A1(n50717), .A2(n52013), .Z(n2061) );
  NOR2_X2 U24148 ( .A1(n17678), .A2(n17677), .ZN(n50717) );
  NOR2_X2 U24155 ( .A1(n15428), .A2(n62674), .ZN(n17977) );
  OR3_X1 U24159 ( .A1(n16013), .A2(n18853), .A3(n965), .Z(n62674) );
  XOR2_X1 U24163 ( .A1(n62675), .A2(n12068), .Z(n38234) );
  XOR2_X1 U24164 ( .A1(n38222), .A2(n38233), .Z(n62675) );
  XOR2_X1 U24165 ( .A1(n62676), .A2(n50475), .Z(Plaintext[41]) );
  NAND4_X2 U24166 ( .A1(n50474), .A2(n50471), .A3(n50473), .A4(n50472), .ZN(
        n62676) );
  NAND2_X1 U24167 ( .A1(n5566), .A2(n5564), .ZN(n62677) );
  AOI21_X2 U24169 ( .A1(n21018), .A2(n35976), .B(n62678), .ZN(n14877) );
  OAI22_X2 U24175 ( .A1(n64024), .A2(n35965), .B1(n35357), .B2(n13769), .ZN(
        n62678) );
  NAND3_X2 U24176 ( .A1(n18144), .A2(n36385), .A3(n36057), .ZN(n35454) );
  XOR2_X1 U24181 ( .A1(n44531), .A2(n57489), .Z(n58692) );
  AOI21_X1 U24182 ( .A1(n48672), .A2(n18498), .B(n63913), .ZN(n25912) );
  XOR2_X1 U24187 ( .A1(n50916), .A2(n14870), .Z(n10953) );
  XOR2_X1 U24188 ( .A1(n50761), .A2(n9619), .Z(n50916) );
  XOR2_X1 U24190 ( .A1(n51035), .A2(n24640), .Z(n63367) );
  NAND3_X2 U24192 ( .A1(n64540), .A2(n64539), .A3(n45176), .ZN(n24640) );
  INV_X2 U24193 ( .I(n62680), .ZN(n3065) );
  NAND2_X2 U24195 ( .A1(n3658), .A2(n49929), .ZN(n62680) );
  NAND3_X1 U24196 ( .A1(n41899), .A2(n62474), .A3(n41096), .ZN(n63371) );
  AND2_X1 U24197 ( .A1(n7541), .A2(n1663), .Z(n9549) );
  NOR3_X2 U24198 ( .A1(n5129), .A2(n1615), .A3(n52126), .ZN(n15820) );
  AND2_X1 U24201 ( .A1(n42140), .A2(n40550), .Z(n41340) );
  NAND2_X2 U24202 ( .A1(n6633), .A2(n1469), .ZN(n48804) );
  BUF_X2 U24204 ( .I(n35653), .Z(n62683) );
  INV_X2 U24205 ( .I(n35340), .ZN(n36200) );
  NAND2_X2 U24210 ( .A1(n26243), .A2(n36202), .ZN(n35340) );
  NOR3_X2 U24211 ( .A1(n60898), .A2(n3661), .A3(n3659), .ZN(n49630) );
  XOR2_X1 U24213 ( .A1(n10952), .A2(n8954), .Z(n13026) );
  NAND2_X1 U24214 ( .A1(n34990), .A2(n30470), .ZN(n30471) );
  NAND2_X1 U24217 ( .A1(n47533), .A2(n48605), .ZN(n62981) );
  XOR2_X1 U24221 ( .A1(n20270), .A2(n22321), .Z(n61226) );
  XOR2_X1 U24222 ( .A1(n31199), .A2(n62684), .Z(n14716) );
  XOR2_X1 U24223 ( .A1(n15840), .A2(n13992), .Z(n62684) );
  NAND4_X2 U24225 ( .A1(n6673), .A2(n6674), .A3(n6672), .A4(n11394), .ZN(
        n62713) );
  AOI21_X2 U24230 ( .A1(n62685), .A2(n28783), .B(n58481), .ZN(n32744) );
  AOI21_X2 U24231 ( .A1(n28776), .A2(n30676), .B(n30242), .ZN(n62685) );
  XOR2_X1 U24234 ( .A1(n3388), .A2(n22332), .Z(n58125) );
  XOR2_X1 U24237 ( .A1(n62687), .A2(n12260), .Z(n62982) );
  XOR2_X1 U24240 ( .A1(n16701), .A2(n62688), .Z(n62687) );
  XOR2_X1 U24246 ( .A1(n57622), .A2(n4440), .Z(n7642) );
  INV_X2 U24247 ( .I(n62689), .ZN(n24645) );
  XOR2_X1 U24248 ( .A1(n7381), .A2(n12380), .Z(n8427) );
  NAND3_X2 U24253 ( .A1(n48267), .A2(n48266), .A3(n49130), .ZN(n2078) );
  XOR2_X1 U24255 ( .A1(n64587), .A2(n65251), .Z(n48404) );
  NAND3_X2 U24258 ( .A1(n34235), .A2(n34234), .A3(n34718), .ZN(n62691) );
  NAND2_X2 U24264 ( .A1(n62859), .A2(n217), .ZN(n14731) );
  OR2_X2 U24265 ( .A1(n24645), .A2(n65089), .Z(n41898) );
  NAND2_X2 U24267 ( .A1(n37677), .A2(n12129), .ZN(n6989) );
  NAND2_X2 U24269 ( .A1(n11227), .A2(n24595), .ZN(n37677) );
  INV_X2 U24270 ( .I(n62693), .ZN(n732) );
  NAND2_X2 U24272 ( .A1(n8203), .A2(n55302), .ZN(n9076) );
  NAND2_X2 U24273 ( .A1(n9076), .A2(n55303), .ZN(n63927) );
  XOR2_X1 U24281 ( .A1(n32637), .A2(n32636), .Z(n62694) );
  NAND2_X2 U24288 ( .A1(n23415), .A2(n13911), .ZN(n9119) );
  NAND2_X2 U24290 ( .A1(n63600), .A2(n26234), .ZN(n23415) );
  AOI22_X1 U24292 ( .A1(n62696), .A2(n30622), .B1(n30617), .B2(n30616), .ZN(
        n30626) );
  INV_X1 U24294 ( .I(n30613), .ZN(n62696) );
  NAND2_X1 U24295 ( .A1(n30348), .A2(n29586), .ZN(n30613) );
  NOR2_X2 U24296 ( .A1(n62697), .A2(n32682), .ZN(n32688) );
  XNOR2_X1 U24299 ( .A1(n32027), .A2(n8262), .ZN(n62792) );
  NAND2_X2 U24300 ( .A1(n8225), .A2(n60241), .ZN(n47834) );
  NOR2_X2 U24305 ( .A1(n21081), .A2(n64850), .ZN(n14879) );
  NOR2_X2 U24307 ( .A1(n12028), .A2(n1237), .ZN(n64850) );
  NAND3_X1 U24309 ( .A1(n59710), .A2(n40), .A3(n21029), .ZN(n29588) );
  OR2_X2 U24311 ( .A1(n39065), .A2(n39064), .Z(n41660) );
  OAI22_X2 U24314 ( .A1(n39059), .A2(n39058), .B1(n59593), .B2(n64040), .ZN(
        n39065) );
  OR2_X1 U24316 ( .A1(n35228), .A2(n62698), .Z(n34410) );
  NAND2_X2 U24326 ( .A1(n19584), .A2(n8266), .ZN(n7253) );
  XOR2_X1 U24327 ( .A1(n51570), .A2(n17127), .Z(n64041) );
  NAND3_X2 U24333 ( .A1(n19324), .A2(n20390), .A3(n20417), .ZN(n51570) );
  INV_X4 U24343 ( .I(n49072), .ZN(n20458) );
  INV_X2 U24345 ( .I(n13667), .ZN(n4312) );
  NAND2_X2 U24350 ( .A1(n52762), .A2(n17012), .ZN(n13667) );
  INV_X4 U24352 ( .I(n42944), .ZN(n25806) );
  NAND3_X2 U24355 ( .A1(n61652), .A2(n13889), .A3(n60533), .ZN(n16653) );
  XOR2_X1 U24359 ( .A1(n62701), .A2(n44885), .Z(n19543) );
  XOR2_X1 U24361 ( .A1(n57759), .A2(n57360), .Z(n62701) );
  AOI21_X2 U24364 ( .A1(n53466), .A2(n53465), .B(n62702), .ZN(n53476) );
  NAND3_X2 U24365 ( .A1(n53511), .A2(n60796), .A3(n53497), .ZN(n62702) );
  XOR2_X1 U24367 ( .A1(n46705), .A2(n21308), .Z(n62834) );
  XOR2_X1 U24368 ( .A1(n21307), .A2(n45875), .Z(n46705) );
  XOR2_X1 U24373 ( .A1(n62703), .A2(n50644), .Z(n59032) );
  XOR2_X1 U24374 ( .A1(n50679), .A2(n51941), .Z(n62703) );
  XOR2_X1 U24375 ( .A1(n57832), .A2(n24458), .Z(n6003) );
  XOR2_X1 U24379 ( .A1(n60661), .A2(n32619), .Z(n24458) );
  AND2_X2 U24381 ( .A1(n23933), .A2(n17133), .Z(n8688) );
  NOR2_X2 U24382 ( .A1(n53383), .A2(n53376), .ZN(n53379) );
  NAND2_X1 U24383 ( .A1(n47126), .A2(n64869), .ZN(n63740) );
  NOR3_X2 U24385 ( .A1(n6629), .A2(n62704), .A3(n38546), .ZN(n6628) );
  NAND2_X1 U24387 ( .A1(n49440), .A2(n1637), .ZN(n49362) );
  AOI21_X2 U24390 ( .A1(n62707), .A2(n62501), .B(n62706), .ZN(n62705) );
  NOR2_X1 U24398 ( .A1(n45434), .A2(n62501), .ZN(n62706) );
  INV_X1 U24399 ( .I(n45433), .ZN(n62707) );
  NAND3_X2 U24401 ( .A1(n10973), .A2(n45894), .A3(n62708), .ZN(n45895) );
  NOR2_X1 U24406 ( .A1(n46763), .A2(n64036), .ZN(n62709) );
  INV_X4 U24407 ( .I(n5055), .ZN(n49014) );
  NOR2_X2 U24408 ( .A1(n19932), .A2(n65215), .ZN(n5055) );
  BUF_X4 U24409 ( .I(n25976), .Z(n64377) );
  NAND2_X2 U24411 ( .A1(n62710), .A2(n44694), .ZN(n22664) );
  OAI21_X2 U24417 ( .A1(n63835), .A2(n63836), .B(n47014), .ZN(n62710) );
  BUF_X2 U24418 ( .I(n55231), .Z(n62711) );
  XOR2_X1 U24419 ( .A1(n62712), .A2(n12177), .Z(n7904) );
  XOR2_X1 U24420 ( .A1(n2578), .A2(n39553), .Z(n62712) );
  NAND3_X2 U24421 ( .A1(n2001), .A2(n53379), .A3(n52845), .ZN(n53606) );
  XOR2_X1 U24424 ( .A1(n5942), .A2(n50785), .Z(n14105) );
  XOR2_X1 U24425 ( .A1(n50615), .A2(n16508), .Z(n50785) );
  NOR2_X2 U24427 ( .A1(n21605), .A2(n24351), .ZN(n2885) );
  INV_X2 U24434 ( .I(n34575), .ZN(n24351) );
  NOR4_X2 U24436 ( .A1(n3720), .A2(n3718), .A3(n684), .A4(n3722), .ZN(n34575)
         );
  NAND2_X2 U24439 ( .A1(n20091), .A2(n12779), .ZN(n22684) );
  NOR2_X2 U24440 ( .A1(n62713), .A2(n6675), .ZN(n11557) );
  INV_X2 U24441 ( .I(n45968), .ZN(n47825) );
  NOR2_X2 U24442 ( .A1(n19645), .A2(n65074), .ZN(n45968) );
  AND2_X1 U24443 ( .A1(n20627), .A2(n62715), .Z(n17743) );
  XOR2_X1 U24445 ( .A1(n33042), .A2(n33032), .Z(n64221) );
  NAND2_X2 U24447 ( .A1(n16402), .A2(n23689), .ZN(n65205) );
  NAND2_X2 U24448 ( .A1(n62716), .A2(n35766), .ZN(n7074) );
  AND3_X1 U24449 ( .A1(n35767), .A2(n10808), .A3(n35768), .Z(n62716) );
  XOR2_X1 U24450 ( .A1(n62717), .A2(n52113), .Z(n11481) );
  XOR2_X1 U24451 ( .A1(n21361), .A2(n62985), .Z(n62717) );
  AOI21_X2 U24453 ( .A1(n7841), .A2(n33003), .B(n62718), .ZN(n14219) );
  NAND2_X2 U24454 ( .A1(n7838), .A2(n7839), .ZN(n62718) );
  NOR3_X1 U24456 ( .A1(n10554), .A2(n40312), .A3(n21207), .ZN(n11048) );
  INV_X2 U24463 ( .I(n25643), .ZN(n26088) );
  NOR2_X2 U24467 ( .A1(n18100), .A2(n19160), .ZN(n1386) );
  INV_X2 U24473 ( .I(n60935), .ZN(n18100) );
  NAND2_X2 U24482 ( .A1(n16943), .A2(n22343), .ZN(n55224) );
  AOI22_X1 U24483 ( .A1(n53111), .A2(n53110), .B1(n53112), .B2(n23830), .ZN(
        n53122) );
  NAND2_X2 U24486 ( .A1(n53078), .A2(n53083), .ZN(n53054) );
  NAND2_X2 U24487 ( .A1(n64816), .A2(n17328), .ZN(n53078) );
  XOR2_X1 U24493 ( .A1(n63723), .A2(n51012), .Z(n62722) );
  XOR2_X1 U24494 ( .A1(Ciphertext[88]), .A2(Key[29]), .Z(n21499) );
  NAND3_X2 U24496 ( .A1(n16603), .A2(n29967), .A3(n29966), .ZN(n16820) );
  NAND2_X1 U24498 ( .A1(n62902), .A2(n64322), .ZN(n3410) );
  NAND3_X2 U24499 ( .A1(n33925), .A2(n35325), .A3(n12184), .ZN(n16726) );
  NAND2_X2 U24500 ( .A1(n31281), .A2(n64998), .ZN(n62725) );
  INV_X2 U24501 ( .I(n62726), .ZN(n55445) );
  AND2_X1 U24505 ( .A1(n52117), .A2(n54998), .Z(n62726) );
  NOR2_X1 U24508 ( .A1(n57461), .A2(n42258), .ZN(n3564) );
  XOR2_X1 U24513 ( .A1(n62727), .A2(n37722), .Z(n8866) );
  XOR2_X1 U24514 ( .A1(n37720), .A2(n37721), .Z(n62727) );
  XOR2_X1 U24516 ( .A1(n9288), .A2(n62729), .Z(n2861) );
  XOR2_X1 U24517 ( .A1(n2952), .A2(n30941), .Z(n62729) );
  NOR3_X2 U24521 ( .A1(n57820), .A2(n5698), .A3(n5696), .ZN(n15065) );
  NOR2_X1 U24524 ( .A1(n62730), .A2(n36168), .ZN(n58942) );
  NAND2_X1 U24532 ( .A1(n25294), .A2(n58938), .ZN(n62730) );
  XOR2_X1 U24537 ( .A1(n62731), .A2(n45866), .Z(n651) );
  XOR2_X1 U24543 ( .A1(n14037), .A2(n63821), .Z(n62731) );
  NOR2_X2 U24545 ( .A1(n61561), .A2(n8942), .ZN(n41476) );
  INV_X2 U24546 ( .I(n40414), .ZN(n8942) );
  NOR2_X2 U24553 ( .A1(n39987), .A2(n38758), .ZN(n40414) );
  XOR2_X1 U24558 ( .A1(n62732), .A2(n50783), .Z(n14178) );
  XOR2_X1 U24565 ( .A1(n14181), .A2(n60914), .Z(n62732) );
  XOR2_X1 U24566 ( .A1(n11091), .A2(n11256), .Z(n11090) );
  AOI21_X2 U24568 ( .A1(n48345), .A2(n14561), .B(n63663), .ZN(n16692) );
  AOI21_X1 U24569 ( .A1(n63265), .A2(n63264), .B(n24856), .ZN(n24855) );
  NAND2_X2 U24570 ( .A1(n12112), .A2(n61383), .ZN(n30231) );
  NAND3_X2 U24571 ( .A1(n31957), .A2(n31958), .A3(n11000), .ZN(n23220) );
  XOR2_X1 U24573 ( .A1(n22573), .A2(n45115), .Z(n61116) );
  NOR2_X2 U24576 ( .A1(n24117), .A2(n22343), .ZN(n58813) );
  NOR2_X2 U24577 ( .A1(n62735), .A2(n64407), .ZN(n17377) );
  NOR2_X2 U24584 ( .A1(n34116), .A2(n34113), .ZN(n64407) );
  AND2_X1 U24585 ( .A1(n32869), .A2(n32870), .Z(n62735) );
  NAND2_X1 U24586 ( .A1(n34441), .A2(n61810), .ZN(n31954) );
  NOR2_X1 U24590 ( .A1(n62736), .A2(n63894), .ZN(n64816) );
  NAND2_X1 U24591 ( .A1(n52885), .A2(n52887), .ZN(n62736) );
  NAND4_X1 U24592 ( .A1(n56169), .A2(n56172), .A3(n56189), .A4(n17606), .ZN(
        n24807) );
  OAI21_X2 U24594 ( .A1(n24628), .A2(n24626), .B(n62737), .ZN(n37821) );
  NAND2_X2 U24597 ( .A1(n62738), .A2(n40884), .ZN(n46305) );
  INV_X4 U24600 ( .I(n7187), .ZN(n41568) );
  NAND2_X2 U24605 ( .A1(n58729), .A2(n58578), .ZN(n7187) );
  NAND2_X1 U24613 ( .A1(n11126), .A2(n63952), .ZN(n11125) );
  BUF_X2 U24614 ( .I(n45991), .Z(n62739) );
  NOR2_X2 U24616 ( .A1(n6129), .A2(n62186), .ZN(n65282) );
  BUF_X2 U24619 ( .I(n20072), .Z(n62740) );
  NOR2_X2 U24622 ( .A1(n27582), .A2(n23737), .ZN(n62784) );
  NAND3_X2 U24623 ( .A1(n58975), .A2(n48847), .A3(n49525), .ZN(n49192) );
  NAND2_X2 U24625 ( .A1(n19646), .A2(n48440), .ZN(n46004) );
  XOR2_X1 U24626 ( .A1(n38304), .A2(n23922), .Z(n7601) );
  NAND4_X2 U24627 ( .A1(n35126), .A2(n35125), .A3(n16955), .A4(n16956), .ZN(
        n38304) );
  OAI21_X2 U24629 ( .A1(n41613), .A2(n41982), .B(n22999), .ZN(n42353) );
  NOR2_X2 U24633 ( .A1(n53888), .A2(n53889), .ZN(n53950) );
  NAND3_X2 U24638 ( .A1(n22718), .A2(n53841), .A3(n62977), .ZN(n53888) );
  NOR2_X2 U24640 ( .A1(n13008), .A2(n13003), .ZN(n58273) );
  OAI21_X1 U24642 ( .A1(n62743), .A2(n62742), .B(n30447), .ZN(n58408) );
  NOR2_X1 U24643 ( .A1(n29428), .A2(n1558), .ZN(n62742) );
  NOR2_X1 U24645 ( .A1(n29427), .A2(n29426), .ZN(n62743) );
  INV_X4 U24646 ( .I(n17223), .ZN(n58572) );
  XOR2_X1 U24647 ( .A1(n62745), .A2(n2886), .Z(n9158) );
  XOR2_X1 U24650 ( .A1(n49719), .A2(n49718), .Z(n62745) );
  NAND3_X2 U24654 ( .A1(n20798), .A2(n12747), .A3(n20799), .ZN(n35109) );
  XOR2_X1 U24659 ( .A1(n9746), .A2(n9745), .Z(n19393) );
  XOR2_X1 U24660 ( .A1(n44839), .A2(n19680), .Z(n44861) );
  NAND2_X1 U24662 ( .A1(n50045), .A2(n18502), .ZN(n63943) );
  INV_X1 U24664 ( .I(n18486), .ZN(n63412) );
  XOR2_X1 U24668 ( .A1(n44733), .A2(n44730), .Z(n64827) );
  XOR2_X1 U24674 ( .A1(n4343), .A2(n14513), .Z(n44733) );
  NOR2_X1 U24684 ( .A1(n12643), .A2(n23488), .ZN(n62970) );
  NAND3_X2 U24685 ( .A1(n13787), .A2(n13785), .A3(n13786), .ZN(n10292) );
  NOR2_X2 U24694 ( .A1(n17144), .A2(n22461), .ZN(n36913) );
  NAND4_X2 U24696 ( .A1(n61614), .A2(n61613), .A3(n56800), .A4(n56799), .ZN(
        n56802) );
  NAND3_X1 U24697 ( .A1(n30050), .A2(n1349), .A3(n30048), .ZN(n2284) );
  NAND2_X1 U24699 ( .A1(n30050), .A2(n1349), .ZN(n2252) );
  XOR2_X1 U24700 ( .A1(n62749), .A2(n21348), .Z(n39001) );
  XOR2_X1 U24702 ( .A1(n5555), .A2(n57096), .Z(n62749) );
  AOI22_X2 U24704 ( .A1(n40289), .A2(n40228), .B1(n40306), .B2(n40287), .ZN(
        n39322) );
  XOR2_X1 U24706 ( .A1(n38276), .A2(n6302), .Z(n39207) );
  NAND2_X2 U24710 ( .A1(n24961), .A2(n24962), .ZN(n38276) );
  NOR2_X2 U24712 ( .A1(n21478), .A2(n20025), .ZN(n27735) );
  NOR2_X2 U24714 ( .A1(n19591), .A2(n39427), .ZN(n43104) );
  NOR2_X2 U24716 ( .A1(n24033), .A2(n37249), .ZN(n37447) );
  OAI21_X2 U24718 ( .A1(n43106), .A2(n20844), .B(n62750), .ZN(n3006) );
  NOR2_X2 U24719 ( .A1(n42425), .A2(n24179), .ZN(n62750) );
  XOR2_X1 U24722 ( .A1(n62751), .A2(n55889), .Z(Plaintext[136]) );
  NAND4_X2 U24723 ( .A1(n11783), .A2(n55901), .A3(n19072), .A4(n11785), .ZN(
        n62751) );
  XOR2_X1 U24725 ( .A1(n58235), .A2(n38856), .Z(n3715) );
  NAND2_X2 U24727 ( .A1(n37600), .A2(n37601), .ZN(n38856) );
  XOR2_X1 U24731 ( .A1(n16688), .A2(n33836), .Z(n58732) );
  NOR3_X2 U24732 ( .A1(n5494), .A2(n28991), .A3(n5493), .ZN(n65193) );
  NAND3_X1 U24733 ( .A1(n22273), .A2(n22643), .A3(n10458), .ZN(n26675) );
  NOR2_X1 U24735 ( .A1(n56883), .A2(n12454), .ZN(n17647) );
  NOR3_X2 U24736 ( .A1(n56881), .A2(n56836), .A3(n21879), .ZN(n56883) );
  BUF_X4 U24737 ( .I(n24210), .Z(n19646) );
  NAND3_X1 U24738 ( .A1(n22273), .A2(n11225), .A3(n27431), .ZN(n26674) );
  NAND2_X2 U24739 ( .A1(n54767), .A2(n19491), .ZN(n54709) );
  BUF_X4 U24745 ( .I(n23284), .Z(n7138) );
  NAND2_X2 U24749 ( .A1(n62784), .A2(n26660), .ZN(n26500) );
  XOR2_X1 U24753 ( .A1(n2410), .A2(n62753), .Z(n21856) );
  XOR2_X1 U24758 ( .A1(n21756), .A2(n51316), .Z(n62753) );
  INV_X2 U24760 ( .I(n58835), .ZN(n19645) );
  XOR2_X1 U24761 ( .A1(n4858), .A2(n13299), .Z(n13298) );
  XOR2_X1 U24762 ( .A1(n62754), .A2(n57408), .Z(n51930) );
  XOR2_X1 U24764 ( .A1(n51595), .A2(n51594), .Z(n62754) );
  XOR2_X1 U24765 ( .A1(n13622), .A2(n10510), .Z(n7540) );
  NAND2_X2 U24766 ( .A1(n56107), .A2(n56084), .ZN(n56103) );
  XOR2_X1 U24767 ( .A1(n15087), .A2(n29070), .Z(n25402) );
  NAND2_X2 U24768 ( .A1(n2144), .A2(n2143), .ZN(n15087) );
  INV_X2 U24771 ( .I(n37234), .ZN(n37455) );
  NAND2_X2 U24772 ( .A1(n20596), .A2(n20597), .ZN(n37234) );
  INV_X4 U24775 ( .I(n24294), .ZN(n43573) );
  XOR2_X1 U24781 ( .A1(n62761), .A2(n18781), .Z(n63127) );
  XOR2_X1 U24782 ( .A1(n38901), .A2(n38144), .Z(n20229) );
  XOR2_X1 U24783 ( .A1(n57757), .A2(n37673), .Z(n38144) );
  NAND3_X2 U24784 ( .A1(n16456), .A2(n15857), .A3(n16455), .ZN(n64477) );
  NOR2_X1 U24793 ( .A1(n3330), .A2(n28005), .ZN(n3382) );
  INV_X2 U24794 ( .I(n53655), .ZN(n63929) );
  AND2_X2 U24795 ( .A1(n5547), .A2(n64481), .Z(n26547) );
  NAND2_X2 U24807 ( .A1(n64579), .A2(n62903), .ZN(n40015) );
  INV_X4 U24813 ( .I(n13622), .ZN(n26022) );
  NOR3_X2 U24816 ( .A1(n1160), .A2(n12000), .A3(n11998), .ZN(n24244) );
  XOR2_X1 U24818 ( .A1(n59752), .A2(n865), .Z(n17384) );
  XOR2_X1 U24819 ( .A1(n7459), .A2(n62757), .Z(n50644) );
  XOR2_X1 U24821 ( .A1(n50549), .A2(n63010), .Z(n62757) );
  INV_X1 U24824 ( .I(n48206), .ZN(n62758) );
  NOR2_X1 U24826 ( .A1(n5704), .A2(n61715), .ZN(n64099) );
  NAND2_X2 U24838 ( .A1(n60467), .A2(n7098), .ZN(n49936) );
  OR2_X1 U24847 ( .A1(n7979), .A2(n28730), .Z(n29845) );
  XOR2_X1 U24850 ( .A1(n62759), .A2(n23455), .Z(Plaintext[71]) );
  NAND3_X1 U24860 ( .A1(n60104), .A2(n54429), .A3(n54428), .ZN(n62759) );
  INV_X1 U24861 ( .I(n35478), .ZN(n62983) );
  NAND2_X2 U24862 ( .A1(n58896), .A2(n54543), .ZN(n23453) );
  XOR2_X1 U24863 ( .A1(n17239), .A2(n62762), .Z(n62761) );
  AOI21_X1 U24864 ( .A1(n47074), .A2(n63923), .B(n49905), .ZN(n47078) );
  AND2_X1 U24867 ( .A1(n52953), .A2(n18145), .Z(n62763) );
  NAND2_X1 U24870 ( .A1(n26983), .A2(n26982), .ZN(n63253) );
  OR2_X1 U24874 ( .A1(n37582), .A2(n62764), .Z(n11793) );
  NOR2_X2 U24876 ( .A1(n35520), .A2(n10096), .ZN(n37582) );
  BUF_X4 U24877 ( .I(n14488), .Z(n64166) );
  NAND3_X1 U24880 ( .A1(n43149), .A2(n43148), .A3(n43147), .ZN(n62765) );
  INV_X2 U24883 ( .I(n24930), .ZN(n52617) );
  NAND3_X2 U24884 ( .A1(n24928), .A2(n1101), .A3(n13259), .ZN(n24930) );
  NAND3_X2 U24885 ( .A1(n16383), .A2(n55218), .A3(n55225), .ZN(n55205) );
  OAI21_X1 U24886 ( .A1(n55788), .A2(n55759), .B(n10736), .ZN(n11687) );
  NAND2_X2 U24887 ( .A1(n24958), .A2(n55812), .ZN(n10736) );
  NOR2_X2 U24889 ( .A1(n62767), .A2(n62766), .ZN(n59316) );
  AOI21_X1 U24895 ( .A1(n47354), .A2(n47353), .B(n4323), .ZN(n47358) );
  BUF_X2 U24897 ( .I(n17211), .Z(n62769) );
  NAND2_X2 U24904 ( .A1(n53247), .A2(n53267), .ZN(n60179) );
  OAI21_X1 U24906 ( .A1(n22907), .A2(n22728), .B(n22727), .ZN(n41208) );
  NAND2_X1 U24907 ( .A1(n43578), .A2(n12154), .ZN(n43584) );
  NOR2_X1 U24909 ( .A1(n26153), .A2(n64596), .ZN(n15203) );
  XOR2_X1 U24911 ( .A1(n62770), .A2(n52026), .Z(n24470) );
  XOR2_X1 U24915 ( .A1(n52024), .A2(n52025), .Z(n62770) );
  NAND2_X1 U24920 ( .A1(n62932), .A2(n42442), .ZN(n24345) );
  NOR2_X1 U24923 ( .A1(n8398), .A2(n58647), .ZN(n63565) );
  NAND3_X2 U24930 ( .A1(n58136), .A2(n48413), .A3(n48823), .ZN(n48061) );
  AOI21_X1 U24936 ( .A1(n62771), .A2(n56814), .B(n5446), .ZN(n5445) );
  NOR3_X2 U24938 ( .A1(n41588), .A2(n43350), .A3(n61198), .ZN(n42749) );
  NOR2_X2 U24939 ( .A1(n61134), .A2(n1494), .ZN(n41588) );
  XOR2_X1 U24942 ( .A1(n31989), .A2(n31993), .Z(n17105) );
  NAND2_X2 U24944 ( .A1(n6058), .A2(n42299), .ZN(n41850) );
  XOR2_X1 U24945 ( .A1(n15755), .A2(n25713), .Z(n60889) );
  INV_X2 U24950 ( .I(n65088), .ZN(n61531) );
  OAI21_X1 U24953 ( .A1(n62774), .A2(n26664), .B(n27569), .ZN(n20875) );
  NAND2_X1 U24954 ( .A1(n457), .A2(n26500), .ZN(n62774) );
  XOR2_X1 U24956 ( .A1(n38770), .A2(n23049), .Z(n16423) );
  XOR2_X1 U24958 ( .A1(n535), .A2(n6597), .Z(n45477) );
  NOR2_X2 U24966 ( .A1(n34306), .A2(n23470), .ZN(n62775) );
  NAND2_X2 U24968 ( .A1(n15882), .A2(n62776), .ZN(n11831) );
  NOR2_X2 U24972 ( .A1(n10577), .A2(n19481), .ZN(n62776) );
  NOR2_X1 U24976 ( .A1(n22293), .A2(n22294), .ZN(n22292) );
  NAND2_X1 U24977 ( .A1(n37327), .A2(n8010), .ZN(n37340) );
  NAND2_X2 U24982 ( .A1(n62777), .A2(n5020), .ZN(n19909) );
  INV_X2 U24984 ( .I(n55956), .ZN(n62777) );
  NAND2_X2 U24988 ( .A1(n61554), .A2(n20737), .ZN(n55956) );
  NOR2_X2 U24992 ( .A1(n43586), .A2(n43585), .ZN(n2691) );
  BUF_X4 U24995 ( .I(n8214), .Z(n64039) );
  XOR2_X1 U25002 ( .A1(n62778), .A2(n46093), .Z(n57899) );
  XOR2_X1 U25010 ( .A1(n59312), .A2(n46092), .Z(n62778) );
  OAI21_X1 U25023 ( .A1(n50804), .A2(n64772), .B(n50807), .ZN(n62779) );
  XOR2_X1 U25026 ( .A1(n63003), .A2(n15096), .Z(n3140) );
  AOI22_X2 U25046 ( .A1(n19077), .A2(n63830), .B1(n1585), .B2(n11782), .ZN(
        n55901) );
  XOR2_X1 U25047 ( .A1(n62780), .A2(n56322), .Z(Plaintext[153]) );
  NAND3_X1 U25049 ( .A1(n11915), .A2(n11919), .A3(n11918), .ZN(n62780) );
  AND2_X2 U25051 ( .A1(n19609), .A2(n33420), .Z(n21106) );
  XOR2_X1 U25053 ( .A1(n8105), .A2(n44116), .Z(n8104) );
  XOR2_X1 U25059 ( .A1(n25243), .A2(n59811), .Z(n8105) );
  INV_X2 U25067 ( .I(n45969), .ZN(n1475) );
  NAND2_X2 U25069 ( .A1(n3510), .A2(n19645), .ZN(n45969) );
  AOI21_X2 U25084 ( .A1(n40810), .A2(n65202), .B(n62781), .ZN(n40839) );
  NAND3_X2 U25085 ( .A1(n40808), .A2(n4367), .A3(n4366), .ZN(n62781) );
  NAND3_X2 U25088 ( .A1(n60142), .A2(n20918), .A3(n30174), .ZN(n30168) );
  NAND2_X2 U25092 ( .A1(n24333), .A2(n17629), .ZN(n24332) );
  NOR2_X2 U25097 ( .A1(n618), .A2(n4095), .ZN(n24333) );
  NOR3_X2 U25104 ( .A1(n62783), .A2(n37962), .A3(n62782), .ZN(n21914) );
  INV_X4 U25106 ( .I(n24210), .ZN(n49109) );
  INV_X4 U25114 ( .I(n5536), .ZN(n10237) );
  AND2_X1 U25115 ( .A1(n41882), .A2(n62785), .Z(n39793) );
  NOR2_X1 U25128 ( .A1(n62786), .A2(n19816), .ZN(n65249) );
  NAND2_X1 U25134 ( .A1(n14728), .A2(n7802), .ZN(n62786) );
  NAND2_X2 U25135 ( .A1(n1782), .A2(n10413), .ZN(n7831) );
  NOR3_X2 U25140 ( .A1(n49832), .A2(n48303), .A3(n23238), .ZN(n64303) );
  XOR2_X1 U25141 ( .A1(n20059), .A2(n64938), .Z(n64131) );
  AOI21_X1 U25145 ( .A1(n56440), .A2(n61368), .B(n56439), .ZN(n63551) );
  NOR3_X1 U25154 ( .A1(n50208), .A2(n50210), .A3(n50209), .ZN(n64981) );
  XOR2_X1 U25155 ( .A1(n59435), .A2(n62787), .Z(n64822) );
  INV_X1 U25156 ( .I(n52408), .ZN(n62787) );
  XOR2_X1 U25159 ( .A1(n32176), .A2(n62831), .Z(n8456) );
  XOR2_X1 U25160 ( .A1(n12504), .A2(n32666), .Z(n32176) );
  NAND3_X2 U25162 ( .A1(n49382), .A2(n49395), .A3(n15753), .ZN(n49322) );
  BUF_X2 U25174 ( .I(n9046), .Z(n62788) );
  INV_X2 U25180 ( .I(n56788), .ZN(n56795) );
  NAND3_X2 U25181 ( .A1(n48149), .A2(n60138), .A3(n62880), .ZN(n48542) );
  XOR2_X1 U25193 ( .A1(n62790), .A2(n45385), .Z(n43748) );
  XOR2_X1 U25197 ( .A1(n43746), .A2(n43745), .Z(n62790) );
  XOR2_X1 U25202 ( .A1(n62791), .A2(n12372), .Z(n12371) );
  XOR2_X1 U25206 ( .A1(n12373), .A2(n60576), .Z(n62791) );
  XOR2_X1 U25209 ( .A1(n3609), .A2(n62792), .Z(n63047) );
  NAND3_X1 U25210 ( .A1(n12359), .A2(n45931), .A3(n45930), .ZN(n45934) );
  INV_X4 U25216 ( .I(n344), .ZN(n47301) );
  NAND2_X1 U25219 ( .A1(n54792), .A2(n63708), .ZN(n63707) );
  XOR2_X1 U25221 ( .A1(n52603), .A2(n5693), .Z(n4041) );
  XOR2_X1 U25222 ( .A1(n26035), .A2(n8562), .Z(n52603) );
  AOI21_X1 U25223 ( .A1(n63542), .A2(n48716), .B(n18608), .ZN(n15131) );
  NAND2_X2 U25228 ( .A1(n39987), .A2(n38758), .ZN(n41473) );
  XOR2_X1 U25229 ( .A1(n20469), .A2(n9108), .Z(n144) );
  NAND3_X1 U25230 ( .A1(n28071), .A2(n28072), .A3(n27044), .ZN(n27045) );
  NAND2_X1 U25235 ( .A1(n41212), .A2(n41210), .ZN(n38939) );
  BUF_X2 U25237 ( .I(n43750), .Z(n47735) );
  NOR2_X1 U25238 ( .A1(n17893), .A2(n26162), .ZN(n56466) );
  NAND2_X2 U25240 ( .A1(n1366), .A2(n9311), .ZN(n17893) );
  NAND2_X2 U25248 ( .A1(n47314), .A2(n10357), .ZN(n2944) );
  NOR2_X2 U25249 ( .A1(n29725), .A2(n22748), .ZN(n29878) );
  NAND2_X2 U25255 ( .A1(n1865), .A2(n13174), .ZN(n29725) );
  INV_X2 U25261 ( .I(n23453), .ZN(n54558) );
  BUF_X2 U25262 ( .I(n25125), .Z(n62794) );
  NAND2_X2 U25265 ( .A1(n1659), .A2(n64634), .ZN(n3221) );
  AND2_X1 U25272 ( .A1(n62999), .A2(n30786), .Z(n30769) );
  BUF_X2 U25274 ( .I(n65222), .Z(n62795) );
  XOR2_X1 U25277 ( .A1(n23222), .A2(n18478), .Z(n6596) );
  NAND3_X2 U25286 ( .A1(n15778), .A2(n18474), .A3(n16187), .ZN(n23222) );
  INV_X2 U25287 ( .I(n62796), .ZN(n18068) );
  XOR2_X1 U25288 ( .A1(n18315), .A2(n37612), .Z(n62796) );
  INV_X2 U25297 ( .I(n20713), .ZN(n42091) );
  NAND3_X2 U25299 ( .A1(n6452), .A2(n6453), .A3(n6451), .ZN(n20713) );
  XOR2_X1 U25301 ( .A1(n22435), .A2(n59250), .Z(n10767) );
  NOR2_X2 U25302 ( .A1(n8394), .A2(n11243), .ZN(n62797) );
  XOR2_X1 U25304 ( .A1(n62798), .A2(n51627), .Z(n65212) );
  XOR2_X1 U25315 ( .A1(n62799), .A2(n24023), .Z(n32184) );
  XOR2_X1 U25322 ( .A1(n2192), .A2(n37761), .Z(n2788) );
  NAND2_X2 U25325 ( .A1(n58030), .A2(n49259), .ZN(n63024) );
  NOR3_X2 U25339 ( .A1(n7553), .A2(n7554), .A3(n19831), .ZN(n58030) );
  NOR2_X2 U25343 ( .A1(n43610), .A2(n42159), .ZN(n21861) );
  NOR2_X2 U25346 ( .A1(n23626), .A2(n60891), .ZN(n35581) );
  NAND2_X2 U25352 ( .A1(n64978), .A2(n53845), .ZN(n54489) );
  NAND3_X1 U25358 ( .A1(n22414), .A2(n56900), .A3(n56899), .ZN(n62805) );
  INV_X2 U25361 ( .I(n24021), .ZN(n58201) );
  NAND3_X2 U25362 ( .A1(n64569), .A2(n58734), .A3(n15494), .ZN(n24021) );
  XOR2_X1 U25366 ( .A1(n22277), .A2(n38848), .Z(n38849) );
  NAND2_X2 U25370 ( .A1(n32451), .A2(n7714), .ZN(n22277) );
  XOR2_X1 U25372 ( .A1(n36298), .A2(n18072), .Z(n18073) );
  XOR2_X1 U25374 ( .A1(n62801), .A2(n39494), .Z(n18316) );
  XOR2_X1 U25375 ( .A1(n37609), .A2(n37698), .Z(n62801) );
  OAI22_X1 U25376 ( .A1(n1070), .A2(n1388), .B1(n1267), .B2(n18361), .ZN(
        n44205) );
  AOI21_X2 U25379 ( .A1(n11312), .A2(n37361), .B(n11311), .ZN(n466) );
  XOR2_X1 U25383 ( .A1(n3244), .A2(n62802), .Z(n4148) );
  XOR2_X1 U25386 ( .A1(n20022), .A2(n19821), .Z(n62802) );
  NOR2_X2 U25388 ( .A1(n57830), .A2(n19231), .ZN(n1903) );
  NOR3_X1 U25389 ( .A1(n7748), .A2(n22541), .A3(n26665), .ZN(n26502) );
  BUF_X2 U25398 ( .I(n1714), .Z(n61171) );
  XNOR2_X1 U25403 ( .A1(n6590), .A2(n65254), .ZN(n15242) );
  XOR2_X1 U25405 ( .A1(n6593), .A2(n63496), .Z(n65254) );
  NOR2_X2 U25407 ( .A1(n15034), .A2(n1531), .ZN(n64753) );
  AOI21_X2 U25416 ( .A1(n57332), .A2(n59660), .B(n62803), .ZN(n7226) );
  NAND2_X2 U25421 ( .A1(n58195), .A2(n12168), .ZN(n62803) );
  AND2_X2 U25429 ( .A1(n54112), .A2(n10969), .Z(n53876) );
  XOR2_X1 U25437 ( .A1(n44905), .A2(n25472), .Z(n25471) );
  NAND2_X2 U25440 ( .A1(n11600), .A2(n12341), .ZN(n11700) );
  NOR2_X2 U25442 ( .A1(n62804), .A2(n61289), .ZN(n11600) );
  OR2_X1 U25445 ( .A1(n11592), .A2(n19051), .Z(n62804) );
  NAND2_X2 U25448 ( .A1(n49678), .A2(n11155), .ZN(n48014) );
  NAND3_X2 U25452 ( .A1(n58645), .A2(n5463), .A3(n17906), .ZN(n49678) );
  XOR2_X1 U25454 ( .A1(n62805), .A2(n56901), .Z(Plaintext[179]) );
  INV_X2 U25455 ( .I(n53118), .ZN(n53083) );
  NAND2_X2 U25465 ( .A1(n13421), .A2(n13230), .ZN(n53118) );
  NAND4_X1 U25480 ( .A1(n63438), .A2(n3085), .A3(n8640), .A4(n60202), .ZN(
        n62806) );
  NOR2_X2 U25488 ( .A1(n24690), .A2(n62807), .ZN(n25953) );
  XOR2_X1 U25489 ( .A1(n18342), .A2(n24065), .Z(n8556) );
  BUF_X2 U25495 ( .I(n51112), .Z(n62808) );
  AND2_X1 U25496 ( .A1(n4723), .A2(n25534), .Z(n42400) );
  NOR2_X2 U25497 ( .A1(n15105), .A2(n62809), .ZN(n15726) );
  NAND3_X2 U25506 ( .A1(n59317), .A2(n59316), .A3(n27994), .ZN(n62809) );
  NAND2_X1 U25507 ( .A1(n7474), .A2(n12876), .ZN(n62812) );
  NAND2_X2 U25512 ( .A1(n62810), .A2(n16698), .ZN(n35882) );
  NOR4_X2 U25513 ( .A1(n60165), .A2(n13251), .A3(n13254), .A4(n60164), .ZN(
        n62810) );
  NOR2_X1 U25518 ( .A1(n63156), .A2(n63154), .ZN(n25767) );
  BUF_X2 U25521 ( .I(n22217), .Z(n4232) );
  NOR2_X1 U25526 ( .A1(n4723), .A2(n19248), .ZN(n41691) );
  NAND2_X1 U25528 ( .A1(n12552), .A2(n56570), .ZN(n64124) );
  NOR2_X2 U25529 ( .A1(n62812), .A2(n38044), .ZN(n21055) );
  AND2_X1 U25542 ( .A1(n1405), .A2(n40713), .Z(n39022) );
  XOR2_X1 U25546 ( .A1(n62813), .A2(n12593), .Z(n4673) );
  XOR2_X1 U25548 ( .A1(n7102), .A2(n4936), .Z(n62813) );
  XOR2_X1 U25551 ( .A1(n59832), .A2(n24776), .Z(n26086) );
  NAND2_X2 U25554 ( .A1(n6411), .A2(n61742), .ZN(n48792) );
  NAND2_X2 U25555 ( .A1(n52723), .A2(n62814), .ZN(n56891) );
  NOR3_X2 U25558 ( .A1(n52715), .A2(n52714), .A3(n52713), .ZN(n62814) );
  NAND2_X2 U25561 ( .A1(n61147), .A2(n53859), .ZN(n9514) );
  XOR2_X1 U25569 ( .A1(n25957), .A2(n3568), .Z(n60261) );
  NAND3_X2 U25571 ( .A1(n62815), .A2(n55041), .A3(n55029), .ZN(n8413) );
  NAND2_X1 U25573 ( .A1(n55033), .A2(n55032), .ZN(n62815) );
  NAND4_X2 U25575 ( .A1(n19738), .A2(n19737), .A3(n45211), .A4(n62817), .ZN(
        n45229) );
  AOI22_X1 U25588 ( .A1(n1663), .A2(n47236), .B1(n47237), .B2(n1069), .ZN(
        n62817) );
  NAND2_X2 U25591 ( .A1(n60129), .A2(n56629), .ZN(n56211) );
  NOR2_X1 U25596 ( .A1(n12760), .A2(n43612), .ZN(n11800) );
  NAND2_X2 U25597 ( .A1(n48068), .A2(n57666), .ZN(n50752) );
  OAI22_X1 U25599 ( .A1(n5713), .A2(n9395), .B1(n49410), .B2(n9164), .ZN(
        n49262) );
  NAND2_X1 U25610 ( .A1(n33415), .A2(n35606), .ZN(n63162) );
  XOR2_X1 U25611 ( .A1(n24730), .A2(n1313), .Z(n8464) );
  NAND4_X1 U25615 ( .A1(n53362), .A2(n9731), .A3(n53334), .A4(n63931), .ZN(
        n52809) );
  NAND2_X2 U25617 ( .A1(n23874), .A2(n52808), .ZN(n63931) );
  NAND2_X2 U25619 ( .A1(n4343), .A2(n44578), .ZN(n3503) );
  NOR2_X2 U25622 ( .A1(n4347), .A2(n4346), .ZN(n4343) );
  OR2_X1 U25625 ( .A1(n5206), .A2(n24233), .Z(n24946) );
  OAI21_X2 U25633 ( .A1(n10167), .A2(n61848), .B(n25417), .ZN(n43319) );
  NOR3_X2 U25649 ( .A1(n9260), .A2(n9261), .A3(n26677), .ZN(n9411) );
  NAND3_X2 U25658 ( .A1(n36353), .A2(n59236), .A3(n36354), .ZN(n39592) );
  NAND3_X2 U25660 ( .A1(n59815), .A2(n33443), .A3(n34649), .ZN(n5937) );
  NAND2_X1 U25676 ( .A1(n21392), .A2(n62820), .ZN(n21391) );
  OR2_X1 U25680 ( .A1(n52949), .A2(n21393), .Z(n62820) );
  NAND3_X2 U25687 ( .A1(n11072), .A2(n35960), .A3(n11493), .ZN(n23949) );
  OAI21_X2 U25689 ( .A1(n2096), .A2(n2095), .B(n7933), .ZN(n11072) );
  OR2_X2 U25702 ( .A1(n33098), .A2(n16857), .Z(n16939) );
  NOR2_X2 U25708 ( .A1(n5959), .A2(n36939), .ZN(n5958) );
  NOR3_X2 U25711 ( .A1(n1559), .A2(n30195), .A3(n30183), .ZN(n29736) );
  NAND2_X1 U25712 ( .A1(n61684), .A2(n55942), .ZN(n63433) );
  XOR2_X1 U25713 ( .A1(n64398), .A2(n2127), .Z(n2126) );
  XOR2_X1 U25715 ( .A1(n3291), .A2(n59648), .Z(n5101) );
  AND2_X1 U25716 ( .A1(n36022), .A2(n36020), .Z(n36027) );
  NAND2_X2 U25717 ( .A1(n56600), .A2(n52683), .ZN(n6991) );
  XOR2_X1 U25719 ( .A1(n62821), .A2(n10688), .Z(n105) );
  NOR2_X2 U25720 ( .A1(n64410), .A2(n35899), .ZN(n35897) );
  NAND2_X2 U25723 ( .A1(n4744), .A2(n30069), .ZN(n32467) );
  NOR2_X2 U25724 ( .A1(n61176), .A2(n62823), .ZN(n50361) );
  OR2_X2 U25729 ( .A1(n40294), .A2(n23477), .Z(n40296) );
  XOR2_X1 U25737 ( .A1(n62825), .A2(n23389), .Z(n31463) );
  XOR2_X1 U25741 ( .A1(n31460), .A2(n19886), .Z(n62825) );
  XOR2_X1 U25743 ( .A1(n62826), .A2(n32544), .Z(n12078) );
  XOR2_X1 U25756 ( .A1(n23706), .A2(n28784), .Z(n62826) );
  NAND3_X2 U25758 ( .A1(n62827), .A2(n8315), .A3(n8314), .ZN(n543) );
  XOR2_X1 U25762 ( .A1(n23726), .A2(n19204), .Z(n65152) );
  NAND3_X2 U25768 ( .A1(n14283), .A2(n15917), .A3(n14281), .ZN(n17409) );
  NAND2_X2 U25770 ( .A1(n12410), .A2(n6748), .ZN(n40987) );
  CLKBUF_X4 U25772 ( .I(n8733), .Z(n4428) );
  NOR3_X2 U25775 ( .A1(n36255), .A2(n62829), .A3(n62828), .ZN(n2684) );
  NOR2_X1 U25784 ( .A1(n36252), .A2(n62794), .ZN(n62828) );
  NOR2_X1 U25794 ( .A1(n36253), .A2(n10067), .ZN(n62829) );
  NAND2_X2 U25797 ( .A1(n61706), .A2(n1226), .ZN(n8853) );
  INV_X2 U25798 ( .I(n47252), .ZN(n59419) );
  NAND2_X1 U25802 ( .A1(n62830), .A2(n56313), .ZN(n56292) );
  XOR2_X1 U25805 ( .A1(n23318), .A2(n11841), .Z(n62830) );
  XOR2_X1 U25806 ( .A1(n31565), .A2(n61946), .Z(n62831) );
  NOR2_X2 U25808 ( .A1(n6284), .A2(n62832), .ZN(n20811) );
  NAND3_X2 U25813 ( .A1(n6282), .A2(n6280), .A3(n6281), .ZN(n62832) );
  NAND3_X2 U25814 ( .A1(n5013), .A2(n34650), .A3(n34651), .ZN(n34695) );
  BUF_X2 U25818 ( .I(n11912), .Z(n23122) );
  OAI21_X1 U25824 ( .A1(n7347), .A2(n7346), .B(n55016), .ZN(n63516) );
  NOR2_X1 U25830 ( .A1(n58199), .A2(n2626), .ZN(n2623) );
  NAND2_X1 U25833 ( .A1(n63184), .A2(n545), .ZN(n60230) );
  NOR2_X1 U25836 ( .A1(n674), .A2(n55015), .ZN(n4087) );
  OR2_X2 U25842 ( .A1(n14039), .A2(n14733), .Z(n65052) );
  NOR3_X2 U25843 ( .A1(n63122), .A2(n21635), .A3(n58083), .ZN(n54239) );
  NOR2_X2 U25844 ( .A1(n62833), .A2(n6053), .ZN(n35140) );
  NAND4_X2 U25845 ( .A1(n12820), .A2(n33679), .A3(n12821), .A4(n33678), .ZN(
        n62833) );
  NOR2_X1 U25846 ( .A1(n62891), .A2(n21491), .ZN(n317) );
  OR2_X2 U25848 ( .A1(n22283), .A2(n16617), .Z(n48249) );
  XOR2_X1 U25850 ( .A1(n62834), .A2(n45877), .Z(n21022) );
  NOR3_X2 U25854 ( .A1(n51905), .A2(n56229), .A3(n56436), .ZN(n25173) );
  XOR2_X1 U25860 ( .A1(n12028), .A2(n12027), .Z(n51905) );
  XOR2_X1 U25862 ( .A1(n62835), .A2(n5247), .Z(n31563) );
  XOR2_X1 U25864 ( .A1(n23690), .A2(n23726), .Z(n62835) );
  XOR2_X1 U25867 ( .A1(n62836), .A2(n2741), .Z(n14878) );
  XOR2_X1 U25881 ( .A1(n37301), .A2(n25965), .Z(n62836) );
  BUF_X2 U25885 ( .I(n38405), .Z(n41158) );
  XOR2_X1 U25888 ( .A1(n62837), .A2(n46386), .Z(n17518) );
  XOR2_X1 U25893 ( .A1(n43763), .A2(n65170), .Z(n62837) );
  INV_X1 U25894 ( .I(n3804), .ZN(n64240) );
  NOR3_X2 U25895 ( .A1(n12220), .A2(n13490), .A3(n60856), .ZN(n6298) );
  INV_X1 U25896 ( .I(n63507), .ZN(n15108) );
  OAI21_X1 U25899 ( .A1(n62838), .A2(n14501), .B(n6311), .ZN(n20414) );
  NOR2_X1 U25903 ( .A1(n6510), .A2(n62768), .ZN(n62838) );
  OAI21_X2 U25907 ( .A1(n58074), .A2(n23778), .B(n58073), .ZN(n37956) );
  OR3_X1 U25908 ( .A1(n53876), .A2(n54107), .A3(n2997), .Z(n12310) );
  OR2_X2 U25910 ( .A1(n6728), .A2(n8170), .Z(n59216) );
  BUF_X4 U25912 ( .I(n46412), .Z(n48135) );
  NAND2_X1 U25915 ( .A1(n62839), .A2(n34014), .ZN(n22495) );
  NOR2_X1 U25917 ( .A1(n4851), .A2(n34632), .ZN(n62839) );
  NAND2_X2 U25919 ( .A1(n25716), .A2(n62840), .ZN(n21470) );
  NAND2_X2 U25920 ( .A1(n24520), .A2(n54259), .ZN(n54213) );
  OR2_X1 U25921 ( .A1(n55644), .A2(n55641), .Z(n63382) );
  AOI21_X1 U25922 ( .A1(n9751), .A2(n8340), .B(n11076), .ZN(n64959) );
  INV_X2 U25930 ( .I(n28409), .ZN(n11076) );
  NOR2_X2 U25932 ( .A1(n58792), .A2(n28004), .ZN(n28409) );
  XOR2_X1 U25933 ( .A1(n62841), .A2(n58432), .Z(n63886) );
  XOR2_X1 U25935 ( .A1(n64511), .A2(n32715), .Z(n62841) );
  NAND4_X2 U25939 ( .A1(n56551), .A2(n62842), .A3(n56549), .A4(n56550), .ZN(
        n56552) );
  AND2_X1 U25940 ( .A1(n14762), .A2(n14761), .Z(n62842) );
  NAND3_X1 U25941 ( .A1(n64665), .A2(n54077), .A3(n54075), .ZN(n62843) );
  XOR2_X1 U25942 ( .A1(n64955), .A2(n24329), .Z(n50716) );
  XOR2_X1 U25945 ( .A1(n16820), .A2(n31345), .Z(n16821) );
  NAND2_X2 U25956 ( .A1(n63313), .A2(n62844), .ZN(n20261) );
  NAND3_X2 U25962 ( .A1(n51568), .A2(n12142), .A3(n62845), .ZN(n5893) );
  NAND3_X2 U25970 ( .A1(n56766), .A2(n65064), .A3(n57212), .ZN(n62845) );
  BUF_X2 U25978 ( .I(n56629), .Z(n62846) );
  BUF_X4 U25980 ( .I(n43898), .Z(n64323) );
  NOR2_X2 U25983 ( .A1(n4724), .A2(n4719), .ZN(n19043) );
  NAND2_X2 U25985 ( .A1(n56803), .A2(n62120), .ZN(n56816) );
  OR2_X1 U25986 ( .A1(n20045), .A2(n55908), .Z(n8969) );
  XOR2_X1 U25990 ( .A1(n1326), .A2(n55909), .Z(n20045) );
  NAND2_X2 U25991 ( .A1(n44786), .A2(n62848), .ZN(n44788) );
  AOI22_X2 U25994 ( .A1(n44777), .A2(n44778), .B1(n44775), .B2(n44776), .ZN(
        n62848) );
  XOR2_X1 U25995 ( .A1(n12918), .A2(n62849), .Z(n3248) );
  XOR2_X1 U25997 ( .A1(n17448), .A2(n12919), .Z(n62849) );
  XNOR2_X1 U26003 ( .A1(n46432), .A2(n45145), .ZN(n25209) );
  NAND3_X2 U26004 ( .A1(n33796), .A2(n33804), .A3(n33803), .ZN(n20254) );
  NOR2_X2 U26005 ( .A1(n21667), .A2(n24179), .ZN(n6563) );
  INV_X4 U26008 ( .I(n1221), .ZN(n62995) );
  INV_X1 U26009 ( .I(n16821), .ZN(n62850) );
  NOR2_X2 U26011 ( .A1(n47554), .A2(n49195), .ZN(n49521) );
  XOR2_X1 U26013 ( .A1(n21580), .A2(n46527), .Z(n60156) );
  NOR2_X2 U26014 ( .A1(n50309), .A2(n3055), .ZN(n4212) );
  INV_X2 U26017 ( .I(n26169), .ZN(n50309) );
  NAND3_X2 U26023 ( .A1(n59980), .A2(n7953), .A3(n5917), .ZN(n26169) );
  NOR2_X2 U26024 ( .A1(n62851), .A2(n3811), .ZN(n25856) );
  NAND3_X2 U26028 ( .A1(n63607), .A2(n3817), .A3(n3818), .ZN(n62851) );
  NAND3_X2 U26046 ( .A1(n40249), .A2(n40248), .A3(n40464), .ZN(n40481) );
  NAND2_X2 U26050 ( .A1(n6052), .A2(n33709), .ZN(n35354) );
  NOR3_X2 U26051 ( .A1(n41706), .A2(n3786), .A3(n22186), .ZN(n59896) );
  AND2_X1 U26059 ( .A1(n28275), .A2(n28281), .Z(n8776) );
  XOR2_X1 U26061 ( .A1(n7187), .A2(n24884), .Z(n42755) );
  OR2_X1 U26069 ( .A1(n36561), .A2(n9273), .Z(n61298) );
  NOR2_X2 U26070 ( .A1(n8356), .A2(n22785), .ZN(n36561) );
  NAND2_X2 U26076 ( .A1(n13745), .A2(n35974), .ZN(n35138) );
  XOR2_X1 U26082 ( .A1(n2452), .A2(n44356), .Z(n19411) );
  NOR2_X2 U26087 ( .A1(n2456), .A2(n2455), .ZN(n2452) );
  NAND4_X1 U26089 ( .A1(n9089), .A2(n54299), .A3(n54487), .A4(n54970), .ZN(
        n54303) );
  NAND3_X1 U26090 ( .A1(n32072), .A2(n10227), .A3(n35811), .ZN(n32073) );
  XOR2_X1 U26091 ( .A1(n2952), .A2(n21172), .Z(n2954) );
  INV_X4 U26093 ( .I(n62853), .ZN(n209) );
  NAND2_X2 U26103 ( .A1(n16617), .A2(n16616), .ZN(n62853) );
  NOR2_X1 U26110 ( .A1(n35669), .A2(n35668), .ZN(n62854) );
  XOR2_X1 U26113 ( .A1(n25995), .A2(n39286), .Z(n38750) );
  NOR2_X2 U26117 ( .A1(n9829), .A2(n26189), .ZN(n62855) );
  NAND2_X2 U26118 ( .A1(n62858), .A2(n36412), .ZN(n36403) );
  NAND2_X2 U26121 ( .A1(n16968), .A2(n36193), .ZN(n3076) );
  NOR2_X2 U26122 ( .A1(n63199), .A2(n63195), .ZN(n62903) );
  NOR2_X2 U26124 ( .A1(n7147), .A2(n60279), .ZN(n62859) );
  OAI22_X2 U26130 ( .A1(n13753), .A2(n62860), .B1(n15120), .B2(n42418), .ZN(
        n15119) );
  BUF_X2 U26135 ( .I(n8298), .Z(n62861) );
  XOR2_X1 U26136 ( .A1(n2153), .A2(n51028), .Z(n6738) );
  NAND3_X2 U26137 ( .A1(n33581), .A2(n33580), .A3(n33582), .ZN(n36410) );
  NAND2_X2 U26142 ( .A1(n47310), .A2(n47329), .ZN(n47327) );
  NOR2_X2 U26144 ( .A1(n45076), .A2(n47307), .ZN(n47310) );
  NAND3_X2 U26150 ( .A1(n37218), .A2(n36986), .A3(n37224), .ZN(n36991) );
  NAND2_X2 U26154 ( .A1(n28093), .A2(n17550), .ZN(n29416) );
  NAND2_X2 U26160 ( .A1(n19649), .A2(n27307), .ZN(n28093) );
  XOR2_X1 U26163 ( .A1(n13964), .A2(n62862), .Z(n24378) );
  XOR2_X1 U26164 ( .A1(n33052), .A2(n26165), .Z(n62862) );
  XOR2_X1 U26167 ( .A1(n62863), .A2(n16511), .Z(n39453) );
  XOR2_X1 U26171 ( .A1(n39270), .A2(n15699), .Z(n62863) );
  INV_X1 U26173 ( .I(n64526), .ZN(n63225) );
  NAND2_X1 U26174 ( .A1(n21570), .A2(n57120), .ZN(n57159) );
  NOR2_X2 U26175 ( .A1(n59180), .A2(n63039), .ZN(n56350) );
  NAND2_X2 U26185 ( .A1(n64652), .A2(n10680), .ZN(n59445) );
  XOR2_X1 U26189 ( .A1(n3717), .A2(n8353), .Z(n63538) );
  OAI21_X2 U26195 ( .A1(n62865), .A2(n23623), .B(n8799), .ZN(n2235) );
  NAND2_X1 U26205 ( .A1(n23622), .A2(n64724), .ZN(n62865) );
  XOR2_X1 U26225 ( .A1(n62866), .A2(n51191), .Z(n50782) );
  XOR2_X1 U26234 ( .A1(n9230), .A2(n9236), .Z(n62866) );
  BUF_X4 U26235 ( .I(n33215), .Z(n35834) );
  XOR2_X1 U26238 ( .A1(n15640), .A2(n16132), .Z(n33116) );
  AND3_X2 U26244 ( .A1(n24141), .A2(n55918), .A3(n55919), .Z(n63591) );
  XOR2_X1 U26253 ( .A1(n62867), .A2(n758), .Z(n9216) );
  XOR2_X1 U26258 ( .A1(n36324), .A2(n64427), .Z(n62867) );
  NAND2_X1 U26259 ( .A1(n60430), .A2(n60429), .ZN(n60004) );
  INV_X1 U26260 ( .I(n101), .ZN(n62868) );
  NOR3_X1 U26262 ( .A1(n39415), .A2(n60113), .A3(n2159), .ZN(n39416) );
  NAND3_X2 U26264 ( .A1(n44289), .A2(n60308), .A3(n44287), .ZN(n48322) );
  INV_X2 U26268 ( .I(n24425), .ZN(n43701) );
  XOR2_X1 U26279 ( .A1(n15722), .A2(n14538), .Z(n8588) );
  INV_X2 U26285 ( .I(n62869), .ZN(n57172) );
  NOR2_X2 U26288 ( .A1(n21699), .A2(n25428), .ZN(n62869) );
  NOR2_X1 U26297 ( .A1(n48488), .A2(n48185), .ZN(n64138) );
  OAI21_X2 U26306 ( .A1(n29236), .A2(n29241), .B(n30815), .ZN(n29928) );
  BUF_X4 U26309 ( .I(n23284), .Z(n5323) );
  NAND2_X1 U26310 ( .A1(n40900), .A2(n40901), .ZN(n62925) );
  NOR2_X1 U26311 ( .A1(n6736), .A2(n16083), .ZN(n6735) );
  NAND3_X1 U26313 ( .A1(n54562), .A2(n62629), .A3(n54570), .ZN(n54528) );
  NAND3_X1 U26314 ( .A1(n50099), .A2(n5282), .A3(n50376), .ZN(n50100) );
  INV_X2 U26315 ( .I(n62871), .ZN(n19142) );
  NAND2_X2 U26317 ( .A1(n18100), .A2(n19160), .ZN(n62871) );
  NAND2_X2 U26321 ( .A1(n60321), .A2(n62872), .ZN(n4002) );
  AOI22_X2 U26324 ( .A1(n59608), .A2(n63583), .B1(n7103), .B2(n36550), .ZN(
        n62872) );
  XOR2_X1 U26333 ( .A1(n43961), .A2(n12654), .Z(n64422) );
  XOR2_X1 U26334 ( .A1(n18993), .A2(n22702), .Z(n43961) );
  INV_X2 U26337 ( .I(n37034), .ZN(n14138) );
  XOR2_X1 U26339 ( .A1(n6906), .A2(n62874), .Z(n13752) );
  XOR2_X1 U26342 ( .A1(n18170), .A2(n62875), .Z(n62874) );
  NOR2_X1 U26344 ( .A1(n26015), .A2(n63473), .ZN(n54764) );
  NAND2_X2 U26358 ( .A1(n18463), .A2(n54695), .ZN(n63473) );
  INV_X2 U26359 ( .I(n18410), .ZN(n64115) );
  NOR2_X2 U26362 ( .A1(n17268), .A2(n29430), .ZN(n13629) );
  AND2_X1 U26366 ( .A1(n41098), .A2(n41097), .Z(n15944) );
  XOR2_X1 U26369 ( .A1(n23619), .A2(n39365), .Z(n3346) );
  NAND3_X2 U26373 ( .A1(n8174), .A2(n8173), .A3(n35948), .ZN(n39365) );
  NAND3_X2 U26374 ( .A1(n12331), .A2(n48005), .A3(n62876), .ZN(n9876) );
  INV_X2 U26382 ( .I(n62877), .ZN(n57405) );
  XOR2_X1 U26383 ( .A1(n2842), .A2(n24908), .Z(n62877) );
  INV_X2 U26384 ( .I(n11620), .ZN(n2147) );
  NAND2_X2 U26386 ( .A1(n348), .A2(n73), .ZN(n11620) );
  NOR2_X2 U26388 ( .A1(n36247), .A2(n34886), .ZN(n12830) );
  NAND3_X2 U26390 ( .A1(n33401), .A2(n33402), .A3(n25230), .ZN(n34886) );
  XOR2_X1 U26391 ( .A1(n10684), .A2(n8506), .Z(n31708) );
  XOR2_X1 U26397 ( .A1(n38921), .A2(n24147), .Z(n38541) );
  XOR2_X1 U26401 ( .A1(n39230), .A2(n24151), .Z(n38921) );
  NAND3_X2 U26402 ( .A1(n49511), .A2(n49525), .A3(n49195), .ZN(n16829) );
  NAND3_X2 U26403 ( .A1(n46880), .A2(n61278), .A3(n46879), .ZN(n48428) );
  NAND4_X2 U26411 ( .A1(n59424), .A2(n56642), .A3(n56640), .A4(n56641), .ZN(
        n56644) );
  XOR2_X1 U26413 ( .A1(n1549), .A2(n32620), .Z(n3519) );
  NAND3_X2 U26416 ( .A1(n15062), .A2(n62879), .A3(n15174), .ZN(n19155) );
  NAND2_X2 U26417 ( .A1(n30537), .A2(n24298), .ZN(n30540) );
  NAND2_X2 U26419 ( .A1(n3065), .A2(n10960), .ZN(n16030) );
  BUF_X2 U26426 ( .I(n48544), .Z(n62880) );
  XOR2_X1 U26432 ( .A1(n11501), .A2(n17863), .Z(n14500) );
  NAND3_X2 U26433 ( .A1(n10040), .A2(n3616), .A3(n62881), .ZN(n56266) );
  NOR2_X2 U26441 ( .A1(n24944), .A2(n56268), .ZN(n62881) );
  INV_X4 U26442 ( .I(n21104), .ZN(n1413) );
  NOR2_X2 U26443 ( .A1(n62882), .A2(n4585), .ZN(n63050) );
  OR2_X1 U26445 ( .A1(n30445), .A2(n30446), .Z(n62882) );
  XOR2_X1 U26450 ( .A1(n62883), .A2(n31941), .Z(n31945) );
  XOR2_X1 U26451 ( .A1(n32013), .A2(n32661), .Z(n62883) );
  BUF_X4 U26453 ( .I(n21830), .Z(n21829) );
  NAND3_X1 U26457 ( .A1(n62887), .A2(n57069), .A3(n62884), .ZN(n57078) );
  INV_X2 U26459 ( .I(n18219), .ZN(n62886) );
  NAND2_X1 U26463 ( .A1(n14091), .A2(n57067), .ZN(n62887) );
  NAND2_X1 U26464 ( .A1(n2287), .A2(n35735), .ZN(n34413) );
  INV_X1 U26469 ( .I(n56891), .ZN(n56863) );
  NAND3_X2 U26477 ( .A1(n62888), .A2(n52496), .A3(n52495), .ZN(n52648) );
  NAND3_X1 U26478 ( .A1(n21391), .A2(n21394), .A3(n55442), .ZN(n62888) );
  NOR3_X2 U26483 ( .A1(n52804), .A2(n52805), .A3(n52803), .ZN(n52794) );
  NOR4_X2 U26500 ( .A1(n61709), .A2(n42898), .A3(n42895), .A4(n42896), .ZN(
        n58918) );
  OR2_X2 U26501 ( .A1(n36020), .A2(n18385), .Z(n35571) );
  XOR2_X1 U26515 ( .A1(n12240), .A2(n62889), .Z(n2290) );
  XOR2_X1 U26520 ( .A1(n12243), .A2(n33870), .Z(n62889) );
  NAND2_X1 U26522 ( .A1(n35578), .A2(n35577), .ZN(n62917) );
  BUF_X4 U26526 ( .I(n56891), .Z(n21879) );
  NAND2_X2 U26527 ( .A1(n26017), .A2(n62890), .ZN(n4743) );
  NAND3_X2 U26528 ( .A1(n26019), .A2(n64428), .A3(n26016), .ZN(n62890) );
  INV_X2 U26540 ( .I(n52409), .ZN(n4513) );
  NAND3_X2 U26543 ( .A1(n48015), .A2(n48016), .A3(n48017), .ZN(n52409) );
  NOR2_X2 U26548 ( .A1(n20996), .A2(n3112), .ZN(n8135) );
  BUF_X4 U26549 ( .I(n36338), .Z(n65234) );
  INV_X2 U26565 ( .I(n52648), .ZN(n55132) );
  NAND2_X1 U26580 ( .A1(n22063), .A2(n34677), .ZN(n34054) );
  NOR2_X2 U26582 ( .A1(n242), .A2(n30832), .ZN(n22063) );
  INV_X2 U26583 ( .I(n23163), .ZN(n21859) );
  XOR2_X1 U26584 ( .A1(n62893), .A2(n37516), .Z(n64299) );
  XOR2_X1 U26585 ( .A1(n62027), .A2(n2032), .Z(n62893) );
  XOR2_X1 U26586 ( .A1(n5101), .A2(n58660), .Z(n63377) );
  NAND2_X2 U26590 ( .A1(n62894), .A2(n14930), .ZN(n11977) );
  INV_X2 U26592 ( .I(n15790), .ZN(n62894) );
  OR2_X1 U26598 ( .A1(n57411), .A2(n28177), .Z(n62895) );
  NAND2_X2 U26600 ( .A1(n36471), .A2(n36584), .ZN(n36582) );
  NAND2_X2 U26603 ( .A1(n31261), .A2(n17978), .ZN(n65051) );
  XOR2_X1 U26604 ( .A1(n3290), .A2(n1050), .Z(n63015) );
  BUF_X2 U26608 ( .I(n46319), .Z(n10552) );
  INV_X2 U26609 ( .I(n61442), .ZN(n25210) );
  INV_X1 U26610 ( .I(n63594), .ZN(n42044) );
  OR2_X1 U26612 ( .A1(n63594), .A2(n61442), .Z(n42638) );
  INV_X2 U26619 ( .I(n62896), .ZN(n34238) );
  XNOR2_X1 U26622 ( .A1(n63383), .A2(n25307), .ZN(n62896) );
  NOR2_X2 U26623 ( .A1(n57685), .A2(n62897), .ZN(n64399) );
  NAND4_X2 U26624 ( .A1(n46472), .A2(n46471), .A3(n46470), .A4(n48480), .ZN(
        n62897) );
  NOR3_X2 U26625 ( .A1(n4166), .A2(n62898), .A3(n4165), .ZN(n16460) );
  AOI21_X2 U26628 ( .A1(n64034), .A2(n4169), .B(n25563), .ZN(n62898) );
  NOR2_X2 U26632 ( .A1(n56775), .A2(n56817), .ZN(n56814) );
  NAND2_X1 U26637 ( .A1(n25556), .A2(n62899), .ZN(n4334) );
  OAI21_X2 U26641 ( .A1(n62901), .A2(n62900), .B(n54344), .ZN(n10527) );
  NOR2_X1 U26642 ( .A1(n4835), .A2(n54340), .ZN(n62901) );
  NOR2_X1 U26645 ( .A1(n55392), .A2(n55391), .ZN(n60421) );
  OAI22_X1 U26649 ( .A1(n3413), .A2(n3414), .B1(n3412), .B2(n18377), .ZN(
        n62902) );
  XOR2_X1 U26651 ( .A1(n62904), .A2(n53772), .Z(Plaintext[42]) );
  NAND3_X1 U26656 ( .A1(n53771), .A2(n7486), .A3(n53770), .ZN(n62904) );
  NOR2_X1 U26657 ( .A1(n3765), .A2(n35947), .ZN(n63995) );
  NAND2_X1 U26658 ( .A1(n23452), .A2(n25386), .ZN(n61539) );
  NAND3_X2 U26659 ( .A1(n55962), .A2(n658), .A3(n55964), .ZN(n56000) );
  NAND2_X2 U26661 ( .A1(n30223), .A2(n23589), .ZN(n29884) );
  OAI22_X1 U26666 ( .A1(n35936), .A2(n16355), .B1(n16354), .B2(n35935), .ZN(
        n16353) );
  XOR2_X1 U26668 ( .A1(n11737), .A2(n12704), .Z(n12703) );
  AND2_X2 U26671 ( .A1(n61742), .A2(n62905), .Z(n49711) );
  NOR2_X2 U26676 ( .A1(n60239), .A2(n11927), .ZN(n58716) );
  XOR2_X1 U26688 ( .A1(n185), .A2(n25869), .Z(n50736) );
  XOR2_X1 U26689 ( .A1(n24930), .A2(n52446), .Z(n185) );
  INV_X2 U26692 ( .I(n51570), .ZN(n64370) );
  XOR2_X1 U26693 ( .A1(n51917), .A2(n16389), .Z(n18512) );
  NAND2_X2 U26698 ( .A1(n46856), .A2(n63136), .ZN(n51917) );
  NAND2_X1 U26701 ( .A1(n12830), .A2(n36256), .ZN(n16054) );
  BUF_X4 U26709 ( .I(n32400), .Z(n34350) );
  NAND2_X1 U26710 ( .A1(n63995), .A2(n595), .ZN(n57509) );
  NAND2_X1 U26712 ( .A1(n63694), .A2(n55933), .ZN(n63023) );
  NAND2_X1 U26713 ( .A1(n28881), .A2(n9138), .ZN(n26694) );
  NAND3_X2 U26714 ( .A1(n9139), .A2(n29351), .A3(n1892), .ZN(n28881) );
  NOR2_X2 U26723 ( .A1(n36196), .A2(n23503), .ZN(n36411) );
  NAND2_X2 U26724 ( .A1(n4263), .A2(n35361), .ZN(n36196) );
  NOR2_X2 U26726 ( .A1(n62906), .A2(n40121), .ZN(n40174) );
  NAND3_X2 U26733 ( .A1(n65238), .A2(n40115), .A3(n40114), .ZN(n62906) );
  NAND3_X2 U26734 ( .A1(n34259), .A2(n62907), .A3(n34257), .ZN(n34288) );
  XOR2_X1 U26737 ( .A1(n62909), .A2(n32545), .Z(n16132) );
  XOR2_X1 U26738 ( .A1(n32554), .A2(n59701), .Z(n62909) );
  XOR2_X1 U26742 ( .A1(n62910), .A2(n63548), .Z(n2703) );
  XOR2_X1 U26743 ( .A1(n16346), .A2(n18426), .Z(n62910) );
  NAND3_X2 U26744 ( .A1(n4468), .A2(n8746), .A3(n9350), .ZN(n8745) );
  NOR2_X2 U26745 ( .A1(n30782), .A2(n29957), .ZN(n28716) );
  XOR2_X1 U26748 ( .A1(n15410), .A2(n62911), .Z(n3556) );
  NOR2_X2 U26755 ( .A1(n6337), .A2(n15411), .ZN(n62911) );
  XOR2_X1 U26758 ( .A1(n62912), .A2(n23641), .Z(n787) );
  XOR2_X1 U26759 ( .A1(n43684), .A2(n20758), .Z(n62912) );
  INV_X4 U26760 ( .I(n1110), .ZN(n19489) );
  OR2_X2 U26762 ( .A1(n58666), .A2(n63472), .Z(n1110) );
  NAND2_X1 U26763 ( .A1(n8408), .A2(n11548), .ZN(n62913) );
  NAND2_X2 U26768 ( .A1(n35986), .A2(n6918), .ZN(n36705) );
  XOR2_X1 U26783 ( .A1(n65270), .A2(n62914), .Z(n60119) );
  XOR2_X1 U26785 ( .A1(n625), .A2(n3604), .Z(n62914) );
  NOR2_X2 U26786 ( .A1(n36715), .A2(n62916), .ZN(n25479) );
  NAND3_X2 U26788 ( .A1(n36712), .A2(n36713), .A3(n36711), .ZN(n62916) );
  NOR3_X2 U26789 ( .A1(n27192), .A2(n27193), .A3(n28112), .ZN(n29456) );
  NAND3_X2 U26790 ( .A1(n25270), .A2(n25272), .A3(n62918), .ZN(n15556) );
  AOI22_X2 U26795 ( .A1(n39115), .A2(n39116), .B1(n39114), .B2(n39113), .ZN(
        n62918) );
  OAI21_X1 U26802 ( .A1(n51903), .A2(n51902), .B(n55704), .ZN(n51904) );
  INV_X4 U26810 ( .I(n16629), .ZN(n24473) );
  NOR2_X2 U26812 ( .A1(n62784), .A2(n26665), .ZN(n12347) );
  BUF_X4 U26816 ( .I(n20280), .Z(n17364) );
  NOR2_X2 U26822 ( .A1(n64595), .A2(n20198), .ZN(n64664) );
  XOR2_X1 U26823 ( .A1(n62919), .A2(n744), .Z(n4813) );
  NOR2_X2 U26824 ( .A1(n11215), .A2(n11216), .ZN(n14372) );
  INV_X2 U26828 ( .I(n62921), .ZN(n39415) );
  NOR2_X2 U26830 ( .A1(n40167), .A2(n8453), .ZN(n62921) );
  INV_X2 U26836 ( .I(n62922), .ZN(n8452) );
  XNOR2_X1 U26846 ( .A1(n7106), .A2(n8454), .ZN(n62922) );
  INV_X4 U26849 ( .I(n15716), .ZN(n55898) );
  NAND3_X1 U26851 ( .A1(n8646), .A2(n8645), .A3(n47238), .ZN(n63472) );
  AOI21_X1 U26852 ( .A1(n61530), .A2(n3738), .B(n60520), .ZN(n49639) );
  NAND2_X1 U26854 ( .A1(n60005), .A2(n60004), .ZN(n62924) );
  BUF_X2 U26859 ( .I(n5140), .Z(n59052) );
  NOR2_X2 U26860 ( .A1(n40902), .A2(n62925), .ZN(n10278) );
  NAND2_X2 U26861 ( .A1(n41665), .A2(n42785), .ZN(n42188) );
  XOR2_X1 U26864 ( .A1(n64297), .A2(n62926), .Z(n63246) );
  XOR2_X1 U26868 ( .A1(n24978), .A2(n18514), .Z(n9948) );
  XOR2_X1 U26879 ( .A1(n16288), .A2(n25021), .Z(n24978) );
  XOR2_X1 U26883 ( .A1(n6302), .A2(n38575), .Z(n38576) );
  INV_X2 U26887 ( .I(n4808), .ZN(n15415) );
  NAND2_X2 U26906 ( .A1(n56815), .A2(n56791), .ZN(n56785) );
  NAND2_X2 U26909 ( .A1(n32868), .A2(n61731), .ZN(n3363) );
  INV_X2 U26914 ( .I(n38405), .ZN(n41161) );
  XOR2_X1 U26915 ( .A1(n62928), .A2(n17940), .Z(n51557) );
  XOR2_X1 U26917 ( .A1(n63819), .A2(n51556), .Z(n62928) );
  XOR2_X1 U26924 ( .A1(n2516), .A2(n51584), .Z(n58843) );
  XOR2_X1 U26929 ( .A1(n11469), .A2(n1617), .Z(n2516) );
  XOR2_X1 U26930 ( .A1(n51689), .A2(n62929), .Z(n54465) );
  XOR2_X1 U26931 ( .A1(n6447), .A2(n65018), .Z(n62929) );
  AND2_X1 U26933 ( .A1(n42990), .A2(n42989), .Z(n22985) );
  NAND3_X2 U26937 ( .A1(n25600), .A2(n1503), .A3(n12677), .ZN(n42989) );
  XOR2_X1 U26944 ( .A1(n8652), .A2(n21172), .Z(n30935) );
  NOR3_X2 U26951 ( .A1(n8476), .A2(n16694), .A3(n27307), .ZN(n28090) );
  NAND2_X2 U26953 ( .A1(n24299), .A2(n1253), .ZN(n8476) );
  XOR2_X1 U26955 ( .A1(n4860), .A2(n33173), .Z(n8567) );
  NAND2_X2 U26956 ( .A1(n14475), .A2(n29527), .ZN(n33173) );
  NAND2_X1 U26957 ( .A1(n10800), .A2(n40154), .ZN(n62930) );
  BUF_X2 U26958 ( .I(n1812), .Z(n62931) );
  AOI21_X1 U26965 ( .A1(n42430), .A2(n42431), .B(n42429), .ZN(n62932) );
  NAND2_X2 U26971 ( .A1(n9598), .A2(n36772), .ZN(n599) );
  XOR2_X1 U26979 ( .A1(n62933), .A2(n64311), .Z(n3879) );
  XOR2_X1 U26987 ( .A1(n3881), .A2(n59539), .Z(n62933) );
  BUF_X2 U26990 ( .I(n53056), .Z(n23243) );
  AND2_X1 U26992 ( .A1(n15616), .A2(n3142), .Z(n59082) );
  XOR2_X1 U26999 ( .A1(n36733), .A2(n64747), .Z(n3354) );
  XOR2_X1 U27000 ( .A1(n6302), .A2(n38999), .Z(n36733) );
  BUF_X2 U27001 ( .I(n58748), .Z(n62934) );
  XOR2_X1 U27002 ( .A1(n62935), .A2(n12727), .Z(n6728) );
  XOR2_X1 U27003 ( .A1(n44821), .A2(n9809), .Z(n62935) );
  XOR2_X1 U27004 ( .A1(n62936), .A2(n44132), .Z(n9926) );
  XOR2_X1 U27006 ( .A1(n18310), .A2(n44128), .Z(n62936) );
  NOR3_X2 U27007 ( .A1(n26160), .A2(n40192), .A3(n57624), .ZN(n22798) );
  NAND3_X2 U27008 ( .A1(n58434), .A2(n24570), .A3(n24568), .ZN(n46521) );
  XOR2_X1 U27014 ( .A1(n46646), .A2(n46202), .Z(n64863) );
  NAND2_X2 U27028 ( .A1(n302), .A2(n62937), .ZN(n30921) );
  INV_X2 U27032 ( .I(n49322), .ZN(n49324) );
  INV_X2 U27038 ( .I(n62938), .ZN(n10909) );
  XNOR2_X1 U27040 ( .A1(n21156), .A2(n16123), .ZN(n62938) );
  NOR2_X2 U27044 ( .A1(n12410), .A2(n6748), .ZN(n40146) );
  INV_X2 U27046 ( .I(n4673), .ZN(n12410) );
  OR2_X1 U27051 ( .A1(n35979), .A2(n8041), .Z(n62939) );
  BUF_X4 U27058 ( .I(n18063), .Z(n18425) );
  XOR2_X1 U27059 ( .A1(n62940), .A2(n17940), .Z(n667) );
  XOR2_X1 U27062 ( .A1(n52600), .A2(n52601), .Z(n62940) );
  NOR3_X2 U27063 ( .A1(n599), .A2(n62941), .A3(n2807), .ZN(n63618) );
  AOI21_X2 U27074 ( .A1(n61832), .A2(n36763), .B(n12031), .ZN(n62941) );
  NAND2_X2 U27077 ( .A1(n62943), .A2(n1171), .ZN(n54758) );
  NOR2_X1 U27083 ( .A1(n3944), .A2(n3945), .ZN(n62943) );
  INV_X2 U27088 ( .I(n62944), .ZN(n55024) );
  NAND2_X2 U27100 ( .A1(n15780), .A2(n667), .ZN(n62944) );
  XOR2_X1 U27104 ( .A1(n15914), .A2(n52585), .Z(n58370) );
  XOR2_X1 U27110 ( .A1(n33849), .A2(n13276), .Z(n4867) );
  INV_X1 U27111 ( .I(n43700), .ZN(n43702) );
  NOR2_X2 U27115 ( .A1(n4275), .A2(n42019), .ZN(n43700) );
  NAND2_X2 U27117 ( .A1(n4042), .A2(n913), .ZN(n58235) );
  OR2_X1 U27118 ( .A1(n34303), .A2(n34302), .Z(n57274) );
  NAND2_X2 U27125 ( .A1(n18989), .A2(n15830), .ZN(n34303) );
  OR2_X1 U27128 ( .A1(n50304), .A2(n50059), .Z(n62946) );
  AOI21_X2 U27130 ( .A1(n4548), .A2(n62947), .B(n34168), .ZN(n60899) );
  INV_X4 U27139 ( .I(n34695), .ZN(n7092) );
  XOR2_X1 U27140 ( .A1(n8381), .A2(n1683), .Z(n58310) );
  NOR2_X2 U27141 ( .A1(n63409), .A2(n61793), .ZN(n62949) );
  XOR2_X1 U27142 ( .A1(n20874), .A2(n58832), .Z(n13430) );
  NAND2_X2 U27143 ( .A1(n8110), .A2(n47064), .ZN(n20874) );
  XOR2_X1 U27145 ( .A1(n59721), .A2(n36903), .Z(n8454) );
  XOR2_X1 U27146 ( .A1(n61011), .A2(n62852), .Z(n36903) );
  NOR2_X2 U27155 ( .A1(n21377), .A2(n9334), .ZN(n21326) );
  INV_X4 U27157 ( .I(n56599), .ZN(n13757) );
  INV_X2 U27158 ( .I(n34649), .ZN(n57999) );
  NAND3_X2 U27163 ( .A1(n5902), .A2(n34631), .A3(n34502), .ZN(n34649) );
  INV_X2 U27164 ( .I(n15337), .ZN(n20632) );
  NAND2_X2 U27167 ( .A1(n42838), .A2(n8912), .ZN(n15337) );
  XOR2_X1 U27168 ( .A1(n14900), .A2(n14901), .Z(n44224) );
  NAND2_X2 U27172 ( .A1(n14899), .A2(n62950), .ZN(n14901) );
  OAI22_X2 U27179 ( .A1(n41482), .A2(n41483), .B1(n1298), .B2(n41481), .ZN(
        n41488) );
  NOR3_X2 U27180 ( .A1(n62954), .A2(n62953), .A3(n30645), .ZN(n30662) );
  OR2_X1 U27186 ( .A1(n30643), .A2(n30646), .Z(n62954) );
  NAND2_X2 U27187 ( .A1(n14894), .A2(n14891), .ZN(n8818) );
  BUF_X2 U27188 ( .I(n55722), .Z(n20653) );
  XOR2_X1 U27193 ( .A1(n21331), .A2(n2788), .Z(n24048) );
  NAND2_X1 U27199 ( .A1(n22738), .A2(n39120), .ZN(n62955) );
  NOR2_X2 U27201 ( .A1(n54961), .A2(n61736), .ZN(n54965) );
  XOR2_X1 U27206 ( .A1(n1907), .A2(n63962), .Z(n11339) );
  OAI22_X1 U27212 ( .A1(n62958), .A2(n62957), .B1(n55831), .B2(n55788), .ZN(
        n55789) );
  NAND2_X1 U27215 ( .A1(n55786), .A2(n55796), .ZN(n62958) );
  XOR2_X1 U27216 ( .A1(n21763), .A2(n21760), .Z(n22739) );
  NOR2_X1 U27222 ( .A1(n57707), .A2(n64409), .ZN(n55746) );
  XOR2_X1 U27225 ( .A1(n62959), .A2(n54126), .Z(Plaintext[54]) );
  NAND4_X1 U27228 ( .A1(n54124), .A2(n54125), .A3(n54122), .A4(n54123), .ZN(
        n62959) );
  NAND2_X2 U27229 ( .A1(n63952), .A2(n58435), .ZN(n40231) );
  NAND4_X2 U27231 ( .A1(n12745), .A2(n12744), .A3(n19147), .A4(n53762), .ZN(
        n63657) );
  XOR2_X1 U27233 ( .A1(n11574), .A2(n18435), .Z(n17237) );
  XOR2_X1 U27236 ( .A1(n11442), .A2(n17597), .Z(n11574) );
  XOR2_X1 U27237 ( .A1(n62964), .A2(n62574), .Z(n13778) );
  XOR2_X1 U27239 ( .A1(n64567), .A2(n21481), .Z(n62964) );
  XOR2_X1 U27241 ( .A1(n14740), .A2(n1888), .Z(n4681) );
  NAND3_X2 U27244 ( .A1(n8702), .A2(n8699), .A3(n8701), .ZN(n14740) );
  NAND2_X2 U27246 ( .A1(n1253), .A2(n15205), .ZN(n3052) );
  XOR2_X1 U27249 ( .A1(n62965), .A2(n4129), .Z(n11026) );
  XOR2_X1 U27250 ( .A1(n32557), .A2(n5433), .Z(n62965) );
  OR2_X1 U27253 ( .A1(n29155), .A2(n22482), .Z(n27263) );
  NAND3_X1 U27259 ( .A1(n49180), .A2(n49178), .A3(n49179), .ZN(n49184) );
  INV_X4 U27260 ( .I(n51863), .ZN(n53035) );
  NAND2_X1 U27263 ( .A1(n22273), .A2(n11761), .ZN(n11760) );
  NAND2_X2 U27270 ( .A1(n41840), .A2(n62969), .ZN(n43487) );
  AOI21_X2 U27271 ( .A1(n16469), .A2(n49932), .B(n53015), .ZN(n49933) );
  NAND2_X2 U27273 ( .A1(n51716), .A2(n53547), .ZN(n16469) );
  AOI22_X1 U27274 ( .A1(n55737), .A2(n52931), .B1(n52932), .B2(n14352), .ZN(
        n23101) );
  NOR2_X2 U27275 ( .A1(n55724), .A2(n55469), .ZN(n55737) );
  XOR2_X1 U27282 ( .A1(n9231), .A2(n14316), .Z(n50952) );
  NOR2_X1 U27287 ( .A1(n62972), .A2(n64538), .ZN(n64537) );
  NAND2_X1 U27288 ( .A1(n27515), .A2(n30720), .ZN(n62972) );
  AND2_X1 U27293 ( .A1(n14635), .A2(n54892), .Z(n57998) );
  NOR2_X2 U27294 ( .A1(n16143), .A2(n24261), .ZN(n18047) );
  XOR2_X1 U27296 ( .A1(n6832), .A2(n18868), .Z(n17404) );
  OAI21_X1 U27297 ( .A1(n42606), .A2(n42605), .B(n2121), .ZN(n42609) );
  XOR2_X1 U27300 ( .A1(n62973), .A2(n52205), .Z(n21598) );
  XOR2_X1 U27301 ( .A1(n52204), .A2(n52203), .Z(n62973) );
  INV_X2 U27302 ( .I(n54259), .ZN(n54266) );
  BUF_X4 U27303 ( .I(n45929), .Z(n344) );
  INV_X2 U27307 ( .I(n10282), .ZN(n64109) );
  NOR2_X2 U27313 ( .A1(n21345), .A2(n35109), .ZN(n18053) );
  NAND2_X2 U27315 ( .A1(n12748), .A2(n12749), .ZN(n21345) );
  INV_X2 U27323 ( .I(n41429), .ZN(n1723) );
  XOR2_X1 U27334 ( .A1(n62976), .A2(n25692), .Z(n45191) );
  XOR2_X1 U27339 ( .A1(n25694), .A2(n45024), .Z(n62976) );
  NAND2_X2 U27340 ( .A1(n19492), .A2(n59051), .ZN(n4316) );
  NAND2_X1 U27343 ( .A1(n64527), .A2(n57742), .ZN(n62977) );
  NAND2_X2 U27344 ( .A1(n40136), .A2(n40303), .ZN(n40220) );
  NAND2_X1 U27350 ( .A1(n12881), .A2(n12884), .ZN(n10484) );
  XOR2_X1 U27355 ( .A1(n22083), .A2(n15306), .Z(n19859) );
  OAI21_X2 U27356 ( .A1(n17952), .A2(n17954), .B(n21789), .ZN(n22083) );
  NAND3_X2 U27360 ( .A1(n24524), .A2(n62980), .A3(n62979), .ZN(n64000) );
  XOR2_X1 U27363 ( .A1(n6364), .A2(n6363), .Z(n19647) );
  XOR2_X1 U27364 ( .A1(n32514), .A2(n32515), .Z(n4650) );
  INV_X2 U27366 ( .I(n25935), .ZN(n32514) );
  NAND4_X2 U27373 ( .A1(n62981), .A2(n47538), .A3(n47537), .A4(n25387), .ZN(
        n12327) );
  XOR2_X1 U27385 ( .A1(n1214), .A2(n1329), .Z(n46268) );
  NOR2_X2 U27395 ( .A1(n37473), .A2(n37268), .ZN(n6632) );
  NAND2_X2 U27400 ( .A1(n36778), .A2(n5740), .ZN(n37473) );
  INV_X2 U27405 ( .I(n62982), .ZN(n16617) );
  NOR2_X1 U27411 ( .A1(n63877), .A2(n56537), .ZN(n56551) );
  INV_X2 U27413 ( .I(n25458), .ZN(n57528) );
  XOR2_X1 U27415 ( .A1(n52408), .A2(n15538), .Z(n15537) );
  NOR2_X2 U27416 ( .A1(n55144), .A2(n55143), .ZN(n21390) );
  NAND2_X1 U27420 ( .A1(n54844), .A2(n1456), .ZN(n52484) );
  NAND2_X2 U27426 ( .A1(n56719), .A2(n13249), .ZN(n56695) );
  XOR2_X1 U27440 ( .A1(n44144), .A2(n14513), .Z(n7699) );
  XOR2_X1 U27447 ( .A1(n46377), .A2(n45093), .Z(n44144) );
  XOR2_X1 U27450 ( .A1(n60050), .A2(n59618), .Z(n58582) );
  NAND4_X2 U27453 ( .A1(n9501), .A2(n9500), .A3(n9499), .A4(n49146), .ZN(
        n52596) );
  NAND2_X2 U27463 ( .A1(n11345), .A2(n64242), .ZN(n40242) );
  NAND2_X2 U27464 ( .A1(n8453), .A2(n8452), .ZN(n64242) );
  INV_X2 U27467 ( .I(n39100), .ZN(n39116) );
  NAND2_X2 U27468 ( .A1(n18032), .A2(n40196), .ZN(n39100) );
  NAND2_X2 U27469 ( .A1(n29292), .A2(n26446), .ZN(n5206) );
  NOR2_X2 U27471 ( .A1(n45596), .A2(n1483), .ZN(n24261) );
  XOR2_X1 U27474 ( .A1(n64454), .A2(n1094), .Z(n8846) );
  NAND2_X2 U27476 ( .A1(n2166), .A2(n40169), .ZN(n64689) );
  NOR2_X2 U27477 ( .A1(n2232), .A2(n1533), .ZN(n11980) );
  NAND2_X2 U27478 ( .A1(n15483), .A2(n351), .ZN(n15481) );
  NAND3_X1 U27482 ( .A1(n24805), .A2(n33811), .A3(n31956), .ZN(n31957) );
  NAND2_X2 U27486 ( .A1(n35312), .A2(n35255), .ZN(n24805) );
  XOR2_X1 U27487 ( .A1(n57908), .A2(n21794), .Z(n6917) );
  NAND4_X2 U27504 ( .A1(n9993), .A2(n48901), .A3(n15625), .A4(n48900), .ZN(
        n21794) );
  XOR2_X1 U27507 ( .A1(n10823), .A2(n5819), .Z(n32357) );
  NAND2_X2 U27511 ( .A1(n9185), .A2(n13823), .ZN(n41538) );
  NAND3_X1 U27513 ( .A1(n54898), .A2(n2474), .A3(n2049), .ZN(n54907) );
  AOI21_X2 U27514 ( .A1(n56797), .A2(n56796), .B(n56807), .ZN(n61614) );
  NAND2_X2 U27523 ( .A1(n1486), .A2(n43750), .ZN(n15421) );
  NAND2_X2 U27528 ( .A1(n16489), .A2(n53732), .ZN(n63449) );
  NOR2_X2 U27531 ( .A1(n31074), .A2(n31077), .ZN(n58931) );
  OAI22_X1 U27534 ( .A1(n63637), .A2(n9112), .B1(n52300), .B2(n52299), .ZN(
        n52304) );
  NAND3_X1 U27535 ( .A1(n41195), .A2(n41191), .A3(n39030), .ZN(n59488) );
  INV_X1 U27540 ( .I(n26248), .ZN(n63102) );
  NOR2_X1 U27542 ( .A1(n34941), .A2(n21467), .ZN(n64818) );
  NAND2_X1 U27546 ( .A1(n42460), .A2(n40360), .ZN(n63385) );
  NOR2_X2 U27558 ( .A1(n43873), .A2(n6144), .ZN(n4511) );
  INV_X4 U27560 ( .I(n12249), .ZN(n23643) );
  NAND3_X2 U27568 ( .A1(n19137), .A2(n18629), .A3(n62648), .ZN(n54098) );
  OAI21_X2 U27574 ( .A1(n36940), .A2(n36945), .B(n20616), .ZN(n36941) );
  NOR2_X2 U27577 ( .A1(n23206), .A2(n25267), .ZN(n3895) );
  NOR2_X2 U27580 ( .A1(n25413), .A2(n51112), .ZN(n56215) );
  NAND2_X2 U27581 ( .A1(n65002), .A2(n42863), .ZN(n65001) );
  NAND3_X2 U27582 ( .A1(n34232), .A2(n32071), .A3(n22797), .ZN(n34234) );
  NOR2_X2 U27584 ( .A1(n59621), .A2(n7868), .ZN(n49815) );
  INV_X2 U27585 ( .I(n1280), .ZN(n24520) );
  INV_X4 U27590 ( .I(n44802), .ZN(n47570) );
  NAND2_X1 U27595 ( .A1(n50547), .A2(n25487), .ZN(n63580) );
  NAND2_X2 U27599 ( .A1(n11912), .A2(n54487), .ZN(n24192) );
  NAND3_X1 U27601 ( .A1(n25119), .A2(n18792), .A3(n43443), .ZN(n65173) );
  NOR2_X1 U27604 ( .A1(n34745), .A2(n34744), .ZN(n64577) );
  NOR2_X2 U27622 ( .A1(n64777), .A2(n43084), .ZN(n5678) );
  BUF_X4 U27623 ( .I(n27507), .Z(n20930) );
  NOR2_X2 U27625 ( .A1(n47260), .A2(n47255), .ZN(n47267) );
  NAND2_X2 U27627 ( .A1(n54006), .A2(n22669), .ZN(n53962) );
  INV_X1 U27632 ( .I(n35970), .ZN(n33669) );
  NOR3_X1 U27646 ( .A1(n56691), .A2(n56690), .A3(n11851), .ZN(n56694) );
  OR2_X1 U27651 ( .A1(n14265), .A2(n47924), .Z(n58892) );
  INV_X1 U27657 ( .I(n47924), .ZN(n49725) );
  NOR2_X1 U27659 ( .A1(n48177), .A2(n48584), .ZN(n48174) );
  AOI21_X1 U27663 ( .A1(n36987), .A2(n37210), .B(n63682), .ZN(n36989) );
  NOR3_X1 U27667 ( .A1(n36987), .A2(n18583), .A3(n37210), .ZN(n36988) );
  OAI22_X1 U27668 ( .A1(n53575), .A2(n64521), .B1(n64522), .B2(n64520), .ZN(
        n53596) );
  OAI21_X1 U27669 ( .A1(n57183), .A2(n53577), .B(n64521), .ZN(n64520) );
  NAND2_X1 U27677 ( .A1(n23895), .A2(n44013), .ZN(n62985) );
  OAI21_X1 U27680 ( .A1(n22412), .A2(n47904), .B(n16162), .ZN(n47908) );
  OR2_X1 U27684 ( .A1(n16227), .A2(n15276), .Z(n64182) );
  INV_X1 U27693 ( .I(n56707), .ZN(n56615) );
  BUF_X2 U27703 ( .I(n61955), .Z(n65170) );
  NAND2_X2 U27708 ( .A1(n26124), .A2(n59230), .ZN(n6337) );
  NAND2_X1 U27717 ( .A1(n34676), .A2(n34675), .ZN(n64904) );
  CLKBUF_X4 U27721 ( .I(n53383), .Z(n23169) );
  NAND3_X1 U27722 ( .A1(n53486), .A2(n53484), .A3(n64671), .ZN(n64670) );
  INV_X1 U27727 ( .I(n58843), .ZN(n62986) );
  INV_X1 U27729 ( .I(n5141), .ZN(n22071) );
  INV_X1 U27741 ( .I(n17173), .ZN(n17172) );
  NAND2_X1 U27742 ( .A1(n64546), .A2(n64545), .ZN(n3386) );
  NAND2_X1 U27751 ( .A1(n49304), .A2(n19043), .ZN(n64546) );
  NAND2_X1 U27753 ( .A1(n60900), .A2(n23556), .ZN(n34236) );
  NOR2_X1 U27756 ( .A1(n54238), .A2(n23756), .ZN(n22315) );
  CLKBUF_X2 U27760 ( .I(n1280), .Z(n19404) );
  NOR2_X1 U27767 ( .A1(n55967), .A2(n55966), .ZN(n55670) );
  NOR2_X1 U27771 ( .A1(n53724), .A2(n17286), .ZN(n53757) );
  OAI21_X1 U27773 ( .A1(n7673), .A2(n47187), .B(n7674), .ZN(n7672) );
  INV_X2 U27777 ( .I(n25854), .ZN(n1463) );
  CLKBUF_X4 U27789 ( .I(n50898), .Z(n1616) );
  NAND2_X1 U27796 ( .A1(n55416), .A2(n65011), .ZN(n52573) );
  NOR2_X1 U27798 ( .A1(n55416), .A2(n55412), .ZN(n55407) );
  NAND3_X1 U27802 ( .A1(n1368), .A2(n54597), .A3(n54589), .ZN(n3884) );
  AOI21_X1 U27805 ( .A1(n54598), .A2(n54597), .B(n54596), .ZN(n54600) );
  NOR2_X1 U27807 ( .A1(n54597), .A2(n54074), .ZN(n54469) );
  NOR2_X1 U27809 ( .A1(n53894), .A2(n54597), .ZN(n22210) );
  NOR2_X1 U27814 ( .A1(n54597), .A2(n54472), .ZN(n54473) );
  INV_X1 U27817 ( .I(n35472), .ZN(n34895) );
  INV_X2 U27819 ( .I(n5172), .ZN(n56174) );
  INV_X2 U27822 ( .I(n52836), .ZN(n53601) );
  BUF_X4 U27824 ( .I(n20621), .Z(n15096) );
  INV_X1 U27825 ( .I(n9022), .ZN(n55714) );
  NAND2_X1 U27830 ( .A1(n56229), .A2(n9022), .ZN(n55988) );
  INV_X1 U27846 ( .I(n17984), .ZN(n7678) );
  AND2_X1 U27854 ( .A1(n54259), .A2(n54272), .Z(n54265) );
  INV_X2 U27856 ( .I(n55133), .ZN(n55170) );
  CLKBUF_X4 U27857 ( .I(n55133), .Z(n1593) );
  CLKBUF_X4 U27864 ( .I(n49281), .Z(n19107) );
  NOR2_X1 U27879 ( .A1(n55416), .A2(n24075), .ZN(n62988) );
  OAI21_X1 U27884 ( .A1(n49710), .A2(n7485), .B(n49709), .ZN(n9051) );
  NAND2_X1 U27888 ( .A1(n48792), .A2(n18469), .ZN(n9052) );
  CLKBUF_X4 U27914 ( .I(n42639), .Z(n1717) );
  NOR2_X1 U27915 ( .A1(n16716), .A2(n53527), .ZN(n53466) );
  NAND2_X1 U27921 ( .A1(n8047), .A2(n25896), .ZN(n5050) );
  INV_X1 U27927 ( .I(n54738), .ZN(n54712) );
  NAND3_X2 U27935 ( .A1(n14042), .A2(n50087), .A3(n14041), .ZN(n62989) );
  INV_X2 U27944 ( .I(n44092), .ZN(n23641) );
  INV_X1 U27947 ( .I(n47670), .ZN(n62990) );
  INV_X1 U27949 ( .I(n55680), .ZN(n62991) );
  CLKBUF_X4 U27955 ( .I(n52007), .Z(n55680) );
  NOR2_X1 U27961 ( .A1(n19307), .A2(n55868), .ZN(n55882) );
  CLKBUF_X2 U27962 ( .I(n53676), .Z(n23935) );
  OR2_X1 U27963 ( .A1(n54447), .A2(n14661), .Z(n54654) );
  INV_X2 U27966 ( .I(n5129), .ZN(n23919) );
  NOR2_X1 U27967 ( .A1(n19637), .A2(n53280), .ZN(n64482) );
  CLKBUF_X2 U27970 ( .I(n52547), .Z(n55400) );
  NOR2_X1 U27971 ( .A1(n56407), .A2(n57203), .ZN(n22387) );
  NAND3_X1 U27973 ( .A1(n52480), .A2(n55277), .A3(n55271), .ZN(n64496) );
  NAND2_X1 U27988 ( .A1(n22933), .A2(n55821), .ZN(n55786) );
  NOR2_X1 U27992 ( .A1(n52482), .A2(n64496), .ZN(n8328) );
  CLKBUF_X2 U28007 ( .I(n55275), .Z(n65101) );
  INV_X2 U28021 ( .I(n5532), .ZN(n1656) );
  NAND2_X1 U28025 ( .A1(n15632), .A2(n20653), .ZN(n55720) );
  AND2_X2 U28026 ( .A1(n7074), .A2(n35852), .Z(n62992) );
  NAND2_X1 U28028 ( .A1(n11869), .A2(n53428), .ZN(n11868) );
  AOI21_X1 U28029 ( .A1(n56089), .A2(n56090), .B(n56110), .ZN(n56094) );
  INV_X4 U28030 ( .I(n55569), .ZN(n55565) );
  INV_X2 U28031 ( .I(n55385), .ZN(n9421) );
  XNOR2_X1 U28033 ( .A1(n46187), .A2(n44909), .ZN(n12755) );
  NOR3_X1 U28035 ( .A1(n54390), .A2(n54354), .A3(n54380), .ZN(n54421) );
  INV_X2 U28047 ( .I(n5323), .ZN(n54380) );
  NAND2_X1 U28049 ( .A1(n7518), .A2(n54966), .ZN(n54630) );
  NOR2_X1 U28052 ( .A1(n16971), .A2(n15126), .ZN(n62994) );
  NAND2_X1 U28059 ( .A1(n16147), .A2(n30362), .ZN(n3169) );
  NOR2_X1 U28062 ( .A1(n62994), .A2(n21159), .ZN(n16147) );
  NAND2_X1 U28064 ( .A1(n61197), .A2(n61196), .ZN(n33359) );
  AOI21_X1 U28065 ( .A1(n25280), .A2(n29930), .B(n10821), .ZN(n25279) );
  NAND3_X1 U28069 ( .A1(n49072), .A2(n23238), .A3(n49835), .ZN(n57574) );
  NAND3_X1 U28070 ( .A1(n35753), .A2(n35764), .A3(n35320), .ZN(n35323) );
  NOR3_X1 U28076 ( .A1(n4658), .A2(n60225), .A3(n57032), .ZN(n57035) );
  NAND2_X1 U28078 ( .A1(n52237), .A2(n4658), .ZN(n52238) );
  OAI22_X1 U28081 ( .A1(n46815), .A2(n46816), .B1(n57463), .B2(n12698), .ZN(
        n12794) );
  AND3_X1 U28092 ( .A1(n12959), .A2(n61361), .A3(n4283), .Z(n62996) );
  NAND3_X1 U28095 ( .A1(n63376), .A2(n24115), .A3(n55206), .ZN(n55207) );
  OAI22_X1 U28099 ( .A1(n55199), .A2(n55198), .B1(n55201), .B2(n55200), .ZN(
        n63376) );
  NAND2_X1 U28102 ( .A1(n7824), .A2(n7588), .ZN(n49343) );
  AOI21_X1 U28105 ( .A1(n61846), .A2(n7824), .B(n50013), .ZN(n25503) );
  INV_X2 U28109 ( .I(n5115), .ZN(n39502) );
  INV_X1 U28114 ( .I(n21364), .ZN(n54472) );
  INV_X2 U28118 ( .I(n2736), .ZN(n22533) );
  INV_X1 U28120 ( .I(n78), .ZN(n63369) );
  NOR2_X1 U28129 ( .A1(n22805), .A2(n78), .ZN(n49254) );
  INV_X1 U28130 ( .I(n56817), .ZN(n20438) );
  NOR2_X1 U28134 ( .A1(n49270), .A2(n49407), .ZN(n22847) );
  OAI21_X1 U28135 ( .A1(n49269), .A2(n49270), .B(n9395), .ZN(n49271) );
  BUF_X4 U28136 ( .I(n51449), .Z(n56817) );
  INV_X1 U28139 ( .I(n306), .ZN(n62998) );
  NAND2_X1 U28142 ( .A1(n42006), .A2(n43094), .ZN(n7401) );
  BUF_X2 U28148 ( .I(n57079), .Z(n64338) );
  NAND3_X1 U28149 ( .A1(n61191), .A2(n23263), .A3(n48642), .ZN(n4213) );
  INV_X1 U28150 ( .I(n61646), .ZN(n33389) );
  NOR2_X1 U28155 ( .A1(n2005), .A2(n1319), .ZN(n62999) );
  NAND3_X1 U28163 ( .A1(n60770), .A2(n35478), .A3(n60771), .ZN(n63000) );
  NOR2_X1 U28166 ( .A1(n2005), .A2(n1319), .ZN(n2921) );
  NAND2_X1 U28190 ( .A1(n1426), .A2(n35774), .ZN(n35786) );
  INV_X2 U28193 ( .I(n29448), .ZN(n14647) );
  NAND2_X1 U28197 ( .A1(n29448), .A2(n63417), .ZN(n29839) );
  INV_X1 U28202 ( .I(n21984), .ZN(n51289) );
  INV_X1 U28203 ( .I(n55425), .ZN(n50932) );
  NAND2_X1 U28208 ( .A1(n63368), .A2(n47458), .ZN(n58980) );
  INV_X1 U28210 ( .I(n22258), .ZN(n64038) );
  INV_X1 U28211 ( .I(n48292), .ZN(n48293) );
  OAI21_X1 U28214 ( .A1(n50291), .A2(n21092), .B(n22867), .ZN(n21790) );
  INV_X1 U28215 ( .I(n5945), .ZN(n57610) );
  NOR2_X1 U28221 ( .A1(n54268), .A2(n24520), .ZN(n54269) );
  INV_X1 U28223 ( .I(n31254), .ZN(n31245) );
  AND2_X2 U28225 ( .A1(n25007), .A2(n2737), .Z(n47860) );
  BUF_X2 U28228 ( .I(n49598), .Z(n25032) );
  INV_X1 U28232 ( .I(n63106), .ZN(n63852) );
  CLKBUF_X8 U28234 ( .I(n47524), .Z(n49195) );
  NOR3_X1 U28235 ( .A1(n12818), .A2(n4658), .A3(n53212), .ZN(n25198) );
  AOI21_X1 U28238 ( .A1(n51265), .A2(n25167), .B(n51268), .ZN(n23377) );
  CLKBUF_X4 U28239 ( .I(n1256), .Z(n63873) );
  NAND4_X1 U28241 ( .A1(n5621), .A2(n52899), .A3(n4601), .A4(n52898), .ZN(n569) );
  CLKBUF_X8 U28259 ( .I(n23863), .Z(n4547) );
  NOR2_X1 U28263 ( .A1(n61343), .A2(n63253), .ZN(n25616) );
  NAND2_X1 U28264 ( .A1(n35570), .A2(n4802), .ZN(n34825) );
  OR2_X1 U28266 ( .A1(n24361), .A2(n8986), .Z(n41651) );
  CLKBUF_X4 U28275 ( .I(n35092), .Z(n35096) );
  INV_X2 U28277 ( .I(n36986), .ZN(n37225) );
  NOR2_X1 U28278 ( .A1(n53297), .A2(n25199), .ZN(n64483) );
  NAND2_X1 U28279 ( .A1(n1164), .A2(n53294), .ZN(n53297) );
  INV_X2 U28281 ( .I(n6342), .ZN(n44948) );
  NOR3_X1 U28284 ( .A1(n48063), .A2(n201), .A3(n19681), .ZN(n59167) );
  NAND2_X1 U28286 ( .A1(n63310), .A2(n63309), .ZN(n9078) );
  NOR2_X1 U28289 ( .A1(n49528), .A2(n49538), .ZN(n48902) );
  AOI22_X1 U28291 ( .A1(n44660), .A2(n6081), .B1(n9972), .B2(n23990), .ZN(
        n4738) );
  INV_X2 U28294 ( .I(n62978), .ZN(n9972) );
  NAND2_X1 U28296 ( .A1(n6360), .A2(n34079), .ZN(n63234) );
  NAND4_X1 U28297 ( .A1(n404), .A2(n40067), .A3(n40068), .A4(n40231), .ZN(
        n25468) );
  INV_X1 U28298 ( .I(n55084), .ZN(n64987) );
  CLKBUF_X2 U28301 ( .I(n2960), .Z(n65058) );
  INV_X1 U28304 ( .I(n52563), .ZN(n59904) );
  OAI22_X1 U28307 ( .A1(n52574), .A2(n55415), .B1(n55416), .B2(n65011), .ZN(
        n7666) );
  NAND2_X1 U28311 ( .A1(n55415), .A2(n55414), .ZN(n55417) );
  OR3_X1 U28313 ( .A1(n56509), .A2(n19827), .A3(n1366), .Z(n59780) );
  CLKBUF_X4 U28315 ( .I(n55884), .Z(n15716) );
  NOR2_X1 U28318 ( .A1(n63170), .A2(n57501), .ZN(n49816) );
  AOI21_X1 U28321 ( .A1(n49814), .A2(n8898), .B(n7868), .ZN(n63170) );
  INV_X1 U28322 ( .I(n59621), .ZN(n50438) );
  CLKBUF_X4 U28330 ( .I(n52174), .Z(n23173) );
  NAND3_X1 U28336 ( .A1(n15202), .A2(n54424), .A3(n1367), .ZN(n54354) );
  AND2_X2 U28339 ( .A1(n55443), .A2(n24166), .Z(n55310) );
  INV_X1 U28340 ( .I(n64263), .ZN(n36249) );
  INV_X2 U28342 ( .I(n55909), .ZN(n18886) );
  NAND2_X2 U28347 ( .A1(n25951), .A2(n57921), .ZN(n63001) );
  OAI21_X1 U28350 ( .A1(n63449), .A2(n53726), .B(n25117), .ZN(n53711) );
  INV_X1 U28355 ( .I(n59831), .ZN(n24111) );
  CLKBUF_X8 U28363 ( .I(n53448), .Z(n53492) );
  INV_X1 U28368 ( .I(n37117), .ZN(n16563) );
  NAND2_X1 U28369 ( .A1(n20269), .A2(n56687), .ZN(n64649) );
  OR2_X2 U28380 ( .A1(n53161), .A2(n23116), .Z(n53148) );
  OR2_X2 U28384 ( .A1(n53161), .A2(n53146), .Z(n53166) );
  AOI21_X1 U28388 ( .A1(n53194), .A2(n11041), .B(n53607), .ZN(n12833) );
  INV_X1 U28390 ( .I(n1196), .ZN(n63003) );
  INV_X2 U28393 ( .I(n1196), .ZN(n1197) );
  NOR2_X1 U28398 ( .A1(n8356), .A2(n19364), .ZN(n35526) );
  CLKBUF_X4 U28406 ( .I(n53905), .Z(n23164) );
  AOI21_X1 U28408 ( .A1(n50274), .A2(n50273), .B(n21835), .ZN(n50281) );
  OR2_X2 U28409 ( .A1(n24596), .A2(n25445), .Z(n63004) );
  INV_X1 U28410 ( .I(n18191), .ZN(n21905) );
  OAI21_X1 U28411 ( .A1(n52944), .A2(n8055), .B(n58283), .ZN(n8054) );
  INV_X1 U28412 ( .I(n2886), .ZN(n63723) );
  INV_X1 U28413 ( .I(n5193), .ZN(n18175) );
  NAND2_X1 U28415 ( .A1(n11716), .A2(n5193), .ZN(n56172) );
  NAND2_X1 U28425 ( .A1(n53214), .A2(n25868), .ZN(n57024) );
  NOR2_X2 U28426 ( .A1(n48804), .A2(n48421), .ZN(n48427) );
  OR2_X2 U28430 ( .A1(n13871), .A2(n13872), .Z(n63005) );
  NAND3_X2 U28433 ( .A1(n52856), .A2(n52855), .A3(n17181), .ZN(n17180) );
  NAND2_X1 U28438 ( .A1(n46885), .A2(n47247), .ZN(n46883) );
  NAND3_X1 U28439 ( .A1(n45922), .A2(n15569), .A3(n25831), .ZN(n25830) );
  NAND2_X1 U28456 ( .A1(n53209), .A2(n53443), .ZN(n53434) );
  NAND2_X1 U28467 ( .A1(n64489), .A2(n25490), .ZN(n12782) );
  XNOR2_X1 U28473 ( .A1(n52569), .A2(n14730), .ZN(n14742) );
  INV_X2 U28476 ( .I(n1486), .ZN(n47736) );
  XOR2_X1 U28481 ( .A1(Key[43]), .A2(Ciphertext[90]), .Z(n63007) );
  BUF_X2 U28482 ( .I(Key[191]), .Z(n57162) );
  NOR2_X1 U28484 ( .A1(n20276), .A2(n43912), .ZN(n12645) );
  NAND2_X1 U28495 ( .A1(n52705), .A2(n56545), .ZN(n52710) );
  NOR2_X1 U28499 ( .A1(n47250), .A2(n59418), .ZN(n46894) );
  NAND3_X1 U28504 ( .A1(n48791), .A2(n48421), .A3(n61742), .ZN(n48347) );
  NOR2_X2 U28505 ( .A1(n51905), .A2(n50882), .ZN(n55709) );
  INV_X1 U28507 ( .I(n14990), .ZN(n59177) );
  NAND2_X1 U28514 ( .A1(n4199), .A2(n5773), .ZN(n42108) );
  INV_X1 U28520 ( .I(n21459), .ZN(n41923) );
  NAND3_X1 U28521 ( .A1(n53342), .A2(n26236), .A3(n64909), .ZN(n63924) );
  NOR2_X1 U28540 ( .A1(n64246), .A2(n56853), .ZN(n56887) );
  INV_X1 U28544 ( .I(n33110), .ZN(n36057) );
  CLKBUF_X4 U28546 ( .I(n15928), .Z(n23206) );
  NAND4_X1 U28547 ( .A1(n55732), .A2(n55731), .A3(n55734), .A4(n55733), .ZN(
        n57707) );
  BUF_X2 U28548 ( .I(n27591), .Z(n7943) );
  INV_X2 U28549 ( .I(n1139), .ZN(n1604) );
  NOR2_X2 U28550 ( .A1(n16868), .A2(n17089), .ZN(n63009) );
  OAI22_X2 U28568 ( .A1(n47980), .A2(n17091), .B1(n47979), .B2(n17090), .ZN(
        n17089) );
  NAND2_X1 U28569 ( .A1(n16675), .A2(n49997), .ZN(n16674) );
  NOR2_X1 U28570 ( .A1(n1377), .A2(n48717), .ZN(n47955) );
  NAND2_X1 U28578 ( .A1(n57182), .A2(n1377), .ZN(n21188) );
  BUF_X2 U28580 ( .I(Key[184]), .Z(n56949) );
  OAI21_X1 U28582 ( .A1(n49511), .A2(n49525), .B(n406), .ZN(n49514) );
  CLKBUF_X2 U28583 ( .I(n52053), .Z(n8006) );
  NAND2_X1 U28590 ( .A1(n49598), .A2(n25320), .ZN(n59086) );
  CLKBUF_X4 U28595 ( .I(n50257), .Z(n21052) );
  INV_X1 U28601 ( .I(n50257), .ZN(n50333) );
  NAND2_X1 U28602 ( .A1(n17896), .A2(n17895), .ZN(n60595) );
  NAND2_X1 U28603 ( .A1(n60651), .A2(n48572), .ZN(n60410) );
  CLKBUF_X4 U28608 ( .I(n37388), .Z(n21881) );
  CLKBUF_X2 U28609 ( .I(n22385), .Z(n59051) );
  AND2_X2 U28613 ( .A1(n61728), .A2(n48074), .Z(n48691) );
  INV_X1 U28614 ( .I(n5277), .ZN(n16846) );
  NAND3_X1 U28615 ( .A1(n53877), .A2(n53876), .A3(n59831), .ZN(n10008) );
  BUF_X2 U28618 ( .I(n10802), .Z(n23277) );
  CLKBUF_X4 U28623 ( .I(n20138), .Z(n61083) );
  NAND3_X1 U28625 ( .A1(n53297), .A2(n53296), .A3(n53295), .ZN(n53298) );
  CLKBUF_X4 U28634 ( .I(n8175), .Z(n8122) );
  NAND2_X1 U28635 ( .A1(n43021), .A2(n43019), .ZN(n64125) );
  NOR2_X1 U28637 ( .A1(n1656), .A2(n2641), .ZN(n16183) );
  NOR2_X1 U28638 ( .A1(n5554), .A2(n2641), .ZN(n9742) );
  NAND3_X1 U28639 ( .A1(n24117), .A2(n16978), .A3(n55222), .ZN(n22497) );
  NAND2_X1 U28646 ( .A1(n15747), .A2(n25522), .ZN(n53577) );
  NAND2_X2 U28647 ( .A1(n13197), .A2(n7431), .ZN(n63010) );
  CLKBUF_X4 U28649 ( .I(n54717), .Z(n22122) );
  INV_X1 U28651 ( .I(n34026), .ZN(n1803) );
  NOR2_X1 U28658 ( .A1(n34026), .A2(n902), .ZN(n15547) );
  NOR3_X1 U28662 ( .A1(n35023), .A2(n34026), .A3(n64499), .ZN(n64498) );
  AOI21_X1 U28663 ( .A1(n51706), .A2(n6211), .B(n59530), .ZN(n65204) );
  INV_X2 U28666 ( .I(n56435), .ZN(n55982) );
  NAND3_X1 U28675 ( .A1(n24551), .A2(n56452), .A3(n56451), .ZN(n56512) );
  INV_X1 U28681 ( .I(n55075), .ZN(n55095) );
  INV_X1 U28682 ( .I(n24181), .ZN(n10562) );
  INV_X1 U28687 ( .I(n46716), .ZN(n48538) );
  INV_X4 U28689 ( .I(n12100), .ZN(n46716) );
  NAND2_X1 U28693 ( .A1(n48232), .A2(n46716), .ZN(n47189) );
  CLKBUF_X2 U28695 ( .I(n52421), .Z(n7343) );
  INV_X1 U28700 ( .I(n36772), .ZN(n34371) );
  BUF_X2 U28702 ( .I(Key[170]), .Z(n56771) );
  AND2_X2 U28709 ( .A1(n9334), .A2(n21377), .Z(n41554) );
  CLKBUF_X4 U28710 ( .I(n19491), .Z(n19492) );
  NAND2_X1 U28714 ( .A1(n58326), .A2(n57072), .ZN(n65187) );
  AOI21_X1 U28715 ( .A1(n50602), .A2(n52255), .B(n57072), .ZN(n50603) );
  BUF_X2 U28716 ( .I(n23415), .Z(n10713) );
  NAND2_X2 U28718 ( .A1(n5109), .A2(n5110), .ZN(n5108) );
  NAND2_X1 U28719 ( .A1(n51887), .A2(n15454), .ZN(n20018) );
  NAND2_X1 U28722 ( .A1(n51887), .A2(n52120), .ZN(n58460) );
  NAND2_X1 U28728 ( .A1(n43995), .A2(n23314), .ZN(n43990) );
  INV_X4 U28729 ( .I(n43995), .ZN(n1334) );
  NAND2_X1 U28734 ( .A1(n6008), .A2(n55971), .ZN(n63012) );
  NAND2_X2 U28735 ( .A1(n6008), .A2(n55971), .ZN(n63013) );
  NAND2_X1 U28739 ( .A1(n6008), .A2(n55971), .ZN(n56085) );
  INV_X2 U28741 ( .I(n54546), .ZN(n54543) );
  INV_X1 U28748 ( .I(n55310), .ZN(n55321) );
  CLKBUF_X4 U28755 ( .I(n52648), .Z(n9550) );
  NOR2_X1 U28757 ( .A1(n41775), .A2(n25126), .ZN(n42177) );
  NAND2_X1 U28760 ( .A1(n56922), .A2(n59853), .ZN(n23832) );
  CLKBUF_X4 U28761 ( .I(n44802), .Z(n47572) );
  NOR3_X1 U28772 ( .A1(n23212), .A2(n53107), .A3(n53108), .ZN(n53117) );
  INV_X2 U28775 ( .I(n53107), .ZN(n53070) );
  BUF_X2 U28782 ( .I(n53077), .Z(n22980) );
  NAND2_X1 U28789 ( .A1(n61673), .A2(n48847), .ZN(n48843) );
  NOR2_X1 U28791 ( .A1(n15101), .A2(n39102), .ZN(n58369) );
  OR2_X2 U28792 ( .A1(n15101), .A2(n24246), .Z(n825) );
  NAND2_X2 U28793 ( .A1(n24174), .A2(n24176), .ZN(n63014) );
  NAND3_X1 U28794 ( .A1(n53926), .A2(n53966), .A3(n54001), .ZN(n53904) );
  OR2_X1 U28795 ( .A1(n1697), .A2(n20922), .Z(n9043) );
  INV_X2 U28796 ( .I(n13166), .ZN(n14773) );
  NAND2_X1 U28797 ( .A1(n25026), .A2(n64548), .ZN(n47723) );
  AND2_X2 U28798 ( .A1(n13393), .A2(n40020), .Z(n42371) );
  NAND2_X1 U28805 ( .A1(n60401), .A2(n41904), .ZN(n5513) );
  INV_X1 U28806 ( .I(n8462), .ZN(n4354) );
  INV_X1 U28810 ( .I(n45333), .ZN(n20413) );
  NOR2_X1 U28815 ( .A1(n55375), .A2(n55376), .ZN(n18134) );
  OAI21_X1 U28816 ( .A1(n54996), .A2(n55270), .B(n18790), .ZN(n52944) );
  OR3_X1 U28817 ( .A1(n54740), .A2(n54741), .A3(n19492), .Z(n54746) );
  NAND4_X1 U28819 ( .A1(n55861), .A2(n55860), .A3(n55858), .A4(n55859), .ZN(
        n55863) );
  INV_X1 U28823 ( .I(n4145), .ZN(n64758) );
  INV_X1 U28835 ( .I(n55734), .ZN(n58553) );
  NAND2_X1 U28837 ( .A1(n56868), .A2(n5658), .ZN(n56843) );
  INV_X1 U28839 ( .I(n29643), .ZN(n28598) );
  INV_X1 U28840 ( .I(n53130), .ZN(n21590) );
  INV_X4 U28841 ( .I(n24287), .ZN(n17283) );
  INV_X1 U28845 ( .I(n41146), .ZN(n1507) );
  NAND2_X1 U28846 ( .A1(n41146), .A2(n5950), .ZN(n41153) );
  NAND2_X1 U28847 ( .A1(n41146), .A2(n23875), .ZN(n13357) );
  CLKBUF_X2 U28848 ( .I(n41146), .Z(n60139) );
  CLKBUF_X4 U28852 ( .I(n20892), .Z(n17774) );
  NAND3_X1 U28853 ( .A1(n55883), .A2(n55898), .A3(n13858), .ZN(n55843) );
  AOI21_X1 U28855 ( .A1(n54268), .A2(n54259), .B(n54281), .ZN(n54210) );
  NAND2_X1 U28857 ( .A1(n56897), .A2(n10507), .ZN(n56853) );
  AND2_X2 U28859 ( .A1(n24420), .A2(n22349), .Z(n61169) );
  CLKBUF_X4 U28868 ( .I(n27233), .Z(n64994) );
  CLKBUF_X12 U28873 ( .I(n38759), .Z(n40748) );
  AOI21_X1 U28874 ( .A1(n52845), .A2(n23974), .B(n53198), .ZN(n23891) );
  OAI22_X1 U28879 ( .A1(n58388), .A2(n58387), .B1(n29233), .B2(n61229), .ZN(
        n19635) );
  XOR2_X1 U28900 ( .A1(n58455), .A2(n3504), .Z(n63016) );
  XOR2_X1 U28902 ( .A1(n65214), .A2(n8864), .Z(n63017) );
  INV_X1 U28905 ( .I(n63712), .ZN(n47918) );
  INV_X1 U28911 ( .I(n11912), .ZN(n54481) );
  INV_X4 U28913 ( .I(n17958), .ZN(n25256) );
  CLKBUF_X4 U28915 ( .I(n34336), .Z(n17958) );
  NOR2_X1 U28919 ( .A1(n20547), .A2(n19434), .ZN(n53178) );
  NOR3_X1 U28921 ( .A1(n55643), .A2(n3307), .A3(n15700), .ZN(n52311) );
  NAND3_X1 U28926 ( .A1(n52298), .A2(n55643), .A3(n55639), .ZN(n63637) );
  NAND2_X1 U28931 ( .A1(n55643), .A2(n59610), .ZN(n52302) );
  NAND2_X1 U28941 ( .A1(n55643), .A2(n19021), .ZN(n55604) );
  NOR2_X1 U28950 ( .A1(n10113), .A2(n13025), .ZN(n19644) );
  NOR2_X1 U28953 ( .A1(n75), .A2(n5178), .ZN(n63130) );
  INV_X1 U28955 ( .I(n24780), .ZN(n63018) );
  XOR2_X1 U28959 ( .A1(n13619), .A2(n13618), .Z(n63019) );
  NAND2_X1 U28960 ( .A1(n55684), .A2(n64019), .ZN(n55686) );
  NAND3_X1 U28964 ( .A1(n47249), .A2(n47248), .A3(n47247), .ZN(n47269) );
  INV_X1 U28970 ( .I(n47260), .ZN(n15568) );
  AND4_X2 U28972 ( .A1(n54832), .A2(n54829), .A3(n54830), .A4(n54831), .Z(
        n63020) );
  NAND3_X1 U28980 ( .A1(n22337), .A2(n54599), .A3(n54601), .ZN(n53892) );
  AOI21_X1 U28982 ( .A1(n16445), .A2(n37420), .B(n16444), .ZN(n16443) );
  OAI21_X1 U28992 ( .A1(n16445), .A2(n35510), .B(n16442), .ZN(n63131) );
  NOR2_X1 U28995 ( .A1(n30437), .A2(n1253), .ZN(n30546) );
  CLKBUF_X8 U28996 ( .I(n24425), .Z(n12034) );
  AOI21_X1 U28998 ( .A1(n39851), .A2(n41399), .B(n39850), .ZN(n64321) );
  NAND3_X1 U28999 ( .A1(n55036), .A2(n55035), .A3(n9067), .ZN(n55039) );
  BUF_X2 U29000 ( .I(n25158), .Z(n16508) );
  INV_X2 U29001 ( .I(n22881), .ZN(n6007) );
  OR2_X2 U29013 ( .A1(n20211), .A2(n16177), .Z(n63021) );
  AND2_X2 U29020 ( .A1(n5215), .A2(n64456), .Z(n63022) );
  NOR2_X2 U29022 ( .A1(n5217), .A2(n5216), .ZN(n5215) );
  NAND4_X2 U29030 ( .A1(n58303), .A2(n64286), .A3(n54307), .A4(n61371), .ZN(
        n18655) );
  INV_X1 U29034 ( .I(n54071), .ZN(n64286) );
  CLKBUF_X2 U29035 ( .I(n19349), .Z(n9416) );
  NAND3_X1 U29038 ( .A1(n18858), .A2(n17467), .A3(n42676), .ZN(n42823) );
  NAND2_X1 U29050 ( .A1(n56539), .A2(n52706), .ZN(n24668) );
  NAND2_X1 U29051 ( .A1(n49458), .A2(n57312), .ZN(n49461) );
  INV_X1 U29052 ( .I(n49458), .ZN(n49229) );
  NAND2_X1 U29062 ( .A1(n49458), .A2(n57610), .ZN(n57609) );
  OAI21_X1 U29064 ( .A1(n47797), .A2(n47700), .B(n47813), .ZN(n44000) );
  CLKBUF_X12 U29066 ( .I(n47017), .Z(n7104) );
  NAND2_X1 U29069 ( .A1(n47017), .A2(n5771), .ZN(n12225) );
  NAND3_X1 U29073 ( .A1(n8203), .A2(n55295), .A3(n55684), .ZN(n17753) );
  AOI21_X1 U29076 ( .A1(n16847), .A2(n6235), .B(n5279), .ZN(n5278) );
  NOR3_X2 U29084 ( .A1(n7763), .A2(n7762), .A3(n7766), .ZN(n10680) );
  NAND2_X1 U29085 ( .A1(n56389), .A2(n11119), .ZN(n56390) );
  CLKBUF_X4 U29089 ( .I(n1487), .Z(n48594) );
  INV_X1 U29095 ( .I(n16886), .ZN(n35567) );
  NAND2_X1 U29096 ( .A1(n6333), .A2(n63569), .ZN(n63568) );
  NAND2_X1 U29097 ( .A1(n60845), .A2(n6333), .ZN(n51775) );
  CLKBUF_X4 U29099 ( .I(n51818), .Z(n22979) );
  NAND3_X1 U29100 ( .A1(n10248), .A2(n55829), .A3(n55828), .ZN(n63177) );
  NAND2_X1 U29113 ( .A1(n10248), .A2(n55772), .ZN(n55826) );
  INV_X1 U29118 ( .I(n10248), .ZN(n55795) );
  NAND2_X1 U29119 ( .A1(n24820), .A2(n5771), .ZN(n8696) );
  NAND2_X1 U29120 ( .A1(n3708), .A2(n54659), .ZN(n59142) );
  NAND2_X1 U29122 ( .A1(n65147), .A2(n61134), .ZN(n38354) );
  NOR2_X1 U29125 ( .A1(n61134), .A2(n42750), .ZN(n43052) );
  NOR2_X1 U29126 ( .A1(n61134), .A2(n8305), .ZN(n43875) );
  NAND3_X1 U29130 ( .A1(n58367), .A2(n4819), .A3(n5675), .ZN(n5674) );
  CLKBUF_X8 U29136 ( .I(n44658), .Z(n49910) );
  CLKBUF_X4 U29138 ( .I(n26245), .Z(n20073) );
  BUF_X2 U29139 ( .I(n9288), .Z(n9040) );
  BUF_X2 U29141 ( .I(n37285), .Z(n38784) );
  INV_X2 U29142 ( .I(n14251), .ZN(n59811) );
  AND2_X2 U29148 ( .A1(n12798), .A2(n7074), .Z(n37168) );
  NAND3_X1 U29152 ( .A1(n36794), .A2(n24351), .A3(n10110), .ZN(n36069) );
  OAI21_X1 U29156 ( .A1(n54767), .A2(n54742), .B(n61057), .ZN(n60688) );
  NAND3_X2 U29160 ( .A1(n27333), .A2(n27332), .A3(n27331), .ZN(n27334) );
  CLKBUF_X12 U29162 ( .I(n30994), .Z(n191) );
  CLKBUF_X4 U29163 ( .I(n24209), .Z(n7271) );
  BUF_X2 U29164 ( .I(n13808), .Z(n9397) );
  BUF_X4 U29165 ( .I(n47055), .Z(n48323) );
  NAND2_X1 U29169 ( .A1(n23581), .A2(n47055), .ZN(n48031) );
  INV_X1 U29173 ( .I(n47055), .ZN(n9853) );
  NAND2_X1 U29174 ( .A1(n20923), .A2(n24287), .ZN(n17282) );
  BUF_X4 U29176 ( .I(n35140), .Z(n35965) );
  CLKBUF_X8 U29177 ( .I(n3864), .Z(n36790) );
  BUF_X4 U29179 ( .I(n34575), .Z(n3864) );
  INV_X4 U29180 ( .I(n47534), .ZN(n5771) );
  CLKBUF_X4 U29185 ( .I(n47534), .Z(n59056) );
  INV_X1 U29188 ( .I(n10618), .ZN(n51097) );
  CLKBUF_X2 U29192 ( .I(n52157), .Z(n2604) );
  INV_X1 U29193 ( .I(n22267), .ZN(n59963) );
  NAND2_X1 U29205 ( .A1(n31357), .A2(n12547), .ZN(n34520) );
  OAI21_X1 U29207 ( .A1(n43089), .A2(n42999), .B(n61864), .ZN(n19193) );
  NOR3_X2 U29208 ( .A1(n15129), .A2(n61392), .A3(n21190), .ZN(n15127) );
  INV_X1 U29219 ( .I(n51119), .ZN(n63025) );
  INV_X1 U29222 ( .I(n63025), .ZN(n63026) );
  NAND2_X1 U29228 ( .A1(n13939), .A2(n53901), .ZN(n53966) );
  INV_X1 U29229 ( .I(n53901), .ZN(n6134) );
  INV_X1 U29237 ( .I(n39935), .ZN(n24002) );
  NAND2_X1 U29240 ( .A1(n25173), .A2(n56431), .ZN(n24555) );
  NAND2_X1 U29249 ( .A1(n16771), .A2(n16768), .ZN(n53326) );
  INV_X1 U29251 ( .I(n26447), .ZN(n1360) );
  BUF_X2 U29265 ( .I(n26447), .Z(n1575) );
  NAND2_X1 U29276 ( .A1(n10986), .A2(n34156), .ZN(n33356) );
  NOR2_X1 U29277 ( .A1(n34150), .A2(n10986), .ZN(n33672) );
  NAND2_X1 U29278 ( .A1(n20923), .A2(n10986), .ZN(n60801) );
  INV_X1 U29279 ( .I(n10986), .ZN(n21020) );
  CLKBUF_X12 U29283 ( .I(n20902), .Z(n10172) );
  NAND2_X1 U29284 ( .A1(n49767), .A2(n49779), .ZN(n4258) );
  OR2_X2 U29292 ( .A1(n49779), .A2(n21623), .Z(n47976) );
  OR2_X2 U29293 ( .A1(n2456), .A2(n2455), .Z(n63027) );
  XOR2_X1 U29299 ( .A1(n25257), .A2(n7711), .Z(n63028) );
  INV_X2 U29301 ( .I(n52828), .ZN(n12777) );
  INV_X1 U29314 ( .I(n32003), .ZN(n63029) );
  INV_X2 U29317 ( .I(n48883), .ZN(n24073) );
  NAND2_X1 U29320 ( .A1(n48883), .A2(n22819), .ZN(n49694) );
  BUF_X2 U29321 ( .I(n48883), .Z(n9863) );
  NAND2_X1 U29330 ( .A1(n48883), .A2(n49701), .ZN(n48897) );
  CLKBUF_X12 U29344 ( .I(n1346), .Z(n23826) );
  OR2_X2 U29345 ( .A1(n54292), .A2(n13184), .Z(n54300) );
  NAND2_X1 U29347 ( .A1(n540), .A2(n54798), .ZN(n58088) );
  NAND2_X1 U29349 ( .A1(n65276), .A2(n49379), .ZN(n2246) );
  INV_X2 U29350 ( .I(n65276), .ZN(n49433) );
  OR2_X2 U29359 ( .A1(n6015), .A2(n47873), .Z(n7622) );
  OR2_X2 U29365 ( .A1(n6015), .A2(n49538), .Z(n49546) );
  CLKBUF_X12 U29367 ( .I(n25111), .Z(n23369) );
  INV_X1 U29371 ( .I(n15414), .ZN(n17633) );
  AOI21_X1 U29384 ( .A1(n30822), .A2(n29238), .B(n58092), .ZN(n26512) );
  NOR2_X1 U29390 ( .A1(n3325), .A2(n34275), .ZN(n34274) );
  NOR2_X1 U29393 ( .A1(n40727), .A2(n57462), .ZN(n40731) );
  BUF_X2 U29403 ( .I(n45015), .Z(n3750) );
  CLKBUF_X4 U29406 ( .I(n25042), .Z(n4901) );
  INV_X1 U29407 ( .I(n22343), .ZN(n17798) );
  NAND3_X1 U29413 ( .A1(n14552), .A2(n54583), .A3(n54581), .ZN(n63155) );
  CLKBUF_X4 U29430 ( .I(n52476), .Z(n54997) );
  NAND2_X1 U29431 ( .A1(n46011), .A2(n20622), .ZN(n63031) );
  AND2_X2 U29436 ( .A1(n46010), .A2(n46009), .Z(n20622) );
  INV_X1 U29439 ( .I(n63031), .ZN(n8063) );
  INV_X1 U29453 ( .I(n50037), .ZN(n65248) );
  NOR2_X2 U29456 ( .A1(n58918), .A2(n42905), .ZN(n42907) );
  NAND2_X1 U29460 ( .A1(n57053), .A2(n57052), .ZN(n57054) );
  INV_X2 U29462 ( .I(n36517), .ZN(n37376) );
  CLKBUF_X4 U29463 ( .I(n36517), .Z(n592) );
  CLKBUF_X4 U29464 ( .I(n22683), .Z(n55225) );
  INV_X2 U29465 ( .I(n48790), .ZN(n18464) );
  CLKBUF_X4 U29468 ( .I(n48790), .Z(n6633) );
  CLKBUF_X4 U29470 ( .I(n18342), .Z(n21142) );
  INV_X1 U29473 ( .I(n20800), .ZN(n64604) );
  INV_X1 U29477 ( .I(n54814), .ZN(n54440) );
  INV_X1 U29483 ( .I(n52596), .ZN(n64628) );
  INV_X2 U29484 ( .I(n23371), .ZN(n50683) );
  NOR2_X1 U29485 ( .A1(n10294), .A2(n41382), .ZN(n41392) );
  NAND2_X1 U29487 ( .A1(n5585), .A2(n56881), .ZN(n56839) );
  NAND2_X1 U29494 ( .A1(n61221), .A2(n60708), .ZN(n56841) );
  NAND2_X1 U29498 ( .A1(n56881), .A2(n56844), .ZN(n56846) );
  NAND2_X1 U29503 ( .A1(n56196), .A2(n56189), .ZN(n56157) );
  NOR2_X1 U29505 ( .A1(n56196), .A2(n56189), .ZN(n56160) );
  NAND2_X1 U29509 ( .A1(n47252), .A2(n47251), .ZN(n47253) );
  CLKBUF_X4 U29514 ( .I(n54317), .Z(n21135) );
  XOR2_X1 U29515 ( .A1(n14128), .A2(n52569), .Z(n63033) );
  XOR2_X1 U29526 ( .A1(n8123), .A2(n63749), .Z(n63034) );
  NAND2_X1 U29530 ( .A1(n54281), .A2(n54272), .ZN(n60742) );
  NAND2_X1 U29539 ( .A1(n54266), .A2(n54272), .ZN(n54232) );
  BUF_X2 U29541 ( .I(n40550), .Z(n42139) );
  AOI21_X1 U29546 ( .A1(n23113), .A2(n63953), .B(n57234), .ZN(n63310) );
  BUF_X2 U29547 ( .I(n38529), .Z(n40971) );
  INV_X1 U29549 ( .I(n57143), .ZN(n18807) );
  NAND4_X1 U29559 ( .A1(n57154), .A2(n57143), .A3(n21569), .A4(n21829), .ZN(
        n63576) );
  BUF_X4 U29563 ( .I(n29392), .Z(n31241) );
  INV_X1 U29573 ( .I(n29392), .ZN(n31246) );
  NOR2_X1 U29574 ( .A1(n33698), .A2(n32808), .ZN(n32812) );
  NAND2_X1 U29580 ( .A1(n43325), .A2(n1298), .ZN(n42772) );
  INV_X1 U29581 ( .I(n3717), .ZN(n25769) );
  INV_X1 U29586 ( .I(n64039), .ZN(n44307) );
  CLKBUF_X4 U29589 ( .I(n11252), .Z(n8214) );
  BUF_X2 U29592 ( .I(Key[116]), .Z(n55546) );
  NAND2_X1 U29599 ( .A1(n60527), .A2(n35705), .ZN(n5999) );
  NOR2_X2 U29600 ( .A1(n7243), .A2(n63509), .ZN(n7242) );
  AND2_X2 U29602 ( .A1(n21385), .A2(n21382), .Z(n63036) );
  XNOR2_X1 U29609 ( .A1(n52623), .A2(n9230), .ZN(n25150) );
  INV_X2 U29613 ( .I(n19770), .ZN(n3246) );
  NAND2_X1 U29614 ( .A1(n49498), .A2(n49496), .ZN(n49482) );
  OR2_X2 U29623 ( .A1(n61728), .A2(n48682), .Z(n47919) );
  NOR2_X1 U29631 ( .A1(n13037), .A2(n43889), .ZN(n13036) );
  INV_X1 U29633 ( .I(n13037), .ZN(n43893) );
  OAI21_X1 U29635 ( .A1(n2797), .A2(n20183), .B(n13037), .ZN(n43236) );
  NAND2_X1 U29640 ( .A1(n57050), .A2(n57039), .ZN(n57041) );
  NAND3_X1 U29644 ( .A1(n52818), .A2(n57051), .A3(n57050), .ZN(n57053) );
  NAND2_X1 U29645 ( .A1(n8195), .A2(n4512), .ZN(n37410) );
  CLKBUF_X4 U29648 ( .I(n4512), .Z(n37404) );
  OR2_X2 U29656 ( .A1(n65222), .A2(n47055), .Z(n49018) );
  NAND2_X1 U29675 ( .A1(n1281), .A2(n53108), .ZN(n23274) );
  NAND2_X1 U29681 ( .A1(n61561), .A2(n14512), .ZN(n14985) );
  OAI21_X1 U29689 ( .A1(n62784), .A2(n26665), .B(n26660), .ZN(n13378) );
  INV_X1 U29690 ( .I(n49076), .ZN(n63200) );
  INV_X2 U29692 ( .I(n49076), .ZN(n8298) );
  CLKBUF_X4 U29697 ( .I(n26014), .Z(n15520) );
  NOR2_X1 U29699 ( .A1(n53165), .A2(n9187), .ZN(n63812) );
  AOI21_X1 U29710 ( .A1(n52229), .A2(n25484), .B(n9187), .ZN(n3537) );
  INV_X1 U29713 ( .I(n26071), .ZN(n13837) );
  OR2_X2 U29716 ( .A1(n26071), .A2(n26070), .Z(n10983) );
  CLKBUF_X12 U29719 ( .I(n26071), .Z(n20738) );
  NAND2_X1 U29722 ( .A1(n41429), .A2(n357), .ZN(n40381) );
  INV_X1 U29730 ( .I(n58896), .ZN(n54537) );
  NOR2_X1 U29732 ( .A1(n58896), .A2(n54546), .ZN(n65013) );
  BUF_X2 U29735 ( .I(n58896), .Z(n54582) );
  NAND2_X1 U29738 ( .A1(n36838), .A2(n36847), .ZN(n36012) );
  INV_X1 U29739 ( .I(n11187), .ZN(n40666) );
  INV_X1 U29740 ( .I(n34588), .ZN(n10134) );
  INV_X2 U29747 ( .I(n35427), .ZN(n1421) );
  NAND4_X1 U29751 ( .A1(n1477), .A2(n13413), .A3(n24367), .A4(n62230), .ZN(
        n63859) );
  OAI21_X1 U29753 ( .A1(n60615), .A2(n30442), .B(n60614), .ZN(n29420) );
  XOR2_X1 U29755 ( .A1(n63096), .A2(n19055), .Z(n63037) );
  XNOR2_X1 U29758 ( .A1(n61077), .A2(n859), .ZN(n63038) );
  NAND3_X2 U29761 ( .A1(n56277), .A2(n25411), .A3(n25410), .ZN(n63039) );
  AOI21_X2 U29762 ( .A1(n56223), .A2(n51110), .B(n56222), .ZN(n56277) );
  CLKBUF_X8 U29767 ( .I(n12960), .Z(n1714) );
  NOR2_X1 U29768 ( .A1(n23108), .A2(n41402), .ZN(n14286) );
  INV_X1 U29776 ( .I(n23108), .ZN(n41235) );
  OAI22_X1 U29781 ( .A1(n41403), .A2(n23108), .B1(n41402), .B2(n41410), .ZN(
        n63839) );
  AND2_X2 U29782 ( .A1(n25677), .A2(n34575), .Z(n36310) );
  INV_X1 U29783 ( .I(n46874), .ZN(n46039) );
  CLKBUF_X4 U29785 ( .I(n6015), .Z(n18769) );
  INV_X1 U29789 ( .I(n48729), .ZN(n63831) );
  NAND2_X1 U29792 ( .A1(n64462), .A2(n43504), .ZN(n42040) );
  INV_X1 U29793 ( .I(n25432), .ZN(n2218) );
  AOI22_X1 U29794 ( .A1(n64935), .A2(n49700), .B1(n58306), .B2(n48350), .ZN(
        n48352) );
  NAND4_X1 U29796 ( .A1(n49703), .A2(n22646), .A3(n49700), .A4(n49702), .ZN(
        n49704) );
  INV_X1 U29797 ( .I(n19049), .ZN(n14333) );
  BUF_X2 U29801 ( .I(n19049), .Z(n14332) );
  XOR2_X1 U29802 ( .A1(n43453), .A2(n46495), .Z(n63040) );
  CLKBUF_X12 U29805 ( .I(n18119), .Z(n58755) );
  XNOR2_X1 U29806 ( .A1(n22922), .A2(n64370), .ZN(n63041) );
  XOR2_X1 U29811 ( .A1(n32488), .A2(n32487), .Z(n63042) );
  BUF_X4 U29814 ( .I(n39081), .Z(n42788) );
  INV_X2 U29815 ( .I(n56215), .ZN(n60129) );
  NOR2_X1 U29817 ( .A1(n61260), .A2(n29187), .ZN(n59883) );
  INV_X2 U29821 ( .I(n29187), .ZN(n27282) );
  BUF_X2 U29828 ( .I(n6721), .Z(n6360) );
  CLKBUF_X2 U29834 ( .I(n27559), .Z(n25807) );
  CLKBUF_X12 U29848 ( .I(n19645), .Z(n58064) );
  INV_X2 U29850 ( .I(n28546), .ZN(n30348) );
  BUF_X4 U29851 ( .I(n28546), .Z(n30343) );
  INV_X2 U29854 ( .I(n1200), .ZN(n23070) );
  AOI21_X2 U29855 ( .A1(n43198), .A2(n43197), .B(n63044), .ZN(n46332) );
  AND2_X1 U29865 ( .A1(n43517), .A2(n43521), .Z(n63044) );
  NAND2_X2 U29866 ( .A1(n48273), .A2(n48272), .ZN(n13387) );
  AOI21_X2 U29867 ( .A1(n63960), .A2(n63961), .B(n51777), .ZN(n58083) );
  NOR2_X2 U29871 ( .A1(n22121), .A2(n17215), .ZN(n8443) );
  BUF_X4 U29873 ( .I(n22903), .Z(n64589) );
  XOR2_X1 U29874 ( .A1(n31911), .A2(n30897), .Z(n33070) );
  NOR2_X1 U29875 ( .A1(n63761), .A2(n58399), .ZN(n57322) );
  INV_X2 U29876 ( .I(n22819), .ZN(n49702) );
  NAND3_X2 U29877 ( .A1(n14235), .A2(n14236), .A3(n45666), .ZN(n22819) );
  NOR2_X2 U29883 ( .A1(n63046), .A2(n63045), .ZN(n11410) );
  NAND2_X2 U29885 ( .A1(n23333), .A2(n35960), .ZN(n63045) );
  INV_X2 U29888 ( .I(n63047), .ZN(n24293) );
  XOR2_X1 U29892 ( .A1(n639), .A2(n43425), .Z(n46668) );
  AND2_X1 U29896 ( .A1(n63048), .A2(n34711), .Z(n21501) );
  AOI22_X2 U29897 ( .A1(n36200), .A2(n36199), .B1(n36198), .B2(n36197), .ZN(
        n63049) );
  AOI21_X1 U29900 ( .A1(n29131), .A2(n29130), .B(n29129), .ZN(n63069) );
  XOR2_X1 U29901 ( .A1(n11442), .A2(n52369), .Z(n52059) );
  XOR2_X1 U29903 ( .A1(n25158), .A2(n61137), .Z(n52369) );
  AND2_X1 U29907 ( .A1(n30832), .A2(n31357), .Z(n34523) );
  NAND2_X2 U29908 ( .A1(n47518), .A2(n44670), .ZN(n47494) );
  XOR2_X1 U29916 ( .A1(n51625), .A2(n50949), .Z(n51662) );
  NAND2_X2 U29919 ( .A1(n12604), .A2(n48827), .ZN(n50949) );
  NAND2_X2 U29924 ( .A1(n56436), .A2(n1616), .ZN(n21081) );
  INV_X1 U29929 ( .I(n61731), .ZN(n25972) );
  INV_X1 U29936 ( .I(n25333), .ZN(n63051) );
  AOI21_X2 U29938 ( .A1(n47776), .A2(n7161), .B(n63052), .ZN(n13840) );
  NAND3_X2 U29939 ( .A1(n44554), .A2(n64296), .A3(n46037), .ZN(n63052) );
  XOR2_X1 U29945 ( .A1(n12578), .A2(n5952), .Z(n5951) );
  NAND2_X2 U29946 ( .A1(n10567), .A2(n1930), .ZN(n63053) );
  AOI22_X2 U29947 ( .A1(n48025), .A2(n63054), .B1(n61083), .B2(n48319), .ZN(
        n13785) );
  XOR2_X1 U29950 ( .A1(n12297), .A2(n12298), .Z(n12296) );
  AND2_X2 U29953 ( .A1(n48338), .A2(n44558), .Z(n48332) );
  NAND2_X2 U29957 ( .A1(n508), .A2(n23643), .ZN(n46941) );
  AND2_X1 U29959 ( .A1(n38201), .A2(n64017), .Z(n63640) );
  NOR3_X2 U29967 ( .A1(n11024), .A2(n33702), .A3(n33693), .ZN(n33567) );
  NAND3_X2 U29972 ( .A1(n10694), .A2(n61853), .A3(n15356), .ZN(n63509) );
  AND2_X1 U29978 ( .A1(n35236), .A2(n63055), .Z(n25450) );
  NAND2_X1 U29980 ( .A1(n35232), .A2(n35837), .ZN(n63055) );
  NAND3_X2 U29981 ( .A1(n31269), .A2(n31159), .A3(n31267), .ZN(n29920) );
  NAND2_X1 U29992 ( .A1(n2851), .A2(n53998), .ZN(n54010) );
  AND2_X1 U29993 ( .A1(n33695), .A2(n63185), .Z(n20761) );
  XOR2_X1 U29996 ( .A1(n63056), .A2(n11650), .Z(n25679) );
  XOR2_X1 U30000 ( .A1(n57714), .A2(n63028), .Z(n63056) );
  AND3_X1 U30001 ( .A1(n46901), .A2(n46902), .A3(n46903), .Z(n63057) );
  OAI21_X1 U30002 ( .A1(n63058), .A2(n5431), .B(n5360), .ZN(n5359) );
  NAND2_X2 U30005 ( .A1(n2036), .A2(n18468), .ZN(n6588) );
  NOR2_X2 U30014 ( .A1(n63059), .A2(n63811), .ZN(n47055) );
  NOR2_X2 U30016 ( .A1(n33702), .A2(n32806), .ZN(n33698) );
  NOR2_X2 U30018 ( .A1(n23064), .A2(n63060), .ZN(n23211) );
  AOI21_X2 U30020 ( .A1(n9167), .A2(n9168), .B(n61942), .ZN(n63060) );
  NOR2_X2 U30030 ( .A1(n58917), .A2(n63061), .ZN(n58368) );
  NAND2_X1 U30032 ( .A1(n33344), .A2(n63064), .ZN(n63063) );
  XOR2_X1 U30036 ( .A1(n63065), .A2(n19228), .Z(n52187) );
  XOR2_X1 U30038 ( .A1(n6725), .A2(n10101), .Z(n63065) );
  XOR2_X1 U30039 ( .A1(n19419), .A2(n63066), .Z(n3178) );
  XOR2_X1 U30040 ( .A1(n61843), .A2(n10654), .Z(n63066) );
  XOR2_X1 U30046 ( .A1(n23451), .A2(n33075), .Z(n33077) );
  XOR2_X1 U30047 ( .A1(n26178), .A2(n63067), .Z(n2975) );
  XOR2_X1 U30051 ( .A1(n8464), .A2(n64593), .Z(n63067) );
  NAND3_X2 U30057 ( .A1(n1393), .A2(n42689), .A3(n42703), .ZN(n41526) );
  NOR2_X2 U30069 ( .A1(n2766), .A2(n47467), .ZN(n65224) );
  NOR2_X1 U30071 ( .A1(n48019), .A2(n49547), .ZN(n64725) );
  NAND2_X2 U30075 ( .A1(n49556), .A2(n49565), .ZN(n49547) );
  NAND2_X1 U30083 ( .A1(n35311), .A2(n18368), .ZN(n60452) );
  NOR2_X2 U30085 ( .A1(n25806), .A2(n43449), .ZN(n42365) );
  NAND2_X2 U30087 ( .A1(n63070), .A2(n10490), .ZN(n49171) );
  NAND2_X1 U30088 ( .A1(n19605), .A2(n47853), .ZN(n63070) );
  XOR2_X1 U30096 ( .A1(n21488), .A2(n63071), .Z(n34317) );
  XOR2_X1 U30099 ( .A1(n23735), .A2(n16360), .Z(n63071) );
  BUF_X2 U30101 ( .I(n2287), .Z(n63072) );
  NAND3_X2 U30102 ( .A1(n45654), .A2(n6248), .A3(n46862), .ZN(n63816) );
  NAND2_X2 U30103 ( .A1(n64563), .A2(n16540), .ZN(n61436) );
  NAND2_X2 U30106 ( .A1(n15740), .A2(n25078), .ZN(n18878) );
  XOR2_X1 U30109 ( .A1(n64165), .A2(n24599), .Z(n25078) );
  NOR2_X2 U30111 ( .A1(n19210), .A2(n63074), .ZN(n40020) );
  NAND4_X2 U30113 ( .A1(n40009), .A2(n40006), .A3(n40008), .A4(n40007), .ZN(
        n63074) );
  XOR2_X1 U30118 ( .A1(n33877), .A2(n2290), .Z(n13195) );
  NAND2_X1 U30119 ( .A1(n41465), .A2(n41464), .ZN(n63674) );
  XOR2_X1 U30120 ( .A1(n52059), .A2(n52055), .Z(n59075) );
  INV_X2 U30125 ( .I(n61572), .ZN(n63075) );
  OR3_X1 U30126 ( .A1(n52696), .A2(n63075), .A3(n22114), .Z(n52263) );
  XOR2_X1 U30127 ( .A1(n13613), .A2(n63040), .Z(n58762) );
  XOR2_X1 U30128 ( .A1(n63076), .A2(n21422), .Z(n25649) );
  XOR2_X1 U30133 ( .A1(n63851), .A2(n1463), .Z(n63076) );
  OR2_X2 U30137 ( .A1(n45551), .A2(n21530), .Z(n47580) );
  NAND4_X2 U30140 ( .A1(n36242), .A2(n60492), .A3(n36240), .A4(n36241), .ZN(
        n39543) );
  NAND2_X1 U30149 ( .A1(n63641), .A2(n17773), .ZN(n3387) );
  NAND4_X2 U30155 ( .A1(n24810), .A2(n56154), .A3(n56153), .A4(n24809), .ZN(
        n64999) );
  NOR2_X2 U30157 ( .A1(n63079), .A2(n63078), .ZN(n63077) );
  NOR2_X1 U30158 ( .A1(n36337), .A2(n24725), .ZN(n24720) );
  INV_X4 U30161 ( .I(n63080), .ZN(n15928) );
  NOR2_X2 U30167 ( .A1(n52994), .A2(n52995), .ZN(n63080) );
  NAND3_X2 U30170 ( .A1(n10515), .A2(n52677), .A3(n52678), .ZN(n52679) );
  NAND2_X1 U30173 ( .A1(n17775), .A2(n9593), .ZN(n36046) );
  NAND2_X2 U30176 ( .A1(n60391), .A2(n64344), .ZN(n17775) );
  NAND3_X1 U30182 ( .A1(n40412), .A2(n8942), .A3(n40411), .ZN(n8941) );
  NOR2_X2 U30185 ( .A1(n23349), .A2(n6615), .ZN(n28776) );
  NOR2_X2 U30186 ( .A1(n13810), .A2(n61383), .ZN(n23349) );
  BUF_X2 U30190 ( .I(n38334), .Z(n63081) );
  XOR2_X1 U30191 ( .A1(n33885), .A2(n33884), .Z(n22661) );
  XOR2_X1 U30195 ( .A1(n33143), .A2(n33142), .Z(n33885) );
  NAND3_X2 U30198 ( .A1(n49025), .A2(n50081), .A3(n20174), .ZN(n46722) );
  NOR2_X2 U30206 ( .A1(n22764), .A2(n25944), .ZN(n49025) );
  NAND2_X2 U30207 ( .A1(n9837), .A2(n46726), .ZN(n25549) );
  NAND3_X1 U30211 ( .A1(n45622), .A2(n45621), .A3(n63294), .ZN(n63698) );
  XOR2_X1 U30217 ( .A1(n46410), .A2(n24798), .Z(n59045) );
  NAND2_X2 U30223 ( .A1(n29211), .A2(n8946), .ZN(n30234) );
  BUF_X2 U30226 ( .I(n50407), .Z(n63084) );
  XOR2_X1 U30228 ( .A1(n22662), .A2(n12872), .Z(n6570) );
  XOR2_X1 U30229 ( .A1(n63102), .A2(n20713), .Z(n12872) );
  BUF_X2 U30232 ( .I(n59138), .Z(n63085) );
  OR2_X2 U30233 ( .A1(n62353), .A2(n41568), .Z(n7877) );
  XOR2_X1 U30234 ( .A1(n63086), .A2(n11233), .Z(n34521) );
  XOR2_X1 U30235 ( .A1(n2892), .A2(n19362), .Z(n63086) );
  XOR2_X1 U30242 ( .A1(n25144), .A2(n25142), .Z(n647) );
  NAND3_X2 U30243 ( .A1(n47079), .A2(n63105), .A3(n2499), .ZN(n47082) );
  NOR2_X2 U30247 ( .A1(n48135), .A2(n22574), .ZN(n63105) );
  NOR2_X2 U30251 ( .A1(n635), .A2(n63087), .ZN(n60884) );
  AND2_X1 U30258 ( .A1(n63089), .A2(n47049), .Z(n21564) );
  OAI21_X1 U30262 ( .A1(n48393), .A2(n48859), .B(n49487), .ZN(n63089) );
  NAND2_X2 U30265 ( .A1(n7165), .A2(n40749), .ZN(n40747) );
  XOR2_X1 U30267 ( .A1(n63090), .A2(n8125), .Z(n4930) );
  XOR2_X1 U30270 ( .A1(n12040), .A2(n58055), .Z(n63090) );
  NAND2_X2 U30271 ( .A1(n3327), .A2(n2557), .ZN(n63091) );
  OAI21_X2 U30272 ( .A1(n63093), .A2(n63092), .B(n39784), .ZN(n18745) );
  XOR2_X1 U30273 ( .A1(n25740), .A2(n61938), .Z(n63505) );
  NOR2_X1 U30277 ( .A1(n64148), .A2(n11864), .ZN(n64763) );
  XOR2_X1 U30279 ( .A1(n62183), .A2(n61137), .Z(n13364) );
  XOR2_X1 U30294 ( .A1(n63096), .A2(n19055), .Z(n20953) );
  XOR2_X1 U30301 ( .A1(n19362), .A2(n13064), .Z(n63096) );
  XOR2_X1 U30311 ( .A1(n32186), .A2(n11485), .Z(n11484) );
  NAND2_X2 U30329 ( .A1(n5877), .A2(n5875), .ZN(n32186) );
  NOR2_X1 U30331 ( .A1(n22957), .A2(n27165), .ZN(n63320) );
  NOR2_X2 U30332 ( .A1(n63097), .A2(n29486), .ZN(n8586) );
  BUF_X2 U30333 ( .I(n20721), .Z(n63100) );
  NAND3_X1 U30334 ( .A1(n43224), .A2(n43223), .A3(n2464), .ZN(n2463) );
  NOR2_X2 U30338 ( .A1(n42407), .A2(n42404), .ZN(n42401) );
  NAND2_X2 U30342 ( .A1(n40347), .A2(n40348), .ZN(n63101) );
  NOR2_X2 U30344 ( .A1(n4317), .A2(n4318), .ZN(n11595) );
  NAND2_X2 U30348 ( .A1(n63103), .A2(n33540), .ZN(n14269) );
  NOR2_X2 U30351 ( .A1(n20461), .A2(n21071), .ZN(n49065) );
  XOR2_X1 U30353 ( .A1(n2364), .A2(n32186), .Z(n59911) );
  NAND2_X2 U30354 ( .A1(n62808), .A2(n25413), .ZN(n56629) );
  NAND2_X2 U30358 ( .A1(n1416), .A2(n21921), .ZN(n63742) );
  XOR2_X1 U30363 ( .A1(n8109), .A2(n59909), .Z(n32615) );
  NAND3_X2 U30367 ( .A1(n64983), .A2(n64982), .A3(n30514), .ZN(n8109) );
  NAND4_X2 U30368 ( .A1(n61620), .A2(n55312), .A3(n55311), .A4(n15100), .ZN(
        n61286) );
  NOR2_X2 U30371 ( .A1(n19000), .A2(n20888), .ZN(n43173) );
  NOR2_X2 U30373 ( .A1(n21570), .A2(n57015), .ZN(n57143) );
  AND2_X1 U30377 ( .A1(n63106), .A2(n17874), .Z(n11171) );
  XOR2_X1 U30378 ( .A1(n38403), .A2(n59751), .Z(n36104) );
  XOR2_X1 U30380 ( .A1(n3717), .A2(n26146), .Z(n38403) );
  OAI21_X2 U30381 ( .A1(n63109), .A2(n17298), .B(n14024), .ZN(n21921) );
  NOR3_X2 U30392 ( .A1(n17297), .A2(n17474), .A3(n21766), .ZN(n63109) );
  NAND3_X2 U30393 ( .A1(n339), .A2(n8120), .A3(n7588), .ZN(n50210) );
  NAND2_X1 U30401 ( .A1(n42195), .A2(n42198), .ZN(n63257) );
  XOR2_X1 U30402 ( .A1(n59926), .A2(n37939), .Z(n11056) );
  XOR2_X1 U30404 ( .A1(n64244), .A2(n37802), .Z(n37939) );
  NAND3_X1 U30412 ( .A1(n45172), .A2(n48894), .A3(n49757), .ZN(n63110) );
  XOR2_X1 U30415 ( .A1(n11426), .A2(n14106), .Z(n4844) );
  XOR2_X1 U30419 ( .A1(n9664), .A2(n12419), .Z(n14106) );
  XOR2_X1 U30421 ( .A1(n63111), .A2(n772), .Z(n6245) );
  XOR2_X1 U30425 ( .A1(n8882), .A2(n4917), .Z(n63111) );
  OR2_X1 U30431 ( .A1(n42936), .A2(n57197), .Z(n24086) );
  NAND3_X1 U30432 ( .A1(n7610), .A2(n33795), .A3(n64272), .ZN(n63313) );
  NOR3_X2 U30433 ( .A1(n30826), .A2(n30827), .A3(n63112), .ZN(n30828) );
  NAND3_X2 U30447 ( .A1(n26138), .A2(n18904), .A3(n18906), .ZN(n63112) );
  NOR3_X2 U30449 ( .A1(n18018), .A2(n18344), .A3(n42408), .ZN(n15117) );
  XOR2_X1 U30451 ( .A1(n8419), .A2(n64837), .Z(n20580) );
  NOR2_X2 U30458 ( .A1(n64396), .A2(n992), .ZN(n57689) );
  NOR2_X2 U30459 ( .A1(n2418), .A2(n21467), .ZN(n36211) );
  XOR2_X1 U30466 ( .A1(n37886), .A2(n63113), .Z(n61478) );
  XOR2_X1 U30468 ( .A1(n64325), .A2(n6703), .Z(n63113) );
  XOR2_X1 U30474 ( .A1(n24152), .A2(n63114), .Z(n26142) );
  NOR2_X2 U30477 ( .A1(n63115), .A2(n37317), .ZN(n37948) );
  OAI21_X1 U30483 ( .A1(n25445), .A2(n24596), .B(n5846), .ZN(n24595) );
  BUF_X2 U30494 ( .I(n10134), .Z(n63116) );
  AOI22_X2 U30497 ( .A1(n17244), .A2(n43565), .B1(n17245), .B2(n17246), .ZN(
        n63117) );
  AND2_X2 U30500 ( .A1(n13195), .A2(n35738), .Z(n35750) );
  INV_X1 U30505 ( .I(n50264), .ZN(n63183) );
  NOR2_X2 U30508 ( .A1(n1815), .A2(n24871), .ZN(n32975) );
  OAI21_X2 U30513 ( .A1(n14550), .A2(n61944), .B(n63118), .ZN(n15189) );
  NOR2_X2 U30515 ( .A1(n16653), .A2(n16652), .ZN(n14550) );
  NAND4_X2 U30516 ( .A1(n18776), .A2(n18775), .A3(n18777), .A4(n63120), .ZN(
        n11311) );
  NOR2_X1 U30517 ( .A1(n34854), .A2(n63121), .ZN(n34006) );
  AND2_X1 U30519 ( .A1(n34009), .A2(n36777), .Z(n63121) );
  AOI21_X1 U30522 ( .A1(n35163), .A2(n7655), .B(n35165), .ZN(n24150) );
  NAND3_X2 U30534 ( .A1(n42100), .A2(n42918), .A3(n42919), .ZN(n41598) );
  XOR2_X1 U30536 ( .A1(n24739), .A2(n51044), .Z(n63149) );
  OAI21_X2 U30537 ( .A1(n9849), .A2(n9850), .B(n62001), .ZN(n42948) );
  XOR2_X1 U30538 ( .A1(n63570), .A2(n63124), .Z(n47819) );
  XOR2_X1 U30539 ( .A1(n24020), .A2(n45004), .Z(n63124) );
  NAND3_X2 U30542 ( .A1(n11987), .A2(n30481), .A3(n60284), .ZN(n27754) );
  AOI21_X1 U30546 ( .A1(n14506), .A2(n42082), .B(n41689), .ZN(n25578) );
  NAND3_X2 U30547 ( .A1(n57495), .A2(n52263), .A3(n52262), .ZN(n20489) );
  NOR2_X1 U30548 ( .A1(n63125), .A2(n20200), .ZN(n63536) );
  AND2_X1 U30553 ( .A1(n20201), .A2(n5684), .Z(n63125) );
  XOR2_X1 U30554 ( .A1(n4041), .A2(n52148), .Z(n57486) );
  XOR2_X1 U30559 ( .A1(n45409), .A2(n14155), .Z(n14154) );
  XOR2_X1 U30560 ( .A1(n15173), .A2(n5358), .Z(n45409) );
  XOR2_X1 U30563 ( .A1(n61672), .A2(n14153), .Z(n45411) );
  NAND2_X1 U30575 ( .A1(n21536), .A2(n23226), .ZN(n37291) );
  INV_X2 U30578 ( .I(n63127), .ZN(n17240) );
  INV_X1 U30585 ( .I(n21983), .ZN(n63128) );
  NOR3_X2 U30587 ( .A1(n10794), .A2(n37293), .A3(n22659), .ZN(n4914) );
  NAND2_X2 U30588 ( .A1(n20124), .A2(n21536), .ZN(n10794) );
  OR2_X1 U30591 ( .A1(n42240), .A2(n41915), .Z(n64972) );
  AOI21_X1 U30592 ( .A1(n30285), .A2(n30264), .B(n30286), .ZN(n63129) );
  NOR2_X1 U30596 ( .A1(n9863), .A2(n49700), .ZN(n1104) );
  NOR2_X2 U30600 ( .A1(n687), .A2(n22962), .ZN(n49700) );
  NAND2_X2 U30601 ( .A1(n39947), .A2(n10395), .ZN(n37663) );
  NAND3_X2 U30605 ( .A1(n23890), .A2(n39510), .A3(n64390), .ZN(n39947) );
  NAND3_X2 U30606 ( .A1(n64588), .A2(n18448), .A3(n18447), .ZN(n17984) );
  NAND2_X1 U30607 ( .A1(n64644), .A2(n48681), .ZN(n22153) );
  NAND2_X2 U30615 ( .A1(n5173), .A2(n63130), .ZN(n5194) );
  NOR2_X2 U30617 ( .A1(n55914), .A2(n14056), .ZN(n55430) );
  XOR2_X1 U30621 ( .A1(n63133), .A2(n1750), .Z(n18578) );
  INV_X2 U30622 ( .I(n58891), .ZN(n63133) );
  AOI21_X2 U30623 ( .A1(n23432), .A2(n36317), .B(n63134), .ZN(n39491) );
  NAND3_X2 U30638 ( .A1(n23320), .A2(n58873), .A3(n36315), .ZN(n63134) );
  XOR2_X1 U30641 ( .A1(n32236), .A2(n1347), .Z(n32665) );
  XOR2_X1 U30644 ( .A1(n33034), .A2(n32089), .Z(n32236) );
  NAND2_X1 U30645 ( .A1(n31606), .A2(n31605), .ZN(n19796) );
  XOR2_X1 U30646 ( .A1(n33069), .A2(n15610), .Z(n10634) );
  XOR2_X1 U30649 ( .A1(n19757), .A2(n25042), .Z(n33069) );
  NAND2_X2 U30650 ( .A1(n57165), .A2(n33972), .ZN(n34186) );
  XOR2_X1 U30651 ( .A1(n3480), .A2(n38364), .Z(n19009) );
  NOR2_X2 U30657 ( .A1(n6469), .A2(n63453), .ZN(n14964) );
  NAND3_X1 U30662 ( .A1(n42316), .A2(n42004), .A3(n43011), .ZN(n39179) );
  XOR2_X1 U30666 ( .A1(n49049), .A2(n3971), .Z(n20709) );
  NAND2_X2 U30667 ( .A1(n48682), .A2(n61728), .ZN(n49049) );
  INV_X2 U30670 ( .I(n58388), .ZN(n29236) );
  NAND2_X1 U30674 ( .A1(n58388), .A2(n65096), .ZN(n25280) );
  NAND2_X2 U30675 ( .A1(n2511), .A2(n3503), .ZN(n8599) );
  XOR2_X1 U30676 ( .A1(n33828), .A2(n15102), .Z(n14945) );
  XOR2_X1 U30685 ( .A1(n13639), .A2(n51540), .Z(n4904) );
  XOR2_X1 U30690 ( .A1(n20232), .A2(n20754), .Z(n8157) );
  BUF_X2 U30691 ( .I(n60146), .Z(n63140) );
  XOR2_X1 U30696 ( .A1(n44922), .A2(n44395), .Z(n63141) );
  NAND2_X2 U30698 ( .A1(n45532), .A2(n13655), .ZN(n45787) );
  OR2_X1 U30704 ( .A1(n42355), .A2(n41987), .Z(n3126) );
  NOR2_X2 U30705 ( .A1(n10277), .A2(n32892), .ZN(n18390) );
  NOR2_X1 U30706 ( .A1(n6162), .A2(n42364), .ZN(n64439) );
  XOR2_X1 U30714 ( .A1(n63142), .A2(n53359), .Z(Plaintext[22]) );
  NAND3_X1 U30715 ( .A1(n53357), .A2(n53358), .A3(n53356), .ZN(n63142) );
  NOR2_X2 U30718 ( .A1(n12459), .A2(n12456), .ZN(n15410) );
  OAI21_X2 U30719 ( .A1(n61438), .A2(n24033), .B(n12797), .ZN(n36969) );
  NOR2_X2 U30722 ( .A1(n10193), .A2(n64573), .ZN(n63144) );
  NAND2_X2 U30724 ( .A1(n63145), .A2(n1093), .ZN(n21623) );
  NAND2_X1 U30731 ( .A1(n57066), .A2(n57065), .ZN(n64731) );
  XOR2_X1 U30733 ( .A1(n63146), .A2(n64448), .Z(n40961) );
  XOR2_X1 U30734 ( .A1(n18966), .A2(n63934), .Z(n63146) );
  OAI21_X1 U30742 ( .A1(n63148), .A2(n20496), .B(n63147), .ZN(n20493) );
  OAI21_X1 U30743 ( .A1(n58635), .A2(n20495), .B(n43518), .ZN(n63147) );
  INV_X1 U30747 ( .I(n63153), .ZN(n4796) );
  NOR2_X2 U30756 ( .A1(n63151), .A2(n60066), .ZN(n61242) );
  NOR2_X2 U30759 ( .A1(n63959), .A2(n58209), .ZN(n63151) );
  NAND2_X2 U30767 ( .A1(n31085), .A2(n31086), .ZN(n30421) );
  AOI22_X2 U30768 ( .A1(n40292), .A2(n40291), .B1(n11940), .B2(n40300), .ZN(
        n26204) );
  NAND2_X2 U30771 ( .A1(n9092), .A2(n9090), .ZN(n40292) );
  XOR2_X1 U30773 ( .A1(n63152), .A2(n39720), .Z(n39781) );
  XOR2_X1 U30779 ( .A1(n58489), .A2(n39719), .Z(n63152) );
  NAND3_X1 U30782 ( .A1(n52676), .A2(n52674), .A3(n52675), .ZN(n52677) );
  INV_X1 U30793 ( .I(n59694), .ZN(n44504) );
  INV_X2 U30794 ( .I(n42365), .ZN(n42367) );
  AND2_X2 U30795 ( .A1(n45140), .A2(n21279), .Z(n47579) );
  INV_X1 U30796 ( .I(n65174), .ZN(n63287) );
  XOR2_X1 U30806 ( .A1(n7750), .A2(n63153), .Z(n52719) );
  NAND2_X1 U30810 ( .A1(n54527), .A2(n54520), .ZN(n63156) );
  INV_X4 U30814 ( .I(n63799), .ZN(n35273) );
  NOR2_X2 U30816 ( .A1(n63159), .A2(n63157), .ZN(n30594) );
  NAND2_X2 U30819 ( .A1(n1316), .A2(n63158), .ZN(n63157) );
  NAND2_X2 U30822 ( .A1(n48386), .A2(n49641), .ZN(n49919) );
  NAND2_X2 U30823 ( .A1(n6130), .A2(n19489), .ZN(n49641) );
  NOR2_X2 U30825 ( .A1(n37114), .A2(n37115), .ZN(n37350) );
  NAND2_X2 U30829 ( .A1(n59011), .A2(n20124), .ZN(n37114) );
  XOR2_X1 U30840 ( .A1(n21025), .A2(n20623), .Z(n33161) );
  NAND2_X2 U30844 ( .A1(n11713), .A2(n63160), .ZN(n56190) );
  NAND2_X2 U30850 ( .A1(n18496), .A2(n38551), .ZN(n19368) );
  INV_X4 U30851 ( .I(n63163), .ZN(n897) );
  NAND2_X2 U30855 ( .A1(n35272), .A2(n17240), .ZN(n63163) );
  NAND2_X2 U30858 ( .A1(n63164), .A2(n15137), .ZN(n22540) );
  NOR2_X2 U30861 ( .A1(n63165), .A2(n7468), .ZN(n63164) );
  NAND2_X2 U30866 ( .A1(n16116), .A2(n26782), .ZN(n63166) );
  NAND4_X2 U30875 ( .A1(n47033), .A2(n47031), .A3(n47030), .A4(n47032), .ZN(
        n47040) );
  NAND2_X2 U30878 ( .A1(n6006), .A2(n22881), .ZN(n6005) );
  XOR2_X1 U30890 ( .A1(n63167), .A2(n31800), .Z(n22440) );
  XOR2_X1 U30891 ( .A1(n31806), .A2(n31805), .Z(n63167) );
  NAND2_X1 U30893 ( .A1(n41194), .A2(n41188), .ZN(n41192) );
  NOR2_X2 U30899 ( .A1(n15215), .A2(n3246), .ZN(n41188) );
  AOI22_X1 U30900 ( .A1(n63168), .A2(n61878), .B1(n20121), .B2(n19887), .ZN(
        n20118) );
  NAND2_X2 U30901 ( .A1(n33573), .A2(n24006), .ZN(n12506) );
  NAND2_X2 U30902 ( .A1(n17885), .A2(n17929), .ZN(n50019) );
  NAND2_X2 U30904 ( .A1(n63169), .A2(n58208), .ZN(n51691) );
  XOR2_X1 U30906 ( .A1(n4521), .A2(n24521), .Z(n63971) );
  INV_X1 U30911 ( .I(n1386), .ZN(n63423) );
  INV_X2 U30913 ( .I(n63173), .ZN(n19935) );
  XOR2_X1 U30915 ( .A1(n19937), .A2(n19936), .Z(n63173) );
  NOR2_X2 U30918 ( .A1(n15695), .A2(n43910), .ZN(n42063) );
  INV_X2 U30922 ( .I(n42226), .ZN(n63435) );
  NAND2_X2 U30926 ( .A1(n6996), .A2(n42224), .ZN(n42226) );
  XOR2_X1 U30929 ( .A1(n61955), .A2(n45019), .Z(n15560) );
  INV_X1 U30938 ( .I(n57983), .ZN(n41513) );
  NAND2_X2 U30941 ( .A1(n61924), .A2(n61826), .ZN(n57983) );
  NOR3_X2 U30944 ( .A1(n27200), .A2(n63175), .A3(n27212), .ZN(n63242) );
  INV_X2 U30954 ( .I(n27196), .ZN(n63175) );
  NAND2_X2 U30955 ( .A1(n7974), .A2(n26682), .ZN(n27196) );
  NOR3_X2 U30956 ( .A1(n39109), .A2(n63176), .A3(n39107), .ZN(n25270) );
  AOI21_X2 U30958 ( .A1(n63483), .A2(n39104), .B(n58599), .ZN(n63176) );
  NAND2_X1 U30963 ( .A1(n57778), .A2(n57553), .ZN(n63728) );
  INV_X2 U30965 ( .I(n26111), .ZN(n64548) );
  XOR2_X1 U30966 ( .A1(n59749), .A2(n61957), .Z(n26111) );
  OAI21_X1 U30967 ( .A1(n42317), .A2(n62389), .B(n5262), .ZN(n42003) );
  NAND2_X1 U30970 ( .A1(n55831), .A2(n63177), .ZN(n12434) );
  NAND2_X2 U30971 ( .A1(n64166), .A2(n13684), .ZN(n50254) );
  XOR2_X1 U30972 ( .A1(n63179), .A2(n23893), .Z(n2275) );
  XOR2_X1 U30976 ( .A1(n12153), .A2(n1268), .Z(n63179) );
  NOR3_X2 U30983 ( .A1(n57881), .A2(n49427), .A3(n18226), .ZN(n6928) );
  NAND2_X2 U30984 ( .A1(n63181), .A2(n63180), .ZN(n24079) );
  NAND3_X1 U30985 ( .A1(n14114), .A2(n63977), .A3(n42783), .ZN(n63184) );
  INV_X4 U30987 ( .I(n63185), .ZN(n33702) );
  NOR2_X2 U30990 ( .A1(n24099), .A2(n48095), .ZN(n46817) );
  NOR2_X2 U30991 ( .A1(n63187), .A2(n29103), .ZN(n5563) );
  OAI21_X2 U30992 ( .A1(n29524), .A2(n30954), .B(n63188), .ZN(n63187) );
  NOR2_X2 U30994 ( .A1(n29102), .A2(n63189), .ZN(n63188) );
  NOR2_X2 U31000 ( .A1(n29100), .A2(n64940), .ZN(n63189) );
  XOR2_X1 U31003 ( .A1(n62455), .A2(n64805), .Z(n2213) );
  XOR2_X1 U31005 ( .A1(n18645), .A2(n11501), .Z(n51812) );
  NOR2_X2 U31009 ( .A1(n65226), .A2(n63190), .ZN(n6342) );
  OR2_X1 U31011 ( .A1(n41603), .A2(n5313), .Z(n63190) );
  NOR2_X1 U31016 ( .A1(n63499), .A2(n19392), .ZN(n45727) );
  NAND3_X2 U31019 ( .A1(n1095), .A2(n8990), .A3(n63192), .ZN(n64372) );
  NAND3_X2 U31020 ( .A1(n22651), .A2(n49841), .A3(n49840), .ZN(n51671) );
  INV_X2 U31028 ( .I(n16943), .ZN(n63193) );
  NAND2_X2 U31029 ( .A1(n17155), .A2(n63193), .ZN(n57295) );
  BUF_X2 U31030 ( .I(n19167), .Z(n63194) );
  OR2_X1 U31032 ( .A1(n39984), .A2(n39983), .Z(n63195) );
  NAND2_X2 U31038 ( .A1(n39525), .A2(n58416), .ZN(n5150) );
  NAND2_X2 U31039 ( .A1(n35484), .A2(n37960), .ZN(n39525) );
  OAI22_X2 U31044 ( .A1(n63196), .A2(n45461), .B1(n45462), .B2(n45463), .ZN(
        n24608) );
  NAND3_X2 U31046 ( .A1(n7194), .A2(n45459), .A3(n25680), .ZN(n63196) );
  INV_X2 U31051 ( .I(n48289), .ZN(n49243) );
  NAND2_X2 U31052 ( .A1(n50426), .A2(n2754), .ZN(n48289) );
  OAI22_X1 U31053 ( .A1(n15207), .A2(n21562), .B1(n27271), .B2(n27270), .ZN(
        n65174) );
  NAND2_X2 U31054 ( .A1(n22461), .A2(n37424), .ZN(n34817) );
  XOR2_X1 U31058 ( .A1(n52604), .A2(n50717), .Z(n14967) );
  NAND3_X2 U31061 ( .A1(n58541), .A2(n45709), .A3(n58540), .ZN(n52604) );
  NAND2_X2 U31068 ( .A1(n63197), .A2(n21565), .ZN(n11742) );
  NOR2_X2 U31070 ( .A1(n63198), .A2(n28095), .ZN(n29976) );
  INV_X2 U31071 ( .I(n28094), .ZN(n63198) );
  NOR2_X2 U31074 ( .A1(n1253), .A2(n15205), .ZN(n28094) );
  INV_X1 U31080 ( .I(n39990), .ZN(n63199) );
  NOR2_X1 U31086 ( .A1(n61806), .A2(n7990), .ZN(n45705) );
  OAI21_X1 U31089 ( .A1(n61521), .A2(n55389), .B(n61763), .ZN(n55391) );
  XOR2_X1 U31090 ( .A1(n2457), .A2(n39722), .Z(n63201) );
  BUF_X4 U31091 ( .I(n16982), .Z(n63205) );
  NAND2_X2 U31095 ( .A1(n38758), .A2(n6237), .ZN(n64655) );
  XOR2_X1 U31098 ( .A1(n51812), .A2(n51813), .Z(n7533) );
  OAI22_X2 U31099 ( .A1(n54225), .A2(n19404), .B1(n54214), .B2(n64075), .ZN(
        n54215) );
  OAI21_X2 U31100 ( .A1(n1309), .A2(n37451), .B(n63207), .ZN(n37452) );
  XOR2_X1 U31102 ( .A1(n46578), .A2(n63208), .Z(n20517) );
  XOR2_X1 U31108 ( .A1(n20516), .A2(n16126), .Z(n63208) );
  XOR2_X1 U31110 ( .A1(n24679), .A2(n14505), .Z(n63681) );
  NOR3_X2 U31126 ( .A1(n11503), .A2(n11504), .A3(n4425), .ZN(n14505) );
  XOR2_X1 U31128 ( .A1(n13355), .A2(n63209), .Z(n25132) );
  XOR2_X1 U31133 ( .A1(n20202), .A2(n39661), .Z(n63209) );
  NOR2_X2 U31134 ( .A1(n1381), .A2(n4174), .ZN(n46729) );
  NOR3_X1 U31138 ( .A1(n27580), .A2(n23071), .A3(n27579), .ZN(n27586) );
  XOR2_X1 U31149 ( .A1(n63210), .A2(n743), .Z(n25517) );
  XOR2_X1 U31150 ( .A1(n60148), .A2(n6035), .Z(n63210) );
  INV_X2 U31152 ( .I(n42370), .ZN(n42940) );
  NOR2_X1 U31160 ( .A1(n42372), .A2(n63211), .ZN(n42375) );
  NAND2_X1 U31171 ( .A1(n42370), .A2(n63212), .ZN(n63211) );
  NAND2_X2 U31174 ( .A1(n57528), .A2(n57197), .ZN(n42370) );
  NOR2_X2 U31175 ( .A1(n48490), .A2(n46468), .ZN(n47161) );
  NAND2_X2 U31179 ( .A1(n10815), .A2(n63214), .ZN(n19261) );
  NOR2_X2 U31186 ( .A1(n10816), .A2(n14445), .ZN(n63214) );
  INV_X2 U31192 ( .I(n63215), .ZN(n34233) );
  NOR2_X2 U31198 ( .A1(n34238), .A2(n24293), .ZN(n63215) );
  XOR2_X1 U31207 ( .A1(n63216), .A2(n63564), .Z(n25405) );
  XOR2_X1 U31209 ( .A1(n25407), .A2(n14157), .Z(n63216) );
  NAND2_X2 U31210 ( .A1(n4211), .A2(n58309), .ZN(n63218) );
  NOR2_X2 U31211 ( .A1(n25262), .A2(n63219), .ZN(n6368) );
  NAND3_X2 U31212 ( .A1(n4452), .A2(n49370), .A3(n2581), .ZN(n63219) );
  OR3_X1 U31213 ( .A1(n8981), .A2(n43105), .A3(n19591), .Z(n20639) );
  BUF_X2 U31214 ( .I(n35765), .Z(n63220) );
  XOR2_X1 U31215 ( .A1(n63221), .A2(n1337), .Z(n14158) );
  XOR2_X1 U31216 ( .A1(n1758), .A2(n39764), .Z(n63221) );
  NAND2_X2 U31217 ( .A1(n18251), .A2(n18754), .ZN(n63485) );
  NAND2_X2 U31223 ( .A1(n43571), .A2(n1397), .ZN(n41966) );
  NOR2_X2 U31225 ( .A1(n5398), .A2(n4547), .ZN(n43571) );
  NAND2_X1 U31226 ( .A1(n61877), .A2(n49205), .ZN(n63526) );
  NOR2_X1 U31227 ( .A1(n63526), .A2(n49206), .ZN(n49207) );
  XOR2_X1 U31238 ( .A1(n12173), .A2(n7557), .Z(n32281) );
  OAI21_X1 U31240 ( .A1(n25357), .A2(n39487), .B(n39504), .ZN(n63972) );
  XOR2_X1 U31247 ( .A1(n11457), .A2(n63223), .Z(n11456) );
  XOR2_X1 U31263 ( .A1(n32293), .A2(n24790), .Z(n63223) );
  NOR2_X2 U31264 ( .A1(n48597), .A2(n61212), .ZN(n63835) );
  XOR2_X1 U31284 ( .A1(n3879), .A2(n16843), .Z(n30944) );
  XOR2_X1 U31292 ( .A1(n11231), .A2(n3878), .Z(n16843) );
  NAND2_X2 U31293 ( .A1(n16937), .A2(n55231), .ZN(n60032) );
  NOR2_X2 U31315 ( .A1(n61702), .A2(n35731), .ZN(n35751) );
  AND2_X2 U31318 ( .A1(n19935), .A2(n9926), .Z(n47529) );
  NOR2_X2 U31327 ( .A1(n55470), .A2(n55728), .ZN(n55739) );
  XOR2_X1 U31343 ( .A1(n2241), .A2(n45269), .Z(n5748) );
  INV_X2 U31348 ( .I(n43998), .ZN(n2241) );
  XOR2_X1 U31349 ( .A1(n2365), .A2(n14313), .Z(n43998) );
  NOR3_X2 U31356 ( .A1(n58119), .A2(n2530), .A3(n55185), .ZN(n525) );
  NOR2_X2 U31357 ( .A1(n3631), .A2(n63226), .ZN(n10894) );
  NOR2_X2 U31360 ( .A1(n7831), .A2(n943), .ZN(n19641) );
  AND2_X1 U31361 ( .A1(n42668), .A2(n9334), .Z(n41784) );
  XOR2_X1 U31367 ( .A1(n3517), .A2(n63227), .Z(n17691) );
  XOR2_X1 U31376 ( .A1(n44957), .A2(n44956), .Z(n63227) );
  NAND2_X1 U31380 ( .A1(n47284), .A2(n63230), .ZN(n3659) );
  NAND2_X2 U31382 ( .A1(n60128), .A2(n40724), .ZN(n63228) );
  OAI21_X2 U31384 ( .A1(n64453), .A2(n24219), .B(n63229), .ZN(n55884) );
  INV_X4 U31385 ( .I(n14330), .ZN(n33642) );
  NAND2_X1 U31387 ( .A1(n48096), .A2(n63231), .ZN(n48100) );
  NAND2_X2 U31391 ( .A1(n15619), .A2(n15620), .ZN(n36394) );
  NOR2_X2 U31415 ( .A1(n10641), .A2(n63234), .ZN(n19240) );
  XOR2_X1 U31417 ( .A1(n39006), .A2(n38707), .Z(n6238) );
  XOR2_X1 U31420 ( .A1(n38828), .A2(n38709), .Z(n39006) );
  NOR2_X2 U31426 ( .A1(n1291), .A2(n60467), .ZN(n50263) );
  XOR2_X1 U31429 ( .A1(n63235), .A2(n23553), .Z(n46409) );
  XOR2_X1 U31432 ( .A1(n46691), .A2(n44627), .Z(n63235) );
  XOR2_X1 U31433 ( .A1(n63277), .A2(n51380), .Z(n7843) );
  NAND3_X2 U31435 ( .A1(n63236), .A2(n16220), .A3(n61780), .ZN(n60476) );
  BUF_X2 U31436 ( .I(n30725), .Z(n63237) );
  NAND3_X1 U31443 ( .A1(n43180), .A2(n63243), .A3(n43181), .ZN(n63239) );
  NAND2_X2 U31446 ( .A1(n440), .A2(n64114), .ZN(n38537) );
  NOR2_X2 U31449 ( .A1(n1081), .A2(n63240), .ZN(n60726) );
  NAND3_X2 U31458 ( .A1(n46962), .A2(n46952), .A3(n9078), .ZN(n63240) );
  XOR2_X1 U31460 ( .A1(n2933), .A2(n61537), .Z(n5406) );
  NOR2_X1 U31462 ( .A1(n51107), .A2(n51106), .ZN(n64227) );
  OR2_X1 U31464 ( .A1(n15040), .A2(n23849), .Z(n54658) );
  NAND3_X2 U31471 ( .A1(n63242), .A2(n24774), .A3(n63241), .ZN(n14759) );
  NAND3_X1 U31482 ( .A1(n43518), .A2(n65262), .A3(n20888), .ZN(n63243) );
  NAND3_X2 U31485 ( .A1(n15008), .A2(n25929), .A3(n15072), .ZN(n42846) );
  NOR2_X2 U31486 ( .A1(n64504), .A2(n64502), .ZN(n15008) );
  OR2_X1 U31491 ( .A1(n57010), .A2(n1153), .Z(n1154) );
  INV_X1 U31494 ( .I(n42782), .ZN(n14115) );
  OR2_X1 U31504 ( .A1(n19142), .A2(n48148), .Z(n20574) );
  NOR3_X2 U31506 ( .A1(n36463), .A2(n12967), .A3(n7933), .ZN(n932) );
  NOR3_X2 U31508 ( .A1(n50366), .A2(n63244), .A3(n50002), .ZN(n16673) );
  INV_X1 U31511 ( .I(n27763), .ZN(n29816) );
  NAND2_X1 U31514 ( .A1(n61162), .A2(n63245), .ZN(n7076) );
  NAND2_X1 U31517 ( .A1(n27763), .A2(n25527), .ZN(n63245) );
  NOR2_X2 U31522 ( .A1(n24728), .A2(n24402), .ZN(n27763) );
  NAND2_X2 U31527 ( .A1(n34984), .A2(n10091), .ZN(n63443) );
  XOR2_X1 U31530 ( .A1(n63246), .A2(n21446), .Z(n63410) );
  AND2_X2 U31531 ( .A1(n15201), .A2(n9971), .Z(n6914) );
  XOR2_X1 U31533 ( .A1(n9885), .A2(n39315), .Z(n3837) );
  NOR2_X2 U31544 ( .A1(n3313), .A2(n3314), .ZN(n39315) );
  OR2_X2 U31545 ( .A1(n40394), .A2(n15078), .Z(n7618) );
  NAND2_X1 U31550 ( .A1(n63576), .A2(n57160), .ZN(n25905) );
  NAND2_X2 U31551 ( .A1(n1663), .A2(n15360), .ZN(n15359) );
  AOI21_X2 U31553 ( .A1(n7865), .A2(n5161), .B(n5158), .ZN(n5160) );
  NOR2_X2 U31561 ( .A1(n63250), .A2(n63248), .ZN(n3432) );
  NAND2_X2 U31563 ( .A1(n2064), .A2(n63249), .ZN(n63248) );
  NOR3_X2 U31568 ( .A1(n342), .A2(n27753), .A3(n63251), .ZN(n21796) );
  AOI21_X2 U31574 ( .A1(n48100), .A2(n48101), .B(n48099), .ZN(n48107) );
  OR2_X2 U31575 ( .A1(n64869), .A2(n64267), .Z(n48575) );
  XOR2_X1 U31581 ( .A1(n45826), .A2(n63514), .Z(n10459) );
  XOR2_X1 U31583 ( .A1(n60859), .A2(n9062), .Z(n9060) );
  XOR2_X1 U31585 ( .A1(n25200), .A2(n18734), .Z(n63263) );
  NOR2_X2 U31589 ( .A1(n23348), .A2(n25685), .ZN(n64734) );
  INV_X2 U31595 ( .I(n13462), .ZN(n23348) );
  XOR2_X1 U31600 ( .A1(n8386), .A2(n19648), .Z(n13462) );
  XOR2_X1 U31601 ( .A1(n25130), .A2(n38812), .Z(n6927) );
  NAND3_X2 U31607 ( .A1(n63477), .A2(n58589), .A3(n25770), .ZN(n38812) );
  NOR2_X2 U31610 ( .A1(n24436), .A2(n24437), .ZN(n25130) );
  NAND2_X2 U31619 ( .A1(n11731), .A2(n15380), .ZN(n13393) );
  OAI22_X1 U31625 ( .A1(n27858), .A2(n13400), .B1(n27857), .B2(n27856), .ZN(
        n63252) );
  NAND2_X2 U31631 ( .A1(n58710), .A2(n60293), .ZN(n12894) );
  INV_X1 U31633 ( .I(n29694), .ZN(n27897) );
  NAND2_X2 U31637 ( .A1(n22214), .A2(n28187), .ZN(n29694) );
  OAI22_X1 U31644 ( .A1(n57001), .A2(n61572), .B1(n57390), .B2(n57002), .ZN(
        n57005) );
  NAND2_X2 U31658 ( .A1(n10237), .A2(n20156), .ZN(n57002) );
  OR2_X1 U31662 ( .A1(n63254), .A2(n21883), .Z(n4972) );
  OR2_X1 U31663 ( .A1(n36394), .A2(n63262), .Z(n36060) );
  OAI21_X1 U31665 ( .A1(n63256), .A2(n27905), .B(n63255), .ZN(n29899) );
  NAND2_X1 U31669 ( .A1(n29896), .A2(n27905), .ZN(n63255) );
  NAND2_X1 U31671 ( .A1(n63257), .A2(n641), .ZN(n63856) );
  NOR3_X2 U31673 ( .A1(n61879), .A2(n36431), .A3(n23975), .ZN(n23977) );
  NAND4_X2 U31674 ( .A1(n39514), .A2(n39515), .A3(n39513), .A4(n39949), .ZN(
        n63258) );
  NAND2_X2 U31681 ( .A1(n34350), .A2(n23281), .ZN(n2064) );
  NAND2_X2 U31682 ( .A1(n8028), .A2(n1701), .ZN(n43129) );
  NOR2_X2 U31685 ( .A1(n19255), .A2(n25349), .ZN(n30883) );
  XOR2_X1 U31688 ( .A1(n63260), .A2(n33051), .Z(n8591) );
  XOR2_X1 U31692 ( .A1(n32206), .A2(n31648), .Z(n63260) );
  NAND2_X2 U31696 ( .A1(n41645), .A2(n40844), .ZN(n41640) );
  NOR2_X2 U31700 ( .A1(n40843), .A2(n41066), .ZN(n41645) );
  NAND2_X2 U31701 ( .A1(n29241), .A2(n30817), .ZN(n30809) );
  NAND2_X2 U31703 ( .A1(n13567), .A2(n57075), .ZN(n52672) );
  XOR2_X1 U31704 ( .A1(n10057), .A2(n9166), .Z(n31456) );
  INV_X2 U31705 ( .I(n63262), .ZN(n8781) );
  XOR2_X1 U31709 ( .A1(n60701), .A2(n16317), .Z(n20886) );
  XOR2_X1 U31710 ( .A1(n25332), .A2(n32234), .Z(n26216) );
  NOR2_X2 U31711 ( .A1(n26712), .A2(n26711), .ZN(n32234) );
  OR2_X2 U31712 ( .A1(n60793), .A2(n32489), .Z(n61522) );
  NOR2_X1 U31713 ( .A1(n9593), .A2(n17775), .ZN(n35418) );
  INV_X1 U31714 ( .I(n16867), .ZN(n63266) );
  OR2_X1 U31716 ( .A1(n57072), .A2(n60934), .Z(n64342) );
  NOR2_X1 U31725 ( .A1(n63267), .A2(n14831), .ZN(n15129) );
  NAND2_X1 U31736 ( .A1(n58414), .A2(n58415), .ZN(n63267) );
  NOR2_X2 U31752 ( .A1(n25456), .A2(n63268), .ZN(n19081) );
  NOR2_X2 U31769 ( .A1(n21459), .A2(n21529), .ZN(n22045) );
  NAND2_X2 U31770 ( .A1(n20552), .A2(n1741), .ZN(n21459) );
  OAI21_X2 U31771 ( .A1(n63914), .A2(n1272), .B(n23484), .ZN(n39968) );
  XOR2_X1 U31779 ( .A1(n18091), .A2(n11323), .Z(n19753) );
  NOR3_X2 U31805 ( .A1(n63628), .A2(n4002), .A3(n4001), .ZN(n63269) );
  XOR2_X1 U31806 ( .A1(n13639), .A2(n52076), .Z(n13643) );
  XOR2_X1 U31809 ( .A1(n7860), .A2(n63024), .Z(n25378) );
  NOR2_X2 U31815 ( .A1(n8723), .A2(n8728), .ZN(n7860) );
  INV_X1 U31824 ( .I(n19206), .ZN(n63582) );
  NAND2_X2 U31829 ( .A1(n8303), .A2(n38345), .ZN(n16526) );
  NAND2_X2 U31834 ( .A1(n37592), .A2(n15731), .ZN(n38345) );
  NOR2_X2 U31835 ( .A1(n12164), .A2(n25698), .ZN(n30055) );
  INV_X2 U31849 ( .I(n18072), .ZN(n18115) );
  XOR2_X1 U31854 ( .A1(n63730), .A2(n37588), .Z(n63271) );
  BUF_X4 U31858 ( .I(n18423), .Z(n64374) );
  BUF_X2 U31859 ( .I(n36540), .Z(n63273) );
  XOR2_X1 U31867 ( .A1(n50549), .A2(n50769), .Z(n10314) );
  OAI21_X2 U31869 ( .A1(n63634), .A2(n44643), .B(n24359), .ZN(n22395) );
  XOR2_X1 U31875 ( .A1(n63274), .A2(n9704), .Z(n13184) );
  XOR2_X1 U31883 ( .A1(n24786), .A2(n52585), .Z(n63274) );
  NOR3_X2 U31892 ( .A1(n57641), .A2(n6669), .A3(n8119), .ZN(n6667) );
  OAI22_X2 U31895 ( .A1(n47783), .A2(n63636), .B1(n49899), .B2(n13839), .ZN(
        n49903) );
  XOR2_X1 U31897 ( .A1(n17442), .A2(n24787), .Z(n17441) );
  NAND4_X2 U31898 ( .A1(n63275), .A2(n54496), .A3(n54494), .A4(n54495), .ZN(
        n54506) );
  NAND3_X2 U31899 ( .A1(n64491), .A2(n59764), .A3(n54490), .ZN(n63275) );
  NOR2_X1 U31900 ( .A1(n63281), .A2(n48799), .ZN(n48807) );
  AND2_X1 U31907 ( .A1(n14988), .A2(n14659), .Z(n64380) );
  NAND2_X2 U31909 ( .A1(n36202), .A2(n35341), .ZN(n59147) );
  NAND3_X2 U31913 ( .A1(n2419), .A2(n18507), .A3(n18505), .ZN(n36202) );
  NAND2_X2 U31915 ( .A1(n8852), .A2(n20817), .ZN(n40899) );
  NAND2_X2 U31917 ( .A1(n1500), .A2(n42355), .ZN(n8852) );
  NAND2_X2 U31926 ( .A1(n61330), .A2(n50678), .ZN(n53161) );
  BUF_X4 U31933 ( .I(n5551), .Z(n63520) );
  XOR2_X1 U31937 ( .A1(n63278), .A2(n51226), .Z(n8844) );
  XOR2_X1 U31941 ( .A1(n8846), .A2(n8847), .Z(n63278) );
  XOR2_X1 U31944 ( .A1(n52372), .A2(n64843), .Z(n59341) );
  XOR2_X1 U31945 ( .A1(n43877), .A2(n11317), .Z(n63279) );
  XOR2_X1 U31948 ( .A1(n23885), .A2(n51943), .Z(n52076) );
  NOR2_X2 U31953 ( .A1(n1450), .A2(n53345), .ZN(n53354) );
  NAND2_X2 U31958 ( .A1(n61812), .A2(n41591), .ZN(n43055) );
  NAND2_X1 U31977 ( .A1(n41592), .A2(n41593), .ZN(n63280) );
  AND2_X1 U31981 ( .A1(n48800), .A2(n48811), .Z(n63281) );
  XOR2_X1 U31982 ( .A1(n32734), .A2(n32636), .Z(n33876) );
  XOR2_X1 U31983 ( .A1(n63282), .A2(n26010), .Z(Plaintext[188]) );
  BUF_X4 U31992 ( .I(n43448), .Z(n65179) );
  NOR2_X2 U31993 ( .A1(n20124), .A2(n37361), .ZN(n37355) );
  NAND2_X2 U31997 ( .A1(n63284), .A2(n35415), .ZN(n25155) );
  NOR3_X2 U32000 ( .A1(n19188), .A2(n35420), .A3(n35419), .ZN(n63284) );
  NAND2_X2 U32001 ( .A1(n63287), .A2(n63286), .ZN(n22997) );
  NOR2_X2 U32018 ( .A1(n61788), .A2(n3553), .ZN(n63286) );
  NAND3_X1 U32021 ( .A1(n46331), .A2(n43502), .A3(n43511), .ZN(n41762) );
  NAND2_X1 U32031 ( .A1(n29787), .A2(n63355), .ZN(n27627) );
  NOR2_X2 U32036 ( .A1(n13320), .A2(n27591), .ZN(n63355) );
  OR2_X2 U32054 ( .A1(n23585), .A2(n6159), .Z(n37112) );
  XOR2_X1 U32055 ( .A1(n45055), .A2(n17159), .Z(n17158) );
  NAND3_X1 U32058 ( .A1(n56178), .A2(n56179), .A3(n63288), .ZN(n56181) );
  AND2_X1 U32062 ( .A1(n18601), .A2(n56177), .Z(n63288) );
  NAND2_X2 U32065 ( .A1(n4205), .A2(n63289), .ZN(n24215) );
  NAND2_X1 U32067 ( .A1(n4202), .A2(n4203), .ZN(n63289) );
  XOR2_X1 U32068 ( .A1(n8000), .A2(n63290), .Z(n9249) );
  XOR2_X1 U32071 ( .A1(n18098), .A2(n19564), .Z(n63290) );
  NOR2_X1 U32075 ( .A1(n9187), .A2(n2820), .ZN(n3526) );
  NOR3_X2 U32077 ( .A1(n63291), .A2(n22308), .A3(n49578), .ZN(n193) );
  XOR2_X1 U32079 ( .A1(n63292), .A2(n3275), .Z(n3272) );
  XOR2_X1 U32095 ( .A1(n3274), .A2(n60264), .Z(n63292) );
  NAND2_X1 U32096 ( .A1(n59950), .A2(n57072), .ZN(n57076) );
  NAND2_X2 U32100 ( .A1(n64338), .A2(n52857), .ZN(n57072) );
  NAND3_X1 U32106 ( .A1(n48601), .A2(n47535), .A3(n47536), .ZN(n4646) );
  NOR2_X2 U32107 ( .A1(n5771), .A2(n24801), .ZN(n48601) );
  AND2_X1 U32108 ( .A1(n18202), .A2(n18464), .Z(n57430) );
  NAND2_X2 U32111 ( .A1(n62905), .A2(n18364), .ZN(n18202) );
  XOR2_X1 U32112 ( .A1(n5105), .A2(n37631), .Z(n14553) );
  NAND2_X2 U32127 ( .A1(n8630), .A2(n13780), .ZN(n37631) );
  NAND2_X2 U32128 ( .A1(n48547), .A2(n48147), .ZN(n21399) );
  NAND2_X2 U32134 ( .A1(n48144), .A2(n48544), .ZN(n48547) );
  NOR2_X2 U32146 ( .A1(n40570), .A2(n40571), .ZN(n4137) );
  XOR2_X1 U32152 ( .A1(n32269), .A2(n32270), .Z(n11634) );
  XOR2_X1 U32157 ( .A1(n6677), .A2(n26245), .Z(n46178) );
  NAND3_X2 U32158 ( .A1(n15109), .A2(n15111), .A3(n27971), .ZN(n60237) );
  INV_X1 U32165 ( .I(n64943), .ZN(n26634) );
  NAND2_X2 U32167 ( .A1(n27565), .A2(n18751), .ZN(n64943) );
  BUF_X2 U32171 ( .I(n11818), .Z(n63293) );
  XOR2_X1 U32173 ( .A1(n22204), .A2(n63295), .Z(n18783) );
  XOR2_X1 U32175 ( .A1(n39473), .A2(n39730), .Z(n63295) );
  OAI21_X2 U32177 ( .A1(n22413), .A2(n19416), .B(n6925), .ZN(n20569) );
  NAND3_X2 U32182 ( .A1(n4439), .A2(n26235), .A3(n60095), .ZN(n25111) );
  INV_X1 U32184 ( .I(n40198), .ZN(n16842) );
  OR2_X1 U32186 ( .A1(n40198), .A2(n2124), .Z(n10374) );
  NAND2_X1 U32190 ( .A1(n64655), .A2(n25131), .ZN(n40763) );
  OAI21_X1 U32195 ( .A1(n14131), .A2(n39972), .B(n16159), .ZN(n39977) );
  NOR2_X2 U32205 ( .A1(n17530), .A2(n48122), .ZN(n64416) );
  NAND3_X1 U32209 ( .A1(n23599), .A2(n12588), .A3(n32899), .ZN(n32903) );
  NAND2_X2 U32210 ( .A1(n59798), .A2(n30195), .ZN(n30181) );
  AOI21_X1 U32211 ( .A1(n40935), .A2(n7201), .B(n63296), .ZN(n40942) );
  NAND2_X1 U32212 ( .A1(n40937), .A2(n57402), .ZN(n63296) );
  NOR2_X1 U32213 ( .A1(n63611), .A2(n61539), .ZN(n25008) );
  XOR2_X1 U32216 ( .A1(n115), .A2(n63297), .Z(n5240) );
  INV_X1 U32220 ( .I(n64945), .ZN(n63297) );
  XOR2_X1 U32222 ( .A1(n58212), .A2(n15125), .Z(n64945) );
  NOR2_X2 U32224 ( .A1(n63300), .A2(n63298), .ZN(n30196) );
  NAND2_X1 U32227 ( .A1(n26289), .A2(n63301), .ZN(n63300) );
  NAND2_X1 U32228 ( .A1(n26284), .A2(n63302), .ZN(n63301) );
  OR2_X2 U32241 ( .A1(n61646), .A2(n57701), .Z(n12768) );
  XOR2_X1 U32250 ( .A1(n22047), .A2(n38912), .Z(n39451) );
  NOR2_X2 U32253 ( .A1(n47422), .A2(n59523), .ZN(n47426) );
  NAND2_X2 U32261 ( .A1(n47683), .A2(n45267), .ZN(n47422) );
  AOI21_X1 U32263 ( .A1(n29786), .A2(n29787), .B(n58237), .ZN(n63304) );
  XOR2_X1 U32270 ( .A1(n13626), .A2(n32403), .Z(n63306) );
  XOR2_X1 U32273 ( .A1(n38794), .A2(n63307), .Z(n37002) );
  XOR2_X1 U32277 ( .A1(n6604), .A2(n15932), .Z(n63307) );
  XOR2_X1 U32280 ( .A1(n9710), .A2(n63308), .Z(n64210) );
  XOR2_X1 U32281 ( .A1(n7034), .A2(n58964), .Z(n9710) );
  XOR2_X1 U32285 ( .A1(n11734), .A2(n57250), .Z(n21027) );
  NAND2_X2 U32295 ( .A1(n33560), .A2(n32807), .ZN(n33349) );
  BUF_X2 U32299 ( .I(n48656), .Z(n63311) );
  NAND3_X2 U32300 ( .A1(n2269), .A2(n61622), .A3(n9047), .ZN(n60146) );
  NAND2_X2 U32301 ( .A1(n35247), .A2(n1221), .ZN(n33798) );
  XOR2_X1 U32305 ( .A1(n32595), .A2(n32596), .Z(n58517) );
  XOR2_X1 U32307 ( .A1(n63314), .A2(n16248), .Z(n23155) );
  XOR2_X1 U32308 ( .A1(n31200), .A2(n63316), .Z(n21488) );
  XOR2_X1 U32309 ( .A1(n19407), .A2(n16952), .Z(n63316) );
  NOR2_X2 U32319 ( .A1(n34784), .A2(n19457), .ZN(n33489) );
  XOR2_X1 U32320 ( .A1(n39586), .A2(n24859), .Z(n58467) );
  NOR3_X2 U32324 ( .A1(n61898), .A2(n63320), .A3(n27166), .ZN(n27241) );
  NOR2_X2 U32336 ( .A1(n3606), .A2(n42803), .ZN(n42975) );
  INV_X2 U32340 ( .I(n63321), .ZN(n25231) );
  XNOR2_X1 U32342 ( .A1(n57708), .A2(n61672), .ZN(n63321) );
  NAND2_X2 U32348 ( .A1(n58561), .A2(n17444), .ZN(n35873) );
  NAND2_X2 U32349 ( .A1(n35876), .A2(n37333), .ZN(n17444) );
  OR2_X1 U32350 ( .A1(n16850), .A2(n41773), .Z(n42344) );
  XOR2_X1 U32352 ( .A1(n63322), .A2(n16952), .Z(n33253) );
  XOR2_X1 U32353 ( .A1(n19407), .A2(n32654), .Z(n63322) );
  NOR2_X2 U32354 ( .A1(n36404), .A2(n21591), .ZN(n36110) );
  NOR2_X2 U32356 ( .A1(n63323), .A2(n16001), .ZN(n34469) );
  INV_X2 U32359 ( .I(n6025), .ZN(n64783) );
  NAND3_X2 U32366 ( .A1(n64304), .A2(n1804), .A3(n34307), .ZN(n6025) );
  XOR2_X1 U32372 ( .A1(n63324), .A2(n38778), .Z(n10703) );
  XOR2_X1 U32377 ( .A1(n23277), .A2(n11239), .Z(n63324) );
  XOR2_X1 U32378 ( .A1(n45844), .A2(n63325), .Z(n10447) );
  XOR2_X1 U32380 ( .A1(n23821), .A2(n63326), .Z(n58527) );
  XOR2_X1 U32385 ( .A1(n39382), .A2(n61802), .Z(n63326) );
  NAND2_X2 U32393 ( .A1(n15530), .A2(n15527), .ZN(n9254) );
  NOR2_X2 U32397 ( .A1(n58386), .A2(n15531), .ZN(n15530) );
  XOR2_X1 U32398 ( .A1(n63327), .A2(n38755), .Z(n4243) );
  XOR2_X1 U32428 ( .A1(n58252), .A2(n38943), .Z(n63327) );
  XOR2_X1 U32430 ( .A1(n63328), .A2(n32496), .Z(n30943) );
  XOR2_X1 U32431 ( .A1(n14380), .A2(n59991), .Z(n63328) );
  NAND2_X2 U32433 ( .A1(n9938), .A2(n60447), .ZN(n11160) );
  CLKBUF_X1 U32439 ( .I(n28444), .Z(n64762) );
  NAND2_X1 U32450 ( .A1(n8189), .A2(n57932), .ZN(n8188) );
  NOR3_X2 U32453 ( .A1(n63884), .A2(n52679), .A3(n52680), .ZN(n59728) );
  NAND2_X2 U32454 ( .A1(n57210), .A2(n8669), .ZN(n35979) );
  AOI21_X2 U32464 ( .A1(n41200), .A2(n22329), .B(n63332), .ZN(n60493) );
  INV_X2 U32465 ( .I(n40734), .ZN(n63332) );
  XOR2_X1 U32467 ( .A1(n25968), .A2(n20883), .Z(n11192) );
  NOR2_X2 U32469 ( .A1(n12941), .A2(n15578), .ZN(n22435) );
  NOR2_X2 U32477 ( .A1(n64459), .A2(n3345), .ZN(n3344) );
  OAI22_X2 U32479 ( .A1(n64657), .A2(n52696), .B1(n1283), .B2(n1602), .ZN(
        n52697) );
  XOR2_X1 U32480 ( .A1(n30977), .A2(n63335), .Z(n30979) );
  XOR2_X1 U32485 ( .A1(n30976), .A2(n30975), .Z(n63335) );
  NAND3_X2 U32486 ( .A1(n24150), .A2(n35164), .A3(n35167), .ZN(n39644) );
  NAND3_X2 U32491 ( .A1(n63336), .A2(n18201), .A3(n993), .ZN(n63649) );
  NAND2_X1 U32499 ( .A1(n11800), .A2(n12759), .ZN(n63336) );
  NOR2_X2 U32502 ( .A1(n63337), .A2(n32541), .ZN(n6723) );
  INV_X2 U32504 ( .I(n37114), .ZN(n36755) );
  BUF_X2 U32506 ( .I(n59020), .Z(n63339) );
  XOR2_X1 U32518 ( .A1(n63340), .A2(n3033), .Z(n17216) );
  XOR2_X1 U32528 ( .A1(n59568), .A2(n46319), .Z(n63340) );
  NAND2_X2 U32531 ( .A1(n9716), .A2(n41898), .ZN(n40802) );
  INV_X2 U32533 ( .I(n3249), .ZN(n58548) );
  NAND2_X2 U32534 ( .A1(n47482), .A2(n24128), .ZN(n3249) );
  NOR2_X2 U32539 ( .A1(n47108), .A2(n47107), .ZN(n24966) );
  NAND4_X2 U32544 ( .A1(n47086), .A2(n3288), .A3(n3287), .A4(n47082), .ZN(
        n47107) );
  XOR2_X1 U32546 ( .A1(n32346), .A2(n59933), .Z(n1313) );
  NAND3_X2 U32547 ( .A1(n14303), .A2(n14302), .A3(n14301), .ZN(n32346) );
  OAI21_X2 U32555 ( .A1(n12050), .A2(n1780), .B(n63638), .ZN(n37083) );
  AND2_X1 U32559 ( .A1(n42273), .A2(n3946), .Z(n57415) );
  XOR2_X1 U32563 ( .A1(n18782), .A2(n496), .Z(n18781) );
  INV_X1 U32566 ( .I(n55944), .ZN(n63432) );
  BUF_X2 U32568 ( .I(n33481), .Z(n63344) );
  AOI22_X2 U32573 ( .A1(n37280), .A2(n11178), .B1(n37278), .B2(n37279), .ZN(
        n37283) );
  NAND2_X2 U32576 ( .A1(n8476), .A2(n16696), .ZN(n28091) );
  XOR2_X1 U32581 ( .A1(n63744), .A2(n51763), .Z(n10618) );
  XOR2_X1 U32582 ( .A1(n50660), .A2(n51097), .Z(n25949) );
  NAND3_X2 U32588 ( .A1(n3594), .A2(n3593), .A3(n3595), .ZN(n22678) );
  XOR2_X1 U32592 ( .A1(n6400), .A2(n63345), .Z(n6404) );
  XOR2_X1 U32597 ( .A1(n6403), .A2(n12533), .Z(n63345) );
  XOR2_X1 U32598 ( .A1(n57507), .A2(n63346), .Z(n63902) );
  XOR2_X1 U32599 ( .A1(n38191), .A2(n37727), .Z(n63346) );
  AOI22_X1 U32603 ( .A1(n4254), .A2(n53381), .B1(n53380), .B2(n63347), .ZN(
        n53390) );
  OAI22_X1 U32605 ( .A1(n53601), .A2(n11041), .B1(n2018), .B2(n53602), .ZN(
        n63347) );
  AOI21_X1 U32606 ( .A1(n12158), .A2(n23112), .B(n41384), .ZN(n41388) );
  NAND2_X2 U32607 ( .A1(n63350), .A2(n61800), .ZN(n63349) );
  NAND2_X2 U32608 ( .A1(n41015), .A2(n60928), .ZN(n63350) );
  NAND2_X2 U32609 ( .A1(n25383), .A2(n24444), .ZN(n50230) );
  OR2_X1 U32616 ( .A1(n61961), .A2(n64347), .Z(n47602) );
  XOR2_X1 U32617 ( .A1(n51041), .A2(n63351), .Z(n7753) );
  XOR2_X1 U32620 ( .A1(n17336), .A2(n63352), .Z(n63351) );
  INV_X2 U32625 ( .I(n51034), .ZN(n63352) );
  INV_X2 U32634 ( .I(n36540), .ZN(n33017) );
  NAND2_X2 U32638 ( .A1(n35687), .A2(n32748), .ZN(n36540) );
  XOR2_X1 U32644 ( .A1(n8526), .A2(n32294), .Z(n11455) );
  XOR2_X1 U32645 ( .A1(n16821), .A2(n63353), .Z(n32294) );
  INV_X2 U32649 ( .I(n22070), .ZN(n63353) );
  NOR3_X2 U32662 ( .A1(n61948), .A2(n15642), .A3(n63354), .ZN(n15619) );
  NAND2_X2 U32663 ( .A1(n33119), .A2(n4266), .ZN(n63354) );
  XOR2_X1 U32683 ( .A1(n44269), .A2(n17919), .Z(n64266) );
  NAND2_X2 U32692 ( .A1(n10862), .A2(n53528), .ZN(n53511) );
  NOR2_X2 U32697 ( .A1(n17225), .A2(n53492), .ZN(n53528) );
  XOR2_X1 U32701 ( .A1(n33048), .A2(n24103), .Z(n13934) );
  XOR2_X1 U32703 ( .A1(n14049), .A2(n18204), .Z(n28983) );
  NOR2_X2 U32705 ( .A1(n8460), .A2(n12896), .ZN(n18204) );
  OAI22_X1 U32715 ( .A1(n27105), .A2(n28381), .B1(n28384), .B2(n15477), .ZN(
        n27108) );
  NAND2_X2 U32717 ( .A1(n28376), .A2(n13704), .ZN(n15477) );
  INV_X2 U32721 ( .I(n28959), .ZN(n25269) );
  NAND2_X2 U32727 ( .A1(n57102), .A2(n57101), .ZN(n63356) );
  NAND4_X1 U32730 ( .A1(n15872), .A2(n56145), .A3(n17961), .A4(n56185), .ZN(
        n22990) );
  NOR2_X2 U32740 ( .A1(n56146), .A2(n56167), .ZN(n56145) );
  NAND2_X1 U32749 ( .A1(n23209), .A2(n27135), .ZN(n28329) );
  OAI21_X1 U32750 ( .A1(n63358), .A2(n19243), .B(n22263), .ZN(n48333) );
  NOR2_X2 U32754 ( .A1(n2024), .A2(n58232), .ZN(n45498) );
  AOI21_X2 U32755 ( .A1(n63362), .A2(n10179), .B(n29738), .ZN(n11430) );
  XOR2_X1 U32756 ( .A1(n46605), .A2(n5029), .Z(n58127) );
  NAND2_X2 U32767 ( .A1(n42907), .A2(n42908), .ZN(n46605) );
  NAND3_X2 U32791 ( .A1(n47400), .A2(n47863), .A3(n47401), .ZN(n63363) );
  NAND2_X2 U32796 ( .A1(n63364), .A2(n4584), .ZN(n58297) );
  NOR3_X2 U32810 ( .A1(n16053), .A2(n57856), .A3(n46074), .ZN(n63364) );
  XOR2_X1 U32815 ( .A1(n63365), .A2(n15644), .Z(n38794) );
  XOR2_X1 U32820 ( .A1(n22949), .A2(n38382), .Z(n63365) );
  XOR2_X1 U32822 ( .A1(n63366), .A2(n45343), .Z(n21303) );
  XOR2_X1 U32825 ( .A1(n45342), .A2(n61564), .Z(n63366) );
  INV_X2 U32832 ( .I(n63367), .ZN(n6988) );
  NOR2_X2 U32833 ( .A1(n63370), .A2(n40746), .ZN(n24174) );
  NAND3_X2 U32834 ( .A1(n40742), .A2(n40741), .A3(n61103), .ZN(n63370) );
  NOR2_X1 U32841 ( .A1(n37022), .A2(n37096), .ZN(n7600) );
  NAND2_X2 U32842 ( .A1(n16750), .A2(n29586), .ZN(n29076) );
  NAND2_X2 U32846 ( .A1(n22755), .A2(n53163), .ZN(n53130) );
  NAND2_X2 U32858 ( .A1(n50484), .A2(n50485), .ZN(n53163) );
  XOR2_X1 U32859 ( .A1(n12293), .A2(n12294), .Z(n38323) );
  NOR3_X2 U32860 ( .A1(n63373), .A2(n47257), .A3(n47264), .ZN(n21684) );
  NAND4_X2 U32863 ( .A1(n5641), .A2(n12500), .A3(n3047), .A4(n35371), .ZN(
        n22048) );
  NOR2_X1 U32864 ( .A1(n65108), .A2(n63374), .ZN(n4284) );
  NAND3_X1 U32865 ( .A1(n2584), .A2(n4078), .A3(n9296), .ZN(n63374) );
  XOR2_X1 U32866 ( .A1(n18941), .A2(n63755), .Z(n38529) );
  XOR2_X1 U32875 ( .A1(n10899), .A2(n59166), .Z(n64055) );
  XOR2_X1 U32880 ( .A1(n3381), .A2(n13705), .Z(n10899) );
  NOR2_X1 U32882 ( .A1(n18116), .A2(n47192), .ZN(n63994) );
  XOR2_X1 U32891 ( .A1(n63377), .A2(n46654), .Z(n60309) );
  NOR3_X2 U32892 ( .A1(n4431), .A2(n39879), .A3(n42011), .ZN(n63378) );
  NOR3_X2 U32895 ( .A1(n48513), .A2(n48254), .A3(n48642), .ZN(n48635) );
  NAND3_X2 U32896 ( .A1(n25766), .A2(n63566), .A3(n54547), .ZN(n25765) );
  OAI21_X2 U32901 ( .A1(n43446), .A2(n43449), .B(n42369), .ZN(n63380) );
  NAND2_X2 U32904 ( .A1(n28398), .A2(n28399), .ZN(n64594) );
  NAND2_X2 U32914 ( .A1(n27087), .A2(n3317), .ZN(n28399) );
  XOR2_X1 U32915 ( .A1(n39757), .A2(n13555), .Z(n60107) );
  XOR2_X1 U32920 ( .A1(n3838), .A2(n37686), .Z(n39757) );
  NAND2_X2 U32922 ( .A1(n59609), .A2(n55625), .ZN(n55654) );
  XOR2_X1 U32924 ( .A1(n14378), .A2(n32356), .Z(n63383) );
  NAND2_X1 U32929 ( .A1(n4312), .A2(n53309), .ZN(n13512) );
  XOR2_X1 U32933 ( .A1(n63384), .A2(n53319), .Z(Plaintext[18]) );
  NOR4_X2 U32939 ( .A1(n53317), .A2(n61469), .A3(n15404), .A4(n16827), .ZN(
        n63384) );
  NAND2_X1 U32942 ( .A1(n28687), .A2(n63589), .ZN(n2417) );
  AOI22_X1 U32950 ( .A1(n63385), .A2(n61916), .B1(n5814), .B2(n5815), .ZN(
        n5813) );
  NAND3_X2 U32951 ( .A1(n10041), .A2(n40557), .A3(n60693), .ZN(n3725) );
  NOR2_X2 U32954 ( .A1(n18333), .A2(n61659), .ZN(n40557) );
  NAND2_X1 U32961 ( .A1(n63470), .A2(n12446), .ZN(n60609) );
  XOR2_X1 U32963 ( .A1(n1189), .A2(n15047), .Z(n64877) );
  NAND2_X2 U32964 ( .A1(n60966), .A2(n5078), .ZN(n15047) );
  XOR2_X1 U32965 ( .A1(n65279), .A2(n52416), .Z(n6255) );
  XOR2_X1 U32981 ( .A1(n51230), .A2(n50743), .Z(n51390) );
  XOR2_X1 U32982 ( .A1(n10344), .A2(n57408), .Z(n51230) );
  XOR2_X1 U32985 ( .A1(n5487), .A2(n6299), .Z(n657) );
  XOR2_X1 U33002 ( .A1(n63390), .A2(n16372), .Z(n16369) );
  XOR2_X1 U33012 ( .A1(n16370), .A2(n39396), .Z(n63390) );
  XOR2_X1 U33017 ( .A1(n6988), .A2(n15047), .Z(n1945) );
  NAND3_X2 U33026 ( .A1(n18325), .A2(n60782), .A3(n61904), .ZN(n63391) );
  NAND2_X2 U33027 ( .A1(n49211), .A2(n17523), .ZN(n44009) );
  NOR2_X2 U33033 ( .A1(n8604), .A2(n359), .ZN(n49211) );
  NOR2_X2 U33039 ( .A1(n13162), .A2(n63393), .ZN(n58734) );
  NAND2_X2 U33040 ( .A1(n42913), .A2(n42912), .ZN(n63393) );
  OAI21_X1 U33042 ( .A1(n21589), .A2(n22726), .B(n27396), .ZN(n18767) );
  NAND2_X2 U33044 ( .A1(n34350), .A2(n32922), .ZN(n63581) );
  BUF_X2 U33053 ( .I(n16491), .Z(n63394) );
  NOR2_X1 U33055 ( .A1(n57676), .A2(n65235), .ZN(n58668) );
  NAND2_X2 U33056 ( .A1(n37268), .A2(n57860), .ZN(n63838) );
  NAND3_X2 U33067 ( .A1(n29932), .A2(n8521), .A3(n162), .ZN(n30802) );
  AOI22_X2 U33071 ( .A1(n41085), .A2(n41086), .B1(n41087), .B2(n64896), .ZN(
        n41088) );
  NAND2_X2 U33073 ( .A1(n61739), .A2(n9663), .ZN(n43318) );
  NAND2_X1 U33080 ( .A1(n63402), .A2(n57716), .ZN(n36844) );
  INV_X2 U33082 ( .I(n49450), .ZN(n49848) );
  OAI22_X1 U33085 ( .A1(n34294), .A2(n34387), .B1(n34293), .B2(n35280), .ZN(
        n11181) );
  XOR2_X1 U33097 ( .A1(n33145), .A2(n14025), .Z(n59923) );
  NOR2_X1 U33099 ( .A1(n1934), .A2(n1941), .ZN(n63397) );
  INV_X4 U33100 ( .I(n59119), .ZN(n15157) );
  NOR2_X2 U33107 ( .A1(n25166), .A2(n8225), .ZN(n59119) );
  NAND2_X2 U33111 ( .A1(n2944), .A2(n45957), .ZN(n3716) );
  XOR2_X1 U33115 ( .A1(n7557), .A2(n5155), .Z(n64419) );
  XOR2_X1 U33118 ( .A1(n6332), .A2(n10295), .Z(n59665) );
  XOR2_X1 U33126 ( .A1(n63400), .A2(n55833), .Z(Plaintext[131]) );
  NAND3_X1 U33128 ( .A1(n12433), .A2(n12430), .A3(n12431), .ZN(n63400) );
  NAND3_X2 U33137 ( .A1(n6655), .A2(n391), .A3(n63401), .ZN(n49012) );
  NOR2_X1 U33141 ( .A1(n63403), .A2(n46809), .ZN(n46812) );
  INV_X2 U33145 ( .I(n47799), .ZN(n63404) );
  NOR2_X2 U33149 ( .A1(n63405), .A2(n16357), .ZN(n58914) );
  XOR2_X1 U33152 ( .A1(n13430), .A2(n7744), .Z(n52094) );
  XOR2_X1 U33161 ( .A1(n63407), .A2(n51506), .Z(n17800) );
  XOR2_X1 U33165 ( .A1(n18091), .A2(n9868), .Z(n63407) );
  NAND2_X2 U33168 ( .A1(n54876), .A2(n54873), .ZN(n54902) );
  AOI22_X2 U33169 ( .A1(n54788), .A2(n54787), .B1(n54789), .B2(n55402), .ZN(
        n54873) );
  NAND3_X2 U33171 ( .A1(n35226), .A2(n35707), .A3(n35228), .ZN(n64464) );
  AOI21_X2 U33172 ( .A1(n64465), .A2(n62598), .B(n64464), .ZN(n59582) );
  XOR2_X1 U33174 ( .A1(n51030), .A2(n23852), .Z(n10416) );
  NAND2_X2 U33178 ( .A1(n2071), .A2(n2076), .ZN(n23852) );
  NAND2_X2 U33183 ( .A1(n9493), .A2(n9495), .ZN(n24257) );
  XOR2_X1 U33186 ( .A1(n52499), .A2(n52498), .Z(n10105) );
  OR2_X1 U33188 ( .A1(n28266), .A2(n63751), .Z(n63750) );
  OR2_X1 U33192 ( .A1(n21073), .A2(n63372), .Z(n4250) );
  NOR2_X2 U33193 ( .A1(n42784), .A2(n41660), .ZN(n42782) );
  XOR2_X1 U33196 ( .A1(n5954), .A2(n61590), .Z(n5953) );
  INV_X2 U33198 ( .I(n63410), .ZN(n19160) );
  INV_X4 U33202 ( .I(n8669), .ZN(n23766) );
  NAND2_X2 U33205 ( .A1(n6919), .A2(n60167), .ZN(n8669) );
  XOR2_X1 U33207 ( .A1(n14055), .A2(n63411), .Z(n6037) );
  XOR2_X1 U33214 ( .A1(n44319), .A2(n23987), .Z(n63411) );
  XOR2_X1 U33215 ( .A1(n12685), .A2(n63413), .Z(n12682) );
  XOR2_X1 U33219 ( .A1(n31673), .A2(n12686), .Z(n63413) );
  NOR2_X1 U33220 ( .A1(n63415), .A2(n63414), .ZN(n64225) );
  INV_X1 U33221 ( .I(n49378), .ZN(n63414) );
  NAND3_X1 U33227 ( .A1(n49380), .A2(n18769), .A3(n49379), .ZN(n63415) );
  OAI22_X1 U33235 ( .A1(n49581), .A2(n20311), .B1(n49572), .B2(n1637), .ZN(
        n48945) );
  NOR3_X1 U33236 ( .A1(n18559), .A2(n63416), .A3(n18558), .ZN(n58394) );
  AOI21_X1 U33237 ( .A1(n18557), .A2(n55897), .B(n60203), .ZN(n63416) );
  AOI21_X1 U33240 ( .A1(n56580), .A2(n56591), .B(n56579), .ZN(n56584) );
  NOR2_X2 U33241 ( .A1(n328), .A2(n6000), .ZN(n5997) );
  NAND2_X2 U33244 ( .A1(n37246), .A2(n37253), .ZN(n16652) );
  NOR2_X2 U33247 ( .A1(n22413), .A2(n12768), .ZN(n5264) );
  NAND3_X2 U33248 ( .A1(n63418), .A2(n14573), .A3(n14571), .ZN(n14570) );
  AOI22_X2 U33249 ( .A1(n63419), .A2(n1740), .B1(n20394), .B2(n39139), .ZN(
        n20393) );
  NAND2_X2 U33251 ( .A1(n20395), .A2(n39137), .ZN(n63419) );
  BUF_X2 U33255 ( .I(n551), .Z(n63421) );
  INV_X1 U33258 ( .I(n57973), .ZN(n63422) );
  XOR2_X1 U33260 ( .A1(n63424), .A2(n51335), .Z(n2256) );
  NOR2_X2 U33264 ( .A1(n9051), .A2(n49715), .ZN(n51335) );
  NAND2_X1 U33267 ( .A1(n57078), .A2(n63425), .ZN(n57084) );
  NAND2_X1 U33268 ( .A1(n57076), .A2(n25435), .ZN(n63425) );
  NAND2_X1 U33269 ( .A1(n46767), .A2(n57398), .ZN(n64881) );
  XOR2_X1 U33283 ( .A1(n38909), .A2(n63426), .Z(n930) );
  XOR2_X1 U33287 ( .A1(n64945), .A2(n64678), .Z(n64297) );
  XOR2_X1 U33294 ( .A1(n10406), .A2(n63427), .Z(n63749) );
  XOR2_X1 U33300 ( .A1(n17801), .A2(n19029), .Z(n63427) );
  NAND3_X2 U33301 ( .A1(n18097), .A2(n60387), .A3(n18095), .ZN(n56812) );
  XOR2_X1 U33309 ( .A1(n32046), .A2(n25025), .Z(n63428) );
  XOR2_X1 U33321 ( .A1(n63429), .A2(n61109), .Z(n2469) );
  AOI22_X1 U33326 ( .A1(n34322), .A2(n17148), .B1(n35306), .B2(n34323), .ZN(
        n34327) );
  XOR2_X1 U33329 ( .A1(n5350), .A2(n5352), .Z(n64260) );
  NOR3_X2 U33330 ( .A1(n63935), .A2(n63433), .A3(n63432), .ZN(n55947) );
  OAI21_X1 U33337 ( .A1(n30468), .A2(n34992), .B(n34982), .ZN(n30472) );
  NAND2_X1 U33343 ( .A1(n57081), .A2(n63781), .ZN(n59954) );
  NAND3_X2 U33350 ( .A1(n59964), .A2(n8578), .A3(n59965), .ZN(n61137) );
  NAND2_X1 U33362 ( .A1(n3561), .A2(n63406), .ZN(n9494) );
  XOR2_X1 U33363 ( .A1(n31773), .A2(n32370), .Z(n58384) );
  AOI22_X2 U33367 ( .A1(n897), .A2(n65225), .B1(n34295), .B2(n13735), .ZN(
        n13404) );
  XOR2_X1 U33374 ( .A1(n13364), .A2(n24953), .Z(n5942) );
  XOR2_X1 U33376 ( .A1(n14960), .A2(n61634), .Z(n63436) );
  NAND2_X2 U33378 ( .A1(n15715), .A2(n1364), .ZN(n26536) );
  NAND2_X2 U33383 ( .A1(n11699), .A2(n11097), .ZN(n19270) );
  NOR2_X2 U33384 ( .A1(n14419), .A2(n47180), .ZN(n47167) );
  NAND3_X2 U33388 ( .A1(n14725), .A2(n31062), .A3(n14724), .ZN(n31985) );
  NAND2_X2 U33389 ( .A1(n38551), .A2(n63430), .ZN(n36778) );
  NAND2_X1 U33391 ( .A1(n8775), .A2(n27965), .ZN(n25302) );
  AOI21_X2 U33392 ( .A1(n58210), .A2(n42842), .B(n42118), .ZN(n63437) );
  INV_X2 U33395 ( .I(n3086), .ZN(n63438) );
  INV_X4 U33397 ( .I(n25096), .ZN(n29566) );
  NAND2_X2 U33398 ( .A1(n14220), .A2(n14221), .ZN(n25096) );
  NOR2_X2 U33401 ( .A1(n52285), .A2(n61724), .ZN(n59722) );
  NOR2_X2 U33402 ( .A1(n52692), .A2(n56239), .ZN(n52285) );
  NOR3_X2 U33403 ( .A1(n11452), .A2(n46757), .A3(n46756), .ZN(n12900) );
  OR2_X2 U33414 ( .A1(n62530), .A2(n43561), .Z(n43566) );
  NAND2_X2 U33417 ( .A1(n1583), .A2(n1257), .ZN(n56967) );
  XOR2_X1 U33421 ( .A1(n11265), .A2(n32470), .Z(n60888) );
  XOR2_X1 U33428 ( .A1(n16821), .A2(n31004), .Z(n13742) );
  XOR2_X1 U33429 ( .A1(n29941), .A2(n17758), .Z(n31004) );
  AND2_X1 U33431 ( .A1(n42393), .A2(n41689), .Z(n42087) );
  NAND2_X2 U33435 ( .A1(n1392), .A2(n19241), .ZN(n42393) );
  NAND2_X1 U33464 ( .A1(n41092), .A2(n41896), .ZN(n41093) );
  NAND3_X2 U33467 ( .A1(n17316), .A2(n18001), .A3(n63439), .ZN(n49226) );
  NAND2_X2 U33468 ( .A1(n16745), .A2(n9346), .ZN(n49272) );
  OR2_X2 U33475 ( .A1(n14662), .A2(n39781), .Z(n41079) );
  XOR2_X1 U33480 ( .A1(n8280), .A2(n63832), .Z(n58392) );
  OAI21_X1 U33481 ( .A1(n40858), .A2(n40857), .B(n40856), .ZN(n64503) );
  INV_X1 U33484 ( .I(n64503), .ZN(n64502) );
  INV_X1 U33488 ( .I(n18214), .ZN(n63440) );
  AOI21_X2 U33496 ( .A1(n9538), .A2(n9539), .B(n63441), .ZN(n9536) );
  NAND2_X1 U33513 ( .A1(n9540), .A2(n9541), .ZN(n63441) );
  NAND4_X2 U33515 ( .A1(n42323), .A2(n42322), .A3(n42321), .A4(n42320), .ZN(
        n63442) );
  OR3_X1 U33517 ( .A1(n18827), .A2(n21960), .A3(n39058), .Z(n38598) );
  NAND2_X2 U33519 ( .A1(n2187), .A2(n63618), .ZN(n2192) );
  NOR2_X1 U33525 ( .A1(n6950), .A2(n6953), .ZN(n7421) );
  BUF_X2 U33533 ( .I(n34989), .Z(n63444) );
  AND2_X1 U33539 ( .A1(n1718), .A2(n42914), .Z(n42911) );
  NOR2_X2 U33543 ( .A1(n63445), .A2(n45745), .ZN(n25870) );
  AOI21_X2 U33544 ( .A1(n22319), .A2(n25691), .B(n4380), .ZN(n63445) );
  NAND2_X1 U33549 ( .A1(n23116), .A2(n53161), .ZN(n9187) );
  NAND3_X2 U33559 ( .A1(n58158), .A2(n12133), .A3(n12134), .ZN(n23116) );
  NOR2_X2 U33562 ( .A1(n49286), .A2(n44788), .ZN(n48768) );
  NAND2_X2 U33563 ( .A1(n16412), .A2(n16418), .ZN(n49277) );
  NAND2_X1 U33564 ( .A1(n3526), .A2(n9533), .ZN(n4645) );
  NAND2_X2 U33572 ( .A1(n41898), .A2(n23145), .ZN(n64659) );
  OR2_X1 U33576 ( .A1(n14872), .A2(n60875), .Z(n34188) );
  INV_X2 U33580 ( .I(n63451), .ZN(n57165) );
  NOR2_X2 U33587 ( .A1(n5147), .A2(n61749), .ZN(n63451) );
  NOR2_X2 U33588 ( .A1(n10000), .A2(n9839), .ZN(n23346) );
  NAND2_X2 U33602 ( .A1(n5203), .A2(n63452), .ZN(n46367) );
  XOR2_X1 U33613 ( .A1(n57408), .A2(n50761), .Z(n12681) );
  BUF_X2 U33614 ( .I(n30953), .Z(n63454) );
  NOR2_X1 U33616 ( .A1(n31245), .A2(n31241), .ZN(n31243) );
  NAND2_X1 U33617 ( .A1(n14090), .A2(n63458), .ZN(n63457) );
  AND2_X1 U33618 ( .A1(n53703), .A2(n53704), .Z(n63458) );
  NAND3_X2 U33619 ( .A1(n36803), .A2(n36312), .A3(n3864), .ZN(n2857) );
  XOR2_X1 U33620 ( .A1(n38741), .A2(n38325), .Z(n39735) );
  NAND2_X2 U33623 ( .A1(n25751), .A2(n34104), .ZN(n38741) );
  NOR2_X1 U33624 ( .A1(n16808), .A2(n23589), .ZN(n25722) );
  NAND2_X1 U33628 ( .A1(n59479), .A2(n63527), .ZN(n59013) );
  XOR2_X1 U33633 ( .A1(n10536), .A2(n64443), .Z(n46383) );
  AND2_X2 U33634 ( .A1(n25999), .A2(n13068), .Z(n33445) );
  XOR2_X1 U33636 ( .A1(n24035), .A2(n39749), .Z(n39786) );
  NAND2_X2 U33637 ( .A1(n9381), .A2(n9382), .ZN(n24953) );
  XOR2_X1 U33639 ( .A1(n46579), .A2(n11879), .Z(n11878) );
  XOR2_X1 U33640 ( .A1(n19226), .A2(n45247), .Z(n46579) );
  NAND2_X2 U33642 ( .A1(n42786), .A2(n42785), .ZN(n43028) );
  NAND2_X2 U33643 ( .A1(n56129), .A2(n63550), .ZN(n64408) );
  NOR2_X2 U33644 ( .A1(n61222), .A2(n51116), .ZN(n56129) );
  NOR2_X1 U33648 ( .A1(n60419), .A2(n63459), .ZN(n64090) );
  NAND4_X1 U33649 ( .A1(n56649), .A2(n56648), .A3(n56646), .A4(n56647), .ZN(
        n63459) );
  AOI22_X2 U33651 ( .A1(n16176), .A2(n63460), .B1(n44874), .B2(n61845), .ZN(
        n14235) );
  INV_X1 U33653 ( .I(n63461), .ZN(n63460) );
  NAND2_X1 U33656 ( .A1(n46900), .A2(n44871), .ZN(n63461) );
  NOR2_X1 U33657 ( .A1(n31789), .A2(n58557), .ZN(n31791) );
  OAI21_X2 U33662 ( .A1(n13593), .A2(n30543), .B(n57526), .ZN(n63462) );
  NOR2_X2 U33666 ( .A1(n63463), .A2(n3666), .ZN(n8660) );
  INV_X2 U33676 ( .I(n3667), .ZN(n63464) );
  NAND2_X2 U33677 ( .A1(n1405), .A2(n58367), .ZN(n41459) );
  XOR2_X1 U33685 ( .A1(n11828), .A2(n11829), .Z(n58147) );
  NAND2_X2 U33688 ( .A1(n36017), .A2(n36016), .ZN(n11829) );
  NAND3_X1 U33689 ( .A1(n5775), .A2(n40656), .A3(n709), .ZN(n40657) );
  INV_X1 U33696 ( .I(n43153), .ZN(n63466) );
  OR2_X2 U33699 ( .A1(n30810), .A2(n25449), .Z(n30804) );
  NAND3_X2 U33700 ( .A1(n61720), .A2(n45267), .A3(n46835), .ZN(n46840) );
  NAND3_X1 U33701 ( .A1(n42019), .A2(n62346), .A3(n43699), .ZN(n63470) );
  INV_X1 U33711 ( .I(n8403), .ZN(n63541) );
  OAI21_X1 U33712 ( .A1(n63468), .A2(n19775), .B(n50292), .ZN(n23614) );
  NAND2_X1 U33715 ( .A1(n18608), .A2(n48717), .ZN(n63468) );
  BUF_X2 U33719 ( .I(n37046), .Z(n63469) );
  AND2_X1 U33722 ( .A1(n17030), .A2(n34836), .Z(n37280) );
  OAI21_X1 U33727 ( .A1(n41689), .A2(n42404), .B(n42407), .ZN(n19807) );
  INV_X2 U33729 ( .I(n58402), .ZN(n41689) );
  NOR2_X2 U33731 ( .A1(n25068), .A2(n13306), .ZN(n58402) );
  INV_X2 U33732 ( .I(n14361), .ZN(n32071) );
  NAND2_X2 U33734 ( .A1(n34238), .A2(n34708), .ZN(n14361) );
  INV_X1 U33735 ( .I(n63471), .ZN(n3433) );
  NAND3_X2 U33743 ( .A1(n29155), .A2(n8528), .A3(n22482), .ZN(n63471) );
  NAND2_X2 U33744 ( .A1(n4926), .A2(n11299), .ZN(n11828) );
  NAND2_X1 U33747 ( .A1(n19853), .A2(n61873), .ZN(n56198) );
  OR2_X2 U33750 ( .A1(n3705), .A2(n41289), .Z(n41294) );
  NAND2_X2 U33772 ( .A1(n29793), .A2(n30078), .ZN(n7736) );
  XOR2_X1 U33777 ( .A1(n36324), .A2(n38847), .Z(n20435) );
  XOR2_X1 U33778 ( .A1(n17845), .A2(n38105), .Z(n36324) );
  NAND2_X2 U33779 ( .A1(n13868), .A2(n13869), .ZN(n15698) );
  XOR2_X1 U33781 ( .A1(n65143), .A2(n4311), .Z(n50680) );
  NAND3_X2 U33788 ( .A1(n63474), .A2(n64792), .A3(n10466), .ZN(n4386) );
  NAND3_X1 U33789 ( .A1(n42560), .A2(n42102), .A3(n42101), .ZN(n63474) );
  OR2_X2 U33790 ( .A1(n29875), .A2(n10079), .Z(n36605) );
  XOR2_X1 U33796 ( .A1(n63475), .A2(n21509), .Z(n18873) );
  XOR2_X1 U33797 ( .A1(n24829), .A2(n18964), .Z(n63475) );
  NAND3_X2 U33798 ( .A1(n63476), .A2(n40814), .A3(n40813), .ZN(n58004) );
  NAND2_X2 U33799 ( .A1(n978), .A2(n42288), .ZN(n42273) );
  NOR2_X1 U33804 ( .A1(n36071), .A2(n36074), .ZN(n63477) );
  AOI21_X2 U33819 ( .A1(n20243), .A2(n41496), .B(n63480), .ZN(n2148) );
  NAND2_X2 U33820 ( .A1(n14214), .A2(n43698), .ZN(n63480) );
  XOR2_X1 U33825 ( .A1(n64837), .A2(n41659), .Z(n58446) );
  NOR2_X2 U33827 ( .A1(n58269), .A2(n2433), .ZN(n49849) );
  NOR3_X2 U33831 ( .A1(n61901), .A2(n15154), .A3(n45612), .ZN(n57471) );
  NAND2_X2 U33832 ( .A1(n25687), .A2(n40911), .ZN(n44238) );
  INV_X2 U33841 ( .I(n40954), .ZN(n63483) );
  NOR2_X2 U33844 ( .A1(n39103), .A2(n40952), .ZN(n40954) );
  BUF_X2 U33848 ( .I(n1787), .Z(n63484) );
  NAND2_X1 U33849 ( .A1(n54976), .A2(n63486), .ZN(n9106) );
  BUF_X2 U33851 ( .I(n59018), .Z(n63487) );
  XOR2_X1 U33856 ( .A1(n24040), .A2(n59854), .Z(n51044) );
  OAI21_X2 U33860 ( .A1(n17865), .A2(n34195), .B(n33710), .ZN(n63488) );
  XOR2_X1 U33871 ( .A1(n51086), .A2(n50942), .Z(n12254) );
  NAND2_X2 U33873 ( .A1(n19242), .A2(n48695), .ZN(n51086) );
  NOR3_X2 U33876 ( .A1(n63489), .A2(n36032), .A3(n36034), .ZN(n36035) );
  NAND2_X2 U33882 ( .A1(n36029), .A2(n36028), .ZN(n63489) );
  NAND2_X1 U33884 ( .A1(n10127), .A2(n63490), .ZN(n36253) );
  OAI21_X1 U33891 ( .A1(n36249), .A2(n61223), .B(n36248), .ZN(n63490) );
  NAND3_X2 U33894 ( .A1(n4232), .A2(n54537), .A3(n54565), .ZN(n54547) );
  NAND2_X1 U33896 ( .A1(n36742), .A2(n36746), .ZN(n36741) );
  NAND2_X2 U33898 ( .A1(n35834), .A2(n33807), .ZN(n8957) );
  XOR2_X1 U33913 ( .A1(n33253), .A2(n63491), .Z(n15381) );
  INV_X1 U33927 ( .I(n31872), .ZN(n63491) );
  OR3_X2 U33949 ( .A1(n63492), .A2(n28638), .A3(n28636), .Z(n7283) );
  OAI22_X1 U33950 ( .A1(n28629), .A2(n28628), .B1(n28626), .B2(n28627), .ZN(
        n63492) );
  NAND2_X2 U33965 ( .A1(n14620), .A2(n11818), .ZN(n42160) );
  AND2_X1 U33986 ( .A1(n19165), .A2(n64015), .Z(n61358) );
  OR2_X1 U33999 ( .A1(n30334), .A2(n11092), .Z(n63497) );
  XOR2_X1 U34009 ( .A1(n33203), .A2(n31425), .Z(n30735) );
  NAND3_X2 U34019 ( .A1(n29852), .A2(n29851), .A3(n29853), .ZN(n33203) );
  XOR2_X1 U34020 ( .A1(n18355), .A2(n39476), .Z(n22204) );
  XOR2_X1 U34021 ( .A1(n13732), .A2(n10898), .Z(n39476) );
  XOR2_X1 U34028 ( .A1(n63498), .A2(n44480), .Z(n44115) );
  XOR2_X1 U34035 ( .A1(n5011), .A2(n44114), .Z(n63498) );
  NAND2_X2 U34040 ( .A1(n27822), .A2(n23825), .ZN(n4848) );
  NAND3_X1 U34058 ( .A1(n63503), .A2(n27836), .A3(n63502), .ZN(n27845) );
  AND2_X1 U34059 ( .A1(n27834), .A2(n27833), .Z(n63502) );
  OAI21_X1 U34063 ( .A1(n27832), .A2(n60541), .B(n27831), .ZN(n63503) );
  XOR2_X1 U34068 ( .A1(n9374), .A2(n30921), .Z(n24292) );
  INV_X2 U34080 ( .I(n63505), .ZN(n63586) );
  NAND3_X1 U34086 ( .A1(n22246), .A2(n59699), .A3(n45676), .ZN(n63508) );
  NOR2_X1 U34088 ( .A1(n63508), .A2(n25002), .ZN(n25001) );
  NAND4_X2 U34090 ( .A1(n17506), .A2(n17505), .A3(n30765), .A4(n30764), .ZN(
        n63507) );
  BUF_X2 U34092 ( .I(n24977), .Z(n63510) );
  NOR2_X2 U34095 ( .A1(n8509), .A2(n8195), .ZN(n37409) );
  NAND2_X2 U34099 ( .A1(n8223), .A2(n4512), .ZN(n8509) );
  XOR2_X1 U34102 ( .A1(n8979), .A2(n2778), .Z(n10300) );
  XOR2_X1 U34111 ( .A1(n1929), .A2(n13359), .Z(n8979) );
  XOR2_X1 U34112 ( .A1(n38630), .A2(n8541), .Z(n24976) );
  NOR3_X2 U34113 ( .A1(n63746), .A2(n20823), .A3(n20822), .ZN(n55423) );
  OR2_X1 U34114 ( .A1(n63621), .A2(n18608), .Z(n58415) );
  NAND2_X2 U34116 ( .A1(n59925), .A2(n63511), .ZN(n1200) );
  AND2_X2 U34124 ( .A1(n55444), .A2(n24165), .Z(n18145) );
  AOI21_X2 U34125 ( .A1(n61912), .A2(n17631), .B(n61215), .ZN(n63513) );
  XOR2_X1 U34127 ( .A1(n39618), .A2(n38711), .Z(n8353) );
  NAND2_X2 U34129 ( .A1(n36103), .A2(n36102), .ZN(n39618) );
  XOR2_X1 U34132 ( .A1(n60570), .A2(n9736), .Z(n63514) );
  NAND2_X2 U34140 ( .A1(n37388), .A2(n16891), .ZN(n6177) );
  NOR2_X2 U34141 ( .A1(n4972), .A2(n11668), .ZN(n37388) );
  NAND2_X1 U34142 ( .A1(n26978), .A2(n28884), .ZN(n63798) );
  AOI21_X2 U34143 ( .A1(n64214), .A2(n9479), .B(n63515), .ZN(n9477) );
  NAND3_X2 U34144 ( .A1(n42061), .A2(n42059), .A3(n42060), .ZN(n63515) );
  NAND2_X1 U34147 ( .A1(n63516), .A2(n55025), .ZN(n14100) );
  NAND2_X2 U34157 ( .A1(n63517), .A2(n63562), .ZN(n54259) );
  OAI22_X2 U34167 ( .A1(n17051), .A2(n51839), .B1(n61694), .B2(n61371), .ZN(
        n63517) );
  NOR2_X2 U34169 ( .A1(n54721), .A2(n57201), .ZN(n54738) );
  NAND2_X2 U34170 ( .A1(n54767), .A2(n26015), .ZN(n54721) );
  AOI21_X2 U34178 ( .A1(n9925), .A2(n9924), .B(n1634), .ZN(n63518) );
  XOR2_X1 U34189 ( .A1(n59341), .A2(n63519), .Z(n61354) );
  XOR2_X1 U34195 ( .A1(n6994), .A2(n11768), .Z(n63519) );
  NOR2_X1 U34201 ( .A1(n60052), .A2(n43836), .ZN(n43076) );
  XOR2_X1 U34202 ( .A1(n63521), .A2(n52630), .Z(n52632) );
  XOR2_X1 U34204 ( .A1(n58989), .A2(n8076), .Z(n63521) );
  NOR3_X2 U34211 ( .A1(n12275), .A2(n12276), .A3(n63522), .ZN(n12273) );
  OAI22_X2 U34221 ( .A1(n27608), .A2(n27607), .B1(n21281), .B2(n9251), .ZN(
        n63522) );
  NOR2_X2 U34223 ( .A1(n40832), .A2(n39950), .ZN(n65110) );
  NAND2_X2 U34234 ( .A1(n41132), .A2(n1407), .ZN(n39950) );
  NAND2_X2 U34240 ( .A1(n23835), .A2(n9548), .ZN(n4998) );
  NOR2_X2 U34243 ( .A1(n64377), .A2(n11855), .ZN(n40703) );
  INV_X2 U34254 ( .I(n56555), .ZN(n52692) );
  NOR2_X2 U34255 ( .A1(n56829), .A2(n12468), .ZN(n56555) );
  NAND2_X2 U34261 ( .A1(n1871), .A2(n19225), .ZN(n29787) );
  NAND2_X2 U34269 ( .A1(n15423), .A2(n15422), .ZN(n1871) );
  XOR2_X1 U34272 ( .A1(n11462), .A2(n57311), .Z(n11460) );
  NAND3_X2 U34284 ( .A1(n46477), .A2(n63523), .A3(n46476), .ZN(n57685) );
  NOR2_X2 U34294 ( .A1(n64372), .A2(n20595), .ZN(n10486) );
  XOR2_X1 U34295 ( .A1(n63524), .A2(n52195), .Z(n52204) );
  XOR2_X1 U34297 ( .A1(n52193), .A2(n19125), .Z(n63524) );
  NAND2_X1 U34299 ( .A1(n29702), .A2(n14212), .ZN(n29708) );
  NOR2_X1 U34300 ( .A1(n29704), .A2(n28620), .ZN(n29702) );
  XOR2_X1 U34307 ( .A1(n19349), .A2(n17171), .Z(n17739) );
  OR2_X1 U34311 ( .A1(n4233), .A2(n46866), .Z(n46037) );
  OAI21_X1 U34313 ( .A1(n19690), .A2(n22595), .B(n19689), .ZN(n63527) );
  XOR2_X1 U34318 ( .A1(n63528), .A2(n7309), .Z(n9989) );
  XOR2_X1 U34328 ( .A1(n2954), .A2(n20789), .Z(n63528) );
  BUF_X2 U34333 ( .I(n3302), .Z(n63529) );
  NAND2_X2 U34335 ( .A1(n1817), .A2(n4560), .ZN(n6206) );
  NAND2_X1 U34343 ( .A1(n3198), .A2(n27879), .ZN(n3197) );
  INV_X2 U34348 ( .I(n63530), .ZN(n30121) );
  NOR2_X2 U34349 ( .A1(n1351), .A2(n29766), .ZN(n63530) );
  BUF_X2 U34353 ( .I(n23508), .Z(n63533) );
  NOR2_X1 U34354 ( .A1(n63534), .A2(n10368), .ZN(n10377) );
  NAND2_X1 U34358 ( .A1(n10375), .A2(n11444), .ZN(n63534) );
  XOR2_X1 U34361 ( .A1(n4370), .A2(n38289), .Z(n64273) );
  XOR2_X1 U34368 ( .A1(n52013), .A2(n51690), .Z(n7246) );
  NAND3_X2 U34373 ( .A1(n15127), .A2(n19782), .A3(n15128), .ZN(n51690) );
  XOR2_X1 U34375 ( .A1(n52436), .A2(n8066), .Z(n5334) );
  XOR2_X1 U34384 ( .A1(n15413), .A2(n8073), .Z(n8074) );
  NOR2_X2 U34386 ( .A1(n64369), .A2(n8093), .ZN(n15413) );
  NAND2_X2 U34387 ( .A1(n42127), .A2(n11883), .ZN(n42129) );
  NAND2_X2 U34395 ( .A1(n46736), .A2(n47434), .ZN(n47752) );
  NOR3_X2 U34396 ( .A1(n63536), .A2(n24424), .A3(n53237), .ZN(n24422) );
  XOR2_X1 U34399 ( .A1(n37967), .A2(n39186), .Z(n5457) );
  NAND2_X2 U34402 ( .A1(n14908), .A2(n14909), .ZN(n37967) );
  XOR2_X1 U34413 ( .A1(n45401), .A2(n44029), .Z(n10746) );
  NAND2_X2 U34414 ( .A1(n58879), .A2(n63539), .ZN(n24425) );
  OR2_X1 U34417 ( .A1(n49884), .A2(n1377), .Z(n63542) );
  XOR2_X1 U34440 ( .A1(n13261), .A2(n14782), .Z(n2963) );
  XOR2_X1 U34445 ( .A1(n25961), .A2(n46691), .Z(n14782) );
  XOR2_X1 U34455 ( .A1(n38191), .A2(n38190), .Z(n38193) );
  XOR2_X1 U34463 ( .A1(n6045), .A2(n1337), .Z(n38191) );
  OAI22_X2 U34467 ( .A1(n6523), .A2(n47583), .B1(n47586), .B2(n47584), .ZN(
        n47589) );
  NOR2_X2 U34473 ( .A1(n63543), .A2(n15548), .ZN(n41232) );
  NAND2_X2 U34478 ( .A1(n11472), .A2(n41400), .ZN(n63543) );
  NOR2_X1 U34499 ( .A1(n57971), .A2(n57972), .ZN(n10815) );
  XOR2_X1 U34505 ( .A1(n63544), .A2(n38959), .Z(n15591) );
  XOR2_X1 U34506 ( .A1(n19249), .A2(n38955), .Z(n63544) );
  XOR2_X1 U34513 ( .A1(n31637), .A2(n63545), .Z(n3522) );
  XOR2_X1 U34516 ( .A1(n31640), .A2(n25652), .Z(n63545) );
  XOR2_X1 U34531 ( .A1(n2741), .A2(n15500), .Z(n14160) );
  BUF_X2 U34544 ( .I(n14314), .Z(n63546) );
  NOR2_X2 U34545 ( .A1(n37424), .A2(n36909), .ZN(n37436) );
  XOR2_X1 U34549 ( .A1(n3523), .A2(n63353), .Z(n31816) );
  INV_X2 U34550 ( .I(n63547), .ZN(n47100) );
  NOR2_X2 U34557 ( .A1(n26032), .A2(n18100), .ZN(n63547) );
  BUF_X2 U34566 ( .I(n38771), .Z(n63548) );
  BUF_X2 U34573 ( .I(n9806), .Z(n63549) );
  XOR2_X1 U34575 ( .A1(n63672), .A2(n57975), .Z(n16558) );
  INV_X1 U34579 ( .I(n34191), .ZN(n63553) );
  NOR3_X2 U34580 ( .A1(n24552), .A2(n63551), .A3(n56443), .ZN(n56522) );
  NOR2_X1 U34588 ( .A1(n3762), .A2(n57339), .ZN(n59479) );
  XOR2_X1 U34594 ( .A1(n7398), .A2(n16983), .Z(n58823) );
  XOR2_X1 U34600 ( .A1(n58822), .A2(n11802), .Z(n7398) );
  OAI21_X1 U34604 ( .A1(n34224), .A2(n34385), .B(n63552), .ZN(n34226) );
  AOI21_X1 U34606 ( .A1(n8631), .A2(n34222), .B(n35802), .ZN(n63552) );
  NOR3_X2 U34611 ( .A1(n15716), .A2(n55893), .A3(n55854), .ZN(n55880) );
  AND2_X1 U34622 ( .A1(n65115), .A2(n8912), .Z(n42684) );
  XOR2_X1 U34629 ( .A1(n63869), .A2(n64319), .Z(n9575) );
  NAND2_X2 U34633 ( .A1(n10064), .A2(n63586), .ZN(n34588) );
  OAI21_X1 U34637 ( .A1(n18134), .A2(n55394), .B(n60421), .ZN(n55396) );
  NAND2_X2 U34639 ( .A1(n17470), .A2(n63554), .ZN(n42822) );
  AND2_X1 U34640 ( .A1(n41208), .A2(n17468), .Z(n63554) );
  OR2_X1 U34642 ( .A1(n54488), .A2(n54487), .Z(n64715) );
  NOR2_X2 U34648 ( .A1(n36075), .A2(n36139), .ZN(n36313) );
  OAI21_X1 U34649 ( .A1(n16103), .A2(n42824), .B(n42823), .ZN(n42830) );
  NAND3_X2 U34661 ( .A1(n11003), .A2(n11001), .A3(n11004), .ZN(n18734) );
  OR2_X1 U34662 ( .A1(n19142), .A2(n1386), .Z(n46798) );
  XOR2_X1 U34668 ( .A1(n63667), .A2(n44507), .Z(n45063) );
  NOR2_X2 U34672 ( .A1(n7828), .A2(n7826), .ZN(n44507) );
  OR3_X1 U34673 ( .A1(n50141), .A2(n62035), .A3(n9646), .Z(n50298) );
  XOR2_X1 U34681 ( .A1(n46353), .A2(n5630), .Z(n44184) );
  NOR2_X2 U34682 ( .A1(n42841), .A2(n42840), .ZN(n46353) );
  NOR2_X2 U34683 ( .A1(n63556), .A2(n13650), .ZN(n21400) );
  NOR2_X2 U34693 ( .A1(n13630), .A2(n43736), .ZN(n42844) );
  NAND3_X2 U34695 ( .A1(n59558), .A2(n16065), .A3(n31219), .ZN(n25455) );
  NAND4_X2 U34697 ( .A1(n40798), .A2(n40789), .A3(n40790), .A4(n40799), .ZN(
        n63556) );
  NAND2_X2 U34698 ( .A1(n63658), .A2(n61664), .ZN(n8767) );
  XOR2_X1 U34702 ( .A1(n3437), .A2(n63558), .Z(n3436) );
  XOR2_X1 U34705 ( .A1(n37901), .A2(n25248), .Z(n63558) );
  NAND2_X2 U34706 ( .A1(n27737), .A2(n27736), .ZN(n4211) );
  NAND2_X2 U34710 ( .A1(n63578), .A2(n63579), .ZN(n34656) );
  NAND2_X2 U34714 ( .A1(n13170), .A2(n26064), .ZN(n39186) );
  XOR2_X1 U34717 ( .A1(n8623), .A2(n8622), .Z(n63559) );
  XOR2_X1 U34718 ( .A1(n63560), .A2(n10320), .Z(n21319) );
  XOR2_X1 U34725 ( .A1(n13324), .A2(n63768), .Z(n63560) );
  NAND2_X1 U34734 ( .A1(n21272), .A2(n1592), .ZN(n55598) );
  XOR2_X1 U34738 ( .A1(n63563), .A2(n32475), .Z(n31414) );
  XOR2_X1 U34742 ( .A1(n17668), .A2(n22227), .Z(n63563) );
  BUF_X4 U34750 ( .I(n40394), .Z(n64459) );
  XOR2_X1 U34751 ( .A1(n46121), .A2(n46122), .Z(n23906) );
  NAND3_X2 U34752 ( .A1(n41707), .A2(n24648), .A3(n25373), .ZN(n46121) );
  XOR2_X1 U34758 ( .A1(n7265), .A2(n24223), .Z(n63564) );
  NAND2_X2 U34765 ( .A1(n14194), .A2(n63565), .ZN(n25677) );
  NAND2_X2 U34773 ( .A1(n54486), .A2(n64715), .ZN(n54507) );
  NAND2_X2 U34779 ( .A1(n19870), .A2(n58349), .ZN(n8287) );
  NOR2_X2 U34784 ( .A1(n98), .A2(n99), .ZN(n911) );
  XOR2_X1 U34792 ( .A1(n24803), .A2(n52325), .Z(n24929) );
  NAND2_X2 U34804 ( .A1(n47650), .A2(n47651), .ZN(n52325) );
  NAND3_X2 U34813 ( .A1(n54558), .A2(n54574), .A3(n54581), .ZN(n63566) );
  NAND2_X2 U34825 ( .A1(n17590), .A2(n29905), .ZN(n30862) );
  OAI22_X2 U34829 ( .A1(n12201), .A2(n47817), .B1(n47820), .B2(n3510), .ZN(
        n64557) );
  INV_X1 U34833 ( .I(n63567), .ZN(n60815) );
  AOI21_X1 U34837 ( .A1(n54630), .A2(n54807), .B(n63568), .ZN(n63567) );
  XOR2_X1 U34851 ( .A1(n44907), .A2(n24019), .Z(n63570) );
  NAND2_X1 U34859 ( .A1(n23617), .A2(n48081), .ZN(n10978) );
  NOR2_X2 U34867 ( .A1(n15823), .A2(n45889), .ZN(n48081) );
  NAND3_X2 U34881 ( .A1(n63573), .A2(n40784), .A3(n40783), .ZN(n46432) );
  AND2_X1 U34884 ( .A1(n40782), .A2(n43199), .Z(n63573) );
  XOR2_X1 U34886 ( .A1(n46543), .A2(n45842), .Z(n10985) );
  NAND2_X1 U34891 ( .A1(n3613), .A2(n56311), .ZN(n56324) );
  XOR2_X1 U34911 ( .A1(n63574), .A2(n65079), .Z(Plaintext[130]) );
  NAND4_X2 U34914 ( .A1(n55808), .A2(n55809), .A3(n55807), .A4(n55806), .ZN(
        n63574) );
  NAND2_X1 U34918 ( .A1(n55665), .A2(n56265), .ZN(n55667) );
  AOI21_X1 U34923 ( .A1(n10486), .A2(n25549), .B(n56905), .ZN(n12765) );
  XOR2_X1 U34926 ( .A1(n46213), .A2(n17059), .Z(n20824) );
  NAND3_X2 U34937 ( .A1(n23107), .A2(n24493), .A3(n24491), .ZN(n46213) );
  NOR2_X1 U34940 ( .A1(n20165), .A2(n4817), .ZN(n63575) );
  NAND3_X1 U34941 ( .A1(n57097), .A2(n57098), .A3(n57115), .ZN(n59920) );
  NAND3_X2 U34951 ( .A1(n17507), .A2(n15108), .A3(n63577), .ZN(n18547) );
  NOR2_X2 U34957 ( .A1(n14526), .A2(n14525), .ZN(n63577) );
  INV_X2 U34958 ( .I(n11643), .ZN(n63578) );
  XOR2_X1 U34962 ( .A1(n1488), .A2(n7698), .Z(n639) );
  XOR2_X1 U34963 ( .A1(n19189), .A2(n24621), .Z(n61524) );
  INV_X2 U34966 ( .I(n33122), .ZN(n63583) );
  NOR2_X2 U34967 ( .A1(n6028), .A2(n60756), .ZN(n3394) );
  NAND2_X2 U34969 ( .A1(n25261), .A2(n36566), .ZN(n4035) );
  NAND2_X2 U34985 ( .A1(n9344), .A2(n24878), .ZN(n27603) );
  XOR2_X1 U34987 ( .A1(n6596), .A2(n63587), .Z(n26148) );
  XOR2_X1 U34989 ( .A1(n51917), .A2(n64507), .Z(n63587) );
  AND2_X1 U34998 ( .A1(n10358), .A2(n22333), .Z(n34596) );
  NAND3_X1 U35007 ( .A1(n21117), .A2(n21114), .A3(n63588), .ZN(n63993) );
  AOI22_X1 U35009 ( .A1(n21124), .A2(n9715), .B1(n24), .B2(n21122), .ZN(n63588) );
  NOR2_X2 U35015 ( .A1(n34078), .A2(n20812), .ZN(n17595) );
  NAND2_X2 U35017 ( .A1(n34032), .A2(n64860), .ZN(n34078) );
  AOI21_X1 U35018 ( .A1(n40752), .A2(n40750), .B(n10611), .ZN(n63590) );
  XOR2_X1 U35021 ( .A1(n5660), .A2(n39658), .Z(n61295) );
  OR2_X1 U35044 ( .A1(n30410), .A2(n30331), .Z(n63592) );
  INV_X2 U35050 ( .I(n40402), .ZN(n41422) );
  NAND2_X2 U35061 ( .A1(n1743), .A2(n38932), .ZN(n40402) );
  XOR2_X1 U35066 ( .A1(n17232), .A2(n32230), .Z(n31966) );
  BUF_X2 U35080 ( .I(n10485), .Z(n63593) );
  XOR2_X1 U35087 ( .A1(n25483), .A2(n63596), .Z(n4514) );
  XOR2_X1 U35093 ( .A1(n63976), .A2(n50905), .Z(n63596) );
  AOI22_X2 U35095 ( .A1(n14118), .A2(n64379), .B1(n42198), .B2(n42197), .ZN(
        n8655) );
  NAND2_X2 U35105 ( .A1(n58148), .A2(n36089), .ZN(n38711) );
  NAND2_X2 U35106 ( .A1(n47304), .A2(n26180), .ZN(n47302) );
  NAND2_X1 U35115 ( .A1(n15514), .A2(n61000), .ZN(n40155) );
  INV_X1 U35116 ( .I(n63597), .ZN(n64581) );
  OAI21_X1 U35123 ( .A1(n39988), .A2(n40759), .B(n41478), .ZN(n63597) );
  NAND3_X2 U35124 ( .A1(n5537), .A2(n57252), .A3(n58017), .ZN(n23067) );
  XOR2_X1 U35130 ( .A1(n11829), .A2(n36994), .Z(n39188) );
  INV_X2 U35142 ( .I(n27442), .ZN(n28798) );
  NAND2_X2 U35145 ( .A1(n27441), .A2(n23800), .ZN(n27442) );
  AND2_X1 U35153 ( .A1(n28803), .A2(n6775), .Z(n26997) );
  AOI21_X2 U35160 ( .A1(n63598), .A2(n11612), .B(n64797), .ZN(n25445) );
  AOI22_X1 U35162 ( .A1(n35999), .A2(n36000), .B1(n57391), .B2(n36608), .ZN(
        n36006) );
  XOR2_X1 U35177 ( .A1(n12596), .A2(n63599), .Z(n5440) );
  XOR2_X1 U35179 ( .A1(n39249), .A2(n36995), .Z(n63599) );
  INV_X1 U35181 ( .I(n48252), .ZN(n48631) );
  NAND2_X2 U35186 ( .A1(n23347), .A2(n25340), .ZN(n45436) );
  AND2_X1 U35189 ( .A1(n42135), .A2(n42136), .Z(n63600) );
  XOR2_X1 U35194 ( .A1(n1684), .A2(n59382), .Z(n60114) );
  NAND2_X2 U35198 ( .A1(n24760), .A2(n42789), .ZN(n59382) );
  XOR2_X1 U35200 ( .A1(n63601), .A2(n12029), .Z(n60176) );
  XOR2_X1 U35208 ( .A1(n9037), .A2(n59625), .Z(n63601) );
  AOI22_X2 U35210 ( .A1(n23925), .A2(n45802), .B1(n22426), .B2(n46758), .ZN(
        n63602) );
  NAND3_X2 U35220 ( .A1(n48788), .A2(n48786), .A3(n48787), .ZN(n52207) );
  XOR2_X1 U35225 ( .A1(n63604), .A2(n18923), .Z(n19010) );
  XOR2_X1 U35234 ( .A1(n38635), .A2(n37509), .Z(n63604) );
  INV_X2 U35243 ( .I(n63606), .ZN(n24274) );
  XNOR2_X1 U35272 ( .A1(n21238), .A2(n21239), .ZN(n63606) );
  NOR3_X2 U35277 ( .A1(n64071), .A2(n22622), .A3(n32801), .ZN(n25366) );
  AOI21_X2 U35302 ( .A1(n29982), .A2(n30549), .B(n29976), .ZN(n63607) );
  NAND2_X1 U35328 ( .A1(n42663), .A2(n42664), .ZN(n43250) );
  NOR4_X2 U35330 ( .A1(n11158), .A2(n15193), .A3(n11159), .A4(n60958), .ZN(
        n24594) );
  AND2_X2 U35339 ( .A1(n26110), .A2(n38134), .Z(n41868) );
  NOR2_X2 U35342 ( .A1(n60476), .A2(n60690), .ZN(n64956) );
  XOR2_X1 U35352 ( .A1(n38300), .A2(n20288), .Z(n37777) );
  NOR2_X2 U35365 ( .A1(n24362), .A2(n10958), .ZN(n18844) );
  NAND2_X2 U35367 ( .A1(n58604), .A2(n47403), .ZN(n23247) );
  XOR2_X1 U35368 ( .A1(n64574), .A2(n5834), .Z(n5833) );
  INV_X2 U35371 ( .I(n63608), .ZN(n22882) );
  XNOR2_X1 U35377 ( .A1(n58479), .A2(n58480), .ZN(n63608) );
  OR2_X1 U35379 ( .A1(n21218), .A2(n20524), .Z(n63609) );
  NAND2_X2 U35398 ( .A1(n55156), .A2(n55164), .ZN(n2784) );
  NAND3_X2 U35401 ( .A1(n11689), .A2(n8212), .A3(n48104), .ZN(n110) );
  INV_X1 U35416 ( .I(n20402), .ZN(n37494) );
  NAND3_X2 U35430 ( .A1(n20382), .A2(n61890), .A3(n5073), .ZN(n20402) );
  NAND2_X2 U35432 ( .A1(n59453), .A2(n61847), .ZN(n57719) );
  NAND2_X1 U35434 ( .A1(n50350), .A2(n50349), .ZN(n21351) );
  XOR2_X1 U35435 ( .A1(n4479), .A2(n17024), .Z(n32133) );
  NAND2_X2 U35437 ( .A1(n24904), .A2(n3567), .ZN(n55674) );
  AOI22_X1 U35439 ( .A1(n2793), .A2(n34930), .B1(n2791), .B2(n34924), .ZN(
        n63611) );
  NOR3_X2 U35442 ( .A1(n60812), .A2(n20969), .A3(n20968), .ZN(n23284) );
  NAND2_X2 U35444 ( .A1(n25507), .A2(n25913), .ZN(n43561) );
  XOR2_X1 U35448 ( .A1(n21535), .A2(n63612), .Z(n59944) );
  XOR2_X1 U35449 ( .A1(n45031), .A2(n63613), .Z(n63612) );
  XOR2_X1 U35461 ( .A1(n1749), .A2(n63614), .Z(n2701) );
  XOR2_X1 U35480 ( .A1(n20367), .A2(n35076), .Z(n63614) );
  NAND3_X2 U35482 ( .A1(n21191), .A2(n21194), .A3(n21193), .ZN(n36080) );
  XOR2_X1 U35494 ( .A1(n63615), .A2(n58338), .Z(n5830) );
  XOR2_X1 U35495 ( .A1(n32294), .A2(n64600), .Z(n63615) );
  INV_X2 U35500 ( .I(n35447), .ZN(n63616) );
  OR2_X1 U35504 ( .A1(n35443), .A2(n63616), .Z(n12570) );
  NAND2_X1 U35505 ( .A1(n14054), .A2(n36965), .ZN(n36963) );
  NAND2_X2 U35506 ( .A1(n52890), .A2(n56993), .ZN(n20634) );
  BUF_X2 U35507 ( .I(n1428), .Z(n63617) );
  NAND4_X2 U35514 ( .A1(n13578), .A2(n20777), .A3(n809), .A4(n58236), .ZN(
        n15155) );
  NAND3_X2 U35517 ( .A1(n40520), .A2(n9314), .A3(n63620), .ZN(n21375) );
  NAND3_X2 U35518 ( .A1(n6112), .A2(n6111), .A3(n6110), .ZN(n23587) );
  XOR2_X1 U35520 ( .A1(n63622), .A2(n31988), .Z(n63991) );
  XOR2_X1 U35523 ( .A1(n6481), .A2(n6483), .Z(n63622) );
  INV_X2 U35533 ( .I(n63623), .ZN(n57239) );
  NAND2_X2 U35538 ( .A1(n56559), .A2(n56829), .ZN(n63623) );
  BUF_X2 U35541 ( .I(n33345), .Z(n63624) );
  XOR2_X1 U35543 ( .A1(n5312), .A2(n15982), .Z(n16582) );
  NOR2_X2 U35553 ( .A1(n29608), .A2(n29619), .ZN(n64145) );
  NAND3_X1 U35554 ( .A1(n40583), .A2(n41898), .A3(n40804), .ZN(n37775) );
  NAND3_X1 U35557 ( .A1(n59271), .A2(n41898), .A3(n42263), .ZN(n63626) );
  XOR2_X1 U35558 ( .A1(n8109), .A2(n23461), .Z(n32292) );
  NOR2_X2 U35565 ( .A1(n7705), .A2(n36224), .ZN(n36456) );
  INV_X1 U35578 ( .I(n3999), .ZN(n63628) );
  OAI21_X2 U35583 ( .A1(n63629), .A2(n28240), .B(n28237), .ZN(n11140) );
  NOR2_X2 U35590 ( .A1(n28069), .A2(n23586), .ZN(n63629) );
  NOR3_X2 U35593 ( .A1(n63630), .A2(n36806), .A3(n36805), .ZN(n36815) );
  AOI21_X2 U35597 ( .A1(n62246), .A2(n36803), .B(n36801), .ZN(n63630) );
  XOR2_X1 U35606 ( .A1(n16458), .A2(n839), .Z(n21503) );
  NOR2_X2 U35610 ( .A1(n59790), .A2(n64976), .ZN(n16458) );
  NAND2_X2 U35626 ( .A1(n1345), .A2(n1545), .ZN(n34957) );
  INV_X2 U35634 ( .I(n3947), .ZN(n22185) );
  XOR2_X1 U35635 ( .A1(n11632), .A2(n63631), .Z(n3947) );
  XOR2_X1 U35642 ( .A1(n63632), .A2(n9637), .Z(n15216) );
  XOR2_X1 U35647 ( .A1(n43665), .A2(n63633), .Z(n63632) );
  NAND2_X1 U35651 ( .A1(n56225), .A2(n63635), .ZN(n55981) );
  INV_X2 U35665 ( .I(n56436), .ZN(n63635) );
  OAI21_X2 U35671 ( .A1(n25812), .A2(n63186), .B(n49908), .ZN(n63636) );
  OAI21_X2 U35674 ( .A1(n63665), .A2(n61887), .B(n37319), .ZN(n6910) );
  INV_X2 U35677 ( .I(n13195), .ZN(n34415) );
  BUF_X2 U35679 ( .I(n13666), .Z(n63638) );
  XOR2_X1 U35685 ( .A1(n63639), .A2(n56915), .Z(Plaintext[182]) );
  NAND3_X1 U35687 ( .A1(n56914), .A2(n56913), .A3(n10233), .ZN(n63639) );
  NAND2_X2 U35689 ( .A1(n2483), .A2(n22892), .ZN(n35996) );
  NOR2_X2 U35695 ( .A1(n15171), .A2(n35508), .ZN(n35950) );
  INV_X4 U35698 ( .I(n24609), .ZN(n35508) );
  NOR2_X2 U35701 ( .A1(n25194), .A2(n22339), .ZN(n24609) );
  NAND2_X2 U35703 ( .A1(n64835), .A2(n63640), .ZN(n21240) );
  NAND3_X1 U35721 ( .A1(n6119), .A2(n6118), .A3(n48392), .ZN(n63641) );
  INV_X1 U35727 ( .I(n10893), .ZN(n11675) );
  XOR2_X1 U35728 ( .A1(n10893), .A2(n63642), .Z(n11647) );
  XOR2_X1 U35732 ( .A1(n46269), .A2(n7365), .Z(n10893) );
  BUF_X2 U35733 ( .I(n1781), .Z(n63643) );
  NAND3_X2 U35739 ( .A1(n17969), .A2(n17968), .A3(n18373), .ZN(n52013) );
  NAND2_X2 U35741 ( .A1(n61574), .A2(n5807), .ZN(n37008) );
  XOR2_X1 U35747 ( .A1(n38591), .A2(n39386), .Z(n21289) );
  NAND3_X2 U35750 ( .A1(n32155), .A2(n32156), .A3(n32157), .ZN(n39386) );
  NOR2_X1 U35766 ( .A1(n55387), .A2(n55389), .ZN(n15310) );
  XOR2_X1 U35770 ( .A1(n39314), .A2(n39315), .Z(n39659) );
  NAND3_X2 U35771 ( .A1(n64754), .A2(n57551), .A3(n63648), .ZN(n56616) );
  NAND3_X2 U35774 ( .A1(n12424), .A2(n64014), .A3(n9599), .ZN(n22396) );
  OAI21_X1 U35777 ( .A1(n40570), .A2(n39836), .B(n59225), .ZN(n4952) );
  NOR2_X1 U35798 ( .A1(n53130), .A2(n53129), .ZN(n2038) );
  NOR2_X2 U35799 ( .A1(n12761), .A2(n63649), .ZN(n20347) );
  NAND3_X1 U35811 ( .A1(n22592), .A2(n57901), .A3(n55463), .ZN(n64841) );
  INV_X2 U35817 ( .I(n63650), .ZN(n65274) );
  XOR2_X1 U35818 ( .A1(n44442), .A2(n3656), .Z(n63650) );
  XOR2_X1 U35819 ( .A1(n59206), .A2(n2666), .Z(n58608) );
  XOR2_X1 U35822 ( .A1(n50863), .A2(n58989), .Z(n51997) );
  XOR2_X1 U35838 ( .A1(n50929), .A2(n54289), .Z(n50863) );
  NOR2_X1 U35843 ( .A1(n17264), .A2(n53181), .ZN(n17263) );
  INV_X1 U35849 ( .I(n53541), .ZN(n17264) );
  NOR2_X2 U35853 ( .A1(n53396), .A2(n62090), .ZN(n53541) );
  AOI21_X2 U35860 ( .A1(n48077), .A2(n48080), .B(n48078), .ZN(n63652) );
  NOR3_X2 U35871 ( .A1(n63654), .A2(n18028), .A3(n63653), .ZN(n18027) );
  NAND2_X2 U35875 ( .A1(n41640), .A2(n40864), .ZN(n63653) );
  NOR3_X2 U35885 ( .A1(n63656), .A2(n63655), .A3(n9323), .ZN(n14676) );
  XOR2_X1 U35900 ( .A1(n63657), .A2(n53764), .Z(Plaintext[40]) );
  NOR3_X1 U35901 ( .A1(n25000), .A2(n24999), .A3(n43215), .ZN(n63658) );
  XOR2_X1 U35920 ( .A1(n63659), .A2(n19202), .Z(n50452) );
  XOR2_X1 U35923 ( .A1(n63660), .A2(n45862), .Z(n57622) );
  XOR2_X1 U35931 ( .A1(n11554), .A2(n42421), .Z(n63660) );
  XOR2_X1 U35932 ( .A1(n2070), .A2(n25150), .Z(n14538) );
  NOR2_X1 U35937 ( .A1(n14127), .A2(n49614), .ZN(n64547) );
  NAND2_X1 U35946 ( .A1(n61814), .A2(n64547), .ZN(n59198) );
  NAND2_X1 U35947 ( .A1(n1628), .A2(n6227), .ZN(n4376) );
  NAND2_X2 U35948 ( .A1(n15632), .A2(n52126), .ZN(n55914) );
  XOR2_X1 U35950 ( .A1(n63662), .A2(n43686), .Z(n64402) );
  XOR2_X1 U35967 ( .A1(n2960), .A2(n60568), .Z(n63662) );
  INV_X1 U35972 ( .I(n49714), .ZN(n48424) );
  NAND2_X2 U35974 ( .A1(n63663), .A2(n48421), .ZN(n49714) );
  XOR2_X1 U35980 ( .A1(n25568), .A2(n24650), .Z(n13156) );
  XOR2_X1 U35984 ( .A1(n22846), .A2(n51956), .Z(n25568) );
  AND2_X1 U35989 ( .A1(n18138), .A2(n47730), .Z(n47745) );
  XOR2_X1 U35999 ( .A1(n37966), .A2(n11665), .Z(n21763) );
  INV_X1 U36000 ( .I(n26046), .ZN(n11665) );
  XOR2_X1 U36001 ( .A1(n18862), .A2(n6832), .Z(n26046) );
  BUF_X2 U36012 ( .I(n18464), .Z(n63664) );
  NOR3_X2 U36013 ( .A1(n4530), .A2(n40913), .A3(n1012), .ZN(n14444) );
  NAND2_X1 U36019 ( .A1(n52254), .A2(n52659), .ZN(n64119) );
  NOR2_X2 U36030 ( .A1(n29824), .A2(n16961), .ZN(n30324) );
  MUX2_X1 U36040 ( .I0(n41663), .I1(n41662), .S(n57283), .Z(n41669) );
  NAND2_X2 U36049 ( .A1(n9608), .A2(n1342), .ZN(n24153) );
  NAND2_X1 U36050 ( .A1(n63668), .A2(n34155), .ZN(n32898) );
  BUF_X2 U36052 ( .I(n15148), .Z(n63671) );
  NAND3_X1 U36072 ( .A1(n42662), .A2(n42127), .A3(n10004), .ZN(n21325) );
  NOR2_X2 U36077 ( .A1(n21549), .A2(n41626), .ZN(n57756) );
  XOR2_X1 U36079 ( .A1(n8196), .A2(n65027), .Z(n7381) );
  XOR2_X1 U36080 ( .A1(n11570), .A2(n13532), .Z(n63672) );
  NAND2_X2 U36082 ( .A1(n63673), .A2(n12135), .ZN(n44735) );
  NOR3_X2 U36084 ( .A1(n58091), .A2(n64411), .A3(n12140), .ZN(n63673) );
  XOR2_X1 U36103 ( .A1(n14910), .A2(n44586), .Z(n61360) );
  XOR2_X1 U36105 ( .A1(n18922), .A2(n9484), .Z(n7872) );
  XOR2_X1 U36114 ( .A1(n4681), .A2(n60717), .Z(n18922) );
  XOR2_X1 U36118 ( .A1(n31597), .A2(n32505), .Z(n17764) );
  NAND2_X2 U36119 ( .A1(n9562), .A2(n27397), .ZN(n65111) );
  OAI21_X1 U36122 ( .A1(n20904), .A2(n63674), .B(n19428), .ZN(n59001) );
  OR2_X1 U36123 ( .A1(n57116), .A2(n63784), .Z(n57088) );
  NAND3_X2 U36129 ( .A1(n63676), .A2(n63675), .A3(n12567), .ZN(n10945) );
  NAND2_X2 U36133 ( .A1(n56377), .A2(n63677), .ZN(n10289) );
  NAND3_X1 U36134 ( .A1(n56373), .A2(n56375), .A3(n56374), .ZN(n63677) );
  NOR2_X2 U36135 ( .A1(n62538), .A2(n64416), .ZN(n50342) );
  AOI21_X2 U36138 ( .A1(n41747), .A2(n41748), .B(n63678), .ZN(n41752) );
  OAI22_X2 U36144 ( .A1(n42940), .A2(n43445), .B1(n41744), .B2(n41745), .ZN(
        n63678) );
  OR2_X2 U36145 ( .A1(n39979), .A2(n39980), .Z(n25458) );
  NAND3_X2 U36148 ( .A1(n18844), .A2(n24692), .A3(n3738), .ZN(n21875) );
  NAND2_X2 U36154 ( .A1(n48189), .A2(n2634), .ZN(n48490) );
  NAND2_X2 U36161 ( .A1(n46148), .A2(n8794), .ZN(n2634) );
  XOR2_X1 U36170 ( .A1(n63680), .A2(n32649), .Z(n18443) );
  XOR2_X1 U36176 ( .A1(n31868), .A2(n22744), .Z(n63680) );
  NAND4_X2 U36185 ( .A1(n5423), .A2(n5424), .A3(n5422), .A4(n30019), .ZN(n5421) );
  XOR2_X1 U36189 ( .A1(n33877), .A2(n4776), .Z(n58407) );
  NAND2_X2 U36191 ( .A1(n23357), .A2(n37227), .ZN(n63682) );
  XOR2_X1 U36199 ( .A1(n32002), .A2(n33856), .Z(n24825) );
  INV_X4 U36215 ( .I(n63683), .ZN(n36979) );
  NAND2_X2 U36216 ( .A1(n43582), .A2(n43573), .ZN(n41963) );
  XOR2_X1 U36221 ( .A1(n11801), .A2(n45249), .Z(n63684) );
  XOR2_X1 U36222 ( .A1(n8384), .A2(n58750), .Z(n63685) );
  NOR3_X2 U36225 ( .A1(n64469), .A2(n64468), .A3(n25290), .ZN(n58524) );
  XOR2_X1 U36230 ( .A1(n51805), .A2(n17370), .Z(n63687) );
  INV_X2 U36237 ( .I(n63688), .ZN(n12924) );
  NOR2_X2 U36238 ( .A1(n20138), .A2(n48742), .ZN(n63688) );
  INV_X2 U36241 ( .I(n65115), .ZN(n16103) );
  XOR2_X1 U36249 ( .A1(n3717), .A2(n38623), .Z(n9219) );
  XOR2_X1 U36250 ( .A1(n23062), .A2(n39618), .Z(n38623) );
  XOR2_X1 U36258 ( .A1(n45320), .A2(n6869), .Z(n6868) );
  XOR2_X1 U36260 ( .A1(n44976), .A2(n60133), .Z(n6869) );
  XOR2_X1 U36263 ( .A1(n24241), .A2(n57931), .Z(n37266) );
  NAND2_X2 U36265 ( .A1(n51863), .A2(n54025), .ZN(n6737) );
  AOI21_X2 U36276 ( .A1(n20268), .A2(n3203), .B(n63692), .ZN(n20266) );
  NOR2_X2 U36280 ( .A1(n59543), .A2(n57280), .ZN(n65056) );
  XOR2_X1 U36281 ( .A1(n11231), .A2(n58859), .Z(n64995) );
  INV_X1 U36283 ( .I(n35898), .ZN(n64410) );
  AND2_X1 U36287 ( .A1(n33570), .A2(n33563), .Z(n33100) );
  XOR2_X1 U36290 ( .A1(n37824), .A2(n63693), .Z(n8516) );
  XOR2_X1 U36295 ( .A1(n15839), .A2(n18132), .Z(n63693) );
  NOR2_X1 U36297 ( .A1(n8248), .A2(n14225), .ZN(n9898) );
  NAND2_X2 U36313 ( .A1(n14226), .A2(n55442), .ZN(n8248) );
  NAND2_X2 U36324 ( .A1(n12497), .A2(n23934), .ZN(n19802) );
  NAND2_X2 U36326 ( .A1(n63694), .A2(n55933), .ZN(n56092) );
  OAI22_X1 U36330 ( .A1(n63696), .A2(n36010), .B1(n35404), .B2(n60374), .ZN(
        n35405) );
  NAND3_X2 U36331 ( .A1(n12272), .A2(n10316), .A3(n43110), .ZN(n45093) );
  NAND3_X2 U36340 ( .A1(n63698), .A2(n46061), .A3(n45624), .ZN(n58987) );
  NAND2_X2 U36351 ( .A1(n59009), .A2(n50674), .ZN(n52751) );
  INV_X2 U36382 ( .I(n7720), .ZN(n43344) );
  NAND2_X2 U36385 ( .A1(n61134), .A2(n43874), .ZN(n7720) );
  XOR2_X1 U36386 ( .A1(n63701), .A2(n12448), .Z(n11973) );
  XOR2_X1 U36388 ( .A1(n24368), .A2(n50632), .Z(n63701) );
  XOR2_X1 U36389 ( .A1(n63702), .A2(n51823), .Z(n23467) );
  XOR2_X1 U36390 ( .A1(n51834), .A2(n51835), .Z(n63702) );
  AOI21_X1 U36391 ( .A1(n55940), .A2(n55939), .B(n12555), .ZN(n63935) );
  NOR2_X2 U36415 ( .A1(n65203), .A2(n43561), .ZN(n43624) );
  NOR2_X2 U36417 ( .A1(n13095), .A2(n13096), .ZN(n24803) );
  OAI21_X2 U36428 ( .A1(n61776), .A2(n50042), .B(n8711), .ZN(n64264) );
  OAI21_X2 U36431 ( .A1(n56992), .A2(n56993), .B(n56991), .ZN(n64829) );
  XOR2_X1 U36438 ( .A1(n1996), .A2(n52441), .Z(n64930) );
  INV_X2 U36443 ( .I(n63704), .ZN(n57408) );
  XOR2_X1 U36452 ( .A1(n61518), .A2(n9155), .Z(n63704) );
  OAI22_X2 U36466 ( .A1(n48597), .A2(n62115), .B1(n47018), .B2(n8012), .ZN(
        n63706) );
  INV_X4 U36469 ( .I(n54902), .ZN(n13671) );
  NOR2_X1 U36472 ( .A1(n54791), .A2(n63707), .ZN(n64008) );
  NOR2_X1 U36473 ( .A1(n63710), .A2(n63709), .ZN(n64310) );
  NAND2_X2 U36475 ( .A1(n21305), .A2(n24099), .ZN(n2743) );
  XNOR2_X1 U36487 ( .A1(n51952), .A2(n1915), .ZN(n57510) );
  XOR2_X1 U36490 ( .A1(n51944), .A2(n7711), .Z(n1915) );
  NAND4_X1 U36497 ( .A1(n56028), .A2(n56027), .A3(n56026), .A4(n56029), .ZN(
        n64140) );
  NOR2_X1 U36500 ( .A1(n56564), .A2(n56397), .ZN(n4943) );
  NAND2_X2 U36510 ( .A1(n25168), .A2(n12605), .ZN(n56397) );
  AOI22_X1 U36513 ( .A1(n54369), .A2(n54393), .B1(n26109), .B2(n54414), .ZN(
        n54372) );
  XOR2_X1 U36514 ( .A1(n63715), .A2(n55340), .Z(Plaintext[109]) );
  NAND3_X2 U36523 ( .A1(n63), .A2(n18284), .A3(n18283), .ZN(n63715) );
  INV_X2 U36524 ( .I(n41904), .ZN(n42269) );
  NOR2_X2 U36539 ( .A1(n25837), .A2(n23155), .ZN(n41904) );
  NAND2_X2 U36556 ( .A1(n2373), .A2(n5402), .ZN(n5401) );
  NOR2_X2 U36572 ( .A1(n2376), .A2(n2378), .ZN(n5402) );
  NAND3_X1 U36585 ( .A1(n62755), .A2(n20140), .A3(n48102), .ZN(n46819) );
  XOR2_X1 U36628 ( .A1(n18889), .A2(n46201), .Z(n63716) );
  NAND3_X1 U36634 ( .A1(n48193), .A2(n18551), .A3(n47490), .ZN(n18550) );
  INV_X2 U36635 ( .I(n56352), .ZN(n1591) );
  NAND3_X2 U36636 ( .A1(n16642), .A2(n17205), .A3(n56232), .ZN(n56352) );
  NAND3_X2 U36653 ( .A1(n19736), .A2(n20352), .A3(n63717), .ZN(n20399) );
  NOR3_X2 U36660 ( .A1(n19460), .A2(n20354), .A3(n53189), .ZN(n63717) );
  NOR2_X1 U36662 ( .A1(n2743), .A2(n6805), .ZN(n59472) );
  XOR2_X1 U36668 ( .A1(n17486), .A2(n63718), .Z(n61546) );
  XOR2_X1 U36671 ( .A1(n37783), .A2(n37782), .Z(n63718) );
  AOI21_X2 U36676 ( .A1(n64495), .A2(n3729), .B(n43269), .ZN(n4329) );
  NAND2_X2 U36684 ( .A1(n8745), .A2(n43124), .ZN(n65217) );
  AOI21_X2 U36690 ( .A1(n16674), .A2(n50364), .B(n63719), .ZN(n24451) );
  NAND2_X2 U36694 ( .A1(n63720), .A2(n24654), .ZN(n49990) );
  AOI21_X2 U36701 ( .A1(n48183), .A2(n58974), .B(n60697), .ZN(n63720) );
  OAI21_X2 U36708 ( .A1(n20598), .A2(n65218), .B(n61796), .ZN(n59543) );
  BUF_X2 U36709 ( .I(n42878), .Z(n63721) );
  OAI21_X2 U36710 ( .A1(n27967), .A2(n57954), .B(n15114), .ZN(n63722) );
  XOR2_X1 U36717 ( .A1(n63903), .A2(n65142), .Z(n51012) );
  NOR2_X2 U36718 ( .A1(n14031), .A2(n14034), .ZN(n24329) );
  BUF_X2 U36734 ( .I(n14643), .Z(n63726) );
  NAND3_X2 U36739 ( .A1(n63727), .A2(n3821), .A3(n3824), .ZN(n29160) );
  NAND3_X1 U36747 ( .A1(n4654), .A2(n62617), .A3(n36751), .ZN(n26017) );
  NAND2_X1 U36763 ( .A1(n32939), .A2(n32937), .ZN(n64469) );
  NAND2_X2 U36774 ( .A1(n63729), .A2(n59918), .ZN(n9532) );
  NOR2_X2 U36779 ( .A1(n59801), .A2(n58450), .ZN(n63729) );
  XOR2_X1 U36781 ( .A1(n46511), .A2(n63731), .Z(n46513) );
  XOR2_X1 U36784 ( .A1(n60740), .A2(n46510), .Z(n63731) );
  XOR2_X1 U36785 ( .A1(n38889), .A2(n65060), .Z(n6291) );
  XOR2_X1 U36790 ( .A1(n38403), .A2(n9930), .Z(n38889) );
  INV_X4 U36810 ( .I(n15784), .ZN(n12962) );
  NAND2_X1 U36811 ( .A1(n63732), .A2(n7), .ZN(n56121) );
  NAND2_X1 U36816 ( .A1(n56118), .A2(n56119), .ZN(n63732) );
  NAND3_X1 U36818 ( .A1(n35436), .A2(n36627), .A3(n1786), .ZN(n35439) );
  XOR2_X1 U36824 ( .A1(n63733), .A2(n50968), .Z(n11166) );
  XOR2_X1 U36825 ( .A1(n51572), .A2(n21133), .Z(n63733) );
  BUF_X2 U36833 ( .I(n6148), .Z(n63734) );
  XOR2_X1 U36841 ( .A1(n63735), .A2(n8033), .Z(n59469) );
  XOR2_X1 U36849 ( .A1(n8035), .A2(n65237), .Z(n63735) );
  OR2_X1 U36850 ( .A1(n64585), .A2(n57015), .Z(n57098) );
  NAND3_X2 U36856 ( .A1(n45454), .A2(n45453), .A3(n15420), .ZN(n2757) );
  OAI22_X1 U36865 ( .A1(n58081), .A2(n61950), .B1(n21471), .B2(n23108), .ZN(
        n41409) );
  NAND2_X2 U36876 ( .A1(n39011), .A2(n17966), .ZN(n23108) );
  NOR2_X2 U36877 ( .A1(n63736), .A2(n39156), .ZN(n41675) );
  XOR2_X1 U36886 ( .A1(n23126), .A2(n15669), .Z(n7991) );
  XOR2_X1 U36889 ( .A1(n21254), .A2(n8737), .Z(n8736) );
  XOR2_X1 U36896 ( .A1(n21253), .A2(n26212), .Z(n21254) );
  XOR2_X1 U36906 ( .A1(n15223), .A2(n63738), .Z(n15257) );
  XOR2_X1 U36909 ( .A1(n18578), .A2(n15222), .Z(n63738) );
  NAND2_X1 U36914 ( .A1(n63741), .A2(n63740), .ZN(n47130) );
  NAND2_X1 U36915 ( .A1(n47125), .A2(n57398), .ZN(n63741) );
  XOR2_X1 U36921 ( .A1(n50570), .A2(n10062), .Z(n17058) );
  INV_X1 U36930 ( .I(n56935), .ZN(n25022) );
  INV_X1 U36931 ( .I(n62987), .ZN(n63744) );
  BUF_X2 U36946 ( .I(n46385), .Z(n63745) );
  OAI22_X1 U36972 ( .A1(n55421), .A2(n55420), .B1(n55418), .B2(n55419), .ZN(
        n63746) );
  OAI21_X2 U36975 ( .A1(n44542), .A2(n44541), .B(n44540), .ZN(n46598) );
  AOI21_X2 U36990 ( .A1(n21173), .A2(n1395), .B(n42685), .ZN(n44542) );
  NAND2_X2 U36997 ( .A1(n22430), .A2(n56342), .ZN(n3613) );
  INV_X2 U37005 ( .I(n43040), .ZN(n42017) );
  NAND2_X2 U37011 ( .A1(n42016), .A2(n63747), .ZN(n43040) );
  INV_X2 U37016 ( .I(n8351), .ZN(n63747) );
  NAND2_X2 U37026 ( .A1(n36150), .A2(n10790), .ZN(n10788) );
  NAND2_X2 U37028 ( .A1(n33522), .A2(n36584), .ZN(n36150) );
  NOR2_X1 U37031 ( .A1(n63748), .A2(n49621), .ZN(n14122) );
  NOR2_X1 U37039 ( .A1(n4190), .A2(n49620), .ZN(n63748) );
  XOR2_X1 U37042 ( .A1(n8123), .A2(n63749), .Z(n8175) );
  AOI22_X2 U37048 ( .A1(n27946), .A2(n28260), .B1(n63750), .B2(n13193), .ZN(
        n27948) );
  NAND2_X1 U37051 ( .A1(n13764), .A2(n27941), .ZN(n63751) );
  XOR2_X1 U37055 ( .A1(n45063), .A2(n22551), .Z(n46630) );
  NAND2_X2 U37070 ( .A1(n42788), .A2(n18847), .ZN(n43023) );
  XOR2_X1 U37072 ( .A1(n2017), .A2(n63753), .Z(n23368) );
  XOR2_X1 U37087 ( .A1(n26142), .A2(n60247), .Z(n63753) );
  NAND4_X2 U37089 ( .A1(n48935), .A2(n48934), .A3(n48936), .A4(n48937), .ZN(
        n18486) );
  NOR2_X2 U37094 ( .A1(n43134), .A2(n43133), .ZN(n57630) );
  NAND2_X2 U37095 ( .A1(n43128), .A2(n4865), .ZN(n43134) );
  NOR2_X2 U37108 ( .A1(n64300), .A2(n63754), .ZN(n60391) );
  XOR2_X1 U37120 ( .A1(n38525), .A2(n64758), .Z(n63755) );
  AOI22_X1 U37128 ( .A1(n42141), .A2(n42142), .B1(n42143), .B2(n42848), .ZN(
        n64526) );
  NOR2_X2 U37133 ( .A1(n42662), .A2(n10004), .ZN(n42848) );
  NOR3_X2 U37143 ( .A1(n65278), .A2(n63757), .A3(n7214), .ZN(n12216) );
  NOR2_X1 U37152 ( .A1(n61674), .A2(n49284), .ZN(n63757) );
  XOR2_X1 U37160 ( .A1(n590), .A2(n63758), .Z(n8293) );
  XOR2_X1 U37168 ( .A1(n39476), .A2(n3975), .Z(n63758) );
  NAND2_X2 U37172 ( .A1(n6379), .A2(n59647), .ZN(n56280) );
  XOR2_X1 U37181 ( .A1(n12586), .A2(n63759), .Z(n32285) );
  XOR2_X1 U37184 ( .A1(n60528), .A2(n602), .Z(n12586) );
  XOR2_X1 U37187 ( .A1(n930), .A2(n23044), .Z(n4145) );
  NAND3_X1 U37197 ( .A1(n14190), .A2(n14191), .A3(n17552), .ZN(n17551) );
  XOR2_X1 U37204 ( .A1(n30828), .A2(n65164), .Z(n24152) );
  XOR2_X1 U37217 ( .A1(n24037), .A2(n50817), .Z(n63763) );
  XNOR2_X1 U37218 ( .A1(n51335), .A2(n52616), .ZN(n51684) );
  NAND3_X2 U37219 ( .A1(n57172), .A2(n59125), .A3(n23086), .ZN(n33531) );
  XOR2_X1 U37226 ( .A1(n26150), .A2(n20593), .Z(n63946) );
  XOR2_X1 U37242 ( .A1(n63764), .A2(n20523), .Z(n64159) );
  XOR2_X1 U37243 ( .A1(n57976), .A2(n57975), .Z(n63764) );
  NAND2_X2 U37258 ( .A1(n24202), .A2(n63765), .ZN(n11034) );
  AOI22_X1 U37260 ( .A1(n46964), .A2(n46963), .B1(n48423), .B2(n48431), .ZN(
        n46967) );
  NAND2_X2 U37261 ( .A1(n14561), .A2(n22570), .ZN(n46963) );
  XOR2_X1 U37286 ( .A1(n63766), .A2(n6963), .Z(n59490) );
  INV_X1 U37291 ( .I(n35470), .ZN(n35469) );
  OAI21_X2 U37294 ( .A1(n6918), .A2(n15720), .B(n61517), .ZN(n35470) );
  NAND2_X1 U37295 ( .A1(n42409), .A2(n42410), .ZN(n63769) );
  XOR2_X1 U37300 ( .A1(n12377), .A2(n45058), .Z(n8285) );
  NAND2_X2 U37302 ( .A1(n41691), .A2(n42401), .ZN(n19490) );
  AND3_X1 U37311 ( .A1(n63772), .A2(n29946), .A3(n29948), .Z(n25371) );
  NAND3_X1 U37312 ( .A1(n8773), .A2(n8522), .A3(n30655), .ZN(n63772) );
  BUF_X2 U37325 ( .I(n1221), .Z(n63773) );
  AOI21_X2 U37331 ( .A1(n1298), .A2(n10882), .B(n63774), .ZN(n42983) );
  NAND3_X1 U37339 ( .A1(n4835), .A2(n25127), .A3(n54344), .ZN(n6672) );
  NAND4_X2 U37343 ( .A1(n6493), .A2(n6496), .A3(n64466), .A4(n6507), .ZN(
        n59299) );
  NAND2_X2 U37357 ( .A1(n6495), .A2(n47233), .ZN(n6507) );
  INV_X1 U37358 ( .I(n5100), .ZN(n63912) );
  NOR2_X2 U37363 ( .A1(n46985), .A2(n46979), .ZN(n47469) );
  XOR2_X1 U37366 ( .A1(n32582), .A2(n3072), .Z(n3071) );
  XOR2_X1 U37370 ( .A1(n13353), .A2(n13464), .Z(n32582) );
  NOR2_X2 U37373 ( .A1(n6130), .A2(n48729), .ZN(n64406) );
  NOR2_X2 U37378 ( .A1(n29456), .A2(n14759), .ZN(n29000) );
  XOR2_X1 U37388 ( .A1(n8021), .A2(n24062), .Z(n44475) );
  NOR2_X2 U37397 ( .A1(n63776), .A2(n58853), .ZN(n64525) );
  INV_X2 U37403 ( .I(n35468), .ZN(n63776) );
  NOR2_X2 U37421 ( .A1(n35986), .A2(n20146), .ZN(n35468) );
  NOR2_X1 U37424 ( .A1(n15539), .A2(n42985), .ZN(n63777) );
  NAND2_X2 U37438 ( .A1(n22228), .A2(n15540), .ZN(n43299) );
  XOR2_X1 U37442 ( .A1(n37555), .A2(n38784), .Z(n38727) );
  XOR2_X1 U37470 ( .A1(n63779), .A2(n7140), .Z(n21792) );
  XOR2_X1 U37472 ( .A1(n44477), .A2(n46252), .Z(n63779) );
  INV_X2 U37481 ( .I(n57845), .ZN(n13412) );
  NAND2_X2 U37485 ( .A1(n63906), .A2(n57937), .ZN(n57845) );
  XOR2_X1 U37494 ( .A1(n63780), .A2(n18849), .Z(n60581) );
  INV_X4 U37505 ( .I(n63968), .ZN(n65283) );
  INV_X2 U37506 ( .I(n14343), .ZN(n1510) );
  NAND2_X2 U37514 ( .A1(n26113), .A2(n59158), .ZN(n14343) );
  NAND2_X1 U37517 ( .A1(n64913), .A2(n64912), .ZN(n15325) );
  AOI21_X2 U37519 ( .A1(n62087), .A2(n48673), .B(n63782), .ZN(n57709) );
  OAI21_X2 U37524 ( .A1(n49358), .A2(n8457), .B(n50046), .ZN(n63782) );
  AND2_X1 U37531 ( .A1(n35552), .A2(n24028), .Z(n64103) );
  NOR2_X2 U37532 ( .A1(n52218), .A2(n22817), .ZN(n55924) );
  NAND2_X2 U37543 ( .A1(n55659), .A2(n23447), .ZN(n52218) );
  XOR2_X1 U37544 ( .A1(n38537), .A2(n39644), .Z(n38729) );
  XOR2_X1 U37547 ( .A1(n63783), .A2(n52530), .Z(n4757) );
  XOR2_X1 U37551 ( .A1(n50615), .A2(n64556), .Z(n63783) );
  XOR2_X1 U37552 ( .A1(n50982), .A2(n50981), .Z(n50983) );
  NAND2_X2 U37553 ( .A1(n10683), .A2(n41469), .ZN(n64308) );
  NAND2_X2 U37554 ( .A1(n63786), .A2(n21324), .ZN(n52248) );
  AND3_X1 U37555 ( .A1(n48477), .A2(n63917), .A3(n63916), .Z(n59980) );
  INV_X2 U37565 ( .I(n63788), .ZN(n35027) );
  XNOR2_X1 U37568 ( .A1(n8558), .A2(n7071), .ZN(n63788) );
  BUF_X2 U37569 ( .I(n46535), .Z(n63789) );
  INV_X1 U37575 ( .I(n58175), .ZN(n56533) );
  NAND2_X1 U37590 ( .A1(n56541), .A2(n2408), .ZN(n58175) );
  NAND4_X2 U37594 ( .A1(n51470), .A2(n51467), .A3(n51469), .A4(n51468), .ZN(
        n63790) );
  INV_X1 U37595 ( .I(n48951), .ZN(n4204) );
  NAND2_X2 U37603 ( .A1(n47977), .A2(n21737), .ZN(n48951) );
  BUF_X2 U37610 ( .I(n33158), .Z(n63791) );
  NAND2_X2 U37611 ( .A1(n60583), .A2(n4689), .ZN(n41347) );
  OR2_X1 U37620 ( .A1(n17744), .A2(n63792), .Z(n10807) );
  NAND3_X1 U37622 ( .A1(n15058), .A2(n33762), .A3(n32958), .ZN(n32959) );
  NAND2_X2 U37636 ( .A1(n23761), .A2(n60960), .ZN(n15058) );
  INV_X4 U37644 ( .I(n22111), .ZN(n57892) );
  NAND2_X2 U37645 ( .A1(n60100), .A2(n5848), .ZN(n22111) );
  AND2_X1 U37647 ( .A1(n43494), .A2(n43926), .Z(n6073) );
  AOI21_X1 U37649 ( .A1(n46884), .A2(n46885), .B(n46894), .ZN(n46886) );
  NAND3_X1 U37651 ( .A1(n46891), .A2(n9730), .A3(n59418), .ZN(n46892) );
  NAND2_X2 U37659 ( .A1(n63796), .A2(n18221), .ZN(n50054) );
  NAND2_X1 U37662 ( .A1(n63798), .A2(n63797), .ZN(n61343) );
  NAND2_X2 U37670 ( .A1(n31842), .A2(n35272), .ZN(n63799) );
  OAI21_X1 U37678 ( .A1(n63801), .A2(n63800), .B(n40260), .ZN(n58139) );
  NAND2_X1 U37685 ( .A1(n52884), .A2(n52886), .ZN(n63894) );
  BUF_X4 U37698 ( .I(n31476), .Z(n37034) );
  NAND2_X2 U37707 ( .A1(n46097), .A2(n8820), .ZN(n47525) );
  NOR2_X2 U37710 ( .A1(n47530), .A2(n48596), .ZN(n46097) );
  XOR2_X1 U37717 ( .A1(n3116), .A2(n61220), .Z(n60383) );
  XOR2_X1 U37738 ( .A1(n18114), .A2(n4890), .Z(n14935) );
  XOR2_X1 U37752 ( .A1(n1749), .A2(n9805), .Z(n6114) );
  XOR2_X1 U37757 ( .A1(n37553), .A2(n103), .Z(n9805) );
  AND2_X1 U37770 ( .A1(n48503), .A2(n48514), .Z(n48510) );
  XOR2_X1 U37815 ( .A1(n6238), .A2(n61657), .Z(n6237) );
  NAND2_X2 U37818 ( .A1(n23746), .A2(n34613), .ZN(n19621) );
  NAND2_X2 U37820 ( .A1(n1281), .A2(n19080), .ZN(n12855) );
  NOR2_X1 U37827 ( .A1(n59927), .A2(n59929), .ZN(n53899) );
  NOR3_X2 U37829 ( .A1(n9947), .A2(n34859), .A3(n1773), .ZN(n3102) );
  NOR2_X2 U37830 ( .A1(n7598), .A2(n22524), .ZN(n9947) );
  NAND2_X1 U37837 ( .A1(n41069), .A2(n40592), .ZN(n63807) );
  NOR2_X2 U37841 ( .A1(n63930), .A2(n42521), .ZN(n25913) );
  NAND3_X2 U37843 ( .A1(n31535), .A2(n31538), .A3(n31534), .ZN(n4515) );
  OAI21_X2 U37845 ( .A1(n31515), .A2(n31516), .B(n1798), .ZN(n31534) );
  AND2_X1 U37859 ( .A1(n54084), .A2(n54589), .Z(n64130) );
  XOR2_X1 U37861 ( .A1(n52407), .A2(n51807), .Z(n12029) );
  XOR2_X1 U37866 ( .A1(n59913), .A2(n20304), .Z(n52407) );
  XOR2_X1 U37867 ( .A1(n63808), .A2(n32422), .Z(n25701) );
  XOR2_X1 U37874 ( .A1(n22440), .A2(n25700), .Z(n63808) );
  XOR2_X1 U37882 ( .A1(n3214), .A2(n63809), .Z(n10311) );
  XOR2_X1 U37883 ( .A1(n6486), .A2(n51644), .Z(n63809) );
  NAND2_X2 U37884 ( .A1(n13163), .A2(n20859), .ZN(n58448) );
  OR2_X1 U37885 ( .A1(n1274), .A2(n41837), .Z(n41871) );
  NOR2_X2 U37889 ( .A1(n9601), .A2(n25849), .ZN(n20978) );
  NAND2_X2 U37891 ( .A1(n6760), .A2(n34622), .ZN(n3560) );
  OAI21_X2 U37895 ( .A1(n44200), .A2(n44199), .B(n44198), .ZN(n63811) );
  OAI21_X1 U37910 ( .A1(n63813), .A2(n63812), .B(n20735), .ZN(n22279) );
  NOR2_X1 U37914 ( .A1(n50740), .A2(n53148), .ZN(n63813) );
  INV_X2 U37915 ( .I(n63814), .ZN(n65271) );
  XOR2_X1 U37916 ( .A1(n6063), .A2(n6062), .Z(n63814) );
  NOR2_X2 U37917 ( .A1(n57369), .A2(n63816), .ZN(n45661) );
  BUF_X2 U37919 ( .I(n23226), .Z(n63817) );
  NAND2_X2 U37920 ( .A1(n56558), .A2(n56369), .ZN(n56377) );
  NOR2_X2 U37923 ( .A1(n56367), .A2(n56368), .ZN(n56558) );
  XOR2_X1 U37925 ( .A1(n51550), .A2(n51549), .Z(n63819) );
  AOI21_X2 U37927 ( .A1(n11221), .A2(n63820), .B(n6491), .ZN(n37851) );
  NOR2_X2 U37930 ( .A1(n1524), .A2(n21536), .ZN(n36292) );
  XOR2_X1 U37939 ( .A1(n51591), .A2(n22455), .Z(n63925) );
  OAI21_X1 U37949 ( .A1(n37404), .A2(n24041), .B(n36818), .ZN(n36823) );
  NAND2_X2 U37956 ( .A1(n35915), .A2(n37405), .ZN(n36818) );
  AND2_X1 U37968 ( .A1(n2962), .A2(n36855), .Z(n15857) );
  NAND3_X1 U37971 ( .A1(n64905), .A2(n35409), .A3(n35408), .ZN(n2962) );
  NAND3_X2 U37976 ( .A1(n44457), .A2(n44456), .A3(n44455), .ZN(n46674) );
  INV_X1 U37983 ( .I(n40356), .ZN(n42460) );
  OR2_X1 U37986 ( .A1(n40356), .A2(n2459), .Z(n42461) );
  NAND4_X1 U37994 ( .A1(n30008), .A2(n18581), .A3(n30760), .A4(n10888), .ZN(
        n30009) );
  XOR2_X1 U38006 ( .A1(n5180), .A2(n7698), .Z(n63821) );
  OAI22_X1 U38009 ( .A1(n14973), .A2(n20432), .B1(n31544), .B2(n31543), .ZN(
        n31549) );
  NOR2_X2 U38012 ( .A1(n7861), .A2(n31533), .ZN(n14973) );
  NOR2_X2 U38015 ( .A1(n1443), .A2(n22498), .ZN(n26765) );
  INV_X2 U38016 ( .I(n7200), .ZN(n55233) );
  NOR2_X1 U38018 ( .A1(n63822), .A2(n7200), .ZN(n15853) );
  NAND2_X2 U38020 ( .A1(n24117), .A2(n22343), .ZN(n7200) );
  NOR2_X2 U38027 ( .A1(n24385), .A2(n63823), .ZN(n24384) );
  OAI22_X2 U38035 ( .A1(n36328), .A2(n36831), .B1(n25339), .B2(n20790), .ZN(
        n63823) );
  NAND2_X1 U38036 ( .A1(n63825), .A2(n63824), .ZN(n45558) );
  NAND2_X1 U38037 ( .A1(n45553), .A2(n47282), .ZN(n63825) );
  NOR2_X2 U38053 ( .A1(n63826), .A2(n906), .ZN(n35266) );
  NAND3_X2 U38055 ( .A1(n13610), .A2(n59873), .A3(n63827), .ZN(n63826) );
  OAI21_X1 U38065 ( .A1(n30610), .A2(n30350), .B(n30616), .ZN(n8267) );
  INV_X1 U38066 ( .I(n41984), .ZN(n63828) );
  NAND2_X1 U38067 ( .A1(n375), .A2(n22370), .ZN(n63877) );
  NAND2_X2 U38068 ( .A1(n43521), .A2(n43508), .ZN(n43199) );
  NAND2_X2 U38081 ( .A1(n28533), .A2(n26431), .ZN(n27249) );
  XOR2_X1 U38088 ( .A1(n59428), .A2(n8285), .Z(n63832) );
  NAND2_X2 U38090 ( .A1(n36838), .A2(n26213), .ZN(n35497) );
  NAND2_X2 U38092 ( .A1(n25205), .A2(n23227), .ZN(n36838) );
  XOR2_X1 U38093 ( .A1(n45358), .A2(n45035), .Z(n61143) );
  XOR2_X1 U38095 ( .A1(n45046), .A2(n46681), .Z(n45358) );
  XOR2_X1 U38096 ( .A1(n57899), .A2(n58921), .Z(n24922) );
  XOR2_X1 U38099 ( .A1(n63833), .A2(n25797), .Z(n666) );
  XOR2_X1 U38102 ( .A1(n60023), .A2(n3072), .Z(n63833) );
  XOR2_X1 U38105 ( .A1(n38838), .A2(n25914), .Z(n59029) );
  XOR2_X1 U38107 ( .A1(n3603), .A2(n38620), .Z(n38838) );
  XOR2_X1 U38108 ( .A1(n63834), .A2(n32354), .Z(n32279) );
  XOR2_X1 U38112 ( .A1(n33143), .A2(n28796), .Z(n63834) );
  NAND2_X1 U38116 ( .A1(n47133), .A2(n47135), .ZN(n64568) );
  NOR2_X1 U38117 ( .A1(n64568), .A2(n61876), .ZN(n25383) );
  NOR2_X2 U38119 ( .A1(n23480), .A2(n46913), .ZN(n57731) );
  BUF_X4 U38121 ( .I(n42619), .Z(n65203) );
  OR2_X1 U38125 ( .A1(n44692), .A2(n63837), .Z(n63836) );
  INV_X1 U38128 ( .I(n40840), .ZN(n41886) );
  XOR2_X1 U38136 ( .A1(n63840), .A2(n61834), .Z(n4413) );
  XOR2_X1 U38139 ( .A1(n5986), .A2(n5987), .Z(n63840) );
  XOR2_X1 U38144 ( .A1(n13156), .A2(n6644), .Z(n52601) );
  NAND2_X1 U38152 ( .A1(n63841), .A2(n11899), .ZN(n11904) );
  XOR2_X1 U38158 ( .A1(n63842), .A2(n53989), .Z(Plaintext[52]) );
  NAND2_X1 U38160 ( .A1(n23685), .A2(n53988), .ZN(n63842) );
  NAND3_X1 U38164 ( .A1(n4188), .A2(n5631), .A3(n30183), .ZN(n10179) );
  NAND2_X2 U38171 ( .A1(n30195), .A2(n21014), .ZN(n4188) );
  INV_X2 U38174 ( .I(n5382), .ZN(n18385) );
  NAND3_X2 U38187 ( .A1(n32839), .A2(n32840), .A3(n32841), .ZN(n5382) );
  OAI22_X2 U38192 ( .A1(n64078), .A2(n1602), .B1(n52266), .B2(n1283), .ZN(
        n19732) );
  NOR2_X2 U38195 ( .A1(n63846), .A2(n23899), .ZN(n41621) );
  NAND3_X2 U38200 ( .A1(n41616), .A2(n41617), .A3(n41615), .ZN(n63846) );
  XOR2_X1 U38206 ( .A1(n22435), .A2(n39714), .Z(n18862) );
  NAND2_X1 U38207 ( .A1(n26253), .A2(n62663), .ZN(n26254) );
  XOR2_X1 U38208 ( .A1(n63881), .A2(n8766), .Z(n65089) );
  BUF_X2 U38211 ( .I(n42262), .Z(n63849) );
  NAND2_X2 U38217 ( .A1(n65057), .A2(n49610), .ZN(n49315) );
  BUF_X2 U38218 ( .I(n1322), .Z(n63850) );
  XOR2_X1 U38220 ( .A1(n59262), .A2(n21339), .Z(n63851) );
  NAND2_X2 U38237 ( .A1(n1838), .A2(n64565), .ZN(n13691) );
  NOR2_X2 U38238 ( .A1(n30343), .A2(n29077), .ZN(n30352) );
  NAND3_X2 U38239 ( .A1(n14359), .A2(n61293), .A3(n55352), .ZN(n18290) );
  BUF_X2 U38241 ( .I(n10428), .Z(n63853) );
  NAND2_X2 U38242 ( .A1(n48107), .A2(n59035), .ZN(n17530) );
  BUF_X2 U38244 ( .I(n23132), .Z(n63854) );
  AND2_X2 U38248 ( .A1(n35629), .A2(n22701), .Z(n8217) );
  NOR2_X2 U38249 ( .A1(n35722), .A2(n25058), .ZN(n63855) );
  AND2_X2 U38264 ( .A1(n56599), .A2(n15536), .Z(n56993) );
  NAND2_X2 U38265 ( .A1(n63857), .A2(n8068), .ZN(n18126) );
  NOR2_X1 U38268 ( .A1(n17043), .A2(n172), .ZN(n63857) );
  NOR2_X2 U38275 ( .A1(n56734), .A2(n56697), .ZN(n56667) );
  NAND2_X1 U38278 ( .A1(n110), .A2(n63859), .ZN(n65063) );
  XOR2_X1 U38280 ( .A1(n38334), .A2(n38160), .Z(n6145) );
  XOR2_X1 U38286 ( .A1(n25995), .A2(n63030), .Z(n38334) );
  XOR2_X1 U38294 ( .A1(n63860), .A2(n30210), .Z(n30291) );
  NAND2_X2 U38296 ( .A1(n16533), .A2(n22436), .ZN(n63913) );
  XOR2_X1 U38300 ( .A1(n63863), .A2(n20435), .Z(n21679) );
  XOR2_X1 U38301 ( .A1(n21344), .A2(n61953), .Z(n63863) );
  OAI21_X1 U38307 ( .A1(n12624), .A2(n50373), .B(n49036), .ZN(n63864) );
  NOR3_X1 U38309 ( .A1(n15617), .A2(n51259), .A3(n18173), .ZN(n22676) );
  OAI22_X2 U38316 ( .A1(n18176), .A2(n56158), .B1(n61697), .B2(n56176), .ZN(
        n15617) );
  NOR2_X2 U38317 ( .A1(n9631), .A2(n63865), .ZN(n13418) );
  NAND2_X2 U38320 ( .A1(n13837), .A2(n55931), .ZN(n55926) );
  NOR2_X2 U38324 ( .A1(n48249), .A2(n44770), .ZN(n46101) );
  BUF_X2 U38332 ( .I(n23086), .Z(n63866) );
  NAND2_X2 U38333 ( .A1(n47382), .A2(n45807), .ZN(n47142) );
  NAND3_X2 U38342 ( .A1(n25064), .A2(n63868), .A3(n48929), .ZN(n23792) );
  XOR2_X1 U38345 ( .A1(n5273), .A2(n63962), .Z(n64319) );
  NAND3_X2 U38347 ( .A1(n1053), .A2(n3001), .A3(n3009), .ZN(n64848) );
  INV_X2 U38351 ( .I(n63870), .ZN(n57701) );
  XOR2_X1 U38352 ( .A1(n59829), .A2(n772), .Z(n63870) );
  OR2_X1 U38353 ( .A1(n3837), .A2(n61851), .Z(n3836) );
  XOR2_X1 U38357 ( .A1(n16632), .A2(n1248), .Z(n4244) );
  XOR2_X1 U38374 ( .A1(n64640), .A2(n7370), .Z(n16632) );
  XOR2_X1 U38384 ( .A1(n22803), .A2(n23264), .Z(n44734) );
  NAND2_X1 U38386 ( .A1(n53754), .A2(n53753), .ZN(n12744) );
  INV_X2 U38396 ( .I(n63874), .ZN(n45591) );
  INV_X2 U38397 ( .I(n63875), .ZN(n14620) );
  AND3_X1 U38410 ( .A1(n14621), .A2(n40587), .A3(n40586), .Z(n63875) );
  BUF_X2 U38425 ( .I(n24007), .Z(n63878) );
  XOR2_X1 U38429 ( .A1(n16025), .A2(n15275), .Z(n7602) );
  NAND2_X1 U38436 ( .A1(n64359), .A2(n38194), .ZN(n4684) );
  NAND2_X2 U38438 ( .A1(n64002), .A2(n3151), .ZN(n7553) );
  NAND3_X2 U38441 ( .A1(n20722), .A2(n5678), .A3(n318), .ZN(n6678) );
  XOR2_X1 U38448 ( .A1(n63925), .A2(n4085), .Z(n63879) );
  OAI21_X2 U38449 ( .A1(n38912), .A2(n19418), .B(n20158), .ZN(n25713) );
  NAND2_X2 U38453 ( .A1(n15594), .A2(n18208), .ZN(n19418) );
  XOR2_X1 U38461 ( .A1(n17231), .A2(n63880), .Z(n17230) );
  XOR2_X1 U38473 ( .A1(n45071), .A2(n45070), .Z(n63880) );
  INV_X2 U38474 ( .I(n56717), .ZN(n56734) );
  NAND3_X2 U38480 ( .A1(n20781), .A2(n56613), .A3(n56614), .ZN(n56717) );
  NAND2_X2 U38483 ( .A1(n18205), .A2(n34203), .ZN(n11020) );
  NOR2_X1 U38488 ( .A1(n59240), .A2(n59534), .ZN(n20887) );
  NAND2_X1 U38491 ( .A1(n5910), .A2(n5909), .ZN(n29463) );
  XOR2_X1 U38492 ( .A1(n31340), .A2(n31341), .Z(n31342) );
  XOR2_X1 U38500 ( .A1(n23204), .A2(n63882), .Z(n63881) );
  BUF_X2 U38507 ( .I(n1575), .Z(n63883) );
  XOR2_X1 U38519 ( .A1(n63887), .A2(n44261), .Z(n60345) );
  XOR2_X1 U38527 ( .A1(n58838), .A2(n11647), .Z(n44261) );
  XOR2_X1 U38528 ( .A1(n63396), .A2(n55242), .Z(n52375) );
  AND2_X1 U38529 ( .A1(n17523), .A2(n359), .Z(n11887) );
  NOR2_X1 U38530 ( .A1(n63023), .A2(n63012), .ZN(n56012) );
  NAND2_X1 U38533 ( .A1(n32952), .A2(n9766), .ZN(n64934) );
  NOR4_X2 U38534 ( .A1(n7718), .A2(n21948), .A3(n21947), .A4(n28284), .ZN(
        n63885) );
  INV_X4 U38535 ( .I(n12287), .ZN(n22169) );
  NAND2_X2 U38536 ( .A1(n12817), .A2(n58943), .ZN(n12287) );
  INV_X2 U38537 ( .I(n63886), .ZN(n24871) );
  XOR2_X1 U38546 ( .A1(n13211), .A2(n11649), .Z(n63887) );
  OR2_X1 U38554 ( .A1(n34783), .A2(n3308), .Z(n12515) );
  NAND2_X1 U38559 ( .A1(n21525), .A2(n17124), .ZN(n64564) );
  NAND2_X2 U38561 ( .A1(n55398), .A2(n55416), .ZN(n55247) );
  INV_X2 U38562 ( .I(n54978), .ZN(n55398) );
  NOR2_X2 U38577 ( .A1(n14919), .A2(n24301), .ZN(n54978) );
  BUF_X2 U38578 ( .I(n11060), .Z(n63888) );
  NOR2_X2 U38581 ( .A1(n10875), .A2(n63889), .ZN(n13862) );
  AND2_X1 U38588 ( .A1(n10878), .A2(n10879), .Z(n63889) );
  BUF_X2 U38599 ( .I(n1562), .Z(n63890) );
  BUF_X2 U38600 ( .I(n29860), .Z(n63891) );
  XOR2_X1 U38603 ( .A1(n23341), .A2(n32183), .Z(n11528) );
  NAND3_X2 U38606 ( .A1(n29923), .A2(n4725), .A3(n29922), .ZN(n32183) );
  NAND4_X2 U38608 ( .A1(n35638), .A2(n35639), .A3(n35637), .A4(n63893), .ZN(
        n44) );
  XOR2_X1 U38610 ( .A1(n63895), .A2(n44261), .Z(n43726) );
  XOR2_X1 U38631 ( .A1(n52331), .A2(n8147), .Z(n49435) );
  NAND2_X2 U38638 ( .A1(n24110), .A2(n47151), .ZN(n52331) );
  NOR2_X2 U38639 ( .A1(n63896), .A2(n5758), .ZN(n5757) );
  BUF_X2 U38650 ( .I(n22431), .Z(n63897) );
  XOR2_X1 U38656 ( .A1(n13555), .A2(n63898), .Z(n4074) );
  XOR2_X1 U38659 ( .A1(n4072), .A2(n38361), .Z(n63898) );
  INV_X1 U38660 ( .I(n37105), .ZN(n63900) );
  NAND2_X2 U38666 ( .A1(n17319), .A2(n47146), .ZN(n21449) );
  XOR2_X1 U38673 ( .A1(n63901), .A2(n53090), .Z(Plaintext[3]) );
  NOR2_X2 U38674 ( .A1(n23759), .A2(n25092), .ZN(n46026) );
  XOR2_X1 U38678 ( .A1(n31485), .A2(n31486), .Z(n31902) );
  XOR2_X1 U38681 ( .A1(n20899), .A2(n23461), .Z(n31485) );
  OR2_X1 U38682 ( .A1(n54343), .A2(n25127), .Z(n6670) );
  NAND3_X2 U38686 ( .A1(n2684), .A2(n2685), .A3(n2683), .ZN(n10351) );
  XOR2_X1 U38703 ( .A1(n63902), .A2(n37849), .Z(n37755) );
  XOR2_X1 U38704 ( .A1(n14424), .A2(n11409), .Z(n63903) );
  XOR2_X1 U38706 ( .A1(n63904), .A2(n32406), .Z(n19879) );
  XOR2_X1 U38710 ( .A1(n33876), .A2(n32204), .Z(n63904) );
  XOR2_X1 U38716 ( .A1(n8606), .A2(n63905), .Z(n58427) );
  NAND2_X2 U38720 ( .A1(n11150), .A2(n24759), .ZN(n15360) );
  NAND4_X2 U38727 ( .A1(n33087), .A2(n33085), .A3(n33086), .A4(n33088), .ZN(
        n33110) );
  NAND3_X2 U38729 ( .A1(n52669), .A2(n61920), .A3(n61516), .ZN(n10515) );
  NAND2_X2 U38731 ( .A1(n58700), .A2(n64461), .ZN(n31356) );
  NOR2_X2 U38735 ( .A1(n1484), .A2(n1666), .ZN(n11183) );
  BUF_X2 U38742 ( .I(n13443), .Z(n63906) );
  CLKBUF_X4 U38743 ( .I(n15237), .Z(n65216) );
  NOR2_X1 U38744 ( .A1(n65114), .A2(n50235), .ZN(n24110) );
  NAND3_X2 U38745 ( .A1(n1000), .A2(n13670), .A3(n63907), .ZN(n4288) );
  NAND2_X1 U38746 ( .A1(n13208), .A2(n43716), .ZN(n63907) );
  XOR2_X1 U38750 ( .A1(n38446), .A2(n63908), .Z(n6711) );
  XOR2_X1 U38766 ( .A1(n6092), .A2(n1412), .Z(n63908) );
  NAND2_X2 U38769 ( .A1(n10869), .A2(n18487), .ZN(n53534) );
  NOR2_X2 U38770 ( .A1(n13370), .A2(n23784), .ZN(n18487) );
  NOR2_X2 U38775 ( .A1(n59043), .A2(n63909), .ZN(n1967) );
  NOR3_X2 U38778 ( .A1(n63911), .A2(n16059), .A3(n63910), .ZN(n20159) );
  NOR2_X2 U38789 ( .A1(n36729), .A2(n22528), .ZN(n63911) );
  AND2_X2 U38791 ( .A1(n4405), .A2(n2974), .Z(n5411) );
  XOR2_X1 U38800 ( .A1(n14626), .A2(n44979), .Z(n60455) );
  OR2_X2 U38801 ( .A1(n22267), .A2(n35490), .Z(n16108) );
  AOI21_X1 U38806 ( .A1(n63912), .A2(n27768), .B(n27767), .ZN(n27770) );
  OAI21_X2 U38813 ( .A1(n4787), .A2(n29530), .B(n60000), .ZN(n5100) );
  INV_X2 U38817 ( .I(n41131), .ZN(n64946) );
  NAND3_X2 U38820 ( .A1(n41090), .A2(n41088), .A3(n41089), .ZN(n41131) );
  OR2_X2 U38821 ( .A1(n59017), .A2(n4570), .Z(n11278) );
  NOR2_X2 U38826 ( .A1(n41289), .A2(n16912), .ZN(n41870) );
  NAND2_X1 U38835 ( .A1(n48473), .A2(n3111), .ZN(n63917) );
  INV_X2 U38844 ( .I(n63918), .ZN(n1094) );
  BUF_X2 U38845 ( .I(n53728), .Z(n63920) );
  NOR2_X2 U38848 ( .A1(n3064), .A2(n63921), .ZN(n65047) );
  XOR2_X1 U38875 ( .A1(n3449), .A2(n59866), .Z(n64403) );
  BUF_X2 U38884 ( .I(n39276), .Z(n63922) );
  NAND3_X2 U38888 ( .A1(n42439), .A2(n42438), .A3(n57208), .ZN(n41823) );
  NOR2_X2 U38889 ( .A1(n41820), .A2(n40314), .ZN(n42439) );
  OAI21_X2 U38890 ( .A1(n42063), .A2(n20219), .B(n43923), .ZN(n20218) );
  XOR2_X1 U38897 ( .A1(n63924), .A2(n53344), .Z(Plaintext[21]) );
  XOR2_X1 U38915 ( .A1(n33067), .A2(n33068), .Z(n15912) );
  OR2_X1 U38917 ( .A1(n60562), .A2(n36436), .Z(n35160) );
  NOR3_X2 U38926 ( .A1(n55350), .A2(n55381), .A3(n61293), .ZN(n55377) );
  OAI21_X2 U38937 ( .A1(n63927), .A2(n9075), .B(n55304), .ZN(n19979) );
  NAND2_X2 U38945 ( .A1(n49521), .A2(n49520), .ZN(n49522) );
  XOR2_X1 U38949 ( .A1(n2522), .A2(n7256), .Z(n65172) );
  AND3_X1 U38952 ( .A1(n63928), .A2(n32361), .A3(n35003), .Z(n32363) );
  NAND3_X1 U38953 ( .A1(n11984), .A2(n25859), .A3(n53665), .ZN(n2837) );
  NAND2_X2 U38954 ( .A1(n53702), .A2(n53690), .ZN(n11984) );
  NAND2_X1 U38992 ( .A1(n63929), .A2(n23935), .ZN(n13372) );
  NAND2_X2 U38995 ( .A1(n53699), .A2(n53672), .ZN(n53655) );
  BUF_X2 U38996 ( .I(n64155), .Z(n63932) );
  NAND2_X2 U39003 ( .A1(n46831), .A2(n21450), .ZN(n46850) );
  INV_X2 U39009 ( .I(n53607), .ZN(n63933) );
  AND2_X1 U39010 ( .A1(n23215), .A2(n36567), .Z(n14093) );
  XOR2_X1 U39023 ( .A1(n45326), .A2(n45145), .Z(n10390) );
  NAND2_X2 U39034 ( .A1(n40689), .A2(n40690), .ZN(n45145) );
  NOR2_X2 U39044 ( .A1(n40971), .A2(n40613), .ZN(n64571) );
  XOR2_X1 U39051 ( .A1(n45426), .A2(n45424), .Z(n14826) );
  XOR2_X1 U39057 ( .A1(n43933), .A2(n45333), .Z(n45426) );
  INV_X1 U39061 ( .I(n60889), .ZN(n63934) );
  XOR2_X1 U39066 ( .A1(n5798), .A2(n2993), .Z(n2992) );
  INV_X2 U39069 ( .I(n31357), .ZN(n34670) );
  NAND2_X1 U39074 ( .A1(n60937), .A2(n21899), .ZN(n31357) );
  INV_X2 U39076 ( .I(n2496), .ZN(n20690) );
  NAND2_X2 U39078 ( .A1(n13389), .A2(n43319), .ZN(n2496) );
  XOR2_X1 U39094 ( .A1(n39658), .A2(n13555), .Z(n2472) );
  AND2_X1 U39095 ( .A1(n56084), .A2(n56106), .Z(n56115) );
  XOR2_X1 U39100 ( .A1(n63936), .A2(n25483), .Z(n6400) );
  XOR2_X1 U39111 ( .A1(n51250), .A2(n8180), .Z(n63936) );
  NOR2_X1 U39119 ( .A1(n58081), .A2(n63937), .ZN(n57245) );
  XOR2_X1 U39129 ( .A1(n63938), .A2(n2131), .Z(n16452) );
  XOR2_X1 U39139 ( .A1(n2132), .A2(n7657), .Z(n63938) );
  INV_X4 U39148 ( .I(n16858), .ZN(n1562) );
  NAND3_X2 U39154 ( .A1(n16860), .A2(n16861), .A3(n16859), .ZN(n16858) );
  NOR2_X2 U39156 ( .A1(n23037), .A2(n25992), .ZN(n64155) );
  NOR3_X2 U39171 ( .A1(n63939), .A2(n30093), .A3(n30193), .ZN(n29742) );
  NOR2_X2 U39173 ( .A1(n63940), .A2(n58863), .ZN(n11069) );
  XOR2_X1 U39176 ( .A1(n14105), .A2(n50614), .Z(n25873) );
  NAND2_X2 U39177 ( .A1(n64430), .A2(n22569), .ZN(n2694) );
  AOI21_X2 U39182 ( .A1(n53455), .A2(n53004), .B(n53003), .ZN(n53012) );
  NAND3_X2 U39190 ( .A1(n13554), .A2(n1644), .A3(n63942), .ZN(n16024) );
  NOR2_X1 U39204 ( .A1(n48070), .A2(n48069), .ZN(n63942) );
  NAND3_X1 U39205 ( .A1(n52748), .A2(n52747), .A3(n52749), .ZN(n25572) );
  OAI21_X1 U39212 ( .A1(n13440), .A2(n50045), .B(n50044), .ZN(n65109) );
  NAND2_X2 U39215 ( .A1(n2068), .A2(n63944), .ZN(n18201) );
  XOR2_X1 U39227 ( .A1(n51818), .A2(n8075), .Z(n4850) );
  NAND2_X2 U39228 ( .A1(n64643), .A2(n7242), .ZN(n8075) );
  NOR2_X2 U39231 ( .A1(n9224), .A2(n25508), .ZN(n59486) );
  BUF_X4 U39233 ( .I(n8305), .Z(n65147) );
  XOR2_X1 U39238 ( .A1(n25395), .A2(n63946), .Z(n2278) );
  XOR2_X1 U39239 ( .A1(n63947), .A2(n23465), .Z(n64026) );
  XOR2_X1 U39241 ( .A1(n16434), .A2(n21369), .Z(n63947) );
  AND2_X1 U39243 ( .A1(n63949), .A2(n59207), .Z(n17004) );
  NAND2_X1 U39248 ( .A1(n48037), .A2(n49010), .ZN(n63949) );
  NOR2_X2 U39261 ( .A1(n9768), .A2(n63950), .ZN(n35341) );
  NAND4_X2 U39264 ( .A1(n34801), .A2(n34802), .A3(n34799), .A4(n34800), .ZN(
        n63950) );
  NAND2_X2 U39265 ( .A1(n63951), .A2(n23910), .ZN(n25193) );
  NAND2_X1 U39271 ( .A1(n20237), .A2(n49827), .ZN(n63951) );
  BUF_X2 U39272 ( .I(n21071), .Z(n63954) );
  OAI22_X1 U39281 ( .A1(n43413), .A2(n43566), .B1(n43418), .B2(n43414), .ZN(
        n43421) );
  NAND3_X2 U39282 ( .A1(n64009), .A2(n60861), .A3(n45903), .ZN(n15866) );
  BUF_X2 U39291 ( .I(n24283), .Z(n63955) );
  NAND3_X1 U39301 ( .A1(n11910), .A2(n62997), .A3(n43626), .ZN(n291) );
  NOR2_X2 U39302 ( .A1(n30623), .A2(n61884), .ZN(n57658) );
  OR2_X2 U39317 ( .A1(n21607), .A2(n6577), .Z(n6576) );
  XOR2_X1 U39330 ( .A1(n18276), .A2(n19145), .Z(n26206) );
  NAND3_X2 U39337 ( .A1(n47792), .A2(n47794), .A3(n47793), .ZN(n51818) );
  NAND2_X2 U39345 ( .A1(n56624), .A2(n56627), .ZN(n56420) );
  NOR2_X1 U39346 ( .A1(n43421), .A2(n63956), .ZN(n6021) );
  OAI22_X1 U39347 ( .A1(n5972), .A2(n43417), .B1(n43418), .B2(n43564), .ZN(
        n63956) );
  NAND2_X1 U39355 ( .A1(n4175), .A2(n63957), .ZN(n8102) );
  NAND2_X2 U39356 ( .A1(n12521), .A2(n1235), .ZN(n4175) );
  NAND2_X2 U39357 ( .A1(n54624), .A2(n54626), .ZN(n63960) );
  INV_X2 U39358 ( .I(n25872), .ZN(n63962) );
  NAND2_X1 U39359 ( .A1(n11327), .A2(n61688), .ZN(n64209) );
  NAND2_X2 U39363 ( .A1(n63963), .A2(n64005), .ZN(n38972) );
  NOR4_X2 U39365 ( .A1(n36989), .A2(n22531), .A3(n36988), .A4(n63964), .ZN(
        n63963) );
  INV_X2 U39381 ( .I(n36991), .ZN(n63964) );
  NOR2_X1 U39382 ( .A1(n10915), .A2(n18202), .ZN(n46965) );
  XOR2_X1 U39385 ( .A1(n59305), .A2(n58330), .Z(n9330) );
  NOR2_X2 U39389 ( .A1(n11229), .A2(n14620), .ZN(n12760) );
  NAND2_X2 U39390 ( .A1(n5323), .A2(n5324), .ZN(n54392) );
  XOR2_X1 U39391 ( .A1(n20668), .A2(n63966), .Z(n24019) );
  INV_X1 U39394 ( .I(n60227), .ZN(n63966) );
  XOR2_X1 U39396 ( .A1(n20905), .A2(n44639), .Z(n60227) );
  NOR3_X2 U39403 ( .A1(n11890), .A2(n11885), .A3(n11891), .ZN(n23895) );
  INV_X2 U39406 ( .I(n63967), .ZN(n57901) );
  XOR2_X1 U39410 ( .A1(n5502), .A2(n58348), .Z(n63967) );
  NOR2_X1 U39417 ( .A1(n46095), .A2(n8696), .ZN(n4773) );
  NOR2_X1 U39425 ( .A1(n21477), .A2(n56907), .ZN(n56914) );
  XOR2_X1 U39429 ( .A1(n23118), .A2(n7971), .Z(n8220) );
  XOR2_X1 U39437 ( .A1(n26246), .A2(n11595), .Z(n23118) );
  AOI21_X1 U39438 ( .A1(n53797), .A2(n53820), .B(n53765), .ZN(n53766) );
  OR2_X2 U39439 ( .A1(n61668), .A2(n47491), .Z(n48194) );
  NOR2_X2 U39445 ( .A1(n24749), .A2(n24748), .ZN(n63968) );
  XOR2_X1 U39468 ( .A1(n63969), .A2(n53805), .Z(Plaintext[44]) );
  AOI21_X1 U39499 ( .A1(n41480), .A2(n41479), .B(n10683), .ZN(n14987) );
  NAND2_X1 U39507 ( .A1(n39982), .A2(n39981), .ZN(n41480) );
  XOR2_X1 U39510 ( .A1(n60616), .A2(n22949), .Z(n12668) );
  OAI21_X2 U39522 ( .A1(n42804), .A2(n13389), .B(n61739), .ZN(n63970) );
  NAND2_X2 U39524 ( .A1(n40301), .A2(n40303), .ZN(n40221) );
  NOR2_X2 U39528 ( .A1(n40304), .A2(n14018), .ZN(n40301) );
  NOR2_X2 U39532 ( .A1(n2925), .A2(n15941), .ZN(n25267) );
  XOR2_X1 U39534 ( .A1(n13016), .A2(n878), .Z(n13015) );
  XOR2_X1 U39542 ( .A1(n2427), .A2(n21369), .Z(n13016) );
  XOR2_X1 U39543 ( .A1(n63971), .A2(n60133), .Z(n4871) );
  XOR2_X1 U39547 ( .A1(n46345), .A2(n8931), .Z(n64021) );
  XOR2_X1 U39553 ( .A1(n7069), .A2(n46655), .Z(n46345) );
  NAND3_X1 U39554 ( .A1(n16748), .A2(n63679), .A3(n1158), .ZN(n14377) );
  AOI21_X2 U39556 ( .A1(n63973), .A2(n24643), .B(n48356), .ZN(n48358) );
  NAND4_X2 U39566 ( .A1(n48354), .A2(n48892), .A3(n48893), .A4(n58306), .ZN(
        n63973) );
  NAND2_X2 U39570 ( .A1(n63974), .A2(n55011), .ZN(n55013) );
  NAND2_X1 U39573 ( .A1(n15681), .A2(n15682), .ZN(n63974) );
  NOR2_X2 U39576 ( .A1(n63975), .A2(n41099), .ZN(n60384) );
  NAND2_X2 U39577 ( .A1(n10434), .A2(n22479), .ZN(n63975) );
  XOR2_X1 U39582 ( .A1(n24731), .A2(n46233), .Z(n44356) );
  NAND2_X2 U39586 ( .A1(n8875), .A2(n8872), .ZN(n46233) );
  NAND3_X1 U39587 ( .A1(n45516), .A2(n45773), .A3(n45515), .ZN(n25457) );
  XOR2_X1 U39600 ( .A1(n50906), .A2(n24621), .Z(n63976) );
  NAND3_X2 U39601 ( .A1(n37204), .A2(n3691), .A3(n18583), .ZN(n37206) );
  XOR2_X1 U39607 ( .A1(n6868), .A2(n63978), .Z(n58404) );
  XOR2_X1 U39612 ( .A1(n6871), .A2(n7880), .Z(n63978) );
  XOR2_X1 U39614 ( .A1(n45387), .A2(n63979), .Z(n17870) );
  XOR2_X1 U39618 ( .A1(n64824), .A2(n58964), .Z(n63979) );
  NAND2_X1 U39621 ( .A1(n53254), .A2(n1164), .ZN(n63980) );
  NOR2_X1 U39622 ( .A1(n19670), .A2(n19671), .ZN(n63981) );
  AND2_X1 U39623 ( .A1(n3907), .A2(n63982), .Z(n36481) );
  NAND2_X2 U39629 ( .A1(n61705), .A2(n26113), .ZN(n42451) );
  NOR2_X2 U39633 ( .A1(n63984), .A2(n61306), .ZN(n3233) );
  NAND3_X2 U39634 ( .A1(n63986), .A2(n2507), .A3(n63985), .ZN(n9274) );
  AND2_X1 U39636 ( .A1(n2508), .A2(n33766), .Z(n63985) );
  INV_X2 U39639 ( .I(n12855), .ZN(n53110) );
  NAND4_X2 U39643 ( .A1(n20361), .A2(n20362), .A3(n63988), .A4(n63987), .ZN(
        n9962) );
  NAND2_X2 U39648 ( .A1(n12100), .A2(n19921), .ZN(n22255) );
  OAI21_X2 U39649 ( .A1(n43563), .A2(n63989), .B(n5001), .ZN(n6784) );
  OAI21_X2 U39650 ( .A1(n3836), .A2(n13505), .B(n3835), .ZN(n13555) );
  XOR2_X1 U39656 ( .A1(n2274), .A2(n8633), .Z(n7063) );
  NAND3_X1 U39658 ( .A1(n518), .A2(n19594), .A3(n4283), .ZN(n53252) );
  AND2_X1 U39662 ( .A1(n28918), .A2(n59710), .Z(n6269) );
  NAND2_X2 U39667 ( .A1(n30343), .A2(n6271), .ZN(n28918) );
  INV_X2 U39670 ( .I(n34836), .ZN(n57860) );
  NAND2_X2 U39672 ( .A1(n17236), .A2(n19007), .ZN(n34836) );
  XOR2_X1 U39677 ( .A1(n63991), .A2(n6484), .Z(n8146) );
  XOR2_X1 U39678 ( .A1(n63992), .A2(n18728), .Z(Plaintext[180]) );
  NOR3_X1 U39693 ( .A1(n12394), .A2(n12399), .A3(n12396), .ZN(n63992) );
  XOR2_X1 U39696 ( .A1(n63993), .A2(n24044), .Z(Plaintext[48]) );
  NAND3_X2 U39699 ( .A1(n61752), .A2(n61897), .A3(n63997), .ZN(n8269) );
  NOR2_X2 U39706 ( .A1(n7252), .A2(n29078), .ZN(n63997) );
  NAND2_X2 U39707 ( .A1(n63998), .A2(n24527), .ZN(n24529) );
  NOR2_X2 U39708 ( .A1(n64000), .A2(n63999), .ZN(n63998) );
  INV_X2 U39712 ( .I(n24530), .ZN(n63999) );
  INV_X1 U39728 ( .I(n47309), .ZN(n64001) );
  NOR2_X1 U39732 ( .A1(n6933), .A2(n64001), .ZN(n6935) );
  NOR3_X2 U39734 ( .A1(n21387), .A2(n25567), .A3(n21386), .ZN(n21385) );
  NOR2_X2 U39752 ( .A1(n11150), .A2(n24759), .ZN(n61601) );
  INV_X2 U39753 ( .I(n19483), .ZN(n11150) );
  XOR2_X1 U39764 ( .A1(n64480), .A2(n8929), .Z(n19483) );
  BUF_X2 U39772 ( .I(n65061), .Z(n64006) );
  NAND3_X2 U39773 ( .A1(n64458), .A2(n35813), .A3(n22797), .ZN(n34718) );
  XOR2_X1 U39774 ( .A1(n38622), .A2(n19145), .Z(n39621) );
  XOR2_X1 U39775 ( .A1(n9255), .A2(n6889), .Z(n38622) );
  NOR3_X2 U39781 ( .A1(n64008), .A2(n64007), .A3(n54797), .ZN(n54876) );
  NOR2_X1 U39785 ( .A1(n19505), .A2(n54794), .ZN(n64007) );
  XOR2_X1 U39789 ( .A1(n26080), .A2(n31587), .Z(n26079) );
  AND2_X1 U39792 ( .A1(n45904), .A2(n45902), .Z(n64009) );
  XOR2_X1 U39794 ( .A1(n45394), .A2(n284), .Z(n64010) );
  AOI21_X2 U39796 ( .A1(n15058), .A2(n58036), .B(n21317), .ZN(n13892) );
  NAND2_X2 U39797 ( .A1(n35055), .A2(n35449), .ZN(n64011) );
  BUF_X2 U39801 ( .I(n1442), .Z(n64012) );
  XOR2_X1 U39805 ( .A1(n15726), .A2(n31327), .Z(n64354) );
  NOR2_X2 U39813 ( .A1(n44226), .A2(n20526), .ZN(n21360) );
  BUF_X2 U39814 ( .I(n45015), .Z(n64013) );
  NOR2_X2 U39818 ( .A1(n7720), .A2(n42750), .ZN(n41596) );
  XOR2_X1 U39819 ( .A1(n64319), .A2(n14720), .Z(n64846) );
  NAND3_X1 U39821 ( .A1(n42560), .A2(n42924), .A3(n57808), .ZN(n64014) );
  NAND2_X2 U39832 ( .A1(n64016), .A2(n7593), .ZN(n36435) );
  NAND2_X1 U39833 ( .A1(n4684), .A2(n4682), .ZN(n64017) );
  NAND2_X1 U39834 ( .A1(n1260), .A2(n55975), .ZN(n55673) );
  NAND2_X2 U39835 ( .A1(n64897), .A2(n17180), .ZN(n53077) );
  XOR2_X1 U39841 ( .A1(n52341), .A2(n19125), .Z(n64769) );
  XOR2_X1 U39843 ( .A1(n52079), .A2(n60857), .Z(n52341) );
  XOR2_X1 U39845 ( .A1(n64018), .A2(n56819), .Z(Plaintext[173]) );
  NAND2_X2 U39851 ( .A1(n48254), .A2(n48642), .ZN(n48253) );
  XOR2_X1 U39853 ( .A1(n64021), .A2(n8929), .Z(n61095) );
  XOR2_X1 U39856 ( .A1(n64022), .A2(n56879), .Z(Plaintext[178]) );
  NAND3_X1 U39857 ( .A1(n56877), .A2(n60956), .A3(n56876), .ZN(n64022) );
  NAND2_X2 U39860 ( .A1(n14905), .A2(n42608), .ZN(n59627) );
  NAND2_X2 U39861 ( .A1(n42600), .A2(n5126), .ZN(n14905) );
  NAND2_X2 U39869 ( .A1(n5335), .A2(n64023), .ZN(n13823) );
  BUF_X2 U39871 ( .I(n35970), .Z(n64024) );
  XOR2_X1 U39873 ( .A1(n4321), .A2(n710), .Z(n64052) );
  NOR2_X2 U39878 ( .A1(n60437), .A2(n36965), .ZN(n35447) );
  XOR2_X1 U39887 ( .A1(n64025), .A2(n38757), .Z(n8196) );
  NAND3_X2 U39890 ( .A1(n30473), .A2(n11495), .A3(n30474), .ZN(n10079) );
  NAND3_X2 U39891 ( .A1(n48809), .A2(n16692), .A3(n17134), .ZN(n2074) );
  INV_X2 U39892 ( .I(n13430), .ZN(n10344) );
  NAND2_X2 U39893 ( .A1(n47786), .A2(n5961), .ZN(n65133) );
  XOR2_X1 U39898 ( .A1(n60174), .A2(n64027), .Z(n25640) );
  XOR2_X1 U39903 ( .A1(n8539), .A2(n61160), .Z(n64027) );
  NOR2_X1 U39916 ( .A1(n21459), .A2(n41914), .ZN(n16151) );
  XOR2_X1 U39922 ( .A1(n64029), .A2(n44907), .Z(n14528) );
  XOR2_X1 U39925 ( .A1(n45004), .A2(n44450), .Z(n64029) );
  AND2_X1 U39931 ( .A1(n31051), .A2(n25112), .Z(n31045) );
  XOR2_X1 U39934 ( .A1(n64032), .A2(n57142), .Z(Plaintext[190]) );
  NAND2_X1 U39937 ( .A1(n59301), .A2(n57140), .ZN(n64032) );
  INV_X2 U39939 ( .I(n64033), .ZN(n24621) );
  XNOR2_X1 U39949 ( .A1(n2950), .A2(n51918), .ZN(n64033) );
  NAND2_X2 U39950 ( .A1(n26522), .A2(n26523), .ZN(n2572) );
  AOI21_X2 U39967 ( .A1(n19789), .A2(n24317), .B(n19791), .ZN(n64034) );
  NAND2_X2 U39970 ( .A1(n50340), .A2(n17900), .ZN(n50348) );
  NAND3_X1 U39972 ( .A1(n16231), .A2(n8343), .A3(n43098), .ZN(n39882) );
  NOR2_X1 U39974 ( .A1(n46014), .A2(n45639), .ZN(n45641) );
  NAND2_X2 U39981 ( .A1(n344), .A2(n47298), .ZN(n46014) );
  OAI21_X2 U39982 ( .A1(n21676), .A2(n21677), .B(n11092), .ZN(n29953) );
  NAND2_X1 U39990 ( .A1(n55009), .A2(n55317), .ZN(n64037) );
  INV_X2 U39992 ( .I(n64041), .ZN(n65279) );
  BUF_X2 U39995 ( .I(n17128), .Z(n64042) );
  NOR3_X2 U39997 ( .A1(n59845), .A2(n64043), .A3(n23620), .ZN(n17873) );
  INV_X1 U40001 ( .I(n64044), .ZN(n64043) );
  OAI21_X1 U40002 ( .A1(n11838), .A2(n15553), .B(n47430), .ZN(n64044) );
  NOR2_X2 U40006 ( .A1(n33109), .A2(n64045), .ZN(n36529) );
  NAND4_X2 U40008 ( .A1(n33107), .A2(n59641), .A3(n33105), .A4(n33108), .ZN(
        n64045) );
  XOR2_X1 U40012 ( .A1(n50923), .A2(n50872), .Z(n57965) );
  XOR2_X1 U40013 ( .A1(n19688), .A2(n20577), .Z(n50923) );
  NAND2_X1 U40014 ( .A1(n18737), .A2(n55262), .ZN(n21249) );
  NAND4_X2 U40021 ( .A1(n32608), .A2(n32609), .A3(n32606), .A4(n64046), .ZN(
        n32610) );
  OAI21_X2 U40024 ( .A1(n32604), .A2(n59174), .B(n32602), .ZN(n64046) );
  OAI21_X2 U40033 ( .A1(n64887), .A2(n48053), .B(n49074), .ZN(n20390) );
  OR2_X2 U40045 ( .A1(n28711), .A2(n63537), .Z(n30659) );
  XOR2_X1 U40048 ( .A1(n44388), .A2(n46377), .Z(n60405) );
  NAND2_X2 U40051 ( .A1(n41374), .A2(n64446), .ZN(n46377) );
  NOR3_X2 U40054 ( .A1(n58529), .A2(n45650), .A3(n58528), .ZN(n64047) );
  NAND3_X1 U40056 ( .A1(n45517), .A2(n58174), .A3(n44680), .ZN(n44066) );
  NOR2_X1 U40061 ( .A1(n49971), .A2(n49970), .ZN(n64433) );
  XOR2_X1 U40070 ( .A1(n64049), .A2(n30599), .Z(n34524) );
  XOR2_X1 U40072 ( .A1(n60755), .A2(n31885), .Z(n64049) );
  XOR2_X1 U40077 ( .A1(n24055), .A2(n64050), .Z(n786) );
  INV_X2 U40079 ( .I(n46164), .ZN(n64050) );
  XOR2_X1 U40087 ( .A1(n64051), .A2(n46628), .Z(n14929) );
  XOR2_X1 U40091 ( .A1(n12769), .A2(n59072), .Z(n64051) );
  OR2_X1 U40101 ( .A1(n12894), .A2(n29254), .Z(n64394) );
  NOR2_X2 U40112 ( .A1(n24682), .A2(n47156), .ZN(n25689) );
  XOR2_X1 U40119 ( .A1(n64052), .A2(n4237), .Z(n4320) );
  XOR2_X1 U40128 ( .A1(n64109), .A2(n23267), .Z(n791) );
  XOR2_X1 U40133 ( .A1(n64054), .A2(n31913), .Z(n10001) );
  XOR2_X1 U40134 ( .A1(n30904), .A2(n30903), .Z(n64054) );
  NAND2_X2 U40135 ( .A1(n20299), .A2(n13655), .ZN(n45536) );
  XOR2_X1 U40153 ( .A1(n64055), .A2(n25324), .Z(n25322) );
  NAND2_X2 U40160 ( .A1(n41306), .A2(n22759), .ZN(n40356) );
  NAND3_X2 U40167 ( .A1(n5308), .A2(n47815), .A3(n5307), .ZN(n5024) );
  OAI22_X1 U40179 ( .A1(n63932), .A2(n28406), .B1(n28007), .B2(n28409), .ZN(
        n64056) );
  BUF_X2 U40195 ( .I(n24987), .Z(n64057) );
  AOI21_X1 U40201 ( .A1(n36366), .A2(n14331), .B(n13557), .ZN(n64058) );
  NOR3_X2 U40213 ( .A1(n64059), .A2(n50157), .A3(n717), .ZN(n50159) );
  NOR2_X1 U40214 ( .A1(n58997), .A2(n52974), .ZN(n64059) );
  NAND3_X2 U40222 ( .A1(n64060), .A2(n14650), .A3(n14651), .ZN(n28948) );
  NAND2_X1 U40227 ( .A1(n27563), .A2(n27564), .ZN(n64060) );
  INV_X2 U40230 ( .I(n7016), .ZN(n32831) );
  AOI21_X2 U40251 ( .A1(n17557), .A2(n41466), .B(n64062), .ZN(n17556) );
  XOR2_X1 U40258 ( .A1(n17781), .A2(n18596), .Z(n32557) );
  INV_X2 U40260 ( .I(n64065), .ZN(n64064) );
  OAI22_X2 U40267 ( .A1(n31281), .A2(n31279), .B1(n31171), .B2(n31284), .ZN(
        n64065) );
  OAI21_X1 U40282 ( .A1(n64066), .A2(n58264), .B(n40143), .ZN(n18714) );
  INV_X2 U40289 ( .I(n48074), .ZN(n48682) );
  NAND2_X2 U40295 ( .A1(n64068), .A2(n1983), .ZN(n33869) );
  OAI21_X2 U40296 ( .A1(n1987), .A2(n1986), .B(n1985), .ZN(n64068) );
  XOR2_X1 U40298 ( .A1(n37792), .A2(n64069), .Z(n8606) );
  XOR2_X1 U40305 ( .A1(n58694), .A2(n13615), .Z(n64069) );
  NAND3_X2 U40311 ( .A1(n1225), .A2(n11727), .A3(n3302), .ZN(n43123) );
  NOR2_X2 U40320 ( .A1(n17199), .A2(n5377), .ZN(n5389) );
  XOR2_X1 U40343 ( .A1(n25245), .A2(n64070), .Z(n58456) );
  XOR2_X1 U40352 ( .A1(n22257), .A2(n32091), .Z(n64070) );
  OR2_X1 U40354 ( .A1(n32791), .A2(n32790), .Z(n64071) );
  NOR2_X2 U40363 ( .A1(n30507), .A2(n64072), .ZN(n19863) );
  NAND4_X2 U40364 ( .A1(n30499), .A2(n30500), .A3(n31252), .A4(n30498), .ZN(
        n64072) );
  XOR2_X1 U40365 ( .A1(n795), .A2(n64073), .Z(n64398) );
  XOR2_X1 U40366 ( .A1(n38976), .A2(n18355), .Z(n64073) );
  NAND3_X2 U40368 ( .A1(n5560), .A2(n5558), .A3(n64074), .ZN(n39254) );
  BUF_X2 U40371 ( .I(n22315), .Z(n64075) );
  XOR2_X1 U40375 ( .A1(n16594), .A2(n9660), .Z(n38891) );
  XOR2_X1 U40376 ( .A1(n32199), .A2(n10057), .Z(n32247) );
  AOI21_X1 U40377 ( .A1(n26831), .A2(n26830), .B(n64079), .ZN(n26832) );
  NAND3_X1 U40378 ( .A1(n26828), .A2(n26901), .A3(n60545), .ZN(n64079) );
  NAND2_X2 U40388 ( .A1(n35267), .A2(n35264), .ZN(n37405) );
  NOR2_X2 U40389 ( .A1(n19198), .A2(n61359), .ZN(n35267) );
  XOR2_X1 U40397 ( .A1(n64081), .A2(n14074), .Z(n14077) );
  XOR2_X1 U40403 ( .A1(n14078), .A2(n14088), .Z(n64081) );
  XOR2_X1 U40405 ( .A1(n18939), .A2(n64082), .Z(n23821) );
  XOR2_X1 U40409 ( .A1(n2191), .A2(n15615), .Z(n18939) );
  INV_X1 U40423 ( .I(n38446), .ZN(n64082) );
  NAND3_X2 U40424 ( .A1(n12650), .A2(n12651), .A3(n57228), .ZN(n54238) );
  OR2_X2 U40428 ( .A1(n15739), .A2(n2665), .Z(n2124) );
  XOR2_X1 U40432 ( .A1(n60173), .A2(n61152), .Z(n15661) );
  NOR2_X2 U40444 ( .A1(n54409), .A2(n11556), .ZN(n54414) );
  INV_X2 U40445 ( .I(n64083), .ZN(n15780) );
  XNOR2_X1 U40450 ( .A1(n58370), .A2(n1132), .ZN(n64083) );
  AOI22_X2 U40452 ( .A1(n20155), .A2(n16152), .B1(n1351), .B2(n64084), .ZN(
        n20153) );
  NOR2_X2 U40455 ( .A1(n40108), .A2(n58351), .ZN(n8479) );
  NAND2_X2 U40456 ( .A1(n64085), .A2(n40943), .ZN(n40108) );
  NAND2_X2 U40458 ( .A1(n57924), .A2(n64086), .ZN(n57922) );
  BUF_X2 U40461 ( .I(n1776), .Z(n64087) );
  NOR2_X2 U40472 ( .A1(n7026), .A2(n19830), .ZN(n17495) );
  NAND2_X1 U40473 ( .A1(n56882), .A2(n56890), .ZN(n64710) );
  XOR2_X1 U40475 ( .A1(n61509), .A2(n10441), .Z(n64088) );
  NAND2_X2 U40476 ( .A1(n65125), .A2(n54966), .ZN(n54624) );
  INV_X4 U40479 ( .I(n6682), .ZN(n9783) );
  NAND2_X2 U40480 ( .A1(n6735), .A2(n5253), .ZN(n6682) );
  AND2_X1 U40488 ( .A1(n499), .A2(n46967), .Z(n15778) );
  NAND3_X1 U40490 ( .A1(n64089), .A2(n18916), .A3(n61992), .ZN(n19113) );
  NAND2_X1 U40494 ( .A1(n17996), .A2(n11850), .ZN(n64089) );
  XOR2_X1 U40502 ( .A1(n64090), .A2(n1576), .Z(Plaintext[162]) );
  OR2_X2 U40505 ( .A1(n20127), .A2(n4054), .Z(n20737) );
  OR2_X2 U40513 ( .A1(n61932), .A2(n20462), .Z(n3641) );
  XOR2_X1 U40526 ( .A1(n25416), .A2(n51067), .Z(n64091) );
  XOR2_X1 U40528 ( .A1(n20899), .A2(n31347), .Z(n31013) );
  NOR2_X2 U40532 ( .A1(n14849), .A2(n14853), .ZN(n20899) );
  NAND3_X1 U40533 ( .A1(n14407), .A2(n12677), .A3(n43958), .ZN(n50) );
  NOR2_X1 U40536 ( .A1(n37364), .A2(n60297), .ZN(n36506) );
  XOR2_X1 U40548 ( .A1(n1617), .A2(n61790), .Z(n64092) );
  NAND3_X2 U40549 ( .A1(n11244), .A2(n40039), .A3(n9798), .ZN(n16643) );
  XOR2_X1 U40551 ( .A1(n9038), .A2(n64094), .Z(n9037) );
  XOR2_X1 U40556 ( .A1(n22338), .A2(n8008), .Z(n52370) );
  BUF_X2 U40557 ( .I(n2876), .Z(n64095) );
  AND2_X1 U40559 ( .A1(n29511), .A2(n2794), .Z(n16161) );
  NOR2_X2 U40560 ( .A1(n12862), .A2(n12861), .ZN(n12879) );
  NAND2_X2 U40563 ( .A1(n64097), .A2(n14487), .ZN(n14335) );
  NOR2_X2 U40565 ( .A1(n58991), .A2(n8133), .ZN(n64097) );
  NOR3_X2 U40569 ( .A1(n48120), .A2(n64099), .A3(n64098), .ZN(n9845) );
  NOR2_X1 U40580 ( .A1(n5705), .A2(n46716), .ZN(n64098) );
  XOR2_X1 U40581 ( .A1(n31581), .A2(n31655), .Z(n31582) );
  BUF_X2 U40601 ( .I(n8006), .Z(n64102) );
  NAND2_X2 U40614 ( .A1(n5090), .A2(n47087), .ZN(n47211) );
  NAND2_X2 U40615 ( .A1(n21231), .A2(n63015), .ZN(n5090) );
  AOI21_X2 U40616 ( .A1(n41316), .A2(n1333), .B(n64104), .ZN(n41318) );
  BUF_X2 U40621 ( .I(n43254), .Z(n64105) );
  XOR2_X1 U40631 ( .A1(n22287), .A2(n24224), .Z(n22286) );
  NAND3_X1 U40639 ( .A1(n49771), .A2(n64107), .A3(n64106), .ZN(n23980) );
  NAND2_X1 U40644 ( .A1(n49769), .A2(n63724), .ZN(n64106) );
  NOR2_X1 U40650 ( .A1(n22022), .A2(n64108), .ZN(n64107) );
  INV_X2 U40657 ( .I(n2817), .ZN(n39258) );
  XOR2_X1 U40663 ( .A1(n64110), .A2(n38088), .Z(n2817) );
  INV_X2 U40665 ( .I(n21348), .ZN(n64110) );
  XOR2_X1 U40675 ( .A1(n64111), .A2(n6872), .Z(n44978) );
  XOR2_X1 U40679 ( .A1(n22975), .A2(n9434), .Z(n64111) );
  OR2_X2 U40681 ( .A1(n20770), .A2(n64518), .Z(n60969) );
  NAND2_X2 U40682 ( .A1(n64943), .A2(n18753), .ZN(n18752) );
  AOI21_X1 U40691 ( .A1(n56971), .A2(n56970), .B(n65163), .ZN(n56972) );
  XOR2_X1 U40692 ( .A1(n23402), .A2(n43731), .Z(n43732) );
  INV_X2 U40719 ( .I(n55295), .ZN(n1458) );
  NAND2_X2 U40722 ( .A1(n23982), .A2(n55494), .ZN(n55295) );
  XOR2_X1 U40723 ( .A1(n32542), .A2(n58440), .Z(n31600) );
  NAND2_X2 U40730 ( .A1(n28694), .A2(n14546), .ZN(n58440) );
  NAND3_X2 U40734 ( .A1(n48577), .A2(n48573), .A3(n46771), .ZN(n48558) );
  NOR2_X2 U40741 ( .A1(n48085), .A2(n46770), .ZN(n48573) );
  XOR2_X1 U40742 ( .A1(n5798), .A2(n32371), .Z(n4887) );
  XOR2_X1 U40747 ( .A1(n31673), .A2(n5342), .Z(n32371) );
  OR3_X1 U40764 ( .A1(n56982), .A2(n7835), .A3(n64113), .Z(n24618) );
  NAND2_X2 U40765 ( .A1(n23901), .A2(n3086), .ZN(n29949) );
  NOR3_X1 U40767 ( .A1(n8776), .A2(n8779), .A3(n27964), .ZN(n8775) );
  OAI21_X2 U40768 ( .A1(n64115), .A2(n18408), .B(n52176), .ZN(n8250) );
  NOR2_X1 U40770 ( .A1(n57084), .A2(n59954), .ZN(n64116) );
  AND2_X1 U40771 ( .A1(n11395), .A2(n63454), .Z(n28749) );
  BUF_X2 U40776 ( .I(n10339), .Z(n64117) );
  XOR2_X1 U40781 ( .A1(n64120), .A2(n15629), .Z(n6688) );
  XOR2_X1 U40785 ( .A1(n62740), .A2(n24347), .Z(n64120) );
  NAND2_X2 U40786 ( .A1(n60202), .A2(n8772), .ZN(n30654) );
  INV_X2 U40791 ( .I(n46097), .ZN(n64122) );
  XOR2_X1 U40794 ( .A1(n15149), .A2(n50718), .Z(n52155) );
  XOR2_X1 U40799 ( .A1(n20621), .A2(n15505), .Z(n15149) );
  NOR2_X2 U40801 ( .A1(n64264), .A2(n48945), .ZN(n8715) );
  XOR2_X1 U40806 ( .A1(n51850), .A2(n51849), .Z(n51853) );
  XOR2_X1 U40821 ( .A1(n22057), .A2(n22056), .Z(n51850) );
  OAI21_X2 U40822 ( .A1(n13729), .A2(n13727), .B(n64123), .ZN(n19891) );
  OAI22_X2 U40829 ( .A1(n13566), .A2(n46872), .B1(n45490), .B2(n45489), .ZN(
        n10910) );
  NAND2_X2 U40831 ( .A1(n64124), .A2(n56394), .ZN(n12550) );
  NOR3_X2 U40833 ( .A1(n41494), .A2(n41492), .A3(n64126), .ZN(n58241) );
  OAI22_X2 U40837 ( .A1(n43703), .A2(n41490), .B1(n43395), .B2(n20242), .ZN(
        n64126) );
  NOR2_X2 U40838 ( .A1(n9551), .A2(n58884), .ZN(n55144) );
  NAND2_X2 U40839 ( .A1(n52131), .A2(n55456), .ZN(n55679) );
  XOR2_X1 U40851 ( .A1(n22141), .A2(n51750), .Z(n24786) );
  XOR2_X1 U40861 ( .A1(n15505), .A2(n6597), .Z(n6595) );
  NOR2_X1 U40864 ( .A1(n54083), .A2(n64130), .ZN(n54085) );
  XOR2_X1 U40865 ( .A1(n64131), .A2(n2550), .Z(n3101) );
  XOR2_X1 U40867 ( .A1(n64749), .A2(n23821), .Z(n15616) );
  BUF_X2 U40868 ( .I(n12539), .Z(n64132) );
  AOI22_X2 U40873 ( .A1(n64133), .A2(n1523), .B1(n5479), .B2(n59154), .ZN(
        n59942) );
  INV_X2 U40876 ( .I(n22081), .ZN(n64133) );
  NAND2_X2 U40877 ( .A1(n24050), .A2(n15247), .ZN(n22081) );
  XOR2_X1 U40878 ( .A1(n64134), .A2(n63035), .Z(n26097) );
  XOR2_X1 U40879 ( .A1(n61082), .A2(n65151), .Z(n65014) );
  XOR2_X1 U40888 ( .A1(n10300), .A2(n64136), .Z(n10600) );
  XOR2_X1 U40889 ( .A1(n8462), .A2(n18956), .Z(n64136) );
  NAND3_X2 U40890 ( .A1(n14772), .A2(n14771), .A3(n48241), .ZN(n14770) );
  NOR2_X1 U40891 ( .A1(n20999), .A2(n49996), .ZN(n60526) );
  NAND2_X2 U40897 ( .A1(n13393), .A2(n43448), .ZN(n8247) );
  NOR3_X2 U40900 ( .A1(n64138), .A2(n64137), .A3(n2633), .ZN(n61577) );
  NOR2_X2 U40902 ( .A1(n48487), .A2(n48584), .ZN(n64137) );
  NAND2_X2 U40904 ( .A1(n5534), .A2(n58169), .ZN(n36401) );
  NAND3_X2 U40908 ( .A1(n12938), .A2(n12936), .A3(n64139), .ZN(n12933) );
  AOI22_X1 U40909 ( .A1(n35195), .A2(n2899), .B1(n19265), .B2(n12935), .ZN(
        n64139) );
  XOR2_X1 U40913 ( .A1(n13999), .A2(n13997), .Z(n46679) );
  XOR2_X1 U40916 ( .A1(n64140), .A2(n60797), .Z(Plaintext[139]) );
  XOR2_X1 U40925 ( .A1(n6717), .A2(n64141), .Z(n64834) );
  XOR2_X1 U40937 ( .A1(n51590), .A2(n64142), .Z(n64141) );
  INV_X2 U40942 ( .I(n51388), .ZN(n64142) );
  XOR2_X1 U40944 ( .A1(n64144), .A2(n741), .Z(n15041) );
  XOR2_X1 U40947 ( .A1(n21105), .A2(n21740), .Z(n64144) );
  OAI21_X1 U40949 ( .A1(n52849), .A2(n52854), .B(n60498), .ZN(n52852) );
  OAI21_X1 U40952 ( .A1(n64146), .A2(n22494), .B(n9304), .ZN(n10279) );
  OR2_X1 U40964 ( .A1(n141), .A2(n36197), .Z(n64146) );
  BUF_X2 U40965 ( .I(n205), .Z(n64147) );
  XOR2_X1 U40971 ( .A1(n64149), .A2(n56008), .Z(Plaintext[138]) );
  NAND4_X2 U40977 ( .A1(n56007), .A2(n56006), .A3(n56004), .A4(n56005), .ZN(
        n64149) );
  XOR2_X1 U40978 ( .A1(n14740), .A2(n8810), .Z(n16581) );
  NAND2_X2 U40983 ( .A1(n8707), .A2(n8704), .ZN(n8810) );
  AND3_X1 U40987 ( .A1(n33391), .A2(n157), .A3(n33654), .Z(n31714) );
  XOR2_X1 U40988 ( .A1(n32720), .A2(n31708), .Z(n64245) );
  NAND2_X2 U41003 ( .A1(n58172), .A2(n64150), .ZN(n35899) );
  AND2_X1 U41015 ( .A1(n25819), .A2(n25820), .Z(n64150) );
  NAND2_X1 U41016 ( .A1(n28101), .A2(n28100), .ZN(n64686) );
  XOR2_X1 U41017 ( .A1(n30907), .A2(n64755), .Z(n59460) );
  NAND4_X2 U41023 ( .A1(n2102), .A2(n60248), .A3(n3108), .A4(n60249), .ZN(
        n30907) );
  XOR2_X1 U41024 ( .A1(n32571), .A2(n64151), .Z(n3275) );
  XOR2_X1 U41030 ( .A1(n8529), .A2(n31555), .Z(n64151) );
  NOR3_X2 U41032 ( .A1(n17655), .A2(n17654), .A3(n56873), .ZN(n64152) );
  XOR2_X1 U41037 ( .A1(n33839), .A2(n31554), .Z(n22361) );
  INV_X2 U41039 ( .I(n8810), .ZN(n33839) );
  NOR3_X2 U41040 ( .A1(n3548), .A2(n64153), .A3(n61842), .ZN(n3547) );
  NOR2_X1 U41047 ( .A1(n35183), .A2(n36262), .ZN(n33413) );
  XOR2_X1 U41049 ( .A1(n2748), .A2(n12835), .Z(n64157) );
  XOR2_X1 U41051 ( .A1(n12569), .A2(n12568), .Z(n25362) );
  XOR2_X1 U41067 ( .A1(n32321), .A2(n32320), .Z(n32726) );
  NAND2_X2 U41070 ( .A1(n45746), .A2(n9299), .ZN(n25691) );
  NOR2_X2 U41073 ( .A1(n45521), .A2(n44064), .ZN(n9299) );
  XOR2_X1 U41083 ( .A1(n39359), .A2(n64159), .Z(n13937) );
  NAND2_X2 U41097 ( .A1(n11279), .A2(n6689), .ZN(n18278) );
  INV_X2 U41101 ( .I(n43203), .ZN(n43059) );
  XOR2_X1 U41110 ( .A1(n11554), .A2(n44807), .Z(n2482) );
  XOR2_X1 U41111 ( .A1(n43209), .A2(n43208), .Z(n44807) );
  XOR2_X1 U41117 ( .A1(n64160), .A2(n32587), .Z(n31405) );
  XOR2_X1 U41119 ( .A1(n63050), .A2(n31401), .Z(n64160) );
  NAND2_X2 U41126 ( .A1(n24318), .A2(n57048), .ZN(n57050) );
  XOR2_X1 U41139 ( .A1(n64163), .A2(n50786), .Z(n9355) );
  XOR2_X1 U41140 ( .A1(n50783), .A2(n50784), .Z(n64163) );
  NAND3_X2 U41143 ( .A1(n35691), .A2(n35688), .A3(n24688), .ZN(n33307) );
  XOR2_X1 U41154 ( .A1(n33031), .A2(n24315), .Z(n64165) );
  NAND2_X2 U41165 ( .A1(n52706), .A2(n56547), .ZN(n21330) );
  OAI21_X2 U41169 ( .A1(n55171), .A2(n26093), .B(n2784), .ZN(n55111) );
  NAND2_X2 U41174 ( .A1(n7890), .A2(n55165), .ZN(n55171) );
  XOR2_X1 U41180 ( .A1(n51331), .A2(n51332), .Z(n51333) );
  AOI22_X1 U41183 ( .A1(n25586), .A2(n29898), .B1(n24556), .B2(n29902), .ZN(
        n11531) );
  NAND4_X1 U41186 ( .A1(n19714), .A2(n19294), .A3(n49049), .A4(n47921), .ZN(
        n17680) );
  BUF_X2 U41187 ( .I(n2810), .Z(n64167) );
  OAI21_X2 U41197 ( .A1(n46042), .A2(n64168), .B(n46041), .ZN(n46044) );
  NAND2_X2 U41214 ( .A1(n40775), .A2(n40774), .ZN(n61442) );
  NOR2_X2 U41231 ( .A1(n1732), .A2(n39957), .ZN(n40439) );
  NAND2_X2 U41232 ( .A1(n25870), .A2(n64171), .ZN(n60830) );
  NAND2_X2 U41233 ( .A1(n43380), .A2(n42630), .ZN(n42760) );
  XOR2_X1 U41234 ( .A1(n3843), .A2(n64173), .Z(n16873) );
  XOR2_X1 U41240 ( .A1(n11506), .A2(n32293), .Z(n64173) );
  BUF_X2 U41242 ( .I(n27114), .Z(n64174) );
  NAND2_X2 U41245 ( .A1(n62391), .A2(n59627), .ZN(n64175) );
  NAND2_X2 U41251 ( .A1(n5317), .A2(n36030), .ZN(n35576) );
  NAND3_X1 U41252 ( .A1(n14230), .A2(n1208), .A3(n28059), .ZN(n30320) );
  XOR2_X1 U41253 ( .A1(n64177), .A2(n13539), .Z(n6816) );
  OR4_X1 U41255 ( .A1(n7618), .A2(n40592), .A3(n63119), .A4(n9790), .Z(n39965)
         );
  OAI21_X2 U41258 ( .A1(n7594), .A2(n29050), .B(n64178), .ZN(n2840) );
  NAND3_X2 U41263 ( .A1(n57496), .A2(n57436), .A3(n30184), .ZN(n64178) );
  NAND3_X2 U41265 ( .A1(n34116), .A2(n32870), .A3(n33953), .ZN(n34126) );
  NOR2_X1 U41270 ( .A1(n64710), .A2(n22276), .ZN(n22274) );
  XOR2_X1 U41274 ( .A1(n37631), .A2(n38145), .Z(n648) );
  NAND2_X1 U41281 ( .A1(n64180), .A2(n64179), .ZN(n58520) );
  NAND2_X1 U41288 ( .A1(n36381), .A2(n36380), .ZN(n64180) );
  AOI21_X2 U41292 ( .A1(n64182), .A2(n46716), .B(n48530), .ZN(n8751) );
  INV_X2 U41293 ( .I(n20879), .ZN(n18483) );
  NOR2_X2 U41307 ( .A1(n61659), .A2(n18068), .ZN(n20879) );
  NOR2_X2 U41318 ( .A1(n15715), .A2(n1364), .ZN(n22110) );
  NAND2_X1 U41323 ( .A1(n40435), .A2(n64184), .ZN(n16929) );
  NAND2_X2 U41324 ( .A1(n36070), .A2(n62934), .ZN(n36308) );
  NOR2_X1 U41338 ( .A1(n4984), .A2(n55021), .ZN(n55027) );
  OAI21_X1 U41339 ( .A1(n8700), .A2(n16695), .B(n24299), .ZN(n8699) );
  XOR2_X1 U41340 ( .A1(n64185), .A2(n55107), .Z(Plaintext[95]) );
  NOR2_X1 U41345 ( .A1(n392), .A2(n55105), .ZN(n64185) );
  NAND2_X2 U41346 ( .A1(n35962), .A2(n35971), .ZN(n33716) );
  XOR2_X1 U41352 ( .A1(n50843), .A2(n16744), .Z(n50898) );
  XOR2_X1 U41367 ( .A1(n22406), .A2(n19029), .Z(n50842) );
  AOI22_X2 U41368 ( .A1(n27263), .A2(n27264), .B1(n27973), .B2(n27981), .ZN(
        n27267) );
  INV_X1 U41376 ( .I(n7499), .ZN(n64191) );
  OR2_X1 U41378 ( .A1(n27974), .A2(n64191), .Z(n57750) );
  NOR2_X2 U41380 ( .A1(n60347), .A2(n57234), .ZN(n22093) );
  INV_X4 U41383 ( .I(n64192), .ZN(n24196) );
  NOR2_X2 U41387 ( .A1(n29160), .A2(n29159), .ZN(n64192) );
  NAND2_X2 U41391 ( .A1(n21738), .A2(n64193), .ZN(n42914) );
  AND3_X1 U41394 ( .A1(n38599), .A2(n38598), .A3(n39137), .Z(n64193) );
  XOR2_X1 U41428 ( .A1(n15647), .A2(n64194), .Z(n59575) );
  XOR2_X1 U41436 ( .A1(n58442), .A2(n37680), .Z(n15647) );
  NAND2_X2 U41438 ( .A1(n5284), .A2(n64195), .ZN(n50378) );
  NOR2_X2 U41443 ( .A1(n61779), .A2(n64196), .ZN(n64195) );
  XOR2_X1 U41446 ( .A1(n64197), .A2(n24392), .Z(n24475) );
  NAND2_X2 U41451 ( .A1(n8044), .A2(n48414), .ZN(n19589) );
  INV_X2 U41456 ( .I(n64198), .ZN(n15870) );
  NOR2_X2 U41471 ( .A1(n35901), .A2(n24118), .ZN(n64198) );
  NOR2_X2 U41475 ( .A1(n33668), .A2(n64199), .ZN(n60758) );
  NAND2_X1 U41476 ( .A1(n59321), .A2(n33666), .ZN(n64199) );
  INV_X1 U41486 ( .I(n31709), .ZN(n64200) );
  AND2_X1 U41487 ( .A1(n12768), .A2(n64200), .Z(n31712) );
  XOR2_X1 U41488 ( .A1(n51389), .A2(n51490), .Z(n23312) );
  XOR2_X1 U41489 ( .A1(n25061), .A2(n50581), .Z(n51389) );
  NOR2_X2 U41492 ( .A1(n26066), .A2(n16294), .ZN(n26065) );
  NOR2_X2 U41509 ( .A1(n25451), .A2(n47070), .ZN(n26066) );
  NAND2_X2 U41519 ( .A1(n33349), .A2(n8780), .ZN(n16957) );
  XOR2_X1 U41521 ( .A1(n17324), .A2(n64201), .Z(n17322) );
  XOR2_X1 U41526 ( .A1(n16252), .A2(n32719), .Z(n64201) );
  AOI21_X1 U41527 ( .A1(n33556), .A2(n64202), .B(n33555), .ZN(n33557) );
  NAND3_X1 U41532 ( .A1(n33551), .A2(n33552), .A3(n8366), .ZN(n64202) );
  XOR2_X1 U41533 ( .A1(n64203), .A2(n38514), .Z(n38516) );
  XOR2_X1 U41537 ( .A1(n39273), .A2(n58473), .Z(n64203) );
  XOR2_X1 U41540 ( .A1(n17980), .A2(n25211), .Z(n19273) );
  XOR2_X1 U41541 ( .A1(n64786), .A2(n18057), .Z(n17980) );
  NAND2_X2 U41547 ( .A1(n1426), .A2(n23717), .ZN(n22835) );
  NAND2_X1 U41554 ( .A1(n10415), .A2(n38684), .ZN(n38685) );
  NOR2_X1 U41560 ( .A1(n4198), .A2(n9190), .ZN(n38684) );
  INV_X4 U41567 ( .I(n43561), .ZN(n43679) );
  XOR2_X1 U41578 ( .A1(n64204), .A2(n52226), .Z(Plaintext[120]) );
  NAND3_X2 U41582 ( .A1(n13386), .A2(n22656), .A3(n13388), .ZN(n15306) );
  NAND2_X1 U41585 ( .A1(n41959), .A2(n22710), .ZN(n64957) );
  NAND3_X1 U41592 ( .A1(n47293), .A2(n47298), .A3(n65095), .ZN(n45637) );
  NOR2_X2 U41595 ( .A1(n32704), .A2(n64205), .ZN(n12110) );
  NAND2_X2 U41596 ( .A1(n7536), .A2(n59298), .ZN(n64205) );
  AOI21_X1 U41599 ( .A1(n25666), .A2(n18869), .B(n61804), .ZN(n57421) );
  NAND2_X2 U41601 ( .A1(n6095), .A2(n54461), .ZN(n9082) );
  NAND3_X2 U41602 ( .A1(n17571), .A2(n17569), .A3(n17567), .ZN(n64599) );
  NAND2_X1 U41603 ( .A1(n49072), .A2(n23532), .ZN(n49077) );
  NOR3_X2 U41610 ( .A1(n57884), .A2(n50225), .A3(n50223), .ZN(n64207) );
  NAND3_X1 U41617 ( .A1(n52685), .A2(n52687), .A3(n56988), .ZN(n51439) );
  XOR2_X1 U41621 ( .A1(n44885), .A2(n44978), .Z(n65094) );
  XOR2_X1 U41631 ( .A1(n21895), .A2(n9861), .Z(n44885) );
  XOR2_X1 U41633 ( .A1(n7688), .A2(n64208), .Z(n7721) );
  XOR2_X1 U41645 ( .A1(n7686), .A2(n24184), .Z(n64208) );
  XOR2_X1 U41652 ( .A1(n3322), .A2(n64210), .Z(n64591) );
  XOR2_X1 U41656 ( .A1(n64211), .A2(n9376), .Z(n3379) );
  XOR2_X1 U41660 ( .A1(n10351), .A2(n39619), .Z(n64211) );
  NAND2_X2 U41675 ( .A1(n64212), .A2(n124), .ZN(n59477) );
  NAND2_X1 U41677 ( .A1(n28585), .A2(n28586), .ZN(n64212) );
  NAND2_X1 U41679 ( .A1(n42571), .A2(n64213), .ZN(n42575) );
  NOR2_X1 U41680 ( .A1(n43147), .A2(n64214), .ZN(n64213) );
  INV_X1 U41688 ( .I(n43161), .ZN(n64214) );
  NOR2_X2 U41689 ( .A1(n20601), .A2(n11179), .ZN(n43147) );
  XOR2_X1 U41690 ( .A1(n64215), .A2(n16561), .Z(n60649) );
  XOR2_X1 U41693 ( .A1(n26088), .A2(n38478), .Z(n64215) );
  NAND2_X2 U41701 ( .A1(n17542), .A2(n61277), .ZN(n10507) );
  NOR2_X2 U41703 ( .A1(n5059), .A2(n4386), .ZN(n25426) );
  NAND2_X2 U41706 ( .A1(n58612), .A2(n65240), .ZN(n5059) );
  NAND2_X2 U41707 ( .A1(n28269), .A2(n64216), .ZN(n58214) );
  NOR2_X2 U41711 ( .A1(n13098), .A2(n27413), .ZN(n64216) );
  XOR2_X1 U41713 ( .A1(n64217), .A2(n31702), .Z(n32307) );
  NOR2_X2 U41724 ( .A1(n64219), .A2(n64218), .ZN(n2736) );
  XOR2_X1 U41728 ( .A1(n64221), .A2(n61837), .Z(n64937) );
  NAND2_X1 U41729 ( .A1(n64222), .A2(n64963), .ZN(n24603) );
  NAND2_X1 U41734 ( .A1(n13690), .A2(n29091), .ZN(n64222) );
  NAND2_X1 U41735 ( .A1(n996), .A2(n11817), .ZN(n42090) );
  NAND2_X1 U41736 ( .A1(n42400), .A2(n42401), .ZN(n64223) );
  NAND3_X1 U41739 ( .A1(n3352), .A2(n3350), .A3(n64414), .ZN(n59336) );
  NAND2_X2 U41741 ( .A1(n56182), .A2(n5172), .ZN(n17961) );
  NOR2_X2 U41744 ( .A1(n30017), .A2(n64228), .ZN(n31433) );
  NAND3_X2 U41745 ( .A1(n30009), .A2(n30011), .A3(n30010), .ZN(n64228) );
  AND3_X1 U41750 ( .A1(n30843), .A2(n63691), .A3(n64229), .Z(n17853) );
  BUF_X2 U41754 ( .I(n56863), .Z(n64230) );
  NAND4_X2 U41755 ( .A1(n3964), .A2(n3963), .A3(n1015), .A4(n5948), .ZN(n3962)
         );
  NOR2_X2 U41756 ( .A1(n64232), .A2(n61797), .ZN(n5196) );
  INV_X1 U41760 ( .I(n64233), .ZN(n64232) );
  OAI21_X1 U41765 ( .A1(n5418), .A2(n56595), .B(n55957), .ZN(n64233) );
  NAND2_X2 U41778 ( .A1(n20129), .A2(n56596), .ZN(n19521) );
  NAND3_X1 U41782 ( .A1(n7485), .A2(n48421), .A3(n18202), .ZN(n17224) );
  BUF_X2 U41785 ( .I(n9608), .Z(n64234) );
  XOR2_X1 U41790 ( .A1(n51317), .A2(n64235), .Z(n20116) );
  XOR2_X1 U41796 ( .A1(n51199), .A2(n51130), .Z(n64235) );
  NAND2_X2 U41802 ( .A1(n60329), .A2(n22894), .ZN(n64462) );
  XOR2_X1 U41807 ( .A1(n10685), .A2(n10197), .Z(n32885) );
  NOR2_X2 U41808 ( .A1(n19793), .A2(n58343), .ZN(n64239) );
  BUF_X2 U41809 ( .I(n38591), .Z(n64241) );
  NAND2_X2 U41813 ( .A1(n6230), .A2(n6231), .ZN(n60259) );
  BUF_X4 U41814 ( .I(n34203), .Z(n35986) );
  INV_X1 U41815 ( .I(n3385), .ZN(n64243) );
  AND2_X2 U41816 ( .A1(n2428), .A2(n64243), .Z(n20734) );
  XOR2_X1 U41821 ( .A1(n64245), .A2(n17821), .Z(n21402) );
  NOR2_X2 U41822 ( .A1(n2435), .A2(n15245), .ZN(n8261) );
  NAND2_X2 U41823 ( .A1(n15310), .A2(n15703), .ZN(n2435) );
  NOR2_X2 U41826 ( .A1(n25201), .A2(n5531), .ZN(n60652) );
  NOR2_X2 U41833 ( .A1(n11590), .A2(n473), .ZN(n40424) );
  XOR2_X1 U41836 ( .A1(n39564), .A2(n920), .Z(n38635) );
  XOR2_X1 U41838 ( .A1(n362), .A2(n12151), .Z(n5586) );
  XOR2_X1 U41841 ( .A1(n64252), .A2(n55603), .Z(Plaintext[119]) );
  NAND4_X1 U41846 ( .A1(n22851), .A2(n55602), .A3(n55600), .A4(n55601), .ZN(
        n64252) );
  OR2_X1 U41848 ( .A1(n47810), .A2(n47797), .Z(n47703) );
  INV_X2 U41850 ( .I(n42803), .ZN(n10897) );
  NAND2_X2 U41854 ( .A1(n13389), .A2(n61739), .ZN(n42803) );
  BUF_X2 U41859 ( .I(n49610), .Z(n64256) );
  NAND3_X2 U41862 ( .A1(n64257), .A2(n14854), .A3(n28999), .ZN(n14853) );
  OAI21_X1 U41863 ( .A1(n29460), .A2(n7403), .B(n28997), .ZN(n64257) );
  OAI21_X1 U41864 ( .A1(n61822), .A2(n55343), .B(n9424), .ZN(n9402) );
  NAND4_X2 U41866 ( .A1(n47909), .A2(n47908), .A3(n47910), .A4(n47907), .ZN(
        n47911) );
  NOR2_X2 U41870 ( .A1(n55595), .A2(n1592), .ZN(n55568) );
  NOR2_X2 U41872 ( .A1(n55485), .A2(n55484), .ZN(n55595) );
  XOR2_X1 U41873 ( .A1(n64260), .A2(n64259), .Z(n64635) );
  OR3_X1 U41879 ( .A1(n64261), .A2(n52494), .A3(n21395), .Z(n21394) );
  NOR2_X1 U41884 ( .A1(n52493), .A2(n52952), .ZN(n64261) );
  INV_X2 U41896 ( .I(n64262), .ZN(n57353) );
  NAND2_X2 U41901 ( .A1(n56370), .A2(n56234), .ZN(n64262) );
  BUF_X2 U41905 ( .I(n34886), .Z(n64263) );
  AOI21_X2 U41912 ( .A1(n48274), .A2(n18690), .B(n64265), .ZN(n13386) );
  NAND2_X2 U41913 ( .A1(n13387), .A2(n48276), .ZN(n64265) );
  BUF_X2 U41918 ( .I(n15246), .Z(n64268) );
  OR2_X2 U41920 ( .A1(n40962), .A2(n40970), .Z(n21960) );
  NAND2_X2 U41922 ( .A1(n60049), .A2(n54046), .ZN(n54053) );
  NOR2_X2 U41926 ( .A1(n14103), .A2(n53915), .ZN(n54046) );
  XOR2_X1 U41930 ( .A1(n1520), .A2(n17846), .Z(n4543) );
  XOR2_X1 U41939 ( .A1(n4727), .A2(n1833), .Z(n31290) );
  XOR2_X1 U41946 ( .A1(n64270), .A2(n61911), .Z(n64575) );
  XOR2_X1 U41949 ( .A1(n11973), .A2(n52570), .Z(n64270) );
  NAND4_X2 U41952 ( .A1(n12210), .A2(n12208), .A3(n53126), .A4(n64271), .ZN(
        n9791) );
  AOI22_X1 U41953 ( .A1(n61690), .A2(n12111), .B1(n23153), .B2(n53145), .ZN(
        n64271) );
  AND2_X1 U41964 ( .A1(n24574), .A2(n33801), .Z(n64272) );
  XOR2_X1 U41972 ( .A1(n64273), .A2(n38290), .Z(n38291) );
  OR3_X1 U41975 ( .A1(n20297), .A2(n20298), .A3(n64274), .Z(n61018) );
  INV_X2 U41984 ( .I(n63853), .ZN(n64274) );
  XOR2_X1 U41985 ( .A1(n64275), .A2(n17340), .Z(n11419) );
  XOR2_X1 U41988 ( .A1(n20334), .A2(n20335), .Z(n64275) );
  OR2_X1 U41993 ( .A1(n23139), .A2(n54504), .Z(n54505) );
  BUF_X2 U41994 ( .I(n34309), .Z(n64276) );
  BUF_X2 U41996 ( .I(n41164), .Z(n64277) );
  NAND2_X1 U41997 ( .A1(n64279), .A2(n46887), .ZN(n64278) );
  OAI22_X1 U41999 ( .A1(n46886), .A2(n9730), .B1(n46885), .B2(n47262), .ZN(
        n64279) );
  INV_X1 U42000 ( .I(n46887), .ZN(n64281) );
  NAND2_X2 U42001 ( .A1(n29516), .A2(n17412), .ZN(n64282) );
  BUF_X2 U42002 ( .I(n23119), .Z(n64283) );
  NAND3_X2 U42005 ( .A1(n64284), .A2(n43556), .A3(n64957), .ZN(n17302) );
  NOR2_X2 U42006 ( .A1(n64477), .A2(n18146), .ZN(n38469) );
  BUF_X2 U42022 ( .I(n37874), .Z(n64285) );
  NOR2_X2 U42025 ( .A1(n15528), .A2(n15529), .ZN(n15527) );
  XOR2_X1 U42027 ( .A1(n64287), .A2(n14873), .Z(n19233) );
  XOR2_X1 U42045 ( .A1(n15074), .A2(n64638), .Z(n64287) );
  NOR2_X1 U42046 ( .A1(n49501), .A2(n49491), .ZN(n19263) );
  OR2_X2 U42047 ( .A1(n63043), .A2(n6055), .Z(n8012) );
  XOR2_X1 U42061 ( .A1(n64289), .A2(n29407), .Z(Plaintext[31]) );
  NOR2_X2 U42068 ( .A1(n20493), .A2(n64290), .ZN(n10939) );
  NAND3_X2 U42074 ( .A1(n20492), .A2(n20468), .A3(n3025), .ZN(n64290) );
  NOR2_X2 U42080 ( .A1(n23877), .A2(n65230), .ZN(n64291) );
  OAI21_X1 U42082 ( .A1(n60730), .A2(n15832), .B(n22263), .ZN(n47077) );
  NOR2_X2 U42085 ( .A1(n14314), .A2(n49910), .ZN(n22263) );
  NOR2_X2 U42092 ( .A1(n65262), .A2(n20619), .ZN(n64292) );
  XOR2_X1 U42096 ( .A1(n23535), .A2(n38433), .Z(n11098) );
  AOI21_X2 U42097 ( .A1(n26222), .A2(n37376), .B(n9992), .ZN(n23535) );
  OR2_X1 U42098 ( .A1(n47152), .A2(n46484), .Z(n64293) );
  INV_X2 U42112 ( .I(n25076), .ZN(n1623) );
  NAND3_X2 U42114 ( .A1(n64294), .A2(n3702), .A3(n3700), .ZN(n25076) );
  AND2_X1 U42123 ( .A1(n3698), .A2(n1100), .Z(n64294) );
  BUF_X2 U42131 ( .I(n18335), .Z(n64295) );
  XOR2_X1 U42141 ( .A1(n46386), .A2(n44938), .Z(n44496) );
  NAND3_X1 U42144 ( .A1(n17013), .A2(n213), .A3(n214), .ZN(n64909) );
  XOR2_X1 U42154 ( .A1(n38836), .A2(n39222), .Z(n37697) );
  NAND2_X2 U42164 ( .A1(n57831), .A2(n5384), .ZN(n38836) );
  XOR2_X1 U42170 ( .A1(n64298), .A2(n50134), .Z(n50150) );
  XOR2_X1 U42173 ( .A1(n50115), .A2(n51011), .Z(n64298) );
  AOI21_X2 U42176 ( .A1(n36645), .A2(n33943), .B(n33942), .ZN(n39670) );
  NOR2_X2 U42182 ( .A1(n4666), .A2(n53570), .ZN(n53676) );
  XOR2_X1 U42184 ( .A1(n64299), .A2(n2028), .Z(n14721) );
  OR2_X2 U42194 ( .A1(n15616), .A2(n39324), .Z(n12592) );
  XOR2_X1 U42201 ( .A1(n50686), .A2(n64301), .Z(n14636) );
  XOR2_X1 U42202 ( .A1(n60312), .A2(n9878), .Z(n64301) );
  OAI22_X1 U42208 ( .A1(n52912), .A2(n52911), .B1(n52914), .B2(n52913), .ZN(
        n61023) );
  NOR3_X2 U42212 ( .A1(n22930), .A2(n49149), .A3(n23242), .ZN(n25951) );
  NOR2_X2 U42220 ( .A1(n23074), .A2(n56863), .ZN(n56882) );
  XOR2_X1 U42224 ( .A1(n60559), .A2(n64305), .Z(n64698) );
  XOR2_X1 U42225 ( .A1(n64306), .A2(n37647), .Z(n64305) );
  NOR3_X2 U42234 ( .A1(n64310), .A2(n15849), .A3(n64309), .ZN(n19870) );
  NAND2_X2 U42240 ( .A1(n9642), .A2(n10450), .ZN(n64309) );
  XOR2_X1 U42249 ( .A1(n14588), .A2(n1757), .Z(n6026) );
  XOR2_X1 U42250 ( .A1(n38573), .A2(n22435), .Z(n12940) );
  XOR2_X1 U42256 ( .A1(n38771), .A2(n4667), .Z(n64973) );
  XOR2_X1 U42261 ( .A1(n61944), .A2(n53284), .Z(n38771) );
  NAND2_X1 U42269 ( .A1(n15493), .A2(n64889), .ZN(n15491) );
  NAND3_X1 U42270 ( .A1(n65129), .A2(n12312), .A3(n1336), .ZN(n43463) );
  XOR2_X1 U42272 ( .A1(n60869), .A2(n31749), .Z(n64311) );
  XOR2_X1 U42274 ( .A1(n10351), .A2(n55624), .Z(n13733) );
  NAND2_X2 U42275 ( .A1(n46840), .A2(n45796), .ZN(n64313) );
  XOR2_X1 U42279 ( .A1(n25326), .A2(n38276), .Z(n38285) );
  AOI21_X2 U42283 ( .A1(n17426), .A2(n34759), .B(n17425), .ZN(n64314) );
  INV_X2 U42288 ( .I(n46843), .ZN(n47418) );
  NAND2_X1 U42292 ( .A1(n23666), .A2(n47680), .ZN(n46843) );
  NOR2_X2 U42297 ( .A1(n10225), .A2(n1387), .ZN(n12648) );
  OR2_X1 U42305 ( .A1(n8047), .A2(n45203), .Z(n47705) );
  INV_X2 U42306 ( .I(n47495), .ZN(n47503) );
  NAND2_X2 U42315 ( .A1(n45484), .A2(n58189), .ZN(n47495) );
  NAND2_X1 U42317 ( .A1(n43257), .A2(n64315), .ZN(n10303) );
  NOR2_X1 U42319 ( .A1(n20526), .A2(n1495), .ZN(n64315) );
  INV_X4 U42323 ( .I(n42914), .ZN(n20180) );
  NAND2_X2 U42330 ( .A1(n46982), .A2(n47472), .ZN(n45746) );
  BUF_X2 U42340 ( .I(n52609), .Z(n64316) );
  OAI21_X1 U42344 ( .A1(n48913), .A2(n48912), .B(n50550), .ZN(n58499) );
  XOR2_X1 U42348 ( .A1(n64317), .A2(n9319), .Z(n24012) );
  XOR2_X1 U42349 ( .A1(n33070), .A2(n12781), .Z(n64317) );
  XOR2_X1 U42355 ( .A1(n11071), .A2(n51541), .Z(n51550) );
  XOR2_X1 U42360 ( .A1(n9416), .A2(n58945), .Z(n51541) );
  NOR2_X1 U42363 ( .A1(n29002), .A2(n2796), .ZN(n64695) );
  NAND3_X1 U42367 ( .A1(n41259), .A2(n41258), .A3(n42251), .ZN(n41260) );
  AOI21_X2 U42372 ( .A1(n2463), .A2(n43230), .B(n64318), .ZN(n43774) );
  NAND4_X2 U42380 ( .A1(n43228), .A2(n16090), .A3(n2197), .A4(n43229), .ZN(
        n64318) );
  XOR2_X1 U42382 ( .A1(n13685), .A2(n13390), .Z(n64320) );
  NOR4_X2 U42384 ( .A1(n39856), .A2(n64321), .A3(n39853), .A4(n39854), .ZN(
        n39859) );
  NAND3_X2 U42387 ( .A1(n49506), .A2(n49507), .A3(n19437), .ZN(n51033) );
  NOR2_X2 U42393 ( .A1(n9293), .A2(n4626), .ZN(n49506) );
  OAI21_X1 U42394 ( .A1(n8471), .A2(n29139), .B(n29138), .ZN(n64322) );
  NAND2_X2 U42396 ( .A1(n24196), .A2(n23589), .ZN(n30213) );
  XOR2_X1 U42397 ( .A1(n14969), .A2(n37885), .Z(n64325) );
  AND2_X1 U42400 ( .A1(n29142), .A2(n27292), .Z(n27931) );
  XOR2_X1 U42402 ( .A1(n25970), .A2(n52174), .Z(n20883) );
  XOR2_X1 U42403 ( .A1(n32619), .A2(n1213), .Z(n32284) );
  XOR2_X1 U42405 ( .A1(n60525), .A2(n32710), .Z(n32619) );
  NOR2_X1 U42407 ( .A1(n64327), .A2(n59630), .ZN(n55861) );
  NAND3_X1 U42408 ( .A1(n55845), .A2(n55843), .A3(n55844), .ZN(n64327) );
  NOR2_X2 U42410 ( .A1(n49858), .A2(n25352), .ZN(n14488) );
  NAND2_X2 U42411 ( .A1(n9845), .A2(n61313), .ZN(n49858) );
  XOR2_X1 U42422 ( .A1(n19647), .A2(n64328), .Z(n22191) );
  XOR2_X1 U42423 ( .A1(n19711), .A2(n6649), .Z(n64328) );
  OAI21_X2 U42427 ( .A1(n65127), .A2(n64329), .B(n58683), .ZN(n3743) );
  NAND2_X2 U42430 ( .A1(n11716), .A2(n64176), .ZN(n17606) );
  NAND4_X2 U42435 ( .A1(n27638), .A2(n7211), .A3(n27639), .A4(n27637), .ZN(
        n10599) );
  OAI21_X2 U42439 ( .A1(n64336), .A2(n64335), .B(n58657), .ZN(n49305) );
  BUF_X2 U42440 ( .I(n27876), .Z(n64337) );
  NAND3_X2 U42442 ( .A1(n33388), .A2(n33386), .A3(n33387), .ZN(n36247) );
  NAND2_X2 U42443 ( .A1(n24948), .A2(n4270), .ZN(n3993) );
  BUF_X2 U42444 ( .I(n49496), .Z(n64341) );
  NAND2_X2 U42445 ( .A1(n12768), .A2(n18884), .ZN(n34134) );
  NAND3_X1 U42447 ( .A1(n19663), .A2(n33663), .A3(n157), .ZN(n18908) );
  INV_X2 U42448 ( .I(n9286), .ZN(n16798) );
  XOR2_X1 U42449 ( .A1(n8864), .A2(n65214), .Z(n9286) );
  NOR3_X2 U42455 ( .A1(n28420), .A2(n64594), .A3(n28403), .ZN(n16861) );
  NAND2_X2 U42465 ( .A1(n10894), .A2(n21347), .ZN(n7365) );
  XOR2_X1 U42467 ( .A1(n31153), .A2(n30950), .Z(n20083) );
  NAND2_X2 U42478 ( .A1(n10824), .A2(n10971), .ZN(n10970) );
  NOR2_X2 U42483 ( .A1(n40151), .A2(n3361), .ZN(n10824) );
  NAND2_X2 U42484 ( .A1(n23976), .A2(n23977), .ZN(n38999) );
  NOR2_X2 U42487 ( .A1(n58988), .A2(n25354), .ZN(n23976) );
  INV_X2 U42489 ( .I(n64343), .ZN(n1929) );
  INV_X2 U42490 ( .I(n49748), .ZN(n49466) );
  NAND2_X2 U42499 ( .A1(n16596), .A2(n15781), .ZN(n49748) );
  NOR3_X2 U42500 ( .A1(n13697), .A2(n17697), .A3(n16257), .ZN(n64344) );
  BUF_X2 U42509 ( .I(n3618), .Z(n64346) );
  NAND2_X1 U42510 ( .A1(n14785), .A2(n14787), .ZN(n14784) );
  NOR2_X2 U42515 ( .A1(n18357), .A2(n65074), .ZN(n64347) );
  XOR2_X1 U42518 ( .A1(n2963), .A2(n64348), .Z(n14087) );
  XOR2_X1 U42522 ( .A1(n12044), .A2(n64349), .Z(n64348) );
  INV_X2 U42523 ( .I(n8021), .ZN(n64349) );
  XOR2_X1 U42526 ( .A1(n64350), .A2(n959), .Z(n3295) );
  XOR2_X1 U42546 ( .A1(n12015), .A2(n58035), .Z(n64350) );
  XOR2_X1 U42550 ( .A1(n64351), .A2(n59619), .Z(n64882) );
  NOR2_X1 U42556 ( .A1(n12768), .A2(n157), .ZN(n33398) );
  OAI22_X1 U42558 ( .A1(n60343), .A2(n59056), .B1(n8012), .B2(n62115), .ZN(
        n64352) );
  NAND2_X2 U42567 ( .A1(n43383), .A2(n11197), .ZN(n42630) );
  NAND2_X1 U42568 ( .A1(n58380), .A2(n56205), .ZN(n56622) );
  NAND2_X2 U42570 ( .A1(n4888), .A2(n49466), .ZN(n49458) );
  BUF_X2 U42575 ( .I(n41289), .Z(n64353) );
  XOR2_X1 U42594 ( .A1(n64354), .A2(n23152), .Z(n33030) );
  XOR2_X1 U42598 ( .A1(n31680), .A2(n32324), .Z(n31681) );
  XOR2_X1 U42606 ( .A1(n64035), .A2(n31344), .Z(n18336) );
  NOR2_X2 U42610 ( .A1(n45698), .A2(n45697), .ZN(n21071) );
  NAND3_X2 U42613 ( .A1(n10195), .A2(n40391), .A3(n40392), .ZN(n42636) );
  OAI21_X2 U42615 ( .A1(n55342), .A2(n58828), .B(n19797), .ZN(n18285) );
  OAI22_X2 U42628 ( .A1(n28565), .A2(n30610), .B1(n28564), .B2(n62495), .ZN(
        n65131) );
  XOR2_X1 U42636 ( .A1(n38744), .A2(n64357), .Z(n18998) );
  XOR2_X1 U42642 ( .A1(n25885), .A2(n39595), .Z(n64357) );
  XOR2_X1 U42650 ( .A1(n51521), .A2(n51057), .Z(n25416) );
  XOR2_X1 U42654 ( .A1(n14500), .A2(n52630), .Z(n51521) );
  OAI22_X1 U42656 ( .A1(n55980), .A2(n14884), .B1(n55981), .B2(n56227), .ZN(
        n55983) );
  NAND2_X2 U42658 ( .A1(n34443), .A2(n33583), .ZN(n35650) );
  NOR3_X2 U42659 ( .A1(n64361), .A2(n35084), .A3(n35083), .ZN(n6907) );
  OR2_X1 U42660 ( .A1(n35082), .A2(n37098), .Z(n64361) );
  XOR2_X1 U42661 ( .A1(n64362), .A2(n25407), .Z(n14997) );
  XOR2_X1 U42668 ( .A1(n60711), .A2(n38726), .Z(n64362) );
  NAND3_X1 U42671 ( .A1(n29153), .A2(n65183), .A3(n29150), .ZN(n26378) );
  NOR2_X2 U42676 ( .A1(n57874), .A2(n58156), .ZN(n23585) );
  BUF_X2 U42692 ( .I(n21791), .Z(n64364) );
  INV_X1 U42702 ( .I(n10292), .ZN(n13831) );
  XOR2_X1 U42704 ( .A1(n12543), .A2(n12540), .Z(n3685) );
  NOR3_X2 U42707 ( .A1(n12794), .A2(n21318), .A3(n46820), .ZN(n5284) );
  NAND3_X2 U42708 ( .A1(n36155), .A2(n15161), .A3(n64368), .ZN(n39714) );
  NAND2_X2 U42729 ( .A1(n57216), .A2(n58537), .ZN(n64369) );
  XOR2_X1 U42746 ( .A1(n64370), .A2(n22922), .Z(n14058) );
  NAND2_X2 U42751 ( .A1(n7075), .A2(n15599), .ZN(n22922) );
  AND2_X2 U42755 ( .A1(n33763), .A2(n13559), .Z(n35004) );
  OR2_X1 U42757 ( .A1(n19231), .A2(n12830), .Z(n35183) );
  NAND4_X2 U42761 ( .A1(n29346), .A2(n29347), .A3(n64376), .A4(n64375), .ZN(
        n29365) );
  OAI21_X2 U42762 ( .A1(n29341), .A2(n29342), .B(n29351), .ZN(n64375) );
  OAI21_X2 U42767 ( .A1(n29336), .A2(n29337), .B(n29335), .ZN(n64376) );
  OR2_X1 U42770 ( .A1(n14212), .A2(n1970), .Z(n28478) );
  INV_X2 U42789 ( .I(n23188), .ZN(n64379) );
  NAND3_X1 U42796 ( .A1(n15775), .A2(n22436), .A3(n16533), .ZN(n48204) );
  NAND2_X2 U42797 ( .A1(n36946), .A2(n34914), .ZN(n130) );
  XOR2_X1 U42805 ( .A1(n64382), .A2(n20614), .Z(n16622) );
  XOR2_X1 U42808 ( .A1(n64383), .A2(n33144), .Z(n29204) );
  XOR2_X1 U42812 ( .A1(n22244), .A2(n29075), .Z(n64383) );
  XNOR2_X1 U42817 ( .A1(n57405), .A2(n3927), .ZN(n64393) );
  XOR2_X1 U42821 ( .A1(n64384), .A2(n17365), .Z(n7862) );
  XOR2_X1 U42829 ( .A1(n62923), .A2(n14085), .Z(n64384) );
  XOR2_X1 U42835 ( .A1(n39497), .A2(n64385), .Z(n57563) );
  XOR2_X1 U42838 ( .A1(n37418), .A2(n18031), .Z(n64385) );
  NAND2_X2 U42841 ( .A1(n45510), .A2(n64386), .ZN(n44775) );
  OR2_X2 U42842 ( .A1(n26105), .A2(n5293), .Z(n20925) );
  NOR2_X2 U42850 ( .A1(n34784), .A2(n64387), .ZN(n7661) );
  INV_X2 U42851 ( .I(n12519), .ZN(n64387) );
  NAND2_X2 U42853 ( .A1(n40203), .A2(n58369), .ZN(n40198) );
  XOR2_X1 U42856 ( .A1(n51507), .A2(n51807), .Z(n26144) );
  XOR2_X1 U42861 ( .A1(n51730), .A2(n51191), .Z(n51507) );
  XOR2_X1 U42870 ( .A1(n44904), .A2(n7385), .Z(n7684) );
  XOR2_X1 U42875 ( .A1(n26191), .A2(n44184), .Z(n44904) );
  AOI21_X1 U42877 ( .A1(n64389), .A2(n27195), .B(n27194), .ZN(n27200) );
  AOI22_X1 U42882 ( .A1(n13047), .A2(n28348), .B1(n296), .B2(n27522), .ZN(
        n64389) );
  BUF_X2 U42895 ( .I(n1742), .Z(n64390) );
  NOR2_X2 U42896 ( .A1(n12152), .A2(n23698), .ZN(n40829) );
  BUF_X2 U42899 ( .I(n13306), .Z(n64391) );
  XOR2_X1 U42900 ( .A1(n9529), .A2(n24794), .Z(n24796) );
  NOR2_X2 U42902 ( .A1(n57698), .A2(n57396), .ZN(n24230) );
  NAND3_X2 U42903 ( .A1(n64392), .A2(n35191), .A3(n35192), .ZN(n37285) );
  OAI21_X1 U42906 ( .A1(n35529), .A2(n19559), .B(n35188), .ZN(n64392) );
  INV_X2 U42920 ( .I(n3925), .ZN(n15552) );
  XOR2_X1 U42921 ( .A1(n3929), .A2(n64393), .Z(n3925) );
  AND3_X1 U42925 ( .A1(n28944), .A2(n64394), .A3(n28945), .Z(n15546) );
  NAND2_X2 U42926 ( .A1(n61225), .A2(n64395), .ZN(n17016) );
  NOR3_X2 U42928 ( .A1(n7436), .A2(n12483), .A3(n12484), .ZN(n64395) );
  NAND2_X2 U42932 ( .A1(n16766), .A2(n7824), .ZN(n8120) );
  NAND2_X1 U42942 ( .A1(n63849), .A2(n42261), .ZN(n3563) );
  NOR2_X2 U42944 ( .A1(n3596), .A2(n5481), .ZN(n6341) );
  NAND3_X2 U42945 ( .A1(n21137), .A2(n21136), .A3(n21139), .ZN(n22108) );
  NAND3_X1 U42949 ( .A1(n33609), .A2(n4263), .A3(n16851), .ZN(n21649) );
  AOI22_X2 U42952 ( .A1(n64397), .A2(n29462), .B1(n29463), .B2(n63315), .ZN(
        n29464) );
  NOR2_X2 U42953 ( .A1(n14647), .A2(n29459), .ZN(n64397) );
  NAND2_X2 U42966 ( .A1(n14964), .A2(n19190), .ZN(n33141) );
  NAND2_X2 U42967 ( .A1(n57467), .A2(n12829), .ZN(n50041) );
  AND2_X2 U42970 ( .A1(n48617), .A2(n48628), .Z(n57467) );
  INV_X2 U42973 ( .I(n43956), .ZN(n1687) );
  NAND2_X2 U42974 ( .A1(n18724), .A2(n43947), .ZN(n43956) );
  NAND2_X2 U42975 ( .A1(n64399), .A2(n58068), .ZN(n50399) );
  XOR2_X1 U42978 ( .A1(n23790), .A2(n23583), .Z(n38976) );
  NAND2_X1 U42984 ( .A1(n43145), .A2(n7490), .ZN(n58288) );
  NOR2_X2 U42988 ( .A1(n41697), .A2(n12195), .ZN(n46122) );
  BUF_X2 U43011 ( .I(n43365), .Z(n64400) );
  XOR2_X1 U43013 ( .A1(n46381), .A2(n64401), .Z(n9437) );
  XOR2_X1 U43015 ( .A1(n5169), .A2(n5170), .Z(n64401) );
  XOR2_X1 U43017 ( .A1(n52157), .A2(n18103), .Z(n50615) );
  XOR2_X1 U43022 ( .A1(n5180), .A2(n64403), .Z(n58289) );
  XOR2_X1 U43023 ( .A1(n3214), .A2(n92), .Z(n24964) );
  INV_X2 U43031 ( .I(n64404), .ZN(n57397) );
  NAND2_X2 U43032 ( .A1(n50123), .A2(n25233), .ZN(n64404) );
  BUF_X2 U43034 ( .I(n32984), .Z(n64405) );
  NOR2_X2 U43037 ( .A1(n57202), .A2(n23756), .ZN(n51878) );
  INV_X4 U43040 ( .I(n64408), .ZN(n56182) );
  NAND2_X1 U43049 ( .A1(n56791), .A2(n23030), .ZN(n56787) );
  NOR3_X2 U43054 ( .A1(n14628), .A2(n14627), .A3(n42983), .ZN(n13801) );
  XOR2_X1 U43055 ( .A1(n7753), .A2(n7752), .Z(n64541) );
  NAND3_X1 U43067 ( .A1(n48556), .A2(n22874), .A3(n48554), .ZN(n15395) );
  NOR2_X1 U43073 ( .A1(n41690), .A2(n42399), .ZN(n64411) );
  XOR2_X1 U43074 ( .A1(n39248), .A2(n65241), .Z(n64412) );
  NOR2_X2 U43076 ( .A1(n7092), .A2(n36853), .ZN(n36850) );
  AOI21_X2 U43077 ( .A1(n42453), .A2(n42452), .B(n10593), .ZN(n41809) );
  NAND2_X2 U43081 ( .A1(n6606), .A2(n35962), .ZN(n35357) );
  XOR2_X1 U43084 ( .A1(n13664), .A2(n64413), .Z(n8078) );
  XOR2_X1 U43101 ( .A1(n64640), .A2(n12356), .Z(n64413) );
  NAND3_X2 U43114 ( .A1(n39944), .A2(n39943), .A3(n39942), .ZN(n4111) );
  NOR2_X2 U43117 ( .A1(n49195), .A2(n61673), .ZN(n60666) );
  NAND4_X2 U43125 ( .A1(n3347), .A2(n50043), .A3(n50044), .A4(n3335), .ZN(
        n64414) );
  NOR2_X1 U43151 ( .A1(n29338), .A2(n58977), .ZN(n29342) );
  NOR2_X2 U43154 ( .A1(n26691), .A2(n27499), .ZN(n58977) );
  INV_X2 U43164 ( .I(n64415), .ZN(n17365) );
  XOR2_X1 U43165 ( .A1(n12880), .A2(n36638), .Z(n64415) );
  NAND2_X2 U43168 ( .A1(n23709), .A2(n57886), .ZN(n16473) );
  NOR2_X1 U43176 ( .A1(n10401), .A2(n33993), .ZN(n33994) );
  BUF_X2 U43180 ( .I(n18339), .Z(n64417) );
  XOR2_X1 U43192 ( .A1(n64419), .A2(n64418), .Z(n849) );
  OAI21_X2 U43194 ( .A1(n43150), .A2(n15214), .B(n23434), .ZN(n43148) );
  XOR2_X1 U43195 ( .A1(n64420), .A2(n400), .Z(n7009) );
  AOI22_X1 U43207 ( .A1(n9600), .A2(n42559), .B1(n42558), .B2(n42910), .ZN(
        n9599) );
  XOR2_X1 U43209 ( .A1(n64422), .A2(n64421), .Z(n20513) );
  XOR2_X1 U43212 ( .A1(n45249), .A2(n44587), .Z(n64421) );
  OR2_X1 U43213 ( .A1(n31355), .A2(n61799), .Z(n21179) );
  INV_X1 U43214 ( .I(n64423), .ZN(n14728) );
  NOR2_X2 U43218 ( .A1(n13297), .A2(n35883), .ZN(n64423) );
  NAND2_X1 U43225 ( .A1(n64426), .A2(n64425), .ZN(n58518) );
  NAND2_X1 U43228 ( .A1(n20855), .A2(n36572), .ZN(n64426) );
  NAND2_X2 U43237 ( .A1(n17829), .A2(n17827), .ZN(n35898) );
  XOR2_X1 U43245 ( .A1(n36323), .A2(n37147), .Z(n64427) );
  NOR2_X2 U43288 ( .A1(n41614), .A2(n17223), .ZN(n64961) );
  NAND2_X2 U43295 ( .A1(n40246), .A2(n40247), .ZN(n41614) );
  AND2_X1 U43303 ( .A1(n35062), .A2(n2460), .Z(n64429) );
  XOR2_X1 U43312 ( .A1(n64432), .A2(n64431), .Z(n4775) );
  XOR2_X1 U43316 ( .A1(n31234), .A2(n31233), .Z(n64432) );
  NAND3_X2 U43336 ( .A1(n61455), .A2(n39838), .A3(n39839), .ZN(n39841) );
  NAND3_X2 U43344 ( .A1(n10578), .A2(n5130), .A3(n34506), .ZN(n58748) );
  BUF_X4 U43355 ( .I(n51703), .Z(n54597) );
  NAND2_X1 U43356 ( .A1(n53147), .A2(n53161), .ZN(n2041) );
  INV_X2 U43364 ( .I(n7302), .ZN(n3029) );
  NAND2_X2 U43366 ( .A1(n18586), .A2(n58944), .ZN(n7302) );
  AOI22_X1 U43373 ( .A1(n36391), .A2(n64434), .B1(n7103), .B2(n36393), .ZN(
        n36398) );
  INV_X1 U43388 ( .I(n36548), .ZN(n64434) );
  NAND2_X2 U43396 ( .A1(n36385), .A2(n36538), .ZN(n36548) );
  INV_X2 U43405 ( .I(n64435), .ZN(n18088) );
  NOR2_X2 U43410 ( .A1(n10737), .A2(n18339), .ZN(n64435) );
  NOR2_X1 U43413 ( .A1(n54280), .A2(n54281), .ZN(n59914) );
  XOR2_X1 U43417 ( .A1(n64436), .A2(n50559), .Z(n2230) );
  XOR2_X1 U43429 ( .A1(n50452), .A2(n19228), .Z(n64436) );
  NOR2_X2 U43435 ( .A1(n15294), .A2(n33312), .ZN(n24249) );
  XOR2_X1 U43458 ( .A1(n64437), .A2(n51068), .Z(n26071) );
  XOR2_X1 U43473 ( .A1(n11166), .A2(n10217), .Z(n64437) );
  XOR2_X1 U43483 ( .A1(n52114), .A2(n51701), .Z(n58131) );
  XOR2_X1 U43498 ( .A1(n63033), .A2(n1196), .Z(n51701) );
  BUF_X2 U43520 ( .I(n56167), .Z(n64438) );
  NOR2_X2 U43539 ( .A1(n64439), .A2(n6164), .ZN(n64714) );
  BUF_X2 U43542 ( .I(n3656), .Z(n64443) );
  NAND2_X2 U43555 ( .A1(n37107), .A2(n37106), .ZN(n6159) );
  OAI21_X2 U43556 ( .A1(n16958), .A2(n16959), .B(n64444), .ZN(n21369) );
  NAND2_X2 U43558 ( .A1(n43601), .A2(n25368), .ZN(n12972) );
  NOR4_X2 U43559 ( .A1(n41371), .A2(n41370), .A3(n41372), .A4(n42148), .ZN(
        n64446) );
  NAND2_X1 U43576 ( .A1(n19209), .A2(n3611), .ZN(n58339) );
  AOI21_X2 U43577 ( .A1(n48173), .A2(n21466), .B(n21465), .ZN(n52623) );
  OAI21_X2 U43583 ( .A1(n23224), .A2(n29453), .B(n7979), .ZN(n28101) );
  NOR2_X2 U43589 ( .A1(n4288), .A2(n12742), .ZN(n12835) );
  NOR2_X1 U43605 ( .A1(n5082), .A2(n59553), .ZN(n6620) );
  INV_X2 U43608 ( .I(n25888), .ZN(n52429) );
  XOR2_X1 U43619 ( .A1(n25888), .A2(n61754), .Z(n50030) );
  NOR2_X2 U43625 ( .A1(n13973), .A2(n13972), .ZN(n25888) );
  XOR2_X1 U43627 ( .A1(n38542), .A2(n38731), .Z(n64448) );
  OAI22_X1 U43638 ( .A1(n6508), .A2(n40958), .B1(n40957), .B2(n40956), .ZN(
        n40960) );
  XOR2_X1 U43643 ( .A1(n64449), .A2(n33868), .Z(n12243) );
  XOR2_X1 U43654 ( .A1(n33873), .A2(n45295), .Z(n64449) );
  BUF_X2 U43660 ( .I(n1407), .Z(n64450) );
  OR2_X1 U43665 ( .A1(n12378), .A2(n42594), .Z(n5044) );
  NOR4_X2 U43671 ( .A1(n23832), .A2(n23831), .A3(n56930), .A4(n56931), .ZN(
        n60870) );
  NAND2_X2 U43672 ( .A1(n40971), .A2(n23787), .ZN(n20374) );
  XOR2_X1 U43680 ( .A1(n64452), .A2(n7639), .Z(n5271) );
  XOR2_X1 U43691 ( .A1(n38630), .A2(n24752), .Z(n64452) );
  NAND2_X2 U43697 ( .A1(n19255), .A2(n25349), .ZN(n29332) );
  NAND2_X2 U43700 ( .A1(n31146), .A2(n14764), .ZN(n29480) );
  OR2_X1 U43705 ( .A1(n847), .A2(n13976), .Z(n31138) );
  XOR2_X1 U43709 ( .A1(n38731), .A2(n39449), .Z(n60714) );
  XOR2_X1 U43712 ( .A1(n38786), .A2(n15308), .Z(n39449) );
  NAND2_X2 U43726 ( .A1(n60901), .A2(n13090), .ZN(n5971) );
  NAND3_X2 U43734 ( .A1(n51864), .A2(n54346), .A3(n6737), .ZN(n54353) );
  XOR2_X1 U43740 ( .A1(n39750), .A2(n64455), .Z(n24035) );
  XOR2_X1 U43743 ( .A1(n39747), .A2(n39746), .Z(n64455) );
  NOR2_X2 U43744 ( .A1(n47186), .A2(n17452), .ZN(n48108) );
  INV_X2 U43745 ( .I(n29461), .ZN(n28117) );
  NAND2_X2 U43758 ( .A1(n29455), .A2(n29456), .ZN(n29461) );
  NAND2_X2 U43760 ( .A1(n5215), .A2(n64456), .ZN(n22486) );
  OAI21_X1 U43764 ( .A1(n59030), .A2(n61698), .B(n62760), .ZN(n64456) );
  OR2_X1 U43782 ( .A1(n16993), .A2(n10863), .Z(n47020) );
  INV_X2 U43801 ( .I(n9082), .ZN(n6635) );
  OAI21_X2 U43803 ( .A1(n48342), .A2(n64457), .B(n48341), .ZN(n61115) );
  NOR2_X2 U43810 ( .A1(n48337), .A2(n63546), .ZN(n64457) );
  XOR2_X1 U43811 ( .A1(n17300), .A2(n25594), .Z(n23089) );
  NOR2_X2 U43816 ( .A1(n5838), .A2(n5839), .ZN(n17300) );
  XOR2_X1 U43823 ( .A1(n9854), .A2(n64460), .Z(n6649) );
  XOR2_X1 U43827 ( .A1(n14316), .A2(n22338), .Z(n64460) );
  XOR2_X1 U43829 ( .A1(n64490), .A2(n59000), .Z(n25134) );
  BUF_X2 U43839 ( .I(n25251), .Z(n64461) );
  NAND2_X1 U43846 ( .A1(n43182), .A2(n22705), .ZN(n20498) );
  NOR2_X2 U43859 ( .A1(n50427), .A2(n50426), .ZN(n50425) );
  AOI21_X1 U43862 ( .A1(n16694), .A2(n1434), .B(n9186), .ZN(n30544) );
  AND2_X1 U43865 ( .A1(n18473), .A2(n42477), .Z(n15921) );
  NOR2_X2 U43877 ( .A1(n14477), .A2(n64463), .ZN(n14498) );
  OR3_X1 U43881 ( .A1(n18137), .A2(n25664), .A3(n60503), .Z(n64463) );
  NOR2_X2 U43885 ( .A1(n57868), .A2(n26687), .ZN(n9543) );
  NAND3_X2 U43886 ( .A1(n53119), .A2(n23243), .A3(n53078), .ZN(n53104) );
  NOR2_X2 U43899 ( .A1(n19080), .A2(n53077), .ZN(n53119) );
  XOR2_X1 U43903 ( .A1(n3182), .A2(n64471), .Z(n15785) );
  XOR2_X1 U43905 ( .A1(n18562), .A2(n19691), .Z(n64471) );
  INV_X1 U43925 ( .I(n12755), .ZN(n5068) );
  OAI21_X2 U43927 ( .A1(n64473), .A2(n64472), .B(n35837), .ZN(n34397) );
  NOR2_X2 U43930 ( .A1(n61764), .A2(n64474), .ZN(n59547) );
  OAI21_X2 U43933 ( .A1(n58881), .A2(n64231), .B(n47102), .ZN(n64474) );
  BUF_X2 U43934 ( .I(n23484), .Z(n64475) );
  NAND2_X1 U43942 ( .A1(n17562), .A2(n5019), .ZN(n64674) );
  NAND2_X2 U43967 ( .A1(n61203), .A2(n46568), .ZN(n50406) );
  NOR3_X2 U43979 ( .A1(n87), .A2(n47848), .A3(n61680), .ZN(n47850) );
  XOR2_X1 U43989 ( .A1(n31686), .A2(n32754), .Z(n31407) );
  NAND2_X2 U43996 ( .A1(n12984), .A2(n3961), .ZN(n32754) );
  NAND2_X2 U44056 ( .A1(n30491), .A2(n18917), .ZN(n30494) );
  XOR2_X1 U44067 ( .A1(n60003), .A2(n15351), .Z(n64480) );
  NOR2_X2 U44087 ( .A1(n3362), .A2(n60774), .ZN(n10971) );
  NAND3_X2 U44124 ( .A1(n11531), .A2(n11532), .A3(n11530), .ZN(n23341) );
  INV_X2 U44181 ( .I(n28375), .ZN(n64481) );
  BUF_X2 U44193 ( .I(n10734), .Z(n64484) );
  NAND3_X1 U44194 ( .A1(n53436), .A2(n53209), .A3(n60475), .ZN(n64489) );
  XOR2_X1 U44200 ( .A1(n43998), .A2(n17762), .Z(n2680) );
  XOR2_X1 U44222 ( .A1(n61347), .A2(n44980), .Z(n17762) );
  XOR2_X1 U44225 ( .A1(n51230), .A2(n25315), .Z(n64490) );
  NOR2_X2 U44230 ( .A1(n54506), .A2(n54505), .ZN(n58896) );
  NAND2_X2 U44234 ( .A1(n32458), .A2(n33614), .ZN(n7838) );
  NAND2_X1 U44240 ( .A1(n11759), .A2(n27430), .ZN(n64494) );
  NAND2_X2 U44243 ( .A1(n6926), .A2(n43268), .ZN(n64495) );
  AND2_X1 U44267 ( .A1(n47077), .A2(n47078), .Z(n65261) );
  XOR2_X1 U44275 ( .A1(n21918), .A2(n21289), .Z(n59551) );
  XOR2_X1 U44325 ( .A1(n37818), .A2(n39223), .Z(n21918) );
  NAND2_X2 U44329 ( .A1(n30731), .A2(n30285), .ZN(n8685) );
  NOR2_X2 U44335 ( .A1(n30265), .A2(n61734), .ZN(n30731) );
  INV_X4 U44429 ( .I(n34078), .ZN(n1417) );
  XOR2_X1 U44442 ( .A1(n46546), .A2(n25926), .Z(n14639) );
  XOR2_X1 U44469 ( .A1(n13180), .A2(n20347), .Z(n25926) );
  NAND2_X2 U44471 ( .A1(n11160), .A2(n15720), .ZN(n3149) );
  OAI21_X2 U44479 ( .A1(n50576), .A2(n52323), .B(n64497), .ZN(n18091) );
  NAND2_X2 U44485 ( .A1(n50576), .A2(n20593), .ZN(n64497) );
  AOI21_X1 U44497 ( .A1(n29869), .A2(n20439), .B(n64498), .ZN(n29873) );
  INV_X2 U44512 ( .I(n23125), .ZN(n64499) );
  XOR2_X1 U44514 ( .A1(n46253), .A2(n22973), .Z(n11252) );
  XOR2_X1 U44591 ( .A1(n44940), .A2(n46553), .Z(n44941) );
  XOR2_X1 U44593 ( .A1(n65170), .A2(n51019), .Z(n44940) );
  XOR2_X1 U44605 ( .A1(n64500), .A2(n31946), .Z(n33810) );
  XOR2_X1 U44622 ( .A1(n31938), .A2(n33079), .Z(n64500) );
  NAND2_X1 U44646 ( .A1(n12798), .A2(n37455), .ZN(n36967) );
  NAND2_X2 U44657 ( .A1(n24459), .A2(n25308), .ZN(n12798) );
  XOR2_X1 U44692 ( .A1(n22478), .A2(n11318), .Z(n50906) );
  XOR2_X1 U44698 ( .A1(n64501), .A2(n17731), .Z(n58272) );
  NAND2_X2 U44708 ( .A1(n24052), .A2(n29613), .ZN(n29616) );
  NAND2_X1 U44709 ( .A1(n64582), .A2(n60278), .ZN(n9631) );
  XOR2_X1 U44748 ( .A1(n64505), .A2(n39715), .Z(n58489) );
  XOR2_X1 U44769 ( .A1(n39716), .A2(n24058), .Z(n64505) );
  NAND2_X2 U44775 ( .A1(n24871), .A2(n24872), .ZN(n15927) );
  XOR2_X1 U44816 ( .A1(n61117), .A2(n12812), .Z(n24872) );
  INV_X2 U44817 ( .I(n64506), .ZN(n27262) );
  NAND3_X2 U44820 ( .A1(n27980), .A2(n64506), .A3(n8528), .ZN(n29158) );
  XOR2_X1 U44833 ( .A1(n3431), .A2(n1213), .Z(n14218) );
  NAND2_X2 U44853 ( .A1(n21290), .A2(n64508), .ZN(n24429) );
  NAND2_X2 U44854 ( .A1(n57247), .A2(n64509), .ZN(n23603) );
  NOR3_X2 U44856 ( .A1(n2987), .A2(n64662), .A3(n57254), .ZN(n64509) );
  XOR2_X1 U44865 ( .A1(n23669), .A2(n33292), .Z(n32069) );
  XOR2_X1 U44868 ( .A1(n8165), .A2(n24018), .Z(n38755) );
  OAI22_X2 U44872 ( .A1(n29768), .A2(n7025), .B1(n26841), .B2(n30126), .ZN(
        n30122) );
  XOR2_X1 U44890 ( .A1(n51945), .A2(n51229), .Z(n50994) );
  OR2_X1 U44927 ( .A1(n3213), .A2(n3436), .Z(n13525) );
  XOR2_X1 U44944 ( .A1(n59678), .A2(n32196), .Z(n64511) );
  XOR2_X1 U44971 ( .A1(n7882), .A2(n7879), .Z(n13836) );
  XOR2_X1 U44988 ( .A1(n64514), .A2(n64513), .Z(n13312) );
  XOR2_X1 U44993 ( .A1(n51990), .A2(n58500), .Z(n64514) );
  XOR2_X1 U44996 ( .A1(n11372), .A2(n64515), .Z(n47653) );
  XOR2_X1 U45015 ( .A1(n44268), .A2(n57785), .Z(n64515) );
  XOR2_X1 U45018 ( .A1(n64516), .A2(n10536), .Z(n41772) );
  XOR2_X1 U45021 ( .A1(n13883), .A2(n41754), .Z(n64516) );
  NOR2_X2 U45037 ( .A1(n64517), .A2(n13075), .ZN(n12905) );
  NAND2_X2 U45040 ( .A1(n5243), .A2(n2572), .ZN(n5242) );
  NAND3_X2 U45043 ( .A1(n26554), .A2(n26556), .A3(n26555), .ZN(n5243) );
  NOR2_X1 U45067 ( .A1(n14904), .A2(n21010), .ZN(n37038) );
  OR2_X1 U45068 ( .A1(n13247), .A2(n35491), .Z(n34866) );
  INV_X2 U45069 ( .I(n10391), .ZN(n59895) );
  NAND2_X2 U45073 ( .A1(n8494), .A2(n22836), .ZN(n10391) );
  XOR2_X1 U45074 ( .A1(n16994), .A2(n10860), .Z(n16993) );
  XOR2_X1 U45075 ( .A1(n38972), .A2(n466), .Z(n39721) );
  INV_X2 U45079 ( .I(n64518), .ZN(n12702) );
  XNOR2_X1 U45115 ( .A1(n57356), .A2(n12703), .ZN(n64518) );
  NOR3_X2 U45126 ( .A1(n18682), .A2(n57388), .A3(n64519), .ZN(n60447) );
  NAND2_X2 U45134 ( .A1(n10930), .A2(n34197), .ZN(n64519) );
  NAND2_X1 U45181 ( .A1(n18915), .A2(n18916), .ZN(n18914) );
  NAND2_X2 U45198 ( .A1(n56411), .A2(n14600), .ZN(n20239) );
  XOR2_X1 U45201 ( .A1(n64523), .A2(n51145), .Z(n51147) );
  NOR3_X2 U45213 ( .A1(n64525), .A2(n35473), .A3(n64524), .ZN(n35478) );
  XOR2_X1 U45225 ( .A1(n15525), .A2(n7145), .Z(n15524) );
  NOR2_X2 U45240 ( .A1(n49673), .A2(n48711), .ZN(n65061) );
  NAND2_X2 U45245 ( .A1(n61223), .A2(n36245), .ZN(n35602) );
  NAND2_X1 U45259 ( .A1(n57744), .A2(n21030), .ZN(n64527) );
  XOR2_X1 U45266 ( .A1(n18191), .A2(n18103), .Z(n6364) );
  NAND2_X2 U45267 ( .A1(n6368), .A2(n6367), .ZN(n18103) );
  XOR2_X1 U45269 ( .A1(n64528), .A2(n38221), .Z(n11644) );
  XOR2_X1 U45278 ( .A1(n3531), .A2(n3529), .Z(n64528) );
  XOR2_X1 U45285 ( .A1(n14299), .A2(n58819), .Z(n11768) );
  NAND2_X2 U45286 ( .A1(n9208), .A2(n9207), .ZN(n14299) );
  NOR2_X2 U45288 ( .A1(n48014), .A2(n64529), .ZN(n48015) );
  NAND3_X1 U45304 ( .A1(n54451), .A2(n55016), .A3(n55022), .ZN(n52640) );
  AND2_X1 U45306 ( .A1(n47607), .A2(n47818), .Z(n64870) );
  NOR2_X2 U45350 ( .A1(n6640), .A2(n10111), .ZN(n64531) );
  NAND2_X1 U45368 ( .A1(n21249), .A2(n15974), .ZN(n54646) );
  XOR2_X1 U45369 ( .A1(n37867), .A2(n38072), .Z(n3397) );
  OAI21_X1 U45382 ( .A1(n22045), .A2(n42252), .B(n60612), .ZN(n58104) );
  NAND2_X2 U45387 ( .A1(n24991), .A2(n3403), .ZN(n60612) );
  BUF_X2 U45398 ( .I(n42127), .Z(n64532) );
  NAND2_X2 U45401 ( .A1(n60364), .A2(n60546), .ZN(n36853) );
  OAI22_X2 U45439 ( .A1(n9119), .A2(n24138), .B1(n45386), .B2(n23415), .ZN(
        n44269) );
  INV_X1 U45468 ( .I(n64810), .ZN(n29359) );
  NAND2_X1 U45469 ( .A1(n21268), .A2(n22947), .ZN(n52943) );
  AND2_X1 U45470 ( .A1(n47646), .A2(n49676), .Z(n49685) );
  OR2_X1 U45481 ( .A1(n43478), .A2(n62686), .Z(n18650) );
  BUF_X2 U45503 ( .I(n22128), .Z(n64534) );
  XOR2_X1 U45506 ( .A1(n31993), .A2(n33269), .Z(n2906) );
  XOR2_X1 U45521 ( .A1(n18516), .A2(n19228), .Z(n60086) );
  XOR2_X1 U45530 ( .A1(n10502), .A2(n23991), .Z(n18516) );
  XOR2_X1 U45531 ( .A1(n64541), .A2(n19753), .Z(n7750) );
  NAND2_X2 U45542 ( .A1(n2951), .A2(n1459), .ZN(n2997) );
  NAND2_X2 U45658 ( .A1(n47901), .A2(n44802), .ZN(n2571) );
  XOR2_X1 U45661 ( .A1(n5363), .A2(n22697), .Z(n38319) );
  XOR2_X1 U45662 ( .A1(n20202), .A2(n64542), .Z(n22060) );
  XOR2_X1 U45663 ( .A1(n22062), .A2(n38320), .Z(n64542) );
  AOI21_X2 U45671 ( .A1(n55961), .A2(n64719), .B(n64543), .ZN(n55962) );
  NAND2_X1 U45695 ( .A1(n46735), .A2(n64544), .ZN(n61389) );
  AND2_X2 U45700 ( .A1(n20953), .A2(n20739), .Z(n9203) );
  NAND2_X2 U45701 ( .A1(n29819), .A2(n7774), .ZN(n28698) );
  NAND2_X2 U45736 ( .A1(n64549), .A2(n64548), .ZN(n20514) );
  INV_X2 U45752 ( .I(n47884), .ZN(n64549) );
  NAND2_X2 U45754 ( .A1(n23976), .A2(n23977), .ZN(n57758) );
  NOR2_X2 U45755 ( .A1(n3432), .A2(n34349), .ZN(n33751) );
  NAND2_X2 U45759 ( .A1(n1408), .A2(n13811), .ZN(n25511) );
  XOR2_X1 U45767 ( .A1(n21546), .A2(n10786), .Z(n4031) );
  NAND2_X2 U45769 ( .A1(n53692), .A2(n53676), .ZN(n25859) );
  XOR2_X1 U45771 ( .A1(n37972), .A2(n64551), .Z(n25142) );
  XOR2_X1 U45775 ( .A1(n37978), .A2(n61791), .Z(n64551) );
  XOR2_X1 U45784 ( .A1(n15292), .A2(n15290), .Z(n15289) );
  NAND4_X2 U45788 ( .A1(n42650), .A2(n22282), .A3(n64400), .A4(n14920), .ZN(
        n11224) );
  NAND2_X2 U45803 ( .A1(n22736), .A2(n23347), .ZN(n47370) );
  OAI21_X2 U45818 ( .A1(n50520), .A2(n50522), .B(n50521), .ZN(n9386) );
  NAND2_X2 U45824 ( .A1(n9387), .A2(n22268), .ZN(n50520) );
  NAND3_X1 U45830 ( .A1(n36561), .A2(n36563), .A3(n36553), .ZN(n35537) );
  NAND2_X1 U45842 ( .A1(n65044), .A2(n49595), .ZN(n49604) );
  NAND2_X1 U45843 ( .A1(n53697), .A2(n53688), .ZN(n2838) );
  XOR2_X1 U45845 ( .A1(n4900), .A2(n58617), .Z(n64552) );
  XOR2_X1 U45853 ( .A1(n52156), .A2(n64553), .Z(n5502) );
  XOR2_X1 U45854 ( .A1(n52166), .A2(n6512), .Z(n64553) );
  INV_X2 U45885 ( .I(n64554), .ZN(n15789) );
  XOR2_X1 U45886 ( .A1(Ciphertext[28]), .A2(Key[185]), .Z(n64554) );
  NOR2_X2 U45888 ( .A1(n17156), .A2(n61646), .ZN(n59398) );
  NAND2_X2 U45909 ( .A1(n64974), .A2(n22117), .ZN(n3862) );
  NAND2_X2 U45913 ( .A1(n46982), .A2(n44680), .ZN(n14875) );
  XOR2_X1 U45914 ( .A1(n64555), .A2(n23093), .Z(Plaintext[69]) );
  NAND3_X1 U45918 ( .A1(n5112), .A2(n6556), .A3(n6562), .ZN(n64555) );
  NAND2_X1 U45941 ( .A1(n16780), .A2(n53327), .ZN(n16779) );
  NOR2_X2 U45943 ( .A1(n40471), .A2(n25118), .ZN(n14004) );
  NAND2_X2 U45957 ( .A1(n39158), .A2(n6276), .ZN(n40471) );
  NAND3_X1 U46092 ( .A1(n27387), .A2(n28239), .A3(n27380), .ZN(n26266) );
  INV_X1 U46108 ( .I(n29578), .ZN(n30300) );
  NAND2_X1 U46214 ( .A1(n29576), .A2(n29269), .ZN(n29578) );
  NAND4_X2 U46217 ( .A1(n44074), .A2(n44071), .A3(n44072), .A4(n44073), .ZN(
        n44075) );
  XOR2_X1 U46220 ( .A1(n2153), .A2(n10594), .Z(n64556) );
  INV_X1 U46224 ( .I(n30398), .ZN(n64694) );
  XOR2_X1 U46225 ( .A1(n61518), .A2(n52453), .Z(n51180) );
  NAND3_X2 U46242 ( .A1(n47056), .A2(n47057), .A3(n49004), .ZN(n61518) );
  AOI21_X2 U46270 ( .A1(n12205), .A2(n47827), .B(n64557), .ZN(n12199) );
  NOR2_X2 U46286 ( .A1(n59198), .A2(n64558), .ZN(n59311) );
  NAND2_X1 U46293 ( .A1(n65048), .A2(n17948), .ZN(n64558) );
  NAND2_X2 U46294 ( .A1(n5563), .A2(n64559), .ZN(n17758) );
  OAI21_X2 U46349 ( .A1(n29095), .A2(n29094), .B(n63891), .ZN(n64559) );
  OAI21_X2 U46359 ( .A1(n55570), .A2(n55569), .B(n55556), .ZN(n55521) );
  NAND2_X2 U46360 ( .A1(n55550), .A2(n21272), .ZN(n55570) );
  XOR2_X1 U46364 ( .A1(n64560), .A2(n50817), .Z(Plaintext[7]) );
  OR2_X1 U46377 ( .A1(n49528), .A2(n64561), .Z(n48778) );
  NAND2_X1 U46411 ( .A1(n16542), .A2(n50355), .ZN(n64563) );
  XOR2_X1 U46433 ( .A1(n52084), .A2(n52085), .Z(n52087) );
  NAND3_X1 U46455 ( .A1(n1177), .A2(n53141), .A3(n53142), .ZN(n65107) );
  NAND2_X2 U46484 ( .A1(n19992), .A2(n17063), .ZN(n64709) );
  INV_X2 U46523 ( .I(n26650), .ZN(n64565) );
  NAND3_X1 U46534 ( .A1(n31145), .A2(n1316), .A3(n30374), .ZN(n29012) );
  BUF_X2 U46550 ( .I(n19990), .Z(n64566) );
  XOR2_X1 U46568 ( .A1(n6384), .A2(n6336), .Z(n64567) );
  XOR2_X1 U46628 ( .A1(n58573), .A2(n44922), .Z(n12373) );
  INV_X2 U46635 ( .I(n1929), .ZN(n58573) );
  NOR2_X2 U46642 ( .A1(n21364), .A2(n23897), .ZN(n54599) );
  NAND3_X2 U46689 ( .A1(n7856), .A2(n7855), .A3(n36609), .ZN(n39343) );
  XOR2_X1 U46692 ( .A1(n23678), .A2(n51503), .Z(n25798) );
  XOR2_X1 U46693 ( .A1(n52604), .A2(n52107), .Z(n51503) );
  XNOR2_X1 U46696 ( .A1(n24254), .A2(n31763), .ZN(n65055) );
  OAI21_X2 U46706 ( .A1(n28437), .A2(n28438), .B(n28436), .ZN(n64572) );
  INV_X1 U46753 ( .I(n15697), .ZN(n64573) );
  OAI21_X2 U46766 ( .A1(n63144), .A2(n46053), .B(n22389), .ZN(n46058) );
  XOR2_X1 U46776 ( .A1(n4294), .A2(n25076), .Z(n7388) );
  NAND2_X2 U46841 ( .A1(n4295), .A2(n4301), .ZN(n4294) );
  XOR2_X1 U46872 ( .A1(n6274), .A2(n58969), .Z(n58968) );
  XOR2_X1 U46873 ( .A1(n59597), .A2(n61263), .Z(n64574) );
  XOR2_X1 U46874 ( .A1(n5154), .A2(n21952), .Z(n31480) );
  INV_X2 U46919 ( .I(n64575), .ZN(n25467) );
  XOR2_X1 U46921 ( .A1(n25713), .A2(n8983), .Z(n37554) );
  NAND3_X1 U46933 ( .A1(n22700), .A2(n47728), .A3(n47736), .ZN(n64576) );
  NOR3_X2 U47095 ( .A1(n64577), .A2(n34738), .A3(n22297), .ZN(n24581) );
  NOR2_X1 U47098 ( .A1(n18510), .A2(n47015), .ZN(n6060) );
  OAI22_X1 U47130 ( .A1(n42245), .A2(n4635), .B1(n60612), .B2(n42240), .ZN(
        n42243) );
  OAI21_X2 U47160 ( .A1(n5963), .A2(n5964), .B(n64578), .ZN(n5968) );
  NAND2_X1 U47167 ( .A1(n1161), .A2(n1581), .ZN(n64578) );
  OAI21_X2 U47246 ( .A1(n5368), .A2(n42355), .B(n20922), .ZN(n41613) );
  NAND3_X2 U47256 ( .A1(n64699), .A2(n6474), .A3(n60803), .ZN(n32541) );
  NOR2_X1 U47257 ( .A1(n41480), .A2(n40753), .ZN(n64580) );
  NAND2_X2 U47323 ( .A1(n12235), .A2(n60507), .ZN(n6138) );
  OR2_X1 U47349 ( .A1(n17414), .A2(n29516), .Z(n28743) );
  NAND4_X2 U47351 ( .A1(n52275), .A2(n52276), .A3(n58789), .A4(n52277), .ZN(
        n52278) );
  INV_X4 U47358 ( .I(n51209), .ZN(n23069) );
  NAND3_X2 U47365 ( .A1(n25039), .A2(n25041), .A3(n17707), .ZN(n51209) );
  NOR2_X2 U47409 ( .A1(n61076), .A2(n35830), .ZN(n35852) );
  INV_X4 U47469 ( .I(n14488), .ZN(n60467) );
  NAND3_X1 U47488 ( .A1(n21434), .A2(n3937), .A3(n57160), .ZN(n21433) );
  INV_X2 U47540 ( .I(n24815), .ZN(n1865) );
  NAND3_X2 U47547 ( .A1(n24813), .A2(n24812), .A3(n16150), .ZN(n24815) );
  NOR2_X1 U47563 ( .A1(n65063), .A2(n11698), .ZN(n64582) );
  INV_X2 U47571 ( .I(n2857), .ZN(n64684) );
  INV_X2 U47576 ( .I(n9504), .ZN(n42058) );
  NAND2_X2 U47589 ( .A1(n61237), .A2(n57886), .ZN(n9504) );
  AOI22_X1 U47592 ( .A1(n57134), .A2(n57107), .B1(n57106), .B2(n57433), .ZN(
        n19195) );
  AND2_X1 U47604 ( .A1(n28762), .A2(n1556), .Z(n755) );
  INV_X2 U47621 ( .I(n28948), .ZN(n13320) );
  XOR2_X1 U47675 ( .A1(n21498), .A2(n21497), .Z(n65045) );
  INV_X2 U47679 ( .I(n64585), .ZN(n57433) );
  XOR2_X1 U47683 ( .A1(n38913), .A2(n58177), .Z(n4816) );
  XOR2_X1 U47684 ( .A1(n37555), .A2(n58281), .Z(n58177) );
  NAND2_X1 U47685 ( .A1(n16801), .A2(n57029), .ZN(n64586) );
  NAND2_X1 U47686 ( .A1(n59724), .A2(n60970), .ZN(n32944) );
  NAND2_X2 U47694 ( .A1(n21878), .A2(n25372), .ZN(n60970) );
  NAND3_X1 U47742 ( .A1(n23110), .A2(n53241), .A3(n57390), .ZN(n52262) );
  AND2_X1 U47743 ( .A1(n52685), .A2(n8597), .Z(n16080) );
  NAND2_X2 U47749 ( .A1(n25261), .A2(n32984), .ZN(n36565) );
  OAI21_X1 U47761 ( .A1(n36093), .A2(n36092), .B(n36576), .ZN(n36094) );
  XOR2_X1 U47774 ( .A1(n6739), .A2(n51120), .Z(n64587) );
  NAND2_X2 U47804 ( .A1(n20160), .A2(n20159), .ZN(n38912) );
  NAND3_X2 U47818 ( .A1(n3710), .A2(n27399), .A3(n64701), .ZN(n65088) );
  NAND3_X2 U47820 ( .A1(n754), .A2(n12343), .A3(n37831), .ZN(n43693) );
  INV_X2 U47821 ( .I(n64591), .ZN(n1203) );
  NAND2_X2 U47824 ( .A1(n19891), .A2(n64711), .ZN(n11037) );
  XOR2_X1 U47832 ( .A1(n15661), .A2(n857), .Z(n64593) );
  XOR2_X1 U47841 ( .A1(n44886), .A2(n44510), .Z(n44550) );
  XOR2_X1 U47854 ( .A1(n9083), .A2(n16932), .Z(n44886) );
  NAND3_X2 U47855 ( .A1(n26630), .A2(n26631), .A3(n27554), .ZN(n64595) );
  NAND4_X2 U47861 ( .A1(n64597), .A2(n48616), .A3(n47169), .A4(n58675), .ZN(
        n47172) );
  NOR2_X2 U47874 ( .A1(n42739), .A2(n61121), .ZN(n42743) );
  NOR2_X2 U47879 ( .A1(n9760), .A2(n33648), .ZN(n33715) );
  INV_X2 U47890 ( .I(n23554), .ZN(n64598) );
  XOR2_X1 U47928 ( .A1(n6592), .A2(n31766), .Z(n57598) );
  NOR2_X2 U47935 ( .A1(n64674), .A2(n64599), .ZN(n3654) );
  NAND2_X2 U47942 ( .A1(n65252), .A2(n2631), .ZN(n2630) );
  XOR2_X1 U47946 ( .A1(n38123), .A2(n38745), .Z(n3438) );
  NOR2_X1 U47954 ( .A1(n40397), .A2(n40398), .ZN(n64924) );
  XOR2_X1 U47959 ( .A1(n6216), .A2(n51508), .Z(n51364) );
  XOR2_X1 U47974 ( .A1(n8002), .A2(n10409), .Z(n64600) );
  XOR2_X1 U47988 ( .A1(n37657), .A2(n64601), .Z(n11527) );
  XOR2_X1 U47994 ( .A1(n37561), .A2(n17321), .Z(n64601) );
  NAND3_X1 U47995 ( .A1(n53068), .A2(n53106), .A3(n22980), .ZN(n53075) );
  XOR2_X1 U48001 ( .A1(n60922), .A2(n10899), .Z(n60194) );
  OAI21_X1 U48005 ( .A1(n42396), .A2(n19809), .B(n1396), .ZN(n19808) );
  NAND2_X2 U48037 ( .A1(n64602), .A2(n59408), .ZN(n7402) );
  BUF_X2 U48040 ( .I(n23331), .Z(n64605) );
  INV_X1 U48067 ( .I(n32107), .ZN(n64607) );
  NOR2_X2 U48085 ( .A1(n30084), .A2(n61729), .ZN(n29798) );
  XOR2_X1 U48087 ( .A1(n64606), .A2(n38874), .Z(n60157) );
  XOR2_X1 U48090 ( .A1(n9803), .A2(n38870), .Z(n64606) );
  AOI22_X1 U48091 ( .A1(n61766), .A2(n64649), .B1(n56716), .B2(n23785), .ZN(
        n56648) );
  NOR2_X2 U48097 ( .A1(n20269), .A2(n56687), .ZN(n56716) );
  NAND4_X2 U48117 ( .A1(n47710), .A2(n47711), .A3(n19422), .A4(n47709), .ZN(
        n47712) );
  INV_X2 U48125 ( .I(n54501), .ZN(n22775) );
  NAND2_X2 U48133 ( .A1(n16797), .A2(n53845), .ZN(n54501) );
  NAND2_X1 U48135 ( .A1(n15716), .A2(n13858), .ZN(n55867) );
  NOR2_X2 U48143 ( .A1(n55469), .A2(n55471), .ZN(n55730) );
  XOR2_X1 U48158 ( .A1(n50861), .A2(n50862), .Z(n24480) );
  XOR2_X1 U48159 ( .A1(n62987), .A2(n52341), .Z(n50862) );
  XOR2_X1 U48169 ( .A1(n13410), .A2(n64611), .Z(n13409) );
  XOR2_X1 U48187 ( .A1(n39313), .A2(n64612), .Z(n64611) );
  BUF_X2 U48188 ( .I(n40295), .Z(n64613) );
  NOR2_X2 U48189 ( .A1(n48913), .A2(n48912), .ZN(n50436) );
  NAND2_X2 U48237 ( .A1(n64737), .A2(n58327), .ZN(n48913) );
  BUF_X2 U48241 ( .I(n25993), .Z(n64614) );
  OR2_X1 U48269 ( .A1(n37034), .A2(n22524), .Z(n59137) );
  NOR2_X2 U48270 ( .A1(n24473), .A2(n56436), .ZN(n24472) );
  NOR2_X2 U48279 ( .A1(n60121), .A2(n9629), .ZN(n10887) );
  NOR2_X2 U48286 ( .A1(n10495), .A2(n23220), .ZN(n32076) );
  XOR2_X1 U48307 ( .A1(n65077), .A2(n64615), .Z(n17891) );
  XOR2_X1 U48310 ( .A1(n45860), .A2(n11725), .Z(n64615) );
  NAND2_X2 U48318 ( .A1(n6121), .A2(n64616), .ZN(n2928) );
  INV_X2 U48326 ( .I(n14759), .ZN(n29455) );
  NAND2_X2 U48333 ( .A1(n28707), .A2(n21159), .ZN(n30364) );
  NAND2_X2 U48334 ( .A1(n3619), .A2(n42868), .ZN(n1908) );
  NAND2_X2 U48337 ( .A1(n59419), .A2(n59418), .ZN(n47260) );
  BUF_X2 U48343 ( .I(n2958), .Z(n64620) );
  NAND3_X2 U48354 ( .A1(n64621), .A2(n28247), .A3(n28246), .ZN(n15094) );
  OR2_X1 U48359 ( .A1(n28241), .A2(n28240), .Z(n64622) );
  XOR2_X1 U48361 ( .A1(n64623), .A2(n10904), .Z(n57832) );
  XOR2_X1 U48366 ( .A1(n33882), .A2(n33881), .Z(n64623) );
  OAI22_X1 U48371 ( .A1(n39420), .A2(n64624), .B1(n21701), .B2(n40242), .ZN(
        n21285) );
  NAND2_X1 U48378 ( .A1(n63952), .A2(n21701), .ZN(n64624) );
  XNOR2_X1 U48393 ( .A1(n15854), .A2(n30070), .ZN(n64632) );
  AOI21_X1 U48396 ( .A1(n36097), .A2(n36098), .B(n36574), .ZN(n36100) );
  NAND2_X2 U48403 ( .A1(n64625), .A2(n9105), .ZN(n55088) );
  XOR2_X1 U48404 ( .A1(n3621), .A2(n51003), .Z(n10406) );
  NOR2_X2 U48405 ( .A1(n16962), .A2(n25921), .ZN(n40052) );
  NOR2_X1 U48410 ( .A1(n64627), .A2(n3545), .ZN(n3544) );
  NAND2_X1 U48411 ( .A1(n59372), .A2(n59373), .ZN(n64627) );
  XOR2_X1 U48414 ( .A1(n64628), .A2(n11070), .Z(n65264) );
  XOR2_X1 U48438 ( .A1(n18452), .A2(n306), .Z(n795) );
  BUF_X2 U48440 ( .I(n41540), .Z(n64629) );
  OR2_X2 U48444 ( .A1(n11413), .A2(n3233), .Z(n17851) );
  XOR2_X1 U48445 ( .A1(n24508), .A2(n2686), .Z(n17618) );
  XOR2_X1 U48461 ( .A1(n64630), .A2(n59417), .Z(n6873) );
  XOR2_X1 U48463 ( .A1(n18308), .A2(n64796), .Z(n64630) );
  NOR2_X2 U48468 ( .A1(n64631), .A2(n61741), .ZN(n65276) );
  NAND3_X2 U48492 ( .A1(n23061), .A2(n18766), .A3(n61756), .ZN(n47813) );
  NAND2_X2 U48493 ( .A1(n10077), .A2(n25495), .ZN(n8673) );
  NOR2_X2 U48509 ( .A1(n32846), .A2(n3272), .ZN(n24287) );
  INV_X2 U48513 ( .I(n17203), .ZN(n34993) );
  XOR2_X1 U48514 ( .A1(n24796), .A2(n64632), .Z(n17203) );
  XOR2_X1 U48537 ( .A1(n8237), .A2(n11922), .Z(n2622) );
  BUF_X2 U48539 ( .I(n60232), .Z(n64634) );
  OAI21_X1 U48546 ( .A1(n2591), .A2(n15011), .B(n2590), .ZN(n2593) );
  INV_X2 U48548 ( .I(n64635), .ZN(n5348) );
  NOR2_X1 U48553 ( .A1(n64636), .A2(n25218), .ZN(n25507) );
  NOR2_X1 U48556 ( .A1(n41869), .A2(n41868), .ZN(n64636) );
  NOR2_X2 U48579 ( .A1(n23941), .A2(n22499), .ZN(n248) );
  NAND2_X2 U48587 ( .A1(n49783), .A2(n21623), .ZN(n48950) );
  XOR2_X1 U48589 ( .A1(n11420), .A2(n24112), .Z(n17340) );
  NOR2_X1 U48591 ( .A1(n24249), .A2(n1769), .ZN(n2592) );
  NAND2_X1 U48592 ( .A1(n52393), .A2(n52394), .ZN(n64637) );
  XOR2_X1 U48593 ( .A1(n44441), .A2(n44596), .Z(n64638) );
  NAND2_X1 U48607 ( .A1(n7076), .A2(n29529), .ZN(n64639) );
  NAND2_X1 U48616 ( .A1(n64927), .A2(n20705), .ZN(n3631) );
  NAND2_X2 U48631 ( .A1(n42140), .A2(n42127), .ZN(n41562) );
  XOR2_X1 U48632 ( .A1(n17691), .A2(n1214), .Z(n45096) );
  OAI21_X1 U48644 ( .A1(n23484), .A2(n41082), .B(n64641), .ZN(n39961) );
  NAND2_X1 U48653 ( .A1(n3344), .A2(n41082), .ZN(n64641) );
  NAND3_X2 U48654 ( .A1(n45313), .A2(n25179), .A3(n45312), .ZN(n50422) );
  NOR3_X1 U48666 ( .A1(n58735), .A2(n8968), .A3(n101), .ZN(n64645) );
  XOR2_X1 U48670 ( .A1(n64642), .A2(n39730), .Z(n60453) );
  AND2_X1 U48674 ( .A1(n55425), .A2(n1324), .Z(n337) );
  NAND2_X2 U48677 ( .A1(n14039), .A2(n14733), .ZN(n10986) );
  OAI21_X1 U48679 ( .A1(n48890), .A2(n24917), .B(n24916), .ZN(n64644) );
  NOR2_X2 U48681 ( .A1(n10958), .A2(n3658), .ZN(n49642) );
  NOR2_X1 U48684 ( .A1(n8965), .A2(n64645), .ZN(n8964) );
  INV_X2 U48691 ( .I(n64647), .ZN(n65270) );
  XOR2_X1 U48694 ( .A1(n3499), .A2(n6207), .Z(n64647) );
  OR2_X1 U48731 ( .A1(n55474), .A2(n58514), .Z(n52925) );
  XOR2_X1 U48737 ( .A1(n25986), .A2(n46288), .Z(n44939) );
  NAND2_X2 U48757 ( .A1(n56191), .A2(n18175), .ZN(n61432) );
  XOR2_X1 U48774 ( .A1(n64650), .A2(n6216), .Z(n6961) );
  XOR2_X1 U48778 ( .A1(n14316), .A2(n23882), .Z(n64650) );
  NAND2_X2 U48783 ( .A1(n57901), .A2(n61354), .ZN(n55287) );
  BUF_X2 U48784 ( .I(n24981), .Z(n64651) );
  XOR2_X1 U48785 ( .A1(n38960), .A2(n38321), .Z(n22061) );
  XOR2_X1 U48786 ( .A1(n19303), .A2(n23882), .Z(n38960) );
  INV_X2 U48787 ( .I(n17059), .ZN(n45246) );
  NAND2_X2 U48789 ( .A1(n14698), .A2(n58406), .ZN(n17059) );
  XOR2_X1 U48811 ( .A1(n4234), .A2(n50797), .Z(n9936) );
  NOR2_X2 U48869 ( .A1(n51263), .A2(n8367), .ZN(n6379) );
  NAND2_X1 U48889 ( .A1(n12212), .A2(n2712), .ZN(n64656) );
  XOR2_X1 U48890 ( .A1(n23957), .A2(n45095), .Z(n64658) );
  NAND2_X2 U48891 ( .A1(n64659), .A2(n2247), .ZN(n41094) );
  AND2_X2 U48909 ( .A1(n5532), .A2(n57603), .Z(n11929) );
  NOR2_X2 U48912 ( .A1(n20588), .A2(n20589), .ZN(n56516) );
  NAND3_X1 U48913 ( .A1(n61246), .A2(n11837), .A3(n11833), .ZN(n64700) );
  OR2_X2 U48929 ( .A1(n47501), .A2(n863), .Z(n9907) );
  NAND3_X2 U48930 ( .A1(n5570), .A2(n54996), .A3(n63194), .ZN(n55277) );
  NOR2_X2 U48931 ( .A1(n5569), .A2(n21169), .ZN(n5570) );
  NAND3_X1 U48948 ( .A1(n43374), .A2(n42755), .A3(n25933), .ZN(n64660) );
  NAND2_X2 U48952 ( .A1(n17364), .A2(n36748), .ZN(n12004) );
  XOR2_X1 U48959 ( .A1(n12478), .A2(n46427), .Z(n22662) );
  NAND2_X2 U48976 ( .A1(n16555), .A2(n16551), .ZN(n46427) );
  NAND2_X1 U48985 ( .A1(n18077), .A2(n34569), .ZN(n10528) );
  NAND2_X2 U48999 ( .A1(n61762), .A2(n64661), .ZN(n45235) );
  NOR2_X2 U49001 ( .A1(n49465), .A2(n4888), .ZN(n49462) );
  INV_X4 U49004 ( .I(n55401), .ZN(n65011) );
  XOR2_X1 U49029 ( .A1(n7811), .A2(n1011), .Z(n59877) );
  NOR2_X1 U49051 ( .A1(n54103), .A2(n54104), .ZN(n64662) );
  XOR2_X1 U49058 ( .A1(n9739), .A2(n44421), .Z(n46202) );
  AND2_X1 U49060 ( .A1(n59936), .A2(n32829), .Z(n64952) );
  NAND3_X2 U49070 ( .A1(n15265), .A2(n44002), .A3(n25899), .ZN(n48868) );
  NAND2_X2 U49094 ( .A1(n12382), .A2(n25141), .ZN(n3505) );
  BUF_X2 U49119 ( .I(n42361), .Z(n64663) );
  XOR2_X1 U49137 ( .A1(n19612), .A2(n19613), .Z(n10455) );
  NAND2_X1 U49138 ( .A1(n12039), .A2(n23119), .ZN(n32893) );
  NOR2_X2 U49142 ( .A1(n31509), .A2(n34627), .ZN(n23119) );
  AND2_X1 U49145 ( .A1(n3654), .A2(n3596), .Z(n3771) );
  BUF_X2 U49146 ( .I(n60285), .Z(n64667) );
  NAND2_X2 U49152 ( .A1(n3745), .A2(n3746), .ZN(n65127) );
  INV_X2 U49246 ( .I(n48868), .ZN(n1292) );
  XOR2_X1 U49247 ( .A1(n31762), .A2(n708), .Z(n7691) );
  XOR2_X1 U49266 ( .A1(n8667), .A2(n31456), .Z(n31762) );
  XOR2_X1 U49271 ( .A1(n64670), .A2(n53487), .Z(Plaintext[26]) );
  AND2_X1 U49305 ( .A1(n53485), .A2(n53513), .Z(n64671) );
  XOR2_X1 U49381 ( .A1(n64673), .A2(n18720), .Z(n2892) );
  XOR2_X1 U49414 ( .A1(n61265), .A2(n8575), .Z(n64673) );
  NOR3_X2 U49424 ( .A1(n8708), .A2(n65168), .A3(n8710), .ZN(n8707) );
  NOR2_X2 U49471 ( .A1(n13714), .A2(n64799), .ZN(n13713) );
  NAND3_X2 U49474 ( .A1(n41972), .A2(n2160), .A3(n20244), .ZN(n42686) );
  AOI21_X2 U49545 ( .A1(n15466), .A2(n34502), .B(n34640), .ZN(n64676) );
  NAND3_X1 U49554 ( .A1(n44454), .A2(n44455), .A3(n54587), .ZN(n7247) );
  XOR2_X1 U49581 ( .A1(n18114), .A2(n46597), .Z(n64678) );
  NOR2_X1 U49617 ( .A1(n34941), .A2(n21489), .ZN(n26170) );
  AOI21_X2 U49652 ( .A1(n50520), .A2(n50521), .B(n50522), .ZN(n52627) );
  OAI21_X1 U49654 ( .A1(n64680), .A2(n18910), .B(n14630), .ZN(n5019) );
  NOR2_X1 U49708 ( .A1(n45559), .A2(n1295), .ZN(n64680) );
  OR2_X1 U49709 ( .A1(n6033), .A2(n60633), .Z(n19924) );
  NAND2_X2 U49736 ( .A1(n19645), .A2(n65074), .ZN(n1652) );
  XOR2_X1 U49794 ( .A1(n52369), .A2(n51645), .Z(n6486) );
  XOR2_X1 U49859 ( .A1(n51028), .A2(n1289), .Z(n51645) );
  BUF_X2 U49866 ( .I(n24873), .Z(n64683) );
  XOR2_X1 U49907 ( .A1(n8021), .A2(n7679), .Z(n4256) );
  NOR2_X1 U49953 ( .A1(n7485), .A2(n18469), .ZN(n48793) );
  NAND2_X2 U49959 ( .A1(n58492), .A2(n58491), .ZN(n54961) );
  XOR2_X1 U49960 ( .A1(n64685), .A2(n18699), .Z(Plaintext[90]) );
  NOR3_X2 U49963 ( .A1(n8406), .A2(n8413), .A3(n8409), .ZN(n64685) );
  NAND3_X2 U49997 ( .A1(n64686), .A2(n14744), .A3(n28102), .ZN(n65168) );
  XOR2_X1 U50151 ( .A1(n64687), .A2(n57301), .Z(n6698) );
  XOR2_X1 U50154 ( .A1(n19680), .A2(n18124), .Z(n64687) );
  NOR2_X2 U50158 ( .A1(n2162), .A2(n64689), .ZN(n2161) );
  NAND3_X1 U50169 ( .A1(n64690), .A2(n540), .A3(n54963), .ZN(n54302) );
  XOR2_X1 U50171 ( .A1(n24005), .A2(n23852), .Z(n2070) );
  INV_X2 U50177 ( .I(n18063), .ZN(n54561) );
  NAND2_X2 U50178 ( .A1(n57857), .A2(n15097), .ZN(n18063) );
  OR2_X2 U50180 ( .A1(n59936), .A2(n32829), .Z(n33995) );
  NOR2_X1 U50191 ( .A1(n1770), .A2(n35142), .ZN(n9933) );
  NOR2_X2 U50192 ( .A1(n64691), .A2(n35977), .ZN(n20132) );
  NAND2_X2 U50201 ( .A1(n258), .A2(n20134), .ZN(n64691) );
  XOR2_X1 U50215 ( .A1(n47757), .A2(n50849), .Z(n64692) );
  OR2_X2 U50232 ( .A1(n3654), .A2(n61716), .Z(n48977) );
  XOR2_X1 U50274 ( .A1(n14086), .A2(n45110), .Z(n4453) );
  INV_X2 U50275 ( .I(n14087), .ZN(n14086) );
  NOR2_X2 U50278 ( .A1(n64695), .A2(n64693), .ZN(n25553) );
  NAND2_X2 U50305 ( .A1(n11882), .A2(n64696), .ZN(n18854) );
  NAND2_X1 U50375 ( .A1(n26007), .A2(n64697), .ZN(n64696) );
  OR2_X1 U50378 ( .A1(n47963), .A2(n47962), .Z(n64697) );
  INV_X2 U50390 ( .I(n64698), .ZN(n8453) );
  XOR2_X1 U50412 ( .A1(n6544), .A2(n14339), .Z(n11733) );
  NAND2_X2 U50425 ( .A1(n6549), .A2(n6548), .ZN(n6544) );
  OR2_X2 U50445 ( .A1(n16631), .A2(n17411), .Z(n21964) );
  NAND4_X2 U50457 ( .A1(n64700), .A2(n15178), .A3(n10115), .A4(n3156), .ZN(
        n23049) );
  NOR2_X1 U50472 ( .A1(n18767), .A2(n58855), .ZN(n64701) );
  NOR4_X2 U50487 ( .A1(n16387), .A2(n16386), .A3(n11280), .A4(n43277), .ZN(
        n10316) );
  XOR2_X1 U50488 ( .A1(n51689), .A2(n64702), .Z(n60744) );
  XOR2_X1 U50501 ( .A1(n18685), .A2(n25316), .Z(n64702) );
  NAND2_X2 U50534 ( .A1(n16338), .A2(n64717), .ZN(n36953) );
  NOR2_X2 U50579 ( .A1(n6435), .A2(n59093), .ZN(n9185) );
  XOR2_X1 U50580 ( .A1(n46150), .A2(n45040), .Z(n10265) );
  NAND2_X2 U50582 ( .A1(n43546), .A2(n43547), .ZN(n45040) );
  NOR2_X2 U50585 ( .A1(n64703), .A2(n41828), .ZN(n61164) );
  NAND3_X2 U50599 ( .A1(n61906), .A2(n41824), .A3(n41822), .ZN(n64703) );
  NOR2_X2 U50603 ( .A1(n65261), .A2(n5599), .ZN(n51687) );
  XOR2_X1 U50611 ( .A1(n17404), .A2(n17405), .Z(n39382) );
  XOR2_X1 U50612 ( .A1(n64705), .A2(n23573), .Z(n36369) );
  XOR2_X1 U50613 ( .A1(n39690), .A2(n36360), .Z(n64705) );
  NAND3_X2 U50616 ( .A1(n36888), .A2(n34914), .A3(n36889), .ZN(n20616) );
  NAND2_X2 U50617 ( .A1(n15552), .A2(n35026), .ZN(n35021) );
  XOR2_X1 U50619 ( .A1(n37777), .A2(n64716), .Z(n59932) );
  XOR2_X1 U50620 ( .A1(n37121), .A2(n24169), .Z(n64716) );
  AOI21_X1 U50621 ( .A1(n21475), .A2(n902), .B(n21473), .ZN(n64717) );
  XOR2_X1 U50630 ( .A1(n7959), .A2(n11957), .Z(n14871) );
  NOR2_X2 U50644 ( .A1(n58826), .A2(n56107), .ZN(n56081) );
  NAND2_X2 U50654 ( .A1(n36264), .A2(n3171), .ZN(n36616) );
  NOR2_X1 U50655 ( .A1(n64720), .A2(n54399), .ZN(n54406) );
  AOI21_X1 U50674 ( .A1(n54396), .A2(n54397), .B(n2676), .ZN(n64720) );
  NOR2_X2 U50677 ( .A1(n64723), .A2(n64721), .ZN(n21565) );
  XOR2_X1 U50682 ( .A1(n51035), .A2(n50717), .Z(n19189) );
  XOR2_X1 U50694 ( .A1(n31323), .A2(n58837), .Z(n64938) );
  OR2_X2 U50700 ( .A1(n24352), .A2(n12772), .Z(n58218) );
  AOI21_X2 U50701 ( .A1(n10178), .A2(n31129), .B(n358), .ZN(n32002) );
  NAND2_X2 U50703 ( .A1(n15319), .A2(n24394), .ZN(n49172) );
  XOR2_X1 U50714 ( .A1(n6961), .A2(n6363), .Z(n6960) );
  XOR2_X1 U50748 ( .A1(n64727), .A2(n25996), .Z(n12307) );
  XOR2_X1 U50754 ( .A1(n39468), .A2(n18056), .Z(n64727) );
  INV_X2 U50755 ( .I(n41060), .ZN(n64728) );
  NAND2_X2 U50763 ( .A1(n64728), .A2(n41889), .ZN(n16220) );
  NOR2_X1 U50766 ( .A1(n9253), .A2(n52817), .ZN(n64729) );
  INV_X1 U50767 ( .I(n9252), .ZN(n64730) );
  AND2_X2 U50784 ( .A1(n24615), .A2(n20826), .Z(n7931) );
  NAND2_X1 U50787 ( .A1(n23689), .A2(n60285), .ZN(n35753) );
  NAND2_X2 U50791 ( .A1(n1533), .A2(n24054), .ZN(n60285) );
  NAND2_X1 U50792 ( .A1(n56570), .A2(n61836), .ZN(n64733) );
  INV_X2 U50801 ( .I(n64734), .ZN(n40832) );
  OAI22_X1 U50809 ( .A1(n32), .A2(n31), .B1(n45563), .B2(n47610), .ZN(n17564)
         );
  XOR2_X1 U50818 ( .A1(n5576), .A2(n43961), .Z(n5575) );
  NOR2_X1 U50819 ( .A1(n25328), .A2(n41131), .ZN(n42339) );
  INV_X2 U50821 ( .I(n5846), .ZN(n703) );
  NAND2_X2 U50843 ( .A1(n58112), .A2(n25963), .ZN(n5846) );
  NOR2_X2 U50859 ( .A1(n5053), .A2(n64735), .ZN(n55099) );
  NAND2_X2 U50867 ( .A1(n21644), .A2(n11039), .ZN(n23838) );
  NAND2_X2 U50879 ( .A1(n2623), .A2(n24732), .ZN(n4546) );
  NOR2_X2 U50884 ( .A1(n64736), .A2(n42010), .ZN(n6112) );
  NAND2_X2 U50889 ( .A1(n43224), .A2(n5103), .ZN(n64736) );
  AND2_X1 U50900 ( .A1(n48903), .A2(n48904), .Z(n64737) );
  NOR2_X2 U50919 ( .A1(n1610), .A2(n54317), .ZN(n64978) );
  AND2_X1 U50921 ( .A1(n54097), .A2(n54096), .Z(n64739) );
  OAI21_X1 U50932 ( .A1(n61851), .A2(n13505), .B(n3837), .ZN(n3835) );
  AND2_X1 U50933 ( .A1(n41193), .A2(n63510), .Z(n17472) );
  AOI22_X1 U50940 ( .A1(n39846), .A2(n22638), .B1(n15441), .B2(n357), .ZN(
        n39848) );
  MUX2_X1 U50947 ( .I0(n47846), .I1(n47847), .S(n23361), .Z(n47848) );
  NOR2_X2 U50952 ( .A1(n8225), .A2(n47832), .ZN(n23361) );
  OR2_X1 U50953 ( .A1(n52950), .A2(n55438), .Z(n64741) );
  XOR2_X1 U50954 ( .A1(n7904), .A2(n39554), .Z(n8260) );
  XOR2_X1 U50979 ( .A1(n50995), .A2(n50994), .Z(n58500) );
  NAND2_X2 U50995 ( .A1(n64742), .A2(n11562), .ZN(n13321) );
  XOR2_X1 U51003 ( .A1(n39193), .A2(n1756), .Z(n39205) );
  XOR2_X1 U51027 ( .A1(n59826), .A2(n24204), .Z(n39193) );
  OR3_X1 U51030 ( .A1(n7241), .A2(n16995), .A3(n55204), .Z(n64743) );
  NAND3_X2 U51031 ( .A1(n42605), .A2(n23928), .A3(n23877), .ZN(n2121) );
  NOR2_X2 U51033 ( .A1(n43634), .A2(n16447), .ZN(n42622) );
  INV_X2 U51046 ( .I(n64744), .ZN(n53443) );
  NOR2_X2 U51052 ( .A1(n24318), .A2(n64750), .ZN(n64744) );
  NAND2_X2 U51063 ( .A1(n64745), .A2(n33515), .ZN(n59988) );
  NOR2_X1 U51067 ( .A1(n10047), .A2(n10046), .ZN(n64745) );
  AND2_X2 U51075 ( .A1(n42224), .A2(n61444), .Z(n41951) );
  INV_X2 U51078 ( .I(n33995), .ZN(n34194) );
  NAND2_X2 U51080 ( .A1(n64746), .A2(n2395), .ZN(n2394) );
  NOR2_X2 U51095 ( .A1(n2402), .A2(n21431), .ZN(n64746) );
  NOR2_X1 U51097 ( .A1(n12400), .A2(n21504), .ZN(n12399) );
  NOR2_X2 U51114 ( .A1(n20531), .A2(n6440), .ZN(n36063) );
  NOR2_X2 U51122 ( .A1(n60866), .A2(n40017), .ZN(n42936) );
  XOR2_X1 U51123 ( .A1(n16594), .A2(n39253), .Z(n64747) );
  NAND3_X2 U51128 ( .A1(n64748), .A2(n64951), .A3(n19805), .ZN(n19950) );
  XOR2_X1 U51138 ( .A1(n673), .A2(n18726), .Z(n45429) );
  XOR2_X1 U51139 ( .A1(n38289), .A2(n3145), .Z(n64749) );
  XOR2_X1 U51144 ( .A1(n31433), .A2(n32283), .Z(n3431) );
  BUF_X2 U51146 ( .I(n7588), .Z(n64751) );
  XOR2_X1 U51155 ( .A1(n59274), .A2(n21660), .Z(n31975) );
  NAND2_X1 U51178 ( .A1(n8840), .A2(n41953), .ZN(n4562) );
  AOI22_X1 U51179 ( .A1(n56569), .A2(n11121), .B1(n56570), .B2(n56571), .ZN(
        n64754) );
  INV_X2 U51184 ( .I(n33058), .ZN(n64755) );
  NAND2_X2 U51188 ( .A1(n33596), .A2(n35680), .ZN(n33300) );
  NOR2_X2 U51197 ( .A1(n23812), .A2(n24688), .ZN(n35680) );
  INV_X1 U51212 ( .I(n64756), .ZN(n60097) );
  OAI21_X1 U51213 ( .A1(n52787), .A2(n52788), .B(n57037), .ZN(n64756) );
  XOR2_X1 U51226 ( .A1(n14002), .A2(n64757), .Z(n22800) );
  XOR2_X1 U51236 ( .A1(n39395), .A2(n39384), .Z(n64757) );
  INV_X2 U51237 ( .I(n64759), .ZN(n50275) );
  NOR2_X2 U51240 ( .A1(n20138), .A2(n1209), .ZN(n64759) );
  XOR2_X1 U51259 ( .A1(n4759), .A2(n39590), .Z(n22719) );
  NAND3_X2 U51275 ( .A1(n64761), .A2(n40906), .A3(n64760), .ZN(n40911) );
  NAND2_X1 U51277 ( .A1(n40903), .A2(n41996), .ZN(n64760) );
  NAND2_X2 U51279 ( .A1(n4995), .A2(n20348), .ZN(n8812) );
  NAND2_X2 U51287 ( .A1(n64763), .A2(n16007), .ZN(n15511) );
  NOR2_X2 U51294 ( .A1(n22664), .A2(n64765), .ZN(n48362) );
  NAND2_X2 U51331 ( .A1(n64767), .A2(n50809), .ZN(n53146) );
  BUF_X2 U51343 ( .I(n1741), .Z(n64768) );
  NAND2_X2 U51351 ( .A1(n59261), .A2(n36422), .ZN(n36171) );
  XOR2_X1 U51381 ( .A1(n64769), .A2(n52344), .Z(n52346) );
  NOR3_X2 U51383 ( .A1(n301), .A2(n3853), .A3(n3852), .ZN(n64770) );
  NAND2_X2 U51419 ( .A1(n64771), .A2(n42170), .ZN(n3854) );
  INV_X2 U51437 ( .I(n41778), .ZN(n64771) );
  NAND2_X2 U51438 ( .A1(n42171), .A2(n64346), .ZN(n41778) );
  NAND2_X2 U51440 ( .A1(n1274), .A2(n38134), .ZN(n42523) );
  XOR2_X1 U51442 ( .A1(n61926), .A2(n31519), .Z(n60247) );
  XOR2_X1 U51450 ( .A1(n2553), .A2(n25203), .Z(n31519) );
  XOR2_X1 U51451 ( .A1(n1111), .A2(n50775), .Z(n64775) );
  NOR2_X2 U51454 ( .A1(n1298), .A2(n24779), .ZN(n43320) );
  NOR2_X1 U51456 ( .A1(n58312), .A2(n64776), .ZN(n58146) );
  NOR2_X2 U51479 ( .A1(n23248), .A2(n7095), .ZN(n64778) );
  NAND4_X1 U51505 ( .A1(n50814), .A2(n53145), .A3(n26135), .A4(n3525), .ZN(
        n60789) );
  NOR2_X2 U51507 ( .A1(n20735), .A2(n4808), .ZN(n53145) );
  NAND3_X2 U51508 ( .A1(n43082), .A2(n43843), .A3(n43081), .ZN(n64777) );
  NAND3_X1 U51516 ( .A1(n50807), .A2(n50806), .A3(n23563), .ZN(n50808) );
  BUF_X2 U51518 ( .I(n4660), .Z(n64779) );
  NAND3_X1 U51534 ( .A1(n17436), .A2(n51877), .A3(n64780), .ZN(n17434) );
  NOR3_X2 U51544 ( .A1(n22545), .A2(n54268), .A3(n54254), .ZN(n54214) );
  NOR3_X2 U51546 ( .A1(n64781), .A2(n2008), .A3(n2006), .ZN(n24334) );
  INV_X2 U51553 ( .I(n27399), .ZN(n64781) );
  NOR2_X2 U51557 ( .A1(n3433), .A2(n27985), .ZN(n27399) );
  NOR2_X2 U51572 ( .A1(n64783), .A2(n64782), .ZN(n31908) );
  NAND2_X2 U51593 ( .A1(n59311), .A2(n64784), .ZN(n12299) );
  NAND2_X1 U51594 ( .A1(n59085), .A2(n58461), .ZN(n64784) );
  INV_X2 U51597 ( .I(n52825), .ZN(n52814) );
  NAND2_X2 U51608 ( .A1(n24318), .A2(n64750), .ZN(n52825) );
  NAND4_X2 U51618 ( .A1(n54967), .A2(n54977), .A3(n54968), .A4(n54975), .ZN(
        n64785) );
  NOR2_X1 U51623 ( .A1(n65020), .A2(n40867), .ZN(n64787) );
  BUF_X2 U51625 ( .I(n14354), .Z(n64788) );
  NAND2_X2 U51626 ( .A1(n64789), .A2(n53523), .ZN(n14020) );
  OAI21_X2 U51627 ( .A1(n14021), .A2(n17101), .B(n53515), .ZN(n64789) );
  NAND2_X1 U51628 ( .A1(n64790), .A2(n1652), .ZN(n12201) );
  NAND2_X2 U51657 ( .A1(n64571), .A2(n40528), .ZN(n39137) );
  NAND4_X2 U51659 ( .A1(n59741), .A2(n18929), .A3(n54098), .A4(n51637), .ZN(
        n58568) );
  BUF_X2 U51690 ( .I(n32058), .Z(n64794) );
  AND2_X2 U51699 ( .A1(n16666), .A2(n10202), .Z(n12497) );
  XOR2_X1 U51700 ( .A1(n64795), .A2(n24822), .Z(n8514) );
  XOR2_X1 U51703 ( .A1(n33911), .A2(n33912), .Z(n64795) );
  OR2_X1 U51706 ( .A1(n45432), .A2(n45411), .Z(n46824) );
  XOR2_X1 U51715 ( .A1(n14825), .A2(n45431), .Z(n45432) );
  XOR2_X1 U51738 ( .A1(n33898), .A2(n33896), .Z(n23463) );
  XOR2_X1 U51753 ( .A1(n13896), .A2(n52637), .Z(n64796) );
  BUF_X2 U51763 ( .I(n35915), .Z(n64797) );
  NOR3_X1 U51777 ( .A1(n18341), .A2(n59531), .A3(n60826), .ZN(n37907) );
  XOR2_X1 U51794 ( .A1(n32668), .A2(n32667), .Z(n32675) );
  XOR2_X1 U51799 ( .A1(n23719), .A2(n14665), .Z(n32668) );
  NAND2_X2 U51831 ( .A1(n36898), .A2(n36533), .ZN(n33122) );
  OAI21_X1 U51832 ( .A1(n36047), .A2(n36048), .B(n20060), .ZN(n11302) );
  NAND2_X1 U51837 ( .A1(n41804), .A2(n40358), .ZN(n13384) );
  INV_X4 U51851 ( .I(n50041), .ZN(n50043) );
  AND3_X1 U51857 ( .A1(n46941), .A2(n9758), .A3(n64800), .Z(n59536) );
  XOR2_X1 U51903 ( .A1(n64801), .A2(n1056), .Z(n6241) );
  XOR2_X1 U51950 ( .A1(n59804), .A2(n6568), .Z(n64801) );
  INV_X2 U51951 ( .I(n64802), .ZN(n22701) );
  XOR2_X1 U51952 ( .A1(n26220), .A2(n26219), .Z(n64802) );
  NAND2_X2 U51958 ( .A1(n17088), .A2(n64803), .ZN(n16868) );
  NAND4_X1 U51976 ( .A1(n53292), .A2(n64804), .A3(n53289), .A4(n53291), .ZN(
        Plaintext[16]) );
  NAND2_X1 U51980 ( .A1(n13238), .A2(n13237), .ZN(n64804) );
  XOR2_X1 U51994 ( .A1(n60497), .A2(n2215), .Z(n64805) );
  AND2_X2 U51996 ( .A1(n10455), .A2(n647), .Z(n12314) );
  XOR2_X1 U52008 ( .A1(n64806), .A2(n38578), .Z(n37978) );
  XOR2_X1 U52017 ( .A1(n23655), .A2(n37975), .Z(n64806) );
  NOR2_X1 U52018 ( .A1(n36551), .A2(n22454), .ZN(n6770) );
  NOR3_X2 U52025 ( .A1(n58366), .A2(n58668), .A3(n28966), .ZN(n28976) );
  XOR2_X1 U52049 ( .A1(n64807), .A2(n53787), .Z(Plaintext[43]) );
  NAND2_X2 U52050 ( .A1(n55982), .A2(n1616), .ZN(n18597) );
  BUF_X2 U52057 ( .I(n56435), .Z(n64808) );
  NAND2_X2 U52079 ( .A1(n35296), .A2(n21464), .ZN(n34733) );
  OR2_X2 U52107 ( .A1(n24890), .A2(n22918), .Z(n8026) );
  BUF_X2 U52123 ( .I(n26431), .Z(n64809) );
  XOR2_X1 U52137 ( .A1(n32486), .A2(n64811), .Z(n8837) );
  XOR2_X1 U52143 ( .A1(n8839), .A2(n32000), .Z(n64811) );
  BUF_X2 U52147 ( .I(n25256), .Z(n64812) );
  BUF_X2 U52170 ( .I(n55397), .Z(n64813) );
  NAND2_X2 U52179 ( .A1(n61237), .A2(n43155), .ZN(n43167) );
  XOR2_X1 U52207 ( .A1(n44634), .A2(n64814), .Z(n31997) );
  XOR2_X1 U52215 ( .A1(n45830), .A2(n39478), .Z(n64814) );
  XOR2_X1 U52216 ( .A1(n44389), .A2(n22650), .Z(n44922) );
  NAND2_X1 U52224 ( .A1(n7469), .A2(n64980), .ZN(n8396) );
  NAND3_X2 U52252 ( .A1(n1838), .A2(n18736), .A3(n17413), .ZN(n29091) );
  XOR2_X1 U52253 ( .A1(n64815), .A2(n61152), .Z(n13475) );
  XOR2_X1 U52254 ( .A1(n17758), .A2(n18467), .Z(n64815) );
  NAND2_X1 U52284 ( .A1(n10279), .A2(n64817), .ZN(n26173) );
  NOR2_X1 U52314 ( .A1(n64819), .A2(n64818), .ZN(n64817) );
  NOR2_X1 U52331 ( .A1(n36722), .A2(n21468), .ZN(n64819) );
  NOR3_X2 U52335 ( .A1(n22000), .A2(n64820), .A3(n16091), .ZN(n21999) );
  NOR2_X2 U52368 ( .A1(n3054), .A2(n3055), .ZN(n50141) );
  INV_X2 U52369 ( .I(n64822), .ZN(n24870) );
  BUF_X2 U52371 ( .I(n49005), .Z(n64823) );
  NAND2_X2 U52393 ( .A1(n5628), .A2(n23738), .ZN(n49020) );
  XOR2_X1 U52396 ( .A1(n44348), .A2(n3941), .Z(n64824) );
  XOR2_X1 U52406 ( .A1(n44732), .A2(n64827), .Z(n16701) );
  XOR2_X1 U52415 ( .A1(n17870), .A2(n17868), .Z(n60283) );
  XOR2_X1 U52416 ( .A1(n23668), .A2(n64828), .Z(n44397) );
  XOR2_X1 U52417 ( .A1(n20073), .A2(n44948), .Z(n64828) );
  AND3_X1 U52419 ( .A1(n64829), .A2(n56995), .A3(n56996), .Z(n22969) );
  XOR2_X1 U52482 ( .A1(n62611), .A2(n10683), .Z(n64831) );
  NAND2_X2 U52491 ( .A1(n54558), .A2(n18425), .ZN(n54548) );
  NAND3_X2 U52507 ( .A1(n7056), .A2(n10108), .A3(n4747), .ZN(n57582) );
  INV_X1 U52548 ( .I(n34186), .ZN(n31417) );
  NOR2_X2 U52554 ( .A1(n21592), .A2(n21346), .ZN(n21699) );
  XOR2_X1 U52563 ( .A1(n2803), .A2(n64834), .Z(n24200) );
  XOR2_X1 U52575 ( .A1(n15225), .A2(n39713), .Z(n61026) );
  NAND2_X2 U52586 ( .A1(n61134), .A2(n17950), .ZN(n15044) );
  NOR2_X1 U52588 ( .A1(n5813), .A2(n4424), .ZN(n64835) );
  OR2_X2 U52596 ( .A1(n28349), .A2(n14903), .Z(n27529) );
  XOR2_X1 U52635 ( .A1(n1752), .A2(n17533), .Z(n38525) );
  NAND2_X2 U52636 ( .A1(n64836), .A2(n57044), .ZN(n57055) );
  BUF_X2 U52637 ( .I(n1542), .Z(n64838) );
  OR2_X2 U52658 ( .A1(n15597), .A2(n47653), .Z(n5145) );
  XOR2_X1 U52669 ( .A1(n14294), .A2(n14293), .Z(n15597) );
  OR2_X2 U52672 ( .A1(n57048), .A2(n24318), .Z(n57037) );
  XOR2_X1 U52703 ( .A1(n44104), .A2(n44105), .Z(n64839) );
  XOR2_X1 U52704 ( .A1(n46202), .A2(n46210), .Z(n18888) );
  NOR3_X2 U52709 ( .A1(n57993), .A2(n19409), .A3(n64840), .ZN(n52216) );
  NAND2_X1 U52740 ( .A1(n52190), .A2(n57720), .ZN(n64842) );
  XOR2_X1 U52745 ( .A1(n52175), .A2(n6141), .Z(n64843) );
  XOR2_X1 U52754 ( .A1(n17438), .A2(n64844), .Z(n59597) );
  XOR2_X1 U52762 ( .A1(n44610), .A2(n57432), .Z(n64844) );
  BUF_X2 U52765 ( .I(n56942), .Z(n64845) );
  XOR2_X1 U52767 ( .A1(n64846), .A2(n114), .Z(n5803) );
  OR2_X1 U52773 ( .A1(n376), .A2(n20138), .Z(n48025) );
  AOI21_X1 U52777 ( .A1(n11652), .A2(n21612), .B(n9899), .ZN(n21611) );
  NAND3_X2 U52797 ( .A1(n28160), .A2(n64847), .A3(n28159), .ZN(n58211) );
  NAND3_X1 U52806 ( .A1(n28158), .A2(n29319), .A3(n29322), .ZN(n64847) );
  NOR2_X2 U52855 ( .A1(n55985), .A2(n14879), .ZN(n51256) );
  NOR2_X2 U52877 ( .A1(n64848), .A2(n2999), .ZN(n2998) );
  BUF_X2 U52931 ( .I(n46863), .Z(n64849) );
  NOR3_X2 U52933 ( .A1(n64853), .A2(n39413), .A3(n64852), .ZN(n43281) );
  NAND2_X2 U52967 ( .A1(n39409), .A2(n39412), .ZN(n64853) );
  NOR2_X1 U52992 ( .A1(n64854), .A2(n11301), .ZN(n4926) );
  NAND2_X1 U53024 ( .A1(n36051), .A2(n18705), .ZN(n64854) );
  NAND3_X1 U53028 ( .A1(n56498), .A2(n56446), .A3(n56492), .ZN(n64855) );
  XOR2_X1 U53046 ( .A1(n38619), .A2(n64856), .Z(n17592) );
  XOR2_X1 U53050 ( .A1(n10360), .A2(n39495), .Z(n64856) );
  XOR2_X1 U53052 ( .A1(n64857), .A2(Key[131]), .Z(n11329) );
  NOR3_X2 U53068 ( .A1(n64858), .A2(n63510), .A3(n60567), .ZN(n40723) );
  INV_X2 U53069 ( .I(n38675), .ZN(n64858) );
  XOR2_X1 U53072 ( .A1(n12773), .A2(n25840), .Z(n39494) );
  AND2_X1 U53086 ( .A1(n34031), .A2(n34030), .Z(n64860) );
  XOR2_X1 U53102 ( .A1(n64861), .A2(n60903), .Z(n21279) );
  XOR2_X1 U53103 ( .A1(n17216), .A2(n6869), .Z(n64861) );
  AOI22_X1 U53104 ( .A1(n5547), .A2(n7109), .B1(n59279), .B2(n20540), .ZN(
        n23251) );
  NAND2_X2 U53116 ( .A1(n1230), .A2(n15477), .ZN(n5547) );
  OR2_X1 U53133 ( .A1(n7219), .A2(n8090), .Z(n8073) );
  XOR2_X1 U53142 ( .A1(n64863), .A2(n23509), .Z(n25403) );
  NAND4_X2 U53143 ( .A1(n11400), .A2(n11397), .A3(n16229), .A4(n64864), .ZN(
        n19322) );
  NAND2_X1 U53144 ( .A1(n57535), .A2(n17419), .ZN(n64864) );
  NOR3_X1 U53150 ( .A1(n42830), .A2(n64865), .A3(n42829), .ZN(n42831) );
  NAND3_X2 U53156 ( .A1(n2097), .A2(n28982), .A3(n19297), .ZN(n33058) );
  BUF_X2 U53157 ( .I(n1317), .Z(n64867) );
  NAND2_X2 U53173 ( .A1(n23924), .A2(n64868), .ZN(n59049) );
  AND3_X1 U53174 ( .A1(n21051), .A2(n7100), .A3(n54442), .Z(n64868) );
  NAND2_X2 U53209 ( .A1(n45889), .A2(n11673), .ZN(n64869) );
  XOR2_X1 U53210 ( .A1(n51617), .A2(n52418), .Z(n22763) );
  XOR2_X1 U53211 ( .A1(n52340), .A2(n11269), .Z(n52418) );
  AOI21_X2 U53228 ( .A1(n18351), .A2(n47821), .B(n64870), .ZN(n16186) );
  XOR2_X1 U53244 ( .A1(n64871), .A2(n60656), .Z(n45826) );
  XOR2_X1 U53245 ( .A1(n12712), .A2(n45822), .Z(n64871) );
  NOR2_X1 U53254 ( .A1(n63683), .A2(n23742), .ZN(n37209) );
  NAND2_X2 U53259 ( .A1(n5997), .A2(n5995), .ZN(n23742) );
  NOR2_X2 U53261 ( .A1(n6419), .A2(n6420), .ZN(n64873) );
  NAND2_X1 U53267 ( .A1(n56001), .A2(n64874), .ZN(n56005) );
  NAND2_X1 U53268 ( .A1(n56082), .A2(n64875), .ZN(n64874) );
  INV_X1 U53282 ( .I(n56081), .ZN(n64875) );
  NAND2_X2 U53296 ( .A1(n56047), .A2(n61740), .ZN(n56082) );
  XOR2_X1 U53297 ( .A1(n15511), .A2(n20308), .Z(n24178) );
  XOR2_X1 U53300 ( .A1(n64877), .A2(n15873), .Z(n2458) );
  BUF_X2 U53313 ( .I(n47773), .Z(n64878) );
  NAND4_X2 U53315 ( .A1(n7876), .A2(n7875), .A3(n20778), .A4(n7874), .ZN(n7581) );
  NOR3_X1 U53318 ( .A1(n54943), .A2(n54944), .A3(n64879), .ZN(n57325) );
  XNOR2_X1 U53353 ( .A1(n16558), .A2(n8450), .ZN(n65027) );
  AOI22_X2 U53355 ( .A1(n5547), .A2(n26625), .B1(n2706), .B2(n26624), .ZN(
        n26631) );
  NAND2_X1 U53357 ( .A1(n47825), .A2(n47611), .ZN(n47612) );
  AOI21_X1 U53361 ( .A1(n11053), .A2(n10574), .B(n18747), .ZN(n11051) );
  XOR2_X1 U53372 ( .A1(n38769), .A2(n1519), .Z(n7102) );
  XOR2_X1 U53375 ( .A1(n57218), .A2(n22160), .Z(n22744) );
  XOR2_X1 U53382 ( .A1(n64882), .A2(n18190), .Z(n13999) );
  BUF_X4 U53385 ( .I(n43989), .Z(n1495) );
  XOR2_X1 U53386 ( .A1(n51522), .A2(n52629), .Z(n5351) );
  OR2_X1 U53395 ( .A1(n40022), .A2(n40023), .Z(n64886) );
  NAND3_X1 U53411 ( .A1(n53397), .A2(n21982), .A3(n53535), .ZN(n50482) );
  OAI21_X1 U53419 ( .A1(n42931), .A2(n42930), .B(n42929), .ZN(n64889) );
  XOR2_X1 U53421 ( .A1(n64890), .A2(n12614), .Z(n9307) );
  XOR2_X1 U53429 ( .A1(n65104), .A2(n64891), .Z(n64890) );
  XNOR2_X1 U53430 ( .A1(n44519), .A2(n44520), .ZN(n65146) );
  AND2_X1 U53438 ( .A1(n54514), .A2(n54527), .Z(n23229) );
  NOR2_X2 U53440 ( .A1(n42843), .A2(n23811), .ZN(n64893) );
  BUF_X2 U53449 ( .I(n61048), .Z(n64894) );
  NOR3_X2 U53453 ( .A1(n26634), .A2(n26552), .A3(n26553), .ZN(n26554) );
  NOR2_X2 U53454 ( .A1(n37400), .A2(n36831), .ZN(n16426) );
  NOR2_X1 U53455 ( .A1(n50419), .A2(n48756), .ZN(n48762) );
  NOR2_X2 U53462 ( .A1(n10063), .A2(n50420), .ZN(n50419) );
  NOR2_X1 U53471 ( .A1(n32984), .A2(n9274), .ZN(n11721) );
  NAND2_X2 U53472 ( .A1(n61746), .A2(n64898), .ZN(n40361) );
  BUF_X2 U53476 ( .I(n1482), .Z(n64899) );
  XOR2_X1 U53487 ( .A1(n7308), .A2(n64900), .Z(n25647) );
  XOR2_X1 U53491 ( .A1(n11254), .A2(n14052), .Z(n64900) );
  OAI22_X1 U53503 ( .A1(n26547), .A2(n20898), .B1(n26311), .B2(n10419), .ZN(
        n26315) );
  NOR2_X2 U53505 ( .A1(n2315), .A2(n64901), .ZN(n2314) );
  AOI21_X2 U53506 ( .A1(n47820), .A2(n45967), .B(n1073), .ZN(n64901) );
  NOR2_X2 U53517 ( .A1(n64902), .A2(n13132), .ZN(n9190) );
  BUF_X2 U53519 ( .I(n28317), .Z(n64903) );
  NOR2_X2 U53522 ( .A1(n56381), .A2(n9555), .ZN(n16645) );
  NAND2_X2 U53523 ( .A1(n56541), .A2(n56539), .ZN(n9555) );
  NAND3_X1 U53525 ( .A1(n64904), .A2(n1813), .A3(n34677), .ZN(n34682) );
  AND2_X1 U53536 ( .A1(n31356), .A2(n2968), .Z(n34689) );
  INV_X1 U53540 ( .I(n65218), .ZN(n57258) );
  NAND2_X1 U53547 ( .A1(n25821), .A2(n64908), .ZN(n19794) );
  AOI22_X1 U53548 ( .A1(n31714), .A2(n31713), .B1(n19416), .B2(n57898), .ZN(
        n64908) );
  NAND2_X2 U53555 ( .A1(n20128), .A2(n15920), .ZN(n8618) );
  NOR2_X2 U53557 ( .A1(n57752), .A2(n57340), .ZN(n57751) );
  NOR2_X1 U53558 ( .A1(n28383), .A2(n28384), .ZN(n28386) );
  BUF_X2 U53565 ( .I(n13292), .Z(n64910) );
  NOR2_X2 U53582 ( .A1(n59753), .A2(n8181), .ZN(n30882) );
  NAND2_X2 U53583 ( .A1(n20869), .A2(n19201), .ZN(n52805) );
  NOR3_X2 U53599 ( .A1(n64911), .A2(n29562), .A3(n29911), .ZN(n24157) );
  OR2_X2 U53603 ( .A1(n32409), .A2(n22355), .Z(n9369) );
  BUF_X2 U53627 ( .I(n11084), .Z(n64914) );
  NAND3_X1 U53629 ( .A1(n32823), .A2(n32822), .A3(n34129), .ZN(n65081) );
  NAND3_X2 U53639 ( .A1(n11807), .A2(n14962), .A3(n11809), .ZN(n11806) );
  XOR2_X1 U53643 ( .A1(n11551), .A2(n24008), .Z(n33884) );
  XOR2_X1 U53644 ( .A1(n5575), .A2(n5572), .Z(n47704) );
  XOR2_X1 U53648 ( .A1(n64915), .A2(n3831), .Z(n3830) );
  XOR2_X1 U53650 ( .A1(n61665), .A2(n60777), .Z(n64915) );
  NOR2_X1 U53657 ( .A1(n2619), .A2(n53664), .ZN(n53671) );
  XOR2_X1 U53658 ( .A1(n64916), .A2(n53685), .Z(Plaintext[34]) );
  NAND2_X1 U53659 ( .A1(n53684), .A2(n53683), .ZN(n64916) );
  NAND3_X2 U53674 ( .A1(n38026), .A2(n40074), .A3(n21701), .ZN(n40068) );
  NAND2_X2 U53695 ( .A1(n64918), .A2(n64917), .ZN(n58949) );
  INV_X2 U53711 ( .I(n29857), .ZN(n64918) );
  XOR2_X1 U53726 ( .A1(n9297), .A2(n51700), .Z(n58157) );
  AOI22_X1 U53727 ( .A1(n2834), .A2(n2835), .B1(n53668), .B2(n53669), .ZN(
        n2833) );
  NAND3_X2 U53743 ( .A1(n5463), .A2(n58645), .A3(n20911), .ZN(n11155) );
  NOR2_X2 U53769 ( .A1(n4780), .A2(n48711), .ZN(n20911) );
  XOR2_X1 U53782 ( .A1(n58692), .A2(n61965), .Z(n24873) );
  XOR2_X1 U53785 ( .A1(n64919), .A2(n19810), .Z(n10367) );
  XOR2_X1 U53790 ( .A1(n11478), .A2(n11481), .Z(n64919) );
  XOR2_X1 U53827 ( .A1(n51629), .A2(n51940), .Z(n50648) );
  NOR3_X2 U53835 ( .A1(n48866), .A2(n22654), .A3(n48865), .ZN(n51629) );
  XOR2_X1 U53841 ( .A1(n52407), .A2(n64920), .Z(n51939) );
  XOR2_X1 U53844 ( .A1(n51936), .A2(n52058), .Z(n64920) );
  NAND2_X2 U53845 ( .A1(n36144), .A2(n60289), .ZN(n25690) );
  NAND2_X2 U53870 ( .A1(n1704), .A2(n41131), .ZN(n42726) );
  XOR2_X1 U53877 ( .A1(n10867), .A2(n64921), .Z(n10868) );
  XOR2_X1 U53878 ( .A1(n50179), .A2(n60642), .Z(n64921) );
  OAI21_X1 U53879 ( .A1(n64923), .A2(n49308), .B(n49318), .ZN(n48994) );
  NAND2_X1 U53885 ( .A1(n49610), .A2(n49602), .ZN(n64923) );
  NOR3_X2 U53894 ( .A1(n64925), .A2(n64924), .A3(n40855), .ZN(n10195) );
  AOI22_X1 U53916 ( .A1(n11170), .A2(n49612), .B1(n64926), .B2(n11171), .ZN(
        n65048) );
  NAND2_X2 U53917 ( .A1(n49610), .A2(n1638), .ZN(n49613) );
  NOR2_X1 U53943 ( .A1(n3633), .A2(n3634), .ZN(n64927) );
  NAND2_X2 U53979 ( .A1(n64928), .A2(n41510), .ZN(n41506) );
  OAI21_X2 U53998 ( .A1(n57983), .A2(n60268), .B(n41516), .ZN(n64928) );
  NAND3_X2 U54016 ( .A1(n40479), .A2(n163), .A3(n40481), .ZN(n40482) );
  NOR3_X1 U54017 ( .A1(n49585), .A2(n49584), .A3(n49586), .ZN(n49587) );
  XOR2_X1 U54048 ( .A1(n64930), .A2(n12258), .Z(n24646) );
  XOR2_X1 U54057 ( .A1(n19859), .A2(n8086), .Z(n59913) );
  AND2_X1 U54064 ( .A1(n57925), .A2(n41402), .Z(n17131) );
  NOR2_X2 U54069 ( .A1(n6685), .A2(n43733), .ZN(n14404) );
  NOR2_X2 U54080 ( .A1(n60516), .A2(n64931), .ZN(n36567) );
  NOR2_X2 U54088 ( .A1(n59541), .A2(n27150), .ZN(n29564) );
  INV_X2 U54111 ( .I(n64937), .ZN(n15740) );
  NAND2_X2 U54112 ( .A1(n8683), .A2(n8794), .ZN(n60232) );
  OAI22_X1 U54115 ( .A1(n20374), .A2(n40524), .B1(n40523), .B2(n40959), .ZN(
        n40525) );
  XOR2_X1 U54122 ( .A1(n4797), .A2(n4796), .Z(n5120) );
  INV_X2 U54123 ( .I(n42693), .ZN(n20244) );
  NAND3_X2 U54124 ( .A1(n20216), .A2(n40138), .A3(n24453), .ZN(n42693) );
  INV_X2 U54125 ( .I(n64939), .ZN(n764) );
  XOR2_X1 U54143 ( .A1(Ciphertext[21]), .A2(Key[40]), .Z(n64939) );
  XOR2_X1 U54145 ( .A1(n10001), .A2(n15393), .Z(n25659) );
  NOR3_X2 U54146 ( .A1(n16665), .A2(n18736), .A3(n64940), .ZN(n60804) );
  INV_X4 U54147 ( .I(n9334), .ZN(n43254) );
  NAND2_X2 U54161 ( .A1(n57427), .A2(n3871), .ZN(n9334) );
  XOR2_X1 U54168 ( .A1(n33054), .A2(n64941), .Z(n12428) );
  XOR2_X1 U54172 ( .A1(n20573), .A2(n61402), .Z(n64941) );
  NOR2_X2 U54173 ( .A1(n19167), .A2(n52475), .ZN(n55264) );
  XOR2_X1 U54203 ( .A1(n12093), .A2(n11914), .Z(n52544) );
  NOR2_X1 U54205 ( .A1(n32824), .A2(n65081), .ZN(n57593) );
  XOR2_X1 U54217 ( .A1(n24343), .A2(n60647), .Z(n65091) );
  XOR2_X1 U54218 ( .A1(n14798), .A2(n39254), .Z(n58891) );
  NOR2_X2 U54225 ( .A1(n54498), .A2(n54492), .ZN(n54316) );
  XOR2_X1 U54237 ( .A1(n18579), .A2(n1412), .Z(n21734) );
  NAND3_X1 U54239 ( .A1(n47189), .A2(n47188), .A3(n48529), .ZN(n7673) );
  XOR2_X1 U54252 ( .A1(n64947), .A2(n8554), .Z(n60003) );
  XOR2_X1 U54255 ( .A1(n11555), .A2(n44966), .Z(n64947) );
  XOR2_X1 U54268 ( .A1(n10709), .A2(n57623), .Z(n38405) );
  BUF_X2 U54269 ( .I(n40167), .Z(n64948) );
  XOR2_X1 U54298 ( .A1(n33054), .A2(n64949), .Z(n33060) );
  NAND2_X2 U54308 ( .A1(n33992), .A2(n5389), .ZN(n64951) );
  OR2_X2 U54309 ( .A1(n64939), .A2(n27559), .Z(n28383) );
  INV_X2 U54322 ( .I(n64952), .ZN(n18277) );
  NOR2_X2 U54326 ( .A1(n16854), .A2(n64953), .ZN(n16853) );
  NAND3_X2 U54329 ( .A1(n25070), .A2(n40341), .A3(n25072), .ZN(n64953) );
  NAND2_X1 U54331 ( .A1(n55429), .A2(n55430), .ZN(n19309) );
  NAND4_X2 U54333 ( .A1(n10113), .A2(n5129), .A3(n20653), .A4(n55721), .ZN(
        n55429) );
  BUF_X2 U54335 ( .I(n23606), .Z(n64960) );
  INV_X2 U54401 ( .I(n64961), .ZN(n1697) );
  NAND2_X2 U54405 ( .A1(n15142), .A2(n15140), .ZN(n20812) );
  NAND3_X2 U54414 ( .A1(n32299), .A2(n34946), .A3(n33757), .ZN(n59237) );
  NOR2_X1 U54425 ( .A1(n40283), .A2(n62656), .ZN(n4649) );
  NOR2_X2 U54429 ( .A1(n34600), .A2(n34599), .ZN(n36851) );
  NOR2_X1 U54438 ( .A1(n65038), .A2(n740), .ZN(n64963) );
  XOR2_X1 U54446 ( .A1(n51687), .A2(n23792), .Z(n3427) );
  AND2_X1 U54470 ( .A1(n56719), .A2(n23785), .Z(n56732) );
  XOR2_X1 U54474 ( .A1(n32420), .A2(n64964), .Z(n58462) );
  XOR2_X1 U54486 ( .A1(n32239), .A2(n32238), .Z(n64964) );
  XOR2_X1 U54496 ( .A1(n38402), .A2(n58135), .Z(n65060) );
  XOR2_X1 U54499 ( .A1(n11211), .A2(n38072), .Z(n38402) );
  XOR2_X1 U54504 ( .A1(n8668), .A2(n22146), .Z(n58841) );
  BUF_X2 U54529 ( .I(n34253), .Z(n64965) );
  NAND2_X2 U54532 ( .A1(n64966), .A2(n30389), .ZN(n19516) );
  OAI21_X2 U54553 ( .A1(n11954), .A2(n30384), .B(n19572), .ZN(n64966) );
  BUF_X2 U54565 ( .I(n36909), .Z(n64967) );
  XOR2_X1 U54568 ( .A1(n59776), .A2(n32418), .Z(n32421) );
  BUF_X2 U54585 ( .I(n33848), .Z(n64968) );
  AND2_X1 U54596 ( .A1(n40446), .A2(n40445), .Z(n64992) );
  BUF_X2 U54598 ( .I(n24091), .Z(n64970) );
  NAND3_X1 U54607 ( .A1(n43654), .A2(n43231), .A3(n2797), .ZN(n43145) );
  NAND2_X2 U54622 ( .A1(n65047), .A2(n3059), .ZN(n43242) );
  XOR2_X1 U54629 ( .A1(n14105), .A2(n57665), .Z(n92) );
  XOR2_X1 U54638 ( .A1(n64973), .A2(n59392), .Z(n59618) );
  NOR2_X2 U54640 ( .A1(n12957), .A2(n24337), .ZN(n64974) );
  AND2_X1 U54641 ( .A1(n42784), .A2(n41660), .Z(n41666) );
  AOI22_X1 U54702 ( .A1(n36293), .A2(n37112), .B1(n36755), .B2(n36756), .ZN(
        n36294) );
  NOR3_X1 U54734 ( .A1(n64975), .A2(n3541), .A3(n3537), .ZN(n3540) );
  AOI21_X1 U54743 ( .A1(n3543), .A2(n9187), .B(n53128), .ZN(n64975) );
  XOR2_X1 U54759 ( .A1(n50649), .A2(n23149), .Z(n50775) );
  XOR2_X1 U54760 ( .A1(n43960), .A2(n46279), .Z(n22803) );
  NAND2_X1 U54767 ( .A1(n27772), .A2(n27771), .ZN(n64976) );
  NAND2_X2 U54772 ( .A1(n48654), .A2(n46106), .ZN(n47489) );
  NAND2_X2 U54775 ( .A1(n57812), .A2(n12865), .ZN(n15539) );
  NAND2_X2 U54785 ( .A1(n19231), .A2(n25125), .ZN(n10127) );
  NAND2_X2 U54794 ( .A1(n36245), .A2(n36246), .ZN(n25125) );
  NAND3_X2 U54807 ( .A1(n23501), .A2(n1274), .A3(n64353), .ZN(n42516) );
  NAND2_X1 U54829 ( .A1(n23757), .A2(n64977), .ZN(n33364) );
  OR2_X1 U54843 ( .A1(n34157), .A2(n61197), .Z(n64977) );
  XOR2_X1 U54880 ( .A1(n9258), .A2(n9257), .Z(n4378) );
  XOR2_X1 U54904 ( .A1(n65025), .A2(n60062), .Z(n39359) );
  NAND3_X1 U54941 ( .A1(n54551), .A2(n18229), .A3(n58810), .ZN(n678) );
  XOR2_X1 U54942 ( .A1(n1945), .A2(n64979), .Z(n12084) );
  XOR2_X1 U54944 ( .A1(n8063), .A2(n5080), .Z(n64979) );
  NAND2_X1 U54945 ( .A1(n57414), .A2(n197), .ZN(n64980) );
  NOR3_X2 U54950 ( .A1(n61273), .A2(n64981), .A3(n5190), .ZN(n5189) );
  NOR2_X2 U54960 ( .A1(n42827), .A2(n6706), .ZN(n41363) );
  NAND2_X2 U54962 ( .A1(n57756), .A2(n4344), .ZN(n4346) );
  NOR2_X2 U54989 ( .A1(n59287), .A2(n4476), .ZN(n64983) );
  XOR2_X1 U54991 ( .A1(n24786), .A2(n52188), .Z(n21060) );
  BUF_X2 U54994 ( .I(n35775), .Z(n64984) );
  XOR2_X1 U54995 ( .A1(n16365), .A2(n64985), .Z(n32109) );
  XOR2_X1 U54996 ( .A1(n2260), .A2(n16367), .Z(n64985) );
  BUF_X2 U54997 ( .I(n42518), .Z(n64986) );
  AOI21_X1 U55000 ( .A1(n57260), .A2(n55082), .B(n64987), .ZN(n60524) );
  INV_X4 U55006 ( .I(n54568), .ZN(n54530) );
  NAND2_X2 U55011 ( .A1(n40695), .A2(n15258), .ZN(n41429) );
  BUF_X2 U55024 ( .I(n54952), .Z(n64989) );
  NAND3_X2 U55025 ( .A1(n8938), .A2(n8933), .A3(n59628), .ZN(n24731) );
  XOR2_X1 U55055 ( .A1(n64993), .A2(n22360), .Z(n59993) );
  XOR2_X1 U55058 ( .A1(n12317), .A2(n51830), .Z(n64993) );
  NOR2_X1 U55079 ( .A1(n61232), .A2(n59409), .ZN(n16824) );
  NAND2_X2 U55081 ( .A1(n548), .A2(n22908), .ZN(n45554) );
  NAND2_X1 U55093 ( .A1(n64996), .A2(n47750), .ZN(n18974) );
  NOR2_X1 U55109 ( .A1(n47747), .A2(n47746), .ZN(n64996) );
  NAND2_X1 U55113 ( .A1(n12521), .A2(n9026), .ZN(n12522) );
  NOR2_X2 U55119 ( .A1(n53901), .A2(n13939), .ZN(n53969) );
  NOR2_X2 U55126 ( .A1(n53900), .A2(n53899), .ZN(n53901) );
  NAND3_X2 U55127 ( .A1(n35923), .A2(n19130), .A3(n35924), .ZN(n24596) );
  OAI22_X1 U55130 ( .A1(n25661), .A2(n11345), .B1(n39418), .B2(n40075), .ZN(
        n38027) );
  NOR2_X2 U55131 ( .A1(n27756), .A2(n23569), .ZN(n28899) );
  NAND2_X2 U55135 ( .A1(n4547), .A2(n64946), .ZN(n43577) );
  NOR2_X2 U55137 ( .A1(n20326), .A2(n34268), .ZN(n35296) );
  AND2_X1 U55139 ( .A1(n40131), .A2(n6702), .Z(n20249) );
  XOR2_X1 U55142 ( .A1(n39758), .A2(n15002), .Z(n15001) );
  XOR2_X1 U55148 ( .A1(n21560), .A2(n16038), .Z(n39758) );
  XOR2_X1 U55155 ( .A1(n10243), .A2(n50493), .Z(n13485) );
  XOR2_X1 U55156 ( .A1(n64999), .A2(n620), .Z(Plaintext[145]) );
  NOR2_X2 U55158 ( .A1(n13169), .A2(n42507), .ZN(n42509) );
  NOR2_X2 U55159 ( .A1(n65001), .A2(n65000), .ZN(n8081) );
  XOR2_X1 U55165 ( .A1(n45111), .A2(n65003), .Z(n45120) );
  XOR2_X1 U55170 ( .A1(n23860), .A2(n46403), .Z(n45111) );
  INV_X2 U55173 ( .I(n7541), .ZN(n45208) );
  NAND2_X2 U55174 ( .A1(n13746), .A2(n24759), .ZN(n7541) );
  NOR2_X2 U55175 ( .A1(n59078), .A2(n61350), .ZN(n33117) );
  XOR2_X1 U55179 ( .A1(n51721), .A2(n65004), .Z(n5353) );
  XOR2_X1 U55180 ( .A1(n64697), .A2(n51527), .Z(n65004) );
  XOR2_X1 U55190 ( .A1(n18829), .A2(n20446), .Z(n39369) );
  XOR2_X1 U55201 ( .A1(n31632), .A2(n65006), .Z(n4631) );
  XOR2_X1 U55212 ( .A1(n64340), .A2(n31072), .Z(n65006) );
  NAND3_X1 U55234 ( .A1(n47734), .A2(n47735), .A3(n47736), .ZN(n47741) );
  OAI22_X1 U55237 ( .A1(n48021), .A2(n8347), .B1(n25128), .B2(n18975), .ZN(
        n48022) );
  NAND2_X2 U55253 ( .A1(n54196), .A2(n54207), .ZN(n65007) );
  OR2_X1 U55258 ( .A1(n49263), .A2(n11795), .Z(n9455) );
  NAND2_X2 U55259 ( .A1(n14676), .A2(n48023), .ZN(n50929) );
  XOR2_X1 U55266 ( .A1(n65008), .A2(n22199), .Z(n14671) );
  XOR2_X1 U55282 ( .A1(n58782), .A2(n59501), .Z(n65008) );
  NAND2_X1 U55290 ( .A1(n54982), .A2(n65009), .ZN(n261) );
  NAND2_X2 U55312 ( .A1(n65011), .A2(n65010), .ZN(n65009) );
  XOR2_X1 U55313 ( .A1(n10992), .A2(n11751), .Z(n38071) );
  NOR3_X2 U55315 ( .A1(n45950), .A2(n65012), .A3(n4713), .ZN(n49106) );
  INV_X2 U55319 ( .I(n65013), .ZN(n54523) );
  NAND2_X2 U55320 ( .A1(n29916), .A2(n14202), .ZN(n29560) );
  XOR2_X1 U55323 ( .A1(n51017), .A2(n51016), .Z(n51018) );
  NAND2_X2 U55336 ( .A1(n10157), .A2(n17017), .ZN(n51017) );
  NAND2_X2 U55350 ( .A1(n14189), .A2(n36749), .ZN(n36335) );
  NOR2_X2 U55375 ( .A1(n24981), .A2(n24250), .ZN(n43003) );
  NAND2_X2 U55397 ( .A1(n2064), .A2(n34725), .ZN(n32924) );
  NAND3_X2 U55412 ( .A1(n24745), .A2(n19979), .A3(n15993), .ZN(n19980) );
  NAND3_X1 U55413 ( .A1(n4175), .A2(n6984), .A3(n8976), .ZN(n12450) );
  XOR2_X1 U55418 ( .A1(n5009), .A2(n23693), .Z(n33880) );
  NAND2_X2 U55427 ( .A1(n19728), .A2(n56477), .ZN(n56462) );
  INV_X2 U55430 ( .I(n19647), .ZN(n17272) );
  XOR2_X1 U55445 ( .A1(n65014), .A2(n1144), .Z(n4403) );
  XOR2_X1 U55446 ( .A1(n6031), .A2(n61220), .Z(n61219) );
  XOR2_X1 U55460 ( .A1(n15401), .A2(n22108), .Z(n254) );
  XOR2_X1 U55471 ( .A1(n65015), .A2(n3334), .Z(n3193) );
  XOR2_X1 U55474 ( .A1(n52412), .A2(n4513), .Z(n65015) );
  BUF_X2 U55501 ( .I(n51030), .Z(n65016) );
  XOR2_X1 U55507 ( .A1(n65017), .A2(n58725), .Z(n7903) );
  XOR2_X1 U55512 ( .A1(n14228), .A2(n50770), .Z(n65017) );
  XOR2_X1 U55513 ( .A1(n3519), .A2(n3520), .Z(n6439) );
  XOR2_X1 U55520 ( .A1(n44919), .A2(n20854), .Z(n26181) );
  XOR2_X1 U55529 ( .A1(n44640), .A2(n46299), .Z(n44919) );
  XOR2_X1 U55538 ( .A1(n52333), .A2(n51792), .Z(n65018) );
  OR2_X2 U55552 ( .A1(n25867), .A2(n10719), .Z(n59523) );
  OAI22_X1 U55564 ( .A1(n58477), .A2(n51529), .B1(n60809), .B2(n61202), .ZN(
        n52694) );
  INV_X2 U55566 ( .I(n65019), .ZN(n57330) );
  NAND2_X1 U55567 ( .A1(n13522), .A2(n13524), .ZN(n65020) );
  NAND2_X1 U55579 ( .A1(n462), .A2(n41997), .ZN(n39175) );
  XOR2_X1 U55632 ( .A1(n17762), .A2(n46695), .Z(n8633) );
  XOR2_X1 U55638 ( .A1(n65023), .A2(n14889), .Z(n686) );
  XOR2_X1 U55641 ( .A1(n60778), .A2(n17466), .Z(n65023) );
  OAI21_X1 U55654 ( .A1(n24114), .A2(n61885), .B(n65024), .ZN(n41979) );
  NOR2_X1 U55655 ( .A1(n15276), .A2(n46716), .ZN(n15903) );
  XOR2_X1 U55657 ( .A1(n8449), .A2(n37724), .Z(n65025) );
  XOR2_X1 U55663 ( .A1(n17340), .A2(n45861), .Z(n25337) );
  NOR2_X2 U55669 ( .A1(n59409), .A2(n41874), .ZN(n41882) );
  OAI22_X1 U55692 ( .A1(n35337), .A2(n37065), .B1(n37068), .B2(n35336), .ZN(
        n35338) );
  OAI21_X1 U55701 ( .A1(n65026), .A2(n28642), .B(n29694), .ZN(n28643) );
  NOR2_X1 U55702 ( .A1(n3749), .A2(n15305), .ZN(n65026) );
  XOR2_X1 U55715 ( .A1(n43218), .A2(n55340), .Z(n1009) );
  NOR2_X2 U55726 ( .A1(n65029), .A2(n65028), .ZN(n21887) );
  NOR2_X2 U55728 ( .A1(n21888), .A2(n20782), .ZN(n65028) );
  NAND4_X2 U55731 ( .A1(n49271), .A2(n65031), .A3(n13783), .A4(n65030), .ZN(
        n50695) );
  NOR2_X2 U55738 ( .A1(n7383), .A2(n12556), .ZN(n65031) );
  INV_X2 U55749 ( .I(n30746), .ZN(n65032) );
  XOR2_X1 U55753 ( .A1(n65033), .A2(n51366), .Z(n25086) );
  XOR2_X1 U55756 ( .A1(n21685), .A2(n5778), .Z(n65033) );
  XOR2_X1 U55757 ( .A1(n60889), .A2(n6065), .Z(n208) );
  NAND4_X2 U55762 ( .A1(n47392), .A2(n47393), .A3(n47395), .A4(n47394), .ZN(
        n47444) );
  NAND2_X2 U55764 ( .A1(n16500), .A2(n65034), .ZN(n55441) );
  AND2_X1 U55768 ( .A1(n55323), .A2(n55442), .Z(n65034) );
  XOR2_X1 U55775 ( .A1(n65035), .A2(n5374), .Z(n36732) );
  XOR2_X1 U55786 ( .A1(n36686), .A2(n39498), .Z(n65035) );
  XOR2_X1 U55790 ( .A1(n24825), .A2(n18748), .Z(n8416) );
  XOR2_X1 U55803 ( .A1(n32242), .A2(n31629), .Z(n18748) );
  XOR2_X1 U55809 ( .A1(n11474), .A2(n38834), .Z(n928) );
  XOR2_X1 U55811 ( .A1(n39299), .A2(n2356), .Z(n11474) );
  NAND3_X2 U55823 ( .A1(n48618), .A2(n48627), .A3(n48616), .ZN(n25486) );
  NAND2_X1 U55824 ( .A1(n55282), .A2(n55283), .ZN(n59038) );
  NAND2_X2 U55827 ( .A1(n3864), .A2(n57211), .ZN(n65036) );
  BUF_X4 U55828 ( .I(n13838), .Z(n65062) );
  BUF_X2 U55831 ( .I(n28383), .Z(n65037) );
  AND2_X1 U55840 ( .A1(n29520), .A2(n15791), .Z(n65038) );
  NAND4_X1 U55848 ( .A1(n52892), .A2(n52883), .A3(n56989), .A4(n56987), .ZN(
        n52884) );
  NAND3_X2 U55850 ( .A1(n42788), .A2(n39087), .A3(n9792), .ZN(n42185) );
  NAND2_X2 U55856 ( .A1(n25807), .A2(n13704), .ZN(n27105) );
  XOR2_X1 U55867 ( .A1(n38070), .A2(n22036), .Z(n4779) );
  XOR2_X1 U55869 ( .A1(n37726), .A2(n24148), .Z(n38070) );
  XOR2_X1 U55870 ( .A1(n58240), .A2(n65040), .Z(n39507) );
  NOR2_X1 U55877 ( .A1(n10833), .A2(n52225), .ZN(n10832) );
  BUF_X2 U55891 ( .I(n31863), .Z(n65041) );
  NOR2_X2 U55905 ( .A1(n47186), .A2(n19361), .ZN(n20878) );
  NAND4_X2 U55925 ( .A1(n7858), .A2(n14973), .A3(n7859), .A4(n917), .ZN(n7857)
         );
  XOR2_X1 U55938 ( .A1(n65042), .A2(n24182), .Z(n51491) );
  XOR2_X1 U55939 ( .A1(n14593), .A2(n14594), .Z(n65042) );
  XOR2_X1 U55946 ( .A1(n65043), .A2(n893), .Z(n21294) );
  XOR2_X1 U55960 ( .A1(n25106), .A2(n8221), .Z(n65043) );
  INV_X1 U55963 ( .I(n11804), .ZN(n56361) );
  NOR2_X1 U55975 ( .A1(n18121), .A2(n25359), .ZN(n11804) );
  OAI21_X1 U55976 ( .A1(n63106), .A2(n8129), .B(n20864), .ZN(n65044) );
  XOR2_X1 U55977 ( .A1(n65045), .A2(n46696), .Z(n60572) );
  XOR2_X1 U55999 ( .A1(n65050), .A2(n54219), .Z(Plaintext[61]) );
  NAND4_X2 U56016 ( .A1(n54218), .A2(n54216), .A3(n54217), .A4(n54215), .ZN(
        n65050) );
  INV_X2 U56017 ( .I(n65051), .ZN(n8182) );
  XOR2_X1 U56018 ( .A1(n65053), .A2(n44896), .Z(n17521) );
  XOR2_X1 U56019 ( .A1(n44969), .A2(n13957), .Z(n65053) );
  XOR2_X1 U56026 ( .A1(n65054), .A2(n55535), .Z(Plaintext[115]) );
  NOR3_X1 U56030 ( .A1(n55533), .A2(n55532), .A3(n55531), .ZN(n65054) );
  NAND2_X2 U56047 ( .A1(n1592), .A2(n21273), .ZN(n55556) );
  NAND3_X2 U56060 ( .A1(n18816), .A2(n60577), .A3(n18815), .ZN(n7249) );
  INV_X2 U56063 ( .I(n17867), .ZN(n24256) );
  XOR2_X1 U56068 ( .A1(n10911), .A2(n65055), .Z(n17867) );
  NAND4_X1 U56070 ( .A1(n43466), .A2(n43465), .A3(n43463), .A4(n58530), .ZN(
        n43481) );
  NOR3_X1 U56095 ( .A1(n17434), .A2(n17437), .A3(n17432), .ZN(n17431) );
  XOR2_X1 U56100 ( .A1(n7703), .A2(n7702), .Z(n65214) );
  INV_X1 U56113 ( .I(n47444), .ZN(n49317) );
  NOR2_X2 U56114 ( .A1(n49496), .A2(n7738), .ZN(n23500) );
  INV_X2 U56119 ( .I(n48852), .ZN(n49496) );
  NAND2_X2 U56142 ( .A1(n60884), .A2(n21257), .ZN(n48852) );
  XOR2_X1 U56145 ( .A1(n1993), .A2(n1995), .Z(n11437) );
  NAND4_X2 U56146 ( .A1(n54530), .A2(n54582), .A3(n54560), .A4(n18425), .ZN(
        n25766) );
  XOR2_X1 U56148 ( .A1(n51584), .A2(n2516), .Z(n5141) );
  XOR2_X1 U56159 ( .A1(n26076), .A2(n31688), .Z(n26075) );
  XOR2_X1 U56184 ( .A1(n7362), .A2(n32516), .Z(n31688) );
  INV_X4 U56221 ( .I(n61601), .ZN(n1069) );
  NOR3_X1 U56254 ( .A1(n56482), .A2(n56510), .A3(n56456), .ZN(n56457) );
  NAND2_X2 U56283 ( .A1(n42804), .A2(n13389), .ZN(n42976) );
  XOR2_X1 U56285 ( .A1(n3104), .A2(n22883), .Z(n7442) );
  NAND3_X2 U56290 ( .A1(n4106), .A2(n1708), .A3(n25368), .ZN(n42158) );
  NOR2_X2 U56295 ( .A1(n4107), .A2(n63293), .ZN(n4106) );
  XOR2_X1 U56298 ( .A1(n38740), .A2(n65065), .Z(n13355) );
  XOR2_X1 U56301 ( .A1(n58926), .A2(n65066), .Z(n65065) );
  INV_X2 U56302 ( .I(n5779), .ZN(n65066) );
  INV_X2 U56309 ( .I(n65067), .ZN(n57400) );
  NOR2_X2 U56332 ( .A1(n46813), .A2(n15728), .ZN(n65067) );
  XOR2_X1 U56336 ( .A1(n65068), .A2(n19224), .Z(n51703) );
  XOR2_X1 U56340 ( .A1(n51850), .A2(n59053), .Z(n65068) );
  XOR2_X1 U56344 ( .A1(n65069), .A2(n23548), .Z(n14055) );
  OAI21_X1 U56349 ( .A1(n3672), .A2(n3966), .B(n3671), .ZN(n65069) );
  NOR2_X2 U56353 ( .A1(n65070), .A2(n20576), .ZN(n19377) );
  NAND2_X2 U56365 ( .A1(n25414), .A2(n21819), .ZN(n65070) );
  OAI21_X2 U56367 ( .A1(n28725), .A2(n30773), .B(n65071), .ZN(n28726) );
  AOI21_X2 U56376 ( .A1(n30771), .A2(n28723), .B(n29744), .ZN(n65071) );
  AOI22_X2 U56377 ( .A1(n65072), .A2(n50278), .B1(n57543), .B2(n50277), .ZN(
        n50280) );
  XOR2_X1 U56379 ( .A1(n57649), .A2(n2816), .Z(n58480) );
  NAND2_X2 U56384 ( .A1(n11078), .A2(n24610), .ZN(n65073) );
  XOR2_X1 U56417 ( .A1(n20471), .A2(n38649), .Z(n9605) );
  XOR2_X1 U56426 ( .A1(n60910), .A2(n9603), .Z(n9606) );
  XOR2_X1 U56431 ( .A1(n18902), .A2(n18903), .Z(n18901) );
  OR3_X1 U56432 ( .A1(n49774), .A2(n48947), .A3(n149), .Z(n57896) );
  NAND2_X2 U56435 ( .A1(n60285), .A2(n1546), .ZN(n35254) );
  NAND2_X1 U56447 ( .A1(n55411), .A2(n55410), .ZN(n20823) );
  NOR2_X2 U56449 ( .A1(n26752), .A2(n65076), .ZN(n29209) );
  XOR2_X1 U56453 ( .A1(n58301), .A2(n45861), .Z(n65077) );
  XOR2_X1 U56465 ( .A1(n8230), .A2(n57187), .Z(n45862) );
  NOR2_X2 U56525 ( .A1(n44075), .A2(n44076), .ZN(n65222) );
  XOR2_X1 U56527 ( .A1(n65078), .A2(n2086), .Z(n2083) );
  XOR2_X1 U56537 ( .A1(n51521), .A2(n5351), .Z(n5350) );
  BUF_X2 U56540 ( .I(n55810), .Z(n65079) );
  AOI21_X2 U56542 ( .A1(n48034), .A2(n48033), .B(n65080), .ZN(n48045) );
  XOR2_X1 U56544 ( .A1(n44269), .A2(n12377), .Z(n6097) );
  OR2_X1 U56546 ( .A1(n40303), .A2(n40304), .Z(n22346) );
  OR2_X1 U56551 ( .A1(n24701), .A2(n3177), .Z(n28008) );
  INV_X2 U56566 ( .I(n40744), .ZN(n41240) );
  NAND2_X2 U56569 ( .A1(n61013), .A2(n15548), .ZN(n40744) );
  BUF_X2 U56578 ( .I(n45281), .Z(n65082) );
  XOR2_X1 U56581 ( .A1(n58751), .A2(n185), .Z(n25315) );
  XOR2_X1 U56582 ( .A1(n65083), .A2(n18963), .Z(n9762) );
  XOR2_X1 U56589 ( .A1(n877), .A2(n18960), .Z(n65083) );
  XOR2_X1 U56590 ( .A1(n13270), .A2(n307), .Z(n8908) );
  XOR2_X1 U56591 ( .A1(n58254), .A2(n22), .Z(n23481) );
  XOR2_X1 U56593 ( .A1(n65087), .A2(n58618), .Z(n60241) );
  XOR2_X1 U56600 ( .A1(n14735), .A2(n6096), .Z(n65087) );
  XOR2_X1 U56601 ( .A1(n21580), .A2(n3036), .Z(n3035) );
  NAND2_X2 U56603 ( .A1(n16108), .A2(n35492), .ZN(n12493) );
  NOR2_X2 U56604 ( .A1(n36442), .A2(n7705), .ZN(n36452) );
  XOR2_X1 U56605 ( .A1(n65090), .A2(n32308), .Z(n21725) );
  XOR2_X1 U56614 ( .A1(n32229), .A2(n18732), .Z(n65090) );
  XOR2_X1 U56615 ( .A1(n65091), .A2(n14737), .Z(n3838) );
  NAND2_X2 U56619 ( .A1(n57310), .A2(n65092), .ZN(n52340) );
  NOR2_X2 U56631 ( .A1(n49855), .A2(n26108), .ZN(n65092) );
  NAND3_X2 U56634 ( .A1(n65093), .A2(n14009), .A3(n14008), .ZN(n14010) );
  XOR2_X1 U56664 ( .A1(n32498), .A2(n19250), .Z(n15611) );
  XOR2_X1 U56689 ( .A1(n7306), .A2(n65094), .Z(n18039) );
  XOR2_X1 U56694 ( .A1(n49938), .A2(n57660), .Z(n59752) );
  XOR2_X1 U56698 ( .A1(n25257), .A2(n7711), .Z(n49938) );
  NAND2_X2 U56717 ( .A1(n18119), .A2(n12058), .ZN(n9410) );
  BUF_X2 U56721 ( .I(n47292), .Z(n65095) );
  NAND2_X2 U56735 ( .A1(n9650), .A2(n54477), .ZN(n54546) );
  XOR2_X1 U56737 ( .A1(n65097), .A2(n49571), .Z(n49625) );
  XOR2_X1 U56743 ( .A1(n4085), .A2(n51592), .Z(n65097) );
  AOI22_X2 U56744 ( .A1(n18876), .A2(n50235), .B1(n50242), .B2(n60622), .ZN(
        n21634) );
  NOR3_X2 U56745 ( .A1(n61487), .A2(n25589), .A3(n61488), .ZN(n18876) );
  AOI21_X2 U56748 ( .A1(n35042), .A2(n35041), .B(n65098), .ZN(n35051) );
  OAI22_X2 U56749 ( .A1(n5186), .A2(n5478), .B1(n35039), .B2(n35038), .ZN(
        n65098) );
  NOR2_X1 U56751 ( .A1(n58594), .A2(n35441), .ZN(n424) );
  XOR2_X1 U56752 ( .A1(n37966), .A2(n65099), .Z(n10709) );
  XOR2_X1 U56757 ( .A1(n25021), .A2(n935), .Z(n65099) );
  XOR2_X1 U56759 ( .A1(n7019), .A2(n17219), .Z(n9737) );
  NAND2_X2 U56765 ( .A1(n34392), .A2(n34402), .ZN(n35228) );
  INV_X4 U56770 ( .I(n59005), .ZN(n35655) );
  XOR2_X1 U56771 ( .A1(n33159), .A2(n65102), .Z(n7708) );
  XOR2_X1 U56772 ( .A1(n33155), .A2(n33157), .Z(n65102) );
  OR3_X1 U56777 ( .A1(n60826), .A2(n41914), .A3(n64768), .Z(n37902) );
  XOR2_X1 U56780 ( .A1(n33264), .A2(n33263), .Z(n33276) );
  XOR2_X1 U56784 ( .A1(n65219), .A2(n21586), .Z(n33264) );
  NAND3_X2 U56792 ( .A1(n31128), .A2(n31127), .A3(n61426), .ZN(n27153) );
  NAND2_X2 U56796 ( .A1(n24265), .A2(n53851), .ZN(n53889) );
  AOI22_X1 U56799 ( .A1(n17901), .A2(n17899), .B1(n49977), .B2(n49976), .ZN(
        n49983) );
  XOR2_X1 U56800 ( .A1(n50203), .A2(n16376), .Z(n65104) );
  NOR4_X2 U56804 ( .A1(n65107), .A2(n53153), .A3(n53150), .A4(n65106), .ZN(
        n53156) );
  NAND2_X1 U56817 ( .A1(n53228), .A2(n9765), .ZN(n65108) );
  OR2_X1 U56822 ( .A1(n36567), .A2(n23215), .Z(n36380) );
  NOR2_X1 U56829 ( .A1(n3338), .A2(n65109), .ZN(n61079) );
  NAND3_X2 U56831 ( .A1(n14170), .A2(n4695), .A3(n14166), .ZN(n49363) );
  XOR2_X1 U56832 ( .A1(n24536), .A2(n60499), .Z(n57534) );
  INV_X2 U56833 ( .I(n23237), .ZN(n29819) );
  XOR2_X1 U56834 ( .A1(n12377), .A2(n46318), .Z(n18903) );
  XOR2_X1 U56835 ( .A1(n38972), .A2(n39543), .Z(n8989) );
  OAI22_X1 U56836 ( .A1(n52909), .A2(n55401), .B1(n52910), .B2(n55244), .ZN(
        n52912) );
  NOR2_X2 U56838 ( .A1(n55400), .A2(n55397), .ZN(n55244) );
  BUF_X2 U56839 ( .I(n18248), .Z(n65112) );
  XOR2_X1 U56842 ( .A1(n65113), .A2(n55242), .Z(Plaintext[107]) );
  NAND4_X2 U56843 ( .A1(n55241), .A2(n55240), .A3(n55239), .A4(n55238), .ZN(
        n65113) );
  OR2_X1 U56851 ( .A1(n47150), .A2(n50448), .Z(n65114) );
  XOR2_X1 U56855 ( .A1(n8833), .A2(n18125), .Z(n7192) );
  NOR2_X2 U56860 ( .A1(n17467), .A2(n42835), .ZN(n65115) );
  NOR3_X2 U56862 ( .A1(n40815), .A2(n65116), .A3(n57387), .ZN(n40824) );
  NAND3_X2 U56863 ( .A1(n51256), .A2(n56432), .A3(n51257), .ZN(n65117) );
  NAND2_X2 U56867 ( .A1(n18423), .A2(n23745), .ZN(n28278) );
  OR2_X1 U56874 ( .A1(n30286), .A2(n14389), .Z(n9167) );
  XOR2_X1 U56879 ( .A1(n57854), .A2(n65118), .Z(n59270) );
  XOR2_X1 U56880 ( .A1(n7937), .A2(n13486), .Z(n65118) );
  INV_X2 U56881 ( .I(n2721), .ZN(n65119) );
  NAND2_X2 U56884 ( .A1(n10086), .A2(n36547), .ZN(n36549) );
  NAND3_X1 U56891 ( .A1(n28727), .A2(n29461), .A3(n65120), .ZN(n16085) );
  OR2_X1 U56896 ( .A1(n30725), .A2(n9426), .Z(n9168) );
  XOR2_X1 U56897 ( .A1(n31674), .A2(n19282), .Z(n59206) );
  XOR2_X1 U56903 ( .A1(n1831), .A2(n60259), .Z(n31674) );
  AOI21_X1 U56905 ( .A1(n38690), .A2(n64858), .B(n65123), .ZN(n24376) );
  NAND2_X1 U56911 ( .A1(n12922), .A2(n38677), .ZN(n65123) );
  INV_X2 U56912 ( .I(n48977), .ZN(n7912) );
  INV_X1 U56914 ( .I(n5944), .ZN(n65125) );
  NAND2_X2 U56918 ( .A1(n3376), .A2(n25213), .ZN(n5944) );
  OAI21_X1 U56929 ( .A1(n53241), .A2(n62515), .B(n21453), .ZN(n25487) );
  NAND2_X2 U56930 ( .A1(n1614), .A2(n1325), .ZN(n21453) );
  NAND2_X2 U56932 ( .A1(n11578), .A2(n65126), .ZN(n26135) );
  INV_X2 U56933 ( .I(n53163), .ZN(n65126) );
  XOR2_X1 U56936 ( .A1(n5349), .A2(n20430), .Z(n4960) );
  XOR2_X1 U56941 ( .A1(n9945), .A2(n61319), .Z(n16930) );
  BUF_X2 U56943 ( .I(n26020), .Z(n65129) );
  XOR2_X1 U56945 ( .A1(n17232), .A2(n31288), .Z(n17908) );
  XOR2_X1 U56947 ( .A1(n15647), .A2(n8719), .Z(n9148) );
  XOR2_X1 U56949 ( .A1(n65130), .A2(n52317), .Z(Plaintext[121]) );
  NAND2_X2 U56950 ( .A1(n44791), .A2(n48917), .ZN(n48929) );
  NOR2_X2 U56959 ( .A1(n57658), .A2(n65131), .ZN(n58537) );
  NOR3_X2 U56965 ( .A1(n5937), .A2(n59602), .A3(n20992), .ZN(n36951) );
  NOR2_X2 U56966 ( .A1(n27620), .A2(n11225), .ZN(n27166) );
  NOR2_X2 U56967 ( .A1(n52756), .A2(n53383), .ZN(n52844) );
  NAND2_X1 U56969 ( .A1(n17917), .A2(n17916), .ZN(n58995) );
  INV_X1 U56982 ( .I(n45319), .ZN(n46522) );
  NAND4_X2 U56989 ( .A1(n4329), .A2(n4327), .A3(n4331), .A4(n4333), .ZN(n45319) );
  NAND3_X2 U56990 ( .A1(n65132), .A2(n59003), .A3(n52876), .ZN(n53056) );
  NOR2_X2 U56996 ( .A1(n65133), .A2(n47790), .ZN(n47792) );
  NOR4_X2 U56997 ( .A1(n10933), .A2(n65134), .A3(n25730), .A4(n10932), .ZN(
        n9938) );
  XOR2_X1 U56998 ( .A1(n65136), .A2(n55840), .Z(Plaintext[132]) );
  NOR2_X1 U56999 ( .A1(n65137), .A2(n15769), .ZN(n17778) );
  NAND2_X1 U57000 ( .A1(n14133), .A2(n14135), .ZN(n65137) );
  NOR2_X1 U57001 ( .A1(n29503), .A2(n59658), .ZN(n65139) );
  OAI22_X1 U57009 ( .A1(n9830), .A2(n65140), .B1(n37327), .B2(n37187), .ZN(
        n34881) );
  BUF_X2 U57010 ( .I(n11883), .Z(n65141) );
  XOR2_X1 U57012 ( .A1(n65142), .A2(n14424), .Z(n10476) );
  INV_X2 U57017 ( .I(n49435), .ZN(n65142) );
  XOR2_X1 U57021 ( .A1(n59402), .A2(n23683), .Z(n31581) );
  INV_X2 U57025 ( .I(n62514), .ZN(n25671) );
  NAND2_X2 U57026 ( .A1(n22157), .A2(n48897), .ZN(n49699) );
  AOI21_X1 U57035 ( .A1(n48734), .A2(n48735), .B(n48733), .ZN(n22690) );
  NOR2_X2 U57036 ( .A1(n23474), .A2(n27486), .ZN(n27542) );
  XOR2_X1 U57037 ( .A1(n65146), .A2(n44511), .Z(n59222) );
  XOR2_X1 U57039 ( .A1(n44371), .A2(n46307), .Z(n44511) );
  NAND3_X2 U57040 ( .A1(n55382), .A2(n9777), .A3(n15703), .ZN(n19797) );
  INV_X2 U57041 ( .I(n2693), .ZN(n12615) );
  NAND2_X2 U57042 ( .A1(n40850), .A2(n41082), .ZN(n2693) );
  OAI21_X1 U57044 ( .A1(n32929), .A2(n32930), .B(n34247), .ZN(n32939) );
  XOR2_X1 U57048 ( .A1(n65148), .A2(n46160), .Z(n2404) );
  XOR2_X1 U57049 ( .A1(n4142), .A2(n46149), .Z(n65148) );
  XOR2_X1 U57059 ( .A1(n17815), .A2(n64039), .Z(n46347) );
  NAND3_X2 U57062 ( .A1(n23794), .A2(n26845), .A3(n26846), .ZN(n61374) );
  NOR2_X2 U57070 ( .A1(n26919), .A2(n19465), .ZN(n23794) );
  NAND2_X1 U57073 ( .A1(n58908), .A2(n54489), .ZN(n65149) );
  INV_X2 U57074 ( .I(n2814), .ZN(n65150) );
  INV_X1 U57075 ( .I(n26843), .ZN(n27925) );
  NAND2_X1 U57078 ( .A1(n57790), .A2(n24987), .ZN(n26843) );
  XOR2_X1 U57083 ( .A1(n13225), .A2(n62998), .Z(n59977) );
  XOR2_X1 U57084 ( .A1(n3190), .A2(n52413), .Z(n65151) );
  XOR2_X1 U57088 ( .A1(n65152), .A2(n32090), .Z(n32092) );
  XOR2_X1 U57089 ( .A1(n65153), .A2(n13285), .Z(n50750) );
  XOR2_X1 U57091 ( .A1(n23375), .A2(n16984), .Z(n65153) );
  NOR2_X2 U57094 ( .A1(n65154), .A2(n42521), .ZN(n57812) );
  BUF_X2 U57096 ( .I(n54349), .Z(n65155) );
  XOR2_X1 U57097 ( .A1(n38099), .A2(n38100), .Z(n38103) );
  NOR3_X2 U57098 ( .A1(n61331), .A2(n61332), .A3(n45543), .ZN(n21320) );
  XOR2_X1 U57099 ( .A1(n19067), .A2(n65156), .Z(n26110) );
  XOR2_X1 U57107 ( .A1(n38525), .A2(n20318), .Z(n65156) );
  NAND2_X1 U57108 ( .A1(n19835), .A2(n53375), .ZN(n65157) );
  NAND2_X2 U57115 ( .A1(n27888), .A2(n1566), .ZN(n28190) );
  XOR2_X1 U57117 ( .A1(n19126), .A2(n26911), .Z(n27888) );
  NAND2_X2 U57118 ( .A1(n20096), .A2(n65158), .ZN(n24056) );
  NOR3_X2 U57121 ( .A1(n20099), .A2(n20098), .A3(n26910), .ZN(n65158) );
  OR2_X2 U57123 ( .A1(n25427), .A2(n5251), .Z(n14330) );
  XOR2_X1 U57125 ( .A1(n13532), .A2(n22266), .Z(n37724) );
  OAI21_X1 U57126 ( .A1(n28030), .A2(n18224), .B(n6222), .ZN(n23498) );
  NOR2_X2 U57127 ( .A1(n33022), .A2(n36539), .ZN(n36536) );
  NAND3_X2 U57129 ( .A1(n58785), .A2(n33021), .A3(n35683), .ZN(n36539) );
  INV_X2 U57132 ( .I(n65159), .ZN(n57436) );
  NOR2_X2 U57140 ( .A1(n30197), .A2(n64950), .ZN(n65159) );
  XOR2_X1 U57149 ( .A1(n8105), .A2(n61958), .Z(n24392) );
  INV_X2 U57151 ( .I(n17617), .ZN(n13962) );
  NAND2_X2 U57152 ( .A1(n67), .A2(n17783), .ZN(n17617) );
  AOI21_X2 U57155 ( .A1(n57949), .A2(n8604), .B(n49395), .ZN(n2889) );
  XOR2_X1 U57163 ( .A1(n65162), .A2(n20113), .Z(n2948) );
  XOR2_X1 U57173 ( .A1(n45366), .A2(n10606), .Z(n65162) );
  INV_X2 U57181 ( .I(n36465), .ZN(n25842) );
  NAND2_X2 U57199 ( .A1(n2362), .A2(n11413), .ZN(n36465) );
  INV_X1 U57208 ( .I(n16458), .ZN(n65164) );
  XOR2_X1 U57209 ( .A1(n10325), .A2(n65165), .Z(n30209) );
  XOR2_X1 U57211 ( .A1(n2952), .A2(n30207), .Z(n65165) );
  NAND2_X2 U57215 ( .A1(n38922), .A2(n40770), .ZN(n61094) );
  NAND2_X2 U57220 ( .A1(n18738), .A2(n18739), .ZN(n7405) );
  NOR2_X2 U57221 ( .A1(n29916), .A2(n25096), .ZN(n28952) );
  NAND2_X1 U57222 ( .A1(n55090), .A2(n65166), .ZN(n23307) );
  NAND3_X1 U57223 ( .A1(n15519), .A2(n55089), .A3(n15520), .ZN(n65166) );
  NOR2_X1 U57224 ( .A1(n3371), .A2(n3372), .ZN(n3370) );
  NAND2_X1 U57225 ( .A1(n53881), .A2(n25127), .ZN(n20610) );
  NAND2_X2 U57226 ( .A1(n53035), .A2(n54025), .ZN(n53881) );
  AND2_X1 U57227 ( .A1(n57119), .A2(n18802), .Z(n65169) );
  NOR2_X2 U57228 ( .A1(n23191), .A2(n23942), .ZN(n22115) );
  NOR4_X2 U57229 ( .A1(n26326), .A2(n15904), .A3(n22932), .A4(n26325), .ZN(
        n11245) );
  XOR2_X1 U57230 ( .A1(n14059), .A2(n14061), .Z(n45046) );
  NOR2_X1 U57231 ( .A1(n26959), .A2(n26960), .ZN(n27218) );
  NAND3_X2 U57232 ( .A1(n5386), .A2(n18277), .A3(n5389), .ZN(n33710) );
  XOR2_X1 U57233 ( .A1(n8157), .A2(n8159), .Z(n59648) );
  XOR2_X1 U57234 ( .A1(n31629), .A2(n20403), .Z(n32244) );
  NOR2_X2 U57235 ( .A1(n2874), .A2(n2872), .ZN(n31629) );
  XOR2_X1 U57236 ( .A1(n65172), .A2(n23204), .Z(n59863) );
  NOR2_X1 U57237 ( .A1(n65173), .A2(n59940), .ZN(n7754) );
  XOR2_X1 U57238 ( .A1(n16458), .A2(n1449), .Z(n33155) );
  NAND2_X2 U57239 ( .A1(n2589), .A2(n4969), .ZN(n2590) );
  NOR2_X2 U57240 ( .A1(n60297), .A2(n1769), .ZN(n2589) );
  XOR2_X1 U57241 ( .A1(n1998), .A2(n1999), .Z(n52441) );
  NOR2_X2 U57242 ( .A1(n58250), .A2(n37224), .ZN(n3171) );
  NOR2_X2 U57243 ( .A1(n40944), .A2(n22593), .ZN(n18032) );
  AOI22_X2 U57244 ( .A1(n57452), .A2(n18115), .B1(n16849), .B2(n18072), .ZN(
        n38159) );
  XOR2_X1 U57245 ( .A1(n65176), .A2(n18971), .Z(n7851) );
  XOR2_X1 U57246 ( .A1(n4395), .A2(n18972), .Z(n65176) );
  XOR2_X1 U57247 ( .A1(n15308), .A2(n23330), .Z(n7575) );
  BUF_X2 U57248 ( .I(n44893), .Z(n65177) );
  NAND2_X2 U57249 ( .A1(n40106), .A2(n65180), .ZN(n40341) );
  AND2_X1 U57250 ( .A1(n38022), .A2(n19611), .Z(n65180) );
  AOI22_X2 U57251 ( .A1(n50367), .A2(n260), .B1(n49476), .B2(n49989), .ZN(
        n49477) );
  NAND2_X2 U57252 ( .A1(n3807), .A2(n3808), .ZN(n13802) );
  BUF_X2 U57253 ( .I(n42825), .Z(n65181) );
  XOR2_X1 U57254 ( .A1(n60731), .A2(n65182), .Z(n2043) );
  XOR2_X1 U57255 ( .A1(n5489), .A2(n32617), .Z(n65182) );
  NOR3_X2 U57256 ( .A1(n58929), .A2(n58019), .A3(n28686), .ZN(n14546) );
  NAND2_X2 U57257 ( .A1(n15181), .A2(n34721), .ZN(n15183) );
  NAND2_X1 U57258 ( .A1(n26588), .A2(n26589), .ZN(n26591) );
  BUF_X2 U57259 ( .I(n9562), .Z(n65183) );
  BUF_X2 U57260 ( .I(n41212), .Z(n65184) );
  BUF_X2 U57261 ( .I(n42676), .Z(n65185) );
  INV_X2 U57262 ( .I(n65186), .ZN(n57424) );
  NAND2_X2 U57263 ( .A1(n26126), .A2(n26192), .ZN(n65186) );
  XOR2_X1 U57264 ( .A1(n12685), .A2(n32371), .Z(n12080) );
  NAND3_X2 U57265 ( .A1(n65190), .A2(n30495), .A3(n30494), .ZN(n11159) );
  XOR2_X1 U57266 ( .A1(n46430), .A2(n44507), .Z(n44155) );
  NAND2_X2 U57267 ( .A1(n42765), .A2(n25398), .ZN(n46430) );
  NAND4_X2 U57268 ( .A1(n34400), .A2(n34397), .A3(n34399), .A4(n34398), .ZN(
        n58156) );
  XOR2_X1 U57269 ( .A1(n6031), .A2(n65191), .Z(n17584) );
  XOR2_X1 U57270 ( .A1(n17586), .A2(n25250), .Z(n65191) );
  NAND2_X2 U57271 ( .A1(n19638), .A2(n18473), .ZN(n18242) );
  NOR2_X2 U57272 ( .A1(n16459), .A2(n65192), .ZN(n8938) );
  NAND2_X2 U57273 ( .A1(n8940), .A2(n16204), .ZN(n65192) );
  INV_X2 U57274 ( .I(n30486), .ZN(n27756) );
  NAND2_X2 U57275 ( .A1(n16791), .A2(n16789), .ZN(n30486) );
  NOR2_X2 U57276 ( .A1(n43733), .A2(n15007), .ZN(n43210) );
  NAND2_X2 U57277 ( .A1(n5490), .A2(n65193), .ZN(n31984) );
  NAND2_X2 U57278 ( .A1(n11197), .A2(n40448), .ZN(n43376) );
  NAND3_X2 U57279 ( .A1(n6880), .A2(n6878), .A3(n6876), .ZN(n11197) );
  XOR2_X1 U57280 ( .A1(n51364), .A2(n51369), .Z(n22101) );
  XOR2_X1 U57281 ( .A1(n50611), .A2(n22102), .Z(n51369) );
  XOR2_X1 U57282 ( .A1(n11847), .A2(n65195), .Z(n11846) );
  BUF_X2 U57283 ( .I(n18138), .Z(n65196) );
  XOR2_X1 U57284 ( .A1(n2576), .A2(n1752), .Z(n12177) );
  NOR2_X2 U57285 ( .A1(n29152), .A2(n21720), .ZN(n27392) );
  INV_X4 U57286 ( .I(n58748), .ZN(n36139) );
  NAND3_X2 U57287 ( .A1(n41932), .A2(n41931), .A3(n41930), .ZN(n57935) );
  XOR2_X1 U57288 ( .A1(n65201), .A2(n51792), .Z(n3402) );
  XOR2_X1 U57289 ( .A1(n51790), .A2(n51789), .Z(n65201) );
  OAI21_X1 U57290 ( .A1(n13496), .A2(n13498), .B(n47420), .ZN(n24952) );
  XOR2_X1 U57291 ( .A1(n24152), .A2(n32084), .Z(n22066) );
  BUF_X2 U57292 ( .I(n40938), .Z(n65206) );
  XOR2_X1 U57293 ( .A1(n65207), .A2(n25804), .Z(n17737) );
  XOR2_X1 U57294 ( .A1(n17739), .A2(n23069), .Z(n65207) );
  NAND3_X2 U57295 ( .A1(n43412), .A2(n43548), .A3(n62997), .ZN(n43559) );
  OR2_X2 U57296 ( .A1(n35427), .A2(n36953), .Z(n36939) );
  BUF_X2 U57297 ( .I(n22842), .Z(n65208) );
  XOR2_X1 U57298 ( .A1(n52419), .A2(n17738), .Z(n51434) );
  NAND2_X1 U57299 ( .A1(n65209), .A2(n17006), .ZN(n16837) );
  OAI21_X1 U57300 ( .A1(n46996), .A2(n46258), .B(n20788), .ZN(n65209) );
  AOI21_X2 U57301 ( .A1(n65211), .A2(n57419), .B(n44410), .ZN(n15467) );
  XOR2_X1 U57302 ( .A1(n17441), .A2(n65212), .Z(n17439) );
  XOR2_X1 U57303 ( .A1(n45343), .A2(n65213), .Z(n5533) );
  XOR2_X1 U57304 ( .A1(n657), .A2(n19691), .Z(n4958) );
  XOR2_X1 U57305 ( .A1(n52066), .A2(n3187), .Z(n19691) );
  XOR2_X1 U57306 ( .A1(n9587), .A2(n9586), .Z(n9607) );
  NOR2_X2 U57307 ( .A1(n9608), .A2(n63586), .ZN(n58702) );
  NAND2_X1 U57308 ( .A1(n33642), .A2(n33538), .ZN(n20092) );
  NOR2_X1 U57309 ( .A1(n19822), .A2(n19826), .ZN(n31777) );
  NOR2_X2 U57310 ( .A1(n1863), .A2(n61383), .ZN(n30681) );
  OR2_X1 U57311 ( .A1(n33630), .A2(n33224), .Z(n20582) );
  XOR2_X1 U57312 ( .A1(n59765), .A2(n59377), .Z(n58385) );
  NAND2_X2 U57313 ( .A1(n59409), .A2(n58587), .ZN(n65218) );
  NOR2_X2 U57314 ( .A1(n60509), .A2(n40578), .ZN(n10500) );
  XOR2_X1 U57315 ( .A1(n65220), .A2(n4933), .Z(n12349) );
  XOR2_X1 U57316 ( .A1(n58715), .A2(n14337), .Z(n65220) );
  XOR2_X1 U57317 ( .A1(n65221), .A2(n26690), .Z(n26692) );
  XOR2_X1 U57318 ( .A1(n55810), .A2(n22691), .Z(n65221) );
  NAND3_X2 U57319 ( .A1(n22395), .A2(n58299), .A3(n44657), .ZN(n44658) );
  XOR2_X1 U57320 ( .A1(n59619), .A2(n59620), .Z(n5574) );
  XOR2_X1 U57321 ( .A1(n12634), .A2(n11213), .Z(n59306) );
  NAND2_X1 U57322 ( .A1(n30944), .A2(n25659), .ZN(n22082) );
  NAND2_X2 U57323 ( .A1(n653), .A2(n1805), .ZN(n65225) );
  XOR2_X1 U57324 ( .A1(n37834), .A2(n61650), .Z(n65227) );
  XOR2_X1 U57325 ( .A1(n38621), .A2(n25249), .Z(n58145) );
  OR2_X1 U57326 ( .A1(n62353), .A2(n7187), .Z(n59150) );
  XNOR2_X1 U57327 ( .A1(n22111), .A2(n46598), .ZN(n46519) );
  XOR2_X1 U57328 ( .A1(n65229), .A2(n39497), .Z(n58113) );
  XOR2_X1 U57329 ( .A1(n39496), .A2(n39495), .Z(n65229) );
  NAND4_X1 U57330 ( .A1(n27218), .A2(n26961), .A3(n5206), .A4(n1882), .ZN(n133) );
  BUF_X2 U57331 ( .I(n60930), .Z(n65230) );
  NAND2_X2 U57332 ( .A1(n29511), .A2(n3908), .ZN(n29002) );
  XOR2_X1 U57333 ( .A1(n65231), .A2(n37072), .Z(n6578) );
  XOR2_X1 U57334 ( .A1(n6437), .A2(n36157), .Z(n65231) );
  XOR2_X1 U57335 ( .A1(n32230), .A2(n60887), .Z(n23246) );
  BUF_X2 U57336 ( .I(n16750), .Z(n65233) );
  NAND2_X2 U57337 ( .A1(n61728), .A2(n2810), .ZN(n6323) );
  OAI21_X2 U57338 ( .A1(n7933), .A2(n1217), .B(n36465), .ZN(n10790) );
  AND2_X1 U57339 ( .A1(n28964), .A2(n29900), .Z(n65235) );
  BUF_X2 U57340 ( .I(n22223), .Z(n65236) );
  XOR2_X1 U57341 ( .A1(n8038), .A2(n14259), .Z(n65237) );
  XOR2_X1 U57342 ( .A1(n22476), .A2(n44263), .Z(n33881) );
  AOI22_X1 U57343 ( .A1(n21248), .A2(n5277), .B1(n5570), .B2(n55275), .ZN(
        n7583) );
  NAND2_X1 U57344 ( .A1(n40112), .A2(n40111), .ZN(n65238) );
  XOR2_X1 U57345 ( .A1(n59932), .A2(n5728), .Z(n65239) );
  XOR2_X1 U57346 ( .A1(n31290), .A2(n31289), .Z(n57869) );
  XOR2_X1 U57347 ( .A1(n25315), .A2(n15079), .Z(n10867) );
  OAI21_X1 U57348 ( .A1(n56462), .A2(n56461), .B(n56502), .ZN(n56469) );
  OR2_X1 U57349 ( .A1(n61194), .A2(n42107), .Z(n65240) );
  XOR2_X1 U57350 ( .A1(n18639), .A2(n50631), .Z(n13289) );
  XOR2_X1 U57351 ( .A1(n39368), .A2(n9120), .Z(n65241) );
  NAND3_X2 U57352 ( .A1(n24503), .A2(n28572), .A3(n65242), .ZN(n28578) );
  NAND4_X1 U57353 ( .A1(n22411), .A2(n28571), .A3(n5267), .A4(n31083), .ZN(
        n65242) );
  NOR2_X2 U57354 ( .A1(n23724), .A2(n65243), .ZN(n23723) );
  NAND3_X2 U57355 ( .A1(n28545), .A2(n61440), .A3(n61439), .ZN(n65243) );
  NAND3_X2 U57356 ( .A1(n27153), .A2(n31131), .A3(n27152), .ZN(n358) );
  AOI21_X1 U57357 ( .A1(n36389), .A2(n36390), .B(n65244), .ZN(n36399) );
  NAND3_X2 U57358 ( .A1(n30154), .A2(n30156), .A3(n30155), .ZN(n25174) );
  AND2_X2 U57359 ( .A1(n20975), .A2(n23286), .Z(n26347) );
  XOR2_X1 U57360 ( .A1(Ciphertext[31]), .A2(Key[110]), .Z(n23286) );
  XOR2_X1 U57361 ( .A1(n44224), .A2(n45047), .Z(n45151) );
  BUF_X2 U57362 ( .I(n59838), .Z(n65245) );
  XOR2_X1 U57363 ( .A1(n60227), .A2(n15734), .Z(n44523) );
  XOR2_X1 U57364 ( .A1(n17233), .A2(n14299), .Z(n61606) );
  XOR2_X1 U57365 ( .A1(n52373), .A2(n17085), .Z(n17233) );
  OR2_X1 U57366 ( .A1(n16974), .A2(n21755), .Z(n44570) );
  NOR3_X2 U57367 ( .A1(n57409), .A2(n19746), .A3(n14843), .ZN(n59389) );
  XOR2_X1 U57368 ( .A1(n15385), .A2(n65247), .Z(n23475) );
  XOR2_X1 U57369 ( .A1(n50371), .A2(n65248), .Z(n65247) );
  XOR2_X1 U57370 ( .A1(n43649), .A2(n22291), .Z(n26166) );
  OR2_X1 U57371 ( .A1(n33610), .A2(n32460), .Z(n7317) );
  NAND2_X2 U57372 ( .A1(n32782), .A2(n64417), .ZN(n33610) );
  XOR2_X1 U57373 ( .A1(n65250), .A2(n46120), .Z(n24201) );
  XOR2_X1 U57374 ( .A1(n5214), .A2(n46288), .Z(n46120) );
  NAND2_X2 U57375 ( .A1(n6841), .A2(n473), .ZN(n6839) );
  NOR2_X2 U57376 ( .A1(n56600), .A2(n24647), .ZN(n52890) );
  XOR2_X1 U57377 ( .A1(n17060), .A2(n48402), .Z(n65251) );
  OAI21_X2 U57378 ( .A1(n49098), .A2(n49099), .B(n49097), .ZN(n65252) );
  XOR2_X1 U57379 ( .A1(n44923), .A2(n791), .Z(n60576) );
  XOR2_X1 U57380 ( .A1(n44460), .A2(n6677), .Z(n44923) );
  INV_X2 U57381 ( .I(n65253), .ZN(n57473) );
  XOR2_X1 U57382 ( .A1(n65255), .A2(n65254), .Z(n31508) );
  XOR2_X1 U57383 ( .A1(n31499), .A2(n31498), .Z(n65255) );
  XOR2_X1 U57384 ( .A1(n65257), .A2(n51722), .Z(n50111) );
  XOR2_X1 U57385 ( .A1(n5724), .A2(n24205), .Z(n65257) );
  XOR2_X1 U57386 ( .A1(n65258), .A2(n61506), .Z(n39268) );
  XOR2_X1 U57387 ( .A1(n15704), .A2(n39265), .Z(n65258) );
  XOR2_X1 U57388 ( .A1(n1676), .A2(n41772), .Z(n44268) );
  NAND2_X1 U57389 ( .A1(n56536), .A2(n65260), .ZN(n56537) );
  NAND3_X1 U57390 ( .A1(n56533), .A2(n56532), .A3(n56534), .ZN(n65260) );
  NOR2_X2 U57391 ( .A1(n20985), .A2(n22401), .ZN(n54400) );
  AND2_X1 U57392 ( .A1(n43508), .A2(n43507), .Z(n15834) );
  NOR2_X2 U57393 ( .A1(n19000), .A2(n61442), .ZN(n43508) );
  NAND2_X2 U57394 ( .A1(n65263), .A2(n18660), .ZN(n18662) );
  NAND2_X1 U57395 ( .A1(n18659), .A2(n18658), .ZN(n65263) );
  INV_X2 U57396 ( .I(n65264), .ZN(n10635) );
  NAND2_X1 U57397 ( .A1(n41983), .A2(n12925), .ZN(n65265) );
  XOR2_X1 U57398 ( .A1(n65266), .A2(n52532), .Z(n25085) );
  XOR2_X1 U57399 ( .A1(n25086), .A2(n22310), .Z(n65266) );
  XOR2_X1 U57400 ( .A1(n65267), .A2(n6040), .Z(n5755) );
  INV_X2 U57401 ( .I(n15844), .ZN(n65267) );
  INV_X1 U57402 ( .I(n22128), .ZN(n33963) );
  INV_X2 U57403 ( .I(n59272), .ZN(n22128) );
  INV_X4 U57404 ( .I(n7253), .ZN(n33144) );
  XNOR2_X1 U57405 ( .A1(n33069), .A2(n15912), .ZN(n65268) );
  INV_X2 U57406 ( .I(n14733), .ZN(n12413) );
  BUF_X4 U57407 ( .I(n37036), .Z(n14904) );
  INV_X2 U57408 ( .I(n34926), .ZN(n1777) );
  INV_X4 U57409 ( .I(n21878), .ZN(n34209) );
  INV_X4 U57410 ( .I(n12412), .ZN(n19435) );
  CLKBUF_X4 U57411 ( .I(n33715), .Z(n35964) );
  INV_X4 U57412 ( .I(n33715), .ZN(n21018) );
  OR2_X1 U57413 ( .A1(n35880), .A2(n57768), .Z(n65269) );
  BUF_X4 U57414 ( .I(n33721), .Z(n36170) );
  INV_X2 U57415 ( .I(n25998), .ZN(n40842) );
  INV_X4 U57416 ( .I(n19291), .ZN(n6170) );
  INV_X2 U57417 ( .I(n8452), .ZN(n40167) );
  AND2_X1 U57418 ( .A1(n38692), .A2(n40623), .Z(n65272) );
  INV_X4 U57419 ( .I(n19466), .ZN(n25816) );
  INV_X1 U57420 ( .I(n64793), .ZN(n40726) );
  INV_X2 U57421 ( .I(n38931), .ZN(n21791) );
  XNOR2_X1 U57422 ( .A1(n24508), .A2(n46497), .ZN(n65273) );
  INV_X2 U57423 ( .I(n6698), .ZN(n14448) );
  INV_X2 U57424 ( .I(n26166), .ZN(n1486) );
  AND2_X2 U57425 ( .A1(n46262), .A2(n58830), .Z(n65275) );
  INV_X2 U57426 ( .I(n47011), .ZN(n20091) );
  INV_X4 U57427 ( .I(n3654), .ZN(n58205) );
  OR2_X1 U57428 ( .A1(n46997), .A2(n48213), .Z(n65277) );
  AND3_X1 U57429 ( .A1(n49275), .A2(n19107), .A3(n49276), .Z(n65278) );
  INV_X4 U57430 ( .I(n6417), .ZN(n18196) );
  XNOR2_X1 U57431 ( .A1(n4451), .A2(n1618), .ZN(n65280) );
  INV_X4 U57432 ( .I(n53384), .ZN(n53198) );
  XOR2_X1 U57433 ( .A1(n50895), .A2(n50896), .Z(n65281) );
  INV_X2 U57434 ( .I(n8517), .ZN(n21877) );
  INV_X2 U57435 ( .I(n14178), .ZN(n22105) );
  INV_X4 U57436 ( .I(n17275), .ZN(n19167) );
  AND2_X2 U57437 ( .A1(n13485), .A2(n26143), .Z(n60710) );
  INV_X2 U57438 ( .I(n54000), .ZN(n2851) );
endmodule


module SPEEDY_Top ( clk, Ciphertext, Key, Plaintext );
  input [191:0] Ciphertext;
  input [191:0] Key;
  output [191:0] Plaintext;
  input clk;

  wire   [191:0] reg_in;
  wire   [191:0] reg_key;
  wire   [191:0] reg_out;

  DFFSNQ_X1 \reg_in_reg[191]  ( .D(Ciphertext[191]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[191]) );
  DFFSNQ_X1 \reg_in_reg[190]  ( .D(Ciphertext[190]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[190]) );
  DFFSNQ_X1 \reg_in_reg[189]  ( .D(Ciphertext[189]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[189]) );
  DFFSNQ_X1 \reg_in_reg[188]  ( .D(Ciphertext[188]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[188]) );
  DFFSNQ_X1 \reg_in_reg[187]  ( .D(Ciphertext[187]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[187]) );
  DFFSNQ_X1 \reg_in_reg[186]  ( .D(Ciphertext[186]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[186]) );
  DFFSNQ_X1 \reg_in_reg[185]  ( .D(Ciphertext[185]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[185]) );
  DFFSNQ_X1 \reg_in_reg[184]  ( .D(Ciphertext[184]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[184]) );
  DFFSNQ_X1 \reg_in_reg[183]  ( .D(Ciphertext[183]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[183]) );
  DFFSNQ_X1 \reg_in_reg[182]  ( .D(Ciphertext[182]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[182]) );
  DFFSNQ_X1 \reg_in_reg[181]  ( .D(Ciphertext[181]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[181]) );
  DFFSNQ_X1 \reg_in_reg[180]  ( .D(Ciphertext[180]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[180]) );
  DFFSNQ_X1 \reg_in_reg[179]  ( .D(Ciphertext[179]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[179]) );
  DFFSNQ_X1 \reg_in_reg[178]  ( .D(Ciphertext[178]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[178]) );
  DFFSNQ_X1 \reg_in_reg[177]  ( .D(Ciphertext[177]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[177]) );
  DFFSNQ_X1 \reg_in_reg[176]  ( .D(Ciphertext[176]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[176]) );
  DFFSNQ_X1 \reg_in_reg[175]  ( .D(Ciphertext[175]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[175]) );
  DFFSNQ_X1 \reg_in_reg[174]  ( .D(Ciphertext[174]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[174]) );
  DFFSNQ_X1 \reg_in_reg[173]  ( .D(Ciphertext[173]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[173]) );
  DFFSNQ_X1 \reg_in_reg[172]  ( .D(Ciphertext[172]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[172]) );
  DFFSNQ_X1 \reg_in_reg[171]  ( .D(Ciphertext[171]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[171]) );
  DFFSNQ_X1 \reg_in_reg[170]  ( .D(Ciphertext[170]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[170]) );
  DFFSNQ_X1 \reg_in_reg[169]  ( .D(Ciphertext[169]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[169]) );
  DFFSNQ_X1 \reg_in_reg[168]  ( .D(Ciphertext[168]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[168]) );
  DFFSNQ_X1 \reg_in_reg[167]  ( .D(Ciphertext[167]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[167]) );
  DFFSNQ_X1 \reg_in_reg[166]  ( .D(Ciphertext[166]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[166]) );
  DFFSNQ_X1 \reg_in_reg[164]  ( .D(Ciphertext[164]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[164]) );
  DFFSNQ_X1 \reg_in_reg[163]  ( .D(Ciphertext[163]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[163]) );
  DFFSNQ_X1 \reg_in_reg[162]  ( .D(Ciphertext[162]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[162]) );
  DFFSNQ_X1 \reg_in_reg[161]  ( .D(Ciphertext[161]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[161]) );
  DFFSNQ_X1 \reg_in_reg[160]  ( .D(Ciphertext[160]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[160]) );
  DFFSNQ_X1 \reg_in_reg[159]  ( .D(Ciphertext[159]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[159]) );
  DFFSNQ_X1 \reg_in_reg[157]  ( .D(Ciphertext[157]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[157]) );
  DFFSNQ_X1 \reg_in_reg[156]  ( .D(Ciphertext[156]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[156]) );
  DFFSNQ_X1 \reg_in_reg[155]  ( .D(Ciphertext[155]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[155]) );
  DFFSNQ_X1 \reg_in_reg[154]  ( .D(Ciphertext[154]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[154]) );
  DFFSNQ_X1 \reg_in_reg[153]  ( .D(Ciphertext[153]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[153]) );
  DFFSNQ_X1 \reg_in_reg[152]  ( .D(Ciphertext[152]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[152]) );
  DFFSNQ_X1 \reg_in_reg[151]  ( .D(Ciphertext[151]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[151]) );
  DFFSNQ_X1 \reg_in_reg[149]  ( .D(Ciphertext[149]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[149]) );
  DFFSNQ_X1 \reg_in_reg[148]  ( .D(Ciphertext[148]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[148]) );
  DFFSNQ_X1 \reg_in_reg[147]  ( .D(Ciphertext[147]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[147]) );
  DFFSNQ_X1 \reg_in_reg[146]  ( .D(Ciphertext[146]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[146]) );
  DFFSNQ_X1 \reg_in_reg[145]  ( .D(Ciphertext[145]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[145]) );
  DFFSNQ_X1 \reg_in_reg[144]  ( .D(Ciphertext[144]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[144]) );
  DFFSNQ_X1 \reg_in_reg[143]  ( .D(Ciphertext[143]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[143]) );
  DFFSNQ_X1 \reg_in_reg[142]  ( .D(Ciphertext[142]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[142]) );
  DFFSNQ_X1 \reg_in_reg[141]  ( .D(Ciphertext[141]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[141]) );
  DFFSNQ_X1 \reg_in_reg[140]  ( .D(Ciphertext[140]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[140]) );
  DFFSNQ_X1 \reg_in_reg[139]  ( .D(Ciphertext[139]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[139]) );
  DFFSNQ_X1 \reg_in_reg[138]  ( .D(Ciphertext[138]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[138]) );
  DFFSNQ_X1 \reg_in_reg[137]  ( .D(Ciphertext[137]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[137]) );
  DFFSNQ_X1 \reg_in_reg[136]  ( .D(Ciphertext[136]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[136]) );
  DFFSNQ_X1 \reg_in_reg[135]  ( .D(Ciphertext[135]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[135]) );
  DFFSNQ_X1 \reg_in_reg[134]  ( .D(Ciphertext[134]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[134]) );
  DFFSNQ_X1 \reg_in_reg[133]  ( .D(Ciphertext[133]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[133]) );
  DFFSNQ_X1 \reg_in_reg[132]  ( .D(Ciphertext[132]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[132]) );
  DFFSNQ_X1 \reg_in_reg[131]  ( .D(Ciphertext[131]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[131]) );
  DFFSNQ_X1 \reg_in_reg[130]  ( .D(Ciphertext[130]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[130]) );
  DFFSNQ_X1 \reg_in_reg[129]  ( .D(Ciphertext[129]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[129]) );
  DFFSNQ_X1 \reg_in_reg[128]  ( .D(Ciphertext[128]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[128]) );
  DFFSNQ_X1 \reg_in_reg[127]  ( .D(Ciphertext[127]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[127]) );
  DFFSNQ_X1 \reg_in_reg[126]  ( .D(Ciphertext[126]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[126]) );
  DFFSNQ_X1 \reg_in_reg[125]  ( .D(Ciphertext[125]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[125]) );
  DFFSNQ_X1 \reg_in_reg[124]  ( .D(Ciphertext[124]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[124]) );
  DFFSNQ_X1 \reg_in_reg[123]  ( .D(Ciphertext[123]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[123]) );
  DFFSNQ_X1 \reg_in_reg[122]  ( .D(Ciphertext[122]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[122]) );
  DFFSNQ_X1 \reg_in_reg[121]  ( .D(Ciphertext[121]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[121]) );
  DFFSNQ_X1 \reg_in_reg[120]  ( .D(Ciphertext[120]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[120]) );
  DFFSNQ_X1 \reg_in_reg[119]  ( .D(Ciphertext[119]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[119]) );
  DFFSNQ_X1 \reg_in_reg[118]  ( .D(Ciphertext[118]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[118]) );
  DFFSNQ_X1 \reg_in_reg[117]  ( .D(Ciphertext[117]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[117]) );
  DFFSNQ_X1 \reg_in_reg[116]  ( .D(Ciphertext[116]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[116]) );
  DFFSNQ_X1 \reg_in_reg[115]  ( .D(Ciphertext[115]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[115]) );
  DFFSNQ_X1 \reg_in_reg[114]  ( .D(Ciphertext[114]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[114]) );
  DFFSNQ_X1 \reg_in_reg[113]  ( .D(Ciphertext[113]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[113]) );
  DFFSNQ_X1 \reg_in_reg[112]  ( .D(Ciphertext[112]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[112]) );
  DFFSNQ_X1 \reg_in_reg[111]  ( .D(Ciphertext[111]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[111]) );
  DFFSNQ_X1 \reg_in_reg[110]  ( .D(Ciphertext[110]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[110]) );
  DFFSNQ_X1 \reg_in_reg[109]  ( .D(Ciphertext[109]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[109]) );
  DFFSNQ_X1 \reg_in_reg[108]  ( .D(Ciphertext[108]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[108]) );
  DFFSNQ_X1 \reg_in_reg[107]  ( .D(Ciphertext[107]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[107]) );
  DFFSNQ_X1 \reg_in_reg[106]  ( .D(Ciphertext[106]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[106]) );
  DFFSNQ_X1 \reg_in_reg[105]  ( .D(Ciphertext[105]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[105]) );
  DFFSNQ_X1 \reg_in_reg[104]  ( .D(Ciphertext[104]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[104]) );
  DFFSNQ_X1 \reg_in_reg[103]  ( .D(Ciphertext[103]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[103]) );
  DFFSNQ_X1 \reg_in_reg[102]  ( .D(Ciphertext[102]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[102]) );
  DFFSNQ_X1 \reg_in_reg[101]  ( .D(Ciphertext[101]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[101]) );
  DFFSNQ_X1 \reg_in_reg[100]  ( .D(Ciphertext[100]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[100]) );
  DFFSNQ_X1 \reg_in_reg[99]  ( .D(Ciphertext[99]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[99]) );
  DFFSNQ_X1 \reg_in_reg[98]  ( .D(Ciphertext[98]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[98]) );
  DFFSNQ_X1 \reg_in_reg[97]  ( .D(Ciphertext[97]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[97]) );
  DFFSNQ_X1 \reg_in_reg[96]  ( .D(Ciphertext[96]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[96]) );
  DFFSNQ_X1 \reg_in_reg[95]  ( .D(Ciphertext[95]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[95]) );
  DFFSNQ_X1 \reg_in_reg[94]  ( .D(Ciphertext[94]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[94]) );
  DFFSNQ_X1 \reg_in_reg[93]  ( .D(Ciphertext[93]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[93]) );
  DFFSNQ_X1 \reg_in_reg[92]  ( .D(Ciphertext[92]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[92]) );
  DFFSNQ_X1 \reg_in_reg[91]  ( .D(Ciphertext[91]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[91]) );
  DFFSNQ_X1 \reg_in_reg[90]  ( .D(Ciphertext[90]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[90]) );
  DFFSNQ_X1 \reg_in_reg[89]  ( .D(Ciphertext[89]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[89]) );
  DFFSNQ_X1 \reg_in_reg[88]  ( .D(Ciphertext[88]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[88]) );
  DFFSNQ_X1 \reg_in_reg[87]  ( .D(Ciphertext[87]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[87]) );
  DFFSNQ_X1 \reg_in_reg[86]  ( .D(Ciphertext[86]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[86]) );
  DFFSNQ_X1 \reg_in_reg[85]  ( .D(Ciphertext[85]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[85]) );
  DFFSNQ_X1 \reg_in_reg[84]  ( .D(Ciphertext[84]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[84]) );
  DFFSNQ_X1 \reg_in_reg[83]  ( .D(Ciphertext[83]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[83]) );
  DFFSNQ_X1 \reg_in_reg[82]  ( .D(Ciphertext[82]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[82]) );
  DFFSNQ_X1 \reg_in_reg[81]  ( .D(Ciphertext[81]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[81]) );
  DFFSNQ_X1 \reg_in_reg[80]  ( .D(Ciphertext[80]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[80]) );
  DFFSNQ_X1 \reg_in_reg[79]  ( .D(Ciphertext[79]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[79]) );
  DFFSNQ_X1 \reg_in_reg[77]  ( .D(Ciphertext[77]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[77]) );
  DFFSNQ_X1 \reg_in_reg[76]  ( .D(Ciphertext[76]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[76]) );
  DFFSNQ_X1 \reg_in_reg[75]  ( .D(Ciphertext[75]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[75]) );
  DFFSNQ_X1 \reg_in_reg[74]  ( .D(Ciphertext[74]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[74]) );
  DFFSNQ_X1 \reg_in_reg[73]  ( .D(Ciphertext[73]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[73]) );
  DFFSNQ_X1 \reg_in_reg[72]  ( .D(Ciphertext[72]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[72]) );
  DFFSNQ_X1 \reg_in_reg[71]  ( .D(Ciphertext[71]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[71]) );
  DFFSNQ_X1 \reg_in_reg[70]  ( .D(Ciphertext[70]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[70]) );
  DFFSNQ_X1 \reg_in_reg[69]  ( .D(Ciphertext[69]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[69]) );
  DFFSNQ_X1 \reg_in_reg[68]  ( .D(Ciphertext[68]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[68]) );
  DFFSNQ_X1 \reg_in_reg[67]  ( .D(Ciphertext[67]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[67]) );
  DFFSNQ_X1 \reg_in_reg[66]  ( .D(Ciphertext[66]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[66]) );
  DFFSNQ_X1 \reg_in_reg[65]  ( .D(Ciphertext[65]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[65]) );
  DFFSNQ_X1 \reg_in_reg[64]  ( .D(Ciphertext[64]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[64]) );
  DFFSNQ_X1 \reg_in_reg[63]  ( .D(Ciphertext[63]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[63]) );
  DFFSNQ_X1 \reg_in_reg[62]  ( .D(Ciphertext[62]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[62]) );
  DFFSNQ_X1 \reg_in_reg[61]  ( .D(Ciphertext[61]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[61]) );
  DFFSNQ_X1 \reg_in_reg[60]  ( .D(Ciphertext[60]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[60]) );
  DFFSNQ_X1 \reg_in_reg[59]  ( .D(Ciphertext[59]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[59]) );
  DFFSNQ_X1 \reg_in_reg[58]  ( .D(Ciphertext[58]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[58]) );
  DFFSNQ_X1 \reg_in_reg[57]  ( .D(Ciphertext[57]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[57]) );
  DFFSNQ_X1 \reg_in_reg[56]  ( .D(Ciphertext[56]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[56]) );
  DFFSNQ_X1 \reg_in_reg[55]  ( .D(Ciphertext[55]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[55]) );
  DFFSNQ_X1 \reg_in_reg[54]  ( .D(Ciphertext[54]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[54]) );
  DFFSNQ_X1 \reg_in_reg[53]  ( .D(Ciphertext[53]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[53]) );
  DFFSNQ_X1 \reg_in_reg[52]  ( .D(Ciphertext[52]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[52]) );
  DFFSNQ_X1 \reg_in_reg[50]  ( .D(Ciphertext[50]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[50]) );
  DFFSNQ_X1 \reg_in_reg[49]  ( .D(Ciphertext[49]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[49]) );
  DFFSNQ_X1 \reg_in_reg[48]  ( .D(Ciphertext[48]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[48]) );
  DFFSNQ_X1 \reg_in_reg[47]  ( .D(Ciphertext[47]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[47]) );
  DFFSNQ_X1 \reg_in_reg[46]  ( .D(Ciphertext[46]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[46]) );
  DFFSNQ_X1 \reg_in_reg[45]  ( .D(Ciphertext[45]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[45]) );
  DFFSNQ_X1 \reg_in_reg[44]  ( .D(Ciphertext[44]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[44]) );
  DFFSNQ_X1 \reg_in_reg[43]  ( .D(Ciphertext[43]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[43]) );
  DFFSNQ_X1 \reg_in_reg[42]  ( .D(Ciphertext[42]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[42]) );
  DFFSNQ_X1 \reg_in_reg[41]  ( .D(Ciphertext[41]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[41]) );
  DFFSNQ_X1 \reg_in_reg[40]  ( .D(Ciphertext[40]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[40]) );
  DFFSNQ_X1 \reg_in_reg[39]  ( .D(Ciphertext[39]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[39]) );
  DFFSNQ_X1 \reg_in_reg[38]  ( .D(Ciphertext[38]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[38]) );
  DFFSNQ_X1 \reg_in_reg[37]  ( .D(Ciphertext[37]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[37]) );
  DFFSNQ_X1 \reg_in_reg[36]  ( .D(Ciphertext[36]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[36]) );
  DFFSNQ_X1 \reg_in_reg[35]  ( .D(Ciphertext[35]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[35]) );
  DFFSNQ_X1 \reg_in_reg[34]  ( .D(Ciphertext[34]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[34]) );
  DFFSNQ_X1 \reg_in_reg[33]  ( .D(Ciphertext[33]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[33]) );
  DFFSNQ_X1 \reg_in_reg[32]  ( .D(Ciphertext[32]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[32]) );
  DFFSNQ_X1 \reg_in_reg[31]  ( .D(Ciphertext[31]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[31]) );
  DFFSNQ_X1 \reg_in_reg[30]  ( .D(Ciphertext[30]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[30]) );
  DFFSNQ_X1 \reg_in_reg[29]  ( .D(Ciphertext[29]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[29]) );
  DFFSNQ_X1 \reg_in_reg[28]  ( .D(Ciphertext[28]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[28]) );
  DFFSNQ_X1 \reg_in_reg[27]  ( .D(Ciphertext[27]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[27]) );
  DFFSNQ_X1 \reg_in_reg[26]  ( .D(Ciphertext[26]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[26]) );
  DFFSNQ_X1 \reg_in_reg[25]  ( .D(Ciphertext[25]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[25]) );
  DFFSNQ_X1 \reg_in_reg[24]  ( .D(Ciphertext[24]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[24]) );
  DFFSNQ_X1 \reg_in_reg[23]  ( .D(Ciphertext[23]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[23]) );
  DFFSNQ_X1 \reg_in_reg[22]  ( .D(Ciphertext[22]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[22]) );
  DFFSNQ_X1 \reg_in_reg[21]  ( .D(Ciphertext[21]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[21]) );
  DFFSNQ_X1 \reg_in_reg[20]  ( .D(Ciphertext[20]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[20]) );
  DFFSNQ_X1 \reg_in_reg[19]  ( .D(Ciphertext[19]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[19]) );
  DFFSNQ_X1 \reg_in_reg[18]  ( .D(Ciphertext[18]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[18]) );
  DFFSNQ_X1 \reg_in_reg[17]  ( .D(Ciphertext[17]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[17]) );
  DFFSNQ_X1 \reg_in_reg[16]  ( .D(Ciphertext[16]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[16]) );
  DFFSNQ_X1 \reg_in_reg[15]  ( .D(Ciphertext[15]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[15]) );
  DFFSNQ_X1 \reg_in_reg[14]  ( .D(Ciphertext[14]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[14]) );
  DFFSNQ_X1 \reg_in_reg[13]  ( .D(Ciphertext[13]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[13]) );
  DFFSNQ_X1 \reg_in_reg[12]  ( .D(Ciphertext[12]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[12]) );
  DFFSNQ_X1 \reg_in_reg[11]  ( .D(Ciphertext[11]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[11]) );
  DFFSNQ_X1 \reg_in_reg[10]  ( .D(Ciphertext[10]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[10]) );
  DFFSNQ_X1 \reg_in_reg[9]  ( .D(Ciphertext[9]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[9]) );
  DFFSNQ_X1 \reg_in_reg[8]  ( .D(Ciphertext[8]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[8]) );
  DFFSNQ_X1 \reg_in_reg[7]  ( .D(Ciphertext[7]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[7]) );
  DFFSNQ_X1 \reg_in_reg[6]  ( .D(Ciphertext[6]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[6]) );
  DFFSNQ_X1 \reg_in_reg[5]  ( .D(Ciphertext[5]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[5]) );
  DFFSNQ_X1 \reg_in_reg[4]  ( .D(Ciphertext[4]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[4]) );
  DFFSNQ_X1 \reg_in_reg[3]  ( .D(Ciphertext[3]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[3]) );
  DFFSNQ_X1 \reg_in_reg[2]  ( .D(Ciphertext[2]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[2]) );
  DFFSNQ_X1 \reg_in_reg[1]  ( .D(Ciphertext[1]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[1]) );
  DFFSNQ_X1 \reg_in_reg[0]  ( .D(Ciphertext[0]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[0]) );
  DFFSNQ_X1 \reg_key_reg[191]  ( .D(Key[191]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[191]) );
  DFFSNQ_X1 \reg_key_reg[190]  ( .D(Key[190]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[190]) );
  DFFSNQ_X1 \reg_key_reg[189]  ( .D(Key[189]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[189]) );
  DFFSNQ_X1 \reg_key_reg[188]  ( .D(Key[188]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[188]) );
  DFFSNQ_X1 \reg_key_reg[187]  ( .D(Key[187]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[187]) );
  DFFSNQ_X1 \reg_key_reg[186]  ( .D(Key[186]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[186]) );
  DFFSNQ_X1 \reg_key_reg[185]  ( .D(Key[185]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[185]) );
  DFFSNQ_X1 \reg_key_reg[184]  ( .D(Key[184]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[184]) );
  DFFSNQ_X1 \reg_key_reg[183]  ( .D(Key[183]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[183]) );
  DFFSNQ_X1 \reg_key_reg[182]  ( .D(Key[182]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[182]) );
  DFFSNQ_X1 \reg_key_reg[181]  ( .D(Key[181]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[181]) );
  DFFSNQ_X1 \reg_key_reg[180]  ( .D(Key[180]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[180]) );
  DFFSNQ_X1 \reg_key_reg[179]  ( .D(Key[179]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[179]) );
  DFFSNQ_X1 \reg_key_reg[178]  ( .D(Key[178]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[178]) );
  DFFSNQ_X1 \reg_key_reg[177]  ( .D(Key[177]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[177]) );
  DFFSNQ_X1 \reg_key_reg[176]  ( .D(Key[176]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[176]) );
  DFFSNQ_X1 \reg_key_reg[175]  ( .D(Key[175]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[175]) );
  DFFSNQ_X1 \reg_key_reg[174]  ( .D(Key[174]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[174]) );
  DFFSNQ_X1 \reg_key_reg[173]  ( .D(Key[173]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[173]) );
  DFFSNQ_X1 \reg_key_reg[172]  ( .D(Key[172]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[172]) );
  DFFSNQ_X1 \reg_key_reg[171]  ( .D(Key[171]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[171]) );
  DFFSNQ_X1 \reg_key_reg[170]  ( .D(Key[170]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[170]) );
  DFFSNQ_X1 \reg_key_reg[169]  ( .D(Key[169]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[169]) );
  DFFSNQ_X1 \reg_key_reg[168]  ( .D(Key[168]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[168]) );
  DFFSNQ_X1 \reg_key_reg[167]  ( .D(Key[167]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[167]) );
  DFFSNQ_X1 \reg_key_reg[166]  ( .D(Key[166]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[166]) );
  DFFSNQ_X1 \reg_key_reg[165]  ( .D(Key[165]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[165]) );
  DFFSNQ_X1 \reg_key_reg[164]  ( .D(Key[164]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[164]) );
  DFFSNQ_X1 \reg_key_reg[163]  ( .D(Key[163]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[163]) );
  DFFSNQ_X1 \reg_key_reg[162]  ( .D(Key[162]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[162]) );
  DFFSNQ_X1 \reg_key_reg[161]  ( .D(Key[161]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[161]) );
  DFFSNQ_X1 \reg_key_reg[160]  ( .D(Key[160]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[160]) );
  DFFSNQ_X1 \reg_key_reg[159]  ( .D(Key[159]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[159]) );
  DFFSNQ_X1 \reg_key_reg[158]  ( .D(Key[158]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[158]) );
  DFFSNQ_X1 \reg_key_reg[157]  ( .D(Key[157]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[157]) );
  DFFSNQ_X1 \reg_key_reg[156]  ( .D(Key[156]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[156]) );
  DFFSNQ_X1 \reg_key_reg[155]  ( .D(Key[155]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[155]) );
  DFFSNQ_X1 \reg_key_reg[154]  ( .D(Key[154]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[154]) );
  DFFSNQ_X1 \reg_key_reg[153]  ( .D(Key[153]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[153]) );
  DFFSNQ_X1 \reg_key_reg[152]  ( .D(Key[152]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[152]) );
  DFFSNQ_X1 \reg_key_reg[151]  ( .D(Key[151]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[151]) );
  DFFSNQ_X1 \reg_key_reg[150]  ( .D(Key[150]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[150]) );
  DFFSNQ_X1 \reg_key_reg[149]  ( .D(Key[149]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[149]) );
  DFFSNQ_X1 \reg_key_reg[148]  ( .D(Key[148]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[148]) );
  DFFSNQ_X1 \reg_key_reg[147]  ( .D(Key[147]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[147]) );
  DFFSNQ_X1 \reg_key_reg[146]  ( .D(Key[146]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[146]) );
  DFFSNQ_X1 \reg_key_reg[145]  ( .D(Key[145]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[145]) );
  DFFSNQ_X1 \reg_key_reg[144]  ( .D(Key[144]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[144]) );
  DFFSNQ_X1 \reg_key_reg[143]  ( .D(Key[143]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[143]) );
  DFFSNQ_X1 \reg_key_reg[142]  ( .D(Key[142]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[142]) );
  DFFSNQ_X1 \reg_key_reg[141]  ( .D(Key[141]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[141]) );
  DFFSNQ_X1 \reg_key_reg[140]  ( .D(Key[140]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[140]) );
  DFFSNQ_X1 \reg_key_reg[139]  ( .D(Key[139]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[139]) );
  DFFSNQ_X1 \reg_key_reg[138]  ( .D(Key[138]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[138]) );
  DFFSNQ_X1 \reg_key_reg[137]  ( .D(Key[137]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[137]) );
  DFFSNQ_X1 \reg_key_reg[136]  ( .D(Key[136]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[136]) );
  DFFSNQ_X1 \reg_key_reg[135]  ( .D(Key[135]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[135]) );
  DFFSNQ_X1 \reg_key_reg[134]  ( .D(Key[134]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[134]) );
  DFFSNQ_X1 \reg_key_reg[133]  ( .D(Key[133]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[133]) );
  DFFSNQ_X1 \reg_key_reg[132]  ( .D(Key[132]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[132]) );
  DFFSNQ_X1 \reg_key_reg[130]  ( .D(Key[130]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[130]) );
  DFFSNQ_X1 \reg_key_reg[129]  ( .D(Key[129]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[129]) );
  DFFSNQ_X1 \reg_key_reg[128]  ( .D(Key[128]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[128]) );
  DFFSNQ_X1 \reg_key_reg[127]  ( .D(Key[127]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[127]) );
  DFFSNQ_X1 \reg_key_reg[126]  ( .D(Key[126]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[126]) );
  DFFSNQ_X1 \reg_key_reg[125]  ( .D(Key[125]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[125]) );
  DFFSNQ_X1 \reg_key_reg[124]  ( .D(Key[124]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[124]) );
  DFFSNQ_X1 \reg_key_reg[123]  ( .D(Key[123]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[123]) );
  DFFSNQ_X1 \reg_key_reg[122]  ( .D(Key[122]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[122]) );
  DFFSNQ_X1 \reg_key_reg[121]  ( .D(Key[121]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[121]) );
  DFFSNQ_X1 \reg_key_reg[120]  ( .D(Key[120]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[120]) );
  DFFSNQ_X1 \reg_key_reg[119]  ( .D(Key[119]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[119]) );
  DFFSNQ_X1 \reg_key_reg[117]  ( .D(Key[117]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[117]) );
  DFFSNQ_X1 \reg_key_reg[116]  ( .D(Key[116]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[116]) );
  DFFSNQ_X1 \reg_key_reg[115]  ( .D(Key[115]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[115]) );
  DFFSNQ_X1 \reg_key_reg[114]  ( .D(Key[114]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[114]) );
  DFFSNQ_X1 \reg_key_reg[113]  ( .D(Key[113]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[113]) );
  DFFSNQ_X1 \reg_key_reg[112]  ( .D(Key[112]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[112]) );
  DFFSNQ_X1 \reg_key_reg[111]  ( .D(Key[111]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[111]) );
  DFFSNQ_X1 \reg_key_reg[110]  ( .D(Key[110]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[110]) );
  DFFSNQ_X1 \reg_key_reg[109]  ( .D(Key[109]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[109]) );
  DFFSNQ_X1 \reg_key_reg[108]  ( .D(Key[108]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[108]) );
  DFFSNQ_X1 \reg_key_reg[107]  ( .D(Key[107]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[107]) );
  DFFSNQ_X1 \reg_key_reg[106]  ( .D(Key[106]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[106]) );
  DFFSNQ_X1 \reg_key_reg[105]  ( .D(Key[105]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[105]) );
  DFFSNQ_X1 \reg_key_reg[104]  ( .D(Key[104]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[104]) );
  DFFSNQ_X1 \reg_key_reg[103]  ( .D(Key[103]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[103]) );
  DFFSNQ_X1 \reg_key_reg[102]  ( .D(Key[102]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[102]) );
  DFFSNQ_X1 \reg_key_reg[101]  ( .D(Key[101]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[101]) );
  DFFSNQ_X1 \reg_key_reg[100]  ( .D(Key[100]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[100]) );
  DFFSNQ_X1 \reg_key_reg[99]  ( .D(Key[99]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[99]) );
  DFFSNQ_X1 \reg_key_reg[98]  ( .D(Key[98]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[98]) );
  DFFSNQ_X1 \reg_key_reg[97]  ( .D(Key[97]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[97]) );
  DFFSNQ_X1 \reg_key_reg[96]  ( .D(Key[96]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[96]) );
  DFFSNQ_X1 \reg_key_reg[95]  ( .D(Key[95]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[95]) );
  DFFSNQ_X1 \reg_key_reg[94]  ( .D(Key[94]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[94]) );
  DFFSNQ_X1 \reg_key_reg[93]  ( .D(Key[93]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[93]) );
  DFFSNQ_X1 \reg_key_reg[92]  ( .D(Key[92]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[92]) );
  DFFSNQ_X1 \reg_key_reg[91]  ( .D(Key[91]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[91]) );
  DFFSNQ_X1 \reg_key_reg[90]  ( .D(Key[90]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[90]) );
  DFFSNQ_X1 \reg_key_reg[89]  ( .D(Key[89]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[89]) );
  DFFSNQ_X1 \reg_key_reg[88]  ( .D(Key[88]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[88]) );
  DFFSNQ_X1 \reg_key_reg[87]  ( .D(Key[87]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[87]) );
  DFFSNQ_X1 \reg_key_reg[86]  ( .D(Key[86]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[86]) );
  DFFSNQ_X1 \reg_key_reg[85]  ( .D(Key[85]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[85]) );
  DFFSNQ_X1 \reg_key_reg[84]  ( .D(Key[84]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[84]) );
  DFFSNQ_X1 \reg_key_reg[83]  ( .D(Key[83]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[83]) );
  DFFSNQ_X1 \reg_key_reg[82]  ( .D(Key[82]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[82]) );
  DFFSNQ_X1 \reg_key_reg[81]  ( .D(Key[81]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[81]) );
  DFFSNQ_X1 \reg_key_reg[80]  ( .D(Key[80]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[80]) );
  DFFSNQ_X1 \reg_key_reg[79]  ( .D(Key[79]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[79]) );
  DFFSNQ_X1 \reg_key_reg[78]  ( .D(Key[78]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[78]) );
  DFFSNQ_X1 \reg_key_reg[77]  ( .D(Key[77]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[77]) );
  DFFSNQ_X1 \reg_key_reg[76]  ( .D(Key[76]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[76]) );
  DFFSNQ_X1 \reg_key_reg[75]  ( .D(Key[75]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[75]) );
  DFFSNQ_X1 \reg_key_reg[74]  ( .D(Key[74]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[74]) );
  DFFSNQ_X1 \reg_key_reg[73]  ( .D(Key[73]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[73]) );
  DFFSNQ_X1 \reg_key_reg[72]  ( .D(Key[72]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[72]) );
  DFFSNQ_X1 \reg_key_reg[71]  ( .D(Key[71]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[71]) );
  DFFSNQ_X1 \reg_key_reg[70]  ( .D(Key[70]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[70]) );
  DFFSNQ_X1 \reg_key_reg[69]  ( .D(Key[69]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[69]) );
  DFFSNQ_X1 \reg_key_reg[68]  ( .D(Key[68]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[68]) );
  DFFSNQ_X1 \reg_key_reg[67]  ( .D(Key[67]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[67]) );
  DFFSNQ_X1 \reg_key_reg[66]  ( .D(Key[66]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[66]) );
  DFFSNQ_X1 \reg_key_reg[65]  ( .D(Key[65]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[65]) );
  DFFSNQ_X1 \reg_key_reg[64]  ( .D(Key[64]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[64]) );
  DFFSNQ_X1 \reg_key_reg[63]  ( .D(Key[63]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[63]) );
  DFFSNQ_X1 \reg_key_reg[62]  ( .D(Key[62]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[62]) );
  DFFSNQ_X1 \reg_key_reg[61]  ( .D(Key[61]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[61]) );
  DFFSNQ_X1 \reg_key_reg[60]  ( .D(Key[60]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[60]) );
  DFFSNQ_X1 \reg_key_reg[59]  ( .D(Key[59]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[59]) );
  DFFSNQ_X1 \reg_key_reg[58]  ( .D(Key[58]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[58]) );
  DFFSNQ_X1 \reg_key_reg[57]  ( .D(Key[57]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[57]) );
  DFFSNQ_X1 \reg_key_reg[56]  ( .D(Key[56]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[56]) );
  DFFSNQ_X1 \reg_key_reg[55]  ( .D(Key[55]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[55]) );
  DFFSNQ_X1 \reg_key_reg[54]  ( .D(Key[54]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[54]) );
  DFFSNQ_X1 \reg_key_reg[53]  ( .D(Key[53]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[53]) );
  DFFSNQ_X1 \reg_key_reg[52]  ( .D(Key[52]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[52]) );
  DFFSNQ_X1 \reg_key_reg[51]  ( .D(Key[51]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[51]) );
  DFFSNQ_X1 \reg_key_reg[50]  ( .D(Key[50]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[50]) );
  DFFSNQ_X1 \reg_key_reg[49]  ( .D(Key[49]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[49]) );
  DFFSNQ_X1 \reg_key_reg[48]  ( .D(Key[48]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[48]) );
  DFFSNQ_X1 \reg_key_reg[47]  ( .D(Key[47]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[47]) );
  DFFSNQ_X1 \reg_key_reg[46]  ( .D(Key[46]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[46]) );
  DFFSNQ_X1 \reg_key_reg[45]  ( .D(Key[45]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[45]) );
  DFFSNQ_X1 \reg_key_reg[44]  ( .D(Key[44]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[44]) );
  DFFSNQ_X1 \reg_key_reg[43]  ( .D(Key[43]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[43]) );
  DFFSNQ_X1 \reg_key_reg[42]  ( .D(Key[42]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[42]) );
  DFFSNQ_X1 \reg_key_reg[41]  ( .D(Key[41]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[41]) );
  DFFSNQ_X1 \reg_key_reg[40]  ( .D(Key[40]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[40]) );
  DFFSNQ_X1 \reg_key_reg[39]  ( .D(Key[39]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[39]) );
  DFFSNQ_X1 \reg_key_reg[38]  ( .D(Key[38]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[38]) );
  DFFSNQ_X1 \reg_key_reg[37]  ( .D(Key[37]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[37]) );
  DFFSNQ_X1 \reg_key_reg[36]  ( .D(Key[36]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[36]) );
  DFFSNQ_X1 \reg_key_reg[35]  ( .D(Key[35]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[35]) );
  DFFSNQ_X1 \reg_key_reg[34]  ( .D(Key[34]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[34]) );
  DFFSNQ_X1 \reg_key_reg[33]  ( .D(Key[33]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[33]) );
  DFFSNQ_X1 \reg_key_reg[32]  ( .D(Key[32]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[32]) );
  DFFSNQ_X1 \reg_key_reg[31]  ( .D(Key[31]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[31]) );
  DFFSNQ_X1 \reg_key_reg[30]  ( .D(Key[30]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[30]) );
  DFFSNQ_X1 \reg_key_reg[29]  ( .D(Key[29]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[29]) );
  DFFSNQ_X1 \reg_key_reg[28]  ( .D(Key[28]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[28]) );
  DFFSNQ_X1 \reg_key_reg[27]  ( .D(Key[27]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[27]) );
  DFFSNQ_X1 \reg_key_reg[26]  ( .D(Key[26]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[26]) );
  DFFSNQ_X1 \reg_key_reg[25]  ( .D(Key[25]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[25]) );
  DFFSNQ_X1 \reg_key_reg[24]  ( .D(Key[24]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[24]) );
  DFFSNQ_X1 \reg_key_reg[23]  ( .D(Key[23]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[23]) );
  DFFSNQ_X1 \reg_key_reg[22]  ( .D(Key[22]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[22]) );
  DFFSNQ_X1 \reg_key_reg[21]  ( .D(Key[21]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[21]) );
  DFFSNQ_X1 \reg_key_reg[20]  ( .D(Key[20]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[20]) );
  DFFSNQ_X1 \reg_key_reg[19]  ( .D(Key[19]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[19]) );
  DFFSNQ_X1 \reg_key_reg[18]  ( .D(Key[18]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[18]) );
  DFFSNQ_X1 \reg_key_reg[17]  ( .D(Key[17]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[17]) );
  DFFSNQ_X1 \reg_key_reg[16]  ( .D(Key[16]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[16]) );
  DFFSNQ_X1 \reg_key_reg[15]  ( .D(Key[15]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[15]) );
  DFFSNQ_X1 \reg_key_reg[14]  ( .D(Key[14]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[14]) );
  DFFSNQ_X1 \reg_key_reg[13]  ( .D(Key[13]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[13]) );
  DFFSNQ_X1 \reg_key_reg[12]  ( .D(Key[12]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[12]) );
  DFFSNQ_X1 \reg_key_reg[11]  ( .D(Key[11]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[11]) );
  DFFSNQ_X1 \reg_key_reg[10]  ( .D(Key[10]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[10]) );
  DFFSNQ_X1 \reg_key_reg[9]  ( .D(Key[9]), .CLK(clk), .SN(1'b1), .Q(reg_key[9]) );
  DFFSNQ_X1 \reg_key_reg[8]  ( .D(Key[8]), .CLK(clk), .SN(1'b1), .Q(reg_key[8]) );
  DFFSNQ_X1 \reg_key_reg[7]  ( .D(Key[7]), .CLK(clk), .SN(1'b1), .Q(reg_key[7]) );
  DFFSNQ_X1 \reg_key_reg[6]  ( .D(Key[6]), .CLK(clk), .SN(1'b1), .Q(reg_key[6]) );
  DFFSNQ_X1 \reg_key_reg[5]  ( .D(Key[5]), .CLK(clk), .SN(1'b1), .Q(reg_key[5]) );
  DFFSNQ_X1 \reg_key_reg[4]  ( .D(Key[4]), .CLK(clk), .SN(1'b1), .Q(reg_key[4]) );
  DFFSNQ_X1 \reg_key_reg[3]  ( .D(Key[3]), .CLK(clk), .SN(1'b1), .Q(reg_key[3]) );
  DFFSNQ_X1 \reg_key_reg[2]  ( .D(Key[2]), .CLK(clk), .SN(1'b1), .Q(reg_key[2]) );
  DFFSNQ_X1 \reg_key_reg[1]  ( .D(Key[1]), .CLK(clk), .SN(1'b1), .Q(reg_key[1]) );
  DFFSNQ_X1 \reg_key_reg[0]  ( .D(Key[0]), .CLK(clk), .SN(1'b1), .Q(reg_key[0]) );
  DFFRNQ_X1 \Plaintext_reg[35]  ( .D(reg_out[35]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[35]) );
  DFFRNQ_X1 \Plaintext_reg[32]  ( .D(reg_out[32]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[32]) );
  DFFRNQ_X1 \Plaintext_reg[30]  ( .D(reg_out[30]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[30]) );
  DFFRNQ_X1 \Plaintext_reg[34]  ( .D(reg_out[34]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[34]) );
  DFFRNQ_X1 \Plaintext_reg[164]  ( .D(reg_out[164]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[164]) );
  DFFRNQ_X1 \Plaintext_reg[26]  ( .D(reg_out[26]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[26]) );
  DFFRNQ_X1 \Plaintext_reg[74]  ( .D(reg_out[74]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[74]) );
  DFFRNQ_X1 \Plaintext_reg[166]  ( .D(reg_out[166]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[166]) );
  DFFRNQ_X1 \Plaintext_reg[75]  ( .D(reg_out[75]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[75]) );
  DFFRNQ_X1 \Plaintext_reg[122]  ( .D(reg_out[122]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[122]) );
  DFFRNQ_X1 \Plaintext_reg[50]  ( .D(reg_out[50]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[50]) );
  DFFRNQ_X1 \Plaintext_reg[170]  ( .D(reg_out[170]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[170]) );
  DFFRNQ_X1 \Plaintext_reg[98]  ( .D(reg_out[98]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[98]) );
  DFFRNQ_X1 \Plaintext_reg[14]  ( .D(reg_out[14]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[14]) );
  DFFRNQ_X1 \Plaintext_reg[31]  ( .D(reg_out[31]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[31]) );
  DFFRNQ_X1 \Plaintext_reg[57]  ( .D(reg_out[57]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[57]) );
  DFFRNQ_X1 \Plaintext_reg[138]  ( .D(reg_out[138]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[138]) );
  DFFRNQ_X1 \Plaintext_reg[167]  ( .D(reg_out[167]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[167]) );
  DFFRNQ_X1 \Plaintext_reg[64]  ( .D(reg_out[64]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[64]) );
  DFFRNQ_X1 \Plaintext_reg[108]  ( .D(reg_out[108]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[108]) );
  DFFRNQ_X1 \Plaintext_reg[124]  ( .D(reg_out[124]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[124]) );
  DFFRNQ_X1 \Plaintext_reg[29]  ( .D(reg_out[29]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[29]) );
  DFFRNQ_X1 \Plaintext_reg[24]  ( .D(reg_out[24]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[24]) );
  DFFRNQ_X1 \Plaintext_reg[110]  ( .D(reg_out[110]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[110]) );
  DFFRNQ_X1 \Plaintext_reg[114]  ( .D(reg_out[114]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[114]) );
  DFFRNQ_X1 \Plaintext_reg[176]  ( .D(reg_out[176]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[176]) );
  DFFRNQ_X1 \Plaintext_reg[27]  ( .D(reg_out[27]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[27]) );
  DFFRNQ_X1 \Plaintext_reg[22]  ( .D(reg_out[22]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[22]) );
  DFFRNQ_X1 \Plaintext_reg[86]  ( .D(reg_out[86]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[86]) );
  DFFRNQ_X1 \Plaintext_reg[58]  ( .D(reg_out[58]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[58]) );
  DFFRNQ_X1 \Plaintext_reg[84]  ( .D(reg_out[84]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[84]) );
  DFFRNQ_X1 \Plaintext_reg[8]  ( .D(reg_out[8]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[8]) );
  DFFRNQ_X1 \Plaintext_reg[152]  ( .D(reg_out[152]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[152]) );
  DFFRNQ_X1 \Plaintext_reg[68]  ( .D(reg_out[68]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[68]) );
  DFFRNQ_X1 \Plaintext_reg[66]  ( .D(reg_out[66]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[66]) );
  DFFRNQ_X1 \Plaintext_reg[88]  ( .D(reg_out[88]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[88]) );
  DFFRNQ_X1 \Plaintext_reg[63]  ( .D(reg_out[63]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[63]) );
  DFFRNQ_X1 \Plaintext_reg[56]  ( .D(reg_out[56]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[56]) );
  DFFRNQ_X1 \Plaintext_reg[140]  ( .D(reg_out[140]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[140]) );
  DFFRNQ_X1 \Plaintext_reg[165]  ( .D(reg_out[165]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[165]) );
  DFFRNQ_X1 \Plaintext_reg[112]  ( .D(reg_out[112]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[112]) );
  DFFRNQ_X1 \Plaintext_reg[134]  ( .D(reg_out[134]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[134]) );
  DFFRNQ_X1 \Plaintext_reg[186]  ( .D(reg_out[186]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[186]) );
  DFFRNQ_X1 \Plaintext_reg[118]  ( .D(reg_out[118]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[118]) );
  DFFRNQ_X1 \Plaintext_reg[83]  ( .D(reg_out[83]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[83]) );
  DFFRNQ_X1 \Plaintext_reg[76]  ( .D(reg_out[76]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[76]) );
  DFFRNQ_X1 \Plaintext_reg[180]  ( .D(reg_out[180]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[180]) );
  DFFRNQ_X1 \Plaintext_reg[139]  ( .D(reg_out[139]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[139]) );
  DFFRNQ_X1 \Plaintext_reg[104]  ( .D(reg_out[104]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[104]) );
  DFFRNQ_X1 \Plaintext_reg[171]  ( .D(reg_out[171]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[171]) );
  DFFRNQ_X1 \Plaintext_reg[119]  ( .D(reg_out[119]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[119]) );
  DFFRNQ_X1 \Plaintext_reg[158]  ( .D(reg_out[158]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[158]) );
  DFFRNQ_X1 \Plaintext_reg[116]  ( .D(reg_out[116]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[116]) );
  DFFRNQ_X1 \Plaintext_reg[149]  ( .D(reg_out[149]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[149]) );
  DFFRNQ_X1 \Plaintext_reg[161]  ( .D(reg_out[161]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[161]) );
  DFFRNQ_X1 \Plaintext_reg[168]  ( .D(reg_out[168]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[168]) );
  DFFRNQ_X1 \Plaintext_reg[142]  ( .D(reg_out[142]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[142]) );
  DFFRNQ_X1 \Plaintext_reg[123]  ( .D(reg_out[123]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[123]) );
  DFFRNQ_X1 \Plaintext_reg[188]  ( .D(reg_out[188]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[188]) );
  DFFRNQ_X1 \Plaintext_reg[159]  ( .D(reg_out[159]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[159]) );
  DFFRNQ_X1 \Plaintext_reg[77]  ( .D(reg_out[77]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[77]) );
  DFFRNQ_X1 \Plaintext_reg[49]  ( .D(reg_out[49]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[49]) );
  DFFRNQ_X1 \Plaintext_reg[85]  ( .D(reg_out[85]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[85]) );
  DFFRNQ_X1 \Plaintext_reg[174]  ( .D(reg_out[174]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[174]) );
  DFFRNQ_X1 \Plaintext_reg[189]  ( .D(reg_out[189]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[189]) );
  DFFRNQ_X1 \Plaintext_reg[51]  ( .D(reg_out[51]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[51]) );
  DFFRNQ_X1 \Plaintext_reg[60]  ( .D(reg_out[60]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[60]) );
  DFFRNQ_X1 \Plaintext_reg[115]  ( .D(reg_out[115]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[115]) );
  DFFRNQ_X1 \Plaintext_reg[135]  ( .D(reg_out[135]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[135]) );
  DFFRNQ_X1 \Plaintext_reg[90]  ( .D(reg_out[90]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[90]) );
  DFFRNQ_X1 \Plaintext_reg[146]  ( .D(reg_out[146]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[146]) );
  DFFRNQ_X1 \Plaintext_reg[183]  ( .D(reg_out[183]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[183]) );
  DFFRNQ_X1 \Plaintext_reg[182]  ( .D(reg_out[182]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[182]) );
  DFFRNQ_X1 \Plaintext_reg[28]  ( .D(reg_out[28]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[28]) );
  DFFRNQ_X1 \Plaintext_reg[21]  ( .D(reg_out[21]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[21]) );
  DFFRNQ_X1 \Plaintext_reg[87]  ( .D(reg_out[87]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[87]) );
  DFFRNQ_X1 \Plaintext_reg[92]  ( .D(reg_out[92]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[92]) );
  DFFRNQ_X1 \Plaintext_reg[101]  ( .D(reg_out[101]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[101]) );
  DFFRNQ_X1 \Plaintext_reg[38]  ( .D(reg_out[38]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[38]) );
  DFFRNQ_X1 \Plaintext_reg[62]  ( .D(reg_out[62]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[62]) );
  DFFRNQ_X1 \Plaintext_reg[154]  ( .D(reg_out[154]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[154]) );
  DFFRNQ_X1 \Plaintext_reg[0]  ( .D(reg_out[0]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[0]) );
  DFFRNQ_X1 \Plaintext_reg[111]  ( .D(reg_out[111]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[111]) );
  DFFRNQ_X1 \Plaintext_reg[39]  ( .D(reg_out[39]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[39]) );
  DFFRNQ_X1 \Plaintext_reg[106]  ( .D(reg_out[106]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[106]) );
  DFFRNQ_X1 \Plaintext_reg[96]  ( .D(reg_out[96]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[96]) );
  DFFRNQ_X1 \Plaintext_reg[80]  ( .D(reg_out[80]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[80]) );
  DFFRNQ_X1 \Plaintext_reg[177]  ( .D(reg_out[177]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[177]) );
  DFFRNQ_X1 \Plaintext_reg[117]  ( .D(reg_out[117]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[117]) );
  DFFRNQ_X1 \Plaintext_reg[82]  ( .D(reg_out[82]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[82]) );
  DFFRNQ_X1 \Plaintext_reg[41]  ( .D(reg_out[41]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[41]) );
  DFFRNQ_X1 \Plaintext_reg[125]  ( .D(reg_out[125]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[125]) );
  DFFRNQ_X1 \Plaintext_reg[6]  ( .D(reg_out[6]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[6]) );
  DFFRNQ_X1 \Plaintext_reg[187]  ( .D(reg_out[187]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[187]) );
  DFFRNQ_X1 \Plaintext_reg[126]  ( .D(reg_out[126]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[126]) );
  DFFRNQ_X1 \Plaintext_reg[93]  ( .D(reg_out[93]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[93]) );
  DFFRNQ_X1 \Plaintext_reg[52]  ( .D(reg_out[52]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[52]) );
  DFFRNQ_X1 \Plaintext_reg[69]  ( .D(reg_out[69]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[69]) );
  DFFRNQ_X1 \Plaintext_reg[136]  ( .D(reg_out[136]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[136]) );
  DFFRNQ_X1 \Plaintext_reg[42]  ( .D(reg_out[42]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[42]) );
  DFFRNQ_X1 \Plaintext_reg[113]  ( .D(reg_out[113]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[113]) );
  DFFRNQ_X1 \Plaintext_reg[15]  ( .D(reg_out[15]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[15]) );
  DFFRNQ_X1 \Plaintext_reg[33]  ( .D(reg_out[33]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[33]) );
  DFFRNQ_X1 \Plaintext_reg[65]  ( .D(reg_out[65]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[65]) );
  DFFRNQ_X1 \Plaintext_reg[7]  ( .D(reg_out[7]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[7]) );
  DFFRNQ_X1 \Plaintext_reg[157]  ( .D(reg_out[157]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[157]) );
  DFFRNQ_X1 \Plaintext_reg[185]  ( .D(reg_out[185]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[185]) );
  DFFRNQ_X1 \Plaintext_reg[163]  ( .D(reg_out[163]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[163]) );
  DFFRNQ_X1 \Plaintext_reg[130]  ( .D(reg_out[130]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[130]) );
  DFFRNQ_X1 \Plaintext_reg[128]  ( .D(reg_out[128]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[128]) );
  DFFRNQ_X1 \Plaintext_reg[129]  ( .D(reg_out[129]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[129]) );
  DFFRNQ_X1 \Plaintext_reg[132]  ( .D(reg_out[132]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[132]) );
  DFFRNQ_X1 \Plaintext_reg[18]  ( .D(reg_out[18]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[18]) );
  DFFRNQ_X1 \Plaintext_reg[148]  ( .D(reg_out[148]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[148]) );
  DFFRNQ_X1 \Plaintext_reg[61]  ( .D(reg_out[61]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[61]) );
  DFFRNQ_X1 \Plaintext_reg[95]  ( .D(reg_out[95]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[95]) );
  DFFRNQ_X1 \Plaintext_reg[72]  ( .D(reg_out[72]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[72]) );
  DFFRNQ_X1 \Plaintext_reg[141]  ( .D(reg_out[141]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[141]) );
  DFFRNQ_X1 \Plaintext_reg[172]  ( .D(reg_out[172]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[172]) );
  DFFRNQ_X1 \Plaintext_reg[25]  ( .D(reg_out[25]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[25]) );
  DFFRNQ_X1 \Plaintext_reg[70]  ( .D(reg_out[70]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[70]) );
  DFFRNQ_X1 \Plaintext_reg[36]  ( .D(reg_out[36]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[36]) );
  DFFRNQ_X1 \Plaintext_reg[99]  ( .D(reg_out[99]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[99]) );
  DFFRNQ_X1 \Plaintext_reg[81]  ( .D(reg_out[81]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[81]) );
  DFFRNQ_X1 \Plaintext_reg[9]  ( .D(reg_out[9]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[9]) );
  DFFRNQ_X1 \Plaintext_reg[79]  ( .D(reg_out[79]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[79]) );
  DFFRNQ_X1 \Plaintext_reg[44]  ( .D(reg_out[44]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[44]) );
  DFFRNQ_X1 \Plaintext_reg[155]  ( .D(reg_out[155]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[155]) );
  DFFRNQ_X1 \Plaintext_reg[10]  ( .D(reg_out[10]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[10]) );
  DFFRNQ_X1 \Plaintext_reg[100]  ( .D(reg_out[100]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[100]) );
  DFFRNQ_X1 \Plaintext_reg[131]  ( .D(reg_out[131]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[131]) );
  DFFRNQ_X1 \Plaintext_reg[133]  ( .D(reg_out[133]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[133]) );
  DFFRNQ_X1 \Plaintext_reg[17]  ( .D(reg_out[17]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[17]) );
  DFFRNQ_X1 \Plaintext_reg[2]  ( .D(reg_out[2]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[2]) );
  DFFRNQ_X1 \Plaintext_reg[19]  ( .D(reg_out[19]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[19]) );
  DFFRNQ_X1 \Plaintext_reg[144]  ( .D(reg_out[144]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[144]) );
  DFFRNQ_X1 \Plaintext_reg[120]  ( .D(reg_out[120]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[120]) );
  DFFRNQ_X1 \Plaintext_reg[13]  ( .D(reg_out[13]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[13]) );
  DFFRNQ_X1 \Plaintext_reg[150]  ( .D(reg_out[150]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[150]) );
  DFFRNQ_X1 \Plaintext_reg[109]  ( .D(reg_out[109]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[109]) );
  DFFRNQ_X1 \Plaintext_reg[40]  ( .D(reg_out[40]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[40]) );
  DFFRNQ_X1 \Plaintext_reg[11]  ( .D(reg_out[11]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[11]) );
  DFFRNQ_X1 \Plaintext_reg[173]  ( .D(reg_out[173]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[173]) );
  DFFRNQ_X1 \Plaintext_reg[23]  ( .D(reg_out[23]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[23]) );
  DFFRNQ_X1 \Plaintext_reg[127]  ( .D(reg_out[127]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[127]) );
  DFFRNQ_X1 \Plaintext_reg[137]  ( .D(reg_out[137]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[137]) );
  DFFRNQ_X1 \Plaintext_reg[3]  ( .D(reg_out[3]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[3]) );
  DFFRNQ_X1 \Plaintext_reg[48]  ( .D(reg_out[48]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[48]) );
  DFFRNQ_X1 \Plaintext_reg[73]  ( .D(reg_out[73]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[73]) );
  DFFRNQ_X1 \Plaintext_reg[53]  ( .D(reg_out[53]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[53]) );
  DFFRNQ_X1 \Plaintext_reg[5]  ( .D(reg_out[5]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[5]) );
  DFFRNQ_X1 \Plaintext_reg[78]  ( .D(reg_out[78]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[78]) );
  DFFRNQ_X1 \Plaintext_reg[153]  ( .D(reg_out[153]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[153]) );
  DFFRNQ_X1 \Plaintext_reg[91]  ( .D(reg_out[91]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[91]) );
  DFFRNQ_X1 \Plaintext_reg[190]  ( .D(reg_out[190]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[190]) );
  DFFRNQ_X1 \Plaintext_reg[102]  ( .D(reg_out[102]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[102]) );
  DFFRNQ_X1 \Plaintext_reg[59]  ( .D(reg_out[59]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[59]) );
  DFFRNQ_X1 \Plaintext_reg[43]  ( .D(reg_out[43]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[43]) );
  DFFRNQ_X1 \Plaintext_reg[151]  ( .D(reg_out[151]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[151]) );
  DFFRNQ_X1 \Plaintext_reg[46]  ( .D(reg_out[46]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[46]) );
  DFFRNQ_X1 \Plaintext_reg[169]  ( .D(reg_out[169]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[169]) );
  DFFRNQ_X1 \Plaintext_reg[16]  ( .D(reg_out[16]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[16]) );
  DFFRNQ_X1 \Plaintext_reg[71]  ( .D(reg_out[71]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[71]) );
  DFFRNQ_X1 \Plaintext_reg[94]  ( .D(reg_out[94]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[94]) );
  DFFRNQ_X1 \Plaintext_reg[54]  ( .D(reg_out[54]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[54]) );
  DFFRNQ_X1 \Plaintext_reg[89]  ( .D(reg_out[89]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[89]) );
  DFFRNQ_X1 \Plaintext_reg[160]  ( .D(reg_out[160]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[160]) );
  DFFRNQ_X1 \Plaintext_reg[105]  ( .D(reg_out[105]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[105]) );
  DFFRNQ_X1 \Plaintext_reg[4]  ( .D(reg_out[4]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[4]) );
  DFFRNQ_X1 \Plaintext_reg[12]  ( .D(reg_out[12]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[12]) );
  DFFRNQ_X1 \Plaintext_reg[178]  ( .D(reg_out[178]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[178]) );
  DFFRNQ_X1 \Plaintext_reg[145]  ( .D(reg_out[145]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[145]) );
  DFFRNQ_X1 \Plaintext_reg[147]  ( .D(reg_out[147]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[147]) );
  DFFRNQ_X1 \Plaintext_reg[179]  ( .D(reg_out[179]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[179]) );
  DFFRNQ_X1 \Plaintext_reg[121]  ( .D(reg_out[121]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[121]) );
  DFFRNQ_X1 \Plaintext_reg[181]  ( .D(reg_out[181]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[181]) );
  DFFRNQ_X1 \Plaintext_reg[97]  ( .D(reg_out[97]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[97]) );
  DFFRNQ_X1 \Plaintext_reg[191]  ( .D(reg_out[191]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[191]) );
  DFFRNQ_X1 \Plaintext_reg[156]  ( .D(reg_out[156]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[156]) );
  DFFRNQ_X1 \Plaintext_reg[67]  ( .D(reg_out[67]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[67]) );
  DFFRNQ_X1 \Plaintext_reg[175]  ( .D(reg_out[175]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[175]) );
  DFFRNQ_X1 \Plaintext_reg[45]  ( .D(reg_out[45]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[45]) );
  DFFRNQ_X1 \Plaintext_reg[143]  ( .D(reg_out[143]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[143]) );
  DFFRNQ_X1 \Plaintext_reg[103]  ( .D(reg_out[103]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[103]) );
  DFFRNQ_X1 \Plaintext_reg[107]  ( .D(reg_out[107]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[107]) );
  DFFRNQ_X1 \Plaintext_reg[1]  ( .D(reg_out[1]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[1]) );
  DFFRNQ_X1 \Plaintext_reg[47]  ( .D(reg_out[47]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[47]) );
  DFFRNQ_X1 \Plaintext_reg[55]  ( .D(reg_out[55]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[55]) );
  DFFRNQ_X1 \reg_in_reg[150]  ( .D(Ciphertext[150]), .CLK(clk), .RN(1'b1), .Q(
        reg_in[150]) );
  DFFRNQ_X1 \Plaintext_reg[37]  ( .D(reg_out[37]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[37]) );
  DFFRNQ_X1 \reg_in_reg[158]  ( .D(Ciphertext[158]), .CLK(clk), .RN(1'b1), .Q(
        reg_in[158]) );
  DFFRNQ_X1 \reg_in_reg[78]  ( .D(Ciphertext[78]), .CLK(clk), .RN(1'b1), .Q(
        reg_in[78]) );
  DFFRNQ_X1 \reg_in_reg[165]  ( .D(Ciphertext[165]), .CLK(clk), .RN(1'b1), .Q(
        reg_in[165]) );
  SPEEDY_Rounds5_0 SPEEDY_instance ( .Ciphertext(reg_in), .Key(reg_key), 
        .Plaintext(reg_out) );
  DFFRNQ_X1 \reg_key_reg[131]  ( .D(Key[131]), .CLK(clk), .RN(1'b1), .Q(
        reg_key[131]) );
  DFFSNQ_X1 \Plaintext_reg[162]  ( .D(reg_out[162]), .CLK(clk), .SN(1'b1), .Q(
        Plaintext[162]) );
  DFFSNQ_X1 \Plaintext_reg[20]  ( .D(reg_out[20]), .CLK(clk), .SN(1'b1), .Q(
        Plaintext[20]) );
  DFFRNQ_X1 \Plaintext_reg[184]  ( .D(reg_out[184]), .CLK(clk), .RN(1'b1), .Q(
        Plaintext[184]) );
  DFFRNQ_X1 \reg_key_reg[118]  ( .D(Key[118]), .CLK(clk), .RN(1'b1), .Q(
        reg_key[118]) );
  DFFRNQ_X1 \reg_in_reg[51]  ( .D(Ciphertext[51]), .CLK(clk), .RN(1'b1), .Q(
        reg_in[51]) );
endmodule

