library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity SB is
    Port ( input : in STD_LOGIC_VECTOR (5 downto 0);
           output : out STD_LOGIC_VECTOR (5 downto 0));
end SB;

architecture Behavioral of SB is

begin

    with input select
    output <= "000001" when "000000",
              "001101" when "000001",
              "100000" when "000010",
              "000011" when "000011",
              "001010" when "000100",
              "011101" when "000101",
              "100001" when "000110",
              "001011" when "000111",
              "000000" when "001000",
              "000010" when "001001",
              "101000" when "001010",
              "100010" when "001011",
              "001000" when "001100",
              "001001" when "001101",
              "101010" when "001110",
              "100011" when "001111",
              "000101" when "010000",
              "101101" when "010001",
              "010001" when "010010",
              "000111" when "010011",
              "011010" when "010100",
              "100111" when "010101",
              "010101" when "010110",
              "100101" when "010111",
              "010010" when "011000",
              "111101" when "011001",
              "010000" when "011010",
              "101001" when "011011",
              "011000" when "011100",
              "011001" when "011101",
              "110101" when "011110",
              "101011" when "011111",
              "001110" when "100000",
              "100110" when "100001",
              "110000" when "100010",
              "001111" when "100011",
              "011110" when "100100",
              "101110" when "100101",
              "110001" when "100110",
              "011111" when "100111",
              "110110" when "101000",
              "000110" when "101001",
              "110010" when "101010",
              "111000" when "101011",
              "010110" when "101100",
              "111110" when "101101",
              "110011" when "101110",
              "111010" when "101111",
              "001100" when "110000",
              "101100" when "110001",
              "010011" when "110010",
              "100100" when "110011",
              "011100" when "110100",
              "101111" when "110101",
              "010111" when "110110",
              "011011" when "110111",
              "000100" when "111000",
              "111100" when "111001",
              "110100" when "111010",
              "111001" when "111011",
              "110111" when "111100",
              "111111" when "111101",
              "010100" when "111110",
              "111011" when others;

end Behavioral;