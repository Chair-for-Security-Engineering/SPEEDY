module SPEEDY_Rounds5_0 ( Plaintext, Key, Ciphertext );
  input [191:0] Plaintext;
  input [191:0] Key;
  output [191:0] Ciphertext;
  wire   \RI1[1][173] , \RI1[1][143] , \RI1[1][71] , \RI1[1][59] ,
         \RI1[1][11] , \RI1[2][167] , \RI1[2][95] , \RI1[2][59] , \RI1[2][47] ,
         \RI1[2][35] , \RI1[2][17] , \RI1[3][167] , \RI1[3][143] ,
         \RI1[3][131] , \RI1[3][89] , \RI1[3][71] , \RI1[3][59] , \RI1[3][41] ,
         \RI1[3][14] , \RI1[3][5] , \RI1[4][179] , \RI1[4][155] ,
         \RI1[4][154] , \RI1[4][143] , \RI1[4][131] , \RI1[4][89] ,
         \RI1[4][87] , \RI1[4][77] , \RI1[4][65] , \RI1[4][59] , \RI1[4][53] ,
         \RI1[4][41] , \RI1[4][29] , \RI1[4][5] , \RI3[0][191] , \RI3[0][190] ,
         \RI3[0][188] , \RI3[0][183] , \RI3[0][182] , \RI3[0][180] ,
         \RI3[0][179] , \RI3[0][178] , \RI3[0][176] , \RI3[0][175] ,
         \RI3[0][172] , \RI3[0][166] , \RI3[0][165] , \RI3[0][164] ,
         \RI3[0][163] , \RI3[0][162] , \RI3[0][161] , \RI3[0][160] ,
         \RI3[0][156] , \RI3[0][155] , \RI3[0][154] , \RI3[0][152] ,
         \RI3[0][149] , \RI3[0][147] , \RI3[0][146] , \RI3[0][142] ,
         \RI3[0][139] , \RI3[0][134] , \RI3[0][131] , \RI3[0][129] ,
         \RI3[0][127] , \RI3[0][126] , \RI3[0][123] , \RI3[0][121] ,
         \RI3[0][118] , \RI3[0][116] , \RI3[0][114] , \RI3[0][113] ,
         \RI3[0][107] , \RI3[0][106] , \RI3[0][105] , \RI3[0][104] ,
         \RI3[0][103] , \RI3[0][100] , \RI3[0][99] , \RI3[0][97] ,
         \RI3[0][96] , \RI3[0][95] , \RI3[0][93] , \RI3[0][92] , \RI3[0][91] ,
         \RI3[0][88] , \RI3[0][86] , \RI3[0][84] , \RI3[0][82] , \RI3[0][81] ,
         \RI3[0][80] , \RI3[0][79] , \RI3[0][76] , \RI3[0][72] , \RI3[0][69] ,
         \RI3[0][68] , \RI3[0][67] , \RI3[0][66] , \RI3[0][63] , \RI3[0][62] ,
         \RI3[0][61] , \RI3[0][58] , \RI3[0][57] , \RI3[0][55] , \RI3[0][54] ,
         \RI3[0][50] , \RI3[0][49] , \RI3[0][48] , \RI3[0][46] , \RI3[0][45] ,
         \RI3[0][44] , \RI3[0][43] , \RI3[0][40] , \RI3[0][39] , \RI3[0][37] ,
         \RI3[0][34] , \RI3[0][33] , \RI3[0][32] , \RI3[0][30] , \RI3[0][27] ,
         \RI3[0][23] , \RI3[0][22] , \RI3[0][20] , \RI3[0][18] , \RI3[0][15] ,
         \RI3[0][10] , \RI3[0][9] , \RI3[0][8] , \RI3[0][7] , \RI3[0][5] ,
         \RI3[0][4] , \RI3[0][3] , \RI3[0][2] , \RI3[0][1] , \RI3[1][182] ,
         \RI3[1][110] , \RI3[1][60] , \RI3[3][35] , \RI3[3][24] , \RI3[3][16] ,
         \RI3[4][105] , \RI3[4][23] , \RI5[0][191] , \RI5[0][190] ,
         \RI5[0][189] , \RI5[0][188] , \RI5[0][187] , \RI5[0][186] ,
         \RI5[0][185] , \RI5[0][184] , \RI5[0][183] , \RI5[0][182] ,
         \RI5[0][181] , \RI5[0][178] , \RI5[0][177] , \RI5[0][176] ,
         \RI5[0][175] , \RI5[0][174] , \RI5[0][173] , \RI5[0][172] ,
         \RI5[0][171] , \RI5[0][170] , \RI5[0][169] , \RI5[0][168] ,
         \RI5[0][164] , \RI5[0][163] , \RI5[0][162] , \RI5[0][161] ,
         \RI5[0][160] , \RI5[0][159] , \RI5[0][158] , \RI5[0][154] ,
         \RI5[0][153] , \RI5[0][152] , \RI5[0][151] , \RI5[0][149] ,
         \RI5[0][148] , \RI5[0][147] , \RI5[0][146] , \RI5[0][145] ,
         \RI5[0][143] , \RI5[0][142] , \RI5[0][140] , \RI5[0][139] ,
         \RI5[0][137] , \RI5[0][136] , \RI5[0][135] , \RI5[0][134] ,
         \RI5[0][133] , \RI5[0][131] , \RI5[0][130] , \RI5[0][129] ,
         \RI5[0][128] , \RI5[0][127] , \RI5[0][126] , \RI5[0][125] ,
         \RI5[0][124] , \RI5[0][123] , \RI5[0][122] , \RI5[0][121] ,
         \RI5[0][120] , \RI5[0][119] , \RI5[0][118] , \RI5[0][117] ,
         \RI5[0][116] , \RI5[0][114] , \RI5[0][113] , \RI5[0][111] ,
         \RI5[0][110] , \RI5[0][108] , \RI5[0][107] , \RI5[0][106] ,
         \RI5[0][104] , \RI5[0][103] , \RI5[0][102] , \RI5[0][101] ,
         \RI5[0][100] , \RI5[0][99] , \RI5[0][98] , \RI5[0][97] , \RI5[0][95] ,
         \RI5[0][94] , \RI5[0][93] , \RI5[0][91] , \RI5[0][89] , \RI5[0][87] ,
         \RI5[0][85] , \RI5[0][84] , \RI5[0][83] , \RI5[0][80] , \RI5[0][77] ,
         \RI5[0][75] , \RI5[0][74] , \RI5[0][72] , \RI5[0][71] , \RI5[0][70] ,
         \RI5[0][68] , \RI5[0][66] , \RI5[0][65] , \RI5[0][64] , \RI5[0][63] ,
         \RI5[0][62] , \RI5[0][60] , \RI5[0][59] , \RI5[0][58] , \RI5[0][57] ,
         \RI5[0][55] , \RI5[0][54] , \RI5[0][53] , \RI5[0][52] , \RI5[0][50] ,
         \RI5[0][47] , \RI5[0][45] , \RI5[0][43] , \RI5[0][41] , \RI5[0][40] ,
         \RI5[0][39] , \RI5[0][38] , \RI5[0][37] , \RI5[0][35] , \RI5[0][34] ,
         \RI5[0][33] , \RI5[0][32] , \RI5[0][31] , \RI5[0][30] , \RI5[0][29] ,
         \RI5[0][28] , \RI5[0][27] , \RI5[0][26] , \RI5[0][25] , \RI5[0][24] ,
         \RI5[0][23] , \RI5[0][20] , \RI5[0][19] , \RI5[0][18] , \RI5[0][17] ,
         \RI5[0][16] , \RI5[0][15] , \RI5[0][14] , \RI5[0][13] , \RI5[0][11] ,
         \RI5[0][10] , \RI5[0][9] , \RI5[0][8] , \RI5[0][6] , \RI5[0][5] ,
         \RI5[0][4] , \RI5[0][3] , \RI5[0][1] , \RI5[0][0] , \RI5[1][191] ,
         \RI5[1][190] , \RI5[1][189] , \RI5[1][188] , \RI5[1][184] ,
         \RI5[1][183] , \RI5[1][182] , \RI5[1][181] , \RI5[1][180] ,
         \RI5[1][178] , \RI5[1][177] , \RI5[1][176] , \RI5[1][175] ,
         \RI5[1][174] , \RI5[1][173] , \RI5[1][172] , \RI5[1][171] ,
         \RI5[1][168] , \RI5[1][167] , \RI5[1][166] , \RI5[1][165] ,
         \RI5[1][164] , \RI5[1][162] , \RI5[1][161] , \RI5[1][158] ,
         \RI5[1][157] , \RI5[1][156] , \RI5[1][154] , \RI5[1][152] ,
         \RI5[1][151] , \RI5[1][150] , \RI5[1][149] , \RI5[1][148] ,
         \RI5[1][147] , \RI5[1][146] , \RI5[1][145] , \RI5[1][144] ,
         \RI5[1][143] , \RI5[1][142] , \RI5[1][141] , \RI5[1][140] ,
         \RI5[1][138] , \RI5[1][137] , \RI5[1][136] , \RI5[1][135] ,
         \RI5[1][134] , \RI5[1][133] , \RI5[1][132] , \RI5[1][131] ,
         \RI5[1][130] , \RI5[1][129] , \RI5[1][128] , \RI5[1][127] ,
         \RI5[1][126] , \RI5[1][125] , \RI5[1][124] , \RI5[1][122] ,
         \RI5[1][121] , \RI5[1][120] , \RI5[1][119] , \RI5[1][118] ,
         \RI5[1][117] , \RI5[1][116] , \RI5[1][115] , \RI5[1][114] ,
         \RI5[1][113] , \RI5[1][112] , \RI5[1][111] , \RI5[1][109] ,
         \RI5[1][108] , \RI5[1][107] , \RI5[1][106] , \RI5[1][104] ,
         \RI5[1][103] , \RI5[1][102] , \RI5[1][98] , \RI5[1][97] ,
         \RI5[1][96] , \RI5[1][94] , \RI5[1][93] , \RI5[1][92] , \RI5[1][91] ,
         \RI5[1][90] , \RI5[1][88] , \RI5[1][87] , \RI5[1][86] , \RI5[1][85] ,
         \RI5[1][83] , \RI5[1][82] , \RI5[1][81] , \RI5[1][79] , \RI5[1][78] ,
         \RI5[1][77] , \RI5[1][76] , \RI5[1][75] , \RI5[1][73] , \RI5[1][72] ,
         \RI5[1][71] , \RI5[1][70] , \RI5[1][69] , \RI5[1][68] , \RI5[1][67] ,
         \RI5[1][65] , \RI5[1][64] , \RI5[1][62] , \RI5[1][61] , \RI5[1][60] ,
         \RI5[1][59] , \RI5[1][58] , \RI5[1][57] , \RI5[1][56] , \RI5[1][55] ,
         \RI5[1][54] , \RI5[1][53] , \RI5[1][52] , \RI5[1][51] , \RI5[1][50] ,
         \RI5[1][49] , \RI5[1][48] , \RI5[1][47] , \RI5[1][46] , \RI5[1][45] ,
         \RI5[1][44] , \RI5[1][43] , \RI5[1][40] , \RI5[1][39] , \RI5[1][37] ,
         \RI5[1][36] , \RI5[1][34] , \RI5[1][32] , \RI5[1][30] , \RI5[1][27] ,
         \RI5[1][26] , \RI5[1][24] , \RI5[1][23] , \RI5[1][21] , \RI5[1][20] ,
         \RI5[1][19] , \RI5[1][18] , \RI5[1][17] , \RI5[1][16] , \RI5[1][15] ,
         \RI5[1][14] , \RI5[1][13] , \RI5[1][12] , \RI5[1][11] , \RI5[1][10] ,
         \RI5[1][8] , \RI5[1][7] , \RI5[1][6] , \RI5[1][5] , \RI5[1][4] ,
         \RI5[1][3] , \RI5[1][2] , \RI5[1][0] , \RI5[2][191] , \RI5[2][190] ,
         \RI5[2][189] , \RI5[2][188] , \RI5[2][187] , \RI5[2][184] ,
         \RI5[2][181] , \RI5[2][180] , \RI5[2][179] , \RI5[2][178] ,
         \RI5[2][176] , \RI5[2][174] , \RI5[2][173] , \RI5[2][172] ,
         \RI5[2][171] , \RI5[2][170] , \RI5[2][169] , \RI5[2][168] ,
         \RI5[2][167] , \RI5[2][166] , \RI5[2][165] , \RI5[2][164] ,
         \RI5[2][163] , \RI5[2][161] , \RI5[2][160] , \RI5[2][159] ,
         \RI5[2][157] , \RI5[2][155] , \RI5[2][154] , \RI5[2][152] ,
         \RI5[2][150] , \RI5[2][147] , \RI5[2][145] , \RI5[2][144] ,
         \RI5[2][143] , \RI5[2][142] , \RI5[2][140] , \RI5[2][139] ,
         \RI5[2][138] , \RI5[2][137] , \RI5[2][135] , \RI5[2][134] ,
         \RI5[2][130] , \RI5[2][126] , \RI5[2][123] , \RI5[2][121] ,
         \RI5[2][120] , \RI5[2][119] , \RI5[2][118] , \RI5[2][114] ,
         \RI5[2][113] , \RI5[2][112] , \RI5[2][111] , \RI5[2][110] ,
         \RI5[2][109] , \RI5[2][108] , \RI5[2][107] , \RI5[2][104] ,
         \RI5[2][103] , \RI5[2][102] , \RI5[2][101] , \RI5[2][100] ,
         \RI5[2][98] , \RI5[2][96] , \RI5[2][94] , \RI5[2][93] , \RI5[2][91] ,
         \RI5[2][90] , \RI5[2][89] , \RI5[2][88] , \RI5[2][87] , \RI5[2][85] ,
         \RI5[2][84] , \RI5[2][80] , \RI5[2][79] , \RI5[2][77] , \RI5[2][75] ,
         \RI5[2][73] , \RI5[2][72] , \RI5[2][71] , \RI5[2][69] , \RI5[2][67] ,
         \RI5[2][66] , \RI5[2][64] , \RI5[2][63] , \RI5[2][62] , \RI5[2][60] ,
         \RI5[2][57] , \RI5[2][55] , \RI5[2][54] , \RI5[2][52] , \RI5[2][51] ,
         \RI5[2][48] , \RI5[2][46] , \RI5[2][44] , \RI5[2][42] , \RI5[2][41] ,
         \RI5[2][40] , \RI5[2][37] , \RI5[2][35] , \RI5[2][33] , \RI5[2][32] ,
         \RI5[2][31] , \RI5[2][28] , \RI5[2][26] , \RI5[2][25] , \RI5[2][24] ,
         \RI5[2][23] , \RI5[2][22] , \RI5[2][21] , \RI5[2][20] , \RI5[2][19] ,
         \RI5[2][18] , \RI5[2][17] , \RI5[2][16] , \RI5[2][15] , \RI5[2][13] ,
         \RI5[2][12] , \RI5[2][11] , \RI5[2][10] , \RI5[2][9] , \RI5[2][8] ,
         \RI5[2][5] , \RI5[2][3] , \RI5[2][1] , \RI5[3][190] , \RI5[3][189] ,
         \RI5[3][188] , \RI5[3][187] , \RI5[3][186] , \RI5[3][185] ,
         \RI5[3][184] , \RI5[3][183] , \RI5[3][181] , \RI5[3][180] ,
         \RI5[3][177] , \RI5[3][175] , \RI5[3][173] , \RI5[3][172] ,
         \RI5[3][171] , \RI5[3][170] , \RI5[3][169] , \RI5[3][164] ,
         \RI5[3][163] , \RI5[3][162] , \RI5[3][161] , \RI5[3][160] ,
         \RI5[3][159] , \RI5[3][158] , \RI5[3][157] , \RI5[3][156] ,
         \RI5[3][153] , \RI5[3][151] , \RI5[3][150] , \RI5[3][149] ,
         \RI5[3][148] , \RI5[3][147] , \RI5[3][146] , \RI5[3][145] ,
         \RI5[3][144] , \RI5[3][143] , \RI5[3][141] , \RI5[3][140] ,
         \RI5[3][139] , \RI5[3][138] , \RI5[3][137] , \RI5[3][136] ,
         \RI5[3][134] , \RI5[3][133] , \RI5[3][131] , \RI5[3][130] ,
         \RI5[3][129] , \RI5[3][128] , \RI5[3][127] , \RI5[3][126] ,
         \RI5[3][125] , \RI5[3][124] , \RI5[3][123] , \RI5[3][121] ,
         \RI5[3][120] , \RI5[3][118] , \RI5[3][117] , \RI5[3][113] ,
         \RI5[3][112] , \RI5[3][108] , \RI5[3][107] , \RI5[3][106] ,
         \RI5[3][105] , \RI5[3][102] , \RI5[3][100] , \RI5[3][99] ,
         \RI5[3][98] , \RI5[3][96] , \RI5[3][95] , \RI5[3][94] , \RI5[3][93] ,
         \RI5[3][92] , \RI5[3][89] , \RI5[3][88] , \RI5[3][87] , \RI5[3][86] ,
         \RI5[3][85] , \RI5[3][84] , \RI5[3][83] , \RI5[3][80] , \RI5[3][79] ,
         \RI5[3][78] , \RI5[3][77] , \RI5[3][76] , \RI5[3][75] , \RI5[3][73] ,
         \RI5[3][72] , \RI5[3][70] , \RI5[3][69] , \RI5[3][68] , \RI5[3][67] ,
         \RI5[3][66] , \RI5[3][65] , \RI5[3][64] , \RI5[3][63] , \RI5[3][62] ,
         \RI5[3][61] , \RI5[3][60] , \RI5[3][59] , \RI5[3][58] , \RI5[3][57] ,
         \RI5[3][55] , \RI5[3][54] , \RI5[3][52] , \RI5[3][50] , \RI5[3][48] ,
         \RI5[3][47] , \RI5[3][46] , \RI5[3][45] , \RI5[3][43] , \RI5[3][42] ,
         \RI5[3][39] , \RI5[3][37] , \RI5[3][35] , \RI5[3][34] , \RI5[3][33] ,
         \RI5[3][32] , \RI5[3][31] , \RI5[3][30] , \RI5[3][29] , \RI5[3][27] ,
         \RI5[3][26] , \RI5[3][25] , \RI5[3][24] , \RI5[3][23] , \RI5[3][21] ,
         \RI5[3][20] , \RI5[3][19] , \RI5[3][18] , \RI5[3][16] , \RI5[3][15] ,
         \RI5[3][13] , \RI5[3][11] , \RI5[3][10] , \RI5[3][9] , \RI5[3][8] ,
         \RI5[3][7] , \RI5[3][4] , \RI5[3][3] , \RI5[3][2] , \RI5[3][1] ,
         \RI5[3][0] , \MC_ARK_ARC_1_0/buf_output[191] ,
         \MC_ARK_ARC_1_0/buf_output[190] , \MC_ARK_ARC_1_0/buf_output[189] ,
         \MC_ARK_ARC_1_0/buf_output[188] , \MC_ARK_ARC_1_0/buf_output[187] ,
         \MC_ARK_ARC_1_0/buf_output[186] , \MC_ARK_ARC_1_0/buf_output[185] ,
         \MC_ARK_ARC_1_0/buf_output[184] , \MC_ARK_ARC_1_0/buf_output[183] ,
         \MC_ARK_ARC_1_0/buf_output[182] , \MC_ARK_ARC_1_0/buf_output[181] ,
         \MC_ARK_ARC_1_0/buf_output[180] , \MC_ARK_ARC_1_0/buf_output[179] ,
         \MC_ARK_ARC_1_0/buf_output[178] , \MC_ARK_ARC_1_0/buf_output[177] ,
         \MC_ARK_ARC_1_0/buf_output[176] , \MC_ARK_ARC_1_0/buf_output[175] ,
         \MC_ARK_ARC_1_0/buf_output[174] , \MC_ARK_ARC_1_0/buf_output[172] ,
         \MC_ARK_ARC_1_0/buf_output[171] , \MC_ARK_ARC_1_0/buf_output[170] ,
         \MC_ARK_ARC_1_0/buf_output[169] , \MC_ARK_ARC_1_0/buf_output[168] ,
         \MC_ARK_ARC_1_0/buf_output[167] , \MC_ARK_ARC_1_0/buf_output[166] ,
         \MC_ARK_ARC_1_0/buf_output[165] , \MC_ARK_ARC_1_0/buf_output[164] ,
         \MC_ARK_ARC_1_0/buf_output[163] , \MC_ARK_ARC_1_0/buf_output[162] ,
         \MC_ARK_ARC_1_0/buf_output[161] , \MC_ARK_ARC_1_0/buf_output[160] ,
         \MC_ARK_ARC_1_0/buf_output[159] , \MC_ARK_ARC_1_0/buf_output[158] ,
         \MC_ARK_ARC_1_0/buf_output[157] , \MC_ARK_ARC_1_0/buf_output[156] ,
         \MC_ARK_ARC_1_0/buf_output[155] , \MC_ARK_ARC_1_0/buf_output[154] ,
         \MC_ARK_ARC_1_0/buf_output[153] , \MC_ARK_ARC_1_0/buf_output[152] ,
         \MC_ARK_ARC_1_0/buf_output[151] , \MC_ARK_ARC_1_0/buf_output[150] ,
         \MC_ARK_ARC_1_0/buf_output[149] , \MC_ARK_ARC_1_0/buf_output[148] ,
         \MC_ARK_ARC_1_0/buf_output[147] , \MC_ARK_ARC_1_0/buf_output[146] ,
         \MC_ARK_ARC_1_0/buf_output[145] , \MC_ARK_ARC_1_0/buf_output[144] ,
         \MC_ARK_ARC_1_0/buf_output[143] , \MC_ARK_ARC_1_0/buf_output[142] ,
         \MC_ARK_ARC_1_0/buf_output[141] , \MC_ARK_ARC_1_0/buf_output[140] ,
         \MC_ARK_ARC_1_0/buf_output[139] , \MC_ARK_ARC_1_0/buf_output[138] ,
         \MC_ARK_ARC_1_0/buf_output[137] , \MC_ARK_ARC_1_0/buf_output[136] ,
         \MC_ARK_ARC_1_0/buf_output[135] , \MC_ARK_ARC_1_0/buf_output[134] ,
         \MC_ARK_ARC_1_0/buf_output[133] , \MC_ARK_ARC_1_0/buf_output[132] ,
         \MC_ARK_ARC_1_0/buf_output[131] , \MC_ARK_ARC_1_0/buf_output[130] ,
         \MC_ARK_ARC_1_0/buf_output[129] , \MC_ARK_ARC_1_0/buf_output[128] ,
         \MC_ARK_ARC_1_0/buf_output[127] , \MC_ARK_ARC_1_0/buf_output[126] ,
         \MC_ARK_ARC_1_0/buf_output[125] , \MC_ARK_ARC_1_0/buf_output[124] ,
         \MC_ARK_ARC_1_0/buf_output[123] , \MC_ARK_ARC_1_0/buf_output[122] ,
         \MC_ARK_ARC_1_0/buf_output[121] , \MC_ARK_ARC_1_0/buf_output[120] ,
         \MC_ARK_ARC_1_0/buf_output[119] , \MC_ARK_ARC_1_0/buf_output[118] ,
         \MC_ARK_ARC_1_0/buf_output[117] , \MC_ARK_ARC_1_0/buf_output[116] ,
         \MC_ARK_ARC_1_0/buf_output[115] , \MC_ARK_ARC_1_0/buf_output[114] ,
         \MC_ARK_ARC_1_0/buf_output[113] , \MC_ARK_ARC_1_0/buf_output[112] ,
         \MC_ARK_ARC_1_0/buf_output[111] , \MC_ARK_ARC_1_0/buf_output[110] ,
         \MC_ARK_ARC_1_0/buf_output[109] , \MC_ARK_ARC_1_0/buf_output[108] ,
         \MC_ARK_ARC_1_0/buf_output[107] , \MC_ARK_ARC_1_0/buf_output[106] ,
         \MC_ARK_ARC_1_0/buf_output[105] , \MC_ARK_ARC_1_0/buf_output[104] ,
         \MC_ARK_ARC_1_0/buf_output[103] , \MC_ARK_ARC_1_0/buf_output[102] ,
         \MC_ARK_ARC_1_0/buf_output[101] , \MC_ARK_ARC_1_0/buf_output[100] ,
         \MC_ARK_ARC_1_0/buf_output[99] , \MC_ARK_ARC_1_0/buf_output[98] ,
         \MC_ARK_ARC_1_0/buf_output[97] , \MC_ARK_ARC_1_0/buf_output[96] ,
         \MC_ARK_ARC_1_0/buf_output[95] , \MC_ARK_ARC_1_0/buf_output[94] ,
         \MC_ARK_ARC_1_0/buf_output[93] , \MC_ARK_ARC_1_0/buf_output[92] ,
         \MC_ARK_ARC_1_0/buf_output[91] , \MC_ARK_ARC_1_0/buf_output[90] ,
         \MC_ARK_ARC_1_0/buf_output[89] , \MC_ARK_ARC_1_0/buf_output[88] ,
         \MC_ARK_ARC_1_0/buf_output[87] , \MC_ARK_ARC_1_0/buf_output[86] ,
         \MC_ARK_ARC_1_0/buf_output[85] , \MC_ARK_ARC_1_0/buf_output[84] ,
         \MC_ARK_ARC_1_0/buf_output[83] , \MC_ARK_ARC_1_0/buf_output[82] ,
         \MC_ARK_ARC_1_0/buf_output[81] , \MC_ARK_ARC_1_0/buf_output[80] ,
         \MC_ARK_ARC_1_0/buf_output[79] , \MC_ARK_ARC_1_0/buf_output[78] ,
         \MC_ARK_ARC_1_0/buf_output[77] , \MC_ARK_ARC_1_0/buf_output[76] ,
         \MC_ARK_ARC_1_0/buf_output[75] , \MC_ARK_ARC_1_0/buf_output[74] ,
         \MC_ARK_ARC_1_0/buf_output[73] , \MC_ARK_ARC_1_0/buf_output[72] ,
         \MC_ARK_ARC_1_0/buf_output[70] , \MC_ARK_ARC_1_0/buf_output[69] ,
         \MC_ARK_ARC_1_0/buf_output[68] , \MC_ARK_ARC_1_0/buf_output[67] ,
         \MC_ARK_ARC_1_0/buf_output[66] , \MC_ARK_ARC_1_0/buf_output[65] ,
         \MC_ARK_ARC_1_0/buf_output[64] , \MC_ARK_ARC_1_0/buf_output[63] ,
         \MC_ARK_ARC_1_0/buf_output[62] , \MC_ARK_ARC_1_0/buf_output[61] ,
         \MC_ARK_ARC_1_0/buf_output[60] , \MC_ARK_ARC_1_0/buf_output[59] ,
         \MC_ARK_ARC_1_0/buf_output[58] , \MC_ARK_ARC_1_0/buf_output[57] ,
         \MC_ARK_ARC_1_0/buf_output[56] , \MC_ARK_ARC_1_0/buf_output[55] ,
         \MC_ARK_ARC_1_0/buf_output[54] , \MC_ARK_ARC_1_0/buf_output[53] ,
         \MC_ARK_ARC_1_0/buf_output[52] , \MC_ARK_ARC_1_0/buf_output[51] ,
         \MC_ARK_ARC_1_0/buf_output[50] , \MC_ARK_ARC_1_0/buf_output[49] ,
         \MC_ARK_ARC_1_0/buf_output[48] , \MC_ARK_ARC_1_0/buf_output[47] ,
         \MC_ARK_ARC_1_0/buf_output[46] , \MC_ARK_ARC_1_0/buf_output[45] ,
         \MC_ARK_ARC_1_0/buf_output[44] , \MC_ARK_ARC_1_0/buf_output[43] ,
         \MC_ARK_ARC_1_0/buf_output[42] , \MC_ARK_ARC_1_0/buf_output[41] ,
         \MC_ARK_ARC_1_0/buf_output[40] , \MC_ARK_ARC_1_0/buf_output[39] ,
         \MC_ARK_ARC_1_0/buf_output[38] , \MC_ARK_ARC_1_0/buf_output[37] ,
         \MC_ARK_ARC_1_0/buf_output[36] , \MC_ARK_ARC_1_0/buf_output[35] ,
         \MC_ARK_ARC_1_0/buf_output[34] , \MC_ARK_ARC_1_0/buf_output[33] ,
         \MC_ARK_ARC_1_0/buf_output[32] , \MC_ARK_ARC_1_0/buf_output[31] ,
         \MC_ARK_ARC_1_0/buf_output[30] , \MC_ARK_ARC_1_0/buf_output[29] ,
         \MC_ARK_ARC_1_0/buf_output[28] , \MC_ARK_ARC_1_0/buf_output[27] ,
         \MC_ARK_ARC_1_0/buf_output[26] , \MC_ARK_ARC_1_0/buf_output[25] ,
         \MC_ARK_ARC_1_0/buf_output[24] , \MC_ARK_ARC_1_0/buf_output[23] ,
         \MC_ARK_ARC_1_0/buf_output[22] , \MC_ARK_ARC_1_0/buf_output[21] ,
         \MC_ARK_ARC_1_0/buf_output[20] , \MC_ARK_ARC_1_0/buf_output[19] ,
         \MC_ARK_ARC_1_0/buf_output[18] , \MC_ARK_ARC_1_0/buf_output[17] ,
         \MC_ARK_ARC_1_0/buf_output[16] , \MC_ARK_ARC_1_0/buf_output[15] ,
         \MC_ARK_ARC_1_0/buf_output[14] , \MC_ARK_ARC_1_0/buf_output[13] ,
         \MC_ARK_ARC_1_0/buf_output[12] , \MC_ARK_ARC_1_0/buf_output[10] ,
         \MC_ARK_ARC_1_0/buf_output[9] , \MC_ARK_ARC_1_0/buf_output[8] ,
         \MC_ARK_ARC_1_0/buf_output[7] , \MC_ARK_ARC_1_0/buf_output[6] ,
         \MC_ARK_ARC_1_0/buf_output[5] , \MC_ARK_ARC_1_0/buf_output[4] ,
         \MC_ARK_ARC_1_0/buf_output[3] , \MC_ARK_ARC_1_0/buf_output[2] ,
         \MC_ARK_ARC_1_0/buf_output[1] , \MC_ARK_ARC_1_0/buf_output[0] ,
         \MC_ARK_ARC_1_0/temp6[185] , \MC_ARK_ARC_1_0/temp6[183] ,
         \MC_ARK_ARC_1_0/temp6[182] , \MC_ARK_ARC_1_0/temp6[181] ,
         \MC_ARK_ARC_1_0/temp6[178] , \MC_ARK_ARC_1_0/temp6[177] ,
         \MC_ARK_ARC_1_0/temp6[175] , \MC_ARK_ARC_1_0/temp6[173] ,
         \MC_ARK_ARC_1_0/temp6[172] , \MC_ARK_ARC_1_0/temp6[171] ,
         \MC_ARK_ARC_1_0/temp6[170] , \MC_ARK_ARC_1_0/temp6[169] ,
         \MC_ARK_ARC_1_0/temp6[163] , \MC_ARK_ARC_1_0/temp6[162] ,
         \MC_ARK_ARC_1_0/temp6[156] , \MC_ARK_ARC_1_0/temp6[155] ,
         \MC_ARK_ARC_1_0/temp6[154] , \MC_ARK_ARC_1_0/temp6[152] ,
         \MC_ARK_ARC_1_0/temp6[150] , \MC_ARK_ARC_1_0/temp6[148] ,
         \MC_ARK_ARC_1_0/temp6[147] , \MC_ARK_ARC_1_0/temp6[142] ,
         \MC_ARK_ARC_1_0/temp6[140] , \MC_ARK_ARC_1_0/temp6[139] ,
         \MC_ARK_ARC_1_0/temp6[130] , \MC_ARK_ARC_1_0/temp6[129] ,
         \MC_ARK_ARC_1_0/temp6[128] , \MC_ARK_ARC_1_0/temp6[125] ,
         \MC_ARK_ARC_1_0/temp6[118] , \MC_ARK_ARC_1_0/temp6[115] ,
         \MC_ARK_ARC_1_0/temp6[112] , \MC_ARK_ARC_1_0/temp6[108] ,
         \MC_ARK_ARC_1_0/temp6[106] , \MC_ARK_ARC_1_0/temp6[105] ,
         \MC_ARK_ARC_1_0/temp6[103] , \MC_ARK_ARC_1_0/temp6[99] ,
         \MC_ARK_ARC_1_0/temp6[97] , \MC_ARK_ARC_1_0/temp6[96] ,
         \MC_ARK_ARC_1_0/temp6[94] , \MC_ARK_ARC_1_0/temp6[91] ,
         \MC_ARK_ARC_1_0/temp6[90] , \MC_ARK_ARC_1_0/temp6[87] ,
         \MC_ARK_ARC_1_0/temp6[83] , \MC_ARK_ARC_1_0/temp6[82] ,
         \MC_ARK_ARC_1_0/temp6[81] , \MC_ARK_ARC_1_0/temp6[78] ,
         \MC_ARK_ARC_1_0/temp6[77] , \MC_ARK_ARC_1_0/temp6[75] ,
         \MC_ARK_ARC_1_0/temp6[74] , \MC_ARK_ARC_1_0/temp6[72] ,
         \MC_ARK_ARC_1_0/temp6[67] , \MC_ARK_ARC_1_0/temp6[65] ,
         \MC_ARK_ARC_1_0/temp6[64] , \MC_ARK_ARC_1_0/temp6[63] ,
         \MC_ARK_ARC_1_0/temp6[62] , \MC_ARK_ARC_1_0/temp6[61] ,
         \MC_ARK_ARC_1_0/temp6[56] , \MC_ARK_ARC_1_0/temp6[54] ,
         \MC_ARK_ARC_1_0/temp6[48] , \MC_ARK_ARC_1_0/temp6[45] ,
         \MC_ARK_ARC_1_0/temp6[43] , \MC_ARK_ARC_1_0/temp6[42] ,
         \MC_ARK_ARC_1_0/temp6[41] , \MC_ARK_ARC_1_0/temp6[40] ,
         \MC_ARK_ARC_1_0/temp6[38] , \MC_ARK_ARC_1_0/temp6[36] ,
         \MC_ARK_ARC_1_0/temp6[33] , \MC_ARK_ARC_1_0/temp6[31] ,
         \MC_ARK_ARC_1_0/temp6[30] , \MC_ARK_ARC_1_0/temp6[29] ,
         \MC_ARK_ARC_1_0/temp6[26] , \MC_ARK_ARC_1_0/temp6[25] ,
         \MC_ARK_ARC_1_0/temp6[19] , \MC_ARK_ARC_1_0/temp6[18] ,
         \MC_ARK_ARC_1_0/temp6[15] , \MC_ARK_ARC_1_0/temp6[14] ,
         \MC_ARK_ARC_1_0/temp6[13] , \MC_ARK_ARC_1_0/temp6[12] ,
         \MC_ARK_ARC_1_0/temp6[11] , \MC_ARK_ARC_1_0/temp6[10] ,
         \MC_ARK_ARC_1_0/temp6[9] , \MC_ARK_ARC_1_0/temp6[6] ,
         \MC_ARK_ARC_1_0/temp6[5] , \MC_ARK_ARC_1_0/temp6[4] ,
         \MC_ARK_ARC_1_0/temp6[3] , \MC_ARK_ARC_1_0/temp6[1] ,
         \MC_ARK_ARC_1_0/temp6[0] , \MC_ARK_ARC_1_0/temp5[190] ,
         \MC_ARK_ARC_1_0/temp5[187] , \MC_ARK_ARC_1_0/temp5[186] ,
         \MC_ARK_ARC_1_0/temp5[181] , \MC_ARK_ARC_1_0/temp5[179] ,
         \MC_ARK_ARC_1_0/temp5[178] , \MC_ARK_ARC_1_0/temp5[177] ,
         \MC_ARK_ARC_1_0/temp5[175] , \MC_ARK_ARC_1_0/temp5[173] ,
         \MC_ARK_ARC_1_0/temp5[171] , \MC_ARK_ARC_1_0/temp5[169] ,
         \MC_ARK_ARC_1_0/temp5[168] , \MC_ARK_ARC_1_0/temp5[167] ,
         \MC_ARK_ARC_1_0/temp5[166] , \MC_ARK_ARC_1_0/temp5[165] ,
         \MC_ARK_ARC_1_0/temp5[163] , \MC_ARK_ARC_1_0/temp5[162] ,
         \MC_ARK_ARC_1_0/temp5[160] , \MC_ARK_ARC_1_0/temp5[155] ,
         \MC_ARK_ARC_1_0/temp5[154] , \MC_ARK_ARC_1_0/temp5[153] ,
         \MC_ARK_ARC_1_0/temp5[152] , \MC_ARK_ARC_1_0/temp5[151] ,
         \MC_ARK_ARC_1_0/temp5[150] , \MC_ARK_ARC_1_0/temp5[147] ,
         \MC_ARK_ARC_1_0/temp5[146] , \MC_ARK_ARC_1_0/temp5[141] ,
         \MC_ARK_ARC_1_0/temp5[137] , \MC_ARK_ARC_1_0/temp5[136] ,
         \MC_ARK_ARC_1_0/temp5[135] , \MC_ARK_ARC_1_0/temp5[132] ,
         \MC_ARK_ARC_1_0/temp5[130] , \MC_ARK_ARC_1_0/temp5[129] ,
         \MC_ARK_ARC_1_0/temp5[128] , \MC_ARK_ARC_1_0/temp5[124] ,
         \MC_ARK_ARC_1_0/temp5[120] , \MC_ARK_ARC_1_0/temp5[118] ,
         \MC_ARK_ARC_1_0/temp5[116] , \MC_ARK_ARC_1_0/temp5[111] ,
         \MC_ARK_ARC_1_0/temp5[109] , \MC_ARK_ARC_1_0/temp5[108] ,
         \MC_ARK_ARC_1_0/temp5[107] , \MC_ARK_ARC_1_0/temp5[106] ,
         \MC_ARK_ARC_1_0/temp5[105] , \MC_ARK_ARC_1_0/temp5[103] ,
         \MC_ARK_ARC_1_0/temp5[102] , \MC_ARK_ARC_1_0/temp5[94] ,
         \MC_ARK_ARC_1_0/temp5[91] , \MC_ARK_ARC_1_0/temp5[90] ,
         \MC_ARK_ARC_1_0/temp5[89] , \MC_ARK_ARC_1_0/temp5[87] ,
         \MC_ARK_ARC_1_0/temp5[84] , \MC_ARK_ARC_1_0/temp5[83] ,
         \MC_ARK_ARC_1_0/temp5[79] , \MC_ARK_ARC_1_0/temp5[78] ,
         \MC_ARK_ARC_1_0/temp5[76] , \MC_ARK_ARC_1_0/temp5[72] ,
         \MC_ARK_ARC_1_0/temp5[70] , \MC_ARK_ARC_1_0/temp5[68] ,
         \MC_ARK_ARC_1_0/temp5[67] , \MC_ARK_ARC_1_0/temp5[64] ,
         \MC_ARK_ARC_1_0/temp5[62] , \MC_ARK_ARC_1_0/temp5[61] ,
         \MC_ARK_ARC_1_0/temp5[58] , \MC_ARK_ARC_1_0/temp5[56] ,
         \MC_ARK_ARC_1_0/temp5[54] , \MC_ARK_ARC_1_0/temp5[49] ,
         \MC_ARK_ARC_1_0/temp5[48] , \MC_ARK_ARC_1_0/temp5[47] ,
         \MC_ARK_ARC_1_0/temp5[46] , \MC_ARK_ARC_1_0/temp5[45] ,
         \MC_ARK_ARC_1_0/temp5[42] , \MC_ARK_ARC_1_0/temp5[38] ,
         \MC_ARK_ARC_1_0/temp5[37] , \MC_ARK_ARC_1_0/temp5[36] ,
         \MC_ARK_ARC_1_0/temp5[33] , \MC_ARK_ARC_1_0/temp5[32] ,
         \MC_ARK_ARC_1_0/temp5[31] , \MC_ARK_ARC_1_0/temp5[29] ,
         \MC_ARK_ARC_1_0/temp5[28] , \MC_ARK_ARC_1_0/temp5[27] ,
         \MC_ARK_ARC_1_0/temp5[25] , \MC_ARK_ARC_1_0/temp5[24] ,
         \MC_ARK_ARC_1_0/temp5[23] , \MC_ARK_ARC_1_0/temp5[21] ,
         \MC_ARK_ARC_1_0/temp5[19] , \MC_ARK_ARC_1_0/temp5[18] ,
         \MC_ARK_ARC_1_0/temp5[16] , \MC_ARK_ARC_1_0/temp5[15] ,
         \MC_ARK_ARC_1_0/temp5[14] , \MC_ARK_ARC_1_0/temp5[13] ,
         \MC_ARK_ARC_1_0/temp5[12] , \MC_ARK_ARC_1_0/temp5[10] ,
         \MC_ARK_ARC_1_0/temp5[9] , \MC_ARK_ARC_1_0/temp5[8] ,
         \MC_ARK_ARC_1_0/temp5[6] , \MC_ARK_ARC_1_0/temp5[4] ,
         \MC_ARK_ARC_1_0/temp5[2] , \MC_ARK_ARC_1_0/temp5[1] ,
         \MC_ARK_ARC_1_0/temp5[0] , \MC_ARK_ARC_1_0/temp4[191] ,
         \MC_ARK_ARC_1_0/temp4[190] , \MC_ARK_ARC_1_0/temp4[189] ,
         \MC_ARK_ARC_1_0/temp4[188] , \MC_ARK_ARC_1_0/temp4[187] ,
         \MC_ARK_ARC_1_0/temp4[186] , \MC_ARK_ARC_1_0/temp4[185] ,
         \MC_ARK_ARC_1_0/temp4[184] , \MC_ARK_ARC_1_0/temp4[183] ,
         \MC_ARK_ARC_1_0/temp4[182] , \MC_ARK_ARC_1_0/temp4[181] ,
         \MC_ARK_ARC_1_0/temp4[180] , \MC_ARK_ARC_1_0/temp4[179] ,
         \MC_ARK_ARC_1_0/temp4[178] , \MC_ARK_ARC_1_0/temp4[177] ,
         \MC_ARK_ARC_1_0/temp4[175] , \MC_ARK_ARC_1_0/temp4[174] ,
         \MC_ARK_ARC_1_0/temp4[173] , \MC_ARK_ARC_1_0/temp4[172] ,
         \MC_ARK_ARC_1_0/temp4[171] , \MC_ARK_ARC_1_0/temp4[170] ,
         \MC_ARK_ARC_1_0/temp4[169] , \MC_ARK_ARC_1_0/temp4[168] ,
         \MC_ARK_ARC_1_0/temp4[167] , \MC_ARK_ARC_1_0/temp4[166] ,
         \MC_ARK_ARC_1_0/temp4[164] , \MC_ARK_ARC_1_0/temp4[163] ,
         \MC_ARK_ARC_1_0/temp4[162] , \MC_ARK_ARC_1_0/temp4[161] ,
         \MC_ARK_ARC_1_0/temp4[160] , \MC_ARK_ARC_1_0/temp4[159] ,
         \MC_ARK_ARC_1_0/temp4[157] , \MC_ARK_ARC_1_0/temp4[156] ,
         \MC_ARK_ARC_1_0/temp4[155] , \MC_ARK_ARC_1_0/temp4[154] ,
         \MC_ARK_ARC_1_0/temp4[153] , \MC_ARK_ARC_1_0/temp4[152] ,
         \MC_ARK_ARC_1_0/temp4[151] , \MC_ARK_ARC_1_0/temp4[150] ,
         \MC_ARK_ARC_1_0/temp4[149] , \MC_ARK_ARC_1_0/temp4[148] ,
         \MC_ARK_ARC_1_0/temp4[147] , \MC_ARK_ARC_1_0/temp4[145] ,
         \MC_ARK_ARC_1_0/temp4[144] , \MC_ARK_ARC_1_0/temp4[142] ,
         \MC_ARK_ARC_1_0/temp4[141] , \MC_ARK_ARC_1_0/temp4[140] ,
         \MC_ARK_ARC_1_0/temp4[139] , \MC_ARK_ARC_1_0/temp4[138] ,
         \MC_ARK_ARC_1_0/temp4[137] , \MC_ARK_ARC_1_0/temp4[136] ,
         \MC_ARK_ARC_1_0/temp4[135] , \MC_ARK_ARC_1_0/temp4[134] ,
         \MC_ARK_ARC_1_0/temp4[133] , \MC_ARK_ARC_1_0/temp4[132] ,
         \MC_ARK_ARC_1_0/temp4[131] , \MC_ARK_ARC_1_0/temp4[130] ,
         \MC_ARK_ARC_1_0/temp4[129] , \MC_ARK_ARC_1_0/temp4[128] ,
         \MC_ARK_ARC_1_0/temp4[127] , \MC_ARK_ARC_1_0/temp4[125] ,
         \MC_ARK_ARC_1_0/temp4[124] , \MC_ARK_ARC_1_0/temp4[123] ,
         \MC_ARK_ARC_1_0/temp4[122] , \MC_ARK_ARC_1_0/temp4[121] ,
         \MC_ARK_ARC_1_0/temp4[120] , \MC_ARK_ARC_1_0/temp4[118] ,
         \MC_ARK_ARC_1_0/temp4[117] , \MC_ARK_ARC_1_0/temp4[116] ,
         \MC_ARK_ARC_1_0/temp4[115] , \MC_ARK_ARC_1_0/temp4[114] ,
         \MC_ARK_ARC_1_0/temp4[113] , \MC_ARK_ARC_1_0/temp4[112] ,
         \MC_ARK_ARC_1_0/temp4[111] , \MC_ARK_ARC_1_0/temp4[110] ,
         \MC_ARK_ARC_1_0/temp4[109] , \MC_ARK_ARC_1_0/temp4[108] ,
         \MC_ARK_ARC_1_0/temp4[107] , \MC_ARK_ARC_1_0/temp4[106] ,
         \MC_ARK_ARC_1_0/temp4[105] , \MC_ARK_ARC_1_0/temp4[104] ,
         \MC_ARK_ARC_1_0/temp4[103] , \MC_ARK_ARC_1_0/temp4[102] ,
         \MC_ARK_ARC_1_0/temp4[100] , \MC_ARK_ARC_1_0/temp4[99] ,
         \MC_ARK_ARC_1_0/temp4[98] , \MC_ARK_ARC_1_0/temp4[97] ,
         \MC_ARK_ARC_1_0/temp4[96] , \MC_ARK_ARC_1_0/temp4[95] ,
         \MC_ARK_ARC_1_0/temp4[94] , \MC_ARK_ARC_1_0/temp4[93] ,
         \MC_ARK_ARC_1_0/temp4[91] , \MC_ARK_ARC_1_0/temp4[90] ,
         \MC_ARK_ARC_1_0/temp4[89] , \MC_ARK_ARC_1_0/temp4[88] ,
         \MC_ARK_ARC_1_0/temp4[87] , \MC_ARK_ARC_1_0/temp4[86] ,
         \MC_ARK_ARC_1_0/temp4[85] , \MC_ARK_ARC_1_0/temp4[84] ,
         \MC_ARK_ARC_1_0/temp4[83] , \MC_ARK_ARC_1_0/temp4[82] ,
         \MC_ARK_ARC_1_0/temp4[81] , \MC_ARK_ARC_1_0/temp4[80] ,
         \MC_ARK_ARC_1_0/temp4[79] , \MC_ARK_ARC_1_0/temp4[78] ,
         \MC_ARK_ARC_1_0/temp4[77] , \MC_ARK_ARC_1_0/temp4[76] ,
         \MC_ARK_ARC_1_0/temp4[75] , \MC_ARK_ARC_1_0/temp4[74] ,
         \MC_ARK_ARC_1_0/temp4[73] , \MC_ARK_ARC_1_0/temp4[72] ,
         \MC_ARK_ARC_1_0/temp4[70] , \MC_ARK_ARC_1_0/temp4[68] ,
         \MC_ARK_ARC_1_0/temp4[67] , \MC_ARK_ARC_1_0/temp4[66] ,
         \MC_ARK_ARC_1_0/temp4[64] , \MC_ARK_ARC_1_0/temp4[63] ,
         \MC_ARK_ARC_1_0/temp4[61] , \MC_ARK_ARC_1_0/temp4[60] ,
         \MC_ARK_ARC_1_0/temp4[59] , \MC_ARK_ARC_1_0/temp4[58] ,
         \MC_ARK_ARC_1_0/temp4[57] , \MC_ARK_ARC_1_0/temp4[56] ,
         \MC_ARK_ARC_1_0/temp4[55] , \MC_ARK_ARC_1_0/temp4[54] ,
         \MC_ARK_ARC_1_0/temp4[53] , \MC_ARK_ARC_1_0/temp4[52] ,
         \MC_ARK_ARC_1_0/temp4[49] , \MC_ARK_ARC_1_0/temp4[48] ,
         \MC_ARK_ARC_1_0/temp4[47] , \MC_ARK_ARC_1_0/temp4[46] ,
         \MC_ARK_ARC_1_0/temp4[45] , \MC_ARK_ARC_1_0/temp4[44] ,
         \MC_ARK_ARC_1_0/temp4[43] , \MC_ARK_ARC_1_0/temp4[42] ,
         \MC_ARK_ARC_1_0/temp4[41] , \MC_ARK_ARC_1_0/temp4[40] ,
         \MC_ARK_ARC_1_0/temp4[39] , \MC_ARK_ARC_1_0/temp4[37] ,
         \MC_ARK_ARC_1_0/temp4[36] , \MC_ARK_ARC_1_0/temp4[35] ,
         \MC_ARK_ARC_1_0/temp4[34] , \MC_ARK_ARC_1_0/temp4[33] ,
         \MC_ARK_ARC_1_0/temp4[32] , \MC_ARK_ARC_1_0/temp4[31] ,
         \MC_ARK_ARC_1_0/temp4[30] , \MC_ARK_ARC_1_0/temp4[29] ,
         \MC_ARK_ARC_1_0/temp4[28] , \MC_ARK_ARC_1_0/temp4[27] ,
         \MC_ARK_ARC_1_0/temp4[26] , \MC_ARK_ARC_1_0/temp4[25] ,
         \MC_ARK_ARC_1_0/temp4[24] , \MC_ARK_ARC_1_0/temp4[23] ,
         \MC_ARK_ARC_1_0/temp4[22] , \MC_ARK_ARC_1_0/temp4[21] ,
         \MC_ARK_ARC_1_0/temp4[20] , \MC_ARK_ARC_1_0/temp4[19] ,
         \MC_ARK_ARC_1_0/temp4[18] , \MC_ARK_ARC_1_0/temp4[17] ,
         \MC_ARK_ARC_1_0/temp4[16] , \MC_ARK_ARC_1_0/temp4[14] ,
         \MC_ARK_ARC_1_0/temp4[13] , \MC_ARK_ARC_1_0/temp4[12] ,
         \MC_ARK_ARC_1_0/temp4[11] , \MC_ARK_ARC_1_0/temp4[10] ,
         \MC_ARK_ARC_1_0/temp4[9] , \MC_ARK_ARC_1_0/temp4[8] ,
         \MC_ARK_ARC_1_0/temp4[7] , \MC_ARK_ARC_1_0/temp4[6] ,
         \MC_ARK_ARC_1_0/temp4[5] , \MC_ARK_ARC_1_0/temp4[4] ,
         \MC_ARK_ARC_1_0/temp4[3] , \MC_ARK_ARC_1_0/temp4[2] ,
         \MC_ARK_ARC_1_0/temp4[1] , \MC_ARK_ARC_1_0/temp4[0] ,
         \MC_ARK_ARC_1_0/temp3[191] , \MC_ARK_ARC_1_0/temp3[190] ,
         \MC_ARK_ARC_1_0/temp3[187] , \MC_ARK_ARC_1_0/temp3[186] ,
         \MC_ARK_ARC_1_0/temp3[185] , \MC_ARK_ARC_1_0/temp3[184] ,
         \MC_ARK_ARC_1_0/temp3[183] , \MC_ARK_ARC_1_0/temp3[182] ,
         \MC_ARK_ARC_1_0/temp3[181] , \MC_ARK_ARC_1_0/temp3[179] ,
         \MC_ARK_ARC_1_0/temp3[178] , \MC_ARK_ARC_1_0/temp3[177] ,
         \MC_ARK_ARC_1_0/temp3[175] , \MC_ARK_ARC_1_0/temp3[174] ,
         \MC_ARK_ARC_1_0/temp3[173] , \MC_ARK_ARC_1_0/temp3[172] ,
         \MC_ARK_ARC_1_0/temp3[169] , \MC_ARK_ARC_1_0/temp3[168] ,
         \MC_ARK_ARC_1_0/temp3[167] , \MC_ARK_ARC_1_0/temp3[166] ,
         \MC_ARK_ARC_1_0/temp3[164] , \MC_ARK_ARC_1_0/temp3[162] ,
         \MC_ARK_ARC_1_0/temp3[161] , \MC_ARK_ARC_1_0/temp3[160] ,
         \MC_ARK_ARC_1_0/temp3[159] , \MC_ARK_ARC_1_0/temp3[157] ,
         \MC_ARK_ARC_1_0/temp3[156] , \MC_ARK_ARC_1_0/temp3[155] ,
         \MC_ARK_ARC_1_0/temp3[154] , \MC_ARK_ARC_1_0/temp3[152] ,
         \MC_ARK_ARC_1_0/temp3[151] , \MC_ARK_ARC_1_0/temp3[150] ,
         \MC_ARK_ARC_1_0/temp3[149] , \MC_ARK_ARC_1_0/temp3[147] ,
         \MC_ARK_ARC_1_0/temp3[145] , \MC_ARK_ARC_1_0/temp3[142] ,
         \MC_ARK_ARC_1_0/temp3[140] , \MC_ARK_ARC_1_0/temp3[139] ,
         \MC_ARK_ARC_1_0/temp3[136] , \MC_ARK_ARC_1_0/temp3[135] ,
         \MC_ARK_ARC_1_0/temp3[133] , \MC_ARK_ARC_1_0/temp3[132] ,
         \MC_ARK_ARC_1_0/temp3[131] , \MC_ARK_ARC_1_0/temp3[129] ,
         \MC_ARK_ARC_1_0/temp3[128] , \MC_ARK_ARC_1_0/temp3[127] ,
         \MC_ARK_ARC_1_0/temp3[124] , \MC_ARK_ARC_1_0/temp3[123] ,
         \MC_ARK_ARC_1_0/temp3[122] , \MC_ARK_ARC_1_0/temp3[120] ,
         \MC_ARK_ARC_1_0/temp3[118] , \MC_ARK_ARC_1_0/temp3[117] ,
         \MC_ARK_ARC_1_0/temp3[115] , \MC_ARK_ARC_1_0/temp3[114] ,
         \MC_ARK_ARC_1_0/temp3[112] , \MC_ARK_ARC_1_0/temp3[109] ,
         \MC_ARK_ARC_1_0/temp3[108] , \MC_ARK_ARC_1_0/temp3[107] ,
         \MC_ARK_ARC_1_0/temp3[106] , \MC_ARK_ARC_1_0/temp3[103] ,
         \MC_ARK_ARC_1_0/temp3[102] , \MC_ARK_ARC_1_0/temp3[100] ,
         \MC_ARK_ARC_1_0/temp3[99] , \MC_ARK_ARC_1_0/temp3[97] ,
         \MC_ARK_ARC_1_0/temp3[96] , \MC_ARK_ARC_1_0/temp3[95] ,
         \MC_ARK_ARC_1_0/temp3[94] , \MC_ARK_ARC_1_0/temp3[93] ,
         \MC_ARK_ARC_1_0/temp3[91] , \MC_ARK_ARC_1_0/temp3[90] ,
         \MC_ARK_ARC_1_0/temp3[89] , \MC_ARK_ARC_1_0/temp3[88] ,
         \MC_ARK_ARC_1_0/temp3[87] , \MC_ARK_ARC_1_0/temp3[85] ,
         \MC_ARK_ARC_1_0/temp3[84] , \MC_ARK_ARC_1_0/temp3[83] ,
         \MC_ARK_ARC_1_0/temp3[82] , \MC_ARK_ARC_1_0/temp3[81] ,
         \MC_ARK_ARC_1_0/temp3[80] , \MC_ARK_ARC_1_0/temp3[79] ,
         \MC_ARK_ARC_1_0/temp3[78] , \MC_ARK_ARC_1_0/temp3[77] ,
         \MC_ARK_ARC_1_0/temp3[76] , \MC_ARK_ARC_1_0/temp3[75] ,
         \MC_ARK_ARC_1_0/temp3[73] , \MC_ARK_ARC_1_0/temp3[72] ,
         \MC_ARK_ARC_1_0/temp3[70] , \MC_ARK_ARC_1_0/temp3[69] ,
         \MC_ARK_ARC_1_0/temp3[68] , \MC_ARK_ARC_1_0/temp3[67] ,
         \MC_ARK_ARC_1_0/temp3[66] , \MC_ARK_ARC_1_0/temp3[63] ,
         \MC_ARK_ARC_1_0/temp3[61] , \MC_ARK_ARC_1_0/temp3[60] ,
         \MC_ARK_ARC_1_0/temp3[59] , \MC_ARK_ARC_1_0/temp3[58] ,
         \MC_ARK_ARC_1_0/temp3[57] , \MC_ARK_ARC_1_0/temp3[54] ,
         \MC_ARK_ARC_1_0/temp3[52] , \MC_ARK_ARC_1_0/temp3[49] ,
         \MC_ARK_ARC_1_0/temp3[48] , \MC_ARK_ARC_1_0/temp3[47] ,
         \MC_ARK_ARC_1_0/temp3[46] , \MC_ARK_ARC_1_0/temp3[45] ,
         \MC_ARK_ARC_1_0/temp3[44] , \MC_ARK_ARC_1_0/temp3[43] ,
         \MC_ARK_ARC_1_0/temp3[42] , \MC_ARK_ARC_1_0/temp3[41] ,
         \MC_ARK_ARC_1_0/temp3[40] , \MC_ARK_ARC_1_0/temp3[39] ,
         \MC_ARK_ARC_1_0/temp3[37] , \MC_ARK_ARC_1_0/temp3[36] ,
         \MC_ARK_ARC_1_0/temp3[35] , \MC_ARK_ARC_1_0/temp3[33] ,
         \MC_ARK_ARC_1_0/temp3[32] , \MC_ARK_ARC_1_0/temp3[31] ,
         \MC_ARK_ARC_1_0/temp3[30] , \MC_ARK_ARC_1_0/temp3[29] ,
         \MC_ARK_ARC_1_0/temp3[28] , \MC_ARK_ARC_1_0/temp3[27] ,
         \MC_ARK_ARC_1_0/temp3[25] , \MC_ARK_ARC_1_0/temp3[24] ,
         \MC_ARK_ARC_1_0/temp3[23] , \MC_ARK_ARC_1_0/temp3[22] ,
         \MC_ARK_ARC_1_0/temp3[20] , \MC_ARK_ARC_1_0/temp3[19] ,
         \MC_ARK_ARC_1_0/temp3[17] , \MC_ARK_ARC_1_0/temp3[16] ,
         \MC_ARK_ARC_1_0/temp3[14] , \MC_ARK_ARC_1_0/temp3[13] ,
         \MC_ARK_ARC_1_0/temp3[12] , \MC_ARK_ARC_1_0/temp3[11] ,
         \MC_ARK_ARC_1_0/temp3[10] , \MC_ARK_ARC_1_0/temp3[9] ,
         \MC_ARK_ARC_1_0/temp3[7] , \MC_ARK_ARC_1_0/temp3[6] ,
         \MC_ARK_ARC_1_0/temp3[5] , \MC_ARK_ARC_1_0/temp3[4] ,
         \MC_ARK_ARC_1_0/temp3[3] , \MC_ARK_ARC_1_0/temp3[2] ,
         \MC_ARK_ARC_1_0/temp3[1] , \MC_ARK_ARC_1_0/temp3[0] ,
         \MC_ARK_ARC_1_0/temp2[191] , \MC_ARK_ARC_1_0/temp2[190] ,
         \MC_ARK_ARC_1_0/temp2[187] , \MC_ARK_ARC_1_0/temp2[185] ,
         \MC_ARK_ARC_1_0/temp2[181] , \MC_ARK_ARC_1_0/temp2[180] ,
         \MC_ARK_ARC_1_0/temp2[179] , \MC_ARK_ARC_1_0/temp2[178] ,
         \MC_ARK_ARC_1_0/temp2[177] , \MC_ARK_ARC_1_0/temp2[176] ,
         \MC_ARK_ARC_1_0/temp2[175] , \MC_ARK_ARC_1_0/temp2[174] ,
         \MC_ARK_ARC_1_0/temp2[173] , \MC_ARK_ARC_1_0/temp2[172] ,
         \MC_ARK_ARC_1_0/temp2[171] , \MC_ARK_ARC_1_0/temp2[170] ,
         \MC_ARK_ARC_1_0/temp2[169] , \MC_ARK_ARC_1_0/temp2[168] ,
         \MC_ARK_ARC_1_0/temp2[167] , \MC_ARK_ARC_1_0/temp2[166] ,
         \MC_ARK_ARC_1_0/temp2[165] , \MC_ARK_ARC_1_0/temp2[164] ,
         \MC_ARK_ARC_1_0/temp2[163] , \MC_ARK_ARC_1_0/temp2[162] ,
         \MC_ARK_ARC_1_0/temp2[161] , \MC_ARK_ARC_1_0/temp2[160] ,
         \MC_ARK_ARC_1_0/temp2[157] , \MC_ARK_ARC_1_0/temp2[156] ,
         \MC_ARK_ARC_1_0/temp2[154] , \MC_ARK_ARC_1_0/temp2[153] ,
         \MC_ARK_ARC_1_0/temp2[151] , \MC_ARK_ARC_1_0/temp2[150] ,
         \MC_ARK_ARC_1_0/temp2[148] , \MC_ARK_ARC_1_0/temp2[146] ,
         \MC_ARK_ARC_1_0/temp2[145] , \MC_ARK_ARC_1_0/temp2[144] ,
         \MC_ARK_ARC_1_0/temp2[142] , \MC_ARK_ARC_1_0/temp2[139] ,
         \MC_ARK_ARC_1_0/temp2[136] , \MC_ARK_ARC_1_0/temp2[135] ,
         \MC_ARK_ARC_1_0/temp2[134] , \MC_ARK_ARC_1_0/temp2[131] ,
         \MC_ARK_ARC_1_0/temp2[130] , \MC_ARK_ARC_1_0/temp2[129] ,
         \MC_ARK_ARC_1_0/temp2[127] , \MC_ARK_ARC_1_0/temp2[124] ,
         \MC_ARK_ARC_1_0/temp2[123] , \MC_ARK_ARC_1_0/temp2[120] ,
         \MC_ARK_ARC_1_0/temp2[118] , \MC_ARK_ARC_1_0/temp2[117] ,
         \MC_ARK_ARC_1_0/temp2[115] , \MC_ARK_ARC_1_0/temp2[114] ,
         \MC_ARK_ARC_1_0/temp2[113] , \MC_ARK_ARC_1_0/temp2[112] ,
         \MC_ARK_ARC_1_0/temp2[110] , \MC_ARK_ARC_1_0/temp2[109] ,
         \MC_ARK_ARC_1_0/temp2[108] , \MC_ARK_ARC_1_0/temp2[107] ,
         \MC_ARK_ARC_1_0/temp2[106] , \MC_ARK_ARC_1_0/temp2[105] ,
         \MC_ARK_ARC_1_0/temp2[104] , \MC_ARK_ARC_1_0/temp2[103] ,
         \MC_ARK_ARC_1_0/temp2[102] , \MC_ARK_ARC_1_0/temp2[101] ,
         \MC_ARK_ARC_1_0/temp2[100] , \MC_ARK_ARC_1_0/temp2[97] ,
         \MC_ARK_ARC_1_0/temp2[96] , \MC_ARK_ARC_1_0/temp2[92] ,
         \MC_ARK_ARC_1_0/temp2[91] , \MC_ARK_ARC_1_0/temp2[90] ,
         \MC_ARK_ARC_1_0/temp2[89] , \MC_ARK_ARC_1_0/temp2[87] ,
         \MC_ARK_ARC_1_0/temp2[86] , \MC_ARK_ARC_1_0/temp2[85] ,
         \MC_ARK_ARC_1_0/temp2[84] , \MC_ARK_ARC_1_0/temp2[81] ,
         \MC_ARK_ARC_1_0/temp2[80] , \MC_ARK_ARC_1_0/temp2[79] ,
         \MC_ARK_ARC_1_0/temp2[78] , \MC_ARK_ARC_1_0/temp2[77] ,
         \MC_ARK_ARC_1_0/temp2[76] , \MC_ARK_ARC_1_0/temp2[71] ,
         \MC_ARK_ARC_1_0/temp2[70] , \MC_ARK_ARC_1_0/temp2[68] ,
         \MC_ARK_ARC_1_0/temp2[67] , \MC_ARK_ARC_1_0/temp2[64] ,
         \MC_ARK_ARC_1_0/temp2[62] , \MC_ARK_ARC_1_0/temp2[61] ,
         \MC_ARK_ARC_1_0/temp2[60] , \MC_ARK_ARC_1_0/temp2[59] ,
         \MC_ARK_ARC_1_0/temp2[58] , \MC_ARK_ARC_1_0/temp2[55] ,
         \MC_ARK_ARC_1_0/temp2[49] , \MC_ARK_ARC_1_0/temp2[47] ,
         \MC_ARK_ARC_1_0/temp2[46] , \MC_ARK_ARC_1_0/temp2[45] ,
         \MC_ARK_ARC_1_0/temp2[44] , \MC_ARK_ARC_1_0/temp2[43] ,
         \MC_ARK_ARC_1_0/temp2[42] , \MC_ARK_ARC_1_0/temp2[41] ,
         \MC_ARK_ARC_1_0/temp2[40] , \MC_ARK_ARC_1_0/temp2[38] ,
         \MC_ARK_ARC_1_0/temp2[37] , \MC_ARK_ARC_1_0/temp2[36] ,
         \MC_ARK_ARC_1_0/temp2[34] , \MC_ARK_ARC_1_0/temp2[32] ,
         \MC_ARK_ARC_1_0/temp2[30] , \MC_ARK_ARC_1_0/temp2[29] ,
         \MC_ARK_ARC_1_0/temp2[27] , \MC_ARK_ARC_1_0/temp2[25] ,
         \MC_ARK_ARC_1_0/temp2[24] , \MC_ARK_ARC_1_0/temp2[23] ,
         \MC_ARK_ARC_1_0/temp2[22] , \MC_ARK_ARC_1_0/temp2[21] ,
         \MC_ARK_ARC_1_0/temp2[20] , \MC_ARK_ARC_1_0/temp2[19] ,
         \MC_ARK_ARC_1_0/temp2[18] , \MC_ARK_ARC_1_0/temp2[17] ,
         \MC_ARK_ARC_1_0/temp2[15] , \MC_ARK_ARC_1_0/temp2[14] ,
         \MC_ARK_ARC_1_0/temp2[13] , \MC_ARK_ARC_1_0/temp2[12] ,
         \MC_ARK_ARC_1_0/temp2[11] , \MC_ARK_ARC_1_0/temp2[10] ,
         \MC_ARK_ARC_1_0/temp2[9] , \MC_ARK_ARC_1_0/temp2[7] ,
         \MC_ARK_ARC_1_0/temp2[6] , \MC_ARK_ARC_1_0/temp2[4] ,
         \MC_ARK_ARC_1_0/temp2[1] , \MC_ARK_ARC_1_0/temp2[0] ,
         \MC_ARK_ARC_1_0/temp1[190] , \MC_ARK_ARC_1_0/temp1[189] ,
         \MC_ARK_ARC_1_0/temp1[187] , \MC_ARK_ARC_1_0/temp1[184] ,
         \MC_ARK_ARC_1_0/temp1[181] , \MC_ARK_ARC_1_0/temp1[180] ,
         \MC_ARK_ARC_1_0/temp1[179] , \MC_ARK_ARC_1_0/temp1[178] ,
         \MC_ARK_ARC_1_0/temp1[176] , \MC_ARK_ARC_1_0/temp1[175] ,
         \MC_ARK_ARC_1_0/temp1[174] , \MC_ARK_ARC_1_0/temp1[173] ,
         \MC_ARK_ARC_1_0/temp1[172] , \MC_ARK_ARC_1_0/temp1[169] ,
         \MC_ARK_ARC_1_0/temp1[168] , \MC_ARK_ARC_1_0/temp1[166] ,
         \MC_ARK_ARC_1_0/temp1[165] , \MC_ARK_ARC_1_0/temp1[162] ,
         \MC_ARK_ARC_1_0/temp1[161] , \MC_ARK_ARC_1_0/temp1[158] ,
         \MC_ARK_ARC_1_0/temp1[156] , \MC_ARK_ARC_1_0/temp1[151] ,
         \MC_ARK_ARC_1_0/temp1[150] , \MC_ARK_ARC_1_0/temp1[148] ,
         \MC_ARK_ARC_1_0/temp1[146] , \MC_ARK_ARC_1_0/temp1[145] ,
         \MC_ARK_ARC_1_0/temp1[144] , \MC_ARK_ARC_1_0/temp1[142] ,
         \MC_ARK_ARC_1_0/temp1[141] , \MC_ARK_ARC_1_0/temp1[139] ,
         \MC_ARK_ARC_1_0/temp1[137] , \MC_ARK_ARC_1_0/temp1[136] ,
         \MC_ARK_ARC_1_0/temp1[135] , \MC_ARK_ARC_1_0/temp1[132] ,
         \MC_ARK_ARC_1_0/temp1[131] , \MC_ARK_ARC_1_0/temp1[130] ,
         \MC_ARK_ARC_1_0/temp1[128] , \MC_ARK_ARC_1_0/temp1[127] ,
         \MC_ARK_ARC_1_0/temp1[125] , \MC_ARK_ARC_1_0/temp1[123] ,
         \MC_ARK_ARC_1_0/temp1[122] , \MC_ARK_ARC_1_0/temp1[121] ,
         \MC_ARK_ARC_1_0/temp1[120] , \MC_ARK_ARC_1_0/temp1[118] ,
         \MC_ARK_ARC_1_0/temp1[116] , \MC_ARK_ARC_1_0/temp1[115] ,
         \MC_ARK_ARC_1_0/temp1[114] , \MC_ARK_ARC_1_0/temp1[112] ,
         \MC_ARK_ARC_1_0/temp1[110] , \MC_ARK_ARC_1_0/temp1[109] ,
         \MC_ARK_ARC_1_0/temp1[108] , \MC_ARK_ARC_1_0/temp1[107] ,
         \MC_ARK_ARC_1_0/temp1[106] , \MC_ARK_ARC_1_0/temp1[105] ,
         \MC_ARK_ARC_1_0/temp1[102] , \MC_ARK_ARC_1_0/temp1[99] ,
         \MC_ARK_ARC_1_0/temp1[97] , \MC_ARK_ARC_1_0/temp1[96] ,
         \MC_ARK_ARC_1_0/temp1[94] , \MC_ARK_ARC_1_0/temp1[90] ,
         \MC_ARK_ARC_1_0/temp1[89] , \MC_ARK_ARC_1_0/temp1[88] ,
         \MC_ARK_ARC_1_0/temp1[85] , \MC_ARK_ARC_1_0/temp1[84] ,
         \MC_ARK_ARC_1_0/temp1[83] , \MC_ARK_ARC_1_0/temp1[82] ,
         \MC_ARK_ARC_1_0/temp1[79] , \MC_ARK_ARC_1_0/temp1[78] ,
         \MC_ARK_ARC_1_0/temp1[77] , \MC_ARK_ARC_1_0/temp1[76] ,
         \MC_ARK_ARC_1_0/temp1[75] , \MC_ARK_ARC_1_0/temp1[72] ,
         \MC_ARK_ARC_1_0/temp1[70] , \MC_ARK_ARC_1_0/temp1[69] ,
         \MC_ARK_ARC_1_0/temp1[66] , \MC_ARK_ARC_1_0/temp1[64] ,
         \MC_ARK_ARC_1_0/temp1[63] , \MC_ARK_ARC_1_0/temp1[62] ,
         \MC_ARK_ARC_1_0/temp1[61] , \MC_ARK_ARC_1_0/temp1[60] ,
         \MC_ARK_ARC_1_0/temp1[58] , \MC_ARK_ARC_1_0/temp1[57] ,
         \MC_ARK_ARC_1_0/temp1[55] , \MC_ARK_ARC_1_0/temp1[54] ,
         \MC_ARK_ARC_1_0/temp1[52] , \MC_ARK_ARC_1_0/temp1[49] ,
         \MC_ARK_ARC_1_0/temp1[48] , \MC_ARK_ARC_1_0/temp1[47] ,
         \MC_ARK_ARC_1_0/temp1[46] , \MC_ARK_ARC_1_0/temp1[45] ,
         \MC_ARK_ARC_1_0/temp1[42] , \MC_ARK_ARC_1_0/temp1[41] ,
         \MC_ARK_ARC_1_0/temp1[40] , \MC_ARK_ARC_1_0/temp1[38] ,
         \MC_ARK_ARC_1_0/temp1[37] , \MC_ARK_ARC_1_0/temp1[36] ,
         \MC_ARK_ARC_1_0/temp1[34] , \MC_ARK_ARC_1_0/temp1[32] ,
         \MC_ARK_ARC_1_0/temp1[31] , \MC_ARK_ARC_1_0/temp1[30] ,
         \MC_ARK_ARC_1_0/temp1[28] , \MC_ARK_ARC_1_0/temp1[26] ,
         \MC_ARK_ARC_1_0/temp1[25] , \MC_ARK_ARC_1_0/temp1[22] ,
         \MC_ARK_ARC_1_0/temp1[20] , \MC_ARK_ARC_1_0/temp1[18] ,
         \MC_ARK_ARC_1_0/temp1[17] , \MC_ARK_ARC_1_0/temp1[16] ,
         \MC_ARK_ARC_1_0/temp1[14] , \MC_ARK_ARC_1_0/temp1[13] ,
         \MC_ARK_ARC_1_0/temp1[12] , \MC_ARK_ARC_1_0/temp1[10] ,
         \MC_ARK_ARC_1_0/temp1[7] , \MC_ARK_ARC_1_0/temp1[6] ,
         \MC_ARK_ARC_1_0/temp1[5] , \MC_ARK_ARC_1_0/temp1[2] ,
         \MC_ARK_ARC_1_0/temp1[1] , \MC_ARK_ARC_1_0/temp1[0] ,
         \MC_ARK_ARC_1_0/buf_datainput[180] ,
         \MC_ARK_ARC_1_0/buf_datainput[179] ,
         \MC_ARK_ARC_1_0/buf_datainput[167] ,
         \MC_ARK_ARC_1_0/buf_datainput[166] ,
         \MC_ARK_ARC_1_0/buf_datainput[165] ,
         \MC_ARK_ARC_1_0/buf_datainput[157] ,
         \MC_ARK_ARC_1_0/buf_datainput[156] ,
         \MC_ARK_ARC_1_0/buf_datainput[155] ,
         \MC_ARK_ARC_1_0/buf_datainput[150] ,
         \MC_ARK_ARC_1_0/buf_datainput[144] ,
         \MC_ARK_ARC_1_0/buf_datainput[141] ,
         \MC_ARK_ARC_1_0/buf_datainput[138] ,
         \MC_ARK_ARC_1_0/buf_datainput[132] ,
         \MC_ARK_ARC_1_0/buf_datainput[115] ,
         \MC_ARK_ARC_1_0/buf_datainput[112] ,
         \MC_ARK_ARC_1_0/buf_datainput[109] ,
         \MC_ARK_ARC_1_0/buf_datainput[105] ,
         \MC_ARK_ARC_1_0/buf_datainput[96] ,
         \MC_ARK_ARC_1_0/buf_datainput[92] ,
         \MC_ARK_ARC_1_0/buf_datainput[90] ,
         \MC_ARK_ARC_1_0/buf_datainput[88] ,
         \MC_ARK_ARC_1_0/buf_datainput[86] ,
         \MC_ARK_ARC_1_0/buf_datainput[82] ,
         \MC_ARK_ARC_1_0/buf_datainput[81] ,
         \MC_ARK_ARC_1_0/buf_datainput[79] ,
         \MC_ARK_ARC_1_0/buf_datainput[78] ,
         \MC_ARK_ARC_1_0/buf_datainput[76] ,
         \MC_ARK_ARC_1_0/buf_datainput[73] ,
         \MC_ARK_ARC_1_0/buf_datainput[69] ,
         \MC_ARK_ARC_1_0/buf_datainput[67] ,
         \MC_ARK_ARC_1_0/buf_datainput[61] ,
         \MC_ARK_ARC_1_0/buf_datainput[56] ,
         \MC_ARK_ARC_1_0/buf_datainput[51] ,
         \MC_ARK_ARC_1_0/buf_datainput[49] ,
         \MC_ARK_ARC_1_0/buf_datainput[48] ,
         \MC_ARK_ARC_1_0/buf_datainput[46] ,
         \MC_ARK_ARC_1_0/buf_datainput[44] ,
         \MC_ARK_ARC_1_0/buf_datainput[42] ,
         \MC_ARK_ARC_1_0/buf_datainput[36] ,
         \MC_ARK_ARC_1_0/buf_datainput[22] ,
         \MC_ARK_ARC_1_0/buf_datainput[21] ,
         \MC_ARK_ARC_1_0/buf_datainput[12] , \MC_ARK_ARC_1_0/buf_datainput[7] ,
         \MC_ARK_ARC_1_0/buf_datainput[2] , \MC_ARK_ARC_1_1/buf_output[191] ,
         \MC_ARK_ARC_1_1/buf_output[190] , \MC_ARK_ARC_1_1/buf_output[189] ,
         \MC_ARK_ARC_1_1/buf_output[188] , \MC_ARK_ARC_1_1/buf_output[187] ,
         \MC_ARK_ARC_1_1/buf_output[186] , \MC_ARK_ARC_1_1/buf_output[185] ,
         \MC_ARK_ARC_1_1/buf_output[184] , \MC_ARK_ARC_1_1/buf_output[183] ,
         \MC_ARK_ARC_1_1/buf_output[182] , \MC_ARK_ARC_1_1/buf_output[181] ,
         \MC_ARK_ARC_1_1/buf_output[180] , \MC_ARK_ARC_1_1/buf_output[179] ,
         \MC_ARK_ARC_1_1/buf_output[178] , \MC_ARK_ARC_1_1/buf_output[177] ,
         \MC_ARK_ARC_1_1/buf_output[176] , \MC_ARK_ARC_1_1/buf_output[175] ,
         \MC_ARK_ARC_1_1/buf_output[174] , \MC_ARK_ARC_1_1/buf_output[173] ,
         \MC_ARK_ARC_1_1/buf_output[172] , \MC_ARK_ARC_1_1/buf_output[171] ,
         \MC_ARK_ARC_1_1/buf_output[170] , \MC_ARK_ARC_1_1/buf_output[169] ,
         \MC_ARK_ARC_1_1/buf_output[168] , \MC_ARK_ARC_1_1/buf_output[166] ,
         \MC_ARK_ARC_1_1/buf_output[165] , \MC_ARK_ARC_1_1/buf_output[164] ,
         \MC_ARK_ARC_1_1/buf_output[163] , \MC_ARK_ARC_1_1/buf_output[162] ,
         \MC_ARK_ARC_1_1/buf_output[161] , \MC_ARK_ARC_1_1/buf_output[160] ,
         \MC_ARK_ARC_1_1/buf_output[159] , \MC_ARK_ARC_1_1/buf_output[158] ,
         \MC_ARK_ARC_1_1/buf_output[157] , \MC_ARK_ARC_1_1/buf_output[156] ,
         \MC_ARK_ARC_1_1/buf_output[155] , \MC_ARK_ARC_1_1/buf_output[154] ,
         \MC_ARK_ARC_1_1/buf_output[153] , \MC_ARK_ARC_1_1/buf_output[152] ,
         \MC_ARK_ARC_1_1/buf_output[151] , \MC_ARK_ARC_1_1/buf_output[150] ,
         \MC_ARK_ARC_1_1/buf_output[149] , \MC_ARK_ARC_1_1/buf_output[148] ,
         \MC_ARK_ARC_1_1/buf_output[147] , \MC_ARK_ARC_1_1/buf_output[146] ,
         \MC_ARK_ARC_1_1/buf_output[145] , \MC_ARK_ARC_1_1/buf_output[144] ,
         \MC_ARK_ARC_1_1/buf_output[143] , \MC_ARK_ARC_1_1/buf_output[141] ,
         \MC_ARK_ARC_1_1/buf_output[140] , \MC_ARK_ARC_1_1/buf_output[139] ,
         \MC_ARK_ARC_1_1/buf_output[138] , \MC_ARK_ARC_1_1/buf_output[137] ,
         \MC_ARK_ARC_1_1/buf_output[136] , \MC_ARK_ARC_1_1/buf_output[135] ,
         \MC_ARK_ARC_1_1/buf_output[134] , \MC_ARK_ARC_1_1/buf_output[133] ,
         \MC_ARK_ARC_1_1/buf_output[132] , \MC_ARK_ARC_1_1/buf_output[131] ,
         \MC_ARK_ARC_1_1/buf_output[130] , \MC_ARK_ARC_1_1/buf_output[129] ,
         \MC_ARK_ARC_1_1/buf_output[128] , \MC_ARK_ARC_1_1/buf_output[127] ,
         \MC_ARK_ARC_1_1/buf_output[126] , \MC_ARK_ARC_1_1/buf_output[125] ,
         \MC_ARK_ARC_1_1/buf_output[124] , \MC_ARK_ARC_1_1/buf_output[123] ,
         \MC_ARK_ARC_1_1/buf_output[122] , \MC_ARK_ARC_1_1/buf_output[121] ,
         \MC_ARK_ARC_1_1/buf_output[120] , \MC_ARK_ARC_1_1/buf_output[119] ,
         \MC_ARK_ARC_1_1/buf_output[118] , \MC_ARK_ARC_1_1/buf_output[117] ,
         \MC_ARK_ARC_1_1/buf_output[116] , \MC_ARK_ARC_1_1/buf_output[115] ,
         \MC_ARK_ARC_1_1/buf_output[114] , \MC_ARK_ARC_1_1/buf_output[113] ,
         \MC_ARK_ARC_1_1/buf_output[112] , \MC_ARK_ARC_1_1/buf_output[111] ,
         \MC_ARK_ARC_1_1/buf_output[110] , \MC_ARK_ARC_1_1/buf_output[109] ,
         \MC_ARK_ARC_1_1/buf_output[108] , \MC_ARK_ARC_1_1/buf_output[107] ,
         \MC_ARK_ARC_1_1/buf_output[106] , \MC_ARK_ARC_1_1/buf_output[105] ,
         \MC_ARK_ARC_1_1/buf_output[104] , \MC_ARK_ARC_1_1/buf_output[103] ,
         \MC_ARK_ARC_1_1/buf_output[102] , \MC_ARK_ARC_1_1/buf_output[101] ,
         \MC_ARK_ARC_1_1/buf_output[100] , \MC_ARK_ARC_1_1/buf_output[99] ,
         \MC_ARK_ARC_1_1/buf_output[98] , \MC_ARK_ARC_1_1/buf_output[97] ,
         \MC_ARK_ARC_1_1/buf_output[96] , \MC_ARK_ARC_1_1/buf_output[95] ,
         \MC_ARK_ARC_1_1/buf_output[94] , \MC_ARK_ARC_1_1/buf_output[93] ,
         \MC_ARK_ARC_1_1/buf_output[92] , \MC_ARK_ARC_1_1/buf_output[91] ,
         \MC_ARK_ARC_1_1/buf_output[90] , \MC_ARK_ARC_1_1/buf_output[89] ,
         \MC_ARK_ARC_1_1/buf_output[88] , \MC_ARK_ARC_1_1/buf_output[87] ,
         \MC_ARK_ARC_1_1/buf_output[86] , \MC_ARK_ARC_1_1/buf_output[85] ,
         \MC_ARK_ARC_1_1/buf_output[84] , \MC_ARK_ARC_1_1/buf_output[83] ,
         \MC_ARK_ARC_1_1/buf_output[82] , \MC_ARK_ARC_1_1/buf_output[81] ,
         \MC_ARK_ARC_1_1/buf_output[80] , \MC_ARK_ARC_1_1/buf_output[79] ,
         \MC_ARK_ARC_1_1/buf_output[78] , \MC_ARK_ARC_1_1/buf_output[77] ,
         \MC_ARK_ARC_1_1/buf_output[76] , \MC_ARK_ARC_1_1/buf_output[75] ,
         \MC_ARK_ARC_1_1/buf_output[74] , \MC_ARK_ARC_1_1/buf_output[73] ,
         \MC_ARK_ARC_1_1/buf_output[72] , \MC_ARK_ARC_1_1/buf_output[71] ,
         \MC_ARK_ARC_1_1/buf_output[70] , \MC_ARK_ARC_1_1/buf_output[69] ,
         \MC_ARK_ARC_1_1/buf_output[68] , \MC_ARK_ARC_1_1/buf_output[67] ,
         \MC_ARK_ARC_1_1/buf_output[66] , \MC_ARK_ARC_1_1/buf_output[64] ,
         \MC_ARK_ARC_1_1/buf_output[63] , \MC_ARK_ARC_1_1/buf_output[62] ,
         \MC_ARK_ARC_1_1/buf_output[61] , \MC_ARK_ARC_1_1/buf_output[60] ,
         \MC_ARK_ARC_1_1/buf_output[58] , \MC_ARK_ARC_1_1/buf_output[57] ,
         \MC_ARK_ARC_1_1/buf_output[56] , \MC_ARK_ARC_1_1/buf_output[55] ,
         \MC_ARK_ARC_1_1/buf_output[54] , \MC_ARK_ARC_1_1/buf_output[53] ,
         \MC_ARK_ARC_1_1/buf_output[52] , \MC_ARK_ARC_1_1/buf_output[51] ,
         \MC_ARK_ARC_1_1/buf_output[50] , \MC_ARK_ARC_1_1/buf_output[49] ,
         \MC_ARK_ARC_1_1/buf_output[48] , \MC_ARK_ARC_1_1/buf_output[47] ,
         \MC_ARK_ARC_1_1/buf_output[46] , \MC_ARK_ARC_1_1/buf_output[45] ,
         \MC_ARK_ARC_1_1/buf_output[44] , \MC_ARK_ARC_1_1/buf_output[43] ,
         \MC_ARK_ARC_1_1/buf_output[42] , \MC_ARK_ARC_1_1/buf_output[41] ,
         \MC_ARK_ARC_1_1/buf_output[40] , \MC_ARK_ARC_1_1/buf_output[39] ,
         \MC_ARK_ARC_1_1/buf_output[38] , \MC_ARK_ARC_1_1/buf_output[37] ,
         \MC_ARK_ARC_1_1/buf_output[36] , \MC_ARK_ARC_1_1/buf_output[35] ,
         \MC_ARK_ARC_1_1/buf_output[34] , \MC_ARK_ARC_1_1/buf_output[33] ,
         \MC_ARK_ARC_1_1/buf_output[32] , \MC_ARK_ARC_1_1/buf_output[31] ,
         \MC_ARK_ARC_1_1/buf_output[30] , \MC_ARK_ARC_1_1/buf_output[29] ,
         \MC_ARK_ARC_1_1/buf_output[28] , \MC_ARK_ARC_1_1/buf_output[27] ,
         \MC_ARK_ARC_1_1/buf_output[26] , \MC_ARK_ARC_1_1/buf_output[25] ,
         \MC_ARK_ARC_1_1/buf_output[24] , \MC_ARK_ARC_1_1/buf_output[23] ,
         \MC_ARK_ARC_1_1/buf_output[22] , \MC_ARK_ARC_1_1/buf_output[21] ,
         \MC_ARK_ARC_1_1/buf_output[20] , \MC_ARK_ARC_1_1/buf_output[19] ,
         \MC_ARK_ARC_1_1/buf_output[18] , \MC_ARK_ARC_1_1/buf_output[17] ,
         \MC_ARK_ARC_1_1/buf_output[16] , \MC_ARK_ARC_1_1/buf_output[15] ,
         \MC_ARK_ARC_1_1/buf_output[14] , \MC_ARK_ARC_1_1/buf_output[13] ,
         \MC_ARK_ARC_1_1/buf_output[12] , \MC_ARK_ARC_1_1/buf_output[11] ,
         \MC_ARK_ARC_1_1/buf_output[10] , \MC_ARK_ARC_1_1/buf_output[9] ,
         \MC_ARK_ARC_1_1/buf_output[8] , \MC_ARK_ARC_1_1/buf_output[7] ,
         \MC_ARK_ARC_1_1/buf_output[6] , \MC_ARK_ARC_1_1/buf_output[5] ,
         \MC_ARK_ARC_1_1/buf_output[4] , \MC_ARK_ARC_1_1/buf_output[3] ,
         \MC_ARK_ARC_1_1/buf_output[2] , \MC_ARK_ARC_1_1/buf_output[1] ,
         \MC_ARK_ARC_1_1/buf_output[0] , \MC_ARK_ARC_1_1/temp6[189] ,
         \MC_ARK_ARC_1_1/temp6[185] , \MC_ARK_ARC_1_1/temp6[183] ,
         \MC_ARK_ARC_1_1/temp6[180] , \MC_ARK_ARC_1_1/temp6[178] ,
         \MC_ARK_ARC_1_1/temp6[176] , \MC_ARK_ARC_1_1/temp6[172] ,
         \MC_ARK_ARC_1_1/temp6[166] , \MC_ARK_ARC_1_1/temp6[162] ,
         \MC_ARK_ARC_1_1/temp6[160] , \MC_ARK_ARC_1_1/temp6[158] ,
         \MC_ARK_ARC_1_1/temp6[156] , \MC_ARK_ARC_1_1/temp6[155] ,
         \MC_ARK_ARC_1_1/temp6[152] , \MC_ARK_ARC_1_1/temp6[150] ,
         \MC_ARK_ARC_1_1/temp6[148] , \MC_ARK_ARC_1_1/temp6[146] ,
         \MC_ARK_ARC_1_1/temp6[144] , \MC_ARK_ARC_1_1/temp6[143] ,
         \MC_ARK_ARC_1_1/temp6[142] , \MC_ARK_ARC_1_1/temp6[140] ,
         \MC_ARK_ARC_1_1/temp6[138] , \MC_ARK_ARC_1_1/temp6[137] ,
         \MC_ARK_ARC_1_1/temp6[134] , \MC_ARK_ARC_1_1/temp6[127] ,
         \MC_ARK_ARC_1_1/temp6[124] , \MC_ARK_ARC_1_1/temp6[118] ,
         \MC_ARK_ARC_1_1/temp6[116] , \MC_ARK_ARC_1_1/temp6[109] ,
         \MC_ARK_ARC_1_1/temp6[108] , \MC_ARK_ARC_1_1/temp6[107] ,
         \MC_ARK_ARC_1_1/temp6[106] , \MC_ARK_ARC_1_1/temp6[105] ,
         \MC_ARK_ARC_1_1/temp6[104] , \MC_ARK_ARC_1_1/temp6[103] ,
         \MC_ARK_ARC_1_1/temp6[102] , \MC_ARK_ARC_1_1/temp6[101] ,
         \MC_ARK_ARC_1_1/temp6[95] , \MC_ARK_ARC_1_1/temp6[94] ,
         \MC_ARK_ARC_1_1/temp6[92] , \MC_ARK_ARC_1_1/temp6[85] ,
         \MC_ARK_ARC_1_1/temp6[82] , \MC_ARK_ARC_1_1/temp6[81] ,
         \MC_ARK_ARC_1_1/temp6[80] , \MC_ARK_ARC_1_1/temp6[78] ,
         \MC_ARK_ARC_1_1/temp6[76] , \MC_ARK_ARC_1_1/temp6[75] ,
         \MC_ARK_ARC_1_1/temp6[73] , \MC_ARK_ARC_1_1/temp6[72] ,
         \MC_ARK_ARC_1_1/temp6[69] , \MC_ARK_ARC_1_1/temp6[65] ,
         \MC_ARK_ARC_1_1/temp6[64] , \MC_ARK_ARC_1_1/temp6[61] ,
         \MC_ARK_ARC_1_1/temp6[59] , \MC_ARK_ARC_1_1/temp6[58] ,
         \MC_ARK_ARC_1_1/temp6[57] , \MC_ARK_ARC_1_1/temp6[56] ,
         \MC_ARK_ARC_1_1/temp6[55] , \MC_ARK_ARC_1_1/temp6[54] ,
         \MC_ARK_ARC_1_1/temp6[51] , \MC_ARK_ARC_1_1/temp6[48] ,
         \MC_ARK_ARC_1_1/temp6[47] , \MC_ARK_ARC_1_1/temp6[45] ,
         \MC_ARK_ARC_1_1/temp6[42] , \MC_ARK_ARC_1_1/temp6[41] ,
         \MC_ARK_ARC_1_1/temp6[39] , \MC_ARK_ARC_1_1/temp6[38] ,
         \MC_ARK_ARC_1_1/temp6[37] , \MC_ARK_ARC_1_1/temp6[36] ,
         \MC_ARK_ARC_1_1/temp6[31] , \MC_ARK_ARC_1_1/temp6[29] ,
         \MC_ARK_ARC_1_1/temp6[28] , \MC_ARK_ARC_1_1/temp6[27] ,
         \MC_ARK_ARC_1_1/temp6[25] , \MC_ARK_ARC_1_1/temp6[24] ,
         \MC_ARK_ARC_1_1/temp6[22] , \MC_ARK_ARC_1_1/temp6[21] ,
         \MC_ARK_ARC_1_1/temp6[19] , \MC_ARK_ARC_1_1/temp6[14] ,
         \MC_ARK_ARC_1_1/temp6[11] , \MC_ARK_ARC_1_1/temp6[6] ,
         \MC_ARK_ARC_1_1/temp6[5] , \MC_ARK_ARC_1_1/temp6[4] ,
         \MC_ARK_ARC_1_1/temp6[1] , \MC_ARK_ARC_1_1/temp6[0] ,
         \MC_ARK_ARC_1_1/temp5[185] , \MC_ARK_ARC_1_1/temp5[184] ,
         \MC_ARK_ARC_1_1/temp5[183] , \MC_ARK_ARC_1_1/temp5[177] ,
         \MC_ARK_ARC_1_1/temp5[175] , \MC_ARK_ARC_1_1/temp5[174] ,
         \MC_ARK_ARC_1_1/temp5[173] , \MC_ARK_ARC_1_1/temp5[172] ,
         \MC_ARK_ARC_1_1/temp5[171] , \MC_ARK_ARC_1_1/temp5[169] ,
         \MC_ARK_ARC_1_1/temp5[168] , \MC_ARK_ARC_1_1/temp5[164] ,
         \MC_ARK_ARC_1_1/temp5[160] , \MC_ARK_ARC_1_1/temp5[159] ,
         \MC_ARK_ARC_1_1/temp5[158] , \MC_ARK_ARC_1_1/temp5[156] ,
         \MC_ARK_ARC_1_1/temp5[154] , \MC_ARK_ARC_1_1/temp5[153] ,
         \MC_ARK_ARC_1_1/temp5[152] , \MC_ARK_ARC_1_1/temp5[151] ,
         \MC_ARK_ARC_1_1/temp5[150] , \MC_ARK_ARC_1_1/temp5[146] ,
         \MC_ARK_ARC_1_1/temp5[145] , \MC_ARK_ARC_1_1/temp5[144] ,
         \MC_ARK_ARC_1_1/temp5[143] , \MC_ARK_ARC_1_1/temp5[142] ,
         \MC_ARK_ARC_1_1/temp5[141] , \MC_ARK_ARC_1_1/temp5[140] ,
         \MC_ARK_ARC_1_1/temp5[138] , \MC_ARK_ARC_1_1/temp5[137] ,
         \MC_ARK_ARC_1_1/temp5[135] , \MC_ARK_ARC_1_1/temp5[133] ,
         \MC_ARK_ARC_1_1/temp5[129] , \MC_ARK_ARC_1_1/temp5[128] ,
         \MC_ARK_ARC_1_1/temp5[127] , \MC_ARK_ARC_1_1/temp5[124] ,
         \MC_ARK_ARC_1_1/temp5[123] , \MC_ARK_ARC_1_1/temp5[121] ,
         \MC_ARK_ARC_1_1/temp5[120] , \MC_ARK_ARC_1_1/temp5[119] ,
         \MC_ARK_ARC_1_1/temp5[118] , \MC_ARK_ARC_1_1/temp5[110] ,
         \MC_ARK_ARC_1_1/temp5[107] , \MC_ARK_ARC_1_1/temp5[105] ,
         \MC_ARK_ARC_1_1/temp5[104] , \MC_ARK_ARC_1_1/temp5[102] ,
         \MC_ARK_ARC_1_1/temp5[101] , \MC_ARK_ARC_1_1/temp5[99] ,
         \MC_ARK_ARC_1_1/temp5[98] , \MC_ARK_ARC_1_1/temp5[97] ,
         \MC_ARK_ARC_1_1/temp5[94] , \MC_ARK_ARC_1_1/temp5[90] ,
         \MC_ARK_ARC_1_1/temp5[87] , \MC_ARK_ARC_1_1/temp5[86] ,
         \MC_ARK_ARC_1_1/temp5[83] , \MC_ARK_ARC_1_1/temp5[82] ,
         \MC_ARK_ARC_1_1/temp5[78] , \MC_ARK_ARC_1_1/temp5[72] ,
         \MC_ARK_ARC_1_1/temp5[71] , \MC_ARK_ARC_1_1/temp5[69] ,
         \MC_ARK_ARC_1_1/temp5[68] , \MC_ARK_ARC_1_1/temp5[66] ,
         \MC_ARK_ARC_1_1/temp5[64] , \MC_ARK_ARC_1_1/temp5[61] ,
         \MC_ARK_ARC_1_1/temp5[57] , \MC_ARK_ARC_1_1/temp5[55] ,
         \MC_ARK_ARC_1_1/temp5[54] , \MC_ARK_ARC_1_1/temp5[52] ,
         \MC_ARK_ARC_1_1/temp5[51] , \MC_ARK_ARC_1_1/temp5[49] ,
         \MC_ARK_ARC_1_1/temp5[48] , \MC_ARK_ARC_1_1/temp5[44] ,
         \MC_ARK_ARC_1_1/temp5[43] , \MC_ARK_ARC_1_1/temp5[42] ,
         \MC_ARK_ARC_1_1/temp5[41] , \MC_ARK_ARC_1_1/temp5[38] ,
         \MC_ARK_ARC_1_1/temp5[37] , \MC_ARK_ARC_1_1/temp5[36] ,
         \MC_ARK_ARC_1_1/temp5[34] , \MC_ARK_ARC_1_1/temp5[32] ,
         \MC_ARK_ARC_1_1/temp5[31] , \MC_ARK_ARC_1_1/temp5[30] ,
         \MC_ARK_ARC_1_1/temp5[28] , \MC_ARK_ARC_1_1/temp5[27] ,
         \MC_ARK_ARC_1_1/temp5[24] , \MC_ARK_ARC_1_1/temp5[22] ,
         \MC_ARK_ARC_1_1/temp5[21] , \MC_ARK_ARC_1_1/temp5[19] ,
         \MC_ARK_ARC_1_1/temp5[18] , \MC_ARK_ARC_1_1/temp5[17] ,
         \MC_ARK_ARC_1_1/temp5[14] , \MC_ARK_ARC_1_1/temp5[12] ,
         \MC_ARK_ARC_1_1/temp5[10] , \MC_ARK_ARC_1_1/temp5[9] ,
         \MC_ARK_ARC_1_1/temp5[6] , \MC_ARK_ARC_1_1/temp5[2] ,
         \MC_ARK_ARC_1_1/temp4[190] , \MC_ARK_ARC_1_1/temp4[189] ,
         \MC_ARK_ARC_1_1/temp4[188] , \MC_ARK_ARC_1_1/temp4[187] ,
         \MC_ARK_ARC_1_1/temp4[186] , \MC_ARK_ARC_1_1/temp4[185] ,
         \MC_ARK_ARC_1_1/temp4[184] , \MC_ARK_ARC_1_1/temp4[183] ,
         \MC_ARK_ARC_1_1/temp4[181] , \MC_ARK_ARC_1_1/temp4[180] ,
         \MC_ARK_ARC_1_1/temp4[179] , \MC_ARK_ARC_1_1/temp4[178] ,
         \MC_ARK_ARC_1_1/temp4[177] , \MC_ARK_ARC_1_1/temp4[176] ,
         \MC_ARK_ARC_1_1/temp4[175] , \MC_ARK_ARC_1_1/temp4[174] ,
         \MC_ARK_ARC_1_1/temp4[173] , \MC_ARK_ARC_1_1/temp4[172] ,
         \MC_ARK_ARC_1_1/temp4[170] , \MC_ARK_ARC_1_1/temp4[169] ,
         \MC_ARK_ARC_1_1/temp4[168] , \MC_ARK_ARC_1_1/temp4[166] ,
         \MC_ARK_ARC_1_1/temp4[165] , \MC_ARK_ARC_1_1/temp4[164] ,
         \MC_ARK_ARC_1_1/temp4[163] , \MC_ARK_ARC_1_1/temp4[162] ,
         \MC_ARK_ARC_1_1/temp4[161] , \MC_ARK_ARC_1_1/temp4[160] ,
         \MC_ARK_ARC_1_1/temp4[159] , \MC_ARK_ARC_1_1/temp4[158] ,
         \MC_ARK_ARC_1_1/temp4[157] , \MC_ARK_ARC_1_1/temp4[156] ,
         \MC_ARK_ARC_1_1/temp4[155] , \MC_ARK_ARC_1_1/temp4[154] ,
         \MC_ARK_ARC_1_1/temp4[151] , \MC_ARK_ARC_1_1/temp4[150] ,
         \MC_ARK_ARC_1_1/temp4[149] , \MC_ARK_ARC_1_1/temp4[148] ,
         \MC_ARK_ARC_1_1/temp4[147] , \MC_ARK_ARC_1_1/temp4[146] ,
         \MC_ARK_ARC_1_1/temp4[145] , \MC_ARK_ARC_1_1/temp4[144] ,
         \MC_ARK_ARC_1_1/temp4[142] , \MC_ARK_ARC_1_1/temp4[141] ,
         \MC_ARK_ARC_1_1/temp4[140] , \MC_ARK_ARC_1_1/temp4[139] ,
         \MC_ARK_ARC_1_1/temp4[138] , \MC_ARK_ARC_1_1/temp4[137] ,
         \MC_ARK_ARC_1_1/temp4[136] , \MC_ARK_ARC_1_1/temp4[135] ,
         \MC_ARK_ARC_1_1/temp4[134] , \MC_ARK_ARC_1_1/temp4[133] ,
         \MC_ARK_ARC_1_1/temp4[132] , \MC_ARK_ARC_1_1/temp4[131] ,
         \MC_ARK_ARC_1_1/temp4[130] , \MC_ARK_ARC_1_1/temp4[129] ,
         \MC_ARK_ARC_1_1/temp4[128] , \MC_ARK_ARC_1_1/temp4[127] ,
         \MC_ARK_ARC_1_1/temp4[126] , \MC_ARK_ARC_1_1/temp4[125] ,
         \MC_ARK_ARC_1_1/temp4[124] , \MC_ARK_ARC_1_1/temp4[123] ,
         \MC_ARK_ARC_1_1/temp4[121] , \MC_ARK_ARC_1_1/temp4[120] ,
         \MC_ARK_ARC_1_1/temp4[119] , \MC_ARK_ARC_1_1/temp4[118] ,
         \MC_ARK_ARC_1_1/temp4[117] , \MC_ARK_ARC_1_1/temp4[114] ,
         \MC_ARK_ARC_1_1/temp4[113] , \MC_ARK_ARC_1_1/temp4[112] ,
         \MC_ARK_ARC_1_1/temp4[111] , \MC_ARK_ARC_1_1/temp4[109] ,
         \MC_ARK_ARC_1_1/temp4[108] , \MC_ARK_ARC_1_1/temp4[106] ,
         \MC_ARK_ARC_1_1/temp4[105] , \MC_ARK_ARC_1_1/temp4[104] ,
         \MC_ARK_ARC_1_1/temp4[103] , \MC_ARK_ARC_1_1/temp4[102] ,
         \MC_ARK_ARC_1_1/temp4[101] , \MC_ARK_ARC_1_1/temp4[100] ,
         \MC_ARK_ARC_1_1/temp4[99] , \MC_ARK_ARC_1_1/temp4[98] ,
         \MC_ARK_ARC_1_1/temp4[97] , \MC_ARK_ARC_1_1/temp4[96] ,
         \MC_ARK_ARC_1_1/temp4[95] , \MC_ARK_ARC_1_1/temp4[94] ,
         \MC_ARK_ARC_1_1/temp4[93] , \MC_ARK_ARC_1_1/temp4[92] ,
         \MC_ARK_ARC_1_1/temp4[91] , \MC_ARK_ARC_1_1/temp4[90] ,
         \MC_ARK_ARC_1_1/temp4[89] , \MC_ARK_ARC_1_1/temp4[88] ,
         \MC_ARK_ARC_1_1/temp4[87] , \MC_ARK_ARC_1_1/temp4[86] ,
         \MC_ARK_ARC_1_1/temp4[85] , \MC_ARK_ARC_1_1/temp4[84] ,
         \MC_ARK_ARC_1_1/temp4[82] , \MC_ARK_ARC_1_1/temp4[81] ,
         \MC_ARK_ARC_1_1/temp4[80] , \MC_ARK_ARC_1_1/temp4[79] ,
         \MC_ARK_ARC_1_1/temp4[78] , \MC_ARK_ARC_1_1/temp4[76] ,
         \MC_ARK_ARC_1_1/temp4[74] , \MC_ARK_ARC_1_1/temp4[73] ,
         \MC_ARK_ARC_1_1/temp4[72] , \MC_ARK_ARC_1_1/temp4[71] ,
         \MC_ARK_ARC_1_1/temp4[70] , \MC_ARK_ARC_1_1/temp4[69] ,
         \MC_ARK_ARC_1_1/temp4[68] , \MC_ARK_ARC_1_1/temp4[67] ,
         \MC_ARK_ARC_1_1/temp4[66] , \MC_ARK_ARC_1_1/temp4[65] ,
         \MC_ARK_ARC_1_1/temp4[64] , \MC_ARK_ARC_1_1/temp4[63] ,
         \MC_ARK_ARC_1_1/temp4[62] , \MC_ARK_ARC_1_1/temp4[61] ,
         \MC_ARK_ARC_1_1/temp4[60] , \MC_ARK_ARC_1_1/temp4[58] ,
         \MC_ARK_ARC_1_1/temp4[57] , \MC_ARK_ARC_1_1/temp4[56] ,
         \MC_ARK_ARC_1_1/temp4[55] , \MC_ARK_ARC_1_1/temp4[54] ,
         \MC_ARK_ARC_1_1/temp4[52] , \MC_ARK_ARC_1_1/temp4[51] ,
         \MC_ARK_ARC_1_1/temp4[50] , \MC_ARK_ARC_1_1/temp4[49] ,
         \MC_ARK_ARC_1_1/temp4[48] , \MC_ARK_ARC_1_1/temp4[47] ,
         \MC_ARK_ARC_1_1/temp4[46] , \MC_ARK_ARC_1_1/temp4[45] ,
         \MC_ARK_ARC_1_1/temp4[43] , \MC_ARK_ARC_1_1/temp4[42] ,
         \MC_ARK_ARC_1_1/temp4[41] , \MC_ARK_ARC_1_1/temp4[39] ,
         \MC_ARK_ARC_1_1/temp4[38] , \MC_ARK_ARC_1_1/temp4[37] ,
         \MC_ARK_ARC_1_1/temp4[36] , \MC_ARK_ARC_1_1/temp4[35] ,
         \MC_ARK_ARC_1_1/temp4[34] , \MC_ARK_ARC_1_1/temp4[33] ,
         \MC_ARK_ARC_1_1/temp4[32] , \MC_ARK_ARC_1_1/temp4[31] ,
         \MC_ARK_ARC_1_1/temp4[30] , \MC_ARK_ARC_1_1/temp4[28] ,
         \MC_ARK_ARC_1_1/temp4[27] , \MC_ARK_ARC_1_1/temp4[26] ,
         \MC_ARK_ARC_1_1/temp4[25] , \MC_ARK_ARC_1_1/temp4[24] ,
         \MC_ARK_ARC_1_1/temp4[22] , \MC_ARK_ARC_1_1/temp4[21] ,
         \MC_ARK_ARC_1_1/temp4[20] , \MC_ARK_ARC_1_1/temp4[19] ,
         \MC_ARK_ARC_1_1/temp4[18] , \MC_ARK_ARC_1_1/temp4[17] ,
         \MC_ARK_ARC_1_1/temp4[16] , \MC_ARK_ARC_1_1/temp4[14] ,
         \MC_ARK_ARC_1_1/temp4[13] , \MC_ARK_ARC_1_1/temp4[12] ,
         \MC_ARK_ARC_1_1/temp4[11] , \MC_ARK_ARC_1_1/temp4[10] ,
         \MC_ARK_ARC_1_1/temp4[9] , \MC_ARK_ARC_1_1/temp4[7] ,
         \MC_ARK_ARC_1_1/temp4[6] , \MC_ARK_ARC_1_1/temp4[5] ,
         \MC_ARK_ARC_1_1/temp4[4] , \MC_ARK_ARC_1_1/temp4[3] ,
         \MC_ARK_ARC_1_1/temp4[2] , \MC_ARK_ARC_1_1/temp4[1] ,
         \MC_ARK_ARC_1_1/temp4[0] , \MC_ARK_ARC_1_1/temp3[191] ,
         \MC_ARK_ARC_1_1/temp3[190] , \MC_ARK_ARC_1_1/temp3[189] ,
         \MC_ARK_ARC_1_1/temp3[186] , \MC_ARK_ARC_1_1/temp3[185] ,
         \MC_ARK_ARC_1_1/temp3[184] , \MC_ARK_ARC_1_1/temp3[183] ,
         \MC_ARK_ARC_1_1/temp3[180] , \MC_ARK_ARC_1_1/temp3[179] ,
         \MC_ARK_ARC_1_1/temp3[178] , \MC_ARK_ARC_1_1/temp3[176] ,
         \MC_ARK_ARC_1_1/temp3[175] , \MC_ARK_ARC_1_1/temp3[174] ,
         \MC_ARK_ARC_1_1/temp3[172] , \MC_ARK_ARC_1_1/temp3[169] ,
         \MC_ARK_ARC_1_1/temp3[168] , \MC_ARK_ARC_1_1/temp3[166] ,
         \MC_ARK_ARC_1_1/temp3[165] , \MC_ARK_ARC_1_1/temp3[164] ,
         \MC_ARK_ARC_1_1/temp3[162] , \MC_ARK_ARC_1_1/temp3[160] ,
         \MC_ARK_ARC_1_1/temp3[158] , \MC_ARK_ARC_1_1/temp3[157] ,
         \MC_ARK_ARC_1_1/temp3[156] , \MC_ARK_ARC_1_1/temp3[155] ,
         \MC_ARK_ARC_1_1/temp3[154] , \MC_ARK_ARC_1_1/temp3[151] ,
         \MC_ARK_ARC_1_1/temp3[150] , \MC_ARK_ARC_1_1/temp3[148] ,
         \MC_ARK_ARC_1_1/temp3[147] , \MC_ARK_ARC_1_1/temp3[145] ,
         \MC_ARK_ARC_1_1/temp3[144] , \MC_ARK_ARC_1_1/temp3[142] ,
         \MC_ARK_ARC_1_1/temp3[141] , \MC_ARK_ARC_1_1/temp3[140] ,
         \MC_ARK_ARC_1_1/temp3[139] , \MC_ARK_ARC_1_1/temp3[137] ,
         \MC_ARK_ARC_1_1/temp3[136] , \MC_ARK_ARC_1_1/temp3[134] ,
         \MC_ARK_ARC_1_1/temp3[133] , \MC_ARK_ARC_1_1/temp3[132] ,
         \MC_ARK_ARC_1_1/temp3[131] , \MC_ARK_ARC_1_1/temp3[130] ,
         \MC_ARK_ARC_1_1/temp3[129] , \MC_ARK_ARC_1_1/temp3[127] ,
         \MC_ARK_ARC_1_1/temp3[125] , \MC_ARK_ARC_1_1/temp3[124] ,
         \MC_ARK_ARC_1_1/temp3[123] , \MC_ARK_ARC_1_1/temp3[121] ,
         \MC_ARK_ARC_1_1/temp3[120] , \MC_ARK_ARC_1_1/temp3[119] ,
         \MC_ARK_ARC_1_1/temp3[118] , \MC_ARK_ARC_1_1/temp3[117] ,
         \MC_ARK_ARC_1_1/temp3[115] , \MC_ARK_ARC_1_1/temp3[114] ,
         \MC_ARK_ARC_1_1/temp3[112] , \MC_ARK_ARC_1_1/temp3[111] ,
         \MC_ARK_ARC_1_1/temp3[110] , \MC_ARK_ARC_1_1/temp3[109] ,
         \MC_ARK_ARC_1_1/temp3[108] , \MC_ARK_ARC_1_1/temp3[106] ,
         \MC_ARK_ARC_1_1/temp3[104] , \MC_ARK_ARC_1_1/temp3[103] ,
         \MC_ARK_ARC_1_1/temp3[102] , \MC_ARK_ARC_1_1/temp3[100] ,
         \MC_ARK_ARC_1_1/temp3[98] , \MC_ARK_ARC_1_1/temp3[96] ,
         \MC_ARK_ARC_1_1/temp3[95] , \MC_ARK_ARC_1_1/temp3[94] ,
         \MC_ARK_ARC_1_1/temp3[91] , \MC_ARK_ARC_1_1/temp3[89] ,
         \MC_ARK_ARC_1_1/temp3[88] , \MC_ARK_ARC_1_1/temp3[86] ,
         \MC_ARK_ARC_1_1/temp3[84] , \MC_ARK_ARC_1_1/temp3[82] ,
         \MC_ARK_ARC_1_1/temp3[81] , \MC_ARK_ARC_1_1/temp3[80] ,
         \MC_ARK_ARC_1_1/temp3[79] , \MC_ARK_ARC_1_1/temp3[78] ,
         \MC_ARK_ARC_1_1/temp3[77] , \MC_ARK_ARC_1_1/temp3[76] ,
         \MC_ARK_ARC_1_1/temp3[73] , \MC_ARK_ARC_1_1/temp3[72] ,
         \MC_ARK_ARC_1_1/temp3[71] , \MC_ARK_ARC_1_1/temp3[70] ,
         \MC_ARK_ARC_1_1/temp3[68] , \MC_ARK_ARC_1_1/temp3[67] ,
         \MC_ARK_ARC_1_1/temp3[66] , \MC_ARK_ARC_1_1/temp3[65] ,
         \MC_ARK_ARC_1_1/temp3[64] , \MC_ARK_ARC_1_1/temp3[63] ,
         \MC_ARK_ARC_1_1/temp3[62] , \MC_ARK_ARC_1_1/temp3[61] ,
         \MC_ARK_ARC_1_1/temp3[60] , \MC_ARK_ARC_1_1/temp3[58] ,
         \MC_ARK_ARC_1_1/temp3[57] , \MC_ARK_ARC_1_1/temp3[56] ,
         \MC_ARK_ARC_1_1/temp3[55] , \MC_ARK_ARC_1_1/temp3[54] ,
         \MC_ARK_ARC_1_1/temp3[51] , \MC_ARK_ARC_1_1/temp3[49] ,
         \MC_ARK_ARC_1_1/temp3[48] , \MC_ARK_ARC_1_1/temp3[47] ,
         \MC_ARK_ARC_1_1/temp3[46] , \MC_ARK_ARC_1_1/temp3[45] ,
         \MC_ARK_ARC_1_1/temp3[43] , \MC_ARK_ARC_1_1/temp3[42] ,
         \MC_ARK_ARC_1_1/temp3[39] , \MC_ARK_ARC_1_1/temp3[38] ,
         \MC_ARK_ARC_1_1/temp3[37] , \MC_ARK_ARC_1_1/temp3[36] ,
         \MC_ARK_ARC_1_1/temp3[33] , \MC_ARK_ARC_1_1/temp3[32] ,
         \MC_ARK_ARC_1_1/temp3[31] , \MC_ARK_ARC_1_1/temp3[28] ,
         \MC_ARK_ARC_1_1/temp3[25] , \MC_ARK_ARC_1_1/temp3[24] ,
         \MC_ARK_ARC_1_1/temp3[21] , \MC_ARK_ARC_1_1/temp3[20] ,
         \MC_ARK_ARC_1_1/temp3[19] , \MC_ARK_ARC_1_1/temp3[18] ,
         \MC_ARK_ARC_1_1/temp3[16] , \MC_ARK_ARC_1_1/temp3[15] ,
         \MC_ARK_ARC_1_1/temp3[13] , \MC_ARK_ARC_1_1/temp3[12] ,
         \MC_ARK_ARC_1_1/temp3[11] , \MC_ARK_ARC_1_1/temp3[10] ,
         \MC_ARK_ARC_1_1/temp3[9] , \MC_ARK_ARC_1_1/temp3[7] ,
         \MC_ARK_ARC_1_1/temp3[6] , \MC_ARK_ARC_1_1/temp3[5] ,
         \MC_ARK_ARC_1_1/temp3[3] , \MC_ARK_ARC_1_1/temp3[2] ,
         \MC_ARK_ARC_1_1/temp3[1] , \MC_ARK_ARC_1_1/temp3[0] ,
         \MC_ARK_ARC_1_1/temp2[190] , \MC_ARK_ARC_1_1/temp2[188] ,
         \MC_ARK_ARC_1_1/temp2[186] , \MC_ARK_ARC_1_1/temp2[184] ,
         \MC_ARK_ARC_1_1/temp2[182] , \MC_ARK_ARC_1_1/temp2[180] ,
         \MC_ARK_ARC_1_1/temp2[179] , \MC_ARK_ARC_1_1/temp2[178] ,
         \MC_ARK_ARC_1_1/temp2[175] , \MC_ARK_ARC_1_1/temp2[173] ,
         \MC_ARK_ARC_1_1/temp2[172] , \MC_ARK_ARC_1_1/temp2[171] ,
         \MC_ARK_ARC_1_1/temp2[168] , \MC_ARK_ARC_1_1/temp2[166] ,
         \MC_ARK_ARC_1_1/temp2[165] , \MC_ARK_ARC_1_1/temp2[163] ,
         \MC_ARK_ARC_1_1/temp2[161] , \MC_ARK_ARC_1_1/temp2[160] ,
         \MC_ARK_ARC_1_1/temp2[159] , \MC_ARK_ARC_1_1/temp2[158] ,
         \MC_ARK_ARC_1_1/temp2[156] , \MC_ARK_ARC_1_1/temp2[155] ,
         \MC_ARK_ARC_1_1/temp2[153] , \MC_ARK_ARC_1_1/temp2[150] ,
         \MC_ARK_ARC_1_1/temp2[149] , \MC_ARK_ARC_1_1/temp2[148] ,
         \MC_ARK_ARC_1_1/temp2[147] , \MC_ARK_ARC_1_1/temp2[145] ,
         \MC_ARK_ARC_1_1/temp2[142] , \MC_ARK_ARC_1_1/temp2[139] ,
         \MC_ARK_ARC_1_1/temp2[138] , \MC_ARK_ARC_1_1/temp2[136] ,
         \MC_ARK_ARC_1_1/temp2[133] , \MC_ARK_ARC_1_1/temp2[130] ,
         \MC_ARK_ARC_1_1/temp2[128] , \MC_ARK_ARC_1_1/temp2[127] ,
         \MC_ARK_ARC_1_1/temp2[126] , \MC_ARK_ARC_1_1/temp2[125] ,
         \MC_ARK_ARC_1_1/temp2[123] , \MC_ARK_ARC_1_1/temp2[120] ,
         \MC_ARK_ARC_1_1/temp2[118] , \MC_ARK_ARC_1_1/temp2[117] ,
         \MC_ARK_ARC_1_1/temp2[116] , \MC_ARK_ARC_1_1/temp2[114] ,
         \MC_ARK_ARC_1_1/temp2[112] , \MC_ARK_ARC_1_1/temp2[109] ,
         \MC_ARK_ARC_1_1/temp2[108] , \MC_ARK_ARC_1_1/temp2[107] ,
         \MC_ARK_ARC_1_1/temp2[106] , \MC_ARK_ARC_1_1/temp2[104] ,
         \MC_ARK_ARC_1_1/temp2[103] , \MC_ARK_ARC_1_1/temp2[102] ,
         \MC_ARK_ARC_1_1/temp2[100] , \MC_ARK_ARC_1_1/temp2[97] ,
         \MC_ARK_ARC_1_1/temp2[96] , \MC_ARK_ARC_1_1/temp2[95] ,
         \MC_ARK_ARC_1_1/temp2[94] , \MC_ARK_ARC_1_1/temp2[93] ,
         \MC_ARK_ARC_1_1/temp2[88] , \MC_ARK_ARC_1_1/temp2[85] ,
         \MC_ARK_ARC_1_1/temp2[84] , \MC_ARK_ARC_1_1/temp2[82] ,
         \MC_ARK_ARC_1_1/temp2[81] , \MC_ARK_ARC_1_1/temp2[78] ,
         \MC_ARK_ARC_1_1/temp2[77] , \MC_ARK_ARC_1_1/temp2[76] ,
         \MC_ARK_ARC_1_1/temp2[75] , \MC_ARK_ARC_1_1/temp2[73] ,
         \MC_ARK_ARC_1_1/temp2[72] , \MC_ARK_ARC_1_1/temp2[71] ,
         \MC_ARK_ARC_1_1/temp2[70] , \MC_ARK_ARC_1_1/temp2[69] ,
         \MC_ARK_ARC_1_1/temp2[68] , \MC_ARK_ARC_1_1/temp2[64] ,
         \MC_ARK_ARC_1_1/temp2[63] , \MC_ARK_ARC_1_1/temp2[62] ,
         \MC_ARK_ARC_1_1/temp2[61] , \MC_ARK_ARC_1_1/temp2[60] ,
         \MC_ARK_ARC_1_1/temp2[58] , \MC_ARK_ARC_1_1/temp2[57] ,
         \MC_ARK_ARC_1_1/temp2[56] , \MC_ARK_ARC_1_1/temp2[55] ,
         \MC_ARK_ARC_1_1/temp2[54] , \MC_ARK_ARC_1_1/temp2[51] ,
         \MC_ARK_ARC_1_1/temp2[49] , \MC_ARK_ARC_1_1/temp2[48] ,
         \MC_ARK_ARC_1_1/temp2[43] , \MC_ARK_ARC_1_1/temp2[42] ,
         \MC_ARK_ARC_1_1/temp2[41] , \MC_ARK_ARC_1_1/temp2[37] ,
         \MC_ARK_ARC_1_1/temp2[34] , \MC_ARK_ARC_1_1/temp2[33] ,
         \MC_ARK_ARC_1_1/temp2[32] , \MC_ARK_ARC_1_1/temp2[30] ,
         \MC_ARK_ARC_1_1/temp2[29] , \MC_ARK_ARC_1_1/temp2[27] ,
         \MC_ARK_ARC_1_1/temp2[25] , \MC_ARK_ARC_1_1/temp2[24] ,
         \MC_ARK_ARC_1_1/temp2[22] , \MC_ARK_ARC_1_1/temp2[21] ,
         \MC_ARK_ARC_1_1/temp2[19] , \MC_ARK_ARC_1_1/temp2[18] ,
         \MC_ARK_ARC_1_1/temp2[13] , \MC_ARK_ARC_1_1/temp2[12] ,
         \MC_ARK_ARC_1_1/temp2[9] , \MC_ARK_ARC_1_1/temp2[7] ,
         \MC_ARK_ARC_1_1/temp2[6] , \MC_ARK_ARC_1_1/temp2[5] ,
         \MC_ARK_ARC_1_1/temp2[4] , \MC_ARK_ARC_1_1/temp2[3] ,
         \MC_ARK_ARC_1_1/temp2[1] , \MC_ARK_ARC_1_1/temp1[190] ,
         \MC_ARK_ARC_1_1/temp1[189] , \MC_ARK_ARC_1_1/temp1[187] ,
         \MC_ARK_ARC_1_1/temp1[186] , \MC_ARK_ARC_1_1/temp1[184] ,
         \MC_ARK_ARC_1_1/temp1[182] , \MC_ARK_ARC_1_1/temp1[179] ,
         \MC_ARK_ARC_1_1/temp1[178] , \MC_ARK_ARC_1_1/temp1[175] ,
         \MC_ARK_ARC_1_1/temp1[174] , \MC_ARK_ARC_1_1/temp1[173] ,
         \MC_ARK_ARC_1_1/temp1[171] , \MC_ARK_ARC_1_1/temp1[168] ,
         \MC_ARK_ARC_1_1/temp1[166] , \MC_ARK_ARC_1_1/temp1[165] ,
         \MC_ARK_ARC_1_1/temp1[160] , \MC_ARK_ARC_1_1/temp1[159] ,
         \MC_ARK_ARC_1_1/temp1[158] , \MC_ARK_ARC_1_1/temp1[156] ,
         \MC_ARK_ARC_1_1/temp1[153] , \MC_ARK_ARC_1_1/temp1[151] ,
         \MC_ARK_ARC_1_1/temp1[149] , \MC_ARK_ARC_1_1/temp1[148] ,
         \MC_ARK_ARC_1_1/temp1[147] , \MC_ARK_ARC_1_1/temp1[146] ,
         \MC_ARK_ARC_1_1/temp1[144] , \MC_ARK_ARC_1_1/temp1[141] ,
         \MC_ARK_ARC_1_1/temp1[139] , \MC_ARK_ARC_1_1/temp1[138] ,
         \MC_ARK_ARC_1_1/temp1[136] , \MC_ARK_ARC_1_1/temp1[134] ,
         \MC_ARK_ARC_1_1/temp1[133] , \MC_ARK_ARC_1_1/temp1[132] ,
         \MC_ARK_ARC_1_1/temp1[127] , \MC_ARK_ARC_1_1/temp1[126] ,
         \MC_ARK_ARC_1_1/temp1[125] , \MC_ARK_ARC_1_1/temp1[123] ,
         \MC_ARK_ARC_1_1/temp1[120] , \MC_ARK_ARC_1_1/temp1[118] ,
         \MC_ARK_ARC_1_1/temp1[114] , \MC_ARK_ARC_1_1/temp1[112] ,
         \MC_ARK_ARC_1_1/temp1[109] , \MC_ARK_ARC_1_1/temp1[106] ,
         \MC_ARK_ARC_1_1/temp1[104] , \MC_ARK_ARC_1_1/temp1[103] ,
         \MC_ARK_ARC_1_1/temp1[102] , \MC_ARK_ARC_1_1/temp1[99] ,
         \MC_ARK_ARC_1_1/temp1[96] , \MC_ARK_ARC_1_1/temp1[94] ,
         \MC_ARK_ARC_1_1/temp1[93] , \MC_ARK_ARC_1_1/temp1[91] ,
         \MC_ARK_ARC_1_1/temp1[90] , \MC_ARK_ARC_1_1/temp1[89] ,
         \MC_ARK_ARC_1_1/temp1[88] , \MC_ARK_ARC_1_1/temp1[83] ,
         \MC_ARK_ARC_1_1/temp1[82] , \MC_ARK_ARC_1_1/temp1[81] ,
         \MC_ARK_ARC_1_1/temp1[78] , \MC_ARK_ARC_1_1/temp1[76] ,
         \MC_ARK_ARC_1_1/temp1[75] , \MC_ARK_ARC_1_1/temp1[74] ,
         \MC_ARK_ARC_1_1/temp1[73] , \MC_ARK_ARC_1_1/temp1[72] ,
         \MC_ARK_ARC_1_1/temp1[71] , \MC_ARK_ARC_1_1/temp1[66] ,
         \MC_ARK_ARC_1_1/temp1[64] , \MC_ARK_ARC_1_1/temp1[63] ,
         \MC_ARK_ARC_1_1/temp1[62] , \MC_ARK_ARC_1_1/temp1[61] ,
         \MC_ARK_ARC_1_1/temp1[60] , \MC_ARK_ARC_1_1/temp1[58] ,
         \MC_ARK_ARC_1_1/temp1[55] , \MC_ARK_ARC_1_1/temp1[54] ,
         \MC_ARK_ARC_1_1/temp1[53] , \MC_ARK_ARC_1_1/temp1[52] ,
         \MC_ARK_ARC_1_1/temp1[51] , \MC_ARK_ARC_1_1/temp1[50] ,
         \MC_ARK_ARC_1_1/temp1[49] , \MC_ARK_ARC_1_1/temp1[48] ,
         \MC_ARK_ARC_1_1/temp1[46] , \MC_ARK_ARC_1_1/temp1[44] ,
         \MC_ARK_ARC_1_1/temp1[43] , \MC_ARK_ARC_1_1/temp1[42] ,
         \MC_ARK_ARC_1_1/temp1[40] , \MC_ARK_ARC_1_1/temp1[39] ,
         \MC_ARK_ARC_1_1/temp1[38] , \MC_ARK_ARC_1_1/temp1[37] ,
         \MC_ARK_ARC_1_1/temp1[36] , \MC_ARK_ARC_1_1/temp1[35] ,
         \MC_ARK_ARC_1_1/temp1[34] , \MC_ARK_ARC_1_1/temp1[33] ,
         \MC_ARK_ARC_1_1/temp1[31] , \MC_ARK_ARC_1_1/temp1[30] ,
         \MC_ARK_ARC_1_1/temp1[29] , \MC_ARK_ARC_1_1/temp1[28] ,
         \MC_ARK_ARC_1_1/temp1[26] , \MC_ARK_ARC_1_1/temp1[25] ,
         \MC_ARK_ARC_1_1/temp1[24] , \MC_ARK_ARC_1_1/temp1[22] ,
         \MC_ARK_ARC_1_1/temp1[21] , \MC_ARK_ARC_1_1/temp1[18] ,
         \MC_ARK_ARC_1_1/temp1[16] , \MC_ARK_ARC_1_1/temp1[14] ,
         \MC_ARK_ARC_1_1/temp1[12] , \MC_ARK_ARC_1_1/temp1[10] ,
         \MC_ARK_ARC_1_1/temp1[7] , \MC_ARK_ARC_1_1/temp1[4] ,
         \MC_ARK_ARC_1_1/temp1[3] , \MC_ARK_ARC_1_1/temp1[1] ,
         \MC_ARK_ARC_1_1/buf_keyinput[51] ,
         \MC_ARK_ARC_1_1/buf_datainput[187] ,
         \MC_ARK_ARC_1_1/buf_datainput[186] ,
         \MC_ARK_ARC_1_1/buf_datainput[185] ,
         \MC_ARK_ARC_1_1/buf_datainput[179] ,
         \MC_ARK_ARC_1_1/buf_datainput[170] ,
         \MC_ARK_ARC_1_1/buf_datainput[169] ,
         \MC_ARK_ARC_1_1/buf_datainput[163] ,
         \MC_ARK_ARC_1_1/buf_datainput[160] ,
         \MC_ARK_ARC_1_1/buf_datainput[159] ,
         \MC_ARK_ARC_1_1/buf_datainput[155] ,
         \MC_ARK_ARC_1_1/buf_datainput[153] ,
         \MC_ARK_ARC_1_1/buf_datainput[139] ,
         \MC_ARK_ARC_1_1/buf_datainput[123] ,
         \MC_ARK_ARC_1_1/buf_datainput[110] ,
         \MC_ARK_ARC_1_1/buf_datainput[105] ,
         \MC_ARK_ARC_1_1/buf_datainput[101] ,
         \MC_ARK_ARC_1_1/buf_datainput[100] ,
         \MC_ARK_ARC_1_1/buf_datainput[99] ,
         \MC_ARK_ARC_1_1/buf_datainput[95] ,
         \MC_ARK_ARC_1_1/buf_datainput[89] ,
         \MC_ARK_ARC_1_1/buf_datainput[84] ,
         \MC_ARK_ARC_1_1/buf_datainput[80] ,
         \MC_ARK_ARC_1_1/buf_datainput[74] ,
         \MC_ARK_ARC_1_1/buf_datainput[66] ,
         \MC_ARK_ARC_1_1/buf_datainput[63] ,
         \MC_ARK_ARC_1_1/buf_datainput[42] ,
         \MC_ARK_ARC_1_1/buf_datainput[41] ,
         \MC_ARK_ARC_1_1/buf_datainput[38] ,
         \MC_ARK_ARC_1_1/buf_datainput[35] ,
         \MC_ARK_ARC_1_1/buf_datainput[31] ,
         \MC_ARK_ARC_1_1/buf_datainput[29] ,
         \MC_ARK_ARC_1_1/buf_datainput[28] ,
         \MC_ARK_ARC_1_1/buf_datainput[25] ,
         \MC_ARK_ARC_1_1/buf_datainput[22] , \MC_ARK_ARC_1_1/buf_datainput[9] ,
         \MC_ARK_ARC_1_1/buf_datainput[1] , \MC_ARK_ARC_1_2/buf_output[191] ,
         \MC_ARK_ARC_1_2/buf_output[190] , \MC_ARK_ARC_1_2/buf_output[189] ,
         \MC_ARK_ARC_1_2/buf_output[188] , \MC_ARK_ARC_1_2/buf_output[187] ,
         \MC_ARK_ARC_1_2/buf_output[186] , \MC_ARK_ARC_1_2/buf_output[185] ,
         \MC_ARK_ARC_1_2/buf_output[184] , \MC_ARK_ARC_1_2/buf_output[183] ,
         \MC_ARK_ARC_1_2/buf_output[182] , \MC_ARK_ARC_1_2/buf_output[181] ,
         \MC_ARK_ARC_1_2/buf_output[180] , \MC_ARK_ARC_1_2/buf_output[179] ,
         \MC_ARK_ARC_1_2/buf_output[178] , \MC_ARK_ARC_1_2/buf_output[177] ,
         \MC_ARK_ARC_1_2/buf_output[176] , \MC_ARK_ARC_1_2/buf_output[175] ,
         \MC_ARK_ARC_1_2/buf_output[174] , \MC_ARK_ARC_1_2/buf_output[173] ,
         \MC_ARK_ARC_1_2/buf_output[172] , \MC_ARK_ARC_1_2/buf_output[171] ,
         \MC_ARK_ARC_1_2/buf_output[170] , \MC_ARK_ARC_1_2/buf_output[169] ,
         \MC_ARK_ARC_1_2/buf_output[168] , \MC_ARK_ARC_1_2/buf_output[166] ,
         \MC_ARK_ARC_1_2/buf_output[165] , \MC_ARK_ARC_1_2/buf_output[164] ,
         \MC_ARK_ARC_1_2/buf_output[163] , \MC_ARK_ARC_1_2/buf_output[162] ,
         \MC_ARK_ARC_1_2/buf_output[161] , \MC_ARK_ARC_1_2/buf_output[160] ,
         \MC_ARK_ARC_1_2/buf_output[159] , \MC_ARK_ARC_1_2/buf_output[158] ,
         \MC_ARK_ARC_1_2/buf_output[157] , \MC_ARK_ARC_1_2/buf_output[156] ,
         \MC_ARK_ARC_1_2/buf_output[155] , \MC_ARK_ARC_1_2/buf_output[154] ,
         \MC_ARK_ARC_1_2/buf_output[153] , \MC_ARK_ARC_1_2/buf_output[152] ,
         \MC_ARK_ARC_1_2/buf_output[151] , \MC_ARK_ARC_1_2/buf_output[150] ,
         \MC_ARK_ARC_1_2/buf_output[149] , \MC_ARK_ARC_1_2/buf_output[148] ,
         \MC_ARK_ARC_1_2/buf_output[147] , \MC_ARK_ARC_1_2/buf_output[146] ,
         \MC_ARK_ARC_1_2/buf_output[145] , \MC_ARK_ARC_1_2/buf_output[144] ,
         \MC_ARK_ARC_1_2/buf_output[142] , \MC_ARK_ARC_1_2/buf_output[141] ,
         \MC_ARK_ARC_1_2/buf_output[140] , \MC_ARK_ARC_1_2/buf_output[139] ,
         \MC_ARK_ARC_1_2/buf_output[138] , \MC_ARK_ARC_1_2/buf_output[137] ,
         \MC_ARK_ARC_1_2/buf_output[136] , \MC_ARK_ARC_1_2/buf_output[134] ,
         \MC_ARK_ARC_1_2/buf_output[133] , \MC_ARK_ARC_1_2/buf_output[132] ,
         \MC_ARK_ARC_1_2/buf_output[131] , \MC_ARK_ARC_1_2/buf_output[130] ,
         \MC_ARK_ARC_1_2/buf_output[129] , \MC_ARK_ARC_1_2/buf_output[128] ,
         \MC_ARK_ARC_1_2/buf_output[127] , \MC_ARK_ARC_1_2/buf_output[126] ,
         \MC_ARK_ARC_1_2/buf_output[125] , \MC_ARK_ARC_1_2/buf_output[124] ,
         \MC_ARK_ARC_1_2/buf_output[123] , \MC_ARK_ARC_1_2/buf_output[122] ,
         \MC_ARK_ARC_1_2/buf_output[121] , \MC_ARK_ARC_1_2/buf_output[120] ,
         \MC_ARK_ARC_1_2/buf_output[119] , \MC_ARK_ARC_1_2/buf_output[118] ,
         \MC_ARK_ARC_1_2/buf_output[117] , \MC_ARK_ARC_1_2/buf_output[116] ,
         \MC_ARK_ARC_1_2/buf_output[115] , \MC_ARK_ARC_1_2/buf_output[114] ,
         \MC_ARK_ARC_1_2/buf_output[113] , \MC_ARK_ARC_1_2/buf_output[112] ,
         \MC_ARK_ARC_1_2/buf_output[111] , \MC_ARK_ARC_1_2/buf_output[110] ,
         \MC_ARK_ARC_1_2/buf_output[109] , \MC_ARK_ARC_1_2/buf_output[108] ,
         \MC_ARK_ARC_1_2/buf_output[106] , \MC_ARK_ARC_1_2/buf_output[105] ,
         \MC_ARK_ARC_1_2/buf_output[104] , \MC_ARK_ARC_1_2/buf_output[103] ,
         \MC_ARK_ARC_1_2/buf_output[102] , \MC_ARK_ARC_1_2/buf_output[101] ,
         \MC_ARK_ARC_1_2/buf_output[100] , \MC_ARK_ARC_1_2/buf_output[99] ,
         \MC_ARK_ARC_1_2/buf_output[98] , \MC_ARK_ARC_1_2/buf_output[97] ,
         \MC_ARK_ARC_1_2/buf_output[96] , \MC_ARK_ARC_1_2/buf_output[95] ,
         \MC_ARK_ARC_1_2/buf_output[94] , \MC_ARK_ARC_1_2/buf_output[93] ,
         \MC_ARK_ARC_1_2/buf_output[92] , \MC_ARK_ARC_1_2/buf_output[91] ,
         \MC_ARK_ARC_1_2/buf_output[90] , \MC_ARK_ARC_1_2/buf_output[88] ,
         \MC_ARK_ARC_1_2/buf_output[87] , \MC_ARK_ARC_1_2/buf_output[86] ,
         \MC_ARK_ARC_1_2/buf_output[85] , \MC_ARK_ARC_1_2/buf_output[84] ,
         \MC_ARK_ARC_1_2/buf_output[83] , \MC_ARK_ARC_1_2/buf_output[82] ,
         \MC_ARK_ARC_1_2/buf_output[81] , \MC_ARK_ARC_1_2/buf_output[80] ,
         \MC_ARK_ARC_1_2/buf_output[79] , \MC_ARK_ARC_1_2/buf_output[78] ,
         \MC_ARK_ARC_1_2/buf_output[77] , \MC_ARK_ARC_1_2/buf_output[76] ,
         \MC_ARK_ARC_1_2/buf_output[75] , \MC_ARK_ARC_1_2/buf_output[74] ,
         \MC_ARK_ARC_1_2/buf_output[73] , \MC_ARK_ARC_1_2/buf_output[72] ,
         \MC_ARK_ARC_1_2/buf_output[70] , \MC_ARK_ARC_1_2/buf_output[69] ,
         \MC_ARK_ARC_1_2/buf_output[68] , \MC_ARK_ARC_1_2/buf_output[67] ,
         \MC_ARK_ARC_1_2/buf_output[66] , \MC_ARK_ARC_1_2/buf_output[65] ,
         \MC_ARK_ARC_1_2/buf_output[64] , \MC_ARK_ARC_1_2/buf_output[63] ,
         \MC_ARK_ARC_1_2/buf_output[62] , \MC_ARK_ARC_1_2/buf_output[61] ,
         \MC_ARK_ARC_1_2/buf_output[60] , \MC_ARK_ARC_1_2/buf_output[58] ,
         \MC_ARK_ARC_1_2/buf_output[57] , \MC_ARK_ARC_1_2/buf_output[56] ,
         \MC_ARK_ARC_1_2/buf_output[55] , \MC_ARK_ARC_1_2/buf_output[54] ,
         \MC_ARK_ARC_1_2/buf_output[53] , \MC_ARK_ARC_1_2/buf_output[51] ,
         \MC_ARK_ARC_1_2/buf_output[50] , \MC_ARK_ARC_1_2/buf_output[49] ,
         \MC_ARK_ARC_1_2/buf_output[48] , \MC_ARK_ARC_1_2/buf_output[47] ,
         \MC_ARK_ARC_1_2/buf_output[46] , \MC_ARK_ARC_1_2/buf_output[45] ,
         \MC_ARK_ARC_1_2/buf_output[44] , \MC_ARK_ARC_1_2/buf_output[43] ,
         \MC_ARK_ARC_1_2/buf_output[42] , \MC_ARK_ARC_1_2/buf_output[40] ,
         \MC_ARK_ARC_1_2/buf_output[39] , \MC_ARK_ARC_1_2/buf_output[38] ,
         \MC_ARK_ARC_1_2/buf_output[37] , \MC_ARK_ARC_1_2/buf_output[36] ,
         \MC_ARK_ARC_1_2/buf_output[35] , \MC_ARK_ARC_1_2/buf_output[34] ,
         \MC_ARK_ARC_1_2/buf_output[33] , \MC_ARK_ARC_1_2/buf_output[32] ,
         \MC_ARK_ARC_1_2/buf_output[31] , \MC_ARK_ARC_1_2/buf_output[30] ,
         \MC_ARK_ARC_1_2/buf_output[29] , \MC_ARK_ARC_1_2/buf_output[28] ,
         \MC_ARK_ARC_1_2/buf_output[27] , \MC_ARK_ARC_1_2/buf_output[26] ,
         \MC_ARK_ARC_1_2/buf_output[25] , \MC_ARK_ARC_1_2/buf_output[24] ,
         \MC_ARK_ARC_1_2/buf_output[23] , \MC_ARK_ARC_1_2/buf_output[22] ,
         \MC_ARK_ARC_1_2/buf_output[21] , \MC_ARK_ARC_1_2/buf_output[20] ,
         \MC_ARK_ARC_1_2/buf_output[19] , \MC_ARK_ARC_1_2/buf_output[18] ,
         \MC_ARK_ARC_1_2/buf_output[16] , \MC_ARK_ARC_1_2/buf_output[15] ,
         \MC_ARK_ARC_1_2/buf_output[14] , \MC_ARK_ARC_1_2/buf_output[13] ,
         \MC_ARK_ARC_1_2/buf_output[12] , \MC_ARK_ARC_1_2/buf_output[11] ,
         \MC_ARK_ARC_1_2/buf_output[10] , \MC_ARK_ARC_1_2/buf_output[9] ,
         \MC_ARK_ARC_1_2/buf_output[8] , \MC_ARK_ARC_1_2/buf_output[7] ,
         \MC_ARK_ARC_1_2/buf_output[6] , \MC_ARK_ARC_1_2/buf_output[4] ,
         \MC_ARK_ARC_1_2/buf_output[3] , \MC_ARK_ARC_1_2/buf_output[2] ,
         \MC_ARK_ARC_1_2/buf_output[1] , \MC_ARK_ARC_1_2/buf_output[0] ,
         \MC_ARK_ARC_1_2/temp6[191] , \MC_ARK_ARC_1_2/temp6[187] ,
         \MC_ARK_ARC_1_2/temp6[186] , \MC_ARK_ARC_1_2/temp6[185] ,
         \MC_ARK_ARC_1_2/temp6[184] , \MC_ARK_ARC_1_2/temp6[182] ,
         \MC_ARK_ARC_1_2/temp6[181] , \MC_ARK_ARC_1_2/temp6[179] ,
         \MC_ARK_ARC_1_2/temp6[178] , \MC_ARK_ARC_1_2/temp6[177] ,
         \MC_ARK_ARC_1_2/temp6[174] , \MC_ARK_ARC_1_2/temp6[172] ,
         \MC_ARK_ARC_1_2/temp6[171] , \MC_ARK_ARC_1_2/temp6[170] ,
         \MC_ARK_ARC_1_2/temp6[169] , \MC_ARK_ARC_1_2/temp6[168] ,
         \MC_ARK_ARC_1_2/temp6[166] , \MC_ARK_ARC_1_2/temp6[162] ,
         \MC_ARK_ARC_1_2/temp6[161] , \MC_ARK_ARC_1_2/temp6[160] ,
         \MC_ARK_ARC_1_2/temp6[156] , \MC_ARK_ARC_1_2/temp6[152] ,
         \MC_ARK_ARC_1_2/temp6[151] , \MC_ARK_ARC_1_2/temp6[150] ,
         \MC_ARK_ARC_1_2/temp6[148] , \MC_ARK_ARC_1_2/temp6[147] ,
         \MC_ARK_ARC_1_2/temp6[145] , \MC_ARK_ARC_1_2/temp6[143] ,
         \MC_ARK_ARC_1_2/temp6[141] , \MC_ARK_ARC_1_2/temp6[140] ,
         \MC_ARK_ARC_1_2/temp6[136] , \MC_ARK_ARC_1_2/temp6[135] ,
         \MC_ARK_ARC_1_2/temp6[131] , \MC_ARK_ARC_1_2/temp6[126] ,
         \MC_ARK_ARC_1_2/temp6[124] , \MC_ARK_ARC_1_2/temp6[123] ,
         \MC_ARK_ARC_1_2/temp6[118] , \MC_ARK_ARC_1_2/temp6[114] ,
         \MC_ARK_ARC_1_2/temp6[113] , \MC_ARK_ARC_1_2/temp6[109] ,
         \MC_ARK_ARC_1_2/temp6[108] , \MC_ARK_ARC_1_2/temp6[106] ,
         \MC_ARK_ARC_1_2/temp6[101] , \MC_ARK_ARC_1_2/temp6[97] ,
         \MC_ARK_ARC_1_2/temp6[96] , \MC_ARK_ARC_1_2/temp6[94] ,
         \MC_ARK_ARC_1_2/temp6[93] , \MC_ARK_ARC_1_2/temp6[88] ,
         \MC_ARK_ARC_1_2/temp6[86] , \MC_ARK_ARC_1_2/temp6[85] ,
         \MC_ARK_ARC_1_2/temp6[84] , \MC_ARK_ARC_1_2/temp6[82] ,
         \MC_ARK_ARC_1_2/temp6[81] , \MC_ARK_ARC_1_2/temp6[80] ,
         \MC_ARK_ARC_1_2/temp6[79] , \MC_ARK_ARC_1_2/temp6[78] ,
         \MC_ARK_ARC_1_2/temp6[77] , \MC_ARK_ARC_1_2/temp6[72] ,
         \MC_ARK_ARC_1_2/temp6[71] , \MC_ARK_ARC_1_2/temp6[70] ,
         \MC_ARK_ARC_1_2/temp6[67] , \MC_ARK_ARC_1_2/temp6[66] ,
         \MC_ARK_ARC_1_2/temp6[65] , \MC_ARK_ARC_1_2/temp6[60] ,
         \MC_ARK_ARC_1_2/temp6[54] , \MC_ARK_ARC_1_2/temp6[53] ,
         \MC_ARK_ARC_1_2/temp6[50] , \MC_ARK_ARC_1_2/temp6[46] ,
         \MC_ARK_ARC_1_2/temp6[45] , \MC_ARK_ARC_1_2/temp6[42] ,
         \MC_ARK_ARC_1_2/temp6[41] , \MC_ARK_ARC_1_2/temp6[40] ,
         \MC_ARK_ARC_1_2/temp6[38] , \MC_ARK_ARC_1_2/temp6[36] ,
         \MC_ARK_ARC_1_2/temp6[28] , \MC_ARK_ARC_1_2/temp6[25] ,
         \MC_ARK_ARC_1_2/temp6[24] , \MC_ARK_ARC_1_2/temp6[21] ,
         \MC_ARK_ARC_1_2/temp6[17] , \MC_ARK_ARC_1_2/temp6[16] ,
         \MC_ARK_ARC_1_2/temp6[14] , \MC_ARK_ARC_1_2/temp6[13] ,
         \MC_ARK_ARC_1_2/temp6[7] , \MC_ARK_ARC_1_2/temp6[2] ,
         \MC_ARK_ARC_1_2/temp6[0] , \MC_ARK_ARC_1_2/temp5[190] ,
         \MC_ARK_ARC_1_2/temp5[189] , \MC_ARK_ARC_1_2/temp5[187] ,
         \MC_ARK_ARC_1_2/temp5[186] , \MC_ARK_ARC_1_2/temp5[184] ,
         \MC_ARK_ARC_1_2/temp5[181] , \MC_ARK_ARC_1_2/temp5[180] ,
         \MC_ARK_ARC_1_2/temp5[178] , \MC_ARK_ARC_1_2/temp5[174] ,
         \MC_ARK_ARC_1_2/temp5[173] , \MC_ARK_ARC_1_2/temp5[172] ,
         \MC_ARK_ARC_1_2/temp5[168] , \MC_ARK_ARC_1_2/temp5[165] ,
         \MC_ARK_ARC_1_2/temp5[164] , \MC_ARK_ARC_1_2/temp5[162] ,
         \MC_ARK_ARC_1_2/temp5[161] , \MC_ARK_ARC_1_2/temp5[160] ,
         \MC_ARK_ARC_1_2/temp5[158] , \MC_ARK_ARC_1_2/temp5[157] ,
         \MC_ARK_ARC_1_2/temp5[154] , \MC_ARK_ARC_1_2/temp5[151] ,
         \MC_ARK_ARC_1_2/temp5[150] , \MC_ARK_ARC_1_2/temp5[145] ,
         \MC_ARK_ARC_1_2/temp5[144] , \MC_ARK_ARC_1_2/temp5[143] ,
         \MC_ARK_ARC_1_2/temp5[142] , \MC_ARK_ARC_1_2/temp5[139] ,
         \MC_ARK_ARC_1_2/temp5[138] , \MC_ARK_ARC_1_2/temp5[136] ,
         \MC_ARK_ARC_1_2/temp5[132] , \MC_ARK_ARC_1_2/temp5[131] ,
         \MC_ARK_ARC_1_2/temp5[127] , \MC_ARK_ARC_1_2/temp5[126] ,
         \MC_ARK_ARC_1_2/temp5[125] , \MC_ARK_ARC_1_2/temp5[124] ,
         \MC_ARK_ARC_1_2/temp5[123] , \MC_ARK_ARC_1_2/temp5[121] ,
         \MC_ARK_ARC_1_2/temp5[115] , \MC_ARK_ARC_1_2/temp5[114] ,
         \MC_ARK_ARC_1_2/temp5[109] , \MC_ARK_ARC_1_2/temp5[108] ,
         \MC_ARK_ARC_1_2/temp5[106] , \MC_ARK_ARC_1_2/temp5[103] ,
         \MC_ARK_ARC_1_2/temp5[102] , \MC_ARK_ARC_1_2/temp5[100] ,
         \MC_ARK_ARC_1_2/temp5[97] , \MC_ARK_ARC_1_2/temp5[92] ,
         \MC_ARK_ARC_1_2/temp5[91] , \MC_ARK_ARC_1_2/temp5[86] ,
         \MC_ARK_ARC_1_2/temp5[84] , \MC_ARK_ARC_1_2/temp5[80] ,
         \MC_ARK_ARC_1_2/temp5[79] , \MC_ARK_ARC_1_2/temp5[78] ,
         \MC_ARK_ARC_1_2/temp5[77] , \MC_ARK_ARC_1_2/temp5[76] ,
         \MC_ARK_ARC_1_2/temp5[74] , \MC_ARK_ARC_1_2/temp5[71] ,
         \MC_ARK_ARC_1_2/temp5[69] , \MC_ARK_ARC_1_2/temp5[66] ,
         \MC_ARK_ARC_1_2/temp5[59] , \MC_ARK_ARC_1_2/temp5[57] ,
         \MC_ARK_ARC_1_2/temp5[56] , \MC_ARK_ARC_1_2/temp5[55] ,
         \MC_ARK_ARC_1_2/temp5[54] , \MC_ARK_ARC_1_2/temp5[52] ,
         \MC_ARK_ARC_1_2/temp5[51] , \MC_ARK_ARC_1_2/temp5[49] ,
         \MC_ARK_ARC_1_2/temp5[48] , \MC_ARK_ARC_1_2/temp5[45] ,
         \MC_ARK_ARC_1_2/temp5[44] , \MC_ARK_ARC_1_2/temp5[40] ,
         \MC_ARK_ARC_1_2/temp5[39] , \MC_ARK_ARC_1_2/temp5[38] ,
         \MC_ARK_ARC_1_2/temp5[37] , \MC_ARK_ARC_1_2/temp5[36] ,
         \MC_ARK_ARC_1_2/temp5[34] , \MC_ARK_ARC_1_2/temp5[30] ,
         \MC_ARK_ARC_1_2/temp5[29] , \MC_ARK_ARC_1_2/temp5[27] ,
         \MC_ARK_ARC_1_2/temp5[25] , \MC_ARK_ARC_1_2/temp5[24] ,
         \MC_ARK_ARC_1_2/temp5[21] , \MC_ARK_ARC_1_2/temp5[20] ,
         \MC_ARK_ARC_1_2/temp5[18] , \MC_ARK_ARC_1_2/temp5[15] ,
         \MC_ARK_ARC_1_2/temp5[14] , \MC_ARK_ARC_1_2/temp5[13] ,
         \MC_ARK_ARC_1_2/temp5[12] , \MC_ARK_ARC_1_2/temp5[10] ,
         \MC_ARK_ARC_1_2/temp5[6] , \MC_ARK_ARC_1_2/temp5[5] ,
         \MC_ARK_ARC_1_2/temp5[4] , \MC_ARK_ARC_1_2/temp5[3] ,
         \MC_ARK_ARC_1_2/temp5[2] , \MC_ARK_ARC_1_2/temp5[0] ,
         \MC_ARK_ARC_1_2/temp4[191] , \MC_ARK_ARC_1_2/temp4[190] ,
         \MC_ARK_ARC_1_2/temp4[189] , \MC_ARK_ARC_1_2/temp4[188] ,
         \MC_ARK_ARC_1_2/temp4[187] , \MC_ARK_ARC_1_2/temp4[186] ,
         \MC_ARK_ARC_1_2/temp4[185] , \MC_ARK_ARC_1_2/temp4[184] ,
         \MC_ARK_ARC_1_2/temp4[183] , \MC_ARK_ARC_1_2/temp4[182] ,
         \MC_ARK_ARC_1_2/temp4[181] , \MC_ARK_ARC_1_2/temp4[180] ,
         \MC_ARK_ARC_1_2/temp4[179] , \MC_ARK_ARC_1_2/temp4[178] ,
         \MC_ARK_ARC_1_2/temp4[177] , \MC_ARK_ARC_1_2/temp4[176] ,
         \MC_ARK_ARC_1_2/temp4[175] , \MC_ARK_ARC_1_2/temp4[174] ,
         \MC_ARK_ARC_1_2/temp4[173] , \MC_ARK_ARC_1_2/temp4[172] ,
         \MC_ARK_ARC_1_2/temp4[171] , \MC_ARK_ARC_1_2/temp4[169] ,
         \MC_ARK_ARC_1_2/temp4[168] , \MC_ARK_ARC_1_2/temp4[166] ,
         \MC_ARK_ARC_1_2/temp4[165] , \MC_ARK_ARC_1_2/temp4[163] ,
         \MC_ARK_ARC_1_2/temp4[162] , \MC_ARK_ARC_1_2/temp4[161] ,
         \MC_ARK_ARC_1_2/temp4[160] , \MC_ARK_ARC_1_2/temp4[159] ,
         \MC_ARK_ARC_1_2/temp4[158] , \MC_ARK_ARC_1_2/temp4[157] ,
         \MC_ARK_ARC_1_2/temp4[156] , \MC_ARK_ARC_1_2/temp4[155] ,
         \MC_ARK_ARC_1_2/temp4[154] , \MC_ARK_ARC_1_2/temp4[153] ,
         \MC_ARK_ARC_1_2/temp4[152] , \MC_ARK_ARC_1_2/temp4[151] ,
         \MC_ARK_ARC_1_2/temp4[150] , \MC_ARK_ARC_1_2/temp4[149] ,
         \MC_ARK_ARC_1_2/temp4[148] , \MC_ARK_ARC_1_2/temp4[147] ,
         \MC_ARK_ARC_1_2/temp4[146] , \MC_ARK_ARC_1_2/temp4[145] ,
         \MC_ARK_ARC_1_2/temp4[144] , \MC_ARK_ARC_1_2/temp4[143] ,
         \MC_ARK_ARC_1_2/temp4[142] , \MC_ARK_ARC_1_2/temp4[141] ,
         \MC_ARK_ARC_1_2/temp4[140] , \MC_ARK_ARC_1_2/temp4[139] ,
         \MC_ARK_ARC_1_2/temp4[138] , \MC_ARK_ARC_1_2/temp4[137] ,
         \MC_ARK_ARC_1_2/temp4[136] , \MC_ARK_ARC_1_2/temp4[135] ,
         \MC_ARK_ARC_1_2/temp4[134] , \MC_ARK_ARC_1_2/temp4[133] ,
         \MC_ARK_ARC_1_2/temp4[132] , \MC_ARK_ARC_1_2/temp4[131] ,
         \MC_ARK_ARC_1_2/temp4[130] , \MC_ARK_ARC_1_2/temp4[129] ,
         \MC_ARK_ARC_1_2/temp4[128] , \MC_ARK_ARC_1_2/temp4[127] ,
         \MC_ARK_ARC_1_2/temp4[126] , \MC_ARK_ARC_1_2/temp4[124] ,
         \MC_ARK_ARC_1_2/temp4[123] , \MC_ARK_ARC_1_2/temp4[121] ,
         \MC_ARK_ARC_1_2/temp4[120] , \MC_ARK_ARC_1_2/temp4[119] ,
         \MC_ARK_ARC_1_2/temp4[118] , \MC_ARK_ARC_1_2/temp4[117] ,
         \MC_ARK_ARC_1_2/temp4[116] , \MC_ARK_ARC_1_2/temp4[115] ,
         \MC_ARK_ARC_1_2/temp4[114] , \MC_ARK_ARC_1_2/temp4[113] ,
         \MC_ARK_ARC_1_2/temp4[112] , \MC_ARK_ARC_1_2/temp4[111] ,
         \MC_ARK_ARC_1_2/temp4[110] , \MC_ARK_ARC_1_2/temp4[109] ,
         \MC_ARK_ARC_1_2/temp4[108] , \MC_ARK_ARC_1_2/temp4[107] ,
         \MC_ARK_ARC_1_2/temp4[106] , \MC_ARK_ARC_1_2/temp4[105] ,
         \MC_ARK_ARC_1_2/temp4[104] , \MC_ARK_ARC_1_2/temp4[103] ,
         \MC_ARK_ARC_1_2/temp4[102] , \MC_ARK_ARC_1_2/temp4[100] ,
         \MC_ARK_ARC_1_2/temp4[99] , \MC_ARK_ARC_1_2/temp4[97] ,
         \MC_ARK_ARC_1_2/temp4[96] , \MC_ARK_ARC_1_2/temp4[95] ,
         \MC_ARK_ARC_1_2/temp4[94] , \MC_ARK_ARC_1_2/temp4[93] ,
         \MC_ARK_ARC_1_2/temp4[92] , \MC_ARK_ARC_1_2/temp4[91] ,
         \MC_ARK_ARC_1_2/temp4[90] , \MC_ARK_ARC_1_2/temp4[89] ,
         \MC_ARK_ARC_1_2/temp4[88] , \MC_ARK_ARC_1_2/temp4[87] ,
         \MC_ARK_ARC_1_2/temp4[86] , \MC_ARK_ARC_1_2/temp4[85] ,
         \MC_ARK_ARC_1_2/temp4[84] , \MC_ARK_ARC_1_2/temp4[83] ,
         \MC_ARK_ARC_1_2/temp4[82] , \MC_ARK_ARC_1_2/temp4[81] ,
         \MC_ARK_ARC_1_2/temp4[80] , \MC_ARK_ARC_1_2/temp4[79] ,
         \MC_ARK_ARC_1_2/temp4[78] , \MC_ARK_ARC_1_2/temp4[77] ,
         \MC_ARK_ARC_1_2/temp4[76] , \MC_ARK_ARC_1_2/temp4[75] ,
         \MC_ARK_ARC_1_2/temp4[74] , \MC_ARK_ARC_1_2/temp4[73] ,
         \MC_ARK_ARC_1_2/temp4[71] , \MC_ARK_ARC_1_2/temp4[70] ,
         \MC_ARK_ARC_1_2/temp4[69] , \MC_ARK_ARC_1_2/temp4[68] ,
         \MC_ARK_ARC_1_2/temp4[67] , \MC_ARK_ARC_1_2/temp4[66] ,
         \MC_ARK_ARC_1_2/temp4[65] , \MC_ARK_ARC_1_2/temp4[64] ,
         \MC_ARK_ARC_1_2/temp4[63] , \MC_ARK_ARC_1_2/temp4[62] ,
         \MC_ARK_ARC_1_2/temp4[61] , \MC_ARK_ARC_1_2/temp4[60] ,
         \MC_ARK_ARC_1_2/temp4[59] , \MC_ARK_ARC_1_2/temp4[58] ,
         \MC_ARK_ARC_1_2/temp4[57] , \MC_ARK_ARC_1_2/temp4[56] ,
         \MC_ARK_ARC_1_2/temp4[55] , \MC_ARK_ARC_1_2/temp4[54] ,
         \MC_ARK_ARC_1_2/temp4[53] , \MC_ARK_ARC_1_2/temp4[51] ,
         \MC_ARK_ARC_1_2/temp4[49] , \MC_ARK_ARC_1_2/temp4[48] ,
         \MC_ARK_ARC_1_2/temp4[47] , \MC_ARK_ARC_1_2/temp4[46] ,
         \MC_ARK_ARC_1_2/temp4[45] , \MC_ARK_ARC_1_2/temp4[44] ,
         \MC_ARK_ARC_1_2/temp4[43] , \MC_ARK_ARC_1_2/temp4[42] ,
         \MC_ARK_ARC_1_2/temp4[41] , \MC_ARK_ARC_1_2/temp4[40] ,
         \MC_ARK_ARC_1_2/temp4[39] , \MC_ARK_ARC_1_2/temp4[37] ,
         \MC_ARK_ARC_1_2/temp4[36] , \MC_ARK_ARC_1_2/temp4[35] ,
         \MC_ARK_ARC_1_2/temp4[34] , \MC_ARK_ARC_1_2/temp4[33] ,
         \MC_ARK_ARC_1_2/temp4[31] , \MC_ARK_ARC_1_2/temp4[30] ,
         \MC_ARK_ARC_1_2/temp4[28] , \MC_ARK_ARC_1_2/temp4[27] ,
         \MC_ARK_ARC_1_2/temp4[26] , \MC_ARK_ARC_1_2/temp4[25] ,
         \MC_ARK_ARC_1_2/temp4[24] , \MC_ARK_ARC_1_2/temp4[23] ,
         \MC_ARK_ARC_1_2/temp4[22] , \MC_ARK_ARC_1_2/temp4[20] ,
         \MC_ARK_ARC_1_2/temp4[19] , \MC_ARK_ARC_1_2/temp4[18] ,
         \MC_ARK_ARC_1_2/temp4[17] , \MC_ARK_ARC_1_2/temp4[16] ,
         \MC_ARK_ARC_1_2/temp4[15] , \MC_ARK_ARC_1_2/temp4[13] ,
         \MC_ARK_ARC_1_2/temp4[12] , \MC_ARK_ARC_1_2/temp4[11] ,
         \MC_ARK_ARC_1_2/temp4[10] , \MC_ARK_ARC_1_2/temp4[9] ,
         \MC_ARK_ARC_1_2/temp4[8] , \MC_ARK_ARC_1_2/temp4[7] ,
         \MC_ARK_ARC_1_2/temp4[6] , \MC_ARK_ARC_1_2/temp4[5] ,
         \MC_ARK_ARC_1_2/temp4[4] , \MC_ARK_ARC_1_2/temp4[3] ,
         \MC_ARK_ARC_1_2/temp4[2] , \MC_ARK_ARC_1_2/temp4[1] ,
         \MC_ARK_ARC_1_2/temp4[0] , \MC_ARK_ARC_1_2/temp3[191] ,
         \MC_ARK_ARC_1_2/temp3[190] , \MC_ARK_ARC_1_2/temp3[189] ,
         \MC_ARK_ARC_1_2/temp3[188] , \MC_ARK_ARC_1_2/temp3[187] ,
         \MC_ARK_ARC_1_2/temp3[186] , \MC_ARK_ARC_1_2/temp3[185] ,
         \MC_ARK_ARC_1_2/temp3[184] , \MC_ARK_ARC_1_2/temp3[183] ,
         \MC_ARK_ARC_1_2/temp3[182] , \MC_ARK_ARC_1_2/temp3[181] ,
         \MC_ARK_ARC_1_2/temp3[180] , \MC_ARK_ARC_1_2/temp3[178] ,
         \MC_ARK_ARC_1_2/temp3[177] , \MC_ARK_ARC_1_2/temp3[176] ,
         \MC_ARK_ARC_1_2/temp3[175] , \MC_ARK_ARC_1_2/temp3[174] ,
         \MC_ARK_ARC_1_2/temp3[173] , \MC_ARK_ARC_1_2/temp3[172] ,
         \MC_ARK_ARC_1_2/temp3[171] , \MC_ARK_ARC_1_2/temp3[169] ,
         \MC_ARK_ARC_1_2/temp3[168] , \MC_ARK_ARC_1_2/temp3[166] ,
         \MC_ARK_ARC_1_2/temp3[163] , \MC_ARK_ARC_1_2/temp3[162] ,
         \MC_ARK_ARC_1_2/temp3[161] , \MC_ARK_ARC_1_2/temp3[160] ,
         \MC_ARK_ARC_1_2/temp3[159] , \MC_ARK_ARC_1_2/temp3[158] ,
         \MC_ARK_ARC_1_2/temp3[156] , \MC_ARK_ARC_1_2/temp3[155] ,
         \MC_ARK_ARC_1_2/temp3[154] , \MC_ARK_ARC_1_2/temp3[153] ,
         \MC_ARK_ARC_1_2/temp3[151] , \MC_ARK_ARC_1_2/temp3[150] ,
         \MC_ARK_ARC_1_2/temp3[148] , \MC_ARK_ARC_1_2/temp3[145] ,
         \MC_ARK_ARC_1_2/temp3[143] , \MC_ARK_ARC_1_2/temp3[142] ,
         \MC_ARK_ARC_1_2/temp3[141] , \MC_ARK_ARC_1_2/temp3[140] ,
         \MC_ARK_ARC_1_2/temp3[139] , \MC_ARK_ARC_1_2/temp3[138] ,
         \MC_ARK_ARC_1_2/temp3[136] , \MC_ARK_ARC_1_2/temp3[135] ,
         \MC_ARK_ARC_1_2/temp3[134] , \MC_ARK_ARC_1_2/temp3[132] ,
         \MC_ARK_ARC_1_2/temp3[130] , \MC_ARK_ARC_1_2/temp3[129] ,
         \MC_ARK_ARC_1_2/temp3[124] , \MC_ARK_ARC_1_2/temp3[120] ,
         \MC_ARK_ARC_1_2/temp3[119] , \MC_ARK_ARC_1_2/temp3[117] ,
         \MC_ARK_ARC_1_2/temp3[115] , \MC_ARK_ARC_1_2/temp3[114] ,
         \MC_ARK_ARC_1_2/temp3[113] , \MC_ARK_ARC_1_2/temp3[111] ,
         \MC_ARK_ARC_1_2/temp3[110] , \MC_ARK_ARC_1_2/temp3[109] ,
         \MC_ARK_ARC_1_2/temp3[108] , \MC_ARK_ARC_1_2/temp3[106] ,
         \MC_ARK_ARC_1_2/temp3[105] , \MC_ARK_ARC_1_2/temp3[103] ,
         \MC_ARK_ARC_1_2/temp3[102] , \MC_ARK_ARC_1_2/temp3[100] ,
         \MC_ARK_ARC_1_2/temp3[97] , \MC_ARK_ARC_1_2/temp3[96] ,
         \MC_ARK_ARC_1_2/temp3[94] , \MC_ARK_ARC_1_2/temp3[93] ,
         \MC_ARK_ARC_1_2/temp3[91] , \MC_ARK_ARC_1_2/temp3[90] ,
         \MC_ARK_ARC_1_2/temp3[88] , \MC_ARK_ARC_1_2/temp3[86] ,
         \MC_ARK_ARC_1_2/temp3[85] , \MC_ARK_ARC_1_2/temp3[84] ,
         \MC_ARK_ARC_1_2/temp3[82] , \MC_ARK_ARC_1_2/temp3[81] ,
         \MC_ARK_ARC_1_2/temp3[80] , \MC_ARK_ARC_1_2/temp3[79] ,
         \MC_ARK_ARC_1_2/temp3[78] , \MC_ARK_ARC_1_2/temp3[77] ,
         \MC_ARK_ARC_1_2/temp3[76] , \MC_ARK_ARC_1_2/temp3[75] ,
         \MC_ARK_ARC_1_2/temp3[74] , \MC_ARK_ARC_1_2/temp3[71] ,
         \MC_ARK_ARC_1_2/temp3[70] , \MC_ARK_ARC_1_2/temp3[69] ,
         \MC_ARK_ARC_1_2/temp3[68] , \MC_ARK_ARC_1_2/temp3[67] ,
         \MC_ARK_ARC_1_2/temp3[66] , \MC_ARK_ARC_1_2/temp3[65] ,
         \MC_ARK_ARC_1_2/temp3[62] , \MC_ARK_ARC_1_2/temp3[61] ,
         \MC_ARK_ARC_1_2/temp3[60] , \MC_ARK_ARC_1_2/temp3[59] ,
         \MC_ARK_ARC_1_2/temp3[57] , \MC_ARK_ARC_1_2/temp3[54] ,
         \MC_ARK_ARC_1_2/temp3[53] , \MC_ARK_ARC_1_2/temp3[51] ,
         \MC_ARK_ARC_1_2/temp3[49] , \MC_ARK_ARC_1_2/temp3[48] ,
         \MC_ARK_ARC_1_2/temp3[46] , \MC_ARK_ARC_1_2/temp3[43] ,
         \MC_ARK_ARC_1_2/temp3[42] , \MC_ARK_ARC_1_2/temp3[41] ,
         \MC_ARK_ARC_1_2/temp3[40] , \MC_ARK_ARC_1_2/temp3[39] ,
         \MC_ARK_ARC_1_2/temp3[36] , \MC_ARK_ARC_1_2/temp3[34] ,
         \MC_ARK_ARC_1_2/temp3[33] , \MC_ARK_ARC_1_2/temp3[31] ,
         \MC_ARK_ARC_1_2/temp3[30] , \MC_ARK_ARC_1_2/temp3[28] ,
         \MC_ARK_ARC_1_2/temp3[27] , \MC_ARK_ARC_1_2/temp3[25] ,
         \MC_ARK_ARC_1_2/temp3[24] , \MC_ARK_ARC_1_2/temp3[23] ,
         \MC_ARK_ARC_1_2/temp3[22] , \MC_ARK_ARC_1_2/temp3[18] ,
         \MC_ARK_ARC_1_2/temp3[17] , \MC_ARK_ARC_1_2/temp3[16] ,
         \MC_ARK_ARC_1_2/temp3[13] , \MC_ARK_ARC_1_2/temp3[11] ,
         \MC_ARK_ARC_1_2/temp3[10] , \MC_ARK_ARC_1_2/temp3[8] ,
         \MC_ARK_ARC_1_2/temp3[7] , \MC_ARK_ARC_1_2/temp3[6] ,
         \MC_ARK_ARC_1_2/temp3[5] , \MC_ARK_ARC_1_2/temp3[4] ,
         \MC_ARK_ARC_1_2/temp3[3] , \MC_ARK_ARC_1_2/temp3[2] ,
         \MC_ARK_ARC_1_2/temp3[1] , \MC_ARK_ARC_1_2/temp3[0] ,
         \MC_ARK_ARC_1_2/temp2[191] , \MC_ARK_ARC_1_2/temp2[190] ,
         \MC_ARK_ARC_1_2/temp2[186] , \MC_ARK_ARC_1_2/temp2[184] ,
         \MC_ARK_ARC_1_2/temp2[183] , \MC_ARK_ARC_1_2/temp2[181] ,
         \MC_ARK_ARC_1_2/temp2[180] , \MC_ARK_ARC_1_2/temp2[179] ,
         \MC_ARK_ARC_1_2/temp2[178] , \MC_ARK_ARC_1_2/temp2[177] ,
         \MC_ARK_ARC_1_2/temp2[176] , \MC_ARK_ARC_1_2/temp2[174] ,
         \MC_ARK_ARC_1_2/temp2[173] , \MC_ARK_ARC_1_2/temp2[172] ,
         \MC_ARK_ARC_1_2/temp2[170] , \MC_ARK_ARC_1_2/temp2[169] ,
         \MC_ARK_ARC_1_2/temp2[167] , \MC_ARK_ARC_1_2/temp2[165] ,
         \MC_ARK_ARC_1_2/temp2[164] , \MC_ARK_ARC_1_2/temp2[162] ,
         \MC_ARK_ARC_1_2/temp2[159] , \MC_ARK_ARC_1_2/temp2[157] ,
         \MC_ARK_ARC_1_2/temp2[154] , \MC_ARK_ARC_1_2/temp2[153] ,
         \MC_ARK_ARC_1_2/temp2[151] , \MC_ARK_ARC_1_2/temp2[150] ,
         \MC_ARK_ARC_1_2/temp2[148] , \MC_ARK_ARC_1_2/temp2[147] ,
         \MC_ARK_ARC_1_2/temp2[145] , \MC_ARK_ARC_1_2/temp2[144] ,
         \MC_ARK_ARC_1_2/temp2[142] , \MC_ARK_ARC_1_2/temp2[139] ,
         \MC_ARK_ARC_1_2/temp2[138] , \MC_ARK_ARC_1_2/temp2[136] ,
         \MC_ARK_ARC_1_2/temp2[133] , \MC_ARK_ARC_1_2/temp2[130] ,
         \MC_ARK_ARC_1_2/temp2[128] , \MC_ARK_ARC_1_2/temp2[126] ,
         \MC_ARK_ARC_1_2/temp2[122] , \MC_ARK_ARC_1_2/temp2[121] ,
         \MC_ARK_ARC_1_2/temp2[118] , \MC_ARK_ARC_1_2/temp2[117] ,
         \MC_ARK_ARC_1_2/temp2[115] , \MC_ARK_ARC_1_2/temp2[114] ,
         \MC_ARK_ARC_1_2/temp2[112] , \MC_ARK_ARC_1_2/temp2[108] ,
         \MC_ARK_ARC_1_2/temp2[106] , \MC_ARK_ARC_1_2/temp2[105] ,
         \MC_ARK_ARC_1_2/temp2[104] , \MC_ARK_ARC_1_2/temp2[103] ,
         \MC_ARK_ARC_1_2/temp2[102] , \MC_ARK_ARC_1_2/temp2[100] ,
         \MC_ARK_ARC_1_2/temp2[97] , \MC_ARK_ARC_1_2/temp2[96] ,
         \MC_ARK_ARC_1_2/temp2[95] , \MC_ARK_ARC_1_2/temp2[94] ,
         \MC_ARK_ARC_1_2/temp2[93] , \MC_ARK_ARC_1_2/temp2[92] ,
         \MC_ARK_ARC_1_2/temp2[88] , \MC_ARK_ARC_1_2/temp2[86] ,
         \MC_ARK_ARC_1_2/temp2[85] , \MC_ARK_ARC_1_2/temp2[84] ,
         \MC_ARK_ARC_1_2/temp2[83] , \MC_ARK_ARC_1_2/temp2[82] ,
         \MC_ARK_ARC_1_2/temp2[80] , \MC_ARK_ARC_1_2/temp2[79] ,
         \MC_ARK_ARC_1_2/temp2[78] , \MC_ARK_ARC_1_2/temp2[76] ,
         \MC_ARK_ARC_1_2/temp2[75] , \MC_ARK_ARC_1_2/temp2[74] ,
         \MC_ARK_ARC_1_2/temp2[73] , \MC_ARK_ARC_1_2/temp2[72] ,
         \MC_ARK_ARC_1_2/temp2[70] , \MC_ARK_ARC_1_2/temp2[69] ,
         \MC_ARK_ARC_1_2/temp2[68] , \MC_ARK_ARC_1_2/temp2[67] ,
         \MC_ARK_ARC_1_2/temp2[66] , \MC_ARK_ARC_1_2/temp2[61] ,
         \MC_ARK_ARC_1_2/temp2[60] , \MC_ARK_ARC_1_2/temp2[55] ,
         \MC_ARK_ARC_1_2/temp2[54] , \MC_ARK_ARC_1_2/temp2[52] ,
         \MC_ARK_ARC_1_2/temp2[49] , \MC_ARK_ARC_1_2/temp2[48] ,
         \MC_ARK_ARC_1_2/temp2[45] , \MC_ARK_ARC_1_2/temp2[44] ,
         \MC_ARK_ARC_1_2/temp2[43] , \MC_ARK_ARC_1_2/temp2[41] ,
         \MC_ARK_ARC_1_2/temp2[40] , \MC_ARK_ARC_1_2/temp2[38] ,
         \MC_ARK_ARC_1_2/temp2[37] , \MC_ARK_ARC_1_2/temp2[36] ,
         \MC_ARK_ARC_1_2/temp2[34] , \MC_ARK_ARC_1_2/temp2[33] ,
         \MC_ARK_ARC_1_2/temp2[31] , \MC_ARK_ARC_1_2/temp2[29] ,
         \MC_ARK_ARC_1_2/temp2[28] , \MC_ARK_ARC_1_2/temp2[27] ,
         \MC_ARK_ARC_1_2/temp2[26] , \MC_ARK_ARC_1_2/temp2[25] ,
         \MC_ARK_ARC_1_2/temp2[24] , \MC_ARK_ARC_1_2/temp2[22] ,
         \MC_ARK_ARC_1_2/temp2[19] , \MC_ARK_ARC_1_2/temp2[18] ,
         \MC_ARK_ARC_1_2/temp2[13] , \MC_ARK_ARC_1_2/temp2[11] ,
         \MC_ARK_ARC_1_2/temp2[8] , \MC_ARK_ARC_1_2/temp2[7] ,
         \MC_ARK_ARC_1_2/temp2[1] , \MC_ARK_ARC_1_2/temp2[0] ,
         \MC_ARK_ARC_1_2/temp1[190] , \MC_ARK_ARC_1_2/temp1[187] ,
         \MC_ARK_ARC_1_2/temp1[186] , \MC_ARK_ARC_1_2/temp1[183] ,
         \MC_ARK_ARC_1_2/temp1[181] , \MC_ARK_ARC_1_2/temp1[180] ,
         \MC_ARK_ARC_1_2/temp1[179] , \MC_ARK_ARC_1_2/temp1[178] ,
         \MC_ARK_ARC_1_2/temp1[177] , \MC_ARK_ARC_1_2/temp1[176] ,
         \MC_ARK_ARC_1_2/temp1[175] , \MC_ARK_ARC_1_2/temp1[174] ,
         \MC_ARK_ARC_1_2/temp1[172] , \MC_ARK_ARC_1_2/temp1[171] ,
         \MC_ARK_ARC_1_2/temp1[169] , \MC_ARK_ARC_1_2/temp1[168] ,
         \MC_ARK_ARC_1_2/temp1[167] , \MC_ARK_ARC_1_2/temp1[165] ,
         \MC_ARK_ARC_1_2/temp1[164] , \MC_ARK_ARC_1_2/temp1[163] ,
         \MC_ARK_ARC_1_2/temp1[162] , \MC_ARK_ARC_1_2/temp1[160] ,
         \MC_ARK_ARC_1_2/temp1[159] , \MC_ARK_ARC_1_2/temp1[157] ,
         \MC_ARK_ARC_1_2/temp1[156] , \MC_ARK_ARC_1_2/temp1[154] ,
         \MC_ARK_ARC_1_2/temp1[153] , \MC_ARK_ARC_1_2/temp1[152] ,
         \MC_ARK_ARC_1_2/temp1[151] , \MC_ARK_ARC_1_2/temp1[150] ,
         \MC_ARK_ARC_1_2/temp1[148] , \MC_ARK_ARC_1_2/temp1[147] ,
         \MC_ARK_ARC_1_2/temp1[145] , \MC_ARK_ARC_1_2/temp1[142] ,
         \MC_ARK_ARC_1_2/temp1[140] , \MC_ARK_ARC_1_2/temp1[139] ,
         \MC_ARK_ARC_1_2/temp1[138] , \MC_ARK_ARC_1_2/temp1[137] ,
         \MC_ARK_ARC_1_2/temp1[136] , \MC_ARK_ARC_1_2/temp1[134] ,
         \MC_ARK_ARC_1_2/temp1[133] , \MC_ARK_ARC_1_2/temp1[130] ,
         \MC_ARK_ARC_1_2/temp1[129] , \MC_ARK_ARC_1_2/temp1[128] ,
         \MC_ARK_ARC_1_2/temp1[127] , \MC_ARK_ARC_1_2/temp1[126] ,
         \MC_ARK_ARC_1_2/temp1[124] , \MC_ARK_ARC_1_2/temp1[121] ,
         \MC_ARK_ARC_1_2/temp1[119] , \MC_ARK_ARC_1_2/temp1[118] ,
         \MC_ARK_ARC_1_2/temp1[115] , \MC_ARK_ARC_1_2/temp1[114] ,
         \MC_ARK_ARC_1_2/temp1[113] , \MC_ARK_ARC_1_2/temp1[112] ,
         \MC_ARK_ARC_1_2/temp1[111] , \MC_ARK_ARC_1_2/temp1[108] ,
         \MC_ARK_ARC_1_2/temp1[106] , \MC_ARK_ARC_1_2/temp1[105] ,
         \MC_ARK_ARC_1_2/temp1[103] , \MC_ARK_ARC_1_2/temp1[102] ,
         \MC_ARK_ARC_1_2/temp1[101] , \MC_ARK_ARC_1_2/temp1[96] ,
         \MC_ARK_ARC_1_2/temp1[95] , \MC_ARK_ARC_1_2/temp1[94] ,
         \MC_ARK_ARC_1_2/temp1[91] , \MC_ARK_ARC_1_2/temp1[88] ,
         \MC_ARK_ARC_1_2/temp1[84] , \MC_ARK_ARC_1_2/temp1[82] ,
         \MC_ARK_ARC_1_2/temp1[81] , \MC_ARK_ARC_1_2/temp1[80] ,
         \MC_ARK_ARC_1_2/temp1[79] , \MC_ARK_ARC_1_2/temp1[78] ,
         \MC_ARK_ARC_1_2/temp1[77] , \MC_ARK_ARC_1_2/temp1[73] ,
         \MC_ARK_ARC_1_2/temp1[72] , \MC_ARK_ARC_1_2/temp1[71] ,
         \MC_ARK_ARC_1_2/temp1[70] , \MC_ARK_ARC_1_2/temp1[67] ,
         \MC_ARK_ARC_1_2/temp1[66] , \MC_ARK_ARC_1_2/temp1[63] ,
         \MC_ARK_ARC_1_2/temp1[61] , \MC_ARK_ARC_1_2/temp1[60] ,
         \MC_ARK_ARC_1_2/temp1[59] , \MC_ARK_ARC_1_2/temp1[58] ,
         \MC_ARK_ARC_1_2/temp1[57] , \MC_ARK_ARC_1_2/temp1[55] ,
         \MC_ARK_ARC_1_2/temp1[54] , \MC_ARK_ARC_1_2/temp1[53] ,
         \MC_ARK_ARC_1_2/temp1[52] , \MC_ARK_ARC_1_2/temp1[51] ,
         \MC_ARK_ARC_1_2/temp1[49] , \MC_ARK_ARC_1_2/temp1[48] ,
         \MC_ARK_ARC_1_2/temp1[46] , \MC_ARK_ARC_1_2/temp1[42] ,
         \MC_ARK_ARC_1_2/temp1[41] , \MC_ARK_ARC_1_2/temp1[40] ,
         \MC_ARK_ARC_1_2/temp1[39] , \MC_ARK_ARC_1_2/temp1[38] ,
         \MC_ARK_ARC_1_2/temp1[37] , \MC_ARK_ARC_1_2/temp1[36] ,
         \MC_ARK_ARC_1_2/temp1[34] , \MC_ARK_ARC_1_2/temp1[32] ,
         \MC_ARK_ARC_1_2/temp1[30] , \MC_ARK_ARC_1_2/temp1[28] ,
         \MC_ARK_ARC_1_2/temp1[27] , \MC_ARK_ARC_1_2/temp1[24] ,
         \MC_ARK_ARC_1_2/temp1[22] , \MC_ARK_ARC_1_2/temp1[20] ,
         \MC_ARK_ARC_1_2/temp1[19] , \MC_ARK_ARC_1_2/temp1[18] ,
         \MC_ARK_ARC_1_2/temp1[17] , \MC_ARK_ARC_1_2/temp1[16] ,
         \MC_ARK_ARC_1_2/temp1[15] , \MC_ARK_ARC_1_2/temp1[14] ,
         \MC_ARK_ARC_1_2/temp1[13] , \MC_ARK_ARC_1_2/temp1[11] ,
         \MC_ARK_ARC_1_2/temp1[10] , \MC_ARK_ARC_1_2/temp1[8] ,
         \MC_ARK_ARC_1_2/temp1[7] , \MC_ARK_ARC_1_2/temp1[4] ,
         \MC_ARK_ARC_1_2/temp1[3] , \MC_ARK_ARC_1_2/temp1[1] ,
         \MC_ARK_ARC_1_2/temp1[0] , \MC_ARK_ARC_1_2/buf_keyinput[54] ,
         \MC_ARK_ARC_1_2/buf_datainput[186] ,
         \MC_ARK_ARC_1_2/buf_datainput[185] ,
         \MC_ARK_ARC_1_2/buf_datainput[183] ,
         \MC_ARK_ARC_1_2/buf_datainput[182] ,
         \MC_ARK_ARC_1_2/buf_datainput[177] ,
         \MC_ARK_ARC_1_2/buf_datainput[175] ,
         \MC_ARK_ARC_1_2/buf_datainput[162] ,
         \MC_ARK_ARC_1_2/buf_datainput[158] ,
         \MC_ARK_ARC_1_2/buf_datainput[156] ,
         \MC_ARK_ARC_1_2/buf_datainput[153] ,
         \MC_ARK_ARC_1_2/buf_datainput[151] ,
         \MC_ARK_ARC_1_2/buf_datainput[149] ,
         \MC_ARK_ARC_1_2/buf_datainput[148] ,
         \MC_ARK_ARC_1_2/buf_datainput[146] ,
         \MC_ARK_ARC_1_2/buf_datainput[141] ,
         \MC_ARK_ARC_1_2/buf_datainput[136] ,
         \MC_ARK_ARC_1_2/buf_datainput[133] ,
         \MC_ARK_ARC_1_2/buf_datainput[132] ,
         \MC_ARK_ARC_1_2/buf_datainput[131] ,
         \MC_ARK_ARC_1_2/buf_datainput[129] ,
         \MC_ARK_ARC_1_2/buf_datainput[128] ,
         \MC_ARK_ARC_1_2/buf_datainput[127] ,
         \MC_ARK_ARC_1_2/buf_datainput[125] ,
         \MC_ARK_ARC_1_2/buf_datainput[124] ,
         \MC_ARK_ARC_1_2/buf_datainput[122] ,
         \MC_ARK_ARC_1_2/buf_datainput[117] ,
         \MC_ARK_ARC_1_2/buf_datainput[116] ,
         \MC_ARK_ARC_1_2/buf_datainput[115] ,
         \MC_ARK_ARC_1_2/buf_datainput[106] ,
         \MC_ARK_ARC_1_2/buf_datainput[105] ,
         \MC_ARK_ARC_1_2/buf_datainput[99] ,
         \MC_ARK_ARC_1_2/buf_datainput[97] ,
         \MC_ARK_ARC_1_2/buf_datainput[95] ,
         \MC_ARK_ARC_1_2/buf_datainput[92] ,
         \MC_ARK_ARC_1_2/buf_datainput[86] ,
         \MC_ARK_ARC_1_2/buf_datainput[83] ,
         \MC_ARK_ARC_1_2/buf_datainput[82] ,
         \MC_ARK_ARC_1_2/buf_datainput[81] ,
         \MC_ARK_ARC_1_2/buf_datainput[78] ,
         \MC_ARK_ARC_1_2/buf_datainput[76] ,
         \MC_ARK_ARC_1_2/buf_datainput[74] ,
         \MC_ARK_ARC_1_2/buf_datainput[70] ,
         \MC_ARK_ARC_1_2/buf_datainput[68] ,
         \MC_ARK_ARC_1_2/buf_datainput[65] ,
         \MC_ARK_ARC_1_2/buf_datainput[61] ,
         \MC_ARK_ARC_1_2/buf_datainput[59] ,
         \MC_ARK_ARC_1_2/buf_datainput[58] ,
         \MC_ARK_ARC_1_2/buf_datainput[56] ,
         \MC_ARK_ARC_1_2/buf_datainput[53] ,
         \MC_ARK_ARC_1_2/buf_datainput[50] ,
         \MC_ARK_ARC_1_2/buf_datainput[49] ,
         \MC_ARK_ARC_1_2/buf_datainput[47] ,
         \MC_ARK_ARC_1_2/buf_datainput[45] ,
         \MC_ARK_ARC_1_2/buf_datainput[43] ,
         \MC_ARK_ARC_1_2/buf_datainput[39] ,
         \MC_ARK_ARC_1_2/buf_datainput[38] ,
         \MC_ARK_ARC_1_2/buf_datainput[36] ,
         \MC_ARK_ARC_1_2/buf_datainput[34] ,
         \MC_ARK_ARC_1_2/buf_datainput[30] ,
         \MC_ARK_ARC_1_2/buf_datainput[29] ,
         \MC_ARK_ARC_1_2/buf_datainput[27] , \MC_ARK_ARC_1_2/buf_datainput[7] ,
         \MC_ARK_ARC_1_2/buf_datainput[6] , \MC_ARK_ARC_1_2/buf_datainput[4] ,
         \MC_ARK_ARC_1_2/buf_datainput[2] , \MC_ARK_ARC_1_2/buf_datainput[0] ,
         \MC_ARK_ARC_1_3/buf_output[191] , \MC_ARK_ARC_1_3/buf_output[190] ,
         \MC_ARK_ARC_1_3/buf_output[189] , \MC_ARK_ARC_1_3/buf_output[188] ,
         \MC_ARK_ARC_1_3/buf_output[187] , \MC_ARK_ARC_1_3/buf_output[186] ,
         \MC_ARK_ARC_1_3/buf_output[185] , \MC_ARK_ARC_1_3/buf_output[184] ,
         \MC_ARK_ARC_1_3/buf_output[183] , \MC_ARK_ARC_1_3/buf_output[182] ,
         \MC_ARK_ARC_1_3/buf_output[181] , \MC_ARK_ARC_1_3/buf_output[180] ,
         \MC_ARK_ARC_1_3/buf_output[178] , \MC_ARK_ARC_1_3/buf_output[177] ,
         \MC_ARK_ARC_1_3/buf_output[176] , \MC_ARK_ARC_1_3/buf_output[175] ,
         \MC_ARK_ARC_1_3/buf_output[174] , \MC_ARK_ARC_1_3/buf_output[173] ,
         \MC_ARK_ARC_1_3/buf_output[172] , \MC_ARK_ARC_1_3/buf_output[171] ,
         \MC_ARK_ARC_1_3/buf_output[170] , \MC_ARK_ARC_1_3/buf_output[169] ,
         \MC_ARK_ARC_1_3/buf_output[168] , \MC_ARK_ARC_1_3/buf_output[167] ,
         \MC_ARK_ARC_1_3/buf_output[166] , \MC_ARK_ARC_1_3/buf_output[165] ,
         \MC_ARK_ARC_1_3/buf_output[164] , \MC_ARK_ARC_1_3/buf_output[163] ,
         \MC_ARK_ARC_1_3/buf_output[162] , \MC_ARK_ARC_1_3/buf_output[161] ,
         \MC_ARK_ARC_1_3/buf_output[160] , \MC_ARK_ARC_1_3/buf_output[159] ,
         \MC_ARK_ARC_1_3/buf_output[158] , \MC_ARK_ARC_1_3/buf_output[157] ,
         \MC_ARK_ARC_1_3/buf_output[156] , \MC_ARK_ARC_1_3/buf_output[155] ,
         \MC_ARK_ARC_1_3/buf_output[154] , \MC_ARK_ARC_1_3/buf_output[153] ,
         \MC_ARK_ARC_1_3/buf_output[152] , \MC_ARK_ARC_1_3/buf_output[151] ,
         \MC_ARK_ARC_1_3/buf_output[150] , \MC_ARK_ARC_1_3/buf_output[149] ,
         \MC_ARK_ARC_1_3/buf_output[148] , \MC_ARK_ARC_1_3/buf_output[147] ,
         \MC_ARK_ARC_1_3/buf_output[146] , \MC_ARK_ARC_1_3/buf_output[145] ,
         \MC_ARK_ARC_1_3/buf_output[144] , \MC_ARK_ARC_1_3/buf_output[142] ,
         \MC_ARK_ARC_1_3/buf_output[141] , \MC_ARK_ARC_1_3/buf_output[140] ,
         \MC_ARK_ARC_1_3/buf_output[139] , \MC_ARK_ARC_1_3/buf_output[138] ,
         \MC_ARK_ARC_1_3/buf_output[137] , \MC_ARK_ARC_1_3/buf_output[136] ,
         \MC_ARK_ARC_1_3/buf_output[135] , \MC_ARK_ARC_1_3/buf_output[134] ,
         \MC_ARK_ARC_1_3/buf_output[133] , \MC_ARK_ARC_1_3/buf_output[132] ,
         \MC_ARK_ARC_1_3/buf_output[130] , \MC_ARK_ARC_1_3/buf_output[129] ,
         \MC_ARK_ARC_1_3/buf_output[128] , \MC_ARK_ARC_1_3/buf_output[127] ,
         \MC_ARK_ARC_1_3/buf_output[126] , \MC_ARK_ARC_1_3/buf_output[124] ,
         \MC_ARK_ARC_1_3/buf_output[123] , \MC_ARK_ARC_1_3/buf_output[122] ,
         \MC_ARK_ARC_1_3/buf_output[121] , \MC_ARK_ARC_1_3/buf_output[120] ,
         \MC_ARK_ARC_1_3/buf_output[119] , \MC_ARK_ARC_1_3/buf_output[118] ,
         \MC_ARK_ARC_1_3/buf_output[117] , \MC_ARK_ARC_1_3/buf_output[116] ,
         \MC_ARK_ARC_1_3/buf_output[115] , \MC_ARK_ARC_1_3/buf_output[114] ,
         \MC_ARK_ARC_1_3/buf_output[113] , \MC_ARK_ARC_1_3/buf_output[112] ,
         \MC_ARK_ARC_1_3/buf_output[111] , \MC_ARK_ARC_1_3/buf_output[110] ,
         \MC_ARK_ARC_1_3/buf_output[109] , \MC_ARK_ARC_1_3/buf_output[108] ,
         \MC_ARK_ARC_1_3/buf_output[107] , \MC_ARK_ARC_1_3/buf_output[106] ,
         \MC_ARK_ARC_1_3/buf_output[105] , \MC_ARK_ARC_1_3/buf_output[104] ,
         \MC_ARK_ARC_1_3/buf_output[103] , \MC_ARK_ARC_1_3/buf_output[102] ,
         \MC_ARK_ARC_1_3/buf_output[101] , \MC_ARK_ARC_1_3/buf_output[100] ,
         \MC_ARK_ARC_1_3/buf_output[99] , \MC_ARK_ARC_1_3/buf_output[98] ,
         \MC_ARK_ARC_1_3/buf_output[97] , \MC_ARK_ARC_1_3/buf_output[96] ,
         \MC_ARK_ARC_1_3/buf_output[95] , \MC_ARK_ARC_1_3/buf_output[94] ,
         \MC_ARK_ARC_1_3/buf_output[93] , \MC_ARK_ARC_1_3/buf_output[92] ,
         \MC_ARK_ARC_1_3/buf_output[91] , \MC_ARK_ARC_1_3/buf_output[90] ,
         \MC_ARK_ARC_1_3/buf_output[88] , \MC_ARK_ARC_1_3/buf_output[86] ,
         \MC_ARK_ARC_1_3/buf_output[85] , \MC_ARK_ARC_1_3/buf_output[84] ,
         \MC_ARK_ARC_1_3/buf_output[83] , \MC_ARK_ARC_1_3/buf_output[82] ,
         \MC_ARK_ARC_1_3/buf_output[81] , \MC_ARK_ARC_1_3/buf_output[80] ,
         \MC_ARK_ARC_1_3/buf_output[79] , \MC_ARK_ARC_1_3/buf_output[78] ,
         \MC_ARK_ARC_1_3/buf_output[76] , \MC_ARK_ARC_1_3/buf_output[75] ,
         \MC_ARK_ARC_1_3/buf_output[74] , \MC_ARK_ARC_1_3/buf_output[73] ,
         \MC_ARK_ARC_1_3/buf_output[72] , \MC_ARK_ARC_1_3/buf_output[71] ,
         \MC_ARK_ARC_1_3/buf_output[70] , \MC_ARK_ARC_1_3/buf_output[69] ,
         \MC_ARK_ARC_1_3/buf_output[68] , \MC_ARK_ARC_1_3/buf_output[67] ,
         \MC_ARK_ARC_1_3/buf_output[66] , \MC_ARK_ARC_1_3/buf_output[65] ,
         \MC_ARK_ARC_1_3/buf_output[64] , \MC_ARK_ARC_1_3/buf_output[63] ,
         \MC_ARK_ARC_1_3/buf_output[62] , \MC_ARK_ARC_1_3/buf_output[61] ,
         \MC_ARK_ARC_1_3/buf_output[60] , \MC_ARK_ARC_1_3/buf_output[58] ,
         \MC_ARK_ARC_1_3/buf_output[57] , \MC_ARK_ARC_1_3/buf_output[56] ,
         \MC_ARK_ARC_1_3/buf_output[55] , \MC_ARK_ARC_1_3/buf_output[54] ,
         \MC_ARK_ARC_1_3/buf_output[52] , \MC_ARK_ARC_1_3/buf_output[51] ,
         \MC_ARK_ARC_1_3/buf_output[49] , \MC_ARK_ARC_1_3/buf_output[48] ,
         \MC_ARK_ARC_1_3/buf_output[47] , \MC_ARK_ARC_1_3/buf_output[46] ,
         \MC_ARK_ARC_1_3/buf_output[45] , \MC_ARK_ARC_1_3/buf_output[44] ,
         \MC_ARK_ARC_1_3/buf_output[43] , \MC_ARK_ARC_1_3/buf_output[42] ,
         \MC_ARK_ARC_1_3/buf_output[40] , \MC_ARK_ARC_1_3/buf_output[39] ,
         \MC_ARK_ARC_1_3/buf_output[38] , \MC_ARK_ARC_1_3/buf_output[37] ,
         \MC_ARK_ARC_1_3/buf_output[36] , \MC_ARK_ARC_1_3/buf_output[35] ,
         \MC_ARK_ARC_1_3/buf_output[34] , \MC_ARK_ARC_1_3/buf_output[33] ,
         \MC_ARK_ARC_1_3/buf_output[32] , \MC_ARK_ARC_1_3/buf_output[31] ,
         \MC_ARK_ARC_1_3/buf_output[30] , \MC_ARK_ARC_1_3/buf_output[28] ,
         \MC_ARK_ARC_1_3/buf_output[27] , \MC_ARK_ARC_1_3/buf_output[26] ,
         \MC_ARK_ARC_1_3/buf_output[25] , \MC_ARK_ARC_1_3/buf_output[24] ,
         \MC_ARK_ARC_1_3/buf_output[23] , \MC_ARK_ARC_1_3/buf_output[22] ,
         \MC_ARK_ARC_1_3/buf_output[21] , \MC_ARK_ARC_1_3/buf_output[20] ,
         \MC_ARK_ARC_1_3/buf_output[19] , \MC_ARK_ARC_1_3/buf_output[18] ,
         \MC_ARK_ARC_1_3/buf_output[17] , \MC_ARK_ARC_1_3/buf_output[16] ,
         \MC_ARK_ARC_1_3/buf_output[15] , \MC_ARK_ARC_1_3/buf_output[14] ,
         \MC_ARK_ARC_1_3/buf_output[13] , \MC_ARK_ARC_1_3/buf_output[12] ,
         \MC_ARK_ARC_1_3/buf_output[10] , \MC_ARK_ARC_1_3/buf_output[9] ,
         \MC_ARK_ARC_1_3/buf_output[8] , \MC_ARK_ARC_1_3/buf_output[7] ,
         \MC_ARK_ARC_1_3/buf_output[6] , \MC_ARK_ARC_1_3/buf_output[4] ,
         \MC_ARK_ARC_1_3/buf_output[3] , \MC_ARK_ARC_1_3/buf_output[2] ,
         \MC_ARK_ARC_1_3/buf_output[1] , \MC_ARK_ARC_1_3/buf_output[0] ,
         \MC_ARK_ARC_1_3/temp6[191] , \MC_ARK_ARC_1_3/temp6[190] ,
         \MC_ARK_ARC_1_3/temp6[187] , \MC_ARK_ARC_1_3/temp6[180] ,
         \MC_ARK_ARC_1_3/temp6[177] , \MC_ARK_ARC_1_3/temp6[176] ,
         \MC_ARK_ARC_1_3/temp6[168] , \MC_ARK_ARC_1_3/temp6[167] ,
         \MC_ARK_ARC_1_3/temp6[166] , \MC_ARK_ARC_1_3/temp6[165] ,
         \MC_ARK_ARC_1_3/temp6[160] , \MC_ARK_ARC_1_3/temp6[157] ,
         \MC_ARK_ARC_1_3/temp6[151] , \MC_ARK_ARC_1_3/temp6[150] ,
         \MC_ARK_ARC_1_3/temp6[149] , \MC_ARK_ARC_1_3/temp6[148] ,
         \MC_ARK_ARC_1_3/temp6[147] , \MC_ARK_ARC_1_3/temp6[145] ,
         \MC_ARK_ARC_1_3/temp6[144] , \MC_ARK_ARC_1_3/temp6[143] ,
         \MC_ARK_ARC_1_3/temp6[142] , \MC_ARK_ARC_1_3/temp6[139] ,
         \MC_ARK_ARC_1_3/temp6[138] , \MC_ARK_ARC_1_3/temp6[135] ,
         \MC_ARK_ARC_1_3/temp6[134] , \MC_ARK_ARC_1_3/temp6[133] ,
         \MC_ARK_ARC_1_3/temp6[132] , \MC_ARK_ARC_1_3/temp6[131] ,
         \MC_ARK_ARC_1_3/temp6[130] , \MC_ARK_ARC_1_3/temp6[128] ,
         \MC_ARK_ARC_1_3/temp6[126] , \MC_ARK_ARC_1_3/temp6[125] ,
         \MC_ARK_ARC_1_3/temp6[123] , \MC_ARK_ARC_1_3/temp6[121] ,
         \MC_ARK_ARC_1_3/temp6[120] , \MC_ARK_ARC_1_3/temp6[119] ,
         \MC_ARK_ARC_1_3/temp6[118] , \MC_ARK_ARC_1_3/temp6[116] ,
         \MC_ARK_ARC_1_3/temp6[113] , \MC_ARK_ARC_1_3/temp6[111] ,
         \MC_ARK_ARC_1_3/temp6[108] , \MC_ARK_ARC_1_3/temp6[106] ,
         \MC_ARK_ARC_1_3/temp6[104] , \MC_ARK_ARC_1_3/temp6[103] ,
         \MC_ARK_ARC_1_3/temp6[102] , \MC_ARK_ARC_1_3/temp6[101] ,
         \MC_ARK_ARC_1_3/temp6[100] , \MC_ARK_ARC_1_3/temp6[99] ,
         \MC_ARK_ARC_1_3/temp6[98] , \MC_ARK_ARC_1_3/temp6[96] ,
         \MC_ARK_ARC_1_3/temp6[91] , \MC_ARK_ARC_1_3/temp6[88] ,
         \MC_ARK_ARC_1_3/temp6[86] , \MC_ARK_ARC_1_3/temp6[81] ,
         \MC_ARK_ARC_1_3/temp6[78] , \MC_ARK_ARC_1_3/temp6[77] ,
         \MC_ARK_ARC_1_3/temp6[75] , \MC_ARK_ARC_1_3/temp6[74] ,
         \MC_ARK_ARC_1_3/temp6[73] , \MC_ARK_ARC_1_3/temp6[72] ,
         \MC_ARK_ARC_1_3/temp6[71] , \MC_ARK_ARC_1_3/temp6[70] ,
         \MC_ARK_ARC_1_3/temp6[69] , \MC_ARK_ARC_1_3/temp6[67] ,
         \MC_ARK_ARC_1_3/temp6[65] , \MC_ARK_ARC_1_3/temp6[64] ,
         \MC_ARK_ARC_1_3/temp6[63] , \MC_ARK_ARC_1_3/temp6[61] ,
         \MC_ARK_ARC_1_3/temp6[60] , \MC_ARK_ARC_1_3/temp6[59] ,
         \MC_ARK_ARC_1_3/temp6[58] , \MC_ARK_ARC_1_3/temp6[57] ,
         \MC_ARK_ARC_1_3/temp6[56] , \MC_ARK_ARC_1_3/temp6[55] ,
         \MC_ARK_ARC_1_3/temp6[54] , \MC_ARK_ARC_1_3/temp6[52] ,
         \MC_ARK_ARC_1_3/temp6[49] , \MC_ARK_ARC_1_3/temp6[47] ,
         \MC_ARK_ARC_1_3/temp6[46] , \MC_ARK_ARC_1_3/temp6[42] ,
         \MC_ARK_ARC_1_3/temp6[40] , \MC_ARK_ARC_1_3/temp6[38] ,
         \MC_ARK_ARC_1_3/temp6[37] , \MC_ARK_ARC_1_3/temp6[36] ,
         \MC_ARK_ARC_1_3/temp6[34] , \MC_ARK_ARC_1_3/temp6[32] ,
         \MC_ARK_ARC_1_3/temp6[30] , \MC_ARK_ARC_1_3/temp6[29] ,
         \MC_ARK_ARC_1_3/temp6[27] , \MC_ARK_ARC_1_3/temp6[24] ,
         \MC_ARK_ARC_1_3/temp6[22] , \MC_ARK_ARC_1_3/temp6[21] ,
         \MC_ARK_ARC_1_3/temp6[20] , \MC_ARK_ARC_1_3/temp6[18] ,
         \MC_ARK_ARC_1_3/temp6[17] , \MC_ARK_ARC_1_3/temp6[16] ,
         \MC_ARK_ARC_1_3/temp6[15] , \MC_ARK_ARC_1_3/temp6[13] ,
         \MC_ARK_ARC_1_3/temp6[12] , \MC_ARK_ARC_1_3/temp6[11] ,
         \MC_ARK_ARC_1_3/temp6[8] , \MC_ARK_ARC_1_3/temp6[5] ,
         \MC_ARK_ARC_1_3/temp6[4] , \MC_ARK_ARC_1_3/temp6[3] ,
         \MC_ARK_ARC_1_3/temp6[2] , \MC_ARK_ARC_1_3/temp6[1] ,
         \MC_ARK_ARC_1_3/temp6[0] , \MC_ARK_ARC_1_3/temp5[190] ,
         \MC_ARK_ARC_1_3/temp5[185] , \MC_ARK_ARC_1_3/temp5[184] ,
         \MC_ARK_ARC_1_3/temp5[183] , \MC_ARK_ARC_1_3/temp5[182] ,
         \MC_ARK_ARC_1_3/temp5[181] , \MC_ARK_ARC_1_3/temp5[178] ,
         \MC_ARK_ARC_1_3/temp5[176] , \MC_ARK_ARC_1_3/temp5[173] ,
         \MC_ARK_ARC_1_3/temp5[172] , \MC_ARK_ARC_1_3/temp5[171] ,
         \MC_ARK_ARC_1_3/temp5[169] , \MC_ARK_ARC_1_3/temp5[168] ,
         \MC_ARK_ARC_1_3/temp5[167] , \MC_ARK_ARC_1_3/temp5[165] ,
         \MC_ARK_ARC_1_3/temp5[164] , \MC_ARK_ARC_1_3/temp5[163] ,
         \MC_ARK_ARC_1_3/temp5[162] , \MC_ARK_ARC_1_3/temp5[161] ,
         \MC_ARK_ARC_1_3/temp5[160] , \MC_ARK_ARC_1_3/temp5[159] ,
         \MC_ARK_ARC_1_3/temp5[157] , \MC_ARK_ARC_1_3/temp5[154] ,
         \MC_ARK_ARC_1_3/temp5[153] , \MC_ARK_ARC_1_3/temp5[152] ,
         \MC_ARK_ARC_1_3/temp5[151] , \MC_ARK_ARC_1_3/temp5[150] ,
         \MC_ARK_ARC_1_3/temp5[149] , \MC_ARK_ARC_1_3/temp5[147] ,
         \MC_ARK_ARC_1_3/temp5[145] , \MC_ARK_ARC_1_3/temp5[144] ,
         \MC_ARK_ARC_1_3/temp5[143] , \MC_ARK_ARC_1_3/temp5[142] ,
         \MC_ARK_ARC_1_3/temp5[141] , \MC_ARK_ARC_1_3/temp5[140] ,
         \MC_ARK_ARC_1_3/temp5[139] , \MC_ARK_ARC_1_3/temp5[137] ,
         \MC_ARK_ARC_1_3/temp5[136] , \MC_ARK_ARC_1_3/temp5[134] ,
         \MC_ARK_ARC_1_3/temp5[133] , \MC_ARK_ARC_1_3/temp5[132] ,
         \MC_ARK_ARC_1_3/temp5[131] , \MC_ARK_ARC_1_3/temp5[130] ,
         \MC_ARK_ARC_1_3/temp5[129] , \MC_ARK_ARC_1_3/temp5[128] ,
         \MC_ARK_ARC_1_3/temp5[126] , \MC_ARK_ARC_1_3/temp5[125] ,
         \MC_ARK_ARC_1_3/temp5[124] , \MC_ARK_ARC_1_3/temp5[123] ,
         \MC_ARK_ARC_1_3/temp5[122] , \MC_ARK_ARC_1_3/temp5[120] ,
         \MC_ARK_ARC_1_3/temp5[119] , \MC_ARK_ARC_1_3/temp5[118] ,
         \MC_ARK_ARC_1_3/temp5[117] , \MC_ARK_ARC_1_3/temp5[116] ,
         \MC_ARK_ARC_1_3/temp5[115] , \MC_ARK_ARC_1_3/temp5[114] ,
         \MC_ARK_ARC_1_3/temp5[112] , \MC_ARK_ARC_1_3/temp5[106] ,
         \MC_ARK_ARC_1_3/temp5[103] , \MC_ARK_ARC_1_3/temp5[101] ,
         \MC_ARK_ARC_1_3/temp5[100] , \MC_ARK_ARC_1_3/temp5[99] ,
         \MC_ARK_ARC_1_3/temp5[98] , \MC_ARK_ARC_1_3/temp5[97] ,
         \MC_ARK_ARC_1_3/temp5[96] , \MC_ARK_ARC_1_3/temp5[95] ,
         \MC_ARK_ARC_1_3/temp5[91] , \MC_ARK_ARC_1_3/temp5[88] ,
         \MC_ARK_ARC_1_3/temp5[86] , \MC_ARK_ARC_1_3/temp5[84] ,
         \MC_ARK_ARC_1_3/temp5[83] , \MC_ARK_ARC_1_3/temp5[82] ,
         \MC_ARK_ARC_1_3/temp5[79] , \MC_ARK_ARC_1_3/temp5[78] ,
         \MC_ARK_ARC_1_3/temp5[76] , \MC_ARK_ARC_1_3/temp5[75] ,
         \MC_ARK_ARC_1_3/temp5[74] , \MC_ARK_ARC_1_3/temp5[73] ,
         \MC_ARK_ARC_1_3/temp5[69] , \MC_ARK_ARC_1_3/temp5[64] ,
         \MC_ARK_ARC_1_3/temp5[62] , \MC_ARK_ARC_1_3/temp5[61] ,
         \MC_ARK_ARC_1_3/temp5[60] , \MC_ARK_ARC_1_3/temp5[59] ,
         \MC_ARK_ARC_1_3/temp5[56] , \MC_ARK_ARC_1_3/temp5[54] ,
         \MC_ARK_ARC_1_3/temp5[51] , \MC_ARK_ARC_1_3/temp5[50] ,
         \MC_ARK_ARC_1_3/temp5[49] , \MC_ARK_ARC_1_3/temp5[47] ,
         \MC_ARK_ARC_1_3/temp5[44] , \MC_ARK_ARC_1_3/temp5[42] ,
         \MC_ARK_ARC_1_3/temp5[41] , \MC_ARK_ARC_1_3/temp5[40] ,
         \MC_ARK_ARC_1_3/temp5[38] , \MC_ARK_ARC_1_3/temp5[37] ,
         \MC_ARK_ARC_1_3/temp5[36] , \MC_ARK_ARC_1_3/temp5[35] ,
         \MC_ARK_ARC_1_3/temp5[34] , \MC_ARK_ARC_1_3/temp5[33] ,
         \MC_ARK_ARC_1_3/temp5[32] , \MC_ARK_ARC_1_3/temp5[30] ,
         \MC_ARK_ARC_1_3/temp5[28] , \MC_ARK_ARC_1_3/temp5[27] ,
         \MC_ARK_ARC_1_3/temp5[25] , \MC_ARK_ARC_1_3/temp5[24] ,
         \MC_ARK_ARC_1_3/temp5[23] , \MC_ARK_ARC_1_3/temp5[22] ,
         \MC_ARK_ARC_1_3/temp5[21] , \MC_ARK_ARC_1_3/temp5[20] ,
         \MC_ARK_ARC_1_3/temp5[19] , \MC_ARK_ARC_1_3/temp5[18] ,
         \MC_ARK_ARC_1_3/temp5[17] , \MC_ARK_ARC_1_3/temp5[15] ,
         \MC_ARK_ARC_1_3/temp5[14] , \MC_ARK_ARC_1_3/temp5[13] ,
         \MC_ARK_ARC_1_3/temp5[11] , \MC_ARK_ARC_1_3/temp5[10] ,
         \MC_ARK_ARC_1_3/temp5[9] , \MC_ARK_ARC_1_3/temp5[7] ,
         \MC_ARK_ARC_1_3/temp5[6] , \MC_ARK_ARC_1_3/temp5[4] ,
         \MC_ARK_ARC_1_3/temp5[3] , \MC_ARK_ARC_1_3/temp4[191] ,
         \MC_ARK_ARC_1_3/temp4[190] , \MC_ARK_ARC_1_3/temp4[189] ,
         \MC_ARK_ARC_1_3/temp4[187] , \MC_ARK_ARC_1_3/temp4[186] ,
         \MC_ARK_ARC_1_3/temp4[184] , \MC_ARK_ARC_1_3/temp4[183] ,
         \MC_ARK_ARC_1_3/temp4[181] , \MC_ARK_ARC_1_3/temp4[180] ,
         \MC_ARK_ARC_1_3/temp4[179] , \MC_ARK_ARC_1_3/temp4[178] ,
         \MC_ARK_ARC_1_3/temp4[177] , \MC_ARK_ARC_1_3/temp4[175] ,
         \MC_ARK_ARC_1_3/temp4[174] , \MC_ARK_ARC_1_3/temp4[173] ,
         \MC_ARK_ARC_1_3/temp4[172] , \MC_ARK_ARC_1_3/temp4[171] ,
         \MC_ARK_ARC_1_3/temp4[170] , \MC_ARK_ARC_1_3/temp4[169] ,
         \MC_ARK_ARC_1_3/temp4[168] , \MC_ARK_ARC_1_3/temp4[167] ,
         \MC_ARK_ARC_1_3/temp4[165] , \MC_ARK_ARC_1_3/temp4[164] ,
         \MC_ARK_ARC_1_3/temp4[162] , \MC_ARK_ARC_1_3/temp4[161] ,
         \MC_ARK_ARC_1_3/temp4[160] , \MC_ARK_ARC_1_3/temp4[159] ,
         \MC_ARK_ARC_1_3/temp4[158] , \MC_ARK_ARC_1_3/temp4[157] ,
         \MC_ARK_ARC_1_3/temp4[156] , \MC_ARK_ARC_1_3/temp4[155] ,
         \MC_ARK_ARC_1_3/temp4[154] , \MC_ARK_ARC_1_3/temp4[152] ,
         \MC_ARK_ARC_1_3/temp4[151] , \MC_ARK_ARC_1_3/temp4[150] ,
         \MC_ARK_ARC_1_3/temp4[149] , \MC_ARK_ARC_1_3/temp4[148] ,
         \MC_ARK_ARC_1_3/temp4[147] , \MC_ARK_ARC_1_3/temp4[146] ,
         \MC_ARK_ARC_1_3/temp4[145] , \MC_ARK_ARC_1_3/temp4[144] ,
         \MC_ARK_ARC_1_3/temp4[143] , \MC_ARK_ARC_1_3/temp4[142] ,
         \MC_ARK_ARC_1_3/temp4[141] , \MC_ARK_ARC_1_3/temp4[140] ,
         \MC_ARK_ARC_1_3/temp4[139] , \MC_ARK_ARC_1_3/temp4[138] ,
         \MC_ARK_ARC_1_3/temp4[137] , \MC_ARK_ARC_1_3/temp4[136] ,
         \MC_ARK_ARC_1_3/temp4[135] , \MC_ARK_ARC_1_3/temp4[134] ,
         \MC_ARK_ARC_1_3/temp4[133] , \MC_ARK_ARC_1_3/temp4[132] ,
         \MC_ARK_ARC_1_3/temp4[131] , \MC_ARK_ARC_1_3/temp4[130] ,
         \MC_ARK_ARC_1_3/temp4[129] , \MC_ARK_ARC_1_3/temp4[128] ,
         \MC_ARK_ARC_1_3/temp4[127] , \MC_ARK_ARC_1_3/temp4[126] ,
         \MC_ARK_ARC_1_3/temp4[125] , \MC_ARK_ARC_1_3/temp4[124] ,
         \MC_ARK_ARC_1_3/temp4[123] , \MC_ARK_ARC_1_3/temp4[122] ,
         \MC_ARK_ARC_1_3/temp4[121] , \MC_ARK_ARC_1_3/temp4[120] ,
         \MC_ARK_ARC_1_3/temp4[119] , \MC_ARK_ARC_1_3/temp4[118] ,
         \MC_ARK_ARC_1_3/temp4[117] , \MC_ARK_ARC_1_3/temp4[116] ,
         \MC_ARK_ARC_1_3/temp4[115] , \MC_ARK_ARC_1_3/temp4[114] ,
         \MC_ARK_ARC_1_3/temp4[113] , \MC_ARK_ARC_1_3/temp4[112] ,
         \MC_ARK_ARC_1_3/temp4[111] , \MC_ARK_ARC_1_3/temp4[110] ,
         \MC_ARK_ARC_1_3/temp4[109] , \MC_ARK_ARC_1_3/temp4[108] ,
         \MC_ARK_ARC_1_3/temp4[106] , \MC_ARK_ARC_1_3/temp4[105] ,
         \MC_ARK_ARC_1_3/temp4[104] , \MC_ARK_ARC_1_3/temp4[102] ,
         \MC_ARK_ARC_1_3/temp4[100] , \MC_ARK_ARC_1_3/temp4[99] ,
         \MC_ARK_ARC_1_3/temp4[98] , \MC_ARK_ARC_1_3/temp4[97] ,
         \MC_ARK_ARC_1_3/temp4[96] , \MC_ARK_ARC_1_3/temp4[95] ,
         \MC_ARK_ARC_1_3/temp4[94] , \MC_ARK_ARC_1_3/temp4[93] ,
         \MC_ARK_ARC_1_3/temp4[92] , \MC_ARK_ARC_1_3/temp4[90] ,
         \MC_ARK_ARC_1_3/temp4[89] , \MC_ARK_ARC_1_3/temp4[88] ,
         \MC_ARK_ARC_1_3/temp4[87] , \MC_ARK_ARC_1_3/temp4[86] ,
         \MC_ARK_ARC_1_3/temp4[85] , \MC_ARK_ARC_1_3/temp4[84] ,
         \MC_ARK_ARC_1_3/temp4[83] , \MC_ARK_ARC_1_3/temp4[82] ,
         \MC_ARK_ARC_1_3/temp4[81] , \MC_ARK_ARC_1_3/temp4[80] ,
         \MC_ARK_ARC_1_3/temp4[79] , \MC_ARK_ARC_1_3/temp4[78] ,
         \MC_ARK_ARC_1_3/temp4[77] , \MC_ARK_ARC_1_3/temp4[76] ,
         \MC_ARK_ARC_1_3/temp4[75] , \MC_ARK_ARC_1_3/temp4[74] ,
         \MC_ARK_ARC_1_3/temp4[73] , \MC_ARK_ARC_1_3/temp4[72] ,
         \MC_ARK_ARC_1_3/temp4[71] , \MC_ARK_ARC_1_3/temp4[70] ,
         \MC_ARK_ARC_1_3/temp4[69] , \MC_ARK_ARC_1_3/temp4[68] ,
         \MC_ARK_ARC_1_3/temp4[67] , \MC_ARK_ARC_1_3/temp4[66] ,
         \MC_ARK_ARC_1_3/temp4[64] , \MC_ARK_ARC_1_3/temp4[63] ,
         \MC_ARK_ARC_1_3/temp4[61] , \MC_ARK_ARC_1_3/temp4[60] ,
         \MC_ARK_ARC_1_3/temp4[59] , \MC_ARK_ARC_1_3/temp4[58] ,
         \MC_ARK_ARC_1_3/temp4[57] , \MC_ARK_ARC_1_3/temp4[56] ,
         \MC_ARK_ARC_1_3/temp4[55] , \MC_ARK_ARC_1_3/temp4[54] ,
         \MC_ARK_ARC_1_3/temp4[53] , \MC_ARK_ARC_1_3/temp4[52] ,
         \MC_ARK_ARC_1_3/temp4[51] , \MC_ARK_ARC_1_3/temp4[50] ,
         \MC_ARK_ARC_1_3/temp4[49] , \MC_ARK_ARC_1_3/temp4[48] ,
         \MC_ARK_ARC_1_3/temp4[46] , \MC_ARK_ARC_1_3/temp4[45] ,
         \MC_ARK_ARC_1_3/temp4[44] , \MC_ARK_ARC_1_3/temp4[43] ,
         \MC_ARK_ARC_1_3/temp4[42] , \MC_ARK_ARC_1_3/temp4[41] ,
         \MC_ARK_ARC_1_3/temp4[40] , \MC_ARK_ARC_1_3/temp4[39] ,
         \MC_ARK_ARC_1_3/temp4[38] , \MC_ARK_ARC_1_3/temp4[37] ,
         \MC_ARK_ARC_1_3/temp4[36] , \MC_ARK_ARC_1_3/temp4[35] ,
         \MC_ARK_ARC_1_3/temp4[34] , \MC_ARK_ARC_1_3/temp4[33] ,
         \MC_ARK_ARC_1_3/temp4[32] , \MC_ARK_ARC_1_3/temp4[31] ,
         \MC_ARK_ARC_1_3/temp4[30] , \MC_ARK_ARC_1_3/temp4[29] ,
         \MC_ARK_ARC_1_3/temp4[28] , \MC_ARK_ARC_1_3/temp4[27] ,
         \MC_ARK_ARC_1_3/temp4[25] , \MC_ARK_ARC_1_3/temp4[24] ,
         \MC_ARK_ARC_1_3/temp4[23] , \MC_ARK_ARC_1_3/temp4[22] ,
         \MC_ARK_ARC_1_3/temp4[21] , \MC_ARK_ARC_1_3/temp4[20] ,
         \MC_ARK_ARC_1_3/temp4[19] , \MC_ARK_ARC_1_3/temp4[18] ,
         \MC_ARK_ARC_1_3/temp4[17] , \MC_ARK_ARC_1_3/temp4[16] ,
         \MC_ARK_ARC_1_3/temp4[15] , \MC_ARK_ARC_1_3/temp4[14] ,
         \MC_ARK_ARC_1_3/temp4[13] , \MC_ARK_ARC_1_3/temp4[12] ,
         \MC_ARK_ARC_1_3/temp4[11] , \MC_ARK_ARC_1_3/temp4[10] ,
         \MC_ARK_ARC_1_3/temp4[9] , \MC_ARK_ARC_1_3/temp4[8] ,
         \MC_ARK_ARC_1_3/temp4[7] , \MC_ARK_ARC_1_3/temp4[6] ,
         \MC_ARK_ARC_1_3/temp4[5] , \MC_ARK_ARC_1_3/temp4[4] ,
         \MC_ARK_ARC_1_3/temp4[3] , \MC_ARK_ARC_1_3/temp4[2] ,
         \MC_ARK_ARC_1_3/temp4[1] , \MC_ARK_ARC_1_3/temp4[0] ,
         \MC_ARK_ARC_1_3/temp3[191] , \MC_ARK_ARC_1_3/temp3[190] ,
         \MC_ARK_ARC_1_3/temp3[188] , \MC_ARK_ARC_1_3/temp3[186] ,
         \MC_ARK_ARC_1_3/temp3[184] , \MC_ARK_ARC_1_3/temp3[181] ,
         \MC_ARK_ARC_1_3/temp3[180] , \MC_ARK_ARC_1_3/temp3[178] ,
         \MC_ARK_ARC_1_3/temp3[177] , \MC_ARK_ARC_1_3/temp3[174] ,
         \MC_ARK_ARC_1_3/temp3[172] , \MC_ARK_ARC_1_3/temp3[171] ,
         \MC_ARK_ARC_1_3/temp3[169] , \MC_ARK_ARC_1_3/temp3[165] ,
         \MC_ARK_ARC_1_3/temp3[160] , \MC_ARK_ARC_1_3/temp3[159] ,
         \MC_ARK_ARC_1_3/temp3[157] , \MC_ARK_ARC_1_3/temp3[155] ,
         \MC_ARK_ARC_1_3/temp3[154] , \MC_ARK_ARC_1_3/temp3[152] ,
         \MC_ARK_ARC_1_3/temp3[151] , \MC_ARK_ARC_1_3/temp3[150] ,
         \MC_ARK_ARC_1_3/temp3[149] , \MC_ARK_ARC_1_3/temp3[148] ,
         \MC_ARK_ARC_1_3/temp3[147] , \MC_ARK_ARC_1_3/temp3[145] ,
         \MC_ARK_ARC_1_3/temp3[144] , \MC_ARK_ARC_1_3/temp3[143] ,
         \MC_ARK_ARC_1_3/temp3[142] , \MC_ARK_ARC_1_3/temp3[141] ,
         \MC_ARK_ARC_1_3/temp3[139] , \MC_ARK_ARC_1_3/temp3[138] ,
         \MC_ARK_ARC_1_3/temp3[137] , \MC_ARK_ARC_1_3/temp3[136] ,
         \MC_ARK_ARC_1_3/temp3[135] , \MC_ARK_ARC_1_3/temp3[133] ,
         \MC_ARK_ARC_1_3/temp3[132] , \MC_ARK_ARC_1_3/temp3[131] ,
         \MC_ARK_ARC_1_3/temp3[130] , \MC_ARK_ARC_1_3/temp3[129] ,
         \MC_ARK_ARC_1_3/temp3[127] , \MC_ARK_ARC_1_3/temp3[126] ,
         \MC_ARK_ARC_1_3/temp3[125] , \MC_ARK_ARC_1_3/temp3[124] ,
         \MC_ARK_ARC_1_3/temp3[122] , \MC_ARK_ARC_1_3/temp3[121] ,
         \MC_ARK_ARC_1_3/temp3[120] , \MC_ARK_ARC_1_3/temp3[119] ,
         \MC_ARK_ARC_1_3/temp3[117] , \MC_ARK_ARC_1_3/temp3[115] ,
         \MC_ARK_ARC_1_3/temp3[114] , \MC_ARK_ARC_1_3/temp3[112] ,
         \MC_ARK_ARC_1_3/temp3[111] , \MC_ARK_ARC_1_3/temp3[110] ,
         \MC_ARK_ARC_1_3/temp3[108] , \MC_ARK_ARC_1_3/temp3[106] ,
         \MC_ARK_ARC_1_3/temp3[105] , \MC_ARK_ARC_1_3/temp3[104] ,
         \MC_ARK_ARC_1_3/temp3[100] , \MC_ARK_ARC_1_3/temp3[98] ,
         \MC_ARK_ARC_1_3/temp3[97] , \MC_ARK_ARC_1_3/temp3[96] ,
         \MC_ARK_ARC_1_3/temp3[95] , \MC_ARK_ARC_1_3/temp3[94] ,
         \MC_ARK_ARC_1_3/temp3[92] , \MC_ARK_ARC_1_3/temp3[90] ,
         \MC_ARK_ARC_1_3/temp3[89] , \MC_ARK_ARC_1_3/temp3[88] ,
         \MC_ARK_ARC_1_3/temp3[86] , \MC_ARK_ARC_1_3/temp3[85] ,
         \MC_ARK_ARC_1_3/temp3[84] , \MC_ARK_ARC_1_3/temp3[82] ,
         \MC_ARK_ARC_1_3/temp3[81] , \MC_ARK_ARC_1_3/temp3[79] ,
         \MC_ARK_ARC_1_3/temp3[77] , \MC_ARK_ARC_1_3/temp3[76] ,
         \MC_ARK_ARC_1_3/temp3[75] , \MC_ARK_ARC_1_3/temp3[74] ,
         \MC_ARK_ARC_1_3/temp3[73] , \MC_ARK_ARC_1_3/temp3[72] ,
         \MC_ARK_ARC_1_3/temp3[71] , \MC_ARK_ARC_1_3/temp3[69] ,
         \MC_ARK_ARC_1_3/temp3[67] , \MC_ARK_ARC_1_3/temp3[66] ,
         \MC_ARK_ARC_1_3/temp3[64] , \MC_ARK_ARC_1_3/temp3[63] ,
         \MC_ARK_ARC_1_3/temp3[61] , \MC_ARK_ARC_1_3/temp3[60] ,
         \MC_ARK_ARC_1_3/temp3[56] , \MC_ARK_ARC_1_3/temp3[55] ,
         \MC_ARK_ARC_1_3/temp3[54] , \MC_ARK_ARC_1_3/temp3[52] ,
         \MC_ARK_ARC_1_3/temp3[51] , \MC_ARK_ARC_1_3/temp3[50] ,
         \MC_ARK_ARC_1_3/temp3[49] , \MC_ARK_ARC_1_3/temp3[46] ,
         \MC_ARK_ARC_1_3/temp3[45] , \MC_ARK_ARC_1_3/temp3[43] ,
         \MC_ARK_ARC_1_3/temp3[42] , \MC_ARK_ARC_1_3/temp3[41] ,
         \MC_ARK_ARC_1_3/temp3[40] , \MC_ARK_ARC_1_3/temp3[39] ,
         \MC_ARK_ARC_1_3/temp3[38] , \MC_ARK_ARC_1_3/temp3[37] ,
         \MC_ARK_ARC_1_3/temp3[36] , \MC_ARK_ARC_1_3/temp3[34] ,
         \MC_ARK_ARC_1_3/temp3[33] , \MC_ARK_ARC_1_3/temp3[32] ,
         \MC_ARK_ARC_1_3/temp3[31] , \MC_ARK_ARC_1_3/temp3[30] ,
         \MC_ARK_ARC_1_3/temp3[28] , \MC_ARK_ARC_1_3/temp3[24] ,
         \MC_ARK_ARC_1_3/temp3[23] , \MC_ARK_ARC_1_3/temp3[22] ,
         \MC_ARK_ARC_1_3/temp3[21] , \MC_ARK_ARC_1_3/temp3[20] ,
         \MC_ARK_ARC_1_3/temp3[19] , \MC_ARK_ARC_1_3/temp3[18] ,
         \MC_ARK_ARC_1_3/temp3[17] , \MC_ARK_ARC_1_3/temp3[16] ,
         \MC_ARK_ARC_1_3/temp3[15] , \MC_ARK_ARC_1_3/temp3[14] ,
         \MC_ARK_ARC_1_3/temp3[13] , \MC_ARK_ARC_1_3/temp3[12] ,
         \MC_ARK_ARC_1_3/temp3[11] , \MC_ARK_ARC_1_3/temp3[10] ,
         \MC_ARK_ARC_1_3/temp3[9] , \MC_ARK_ARC_1_3/temp3[7] ,
         \MC_ARK_ARC_1_3/temp3[6] , \MC_ARK_ARC_1_3/temp3[5] ,
         \MC_ARK_ARC_1_3/temp3[4] , \MC_ARK_ARC_1_3/temp3[3] ,
         \MC_ARK_ARC_1_3/temp3[2] , \MC_ARK_ARC_1_3/temp3[1] ,
         \MC_ARK_ARC_1_3/temp3[0] , \MC_ARK_ARC_1_3/temp2[191] ,
         \MC_ARK_ARC_1_3/temp2[187] , \MC_ARK_ARC_1_3/temp2[186] ,
         \MC_ARK_ARC_1_3/temp2[185] , \MC_ARK_ARC_1_3/temp2[184] ,
         \MC_ARK_ARC_1_3/temp2[183] , \MC_ARK_ARC_1_3/temp2[181] ,
         \MC_ARK_ARC_1_3/temp2[180] , \MC_ARK_ARC_1_3/temp2[178] ,
         \MC_ARK_ARC_1_3/temp2[177] , \MC_ARK_ARC_1_3/temp2[176] ,
         \MC_ARK_ARC_1_3/temp2[175] , \MC_ARK_ARC_1_3/temp2[173] ,
         \MC_ARK_ARC_1_3/temp2[172] , \MC_ARK_ARC_1_3/temp2[170] ,
         \MC_ARK_ARC_1_3/temp2[166] , \MC_ARK_ARC_1_3/temp2[165] ,
         \MC_ARK_ARC_1_3/temp2[163] , \MC_ARK_ARC_1_3/temp2[161] ,
         \MC_ARK_ARC_1_3/temp2[159] , \MC_ARK_ARC_1_3/temp2[156] ,
         \MC_ARK_ARC_1_3/temp2[155] , \MC_ARK_ARC_1_3/temp2[154] ,
         \MC_ARK_ARC_1_3/temp2[153] , \MC_ARK_ARC_1_3/temp2[152] ,
         \MC_ARK_ARC_1_3/temp2[150] , \MC_ARK_ARC_1_3/temp2[149] ,
         \MC_ARK_ARC_1_3/temp2[148] , \MC_ARK_ARC_1_3/temp2[147] ,
         \MC_ARK_ARC_1_3/temp2[146] , \MC_ARK_ARC_1_3/temp2[144] ,
         \MC_ARK_ARC_1_3/temp2[142] , \MC_ARK_ARC_1_3/temp2[141] ,
         \MC_ARK_ARC_1_3/temp2[140] , \MC_ARK_ARC_1_3/temp2[139] ,
         \MC_ARK_ARC_1_3/temp2[137] , \MC_ARK_ARC_1_3/temp2[136] ,
         \MC_ARK_ARC_1_3/temp2[135] , \MC_ARK_ARC_1_3/temp2[134] ,
         \MC_ARK_ARC_1_3/temp2[133] , \MC_ARK_ARC_1_3/temp2[132] ,
         \MC_ARK_ARC_1_3/temp2[130] , \MC_ARK_ARC_1_3/temp2[128] ,
         \MC_ARK_ARC_1_3/temp2[126] , \MC_ARK_ARC_1_3/temp2[125] ,
         \MC_ARK_ARC_1_3/temp2[124] , \MC_ARK_ARC_1_3/temp2[123] ,
         \MC_ARK_ARC_1_3/temp2[122] , \MC_ARK_ARC_1_3/temp2[120] ,
         \MC_ARK_ARC_1_3/temp2[118] , \MC_ARK_ARC_1_3/temp2[116] ,
         \MC_ARK_ARC_1_3/temp2[114] , \MC_ARK_ARC_1_3/temp2[113] ,
         \MC_ARK_ARC_1_3/temp2[111] , \MC_ARK_ARC_1_3/temp2[110] ,
         \MC_ARK_ARC_1_3/temp2[109] , \MC_ARK_ARC_1_3/temp2[108] ,
         \MC_ARK_ARC_1_3/temp2[107] , \MC_ARK_ARC_1_3/temp2[106] ,
         \MC_ARK_ARC_1_3/temp2[103] , \MC_ARK_ARC_1_3/temp2[102] ,
         \MC_ARK_ARC_1_3/temp2[100] , \MC_ARK_ARC_1_3/temp2[99] ,
         \MC_ARK_ARC_1_3/temp2[98] , \MC_ARK_ARC_1_3/temp2[97] ,
         \MC_ARK_ARC_1_3/temp2[96] , \MC_ARK_ARC_1_3/temp2[92] ,
         \MC_ARK_ARC_1_3/temp2[88] , \MC_ARK_ARC_1_3/temp2[86] ,
         \MC_ARK_ARC_1_3/temp2[85] , \MC_ARK_ARC_1_3/temp2[82] ,
         \MC_ARK_ARC_1_3/temp2[76] , \MC_ARK_ARC_1_3/temp2[74] ,
         \MC_ARK_ARC_1_3/temp2[73] , \MC_ARK_ARC_1_3/temp2[72] ,
         \MC_ARK_ARC_1_3/temp2[70] , \MC_ARK_ARC_1_3/temp2[67] ,
         \MC_ARK_ARC_1_3/temp2[66] , \MC_ARK_ARC_1_3/temp2[64] ,
         \MC_ARK_ARC_1_3/temp2[63] , \MC_ARK_ARC_1_3/temp2[62] ,
         \MC_ARK_ARC_1_3/temp2[61] , \MC_ARK_ARC_1_3/temp2[60] ,
         \MC_ARK_ARC_1_3/temp2[59] , \MC_ARK_ARC_1_3/temp2[58] ,
         \MC_ARK_ARC_1_3/temp2[57] , \MC_ARK_ARC_1_3/temp2[56] ,
         \MC_ARK_ARC_1_3/temp2[55] , \MC_ARK_ARC_1_3/temp2[54] ,
         \MC_ARK_ARC_1_3/temp2[53] , \MC_ARK_ARC_1_3/temp2[52] ,
         \MC_ARK_ARC_1_3/temp2[51] , \MC_ARK_ARC_1_3/temp2[49] ,
         \MC_ARK_ARC_1_3/temp2[48] , \MC_ARK_ARC_1_3/temp2[46] ,
         \MC_ARK_ARC_1_3/temp2[45] , \MC_ARK_ARC_1_3/temp2[43] ,
         \MC_ARK_ARC_1_3/temp2[42] , \MC_ARK_ARC_1_3/temp2[40] ,
         \MC_ARK_ARC_1_3/temp2[39] , \MC_ARK_ARC_1_3/temp2[38] ,
         \MC_ARK_ARC_1_3/temp2[37] , \MC_ARK_ARC_1_3/temp2[36] ,
         \MC_ARK_ARC_1_3/temp2[34] , \MC_ARK_ARC_1_3/temp2[33] ,
         \MC_ARK_ARC_1_3/temp2[30] , \MC_ARK_ARC_1_3/temp2[28] ,
         \MC_ARK_ARC_1_3/temp2[25] , \MC_ARK_ARC_1_3/temp2[24] ,
         \MC_ARK_ARC_1_3/temp2[22] , \MC_ARK_ARC_1_3/temp2[21] ,
         \MC_ARK_ARC_1_3/temp2[20] , \MC_ARK_ARC_1_3/temp2[19] ,
         \MC_ARK_ARC_1_3/temp2[18] , \MC_ARK_ARC_1_3/temp2[16] ,
         \MC_ARK_ARC_1_3/temp2[15] , \MC_ARK_ARC_1_3/temp2[14] ,
         \MC_ARK_ARC_1_3/temp2[13] , \MC_ARK_ARC_1_3/temp2[12] ,
         \MC_ARK_ARC_1_3/temp2[9] , \MC_ARK_ARC_1_3/temp2[7] ,
         \MC_ARK_ARC_1_3/temp2[4] , \MC_ARK_ARC_1_3/temp2[3] ,
         \MC_ARK_ARC_1_3/temp2[2] , \MC_ARK_ARC_1_3/temp2[1] ,
         \MC_ARK_ARC_1_3/temp2[0] , \MC_ARK_ARC_1_3/temp1[190] ,
         \MC_ARK_ARC_1_3/temp1[187] , \MC_ARK_ARC_1_3/temp1[186] ,
         \MC_ARK_ARC_1_3/temp1[184] , \MC_ARK_ARC_1_3/temp1[183] ,
         \MC_ARK_ARC_1_3/temp1[181] , \MC_ARK_ARC_1_3/temp1[180] ,
         \MC_ARK_ARC_1_3/temp1[178] , \MC_ARK_ARC_1_3/temp1[177] ,
         \MC_ARK_ARC_1_3/temp1[176] , \MC_ARK_ARC_1_3/temp1[175] ,
         \MC_ARK_ARC_1_3/temp1[174] , \MC_ARK_ARC_1_3/temp1[172] ,
         \MC_ARK_ARC_1_3/temp1[171] , \MC_ARK_ARC_1_3/temp1[169] ,
         \MC_ARK_ARC_1_3/temp1[168] , \MC_ARK_ARC_1_3/temp1[164] ,
         \MC_ARK_ARC_1_3/temp1[162] , \MC_ARK_ARC_1_3/temp1[157] ,
         \MC_ARK_ARC_1_3/temp1[156] , \MC_ARK_ARC_1_3/temp1[154] ,
         \MC_ARK_ARC_1_3/temp1[153] , \MC_ARK_ARC_1_3/temp1[152] ,
         \MC_ARK_ARC_1_3/temp1[151] , \MC_ARK_ARC_1_3/temp1[150] ,
         \MC_ARK_ARC_1_3/temp1[149] , \MC_ARK_ARC_1_3/temp1[148] ,
         \MC_ARK_ARC_1_3/temp1[146] , \MC_ARK_ARC_1_3/temp1[145] ,
         \MC_ARK_ARC_1_3/temp1[144] , \MC_ARK_ARC_1_3/temp1[143] ,
         \MC_ARK_ARC_1_3/temp1[139] , \MC_ARK_ARC_1_3/temp1[137] ,
         \MC_ARK_ARC_1_3/temp1[136] , \MC_ARK_ARC_1_3/temp1[135] ,
         \MC_ARK_ARC_1_3/temp1[134] , \MC_ARK_ARC_1_3/temp1[133] ,
         \MC_ARK_ARC_1_3/temp1[132] , \MC_ARK_ARC_1_3/temp1[131] ,
         \MC_ARK_ARC_1_3/temp1[130] , \MC_ARK_ARC_1_3/temp1[129] ,
         \MC_ARK_ARC_1_3/temp1[127] , \MC_ARK_ARC_1_3/temp1[126] ,
         \MC_ARK_ARC_1_3/temp1[125] , \MC_ARK_ARC_1_3/temp1[124] ,
         \MC_ARK_ARC_1_3/temp1[121] , \MC_ARK_ARC_1_3/temp1[118] ,
         \MC_ARK_ARC_1_3/temp1[115] , \MC_ARK_ARC_1_3/temp1[112] ,
         \MC_ARK_ARC_1_3/temp1[111] , \MC_ARK_ARC_1_3/temp1[110] ,
         \MC_ARK_ARC_1_3/temp1[109] , \MC_ARK_ARC_1_3/temp1[108] ,
         \MC_ARK_ARC_1_3/temp1[106] , \MC_ARK_ARC_1_3/temp1[104] ,
         \MC_ARK_ARC_1_3/temp1[103] , \MC_ARK_ARC_1_3/temp1[102] ,
         \MC_ARK_ARC_1_3/temp1[101] , \MC_ARK_ARC_1_3/temp1[100] ,
         \MC_ARK_ARC_1_3/temp1[99] , \MC_ARK_ARC_1_3/temp1[98] ,
         \MC_ARK_ARC_1_3/temp1[97] , \MC_ARK_ARC_1_3/temp1[96] ,
         \MC_ARK_ARC_1_3/temp1[94] , \MC_ARK_ARC_1_3/temp1[92] ,
         \MC_ARK_ARC_1_3/temp1[91] , \MC_ARK_ARC_1_3/temp1[90] ,
         \MC_ARK_ARC_1_3/temp1[89] , \MC_ARK_ARC_1_3/temp1[88] ,
         \MC_ARK_ARC_1_3/temp1[87] , \MC_ARK_ARC_1_3/temp1[85] ,
         \MC_ARK_ARC_1_3/temp1[84] , \MC_ARK_ARC_1_3/temp1[81] ,
         \MC_ARK_ARC_1_3/temp1[79] , \MC_ARK_ARC_1_3/temp1[76] ,
         \MC_ARK_ARC_1_3/temp1[75] , \MC_ARK_ARC_1_3/temp1[73] ,
         \MC_ARK_ARC_1_3/temp1[72] , \MC_ARK_ARC_1_3/temp1[70] ,
         \MC_ARK_ARC_1_3/temp1[67] , \MC_ARK_ARC_1_3/temp1[66] ,
         \MC_ARK_ARC_1_3/temp1[64] , \MC_ARK_ARC_1_3/temp1[62] ,
         \MC_ARK_ARC_1_3/temp1[61] , \MC_ARK_ARC_1_3/temp1[60] ,
         \MC_ARK_ARC_1_3/temp1[58] , \MC_ARK_ARC_1_3/temp1[57] ,
         \MC_ARK_ARC_1_3/temp1[55] , \MC_ARK_ARC_1_3/temp1[54] ,
         \MC_ARK_ARC_1_3/temp1[52] , \MC_ARK_ARC_1_3/temp1[51] ,
         \MC_ARK_ARC_1_3/temp1[49] , \MC_ARK_ARC_1_3/temp1[45] ,
         \MC_ARK_ARC_1_3/temp1[42] , \MC_ARK_ARC_1_3/temp1[41] ,
         \MC_ARK_ARC_1_3/temp1[40] , \MC_ARK_ARC_1_3/temp1[38] ,
         \MC_ARK_ARC_1_3/temp1[37] , \MC_ARK_ARC_1_3/temp1[36] ,
         \MC_ARK_ARC_1_3/temp1[35] , \MC_ARK_ARC_1_3/temp1[34] ,
         \MC_ARK_ARC_1_3/temp1[33] , \MC_ARK_ARC_1_3/temp1[32] ,
         \MC_ARK_ARC_1_3/temp1[31] , \MC_ARK_ARC_1_3/temp1[30] ,
         \MC_ARK_ARC_1_3/temp1[29] , \MC_ARK_ARC_1_3/temp1[28] ,
         \MC_ARK_ARC_1_3/temp1[27] , \MC_ARK_ARC_1_3/temp1[25] ,
         \MC_ARK_ARC_1_3/temp1[24] , \MC_ARK_ARC_1_3/temp1[23] ,
         \MC_ARK_ARC_1_3/temp1[22] , \MC_ARK_ARC_1_3/temp1[21] ,
         \MC_ARK_ARC_1_3/temp1[20] , \MC_ARK_ARC_1_3/temp1[19] ,
         \MC_ARK_ARC_1_3/temp1[18] , \MC_ARK_ARC_1_3/temp1[17] ,
         \MC_ARK_ARC_1_3/temp1[15] , \MC_ARK_ARC_1_3/temp1[13] ,
         \MC_ARK_ARC_1_3/temp1[12] , \MC_ARK_ARC_1_3/temp1[9] ,
         \MC_ARK_ARC_1_3/temp1[7] , \MC_ARK_ARC_1_3/temp1[6] ,
         \MC_ARK_ARC_1_3/temp1[4] , \MC_ARK_ARC_1_3/temp1[2] ,
         \MC_ARK_ARC_1_3/temp1[0] , \MC_ARK_ARC_1_3/buf_datainput[191] ,
         \MC_ARK_ARC_1_3/buf_datainput[182] ,
         \MC_ARK_ARC_1_3/buf_datainput[179] ,
         \MC_ARK_ARC_1_3/buf_datainput[178] ,
         \MC_ARK_ARC_1_3/buf_datainput[176] ,
         \MC_ARK_ARC_1_3/buf_datainput[174] ,
         \MC_ARK_ARC_1_3/buf_datainput[168] ,
         \MC_ARK_ARC_1_3/buf_datainput[166] ,
         \MC_ARK_ARC_1_3/buf_datainput[165] ,
         \MC_ARK_ARC_1_3/buf_datainput[155] ,
         \MC_ARK_ARC_1_3/buf_datainput[154] ,
         \MC_ARK_ARC_1_3/buf_datainput[152] ,
         \MC_ARK_ARC_1_3/buf_datainput[142] ,
         \MC_ARK_ARC_1_3/buf_datainput[135] ,
         \MC_ARK_ARC_1_3/buf_datainput[132] ,
         \MC_ARK_ARC_1_3/buf_datainput[122] ,
         \MC_ARK_ARC_1_3/buf_datainput[119] ,
         \MC_ARK_ARC_1_3/buf_datainput[116] ,
         \MC_ARK_ARC_1_3/buf_datainput[115] ,
         \MC_ARK_ARC_1_3/buf_datainput[114] ,
         \MC_ARK_ARC_1_3/buf_datainput[110] ,
         \MC_ARK_ARC_1_3/buf_datainput[109] ,
         \MC_ARK_ARC_1_3/buf_datainput[104] ,
         \MC_ARK_ARC_1_3/buf_datainput[103] ,
         \MC_ARK_ARC_1_3/buf_datainput[101] ,
         \MC_ARK_ARC_1_3/buf_datainput[97] ,
         \MC_ARK_ARC_1_3/buf_datainput[91] ,
         \MC_ARK_ARC_1_3/buf_datainput[90] ,
         \MC_ARK_ARC_1_3/buf_datainput[82] ,
         \MC_ARK_ARC_1_3/buf_datainput[81] ,
         \MC_ARK_ARC_1_3/buf_datainput[74] ,
         \MC_ARK_ARC_1_3/buf_datainput[71] ,
         \MC_ARK_ARC_1_3/buf_datainput[56] ,
         \MC_ARK_ARC_1_3/buf_datainput[53] ,
         \MC_ARK_ARC_1_3/buf_datainput[51] ,
         \MC_ARK_ARC_1_3/buf_datainput[49] ,
         \MC_ARK_ARC_1_3/buf_datainput[44] ,
         \MC_ARK_ARC_1_3/buf_datainput[41] ,
         \MC_ARK_ARC_1_3/buf_datainput[40] ,
         \MC_ARK_ARC_1_3/buf_datainput[38] ,
         \MC_ARK_ARC_1_3/buf_datainput[36] ,
         \MC_ARK_ARC_1_3/buf_datainput[28] ,
         \MC_ARK_ARC_1_3/buf_datainput[22] ,
         \MC_ARK_ARC_1_3/buf_datainput[17] ,
         \MC_ARK_ARC_1_3/buf_datainput[14] ,
         \MC_ARK_ARC_1_3/buf_datainput[12] , \MC_ARK_ARC_1_3/buf_datainput[6] ,
         \MC_ARK_ARC_1_3/buf_datainput[5] , \SB1_0_0/buf_output[5] ,
         \SB1_0_0/buf_output[4] , \SB1_0_0/buf_output[2] ,
         \SB1_0_0/buf_output[1] , \SB1_0_0/i3[0] , \SB1_0_0/i1_5 ,
         \SB1_0_0/i1_7 , \SB1_0_0/i1[9] , \SB1_0_0/i0_0 , \SB1_0_0/i0_3 ,
         \SB1_0_0/i0_4 , \SB1_0_0/i0[10] , \SB1_0_0/i0[9] , \SB1_0_0/i0[8] ,
         \SB1_0_0/i0[7] , \SB1_0_1/buf_output[5] , \SB1_0_1/buf_output[4] ,
         \SB1_0_1/buf_output[1] , \SB1_0_1/buf_output[0] , \SB1_0_1/i3[0] ,
         \SB1_0_1/i1_5 , \SB1_0_1/i1_7 , \SB1_0_1/i1[9] , \SB1_0_1/i0_0 ,
         \SB1_0_1/i0_3 , \SB1_0_1/i0_4 , \SB1_0_1/i0[10] , \SB1_0_1/i0[9] ,
         \SB1_0_1/i0[8] , \SB1_0_1/i0[7] , \SB1_0_1/i0[6] ,
         \SB1_0_2/buf_output[3] , \SB1_0_2/i3[0] , \SB1_0_2/i1_5 ,
         \SB1_0_2/i1_7 , \SB1_0_2/i1[9] , \SB1_0_2/i0_0 , \SB1_0_2/i0_3 ,
         \SB1_0_2/i0_4 , \SB1_0_2/i0[10] , \SB1_0_2/i0[9] , \SB1_0_2/i0[8] ,
         \SB1_0_2/i0[7] , \SB1_0_2/i0[6] , \SB1_0_3/buf_output[5] ,
         \SB1_0_3/buf_output[0] , \SB1_0_3/i3[0] , \SB1_0_3/i1_5 ,
         \SB1_0_3/i1_7 , \SB1_0_3/i1[9] , \SB1_0_3/i0_0 , \SB1_0_3/i0_3 ,
         \SB1_0_3/i0_4 , \SB1_0_3/i0[10] , \SB1_0_3/i0[9] , \SB1_0_3/i0[8] ,
         \SB1_0_3/i0[7] , \SB1_0_3/i0[6] , \SB1_0_4/buf_output[5] ,
         \SB1_0_4/buf_output[4] , \SB1_0_4/buf_output[1] ,
         \SB1_0_4/buf_output[0] , \SB1_0_4/i3[0] , \SB1_0_4/i1_5 ,
         \SB1_0_4/i1_7 , \SB1_0_4/i1[9] , \SB1_0_4/i0_0 , \SB1_0_4/i0_3 ,
         \SB1_0_4/i0_4 , \SB1_0_4/i0[10] , \SB1_0_4/i0[9] , \SB1_0_4/i0[8] ,
         \SB1_0_4/i0[7] , \SB1_0_4/i0[6] , \SB1_0_5/buf_output[4] ,
         \SB1_0_5/buf_output[3] , \SB1_0_5/buf_output[2] ,
         \SB1_0_5/buf_output[1] , \SB1_0_5/buf_output[0] , \SB1_0_5/i3[0] ,
         \SB1_0_5/i1_5 , \SB1_0_5/i1_7 , \SB1_0_5/i1[9] , \SB1_0_5/i0_0 ,
         \SB1_0_5/i0_3 , \SB1_0_5/i0_4 , \SB1_0_5/i0[10] , \SB1_0_5/i0[9] ,
         \SB1_0_5/i0[8] , \SB1_0_5/i0[7] , \SB1_0_5/i0[6] ,
         \SB1_0_6/buf_output[5] , \SB1_0_6/buf_output[2] , \SB1_0_6/i3[0] ,
         \SB1_0_6/i1_5 , \SB1_0_6/i1_7 , \SB1_0_6/i1[9] , \SB1_0_6/i0_0 ,
         \SB1_0_6/i0_3 , \SB1_0_6/i0_4 , \SB1_0_6/i0[10] , \SB1_0_6/i0[9] ,
         \SB1_0_6/i0[8] , \SB1_0_6/i0[7] , \SB1_0_6/i0[6] ,
         \SB1_0_7/buf_output[3] , \SB1_0_7/buf_output[1] ,
         \SB1_0_7/buf_output[0] , \SB1_0_7/i3[0] , \SB1_0_7/i1_5 ,
         \SB1_0_7/i1_7 , \SB1_0_7/i1[9] , \SB1_0_7/i0_0 , \SB1_0_7/i0_3 ,
         \SB1_0_7/i0[10] , \SB1_0_7/i0[9] , \SB1_0_7/i0[8] , \SB1_0_7/i0[7] ,
         \SB1_0_7/i0[6] , \SB1_0_8/buf_output[5] , \SB1_0_8/buf_output[4] ,
         \SB1_0_8/buf_output[0] , \SB1_0_8/i3[0] , \SB1_0_8/i1_5 ,
         \SB1_0_8/i1_7 , \SB1_0_8/i1[9] , \SB1_0_8/i0_0 , \SB1_0_8/i0_3 ,
         \SB1_0_8/i0_4 , \SB1_0_8/i0[10] , \SB1_0_8/i0[9] , \SB1_0_8/i0[8] ,
         \SB1_0_8/i0[7] , \SB1_0_8/i0[6] , \SB1_0_9/buf_output[5] ,
         \SB1_0_9/buf_output[4] , \SB1_0_9/buf_output[1] , \SB1_0_9/i3[0] ,
         \SB1_0_9/i1_5 , \SB1_0_9/i1_7 , \SB1_0_9/i1[9] , \SB1_0_9/i0_0 ,
         \SB1_0_9/i0_3 , \SB1_0_9/i0_4 , \SB1_0_9/i0[10] , \SB1_0_9/i0[9] ,
         \SB1_0_9/i0[8] , \SB1_0_9/i0[7] , \SB1_0_9/i0[6] ,
         \SB1_0_10/buf_output[3] , \SB1_0_10/buf_output[1] ,
         \SB1_0_10/buf_output[0] , \SB1_0_10/i3[0] , \SB1_0_10/i1_5 ,
         \SB1_0_10/i1_7 , \SB1_0_10/i1[9] , \SB1_0_10/i0_0 , \SB1_0_10/i0_3 ,
         \SB1_0_10/i0_4 , \SB1_0_10/i0[10] , \SB1_0_10/i0[9] ,
         \SB1_0_10/i0[8] , \SB1_0_10/i0[7] , \SB1_0_10/i0[6] ,
         \SB1_0_11/buf_output[5] , \SB1_0_11/buf_output[3] ,
         \SB1_0_11/buf_output[2] , \SB1_0_11/buf_output[0] , \SB1_0_11/i3[0] ,
         \SB1_0_11/i1_5 , \SB1_0_11/i1_7 , \SB1_0_11/i1[9] , \SB1_0_11/i0_0 ,
         \SB1_0_11/i0_3 , \SB1_0_11/i0_4 , \SB1_0_11/i0[10] , \SB1_0_11/i0[9] ,
         \SB1_0_11/i0[8] , \SB1_0_11/i0[7] , \SB1_0_11/i0[6] ,
         \SB1_0_12/buf_output[5] , \SB1_0_12/buf_output[2] ,
         \SB1_0_12/buf_output[0] , \SB1_0_12/i3[0] , \SB1_0_12/i1_5 ,
         \SB1_0_12/i1_7 , \SB1_0_12/i1[9] , \SB1_0_12/i0_0 , \SB1_0_12/i0_3 ,
         \SB1_0_12/i0_4 , \SB1_0_12/i0[10] , \SB1_0_12/i0[9] ,
         \SB1_0_12/i0[8] , \SB1_0_12/i0[7] , \SB1_0_12/i0[6] ,
         \SB1_0_13/buf_output[2] , \SB1_0_13/buf_output[1] ,
         \SB1_0_13/buf_output[0] , \SB1_0_13/i3[0] , \SB1_0_13/i1_5 ,
         \SB1_0_13/i1_7 , \SB1_0_13/i1[9] , \SB1_0_13/i0_0 , \SB1_0_13/i0_3 ,
         \SB1_0_13/i0_4 , \SB1_0_13/i0[10] , \SB1_0_13/i0[9] ,
         \SB1_0_13/i0[8] , \SB1_0_13/i0[7] , \SB1_0_13/i0[6] ,
         \SB1_0_14/buf_output[3] , \SB1_0_14/buf_output[2] ,
         \SB1_0_14/buf_output[0] , \SB1_0_14/i3[0] , \SB1_0_14/i1_5 ,
         \SB1_0_14/i1_7 , \SB1_0_14/i1[9] , \SB1_0_14/i0_0 , \SB1_0_14/i0_3 ,
         \SB1_0_14/i0_4 , \SB1_0_14/i0[10] , \SB1_0_14/i0[9] ,
         \SB1_0_14/i0[8] , \SB1_0_14/i0[7] , \SB1_0_14/i0[6] ,
         \SB1_0_15/buf_output[5] , \SB1_0_15/buf_output[4] ,
         \SB1_0_15/buf_output[3] , \SB1_0_15/i3[0] , \SB1_0_15/i1_5 ,
         \SB1_0_15/i1_7 , \SB1_0_15/i1[9] , \SB1_0_15/i0_0 , \SB1_0_15/i0_3 ,
         \SB1_0_15/i0_4 , \SB1_0_15/i0[10] , \SB1_0_15/i0[9] ,
         \SB1_0_15/i0[8] , \SB1_0_15/i0[7] , \SB1_0_15/i0[6] ,
         \SB1_0_16/buf_output[4] , \SB1_0_16/buf_output[3] ,
         \SB1_0_16/buf_output[2] , \SB1_0_16/buf_output[1] , \SB1_0_16/i3[0] ,
         \SB1_0_16/i1_5 , \SB1_0_16/i1_7 , \SB1_0_16/i1[9] , \SB1_0_16/i0_0 ,
         \SB1_0_16/i0_3 , \SB1_0_16/i0[10] , \SB1_0_16/i0[9] ,
         \SB1_0_16/i0[8] , \SB1_0_16/i0[7] , \SB1_0_16/i0[6] ,
         \SB1_0_17/buf_output[5] , \SB1_0_17/buf_output[2] ,
         \SB1_0_17/buf_output[1] , \SB1_0_17/i3[0] , \SB1_0_17/i1_5 ,
         \SB1_0_17/i1_7 , \SB1_0_17/i1[9] , \SB1_0_17/i0_0 , \SB1_0_17/i0_3 ,
         \SB1_0_17/i0[10] , \SB1_0_17/i0[9] , \SB1_0_17/i0[8] ,
         \SB1_0_17/i0[7] , \SB1_0_17/i0[6] , \SB1_0_18/buf_output[5] ,
         \SB1_0_18/buf_output[4] , \SB1_0_18/buf_output[2] ,
         \SB1_0_18/buf_output[0] , \SB1_0_18/i3[0] , \SB1_0_18/i1_5 ,
         \SB1_0_18/i1_7 , \SB1_0_18/i1[9] , \SB1_0_18/i0_0 , \SB1_0_18/i0_3 ,
         \SB1_0_18/i0[9] , \SB1_0_18/i0[8] , \SB1_0_18/i0[7] ,
         \SB1_0_18/i0[6] , \SB1_0_19/buf_output[5] , \SB1_0_19/buf_output[4] ,
         \SB1_0_19/buf_output[3] , \SB1_0_19/buf_output[0] , \SB1_0_19/i3[0] ,
         \SB1_0_19/i1_5 , \SB1_0_19/i1_7 , \SB1_0_19/i1[9] , \SB1_0_19/i0_0 ,
         \SB1_0_19/i0_3 , \SB1_0_19/i0_4 , \SB1_0_19/i0[10] , \SB1_0_19/i0[9] ,
         \SB1_0_19/i0[8] , \SB1_0_19/i0[7] , \SB1_0_19/i0[6] ,
         \SB1_0_20/buf_output[5] , \SB1_0_20/i3[0] , \SB1_0_20/i1_5 ,
         \SB1_0_20/i1_7 , \SB1_0_20/i1[9] , \SB1_0_20/i0_0 , \SB1_0_20/i0_3 ,
         \SB1_0_20/i0_4 , \SB1_0_20/i0[10] , \SB1_0_20/i0[9] ,
         \SB1_0_20/i0[8] , \SB1_0_20/i0[7] , \SB1_0_20/i0[6] ,
         \SB1_0_21/buf_output[5] , \SB1_0_21/buf_output[1] ,
         \SB1_0_21/buf_output[0] , \SB1_0_21/i3[0] , \SB1_0_21/i1_5 ,
         \SB1_0_21/i1_7 , \SB1_0_21/i1[9] , \SB1_0_21/i0_0 , \SB1_0_21/i0_3 ,
         \SB1_0_21/i0_4 , \SB1_0_21/i0[10] , \SB1_0_21/i0[9] ,
         \SB1_0_21/i0[8] , \SB1_0_21/i0[7] , \SB1_0_21/i0[6] ,
         \SB1_0_22/buf_output[5] , \SB1_0_22/buf_output[4] ,
         \SB1_0_22/buf_output[2] , \SB1_0_22/i3[0] , \SB1_0_22/i1_5 ,
         \SB1_0_22/i1_7 , \SB1_0_22/i1[9] , \SB1_0_22/i0_0 , \SB1_0_22/i0_3 ,
         \SB1_0_22/i0_4 , \SB1_0_22/i0[10] , \SB1_0_22/i0[9] ,
         \SB1_0_22/i0[8] , \SB1_0_22/i0[7] , \SB1_0_22/i0[6] ,
         \SB1_0_23/buf_output[5] , \SB1_0_23/buf_output[1] ,
         \SB1_0_23/buf_output[0] , \SB1_0_23/i3[0] , \SB1_0_23/i1_5 ,
         \SB1_0_23/i1_7 , \SB1_0_23/i1[9] , \SB1_0_23/i0_0 , \SB1_0_23/i0_3 ,
         \SB1_0_23/i0_4 , \SB1_0_23/i0[10] , \SB1_0_23/i0[9] ,
         \SB1_0_23/i0[8] , \SB1_0_23/i0[7] , \SB1_0_23/i0[6] ,
         \SB1_0_24/buf_output[5] , \SB1_0_24/i3[0] , \SB1_0_24/i1_5 ,
         \SB1_0_24/i1_7 , \SB1_0_24/i1[9] , \SB1_0_24/i0_0 , \SB1_0_24/i0_3 ,
         \SB1_0_24/i0_4 , \SB1_0_24/i0[10] , \SB1_0_24/i0[9] ,
         \SB1_0_24/i0[8] , \SB1_0_24/i0[7] , \SB1_0_24/i0[6] ,
         \SB1_0_25/buf_output[5] , \SB1_0_25/buf_output[3] ,
         \SB1_0_25/buf_output[2] , \SB1_0_25/i3[0] , \SB1_0_25/i1_5 ,
         \SB1_0_25/i1_7 , \SB1_0_25/i1[9] , \SB1_0_25/i0_0 , \SB1_0_25/i0_3 ,
         \SB1_0_25/i0_4 , \SB1_0_25/i0[10] , \SB1_0_25/i0[9] ,
         \SB1_0_25/i0[8] , \SB1_0_25/i0[7] , \SB1_0_25/i0[6] ,
         \SB1_0_26/buf_output[5] , \SB1_0_26/buf_output[4] ,
         \SB1_0_26/buf_output[0] , \SB1_0_26/i3[0] , \SB1_0_26/i1_5 ,
         \SB1_0_26/i1_7 , \SB1_0_26/i1[9] , \SB1_0_26/i0_0 , \SB1_0_26/i0_3 ,
         \SB1_0_26/i0_4 , \SB1_0_26/i0[10] , \SB1_0_26/i0[9] ,
         \SB1_0_26/i0[8] , \SB1_0_26/i0[7] , \SB1_0_26/i0[6] ,
         \SB1_0_27/buf_output[5] , \SB1_0_27/buf_output[4] ,
         \SB1_0_27/buf_output[0] , \SB1_0_27/i3[0] , \SB1_0_27/i1_5 ,
         \SB1_0_27/i1_7 , \SB1_0_27/i1[9] , \SB1_0_27/i0_0 , \SB1_0_27/i0_3 ,
         \SB1_0_27/i0_4 , \SB1_0_27/i0[10] , \SB1_0_27/i0[9] ,
         \SB1_0_27/i0[8] , \SB1_0_27/i0[7] , \SB1_0_27/i0[6] ,
         \SB1_0_28/buf_output[2] , \SB1_0_28/buf_output[1] , \SB1_0_28/i3[0] ,
         \SB1_0_28/i1_5 , \SB1_0_28/i1_7 , \SB1_0_28/i1[9] , \SB1_0_28/i0_0 ,
         \SB1_0_28/i0_3 , \SB1_0_28/i0_4 , \SB1_0_28/i0[10] , \SB1_0_28/i0[9] ,
         \SB1_0_28/i0[8] , \SB1_0_28/i0[7] , \SB1_0_28/i0[6] ,
         \SB1_0_29/buf_output[5] , \SB1_0_29/buf_output[1] ,
         \SB1_0_29/buf_output[0] , \SB1_0_29/i3[0] , \SB1_0_29/i1_5 ,
         \SB1_0_29/i1_7 , \SB1_0_29/i1[9] , \SB1_0_29/i0_0 , \SB1_0_29/i0_3 ,
         \SB1_0_29/i0_4 , \SB1_0_29/i0[10] , \SB1_0_29/i0[9] ,
         \SB1_0_29/i0[8] , \SB1_0_29/i0[7] , \SB1_0_29/i0[6] ,
         \SB1_0_30/buf_output[5] , \SB1_0_30/buf_output[4] ,
         \SB1_0_30/buf_output[3] , \SB1_0_30/buf_output[2] ,
         \SB1_0_30/buf_output[1] , \SB1_0_30/buf_output[0] , \SB1_0_30/i3[0] ,
         \SB1_0_30/i1_5 , \SB1_0_30/i1_7 , \SB1_0_30/i1[9] , \SB1_0_30/i0_0 ,
         \SB1_0_30/i0_3 , \SB1_0_30/i0_4 , \SB1_0_30/i0[10] , \SB1_0_30/i0[9] ,
         \SB1_0_30/i0[8] , \SB1_0_30/i0[7] , \SB1_0_30/i0[6] ,
         \SB1_0_31/buf_output[3] , \SB1_0_31/buf_output[1] , \SB1_0_31/i3[0] ,
         \SB1_0_31/i1_5 , \SB1_0_31/i1_7 , \SB1_0_31/i1[9] , \SB1_0_31/i0_0 ,
         \SB1_0_31/i0_3 , \SB1_0_31/i0_4 , \SB1_0_31/i0[10] , \SB1_0_31/i0[9] ,
         \SB1_0_31/i0[8] , \SB1_0_31/i0[7] , \SB1_0_31/i0[6] ,
         \SB2_0_0/buf_output[5] , \SB2_0_0/buf_output[4] ,
         \SB2_0_0/buf_output[3] , \SB2_0_0/buf_output[2] ,
         \SB2_0_0/buf_output[1] , \SB2_0_0/buf_output[0] , \SB2_0_0/i3[0] ,
         \SB2_0_0/i1_5 , \SB2_0_0/i1_7 , \SB2_0_0/i1[9] , \SB2_0_0/i0_0 ,
         \SB2_0_0/i0[10] , \SB2_0_0/i0[9] , \SB2_0_0/i0[8] , \SB2_0_0/i0[7] ,
         \SB2_0_0/i0[6] , \SB2_0_1/buf_output[5] , \SB2_0_1/buf_output[4] ,
         \SB2_0_1/buf_output[3] , \SB2_0_1/buf_output[2] ,
         \SB2_0_1/buf_output[1] , \SB2_0_1/buf_output[0] , \SB2_0_1/i3[0] ,
         \SB2_0_1/i1_5 , \SB2_0_1/i1_7 , \SB2_0_1/i1[9] , \SB2_0_1/i0_0 ,
         \SB2_0_1/i0_3 , \SB2_0_1/i0_4 , \SB2_0_1/i0[10] , \SB2_0_1/i0[9] ,
         \SB2_0_1/i0[8] , \SB2_0_1/i0[6] , \SB2_0_2/buf_output[5] ,
         \SB2_0_2/buf_output[4] , \SB2_0_2/buf_output[3] ,
         \SB2_0_2/buf_output[2] , \SB2_0_2/buf_output[1] ,
         \SB2_0_2/buf_output[0] , \SB2_0_2/i3[0] , \SB2_0_2/i1_5 ,
         \SB2_0_2/i1_7 , \SB2_0_2/i1[9] , \SB2_0_2/i0_3 , \SB2_0_2/i0[10] ,
         \SB2_0_2/i0[9] , \SB2_0_2/i0[8] , \SB2_0_2/i0[7] , \SB2_0_2/i0[6] ,
         \SB2_0_3/buf_output[5] , \SB2_0_3/buf_output[4] ,
         \SB2_0_3/buf_output[3] , \SB2_0_3/buf_output[2] ,
         \SB2_0_3/buf_output[1] , \SB2_0_3/buf_output[0] , \SB2_0_3/i3[0] ,
         \SB2_0_3/i1_5 , \SB2_0_3/i1_7 , \SB2_0_3/i1[9] , \SB2_0_3/i0_0 ,
         \SB2_0_3/i0_3 , \SB2_0_3/i0[10] , \SB2_0_3/i0[9] , \SB2_0_3/i0[8] ,
         \SB2_0_3/i0[7] , \SB2_0_3/i0[6] , \SB2_0_4/buf_output[5] ,
         \SB2_0_4/buf_output[4] , \SB2_0_4/buf_output[3] ,
         \SB2_0_4/buf_output[2] , \SB2_0_4/buf_output[1] ,
         \SB2_0_4/buf_output[0] , \SB2_0_4/i3[0] , \SB2_0_4/i1_5 ,
         \SB2_0_4/i1_7 , \SB2_0_4/i1[9] , \SB2_0_4/i0_0 , \SB2_0_4/i0_3 ,
         \SB2_0_4/i0[10] , \SB2_0_4/i0[9] , \SB2_0_4/i0[8] , \SB2_0_4/i0[7] ,
         \SB2_0_4/i0[6] , \SB2_0_5/buf_output[5] , \SB2_0_5/buf_output[4] ,
         \SB2_0_5/buf_output[3] , \SB2_0_5/buf_output[2] ,
         \SB2_0_5/buf_output[1] , \SB2_0_5/buf_output[0] , \SB2_0_5/i3[0] ,
         \SB2_0_5/i1_5 , \SB2_0_5/i1_7 , \SB2_0_5/i0_0 , \SB2_0_5/i0_3 ,
         \SB2_0_5/i0[10] , \SB2_0_5/i0[8] , \SB2_0_5/i0[7] , \SB2_0_5/i0[6] ,
         \SB2_0_6/buf_output[5] , \SB2_0_6/buf_output[4] ,
         \SB2_0_6/buf_output[3] , \SB2_0_6/buf_output[2] ,
         \SB2_0_6/buf_output[1] , \SB2_0_6/buf_output[0] , \SB2_0_6/i3[0] ,
         \SB2_0_6/i1_5 , \SB2_0_6/i1_7 , \SB2_0_6/i1[9] , \SB2_0_6/i0_0 ,
         \SB2_0_6/i0[10] , \SB2_0_6/i0[9] , \SB2_0_6/i0[8] , \SB2_0_6/i0[7] ,
         \SB2_0_6/i0[6] , \SB2_0_7/buf_output[5] , \SB2_0_7/buf_output[4] ,
         \SB2_0_7/buf_output[3] , \SB2_0_7/buf_output[2] ,
         \SB2_0_7/buf_output[1] , \SB2_0_7/buf_output[0] , \SB2_0_7/i3[0] ,
         \SB2_0_7/i1_5 , \SB2_0_7/i1_7 , \SB2_0_7/i1[9] , \SB2_0_7/i0_0 ,
         \SB2_0_7/i0_3 , \SB2_0_7/i0[10] , \SB2_0_7/i0[9] , \SB2_0_7/i0[8] ,
         \SB2_0_7/i0[7] , \SB2_0_7/i0[6] , \SB2_0_8/buf_output[5] ,
         \SB2_0_8/buf_output[4] , \SB2_0_8/buf_output[3] ,
         \SB2_0_8/buf_output[2] , \SB2_0_8/buf_output[1] ,
         \SB2_0_8/buf_output[0] , \SB2_0_8/i3[0] , \SB2_0_8/i1_5 ,
         \SB2_0_8/i1_7 , \SB2_0_8/i1[9] , \SB2_0_8/i0_0 , \SB2_0_8/i0_3 ,
         \SB2_0_8/i0[10] , \SB2_0_8/i0[9] , \SB2_0_8/i0[8] , \SB2_0_8/i0[7] ,
         \SB2_0_8/i0[6] , \SB2_0_9/buf_output[5] , \SB2_0_9/buf_output[4] ,
         \SB2_0_9/buf_output[3] , \SB2_0_9/buf_output[2] ,
         \SB2_0_9/buf_output[1] , \SB2_0_9/buf_output[0] , \SB2_0_9/i3[0] ,
         \SB2_0_9/i1_7 , \SB2_0_9/i1[9] , \SB2_0_9/i0_3 , \SB2_0_9/i0_4 ,
         \SB2_0_9/i0[10] , \SB2_0_9/i0[9] , \SB2_0_9/i0[8] , \SB2_0_9/i0[7] ,
         \SB2_0_9/i0[6] , \SB2_0_10/buf_output[5] , \SB2_0_10/buf_output[4] ,
         \SB2_0_10/buf_output[3] , \SB2_0_10/buf_output[2] ,
         \SB2_0_10/buf_output[1] , \SB2_0_10/buf_output[0] , \SB2_0_10/i3[0] ,
         \SB2_0_10/i1_5 , \SB2_0_10/i1_7 , \SB2_0_10/i1[9] , \SB2_0_10/i0_0 ,
         \SB2_0_10/i0_3 , \SB2_0_10/i0_4 , \SB2_0_10/i0[10] , \SB2_0_10/i0[8] ,
         \SB2_0_10/i0[6] , \SB2_0_11/buf_output[5] , \SB2_0_11/buf_output[4] ,
         \SB2_0_11/buf_output[3] , \SB2_0_11/buf_output[2] ,
         \SB2_0_11/buf_output[1] , \SB2_0_11/buf_output[0] , \SB2_0_11/i3[0] ,
         \SB2_0_11/i1_5 , \SB2_0_11/i1_7 , \SB2_0_11/i1[9] , \SB2_0_11/i0_0 ,
         \SB2_0_11/i0_3 , \SB2_0_11/i0_4 , \SB2_0_11/i0[10] , \SB2_0_11/i0[9] ,
         \SB2_0_11/i0[8] , \SB2_0_11/i0[7] , \SB2_0_11/i0[6] ,
         \SB2_0_12/buf_output[5] , \SB2_0_12/buf_output[4] ,
         \SB2_0_12/buf_output[3] , \SB2_0_12/buf_output[2] ,
         \SB2_0_12/buf_output[1] , \SB2_0_12/buf_output[0] , \SB2_0_12/i3[0] ,
         \SB2_0_12/i1_5 , \SB2_0_12/i1_7 , \SB2_0_12/i1[9] , \SB2_0_12/i0_0 ,
         \SB2_0_12/i0_3 , \SB2_0_12/i0_4 , \SB2_0_12/i0[10] , \SB2_0_12/i0[9] ,
         \SB2_0_12/i0[8] , \SB2_0_12/i0[7] , \SB2_0_12/i0[6] ,
         \SB2_0_13/buf_output[5] , \SB2_0_13/buf_output[4] ,
         \SB2_0_13/buf_output[3] , \SB2_0_13/buf_output[2] ,
         \SB2_0_13/buf_output[1] , \SB2_0_13/buf_output[0] , \SB2_0_13/i3[0] ,
         \SB2_0_13/i1_7 , \SB2_0_13/i1[9] , \SB2_0_13/i0_0 , \SB2_0_13/i0_3 ,
         \SB2_0_13/i0_4 , \SB2_0_13/i0[10] , \SB2_0_13/i0[9] ,
         \SB2_0_13/i0[6] , \SB2_0_14/buf_output[5] , \SB2_0_14/buf_output[4] ,
         \SB2_0_14/buf_output[3] , \SB2_0_14/buf_output[2] ,
         \SB2_0_14/buf_output[1] , \SB2_0_14/buf_output[0] , \SB2_0_14/i3[0] ,
         \SB2_0_14/i1_5 , \SB2_0_14/i1_7 , \SB2_0_14/i1[9] , \SB2_0_14/i0_3 ,
         \SB2_0_14/i0[9] , \SB2_0_14/i0[8] , \SB2_0_14/i0[7] ,
         \SB2_0_14/i0[6] , \SB2_0_15/buf_output[5] , \SB2_0_15/buf_output[4] ,
         \SB2_0_15/buf_output[3] , \SB2_0_15/buf_output[2] ,
         \SB2_0_15/buf_output[1] , \SB2_0_15/buf_output[0] , \SB2_0_15/i3[0] ,
         \SB2_0_15/i1_5 , \SB2_0_15/i1_7 , \SB2_0_15/i1[9] , \SB2_0_15/i0_0 ,
         \SB2_0_15/i0_3 , \SB2_0_15/i0[10] , \SB2_0_15/i0[9] ,
         \SB2_0_15/i0[8] , \SB2_0_15/i0[7] , \SB2_0_15/i0[6] ,
         \SB2_0_16/buf_output[5] , \SB2_0_16/buf_output[4] ,
         \SB2_0_16/buf_output[3] , \SB2_0_16/buf_output[2] ,
         \SB2_0_16/buf_output[1] , \SB2_0_16/buf_output[0] , \SB2_0_16/i3[0] ,
         \SB2_0_16/i1_5 , \SB2_0_16/i1_7 , \SB2_0_16/i1[9] , \SB2_0_16/i0_0 ,
         \SB2_0_16/i0_3 , \SB2_0_16/i0_4 , \SB2_0_16/i0[10] , \SB2_0_16/i0[9] ,
         \SB2_0_16/i0[8] , \SB2_0_16/i0[6] , \SB2_0_17/buf_output[5] ,
         \SB2_0_17/buf_output[4] , \SB2_0_17/buf_output[3] ,
         \SB2_0_17/buf_output[2] , \SB2_0_17/buf_output[1] ,
         \SB2_0_17/buf_output[0] , \SB2_0_17/i3[0] , \SB2_0_17/i1_5 ,
         \SB2_0_17/i1_7 , \SB2_0_17/i1[9] , \SB2_0_17/i0_0 , \SB2_0_17/i0_3 ,
         \SB2_0_17/i0[10] , \SB2_0_17/i0[9] , \SB2_0_17/i0[8] ,
         \SB2_0_17/i0[7] , \SB2_0_17/i0[6] , \SB2_0_18/buf_output[5] ,
         \SB2_0_18/buf_output[4] , \SB2_0_18/buf_output[3] ,
         \SB2_0_18/buf_output[2] , \SB2_0_18/buf_output[1] ,
         \SB2_0_18/buf_output[0] , \SB2_0_18/i3[0] , \SB2_0_18/i1_5 ,
         \SB2_0_18/i1_7 , \SB2_0_18/i1[9] , \SB2_0_18/i0_0 , \SB2_0_18/i0_3 ,
         \SB2_0_18/i0[10] , \SB2_0_18/i0[9] , \SB2_0_18/i0[8] ,
         \SB2_0_18/i0[7] , \SB2_0_18/i0[6] , \SB2_0_19/buf_output[5] ,
         \SB2_0_19/buf_output[4] , \SB2_0_19/buf_output[3] ,
         \SB2_0_19/buf_output[2] , \SB2_0_19/buf_output[1] ,
         \SB2_0_19/buf_output[0] , \SB2_0_19/i3[0] , \SB2_0_19/i1_5 ,
         \SB2_0_19/i1_7 , \SB2_0_19/i1[9] , \SB2_0_19/i0_0 , \SB2_0_19/i0_3 ,
         \SB2_0_19/i0[10] , \SB2_0_19/i0[9] , \SB2_0_19/i0[8] ,
         \SB2_0_19/i0[7] , \SB2_0_19/i0[6] , \SB2_0_20/buf_output[5] ,
         \SB2_0_20/buf_output[4] , \SB2_0_20/buf_output[3] ,
         \SB2_0_20/buf_output[2] , \SB2_0_20/buf_output[1] ,
         \SB2_0_20/buf_output[0] , \SB2_0_20/i3[0] , \SB2_0_20/i1_5 ,
         \SB2_0_20/i1_7 , \SB2_0_20/i1[9] , \SB2_0_20/i0_0 , \SB2_0_20/i0_3 ,
         \SB2_0_20/i0_4 , \SB2_0_20/i0[10] , \SB2_0_20/i0[9] ,
         \SB2_0_20/i0[8] , \SB2_0_20/i0[7] , \SB2_0_20/i0[6] ,
         \SB2_0_21/buf_output[5] , \SB2_0_21/buf_output[4] ,
         \SB2_0_21/buf_output[3] , \SB2_0_21/buf_output[2] ,
         \SB2_0_21/buf_output[1] , \SB2_0_21/buf_output[0] , \SB2_0_21/i3[0] ,
         \SB2_0_21/i1_5 , \SB2_0_21/i1_7 , \SB2_0_21/i1[9] , \SB2_0_21/i0_0 ,
         \SB2_0_21/i0_3 , \SB2_0_21/i0_4 , \SB2_0_21/i0[10] , \SB2_0_21/i0[9] ,
         \SB2_0_21/i0[8] , \SB2_0_21/i0[7] , \SB2_0_21/i0[6] ,
         \SB2_0_22/buf_output[5] , \SB2_0_22/buf_output[4] ,
         \SB2_0_22/buf_output[3] , \SB2_0_22/buf_output[2] ,
         \SB2_0_22/buf_output[1] , \SB2_0_22/buf_output[0] , \SB2_0_22/i3[0] ,
         \SB2_0_22/i1_5 , \SB2_0_22/i1_7 , \SB2_0_22/i1[9] , \SB2_0_22/i0_0 ,
         \SB2_0_22/i0_3 , \SB2_0_22/i0_4 , \SB2_0_22/i0[10] , \SB2_0_22/i0[8] ,
         \SB2_0_22/i0[7] , \SB2_0_22/i0[6] , \SB2_0_23/buf_output[5] ,
         \SB2_0_23/buf_output[4] , \SB2_0_23/buf_output[3] ,
         \SB2_0_23/buf_output[2] , \SB2_0_23/buf_output[1] ,
         \SB2_0_23/buf_output[0] , \SB2_0_23/i3[0] , \SB2_0_23/i1_5 ,
         \SB2_0_23/i1_7 , \SB2_0_23/i1[9] , \SB2_0_23/i0_0 , \SB2_0_23/i0_3 ,
         \SB2_0_23/i0_4 , \SB2_0_23/i0[10] , \SB2_0_23/i0[9] ,
         \SB2_0_23/i0[8] , \SB2_0_23/i0[6] , \SB2_0_24/buf_output[5] ,
         \SB2_0_24/buf_output[4] , \SB2_0_24/buf_output[3] ,
         \SB2_0_24/buf_output[2] , \SB2_0_24/buf_output[1] ,
         \SB2_0_24/buf_output[0] , \SB2_0_24/i3[0] , \SB2_0_24/i1_5 ,
         \SB2_0_24/i1_7 , \SB2_0_24/i1[9] , \SB2_0_24/i0_0 , \SB2_0_24/i0_3 ,
         \SB2_0_24/i0[10] , \SB2_0_24/i0[9] , \SB2_0_24/i0[8] ,
         \SB2_0_24/i0[7] , \SB2_0_25/buf_output[5] , \SB2_0_25/buf_output[4] ,
         \SB2_0_25/buf_output[3] , \SB2_0_25/buf_output[2] ,
         \SB2_0_25/buf_output[1] , \SB2_0_25/buf_output[0] , \SB2_0_25/i3[0] ,
         \SB2_0_25/i1_5 , \SB2_0_25/i1_7 , \SB2_0_25/i1[9] , \SB2_0_25/i0_0 ,
         \SB2_0_25/i0_3 , \SB2_0_25/i0[9] , \SB2_0_25/i0[8] , \SB2_0_25/i0[7] ,
         \SB2_0_26/buf_output[5] , \SB2_0_26/buf_output[4] ,
         \SB2_0_26/buf_output[3] , \SB2_0_26/buf_output[2] ,
         \SB2_0_26/buf_output[1] , \SB2_0_26/buf_output[0] , \SB2_0_26/i3[0] ,
         \SB2_0_26/i1_5 , \SB2_0_26/i1_7 , \SB2_0_26/i1[9] , \SB2_0_26/i0_0 ,
         \SB2_0_26/i0_3 , \SB2_0_26/i0[10] , \SB2_0_26/i0[9] ,
         \SB2_0_26/i0[8] , \SB2_0_26/i0[7] , \SB2_0_26/i0[6] ,
         \SB2_0_27/buf_output[5] , \SB2_0_27/buf_output[4] ,
         \SB2_0_27/buf_output[3] , \SB2_0_27/buf_output[2] ,
         \SB2_0_27/buf_output[1] , \SB2_0_27/buf_output[0] , \SB2_0_27/i3[0] ,
         \SB2_0_27/i1_5 , \SB2_0_27/i1_7 , \SB2_0_27/i1[9] , \SB2_0_27/i0_0 ,
         \SB2_0_27/i0_3 , \SB2_0_27/i0_4 , \SB2_0_27/i0[10] , \SB2_0_27/i0[9] ,
         \SB2_0_27/i0[8] , \SB2_0_27/i0[6] , \SB2_0_28/buf_output[5] ,
         \SB2_0_28/buf_output[4] , \SB2_0_28/buf_output[3] ,
         \SB2_0_28/buf_output[2] , \SB2_0_28/buf_output[1] ,
         \SB2_0_28/buf_output[0] , \SB2_0_28/i3[0] , \SB2_0_28/i1_5 ,
         \SB2_0_28/i1_7 , \SB2_0_28/i1[9] , \SB2_0_28/i0_0 , \SB2_0_28/i0_3 ,
         \SB2_0_28/i0[10] , \SB2_0_28/i0[8] , \SB2_0_28/i0[7] ,
         \SB2_0_28/i0[6] , \SB2_0_29/buf_output[5] , \SB2_0_29/buf_output[4] ,
         \SB2_0_29/buf_output[3] , \SB2_0_29/buf_output[2] ,
         \SB2_0_29/buf_output[1] , \SB2_0_29/buf_output[0] , \SB2_0_29/i3[0] ,
         \SB2_0_29/i1_5 , \SB2_0_29/i1_7 , \SB2_0_29/i1[9] , \SB2_0_29/i0_0 ,
         \SB2_0_29/i0_3 , \SB2_0_29/i0_4 , \SB2_0_29/i0[9] , \SB2_0_29/i0[8] ,
         \SB2_0_29/i0[7] , \SB2_0_29/i0[6] , \SB2_0_30/buf_output[5] ,
         \SB2_0_30/buf_output[4] , \SB2_0_30/buf_output[3] ,
         \SB2_0_30/buf_output[2] , \SB2_0_30/buf_output[1] ,
         \SB2_0_30/buf_output[0] , \SB2_0_30/i3[0] , \SB2_0_30/i1_5 ,
         \SB2_0_30/i1_7 , \SB2_0_30/i1[9] , \SB2_0_30/i0_0 , \SB2_0_30/i0_3 ,
         \SB2_0_30/i0[10] , \SB2_0_30/i0[9] , \SB2_0_30/i0[8] ,
         \SB2_0_30/i0[7] , \SB2_0_30/i0[6] , \SB2_0_31/buf_output[5] ,
         \SB2_0_31/buf_output[4] , \SB2_0_31/buf_output[3] ,
         \SB2_0_31/buf_output[2] , \SB2_0_31/buf_output[1] ,
         \SB2_0_31/buf_output[0] , \SB2_0_31/i3[0] , \SB2_0_31/i1_5 ,
         \SB2_0_31/i1_7 , \SB2_0_31/i1[9] , \SB2_0_31/i0_0 , \SB2_0_31/i0_3 ,
         \SB2_0_31/i0[10] , \SB2_0_31/i0[9] , \SB2_0_31/i0[8] ,
         \SB2_0_31/i0[7] , \SB2_0_31/i0[6] , \SB1_1_0/buf_output[5] ,
         \SB1_1_0/buf_output[3] , \SB1_1_0/buf_output[2] ,
         \SB1_1_0/buf_output[1] , \SB1_1_0/buf_output[0] , \SB1_1_0/i3[0] ,
         \SB1_1_0/i1_5 , \SB1_1_0/i1_7 , \SB1_1_0/i1[9] , \SB1_1_0/i0_0 ,
         \SB1_1_0/i0_3 , \SB1_1_0/i0_4 , \SB1_1_0/i0[10] , \SB1_1_0/i0[9] ,
         \SB1_1_0/i0[8] , \SB1_1_0/i0[7] , \SB1_1_0/i0[6] ,
         \SB1_1_1/buf_output[5] , \SB1_1_1/buf_output[3] ,
         \SB1_1_1/buf_output[2] , \SB1_1_1/buf_output[1] ,
         \SB1_1_1/buf_output[0] , \SB1_1_1/i3[0] , \SB1_1_1/i1_5 ,
         \SB1_1_1/i1_7 , \SB1_1_1/i1[9] , \SB1_1_1/i0_0 , \SB1_1_1/i0_3 ,
         \SB1_1_1/i0_4 , \SB1_1_1/i0[10] , \SB1_1_1/i0[9] , \SB1_1_1/i0[8] ,
         \SB1_1_1/i0[7] , \SB1_1_1/i0[6] , \SB1_1_2/buf_output[5] ,
         \SB1_1_2/buf_output[4] , \SB1_1_2/buf_output[3] ,
         \SB1_1_2/buf_output[2] , \SB1_1_2/buf_output[1] ,
         \SB1_1_2/buf_output[0] , \SB1_1_2/i3[0] , \SB1_1_2/i1_5 ,
         \SB1_1_2/i1_7 , \SB1_1_2/i1[9] , \SB1_1_2/i0_0 , \SB1_1_2/i0_3 ,
         \SB1_1_2/i0_4 , \SB1_1_2/i0[10] , \SB1_1_2/i0[9] , \SB1_1_2/i0[8] ,
         \SB1_1_2/i0[7] , \SB1_1_2/i0[6] , \SB1_1_3/buf_output[5] ,
         \SB1_1_3/buf_output[4] , \SB1_1_3/buf_output[3] ,
         \SB1_1_3/buf_output[2] , \SB1_1_3/buf_output[1] ,
         \SB1_1_3/buf_output[0] , \SB1_1_3/i3[0] , \SB1_1_3/i1_5 ,
         \SB1_1_3/i1_7 , \SB1_1_3/i1[9] , \SB1_1_3/i0_0 , \SB1_1_3/i0_3 ,
         \SB1_1_3/i0_4 , \SB1_1_3/i0[10] , \SB1_1_3/i0[9] , \SB1_1_3/i0[8] ,
         \SB1_1_3/i0[7] , \SB1_1_3/i0[6] , \SB1_1_4/buf_output[5] ,
         \SB1_1_4/buf_output[3] , \SB1_1_4/buf_output[1] ,
         \SB1_1_4/buf_output[0] , \SB1_1_4/i3[0] , \SB1_1_4/i1_5 ,
         \SB1_1_4/i1_7 , \SB1_1_4/i1[9] , \SB1_1_4/i0_0 , \SB1_1_4/i0_3 ,
         \SB1_1_4/i0_4 , \SB1_1_4/i0[10] , \SB1_1_4/i0[9] , \SB1_1_4/i0[8] ,
         \SB1_1_4/i0[7] , \SB1_1_4/i0[6] , \SB1_1_5/buf_output[5] ,
         \SB1_1_5/buf_output[4] , \SB1_1_5/buf_output[3] ,
         \SB1_1_5/buf_output[2] , \SB1_1_5/buf_output[1] ,
         \SB1_1_5/buf_output[0] , \SB1_1_5/i3[0] , \SB1_1_5/i1_5 ,
         \SB1_1_5/i1_7 , \SB1_1_5/i1[9] , \SB1_1_5/i0_0 , \SB1_1_5/i0_3 ,
         \SB1_1_5/i0_4 , \SB1_1_5/i0[10] , \SB1_1_5/i0[9] , \SB1_1_5/i0[8] ,
         \SB1_1_5/i0[7] , \SB1_1_5/i0[6] , \SB1_1_6/buf_output[5] ,
         \SB1_1_6/buf_output[4] , \SB1_1_6/buf_output[3] ,
         \SB1_1_6/buf_output[2] , \SB1_1_6/buf_output[1] ,
         \SB1_1_6/buf_output[0] , \SB1_1_6/i3[0] , \SB1_1_6/i1_5 ,
         \SB1_1_6/i1_7 , \SB1_1_6/i1[9] , \SB1_1_6/i0_0 , \SB1_1_6/i0_3 ,
         \SB1_1_6/i0_4 , \SB1_1_6/i0[10] , \SB1_1_6/i0[9] , \SB1_1_6/i0[8] ,
         \SB1_1_6/i0[7] , \SB1_1_6/i0[6] , \SB1_1_7/buf_output[5] ,
         \SB1_1_7/buf_output[4] , \SB1_1_7/buf_output[3] ,
         \SB1_1_7/buf_output[2] , \SB1_1_7/buf_output[1] ,
         \SB1_1_7/buf_output[0] , \SB1_1_7/i3[0] , \SB1_1_7/i1_5 ,
         \SB1_1_7/i1_7 , \SB1_1_7/i1[9] , \SB1_1_7/i0_0 , \SB1_1_7/i0_3 ,
         \SB1_1_7/i0_4 , \SB1_1_7/i0[10] , \SB1_1_7/i0[9] , \SB1_1_7/i0[8] ,
         \SB1_1_7/i0[7] , \SB1_1_7/i0[6] , \SB1_1_8/buf_output[5] ,
         \SB1_1_8/buf_output[3] , \SB1_1_8/buf_output[2] ,
         \SB1_1_8/buf_output[1] , \SB1_1_8/buf_output[0] , \SB1_1_8/i3[0] ,
         \SB1_1_8/i1_7 , \SB1_1_8/i1[9] , \SB1_1_8/i0_0 , \SB1_1_8/i0_4 ,
         \SB1_1_8/i0[10] , \SB1_1_8/i0[9] , \SB1_1_8/i0[8] , \SB1_1_8/i0[7] ,
         \SB1_1_8/i0[6] , \SB1_1_9/buf_output[5] , \SB1_1_9/buf_output[4] ,
         \SB1_1_9/buf_output[3] , \SB1_1_9/buf_output[2] ,
         \SB1_1_9/buf_output[1] , \SB1_1_9/buf_output[0] , \SB1_1_9/i3[0] ,
         \SB1_1_9/i1_5 , \SB1_1_9/i1_7 , \SB1_1_9/i1[9] , \SB1_1_9/i0_0 ,
         \SB1_1_9/i0_3 , \SB1_1_9/i0_4 , \SB1_1_9/i0[10] , \SB1_1_9/i0[9] ,
         \SB1_1_9/i0[8] , \SB1_1_9/i0[7] , \SB1_1_9/i0[6] ,
         \SB1_1_10/buf_output[5] , \SB1_1_10/buf_output[4] ,
         \SB1_1_10/buf_output[3] , \SB1_1_10/buf_output[2] ,
         \SB1_1_10/buf_output[1] , \SB1_1_10/buf_output[0] , \SB1_1_10/i3[0] ,
         \SB1_1_10/i1_5 , \SB1_1_10/i1_7 , \SB1_1_10/i1[9] , \SB1_1_10/i0_0 ,
         \SB1_1_10/i0_3 , \SB1_1_10/i0_4 , \SB1_1_10/i0[10] , \SB1_1_10/i0[9] ,
         \SB1_1_10/i0[8] , \SB1_1_10/i0[7] , \SB1_1_10/i0[6] ,
         \SB1_1_11/buf_output[5] , \SB1_1_11/buf_output[4] ,
         \SB1_1_11/buf_output[3] , \SB1_1_11/buf_output[2] ,
         \SB1_1_11/buf_output[1] , \SB1_1_11/buf_output[0] , \SB1_1_11/i3[0] ,
         \SB1_1_11/i1_5 , \SB1_1_11/i1_7 , \SB1_1_11/i1[9] , \SB1_1_11/i0_0 ,
         \SB1_1_11/i0_3 , \SB1_1_11/i0_4 , \SB1_1_11/i0[10] , \SB1_1_11/i0[9] ,
         \SB1_1_11/i0[8] , \SB1_1_11/i0[7] , \SB1_1_11/i0[6] ,
         \SB1_1_12/buf_output[5] , \SB1_1_12/buf_output[4] ,
         \SB1_1_12/buf_output[3] , \SB1_1_12/buf_output[2] ,
         \SB1_1_12/buf_output[1] , \SB1_1_12/buf_output[0] , \SB1_1_12/i3[0] ,
         \SB1_1_12/i1_5 , \SB1_1_12/i1_7 , \SB1_1_12/i1[9] , \SB1_1_12/i0_0 ,
         \SB1_1_12/i0_3 , \SB1_1_12/i0_4 , \SB1_1_12/i0[10] , \SB1_1_12/i0[9] ,
         \SB1_1_12/i0[8] , \SB1_1_12/i0[7] , \SB1_1_12/i0[6] ,
         \SB1_1_13/buf_output[5] , \SB1_1_13/buf_output[4] ,
         \SB1_1_13/buf_output[3] , \SB1_1_13/buf_output[2] ,
         \SB1_1_13/buf_output[1] , \SB1_1_13/buf_output[0] , \SB1_1_13/i3[0] ,
         \SB1_1_13/i1_5 , \SB1_1_13/i1_7 , \SB1_1_13/i1[9] , \SB1_1_13/i0_0 ,
         \SB1_1_13/i0_3 , \SB1_1_13/i0_4 , \SB1_1_13/i0[10] , \SB1_1_13/i0[9] ,
         \SB1_1_13/i0[8] , \SB1_1_13/i0[7] , \SB1_1_13/i0[6] ,
         \SB1_1_14/buf_output[5] , \SB1_1_14/buf_output[4] ,
         \SB1_1_14/buf_output[3] , \SB1_1_14/buf_output[2] ,
         \SB1_1_14/buf_output[1] , \SB1_1_14/buf_output[0] , \SB1_1_14/i3[0] ,
         \SB1_1_14/i1_5 , \SB1_1_14/i1_7 , \SB1_1_14/i1[9] , \SB1_1_14/i0_0 ,
         \SB1_1_14/i0_3 , \SB1_1_14/i0_4 , \SB1_1_14/i0[10] , \SB1_1_14/i0[9] ,
         \SB1_1_14/i0[8] , \SB1_1_14/i0[7] , \SB1_1_14/i0[6] ,
         \SB1_1_15/buf_output[5] , \SB1_1_15/buf_output[4] ,
         \SB1_1_15/buf_output[3] , \SB1_1_15/buf_output[2] ,
         \SB1_1_15/buf_output[1] , \SB1_1_15/buf_output[0] , \SB1_1_15/i3[0] ,
         \SB1_1_15/i1_5 , \SB1_1_15/i1_7 , \SB1_1_15/i1[9] , \SB1_1_15/i0_0 ,
         \SB1_1_15/i0_3 , \SB1_1_15/i0_4 , \SB1_1_15/i0[10] , \SB1_1_15/i0[9] ,
         \SB1_1_15/i0[8] , \SB1_1_15/i0[7] , \SB1_1_15/i0[6] ,
         \SB1_1_16/buf_output[5] , \SB1_1_16/buf_output[3] ,
         \SB1_1_16/buf_output[1] , \SB1_1_16/buf_output[0] , \SB1_1_16/i3[0] ,
         \SB1_1_16/i1_5 , \SB1_1_16/i1_7 , \SB1_1_16/i1[9] , \SB1_1_16/i0_0 ,
         \SB1_1_16/i0_3 , \SB1_1_16/i0_4 , \SB1_1_16/i0[10] , \SB1_1_16/i0[9] ,
         \SB1_1_16/i0[8] , \SB1_1_16/i0[7] , \SB1_1_16/i0[6] ,
         \SB1_1_17/buf_output[5] , \SB1_1_17/buf_output[4] ,
         \SB1_1_17/buf_output[3] , \SB1_1_17/buf_output[2] ,
         \SB1_1_17/buf_output[1] , \SB1_1_17/buf_output[0] , \SB1_1_17/i3[0] ,
         \SB1_1_17/i1_5 , \SB1_1_17/i1_7 , \SB1_1_17/i1[9] , \SB1_1_17/i0_0 ,
         \SB1_1_17/i0_3 , \SB1_1_17/i0_4 , \SB1_1_17/i0[10] , \SB1_1_17/i0[9] ,
         \SB1_1_17/i0[8] , \SB1_1_17/i0[7] , \SB1_1_17/i0[6] ,
         \SB1_1_18/buf_output[5] , \SB1_1_18/buf_output[4] ,
         \SB1_1_18/buf_output[3] , \SB1_1_18/buf_output[2] ,
         \SB1_1_18/buf_output[1] , \SB1_1_18/buf_output[0] , \SB1_1_18/i3[0] ,
         \SB1_1_18/i1_5 , \SB1_1_18/i1_7 , \SB1_1_18/i1[9] , \SB1_1_18/i0_0 ,
         \SB1_1_18/i0_3 , \SB1_1_18/i0_4 , \SB1_1_18/i0[10] , \SB1_1_18/i0[9] ,
         \SB1_1_18/i0[8] , \SB1_1_18/i0[7] , \SB1_1_18/i0[6] ,
         \SB1_1_19/buf_output[5] , \SB1_1_19/buf_output[4] ,
         \SB1_1_19/buf_output[3] , \SB1_1_19/buf_output[2] ,
         \SB1_1_19/buf_output[1] , \SB1_1_19/buf_output[0] , \SB1_1_19/i3[0] ,
         \SB1_1_19/i1_5 , \SB1_1_19/i1_7 , \SB1_1_19/i1[9] , \SB1_1_19/i0_0 ,
         \SB1_1_19/i0_3 , \SB1_1_19/i0_4 , \SB1_1_19/i0[10] , \SB1_1_19/i0[9] ,
         \SB1_1_19/i0[8] , \SB1_1_19/i0[7] , \SB1_1_19/i0[6] ,
         \SB1_1_20/buf_output[5] , \SB1_1_20/buf_output[3] ,
         \SB1_1_20/buf_output[2] , \SB1_1_20/buf_output[1] ,
         \SB1_1_20/buf_output[0] , \SB1_1_20/i3[0] , \SB1_1_20/i1_5 ,
         \SB1_1_20/i1_7 , \SB1_1_20/i1[9] , \SB1_1_20/i0_0 , \SB1_1_20/i0_3 ,
         \SB1_1_20/i0_4 , \SB1_1_20/i0[10] , \SB1_1_20/i0[9] ,
         \SB1_1_20/i0[8] , \SB1_1_20/i0[7] , \SB1_1_20/i0[6] ,
         \SB1_1_21/buf_output[5] , \SB1_1_21/buf_output[4] ,
         \SB1_1_21/buf_output[3] , \SB1_1_21/buf_output[2] ,
         \SB1_1_21/buf_output[1] , \SB1_1_21/buf_output[0] , \SB1_1_21/i3[0] ,
         \SB1_1_21/i1_5 , \SB1_1_21/i1_7 , \SB1_1_21/i1[9] , \SB1_1_21/i0_0 ,
         \SB1_1_21/i0_3 , \SB1_1_21/i0_4 , \SB1_1_21/i0[10] , \SB1_1_21/i0[9] ,
         \SB1_1_21/i0[8] , \SB1_1_21/i0[7] , \SB1_1_21/i0[6] ,
         \SB1_1_22/buf_output[5] , \SB1_1_22/buf_output[4] ,
         \SB1_1_22/buf_output[3] , \SB1_1_22/buf_output[2] ,
         \SB1_1_22/buf_output[1] , \SB1_1_22/buf_output[0] , \SB1_1_22/i3[0] ,
         \SB1_1_22/i1_5 , \SB1_1_22/i1_7 , \SB1_1_22/i1[9] , \SB1_1_22/i0_0 ,
         \SB1_1_22/i0_4 , \SB1_1_22/i0[10] , \SB1_1_22/i0[9] ,
         \SB1_1_22/i0[8] , \SB1_1_22/i0[7] , \SB1_1_22/i0[6] ,
         \SB1_1_23/buf_output[5] , \SB1_1_23/buf_output[4] ,
         \SB1_1_23/buf_output[3] , \SB1_1_23/buf_output[2] ,
         \SB1_1_23/buf_output[1] , \SB1_1_23/buf_output[0] , \SB1_1_23/i3[0] ,
         \SB1_1_23/i1_5 , \SB1_1_23/i1_7 , \SB1_1_23/i1[9] , \SB1_1_23/i0_0 ,
         \SB1_1_23/i0_3 , \SB1_1_23/i0_4 , \SB1_1_23/i0[10] , \SB1_1_23/i0[9] ,
         \SB1_1_23/i0[8] , \SB1_1_23/i0[7] , \SB1_1_23/i0[6] ,
         \SB1_1_24/buf_output[5] , \SB1_1_24/buf_output[4] ,
         \SB1_1_24/buf_output[3] , \SB1_1_24/buf_output[2] ,
         \SB1_1_24/buf_output[1] , \SB1_1_24/buf_output[0] , \SB1_1_24/i3[0] ,
         \SB1_1_24/i1_5 , \SB1_1_24/i1_7 , \SB1_1_24/i1[9] , \SB1_1_24/i0_0 ,
         \SB1_1_24/i0_3 , \SB1_1_24/i0_4 , \SB1_1_24/i0[10] , \SB1_1_24/i0[9] ,
         \SB1_1_24/i0[8] , \SB1_1_24/i0[7] , \SB1_1_24/i0[6] ,
         \SB1_1_25/buf_output[5] , \SB1_1_25/buf_output[4] ,
         \SB1_1_25/buf_output[3] , \SB1_1_25/buf_output[2] ,
         \SB1_1_25/buf_output[1] , \SB1_1_25/buf_output[0] , \SB1_1_25/i3[0] ,
         \SB1_1_25/i1_5 , \SB1_1_25/i1_7 , \SB1_1_25/i1[9] , \SB1_1_25/i0_0 ,
         \SB1_1_25/i0_3 , \SB1_1_25/i0_4 , \SB1_1_25/i0[10] , \SB1_1_25/i0[9] ,
         \SB1_1_25/i0[8] , \SB1_1_25/i0[7] , \SB1_1_25/i0[6] ,
         \SB1_1_26/buf_output[5] , \SB1_1_26/buf_output[4] ,
         \SB1_1_26/buf_output[3] , \SB1_1_26/buf_output[2] ,
         \SB1_1_26/buf_output[1] , \SB1_1_26/i3[0] , \SB1_1_26/i1_5 ,
         \SB1_1_26/i1_7 , \SB1_1_26/i1[9] , \SB1_1_26/i0_0 , \SB1_1_26/i0_3 ,
         \SB1_1_26/i0_4 , \SB1_1_26/i0[10] , \SB1_1_26/i0[9] ,
         \SB1_1_26/i0[8] , \SB1_1_26/i0[7] , \SB1_1_26/i0[6] ,
         \SB1_1_27/buf_output[5] , \SB1_1_27/buf_output[4] ,
         \SB1_1_27/buf_output[3] , \SB1_1_27/buf_output[2] ,
         \SB1_1_27/buf_output[1] , \SB1_1_27/buf_output[0] , \SB1_1_27/i3[0] ,
         \SB1_1_27/i1_5 , \SB1_1_27/i1_7 , \SB1_1_27/i1[9] , \SB1_1_27/i0_0 ,
         \SB1_1_27/i0_3 , \SB1_1_27/i0_4 , \SB1_1_27/i0[10] , \SB1_1_27/i0[9] ,
         \SB1_1_27/i0[8] , \SB1_1_27/i0[7] , \SB1_1_27/i0[6] ,
         \SB1_1_28/buf_output[5] , \SB1_1_28/buf_output[4] ,
         \SB1_1_28/buf_output[3] , \SB1_1_28/buf_output[2] ,
         \SB1_1_28/buf_output[1] , \SB1_1_28/buf_output[0] , \SB1_1_28/i3[0] ,
         \SB1_1_28/i1_5 , \SB1_1_28/i1_7 , \SB1_1_28/i1[9] , \SB1_1_28/i0_0 ,
         \SB1_1_28/i0_3 , \SB1_1_28/i0_4 , \SB1_1_28/i0[10] , \SB1_1_28/i0[9] ,
         \SB1_1_28/i0[8] , \SB1_1_28/i0[7] , \SB1_1_28/i0[6] ,
         \SB1_1_29/buf_output[5] , \SB1_1_29/buf_output[4] ,
         \SB1_1_29/buf_output[3] , \SB1_1_29/buf_output[2] ,
         \SB1_1_29/buf_output[1] , \SB1_1_29/buf_output[0] , \SB1_1_29/i3[0] ,
         \SB1_1_29/i1_5 , \SB1_1_29/i1_7 , \SB1_1_29/i1[9] , \SB1_1_29/i0_0 ,
         \SB1_1_29/i0_3 , \SB1_1_29/i0_4 , \SB1_1_29/i0[10] , \SB1_1_29/i0[9] ,
         \SB1_1_29/i0[8] , \SB1_1_29/i0[7] , \SB1_1_29/i0[6] ,
         \SB1_1_30/buf_output[5] , \SB1_1_30/buf_output[3] ,
         \SB1_1_30/buf_output[2] , \SB1_1_30/buf_output[1] ,
         \SB1_1_30/buf_output[0] , \SB1_1_30/i3[0] , \SB1_1_30/i1_5 ,
         \SB1_1_30/i1_7 , \SB1_1_30/i1[9] , \SB1_1_30/i0_0 , \SB1_1_30/i0_3 ,
         \SB1_1_30/i0_4 , \SB1_1_30/i0[10] , \SB1_1_30/i0[9] ,
         \SB1_1_30/i0[8] , \SB1_1_30/i0[7] , \SB1_1_30/i0[6] ,
         \SB1_1_31/buf_output[5] , \SB1_1_31/buf_output[3] ,
         \SB1_1_31/buf_output[2] , \SB1_1_31/buf_output[1] ,
         \SB1_1_31/buf_output[0] , \SB1_1_31/i3[0] , \SB1_1_31/i1_5 ,
         \SB1_1_31/i1_7 , \SB1_1_31/i1[9] , \SB1_1_31/i0_0 , \SB1_1_31/i0_3 ,
         \SB1_1_31/i0_4 , \SB1_1_31/i0[10] , \SB1_1_31/i0[9] ,
         \SB1_1_31/i0[8] , \SB1_1_31/i0[7] , \SB1_1_31/i0[6] ,
         \SB2_1_0/buf_output[5] , \SB2_1_0/buf_output[4] ,
         \SB2_1_0/buf_output[3] , \SB2_1_0/buf_output[2] ,
         \SB2_1_0/buf_output[1] , \SB2_1_0/buf_output[0] , \SB2_1_0/i3[0] ,
         \SB2_1_0/i1_5 , \SB2_1_0/i1_7 , \SB2_1_0/i1[9] , \SB2_1_0/i0_0 ,
         \SB2_1_0/i0_3 , \SB2_1_0/i0[10] , \SB2_1_0/i0[9] , \SB2_1_0/i0[8] ,
         \SB2_1_0/i0[7] , \SB2_1_0/i0[6] , \SB2_1_1/buf_output[5] ,
         \SB2_1_1/buf_output[4] , \SB2_1_1/buf_output[3] ,
         \SB2_1_1/buf_output[2] , \SB2_1_1/buf_output[1] ,
         \SB2_1_1/buf_output[0] , \SB2_1_1/i3[0] , \SB2_1_1/i1_5 ,
         \SB2_1_1/i1_7 , \SB2_1_1/i1[9] , \SB2_1_1/i0_0 , \SB2_1_1/i0_3 ,
         \SB2_1_1/i0_4 , \SB2_1_1/i0[10] , \SB2_1_1/i0[9] , \SB2_1_1/i0[8] ,
         \SB2_1_1/i0[7] , \SB2_1_1/i0[6] , \SB2_1_2/buf_output[5] ,
         \SB2_1_2/buf_output[4] , \SB2_1_2/buf_output[3] ,
         \SB2_1_2/buf_output[2] , \SB2_1_2/buf_output[1] ,
         \SB2_1_2/buf_output[0] , \SB2_1_2/i3[0] , \SB2_1_2/i1_5 ,
         \SB2_1_2/i1_7 , \SB2_1_2/i1[9] , \SB2_1_2/i0_0 , \SB2_1_2/i0_3 ,
         \SB2_1_2/i0_4 , \SB2_1_2/i0[10] , \SB2_1_2/i0[9] , \SB2_1_2/i0[8] ,
         \SB2_1_2/i0[7] , \SB2_1_2/i0[6] , \SB2_1_3/buf_output[5] ,
         \SB2_1_3/buf_output[4] , \SB2_1_3/buf_output[3] ,
         \SB2_1_3/buf_output[2] , \SB2_1_3/buf_output[1] ,
         \SB2_1_3/buf_output[0] , \SB2_1_3/i3[0] , \SB2_1_3/i1_5 ,
         \SB2_1_3/i1_7 , \SB2_1_3/i1[9] , \SB2_1_3/i0_0 , \SB2_1_3/i0_3 ,
         \SB2_1_3/i0_4 , \SB2_1_3/i0[10] , \SB2_1_3/i0[9] , \SB2_1_3/i0[8] ,
         \SB2_1_3/i0[7] , \SB2_1_3/i0[6] , \SB2_1_4/buf_output[5] ,
         \SB2_1_4/buf_output[4] , \SB2_1_4/buf_output[3] ,
         \SB2_1_4/buf_output[2] , \SB2_1_4/buf_output[1] ,
         \SB2_1_4/buf_output[0] , \SB2_1_4/i3[0] , \SB2_1_4/i1_5 ,
         \SB2_1_4/i1_7 , \SB2_1_4/i0_3 , \SB2_1_4/i0[10] , \SB2_1_4/i0[9] ,
         \SB2_1_4/i0[8] , \SB2_1_4/i0[7] , \SB2_1_4/i0[6] ,
         \SB2_1_5/buf_output[5] , \SB2_1_5/buf_output[4] ,
         \SB2_1_5/buf_output[2] , \SB2_1_5/buf_output[1] ,
         \SB2_1_5/buf_output[0] , \SB2_1_5/i3[0] , \SB2_1_5/i1_5 ,
         \SB2_1_5/i1_7 , \SB2_1_5/i1[9] , \SB2_1_5/i0_0 , \SB2_1_5/i0_3 ,
         \SB2_1_5/i0[10] , \SB2_1_5/i0[9] , \SB2_1_5/i0[8] , \SB2_1_5/i0[6] ,
         \SB2_1_6/buf_output[5] , \SB2_1_6/buf_output[4] ,
         \SB2_1_6/buf_output[3] , \SB2_1_6/buf_output[2] ,
         \SB2_1_6/buf_output[1] , \SB2_1_6/buf_output[0] , \SB2_1_6/i3[0] ,
         \SB2_1_6/i1_5 , \SB2_1_6/i1_7 , \SB2_1_6/i1[9] , \SB2_1_6/i0_0 ,
         \SB2_1_6/i0_3 , \SB2_1_6/i0_4 , \SB2_1_6/i0[10] , \SB2_1_6/i0[9] ,
         \SB2_1_6/i0[8] , \SB2_1_6/i0[7] , \SB2_1_6/i0[6] ,
         \SB2_1_7/buf_output[5] , \SB2_1_7/buf_output[4] ,
         \SB2_1_7/buf_output[3] , \SB2_1_7/buf_output[2] ,
         \SB2_1_7/buf_output[1] , \SB2_1_7/buf_output[0] , \SB2_1_7/i3[0] ,
         \SB2_1_7/i1_5 , \SB2_1_7/i1_7 , \SB2_1_7/i1[9] , \SB2_1_7/i0_0 ,
         \SB2_1_7/i0_3 , \SB2_1_7/i0_4 , \SB2_1_7/i0[10] , \SB2_1_7/i0[9] ,
         \SB2_1_7/i0[8] , \SB2_1_7/i0[7] , \SB2_1_8/buf_output[5] ,
         \SB2_1_8/buf_output[4] , \SB2_1_8/buf_output[3] ,
         \SB2_1_8/buf_output[2] , \SB2_1_8/buf_output[0] , \SB2_1_8/i3[0] ,
         \SB2_1_8/i1_5 , \SB2_1_8/i1_7 , \SB2_1_8/i1[9] , \SB2_1_8/i0_0 ,
         \SB2_1_8/i0_3 , \SB2_1_8/i0_4 , \SB2_1_8/i0[10] , \SB2_1_8/i0[8] ,
         \SB2_1_8/i0[7] , \SB2_1_8/i0[6] , \SB2_1_9/buf_output[5] ,
         \SB2_1_9/buf_output[4] , \SB2_1_9/buf_output[2] ,
         \SB2_1_9/buf_output[1] , \SB2_1_9/buf_output[0] , \SB2_1_9/i3[0] ,
         \SB2_1_9/i1_5 , \SB2_1_9/i1_7 , \SB2_1_9/i1[9] , \SB2_1_9/i0_0 ,
         \SB2_1_9/i0_3 , \SB2_1_9/i0_4 , \SB2_1_9/i0[10] , \SB2_1_9/i0[9] ,
         \SB2_1_9/i0[8] , \SB2_1_9/i0[7] , \SB2_1_9/i0[6] ,
         \SB2_1_10/buf_output[5] , \SB2_1_10/buf_output[4] ,
         \SB2_1_10/buf_output[3] , \SB2_1_10/buf_output[2] ,
         \SB2_1_10/buf_output[1] , \SB2_1_10/buf_output[0] , \SB2_1_10/i3[0] ,
         \SB2_1_10/i1_5 , \SB2_1_10/i1_7 , \SB2_1_10/i1[9] , \SB2_1_10/i0_0 ,
         \SB2_1_10/i0_3 , \SB2_1_10/i0[10] , \SB2_1_10/i0[9] ,
         \SB2_1_10/i0[8] , \SB2_1_10/i0[7] , \SB2_1_10/i0[6] ,
         \SB2_1_11/buf_output[5] , \SB2_1_11/buf_output[4] ,
         \SB2_1_11/buf_output[3] , \SB2_1_11/buf_output[2] ,
         \SB2_1_11/buf_output[1] , \SB2_1_11/buf_output[0] , \SB2_1_11/i3[0] ,
         \SB2_1_11/i1_5 , \SB2_1_11/i1_7 , \SB2_1_11/i1[9] , \SB2_1_11/i0_0 ,
         \SB2_1_11/i0_3 , \SB2_1_11/i0[10] , \SB2_1_11/i0[9] ,
         \SB2_1_11/i0[8] , \SB2_1_11/i0[7] , \SB2_1_11/i0[6] ,
         \SB2_1_12/buf_output[5] , \SB2_1_12/buf_output[4] ,
         \SB2_1_12/buf_output[3] , \SB2_1_12/buf_output[2] ,
         \SB2_1_12/buf_output[1] , \SB2_1_12/buf_output[0] , \SB2_1_12/i3[0] ,
         \SB2_1_12/i1_5 , \SB2_1_12/i1_7 , \SB2_1_12/i1[9] , \SB2_1_12/i0_0 ,
         \SB2_1_12/i0_3 , \SB2_1_12/i0_4 , \SB2_1_12/i0[10] , \SB2_1_12/i0[9] ,
         \SB2_1_12/i0[8] , \SB2_1_12/i0[7] , \SB2_1_12/i0[6] ,
         \SB2_1_13/buf_output[5] , \SB2_1_13/buf_output[4] ,
         \SB2_1_13/buf_output[3] , \SB2_1_13/buf_output[2] ,
         \SB2_1_13/buf_output[1] , \SB2_1_13/buf_output[0] , \SB2_1_13/i1_5 ,
         \SB2_1_13/i1_7 , \SB2_1_13/i1[9] , \SB2_1_13/i0_0 , \SB2_1_13/i0_3 ,
         \SB2_1_13/i0_4 , \SB2_1_13/i0[10] , \SB2_1_13/i0[8] ,
         \SB2_1_13/i0[7] , \SB2_1_13/i0[6] , \SB2_1_14/buf_output[5] ,
         \SB2_1_14/buf_output[4] , \SB2_1_14/buf_output[3] ,
         \SB2_1_14/buf_output[2] , \SB2_1_14/buf_output[1] ,
         \SB2_1_14/buf_output[0] , \SB2_1_14/i3[0] , \SB2_1_14/i1_5 ,
         \SB2_1_14/i1_7 , \SB2_1_14/i1[9] , \SB2_1_14/i0_0 , \SB2_1_14/i0_3 ,
         \SB2_1_14/i0_4 , \SB2_1_14/i0[10] , \SB2_1_14/i0[9] ,
         \SB2_1_14/i0[8] , \SB2_1_14/i0[7] , \SB2_1_14/i0[6] ,
         \SB2_1_15/buf_output[5] , \SB2_1_15/buf_output[4] ,
         \SB2_1_15/buf_output[3] , \SB2_1_15/buf_output[2] ,
         \SB2_1_15/buf_output[1] , \SB2_1_15/buf_output[0] , \SB2_1_15/i3[0] ,
         \SB2_1_15/i1_5 , \SB2_1_15/i1_7 , \SB2_1_15/i1[9] , \SB2_1_15/i0_0 ,
         \SB2_1_15/i0_3 , \SB2_1_15/i0_4 , \SB2_1_15/i0[10] , \SB2_1_15/i0[9] ,
         \SB2_1_15/i0[8] , \SB2_1_15/i0[6] , \SB2_1_16/buf_output[5] ,
         \SB2_1_16/buf_output[4] , \SB2_1_16/buf_output[3] ,
         \SB2_1_16/buf_output[2] , \SB2_1_16/buf_output[1] ,
         \SB2_1_16/buf_output[0] , \SB2_1_16/i3[0] , \SB2_1_16/i1_5 ,
         \SB2_1_16/i1_7 , \SB2_1_16/i1[9] , \SB2_1_16/i0_0 , \SB2_1_16/i0_3 ,
         \SB2_1_16/i0_4 , \SB2_1_16/i0[10] , \SB2_1_16/i0[9] ,
         \SB2_1_16/i0[8] , \SB2_1_16/i0[7] , \SB2_1_16/i0[6] ,
         \SB2_1_17/buf_output[5] , \SB2_1_17/buf_output[4] ,
         \SB2_1_17/buf_output[3] , \SB2_1_17/buf_output[2] ,
         \SB2_1_17/buf_output[1] , \SB2_1_17/buf_output[0] , \SB2_1_17/i3[0] ,
         \SB2_1_17/i1_5 , \SB2_1_17/i1_7 , \SB2_1_17/i1[9] , \SB2_1_17/i0_0 ,
         \SB2_1_17/i0_3 , \SB2_1_17/i0_4 , \SB2_1_17/i0[10] , \SB2_1_17/i0[9] ,
         \SB2_1_17/i0[8] , \SB2_1_17/i0[7] , \SB2_1_17/i0[6] ,
         \SB2_1_18/buf_output[5] , \SB2_1_18/buf_output[4] ,
         \SB2_1_18/buf_output[3] , \SB2_1_18/buf_output[2] ,
         \SB2_1_18/buf_output[1] , \SB2_1_18/buf_output[0] , \SB2_1_18/i3[0] ,
         \SB2_1_18/i1_5 , \SB2_1_18/i1_7 , \SB2_1_18/i1[9] , \SB2_1_18/i0_0 ,
         \SB2_1_18/i0_3 , \SB2_1_18/i0_4 , \SB2_1_18/i0[10] , \SB2_1_18/i0[9] ,
         \SB2_1_18/i0[8] , \SB2_1_19/buf_output[5] , \SB2_1_19/buf_output[4] ,
         \SB2_1_19/buf_output[3] , \SB2_1_19/buf_output[2] ,
         \SB2_1_19/buf_output[1] , \SB2_1_19/buf_output[0] , \SB2_1_19/i3[0] ,
         \SB2_1_19/i1_5 , \SB2_1_19/i1_7 , \SB2_1_19/i0_3 , \SB2_1_19/i0[10] ,
         \SB2_1_19/i0[9] , \SB2_1_19/i0[8] , \SB2_1_19/i0[6] ,
         \SB2_1_20/buf_output[5] , \SB2_1_20/buf_output[4] ,
         \SB2_1_20/buf_output[3] , \SB2_1_20/buf_output[2] ,
         \SB2_1_20/buf_output[1] , \SB2_1_20/buf_output[0] , \SB2_1_20/i3[0] ,
         \SB2_1_20/i1_5 , \SB2_1_20/i1_7 , \SB2_1_20/i1[9] , \SB2_1_20/i0_0 ,
         \SB2_1_20/i0_3 , \SB2_1_20/i0_4 , \SB2_1_20/i0[10] , \SB2_1_20/i0[9] ,
         \SB2_1_20/i0[8] , \SB2_1_20/i0[7] , \SB2_1_20/i0[6] ,
         \SB2_1_21/buf_output[5] , \SB2_1_21/buf_output[4] ,
         \SB2_1_21/buf_output[3] , \SB2_1_21/buf_output[2] ,
         \SB2_1_21/buf_output[1] , \SB2_1_21/buf_output[0] , \SB2_1_21/i3[0] ,
         \SB2_1_21/i1_5 , \SB2_1_21/i1_7 , \SB2_1_21/i1[9] , \SB2_1_21/i0_0 ,
         \SB2_1_21/i0_3 , \SB2_1_21/i0_4 , \SB2_1_21/i0[10] , \SB2_1_21/i0[8] ,
         \SB2_1_21/i0[7] , \SB2_1_21/i0[6] , \SB2_1_22/buf_output[5] ,
         \SB2_1_22/buf_output[4] , \SB2_1_22/buf_output[3] ,
         \SB2_1_22/buf_output[2] , \SB2_1_22/buf_output[1] ,
         \SB2_1_22/buf_output[0] , \SB2_1_22/i3[0] , \SB2_1_22/i1_5 ,
         \SB2_1_22/i1_7 , \SB2_1_22/i1[9] , \SB2_1_22/i0_0 , \SB2_1_22/i0_3 ,
         \SB2_1_22/i0_4 , \SB2_1_22/i0[10] , \SB2_1_22/i0[9] ,
         \SB2_1_22/i0[8] , \SB2_1_22/i0[7] , \SB2_1_22/i0[6] ,
         \SB2_1_23/buf_output[5] , \SB2_1_23/buf_output[4] ,
         \SB2_1_23/buf_output[3] , \SB2_1_23/buf_output[2] ,
         \SB2_1_23/buf_output[1] , \SB2_1_23/buf_output[0] , \SB2_1_23/i3[0] ,
         \SB2_1_23/i1_5 , \SB2_1_23/i1_7 , \SB2_1_23/i1[9] , \SB2_1_23/i0_0 ,
         \SB2_1_23/i0_3 , \SB2_1_23/i0_4 , \SB2_1_23/i0[10] , \SB2_1_23/i0[9] ,
         \SB2_1_23/i0[8] , \SB2_1_23/i0[7] , \SB2_1_23/i0[6] ,
         \SB2_1_24/buf_output[5] , \SB2_1_24/buf_output[4] ,
         \SB2_1_24/buf_output[3] , \SB2_1_24/buf_output[2] ,
         \SB2_1_24/buf_output[1] , \SB2_1_24/buf_output[0] , \SB2_1_24/i3[0] ,
         \SB2_1_24/i1_5 , \SB2_1_24/i1_7 , \SB2_1_24/i1[9] , \SB2_1_24/i0_0 ,
         \SB2_1_24/i0_3 , \SB2_1_24/i0_4 , \SB2_1_24/i0[10] , \SB2_1_24/i0[9] ,
         \SB2_1_24/i0[8] , \SB2_1_24/i0[7] , \SB2_1_24/i0[6] ,
         \SB2_1_25/buf_output[5] , \SB2_1_25/buf_output[4] ,
         \SB2_1_25/buf_output[3] , \SB2_1_25/buf_output[2] ,
         \SB2_1_25/buf_output[1] , \SB2_1_25/buf_output[0] , \SB2_1_25/i3[0] ,
         \SB2_1_25/i1_5 , \SB2_1_25/i1_7 , \SB2_1_25/i1[9] , \SB2_1_25/i0_0 ,
         \SB2_1_25/i0_3 , \SB2_1_25/i0[10] , \SB2_1_25/i0[9] ,
         \SB2_1_25/i0[8] , \SB2_1_25/i0[7] , \SB2_1_25/i0[6] ,
         \SB2_1_26/buf_output[5] , \SB2_1_26/buf_output[4] ,
         \SB2_1_26/buf_output[3] , \SB2_1_26/buf_output[2] ,
         \SB2_1_26/buf_output[1] , \SB2_1_26/buf_output[0] , \SB2_1_26/i3[0] ,
         \SB2_1_26/i1_5 , \SB2_1_26/i1_7 , \SB2_1_26/i1[9] , \SB2_1_26/i0_0 ,
         \SB2_1_26/i0_3 , \SB2_1_26/i0_4 , \SB2_1_26/i0[10] , \SB2_1_26/i0[9] ,
         \SB2_1_26/i0[8] , \SB2_1_26/i0[7] , \SB2_1_26/i0[6] ,
         \SB2_1_27/buf_output[5] , \SB2_1_27/buf_output[4] ,
         \SB2_1_27/buf_output[3] , \SB2_1_27/buf_output[2] ,
         \SB2_1_27/buf_output[1] , \SB2_1_27/buf_output[0] , \SB2_1_27/i3[0] ,
         \SB2_1_27/i1_5 , \SB2_1_27/i1_7 , \SB2_1_27/i1[9] , \SB2_1_27/i0_0 ,
         \SB2_1_27/i0_3 , \SB2_1_27/i0_4 , \SB2_1_27/i0[10] , \SB2_1_27/i0[9] ,
         \SB2_1_27/i0[8] , \SB2_1_27/i0[7] , \SB2_1_27/i0[6] ,
         \SB2_1_28/buf_output[5] , \SB2_1_28/buf_output[4] ,
         \SB2_1_28/buf_output[3] , \SB2_1_28/buf_output[2] ,
         \SB2_1_28/buf_output[1] , \SB2_1_28/buf_output[0] , \SB2_1_28/i3[0] ,
         \SB2_1_28/i1_5 , \SB2_1_28/i1_7 , \SB2_1_28/i1[9] , \SB2_1_28/i0_0 ,
         \SB2_1_28/i0_3 , \SB2_1_28/i0_4 , \SB2_1_28/i0[10] , \SB2_1_28/i0[9] ,
         \SB2_1_28/i0[8] , \SB2_1_28/i0[7] , \SB2_1_28/i0[6] ,
         \SB2_1_29/buf_output[5] , \SB2_1_29/buf_output[4] ,
         \SB2_1_29/buf_output[3] , \SB2_1_29/buf_output[2] ,
         \SB2_1_29/buf_output[1] , \SB2_1_29/buf_output[0] , \SB2_1_29/i3[0] ,
         \SB2_1_29/i1_5 , \SB2_1_29/i1_7 , \SB2_1_29/i1[9] , \SB2_1_29/i0_0 ,
         \SB2_1_29/i0_3 , \SB2_1_29/i0_4 , \SB2_1_29/i0[10] , \SB2_1_29/i0[9] ,
         \SB2_1_29/i0[8] , \SB2_1_29/i0[7] , \SB2_1_29/i0[6] ,
         \SB2_1_30/buf_output[5] , \SB2_1_30/buf_output[4] ,
         \SB2_1_30/buf_output[3] , \SB2_1_30/buf_output[2] ,
         \SB2_1_30/buf_output[1] , \SB2_1_30/buf_output[0] , \SB2_1_30/i3[0] ,
         \SB2_1_30/i1_5 , \SB2_1_30/i1_7 , \SB2_1_30/i1[9] , \SB2_1_30/i0_0 ,
         \SB2_1_30/i0_3 , \SB2_1_30/i0_4 , \SB2_1_30/i0[9] , \SB2_1_30/i0[8] ,
         \SB2_1_30/i0[6] , \SB2_1_31/buf_output[5] , \SB2_1_31/buf_output[4] ,
         \SB2_1_31/buf_output[3] , \SB2_1_31/buf_output[2] ,
         \SB2_1_31/buf_output[1] , \SB2_1_31/buf_output[0] , \SB2_1_31/i3[0] ,
         \SB2_1_31/i1_7 , \SB2_1_31/i1[9] , \SB2_1_31/i0_0 , \SB2_1_31/i0_3 ,
         \SB2_1_31/i0_4 , \SB2_1_31/i0[10] , \SB2_1_31/i0[9] ,
         \SB2_1_31/i0[8] , \SB2_1_31/i0[7] , \SB2_1_31/i0[6] ,
         \SB1_2_0/buf_output[5] , \SB1_2_0/buf_output[3] ,
         \SB1_2_0/buf_output[2] , \SB1_2_0/buf_output[1] ,
         \SB1_2_0/buf_output[0] , \SB1_2_0/i3[0] , \SB1_2_0/i1_5 ,
         \SB1_2_0/i1_7 , \SB1_2_0/i1[9] , \SB1_2_0/i0_0 , \SB1_2_0/i0_3 ,
         \SB1_2_0/i0_4 , \SB1_2_0/i0[10] , \SB1_2_0/i0[9] , \SB1_2_0/i0[8] ,
         \SB1_2_0/i0[7] , \SB1_2_0/i0[6] , \SB1_2_1/buf_output[5] ,
         \SB1_2_1/buf_output[4] , \SB1_2_1/buf_output[3] ,
         \SB1_2_1/buf_output[2] , \SB1_2_1/buf_output[1] ,
         \SB1_2_1/buf_output[0] , \SB1_2_1/i3[0] , \SB1_2_1/i1_5 ,
         \SB1_2_1/i1_7 , \SB1_2_1/i1[9] , \SB1_2_1/i0_0 , \SB1_2_1/i0_3 ,
         \SB1_2_1/i0_4 , \SB1_2_1/i0[10] , \SB1_2_1/i0[9] , \SB1_2_1/i0[8] ,
         \SB1_2_1/i0[7] , \SB1_2_1/i0[6] , \SB1_2_2/buf_output[5] ,
         \SB1_2_2/buf_output[3] , \SB1_2_2/buf_output[2] ,
         \SB1_2_2/buf_output[1] , \SB1_2_2/buf_output[0] , \SB1_2_2/i3[0] ,
         \SB1_2_2/i1_5 , \SB1_2_2/i1_7 , \SB1_2_2/i1[9] , \SB1_2_2/i0_0 ,
         \SB1_2_2/i0_3 , \SB1_2_2/i0_4 , \SB1_2_2/i0[10] , \SB1_2_2/i0[9] ,
         \SB1_2_2/i0[8] , \SB1_2_2/i0[7] , \SB1_2_2/i0[6] ,
         \SB1_2_3/buf_output[5] , \SB1_2_3/buf_output[4] ,
         \SB1_2_3/buf_output[3] , \SB1_2_3/buf_output[2] ,
         \SB1_2_3/buf_output[1] , \SB1_2_3/buf_output[0] , \SB1_2_3/i3[0] ,
         \SB1_2_3/i1_5 , \SB1_2_3/i1_7 , \SB1_2_3/i1[9] , \SB1_2_3/i0_0 ,
         \SB1_2_3/i0_3 , \SB1_2_3/i0_4 , \SB1_2_3/i0[10] , \SB1_2_3/i0[9] ,
         \SB1_2_3/i0[8] , \SB1_2_3/i0[7] , \SB1_2_3/i0[6] ,
         \SB1_2_4/buf_output[5] , \SB1_2_4/buf_output[4] ,
         \SB1_2_4/buf_output[3] , \SB1_2_4/buf_output[2] ,
         \SB1_2_4/buf_output[1] , \SB1_2_4/buf_output[0] , \SB1_2_4/i3[0] ,
         \SB1_2_4/i1_5 , \SB1_2_4/i1_7 , \SB1_2_4/i1[9] , \SB1_2_4/i0_0 ,
         \SB1_2_4/i0_3 , \SB1_2_4/i0_4 , \SB1_2_4/i0[10] , \SB1_2_4/i0[9] ,
         \SB1_2_4/i0[8] , \SB1_2_4/i0[7] , \SB1_2_4/i0[6] ,
         \SB1_2_5/buf_output[5] , \SB1_2_5/buf_output[3] ,
         \SB1_2_5/buf_output[2] , \SB1_2_5/buf_output[1] ,
         \SB1_2_5/buf_output[0] , \SB1_2_5/i3[0] , \SB1_2_5/i1_5 ,
         \SB1_2_5/i1_7 , \SB1_2_5/i1[9] , \SB1_2_5/i0_0 , \SB1_2_5/i0_3 ,
         \SB1_2_5/i0_4 , \SB1_2_5/i0[10] , \SB1_2_5/i0[9] , \SB1_2_5/i0[8] ,
         \SB1_2_5/i0[7] , \SB1_2_5/i0[6] , \SB1_2_6/buf_output[5] ,
         \SB1_2_6/buf_output[4] , \SB1_2_6/buf_output[3] ,
         \SB1_2_6/buf_output[2] , \SB1_2_6/buf_output[1] ,
         \SB1_2_6/buf_output[0] , \SB1_2_6/i3[0] , \SB1_2_6/i1_5 ,
         \SB1_2_6/i1_7 , \SB1_2_6/i1[9] , \SB1_2_6/i0_0 , \SB1_2_6/i0_3 ,
         \SB1_2_6/i0_4 , \SB1_2_6/i0[10] , \SB1_2_6/i0[9] , \SB1_2_6/i0[8] ,
         \SB1_2_6/i0[7] , \SB1_2_6/i0[6] , \SB1_2_7/buf_output[5] ,
         \SB1_2_7/buf_output[4] , \SB1_2_7/buf_output[3] ,
         \SB1_2_7/buf_output[2] , \SB1_2_7/buf_output[1] ,
         \SB1_2_7/buf_output[0] , \SB1_2_7/i3[0] , \SB1_2_7/i1_5 ,
         \SB1_2_7/i1_7 , \SB1_2_7/i1[9] , \SB1_2_7/i0_0 , \SB1_2_7/i0_3 ,
         \SB1_2_7/i0_4 , \SB1_2_7/i0[10] , \SB1_2_7/i0[9] , \SB1_2_7/i0[8] ,
         \SB1_2_7/i0[7] , \SB1_2_7/i0[6] , \SB1_2_8/buf_output[5] ,
         \SB1_2_8/buf_output[4] , \SB1_2_8/buf_output[3] ,
         \SB1_2_8/buf_output[2] , \SB1_2_8/buf_output[1] ,
         \SB1_2_8/buf_output[0] , \SB1_2_8/i3[0] , \SB1_2_8/i1_5 ,
         \SB1_2_8/i1_7 , \SB1_2_8/i1[9] , \SB1_2_8/i0_0 , \SB1_2_8/i0_3 ,
         \SB1_2_8/i0_4 , \SB1_2_8/i0[10] , \SB1_2_8/i0[9] , \SB1_2_8/i0[8] ,
         \SB1_2_8/i0[7] , \SB1_2_8/i0[6] , \SB1_2_9/buf_output[5] ,
         \SB1_2_9/buf_output[3] , \SB1_2_9/buf_output[2] ,
         \SB1_2_9/buf_output[1] , \SB1_2_9/buf_output[0] , \SB1_2_9/i3[0] ,
         \SB1_2_9/i1_5 , \SB1_2_9/i1_7 , \SB1_2_9/i1[9] , \SB1_2_9/i0_0 ,
         \SB1_2_9/i0_3 , \SB1_2_9/i0_4 , \SB1_2_9/i0[10] , \SB1_2_9/i0[9] ,
         \SB1_2_9/i0[8] , \SB1_2_9/i0[7] , \SB1_2_9/i0[6] ,
         \SB1_2_10/buf_output[5] , \SB1_2_10/buf_output[3] ,
         \SB1_2_10/buf_output[2] , \SB1_2_10/buf_output[1] ,
         \SB1_2_10/buf_output[0] , \SB1_2_10/i3[0] , \SB1_2_10/i1_5 ,
         \SB1_2_10/i1_7 , \SB1_2_10/i1[9] , \SB1_2_10/i0_0 , \SB1_2_10/i0_3 ,
         \SB1_2_10/i0_4 , \SB1_2_10/i0[10] , \SB1_2_10/i0[9] ,
         \SB1_2_10/i0[8] , \SB1_2_10/i0[7] , \SB1_2_10/i0[6] ,
         \SB1_2_11/buf_output[5] , \SB1_2_11/buf_output[3] ,
         \SB1_2_11/buf_output[2] , \SB1_2_11/buf_output[1] ,
         \SB1_2_11/buf_output[0] , \SB1_2_11/i3[0] , \SB1_2_11/i1_5 ,
         \SB1_2_11/i1_7 , \SB1_2_11/i1[9] , \SB1_2_11/i0_0 , \SB1_2_11/i0_3 ,
         \SB1_2_11/i0_4 , \SB1_2_11/i0[10] , \SB1_2_11/i0[9] ,
         \SB1_2_11/i0[8] , \SB1_2_11/i0[7] , \SB1_2_11/i0[6] ,
         \SB1_2_12/buf_output[5] , \SB1_2_12/buf_output[4] ,
         \SB1_2_12/buf_output[3] , \SB1_2_12/buf_output[2] ,
         \SB1_2_12/buf_output[1] , \SB1_2_12/buf_output[0] , \SB1_2_12/i3[0] ,
         \SB1_2_12/i1_5 , \SB1_2_12/i1_7 , \SB1_2_12/i1[9] , \SB1_2_12/i0_0 ,
         \SB1_2_12/i0_3 , \SB1_2_12/i0_4 , \SB1_2_12/i0[10] , \SB1_2_12/i0[9] ,
         \SB1_2_12/i0[8] , \SB1_2_12/i0[7] , \SB1_2_12/i0[6] ,
         \SB1_2_13/buf_output[5] , \SB1_2_13/buf_output[4] ,
         \SB1_2_13/buf_output[3] , \SB1_2_13/buf_output[2] ,
         \SB1_2_13/buf_output[1] , \SB1_2_13/buf_output[0] , \SB1_2_13/i3[0] ,
         \SB1_2_13/i1_5 , \SB1_2_13/i1_7 , \SB1_2_13/i1[9] , \SB1_2_13/i0_0 ,
         \SB1_2_13/i0_3 , \SB1_2_13/i0_4 , \SB1_2_13/i0[10] , \SB1_2_13/i0[9] ,
         \SB1_2_13/i0[8] , \SB1_2_13/i0[7] , \SB1_2_13/i0[6] ,
         \SB1_2_14/buf_output[5] , \SB1_2_14/buf_output[3] ,
         \SB1_2_14/buf_output[2] , \SB1_2_14/buf_output[1] ,
         \SB1_2_14/buf_output[0] , \SB1_2_14/i3[0] , \SB1_2_14/i1_5 ,
         \SB1_2_14/i1_7 , \SB1_2_14/i1[9] , \SB1_2_14/i0_0 , \SB1_2_14/i0_3 ,
         \SB1_2_14/i0_4 , \SB1_2_14/i0[10] , \SB1_2_14/i0[9] ,
         \SB1_2_14/i0[8] , \SB1_2_14/i0[7] , \SB1_2_14/i0[6] ,
         \SB1_2_15/buf_output[5] , \SB1_2_15/buf_output[3] ,
         \SB1_2_15/buf_output[2] , \SB1_2_15/buf_output[1] ,
         \SB1_2_15/buf_output[0] , \SB1_2_15/i3[0] , \SB1_2_15/i1_5 ,
         \SB1_2_15/i1_7 , \SB1_2_15/i1[9] , \SB1_2_15/i0_0 , \SB1_2_15/i0_3 ,
         \SB1_2_15/i0_4 , \SB1_2_15/i0[10] , \SB1_2_15/i0[9] ,
         \SB1_2_15/i0[8] , \SB1_2_15/i0[7] , \SB1_2_15/i0[6] ,
         \SB1_2_16/buf_output[5] , \SB1_2_16/buf_output[3] ,
         \SB1_2_16/buf_output[2] , \SB1_2_16/buf_output[1] ,
         \SB1_2_16/buf_output[0] , \SB1_2_16/i3[0] , \SB1_2_16/i1_5 ,
         \SB1_2_16/i1_7 , \SB1_2_16/i1[9] , \SB1_2_16/i0_0 , \SB1_2_16/i0_4 ,
         \SB1_2_16/i0[10] , \SB1_2_16/i0[9] , \SB1_2_16/i0[8] ,
         \SB1_2_16/i0[7] , \SB1_2_16/i0[6] , \SB1_2_17/buf_output[5] ,
         \SB1_2_17/buf_output[4] , \SB1_2_17/buf_output[3] ,
         \SB1_2_17/buf_output[2] , \SB1_2_17/buf_output[1] ,
         \SB1_2_17/buf_output[0] , \SB1_2_17/i3[0] , \SB1_2_17/i1_5 ,
         \SB1_2_17/i1_7 , \SB1_2_17/i1[9] , \SB1_2_17/i0_0 , \SB1_2_17/i0_3 ,
         \SB1_2_17/i0_4 , \SB1_2_17/i0[10] , \SB1_2_17/i0[9] ,
         \SB1_2_17/i0[8] , \SB1_2_17/i0[7] , \SB1_2_17/i0[6] ,
         \SB1_2_18/buf_output[5] , \SB1_2_18/buf_output[4] ,
         \SB1_2_18/buf_output[3] , \SB1_2_18/buf_output[2] ,
         \SB1_2_18/buf_output[1] , \SB1_2_18/buf_output[0] , \SB1_2_18/i3[0] ,
         \SB1_2_18/i1_5 , \SB1_2_18/i1_7 , \SB1_2_18/i1[9] , \SB1_2_18/i0_0 ,
         \SB1_2_18/i0_3 , \SB1_2_18/i0_4 , \SB1_2_18/i0[10] , \SB1_2_18/i0[9] ,
         \SB1_2_18/i0[7] , \SB1_2_18/i0[6] , \SB1_2_19/buf_output[5] ,
         \SB1_2_19/buf_output[4] , \SB1_2_19/buf_output[3] ,
         \SB1_2_19/buf_output[2] , \SB1_2_19/buf_output[1] ,
         \SB1_2_19/buf_output[0] , \SB1_2_19/i3[0] , \SB1_2_19/i1_5 ,
         \SB1_2_19/i1_7 , \SB1_2_19/i1[9] , \SB1_2_19/i0_0 , \SB1_2_19/i0_3 ,
         \SB1_2_19/i0_4 , \SB1_2_19/i0[10] , \SB1_2_19/i0[9] ,
         \SB1_2_19/i0[8] , \SB1_2_19/i0[7] , \SB1_2_19/i0[6] ,
         \SB1_2_20/buf_output[5] , \SB1_2_20/buf_output[4] ,
         \SB1_2_20/buf_output[3] , \SB1_2_20/buf_output[2] ,
         \SB1_2_20/buf_output[1] , \SB1_2_20/buf_output[0] , \SB1_2_20/i3[0] ,
         \SB1_2_20/i1_7 , \SB1_2_20/i1[9] , \SB1_2_20/i0_0 , \SB1_2_20/i0_3 ,
         \SB1_2_20/i0_4 , \SB1_2_20/i0[10] , \SB1_2_20/i0[9] ,
         \SB1_2_20/i0[7] , \SB1_2_20/i0[6] , \SB1_2_21/buf_output[5] ,
         \SB1_2_21/buf_output[4] , \SB1_2_21/buf_output[3] ,
         \SB1_2_21/buf_output[2] , \SB1_2_21/buf_output[1] ,
         \SB1_2_21/buf_output[0] , \SB1_2_21/i3[0] , \SB1_2_21/i1_5 ,
         \SB1_2_21/i1_7 , \SB1_2_21/i1[9] , \SB1_2_21/i0_0 , \SB1_2_21/i0_3 ,
         \SB1_2_21/i0_4 , \SB1_2_21/i0[10] , \SB1_2_21/i0[9] ,
         \SB1_2_21/i0[8] , \SB1_2_21/i0[7] , \SB1_2_21/i0[6] ,
         \SB1_2_22/buf_output[5] , \SB1_2_22/buf_output[4] ,
         \SB1_2_22/buf_output[3] , \SB1_2_22/buf_output[2] ,
         \SB1_2_22/buf_output[1] , \SB1_2_22/buf_output[0] , \SB1_2_22/i3[0] ,
         \SB1_2_22/i1_5 , \SB1_2_22/i1_7 , \SB1_2_22/i1[9] , \SB1_2_22/i0_0 ,
         \SB1_2_22/i0_3 , \SB1_2_22/i0_4 , \SB1_2_22/i0[10] , \SB1_2_22/i0[9] ,
         \SB1_2_22/i0[8] , \SB1_2_22/i0[7] , \SB1_2_22/i0[6] ,
         \SB1_2_23/buf_output[5] , \SB1_2_23/buf_output[4] ,
         \SB1_2_23/buf_output[3] , \SB1_2_23/buf_output[2] ,
         \SB1_2_23/buf_output[1] , \SB1_2_23/buf_output[0] , \SB1_2_23/i3[0] ,
         \SB1_2_23/i1_5 , \SB1_2_23/i1_7 , \SB1_2_23/i1[9] , \SB1_2_23/i0_0 ,
         \SB1_2_23/i0_3 , \SB1_2_23/i0_4 , \SB1_2_23/i0[10] , \SB1_2_23/i0[9] ,
         \SB1_2_23/i0[8] , \SB1_2_23/i0[7] , \SB1_2_23/i0[6] ,
         \SB1_2_24/buf_output[5] , \SB1_2_24/buf_output[4] ,
         \SB1_2_24/buf_output[3] , \SB1_2_24/buf_output[2] ,
         \SB1_2_24/buf_output[1] , \SB1_2_24/buf_output[0] , \SB1_2_24/i3[0] ,
         \SB1_2_24/i1_5 , \SB1_2_24/i1_7 , \SB1_2_24/i1[9] , \SB1_2_24/i0_0 ,
         \SB1_2_24/i0_4 , \SB1_2_24/i0[10] , \SB1_2_24/i0[9] ,
         \SB1_2_24/i0[8] , \SB1_2_24/i0[7] , \SB1_2_24/i0[6] ,
         \SB1_2_25/buf_output[5] , \SB1_2_25/buf_output[4] ,
         \SB1_2_25/buf_output[3] , \SB1_2_25/buf_output[2] ,
         \SB1_2_25/buf_output[1] , \SB1_2_25/buf_output[0] , \SB1_2_25/i3[0] ,
         \SB1_2_25/i1_5 , \SB1_2_25/i1_7 , \SB1_2_25/i1[9] , \SB1_2_25/i0_0 ,
         \SB1_2_25/i0_3 , \SB1_2_25/i0_4 , \SB1_2_25/i0[10] , \SB1_2_25/i0[9] ,
         \SB1_2_25/i0[8] , \SB1_2_25/i0[7] , \SB1_2_25/i0[6] ,
         \SB1_2_26/buf_output[5] , \SB1_2_26/buf_output[4] ,
         \SB1_2_26/buf_output[3] , \SB1_2_26/buf_output[2] ,
         \SB1_2_26/buf_output[1] , \SB1_2_26/buf_output[0] , \SB1_2_26/i3[0] ,
         \SB1_2_26/i1_5 , \SB1_2_26/i1_7 , \SB1_2_26/i1[9] , \SB1_2_26/i0_0 ,
         \SB1_2_26/i0_4 , \SB1_2_26/i0[10] , \SB1_2_26/i0[9] ,
         \SB1_2_26/i0[8] , \SB1_2_26/i0[7] , \SB1_2_26/i0[6] ,
         \SB1_2_27/buf_output[5] , \SB1_2_27/buf_output[4] ,
         \SB1_2_27/buf_output[3] , \SB1_2_27/buf_output[2] ,
         \SB1_2_27/buf_output[1] , \SB1_2_27/buf_output[0] , \SB1_2_27/i3[0] ,
         \SB1_2_27/i1_5 , \SB1_2_27/i1_7 , \SB1_2_27/i1[9] , \SB1_2_27/i0_0 ,
         \SB1_2_27/i0_3 , \SB1_2_27/i0_4 , \SB1_2_27/i0[10] , \SB1_2_27/i0[9] ,
         \SB1_2_27/i0[8] , \SB1_2_27/i0[7] , \SB1_2_27/i0[6] ,
         \SB1_2_28/buf_output[5] , \SB1_2_28/buf_output[4] ,
         \SB1_2_28/buf_output[3] , \SB1_2_28/buf_output[2] ,
         \SB1_2_28/buf_output[1] , \SB1_2_28/buf_output[0] , \SB1_2_28/i3[0] ,
         \SB1_2_28/i1_5 , \SB1_2_28/i1_7 , \SB1_2_28/i1[9] , \SB1_2_28/i0_0 ,
         \SB1_2_28/i0_3 , \SB1_2_28/i0_4 , \SB1_2_28/i0[10] , \SB1_2_28/i0[9] ,
         \SB1_2_28/i0[8] , \SB1_2_28/i0[7] , \SB1_2_28/i0[6] ,
         \SB1_2_29/buf_output[5] , \SB1_2_29/buf_output[3] ,
         \SB1_2_29/buf_output[2] , \SB1_2_29/buf_output[1] ,
         \SB1_2_29/buf_output[0] , \SB1_2_29/i3[0] , \SB1_2_29/i1_5 ,
         \SB1_2_29/i1_7 , \SB1_2_29/i1[9] , \SB1_2_29/i0_0 , \SB1_2_29/i0_4 ,
         \SB1_2_29/i0[10] , \SB1_2_29/i0[9] , \SB1_2_29/i0[8] ,
         \SB1_2_29/i0[7] , \SB1_2_29/i0[6] , \SB1_2_30/buf_output[5] ,
         \SB1_2_30/buf_output[3] , \SB1_2_30/buf_output[2] ,
         \SB1_2_30/buf_output[1] , \SB1_2_30/buf_output[0] , \SB1_2_30/i3[0] ,
         \SB1_2_30/i1_5 , \SB1_2_30/i1_7 , \SB1_2_30/i1[9] , \SB1_2_30/i0_0 ,
         \SB1_2_30/i0_3 , \SB1_2_30/i0_4 , \SB1_2_30/i0[10] , \SB1_2_30/i0[9] ,
         \SB1_2_30/i0[8] , \SB1_2_30/i0[7] , \SB1_2_30/i0[6] ,
         \SB1_2_31/buf_output[5] , \SB1_2_31/buf_output[3] ,
         \SB1_2_31/buf_output[2] , \SB1_2_31/buf_output[1] ,
         \SB1_2_31/buf_output[0] , \SB1_2_31/i3[0] , \SB1_2_31/i1_5 ,
         \SB1_2_31/i1_7 , \SB1_2_31/i1[9] , \SB1_2_31/i0_0 , \SB1_2_31/i0_3 ,
         \SB1_2_31/i0_4 , \SB1_2_31/i0[10] , \SB1_2_31/i0[9] ,
         \SB1_2_31/i0[8] , \SB1_2_31/i0[7] , \SB1_2_31/i0[6] ,
         \SB2_2_0/buf_output[5] , \SB2_2_0/buf_output[4] ,
         \SB2_2_0/buf_output[3] , \SB2_2_0/buf_output[2] ,
         \SB2_2_0/buf_output[1] , \SB2_2_0/buf_output[0] , \SB2_2_0/i3[0] ,
         \SB2_2_0/i1_5 , \SB2_2_0/i1_7 , \SB2_2_0/i1[9] , \SB2_2_0/i0_0 ,
         \SB2_2_0/i0_3 , \SB2_2_0/i0_4 , \SB2_2_0/i0[10] , \SB2_2_0/i0[9] ,
         \SB2_2_0/i0[8] , \SB2_2_0/i0[7] , \SB2_2_0/i0[6] ,
         \SB2_2_1/buf_output[5] , \SB2_2_1/buf_output[4] ,
         \SB2_2_1/buf_output[3] , \SB2_2_1/buf_output[2] ,
         \SB2_2_1/buf_output[1] , \SB2_2_1/buf_output[0] , \SB2_2_1/i3[0] ,
         \SB2_2_1/i1_5 , \SB2_2_1/i1_7 , \SB2_2_1/i1[9] , \SB2_2_1/i0_0 ,
         \SB2_2_1/i0_3 , \SB2_2_1/i0_4 , \SB2_2_1/i0[10] , \SB2_2_1/i0[9] ,
         \SB2_2_1/i0[8] , \SB2_2_1/i0[7] , \SB2_2_1/i0[6] ,
         \SB2_2_2/buf_output[5] , \SB2_2_2/buf_output[4] ,
         \SB2_2_2/buf_output[3] , \SB2_2_2/buf_output[2] ,
         \SB2_2_2/buf_output[1] , \SB2_2_2/buf_output[0] , \SB2_2_2/i3[0] ,
         \SB2_2_2/i1_5 , \SB2_2_2/i1_7 , \SB2_2_2/i1[9] , \SB2_2_2/i0_0 ,
         \SB2_2_2/i0_3 , \SB2_2_2/i0_4 , \SB2_2_2/i0[10] , \SB2_2_2/i0[9] ,
         \SB2_2_2/i0[8] , \SB2_2_2/i0[7] , \SB2_2_2/i0[6] ,
         \SB2_2_3/buf_output[5] , \SB2_2_3/buf_output[4] ,
         \SB2_2_3/buf_output[3] , \SB2_2_3/buf_output[2] ,
         \SB2_2_3/buf_output[1] , \SB2_2_3/buf_output[0] , \SB2_2_3/i3[0] ,
         \SB2_2_3/i1_5 , \SB2_2_3/i1_7 , \SB2_2_3/i1[9] , \SB2_2_3/i0_0 ,
         \SB2_2_3/i0_3 , \SB2_2_3/i0[10] , \SB2_2_3/i0[9] , \SB2_2_3/i0[8] ,
         \SB2_2_3/i0[6] , \SB2_2_4/buf_output[5] , \SB2_2_4/buf_output[4] ,
         \SB2_2_4/buf_output[3] , \SB2_2_4/buf_output[2] ,
         \SB2_2_4/buf_output[1] , \SB2_2_4/buf_output[0] , \SB2_2_4/i3[0] ,
         \SB2_2_4/i1_5 , \SB2_2_4/i1_7 , \SB2_2_4/i1[9] , \SB2_2_4/i0_0 ,
         \SB2_2_4/i0_3 , \SB2_2_4/i0_4 , \SB2_2_4/i0[10] , \SB2_2_4/i0[9] ,
         \SB2_2_4/i0[8] , \SB2_2_4/i0[7] , \SB2_2_4/i0[6] ,
         \SB2_2_5/buf_output[5] , \SB2_2_5/buf_output[4] ,
         \SB2_2_5/buf_output[3] , \SB2_2_5/buf_output[2] ,
         \SB2_2_5/buf_output[1] , \SB2_2_5/buf_output[0] , \SB2_2_5/i3[0] ,
         \SB2_2_5/i1_5 , \SB2_2_5/i1_7 , \SB2_2_5/i1[9] , \SB2_2_5/i0_0 ,
         \SB2_2_5/i0_3 , \SB2_2_5/i0_4 , \SB2_2_5/i0[10] , \SB2_2_5/i0[9] ,
         \SB2_2_5/i0[8] , \SB2_2_5/i0[7] , \SB2_2_5/i0[6] ,
         \SB2_2_6/buf_output[5] , \SB2_2_6/buf_output[4] ,
         \SB2_2_6/buf_output[3] , \SB2_2_6/buf_output[2] ,
         \SB2_2_6/buf_output[1] , \SB2_2_6/buf_output[0] , \SB2_2_6/i3[0] ,
         \SB2_2_6/i1_5 , \SB2_2_6/i1_7 , \SB2_2_6/i1[9] , \SB2_2_6/i0_0 ,
         \SB2_2_6/i0_3 , \SB2_2_6/i0[10] , \SB2_2_6/i0[9] , \SB2_2_6/i0[8] ,
         \SB2_2_6/i0[7] , \SB2_2_6/i0[6] , \SB2_2_7/buf_output[5] ,
         \SB2_2_7/buf_output[4] , \SB2_2_7/buf_output[3] ,
         \SB2_2_7/buf_output[2] , \SB2_2_7/buf_output[1] ,
         \SB2_2_7/buf_output[0] , \SB2_2_7/i3[0] , \SB2_2_7/i1_5 ,
         \SB2_2_7/i1_7 , \SB2_2_7/i1[9] , \SB2_2_7/i0_0 , \SB2_2_7/i0_3 ,
         \SB2_2_7/i0[10] , \SB2_2_7/i0[9] , \SB2_2_7/i0[8] , \SB2_2_7/i0[7] ,
         \SB2_2_7/i0[6] , \SB2_2_8/buf_output[5] , \SB2_2_8/buf_output[4] ,
         \SB2_2_8/buf_output[3] , \SB2_2_8/buf_output[2] ,
         \SB2_2_8/buf_output[1] , \SB2_2_8/buf_output[0] , \SB2_2_8/i3[0] ,
         \SB2_2_8/i1_5 , \SB2_2_8/i1_7 , \SB2_2_8/i1[9] , \SB2_2_8/i0_0 ,
         \SB2_2_8/i0_3 , \SB2_2_8/i0_4 , \SB2_2_8/i0[10] , \SB2_2_8/i0[9] ,
         \SB2_2_8/i0[8] , \SB2_2_8/i0[7] , \SB2_2_8/i0[6] ,
         \SB2_2_9/buf_output[5] , \SB2_2_9/buf_output[4] ,
         \SB2_2_9/buf_output[3] , \SB2_2_9/buf_output[2] ,
         \SB2_2_9/buf_output[0] , \SB2_2_9/i3[0] , \SB2_2_9/i1_7 ,
         \SB2_2_9/i1[9] , \SB2_2_9/i0_0 , \SB2_2_9/i0_3 , \SB2_2_9/i0_4 ,
         \SB2_2_9/i0[10] , \SB2_2_9/i0[9] , \SB2_2_9/i0[8] , \SB2_2_9/i0[6] ,
         \SB2_2_10/buf_output[5] , \SB2_2_10/buf_output[4] ,
         \SB2_2_10/buf_output[3] , \SB2_2_10/buf_output[2] ,
         \SB2_2_10/buf_output[1] , \SB2_2_10/buf_output[0] , \SB2_2_10/i3[0] ,
         \SB2_2_10/i1_5 , \SB2_2_10/i1_7 , \SB2_2_10/i1[9] , \SB2_2_10/i0_0 ,
         \SB2_2_10/i0_3 , \SB2_2_10/i0[10] , \SB2_2_10/i0[9] ,
         \SB2_2_10/i0[8] , \SB2_2_10/i0[7] , \SB2_2_10/i0[6] ,
         \SB2_2_11/buf_output[5] , \SB2_2_11/buf_output[4] ,
         \SB2_2_11/buf_output[3] , \SB2_2_11/buf_output[2] ,
         \SB2_2_11/buf_output[1] , \SB2_2_11/buf_output[0] , \SB2_2_11/i3[0] ,
         \SB2_2_11/i1_5 , \SB2_2_11/i1_7 , \SB2_2_11/i0_0 , \SB2_2_11/i0_3 ,
         \SB2_2_11/i0_4 , \SB2_2_11/i0[9] , \SB2_2_11/i0[8] , \SB2_2_11/i0[7] ,
         \SB2_2_11/i0[6] , \SB2_2_12/buf_output[5] , \SB2_2_12/buf_output[4] ,
         \SB2_2_12/buf_output[3] , \SB2_2_12/buf_output[2] ,
         \SB2_2_12/buf_output[0] , \SB2_2_12/i3[0] , \SB2_2_12/i1_5 ,
         \SB2_2_12/i1_7 , \SB2_2_12/i1[9] , \SB2_2_12/i0_0 , \SB2_2_12/i0_3 ,
         \SB2_2_12/i0_4 , \SB2_2_12/i0[10] , \SB2_2_12/i0[9] ,
         \SB2_2_12/i0[8] , \SB2_2_12/i0[7] , \SB2_2_12/i0[6] ,
         \SB2_2_13/buf_output[5] , \SB2_2_13/buf_output[4] ,
         \SB2_2_13/buf_output[3] , \SB2_2_13/buf_output[2] ,
         \SB2_2_13/buf_output[1] , \SB2_2_13/buf_output[0] , \SB2_2_13/i3[0] ,
         \SB2_2_13/i1_7 , \SB2_2_13/i1[9] , \SB2_2_13/i0_0 , \SB2_2_13/i0_3 ,
         \SB2_2_13/i0[10] , \SB2_2_13/i0[9] , \SB2_2_13/i0[8] ,
         \SB2_2_13/i0[7] , \SB2_2_13/i0[6] , \SB2_2_14/buf_output[5] ,
         \SB2_2_14/buf_output[4] , \SB2_2_14/buf_output[3] ,
         \SB2_2_14/buf_output[2] , \SB2_2_14/buf_output[1] ,
         \SB2_2_14/buf_output[0] , \SB2_2_14/i3[0] , \SB2_2_14/i1_5 ,
         \SB2_2_14/i1_7 , \SB2_2_14/i1[9] , \SB2_2_14/i0_0 , \SB2_2_14/i0_3 ,
         \SB2_2_14/i0_4 , \SB2_2_14/i0[10] , \SB2_2_14/i0[9] ,
         \SB2_2_14/i0[8] , \SB2_2_14/i0[7] , \SB2_2_14/i0[6] ,
         \SB2_2_15/buf_output[5] , \SB2_2_15/buf_output[4] ,
         \SB2_2_15/buf_output[3] , \SB2_2_15/buf_output[2] ,
         \SB2_2_15/buf_output[1] , \SB2_2_15/buf_output[0] , \SB2_2_15/i3[0] ,
         \SB2_2_15/i1_5 , \SB2_2_15/i1_7 , \SB2_2_15/i1[9] , \SB2_2_15/i0_0 ,
         \SB2_2_15/i0_3 , \SB2_2_15/i0_4 , \SB2_2_15/i0[10] , \SB2_2_15/i0[9] ,
         \SB2_2_15/i0[8] , \SB2_2_15/i0[6] , \SB2_2_16/buf_output[5] ,
         \SB2_2_16/buf_output[4] , \SB2_2_16/buf_output[3] ,
         \SB2_2_16/buf_output[2] , \SB2_2_16/buf_output[1] ,
         \SB2_2_16/buf_output[0] , \SB2_2_16/i3[0] , \SB2_2_16/i1_5 ,
         \SB2_2_16/i1_7 , \SB2_2_16/i1[9] , \SB2_2_16/i0_0 , \SB2_2_16/i0_3 ,
         \SB2_2_16/i0_4 , \SB2_2_16/i0[10] , \SB2_2_16/i0[9] ,
         \SB2_2_16/i0[8] , \SB2_2_16/i0[7] , \SB2_2_16/i0[6] ,
         \SB2_2_17/buf_output[5] , \SB2_2_17/buf_output[4] ,
         \SB2_2_17/buf_output[3] , \SB2_2_17/buf_output[2] ,
         \SB2_2_17/buf_output[1] , \SB2_2_17/buf_output[0] , \SB2_2_17/i3[0] ,
         \SB2_2_17/i1_5 , \SB2_2_17/i1_7 , \SB2_2_17/i1[9] , \SB2_2_17/i0_0 ,
         \SB2_2_17/i0_3 , \SB2_2_17/i0_4 , \SB2_2_17/i0[10] , \SB2_2_17/i0[9] ,
         \SB2_2_17/i0[8] , \SB2_2_17/i0[7] , \SB2_2_17/i0[6] ,
         \SB2_2_18/buf_output[5] , \SB2_2_18/buf_output[4] ,
         \SB2_2_18/buf_output[3] , \SB2_2_18/buf_output[2] ,
         \SB2_2_18/buf_output[1] , \SB2_2_18/buf_output[0] , \SB2_2_18/i3[0] ,
         \SB2_2_18/i1_7 , \SB2_2_18/i1[9] , \SB2_2_18/i0_0 , \SB2_2_18/i0_3 ,
         \SB2_2_18/i0_4 , \SB2_2_18/i0[10] , \SB2_2_18/i0[9] ,
         \SB2_2_18/i0[8] , \SB2_2_18/i0[7] , \SB2_2_18/i0[6] ,
         \SB2_2_19/buf_output[5] , \SB2_2_19/buf_output[4] ,
         \SB2_2_19/buf_output[3] , \SB2_2_19/buf_output[2] ,
         \SB2_2_19/buf_output[1] , \SB2_2_19/buf_output[0] , \SB2_2_19/i3[0] ,
         \SB2_2_19/i1_5 , \SB2_2_19/i1_7 , \SB2_2_19/i1[9] , \SB2_2_19/i0_0 ,
         \SB2_2_19/i0_3 , \SB2_2_19/i0_4 , \SB2_2_19/i0[10] , \SB2_2_19/i0[9] ,
         \SB2_2_19/i0[8] , \SB2_2_19/i0[7] , \SB2_2_19/i0[6] ,
         \SB2_2_20/buf_output[5] , \SB2_2_20/buf_output[4] ,
         \SB2_2_20/buf_output[3] , \SB2_2_20/buf_output[2] ,
         \SB2_2_20/buf_output[1] , \SB2_2_20/buf_output[0] , \SB2_2_20/i3[0] ,
         \SB2_2_20/i1_5 , \SB2_2_20/i1_7 , \SB2_2_20/i1[9] , \SB2_2_20/i0_0 ,
         \SB2_2_20/i0_3 , \SB2_2_20/i0_4 , \SB2_2_20/i0[10] , \SB2_2_20/i0[9] ,
         \SB2_2_20/i0[8] , \SB2_2_20/i0[7] , \SB2_2_20/i0[6] ,
         \SB2_2_21/buf_output[5] , \SB2_2_21/buf_output[4] ,
         \SB2_2_21/buf_output[3] , \SB2_2_21/buf_output[2] ,
         \SB2_2_21/buf_output[1] , \SB2_2_21/buf_output[0] , \SB2_2_21/i3[0] ,
         \SB2_2_21/i1_5 , \SB2_2_21/i1_7 , \SB2_2_21/i1[9] , \SB2_2_21/i0_0 ,
         \SB2_2_21/i0_3 , \SB2_2_21/i0_4 , \SB2_2_21/i0[10] , \SB2_2_21/i0[9] ,
         \SB2_2_21/i0[8] , \SB2_2_21/i0[7] , \SB2_2_21/i0[6] ,
         \SB2_2_22/buf_output[5] , \SB2_2_22/buf_output[4] ,
         \SB2_2_22/buf_output[3] , \SB2_2_22/buf_output[2] ,
         \SB2_2_22/buf_output[1] , \SB2_2_22/buf_output[0] , \SB2_2_22/i3[0] ,
         \SB2_2_22/i1_5 , \SB2_2_22/i1_7 , \SB2_2_22/i1[9] , \SB2_2_22/i0_0 ,
         \SB2_2_22/i0_3 , \SB2_2_22/i0_4 , \SB2_2_22/i0[10] , \SB2_2_22/i0[9] ,
         \SB2_2_22/i0[8] , \SB2_2_22/i0[7] , \SB2_2_22/i0[6] ,
         \SB2_2_23/buf_output[5] , \SB2_2_23/buf_output[4] ,
         \SB2_2_23/buf_output[3] , \SB2_2_23/buf_output[2] ,
         \SB2_2_23/buf_output[1] , \SB2_2_23/buf_output[0] , \SB2_2_23/i3[0] ,
         \SB2_2_23/i1_5 , \SB2_2_23/i1_7 , \SB2_2_23/i1[9] , \SB2_2_23/i0_0 ,
         \SB2_2_23/i0_3 , \SB2_2_23/i0_4 , \SB2_2_23/i0[10] , \SB2_2_23/i0[9] ,
         \SB2_2_23/i0[8] , \SB2_2_23/i0[7] , \SB2_2_23/i0[6] ,
         \SB2_2_24/buf_output[5] , \SB2_2_24/buf_output[4] ,
         \SB2_2_24/buf_output[3] , \SB2_2_24/buf_output[2] ,
         \SB2_2_24/buf_output[1] , \SB2_2_24/buf_output[0] , \SB2_2_24/i3[0] ,
         \SB2_2_24/i1_5 , \SB2_2_24/i1_7 , \SB2_2_24/i1[9] , \SB2_2_24/i0_0 ,
         \SB2_2_24/i0_3 , \SB2_2_24/i0_4 , \SB2_2_24/i0[10] , \SB2_2_24/i0[9] ,
         \SB2_2_24/i0[8] , \SB2_2_24/i0[7] , \SB2_2_24/i0[6] ,
         \SB2_2_25/buf_output[5] , \SB2_2_25/buf_output[4] ,
         \SB2_2_25/buf_output[3] , \SB2_2_25/buf_output[2] ,
         \SB2_2_25/buf_output[1] , \SB2_2_25/buf_output[0] , \SB2_2_25/i3[0] ,
         \SB2_2_25/i1_5 , \SB2_2_25/i1_7 , \SB2_2_25/i1[9] , \SB2_2_25/i0_0 ,
         \SB2_2_25/i0_3 , \SB2_2_25/i0_4 , \SB2_2_25/i0[10] , \SB2_2_25/i0[9] ,
         \SB2_2_25/i0[8] , \SB2_2_25/i0[7] , \SB2_2_25/i0[6] ,
         \SB2_2_26/buf_output[5] , \SB2_2_26/buf_output[4] ,
         \SB2_2_26/buf_output[3] , \SB2_2_26/buf_output[2] ,
         \SB2_2_26/buf_output[1] , \SB2_2_26/buf_output[0] , \SB2_2_26/i3[0] ,
         \SB2_2_26/i1_5 , \SB2_2_26/i1_7 , \SB2_2_26/i1[9] , \SB2_2_26/i0_0 ,
         \SB2_2_26/i0_3 , \SB2_2_26/i0_4 , \SB2_2_26/i0[10] , \SB2_2_26/i0[9] ,
         \SB2_2_26/i0[8] , \SB2_2_26/i0[7] , \SB2_2_26/i0[6] ,
         \SB2_2_27/buf_output[5] , \SB2_2_27/buf_output[4] ,
         \SB2_2_27/buf_output[3] , \SB2_2_27/buf_output[2] ,
         \SB2_2_27/buf_output[1] , \SB2_2_27/buf_output[0] , \SB2_2_27/i3[0] ,
         \SB2_2_27/i1_5 , \SB2_2_27/i1_7 , \SB2_2_27/i1[9] , \SB2_2_27/i0_0 ,
         \SB2_2_27/i0_3 , \SB2_2_27/i0[10] , \SB2_2_27/i0[9] ,
         \SB2_2_27/i0[8] , \SB2_2_27/i0[6] , \SB2_2_28/buf_output[5] ,
         \SB2_2_28/buf_output[4] , \SB2_2_28/buf_output[3] ,
         \SB2_2_28/buf_output[2] , \SB2_2_28/buf_output[1] ,
         \SB2_2_28/buf_output[0] , \SB2_2_28/i3[0] , \SB2_2_28/i1_5 ,
         \SB2_2_28/i1_7 , \SB2_2_28/i1[9] , \SB2_2_28/i0_0 , \SB2_2_28/i0_3 ,
         \SB2_2_28/i0_4 , \SB2_2_28/i0[10] , \SB2_2_28/i0[9] ,
         \SB2_2_28/i0[8] , \SB2_2_28/i0[7] , \SB2_2_28/i0[6] ,
         \SB2_2_29/buf_output[5] , \SB2_2_29/buf_output[4] ,
         \SB2_2_29/buf_output[3] , \SB2_2_29/buf_output[2] ,
         \SB2_2_29/buf_output[1] , \SB2_2_29/buf_output[0] , \SB2_2_29/i3[0] ,
         \SB2_2_29/i1_5 , \SB2_2_29/i1_7 , \SB2_2_29/i1[9] , \SB2_2_29/i0_0 ,
         \SB2_2_29/i0_3 , \SB2_2_29/i0_4 , \SB2_2_29/i0[10] , \SB2_2_29/i0[9] ,
         \SB2_2_29/i0[8] , \SB2_2_29/i0[7] , \SB2_2_29/i0[6] ,
         \SB2_2_30/buf_output[5] , \SB2_2_30/buf_output[4] ,
         \SB2_2_30/buf_output[3] , \SB2_2_30/buf_output[2] ,
         \SB2_2_30/buf_output[1] , \SB2_2_30/buf_output[0] , \SB2_2_30/i3[0] ,
         \SB2_2_30/i1_5 , \SB2_2_30/i1_7 , \SB2_2_30/i1[9] , \SB2_2_30/i0_0 ,
         \SB2_2_30/i0_3 , \SB2_2_30/i0_4 , \SB2_2_30/i0[10] , \SB2_2_30/i0[9] ,
         \SB2_2_30/i0[8] , \SB2_2_30/i0[7] , \SB2_2_30/i0[6] ,
         \SB2_2_31/buf_output[5] , \SB2_2_31/buf_output[4] ,
         \SB2_2_31/buf_output[3] , \SB2_2_31/buf_output[2] ,
         \SB2_2_31/buf_output[1] , \SB2_2_31/buf_output[0] , \SB2_2_31/i3[0] ,
         \SB2_2_31/i1_5 , \SB2_2_31/i1_7 , \SB2_2_31/i1[9] , \SB2_2_31/i0_0 ,
         \SB2_2_31/i0_3 , \SB2_2_31/i0[10] , \SB2_2_31/i0[9] ,
         \SB2_2_31/i0[8] , \SB2_2_31/i0[7] , \SB2_2_31/i0[6] ,
         \SB1_3_0/buf_output[5] , \SB1_3_0/buf_output[4] ,
         \SB1_3_0/buf_output[3] , \SB1_3_0/buf_output[2] ,
         \SB1_3_0/buf_output[1] , \SB1_3_0/buf_output[0] , \SB1_3_0/i3[0] ,
         \SB1_3_0/i1_5 , \SB1_3_0/i1_7 , \SB1_3_0/i1[9] , \SB1_3_0/i0_0 ,
         \SB1_3_0/i0_3 , \SB1_3_0/i0_4 , \SB1_3_0/i0[10] , \SB1_3_0/i0[9] ,
         \SB1_3_0/i0[8] , \SB1_3_0/i0[7] , \SB1_3_0/i0[6] ,
         \SB1_3_1/buf_output[5] , \SB1_3_1/buf_output[4] ,
         \SB1_3_1/buf_output[3] , \SB1_3_1/buf_output[2] ,
         \SB1_3_1/buf_output[1] , \SB1_3_1/buf_output[0] , \SB1_3_1/i3[0] ,
         \SB1_3_1/i1_5 , \SB1_3_1/i1_7 , \SB1_3_1/i1[9] , \SB1_3_1/i0_0 ,
         \SB1_3_1/i0_3 , \SB1_3_1/i0_4 , \SB1_3_1/i0[10] , \SB1_3_1/i0[9] ,
         \SB1_3_1/i0[8] , \SB1_3_1/i0[7] , \SB1_3_1/i0[6] ,
         \SB1_3_2/buf_output[5] , \SB1_3_2/buf_output[4] ,
         \SB1_3_2/buf_output[3] , \SB1_3_2/buf_output[2] ,
         \SB1_3_2/buf_output[1] , \SB1_3_2/buf_output[0] , \SB1_3_2/i3[0] ,
         \SB1_3_2/i1_5 , \SB1_3_2/i1_7 , \SB1_3_2/i1[9] , \SB1_3_2/i0_0 ,
         \SB1_3_2/i0_3 , \SB1_3_2/i0_4 , \SB1_3_2/i0[10] , \SB1_3_2/i0[9] ,
         \SB1_3_2/i0[8] , \SB1_3_2/i0[7] , \SB1_3_2/i0[6] ,
         \SB1_3_3/buf_output[5] , \SB1_3_3/buf_output[4] ,
         \SB1_3_3/buf_output[3] , \SB1_3_3/buf_output[2] ,
         \SB1_3_3/buf_output[1] , \SB1_3_3/buf_output[0] , \SB1_3_3/i3[0] ,
         \SB1_3_3/i1_5 , \SB1_3_3/i1_7 , \SB1_3_3/i1[9] , \SB1_3_3/i0_0 ,
         \SB1_3_3/i0_3 , \SB1_3_3/i0_4 , \SB1_3_3/i0[10] , \SB1_3_3/i0[9] ,
         \SB1_3_3/i0[8] , \SB1_3_3/i0[7] , \SB1_3_3/i0[6] ,
         \SB1_3_4/buf_output[5] , \SB1_3_4/buf_output[4] ,
         \SB1_3_4/buf_output[3] , \SB1_3_4/buf_output[2] ,
         \SB1_3_4/buf_output[1] , \SB1_3_4/buf_output[0] , \SB1_3_4/i3[0] ,
         \SB1_3_4/i1_5 , \SB1_3_4/i1_7 , \SB1_3_4/i1[9] , \SB1_3_4/i0_0 ,
         \SB1_3_4/i0_3 , \SB1_3_4/i0_4 , \SB1_3_4/i0[10] , \SB1_3_4/i0[9] ,
         \SB1_3_4/i0[8] , \SB1_3_4/i0[7] , \SB1_3_4/i0[6] ,
         \SB1_3_5/buf_output[5] , \SB1_3_5/buf_output[4] ,
         \SB1_3_5/buf_output[3] , \SB1_3_5/buf_output[2] ,
         \SB1_3_5/buf_output[1] , \SB1_3_5/buf_output[0] , \SB1_3_5/i3[0] ,
         \SB1_3_5/i1_5 , \SB1_3_5/i1_7 , \SB1_3_5/i1[9] , \SB1_3_5/i0_0 ,
         \SB1_3_5/i0_3 , \SB1_3_5/i0_4 , \SB1_3_5/i0[10] , \SB1_3_5/i0[9] ,
         \SB1_3_5/i0[8] , \SB1_3_5/i0[7] , \SB1_3_5/i0[6] ,
         \SB1_3_6/buf_output[5] , \SB1_3_6/buf_output[4] ,
         \SB1_3_6/buf_output[3] , \SB1_3_6/buf_output[2] ,
         \SB1_3_6/buf_output[1] , \SB1_3_6/buf_output[0] , \SB1_3_6/i3[0] ,
         \SB1_3_6/i1_5 , \SB1_3_6/i1_7 , \SB1_3_6/i1[9] , \SB1_3_6/i0_0 ,
         \SB1_3_6/i0_3 , \SB1_3_6/i0_4 , \SB1_3_6/i0[10] , \SB1_3_6/i0[9] ,
         \SB1_3_6/i0[8] , \SB1_3_6/i0[7] , \SB1_3_6/i0[6] ,
         \SB1_3_7/buf_output[5] , \SB1_3_7/buf_output[4] ,
         \SB1_3_7/buf_output[3] , \SB1_3_7/buf_output[2] ,
         \SB1_3_7/buf_output[1] , \SB1_3_7/buf_output[0] , \SB1_3_7/i3[0] ,
         \SB1_3_7/i1_5 , \SB1_3_7/i1_7 , \SB1_3_7/i1[9] , \SB1_3_7/i0_0 ,
         \SB1_3_7/i0_3 , \SB1_3_7/i0_4 , \SB1_3_7/i0[10] , \SB1_3_7/i0[9] ,
         \SB1_3_7/i0[8] , \SB1_3_7/i0[7] , \SB1_3_7/i0[6] ,
         \SB1_3_8/buf_output[5] , \SB1_3_8/buf_output[4] ,
         \SB1_3_8/buf_output[3] , \SB1_3_8/buf_output[2] ,
         \SB1_3_8/buf_output[1] , \SB1_3_8/buf_output[0] , \SB1_3_8/i3[0] ,
         \SB1_3_8/i1_5 , \SB1_3_8/i1_7 , \SB1_3_8/i1[9] , \SB1_3_8/i0_0 ,
         \SB1_3_8/i0_3 , \SB1_3_8/i0_4 , \SB1_3_8/i0[10] , \SB1_3_8/i0[9] ,
         \SB1_3_8/i0[8] , \SB1_3_8/i0[7] , \SB1_3_8/i0[6] ,
         \SB1_3_9/buf_output[5] , \SB1_3_9/buf_output[4] ,
         \SB1_3_9/buf_output[3] , \SB1_3_9/buf_output[2] ,
         \SB1_3_9/buf_output[1] , \SB1_3_9/buf_output[0] , \SB1_3_9/i3[0] ,
         \SB1_3_9/i1_5 , \SB1_3_9/i1_7 , \SB1_3_9/i1[9] , \SB1_3_9/i0_0 ,
         \SB1_3_9/i0_3 , \SB1_3_9/i0_4 , \SB1_3_9/i0[10] , \SB1_3_9/i0[9] ,
         \SB1_3_9/i0[8] , \SB1_3_9/i0[7] , \SB1_3_9/i0[6] ,
         \SB1_3_10/buf_output[5] , \SB1_3_10/buf_output[4] ,
         \SB1_3_10/buf_output[3] , \SB1_3_10/buf_output[2] ,
         \SB1_3_10/buf_output[1] , \SB1_3_10/buf_output[0] , \SB1_3_10/i3[0] ,
         \SB1_3_10/i1_5 , \SB1_3_10/i1_7 , \SB1_3_10/i1[9] , \SB1_3_10/i0_0 ,
         \SB1_3_10/i0_3 , \SB1_3_10/i0_4 , \SB1_3_10/i0[10] , \SB1_3_10/i0[9] ,
         \SB1_3_10/i0[8] , \SB1_3_10/i0[7] , \SB1_3_10/i0[6] ,
         \SB1_3_11/buf_output[5] , \SB1_3_11/buf_output[4] ,
         \SB1_3_11/buf_output[3] , \SB1_3_11/buf_output[2] ,
         \SB1_3_11/buf_output[1] , \SB1_3_11/buf_output[0] , \SB1_3_11/i3[0] ,
         \SB1_3_11/i1_7 , \SB1_3_11/i1[9] , \SB1_3_11/i0_0 , \SB1_3_11/i0_3 ,
         \SB1_3_11/i0_4 , \SB1_3_11/i0[10] , \SB1_3_11/i0[9] ,
         \SB1_3_11/i0[8] , \SB1_3_11/i0[6] , \SB1_3_12/buf_output[5] ,
         \SB1_3_12/buf_output[3] , \SB1_3_12/buf_output[2] ,
         \SB1_3_12/buf_output[1] , \SB1_3_12/buf_output[0] , \SB1_3_12/i3[0] ,
         \SB1_3_12/i1_5 , \SB1_3_12/i1_7 , \SB1_3_12/i1[9] , \SB1_3_12/i0_0 ,
         \SB1_3_12/i0_3 , \SB1_3_12/i0_4 , \SB1_3_12/i0[10] , \SB1_3_12/i0[9] ,
         \SB1_3_12/i0[8] , \SB1_3_12/i0[7] , \SB1_3_12/i0[6] ,
         \SB1_3_13/buf_output[5] , \SB1_3_13/buf_output[4] ,
         \SB1_3_13/buf_output[3] , \SB1_3_13/buf_output[2] ,
         \SB1_3_13/buf_output[1] , \SB1_3_13/buf_output[0] , \SB1_3_13/i3[0] ,
         \SB1_3_13/i1_5 , \SB1_3_13/i1_7 , \SB1_3_13/i1[9] , \SB1_3_13/i0_0 ,
         \SB1_3_13/i0_3 , \SB1_3_13/i0_4 , \SB1_3_13/i0[10] , \SB1_3_13/i0[9] ,
         \SB1_3_13/i0[8] , \SB1_3_13/i0[7] , \SB1_3_13/i0[6] ,
         \SB1_3_14/buf_output[5] , \SB1_3_14/buf_output[4] ,
         \SB1_3_14/buf_output[3] , \SB1_3_14/buf_output[2] ,
         \SB1_3_14/buf_output[1] , \SB1_3_14/buf_output[0] , \SB1_3_14/i3[0] ,
         \SB1_3_14/i1_5 , \SB1_3_14/i1_7 , \SB1_3_14/i1[9] , \SB1_3_14/i0_0 ,
         \SB1_3_14/i0_3 , \SB1_3_14/i0_4 , \SB1_3_14/i0[10] , \SB1_3_14/i0[9] ,
         \SB1_3_14/i0[8] , \SB1_3_14/i0[7] , \SB1_3_14/i0[6] ,
         \SB1_3_15/buf_output[5] , \SB1_3_15/buf_output[4] ,
         \SB1_3_15/buf_output[3] , \SB1_3_15/buf_output[2] ,
         \SB1_3_15/buf_output[1] , \SB1_3_15/buf_output[0] , \SB1_3_15/i3[0] ,
         \SB1_3_15/i1_5 , \SB1_3_15/i1_7 , \SB1_3_15/i1[9] , \SB1_3_15/i0_0 ,
         \SB1_3_15/i0_3 , \SB1_3_15/i0_4 , \SB1_3_15/i0[10] , \SB1_3_15/i0[9] ,
         \SB1_3_15/i0[8] , \SB1_3_15/i0[7] , \SB1_3_15/i0[6] ,
         \SB1_3_16/buf_output[5] , \SB1_3_16/buf_output[4] ,
         \SB1_3_16/buf_output[3] , \SB1_3_16/buf_output[2] ,
         \SB1_3_16/buf_output[1] , \SB1_3_16/buf_output[0] , \SB1_3_16/i3[0] ,
         \SB1_3_16/i1_5 , \SB1_3_16/i1_7 , \SB1_3_16/i1[9] , \SB1_3_16/i0_0 ,
         \SB1_3_16/i0_3 , \SB1_3_16/i0_4 , \SB1_3_16/i0[10] , \SB1_3_16/i0[9] ,
         \SB1_3_16/i0[8] , \SB1_3_16/i0[7] , \SB1_3_16/i0[6] ,
         \SB1_3_17/buf_output[5] , \SB1_3_17/buf_output[4] ,
         \SB1_3_17/buf_output[3] , \SB1_3_17/buf_output[2] ,
         \SB1_3_17/buf_output[1] , \SB1_3_17/i3[0] , \SB1_3_17/i1_5 ,
         \SB1_3_17/i1_7 , \SB1_3_17/i1[9] , \SB1_3_17/i0_0 , \SB1_3_17/i0_3 ,
         \SB1_3_17/i0_4 , \SB1_3_17/i0[10] , \SB1_3_17/i0[9] ,
         \SB1_3_17/i0[8] , \SB1_3_17/i0[7] , \SB1_3_17/i0[6] ,
         \SB1_3_18/buf_output[5] , \SB1_3_18/buf_output[4] ,
         \SB1_3_18/buf_output[3] , \SB1_3_18/buf_output[2] ,
         \SB1_3_18/buf_output[1] , \SB1_3_18/buf_output[0] , \SB1_3_18/i3[0] ,
         \SB1_3_18/i1_5 , \SB1_3_18/i1_7 , \SB1_3_18/i1[9] , \SB1_3_18/i0_0 ,
         \SB1_3_18/i0_3 , \SB1_3_18/i0_4 , \SB1_3_18/i0[10] , \SB1_3_18/i0[9] ,
         \SB1_3_18/i0[8] , \SB1_3_18/i0[7] , \SB1_3_18/i0[6] ,
         \SB1_3_19/buf_output[5] , \SB1_3_19/buf_output[4] ,
         \SB1_3_19/buf_output[3] , \SB1_3_19/buf_output[2] ,
         \SB1_3_19/buf_output[1] , \SB1_3_19/buf_output[0] , \SB1_3_19/i3[0] ,
         \SB1_3_19/i1_5 , \SB1_3_19/i1_7 , \SB1_3_19/i1[9] , \SB1_3_19/i0_0 ,
         \SB1_3_19/i0_3 , \SB1_3_19/i0_4 , \SB1_3_19/i0[10] , \SB1_3_19/i0[9] ,
         \SB1_3_19/i0[8] , \SB1_3_19/i0[7] , \SB1_3_19/i0[6] ,
         \SB1_3_20/buf_output[5] , \SB1_3_20/buf_output[4] ,
         \SB1_3_20/buf_output[3] , \SB1_3_20/buf_output[2] ,
         \SB1_3_20/buf_output[1] , \SB1_3_20/buf_output[0] , \SB1_3_20/i3[0] ,
         \SB1_3_20/i1_5 , \SB1_3_20/i1_7 , \SB1_3_20/i1[9] , \SB1_3_20/i0_0 ,
         \SB1_3_20/i0_3 , \SB1_3_20/i0_4 , \SB1_3_20/i0[10] , \SB1_3_20/i0[9] ,
         \SB1_3_20/i0[8] , \SB1_3_20/i0[7] , \SB1_3_20/i0[6] ,
         \SB1_3_21/buf_output[5] , \SB1_3_21/buf_output[3] ,
         \SB1_3_21/buf_output[2] , \SB1_3_21/buf_output[1] ,
         \SB1_3_21/buf_output[0] , \SB1_3_21/i3[0] , \SB1_3_21/i1_5 ,
         \SB1_3_21/i1_7 , \SB1_3_21/i1[9] , \SB1_3_21/i0_0 , \SB1_3_21/i0_3 ,
         \SB1_3_21/i0_4 , \SB1_3_21/i0[10] , \SB1_3_21/i0[9] ,
         \SB1_3_21/i0[8] , \SB1_3_21/i0[7] , \SB1_3_21/i0[6] ,
         \SB1_3_22/buf_output[5] , \SB1_3_22/buf_output[4] ,
         \SB1_3_22/buf_output[3] , \SB1_3_22/buf_output[2] ,
         \SB1_3_22/buf_output[1] , \SB1_3_22/buf_output[0] , \SB1_3_22/i3[0] ,
         \SB1_3_22/i1_5 , \SB1_3_22/i1_7 , \SB1_3_22/i1[9] , \SB1_3_22/i0_0 ,
         \SB1_3_22/i0_3 , \SB1_3_22/i0_4 , \SB1_3_22/i0[10] , \SB1_3_22/i0[9] ,
         \SB1_3_22/i0[8] , \SB1_3_22/i0[7] , \SB1_3_22/i0[6] ,
         \SB1_3_23/buf_output[5] , \SB1_3_23/buf_output[4] ,
         \SB1_3_23/buf_output[3] , \SB1_3_23/buf_output[1] ,
         \SB1_3_23/buf_output[0] , \SB1_3_23/i3[0] , \SB1_3_23/i1_5 ,
         \SB1_3_23/i1_7 , \SB1_3_23/i1[9] , \SB1_3_23/i0_0 , \SB1_3_23/i0_3 ,
         \SB1_3_23/i0_4 , \SB1_3_23/i0[10] , \SB1_3_23/i0[9] ,
         \SB1_3_23/i0[8] , \SB1_3_23/i0[7] , \SB1_3_23/i0[6] ,
         \SB1_3_24/buf_output[5] , \SB1_3_24/buf_output[4] ,
         \SB1_3_24/buf_output[3] , \SB1_3_24/buf_output[2] ,
         \SB1_3_24/buf_output[1] , \SB1_3_24/buf_output[0] , \SB1_3_24/i3[0] ,
         \SB1_3_24/i1_5 , \SB1_3_24/i1_7 , \SB1_3_24/i1[9] , \SB1_3_24/i0_0 ,
         \SB1_3_24/i0_3 , \SB1_3_24/i0_4 , \SB1_3_24/i0[10] , \SB1_3_24/i0[9] ,
         \SB1_3_24/i0[8] , \SB1_3_24/i0[7] , \SB1_3_24/i0[6] ,
         \SB1_3_25/buf_output[5] , \SB1_3_25/buf_output[3] ,
         \SB1_3_25/buf_output[2] , \SB1_3_25/buf_output[1] ,
         \SB1_3_25/buf_output[0] , \SB1_3_25/i3[0] , \SB1_3_25/i1_5 ,
         \SB1_3_25/i1_7 , \SB1_3_25/i1[9] , \SB1_3_25/i0_0 , \SB1_3_25/i0_3 ,
         \SB1_3_25/i0_4 , \SB1_3_25/i0[10] , \SB1_3_25/i0[9] ,
         \SB1_3_25/i0[8] , \SB1_3_25/i0[7] , \SB1_3_25/i0[6] ,
         \SB1_3_26/buf_output[4] , \SB1_3_26/buf_output[3] ,
         \SB1_3_26/buf_output[2] , \SB1_3_26/buf_output[1] ,
         \SB1_3_26/buf_output[0] , \SB1_3_26/i3[0] , \SB1_3_26/i1_5 ,
         \SB1_3_26/i1_7 , \SB1_3_26/i1[9] , \SB1_3_26/i0_0 , \SB1_3_26/i0_3 ,
         \SB1_3_26/i0_4 , \SB1_3_26/i0[10] , \SB1_3_26/i0[9] ,
         \SB1_3_26/i0[8] , \SB1_3_26/i0[7] , \SB1_3_26/i0[6] ,
         \SB1_3_27/buf_output[5] , \SB1_3_27/buf_output[3] ,
         \SB1_3_27/buf_output[2] , \SB1_3_27/buf_output[1] ,
         \SB1_3_27/buf_output[0] , \SB1_3_27/i3[0] , \SB1_3_27/i1_5 ,
         \SB1_3_27/i1_7 , \SB1_3_27/i1[9] , \SB1_3_27/i0_0 , \SB1_3_27/i0_3 ,
         \SB1_3_27/i0_4 , \SB1_3_27/i0[10] , \SB1_3_27/i0[9] ,
         \SB1_3_27/i0[8] , \SB1_3_27/i0[7] , \SB1_3_27/i0[6] ,
         \SB1_3_28/buf_output[5] , \SB1_3_28/buf_output[4] ,
         \SB1_3_28/buf_output[3] , \SB1_3_28/buf_output[2] ,
         \SB1_3_28/buf_output[1] , \SB1_3_28/buf_output[0] , \SB1_3_28/i3[0] ,
         \SB1_3_28/i1_5 , \SB1_3_28/i1_7 , \SB1_3_28/i1[9] , \SB1_3_28/i0_0 ,
         \SB1_3_28/i0_3 , \SB1_3_28/i0_4 , \SB1_3_28/i0[10] , \SB1_3_28/i0[9] ,
         \SB1_3_28/i0[8] , \SB1_3_28/i0[7] , \SB1_3_28/i0[6] ,
         \SB1_3_29/buf_output[5] , \SB1_3_29/buf_output[3] ,
         \SB1_3_29/buf_output[2] , \SB1_3_29/buf_output[1] ,
         \SB1_3_29/buf_output[0] , \SB1_3_29/i3[0] , \SB1_3_29/i1_5 ,
         \SB1_3_29/i1_7 , \SB1_3_29/i1[9] , \SB1_3_29/i0_3 , \SB1_3_29/i0_4 ,
         \SB1_3_29/i0[10] , \SB1_3_29/i0[9] , \SB1_3_29/i0[8] ,
         \SB1_3_29/i0[7] , \SB1_3_29/i0[6] , \SB1_3_30/buf_output[5] ,
         \SB1_3_30/buf_output[3] , \SB1_3_30/buf_output[2] ,
         \SB1_3_30/buf_output[1] , \SB1_3_30/buf_output[0] , \SB1_3_30/i3[0] ,
         \SB1_3_30/i1_5 , \SB1_3_30/i1_7 , \SB1_3_30/i1[9] , \SB1_3_30/i0_0 ,
         \SB1_3_30/i0_3 , \SB1_3_30/i0_4 , \SB1_3_30/i0[10] , \SB1_3_30/i0[9] ,
         \SB1_3_30/i0[8] , \SB1_3_30/i0[7] , \SB1_3_30/i0[6] ,
         \SB1_3_31/buf_output[5] , \SB1_3_31/buf_output[4] ,
         \SB1_3_31/buf_output[3] , \SB1_3_31/buf_output[1] ,
         \SB1_3_31/buf_output[0] , \SB1_3_31/i3[0] , \SB1_3_31/i1_5 ,
         \SB1_3_31/i1_7 , \SB1_3_31/i1[9] , \SB1_3_31/i0_0 , \SB1_3_31/i0_3 ,
         \SB1_3_31/i0_4 , \SB1_3_31/i0[10] , \SB1_3_31/i0[9] ,
         \SB1_3_31/i0[8] , \SB1_3_31/i0[7] , \SB1_3_31/i0[6] ,
         \SB2_3_0/buf_output[5] , \SB2_3_0/buf_output[4] ,
         \SB2_3_0/buf_output[3] , \SB2_3_0/buf_output[2] ,
         \SB2_3_0/buf_output[1] , \SB2_3_0/buf_output[0] , \SB2_3_0/i3[0] ,
         \SB2_3_0/i1_5 , \SB2_3_0/i1_7 , \SB2_3_0/i1[9] , \SB2_3_0/i0_0 ,
         \SB2_3_0/i0_3 , \SB2_3_0/i0[10] , \SB2_3_0/i0[9] , \SB2_3_0/i0[6] ,
         \SB2_3_1/buf_output[5] , \SB2_3_1/buf_output[4] ,
         \SB2_3_1/buf_output[3] , \SB2_3_1/buf_output[1] ,
         \SB2_3_1/buf_output[0] , \SB2_3_1/i3[0] , \SB2_3_1/i1_5 ,
         \SB2_3_1/i1_7 , \SB2_3_1/i1[9] , \SB2_3_1/i0_0 , \SB2_3_1/i0_3 ,
         \SB2_3_1/i0_4 , \SB2_3_1/i0[10] , \SB2_3_1/i0[9] , \SB2_3_1/i0[8] ,
         \SB2_3_1/i0[7] , \SB2_3_1/i0[6] , \SB2_3_2/buf_output[5] ,
         \SB2_3_2/buf_output[4] , \SB2_3_2/buf_output[3] ,
         \SB2_3_2/buf_output[2] , \SB2_3_2/buf_output[1] ,
         \SB2_3_2/buf_output[0] , \SB2_3_2/i3[0] , \SB2_3_2/i1_5 ,
         \SB2_3_2/i1_7 , \SB2_3_2/i1[9] , \SB2_3_2/i0_0 , \SB2_3_2/i0_3 ,
         \SB2_3_2/i0_4 , \SB2_3_2/i0[10] , \SB2_3_2/i0[9] , \SB2_3_2/i0[7] ,
         \SB2_3_2/i0[6] , \SB2_3_3/buf_output[5] , \SB2_3_3/buf_output[4] ,
         \SB2_3_3/buf_output[3] , \SB2_3_3/buf_output[2] ,
         \SB2_3_3/buf_output[0] , \SB2_3_3/i3[0] , \SB2_3_3/i1_5 ,
         \SB2_3_3/i1_7 , \SB2_3_3/i1[9] , \SB2_3_3/i0_0 , \SB2_3_3/i0_3 ,
         \SB2_3_3/i0_4 , \SB2_3_3/i0[10] , \SB2_3_3/i0[9] , \SB2_3_3/i0[8] ,
         \SB2_3_3/i0[7] , \SB2_3_3/i0[6] , \SB2_3_4/buf_output[5] ,
         \SB2_3_4/buf_output[4] , \SB2_3_4/buf_output[3] ,
         \SB2_3_4/buf_output[2] , \SB2_3_4/buf_output[1] ,
         \SB2_3_4/buf_output[0] , \SB2_3_4/i3[0] , \SB2_3_4/i1_7 ,
         \SB2_3_4/i1[9] , \SB2_3_4/i0_0 , \SB2_3_4/i0_3 , \SB2_3_4/i0_4 ,
         \SB2_3_4/i0[10] , \SB2_3_4/i0[9] , \SB2_3_4/i0[8] , \SB2_3_4/i0[7] ,
         \SB2_3_4/i0[6] , \SB2_3_5/buf_output[5] , \SB2_3_5/buf_output[4] ,
         \SB2_3_5/buf_output[3] , \SB2_3_5/buf_output[2] ,
         \SB2_3_5/buf_output[1] , \SB2_3_5/buf_output[0] , \SB2_3_5/i3[0] ,
         \SB2_3_5/i1_5 , \SB2_3_5/i1_7 , \SB2_3_5/i0_0 , \SB2_3_5/i0_3 ,
         \SB2_3_5/i0_4 , \SB2_3_5/i0[10] , \SB2_3_5/i0[9] , \SB2_3_5/i0[8] ,
         \SB2_3_5/i0[7] , \SB2_3_5/i0[6] , \SB2_3_6/buf_output[5] ,
         \SB2_3_6/buf_output[3] , \SB2_3_6/buf_output[2] ,
         \SB2_3_6/buf_output[1] , \SB2_3_6/buf_output[0] , \SB2_3_6/i3[0] ,
         \SB2_3_6/i1_5 , \SB2_3_6/i1_7 , \SB2_3_6/i1[9] , \SB2_3_6/i0_0 ,
         \SB2_3_6/i0_3 , \SB2_3_6/i0_4 , \SB2_3_6/i0[10] , \SB2_3_6/i0[9] ,
         \SB2_3_6/i0[8] , \SB2_3_6/i0[7] , \SB2_3_6/i0[6] ,
         \SB2_3_7/buf_output[5] , \SB2_3_7/buf_output[4] ,
         \SB2_3_7/buf_output[3] , \SB2_3_7/buf_output[2] ,
         \SB2_3_7/buf_output[1] , \SB2_3_7/buf_output[0] , \SB2_3_7/i3[0] ,
         \SB2_3_7/i1_5 , \SB2_3_7/i1_7 , \SB2_3_7/i1[9] , \SB2_3_7/i0_0 ,
         \SB2_3_7/i0_3 , \SB2_3_7/i0[10] , \SB2_3_7/i0[9] , \SB2_3_7/i0[8] ,
         \SB2_3_8/buf_output[5] , \SB2_3_8/buf_output[4] ,
         \SB2_3_8/buf_output[3] , \SB2_3_8/buf_output[2] ,
         \SB2_3_8/buf_output[1] , \SB2_3_8/buf_output[0] , \SB2_3_8/i3[0] ,
         \SB2_3_8/i1_5 , \SB2_3_8/i1_7 , \SB2_3_8/i0_0 , \SB2_3_8/i0_3 ,
         \SB2_3_8/i0[10] , \SB2_3_8/i0[9] , \SB2_3_8/i0[8] , \SB2_3_8/i0[7] ,
         \SB2_3_8/i0[6] , \SB2_3_9/buf_output[5] , \SB2_3_9/buf_output[4] ,
         \SB2_3_9/buf_output[3] , \SB2_3_9/buf_output[2] ,
         \SB2_3_9/buf_output[1] , \SB2_3_9/buf_output[0] , \SB2_3_9/i3[0] ,
         \SB2_3_9/i1_5 , \SB2_3_9/i1_7 , \SB2_3_9/i1[9] , \SB2_3_9/i0_0 ,
         \SB2_3_9/i0_3 , \SB2_3_9/i0_4 , \SB2_3_9/i0[10] , \SB2_3_9/i0[9] ,
         \SB2_3_9/i0[8] , \SB2_3_9/i0[7] , \SB2_3_9/i0[6] ,
         \SB2_3_10/buf_output[5] , \SB2_3_10/buf_output[4] ,
         \SB2_3_10/buf_output[3] , \SB2_3_10/buf_output[2] ,
         \SB2_3_10/buf_output[1] , \SB2_3_10/buf_output[0] , \SB2_3_10/i3[0] ,
         \SB2_3_10/i1_5 , \SB2_3_10/i1_7 , \SB2_3_10/i1[9] , \SB2_3_10/i0_0 ,
         \SB2_3_10/i0_3 , \SB2_3_10/i0_4 , \SB2_3_10/i0[10] , \SB2_3_10/i0[9] ,
         \SB2_3_10/i0[8] , \SB2_3_10/i0[7] , \SB2_3_10/i0[6] ,
         \SB2_3_11/buf_output[5] , \SB2_3_11/buf_output[4] ,
         \SB2_3_11/buf_output[3] , \SB2_3_11/buf_output[2] ,
         \SB2_3_11/buf_output[1] , \SB2_3_11/buf_output[0] , \SB2_3_11/i3[0] ,
         \SB2_3_11/i1_7 , \SB2_3_11/i1[9] , \SB2_3_11/i0_0 , \SB2_3_11/i0_3 ,
         \SB2_3_11/i0[10] , \SB2_3_11/i0[9] , \SB2_3_11/i0[8] ,
         \SB2_3_11/i0[6] , \SB2_3_12/buf_output[5] , \SB2_3_12/buf_output[4] ,
         \SB2_3_12/buf_output[3] , \SB2_3_12/buf_output[2] ,
         \SB2_3_12/buf_output[1] , \SB2_3_12/buf_output[0] , \SB2_3_12/i3[0] ,
         \SB2_3_12/i1_5 , \SB2_3_12/i1_7 , \SB2_3_12/i1[9] , \SB2_3_12/i0_0 ,
         \SB2_3_12/i0_3 , \SB2_3_12/i0_4 , \SB2_3_12/i0[10] , \SB2_3_12/i0[7] ,
         \SB2_3_12/i0[6] , \SB2_3_13/buf_output[5] , \SB2_3_13/buf_output[4] ,
         \SB2_3_13/buf_output[3] , \SB2_3_13/buf_output[2] ,
         \SB2_3_13/buf_output[1] , \SB2_3_13/buf_output[0] , \SB2_3_13/i3[0] ,
         \SB2_3_13/i1_5 , \SB2_3_13/i1_7 , \SB2_3_13/i1[9] , \SB2_3_13/i0_0 ,
         \SB2_3_13/i0_3 , \SB2_3_13/i0[10] , \SB2_3_13/i0[9] ,
         \SB2_3_13/i0[8] , \SB2_3_13/i0[7] , \SB2_3_13/i0[6] ,
         \SB2_3_14/buf_output[5] , \SB2_3_14/buf_output[4] ,
         \SB2_3_14/buf_output[3] , \SB2_3_14/buf_output[2] ,
         \SB2_3_14/buf_output[1] , \SB2_3_14/buf_output[0] , \SB2_3_14/i3[0] ,
         \SB2_3_14/i1_5 , \SB2_3_14/i1_7 , \SB2_3_14/i1[9] , \SB2_3_14/i0_0 ,
         \SB2_3_14/i0_3 , \SB2_3_14/i0_4 , \SB2_3_14/i0[10] , \SB2_3_14/i0[9] ,
         \SB2_3_14/i0[8] , \SB2_3_14/i0[7] , \SB2_3_14/i0[6] ,
         \SB2_3_15/buf_output[5] , \SB2_3_15/buf_output[4] ,
         \SB2_3_15/buf_output[3] , \SB2_3_15/buf_output[2] ,
         \SB2_3_15/buf_output[1] , \SB2_3_15/buf_output[0] , \SB2_3_15/i3[0] ,
         \SB2_3_15/i1_5 , \SB2_3_15/i1_7 , \SB2_3_15/i1[9] , \SB2_3_15/i0_0 ,
         \SB2_3_15/i0_3 , \SB2_3_15/i0[10] , \SB2_3_15/i0[9] ,
         \SB2_3_15/i0[7] , \SB2_3_15/i0[6] , \SB2_3_16/buf_output[5] ,
         \SB2_3_16/buf_output[4] , \SB2_3_16/buf_output[3] ,
         \SB2_3_16/buf_output[2] , \SB2_3_16/buf_output[1] ,
         \SB2_3_16/buf_output[0] , \SB2_3_16/i3[0] , \SB2_3_16/i1_5 ,
         \SB2_3_16/i1_7 , \SB2_3_16/i1[9] , \SB2_3_16/i0_0 , \SB2_3_16/i0_3 ,
         \SB2_3_16/i0_4 , \SB2_3_16/i0[10] , \SB2_3_16/i0[9] ,
         \SB2_3_16/i0[8] , \SB2_3_16/i0[7] , \SB2_3_16/i0[6] ,
         \SB2_3_17/buf_output[5] , \SB2_3_17/buf_output[4] ,
         \SB2_3_17/buf_output[3] , \SB2_3_17/buf_output[2] ,
         \SB2_3_17/buf_output[1] , \SB2_3_17/buf_output[0] , \SB2_3_17/i3[0] ,
         \SB2_3_17/i1_7 , \SB2_3_17/i1[9] , \SB2_3_17/i0_0 , \SB2_3_17/i0_3 ,
         \SB2_3_17/i0_4 , \SB2_3_17/i0[10] , \SB2_3_17/i0[9] ,
         \SB2_3_17/i0[8] , \SB2_3_17/i0[7] , \SB2_3_17/i0[6] ,
         \SB2_3_18/buf_output[5] , \SB2_3_18/buf_output[4] ,
         \SB2_3_18/buf_output[3] , \SB2_3_18/buf_output[2] ,
         \SB2_3_18/buf_output[1] , \SB2_3_18/buf_output[0] , \SB2_3_18/i3[0] ,
         \SB2_3_18/i1_5 , \SB2_3_18/i1_7 , \SB2_3_18/i1[9] , \SB2_3_18/i0_0 ,
         \SB2_3_18/i0_3 , \SB2_3_18/i0_4 , \SB2_3_18/i0[10] , \SB2_3_18/i0[9] ,
         \SB2_3_18/i0[8] , \SB2_3_18/i0[7] , \SB2_3_18/i0[6] ,
         \SB2_3_19/buf_output[5] , \SB2_3_19/buf_output[4] ,
         \SB2_3_19/buf_output[3] , \SB2_3_19/buf_output[2] ,
         \SB2_3_19/buf_output[1] , \SB2_3_19/i3[0] , \SB2_3_19/i1_5 ,
         \SB2_3_19/i1_7 , \SB2_3_19/i0_0 , \SB2_3_19/i0_3 , \SB2_3_19/i0_4 ,
         \SB2_3_19/i0[10] , \SB2_3_19/i0[9] , \SB2_3_19/i0[8] ,
         \SB2_3_19/i0[7] , \SB2_3_19/i0[6] , \SB2_3_20/buf_output[5] ,
         \SB2_3_20/buf_output[4] , \SB2_3_20/buf_output[3] ,
         \SB2_3_20/buf_output[2] , \SB2_3_20/buf_output[1] ,
         \SB2_3_20/buf_output[0] , \SB2_3_20/i3[0] , \SB2_3_20/i1_5 ,
         \SB2_3_20/i1_7 , \SB2_3_20/i1[9] , \SB2_3_20/i0_0 , \SB2_3_20/i0_3 ,
         \SB2_3_20/i0_4 , \SB2_3_20/i0[10] , \SB2_3_20/i0[9] ,
         \SB2_3_20/i0[8] , \SB2_3_20/i0[7] , \SB2_3_20/i0[6] ,
         \SB2_3_21/buf_output[5] , \SB2_3_21/buf_output[4] ,
         \SB2_3_21/buf_output[3] , \SB2_3_21/buf_output[2] ,
         \SB2_3_21/buf_output[1] , \SB2_3_21/i3[0] , \SB2_3_21/i1_5 ,
         \SB2_3_21/i1_7 , \SB2_3_21/i1[9] , \SB2_3_21/i0_0 , \SB2_3_21/i0_3 ,
         \SB2_3_21/i0[10] , \SB2_3_21/i0[9] , \SB2_3_21/i0[8] ,
         \SB2_3_21/i0[7] , \SB2_3_21/i0[6] , \SB2_3_22/buf_output[5] ,
         \SB2_3_22/buf_output[4] , \SB2_3_22/buf_output[3] ,
         \SB2_3_22/buf_output[2] , \SB2_3_22/buf_output[1] ,
         \SB2_3_22/buf_output[0] , \SB2_3_22/i3[0] , \SB2_3_22/i1_5 ,
         \SB2_3_22/i1_7 , \SB2_3_22/i1[9] , \SB2_3_22/i0_0 , \SB2_3_22/i0_3 ,
         \SB2_3_22/i0_4 , \SB2_3_22/i0[10] , \SB2_3_22/i0[9] ,
         \SB2_3_22/i0[8] , \SB2_3_22/i0[7] , \SB2_3_22/i0[6] ,
         \SB2_3_23/buf_output[5] , \SB2_3_23/buf_output[4] ,
         \SB2_3_23/buf_output[3] , \SB2_3_23/buf_output[2] ,
         \SB2_3_23/buf_output[1] , \SB2_3_23/buf_output[0] , \SB2_3_23/i3[0] ,
         \SB2_3_23/i1_5 , \SB2_3_23/i1_7 , \SB2_3_23/i1[9] , \SB2_3_23/i0_0 ,
         \SB2_3_23/i0_3 , \SB2_3_23/i0_4 , \SB2_3_23/i0[10] , \SB2_3_23/i0[9] ,
         \SB2_3_23/i0[8] , \SB2_3_23/i0[7] , \SB2_3_23/i0[6] ,
         \SB2_3_24/buf_output[5] , \SB2_3_24/buf_output[4] ,
         \SB2_3_24/buf_output[3] , \SB2_3_24/buf_output[2] ,
         \SB2_3_24/buf_output[1] , \SB2_3_24/buf_output[0] , \SB2_3_24/i3[0] ,
         \SB2_3_24/i1_5 , \SB2_3_24/i1_7 , \SB2_3_24/i1[9] , \SB2_3_24/i0_0 ,
         \SB2_3_24/i0_3 , \SB2_3_24/i0_4 , \SB2_3_24/i0[9] , \SB2_3_24/i0[6] ,
         \SB2_3_25/buf_output[5] , \SB2_3_25/buf_output[4] ,
         \SB2_3_25/buf_output[3] , \SB2_3_25/buf_output[2] ,
         \SB2_3_25/buf_output[1] , \SB2_3_25/buf_output[0] , \SB2_3_25/i3[0] ,
         \SB2_3_25/i1_5 , \SB2_3_25/i1_7 , \SB2_3_25/i1[9] , \SB2_3_25/i0_0 ,
         \SB2_3_25/i0_3 , \SB2_3_25/i0[10] , \SB2_3_25/i0[9] ,
         \SB2_3_25/i0[8] , \SB2_3_25/i0[7] , \SB2_3_25/i0[6] ,
         \SB2_3_26/buf_output[5] , \SB2_3_26/buf_output[4] ,
         \SB2_3_26/buf_output[3] , \SB2_3_26/buf_output[2] ,
         \SB2_3_26/buf_output[1] , \SB2_3_26/buf_output[0] , \SB2_3_26/i3[0] ,
         \SB2_3_26/i1_5 , \SB2_3_26/i1_7 , \SB2_3_26/i1[9] , \SB2_3_26/i0_0 ,
         \SB2_3_26/i0_3 , \SB2_3_26/i0_4 , \SB2_3_26/i0[9] , \SB2_3_26/i0[7] ,
         \SB2_3_26/i0[6] , \SB2_3_27/buf_output[5] , \SB2_3_27/buf_output[4] ,
         \SB2_3_27/buf_output[3] , \SB2_3_27/buf_output[2] ,
         \SB2_3_27/buf_output[1] , \SB2_3_27/buf_output[0] , \SB2_3_27/i3[0] ,
         \SB2_3_27/i1_5 , \SB2_3_27/i1_7 , \SB2_3_27/i1[9] , \SB2_3_27/i0_0 ,
         \SB2_3_27/i0_3 , \SB2_3_27/i0_4 , \SB2_3_27/i0[10] , \SB2_3_27/i0[8] ,
         \SB2_3_27/i0[7] , \SB2_3_28/buf_output[5] , \SB2_3_28/buf_output[4] ,
         \SB2_3_28/buf_output[3] , \SB2_3_28/buf_output[2] ,
         \SB2_3_28/buf_output[1] , \SB2_3_28/buf_output[0] , \SB2_3_28/i3[0] ,
         \SB2_3_28/i1_5 , \SB2_3_28/i1_7 , \SB2_3_28/i0_0 , \SB2_3_28/i0_3 ,
         \SB2_3_28/i0[9] , \SB2_3_28/i0[8] , \SB2_3_28/i0[7] ,
         \SB2_3_28/i0[6] , \SB2_3_29/buf_output[5] , \SB2_3_29/buf_output[4] ,
         \SB2_3_29/buf_output[3] , \SB2_3_29/buf_output[2] ,
         \SB2_3_29/buf_output[1] , \SB2_3_29/buf_output[0] , \SB2_3_29/i3[0] ,
         \SB2_3_29/i1_5 , \SB2_3_29/i1_7 , \SB2_3_29/i1[9] , \SB2_3_29/i0_0 ,
         \SB2_3_29/i0_3 , \SB2_3_29/i0[10] , \SB2_3_29/i0[9] ,
         \SB2_3_29/i0[8] , \SB2_3_29/i0[7] , \SB2_3_29/i0[6] ,
         \SB2_3_30/buf_output[5] , \SB2_3_30/buf_output[4] ,
         \SB2_3_30/buf_output[3] , \SB2_3_30/buf_output[2] ,
         \SB2_3_30/buf_output[1] , \SB2_3_30/buf_output[0] , \SB2_3_30/i3[0] ,
         \SB2_3_30/i1_5 , \SB2_3_30/i1_7 , \SB2_3_30/i1[9] , \SB2_3_30/i0_0 ,
         \SB2_3_30/i0_3 , \SB2_3_30/i0_4 , \SB2_3_30/i0[10] , \SB2_3_30/i0[9] ,
         \SB2_3_30/i0[8] , \SB2_3_30/i0[7] , \SB2_3_30/i0[6] ,
         \SB2_3_31/buf_output[5] , \SB2_3_31/buf_output[4] ,
         \SB2_3_31/buf_output[3] , \SB2_3_31/buf_output[2] ,
         \SB2_3_31/buf_output[1] , \SB2_3_31/buf_output[0] , \SB2_3_31/i3[0] ,
         \SB2_3_31/i1_5 , \SB2_3_31/i1_7 , \SB2_3_31/i1[9] , \SB2_3_31/i0_0 ,
         \SB2_3_31/i0_3 , \SB2_3_31/i0_4 , \SB2_3_31/i0[10] , \SB2_3_31/i0[9] ,
         \SB2_3_31/i0[8] , \SB2_3_31/i0[7] , \SB2_3_31/i0[6] ,
         \SB3_0/buf_output[5] , \SB3_0/buf_output[4] , \SB3_0/buf_output[3] ,
         \SB3_0/buf_output[2] , \SB3_0/buf_output[1] , \SB3_0/buf_output[0] ,
         \SB3_0/i3[0] , \SB3_0/i1_5 , \SB3_0/i1_7 , \SB3_0/i1[9] ,
         \SB3_0/i0_0 , \SB3_0/i0_3 , \SB3_0/i0_4 , \SB3_0/i0[10] ,
         \SB3_0/i0[9] , \SB3_0/i0[8] , \SB3_0/i0[7] , \SB3_0/i0[6] ,
         \SB3_1/buf_output[5] , \SB3_1/buf_output[4] , \SB3_1/buf_output[2] ,
         \SB3_1/buf_output[1] , \SB3_1/buf_output[0] , \SB3_1/i3[0] ,
         \SB3_1/i1_5 , \SB3_1/i1_7 , \SB3_1/i0_0 , \SB3_1/i0_3 , \SB3_1/i0_4 ,
         \SB3_1/i0[10] , \SB3_1/i0[9] , \SB3_1/i0[8] , \SB3_1/i0[7] ,
         \SB3_1/i0[6] , \SB3_2/buf_output[5] , \SB3_2/buf_output[4] ,
         \SB3_2/buf_output[3] , \SB3_2/buf_output[2] , \SB3_2/buf_output[1] ,
         \SB3_2/buf_output[0] , \SB3_2/i3[0] , \SB3_2/i1_5 , \SB3_2/i1_7 ,
         \SB3_2/i1[9] , \SB3_2/i0_0 , \SB3_2/i0_3 , \SB3_2/i0_4 ,
         \SB3_2/i0[10] , \SB3_2/i0[9] , \SB3_2/i0[8] , \SB3_2/i0[7] ,
         \SB3_2/i0[6] , \SB3_3/buf_output[5] , \SB3_3/buf_output[4] ,
         \SB3_3/buf_output[3] , \SB3_3/buf_output[2] , \SB3_3/buf_output[1] ,
         \SB3_3/buf_output[0] , \SB3_3/i3[0] , \SB3_3/i1_5 , \SB3_3/i1_7 ,
         \SB3_3/i1[9] , \SB3_3/i0_0 , \SB3_3/i0_3 , \SB3_3/i0_4 ,
         \SB3_3/i0[10] , \SB3_3/i0[9] , \SB3_3/i0[8] , \SB3_3/i0[7] ,
         \SB3_3/i0[6] , \SB3_4/buf_output[5] , \SB3_4/buf_output[4] ,
         \SB3_4/buf_output[3] , \SB3_4/buf_output[2] , \SB3_4/buf_output[1] ,
         \SB3_4/buf_output[0] , \SB3_4/i3[0] , \SB3_4/i1_7 , \SB3_4/i1[9] ,
         \SB3_4/i0_0 , \SB3_4/i0_3 , \SB3_4/i0_4 , \SB3_4/i0[10] ,
         \SB3_4/i0[9] , \SB3_4/i0[8] , \SB3_4/i0[7] , \SB3_4/i0[6] ,
         \SB3_5/buf_output[5] , \SB3_5/buf_output[4] , \SB3_5/buf_output[3] ,
         \SB3_5/buf_output[2] , \SB3_5/buf_output[1] , \SB3_5/buf_output[0] ,
         \SB3_5/i3[0] , \SB3_5/i1_5 , \SB3_5/i1_7 , \SB3_5/i1[9] ,
         \SB3_5/i0_0 , \SB3_5/i0_3 , \SB3_5/i0_4 , \SB3_5/i0[10] ,
         \SB3_5/i0[9] , \SB3_5/i0[8] , \SB3_5/i0[7] , \SB3_5/i0[6] ,
         \SB3_6/buf_output[5] , \SB3_6/buf_output[4] , \SB3_6/buf_output[3] ,
         \SB3_6/buf_output[2] , \SB3_6/buf_output[1] , \SB3_6/buf_output[0] ,
         \SB3_6/i3[0] , \SB3_6/i1_5 , \SB3_6/i1_7 , \SB3_6/i1[9] ,
         \SB3_6/i0_0 , \SB3_6/i0[10] , \SB3_6/i0[9] , \SB3_6/i0[8] ,
         \SB3_6/i0[7] , \SB3_6/i0[6] , \SB3_7/buf_output[5] ,
         \SB3_7/buf_output[4] , \SB3_7/buf_output[3] , \SB3_7/buf_output[2] ,
         \SB3_7/buf_output[1] , \SB3_7/buf_output[0] , \SB3_7/i3[0] ,
         \SB3_7/i1_7 , \SB3_7/i1[9] , \SB3_7/i0_0 , \SB3_7/i0_3 , \SB3_7/i0_4 ,
         \SB3_7/i0[10] , \SB3_7/i0[9] , \SB3_7/i0[8] , \SB3_7/i0[7] ,
         \SB3_7/i0[6] , \SB3_8/buf_output[5] , \SB3_8/buf_output[4] ,
         \SB3_8/buf_output[2] , \SB3_8/buf_output[1] , \SB3_8/buf_output[0] ,
         \SB3_8/i3[0] , \SB3_8/i1_5 , \SB3_8/i1_7 , \SB3_8/i1[9] ,
         \SB3_8/i0_0 , \SB3_8/i0_3 , \SB3_8/i0_4 , \SB3_8/i0[10] ,
         \SB3_8/i0[9] , \SB3_8/i0[8] , \SB3_8/i0[7] , \SB3_8/i0[6] ,
         \SB3_9/buf_output[5] , \SB3_9/buf_output[4] , \SB3_9/buf_output[3] ,
         \SB3_9/buf_output[2] , \SB3_9/buf_output[1] , \SB3_9/buf_output[0] ,
         \SB3_9/i3[0] , \SB3_9/i1_5 , \SB3_9/i1_7 , \SB3_9/i1[9] ,
         \SB3_9/i0_0 , \SB3_9/i0_3 , \SB3_9/i0_4 , \SB3_9/i0[10] ,
         \SB3_9/i0[9] , \SB3_9/i0[8] , \SB3_9/i0[7] , \SB3_9/i0[6] ,
         \SB3_10/buf_output[5] , \SB3_10/buf_output[4] ,
         \SB3_10/buf_output[3] , \SB3_10/buf_output[2] ,
         \SB3_10/buf_output[1] , \SB3_10/buf_output[0] , \SB3_10/i3[0] ,
         \SB3_10/i1_5 , \SB3_10/i1_7 , \SB3_10/i1[9] , \SB3_10/i0_0 ,
         \SB3_10/i0_3 , \SB3_10/i0_4 , \SB3_10/i0[10] , \SB3_10/i0[9] ,
         \SB3_10/i0[8] , \SB3_10/i0[7] , \SB3_10/i0[6] ,
         \SB3_11/buf_output[5] , \SB3_11/buf_output[4] ,
         \SB3_11/buf_output[3] , \SB3_11/buf_output[2] ,
         \SB3_11/buf_output[1] , \SB3_11/buf_output[0] , \SB3_11/i3[0] ,
         \SB3_11/i1_7 , \SB3_11/i1[9] , \SB3_11/i0_0 , \SB3_11/i0_3 ,
         \SB3_11/i0_4 , \SB3_11/i0[10] , \SB3_11/i0[9] , \SB3_11/i0[8] ,
         \SB3_11/i0[7] , \SB3_11/i0[6] , \SB3_12/buf_output[5] ,
         \SB3_12/buf_output[4] , \SB3_12/buf_output[3] ,
         \SB3_12/buf_output[2] , \SB3_12/buf_output[1] ,
         \SB3_12/buf_output[0] , \SB3_12/i3[0] , \SB3_12/i1_5 , \SB3_12/i1_7 ,
         \SB3_12/i1[9] , \SB3_12/i0_0 , \SB3_12/i0_3 , \SB3_12/i0_4 ,
         \SB3_12/i0[10] , \SB3_12/i0[9] , \SB3_12/i0[8] , \SB3_12/i0[7] ,
         \SB3_12/i0[6] , \SB3_13/buf_output[5] , \SB3_13/buf_output[4] ,
         \SB3_13/buf_output[3] , \SB3_13/buf_output[2] ,
         \SB3_13/buf_output[1] , \SB3_13/buf_output[0] , \SB3_13/i3[0] ,
         \SB3_13/i1_5 , \SB3_13/i1_7 , \SB3_13/i1[9] , \SB3_13/i0_3 ,
         \SB3_13/i0_4 , \SB3_13/i0[10] , \SB3_13/i0[9] , \SB3_13/i0[8] ,
         \SB3_13/i0[7] , \SB3_13/i0[6] , \SB3_14/buf_output[5] ,
         \SB3_14/buf_output[4] , \SB3_14/buf_output[3] ,
         \SB3_14/buf_output[2] , \SB3_14/buf_output[1] ,
         \SB3_14/buf_output[0] , \SB3_14/i3[0] , \SB3_14/i1_5 , \SB3_14/i1_7 ,
         \SB3_14/i1[9] , \SB3_14/i0_0 , \SB3_14/i0_3 , \SB3_14/i0_4 ,
         \SB3_14/i0[10] , \SB3_14/i0[9] , \SB3_14/i0[8] , \SB3_14/i0[7] ,
         \SB3_14/i0[6] , \SB3_15/buf_output[5] , \SB3_15/buf_output[4] ,
         \SB3_15/buf_output[3] , \SB3_15/buf_output[2] ,
         \SB3_15/buf_output[1] , \SB3_15/buf_output[0] , \SB3_15/i3[0] ,
         \SB3_15/i1_5 , \SB3_15/i1_7 , \SB3_15/i1[9] , \SB3_15/i0_0 ,
         \SB3_15/i0_3 , \SB3_15/i0_4 , \SB3_15/i0[10] , \SB3_15/i0[9] ,
         \SB3_15/i0[8] , \SB3_15/i0[7] , \SB3_15/i0[6] ,
         \SB3_16/buf_output[5] , \SB3_16/buf_output[4] ,
         \SB3_16/buf_output[2] , \SB3_16/buf_output[1] ,
         \SB3_16/buf_output[0] , \SB3_16/i3[0] , \SB3_16/i1_5 , \SB3_16/i1_7 ,
         \SB3_16/i1[9] , \SB3_16/i0_0 , \SB3_16/i0_3 , \SB3_16/i0_4 ,
         \SB3_16/i0[10] , \SB3_16/i0[9] , \SB3_16/i0[8] , \SB3_16/i0[7] ,
         \SB3_16/i0[6] , \SB3_17/buf_output[5] , \SB3_17/buf_output[4] ,
         \SB3_17/buf_output[3] , \SB3_17/buf_output[2] ,
         \SB3_17/buf_output[1] , \SB3_17/buf_output[0] , \SB3_17/i3[0] ,
         \SB3_17/i1_5 , \SB3_17/i1_7 , \SB3_17/i1[9] , \SB3_17/i0_0 ,
         \SB3_17/i0_3 , \SB3_17/i0_4 , \SB3_17/i0[10] , \SB3_17/i0[9] ,
         \SB3_17/i0[8] , \SB3_17/i0[7] , \SB3_17/i0[6] ,
         \SB3_18/buf_output[5] , \SB3_18/buf_output[4] ,
         \SB3_18/buf_output[3] , \SB3_18/buf_output[2] ,
         \SB3_18/buf_output[1] , \SB3_18/buf_output[0] , \SB3_18/i3[0] ,
         \SB3_18/i1_5 , \SB3_18/i1_7 , \SB3_18/i1[9] , \SB3_18/i0_0 ,
         \SB3_18/i0_3 , \SB3_18/i0_4 , \SB3_18/i0[10] , \SB3_18/i0[9] ,
         \SB3_18/i0[8] , \SB3_18/i0[7] , \SB3_18/i0[6] ,
         \SB3_19/buf_output[5] , \SB3_19/buf_output[4] ,
         \SB3_19/buf_output[3] , \SB3_19/buf_output[2] ,
         \SB3_19/buf_output[1] , \SB3_19/buf_output[0] , \SB3_19/i3[0] ,
         \SB3_19/i1_5 , \SB3_19/i1_7 , \SB3_19/i1[9] , \SB3_19/i0_0 ,
         \SB3_19/i0_3 , \SB3_19/i0_4 , \SB3_19/i0[10] , \SB3_19/i0[9] ,
         \SB3_19/i0[8] , \SB3_19/i0[7] , \SB3_19/i0[6] ,
         \SB3_20/buf_output[5] , \SB3_20/buf_output[4] ,
         \SB3_20/buf_output[3] , \SB3_20/buf_output[2] ,
         \SB3_20/buf_output[1] , \SB3_20/buf_output[0] , \SB3_20/i3[0] ,
         \SB3_20/i1_5 , \SB3_20/i1_7 , \SB3_20/i1[9] , \SB3_20/i0_0 ,
         \SB3_20/i0_3 , \SB3_20/i0_4 , \SB3_20/i0[10] , \SB3_20/i0[9] ,
         \SB3_20/i0[8] , \SB3_20/i0[7] , \SB3_20/i0[6] ,
         \SB3_21/buf_output[4] , \SB3_21/buf_output[3] ,
         \SB3_21/buf_output[2] , \SB3_21/buf_output[1] ,
         \SB3_21/buf_output[0] , \SB3_21/i3[0] , \SB3_21/i1_5 , \SB3_21/i1_7 ,
         \SB3_21/i1[9] , \SB3_21/i0_0 , \SB3_21/i0_3 , \SB3_21/i0_4 ,
         \SB3_21/i0[10] , \SB3_21/i0[9] , \SB3_21/i0[8] , \SB3_21/i0[7] ,
         \SB3_21/i0[6] , \SB3_22/buf_output[5] , \SB3_22/buf_output[4] ,
         \SB3_22/buf_output[3] , \SB3_22/buf_output[2] ,
         \SB3_22/buf_output[1] , \SB3_22/buf_output[0] , \SB3_22/i3[0] ,
         \SB3_22/i1_5 , \SB3_22/i1_7 , \SB3_22/i1[9] , \SB3_22/i0_0 ,
         \SB3_22/i0_3 , \SB3_22/i0_4 , \SB3_22/i0[10] , \SB3_22/i0[9] ,
         \SB3_22/i0[8] , \SB3_22/i0[7] , \SB3_22/i0[6] ,
         \SB3_23/buf_output[5] , \SB3_23/buf_output[4] ,
         \SB3_23/buf_output[3] , \SB3_23/buf_output[2] ,
         \SB3_23/buf_output[1] , \SB3_23/buf_output[0] , \SB3_23/i3[0] ,
         \SB3_23/i1_5 , \SB3_23/i1_7 , \SB3_23/i1[9] , \SB3_23/i0_0 ,
         \SB3_23/i0_3 , \SB3_23/i0_4 , \SB3_23/i0[10] , \SB3_23/i0[9] ,
         \SB3_23/i0[8] , \SB3_23/i0[7] , \SB3_23/i0[6] ,
         \SB3_24/buf_output[5] , \SB3_24/buf_output[4] ,
         \SB3_24/buf_output[3] , \SB3_24/buf_output[2] ,
         \SB3_24/buf_output[1] , \SB3_24/buf_output[0] , \SB3_24/i3[0] ,
         \SB3_24/i1_5 , \SB3_24/i1_7 , \SB3_24/i1[9] , \SB3_24/i0_0 ,
         \SB3_24/i0_3 , \SB3_24/i0_4 , \SB3_24/i0[10] , \SB3_24/i0[9] ,
         \SB3_24/i0[8] , \SB3_24/i0[7] , \SB3_24/i0[6] ,
         \SB3_25/buf_output[5] , \SB3_25/buf_output[4] ,
         \SB3_25/buf_output[3] , \SB3_25/buf_output[2] ,
         \SB3_25/buf_output[1] , \SB3_25/buf_output[0] , \SB3_25/i3[0] ,
         \SB3_25/i1_5 , \SB3_25/i1_7 , \SB3_25/i1[9] , \SB3_25/i0_0 ,
         \SB3_25/i0_3 , \SB3_25/i0_4 , \SB3_25/i0[10] , \SB3_25/i0[9] ,
         \SB3_25/i0[8] , \SB3_25/i0[7] , \SB3_25/i0[6] ,
         \SB3_26/buf_output[5] , \SB3_26/buf_output[4] ,
         \SB3_26/buf_output[3] , \SB3_26/buf_output[2] ,
         \SB3_26/buf_output[1] , \SB3_26/buf_output[0] , \SB3_26/i3[0] ,
         \SB3_26/i1_5 , \SB3_26/i1_7 , \SB3_26/i1[9] , \SB3_26/i0_0 ,
         \SB3_26/i0_3 , \SB3_26/i0_4 , \SB3_26/i0[10] , \SB3_26/i0[9] ,
         \SB3_26/i0[8] , \SB3_26/i0[7] , \SB3_26/i0[6] ,
         \SB3_27/buf_output[5] , \SB3_27/buf_output[4] ,
         \SB3_27/buf_output[3] , \SB3_27/buf_output[2] ,
         \SB3_27/buf_output[1] , \SB3_27/buf_output[0] , \SB3_27/i3[0] ,
         \SB3_27/i1_5 , \SB3_27/i1_7 , \SB3_27/i0_0 , \SB3_27/i0_3 ,
         \SB3_27/i0_4 , \SB3_27/i0[10] , \SB3_27/i0[9] , \SB3_27/i0[8] ,
         \SB3_27/i0[7] , \SB3_27/i0[6] , \SB3_28/buf_output[4] ,
         \SB3_28/buf_output[3] , \SB3_28/buf_output[2] ,
         \SB3_28/buf_output[1] , \SB3_28/buf_output[0] , \SB3_28/i3[0] ,
         \SB3_28/i1_5 , \SB3_28/i1_7 , \SB3_28/i1[9] , \SB3_28/i0_0 ,
         \SB3_28/i0_3 , \SB3_28/i0_4 , \SB3_28/i0[10] , \SB3_28/i0[9] ,
         \SB3_28/i0[8] , \SB3_28/i0[7] , \SB3_28/i0[6] ,
         \SB3_29/buf_output[5] , \SB3_29/buf_output[4] ,
         \SB3_29/buf_output[3] , \SB3_29/buf_output[2] ,
         \SB3_29/buf_output[1] , \SB3_29/buf_output[0] , \SB3_29/i3[0] ,
         \SB3_29/i1_5 , \SB3_29/i1_7 , \SB3_29/i1[9] , \SB3_29/i0_0 ,
         \SB3_29/i0_3 , \SB3_29/i0_4 , \SB3_29/i0[10] , \SB3_29/i0[9] ,
         \SB3_29/i0[8] , \SB3_29/i0[7] , \SB3_29/i0[6] ,
         \SB3_30/buf_output[5] , \SB3_30/buf_output[3] ,
         \SB3_30/buf_output[2] , \SB3_30/buf_output[1] ,
         \SB3_30/buf_output[0] , \SB3_30/i3[0] , \SB3_30/i1_5 , \SB3_30/i1_7 ,
         \SB3_30/i1[9] , \SB3_30/i0_0 , \SB3_30/i0_3 , \SB3_30/i0_4 ,
         \SB3_30/i0[10] , \SB3_30/i0[9] , \SB3_30/i0[8] , \SB3_30/i0[7] ,
         \SB3_30/i0[6] , \SB3_31/buf_output[5] , \SB3_31/buf_output[4] ,
         \SB3_31/buf_output[3] , \SB3_31/buf_output[2] ,
         \SB3_31/buf_output[1] , \SB3_31/buf_output[0] , \SB3_31/i3[0] ,
         \SB3_31/i1_5 , \SB3_31/i1_7 , \SB3_31/i1[9] , \SB3_31/i0_0 ,
         \SB3_31/i0_3 , \SB3_31/i0_4 , \SB3_31/i0[10] , \SB3_31/i0[9] ,
         \SB3_31/i0[8] , \SB3_31/i0[7] , \SB3_31/i0[6] , \SB4_0/i3[0] ,
         \SB4_0/i1_5 , \SB4_0/i1_7 , \SB4_0/i0_3 , \SB4_0/i0_4 ,
         \SB4_0/i0[10] , \SB4_0/i0[9] , \SB4_0/i0[8] , \SB4_0/i0[7] ,
         \SB4_0/i0[6] , \SB4_1/i3[0] , \SB4_1/i1_5 , \SB4_1/i1_7 ,
         \SB4_1/i1[9] , \SB4_1/i0_0 , \SB4_1/i0_3 , \SB4_1/i0_4 ,
         \SB4_1/i0[10] , \SB4_1/i0[9] , \SB4_1/i0[8] , \SB4_1/i0[7] ,
         \SB4_1/i0[6] , \SB4_2/i3[0] , \SB4_2/i1_5 , \SB4_2/i1_7 ,
         \SB4_2/i1[9] , \SB4_2/i0_0 , \SB4_2/i0_3 , \SB4_2/i0_4 ,
         \SB4_2/i0[10] , \SB4_2/i0[9] , \SB4_2/i0[8] , \SB4_2/i0[7] ,
         \SB4_2/i0[6] , \SB4_3/i3[0] , \SB4_3/i1_5 , \SB4_3/i1_7 ,
         \SB4_3/i0_3 , \SB4_3/i0_4 , \SB4_3/i0[9] , \SB4_3/i0[7] ,
         \SB4_3/i0[6] , \SB4_4/i3[0] , \SB4_4/i1_5 , \SB4_4/i1_7 ,
         \SB4_4/i0_3 , \SB4_4/i0_4 , \SB4_4/i0[10] , \SB4_4/i0[9] ,
         \SB4_4/i0[8] , \SB4_4/i0[7] , \SB4_4/i0[6] , \SB4_5/i3[0] ,
         \SB4_5/i1_5 , \SB4_5/i1_7 , \SB4_5/i1[9] , \SB4_5/i0_0 , \SB4_5/i0_3 ,
         \SB4_5/i0_4 , \SB4_5/i0[10] , \SB4_5/i0[9] , \SB4_5/i0[8] ,
         \SB4_5/i0[7] , \SB4_5/i0[6] , \SB4_6/i3[0] , \SB4_6/i1_5 ,
         \SB4_6/i1_7 , \SB4_6/i1[9] , \SB4_6/i0_0 , \SB4_6/i0_3 , \SB4_6/i0_4 ,
         \SB4_6/i0[10] , \SB4_6/i0[9] , \SB4_6/i0[7] , \SB4_6/i0[6] ,
         \SB4_7/i3[0] , \SB4_7/i1_5 , \SB4_7/i1_7 , \SB4_7/i1[9] ,
         \SB4_7/i0_0 , \SB4_7/i0_3 , \SB4_7/i0_4 , \SB4_7/i0[10] ,
         \SB4_7/i0[9] , \SB4_7/i0[8] , \SB4_7/i0[7] , \SB4_7/i0[6] ,
         \SB4_8/i3[0] , \SB4_8/i1_5 , \SB4_8/i1_7 , \SB4_8/i1[9] ,
         \SB4_8/i0_0 , \SB4_8/i0_3 , \SB4_8/i0_4 , \SB4_8/i0[10] ,
         \SB4_8/i0[9] , \SB4_8/i0[8] , \SB4_8/i0[7] , \SB4_8/i0[6] ,
         \SB4_9/i3[0] , \SB4_9/i1_5 , \SB4_9/i1_7 , \SB4_9/i1[9] ,
         \SB4_9/i0_0 , \SB4_9/i0_3 , \SB4_9/i0_4 , \SB4_9/i0[10] ,
         \SB4_9/i0[9] , \SB4_9/i0[8] , \SB4_9/i0[7] , \SB4_9/i0[6] ,
         \SB4_10/i3[0] , \SB4_10/i1_5 , \SB4_10/i1_7 , \SB4_10/i0_3 ,
         \SB4_10/i0_4 , \SB4_10/i0[10] , \SB4_10/i0[9] , \SB4_10/i0[8] ,
         \SB4_10/i0[7] , \SB4_10/i0[6] , \SB4_11/i3[0] , \SB4_11/i1_7 ,
         \SB4_11/i1[9] , \SB4_11/i0_0 , \SB4_11/i0_3 , \SB4_11/i0_4 ,
         \SB4_11/i0[10] , \SB4_11/i0[9] , \SB4_11/i0[8] , \SB4_11/i0[7] ,
         \SB4_11/i0[6] , \SB4_12/i3[0] , \SB4_12/i1_5 , \SB4_12/i1_7 ,
         \SB4_12/i1[9] , \SB4_12/i0_0 , \SB4_12/i0_3 , \SB4_12/i0_4 ,
         \SB4_12/i0[10] , \SB4_12/i0[9] , \SB4_12/i0[8] , \SB4_12/i0[7] ,
         \SB4_12/i0[6] , \SB4_13/i3[0] , \SB4_13/i1_5 , \SB4_13/i1_7 ,
         \SB4_13/i1[9] , \SB4_13/i0_0 , \SB4_13/i0_3 , \SB4_13/i0_4 ,
         \SB4_13/i0[10] , \SB4_13/i0[9] , \SB4_13/i0[7] , \SB4_13/i0[6] ,
         \SB4_14/i3[0] , \SB4_14/i1_5 , \SB4_14/i1_7 , \SB4_14/i1[9] ,
         \SB4_14/i0_0 , \SB4_14/i0_3 , \SB4_14/i0_4 , \SB4_14/i0[10] ,
         \SB4_14/i0[9] , \SB4_14/i0[8] , \SB4_14/i0[7] , \SB4_14/i0[6] ,
         \SB4_15/i3[0] , \SB4_15/i1_5 , \SB4_15/i1_7 , \SB4_15/i1[9] ,
         \SB4_15/i0_0 , \SB4_15/i0_3 , \SB4_15/i0_4 , \SB4_15/i0[10] ,
         \SB4_15/i0[9] , \SB4_15/i0[8] , \SB4_15/i0[7] , \SB4_15/i0[6] ,
         \SB4_16/i3[0] , \SB4_16/i1_5 , \SB4_16/i1_7 , \SB4_16/i1[9] ,
         \SB4_16/i0_0 , \SB4_16/i0_3 , \SB4_16/i0_4 , \SB4_16/i0[10] ,
         \SB4_16/i0[9] , \SB4_16/i0[8] , \SB4_16/i0[7] , \SB4_16/i0[6] ,
         \SB4_17/i3[0] , \SB4_17/i1_5 , \SB4_17/i1_7 , \SB4_17/i1[9] ,
         \SB4_17/i0_0 , \SB4_17/i0_3 , \SB4_17/i0_4 , \SB4_17/i0[10] ,
         \SB4_17/i0[9] , \SB4_17/i0[7] , \SB4_17/i0[6] , \SB4_18/i3[0] ,
         \SB4_18/i1_5 , \SB4_18/i1_7 , \SB4_18/i1[9] , \SB4_18/i0_0 ,
         \SB4_18/i0_3 , \SB4_18/i0_4 , \SB4_18/i0[10] , \SB4_18/i0[9] ,
         \SB4_18/i0[7] , \SB4_18/i0[6] , \SB4_19/i3[0] , \SB4_19/i1_5 ,
         \SB4_19/i1_7 , \SB4_19/i1[9] , \SB4_19/i0_0 , \SB4_19/i0_3 ,
         \SB4_19/i0_4 , \SB4_19/i0[9] , \SB4_19/i0[7] , \SB4_19/i0[6] ,
         \SB4_20/i3[0] , \SB4_20/i1_7 , \SB4_20/i1[9] , \SB4_20/i0_0 ,
         \SB4_20/i0_3 , \SB4_20/i0_4 , \SB4_20/i0[10] , \SB4_20/i0[9] ,
         \SB4_20/i0[8] , \SB4_20/i0[7] , \SB4_20/i0[6] , \SB4_21/i3[0] ,
         \SB4_21/i1_5 , \SB4_21/i1_7 , \SB4_21/i0_3 , \SB4_21/i0_4 ,
         \SB4_21/i0[10] , \SB4_21/i0[9] , \SB4_21/i0[8] , \SB4_21/i0[7] ,
         \SB4_21/i0[6] , \SB4_22/i3[0] , \SB4_22/i1_5 , \SB4_22/i1_7 ,
         \SB4_22/i1[9] , \SB4_22/i0_0 , \SB4_22/i0_3 , \SB4_22/i0_4 ,
         \SB4_22/i0[10] , \SB4_22/i0[9] , \SB4_22/i0[8] , \SB4_22/i0[7] ,
         \SB4_22/i0[6] , \SB4_23/i3[0] , \SB4_23/i1_5 , \SB4_23/i1_7 ,
         \SB4_23/i1[9] , \SB4_23/i0_0 , \SB4_23/i0_3 , \SB4_23/i0_4 ,
         \SB4_23/i0[10] , \SB4_23/i0[9] , \SB4_23/i0[8] , \SB4_23/i0[7] ,
         \SB4_23/i0[6] , \SB4_24/i3[0] , \SB4_24/i1_5 , \SB4_24/i1_7 ,
         \SB4_24/i1[9] , \SB4_24/i0_0 , \SB4_24/i0_3 , \SB4_24/i0_4 ,
         \SB4_24/i0[10] , \SB4_24/i0[9] , \SB4_24/i0[8] , \SB4_24/i0[7] ,
         \SB4_24/i0[6] , \SB4_25/i3[0] , \SB4_25/i1_5 , \SB4_25/i1_7 ,
         \SB4_25/i1[9] , \SB4_25/i0_0 , \SB4_25/i0_3 , \SB4_25/i0_4 ,
         \SB4_25/i0[10] , \SB4_25/i0[9] , \SB4_25/i0[8] , \SB4_25/i0[7] ,
         \SB4_25/i0[6] , \SB4_26/i3[0] , \SB4_26/i1_5 , \SB4_26/i1_7 ,
         \SB4_26/i1[9] , \SB4_26/i0_0 , \SB4_26/i0_3 , \SB4_26/i0_4 ,
         \SB4_26/i0[10] , \SB4_26/i0[9] , \SB4_26/i0[8] , \SB4_26/i0[7] ,
         \SB4_26/i0[6] , \SB4_27/i3[0] , \SB4_27/i1_5 , \SB4_27/i1_7 ,
         \SB4_27/i0_3 , \SB4_27/i0_4 , \SB4_27/i0[10] , \SB4_27/i0[9] ,
         \SB4_27/i0[8] , \SB4_27/i0[7] , \SB4_27/i0[6] , \SB4_28/i3[0] ,
         \SB4_28/i1_5 , \SB4_28/i1_7 , \SB4_28/i0_0 , \SB4_28/i0_3 ,
         \SB4_28/i0_4 , \SB4_28/i0[10] , \SB4_28/i0[9] , \SB4_28/i0[8] ,
         \SB4_28/i0[7] , \SB4_28/i0[6] , \SB4_29/i3[0] , \SB4_29/i1_5 ,
         \SB4_29/i1_7 , \SB4_29/i1[9] , \SB4_29/i0_0 , \SB4_29/i0_3 ,
         \SB4_29/i0_4 , \SB4_29/i0[10] , \SB4_29/i0[9] , \SB4_29/i0[8] ,
         \SB4_29/i0[7] , \SB4_29/i0[6] , \SB4_30/i3[0] , \SB4_30/i1_7 ,
         \SB4_30/i0_0 , \SB4_30/i0_3 , \SB4_30/i0_4 , \SB4_30/i0[10] ,
         \SB4_30/i0[9] , \SB4_30/i0[8] , \SB4_30/i0[7] , \SB4_30/i0[6] ,
         \SB4_31/i3[0] , \SB4_31/i1_5 , \SB4_31/i1_7 , \SB4_31/i1[9] ,
         \SB4_31/i0_0 , \SB4_31/i0_3 , \SB4_31/i0_4 , \SB4_31/i0[10] ,
         \SB4_31/i0[9] , \SB4_31/i0[7] , \SB4_31/i0[6] ,
         \SB1_0_0/Component_Function_2/NAND4_in[2] ,
         \SB1_0_0/Component_Function_2/NAND4_in[1] ,
         \SB1_0_0/Component_Function_2/NAND4_in[0] ,
         \SB1_0_0/Component_Function_3/NAND4_in[3] ,
         \SB1_0_0/Component_Function_3/NAND4_in[2] ,
         \SB1_0_0/Component_Function_3/NAND4_in[1] ,
         \SB1_0_0/Component_Function_4/NAND4_in[3] ,
         \SB1_0_0/Component_Function_4/NAND4_in[1] ,
         \SB1_0_0/Component_Function_4/NAND4_in[0] ,
         \SB1_0_1/Component_Function_2/NAND4_in[3] ,
         \SB1_0_1/Component_Function_2/NAND4_in[2] ,
         \SB1_0_1/Component_Function_2/NAND4_in[1] ,
         \SB1_0_1/Component_Function_2/NAND4_in[0] ,
         \SB1_0_1/Component_Function_3/NAND4_in[2] ,
         \SB1_0_1/Component_Function_3/NAND4_in[1] ,
         \SB1_0_1/Component_Function_3/NAND4_in[0] ,
         \SB1_0_1/Component_Function_4/NAND4_in[3] ,
         \SB1_0_1/Component_Function_4/NAND4_in[2] ,
         \SB1_0_1/Component_Function_4/NAND4_in[1] ,
         \SB1_0_1/Component_Function_4/NAND4_in[0] ,
         \SB1_0_2/Component_Function_2/NAND4_in[2] ,
         \SB1_0_2/Component_Function_2/NAND4_in[0] ,
         \SB1_0_2/Component_Function_3/NAND4_in[3] ,
         \SB1_0_2/Component_Function_3/NAND4_in[2] ,
         \SB1_0_2/Component_Function_3/NAND4_in[1] ,
         \SB1_0_2/Component_Function_3/NAND4_in[0] ,
         \SB1_0_2/Component_Function_4/NAND4_in[3] ,
         \SB1_0_2/Component_Function_4/NAND4_in[2] ,
         \SB1_0_2/Component_Function_4/NAND4_in[1] ,
         \SB1_0_3/Component_Function_2/NAND4_in[3] ,
         \SB1_0_3/Component_Function_2/NAND4_in[2] ,
         \SB1_0_3/Component_Function_2/NAND4_in[0] ,
         \SB1_0_3/Component_Function_3/NAND4_in[3] ,
         \SB1_0_3/Component_Function_3/NAND4_in[1] ,
         \SB1_0_3/Component_Function_4/NAND4_in[3] ,
         \SB1_0_3/Component_Function_4/NAND4_in[2] ,
         \SB1_0_3/Component_Function_4/NAND4_in[1] ,
         \SB1_0_4/Component_Function_2/NAND4_in[3] ,
         \SB1_0_4/Component_Function_2/NAND4_in[2] ,
         \SB1_0_4/Component_Function_2/NAND4_in[1] ,
         \SB1_0_4/Component_Function_2/NAND4_in[0] ,
         \SB1_0_4/Component_Function_3/NAND4_in[3] ,
         \SB1_0_4/Component_Function_3/NAND4_in[1] ,
         \SB1_0_4/Component_Function_4/NAND4_in[3] ,
         \SB1_0_4/Component_Function_4/NAND4_in[2] ,
         \SB1_0_4/Component_Function_4/NAND4_in[1] ,
         \SB1_0_4/Component_Function_4/NAND4_in[0] ,
         \SB1_0_5/Component_Function_2/NAND4_in[2] ,
         \SB1_0_5/Component_Function_2/NAND4_in[0] ,
         \SB1_0_5/Component_Function_3/NAND4_in[3] ,
         \SB1_0_5/Component_Function_3/NAND4_in[1] ,
         \SB1_0_5/Component_Function_3/NAND4_in[0] ,
         \SB1_0_5/Component_Function_4/NAND4_in[3] ,
         \SB1_0_5/Component_Function_4/NAND4_in[1] ,
         \SB1_0_5/Component_Function_4/NAND4_in[0] ,
         \SB1_0_6/Component_Function_2/NAND4_in[2] ,
         \SB1_0_6/Component_Function_2/NAND4_in[1] ,
         \SB1_0_6/Component_Function_2/NAND4_in[0] ,
         \SB1_0_6/Component_Function_3/NAND4_in[2] ,
         \SB1_0_6/Component_Function_3/NAND4_in[0] ,
         \SB1_0_6/Component_Function_4/NAND4_in[3] ,
         \SB1_0_6/Component_Function_4/NAND4_in[0] ,
         \SB1_0_7/Component_Function_2/NAND4_in[3] ,
         \SB1_0_7/Component_Function_2/NAND4_in[2] ,
         \SB1_0_7/Component_Function_2/NAND4_in[1] ,
         \SB1_0_7/Component_Function_2/NAND4_in[0] ,
         \SB1_0_7/Component_Function_3/NAND4_in[3] ,
         \SB1_0_7/Component_Function_3/NAND4_in[2] ,
         \SB1_0_7/Component_Function_3/NAND4_in[1] ,
         \SB1_0_7/Component_Function_3/NAND4_in[0] ,
         \SB1_0_7/Component_Function_4/NAND4_in[1] ,
         \SB1_0_7/Component_Function_4/NAND4_in[0] ,
         \SB1_0_8/Component_Function_2/NAND4_in[2] ,
         \SB1_0_8/Component_Function_2/NAND4_in[1] ,
         \SB1_0_8/Component_Function_2/NAND4_in[0] ,
         \SB1_0_8/Component_Function_3/NAND4_in[2] ,
         \SB1_0_8/Component_Function_3/NAND4_in[0] ,
         \SB1_0_8/Component_Function_4/NAND4_in[3] ,
         \SB1_0_8/Component_Function_4/NAND4_in[2] ,
         \SB1_0_8/Component_Function_4/NAND4_in[1] ,
         \SB1_0_8/Component_Function_4/NAND4_in[0] ,
         \SB1_0_9/Component_Function_2/NAND4_in[3] ,
         \SB1_0_9/Component_Function_2/NAND4_in[2] ,
         \SB1_0_9/Component_Function_2/NAND4_in[0] ,
         \SB1_0_9/Component_Function_3/NAND4_in[3] ,
         \SB1_0_9/Component_Function_3/NAND4_in[1] ,
         \SB1_0_9/Component_Function_3/NAND4_in[0] ,
         \SB1_0_9/Component_Function_4/NAND4_in[3] ,
         \SB1_0_9/Component_Function_4/NAND4_in[2] ,
         \SB1_0_9/Component_Function_4/NAND4_in[1] ,
         \SB1_0_9/Component_Function_4/NAND4_in[0] ,
         \SB1_0_10/Component_Function_2/NAND4_in[2] ,
         \SB1_0_10/Component_Function_2/NAND4_in[0] ,
         \SB1_0_10/Component_Function_3/NAND4_in[3] ,
         \SB1_0_10/Component_Function_3/NAND4_in[2] ,
         \SB1_0_10/Component_Function_3/NAND4_in[1] ,
         \SB1_0_10/Component_Function_3/NAND4_in[0] ,
         \SB1_0_10/Component_Function_4/NAND4_in[3] ,
         \SB1_0_10/Component_Function_4/NAND4_in[2] ,
         \SB1_0_10/Component_Function_4/NAND4_in[0] ,
         \SB1_0_11/Component_Function_2/NAND4_in[2] ,
         \SB1_0_11/Component_Function_2/NAND4_in[1] ,
         \SB1_0_11/Component_Function_3/NAND4_in[3] ,
         \SB1_0_11/Component_Function_3/NAND4_in[1] ,
         \SB1_0_11/Component_Function_3/NAND4_in[0] ,
         \SB1_0_11/Component_Function_4/NAND4_in[3] ,
         \SB1_0_11/Component_Function_4/NAND4_in[1] ,
         \SB1_0_11/Component_Function_4/NAND4_in[0] ,
         \SB1_0_12/Component_Function_2/NAND4_in[2] ,
         \SB1_0_12/Component_Function_2/NAND4_in[0] ,
         \SB1_0_12/Component_Function_3/NAND4_in[3] ,
         \SB1_0_12/Component_Function_3/NAND4_in[1] ,
         \SB1_0_12/Component_Function_4/NAND4_in[3] ,
         \SB1_0_12/Component_Function_4/NAND4_in[1] ,
         \SB1_0_12/Component_Function_4/NAND4_in[0] ,
         \SB1_0_13/Component_Function_2/NAND4_in[2] ,
         \SB1_0_13/Component_Function_2/NAND4_in[1] ,
         \SB1_0_13/Component_Function_2/NAND4_in[0] ,
         \SB1_0_13/Component_Function_3/NAND4_in[3] ,
         \SB1_0_13/Component_Function_3/NAND4_in[2] ,
         \SB1_0_13/Component_Function_3/NAND4_in[0] ,
         \SB1_0_13/Component_Function_4/NAND4_in[3] ,
         \SB1_0_13/Component_Function_4/NAND4_in[1] ,
         \SB1_0_13/Component_Function_4/NAND4_in[0] ,
         \SB1_0_14/Component_Function_2/NAND4_in[3] ,
         \SB1_0_14/Component_Function_2/NAND4_in[1] ,
         \SB1_0_14/Component_Function_2/NAND4_in[0] ,
         \SB1_0_14/Component_Function_3/NAND4_in[3] ,
         \SB1_0_14/Component_Function_3/NAND4_in[2] ,
         \SB1_0_14/Component_Function_3/NAND4_in[1] ,
         \SB1_0_14/Component_Function_3/NAND4_in[0] ,
         \SB1_0_14/Component_Function_4/NAND4_in[3] ,
         \SB1_0_14/Component_Function_4/NAND4_in[2] ,
         \SB1_0_14/Component_Function_4/NAND4_in[1] ,
         \SB1_0_15/Component_Function_2/NAND4_in[3] ,
         \SB1_0_15/Component_Function_2/NAND4_in[1] ,
         \SB1_0_15/Component_Function_2/NAND4_in[0] ,
         \SB1_0_15/Component_Function_3/NAND4_in[3] ,
         \SB1_0_15/Component_Function_3/NAND4_in[1] ,
         \SB1_0_15/Component_Function_3/NAND4_in[0] ,
         \SB1_0_15/Component_Function_4/NAND4_in[3] ,
         \SB1_0_15/Component_Function_4/NAND4_in[1] ,
         \SB1_0_15/Component_Function_4/NAND4_in[0] ,
         \SB1_0_16/Component_Function_2/NAND4_in[1] ,
         \SB1_0_16/Component_Function_2/NAND4_in[0] ,
         \SB1_0_16/Component_Function_3/NAND4_in[2] ,
         \SB1_0_16/Component_Function_3/NAND4_in[1] ,
         \SB1_0_16/Component_Function_3/NAND4_in[0] ,
         \SB1_0_16/Component_Function_4/NAND4_in[3] ,
         \SB1_0_16/Component_Function_4/NAND4_in[2] ,
         \SB1_0_16/Component_Function_4/NAND4_in[1] ,
         \SB1_0_17/Component_Function_2/NAND4_in[2] ,
         \SB1_0_17/Component_Function_2/NAND4_in[1] ,
         \SB1_0_17/Component_Function_2/NAND4_in[0] ,
         \SB1_0_17/Component_Function_3/NAND4_in[3] ,
         \SB1_0_17/Component_Function_3/NAND4_in[2] ,
         \SB1_0_17/Component_Function_3/NAND4_in[0] ,
         \SB1_0_17/Component_Function_4/NAND4_in[3] ,
         \SB1_0_17/Component_Function_4/NAND4_in[1] ,
         \SB1_0_18/Component_Function_2/NAND4_in[3] ,
         \SB1_0_18/Component_Function_2/NAND4_in[2] ,
         \SB1_0_18/Component_Function_2/NAND4_in[0] ,
         \SB1_0_18/Component_Function_3/NAND4_in[3] ,
         \SB1_0_18/Component_Function_3/NAND4_in[2] ,
         \SB1_0_18/Component_Function_3/NAND4_in[1] ,
         \SB1_0_18/Component_Function_3/NAND4_in[0] ,
         \SB1_0_18/Component_Function_4/NAND4_in[3] ,
         \SB1_0_18/Component_Function_4/NAND4_in[1] ,
         \SB1_0_18/Component_Function_4/NAND4_in[0] ,
         \SB1_0_19/Component_Function_2/NAND4_in[3] ,
         \SB1_0_19/Component_Function_2/NAND4_in[2] ,
         \SB1_0_19/Component_Function_2/NAND4_in[0] ,
         \SB1_0_19/Component_Function_3/NAND4_in[3] ,
         \SB1_0_19/Component_Function_3/NAND4_in[2] ,
         \SB1_0_19/Component_Function_3/NAND4_in[1] ,
         \SB1_0_19/Component_Function_3/NAND4_in[0] ,
         \SB1_0_19/Component_Function_4/NAND4_in[3] ,
         \SB1_0_19/Component_Function_4/NAND4_in[2] ,
         \SB1_0_19/Component_Function_4/NAND4_in[1] ,
         \SB1_0_19/Component_Function_4/NAND4_in[0] ,
         \SB1_0_20/Component_Function_2/NAND4_in[3] ,
         \SB1_0_20/Component_Function_2/NAND4_in[2] ,
         \SB1_0_20/Component_Function_2/NAND4_in[0] ,
         \SB1_0_20/Component_Function_3/NAND4_in[2] ,
         \SB1_0_20/Component_Function_3/NAND4_in[1] ,
         \SB1_0_20/Component_Function_3/NAND4_in[0] ,
         \SB1_0_20/Component_Function_4/NAND4_in[2] ,
         \SB1_0_20/Component_Function_4/NAND4_in[1] ,
         \SB1_0_21/Component_Function_2/NAND4_in[2] ,
         \SB1_0_21/Component_Function_2/NAND4_in[0] ,
         \SB1_0_21/Component_Function_3/NAND4_in[3] ,
         \SB1_0_21/Component_Function_4/NAND4_in[3] ,
         \SB1_0_21/Component_Function_4/NAND4_in[2] ,
         \SB1_0_21/Component_Function_4/NAND4_in[1] ,
         \SB1_0_22/Component_Function_2/NAND4_in[3] ,
         \SB1_0_22/Component_Function_2/NAND4_in[2] ,
         \SB1_0_22/Component_Function_3/NAND4_in[3] ,
         \SB1_0_22/Component_Function_3/NAND4_in[1] ,
         \SB1_0_22/Component_Function_3/NAND4_in[0] ,
         \SB1_0_22/Component_Function_4/NAND4_in[3] ,
         \SB1_0_22/Component_Function_4/NAND4_in[1] ,
         \SB1_0_22/Component_Function_4/NAND4_in[0] ,
         \SB1_0_23/Component_Function_2/NAND4_in[3] ,
         \SB1_0_23/Component_Function_2/NAND4_in[0] ,
         \SB1_0_23/Component_Function_3/NAND4_in[3] ,
         \SB1_0_23/Component_Function_3/NAND4_in[1] ,
         \SB1_0_23/Component_Function_3/NAND4_in[0] ,
         \SB1_0_23/Component_Function_4/NAND4_in[3] ,
         \SB1_0_23/Component_Function_4/NAND4_in[2] ,
         \SB1_0_23/Component_Function_4/NAND4_in[1] ,
         \SB1_0_23/Component_Function_4/NAND4_in[0] ,
         \SB1_0_24/Component_Function_2/NAND4_in[2] ,
         \SB1_0_24/Component_Function_2/NAND4_in[1] ,
         \SB1_0_24/Component_Function_2/NAND4_in[0] ,
         \SB1_0_24/Component_Function_3/NAND4_in[3] ,
         \SB1_0_24/Component_Function_3/NAND4_in[2] ,
         \SB1_0_24/Component_Function_3/NAND4_in[1] ,
         \SB1_0_24/Component_Function_3/NAND4_in[0] ,
         \SB1_0_24/Component_Function_4/NAND4_in[3] ,
         \SB1_0_24/Component_Function_4/NAND4_in[2] ,
         \SB1_0_24/Component_Function_4/NAND4_in[0] ,
         \SB1_0_25/Component_Function_2/NAND4_in[2] ,
         \SB1_0_25/Component_Function_2/NAND4_in[1] ,
         \SB1_0_25/Component_Function_2/NAND4_in[0] ,
         \SB1_0_25/Component_Function_3/NAND4_in[2] ,
         \SB1_0_25/Component_Function_3/NAND4_in[1] ,
         \SB1_0_25/Component_Function_3/NAND4_in[0] ,
         \SB1_0_25/Component_Function_4/NAND4_in[2] ,
         \SB1_0_25/Component_Function_4/NAND4_in[1] ,
         \SB1_0_25/Component_Function_4/NAND4_in[0] ,
         \SB1_0_26/Component_Function_2/NAND4_in[3] ,
         \SB1_0_26/Component_Function_2/NAND4_in[2] ,
         \SB1_0_26/Component_Function_2/NAND4_in[1] ,
         \SB1_0_26/Component_Function_3/NAND4_in[3] ,
         \SB1_0_26/Component_Function_3/NAND4_in[2] ,
         \SB1_0_26/Component_Function_3/NAND4_in[1] ,
         \SB1_0_26/Component_Function_3/NAND4_in[0] ,
         \SB1_0_26/Component_Function_4/NAND4_in[3] ,
         \SB1_0_26/Component_Function_4/NAND4_in[2] ,
         \SB1_0_26/Component_Function_4/NAND4_in[1] ,
         \SB1_0_26/Component_Function_4/NAND4_in[0] ,
         \SB1_0_27/Component_Function_2/NAND4_in[3] ,
         \SB1_0_27/Component_Function_2/NAND4_in[2] ,
         \SB1_0_27/Component_Function_2/NAND4_in[1] ,
         \SB1_0_27/Component_Function_2/NAND4_in[0] ,
         \SB1_0_27/Component_Function_3/NAND4_in[3] ,
         \SB1_0_27/Component_Function_3/NAND4_in[1] ,
         \SB1_0_27/Component_Function_4/NAND4_in[3] ,
         \SB1_0_27/Component_Function_4/NAND4_in[2] ,
         \SB1_0_27/Component_Function_4/NAND4_in[1] ,
         \SB1_0_27/Component_Function_4/NAND4_in[0] ,
         \SB1_0_28/Component_Function_2/NAND4_in[2] ,
         \SB1_0_28/Component_Function_2/NAND4_in[1] ,
         \SB1_0_28/Component_Function_2/NAND4_in[0] ,
         \SB1_0_28/Component_Function_3/NAND4_in[3] ,
         \SB1_0_28/Component_Function_3/NAND4_in[2] ,
         \SB1_0_28/Component_Function_3/NAND4_in[1] ,
         \SB1_0_28/Component_Function_4/NAND4_in[3] ,
         \SB1_0_28/Component_Function_4/NAND4_in[1] ,
         \SB1_0_28/Component_Function_4/NAND4_in[0] ,
         \SB1_0_29/Component_Function_3/NAND4_in[3] ,
         \SB1_0_29/Component_Function_3/NAND4_in[1] ,
         \SB1_0_29/Component_Function_4/NAND4_in[3] ,
         \SB1_0_29/Component_Function_4/NAND4_in[1] ,
         \SB1_0_30/Component_Function_2/NAND4_in[3] ,
         \SB1_0_30/Component_Function_2/NAND4_in[2] ,
         \SB1_0_30/Component_Function_2/NAND4_in[1] ,
         \SB1_0_30/Component_Function_2/NAND4_in[0] ,
         \SB1_0_30/Component_Function_3/NAND4_in[3] ,
         \SB1_0_30/Component_Function_3/NAND4_in[1] ,
         \SB1_0_30/Component_Function_3/NAND4_in[0] ,
         \SB1_0_30/Component_Function_4/NAND4_in[3] ,
         \SB1_0_30/Component_Function_4/NAND4_in[2] ,
         \SB1_0_30/Component_Function_4/NAND4_in[1] ,
         \SB1_0_30/Component_Function_4/NAND4_in[0] ,
         \SB1_0_31/Component_Function_2/NAND4_in[3] ,
         \SB1_0_31/Component_Function_2/NAND4_in[2] ,
         \SB1_0_31/Component_Function_2/NAND4_in[1] ,
         \SB1_0_31/Component_Function_2/NAND4_in[0] ,
         \SB1_0_31/Component_Function_3/NAND4_in[3] ,
         \SB1_0_31/Component_Function_3/NAND4_in[1] ,
         \SB1_0_31/Component_Function_3/NAND4_in[0] ,
         \SB1_0_31/Component_Function_4/NAND4_in[3] ,
         \SB1_0_31/Component_Function_4/NAND4_in[2] ,
         \SB1_0_31/Component_Function_4/NAND4_in[1] ,
         \SB1_0_31/Component_Function_4/NAND4_in[0] ,
         \SB2_0_0/Component_Function_2/NAND4_in[3] ,
         \SB2_0_0/Component_Function_2/NAND4_in[2] ,
         \SB2_0_0/Component_Function_2/NAND4_in[1] ,
         \SB2_0_0/Component_Function_2/NAND4_in[0] ,
         \SB2_0_0/Component_Function_3/NAND4_in[3] ,
         \SB2_0_0/Component_Function_4/NAND4_in[3] ,
         \SB2_0_0/Component_Function_4/NAND4_in[0] ,
         \SB2_0_1/Component_Function_2/NAND4_in[0] ,
         \SB2_0_1/Component_Function_3/NAND4_in[2] ,
         \SB2_0_1/Component_Function_3/NAND4_in[1] ,
         \SB2_0_1/Component_Function_3/NAND4_in[0] ,
         \SB2_0_1/Component_Function_4/NAND4_in[3] ,
         \SB2_0_1/Component_Function_4/NAND4_in[2] ,
         \SB2_0_1/Component_Function_4/NAND4_in[1] ,
         \SB2_0_1/Component_Function_4/NAND4_in[0] ,
         \SB2_0_2/Component_Function_2/NAND4_in[3] ,
         \SB2_0_2/Component_Function_2/NAND4_in[1] ,
         \SB2_0_2/Component_Function_2/NAND4_in[0] ,
         \SB2_0_2/Component_Function_3/NAND4_in[3] ,
         \SB2_0_2/Component_Function_4/NAND4_in[3] ,
         \SB2_0_2/Component_Function_4/NAND4_in[1] ,
         \SB2_0_2/Component_Function_4/NAND4_in[0] ,
         \SB2_0_3/Component_Function_2/NAND4_in[2] ,
         \SB2_0_3/Component_Function_2/NAND4_in[1] ,
         \SB2_0_3/Component_Function_2/NAND4_in[0] ,
         \SB2_0_3/Component_Function_3/NAND4_in[3] ,
         \SB2_0_3/Component_Function_3/NAND4_in[2] ,
         \SB2_0_3/Component_Function_3/NAND4_in[1] ,
         \SB2_0_3/Component_Function_3/NAND4_in[0] ,
         \SB2_0_3/Component_Function_4/NAND4_in[3] ,
         \SB2_0_3/Component_Function_4/NAND4_in[2] ,
         \SB2_0_3/Component_Function_4/NAND4_in[1] ,
         \SB2_0_3/Component_Function_4/NAND4_in[0] ,
         \SB2_0_4/Component_Function_2/NAND4_in[3] ,
         \SB2_0_4/Component_Function_2/NAND4_in[2] ,
         \SB2_0_4/Component_Function_2/NAND4_in[1] ,
         \SB2_0_4/Component_Function_2/NAND4_in[0] ,
         \SB2_0_4/Component_Function_3/NAND4_in[3] ,
         \SB2_0_4/Component_Function_3/NAND4_in[2] ,
         \SB2_0_4/Component_Function_4/NAND4_in[3] ,
         \SB2_0_4/Component_Function_4/NAND4_in[1] ,
         \SB2_0_4/Component_Function_4/NAND4_in[0] ,
         \SB2_0_5/Component_Function_2/NAND4_in[3] ,
         \SB2_0_5/Component_Function_2/NAND4_in[2] ,
         \SB2_0_5/Component_Function_2/NAND4_in[0] ,
         \SB2_0_5/Component_Function_3/NAND4_in[3] ,
         \SB2_0_5/Component_Function_3/NAND4_in[1] ,
         \SB2_0_5/Component_Function_4/NAND4_in[2] ,
         \SB2_0_5/Component_Function_4/NAND4_in[1] ,
         \SB2_0_5/Component_Function_4/NAND4_in[0] ,
         \SB2_0_6/Component_Function_2/NAND4_in[2] ,
         \SB2_0_6/Component_Function_2/NAND4_in[1] ,
         \SB2_0_6/Component_Function_2/NAND4_in[0] ,
         \SB2_0_6/Component_Function_3/NAND4_in[3] ,
         \SB2_0_6/Component_Function_3/NAND4_in[2] ,
         \SB2_0_6/Component_Function_3/NAND4_in[1] ,
         \SB2_0_6/Component_Function_3/NAND4_in[0] ,
         \SB2_0_6/Component_Function_4/NAND4_in[3] ,
         \SB2_0_6/Component_Function_4/NAND4_in[1] ,
         \SB2_0_6/Component_Function_4/NAND4_in[0] ,
         \SB2_0_7/Component_Function_2/NAND4_in[1] ,
         \SB2_0_7/Component_Function_2/NAND4_in[0] ,
         \SB2_0_7/Component_Function_3/NAND4_in[3] ,
         \SB2_0_7/Component_Function_3/NAND4_in[2] ,
         \SB2_0_7/Component_Function_3/NAND4_in[1] ,
         \SB2_0_7/Component_Function_3/NAND4_in[0] ,
         \SB2_0_7/Component_Function_4/NAND4_in[3] ,
         \SB2_0_7/Component_Function_4/NAND4_in[1] ,
         \SB2_0_7/Component_Function_4/NAND4_in[0] ,
         \SB2_0_8/Component_Function_2/NAND4_in[3] ,
         \SB2_0_8/Component_Function_2/NAND4_in[2] ,
         \SB2_0_8/Component_Function_2/NAND4_in[1] ,
         \SB2_0_8/Component_Function_2/NAND4_in[0] ,
         \SB2_0_8/Component_Function_3/NAND4_in[3] ,
         \SB2_0_8/Component_Function_3/NAND4_in[2] ,
         \SB2_0_8/Component_Function_3/NAND4_in[0] ,
         \SB2_0_8/Component_Function_4/NAND4_in[3] ,
         \SB2_0_8/Component_Function_4/NAND4_in[2] ,
         \SB2_0_8/Component_Function_4/NAND4_in[1] ,
         \SB2_0_8/Component_Function_4/NAND4_in[0] ,
         \SB2_0_9/Component_Function_2/NAND4_in[3] ,
         \SB2_0_9/Component_Function_2/NAND4_in[0] ,
         \SB2_0_9/Component_Function_3/NAND4_in[3] ,
         \SB2_0_9/Component_Function_3/NAND4_in[1] ,
         \SB2_0_9/Component_Function_3/NAND4_in[0] ,
         \SB2_0_9/Component_Function_4/NAND4_in[3] ,
         \SB2_0_9/Component_Function_4/NAND4_in[1] ,
         \SB2_0_9/Component_Function_4/NAND4_in[0] ,
         \SB2_0_10/Component_Function_2/NAND4_in[3] ,
         \SB2_0_10/Component_Function_2/NAND4_in[0] ,
         \SB2_0_10/Component_Function_3/NAND4_in[3] ,
         \SB2_0_10/Component_Function_3/NAND4_in[1] ,
         \SB2_0_10/Component_Function_3/NAND4_in[0] ,
         \SB2_0_10/Component_Function_4/NAND4_in[3] ,
         \SB2_0_10/Component_Function_4/NAND4_in[1] ,
         \SB2_0_10/Component_Function_4/NAND4_in[0] ,
         \SB2_0_11/Component_Function_2/NAND4_in[3] ,
         \SB2_0_11/Component_Function_2/NAND4_in[2] ,
         \SB2_0_11/Component_Function_2/NAND4_in[1] ,
         \SB2_0_11/Component_Function_2/NAND4_in[0] ,
         \SB2_0_11/Component_Function_3/NAND4_in[2] ,
         \SB2_0_11/Component_Function_3/NAND4_in[0] ,
         \SB2_0_11/Component_Function_4/NAND4_in[3] ,
         \SB2_0_11/Component_Function_4/NAND4_in[2] ,
         \SB2_0_11/Component_Function_4/NAND4_in[1] ,
         \SB2_0_11/Component_Function_4/NAND4_in[0] ,
         \SB2_0_12/Component_Function_2/NAND4_in[2] ,
         \SB2_0_12/Component_Function_2/NAND4_in[1] ,
         \SB2_0_12/Component_Function_2/NAND4_in[0] ,
         \SB2_0_12/Component_Function_3/NAND4_in[2] ,
         \SB2_0_12/Component_Function_3/NAND4_in[1] ,
         \SB2_0_12/Component_Function_3/NAND4_in[0] ,
         \SB2_0_12/Component_Function_4/NAND4_in[3] ,
         \SB2_0_12/Component_Function_4/NAND4_in[2] ,
         \SB2_0_12/Component_Function_4/NAND4_in[1] ,
         \SB2_0_12/Component_Function_4/NAND4_in[0] ,
         \SB2_0_13/Component_Function_2/NAND4_in[2] ,
         \SB2_0_13/Component_Function_2/NAND4_in[1] ,
         \SB2_0_13/Component_Function_2/NAND4_in[0] ,
         \SB2_0_13/Component_Function_3/NAND4_in[3] ,
         \SB2_0_13/Component_Function_3/NAND4_in[2] ,
         \SB2_0_13/Component_Function_3/NAND4_in[1] ,
         \SB2_0_13/Component_Function_3/NAND4_in[0] ,
         \SB2_0_13/Component_Function_4/NAND4_in[3] ,
         \SB2_0_13/Component_Function_4/NAND4_in[2] ,
         \SB2_0_13/Component_Function_4/NAND4_in[1] ,
         \SB2_0_13/Component_Function_4/NAND4_in[0] ,
         \SB2_0_14/Component_Function_2/NAND4_in[3] ,
         \SB2_0_14/Component_Function_2/NAND4_in[2] ,
         \SB2_0_14/Component_Function_2/NAND4_in[1] ,
         \SB2_0_14/Component_Function_2/NAND4_in[0] ,
         \SB2_0_14/Component_Function_3/NAND4_in[3] ,
         \SB2_0_14/Component_Function_3/NAND4_in[2] ,
         \SB2_0_14/Component_Function_3/NAND4_in[1] ,
         \SB2_0_14/Component_Function_3/NAND4_in[0] ,
         \SB2_0_14/Component_Function_4/NAND4_in[3] ,
         \SB2_0_14/Component_Function_4/NAND4_in[1] ,
         \SB2_0_14/Component_Function_4/NAND4_in[0] ,
         \SB2_0_15/Component_Function_2/NAND4_in[2] ,
         \SB2_0_15/Component_Function_2/NAND4_in[1] ,
         \SB2_0_15/Component_Function_2/NAND4_in[0] ,
         \SB2_0_15/Component_Function_3/NAND4_in[3] ,
         \SB2_0_15/Component_Function_3/NAND4_in[1] ,
         \SB2_0_15/Component_Function_3/NAND4_in[0] ,
         \SB2_0_15/Component_Function_4/NAND4_in[3] ,
         \SB2_0_15/Component_Function_4/NAND4_in[1] ,
         \SB2_0_15/Component_Function_4/NAND4_in[0] ,
         \SB2_0_16/Component_Function_2/NAND4_in[3] ,
         \SB2_0_16/Component_Function_2/NAND4_in[1] ,
         \SB2_0_16/Component_Function_2/NAND4_in[0] ,
         \SB2_0_16/Component_Function_3/NAND4_in[3] ,
         \SB2_0_16/Component_Function_3/NAND4_in[1] ,
         \SB2_0_16/Component_Function_3/NAND4_in[0] ,
         \SB2_0_16/Component_Function_4/NAND4_in[3] ,
         \SB2_0_16/Component_Function_4/NAND4_in[1] ,
         \SB2_0_16/Component_Function_4/NAND4_in[0] ,
         \SB2_0_17/Component_Function_2/NAND4_in[2] ,
         \SB2_0_17/Component_Function_2/NAND4_in[1] ,
         \SB2_0_17/Component_Function_2/NAND4_in[0] ,
         \SB2_0_17/Component_Function_3/NAND4_in[3] ,
         \SB2_0_17/Component_Function_3/NAND4_in[2] ,
         \SB2_0_17/Component_Function_3/NAND4_in[1] ,
         \SB2_0_17/Component_Function_4/NAND4_in[3] ,
         \SB2_0_17/Component_Function_4/NAND4_in[1] ,
         \SB2_0_17/Component_Function_4/NAND4_in[0] ,
         \SB2_0_18/Component_Function_2/NAND4_in[0] ,
         \SB2_0_18/Component_Function_3/NAND4_in[3] ,
         \SB2_0_18/Component_Function_3/NAND4_in[2] ,
         \SB2_0_18/Component_Function_3/NAND4_in[1] ,
         \SB2_0_18/Component_Function_4/NAND4_in[3] ,
         \SB2_0_18/Component_Function_4/NAND4_in[2] ,
         \SB2_0_18/Component_Function_4/NAND4_in[1] ,
         \SB2_0_18/Component_Function_4/NAND4_in[0] ,
         \SB2_0_19/Component_Function_2/NAND4_in[3] ,
         \SB2_0_19/Component_Function_2/NAND4_in[1] ,
         \SB2_0_19/Component_Function_2/NAND4_in[0] ,
         \SB2_0_19/Component_Function_3/NAND4_in[2] ,
         \SB2_0_19/Component_Function_3/NAND4_in[0] ,
         \SB2_0_19/Component_Function_4/NAND4_in[3] ,
         \SB2_0_19/Component_Function_4/NAND4_in[2] ,
         \SB2_0_19/Component_Function_4/NAND4_in[1] ,
         \SB2_0_19/Component_Function_4/NAND4_in[0] ,
         \SB2_0_20/Component_Function_2/NAND4_in[2] ,
         \SB2_0_20/Component_Function_2/NAND4_in[1] ,
         \SB2_0_20/Component_Function_2/NAND4_in[0] ,
         \SB2_0_20/Component_Function_3/NAND4_in[3] ,
         \SB2_0_20/Component_Function_3/NAND4_in[1] ,
         \SB2_0_20/Component_Function_3/NAND4_in[0] ,
         \SB2_0_20/Component_Function_4/NAND4_in[1] ,
         \SB2_0_20/Component_Function_4/NAND4_in[0] ,
         \SB2_0_21/Component_Function_2/NAND4_in[3] ,
         \SB2_0_21/Component_Function_2/NAND4_in[1] ,
         \SB2_0_21/Component_Function_2/NAND4_in[0] ,
         \SB2_0_21/Component_Function_3/NAND4_in[3] ,
         \SB2_0_21/Component_Function_4/NAND4_in[3] ,
         \SB2_0_21/Component_Function_4/NAND4_in[2] ,
         \SB2_0_21/Component_Function_4/NAND4_in[1] ,
         \SB2_0_21/Component_Function_4/NAND4_in[0] ,
         \SB2_0_22/Component_Function_2/NAND4_in[2] ,
         \SB2_0_22/Component_Function_2/NAND4_in[1] ,
         \SB2_0_22/Component_Function_2/NAND4_in[0] ,
         \SB2_0_22/Component_Function_3/NAND4_in[2] ,
         \SB2_0_22/Component_Function_3/NAND4_in[0] ,
         \SB2_0_22/Component_Function_4/NAND4_in[3] ,
         \SB2_0_22/Component_Function_4/NAND4_in[2] ,
         \SB2_0_22/Component_Function_4/NAND4_in[1] ,
         \SB2_0_22/Component_Function_4/NAND4_in[0] ,
         \SB2_0_23/Component_Function_2/NAND4_in[3] ,
         \SB2_0_23/Component_Function_2/NAND4_in[1] ,
         \SB2_0_23/Component_Function_2/NAND4_in[0] ,
         \SB2_0_23/Component_Function_3/NAND4_in[2] ,
         \SB2_0_23/Component_Function_3/NAND4_in[0] ,
         \SB2_0_23/Component_Function_4/NAND4_in[3] ,
         \SB2_0_23/Component_Function_4/NAND4_in[1] ,
         \SB2_0_23/Component_Function_4/NAND4_in[0] ,
         \SB2_0_24/Component_Function_2/NAND4_in[3] ,
         \SB2_0_24/Component_Function_2/NAND4_in[2] ,
         \SB2_0_24/Component_Function_3/NAND4_in[3] ,
         \SB2_0_24/Component_Function_3/NAND4_in[0] ,
         \SB2_0_24/Component_Function_4/NAND4_in[3] ,
         \SB2_0_24/Component_Function_4/NAND4_in[2] ,
         \SB2_0_24/Component_Function_4/NAND4_in[1] ,
         \SB2_0_24/Component_Function_4/NAND4_in[0] ,
         \SB2_0_25/Component_Function_2/NAND4_in[2] ,
         \SB2_0_25/Component_Function_2/NAND4_in[0] ,
         \SB2_0_25/Component_Function_3/NAND4_in[2] ,
         \SB2_0_25/Component_Function_3/NAND4_in[0] ,
         \SB2_0_25/Component_Function_4/NAND4_in[3] ,
         \SB2_0_25/Component_Function_4/NAND4_in[2] ,
         \SB2_0_25/Component_Function_4/NAND4_in[0] ,
         \SB2_0_26/Component_Function_2/NAND4_in[3] ,
         \SB2_0_26/Component_Function_2/NAND4_in[2] ,
         \SB2_0_26/Component_Function_2/NAND4_in[1] ,
         \SB2_0_26/Component_Function_2/NAND4_in[0] ,
         \SB2_0_26/Component_Function_3/NAND4_in[3] ,
         \SB2_0_26/Component_Function_3/NAND4_in[2] ,
         \SB2_0_26/Component_Function_3/NAND4_in[1] ,
         \SB2_0_26/Component_Function_3/NAND4_in[0] ,
         \SB2_0_26/Component_Function_4/NAND4_in[3] ,
         \SB2_0_26/Component_Function_4/NAND4_in[1] ,
         \SB2_0_26/Component_Function_4/NAND4_in[0] ,
         \SB2_0_27/Component_Function_2/NAND4_in[3] ,
         \SB2_0_27/Component_Function_2/NAND4_in[2] ,
         \SB2_0_27/Component_Function_2/NAND4_in[1] ,
         \SB2_0_27/Component_Function_2/NAND4_in[0] ,
         \SB2_0_27/Component_Function_3/NAND4_in[3] ,
         \SB2_0_27/Component_Function_3/NAND4_in[2] ,
         \SB2_0_27/Component_Function_3/NAND4_in[1] ,
         \SB2_0_27/Component_Function_3/NAND4_in[0] ,
         \SB2_0_27/Component_Function_4/NAND4_in[3] ,
         \SB2_0_27/Component_Function_4/NAND4_in[1] ,
         \SB2_0_27/Component_Function_4/NAND4_in[0] ,
         \SB2_0_28/Component_Function_2/NAND4_in[2] ,
         \SB2_0_28/Component_Function_2/NAND4_in[1] ,
         \SB2_0_28/Component_Function_2/NAND4_in[0] ,
         \SB2_0_28/Component_Function_3/NAND4_in[3] ,
         \SB2_0_28/Component_Function_3/NAND4_in[2] ,
         \SB2_0_28/Component_Function_3/NAND4_in[1] ,
         \SB2_0_28/Component_Function_3/NAND4_in[0] ,
         \SB2_0_28/Component_Function_4/NAND4_in[3] ,
         \SB2_0_28/Component_Function_4/NAND4_in[2] ,
         \SB2_0_28/Component_Function_4/NAND4_in[1] ,
         \SB2_0_28/Component_Function_4/NAND4_in[0] ,
         \SB2_0_29/Component_Function_2/NAND4_in[3] ,
         \SB2_0_29/Component_Function_2/NAND4_in[0] ,
         \SB2_0_29/Component_Function_3/NAND4_in[2] ,
         \SB2_0_29/Component_Function_3/NAND4_in[1] ,
         \SB2_0_29/Component_Function_3/NAND4_in[0] ,
         \SB2_0_29/Component_Function_4/NAND4_in[3] ,
         \SB2_0_29/Component_Function_4/NAND4_in[2] ,
         \SB2_0_29/Component_Function_4/NAND4_in[1] ,
         \SB2_0_29/Component_Function_4/NAND4_in[0] ,
         \SB2_0_30/Component_Function_2/NAND4_in[3] ,
         \SB2_0_30/Component_Function_2/NAND4_in[1] ,
         \SB2_0_30/Component_Function_3/NAND4_in[3] ,
         \SB2_0_30/Component_Function_3/NAND4_in[2] ,
         \SB2_0_30/Component_Function_3/NAND4_in[1] ,
         \SB2_0_30/Component_Function_3/NAND4_in[0] ,
         \SB2_0_30/Component_Function_4/NAND4_in[3] ,
         \SB2_0_30/Component_Function_4/NAND4_in[2] ,
         \SB2_0_30/Component_Function_4/NAND4_in[1] ,
         \SB2_0_30/Component_Function_4/NAND4_in[0] ,
         \SB2_0_31/Component_Function_2/NAND4_in[2] ,
         \SB2_0_31/Component_Function_2/NAND4_in[1] ,
         \SB2_0_31/Component_Function_2/NAND4_in[0] ,
         \SB2_0_31/Component_Function_3/NAND4_in[3] ,
         \SB2_0_31/Component_Function_3/NAND4_in[2] ,
         \SB2_0_31/Component_Function_3/NAND4_in[0] ,
         \SB2_0_31/Component_Function_4/NAND4_in[2] ,
         \SB2_0_31/Component_Function_4/NAND4_in[1] ,
         \SB2_0_31/Component_Function_4/NAND4_in[0] ,
         \SB1_1_0/Component_Function_2/NAND4_in[3] ,
         \SB1_1_0/Component_Function_2/NAND4_in[0] ,
         \SB1_1_0/Component_Function_3/NAND4_in[1] ,
         \SB1_1_0/Component_Function_3/NAND4_in[0] ,
         \SB1_1_0/Component_Function_4/NAND4_in[3] ,
         \SB1_1_0/Component_Function_4/NAND4_in[1] ,
         \SB1_1_1/Component_Function_2/NAND4_in[2] ,
         \SB1_1_1/Component_Function_2/NAND4_in[0] ,
         \SB1_1_1/Component_Function_3/NAND4_in[3] ,
         \SB1_1_1/Component_Function_3/NAND4_in[2] ,
         \SB1_1_1/Component_Function_3/NAND4_in[1] ,
         \SB1_1_1/Component_Function_3/NAND4_in[0] ,
         \SB1_1_1/Component_Function_4/NAND4_in[3] ,
         \SB1_1_1/Component_Function_4/NAND4_in[2] ,
         \SB1_1_1/Component_Function_4/NAND4_in[1] ,
         \SB1_1_2/Component_Function_2/NAND4_in[3] ,
         \SB1_1_2/Component_Function_2/NAND4_in[1] ,
         \SB1_1_2/Component_Function_2/NAND4_in[0] ,
         \SB1_1_2/Component_Function_3/NAND4_in[2] ,
         \SB1_1_2/Component_Function_3/NAND4_in[1] ,
         \SB1_1_2/Component_Function_4/NAND4_in[3] ,
         \SB1_1_2/Component_Function_4/NAND4_in[2] ,
         \SB1_1_2/Component_Function_4/NAND4_in[1] ,
         \SB1_1_2/Component_Function_4/NAND4_in[0] ,
         \SB1_1_3/Component_Function_2/NAND4_in[2] ,
         \SB1_1_3/Component_Function_2/NAND4_in[0] ,
         \SB1_1_3/Component_Function_3/NAND4_in[3] ,
         \SB1_1_3/Component_Function_3/NAND4_in[2] ,
         \SB1_1_3/Component_Function_3/NAND4_in[1] ,
         \SB1_1_3/Component_Function_3/NAND4_in[0] ,
         \SB1_1_3/Component_Function_4/NAND4_in[1] ,
         \SB1_1_3/Component_Function_4/NAND4_in[0] ,
         \SB1_1_4/Component_Function_2/NAND4_in[3] ,
         \SB1_1_4/Component_Function_2/NAND4_in[2] ,
         \SB1_1_4/Component_Function_2/NAND4_in[0] ,
         \SB1_1_4/Component_Function_3/NAND4_in[3] ,
         \SB1_1_4/Component_Function_3/NAND4_in[1] ,
         \SB1_1_4/Component_Function_3/NAND4_in[0] ,
         \SB1_1_4/Component_Function_4/NAND4_in[2] ,
         \SB1_1_5/Component_Function_2/NAND4_in[3] ,
         \SB1_1_5/Component_Function_2/NAND4_in[2] ,
         \SB1_1_5/Component_Function_2/NAND4_in[1] ,
         \SB1_1_5/Component_Function_2/NAND4_in[0] ,
         \SB1_1_5/Component_Function_3/NAND4_in[2] ,
         \SB1_1_5/Component_Function_3/NAND4_in[1] ,
         \SB1_1_5/Component_Function_4/NAND4_in[3] ,
         \SB1_1_5/Component_Function_4/NAND4_in[2] ,
         \SB1_1_6/Component_Function_2/NAND4_in[1] ,
         \SB1_1_6/Component_Function_2/NAND4_in[0] ,
         \SB1_1_6/Component_Function_3/NAND4_in[1] ,
         \SB1_1_6/Component_Function_4/NAND4_in[3] ,
         \SB1_1_6/Component_Function_4/NAND4_in[2] ,
         \SB1_1_6/Component_Function_4/NAND4_in[1] ,
         \SB1_1_7/Component_Function_2/NAND4_in[3] ,
         \SB1_1_7/Component_Function_2/NAND4_in[2] ,
         \SB1_1_7/Component_Function_2/NAND4_in[1] ,
         \SB1_1_7/Component_Function_2/NAND4_in[0] ,
         \SB1_1_7/Component_Function_3/NAND4_in[2] ,
         \SB1_1_7/Component_Function_3/NAND4_in[1] ,
         \SB1_1_7/Component_Function_3/NAND4_in[0] ,
         \SB1_1_7/Component_Function_4/NAND4_in[3] ,
         \SB1_1_7/Component_Function_4/NAND4_in[1] ,
         \SB1_1_8/Component_Function_2/NAND4_in[3] ,
         \SB1_1_8/Component_Function_2/NAND4_in[2] ,
         \SB1_1_8/Component_Function_3/NAND4_in[3] ,
         \SB1_1_8/Component_Function_3/NAND4_in[2] ,
         \SB1_1_8/Component_Function_3/NAND4_in[1] ,
         \SB1_1_8/Component_Function_3/NAND4_in[0] ,
         \SB1_1_8/Component_Function_4/NAND4_in[1] ,
         \SB1_1_8/Component_Function_4/NAND4_in[0] ,
         \SB1_1_9/Component_Function_2/NAND4_in[2] ,
         \SB1_1_9/Component_Function_2/NAND4_in[1] ,
         \SB1_1_9/Component_Function_3/NAND4_in[2] ,
         \SB1_1_9/Component_Function_3/NAND4_in[1] ,
         \SB1_1_9/Component_Function_3/NAND4_in[0] ,
         \SB1_1_9/Component_Function_4/NAND4_in[3] ,
         \SB1_1_9/Component_Function_4/NAND4_in[2] ,
         \SB1_1_9/Component_Function_4/NAND4_in[1] ,
         \SB1_1_9/Component_Function_4/NAND4_in[0] ,
         \SB1_1_10/Component_Function_2/NAND4_in[3] ,
         \SB1_1_10/Component_Function_2/NAND4_in[1] ,
         \SB1_1_10/Component_Function_2/NAND4_in[0] ,
         \SB1_1_10/Component_Function_3/NAND4_in[2] ,
         \SB1_1_10/Component_Function_3/NAND4_in[1] ,
         \SB1_1_10/Component_Function_3/NAND4_in[0] ,
         \SB1_1_10/Component_Function_4/NAND4_in[1] ,
         \SB1_1_10/Component_Function_4/NAND4_in[0] ,
         \SB1_1_11/Component_Function_2/NAND4_in[2] ,
         \SB1_1_11/Component_Function_2/NAND4_in[0] ,
         \SB1_1_11/Component_Function_3/NAND4_in[1] ,
         \SB1_1_11/Component_Function_4/NAND4_in[3] ,
         \SB1_1_11/Component_Function_4/NAND4_in[2] ,
         \SB1_1_11/Component_Function_4/NAND4_in[0] ,
         \SB1_1_12/Component_Function_2/NAND4_in[1] ,
         \SB1_1_12/Component_Function_2/NAND4_in[0] ,
         \SB1_1_12/Component_Function_3/NAND4_in[2] ,
         \SB1_1_12/Component_Function_3/NAND4_in[1] ,
         \SB1_1_12/Component_Function_4/NAND4_in[2] ,
         \SB1_1_13/Component_Function_2/NAND4_in[1] ,
         \SB1_1_13/Component_Function_2/NAND4_in[0] ,
         \SB1_1_13/Component_Function_3/NAND4_in[2] ,
         \SB1_1_13/Component_Function_3/NAND4_in[1] ,
         \SB1_1_13/Component_Function_3/NAND4_in[0] ,
         \SB1_1_13/Component_Function_4/NAND4_in[0] ,
         \SB1_1_14/Component_Function_2/NAND4_in[3] ,
         \SB1_1_14/Component_Function_2/NAND4_in[2] ,
         \SB1_1_14/Component_Function_3/NAND4_in[3] ,
         \SB1_1_14/Component_Function_3/NAND4_in[1] ,
         \SB1_1_14/Component_Function_4/NAND4_in[3] ,
         \SB1_1_14/Component_Function_4/NAND4_in[2] ,
         \SB1_1_14/Component_Function_4/NAND4_in[1] ,
         \SB1_1_14/Component_Function_4/NAND4_in[0] ,
         \SB1_1_15/Component_Function_2/NAND4_in[3] ,
         \SB1_1_15/Component_Function_2/NAND4_in[2] ,
         \SB1_1_15/Component_Function_2/NAND4_in[1] ,
         \SB1_1_15/Component_Function_2/NAND4_in[0] ,
         \SB1_1_15/Component_Function_3/NAND4_in[2] ,
         \SB1_1_15/Component_Function_3/NAND4_in[1] ,
         \SB1_1_15/Component_Function_3/NAND4_in[0] ,
         \SB1_1_15/Component_Function_4/NAND4_in[3] ,
         \SB1_1_15/Component_Function_4/NAND4_in[2] ,
         \SB1_1_15/Component_Function_4/NAND4_in[1] ,
         \SB1_1_15/Component_Function_4/NAND4_in[0] ,
         \SB1_1_16/Component_Function_2/NAND4_in[1] ,
         \SB1_1_16/Component_Function_3/NAND4_in[2] ,
         \SB1_1_16/Component_Function_3/NAND4_in[1] ,
         \SB1_1_16/Component_Function_3/NAND4_in[0] ,
         \SB1_1_16/Component_Function_4/NAND4_in[3] ,
         \SB1_1_17/Component_Function_2/NAND4_in[2] ,
         \SB1_1_17/Component_Function_2/NAND4_in[0] ,
         \SB1_1_17/Component_Function_3/NAND4_in[3] ,
         \SB1_1_17/Component_Function_3/NAND4_in[2] ,
         \SB1_1_17/Component_Function_3/NAND4_in[1] ,
         \SB1_1_17/Component_Function_3/NAND4_in[0] ,
         \SB1_1_17/Component_Function_4/NAND4_in[2] ,
         \SB1_1_17/Component_Function_4/NAND4_in[1] ,
         \SB1_1_17/Component_Function_4/NAND4_in[0] ,
         \SB1_1_18/Component_Function_2/NAND4_in[2] ,
         \SB1_1_18/Component_Function_2/NAND4_in[1] ,
         \SB1_1_18/Component_Function_2/NAND4_in[0] ,
         \SB1_1_18/Component_Function_3/NAND4_in[2] ,
         \SB1_1_18/Component_Function_3/NAND4_in[1] ,
         \SB1_1_18/Component_Function_3/NAND4_in[0] ,
         \SB1_1_18/Component_Function_4/NAND4_in[2] ,
         \SB1_1_18/Component_Function_4/NAND4_in[1] ,
         \SB1_1_18/Component_Function_4/NAND4_in[0] ,
         \SB1_1_19/Component_Function_2/NAND4_in[3] ,
         \SB1_1_19/Component_Function_2/NAND4_in[1] ,
         \SB1_1_19/Component_Function_2/NAND4_in[0] ,
         \SB1_1_19/Component_Function_3/NAND4_in[3] ,
         \SB1_1_19/Component_Function_3/NAND4_in[1] ,
         \SB1_1_19/Component_Function_3/NAND4_in[0] ,
         \SB1_1_19/Component_Function_4/NAND4_in[1] ,
         \SB1_1_19/Component_Function_4/NAND4_in[0] ,
         \SB1_1_20/Component_Function_2/NAND4_in[3] ,
         \SB1_1_20/Component_Function_2/NAND4_in[2] ,
         \SB1_1_20/Component_Function_2/NAND4_in[1] ,
         \SB1_1_20/Component_Function_2/NAND4_in[0] ,
         \SB1_1_20/Component_Function_3/NAND4_in[3] ,
         \SB1_1_20/Component_Function_3/NAND4_in[2] ,
         \SB1_1_20/Component_Function_3/NAND4_in[1] ,
         \SB1_1_20/Component_Function_3/NAND4_in[0] ,
         \SB1_1_20/Component_Function_4/NAND4_in[3] ,
         \SB1_1_20/Component_Function_4/NAND4_in[1] ,
         \SB1_1_20/Component_Function_4/NAND4_in[0] ,
         \SB1_1_21/Component_Function_2/NAND4_in[3] ,
         \SB1_1_21/Component_Function_2/NAND4_in[1] ,
         \SB1_1_21/Component_Function_3/NAND4_in[0] ,
         \SB1_1_21/Component_Function_4/NAND4_in[3] ,
         \SB1_1_21/Component_Function_4/NAND4_in[1] ,
         \SB1_1_21/Component_Function_4/NAND4_in[0] ,
         \SB1_1_22/Component_Function_2/NAND4_in[3] ,
         \SB1_1_22/Component_Function_2/NAND4_in[2] ,
         \SB1_1_22/Component_Function_2/NAND4_in[1] ,
         \SB1_1_22/Component_Function_3/NAND4_in[3] ,
         \SB1_1_22/Component_Function_3/NAND4_in[1] ,
         \SB1_1_22/Component_Function_3/NAND4_in[0] ,
         \SB1_1_22/Component_Function_4/NAND4_in[3] ,
         \SB1_1_22/Component_Function_4/NAND4_in[1] ,
         \SB1_1_23/Component_Function_2/NAND4_in[1] ,
         \SB1_1_23/Component_Function_3/NAND4_in[2] ,
         \SB1_1_23/Component_Function_3/NAND4_in[1] ,
         \SB1_1_23/Component_Function_3/NAND4_in[0] ,
         \SB1_1_23/Component_Function_4/NAND4_in[2] ,
         \SB1_1_23/Component_Function_4/NAND4_in[1] ,
         \SB1_1_23/Component_Function_4/NAND4_in[0] ,
         \SB1_1_24/Component_Function_2/NAND4_in[3] ,
         \SB1_1_24/Component_Function_2/NAND4_in[2] ,
         \SB1_1_24/Component_Function_2/NAND4_in[1] ,
         \SB1_1_24/Component_Function_2/NAND4_in[0] ,
         \SB1_1_24/Component_Function_3/NAND4_in[1] ,
         \SB1_1_24/Component_Function_3/NAND4_in[0] ,
         \SB1_1_24/Component_Function_4/NAND4_in[3] ,
         \SB1_1_24/Component_Function_4/NAND4_in[2] ,
         \SB1_1_24/Component_Function_4/NAND4_in[1] ,
         \SB1_1_24/Component_Function_4/NAND4_in[0] ,
         \SB1_1_25/Component_Function_2/NAND4_in[2] ,
         \SB1_1_25/Component_Function_2/NAND4_in[1] ,
         \SB1_1_25/Component_Function_2/NAND4_in[0] ,
         \SB1_1_25/Component_Function_3/NAND4_in[1] ,
         \SB1_1_25/Component_Function_3/NAND4_in[0] ,
         \SB1_1_25/Component_Function_4/NAND4_in[3] ,
         \SB1_1_25/Component_Function_4/NAND4_in[2] ,
         \SB1_1_25/Component_Function_4/NAND4_in[1] ,
         \SB1_1_25/Component_Function_4/NAND4_in[0] ,
         \SB1_1_26/Component_Function_2/NAND4_in[2] ,
         \SB1_1_26/Component_Function_3/NAND4_in[1] ,
         \SB1_1_26/Component_Function_3/NAND4_in[0] ,
         \SB1_1_26/Component_Function_4/NAND4_in[3] ,
         \SB1_1_26/Component_Function_4/NAND4_in[1] ,
         \SB1_1_26/Component_Function_4/NAND4_in[0] ,
         \SB1_1_27/Component_Function_2/NAND4_in[1] ,
         \SB1_1_27/Component_Function_2/NAND4_in[0] ,
         \SB1_1_27/Component_Function_3/NAND4_in[2] ,
         \SB1_1_27/Component_Function_3/NAND4_in[1] ,
         \SB1_1_27/Component_Function_3/NAND4_in[0] ,
         \SB1_1_27/Component_Function_4/NAND4_in[3] ,
         \SB1_1_27/Component_Function_4/NAND4_in[2] ,
         \SB1_1_27/Component_Function_4/NAND4_in[1] ,
         \SB1_1_27/Component_Function_4/NAND4_in[0] ,
         \SB1_1_28/Component_Function_2/NAND4_in[2] ,
         \SB1_1_28/Component_Function_2/NAND4_in[1] ,
         \SB1_1_28/Component_Function_3/NAND4_in[2] ,
         \SB1_1_28/Component_Function_3/NAND4_in[0] ,
         \SB1_1_28/Component_Function_4/NAND4_in[3] ,
         \SB1_1_28/Component_Function_4/NAND4_in[2] ,
         \SB1_1_28/Component_Function_4/NAND4_in[1] ,
         \SB1_1_28/Component_Function_4/NAND4_in[0] ,
         \SB1_1_29/Component_Function_2/NAND4_in[1] ,
         \SB1_1_29/Component_Function_2/NAND4_in[0] ,
         \SB1_1_29/Component_Function_3/NAND4_in[3] ,
         \SB1_1_29/Component_Function_3/NAND4_in[2] ,
         \SB1_1_29/Component_Function_3/NAND4_in[1] ,
         \SB1_1_29/Component_Function_3/NAND4_in[0] ,
         \SB1_1_29/Component_Function_4/NAND4_in[3] ,
         \SB1_1_29/Component_Function_4/NAND4_in[2] ,
         \SB1_1_29/Component_Function_4/NAND4_in[1] ,
         \SB1_1_29/Component_Function_4/NAND4_in[0] ,
         \SB1_1_30/Component_Function_2/NAND4_in[2] ,
         \SB1_1_30/Component_Function_2/NAND4_in[1] ,
         \SB1_1_30/Component_Function_3/NAND4_in[2] ,
         \SB1_1_30/Component_Function_3/NAND4_in[1] ,
         \SB1_1_30/Component_Function_3/NAND4_in[0] ,
         \SB1_1_30/Component_Function_4/NAND4_in[2] ,
         \SB1_1_31/Component_Function_2/NAND4_in[3] ,
         \SB1_1_31/Component_Function_2/NAND4_in[1] ,
         \SB1_1_31/Component_Function_2/NAND4_in[0] ,
         \SB1_1_31/Component_Function_3/NAND4_in[3] ,
         \SB1_1_31/Component_Function_3/NAND4_in[2] ,
         \SB1_1_31/Component_Function_3/NAND4_in[1] ,
         \SB1_1_31/Component_Function_3/NAND4_in[0] ,
         \SB1_1_31/Component_Function_4/NAND4_in[3] ,
         \SB1_1_31/Component_Function_4/NAND4_in[2] ,
         \SB1_1_31/Component_Function_4/NAND4_in[1] ,
         \SB2_1_0/Component_Function_2/NAND4_in[3] ,
         \SB2_1_0/Component_Function_2/NAND4_in[2] ,
         \SB2_1_0/Component_Function_2/NAND4_in[0] ,
         \SB2_1_0/Component_Function_3/NAND4_in[2] ,
         \SB2_1_0/Component_Function_3/NAND4_in[1] ,
         \SB2_1_0/Component_Function_3/NAND4_in[0] ,
         \SB2_1_0/Component_Function_4/NAND4_in[3] ,
         \SB2_1_0/Component_Function_4/NAND4_in[1] ,
         \SB2_1_0/Component_Function_4/NAND4_in[0] ,
         \SB2_1_1/Component_Function_2/NAND4_in[0] ,
         \SB2_1_1/Component_Function_3/NAND4_in[3] ,
         \SB2_1_1/Component_Function_3/NAND4_in[1] ,
         \SB2_1_1/Component_Function_4/NAND4_in[3] ,
         \SB2_1_1/Component_Function_4/NAND4_in[1] ,
         \SB2_1_1/Component_Function_4/NAND4_in[0] ,
         \SB2_1_2/Component_Function_2/NAND4_in[2] ,
         \SB2_1_2/Component_Function_2/NAND4_in[1] ,
         \SB2_1_2/Component_Function_2/NAND4_in[0] ,
         \SB2_1_2/Component_Function_3/NAND4_in[3] ,
         \SB2_1_2/Component_Function_3/NAND4_in[2] ,
         \SB2_1_2/Component_Function_3/NAND4_in[1] ,
         \SB2_1_2/Component_Function_4/NAND4_in[2] ,
         \SB2_1_2/Component_Function_4/NAND4_in[1] ,
         \SB2_1_2/Component_Function_4/NAND4_in[0] ,
         \SB2_1_3/Component_Function_2/NAND4_in[2] ,
         \SB2_1_3/Component_Function_2/NAND4_in[1] ,
         \SB2_1_3/Component_Function_2/NAND4_in[0] ,
         \SB2_1_3/Component_Function_3/NAND4_in[3] ,
         \SB2_1_3/Component_Function_3/NAND4_in[1] ,
         \SB2_1_3/Component_Function_3/NAND4_in[0] ,
         \SB2_1_3/Component_Function_4/NAND4_in[2] ,
         \SB2_1_3/Component_Function_4/NAND4_in[1] ,
         \SB2_1_3/Component_Function_4/NAND4_in[0] ,
         \SB2_1_4/Component_Function_2/NAND4_in[3] ,
         \SB2_1_4/Component_Function_2/NAND4_in[1] ,
         \SB2_1_4/Component_Function_2/NAND4_in[0] ,
         \SB2_1_4/Component_Function_3/NAND4_in[3] ,
         \SB2_1_4/Component_Function_3/NAND4_in[2] ,
         \SB2_1_4/Component_Function_3/NAND4_in[0] ,
         \SB2_1_4/Component_Function_4/NAND4_in[3] ,
         \SB2_1_4/Component_Function_4/NAND4_in[2] ,
         \SB2_1_4/Component_Function_4/NAND4_in[1] ,
         \SB2_1_4/Component_Function_4/NAND4_in[0] ,
         \SB2_1_5/Component_Function_2/NAND4_in[2] ,
         \SB2_1_5/Component_Function_2/NAND4_in[0] ,
         \SB2_1_5/Component_Function_3/NAND4_in[3] ,
         \SB2_1_5/Component_Function_4/NAND4_in[3] ,
         \SB2_1_5/Component_Function_4/NAND4_in[1] ,
         \SB2_1_5/Component_Function_4/NAND4_in[0] ,
         \SB2_1_6/Component_Function_2/NAND4_in[1] ,
         \SB2_1_6/Component_Function_2/NAND4_in[0] ,
         \SB2_1_6/Component_Function_3/NAND4_in[3] ,
         \SB2_1_6/Component_Function_3/NAND4_in[2] ,
         \SB2_1_6/Component_Function_3/NAND4_in[1] ,
         \SB2_1_6/Component_Function_3/NAND4_in[0] ,
         \SB2_1_6/Component_Function_4/NAND4_in[3] ,
         \SB2_1_6/Component_Function_4/NAND4_in[2] ,
         \SB2_1_6/Component_Function_4/NAND4_in[1] ,
         \SB2_1_6/Component_Function_4/NAND4_in[0] ,
         \SB2_1_7/Component_Function_2/NAND4_in[2] ,
         \SB2_1_7/Component_Function_2/NAND4_in[1] ,
         \SB2_1_7/Component_Function_2/NAND4_in[0] ,
         \SB2_1_7/Component_Function_3/NAND4_in[3] ,
         \SB2_1_7/Component_Function_3/NAND4_in[2] ,
         \SB2_1_7/Component_Function_3/NAND4_in[0] ,
         \SB2_1_7/Component_Function_4/NAND4_in[2] ,
         \SB2_1_7/Component_Function_4/NAND4_in[1] ,
         \SB2_1_7/Component_Function_4/NAND4_in[0] ,
         \SB2_1_8/Component_Function_2/NAND4_in[2] ,
         \SB2_1_8/Component_Function_2/NAND4_in[0] ,
         \SB2_1_8/Component_Function_3/NAND4_in[3] ,
         \SB2_1_8/Component_Function_3/NAND4_in[0] ,
         \SB2_1_8/Component_Function_4/NAND4_in[2] ,
         \SB2_1_8/Component_Function_4/NAND4_in[1] ,
         \SB2_1_8/Component_Function_4/NAND4_in[0] ,
         \SB2_1_9/Component_Function_2/NAND4_in[2] ,
         \SB2_1_9/Component_Function_3/NAND4_in[3] ,
         \SB2_1_9/Component_Function_3/NAND4_in[2] ,
         \SB2_1_9/Component_Function_4/NAND4_in[3] ,
         \SB2_1_9/Component_Function_4/NAND4_in[2] ,
         \SB2_1_9/Component_Function_4/NAND4_in[1] ,
         \SB2_1_10/Component_Function_2/NAND4_in[2] ,
         \SB2_1_10/Component_Function_2/NAND4_in[1] ,
         \SB2_1_10/Component_Function_2/NAND4_in[0] ,
         \SB2_1_10/Component_Function_3/NAND4_in[3] ,
         \SB2_1_10/Component_Function_3/NAND4_in[2] ,
         \SB2_1_10/Component_Function_3/NAND4_in[0] ,
         \SB2_1_10/Component_Function_4/NAND4_in[3] ,
         \SB2_1_11/Component_Function_2/NAND4_in[3] ,
         \SB2_1_11/Component_Function_2/NAND4_in[2] ,
         \SB2_1_11/Component_Function_2/NAND4_in[1] ,
         \SB2_1_11/Component_Function_3/NAND4_in[3] ,
         \SB2_1_11/Component_Function_3/NAND4_in[2] ,
         \SB2_1_11/Component_Function_3/NAND4_in[1] ,
         \SB2_1_11/Component_Function_3/NAND4_in[0] ,
         \SB2_1_11/Component_Function_4/NAND4_in[3] ,
         \SB2_1_11/Component_Function_4/NAND4_in[1] ,
         \SB2_1_11/Component_Function_4/NAND4_in[0] ,
         \SB2_1_12/Component_Function_2/NAND4_in[2] ,
         \SB2_1_12/Component_Function_2/NAND4_in[1] ,
         \SB2_1_12/Component_Function_2/NAND4_in[0] ,
         \SB2_1_12/Component_Function_3/NAND4_in[3] ,
         \SB2_1_12/Component_Function_3/NAND4_in[2] ,
         \SB2_1_12/Component_Function_3/NAND4_in[1] ,
         \SB2_1_12/Component_Function_3/NAND4_in[0] ,
         \SB2_1_12/Component_Function_4/NAND4_in[3] ,
         \SB2_1_12/Component_Function_4/NAND4_in[1] ,
         \SB2_1_12/Component_Function_4/NAND4_in[0] ,
         \SB2_1_13/Component_Function_2/NAND4_in[2] ,
         \SB2_1_13/Component_Function_2/NAND4_in[1] ,
         \SB2_1_13/Component_Function_2/NAND4_in[0] ,
         \SB2_1_13/Component_Function_3/NAND4_in[2] ,
         \SB2_1_13/Component_Function_3/NAND4_in[1] ,
         \SB2_1_13/Component_Function_3/NAND4_in[0] ,
         \SB2_1_13/Component_Function_4/NAND4_in[3] ,
         \SB2_1_13/Component_Function_4/NAND4_in[1] ,
         \SB2_1_13/Component_Function_4/NAND4_in[0] ,
         \SB2_1_14/Component_Function_2/NAND4_in[2] ,
         \SB2_1_14/Component_Function_3/NAND4_in[2] ,
         \SB2_1_14/Component_Function_3/NAND4_in[1] ,
         \SB2_1_14/Component_Function_3/NAND4_in[0] ,
         \SB2_1_14/Component_Function_4/NAND4_in[3] ,
         \SB2_1_14/Component_Function_4/NAND4_in[1] ,
         \SB2_1_14/Component_Function_4/NAND4_in[0] ,
         \SB2_1_15/Component_Function_2/NAND4_in[0] ,
         \SB2_1_15/Component_Function_3/NAND4_in[3] ,
         \SB2_1_15/Component_Function_3/NAND4_in[2] ,
         \SB2_1_15/Component_Function_3/NAND4_in[1] ,
         \SB2_1_15/Component_Function_4/NAND4_in[2] ,
         \SB2_1_15/Component_Function_4/NAND4_in[1] ,
         \SB2_1_15/Component_Function_4/NAND4_in[0] ,
         \SB2_1_16/Component_Function_2/NAND4_in[1] ,
         \SB2_1_16/Component_Function_2/NAND4_in[0] ,
         \SB2_1_16/Component_Function_3/NAND4_in[3] ,
         \SB2_1_16/Component_Function_3/NAND4_in[1] ,
         \SB2_1_16/Component_Function_3/NAND4_in[0] ,
         \SB2_1_16/Component_Function_4/NAND4_in[3] ,
         \SB2_1_16/Component_Function_4/NAND4_in[2] ,
         \SB2_1_16/Component_Function_4/NAND4_in[1] ,
         \SB2_1_16/Component_Function_4/NAND4_in[0] ,
         \SB2_1_17/Component_Function_2/NAND4_in[3] ,
         \SB2_1_17/Component_Function_2/NAND4_in[2] ,
         \SB2_1_17/Component_Function_2/NAND4_in[0] ,
         \SB2_1_17/Component_Function_3/NAND4_in[3] ,
         \SB2_1_17/Component_Function_3/NAND4_in[1] ,
         \SB2_1_17/Component_Function_3/NAND4_in[0] ,
         \SB2_1_17/Component_Function_4/NAND4_in[3] ,
         \SB2_1_17/Component_Function_4/NAND4_in[0] ,
         \SB2_1_18/Component_Function_2/NAND4_in[3] ,
         \SB2_1_18/Component_Function_2/NAND4_in[2] ,
         \SB2_1_18/Component_Function_2/NAND4_in[0] ,
         \SB2_1_18/Component_Function_3/NAND4_in[1] ,
         \SB2_1_18/Component_Function_3/NAND4_in[0] ,
         \SB2_1_18/Component_Function_4/NAND4_in[3] ,
         \SB2_1_18/Component_Function_4/NAND4_in[2] ,
         \SB2_1_18/Component_Function_4/NAND4_in[1] ,
         \SB2_1_18/Component_Function_4/NAND4_in[0] ,
         \SB2_1_19/Component_Function_2/NAND4_in[2] ,
         \SB2_1_19/Component_Function_2/NAND4_in[1] ,
         \SB2_1_19/Component_Function_3/NAND4_in[2] ,
         \SB2_1_19/Component_Function_3/NAND4_in[1] ,
         \SB2_1_19/Component_Function_3/NAND4_in[0] ,
         \SB2_1_19/Component_Function_4/NAND4_in[1] ,
         \SB2_1_19/Component_Function_4/NAND4_in[0] ,
         \SB2_1_20/Component_Function_2/NAND4_in[3] ,
         \SB2_1_20/Component_Function_2/NAND4_in[2] ,
         \SB2_1_20/Component_Function_2/NAND4_in[0] ,
         \SB2_1_20/Component_Function_3/NAND4_in[3] ,
         \SB2_1_20/Component_Function_3/NAND4_in[0] ,
         \SB2_1_20/Component_Function_4/NAND4_in[3] ,
         \SB2_1_20/Component_Function_4/NAND4_in[1] ,
         \SB2_1_20/Component_Function_4/NAND4_in[0] ,
         \SB2_1_21/Component_Function_2/NAND4_in[2] ,
         \SB2_1_21/Component_Function_2/NAND4_in[0] ,
         \SB2_1_21/Component_Function_3/NAND4_in[2] ,
         \SB2_1_21/Component_Function_4/NAND4_in[3] ,
         \SB2_1_21/Component_Function_4/NAND4_in[1] ,
         \SB2_1_21/Component_Function_4/NAND4_in[0] ,
         \SB2_1_22/Component_Function_2/NAND4_in[2] ,
         \SB2_1_22/Component_Function_2/NAND4_in[1] ,
         \SB2_1_22/Component_Function_2/NAND4_in[0] ,
         \SB2_1_22/Component_Function_3/NAND4_in[3] ,
         \SB2_1_22/Component_Function_3/NAND4_in[2] ,
         \SB2_1_22/Component_Function_3/NAND4_in[1] ,
         \SB2_1_22/Component_Function_3/NAND4_in[0] ,
         \SB2_1_22/Component_Function_4/NAND4_in[3] ,
         \SB2_1_22/Component_Function_4/NAND4_in[1] ,
         \SB2_1_22/Component_Function_4/NAND4_in[0] ,
         \SB2_1_23/Component_Function_2/NAND4_in[2] ,
         \SB2_1_23/Component_Function_2/NAND4_in[1] ,
         \SB2_1_23/Component_Function_3/NAND4_in[3] ,
         \SB2_1_23/Component_Function_3/NAND4_in[2] ,
         \SB2_1_23/Component_Function_3/NAND4_in[1] ,
         \SB2_1_23/Component_Function_3/NAND4_in[0] ,
         \SB2_1_23/Component_Function_4/NAND4_in[3] ,
         \SB2_1_23/Component_Function_4/NAND4_in[2] ,
         \SB2_1_23/Component_Function_4/NAND4_in[1] ,
         \SB2_1_23/Component_Function_4/NAND4_in[0] ,
         \SB2_1_24/Component_Function_2/NAND4_in[3] ,
         \SB2_1_24/Component_Function_2/NAND4_in[2] ,
         \SB2_1_24/Component_Function_2/NAND4_in[1] ,
         \SB2_1_24/Component_Function_2/NAND4_in[0] ,
         \SB2_1_24/Component_Function_3/NAND4_in[3] ,
         \SB2_1_24/Component_Function_3/NAND4_in[1] ,
         \SB2_1_24/Component_Function_3/NAND4_in[0] ,
         \SB2_1_24/Component_Function_4/NAND4_in[3] ,
         \SB2_1_24/Component_Function_4/NAND4_in[1] ,
         \SB2_1_24/Component_Function_4/NAND4_in[0] ,
         \SB2_1_25/Component_Function_2/NAND4_in[1] ,
         \SB2_1_25/Component_Function_3/NAND4_in[3] ,
         \SB2_1_25/Component_Function_3/NAND4_in[0] ,
         \SB2_1_25/Component_Function_4/NAND4_in[2] ,
         \SB2_1_25/Component_Function_4/NAND4_in[1] ,
         \SB2_1_25/Component_Function_4/NAND4_in[0] ,
         \SB2_1_26/Component_Function_2/NAND4_in[2] ,
         \SB2_1_26/Component_Function_2/NAND4_in[0] ,
         \SB2_1_26/Component_Function_3/NAND4_in[3] ,
         \SB2_1_26/Component_Function_3/NAND4_in[2] ,
         \SB2_1_26/Component_Function_3/NAND4_in[1] ,
         \SB2_1_26/Component_Function_3/NAND4_in[0] ,
         \SB2_1_26/Component_Function_4/NAND4_in[3] ,
         \SB2_1_26/Component_Function_4/NAND4_in[1] ,
         \SB2_1_26/Component_Function_4/NAND4_in[0] ,
         \SB2_1_27/Component_Function_2/NAND4_in[2] ,
         \SB2_1_27/Component_Function_2/NAND4_in[0] ,
         \SB2_1_27/Component_Function_3/NAND4_in[3] ,
         \SB2_1_27/Component_Function_3/NAND4_in[1] ,
         \SB2_1_27/Component_Function_3/NAND4_in[0] ,
         \SB2_1_27/Component_Function_4/NAND4_in[3] ,
         \SB2_1_27/Component_Function_4/NAND4_in[1] ,
         \SB2_1_27/Component_Function_4/NAND4_in[0] ,
         \SB2_1_28/Component_Function_2/NAND4_in[1] ,
         \SB2_1_28/Component_Function_2/NAND4_in[0] ,
         \SB2_1_28/Component_Function_3/NAND4_in[2] ,
         \SB2_1_28/Component_Function_3/NAND4_in[1] ,
         \SB2_1_28/Component_Function_3/NAND4_in[0] ,
         \SB2_1_28/Component_Function_4/NAND4_in[3] ,
         \SB2_1_28/Component_Function_4/NAND4_in[2] ,
         \SB2_1_28/Component_Function_4/NAND4_in[1] ,
         \SB2_1_28/Component_Function_4/NAND4_in[0] ,
         \SB2_1_29/Component_Function_2/NAND4_in[2] ,
         \SB2_1_29/Component_Function_2/NAND4_in[1] ,
         \SB2_1_29/Component_Function_2/NAND4_in[0] ,
         \SB2_1_29/Component_Function_3/NAND4_in[3] ,
         \SB2_1_29/Component_Function_3/NAND4_in[1] ,
         \SB2_1_29/Component_Function_3/NAND4_in[0] ,
         \SB2_1_29/Component_Function_4/NAND4_in[3] ,
         \SB2_1_29/Component_Function_4/NAND4_in[1] ,
         \SB2_1_29/Component_Function_4/NAND4_in[0] ,
         \SB2_1_30/Component_Function_2/NAND4_in[2] ,
         \SB2_1_30/Component_Function_2/NAND4_in[1] ,
         \SB2_1_30/Component_Function_2/NAND4_in[0] ,
         \SB2_1_30/Component_Function_3/NAND4_in[3] ,
         \SB2_1_30/Component_Function_3/NAND4_in[2] ,
         \SB2_1_30/Component_Function_3/NAND4_in[1] ,
         \SB2_1_30/Component_Function_3/NAND4_in[0] ,
         \SB2_1_30/Component_Function_4/NAND4_in[3] ,
         \SB2_1_30/Component_Function_4/NAND4_in[2] ,
         \SB2_1_30/Component_Function_4/NAND4_in[1] ,
         \SB2_1_30/Component_Function_4/NAND4_in[0] ,
         \SB2_1_31/Component_Function_2/NAND4_in[1] ,
         \SB2_1_31/Component_Function_2/NAND4_in[0] ,
         \SB2_1_31/Component_Function_3/NAND4_in[3] ,
         \SB2_1_31/Component_Function_3/NAND4_in[2] ,
         \SB2_1_31/Component_Function_3/NAND4_in[1] ,
         \SB2_1_31/Component_Function_3/NAND4_in[0] ,
         \SB2_1_31/Component_Function_4/NAND4_in[2] ,
         \SB2_1_31/Component_Function_4/NAND4_in[1] ,
         \SB1_2_0/Component_Function_2/NAND4_in[1] ,
         \SB1_2_0/Component_Function_2/NAND4_in[0] ,
         \SB1_2_0/Component_Function_3/NAND4_in[2] ,
         \SB1_2_0/Component_Function_3/NAND4_in[0] ,
         \SB1_2_0/Component_Function_4/NAND4_in[2] ,
         \SB1_2_0/Component_Function_4/NAND4_in[1] ,
         \SB1_2_0/Component_Function_4/NAND4_in[0] ,
         \SB1_2_1/Component_Function_2/NAND4_in[3] ,
         \SB1_2_1/Component_Function_2/NAND4_in[2] ,
         \SB1_2_1/Component_Function_2/NAND4_in[0] ,
         \SB1_2_1/Component_Function_3/NAND4_in[3] ,
         \SB1_2_1/Component_Function_3/NAND4_in[1] ,
         \SB1_2_1/Component_Function_3/NAND4_in[0] ,
         \SB1_2_1/Component_Function_4/NAND4_in[2] ,
         \SB1_2_1/Component_Function_4/NAND4_in[1] ,
         \SB1_2_1/Component_Function_4/NAND4_in[0] ,
         \SB1_2_2/Component_Function_2/NAND4_in[3] ,
         \SB1_2_2/Component_Function_2/NAND4_in[2] ,
         \SB1_2_2/Component_Function_2/NAND4_in[0] ,
         \SB1_2_2/Component_Function_3/NAND4_in[2] ,
         \SB1_2_2/Component_Function_3/NAND4_in[1] ,
         \SB1_2_2/Component_Function_3/NAND4_in[0] ,
         \SB1_2_2/Component_Function_4/NAND4_in[3] ,
         \SB1_2_2/Component_Function_4/NAND4_in[2] ,
         \SB1_2_2/Component_Function_4/NAND4_in[1] ,
         \SB1_2_3/Component_Function_2/NAND4_in[3] ,
         \SB1_2_3/Component_Function_2/NAND4_in[1] ,
         \SB1_2_3/Component_Function_3/NAND4_in[2] ,
         \SB1_2_3/Component_Function_3/NAND4_in[1] ,
         \SB1_2_3/Component_Function_3/NAND4_in[0] ,
         \SB1_2_3/Component_Function_4/NAND4_in[3] ,
         \SB1_2_3/Component_Function_4/NAND4_in[2] ,
         \SB1_2_3/Component_Function_4/NAND4_in[0] ,
         \SB1_2_4/Component_Function_2/NAND4_in[2] ,
         \SB1_2_4/Component_Function_2/NAND4_in[0] ,
         \SB1_2_4/Component_Function_3/NAND4_in[0] ,
         \SB1_2_4/Component_Function_4/NAND4_in[3] ,
         \SB1_2_4/Component_Function_4/NAND4_in[2] ,
         \SB1_2_5/Component_Function_2/NAND4_in[3] ,
         \SB1_2_5/Component_Function_2/NAND4_in[2] ,
         \SB1_2_5/Component_Function_2/NAND4_in[1] ,
         \SB1_2_5/Component_Function_3/NAND4_in[1] ,
         \SB1_2_5/Component_Function_3/NAND4_in[0] ,
         \SB1_2_5/Component_Function_4/NAND4_in[3] ,
         \SB1_2_5/Component_Function_4/NAND4_in[2] ,
         \SB1_2_5/Component_Function_4/NAND4_in[1] ,
         \SB1_2_5/Component_Function_4/NAND4_in[0] ,
         \SB1_2_6/Component_Function_2/NAND4_in[3] ,
         \SB1_2_6/Component_Function_3/NAND4_in[2] ,
         \SB1_2_6/Component_Function_3/NAND4_in[1] ,
         \SB1_2_6/Component_Function_3/NAND4_in[0] ,
         \SB1_2_6/Component_Function_4/NAND4_in[3] ,
         \SB1_2_6/Component_Function_4/NAND4_in[2] ,
         \SB1_2_6/Component_Function_4/NAND4_in[1] ,
         \SB1_2_6/Component_Function_4/NAND4_in[0] ,
         \SB1_2_7/Component_Function_2/NAND4_in[1] ,
         \SB1_2_7/Component_Function_2/NAND4_in[0] ,
         \SB1_2_7/Component_Function_3/NAND4_in[1] ,
         \SB1_2_7/Component_Function_3/NAND4_in[0] ,
         \SB1_2_7/Component_Function_4/NAND4_in[3] ,
         \SB1_2_7/Component_Function_4/NAND4_in[1] ,
         \SB1_2_7/Component_Function_4/NAND4_in[0] ,
         \SB1_2_8/Component_Function_2/NAND4_in[2] ,
         \SB1_2_8/Component_Function_2/NAND4_in[1] ,
         \SB1_2_8/Component_Function_3/NAND4_in[3] ,
         \SB1_2_8/Component_Function_3/NAND4_in[1] ,
         \SB1_2_8/Component_Function_3/NAND4_in[0] ,
         \SB1_2_8/Component_Function_4/NAND4_in[3] ,
         \SB1_2_8/Component_Function_4/NAND4_in[0] ,
         \SB1_2_9/Component_Function_2/NAND4_in[2] ,
         \SB1_2_9/Component_Function_2/NAND4_in[1] ,
         \SB1_2_9/Component_Function_3/NAND4_in[1] ,
         \SB1_2_9/Component_Function_3/NAND4_in[0] ,
         \SB1_2_9/Component_Function_4/NAND4_in[3] ,
         \SB1_2_10/Component_Function_2/NAND4_in[2] ,
         \SB1_2_10/Component_Function_2/NAND4_in[1] ,
         \SB1_2_10/Component_Function_3/NAND4_in[2] ,
         \SB1_2_10/Component_Function_3/NAND4_in[1] ,
         \SB1_2_10/Component_Function_3/NAND4_in[0] ,
         \SB1_2_10/Component_Function_4/NAND4_in[3] ,
         \SB1_2_11/Component_Function_2/NAND4_in[2] ,
         \SB1_2_11/Component_Function_2/NAND4_in[1] ,
         \SB1_2_11/Component_Function_2/NAND4_in[0] ,
         \SB1_2_11/Component_Function_3/NAND4_in[3] ,
         \SB1_2_11/Component_Function_3/NAND4_in[2] ,
         \SB1_2_11/Component_Function_3/NAND4_in[1] ,
         \SB1_2_11/Component_Function_3/NAND4_in[0] ,
         \SB1_2_12/Component_Function_2/NAND4_in[2] ,
         \SB1_2_12/Component_Function_2/NAND4_in[0] ,
         \SB1_2_12/Component_Function_3/NAND4_in[2] ,
         \SB1_2_12/Component_Function_3/NAND4_in[1] ,
         \SB1_2_12/Component_Function_4/NAND4_in[3] ,
         \SB1_2_12/Component_Function_4/NAND4_in[2] ,
         \SB1_2_12/Component_Function_4/NAND4_in[0] ,
         \SB1_2_13/Component_Function_2/NAND4_in[1] ,
         \SB1_2_13/Component_Function_2/NAND4_in[0] ,
         \SB1_2_13/Component_Function_3/NAND4_in[3] ,
         \SB1_2_13/Component_Function_3/NAND4_in[1] ,
         \SB1_2_13/Component_Function_4/NAND4_in[3] ,
         \SB1_2_13/Component_Function_4/NAND4_in[1] ,
         \SB1_2_13/Component_Function_4/NAND4_in[0] ,
         \SB1_2_14/Component_Function_2/NAND4_in[2] ,
         \SB1_2_14/Component_Function_2/NAND4_in[1] ,
         \SB1_2_14/Component_Function_2/NAND4_in[0] ,
         \SB1_2_14/Component_Function_3/NAND4_in[3] ,
         \SB1_2_14/Component_Function_3/NAND4_in[1] ,
         \SB1_2_14/Component_Function_3/NAND4_in[0] ,
         \SB1_2_14/Component_Function_4/NAND4_in[2] ,
         \SB1_2_14/Component_Function_4/NAND4_in[0] ,
         \SB1_2_15/Component_Function_2/NAND4_in[2] ,
         \SB1_2_15/Component_Function_2/NAND4_in[1] ,
         \SB1_2_15/Component_Function_2/NAND4_in[0] ,
         \SB1_2_15/Component_Function_3/NAND4_in[1] ,
         \SB1_2_15/Component_Function_3/NAND4_in[0] ,
         \SB1_2_15/Component_Function_4/NAND4_in[3] ,
         \SB1_2_16/Component_Function_2/NAND4_in[2] ,
         \SB1_2_16/Component_Function_2/NAND4_in[1] ,
         \SB1_2_16/Component_Function_2/NAND4_in[0] ,
         \SB1_2_16/Component_Function_3/NAND4_in[3] ,
         \SB1_2_16/Component_Function_3/NAND4_in[1] ,
         \SB1_2_16/Component_Function_4/NAND4_in[3] ,
         \SB1_2_16/Component_Function_4/NAND4_in[2] ,
         \SB1_2_16/Component_Function_4/NAND4_in[1] ,
         \SB1_2_16/Component_Function_4/NAND4_in[0] ,
         \SB1_2_17/Component_Function_2/NAND4_in[3] ,
         \SB1_2_17/Component_Function_2/NAND4_in[2] ,
         \SB1_2_17/Component_Function_2/NAND4_in[0] ,
         \SB1_2_17/Component_Function_3/NAND4_in[2] ,
         \SB1_2_17/Component_Function_3/NAND4_in[1] ,
         \SB1_2_17/Component_Function_3/NAND4_in[0] ,
         \SB1_2_17/Component_Function_4/NAND4_in[3] ,
         \SB1_2_17/Component_Function_4/NAND4_in[1] ,
         \SB1_2_17/Component_Function_4/NAND4_in[0] ,
         \SB1_2_18/Component_Function_2/NAND4_in[3] ,
         \SB1_2_18/Component_Function_2/NAND4_in[2] ,
         \SB1_2_18/Component_Function_2/NAND4_in[0] ,
         \SB1_2_18/Component_Function_3/NAND4_in[2] ,
         \SB1_2_18/Component_Function_3/NAND4_in[1] ,
         \SB1_2_18/Component_Function_4/NAND4_in[3] ,
         \SB1_2_18/Component_Function_4/NAND4_in[2] ,
         \SB1_2_18/Component_Function_4/NAND4_in[1] ,
         \SB1_2_18/Component_Function_4/NAND4_in[0] ,
         \SB1_2_19/Component_Function_2/NAND4_in[3] ,
         \SB1_2_19/Component_Function_2/NAND4_in[1] ,
         \SB1_2_19/Component_Function_2/NAND4_in[0] ,
         \SB1_2_19/Component_Function_3/NAND4_in[3] ,
         \SB1_2_19/Component_Function_3/NAND4_in[1] ,
         \SB1_2_19/Component_Function_3/NAND4_in[0] ,
         \SB1_2_19/Component_Function_4/NAND4_in[3] ,
         \SB1_2_19/Component_Function_4/NAND4_in[2] ,
         \SB1_2_19/Component_Function_4/NAND4_in[1] ,
         \SB1_2_19/Component_Function_4/NAND4_in[0] ,
         \SB1_2_20/Component_Function_2/NAND4_in[1] ,
         \SB1_2_20/Component_Function_3/NAND4_in[3] ,
         \SB1_2_20/Component_Function_3/NAND4_in[1] ,
         \SB1_2_20/Component_Function_3/NAND4_in[0] ,
         \SB1_2_20/Component_Function_4/NAND4_in[3] ,
         \SB1_2_20/Component_Function_4/NAND4_in[2] ,
         \SB1_2_20/Component_Function_4/NAND4_in[1] ,
         \SB1_2_20/Component_Function_4/NAND4_in[0] ,
         \SB1_2_21/Component_Function_2/NAND4_in[3] ,
         \SB1_2_21/Component_Function_2/NAND4_in[2] ,
         \SB1_2_21/Component_Function_2/NAND4_in[0] ,
         \SB1_2_21/Component_Function_3/NAND4_in[3] ,
         \SB1_2_21/Component_Function_3/NAND4_in[1] ,
         \SB1_2_21/Component_Function_3/NAND4_in[0] ,
         \SB1_2_21/Component_Function_4/NAND4_in[3] ,
         \SB1_2_21/Component_Function_4/NAND4_in[0] ,
         \SB1_2_22/Component_Function_2/NAND4_in[2] ,
         \SB1_2_22/Component_Function_2/NAND4_in[1] ,
         \SB1_2_22/Component_Function_2/NAND4_in[0] ,
         \SB1_2_22/Component_Function_3/NAND4_in[3] ,
         \SB1_2_22/Component_Function_3/NAND4_in[1] ,
         \SB1_2_22/Component_Function_3/NAND4_in[0] ,
         \SB1_2_22/Component_Function_4/NAND4_in[3] ,
         \SB1_2_22/Component_Function_4/NAND4_in[2] ,
         \SB1_2_22/Component_Function_4/NAND4_in[1] ,
         \SB1_2_22/Component_Function_4/NAND4_in[0] ,
         \SB1_2_23/Component_Function_2/NAND4_in[3] ,
         \SB1_2_23/Component_Function_2/NAND4_in[2] ,
         \SB1_2_23/Component_Function_2/NAND4_in[1] ,
         \SB1_2_23/Component_Function_2/NAND4_in[0] ,
         \SB1_2_23/Component_Function_3/NAND4_in[2] ,
         \SB1_2_23/Component_Function_3/NAND4_in[0] ,
         \SB1_2_23/Component_Function_4/NAND4_in[3] ,
         \SB1_2_23/Component_Function_4/NAND4_in[2] ,
         \SB1_2_23/Component_Function_4/NAND4_in[1] ,
         \SB1_2_23/Component_Function_4/NAND4_in[0] ,
         \SB1_2_24/Component_Function_2/NAND4_in[3] ,
         \SB1_2_24/Component_Function_2/NAND4_in[2] ,
         \SB1_2_24/Component_Function_2/NAND4_in[0] ,
         \SB1_2_24/Component_Function_3/NAND4_in[1] ,
         \SB1_2_24/Component_Function_3/NAND4_in[0] ,
         \SB1_2_24/Component_Function_4/NAND4_in[2] ,
         \SB1_2_24/Component_Function_4/NAND4_in[1] ,
         \SB1_2_24/Component_Function_4/NAND4_in[0] ,
         \SB1_2_25/Component_Function_2/NAND4_in[2] ,
         \SB1_2_25/Component_Function_2/NAND4_in[1] ,
         \SB1_2_25/Component_Function_2/NAND4_in[0] ,
         \SB1_2_25/Component_Function_3/NAND4_in[2] ,
         \SB1_2_25/Component_Function_3/NAND4_in[1] ,
         \SB1_2_25/Component_Function_3/NAND4_in[0] ,
         \SB1_2_25/Component_Function_4/NAND4_in[3] ,
         \SB1_2_25/Component_Function_4/NAND4_in[1] ,
         \SB1_2_25/Component_Function_4/NAND4_in[0] ,
         \SB1_2_26/Component_Function_2/NAND4_in[2] ,
         \SB1_2_26/Component_Function_2/NAND4_in[1] ,
         \SB1_2_26/Component_Function_2/NAND4_in[0] ,
         \SB1_2_26/Component_Function_3/NAND4_in[3] ,
         \SB1_2_26/Component_Function_3/NAND4_in[0] ,
         \SB1_2_26/Component_Function_4/NAND4_in[1] ,
         \SB1_2_26/Component_Function_4/NAND4_in[0] ,
         \SB1_2_27/Component_Function_2/NAND4_in[2] ,
         \SB1_2_27/Component_Function_2/NAND4_in[1] ,
         \SB1_2_27/Component_Function_2/NAND4_in[0] ,
         \SB1_2_27/Component_Function_3/NAND4_in[3] ,
         \SB1_2_27/Component_Function_3/NAND4_in[1] ,
         \SB1_2_27/Component_Function_3/NAND4_in[0] ,
         \SB1_2_27/Component_Function_4/NAND4_in[2] ,
         \SB1_2_27/Component_Function_4/NAND4_in[1] ,
         \SB1_2_27/Component_Function_4/NAND4_in[0] ,
         \SB1_2_28/Component_Function_2/NAND4_in[2] ,
         \SB1_2_28/Component_Function_2/NAND4_in[1] ,
         \SB1_2_28/Component_Function_2/NAND4_in[0] ,
         \SB1_2_28/Component_Function_3/NAND4_in[3] ,
         \SB1_2_28/Component_Function_3/NAND4_in[1] ,
         \SB1_2_28/Component_Function_3/NAND4_in[0] ,
         \SB1_2_28/Component_Function_4/NAND4_in[3] ,
         \SB1_2_28/Component_Function_4/NAND4_in[2] ,
         \SB1_2_28/Component_Function_4/NAND4_in[0] ,
         \SB1_2_29/Component_Function_2/NAND4_in[1] ,
         \SB1_2_29/Component_Function_2/NAND4_in[0] ,
         \SB1_2_29/Component_Function_3/NAND4_in[2] ,
         \SB1_2_29/Component_Function_3/NAND4_in[0] ,
         \SB1_2_29/Component_Function_4/NAND4_in[3] ,
         \SB1_2_29/Component_Function_4/NAND4_in[2] ,
         \SB1_2_30/Component_Function_2/NAND4_in[2] ,
         \SB1_2_30/Component_Function_2/NAND4_in[1] ,
         \SB1_2_30/Component_Function_2/NAND4_in[0] ,
         \SB1_2_30/Component_Function_3/NAND4_in[1] ,
         \SB1_2_30/Component_Function_3/NAND4_in[0] ,
         \SB1_2_30/Component_Function_4/NAND4_in[1] ,
         \SB1_2_30/Component_Function_4/NAND4_in[0] ,
         \SB1_2_31/Component_Function_2/NAND4_in[3] ,
         \SB1_2_31/Component_Function_2/NAND4_in[1] ,
         \SB1_2_31/Component_Function_2/NAND4_in[0] ,
         \SB1_2_31/Component_Function_3/NAND4_in[2] ,
         \SB1_2_31/Component_Function_3/NAND4_in[0] ,
         \SB1_2_31/Component_Function_4/NAND4_in[3] ,
         \SB1_2_31/Component_Function_4/NAND4_in[2] ,
         \SB1_2_31/Component_Function_4/NAND4_in[1] ,
         \SB2_2_0/Component_Function_2/NAND4_in[3] ,
         \SB2_2_0/Component_Function_2/NAND4_in[2] ,
         \SB2_2_0/Component_Function_2/NAND4_in[1] ,
         \SB2_2_0/Component_Function_2/NAND4_in[0] ,
         \SB2_2_0/Component_Function_3/NAND4_in[3] ,
         \SB2_2_0/Component_Function_3/NAND4_in[1] ,
         \SB2_2_0/Component_Function_4/NAND4_in[3] ,
         \SB2_2_0/Component_Function_4/NAND4_in[2] ,
         \SB2_2_0/Component_Function_4/NAND4_in[1] ,
         \SB2_2_0/Component_Function_4/NAND4_in[0] ,
         \SB2_2_1/Component_Function_2/NAND4_in[2] ,
         \SB2_2_1/Component_Function_2/NAND4_in[1] ,
         \SB2_2_1/Component_Function_2/NAND4_in[0] ,
         \SB2_2_1/Component_Function_3/NAND4_in[3] ,
         \SB2_2_1/Component_Function_3/NAND4_in[2] ,
         \SB2_2_1/Component_Function_3/NAND4_in[0] ,
         \SB2_2_1/Component_Function_4/NAND4_in[1] ,
         \SB2_2_1/Component_Function_4/NAND4_in[0] ,
         \SB2_2_2/Component_Function_2/NAND4_in[2] ,
         \SB2_2_2/Component_Function_3/NAND4_in[3] ,
         \SB2_2_2/Component_Function_3/NAND4_in[2] ,
         \SB2_2_2/Component_Function_3/NAND4_in[1] ,
         \SB2_2_2/Component_Function_3/NAND4_in[0] ,
         \SB2_2_2/Component_Function_4/NAND4_in[2] ,
         \SB2_2_2/Component_Function_4/NAND4_in[1] ,
         \SB2_2_2/Component_Function_4/NAND4_in[0] ,
         \SB2_2_3/Component_Function_2/NAND4_in[3] ,
         \SB2_2_3/Component_Function_2/NAND4_in[2] ,
         \SB2_2_3/Component_Function_3/NAND4_in[3] ,
         \SB2_2_3/Component_Function_3/NAND4_in[1] ,
         \SB2_2_3/Component_Function_3/NAND4_in[0] ,
         \SB2_2_3/Component_Function_4/NAND4_in[1] ,
         \SB2_2_3/Component_Function_4/NAND4_in[0] ,
         \SB2_2_4/Component_Function_2/NAND4_in[3] ,
         \SB2_2_4/Component_Function_2/NAND4_in[0] ,
         \SB2_2_4/Component_Function_3/NAND4_in[3] ,
         \SB2_2_4/Component_Function_3/NAND4_in[2] ,
         \SB2_2_4/Component_Function_3/NAND4_in[1] ,
         \SB2_2_4/Component_Function_3/NAND4_in[0] ,
         \SB2_2_4/Component_Function_4/NAND4_in[3] ,
         \SB2_2_4/Component_Function_4/NAND4_in[2] ,
         \SB2_2_4/Component_Function_4/NAND4_in[1] ,
         \SB2_2_4/Component_Function_4/NAND4_in[0] ,
         \SB2_2_5/Component_Function_2/NAND4_in[2] ,
         \SB2_2_5/Component_Function_2/NAND4_in[1] ,
         \SB2_2_5/Component_Function_2/NAND4_in[0] ,
         \SB2_2_5/Component_Function_3/NAND4_in[3] ,
         \SB2_2_5/Component_Function_3/NAND4_in[2] ,
         \SB2_2_5/Component_Function_4/NAND4_in[3] ,
         \SB2_2_5/Component_Function_4/NAND4_in[1] ,
         \SB2_2_5/Component_Function_4/NAND4_in[0] ,
         \SB2_2_6/Component_Function_2/NAND4_in[2] ,
         \SB2_2_6/Component_Function_3/NAND4_in[3] ,
         \SB2_2_6/Component_Function_3/NAND4_in[2] ,
         \SB2_2_6/Component_Function_3/NAND4_in[1] ,
         \SB2_2_6/Component_Function_3/NAND4_in[0] ,
         \SB2_2_6/Component_Function_4/NAND4_in[3] ,
         \SB2_2_6/Component_Function_4/NAND4_in[1] ,
         \SB2_2_7/Component_Function_2/NAND4_in[3] ,
         \SB2_2_7/Component_Function_2/NAND4_in[2] ,
         \SB2_2_7/Component_Function_3/NAND4_in[2] ,
         \SB2_2_7/Component_Function_3/NAND4_in[1] ,
         \SB2_2_7/Component_Function_3/NAND4_in[0] ,
         \SB2_2_7/Component_Function_4/NAND4_in[3] ,
         \SB2_2_7/Component_Function_4/NAND4_in[1] ,
         \SB2_2_7/Component_Function_4/NAND4_in[0] ,
         \SB2_2_8/Component_Function_2/NAND4_in[3] ,
         \SB2_2_8/Component_Function_2/NAND4_in[2] ,
         \SB2_2_8/Component_Function_2/NAND4_in[0] ,
         \SB2_2_8/Component_Function_3/NAND4_in[3] ,
         \SB2_2_8/Component_Function_3/NAND4_in[2] ,
         \SB2_2_8/Component_Function_3/NAND4_in[1] ,
         \SB2_2_8/Component_Function_3/NAND4_in[0] ,
         \SB2_2_8/Component_Function_4/NAND4_in[2] ,
         \SB2_2_8/Component_Function_4/NAND4_in[1] ,
         \SB2_2_8/Component_Function_4/NAND4_in[0] ,
         \SB2_2_9/Component_Function_2/NAND4_in[3] ,
         \SB2_2_9/Component_Function_2/NAND4_in[2] ,
         \SB2_2_9/Component_Function_2/NAND4_in[1] ,
         \SB2_2_9/Component_Function_2/NAND4_in[0] ,
         \SB2_2_9/Component_Function_3/NAND4_in[2] ,
         \SB2_2_9/Component_Function_3/NAND4_in[0] ,
         \SB2_2_9/Component_Function_4/NAND4_in[3] ,
         \SB2_2_9/Component_Function_4/NAND4_in[1] ,
         \SB2_2_9/Component_Function_4/NAND4_in[0] ,
         \SB2_2_10/Component_Function_2/NAND4_in[2] ,
         \SB2_2_10/Component_Function_2/NAND4_in[0] ,
         \SB2_2_10/Component_Function_3/NAND4_in[3] ,
         \SB2_2_10/Component_Function_3/NAND4_in[2] ,
         \SB2_2_10/Component_Function_3/NAND4_in[1] ,
         \SB2_2_10/Component_Function_3/NAND4_in[0] ,
         \SB2_2_10/Component_Function_4/NAND4_in[3] ,
         \SB2_2_10/Component_Function_4/NAND4_in[1] ,
         \SB2_2_10/Component_Function_4/NAND4_in[0] ,
         \SB2_2_11/Component_Function_3/NAND4_in[2] ,
         \SB2_2_11/Component_Function_3/NAND4_in[0] ,
         \SB2_2_11/Component_Function_4/NAND4_in[3] ,
         \SB2_2_11/Component_Function_4/NAND4_in[1] ,
         \SB2_2_11/Component_Function_4/NAND4_in[0] ,
         \SB2_2_12/Component_Function_2/NAND4_in[2] ,
         \SB2_2_12/Component_Function_2/NAND4_in[0] ,
         \SB2_2_12/Component_Function_3/NAND4_in[3] ,
         \SB2_2_12/Component_Function_3/NAND4_in[2] ,
         \SB2_2_12/Component_Function_3/NAND4_in[1] ,
         \SB2_2_12/Component_Function_3/NAND4_in[0] ,
         \SB2_2_12/Component_Function_4/NAND4_in[3] ,
         \SB2_2_12/Component_Function_4/NAND4_in[1] ,
         \SB2_2_12/Component_Function_4/NAND4_in[0] ,
         \SB2_2_13/Component_Function_2/NAND4_in[2] ,
         \SB2_2_13/Component_Function_3/NAND4_in[2] ,
         \SB2_2_13/Component_Function_4/NAND4_in[3] ,
         \SB2_2_13/Component_Function_4/NAND4_in[1] ,
         \SB2_2_14/Component_Function_2/NAND4_in[0] ,
         \SB2_2_14/Component_Function_3/NAND4_in[3] ,
         \SB2_2_14/Component_Function_3/NAND4_in[2] ,
         \SB2_2_14/Component_Function_3/NAND4_in[0] ,
         \SB2_2_14/Component_Function_4/NAND4_in[3] ,
         \SB2_2_14/Component_Function_4/NAND4_in[1] ,
         \SB2_2_14/Component_Function_4/NAND4_in[0] ,
         \SB2_2_15/Component_Function_2/NAND4_in[3] ,
         \SB2_2_15/Component_Function_2/NAND4_in[0] ,
         \SB2_2_15/Component_Function_3/NAND4_in[2] ,
         \SB2_2_15/Component_Function_3/NAND4_in[0] ,
         \SB2_2_15/Component_Function_4/NAND4_in[3] ,
         \SB2_2_15/Component_Function_4/NAND4_in[1] ,
         \SB2_2_15/Component_Function_4/NAND4_in[0] ,
         \SB2_2_16/Component_Function_2/NAND4_in[2] ,
         \SB2_2_16/Component_Function_2/NAND4_in[1] ,
         \SB2_2_16/Component_Function_2/NAND4_in[0] ,
         \SB2_2_16/Component_Function_3/NAND4_in[3] ,
         \SB2_2_16/Component_Function_3/NAND4_in[2] ,
         \SB2_2_16/Component_Function_3/NAND4_in[0] ,
         \SB2_2_16/Component_Function_4/NAND4_in[3] ,
         \SB2_2_16/Component_Function_4/NAND4_in[2] ,
         \SB2_2_16/Component_Function_4/NAND4_in[1] ,
         \SB2_2_16/Component_Function_4/NAND4_in[0] ,
         \SB2_2_17/Component_Function_2/NAND4_in[3] ,
         \SB2_2_17/Component_Function_2/NAND4_in[2] ,
         \SB2_2_17/Component_Function_2/NAND4_in[1] ,
         \SB2_2_17/Component_Function_2/NAND4_in[0] ,
         \SB2_2_17/Component_Function_3/NAND4_in[3] ,
         \SB2_2_17/Component_Function_3/NAND4_in[1] ,
         \SB2_2_17/Component_Function_3/NAND4_in[0] ,
         \SB2_2_17/Component_Function_4/NAND4_in[1] ,
         \SB2_2_17/Component_Function_4/NAND4_in[0] ,
         \SB2_2_18/Component_Function_2/NAND4_in[2] ,
         \SB2_2_18/Component_Function_2/NAND4_in[0] ,
         \SB2_2_18/Component_Function_3/NAND4_in[3] ,
         \SB2_2_18/Component_Function_3/NAND4_in[2] ,
         \SB2_2_18/Component_Function_3/NAND4_in[1] ,
         \SB2_2_18/Component_Function_3/NAND4_in[0] ,
         \SB2_2_18/Component_Function_4/NAND4_in[2] ,
         \SB2_2_18/Component_Function_4/NAND4_in[1] ,
         \SB2_2_18/Component_Function_4/NAND4_in[0] ,
         \SB2_2_19/Component_Function_2/NAND4_in[2] ,
         \SB2_2_19/Component_Function_2/NAND4_in[1] ,
         \SB2_2_19/Component_Function_2/NAND4_in[0] ,
         \SB2_2_19/Component_Function_3/NAND4_in[3] ,
         \SB2_2_19/Component_Function_3/NAND4_in[1] ,
         \SB2_2_19/Component_Function_3/NAND4_in[0] ,
         \SB2_2_19/Component_Function_4/NAND4_in[3] ,
         \SB2_2_19/Component_Function_4/NAND4_in[1] ,
         \SB2_2_19/Component_Function_4/NAND4_in[0] ,
         \SB2_2_20/Component_Function_2/NAND4_in[2] ,
         \SB2_2_20/Component_Function_2/NAND4_in[0] ,
         \SB2_2_20/Component_Function_3/NAND4_in[3] ,
         \SB2_2_20/Component_Function_4/NAND4_in[3] ,
         \SB2_2_20/Component_Function_4/NAND4_in[1] ,
         \SB2_2_20/Component_Function_4/NAND4_in[0] ,
         \SB2_2_21/Component_Function_2/NAND4_in[2] ,
         \SB2_2_21/Component_Function_2/NAND4_in[1] ,
         \SB2_2_21/Component_Function_2/NAND4_in[0] ,
         \SB2_2_21/Component_Function_3/NAND4_in[3] ,
         \SB2_2_21/Component_Function_3/NAND4_in[2] ,
         \SB2_2_21/Component_Function_3/NAND4_in[0] ,
         \SB2_2_21/Component_Function_4/NAND4_in[3] ,
         \SB2_2_22/Component_Function_2/NAND4_in[2] ,
         \SB2_2_22/Component_Function_2/NAND4_in[0] ,
         \SB2_2_22/Component_Function_3/NAND4_in[1] ,
         \SB2_2_22/Component_Function_3/NAND4_in[0] ,
         \SB2_2_22/Component_Function_4/NAND4_in[3] ,
         \SB2_2_22/Component_Function_4/NAND4_in[1] ,
         \SB2_2_22/Component_Function_4/NAND4_in[0] ,
         \SB2_2_23/Component_Function_2/NAND4_in[2] ,
         \SB2_2_23/Component_Function_2/NAND4_in[1] ,
         \SB2_2_23/Component_Function_2/NAND4_in[0] ,
         \SB2_2_23/Component_Function_3/NAND4_in[3] ,
         \SB2_2_23/Component_Function_3/NAND4_in[2] ,
         \SB2_2_23/Component_Function_3/NAND4_in[0] ,
         \SB2_2_23/Component_Function_4/NAND4_in[3] ,
         \SB2_2_23/Component_Function_4/NAND4_in[1] ,
         \SB2_2_23/Component_Function_4/NAND4_in[0] ,
         \SB2_2_24/Component_Function_2/NAND4_in[2] ,
         \SB2_2_24/Component_Function_2/NAND4_in[0] ,
         \SB2_2_24/Component_Function_3/NAND4_in[3] ,
         \SB2_2_24/Component_Function_3/NAND4_in[0] ,
         \SB2_2_24/Component_Function_4/NAND4_in[3] ,
         \SB2_2_24/Component_Function_4/NAND4_in[1] ,
         \SB2_2_24/Component_Function_4/NAND4_in[0] ,
         \SB2_2_25/Component_Function_2/NAND4_in[3] ,
         \SB2_2_25/Component_Function_2/NAND4_in[2] ,
         \SB2_2_25/Component_Function_2/NAND4_in[1] ,
         \SB2_2_25/Component_Function_2/NAND4_in[0] ,
         \SB2_2_25/Component_Function_3/NAND4_in[3] ,
         \SB2_2_25/Component_Function_3/NAND4_in[2] ,
         \SB2_2_25/Component_Function_3/NAND4_in[1] ,
         \SB2_2_25/Component_Function_3/NAND4_in[0] ,
         \SB2_2_25/Component_Function_4/NAND4_in[2] ,
         \SB2_2_25/Component_Function_4/NAND4_in[1] ,
         \SB2_2_25/Component_Function_4/NAND4_in[0] ,
         \SB2_2_26/Component_Function_2/NAND4_in[3] ,
         \SB2_2_26/Component_Function_2/NAND4_in[2] ,
         \SB2_2_26/Component_Function_2/NAND4_in[1] ,
         \SB2_2_26/Component_Function_2/NAND4_in[0] ,
         \SB2_2_26/Component_Function_3/NAND4_in[3] ,
         \SB2_2_26/Component_Function_3/NAND4_in[1] ,
         \SB2_2_26/Component_Function_4/NAND4_in[2] ,
         \SB2_2_26/Component_Function_4/NAND4_in[1] ,
         \SB2_2_26/Component_Function_4/NAND4_in[0] ,
         \SB2_2_27/Component_Function_2/NAND4_in[2] ,
         \SB2_2_27/Component_Function_2/NAND4_in[0] ,
         \SB2_2_27/Component_Function_3/NAND4_in[3] ,
         \SB2_2_27/Component_Function_3/NAND4_in[0] ,
         \SB2_2_27/Component_Function_4/NAND4_in[3] ,
         \SB2_2_27/Component_Function_4/NAND4_in[1] ,
         \SB2_2_28/Component_Function_2/NAND4_in[3] ,
         \SB2_2_28/Component_Function_2/NAND4_in[2] ,
         \SB2_2_28/Component_Function_2/NAND4_in[0] ,
         \SB2_2_28/Component_Function_3/NAND4_in[1] ,
         \SB2_2_28/Component_Function_3/NAND4_in[0] ,
         \SB2_2_28/Component_Function_4/NAND4_in[3] ,
         \SB2_2_28/Component_Function_4/NAND4_in[1] ,
         \SB2_2_28/Component_Function_4/NAND4_in[0] ,
         \SB2_2_29/Component_Function_2/NAND4_in[1] ,
         \SB2_2_29/Component_Function_2/NAND4_in[0] ,
         \SB2_2_29/Component_Function_3/NAND4_in[1] ,
         \SB2_2_29/Component_Function_3/NAND4_in[0] ,
         \SB2_2_29/Component_Function_4/NAND4_in[3] ,
         \SB2_2_29/Component_Function_4/NAND4_in[2] ,
         \SB2_2_29/Component_Function_4/NAND4_in[1] ,
         \SB2_2_29/Component_Function_4/NAND4_in[0] ,
         \SB2_2_30/Component_Function_2/NAND4_in[3] ,
         \SB2_2_30/Component_Function_2/NAND4_in[2] ,
         \SB2_2_30/Component_Function_2/NAND4_in[0] ,
         \SB2_2_30/Component_Function_3/NAND4_in[3] ,
         \SB2_2_30/Component_Function_3/NAND4_in[1] ,
         \SB2_2_30/Component_Function_3/NAND4_in[0] ,
         \SB2_2_30/Component_Function_4/NAND4_in[3] ,
         \SB2_2_30/Component_Function_4/NAND4_in[1] ,
         \SB2_2_30/Component_Function_4/NAND4_in[0] ,
         \SB2_2_31/Component_Function_2/NAND4_in[3] ,
         \SB2_2_31/Component_Function_2/NAND4_in[2] ,
         \SB2_2_31/Component_Function_2/NAND4_in[1] ,
         \SB2_2_31/Component_Function_2/NAND4_in[0] ,
         \SB2_2_31/Component_Function_3/NAND4_in[3] ,
         \SB2_2_31/Component_Function_3/NAND4_in[2] ,
         \SB2_2_31/Component_Function_3/NAND4_in[1] ,
         \SB2_2_31/Component_Function_3/NAND4_in[0] ,
         \SB2_2_31/Component_Function_4/NAND4_in[3] ,
         \SB2_2_31/Component_Function_4/NAND4_in[1] ,
         \SB2_2_31/Component_Function_4/NAND4_in[0] ,
         \SB1_3_0/Component_Function_2/NAND4_in[2] ,
         \SB1_3_0/Component_Function_2/NAND4_in[1] ,
         \SB1_3_0/Component_Function_2/NAND4_in[0] ,
         \SB1_3_0/Component_Function_3/NAND4_in[3] ,
         \SB1_3_0/Component_Function_3/NAND4_in[1] ,
         \SB1_3_0/Component_Function_3/NAND4_in[0] ,
         \SB1_3_0/Component_Function_4/NAND4_in[3] ,
         \SB1_3_0/Component_Function_4/NAND4_in[1] ,
         \SB1_3_0/Component_Function_4/NAND4_in[0] ,
         \SB1_3_1/Component_Function_2/NAND4_in[2] ,
         \SB1_3_1/Component_Function_2/NAND4_in[1] ,
         \SB1_3_1/Component_Function_2/NAND4_in[0] ,
         \SB1_3_1/Component_Function_3/NAND4_in[1] ,
         \SB1_3_1/Component_Function_3/NAND4_in[0] ,
         \SB1_3_1/Component_Function_4/NAND4_in[3] ,
         \SB1_3_1/Component_Function_4/NAND4_in[0] ,
         \SB1_3_2/Component_Function_2/NAND4_in[3] ,
         \SB1_3_2/Component_Function_2/NAND4_in[2] ,
         \SB1_3_2/Component_Function_2/NAND4_in[0] ,
         \SB1_3_2/Component_Function_3/NAND4_in[1] ,
         \SB1_3_2/Component_Function_3/NAND4_in[0] ,
         \SB1_3_2/Component_Function_4/NAND4_in[3] ,
         \SB1_3_2/Component_Function_4/NAND4_in[2] ,
         \SB1_3_2/Component_Function_4/NAND4_in[1] ,
         \SB1_3_2/Component_Function_4/NAND4_in[0] ,
         \SB1_3_3/Component_Function_2/NAND4_in[3] ,
         \SB1_3_3/Component_Function_2/NAND4_in[1] ,
         \SB1_3_3/Component_Function_2/NAND4_in[0] ,
         \SB1_3_3/Component_Function_3/NAND4_in[1] ,
         \SB1_3_3/Component_Function_4/NAND4_in[3] ,
         \SB1_3_3/Component_Function_4/NAND4_in[2] ,
         \SB1_3_3/Component_Function_4/NAND4_in[1] ,
         \SB1_3_3/Component_Function_4/NAND4_in[0] ,
         \SB1_3_4/Component_Function_2/NAND4_in[2] ,
         \SB1_3_4/Component_Function_2/NAND4_in[1] ,
         \SB1_3_4/Component_Function_3/NAND4_in[1] ,
         \SB1_3_4/Component_Function_4/NAND4_in[0] ,
         \SB1_3_5/Component_Function_2/NAND4_in[0] ,
         \SB1_3_5/Component_Function_3/NAND4_in[2] ,
         \SB1_3_5/Component_Function_3/NAND4_in[1] ,
         \SB1_3_5/Component_Function_3/NAND4_in[0] ,
         \SB1_3_5/Component_Function_4/NAND4_in[3] ,
         \SB1_3_5/Component_Function_4/NAND4_in[2] ,
         \SB1_3_5/Component_Function_4/NAND4_in[1] ,
         \SB1_3_5/Component_Function_4/NAND4_in[0] ,
         \SB1_3_6/Component_Function_2/NAND4_in[2] ,
         \SB1_3_6/Component_Function_2/NAND4_in[1] ,
         \SB1_3_6/Component_Function_2/NAND4_in[0] ,
         \SB1_3_6/Component_Function_3/NAND4_in[1] ,
         \SB1_3_6/Component_Function_3/NAND4_in[0] ,
         \SB1_3_6/Component_Function_4/NAND4_in[3] ,
         \SB1_3_6/Component_Function_4/NAND4_in[2] ,
         \SB1_3_6/Component_Function_4/NAND4_in[1] ,
         \SB1_3_6/Component_Function_4/NAND4_in[0] ,
         \SB1_3_7/Component_Function_2/NAND4_in[1] ,
         \SB1_3_7/Component_Function_2/NAND4_in[0] ,
         \SB1_3_7/Component_Function_3/NAND4_in[3] ,
         \SB1_3_7/Component_Function_3/NAND4_in[1] ,
         \SB1_3_7/Component_Function_4/NAND4_in[3] ,
         \SB1_3_7/Component_Function_4/NAND4_in[2] ,
         \SB1_3_7/Component_Function_4/NAND4_in[1] ,
         \SB1_3_7/Component_Function_4/NAND4_in[0] ,
         \SB1_3_8/Component_Function_2/NAND4_in[3] ,
         \SB1_3_8/Component_Function_2/NAND4_in[2] ,
         \SB1_3_8/Component_Function_2/NAND4_in[1] ,
         \SB1_3_8/Component_Function_2/NAND4_in[0] ,
         \SB1_3_8/Component_Function_3/NAND4_in[2] ,
         \SB1_3_8/Component_Function_3/NAND4_in[1] ,
         \SB1_3_8/Component_Function_3/NAND4_in[0] ,
         \SB1_3_8/Component_Function_4/NAND4_in[0] ,
         \SB1_3_9/Component_Function_2/NAND4_in[3] ,
         \SB1_3_9/Component_Function_2/NAND4_in[1] ,
         \SB1_3_9/Component_Function_3/NAND4_in[1] ,
         \SB1_3_9/Component_Function_3/NAND4_in[0] ,
         \SB1_3_9/Component_Function_4/NAND4_in[3] ,
         \SB1_3_9/Component_Function_4/NAND4_in[1] ,
         \SB1_3_10/Component_Function_2/NAND4_in[3] ,
         \SB1_3_10/Component_Function_2/NAND4_in[1] ,
         \SB1_3_10/Component_Function_3/NAND4_in[3] ,
         \SB1_3_10/Component_Function_3/NAND4_in[0] ,
         \SB1_3_10/Component_Function_4/NAND4_in[3] ,
         \SB1_3_10/Component_Function_4/NAND4_in[2] ,
         \SB1_3_10/Component_Function_4/NAND4_in[1] ,
         \SB1_3_10/Component_Function_4/NAND4_in[0] ,
         \SB1_3_11/Component_Function_2/NAND4_in[2] ,
         \SB1_3_11/Component_Function_2/NAND4_in[1] ,
         \SB1_3_11/Component_Function_2/NAND4_in[0] ,
         \SB1_3_11/Component_Function_3/NAND4_in[2] ,
         \SB1_3_11/Component_Function_3/NAND4_in[1] ,
         \SB1_3_11/Component_Function_3/NAND4_in[0] ,
         \SB1_3_11/Component_Function_4/NAND4_in[3] ,
         \SB1_3_11/Component_Function_4/NAND4_in[1] ,
         \SB1_3_11/Component_Function_4/NAND4_in[0] ,
         \SB1_3_12/Component_Function_2/NAND4_in[2] ,
         \SB1_3_12/Component_Function_2/NAND4_in[1] ,
         \SB1_3_12/Component_Function_2/NAND4_in[0] ,
         \SB1_3_12/Component_Function_3/NAND4_in[3] ,
         \SB1_3_12/Component_Function_3/NAND4_in[2] ,
         \SB1_3_12/Component_Function_4/NAND4_in[1] ,
         \SB1_3_13/Component_Function_2/NAND4_in[3] ,
         \SB1_3_13/Component_Function_2/NAND4_in[2] ,
         \SB1_3_13/Component_Function_2/NAND4_in[1] ,
         \SB1_3_13/Component_Function_2/NAND4_in[0] ,
         \SB1_3_13/Component_Function_3/NAND4_in[2] ,
         \SB1_3_13/Component_Function_3/NAND4_in[0] ,
         \SB1_3_13/Component_Function_4/NAND4_in[3] ,
         \SB1_3_13/Component_Function_4/NAND4_in[1] ,
         \SB1_3_13/Component_Function_4/NAND4_in[0] ,
         \SB1_3_14/Component_Function_2/NAND4_in[2] ,
         \SB1_3_14/Component_Function_2/NAND4_in[1] ,
         \SB1_3_14/Component_Function_3/NAND4_in[1] ,
         \SB1_3_14/Component_Function_3/NAND4_in[0] ,
         \SB1_3_14/Component_Function_4/NAND4_in[3] ,
         \SB1_3_14/Component_Function_4/NAND4_in[2] ,
         \SB1_3_15/Component_Function_2/NAND4_in[3] ,
         \SB1_3_15/Component_Function_2/NAND4_in[1] ,
         \SB1_3_15/Component_Function_2/NAND4_in[0] ,
         \SB1_3_15/Component_Function_3/NAND4_in[1] ,
         \SB1_3_15/Component_Function_3/NAND4_in[0] ,
         \SB1_3_15/Component_Function_4/NAND4_in[3] ,
         \SB1_3_15/Component_Function_4/NAND4_in[1] ,
         \SB1_3_15/Component_Function_4/NAND4_in[0] ,
         \SB1_3_16/Component_Function_2/NAND4_in[1] ,
         \SB1_3_16/Component_Function_2/NAND4_in[0] ,
         \SB1_3_16/Component_Function_3/NAND4_in[3] ,
         \SB1_3_16/Component_Function_3/NAND4_in[1] ,
         \SB1_3_16/Component_Function_4/NAND4_in[3] ,
         \SB1_3_17/Component_Function_2/NAND4_in[2] ,
         \SB1_3_17/Component_Function_2/NAND4_in[0] ,
         \SB1_3_17/Component_Function_3/NAND4_in[3] ,
         \SB1_3_17/Component_Function_3/NAND4_in[1] ,
         \SB1_3_17/Component_Function_3/NAND4_in[0] ,
         \SB1_3_17/Component_Function_4/NAND4_in[1] ,
         \SB1_3_18/Component_Function_2/NAND4_in[2] ,
         \SB1_3_18/Component_Function_2/NAND4_in[1] ,
         \SB1_3_18/Component_Function_2/NAND4_in[0] ,
         \SB1_3_18/Component_Function_3/NAND4_in[2] ,
         \SB1_3_18/Component_Function_3/NAND4_in[1] ,
         \SB1_3_18/Component_Function_4/NAND4_in[3] ,
         \SB1_3_18/Component_Function_4/NAND4_in[2] ,
         \SB1_3_18/Component_Function_4/NAND4_in[1] ,
         \SB1_3_18/Component_Function_4/NAND4_in[0] ,
         \SB1_3_19/Component_Function_2/NAND4_in[2] ,
         \SB1_3_19/Component_Function_2/NAND4_in[1] ,
         \SB1_3_19/Component_Function_2/NAND4_in[0] ,
         \SB1_3_19/Component_Function_3/NAND4_in[1] ,
         \SB1_3_19/Component_Function_4/NAND4_in[3] ,
         \SB1_3_19/Component_Function_4/NAND4_in[2] ,
         \SB1_3_19/Component_Function_4/NAND4_in[1] ,
         \SB1_3_19/Component_Function_4/NAND4_in[0] ,
         \SB1_3_20/Component_Function_2/NAND4_in[3] ,
         \SB1_3_20/Component_Function_2/NAND4_in[2] ,
         \SB1_3_20/Component_Function_2/NAND4_in[1] ,
         \SB1_3_20/Component_Function_2/NAND4_in[0] ,
         \SB1_3_20/Component_Function_3/NAND4_in[2] ,
         \SB1_3_20/Component_Function_3/NAND4_in[1] ,
         \SB1_3_20/Component_Function_3/NAND4_in[0] ,
         \SB1_3_20/Component_Function_4/NAND4_in[3] ,
         \SB1_3_20/Component_Function_4/NAND4_in[1] ,
         \SB1_3_20/Component_Function_4/NAND4_in[0] ,
         \SB1_3_21/Component_Function_2/NAND4_in[2] ,
         \SB1_3_21/Component_Function_2/NAND4_in[1] ,
         \SB1_3_21/Component_Function_3/NAND4_in[0] ,
         \SB1_3_22/Component_Function_2/NAND4_in[2] ,
         \SB1_3_22/Component_Function_2/NAND4_in[0] ,
         \SB1_3_22/Component_Function_3/NAND4_in[2] ,
         \SB1_3_22/Component_Function_3/NAND4_in[1] ,
         \SB1_3_22/Component_Function_3/NAND4_in[0] ,
         \SB1_3_22/Component_Function_4/NAND4_in[3] ,
         \SB1_3_23/Component_Function_2/NAND4_in[1] ,
         \SB1_3_23/Component_Function_2/NAND4_in[0] ,
         \SB1_3_23/Component_Function_3/NAND4_in[2] ,
         \SB1_3_23/Component_Function_3/NAND4_in[1] ,
         \SB1_3_23/Component_Function_3/NAND4_in[0] ,
         \SB1_3_23/Component_Function_4/NAND4_in[3] ,
         \SB1_3_23/Component_Function_4/NAND4_in[0] ,
         \SB1_3_24/Component_Function_2/NAND4_in[2] ,
         \SB1_3_24/Component_Function_2/NAND4_in[1] ,
         \SB1_3_24/Component_Function_3/NAND4_in[3] ,
         \SB1_3_24/Component_Function_3/NAND4_in[2] ,
         \SB1_3_24/Component_Function_3/NAND4_in[0] ,
         \SB1_3_24/Component_Function_4/NAND4_in[2] ,
         \SB1_3_24/Component_Function_4/NAND4_in[1] ,
         \SB1_3_24/Component_Function_4/NAND4_in[0] ,
         \SB1_3_25/Component_Function_2/NAND4_in[2] ,
         \SB1_3_25/Component_Function_2/NAND4_in[1] ,
         \SB1_3_25/Component_Function_3/NAND4_in[2] ,
         \SB1_3_25/Component_Function_3/NAND4_in[1] ,
         \SB1_3_25/Component_Function_3/NAND4_in[0] ,
         \SB1_3_25/Component_Function_4/NAND4_in[3] ,
         \SB1_3_25/Component_Function_4/NAND4_in[2] ,
         \SB1_3_25/Component_Function_4/NAND4_in[0] ,
         \SB1_3_26/Component_Function_2/NAND4_in[1] ,
         \SB1_3_26/Component_Function_3/NAND4_in[1] ,
         \SB1_3_26/Component_Function_3/NAND4_in[0] ,
         \SB1_3_26/Component_Function_4/NAND4_in[3] ,
         \SB1_3_26/Component_Function_4/NAND4_in[2] ,
         \SB1_3_26/Component_Function_4/NAND4_in[0] ,
         \SB1_3_27/Component_Function_2/NAND4_in[1] ,
         \SB1_3_27/Component_Function_2/NAND4_in[0] ,
         \SB1_3_27/Component_Function_3/NAND4_in[1] ,
         \SB1_3_27/Component_Function_4/NAND4_in[3] ,
         \SB1_3_27/Component_Function_4/NAND4_in[2] ,
         \SB1_3_27/Component_Function_4/NAND4_in[1] ,
         \SB1_3_28/Component_Function_2/NAND4_in[1] ,
         \SB1_3_28/Component_Function_2/NAND4_in[0] ,
         \SB1_3_28/Component_Function_3/NAND4_in[3] ,
         \SB1_3_28/Component_Function_3/NAND4_in[1] ,
         \SB1_3_28/Component_Function_3/NAND4_in[0] ,
         \SB1_3_28/Component_Function_4/NAND4_in[3] ,
         \SB1_3_28/Component_Function_4/NAND4_in[1] ,
         \SB1_3_28/Component_Function_4/NAND4_in[0] ,
         \SB1_3_29/Component_Function_2/NAND4_in[2] ,
         \SB1_3_29/Component_Function_2/NAND4_in[0] ,
         \SB1_3_29/Component_Function_3/NAND4_in[3] ,
         \SB1_3_29/Component_Function_3/NAND4_in[2] ,
         \SB1_3_29/Component_Function_3/NAND4_in[1] ,
         \SB1_3_29/Component_Function_3/NAND4_in[0] ,
         \SB1_3_29/Component_Function_4/NAND4_in[1] ,
         \SB1_3_29/Component_Function_4/NAND4_in[0] ,
         \SB1_3_30/Component_Function_2/NAND4_in[0] ,
         \SB1_3_30/Component_Function_3/NAND4_in[1] ,
         \SB1_3_30/Component_Function_4/NAND4_in[3] ,
         \SB1_3_30/Component_Function_4/NAND4_in[2] ,
         \SB1_3_30/Component_Function_4/NAND4_in[1] ,
         \SB1_3_30/Component_Function_4/NAND4_in[0] ,
         \SB1_3_31/Component_Function_2/NAND4_in[2] ,
         \SB1_3_31/Component_Function_2/NAND4_in[1] ,
         \SB1_3_31/Component_Function_2/NAND4_in[0] ,
         \SB1_3_31/Component_Function_3/NAND4_in[0] ,
         \SB1_3_31/Component_Function_4/NAND4_in[3] ,
         \SB1_3_31/Component_Function_4/NAND4_in[1] ,
         \SB1_3_31/Component_Function_4/NAND4_in[0] ,
         \SB2_3_0/Component_Function_2/NAND4_in[2] ,
         \SB2_3_0/Component_Function_3/NAND4_in[3] ,
         \SB2_3_0/Component_Function_3/NAND4_in[1] ,
         \SB2_3_0/Component_Function_3/NAND4_in[0] ,
         \SB2_3_0/Component_Function_4/NAND4_in[3] ,
         \SB2_3_0/Component_Function_4/NAND4_in[1] ,
         \SB2_3_0/Component_Function_4/NAND4_in[0] ,
         \SB2_3_1/Component_Function_2/NAND4_in[3] ,
         \SB2_3_1/Component_Function_2/NAND4_in[0] ,
         \SB2_3_1/Component_Function_3/NAND4_in[1] ,
         \SB2_3_1/Component_Function_3/NAND4_in[0] ,
         \SB2_3_1/Component_Function_4/NAND4_in[3] ,
         \SB2_3_1/Component_Function_4/NAND4_in[2] ,
         \SB2_3_1/Component_Function_4/NAND4_in[1] ,
         \SB2_3_1/Component_Function_4/NAND4_in[0] ,
         \SB2_3_2/Component_Function_2/NAND4_in[3] ,
         \SB2_3_2/Component_Function_2/NAND4_in[1] ,
         \SB2_3_2/Component_Function_2/NAND4_in[0] ,
         \SB2_3_2/Component_Function_3/NAND4_in[2] ,
         \SB2_3_2/Component_Function_3/NAND4_in[0] ,
         \SB2_3_2/Component_Function_4/NAND4_in[3] ,
         \SB2_3_2/Component_Function_4/NAND4_in[0] ,
         \SB2_3_3/Component_Function_2/NAND4_in[3] ,
         \SB2_3_3/Component_Function_2/NAND4_in[1] ,
         \SB2_3_3/Component_Function_2/NAND4_in[0] ,
         \SB2_3_3/Component_Function_3/NAND4_in[3] ,
         \SB2_3_3/Component_Function_3/NAND4_in[2] ,
         \SB2_3_3/Component_Function_3/NAND4_in[1] ,
         \SB2_3_3/Component_Function_3/NAND4_in[0] ,
         \SB2_3_3/Component_Function_4/NAND4_in[2] ,
         \SB2_3_3/Component_Function_4/NAND4_in[1] ,
         \SB2_3_3/Component_Function_4/NAND4_in[0] ,
         \SB2_3_4/Component_Function_2/NAND4_in[1] ,
         \SB2_3_4/Component_Function_3/NAND4_in[3] ,
         \SB2_3_4/Component_Function_3/NAND4_in[2] ,
         \SB2_3_4/Component_Function_4/NAND4_in[3] ,
         \SB2_3_4/Component_Function_4/NAND4_in[1] ,
         \SB2_3_4/Component_Function_4/NAND4_in[0] ,
         \SB2_3_5/Component_Function_2/NAND4_in[2] ,
         \SB2_3_5/Component_Function_2/NAND4_in[1] ,
         \SB2_3_5/Component_Function_2/NAND4_in[0] ,
         \SB2_3_5/Component_Function_3/NAND4_in[3] ,
         \SB2_3_5/Component_Function_3/NAND4_in[2] ,
         \SB2_3_5/Component_Function_3/NAND4_in[1] ,
         \SB2_3_5/Component_Function_3/NAND4_in[0] ,
         \SB2_3_5/Component_Function_4/NAND4_in[3] ,
         \SB2_3_5/Component_Function_4/NAND4_in[1] ,
         \SB2_3_5/Component_Function_4/NAND4_in[0] ,
         \SB2_3_6/Component_Function_2/NAND4_in[2] ,
         \SB2_3_6/Component_Function_2/NAND4_in[1] ,
         \SB2_3_6/Component_Function_2/NAND4_in[0] ,
         \SB2_3_6/Component_Function_3/NAND4_in[3] ,
         \SB2_3_6/Component_Function_3/NAND4_in[0] ,
         \SB2_3_6/Component_Function_4/NAND4_in[3] ,
         \SB2_3_6/Component_Function_4/NAND4_in[2] ,
         \SB2_3_7/Component_Function_2/NAND4_in[0] ,
         \SB2_3_7/Component_Function_3/NAND4_in[3] ,
         \SB2_3_7/Component_Function_3/NAND4_in[2] ,
         \SB2_3_7/Component_Function_4/NAND4_in[3] ,
         \SB2_3_7/Component_Function_4/NAND4_in[1] ,
         \SB2_3_7/Component_Function_4/NAND4_in[0] ,
         \SB2_3_8/Component_Function_2/NAND4_in[2] ,
         \SB2_3_8/Component_Function_2/NAND4_in[1] ,
         \SB2_3_8/Component_Function_3/NAND4_in[1] ,
         \SB2_3_8/Component_Function_3/NAND4_in[0] ,
         \SB2_3_8/Component_Function_4/NAND4_in[3] ,
         \SB2_3_8/Component_Function_4/NAND4_in[0] ,
         \SB2_3_9/Component_Function_2/NAND4_in[2] ,
         \SB2_3_9/Component_Function_2/NAND4_in[0] ,
         \SB2_3_9/Component_Function_3/NAND4_in[3] ,
         \SB2_3_9/Component_Function_3/NAND4_in[2] ,
         \SB2_3_9/Component_Function_3/NAND4_in[1] ,
         \SB2_3_9/Component_Function_3/NAND4_in[0] ,
         \SB2_3_9/Component_Function_4/NAND4_in[2] ,
         \SB2_3_9/Component_Function_4/NAND4_in[1] ,
         \SB2_3_9/Component_Function_4/NAND4_in[0] ,
         \SB2_3_10/Component_Function_2/NAND4_in[2] ,
         \SB2_3_10/Component_Function_2/NAND4_in[1] ,
         \SB2_3_10/Component_Function_3/NAND4_in[3] ,
         \SB2_3_10/Component_Function_3/NAND4_in[2] ,
         \SB2_3_10/Component_Function_3/NAND4_in[0] ,
         \SB2_3_10/Component_Function_4/NAND4_in[3] ,
         \SB2_3_10/Component_Function_4/NAND4_in[1] ,
         \SB2_3_10/Component_Function_4/NAND4_in[0] ,
         \SB2_3_11/Component_Function_2/NAND4_in[3] ,
         \SB2_3_11/Component_Function_2/NAND4_in[1] ,
         \SB2_3_11/Component_Function_2/NAND4_in[0] ,
         \SB2_3_11/Component_Function_3/NAND4_in[3] ,
         \SB2_3_11/Component_Function_3/NAND4_in[1] ,
         \SB2_3_11/Component_Function_3/NAND4_in[0] ,
         \SB2_3_11/Component_Function_4/NAND4_in[3] ,
         \SB2_3_11/Component_Function_4/NAND4_in[1] ,
         \SB2_3_11/Component_Function_4/NAND4_in[0] ,
         \SB2_3_12/Component_Function_2/NAND4_in[2] ,
         \SB2_3_12/Component_Function_2/NAND4_in[0] ,
         \SB2_3_12/Component_Function_3/NAND4_in[3] ,
         \SB2_3_12/Component_Function_3/NAND4_in[2] ,
         \SB2_3_12/Component_Function_3/NAND4_in[1] ,
         \SB2_3_12/Component_Function_3/NAND4_in[0] ,
         \SB2_3_12/Component_Function_4/NAND4_in[3] ,
         \SB2_3_12/Component_Function_4/NAND4_in[1] ,
         \SB2_3_12/Component_Function_4/NAND4_in[0] ,
         \SB2_3_13/Component_Function_2/NAND4_in[3] ,
         \SB2_3_13/Component_Function_2/NAND4_in[2] ,
         \SB2_3_13/Component_Function_2/NAND4_in[0] ,
         \SB2_3_13/Component_Function_3/NAND4_in[3] ,
         \SB2_3_13/Component_Function_3/NAND4_in[2] ,
         \SB2_3_13/Component_Function_3/NAND4_in[1] ,
         \SB2_3_13/Component_Function_3/NAND4_in[0] ,
         \SB2_3_13/Component_Function_4/NAND4_in[2] ,
         \SB2_3_13/Component_Function_4/NAND4_in[1] ,
         \SB2_3_13/Component_Function_4/NAND4_in[0] ,
         \SB2_3_14/Component_Function_2/NAND4_in[2] ,
         \SB2_3_14/Component_Function_2/NAND4_in[1] ,
         \SB2_3_14/Component_Function_2/NAND4_in[0] ,
         \SB2_3_14/Component_Function_3/NAND4_in[3] ,
         \SB2_3_14/Component_Function_3/NAND4_in[1] ,
         \SB2_3_14/Component_Function_3/NAND4_in[0] ,
         \SB2_3_14/Component_Function_4/NAND4_in[2] ,
         \SB2_3_14/Component_Function_4/NAND4_in[1] ,
         \SB2_3_14/Component_Function_4/NAND4_in[0] ,
         \SB2_3_15/Component_Function_2/NAND4_in[3] ,
         \SB2_3_15/Component_Function_2/NAND4_in[1] ,
         \SB2_3_15/Component_Function_2/NAND4_in[0] ,
         \SB2_3_15/Component_Function_3/NAND4_in[3] ,
         \SB2_3_15/Component_Function_3/NAND4_in[1] ,
         \SB2_3_15/Component_Function_3/NAND4_in[0] ,
         \SB2_3_15/Component_Function_4/NAND4_in[3] ,
         \SB2_3_15/Component_Function_4/NAND4_in[1] ,
         \SB2_3_15/Component_Function_4/NAND4_in[0] ,
         \SB2_3_16/Component_Function_2/NAND4_in[3] ,
         \SB2_3_16/Component_Function_2/NAND4_in[2] ,
         \SB2_3_16/Component_Function_2/NAND4_in[1] ,
         \SB2_3_16/Component_Function_2/NAND4_in[0] ,
         \SB2_3_16/Component_Function_3/NAND4_in[3] ,
         \SB2_3_16/Component_Function_3/NAND4_in[2] ,
         \SB2_3_16/Component_Function_3/NAND4_in[1] ,
         \SB2_3_16/Component_Function_3/NAND4_in[0] ,
         \SB2_3_16/Component_Function_4/NAND4_in[3] ,
         \SB2_3_16/Component_Function_4/NAND4_in[2] ,
         \SB2_3_16/Component_Function_4/NAND4_in[1] ,
         \SB2_3_16/Component_Function_4/NAND4_in[0] ,
         \SB2_3_17/Component_Function_2/NAND4_in[3] ,
         \SB2_3_17/Component_Function_2/NAND4_in[2] ,
         \SB2_3_17/Component_Function_2/NAND4_in[1] ,
         \SB2_3_17/Component_Function_3/NAND4_in[3] ,
         \SB2_3_17/Component_Function_3/NAND4_in[1] ,
         \SB2_3_17/Component_Function_3/NAND4_in[0] ,
         \SB2_3_17/Component_Function_4/NAND4_in[3] ,
         \SB2_3_17/Component_Function_4/NAND4_in[1] ,
         \SB2_3_17/Component_Function_4/NAND4_in[0] ,
         \SB2_3_18/Component_Function_2/NAND4_in[1] ,
         \SB2_3_18/Component_Function_2/NAND4_in[0] ,
         \SB2_3_18/Component_Function_3/NAND4_in[2] ,
         \SB2_3_18/Component_Function_3/NAND4_in[0] ,
         \SB2_3_18/Component_Function_4/NAND4_in[2] ,
         \SB2_3_18/Component_Function_4/NAND4_in[1] ,
         \SB2_3_18/Component_Function_4/NAND4_in[0] ,
         \SB2_3_19/Component_Function_2/NAND4_in[2] ,
         \SB2_3_19/Component_Function_2/NAND4_in[0] ,
         \SB2_3_19/Component_Function_3/NAND4_in[3] ,
         \SB2_3_19/Component_Function_3/NAND4_in[2] ,
         \SB2_3_19/Component_Function_3/NAND4_in[1] ,
         \SB2_3_19/Component_Function_3/NAND4_in[0] ,
         \SB2_3_19/Component_Function_4/NAND4_in[3] ,
         \SB2_3_19/Component_Function_4/NAND4_in[1] ,
         \SB2_3_19/Component_Function_4/NAND4_in[0] ,
         \SB2_3_20/Component_Function_2/NAND4_in[2] ,
         \SB2_3_20/Component_Function_2/NAND4_in[1] ,
         \SB2_3_20/Component_Function_2/NAND4_in[0] ,
         \SB2_3_20/Component_Function_3/NAND4_in[3] ,
         \SB2_3_20/Component_Function_3/NAND4_in[1] ,
         \SB2_3_20/Component_Function_3/NAND4_in[0] ,
         \SB2_3_20/Component_Function_4/NAND4_in[3] ,
         \SB2_3_20/Component_Function_4/NAND4_in[1] ,
         \SB2_3_20/Component_Function_4/NAND4_in[0] ,
         \SB2_3_21/Component_Function_2/NAND4_in[0] ,
         \SB2_3_21/Component_Function_3/NAND4_in[3] ,
         \SB2_3_21/Component_Function_3/NAND4_in[0] ,
         \SB2_3_21/Component_Function_4/NAND4_in[2] ,
         \SB2_3_21/Component_Function_4/NAND4_in[1] ,
         \SB2_3_21/Component_Function_4/NAND4_in[0] ,
         \SB2_3_22/Component_Function_2/NAND4_in[2] ,
         \SB2_3_22/Component_Function_2/NAND4_in[0] ,
         \SB2_3_22/Component_Function_3/NAND4_in[3] ,
         \SB2_3_22/Component_Function_3/NAND4_in[2] ,
         \SB2_3_22/Component_Function_3/NAND4_in[1] ,
         \SB2_3_22/Component_Function_3/NAND4_in[0] ,
         \SB2_3_22/Component_Function_4/NAND4_in[3] ,
         \SB2_3_22/Component_Function_4/NAND4_in[1] ,
         \SB2_3_22/Component_Function_4/NAND4_in[0] ,
         \SB2_3_23/Component_Function_2/NAND4_in[0] ,
         \SB2_3_23/Component_Function_3/NAND4_in[3] ,
         \SB2_3_23/Component_Function_3/NAND4_in[2] ,
         \SB2_3_23/Component_Function_3/NAND4_in[1] ,
         \SB2_3_23/Component_Function_3/NAND4_in[0] ,
         \SB2_3_23/Component_Function_4/NAND4_in[2] ,
         \SB2_3_23/Component_Function_4/NAND4_in[1] ,
         \SB2_3_23/Component_Function_4/NAND4_in[0] ,
         \SB2_3_24/Component_Function_2/NAND4_in[3] ,
         \SB2_3_24/Component_Function_2/NAND4_in[1] ,
         \SB2_3_24/Component_Function_2/NAND4_in[0] ,
         \SB2_3_24/Component_Function_3/NAND4_in[1] ,
         \SB2_3_24/Component_Function_3/NAND4_in[0] ,
         \SB2_3_24/Component_Function_4/NAND4_in[3] ,
         \SB2_3_24/Component_Function_4/NAND4_in[1] ,
         \SB2_3_24/Component_Function_4/NAND4_in[0] ,
         \SB2_3_25/Component_Function_2/NAND4_in[3] ,
         \SB2_3_25/Component_Function_2/NAND4_in[0] ,
         \SB2_3_25/Component_Function_3/NAND4_in[3] ,
         \SB2_3_25/Component_Function_3/NAND4_in[1] ,
         \SB2_3_25/Component_Function_3/NAND4_in[0] ,
         \SB2_3_25/Component_Function_4/NAND4_in[1] ,
         \SB2_3_25/Component_Function_4/NAND4_in[0] ,
         \SB2_3_26/Component_Function_2/NAND4_in[1] ,
         \SB2_3_26/Component_Function_2/NAND4_in[0] ,
         \SB2_3_26/Component_Function_3/NAND4_in[3] ,
         \SB2_3_26/Component_Function_3/NAND4_in[2] ,
         \SB2_3_26/Component_Function_3/NAND4_in[1] ,
         \SB2_3_26/Component_Function_3/NAND4_in[0] ,
         \SB2_3_26/Component_Function_4/NAND4_in[3] ,
         \SB2_3_26/Component_Function_4/NAND4_in[1] ,
         \SB2_3_26/Component_Function_4/NAND4_in[0] ,
         \SB2_3_27/Component_Function_2/NAND4_in[2] ,
         \SB2_3_27/Component_Function_2/NAND4_in[0] ,
         \SB2_3_27/Component_Function_3/NAND4_in[3] ,
         \SB2_3_27/Component_Function_3/NAND4_in[2] ,
         \SB2_3_27/Component_Function_3/NAND4_in[1] ,
         \SB2_3_27/Component_Function_3/NAND4_in[0] ,
         \SB2_3_27/Component_Function_4/NAND4_in[3] ,
         \SB2_3_27/Component_Function_4/NAND4_in[1] ,
         \SB2_3_27/Component_Function_4/NAND4_in[0] ,
         \SB2_3_28/Component_Function_3/NAND4_in[3] ,
         \SB2_3_28/Component_Function_3/NAND4_in[2] ,
         \SB2_3_28/Component_Function_3/NAND4_in[1] ,
         \SB2_3_28/Component_Function_3/NAND4_in[0] ,
         \SB2_3_28/Component_Function_4/NAND4_in[2] ,
         \SB2_3_28/Component_Function_4/NAND4_in[1] ,
         \SB2_3_28/Component_Function_4/NAND4_in[0] ,
         \SB2_3_29/Component_Function_2/NAND4_in[3] ,
         \SB2_3_29/Component_Function_2/NAND4_in[2] ,
         \SB2_3_29/Component_Function_2/NAND4_in[0] ,
         \SB2_3_29/Component_Function_3/NAND4_in[2] ,
         \SB2_3_29/Component_Function_3/NAND4_in[1] ,
         \SB2_3_29/Component_Function_3/NAND4_in[0] ,
         \SB2_3_29/Component_Function_4/NAND4_in[2] ,
         \SB2_3_29/Component_Function_4/NAND4_in[1] ,
         \SB2_3_29/Component_Function_4/NAND4_in[0] ,
         \SB2_3_30/Component_Function_2/NAND4_in[3] ,
         \SB2_3_30/Component_Function_2/NAND4_in[2] ,
         \SB2_3_30/Component_Function_2/NAND4_in[1] ,
         \SB2_3_30/Component_Function_2/NAND4_in[0] ,
         \SB2_3_30/Component_Function_3/NAND4_in[3] ,
         \SB2_3_30/Component_Function_3/NAND4_in[1] ,
         \SB2_3_30/Component_Function_3/NAND4_in[0] ,
         \SB2_3_30/Component_Function_4/NAND4_in[2] ,
         \SB2_3_30/Component_Function_4/NAND4_in[1] ,
         \SB2_3_30/Component_Function_4/NAND4_in[0] ,
         \SB2_3_31/Component_Function_2/NAND4_in[2] ,
         \SB2_3_31/Component_Function_2/NAND4_in[1] ,
         \SB2_3_31/Component_Function_2/NAND4_in[0] ,
         \SB2_3_31/Component_Function_3/NAND4_in[3] ,
         \SB2_3_31/Component_Function_3/NAND4_in[2] ,
         \SB2_3_31/Component_Function_3/NAND4_in[0] ,
         \SB2_3_31/Component_Function_4/NAND4_in[3] ,
         \SB2_3_31/Component_Function_4/NAND4_in[2] ,
         \SB3_0/Component_Function_2/NAND4_in[3] ,
         \SB3_0/Component_Function_3/NAND4_in[1] ,
         \SB3_0/Component_Function_4/NAND4_in[3] ,
         \SB3_0/Component_Function_4/NAND4_in[2] ,
         \SB3_0/Component_Function_4/NAND4_in[1] ,
         \SB3_0/Component_Function_4/NAND4_in[0] ,
         \SB3_1/Component_Function_2/NAND4_in[2] ,
         \SB3_1/Component_Function_2/NAND4_in[1] ,
         \SB3_1/Component_Function_2/NAND4_in[0] ,
         \SB3_1/Component_Function_3/NAND4_in[1] ,
         \SB3_1/Component_Function_3/NAND4_in[0] ,
         \SB3_1/Component_Function_4/NAND4_in[3] ,
         \SB3_1/Component_Function_4/NAND4_in[2] ,
         \SB3_1/Component_Function_4/NAND4_in[1] ,
         \SB3_1/Component_Function_4/NAND4_in[0] ,
         \SB3_2/Component_Function_2/NAND4_in[1] ,
         \SB3_2/Component_Function_3/NAND4_in[2] ,
         \SB3_2/Component_Function_3/NAND4_in[1] ,
         \SB3_2/Component_Function_3/NAND4_in[0] ,
         \SB3_2/Component_Function_4/NAND4_in[3] ,
         \SB3_2/Component_Function_4/NAND4_in[0] ,
         \SB3_3/Component_Function_2/NAND4_in[2] ,
         \SB3_3/Component_Function_2/NAND4_in[0] ,
         \SB3_3/Component_Function_3/NAND4_in[0] ,
         \SB3_3/Component_Function_4/NAND4_in[3] ,
         \SB3_3/Component_Function_4/NAND4_in[1] ,
         \SB3_3/Component_Function_4/NAND4_in[0] ,
         \SB3_4/Component_Function_2/NAND4_in[3] ,
         \SB3_4/Component_Function_2/NAND4_in[1] ,
         \SB3_4/Component_Function_2/NAND4_in[0] ,
         \SB3_4/Component_Function_3/NAND4_in[1] ,
         \SB3_4/Component_Function_3/NAND4_in[0] ,
         \SB3_4/Component_Function_4/NAND4_in[3] ,
         \SB3_4/Component_Function_4/NAND4_in[2] ,
         \SB3_4/Component_Function_4/NAND4_in[1] ,
         \SB3_4/Component_Function_4/NAND4_in[0] ,
         \SB3_5/Component_Function_2/NAND4_in[3] ,
         \SB3_5/Component_Function_2/NAND4_in[2] ,
         \SB3_5/Component_Function_3/NAND4_in[3] ,
         \SB3_5/Component_Function_3/NAND4_in[2] ,
         \SB3_5/Component_Function_3/NAND4_in[1] ,
         \SB3_5/Component_Function_4/NAND4_in[3] ,
         \SB3_5/Component_Function_4/NAND4_in[1] ,
         \SB3_5/Component_Function_4/NAND4_in[0] ,
         \SB3_6/Component_Function_2/NAND4_in[3] ,
         \SB3_6/Component_Function_2/NAND4_in[2] ,
         \SB3_6/Component_Function_2/NAND4_in[1] ,
         \SB3_6/Component_Function_2/NAND4_in[0] ,
         \SB3_6/Component_Function_3/NAND4_in[2] ,
         \SB3_6/Component_Function_3/NAND4_in[1] ,
         \SB3_6/Component_Function_3/NAND4_in[0] ,
         \SB3_6/Component_Function_4/NAND4_in[0] ,
         \SB3_7/Component_Function_2/NAND4_in[3] ,
         \SB3_7/Component_Function_2/NAND4_in[1] ,
         \SB3_7/Component_Function_2/NAND4_in[0] ,
         \SB3_7/Component_Function_3/NAND4_in[1] ,
         \SB3_7/Component_Function_3/NAND4_in[0] ,
         \SB3_7/Component_Function_4/NAND4_in[3] ,
         \SB3_7/Component_Function_4/NAND4_in[1] ,
         \SB3_7/Component_Function_4/NAND4_in[0] ,
         \SB3_8/Component_Function_2/NAND4_in[3] ,
         \SB3_8/Component_Function_2/NAND4_in[2] ,
         \SB3_8/Component_Function_2/NAND4_in[1] ,
         \SB3_8/Component_Function_2/NAND4_in[0] ,
         \SB3_8/Component_Function_3/NAND4_in[2] ,
         \SB3_8/Component_Function_3/NAND4_in[1] ,
         \SB3_8/Component_Function_3/NAND4_in[0] ,
         \SB3_8/Component_Function_4/NAND4_in[3] ,
         \SB3_8/Component_Function_4/NAND4_in[1] ,
         \SB3_8/Component_Function_4/NAND4_in[0] ,
         \SB3_9/Component_Function_2/NAND4_in[2] ,
         \SB3_9/Component_Function_2/NAND4_in[1] ,
         \SB3_9/Component_Function_2/NAND4_in[0] ,
         \SB3_9/Component_Function_3/NAND4_in[2] ,
         \SB3_9/Component_Function_3/NAND4_in[1] ,
         \SB3_9/Component_Function_3/NAND4_in[0] ,
         \SB3_9/Component_Function_4/NAND4_in[3] ,
         \SB3_9/Component_Function_4/NAND4_in[2] ,
         \SB3_9/Component_Function_4/NAND4_in[1] ,
         \SB3_9/Component_Function_4/NAND4_in[0] ,
         \SB3_10/Component_Function_2/NAND4_in[3] ,
         \SB3_10/Component_Function_2/NAND4_in[1] ,
         \SB3_10/Component_Function_2/NAND4_in[0] ,
         \SB3_10/Component_Function_3/NAND4_in[1] ,
         \SB3_10/Component_Function_4/NAND4_in[3] ,
         \SB3_10/Component_Function_4/NAND4_in[2] ,
         \SB3_10/Component_Function_4/NAND4_in[1] ,
         \SB3_10/Component_Function_4/NAND4_in[0] ,
         \SB3_11/Component_Function_2/NAND4_in[2] ,
         \SB3_11/Component_Function_2/NAND4_in[1] ,
         \SB3_11/Component_Function_3/NAND4_in[3] ,
         \SB3_11/Component_Function_3/NAND4_in[1] ,
         \SB3_11/Component_Function_3/NAND4_in[0] ,
         \SB3_11/Component_Function_4/NAND4_in[3] ,
         \SB3_11/Component_Function_4/NAND4_in[1] ,
         \SB3_12/Component_Function_2/NAND4_in[2] ,
         \SB3_12/Component_Function_2/NAND4_in[1] ,
         \SB3_12/Component_Function_2/NAND4_in[0] ,
         \SB3_12/Component_Function_3/NAND4_in[2] ,
         \SB3_12/Component_Function_3/NAND4_in[0] ,
         \SB3_12/Component_Function_4/NAND4_in[2] ,
         \SB3_12/Component_Function_4/NAND4_in[0] ,
         \SB3_13/Component_Function_2/NAND4_in[3] ,
         \SB3_13/Component_Function_2/NAND4_in[1] ,
         \SB3_13/Component_Function_2/NAND4_in[0] ,
         \SB3_13/Component_Function_3/NAND4_in[0] ,
         \SB3_13/Component_Function_4/NAND4_in[2] ,
         \SB3_13/Component_Function_4/NAND4_in[1] ,
         \SB3_14/Component_Function_2/NAND4_in[3] ,
         \SB3_14/Component_Function_2/NAND4_in[2] ,
         \SB3_14/Component_Function_2/NAND4_in[0] ,
         \SB3_14/Component_Function_3/NAND4_in[1] ,
         \SB3_14/Component_Function_3/NAND4_in[0] ,
         \SB3_14/Component_Function_4/NAND4_in[3] ,
         \SB3_14/Component_Function_4/NAND4_in[1] ,
         \SB3_15/Component_Function_2/NAND4_in[3] ,
         \SB3_15/Component_Function_2/NAND4_in[2] ,
         \SB3_15/Component_Function_2/NAND4_in[1] ,
         \SB3_15/Component_Function_2/NAND4_in[0] ,
         \SB3_15/Component_Function_3/NAND4_in[1] ,
         \SB3_15/Component_Function_3/NAND4_in[0] ,
         \SB3_15/Component_Function_4/NAND4_in[3] ,
         \SB3_15/Component_Function_4/NAND4_in[2] ,
         \SB3_15/Component_Function_4/NAND4_in[1] ,
         \SB3_15/Component_Function_4/NAND4_in[0] ,
         \SB3_16/Component_Function_2/NAND4_in[1] ,
         \SB3_16/Component_Function_3/NAND4_in[1] ,
         \SB3_16/Component_Function_3/NAND4_in[0] ,
         \SB3_16/Component_Function_4/NAND4_in[2] ,
         \SB3_16/Component_Function_4/NAND4_in[1] ,
         \SB3_16/Component_Function_4/NAND4_in[0] ,
         \SB3_17/Component_Function_2/NAND4_in[3] ,
         \SB3_17/Component_Function_2/NAND4_in[2] ,
         \SB3_17/Component_Function_2/NAND4_in[0] ,
         \SB3_17/Component_Function_3/NAND4_in[0] ,
         \SB3_17/Component_Function_4/NAND4_in[2] ,
         \SB3_17/Component_Function_4/NAND4_in[1] ,
         \SB3_17/Component_Function_4/NAND4_in[0] ,
         \SB3_18/Component_Function_2/NAND4_in[2] ,
         \SB3_18/Component_Function_2/NAND4_in[0] ,
         \SB3_18/Component_Function_3/NAND4_in[1] ,
         \SB3_18/Component_Function_3/NAND4_in[0] ,
         \SB3_18/Component_Function_4/NAND4_in[3] ,
         \SB3_18/Component_Function_4/NAND4_in[2] ,
         \SB3_18/Component_Function_4/NAND4_in[1] ,
         \SB3_18/Component_Function_4/NAND4_in[0] ,
         \SB3_19/Component_Function_2/NAND4_in[2] ,
         \SB3_19/Component_Function_2/NAND4_in[0] ,
         \SB3_19/Component_Function_3/NAND4_in[0] ,
         \SB3_19/Component_Function_4/NAND4_in[2] ,
         \SB3_19/Component_Function_4/NAND4_in[1] ,
         \SB3_19/Component_Function_4/NAND4_in[0] ,
         \SB3_20/Component_Function_2/NAND4_in[3] ,
         \SB3_20/Component_Function_2/NAND4_in[0] ,
         \SB3_20/Component_Function_3/NAND4_in[1] ,
         \SB3_20/Component_Function_4/NAND4_in[2] ,
         \SB3_20/Component_Function_4/NAND4_in[1] ,
         \SB3_20/Component_Function_4/NAND4_in[0] ,
         \SB3_21/Component_Function_2/NAND4_in[0] ,
         \SB3_21/Component_Function_3/NAND4_in[1] ,
         \SB3_21/Component_Function_3/NAND4_in[0] ,
         \SB3_21/Component_Function_4/NAND4_in[3] ,
         \SB3_21/Component_Function_4/NAND4_in[1] ,
         \SB3_21/Component_Function_4/NAND4_in[0] ,
         \SB3_22/Component_Function_2/NAND4_in[2] ,
         \SB3_22/Component_Function_2/NAND4_in[1] ,
         \SB3_22/Component_Function_2/NAND4_in[0] ,
         \SB3_22/Component_Function_3/NAND4_in[2] ,
         \SB3_22/Component_Function_3/NAND4_in[1] ,
         \SB3_22/Component_Function_3/NAND4_in[0] ,
         \SB3_22/Component_Function_4/NAND4_in[3] ,
         \SB3_22/Component_Function_4/NAND4_in[2] ,
         \SB3_22/Component_Function_4/NAND4_in[1] ,
         \SB3_22/Component_Function_4/NAND4_in[0] ,
         \SB3_23/Component_Function_2/NAND4_in[1] ,
         \SB3_23/Component_Function_2/NAND4_in[0] ,
         \SB3_23/Component_Function_3/NAND4_in[2] ,
         \SB3_23/Component_Function_3/NAND4_in[1] ,
         \SB3_23/Component_Function_4/NAND4_in[2] ,
         \SB3_23/Component_Function_4/NAND4_in[1] ,
         \SB3_23/Component_Function_4/NAND4_in[0] ,
         \SB3_24/Component_Function_2/NAND4_in[3] ,
         \SB3_24/Component_Function_2/NAND4_in[1] ,
         \SB3_24/Component_Function_3/NAND4_in[1] ,
         \SB3_24/Component_Function_4/NAND4_in[2] ,
         \SB3_24/Component_Function_4/NAND4_in[1] ,
         \SB3_25/Component_Function_2/NAND4_in[2] ,
         \SB3_25/Component_Function_2/NAND4_in[0] ,
         \SB3_25/Component_Function_3/NAND4_in[1] ,
         \SB3_25/Component_Function_4/NAND4_in[2] ,
         \SB3_25/Component_Function_4/NAND4_in[1] ,
         \SB3_25/Component_Function_4/NAND4_in[0] ,
         \SB3_26/Component_Function_2/NAND4_in[2] ,
         \SB3_26/Component_Function_2/NAND4_in[0] ,
         \SB3_26/Component_Function_3/NAND4_in[3] ,
         \SB3_26/Component_Function_3/NAND4_in[0] ,
         \SB3_26/Component_Function_4/NAND4_in[2] ,
         \SB3_26/Component_Function_4/NAND4_in[1] ,
         \SB3_26/Component_Function_4/NAND4_in[0] ,
         \SB3_27/Component_Function_2/NAND4_in[0] ,
         \SB3_27/Component_Function_3/NAND4_in[2] ,
         \SB3_27/Component_Function_3/NAND4_in[1] ,
         \SB3_27/Component_Function_4/NAND4_in[3] ,
         \SB3_27/Component_Function_4/NAND4_in[2] ,
         \SB3_27/Component_Function_4/NAND4_in[1] ,
         \SB3_27/Component_Function_4/NAND4_in[0] ,
         \SB3_28/Component_Function_2/NAND4_in[3] ,
         \SB3_28/Component_Function_2/NAND4_in[2] ,
         \SB3_28/Component_Function_2/NAND4_in[1] ,
         \SB3_28/Component_Function_2/NAND4_in[0] ,
         \SB3_28/Component_Function_3/NAND4_in[2] ,
         \SB3_28/Component_Function_3/NAND4_in[1] ,
         \SB3_28/Component_Function_3/NAND4_in[0] ,
         \SB3_28/Component_Function_4/NAND4_in[3] ,
         \SB3_28/Component_Function_4/NAND4_in[2] ,
         \SB3_28/Component_Function_4/NAND4_in[1] ,
         \SB3_28/Component_Function_4/NAND4_in[0] ,
         \SB3_29/Component_Function_2/NAND4_in[3] ,
         \SB3_29/Component_Function_2/NAND4_in[2] ,
         \SB3_29/Component_Function_2/NAND4_in[0] ,
         \SB3_29/Component_Function_3/NAND4_in[3] ,
         \SB3_29/Component_Function_3/NAND4_in[1] ,
         \SB3_29/Component_Function_3/NAND4_in[0] ,
         \SB3_29/Component_Function_4/NAND4_in[3] ,
         \SB3_29/Component_Function_4/NAND4_in[2] ,
         \SB3_29/Component_Function_4/NAND4_in[1] ,
         \SB3_29/Component_Function_4/NAND4_in[0] ,
         \SB3_30/Component_Function_2/NAND4_in[2] ,
         \SB3_30/Component_Function_2/NAND4_in[1] ,
         \SB3_30/Component_Function_2/NAND4_in[0] ,
         \SB3_30/Component_Function_3/NAND4_in[1] ,
         \SB3_30/Component_Function_4/NAND4_in[3] ,
         \SB3_30/Component_Function_4/NAND4_in[2] ,
         \SB3_30/Component_Function_4/NAND4_in[1] ,
         \SB3_31/Component_Function_2/NAND4_in[3] ,
         \SB3_31/Component_Function_2/NAND4_in[2] ,
         \SB3_31/Component_Function_2/NAND4_in[1] ,
         \SB3_31/Component_Function_2/NAND4_in[0] ,
         \SB3_31/Component_Function_3/NAND4_in[3] ,
         \SB3_31/Component_Function_3/NAND4_in[1] ,
         \SB3_31/Component_Function_3/NAND4_in[0] ,
         \SB3_31/Component_Function_4/NAND4_in[3] ,
         \SB3_31/Component_Function_4/NAND4_in[2] ,
         \SB3_31/Component_Function_4/NAND4_in[1] ,
         \SB4_0/Component_Function_3/NAND4_in[3] ,
         \SB4_0/Component_Function_3/NAND4_in[1] ,
         \SB4_0/Component_Function_4/NAND4_in[2] ,
         \SB4_0/Component_Function_4/NAND4_in[0] ,
         \SB4_1/Component_Function_3/NAND4_in[3] ,
         \SB4_1/Component_Function_4/NAND4_in[3] ,
         \SB4_2/Component_Function_2/NAND4_in[3] ,
         \SB4_2/Component_Function_2/NAND4_in[2] ,
         \SB4_2/Component_Function_3/NAND4_in[3] ,
         \SB4_2/Component_Function_3/NAND4_in[2] ,
         \SB4_2/Component_Function_3/NAND4_in[1] ,
         \SB4_2/Component_Function_3/NAND4_in[0] ,
         \SB4_2/Component_Function_4/NAND4_in[1] ,
         \SB4_2/Component_Function_4/NAND4_in[0] ,
         \SB4_3/Component_Function_2/NAND4_in[2] ,
         \SB4_3/Component_Function_2/NAND4_in[0] ,
         \SB4_3/Component_Function_3/NAND4_in[3] ,
         \SB4_3/Component_Function_3/NAND4_in[2] ,
         \SB4_3/Component_Function_4/NAND4_in[1] ,
         \SB4_3/Component_Function_4/NAND4_in[0] ,
         \SB4_4/Component_Function_2/NAND4_in[3] ,
         \SB4_4/Component_Function_3/NAND4_in[3] ,
         \SB4_4/Component_Function_3/NAND4_in[2] ,
         \SB4_4/Component_Function_4/NAND4_in[1] ,
         \SB4_4/Component_Function_4/NAND4_in[0] ,
         \SB4_5/Component_Function_2/NAND4_in[0] ,
         \SB4_5/Component_Function_3/NAND4_in[3] ,
         \SB4_5/Component_Function_4/NAND4_in[2] ,
         \SB4_5/Component_Function_4/NAND4_in[0] ,
         \SB4_6/Component_Function_2/NAND4_in[3] ,
         \SB4_6/Component_Function_2/NAND4_in[0] ,
         \SB4_6/Component_Function_3/NAND4_in[3] ,
         \SB4_6/Component_Function_3/NAND4_in[2] ,
         \SB4_6/Component_Function_3/NAND4_in[1] ,
         \SB4_6/Component_Function_4/NAND4_in[3] ,
         \SB4_6/Component_Function_4/NAND4_in[2] ,
         \SB4_6/Component_Function_4/NAND4_in[0] ,
         \SB4_7/Component_Function_2/NAND4_in[1] ,
         \SB4_7/Component_Function_2/NAND4_in[0] ,
         \SB4_7/Component_Function_3/NAND4_in[3] ,
         \SB4_7/Component_Function_3/NAND4_in[1] ,
         \SB4_7/Component_Function_4/NAND4_in[2] ,
         \SB4_8/Component_Function_2/NAND4_in[3] ,
         \SB4_8/Component_Function_2/NAND4_in[2] ,
         \SB4_8/Component_Function_2/NAND4_in[0] ,
         \SB4_8/Component_Function_3/NAND4_in[3] ,
         \SB4_8/Component_Function_3/NAND4_in[2] ,
         \SB4_8/Component_Function_4/NAND4_in[3] ,
         \SB4_9/Component_Function_3/NAND4_in[3] ,
         \SB4_9/Component_Function_4/NAND4_in[3] ,
         \SB4_10/Component_Function_2/NAND4_in[0] ,
         \SB4_10/Component_Function_3/NAND4_in[3] ,
         \SB4_10/Component_Function_3/NAND4_in[2] ,
         \SB4_10/Component_Function_4/NAND4_in[3] ,
         \SB4_10/Component_Function_4/NAND4_in[2] ,
         \SB4_10/Component_Function_4/NAND4_in[1] ,
         \SB4_10/Component_Function_4/NAND4_in[0] ,
         \SB4_11/Component_Function_2/NAND4_in[3] ,
         \SB4_11/Component_Function_2/NAND4_in[2] ,
         \SB4_11/Component_Function_3/NAND4_in[3] ,
         \SB4_11/Component_Function_3/NAND4_in[2] ,
         \SB4_11/Component_Function_3/NAND4_in[1] ,
         \SB4_11/Component_Function_3/NAND4_in[0] ,
         \SB4_11/Component_Function_4/NAND4_in[3] ,
         \SB4_12/Component_Function_2/NAND4_in[2] ,
         \SB4_12/Component_Function_2/NAND4_in[0] ,
         \SB4_12/Component_Function_3/NAND4_in[3] ,
         \SB4_12/Component_Function_4/NAND4_in[3] ,
         \SB4_12/Component_Function_4/NAND4_in[0] ,
         \SB4_13/Component_Function_2/NAND4_in[2] ,
         \SB4_13/Component_Function_2/NAND4_in[1] ,
         \SB4_13/Component_Function_2/NAND4_in[0] ,
         \SB4_13/Component_Function_3/NAND4_in[3] ,
         \SB4_13/Component_Function_3/NAND4_in[0] ,
         \SB4_13/Component_Function_4/NAND4_in[1] ,
         \SB4_13/Component_Function_4/NAND4_in[0] ,
         \SB4_14/Component_Function_2/NAND4_in[2] ,
         \SB4_14/Component_Function_2/NAND4_in[1] ,
         \SB4_14/Component_Function_3/NAND4_in[3] ,
         \SB4_14/Component_Function_4/NAND4_in[3] ,
         \SB4_14/Component_Function_4/NAND4_in[2] ,
         \SB4_14/Component_Function_4/NAND4_in[0] ,
         \SB4_15/Component_Function_2/NAND4_in[1] ,
         \SB4_15/Component_Function_2/NAND4_in[0] ,
         \SB4_15/Component_Function_3/NAND4_in[3] ,
         \SB4_15/Component_Function_4/NAND4_in[3] ,
         \SB4_16/Component_Function_2/NAND4_in[3] ,
         \SB4_16/Component_Function_2/NAND4_in[2] ,
         \SB4_16/Component_Function_2/NAND4_in[0] ,
         \SB4_16/Component_Function_3/NAND4_in[3] ,
         \SB4_16/Component_Function_3/NAND4_in[2] ,
         \SB4_16/Component_Function_4/NAND4_in[0] ,
         \SB4_17/Component_Function_2/NAND4_in[2] ,
         \SB4_17/Component_Function_2/NAND4_in[1] ,
         \SB4_17/Component_Function_3/NAND4_in[3] ,
         \SB4_17/Component_Function_3/NAND4_in[2] ,
         \SB4_17/Component_Function_4/NAND4_in[0] ,
         \SB4_18/Component_Function_2/NAND4_in[2] ,
         \SB4_18/Component_Function_3/NAND4_in[3] ,
         \SB4_18/Component_Function_3/NAND4_in[2] ,
         \SB4_18/Component_Function_3/NAND4_in[1] ,
         \SB4_18/Component_Function_4/NAND4_in[3] ,
         \SB4_19/Component_Function_2/NAND4_in[2] ,
         \SB4_19/Component_Function_2/NAND4_in[1] ,
         \SB4_19/Component_Function_2/NAND4_in[0] ,
         \SB4_19/Component_Function_3/NAND4_in[3] ,
         \SB4_19/Component_Function_3/NAND4_in[1] ,
         \SB4_19/Component_Function_4/NAND4_in[3] ,
         \SB4_19/Component_Function_4/NAND4_in[2] ,
         \SB4_19/Component_Function_4/NAND4_in[1] ,
         \SB4_19/Component_Function_4/NAND4_in[0] ,
         \SB4_20/Component_Function_2/NAND4_in[2] ,
         \SB4_20/Component_Function_2/NAND4_in[1] ,
         \SB4_20/Component_Function_2/NAND4_in[0] ,
         \SB4_20/Component_Function_3/NAND4_in[2] ,
         \SB4_20/Component_Function_3/NAND4_in[0] ,
         \SB4_20/Component_Function_4/NAND4_in[3] ,
         \SB4_20/Component_Function_4/NAND4_in[1] ,
         \SB4_20/Component_Function_4/NAND4_in[0] ,
         \SB4_21/Component_Function_2/NAND4_in[2] ,
         \SB4_21/Component_Function_3/NAND4_in[3] ,
         \SB4_21/Component_Function_3/NAND4_in[1] ,
         \SB4_21/Component_Function_4/NAND4_in[3] ,
         \SB4_21/Component_Function_4/NAND4_in[1] ,
         \SB4_22/Component_Function_2/NAND4_in[3] ,
         \SB4_22/Component_Function_2/NAND4_in[1] ,
         \SB4_22/Component_Function_3/NAND4_in[2] ,
         \SB4_22/Component_Function_3/NAND4_in[0] ,
         \SB4_22/Component_Function_4/NAND4_in[3] ,
         \SB4_22/Component_Function_4/NAND4_in[0] ,
         \SB4_23/Component_Function_2/NAND4_in[2] ,
         \SB4_23/Component_Function_2/NAND4_in[0] ,
         \SB4_23/Component_Function_3/NAND4_in[3] ,
         \SB4_23/Component_Function_3/NAND4_in[2] ,
         \SB4_23/Component_Function_3/NAND4_in[1] ,
         \SB4_23/Component_Function_3/NAND4_in[0] ,
         \SB4_23/Component_Function_4/NAND4_in[2] ,
         \SB4_24/Component_Function_2/NAND4_in[3] ,
         \SB4_24/Component_Function_2/NAND4_in[2] ,
         \SB4_24/Component_Function_2/NAND4_in[1] ,
         \SB4_24/Component_Function_2/NAND4_in[0] ,
         \SB4_24/Component_Function_3/NAND4_in[3] ,
         \SB4_24/Component_Function_3/NAND4_in[2] ,
         \SB4_24/Component_Function_3/NAND4_in[1] ,
         \SB4_24/Component_Function_3/NAND4_in[0] ,
         \SB4_24/Component_Function_4/NAND4_in[3] ,
         \SB4_24/Component_Function_4/NAND4_in[0] ,
         \SB4_25/Component_Function_2/NAND4_in[3] ,
         \SB4_25/Component_Function_2/NAND4_in[2] ,
         \SB4_25/Component_Function_2/NAND4_in[1] ,
         \SB4_25/Component_Function_3/NAND4_in[3] ,
         \SB4_25/Component_Function_3/NAND4_in[2] ,
         \SB4_25/Component_Function_3/NAND4_in[1] ,
         \SB4_25/Component_Function_4/NAND4_in[3] ,
         \SB4_25/Component_Function_4/NAND4_in[1] ,
         \SB4_25/Component_Function_4/NAND4_in[0] ,
         \SB4_26/Component_Function_2/NAND4_in[3] ,
         \SB4_26/Component_Function_2/NAND4_in[1] ,
         \SB4_26/Component_Function_2/NAND4_in[0] ,
         \SB4_26/Component_Function_3/NAND4_in[3] ,
         \SB4_26/Component_Function_3/NAND4_in[1] ,
         \SB4_26/Component_Function_4/NAND4_in[1] ,
         \SB4_27/Component_Function_2/NAND4_in[1] ,
         \SB4_27/Component_Function_2/NAND4_in[0] ,
         \SB4_27/Component_Function_3/NAND4_in[3] ,
         \SB4_27/Component_Function_3/NAND4_in[2] ,
         \SB4_27/Component_Function_3/NAND4_in[1] ,
         \SB4_27/Component_Function_3/NAND4_in[0] ,
         \SB4_27/Component_Function_4/NAND4_in[1] ,
         \SB4_28/Component_Function_2/NAND4_in[2] ,
         \SB4_28/Component_Function_2/NAND4_in[0] ,
         \SB4_28/Component_Function_3/NAND4_in[3] ,
         \SB4_28/Component_Function_3/NAND4_in[2] ,
         \SB4_29/Component_Function_2/NAND4_in[3] ,
         \SB4_29/Component_Function_2/NAND4_in[2] ,
         \SB4_29/Component_Function_2/NAND4_in[0] ,
         \SB4_29/Component_Function_3/NAND4_in[3] ,
         \SB4_29/Component_Function_4/NAND4_in[3] ,
         \SB4_29/Component_Function_4/NAND4_in[1] ,
         \SB4_29/Component_Function_4/NAND4_in[0] ,
         \SB4_30/Component_Function_2/NAND4_in[2] ,
         \SB4_30/Component_Function_2/NAND4_in[0] ,
         \SB4_30/Component_Function_3/NAND4_in[3] ,
         \SB4_30/Component_Function_3/NAND4_in[2] ,
         \SB4_30/Component_Function_4/NAND4_in[3] ,
         \SB4_30/Component_Function_4/NAND4_in[1] ,
         \SB4_31/Component_Function_2/NAND4_in[2] ,
         \SB4_31/Component_Function_3/NAND4_in[3] ,
         \SB4_31/Component_Function_3/NAND4_in[2] ,
         \SB4_31/Component_Function_3/NAND4_in[1] ,
         \SB4_31/Component_Function_4/NAND4_in[3] ,
         \SB1_0_0/Component_Function_0/NAND4_in[3] ,
         \SB1_0_0/Component_Function_0/NAND4_in[2] ,
         \SB1_0_0/Component_Function_0/NAND4_in[1] ,
         \SB1_0_0/Component_Function_0/NAND4_in[0] ,
         \SB1_0_0/Component_Function_1/NAND4_in[3] ,
         \SB1_0_0/Component_Function_1/NAND4_in[2] ,
         \SB1_0_0/Component_Function_1/NAND4_in[1] ,
         \SB1_0_0/Component_Function_1/NAND4_in[0] ,
         \SB1_0_0/Component_Function_5/NAND4_in[2] ,
         \SB1_0_0/Component_Function_5/NAND4_in[0] ,
         \SB1_0_1/Component_Function_0/NAND4_in[3] ,
         \SB1_0_1/Component_Function_0/NAND4_in[1] ,
         \SB1_0_1/Component_Function_0/NAND4_in[0] ,
         \SB1_0_1/Component_Function_1/NAND4_in[3] ,
         \SB1_0_1/Component_Function_1/NAND4_in[2] ,
         \SB1_0_1/Component_Function_1/NAND4_in[1] ,
         \SB1_0_1/Component_Function_1/NAND4_in[0] ,
         \SB1_0_1/Component_Function_5/NAND4_in[3] ,
         \SB1_0_1/Component_Function_5/NAND4_in[2] ,
         \SB1_0_1/Component_Function_5/NAND4_in[1] ,
         \SB1_0_2/Component_Function_0/NAND4_in[3] ,
         \SB1_0_2/Component_Function_0/NAND4_in[2] ,
         \SB1_0_2/Component_Function_0/NAND4_in[1] ,
         \SB1_0_2/Component_Function_0/NAND4_in[0] ,
         \SB1_0_2/Component_Function_1/NAND4_in[3] ,
         \SB1_0_2/Component_Function_1/NAND4_in[2] ,
         \SB1_0_2/Component_Function_1/NAND4_in[1] ,
         \SB1_0_2/Component_Function_5/NAND4_in[2] ,
         \SB1_0_2/Component_Function_5/NAND4_in[1] ,
         \SB1_0_3/Component_Function_0/NAND4_in[3] ,
         \SB1_0_3/Component_Function_0/NAND4_in[2] ,
         \SB1_0_3/Component_Function_0/NAND4_in[1] ,
         \SB1_0_3/Component_Function_0/NAND4_in[0] ,
         \SB1_0_3/Component_Function_1/NAND4_in[3] ,
         \SB1_0_3/Component_Function_1/NAND4_in[2] ,
         \SB1_0_3/Component_Function_1/NAND4_in[1] ,
         \SB1_0_3/Component_Function_1/NAND4_in[0] ,
         \SB1_0_3/Component_Function_5/NAND4_in[3] ,
         \SB1_0_3/Component_Function_5/NAND4_in[2] ,
         \SB1_0_3/Component_Function_5/NAND4_in[1] ,
         \SB1_0_3/Component_Function_5/NAND4_in[0] ,
         \SB1_0_4/Component_Function_0/NAND4_in[3] ,
         \SB1_0_4/Component_Function_0/NAND4_in[2] ,
         \SB1_0_4/Component_Function_0/NAND4_in[1] ,
         \SB1_0_4/Component_Function_0/NAND4_in[0] ,
         \SB1_0_4/Component_Function_1/NAND4_in[3] ,
         \SB1_0_4/Component_Function_1/NAND4_in[2] ,
         \SB1_0_4/Component_Function_1/NAND4_in[1] ,
         \SB1_0_4/Component_Function_1/NAND4_in[0] ,
         \SB1_0_4/Component_Function_5/NAND4_in[3] ,
         \SB1_0_4/Component_Function_5/NAND4_in[2] ,
         \SB1_0_4/Component_Function_5/NAND4_in[1] ,
         \SB1_0_4/Component_Function_5/NAND4_in[0] ,
         \SB1_0_5/Component_Function_0/NAND4_in[3] ,
         \SB1_0_5/Component_Function_0/NAND4_in[2] ,
         \SB1_0_5/Component_Function_0/NAND4_in[1] ,
         \SB1_0_5/Component_Function_0/NAND4_in[0] ,
         \SB1_0_5/Component_Function_1/NAND4_in[2] ,
         \SB1_0_5/Component_Function_1/NAND4_in[1] ,
         \SB1_0_5/Component_Function_5/NAND4_in[3] ,
         \SB1_0_5/Component_Function_5/NAND4_in[2] ,
         \SB1_0_5/Component_Function_5/NAND4_in[1] ,
         \SB1_0_5/Component_Function_5/NAND4_in[0] ,
         \SB1_0_6/Component_Function_0/NAND4_in[3] ,
         \SB1_0_6/Component_Function_0/NAND4_in[2] ,
         \SB1_0_6/Component_Function_0/NAND4_in[1] ,
         \SB1_0_6/Component_Function_0/NAND4_in[0] ,
         \SB1_0_6/Component_Function_1/NAND4_in[3] ,
         \SB1_0_6/Component_Function_1/NAND4_in[1] ,
         \SB1_0_6/Component_Function_1/NAND4_in[0] ,
         \SB1_0_6/Component_Function_5/NAND4_in[3] ,
         \SB1_0_6/Component_Function_5/NAND4_in[1] ,
         \SB1_0_6/Component_Function_5/NAND4_in[0] ,
         \SB1_0_7/Component_Function_0/NAND4_in[1] ,
         \SB1_0_7/Component_Function_0/NAND4_in[0] ,
         \SB1_0_7/Component_Function_1/NAND4_in[3] ,
         \SB1_0_7/Component_Function_1/NAND4_in[2] ,
         \SB1_0_7/Component_Function_1/NAND4_in[1] ,
         \SB1_0_7/Component_Function_1/NAND4_in[0] ,
         \SB1_0_7/Component_Function_5/NAND4_in[3] ,
         \SB1_0_7/Component_Function_5/NAND4_in[2] ,
         \SB1_0_7/Component_Function_5/NAND4_in[1] ,
         \SB1_0_7/Component_Function_5/NAND4_in[0] ,
         \SB1_0_8/Component_Function_0/NAND4_in[3] ,
         \SB1_0_8/Component_Function_0/NAND4_in[2] ,
         \SB1_0_8/Component_Function_0/NAND4_in[1] ,
         \SB1_0_8/Component_Function_0/NAND4_in[0] ,
         \SB1_0_8/Component_Function_1/NAND4_in[3] ,
         \SB1_0_8/Component_Function_1/NAND4_in[2] ,
         \SB1_0_8/Component_Function_1/NAND4_in[1] ,
         \SB1_0_8/Component_Function_1/NAND4_in[0] ,
         \SB1_0_8/Component_Function_5/NAND4_in[1] ,
         \SB1_0_8/Component_Function_5/NAND4_in[0] ,
         \SB1_0_9/Component_Function_0/NAND4_in[3] ,
         \SB1_0_9/Component_Function_0/NAND4_in[2] ,
         \SB1_0_9/Component_Function_0/NAND4_in[1] ,
         \SB1_0_9/Component_Function_0/NAND4_in[0] ,
         \SB1_0_9/Component_Function_1/NAND4_in[3] ,
         \SB1_0_9/Component_Function_1/NAND4_in[2] ,
         \SB1_0_9/Component_Function_1/NAND4_in[1] ,
         \SB1_0_9/Component_Function_1/NAND4_in[0] ,
         \SB1_0_9/Component_Function_5/NAND4_in[3] ,
         \SB1_0_9/Component_Function_5/NAND4_in[1] ,
         \SB1_0_9/Component_Function_5/NAND4_in[0] ,
         \SB1_0_10/Component_Function_0/NAND4_in[3] ,
         \SB1_0_10/Component_Function_0/NAND4_in[2] ,
         \SB1_0_10/Component_Function_0/NAND4_in[1] ,
         \SB1_0_10/Component_Function_0/NAND4_in[0] ,
         \SB1_0_10/Component_Function_1/NAND4_in[3] ,
         \SB1_0_10/Component_Function_1/NAND4_in[2] ,
         \SB1_0_10/Component_Function_1/NAND4_in[1] ,
         \SB1_0_10/Component_Function_1/NAND4_in[0] ,
         \SB1_0_10/Component_Function_5/NAND4_in[3] ,
         \SB1_0_10/Component_Function_5/NAND4_in[2] ,
         \SB1_0_10/Component_Function_5/NAND4_in[0] ,
         \SB1_0_11/Component_Function_0/NAND4_in[3] ,
         \SB1_0_11/Component_Function_0/NAND4_in[2] ,
         \SB1_0_11/Component_Function_0/NAND4_in[1] ,
         \SB1_0_11/Component_Function_0/NAND4_in[0] ,
         \SB1_0_11/Component_Function_1/NAND4_in[3] ,
         \SB1_0_11/Component_Function_1/NAND4_in[2] ,
         \SB1_0_11/Component_Function_1/NAND4_in[1] ,
         \SB1_0_11/Component_Function_1/NAND4_in[0] ,
         \SB1_0_11/Component_Function_5/NAND4_in[3] ,
         \SB1_0_11/Component_Function_5/NAND4_in[1] ,
         \SB1_0_11/Component_Function_5/NAND4_in[0] ,
         \SB1_0_12/Component_Function_0/NAND4_in[3] ,
         \SB1_0_12/Component_Function_0/NAND4_in[1] ,
         \SB1_0_12/Component_Function_0/NAND4_in[0] ,
         \SB1_0_12/Component_Function_1/NAND4_in[3] ,
         \SB1_0_12/Component_Function_1/NAND4_in[2] ,
         \SB1_0_12/Component_Function_1/NAND4_in[1] ,
         \SB1_0_12/Component_Function_5/NAND4_in[2] ,
         \SB1_0_12/Component_Function_5/NAND4_in[1] ,
         \SB1_0_12/Component_Function_5/NAND4_in[0] ,
         \SB1_0_13/Component_Function_0/NAND4_in[1] ,
         \SB1_0_13/Component_Function_0/NAND4_in[0] ,
         \SB1_0_13/Component_Function_1/NAND4_in[3] ,
         \SB1_0_13/Component_Function_1/NAND4_in[2] ,
         \SB1_0_13/Component_Function_1/NAND4_in[1] ,
         \SB1_0_13/Component_Function_1/NAND4_in[0] ,
         \SB1_0_13/Component_Function_5/NAND4_in[2] ,
         \SB1_0_13/Component_Function_5/NAND4_in[1] ,
         \SB1_0_13/Component_Function_5/NAND4_in[0] ,
         \SB1_0_14/Component_Function_0/NAND4_in[3] ,
         \SB1_0_14/Component_Function_0/NAND4_in[2] ,
         \SB1_0_14/Component_Function_0/NAND4_in[1] ,
         \SB1_0_14/Component_Function_0/NAND4_in[0] ,
         \SB1_0_14/Component_Function_1/NAND4_in[3] ,
         \SB1_0_14/Component_Function_1/NAND4_in[2] ,
         \SB1_0_14/Component_Function_1/NAND4_in[1] ,
         \SB1_0_14/Component_Function_1/NAND4_in[0] ,
         \SB1_0_14/Component_Function_5/NAND4_in[3] ,
         \SB1_0_14/Component_Function_5/NAND4_in[2] ,
         \SB1_0_14/Component_Function_5/NAND4_in[1] ,
         \SB1_0_14/Component_Function_5/NAND4_in[0] ,
         \SB1_0_15/Component_Function_0/NAND4_in[3] ,
         \SB1_0_15/Component_Function_0/NAND4_in[2] ,
         \SB1_0_15/Component_Function_0/NAND4_in[1] ,
         \SB1_0_15/Component_Function_0/NAND4_in[0] ,
         \SB1_0_15/Component_Function_1/NAND4_in[3] ,
         \SB1_0_15/Component_Function_1/NAND4_in[2] ,
         \SB1_0_15/Component_Function_1/NAND4_in[1] ,
         \SB1_0_15/Component_Function_1/NAND4_in[0] ,
         \SB1_0_15/Component_Function_5/NAND4_in[3] ,
         \SB1_0_15/Component_Function_5/NAND4_in[2] ,
         \SB1_0_15/Component_Function_5/NAND4_in[1] ,
         \SB1_0_15/Component_Function_5/NAND4_in[0] ,
         \SB1_0_16/Component_Function_0/NAND4_in[3] ,
         \SB1_0_16/Component_Function_0/NAND4_in[2] ,
         \SB1_0_16/Component_Function_0/NAND4_in[1] ,
         \SB1_0_16/Component_Function_0/NAND4_in[0] ,
         \SB1_0_16/Component_Function_1/NAND4_in[2] ,
         \SB1_0_16/Component_Function_1/NAND4_in[1] ,
         \SB1_0_16/Component_Function_1/NAND4_in[0] ,
         \SB1_0_16/Component_Function_5/NAND4_in[2] ,
         \SB1_0_16/Component_Function_5/NAND4_in[0] ,
         \SB1_0_17/Component_Function_0/NAND4_in[3] ,
         \SB1_0_17/Component_Function_0/NAND4_in[2] ,
         \SB1_0_17/Component_Function_0/NAND4_in[1] ,
         \SB1_0_17/Component_Function_0/NAND4_in[0] ,
         \SB1_0_17/Component_Function_1/NAND4_in[3] ,
         \SB1_0_17/Component_Function_1/NAND4_in[2] ,
         \SB1_0_17/Component_Function_1/NAND4_in[1] ,
         \SB1_0_17/Component_Function_5/NAND4_in[2] ,
         \SB1_0_17/Component_Function_5/NAND4_in[0] ,
         \SB1_0_18/Component_Function_0/NAND4_in[2] ,
         \SB1_0_18/Component_Function_0/NAND4_in[1] ,
         \SB1_0_18/Component_Function_0/NAND4_in[0] ,
         \SB1_0_18/Component_Function_1/NAND4_in[3] ,
         \SB1_0_18/Component_Function_1/NAND4_in[2] ,
         \SB1_0_18/Component_Function_1/NAND4_in[1] ,
         \SB1_0_18/Component_Function_5/NAND4_in[2] ,
         \SB1_0_18/Component_Function_5/NAND4_in[1] ,
         \SB1_0_18/Component_Function_5/NAND4_in[0] ,
         \SB1_0_19/Component_Function_0/NAND4_in[2] ,
         \SB1_0_19/Component_Function_0/NAND4_in[1] ,
         \SB1_0_19/Component_Function_0/NAND4_in[0] ,
         \SB1_0_19/Component_Function_1/NAND4_in[3] ,
         \SB1_0_19/Component_Function_1/NAND4_in[2] ,
         \SB1_0_19/Component_Function_1/NAND4_in[1] ,
         \SB1_0_19/Component_Function_5/NAND4_in[3] ,
         \SB1_0_19/Component_Function_5/NAND4_in[1] ,
         \SB1_0_19/Component_Function_5/NAND4_in[0] ,
         \SB1_0_20/Component_Function_0/NAND4_in[3] ,
         \SB1_0_20/Component_Function_0/NAND4_in[2] ,
         \SB1_0_20/Component_Function_0/NAND4_in[1] ,
         \SB1_0_20/Component_Function_0/NAND4_in[0] ,
         \SB1_0_20/Component_Function_1/NAND4_in[2] ,
         \SB1_0_20/Component_Function_1/NAND4_in[1] ,
         \SB1_0_20/Component_Function_1/NAND4_in[0] ,
         \SB1_0_20/Component_Function_5/NAND4_in[3] ,
         \SB1_0_20/Component_Function_5/NAND4_in[1] ,
         \SB1_0_20/Component_Function_5/NAND4_in[0] ,
         \SB1_0_21/Component_Function_0/NAND4_in[2] ,
         \SB1_0_21/Component_Function_0/NAND4_in[1] ,
         \SB1_0_21/Component_Function_0/NAND4_in[0] ,
         \SB1_0_21/Component_Function_1/NAND4_in[3] ,
         \SB1_0_21/Component_Function_1/NAND4_in[2] ,
         \SB1_0_21/Component_Function_1/NAND4_in[1] ,
         \SB1_0_21/Component_Function_1/NAND4_in[0] ,
         \SB1_0_21/Component_Function_5/NAND4_in[3] ,
         \SB1_0_21/Component_Function_5/NAND4_in[2] ,
         \SB1_0_21/Component_Function_5/NAND4_in[0] ,
         \SB1_0_22/Component_Function_0/NAND4_in[3] ,
         \SB1_0_22/Component_Function_0/NAND4_in[2] ,
         \SB1_0_22/Component_Function_0/NAND4_in[1] ,
         \SB1_0_22/Component_Function_0/NAND4_in[0] ,
         \SB1_0_22/Component_Function_1/NAND4_in[3] ,
         \SB1_0_22/Component_Function_1/NAND4_in[2] ,
         \SB1_0_22/Component_Function_1/NAND4_in[1] ,
         \SB1_0_22/Component_Function_1/NAND4_in[0] ,
         \SB1_0_22/Component_Function_5/NAND4_in[2] ,
         \SB1_0_22/Component_Function_5/NAND4_in[0] ,
         \SB1_0_23/Component_Function_0/NAND4_in[3] ,
         \SB1_0_23/Component_Function_0/NAND4_in[1] ,
         \SB1_0_23/Component_Function_0/NAND4_in[0] ,
         \SB1_0_23/Component_Function_1/NAND4_in[3] ,
         \SB1_0_23/Component_Function_1/NAND4_in[2] ,
         \SB1_0_23/Component_Function_1/NAND4_in[1] ,
         \SB1_0_23/Component_Function_1/NAND4_in[0] ,
         \SB1_0_23/Component_Function_5/NAND4_in[2] ,
         \SB1_0_23/Component_Function_5/NAND4_in[1] ,
         \SB1_0_23/Component_Function_5/NAND4_in[0] ,
         \SB1_0_24/Component_Function_0/NAND4_in[3] ,
         \SB1_0_24/Component_Function_0/NAND4_in[2] ,
         \SB1_0_24/Component_Function_0/NAND4_in[1] ,
         \SB1_0_24/Component_Function_0/NAND4_in[0] ,
         \SB1_0_24/Component_Function_1/NAND4_in[2] ,
         \SB1_0_24/Component_Function_1/NAND4_in[1] ,
         \SB1_0_24/Component_Function_1/NAND4_in[0] ,
         \SB1_0_24/Component_Function_5/NAND4_in[2] ,
         \SB1_0_24/Component_Function_5/NAND4_in[1] ,
         \SB1_0_24/Component_Function_5/NAND4_in[0] ,
         \SB1_0_25/Component_Function_0/NAND4_in[3] ,
         \SB1_0_25/Component_Function_0/NAND4_in[1] ,
         \SB1_0_25/Component_Function_0/NAND4_in[0] ,
         \SB1_0_25/Component_Function_1/NAND4_in[3] ,
         \SB1_0_25/Component_Function_1/NAND4_in[2] ,
         \SB1_0_25/Component_Function_1/NAND4_in[1] ,
         \SB1_0_25/Component_Function_1/NAND4_in[0] ,
         \SB1_0_25/Component_Function_5/NAND4_in[2] ,
         \SB1_0_25/Component_Function_5/NAND4_in[1] ,
         \SB1_0_25/Component_Function_5/NAND4_in[0] ,
         \SB1_0_26/Component_Function_0/NAND4_in[3] ,
         \SB1_0_26/Component_Function_0/NAND4_in[1] ,
         \SB1_0_26/Component_Function_0/NAND4_in[0] ,
         \SB1_0_26/Component_Function_1/NAND4_in[3] ,
         \SB1_0_26/Component_Function_1/NAND4_in[2] ,
         \SB1_0_26/Component_Function_1/NAND4_in[1] ,
         \SB1_0_26/Component_Function_1/NAND4_in[0] ,
         \SB1_0_26/Component_Function_5/NAND4_in[3] ,
         \SB1_0_26/Component_Function_5/NAND4_in[2] ,
         \SB1_0_26/Component_Function_5/NAND4_in[1] ,
         \SB1_0_26/Component_Function_5/NAND4_in[0] ,
         \SB1_0_27/Component_Function_0/NAND4_in[2] ,
         \SB1_0_27/Component_Function_0/NAND4_in[1] ,
         \SB1_0_27/Component_Function_0/NAND4_in[0] ,
         \SB1_0_27/Component_Function_1/NAND4_in[3] ,
         \SB1_0_27/Component_Function_1/NAND4_in[2] ,
         \SB1_0_27/Component_Function_1/NAND4_in[1] ,
         \SB1_0_27/Component_Function_1/NAND4_in[0] ,
         \SB1_0_27/Component_Function_5/NAND4_in[3] ,
         \SB1_0_27/Component_Function_5/NAND4_in[1] ,
         \SB1_0_27/Component_Function_5/NAND4_in[0] ,
         \SB1_0_28/Component_Function_0/NAND4_in[3] ,
         \SB1_0_28/Component_Function_0/NAND4_in[2] ,
         \SB1_0_28/Component_Function_0/NAND4_in[1] ,
         \SB1_0_28/Component_Function_0/NAND4_in[0] ,
         \SB1_0_28/Component_Function_1/NAND4_in[3] ,
         \SB1_0_28/Component_Function_1/NAND4_in[2] ,
         \SB1_0_28/Component_Function_1/NAND4_in[1] ,
         \SB1_0_28/Component_Function_1/NAND4_in[0] ,
         \SB1_0_28/Component_Function_5/NAND4_in[3] ,
         \SB1_0_28/Component_Function_5/NAND4_in[1] ,
         \SB1_0_28/Component_Function_5/NAND4_in[0] ,
         \SB1_0_29/Component_Function_0/NAND4_in[3] ,
         \SB1_0_29/Component_Function_0/NAND4_in[1] ,
         \SB1_0_29/Component_Function_0/NAND4_in[0] ,
         \SB1_0_29/Component_Function_1/NAND4_in[2] ,
         \SB1_0_29/Component_Function_1/NAND4_in[1] ,
         \SB1_0_29/Component_Function_1/NAND4_in[0] ,
         \SB1_0_29/Component_Function_5/NAND4_in[2] ,
         \SB1_0_29/Component_Function_5/NAND4_in[0] ,
         \SB1_0_30/Component_Function_0/NAND4_in[3] ,
         \SB1_0_30/Component_Function_0/NAND4_in[2] ,
         \SB1_0_30/Component_Function_0/NAND4_in[1] ,
         \SB1_0_30/Component_Function_0/NAND4_in[0] ,
         \SB1_0_30/Component_Function_1/NAND4_in[3] ,
         \SB1_0_30/Component_Function_1/NAND4_in[2] ,
         \SB1_0_30/Component_Function_1/NAND4_in[1] ,
         \SB1_0_30/Component_Function_1/NAND4_in[0] ,
         \SB1_0_30/Component_Function_5/NAND4_in[3] ,
         \SB1_0_30/Component_Function_5/NAND4_in[1] ,
         \SB1_0_30/Component_Function_5/NAND4_in[0] ,
         \SB1_0_31/Component_Function_0/NAND4_in[3] ,
         \SB1_0_31/Component_Function_0/NAND4_in[2] ,
         \SB1_0_31/Component_Function_0/NAND4_in[1] ,
         \SB1_0_31/Component_Function_0/NAND4_in[0] ,
         \SB1_0_31/Component_Function_1/NAND4_in[3] ,
         \SB1_0_31/Component_Function_1/NAND4_in[2] ,
         \SB1_0_31/Component_Function_1/NAND4_in[1] ,
         \SB1_0_31/Component_Function_1/NAND4_in[0] ,
         \SB1_0_31/Component_Function_5/NAND4_in[3] ,
         \SB1_0_31/Component_Function_5/NAND4_in[2] ,
         \SB1_0_31/Component_Function_5/NAND4_in[1] ,
         \SB2_0_0/Component_Function_0/NAND4_in[2] ,
         \SB2_0_0/Component_Function_0/NAND4_in[1] ,
         \SB2_0_0/Component_Function_0/NAND4_in[0] ,
         \SB2_0_0/Component_Function_1/NAND4_in[3] ,
         \SB2_0_0/Component_Function_1/NAND4_in[2] ,
         \SB2_0_0/Component_Function_1/NAND4_in[1] ,
         \SB2_0_0/Component_Function_1/NAND4_in[0] ,
         \SB2_0_0/Component_Function_5/NAND4_in[3] ,
         \SB2_0_0/Component_Function_5/NAND4_in[2] ,
         \SB2_0_0/Component_Function_5/NAND4_in[0] ,
         \SB2_0_1/Component_Function_0/NAND4_in[2] ,
         \SB2_0_1/Component_Function_0/NAND4_in[0] ,
         \SB2_0_1/Component_Function_1/NAND4_in[3] ,
         \SB2_0_1/Component_Function_1/NAND4_in[1] ,
         \SB2_0_1/Component_Function_1/NAND4_in[0] ,
         \SB2_0_1/Component_Function_5/NAND4_in[3] ,
         \SB2_0_1/Component_Function_5/NAND4_in[2] ,
         \SB2_0_1/Component_Function_5/NAND4_in[1] ,
         \SB2_0_1/Component_Function_5/NAND4_in[0] ,
         \SB2_0_2/Component_Function_0/NAND4_in[3] ,
         \SB2_0_2/Component_Function_0/NAND4_in[1] ,
         \SB2_0_2/Component_Function_0/NAND4_in[0] ,
         \SB2_0_2/Component_Function_1/NAND4_in[3] ,
         \SB2_0_2/Component_Function_1/NAND4_in[2] ,
         \SB2_0_2/Component_Function_1/NAND4_in[1] ,
         \SB2_0_2/Component_Function_1/NAND4_in[0] ,
         \SB2_0_2/Component_Function_5/NAND4_in[2] ,
         \SB2_0_2/Component_Function_5/NAND4_in[1] ,
         \SB2_0_2/Component_Function_5/NAND4_in[0] ,
         \SB2_0_3/Component_Function_0/NAND4_in[3] ,
         \SB2_0_3/Component_Function_0/NAND4_in[2] ,
         \SB2_0_3/Component_Function_0/NAND4_in[1] ,
         \SB2_0_3/Component_Function_0/NAND4_in[0] ,
         \SB2_0_3/Component_Function_1/NAND4_in[3] ,
         \SB2_0_3/Component_Function_1/NAND4_in[2] ,
         \SB2_0_3/Component_Function_1/NAND4_in[1] ,
         \SB2_0_3/Component_Function_1/NAND4_in[0] ,
         \SB2_0_3/Component_Function_5/NAND4_in[1] ,
         \SB2_0_3/Component_Function_5/NAND4_in[0] ,
         \SB2_0_4/Component_Function_0/NAND4_in[3] ,
         \SB2_0_4/Component_Function_0/NAND4_in[2] ,
         \SB2_0_4/Component_Function_0/NAND4_in[1] ,
         \SB2_0_4/Component_Function_0/NAND4_in[0] ,
         \SB2_0_4/Component_Function_1/NAND4_in[2] ,
         \SB2_0_4/Component_Function_1/NAND4_in[1] ,
         \SB2_0_4/Component_Function_5/NAND4_in[2] ,
         \SB2_0_4/Component_Function_5/NAND4_in[0] ,
         \SB2_0_5/Component_Function_0/NAND4_in[3] ,
         \SB2_0_5/Component_Function_0/NAND4_in[2] ,
         \SB2_0_5/Component_Function_0/NAND4_in[0] ,
         \SB2_0_5/Component_Function_1/NAND4_in[3] ,
         \SB2_0_5/Component_Function_1/NAND4_in[2] ,
         \SB2_0_5/Component_Function_1/NAND4_in[1] ,
         \SB2_0_5/Component_Function_1/NAND4_in[0] ,
         \SB2_0_5/Component_Function_5/NAND4_in[3] ,
         \SB2_0_5/Component_Function_5/NAND4_in[2] ,
         \SB2_0_5/Component_Function_5/NAND4_in[1] ,
         \SB2_0_5/Component_Function_5/NAND4_in[0] ,
         \SB2_0_6/Component_Function_0/NAND4_in[3] ,
         \SB2_0_6/Component_Function_0/NAND4_in[2] ,
         \SB2_0_6/Component_Function_0/NAND4_in[1] ,
         \SB2_0_6/Component_Function_0/NAND4_in[0] ,
         \SB2_0_6/Component_Function_1/NAND4_in[3] ,
         \SB2_0_6/Component_Function_1/NAND4_in[1] ,
         \SB2_0_6/Component_Function_1/NAND4_in[0] ,
         \SB2_0_6/Component_Function_5/NAND4_in[3] ,
         \SB2_0_6/Component_Function_5/NAND4_in[1] ,
         \SB2_0_6/Component_Function_5/NAND4_in[0] ,
         \SB2_0_7/Component_Function_0/NAND4_in[3] ,
         \SB2_0_7/Component_Function_0/NAND4_in[1] ,
         \SB2_0_7/Component_Function_0/NAND4_in[0] ,
         \SB2_0_7/Component_Function_1/NAND4_in[3] ,
         \SB2_0_7/Component_Function_1/NAND4_in[2] ,
         \SB2_0_7/Component_Function_1/NAND4_in[1] ,
         \SB2_0_7/Component_Function_1/NAND4_in[0] ,
         \SB2_0_7/Component_Function_5/NAND4_in[1] ,
         \SB2_0_7/Component_Function_5/NAND4_in[0] ,
         \SB2_0_8/Component_Function_0/NAND4_in[3] ,
         \SB2_0_8/Component_Function_0/NAND4_in[2] ,
         \SB2_0_8/Component_Function_0/NAND4_in[1] ,
         \SB2_0_8/Component_Function_0/NAND4_in[0] ,
         \SB2_0_8/Component_Function_1/NAND4_in[3] ,
         \SB2_0_8/Component_Function_1/NAND4_in[2] ,
         \SB2_0_8/Component_Function_1/NAND4_in[1] ,
         \SB2_0_8/Component_Function_1/NAND4_in[0] ,
         \SB2_0_8/Component_Function_5/NAND4_in[3] ,
         \SB2_0_8/Component_Function_5/NAND4_in[2] ,
         \SB2_0_8/Component_Function_5/NAND4_in[0] ,
         \SB2_0_9/Component_Function_0/NAND4_in[3] ,
         \SB2_0_9/Component_Function_0/NAND4_in[2] ,
         \SB2_0_9/Component_Function_0/NAND4_in[1] ,
         \SB2_0_9/Component_Function_0/NAND4_in[0] ,
         \SB2_0_9/Component_Function_1/NAND4_in[3] ,
         \SB2_0_9/Component_Function_1/NAND4_in[2] ,
         \SB2_0_9/Component_Function_1/NAND4_in[1] ,
         \SB2_0_9/Component_Function_1/NAND4_in[0] ,
         \SB2_0_9/Component_Function_5/NAND4_in[0] ,
         \SB2_0_10/Component_Function_0/NAND4_in[2] ,
         \SB2_0_10/Component_Function_0/NAND4_in[1] ,
         \SB2_0_10/Component_Function_0/NAND4_in[0] ,
         \SB2_0_10/Component_Function_1/NAND4_in[3] ,
         \SB2_0_10/Component_Function_1/NAND4_in[2] ,
         \SB2_0_10/Component_Function_1/NAND4_in[1] ,
         \SB2_0_10/Component_Function_1/NAND4_in[0] ,
         \SB2_0_10/Component_Function_5/NAND4_in[3] ,
         \SB2_0_10/Component_Function_5/NAND4_in[2] ,
         \SB2_0_10/Component_Function_5/NAND4_in[1] ,
         \SB2_0_11/Component_Function_0/NAND4_in[2] ,
         \SB2_0_11/Component_Function_0/NAND4_in[1] ,
         \SB2_0_11/Component_Function_0/NAND4_in[0] ,
         \SB2_0_11/Component_Function_1/NAND4_in[2] ,
         \SB2_0_11/Component_Function_1/NAND4_in[1] ,
         \SB2_0_11/Component_Function_1/NAND4_in[0] ,
         \SB2_0_11/Component_Function_5/NAND4_in[3] ,
         \SB2_0_11/Component_Function_5/NAND4_in[1] ,
         \SB2_0_11/Component_Function_5/NAND4_in[0] ,
         \SB2_0_12/Component_Function_0/NAND4_in[3] ,
         \SB2_0_12/Component_Function_0/NAND4_in[2] ,
         \SB2_0_12/Component_Function_0/NAND4_in[1] ,
         \SB2_0_12/Component_Function_0/NAND4_in[0] ,
         \SB2_0_12/Component_Function_1/NAND4_in[3] ,
         \SB2_0_12/Component_Function_1/NAND4_in[2] ,
         \SB2_0_12/Component_Function_1/NAND4_in[1] ,
         \SB2_0_12/Component_Function_1/NAND4_in[0] ,
         \SB2_0_12/Component_Function_5/NAND4_in[1] ,
         \SB2_0_12/Component_Function_5/NAND4_in[0] ,
         \SB2_0_13/Component_Function_0/NAND4_in[2] ,
         \SB2_0_13/Component_Function_0/NAND4_in[1] ,
         \SB2_0_13/Component_Function_0/NAND4_in[0] ,
         \SB2_0_13/Component_Function_1/NAND4_in[2] ,
         \SB2_0_13/Component_Function_1/NAND4_in[1] ,
         \SB2_0_13/Component_Function_1/NAND4_in[0] ,
         \SB2_0_13/Component_Function_5/NAND4_in[2] ,
         \SB2_0_13/Component_Function_5/NAND4_in[0] ,
         \SB2_0_14/Component_Function_0/NAND4_in[3] ,
         \SB2_0_14/Component_Function_0/NAND4_in[2] ,
         \SB2_0_14/Component_Function_0/NAND4_in[0] ,
         \SB2_0_14/Component_Function_1/NAND4_in[3] ,
         \SB2_0_14/Component_Function_1/NAND4_in[1] ,
         \SB2_0_14/Component_Function_1/NAND4_in[0] ,
         \SB2_0_14/Component_Function_5/NAND4_in[1] ,
         \SB2_0_14/Component_Function_5/NAND4_in[0] ,
         \SB2_0_15/Component_Function_0/NAND4_in[3] ,
         \SB2_0_15/Component_Function_0/NAND4_in[0] ,
         \SB2_0_15/Component_Function_1/NAND4_in[3] ,
         \SB2_0_15/Component_Function_1/NAND4_in[2] ,
         \SB2_0_15/Component_Function_1/NAND4_in[1] ,
         \SB2_0_15/Component_Function_1/NAND4_in[0] ,
         \SB2_0_15/Component_Function_5/NAND4_in[3] ,
         \SB2_0_15/Component_Function_5/NAND4_in[0] ,
         \SB2_0_16/Component_Function_0/NAND4_in[3] ,
         \SB2_0_16/Component_Function_0/NAND4_in[1] ,
         \SB2_0_16/Component_Function_0/NAND4_in[0] ,
         \SB2_0_16/Component_Function_1/NAND4_in[3] ,
         \SB2_0_16/Component_Function_1/NAND4_in[2] ,
         \SB2_0_16/Component_Function_1/NAND4_in[1] ,
         \SB2_0_16/Component_Function_1/NAND4_in[0] ,
         \SB2_0_16/Component_Function_5/NAND4_in[2] ,
         \SB2_0_16/Component_Function_5/NAND4_in[0] ,
         \SB2_0_17/Component_Function_0/NAND4_in[3] ,
         \SB2_0_17/Component_Function_0/NAND4_in[2] ,
         \SB2_0_17/Component_Function_0/NAND4_in[0] ,
         \SB2_0_17/Component_Function_1/NAND4_in[2] ,
         \SB2_0_17/Component_Function_1/NAND4_in[1] ,
         \SB2_0_17/Component_Function_1/NAND4_in[0] ,
         \SB2_0_17/Component_Function_5/NAND4_in[2] ,
         \SB2_0_17/Component_Function_5/NAND4_in[0] ,
         \SB2_0_18/Component_Function_0/NAND4_in[2] ,
         \SB2_0_18/Component_Function_0/NAND4_in[1] ,
         \SB2_0_18/Component_Function_1/NAND4_in[3] ,
         \SB2_0_18/Component_Function_1/NAND4_in[2] ,
         \SB2_0_18/Component_Function_1/NAND4_in[1] ,
         \SB2_0_18/Component_Function_1/NAND4_in[0] ,
         \SB2_0_18/Component_Function_5/NAND4_in[2] ,
         \SB2_0_18/Component_Function_5/NAND4_in[1] ,
         \SB2_0_18/Component_Function_5/NAND4_in[0] ,
         \SB2_0_19/Component_Function_0/NAND4_in[3] ,
         \SB2_0_19/Component_Function_0/NAND4_in[2] ,
         \SB2_0_19/Component_Function_0/NAND4_in[1] ,
         \SB2_0_19/Component_Function_0/NAND4_in[0] ,
         \SB2_0_19/Component_Function_1/NAND4_in[3] ,
         \SB2_0_19/Component_Function_1/NAND4_in[2] ,
         \SB2_0_19/Component_Function_1/NAND4_in[1] ,
         \SB2_0_19/Component_Function_1/NAND4_in[0] ,
         \SB2_0_19/Component_Function_5/NAND4_in[3] ,
         \SB2_0_19/Component_Function_5/NAND4_in[0] ,
         \SB2_0_20/Component_Function_0/NAND4_in[3] ,
         \SB2_0_20/Component_Function_0/NAND4_in[2] ,
         \SB2_0_20/Component_Function_0/NAND4_in[0] ,
         \SB2_0_20/Component_Function_1/NAND4_in[3] ,
         \SB2_0_20/Component_Function_1/NAND4_in[2] ,
         \SB2_0_20/Component_Function_1/NAND4_in[1] ,
         \SB2_0_20/Component_Function_1/NAND4_in[0] ,
         \SB2_0_20/Component_Function_5/NAND4_in[3] ,
         \SB2_0_20/Component_Function_5/NAND4_in[2] ,
         \SB2_0_20/Component_Function_5/NAND4_in[1] ,
         \SB2_0_20/Component_Function_5/NAND4_in[0] ,
         \SB2_0_21/Component_Function_0/NAND4_in[3] ,
         \SB2_0_21/Component_Function_0/NAND4_in[1] ,
         \SB2_0_21/Component_Function_0/NAND4_in[0] ,
         \SB2_0_21/Component_Function_1/NAND4_in[3] ,
         \SB2_0_21/Component_Function_1/NAND4_in[2] ,
         \SB2_0_21/Component_Function_1/NAND4_in[1] ,
         \SB2_0_21/Component_Function_1/NAND4_in[0] ,
         \SB2_0_21/Component_Function_5/NAND4_in[0] ,
         \SB2_0_22/Component_Function_0/NAND4_in[2] ,
         \SB2_0_22/Component_Function_0/NAND4_in[1] ,
         \SB2_0_22/Component_Function_0/NAND4_in[0] ,
         \SB2_0_22/Component_Function_1/NAND4_in[3] ,
         \SB2_0_22/Component_Function_1/NAND4_in[2] ,
         \SB2_0_22/Component_Function_1/NAND4_in[1] ,
         \SB2_0_22/Component_Function_1/NAND4_in[0] ,
         \SB2_0_22/Component_Function_5/NAND4_in[0] ,
         \SB2_0_23/Component_Function_0/NAND4_in[3] ,
         \SB2_0_23/Component_Function_0/NAND4_in[1] ,
         \SB2_0_23/Component_Function_0/NAND4_in[0] ,
         \SB2_0_23/Component_Function_1/NAND4_in[3] ,
         \SB2_0_23/Component_Function_1/NAND4_in[2] ,
         \SB2_0_23/Component_Function_1/NAND4_in[1] ,
         \SB2_0_23/Component_Function_1/NAND4_in[0] ,
         \SB2_0_23/Component_Function_5/NAND4_in[2] ,
         \SB2_0_23/Component_Function_5/NAND4_in[0] ,
         \SB2_0_24/Component_Function_0/NAND4_in[3] ,
         \SB2_0_24/Component_Function_0/NAND4_in[2] ,
         \SB2_0_24/Component_Function_0/NAND4_in[0] ,
         \SB2_0_24/Component_Function_1/NAND4_in[3] ,
         \SB2_0_24/Component_Function_1/NAND4_in[2] ,
         \SB2_0_24/Component_Function_1/NAND4_in[0] ,
         \SB2_0_24/Component_Function_5/NAND4_in[3] ,
         \SB2_0_24/Component_Function_5/NAND4_in[0] ,
         \SB2_0_25/Component_Function_0/NAND4_in[1] ,
         \SB2_0_25/Component_Function_0/NAND4_in[0] ,
         \SB2_0_25/Component_Function_1/NAND4_in[3] ,
         \SB2_0_25/Component_Function_1/NAND4_in[2] ,
         \SB2_0_25/Component_Function_1/NAND4_in[0] ,
         \SB2_0_25/Component_Function_5/NAND4_in[3] ,
         \SB2_0_25/Component_Function_5/NAND4_in[1] ,
         \SB2_0_25/Component_Function_5/NAND4_in[0] ,
         \SB2_0_26/Component_Function_0/NAND4_in[3] ,
         \SB2_0_26/Component_Function_0/NAND4_in[2] ,
         \SB2_0_26/Component_Function_0/NAND4_in[1] ,
         \SB2_0_26/Component_Function_0/NAND4_in[0] ,
         \SB2_0_26/Component_Function_1/NAND4_in[3] ,
         \SB2_0_26/Component_Function_1/NAND4_in[2] ,
         \SB2_0_26/Component_Function_1/NAND4_in[1] ,
         \SB2_0_26/Component_Function_5/NAND4_in[3] ,
         \SB2_0_27/Component_Function_0/NAND4_in[3] ,
         \SB2_0_27/Component_Function_0/NAND4_in[0] ,
         \SB2_0_27/Component_Function_1/NAND4_in[3] ,
         \SB2_0_27/Component_Function_1/NAND4_in[2] ,
         \SB2_0_27/Component_Function_1/NAND4_in[1] ,
         \SB2_0_27/Component_Function_1/NAND4_in[0] ,
         \SB2_0_27/Component_Function_5/NAND4_in[2] ,
         \SB2_0_27/Component_Function_5/NAND4_in[0] ,
         \SB2_0_28/Component_Function_0/NAND4_in[2] ,
         \SB2_0_28/Component_Function_0/NAND4_in[1] ,
         \SB2_0_28/Component_Function_0/NAND4_in[0] ,
         \SB2_0_28/Component_Function_1/NAND4_in[3] ,
         \SB2_0_28/Component_Function_1/NAND4_in[1] ,
         \SB2_0_28/Component_Function_1/NAND4_in[0] ,
         \SB2_0_28/Component_Function_5/NAND4_in[1] ,
         \SB2_0_28/Component_Function_5/NAND4_in[0] ,
         \SB2_0_29/Component_Function_0/NAND4_in[3] ,
         \SB2_0_29/Component_Function_0/NAND4_in[2] ,
         \SB2_0_29/Component_Function_0/NAND4_in[1] ,
         \SB2_0_29/Component_Function_0/NAND4_in[0] ,
         \SB2_0_29/Component_Function_1/NAND4_in[3] ,
         \SB2_0_29/Component_Function_1/NAND4_in[2] ,
         \SB2_0_29/Component_Function_1/NAND4_in[1] ,
         \SB2_0_29/Component_Function_1/NAND4_in[0] ,
         \SB2_0_29/Component_Function_5/NAND4_in[1] ,
         \SB2_0_29/Component_Function_5/NAND4_in[0] ,
         \SB2_0_30/Component_Function_0/NAND4_in[3] ,
         \SB2_0_30/Component_Function_0/NAND4_in[2] ,
         \SB2_0_30/Component_Function_0/NAND4_in[0] ,
         \SB2_0_30/Component_Function_1/NAND4_in[2] ,
         \SB2_0_30/Component_Function_1/NAND4_in[1] ,
         \SB2_0_30/Component_Function_1/NAND4_in[0] ,
         \SB2_0_30/Component_Function_5/NAND4_in[2] ,
         \SB2_0_30/Component_Function_5/NAND4_in[0] ,
         \SB2_0_31/Component_Function_0/NAND4_in[3] ,
         \SB2_0_31/Component_Function_0/NAND4_in[2] ,
         \SB2_0_31/Component_Function_0/NAND4_in[1] ,
         \SB2_0_31/Component_Function_0/NAND4_in[0] ,
         \SB2_0_31/Component_Function_1/NAND4_in[3] ,
         \SB2_0_31/Component_Function_1/NAND4_in[2] ,
         \SB2_0_31/Component_Function_1/NAND4_in[1] ,
         \SB2_0_31/Component_Function_1/NAND4_in[0] ,
         \SB2_0_31/Component_Function_5/NAND4_in[1] ,
         \SB2_0_31/Component_Function_5/NAND4_in[0] ,
         \SB1_1_0/Component_Function_0/NAND4_in[2] ,
         \SB1_1_0/Component_Function_0/NAND4_in[1] ,
         \SB1_1_0/Component_Function_0/NAND4_in[0] ,
         \SB1_1_0/Component_Function_1/NAND4_in[3] ,
         \SB1_1_0/Component_Function_5/NAND4_in[2] ,
         \SB1_1_0/Component_Function_5/NAND4_in[0] ,
         \SB1_1_1/Component_Function_0/NAND4_in[2] ,
         \SB1_1_1/Component_Function_0/NAND4_in[1] ,
         \SB1_1_1/Component_Function_0/NAND4_in[0] ,
         \SB1_1_1/Component_Function_1/NAND4_in[2] ,
         \SB1_1_1/Component_Function_1/NAND4_in[1] ,
         \SB1_1_1/Component_Function_1/NAND4_in[0] ,
         \SB1_1_1/Component_Function_5/NAND4_in[1] ,
         \SB1_1_1/Component_Function_5/NAND4_in[0] ,
         \SB1_1_2/Component_Function_0/NAND4_in[3] ,
         \SB1_1_2/Component_Function_0/NAND4_in[2] ,
         \SB1_1_2/Component_Function_0/NAND4_in[1] ,
         \SB1_1_2/Component_Function_0/NAND4_in[0] ,
         \SB1_1_2/Component_Function_1/NAND4_in[2] ,
         \SB1_1_2/Component_Function_1/NAND4_in[1] ,
         \SB1_1_2/Component_Function_1/NAND4_in[0] ,
         \SB1_1_2/Component_Function_5/NAND4_in[3] ,
         \SB1_1_2/Component_Function_5/NAND4_in[0] ,
         \SB1_1_3/Component_Function_0/NAND4_in[2] ,
         \SB1_1_3/Component_Function_0/NAND4_in[1] ,
         \SB1_1_3/Component_Function_0/NAND4_in[0] ,
         \SB1_1_3/Component_Function_1/NAND4_in[3] ,
         \SB1_1_3/Component_Function_1/NAND4_in[2] ,
         \SB1_1_3/Component_Function_1/NAND4_in[1] ,
         \SB1_1_3/Component_Function_1/NAND4_in[0] ,
         \SB1_1_3/Component_Function_5/NAND4_in[2] ,
         \SB1_1_3/Component_Function_5/NAND4_in[1] ,
         \SB1_1_3/Component_Function_5/NAND4_in[0] ,
         \SB1_1_4/Component_Function_0/NAND4_in[3] ,
         \SB1_1_4/Component_Function_0/NAND4_in[2] ,
         \SB1_1_4/Component_Function_0/NAND4_in[1] ,
         \SB1_1_4/Component_Function_0/NAND4_in[0] ,
         \SB1_1_4/Component_Function_1/NAND4_in[3] ,
         \SB1_1_4/Component_Function_1/NAND4_in[1] ,
         \SB1_1_4/Component_Function_1/NAND4_in[0] ,
         \SB1_1_4/Component_Function_5/NAND4_in[2] ,
         \SB1_1_4/Component_Function_5/NAND4_in[1] ,
         \SB1_1_4/Component_Function_5/NAND4_in[0] ,
         \SB1_1_5/Component_Function_0/NAND4_in[3] ,
         \SB1_1_5/Component_Function_0/NAND4_in[2] ,
         \SB1_1_5/Component_Function_0/NAND4_in[1] ,
         \SB1_1_5/Component_Function_0/NAND4_in[0] ,
         \SB1_1_5/Component_Function_1/NAND4_in[3] ,
         \SB1_1_5/Component_Function_1/NAND4_in[2] ,
         \SB1_1_5/Component_Function_1/NAND4_in[1] ,
         \SB1_1_5/Component_Function_1/NAND4_in[0] ,
         \SB1_1_5/Component_Function_5/NAND4_in[3] ,
         \SB1_1_5/Component_Function_5/NAND4_in[1] ,
         \SB1_1_5/Component_Function_5/NAND4_in[0] ,
         \SB1_1_6/Component_Function_0/NAND4_in[3] ,
         \SB1_1_6/Component_Function_0/NAND4_in[2] ,
         \SB1_1_6/Component_Function_0/NAND4_in[1] ,
         \SB1_1_6/Component_Function_0/NAND4_in[0] ,
         \SB1_1_6/Component_Function_1/NAND4_in[3] ,
         \SB1_1_6/Component_Function_1/NAND4_in[2] ,
         \SB1_1_6/Component_Function_1/NAND4_in[1] ,
         \SB1_1_6/Component_Function_1/NAND4_in[0] ,
         \SB1_1_6/Component_Function_5/NAND4_in[0] ,
         \SB1_1_7/Component_Function_0/NAND4_in[3] ,
         \SB1_1_7/Component_Function_0/NAND4_in[2] ,
         \SB1_1_7/Component_Function_0/NAND4_in[1] ,
         \SB1_1_7/Component_Function_0/NAND4_in[0] ,
         \SB1_1_7/Component_Function_1/NAND4_in[3] ,
         \SB1_1_7/Component_Function_1/NAND4_in[1] ,
         \SB1_1_7/Component_Function_1/NAND4_in[0] ,
         \SB1_1_7/Component_Function_5/NAND4_in[3] ,
         \SB1_1_7/Component_Function_5/NAND4_in[2] ,
         \SB1_1_7/Component_Function_5/NAND4_in[1] ,
         \SB1_1_7/Component_Function_5/NAND4_in[0] ,
         \SB1_1_8/Component_Function_0/NAND4_in[3] ,
         \SB1_1_8/Component_Function_0/NAND4_in[1] ,
         \SB1_1_8/Component_Function_0/NAND4_in[0] ,
         \SB1_1_8/Component_Function_1/NAND4_in[3] ,
         \SB1_1_8/Component_Function_1/NAND4_in[2] ,
         \SB1_1_8/Component_Function_1/NAND4_in[1] ,
         \SB1_1_8/Component_Function_1/NAND4_in[0] ,
         \SB1_1_8/Component_Function_5/NAND4_in[3] ,
         \SB1_1_8/Component_Function_5/NAND4_in[2] ,
         \SB1_1_8/Component_Function_5/NAND4_in[1] ,
         \SB1_1_8/Component_Function_5/NAND4_in[0] ,
         \SB1_1_9/Component_Function_0/NAND4_in[2] ,
         \SB1_1_9/Component_Function_0/NAND4_in[1] ,
         \SB1_1_9/Component_Function_0/NAND4_in[0] ,
         \SB1_1_9/Component_Function_1/NAND4_in[3] ,
         \SB1_1_9/Component_Function_1/NAND4_in[2] ,
         \SB1_1_9/Component_Function_1/NAND4_in[1] ,
         \SB1_1_9/Component_Function_1/NAND4_in[0] ,
         \SB1_1_9/Component_Function_5/NAND4_in[1] ,
         \SB1_1_9/Component_Function_5/NAND4_in[0] ,
         \SB1_1_10/Component_Function_0/NAND4_in[2] ,
         \SB1_1_10/Component_Function_0/NAND4_in[1] ,
         \SB1_1_10/Component_Function_0/NAND4_in[0] ,
         \SB1_1_10/Component_Function_1/NAND4_in[3] ,
         \SB1_1_10/Component_Function_1/NAND4_in[2] ,
         \SB1_1_10/Component_Function_1/NAND4_in[1] ,
         \SB1_1_10/Component_Function_1/NAND4_in[0] ,
         \SB1_1_10/Component_Function_5/NAND4_in[1] ,
         \SB1_1_10/Component_Function_5/NAND4_in[0] ,
         \SB1_1_11/Component_Function_0/NAND4_in[3] ,
         \SB1_1_11/Component_Function_0/NAND4_in[2] ,
         \SB1_1_11/Component_Function_0/NAND4_in[1] ,
         \SB1_1_11/Component_Function_0/NAND4_in[0] ,
         \SB1_1_11/Component_Function_1/NAND4_in[2] ,
         \SB1_1_11/Component_Function_1/NAND4_in[1] ,
         \SB1_1_11/Component_Function_1/NAND4_in[0] ,
         \SB1_1_11/Component_Function_5/NAND4_in[2] ,
         \SB1_1_11/Component_Function_5/NAND4_in[1] ,
         \SB1_1_11/Component_Function_5/NAND4_in[0] ,
         \SB1_1_12/Component_Function_0/NAND4_in[2] ,
         \SB1_1_12/Component_Function_0/NAND4_in[1] ,
         \SB1_1_12/Component_Function_0/NAND4_in[0] ,
         \SB1_1_12/Component_Function_1/NAND4_in[3] ,
         \SB1_1_12/Component_Function_1/NAND4_in[2] ,
         \SB1_1_12/Component_Function_1/NAND4_in[1] ,
         \SB1_1_12/Component_Function_1/NAND4_in[0] ,
         \SB1_1_12/Component_Function_5/NAND4_in[3] ,
         \SB1_1_12/Component_Function_5/NAND4_in[1] ,
         \SB1_1_13/Component_Function_0/NAND4_in[3] ,
         \SB1_1_13/Component_Function_0/NAND4_in[2] ,
         \SB1_1_13/Component_Function_0/NAND4_in[1] ,
         \SB1_1_13/Component_Function_0/NAND4_in[0] ,
         \SB1_1_13/Component_Function_1/NAND4_in[3] ,
         \SB1_1_13/Component_Function_1/NAND4_in[2] ,
         \SB1_1_13/Component_Function_1/NAND4_in[1] ,
         \SB1_1_13/Component_Function_1/NAND4_in[0] ,
         \SB1_1_13/Component_Function_5/NAND4_in[3] ,
         \SB1_1_13/Component_Function_5/NAND4_in[1] ,
         \SB1_1_14/Component_Function_0/NAND4_in[3] ,
         \SB1_1_14/Component_Function_0/NAND4_in[2] ,
         \SB1_1_14/Component_Function_0/NAND4_in[1] ,
         \SB1_1_14/Component_Function_0/NAND4_in[0] ,
         \SB1_1_14/Component_Function_1/NAND4_in[2] ,
         \SB1_1_14/Component_Function_1/NAND4_in[1] ,
         \SB1_1_14/Component_Function_1/NAND4_in[0] ,
         \SB1_1_14/Component_Function_5/NAND4_in[2] ,
         \SB1_1_14/Component_Function_5/NAND4_in[1] ,
         \SB1_1_14/Component_Function_5/NAND4_in[0] ,
         \SB1_1_15/Component_Function_0/NAND4_in[2] ,
         \SB1_1_15/Component_Function_0/NAND4_in[1] ,
         \SB1_1_15/Component_Function_0/NAND4_in[0] ,
         \SB1_1_15/Component_Function_1/NAND4_in[1] ,
         \SB1_1_15/Component_Function_1/NAND4_in[0] ,
         \SB1_1_15/Component_Function_5/NAND4_in[1] ,
         \SB1_1_15/Component_Function_5/NAND4_in[0] ,
         \SB1_1_16/Component_Function_0/NAND4_in[3] ,
         \SB1_1_16/Component_Function_0/NAND4_in[2] ,
         \SB1_1_16/Component_Function_0/NAND4_in[1] ,
         \SB1_1_16/Component_Function_0/NAND4_in[0] ,
         \SB1_1_16/Component_Function_1/NAND4_in[2] ,
         \SB1_1_16/Component_Function_1/NAND4_in[1] ,
         \SB1_1_16/Component_Function_1/NAND4_in[0] ,
         \SB1_1_16/Component_Function_5/NAND4_in[2] ,
         \SB1_1_16/Component_Function_5/NAND4_in[1] ,
         \SB1_1_16/Component_Function_5/NAND4_in[0] ,
         \SB1_1_17/Component_Function_0/NAND4_in[3] ,
         \SB1_1_17/Component_Function_0/NAND4_in[2] ,
         \SB1_1_17/Component_Function_0/NAND4_in[1] ,
         \SB1_1_17/Component_Function_0/NAND4_in[0] ,
         \SB1_1_17/Component_Function_1/NAND4_in[3] ,
         \SB1_1_17/Component_Function_1/NAND4_in[0] ,
         \SB1_1_17/Component_Function_5/NAND4_in[2] ,
         \SB1_1_17/Component_Function_5/NAND4_in[1] ,
         \SB1_1_17/Component_Function_5/NAND4_in[0] ,
         \SB1_1_18/Component_Function_0/NAND4_in[3] ,
         \SB1_1_18/Component_Function_0/NAND4_in[1] ,
         \SB1_1_18/Component_Function_0/NAND4_in[0] ,
         \SB1_1_18/Component_Function_1/NAND4_in[3] ,
         \SB1_1_18/Component_Function_1/NAND4_in[2] ,
         \SB1_1_18/Component_Function_1/NAND4_in[1] ,
         \SB1_1_18/Component_Function_1/NAND4_in[0] ,
         \SB1_1_18/Component_Function_5/NAND4_in[3] ,
         \SB1_1_18/Component_Function_5/NAND4_in[2] ,
         \SB1_1_18/Component_Function_5/NAND4_in[1] ,
         \SB1_1_18/Component_Function_5/NAND4_in[0] ,
         \SB1_1_19/Component_Function_0/NAND4_in[3] ,
         \SB1_1_19/Component_Function_0/NAND4_in[2] ,
         \SB1_1_19/Component_Function_0/NAND4_in[1] ,
         \SB1_1_19/Component_Function_0/NAND4_in[0] ,
         \SB1_1_19/Component_Function_1/NAND4_in[3] ,
         \SB1_1_19/Component_Function_1/NAND4_in[1] ,
         \SB1_1_19/Component_Function_1/NAND4_in[0] ,
         \SB1_1_19/Component_Function_5/NAND4_in[2] ,
         \SB1_1_19/Component_Function_5/NAND4_in[0] ,
         \SB1_1_20/Component_Function_0/NAND4_in[2] ,
         \SB1_1_20/Component_Function_0/NAND4_in[1] ,
         \SB1_1_20/Component_Function_1/NAND4_in[3] ,
         \SB1_1_20/Component_Function_1/NAND4_in[1] ,
         \SB1_1_20/Component_Function_1/NAND4_in[0] ,
         \SB1_1_20/Component_Function_5/NAND4_in[1] ,
         \SB1_1_20/Component_Function_5/NAND4_in[0] ,
         \SB1_1_21/Component_Function_0/NAND4_in[3] ,
         \SB1_1_21/Component_Function_0/NAND4_in[1] ,
         \SB1_1_21/Component_Function_1/NAND4_in[3] ,
         \SB1_1_21/Component_Function_1/NAND4_in[2] ,
         \SB1_1_21/Component_Function_1/NAND4_in[1] ,
         \SB1_1_21/Component_Function_1/NAND4_in[0] ,
         \SB1_1_21/Component_Function_5/NAND4_in[2] ,
         \SB1_1_21/Component_Function_5/NAND4_in[1] ,
         \SB1_1_21/Component_Function_5/NAND4_in[0] ,
         \SB1_1_22/Component_Function_0/NAND4_in[3] ,
         \SB1_1_22/Component_Function_0/NAND4_in[2] ,
         \SB1_1_22/Component_Function_0/NAND4_in[1] ,
         \SB1_1_22/Component_Function_0/NAND4_in[0] ,
         \SB1_1_22/Component_Function_1/NAND4_in[2] ,
         \SB1_1_22/Component_Function_1/NAND4_in[1] ,
         \SB1_1_22/Component_Function_1/NAND4_in[0] ,
         \SB1_1_22/Component_Function_5/NAND4_in[3] ,
         \SB1_1_23/Component_Function_0/NAND4_in[2] ,
         \SB1_1_23/Component_Function_0/NAND4_in[1] ,
         \SB1_1_23/Component_Function_0/NAND4_in[0] ,
         \SB1_1_23/Component_Function_1/NAND4_in[2] ,
         \SB1_1_23/Component_Function_1/NAND4_in[1] ,
         \SB1_1_23/Component_Function_1/NAND4_in[0] ,
         \SB1_1_23/Component_Function_5/NAND4_in[3] ,
         \SB1_1_23/Component_Function_5/NAND4_in[1] ,
         \SB1_1_23/Component_Function_5/NAND4_in[0] ,
         \SB1_1_24/Component_Function_0/NAND4_in[3] ,
         \SB1_1_24/Component_Function_0/NAND4_in[2] ,
         \SB1_1_24/Component_Function_0/NAND4_in[1] ,
         \SB1_1_24/Component_Function_0/NAND4_in[0] ,
         \SB1_1_24/Component_Function_1/NAND4_in[3] ,
         \SB1_1_24/Component_Function_1/NAND4_in[2] ,
         \SB1_1_24/Component_Function_5/NAND4_in[3] ,
         \SB1_1_24/Component_Function_5/NAND4_in[2] ,
         \SB1_1_24/Component_Function_5/NAND4_in[0] ,
         \SB1_1_25/Component_Function_0/NAND4_in[3] ,
         \SB1_1_25/Component_Function_0/NAND4_in[2] ,
         \SB1_1_25/Component_Function_0/NAND4_in[1] ,
         \SB1_1_25/Component_Function_0/NAND4_in[0] ,
         \SB1_1_25/Component_Function_1/NAND4_in[2] ,
         \SB1_1_25/Component_Function_5/NAND4_in[3] ,
         \SB1_1_25/Component_Function_5/NAND4_in[1] ,
         \SB1_1_26/Component_Function_0/NAND4_in[2] ,
         \SB1_1_26/Component_Function_0/NAND4_in[1] ,
         \SB1_1_26/Component_Function_0/NAND4_in[0] ,
         \SB1_1_26/Component_Function_1/NAND4_in[2] ,
         \SB1_1_26/Component_Function_1/NAND4_in[1] ,
         \SB1_1_26/Component_Function_1/NAND4_in[0] ,
         \SB1_1_26/Component_Function_5/NAND4_in[3] ,
         \SB1_1_26/Component_Function_5/NAND4_in[1] ,
         \SB1_1_26/Component_Function_5/NAND4_in[0] ,
         \SB1_1_27/Component_Function_0/NAND4_in[3] ,
         \SB1_1_27/Component_Function_0/NAND4_in[2] ,
         \SB1_1_27/Component_Function_0/NAND4_in[1] ,
         \SB1_1_27/Component_Function_0/NAND4_in[0] ,
         \SB1_1_27/Component_Function_1/NAND4_in[2] ,
         \SB1_1_27/Component_Function_1/NAND4_in[1] ,
         \SB1_1_27/Component_Function_1/NAND4_in[0] ,
         \SB1_1_27/Component_Function_5/NAND4_in[1] ,
         \SB1_1_27/Component_Function_5/NAND4_in[0] ,
         \SB1_1_28/Component_Function_0/NAND4_in[3] ,
         \SB1_1_28/Component_Function_0/NAND4_in[2] ,
         \SB1_1_28/Component_Function_0/NAND4_in[1] ,
         \SB1_1_28/Component_Function_0/NAND4_in[0] ,
         \SB1_1_28/Component_Function_1/NAND4_in[3] ,
         \SB1_1_28/Component_Function_1/NAND4_in[2] ,
         \SB1_1_28/Component_Function_1/NAND4_in[1] ,
         \SB1_1_28/Component_Function_1/NAND4_in[0] ,
         \SB1_1_28/Component_Function_5/NAND4_in[2] ,
         \SB1_1_28/Component_Function_5/NAND4_in[1] ,
         \SB1_1_28/Component_Function_5/NAND4_in[0] ,
         \SB1_1_29/Component_Function_0/NAND4_in[3] ,
         \SB1_1_29/Component_Function_0/NAND4_in[2] ,
         \SB1_1_29/Component_Function_0/NAND4_in[1] ,
         \SB1_1_29/Component_Function_0/NAND4_in[0] ,
         \SB1_1_29/Component_Function_1/NAND4_in[3] ,
         \SB1_1_29/Component_Function_1/NAND4_in[0] ,
         \SB1_1_29/Component_Function_5/NAND4_in[2] ,
         \SB1_1_29/Component_Function_5/NAND4_in[1] ,
         \SB1_1_29/Component_Function_5/NAND4_in[0] ,
         \SB1_1_30/Component_Function_0/NAND4_in[2] ,
         \SB1_1_30/Component_Function_0/NAND4_in[1] ,
         \SB1_1_30/Component_Function_0/NAND4_in[0] ,
         \SB1_1_30/Component_Function_1/NAND4_in[2] ,
         \SB1_1_30/Component_Function_1/NAND4_in[1] ,
         \SB1_1_30/Component_Function_1/NAND4_in[0] ,
         \SB1_1_30/Component_Function_5/NAND4_in[2] ,
         \SB1_1_30/Component_Function_5/NAND4_in[1] ,
         \SB1_1_30/Component_Function_5/NAND4_in[0] ,
         \SB1_1_31/Component_Function_0/NAND4_in[2] ,
         \SB1_1_31/Component_Function_0/NAND4_in[1] ,
         \SB1_1_31/Component_Function_0/NAND4_in[0] ,
         \SB1_1_31/Component_Function_1/NAND4_in[2] ,
         \SB1_1_31/Component_Function_1/NAND4_in[1] ,
         \SB1_1_31/Component_Function_1/NAND4_in[0] ,
         \SB1_1_31/Component_Function_5/NAND4_in[3] ,
         \SB1_1_31/Component_Function_5/NAND4_in[1] ,
         \SB1_1_31/Component_Function_5/NAND4_in[0] ,
         \SB2_1_0/Component_Function_0/NAND4_in[1] ,
         \SB2_1_0/Component_Function_0/NAND4_in[0] ,
         \SB2_1_0/Component_Function_1/NAND4_in[2] ,
         \SB2_1_0/Component_Function_1/NAND4_in[1] ,
         \SB2_1_0/Component_Function_1/NAND4_in[0] ,
         \SB2_1_0/Component_Function_5/NAND4_in[2] ,
         \SB2_1_0/Component_Function_5/NAND4_in[0] ,
         \SB2_1_1/Component_Function_0/NAND4_in[3] ,
         \SB2_1_1/Component_Function_0/NAND4_in[1] ,
         \SB2_1_1/Component_Function_0/NAND4_in[0] ,
         \SB2_1_1/Component_Function_1/NAND4_in[2] ,
         \SB2_1_1/Component_Function_1/NAND4_in[1] ,
         \SB2_1_1/Component_Function_1/NAND4_in[0] ,
         \SB2_1_1/Component_Function_5/NAND4_in[1] ,
         \SB2_1_1/Component_Function_5/NAND4_in[0] ,
         \SB2_1_2/Component_Function_0/NAND4_in[1] ,
         \SB2_1_2/Component_Function_0/NAND4_in[0] ,
         \SB2_1_2/Component_Function_1/NAND4_in[3] ,
         \SB2_1_2/Component_Function_1/NAND4_in[2] ,
         \SB2_1_2/Component_Function_5/NAND4_in[2] ,
         \SB2_1_2/Component_Function_5/NAND4_in[0] ,
         \SB2_1_3/Component_Function_0/NAND4_in[3] ,
         \SB2_1_3/Component_Function_0/NAND4_in[2] ,
         \SB2_1_3/Component_Function_0/NAND4_in[0] ,
         \SB2_1_3/Component_Function_1/NAND4_in[3] ,
         \SB2_1_3/Component_Function_1/NAND4_in[1] ,
         \SB2_1_3/Component_Function_1/NAND4_in[0] ,
         \SB2_1_3/Component_Function_5/NAND4_in[2] ,
         \SB2_1_4/Component_Function_0/NAND4_in[3] ,
         \SB2_1_4/Component_Function_0/NAND4_in[1] ,
         \SB2_1_4/Component_Function_0/NAND4_in[0] ,
         \SB2_1_4/Component_Function_1/NAND4_in[2] ,
         \SB2_1_4/Component_Function_1/NAND4_in[1] ,
         \SB2_1_4/Component_Function_1/NAND4_in[0] ,
         \SB2_1_4/Component_Function_5/NAND4_in[2] ,
         \SB2_1_4/Component_Function_5/NAND4_in[0] ,
         \SB2_1_5/Component_Function_0/NAND4_in[3] ,
         \SB2_1_5/Component_Function_0/NAND4_in[0] ,
         \SB2_1_5/Component_Function_1/NAND4_in[3] ,
         \SB2_1_5/Component_Function_1/NAND4_in[2] ,
         \SB2_1_5/Component_Function_1/NAND4_in[1] ,
         \SB2_1_5/Component_Function_5/NAND4_in[3] ,
         \SB2_1_5/Component_Function_5/NAND4_in[2] ,
         \SB2_1_6/Component_Function_0/NAND4_in[3] ,
         \SB2_1_6/Component_Function_0/NAND4_in[1] ,
         \SB2_1_6/Component_Function_0/NAND4_in[0] ,
         \SB2_1_6/Component_Function_1/NAND4_in[3] ,
         \SB2_1_6/Component_Function_1/NAND4_in[1] ,
         \SB2_1_6/Component_Function_1/NAND4_in[0] ,
         \SB2_1_6/Component_Function_5/NAND4_in[1] ,
         \SB2_1_6/Component_Function_5/NAND4_in[0] ,
         \SB2_1_7/Component_Function_0/NAND4_in[3] ,
         \SB2_1_7/Component_Function_0/NAND4_in[2] ,
         \SB2_1_7/Component_Function_0/NAND4_in[1] ,
         \SB2_1_7/Component_Function_0/NAND4_in[0] ,
         \SB2_1_7/Component_Function_1/NAND4_in[2] ,
         \SB2_1_7/Component_Function_1/NAND4_in[1] ,
         \SB2_1_7/Component_Function_1/NAND4_in[0] ,
         \SB2_1_7/Component_Function_5/NAND4_in[2] ,
         \SB2_1_7/Component_Function_5/NAND4_in[0] ,
         \SB2_1_8/Component_Function_0/NAND4_in[3] ,
         \SB2_1_8/Component_Function_0/NAND4_in[1] ,
         \SB2_1_8/Component_Function_1/NAND4_in[2] ,
         \SB2_1_8/Component_Function_1/NAND4_in[1] ,
         \SB2_1_8/Component_Function_1/NAND4_in[0] ,
         \SB2_1_8/Component_Function_5/NAND4_in[2] ,
         \SB2_1_8/Component_Function_5/NAND4_in[0] ,
         \SB2_1_9/Component_Function_0/NAND4_in[3] ,
         \SB2_1_9/Component_Function_0/NAND4_in[2] ,
         \SB2_1_9/Component_Function_0/NAND4_in[1] ,
         \SB2_1_9/Component_Function_1/NAND4_in[3] ,
         \SB2_1_9/Component_Function_1/NAND4_in[2] ,
         \SB2_1_9/Component_Function_5/NAND4_in[1] ,
         \SB2_1_9/Component_Function_5/NAND4_in[0] ,
         \SB2_1_10/Component_Function_0/NAND4_in[3] ,
         \SB2_1_10/Component_Function_0/NAND4_in[1] ,
         \SB2_1_10/Component_Function_1/NAND4_in[3] ,
         \SB2_1_10/Component_Function_1/NAND4_in[2] ,
         \SB2_1_10/Component_Function_1/NAND4_in[1] ,
         \SB2_1_10/Component_Function_1/NAND4_in[0] ,
         \SB2_1_10/Component_Function_5/NAND4_in[3] ,
         \SB2_1_11/Component_Function_0/NAND4_in[2] ,
         \SB2_1_11/Component_Function_0/NAND4_in[1] ,
         \SB2_1_11/Component_Function_0/NAND4_in[0] ,
         \SB2_1_11/Component_Function_1/NAND4_in[3] ,
         \SB2_1_11/Component_Function_1/NAND4_in[2] ,
         \SB2_1_11/Component_Function_1/NAND4_in[1] ,
         \SB2_1_11/Component_Function_1/NAND4_in[0] ,
         \SB2_1_11/Component_Function_5/NAND4_in[2] ,
         \SB2_1_11/Component_Function_5/NAND4_in[0] ,
         \SB2_1_12/Component_Function_0/NAND4_in[3] ,
         \SB2_1_12/Component_Function_0/NAND4_in[1] ,
         \SB2_1_12/Component_Function_0/NAND4_in[0] ,
         \SB2_1_12/Component_Function_1/NAND4_in[2] ,
         \SB2_1_12/Component_Function_1/NAND4_in[1] ,
         \SB2_1_12/Component_Function_1/NAND4_in[0] ,
         \SB2_1_12/Component_Function_5/NAND4_in[2] ,
         \SB2_1_12/Component_Function_5/NAND4_in[1] ,
         \SB2_1_12/Component_Function_5/NAND4_in[0] ,
         \SB2_1_13/Component_Function_0/NAND4_in[1] ,
         \SB2_1_13/Component_Function_0/NAND4_in[0] ,
         \SB2_1_13/Component_Function_1/NAND4_in[2] ,
         \SB2_1_13/Component_Function_1/NAND4_in[1] ,
         \SB2_1_13/Component_Function_1/NAND4_in[0] ,
         \SB2_1_13/Component_Function_5/NAND4_in[3] ,
         \SB2_1_13/Component_Function_5/NAND4_in[1] ,
         \SB2_1_13/Component_Function_5/NAND4_in[0] ,
         \SB2_1_14/Component_Function_0/NAND4_in[2] ,
         \SB2_1_14/Component_Function_0/NAND4_in[1] ,
         \SB2_1_14/Component_Function_0/NAND4_in[0] ,
         \SB2_1_14/Component_Function_1/NAND4_in[3] ,
         \SB2_1_14/Component_Function_1/NAND4_in[2] ,
         \SB2_1_14/Component_Function_1/NAND4_in[1] ,
         \SB2_1_14/Component_Function_1/NAND4_in[0] ,
         \SB2_1_14/Component_Function_5/NAND4_in[2] ,
         \SB2_1_14/Component_Function_5/NAND4_in[1] ,
         \SB2_1_14/Component_Function_5/NAND4_in[0] ,
         \SB2_1_15/Component_Function_0/NAND4_in[3] ,
         \SB2_1_15/Component_Function_0/NAND4_in[2] ,
         \SB2_1_15/Component_Function_0/NAND4_in[1] ,
         \SB2_1_15/Component_Function_0/NAND4_in[0] ,
         \SB2_1_15/Component_Function_1/NAND4_in[3] ,
         \SB2_1_15/Component_Function_1/NAND4_in[2] ,
         \SB2_1_15/Component_Function_1/NAND4_in[1] ,
         \SB2_1_15/Component_Function_1/NAND4_in[0] ,
         \SB2_1_15/Component_Function_5/NAND4_in[1] ,
         \SB2_1_15/Component_Function_5/NAND4_in[0] ,
         \SB2_1_16/Component_Function_0/NAND4_in[3] ,
         \SB2_1_16/Component_Function_0/NAND4_in[2] ,
         \SB2_1_16/Component_Function_0/NAND4_in[1] ,
         \SB2_1_16/Component_Function_0/NAND4_in[0] ,
         \SB2_1_16/Component_Function_1/NAND4_in[2] ,
         \SB2_1_16/Component_Function_1/NAND4_in[1] ,
         \SB2_1_16/Component_Function_1/NAND4_in[0] ,
         \SB2_1_16/Component_Function_5/NAND4_in[1] ,
         \SB2_1_16/Component_Function_5/NAND4_in[0] ,
         \SB2_1_17/Component_Function_0/NAND4_in[3] ,
         \SB2_1_17/Component_Function_0/NAND4_in[2] ,
         \SB2_1_17/Component_Function_0/NAND4_in[1] ,
         \SB2_1_17/Component_Function_1/NAND4_in[3] ,
         \SB2_1_17/Component_Function_1/NAND4_in[1] ,
         \SB2_1_17/Component_Function_1/NAND4_in[0] ,
         \SB2_1_17/Component_Function_5/NAND4_in[0] ,
         \SB2_1_18/Component_Function_0/NAND4_in[2] ,
         \SB2_1_18/Component_Function_0/NAND4_in[1] ,
         \SB2_1_18/Component_Function_0/NAND4_in[0] ,
         \SB2_1_18/Component_Function_1/NAND4_in[3] ,
         \SB2_1_18/Component_Function_1/NAND4_in[2] ,
         \SB2_1_18/Component_Function_1/NAND4_in[1] ,
         \SB2_1_18/Component_Function_1/NAND4_in[0] ,
         \SB2_1_18/Component_Function_5/NAND4_in[2] ,
         \SB2_1_18/Component_Function_5/NAND4_in[0] ,
         \SB2_1_19/Component_Function_0/NAND4_in[3] ,
         \SB2_1_19/Component_Function_0/NAND4_in[2] ,
         \SB2_1_19/Component_Function_0/NAND4_in[1] ,
         \SB2_1_19/Component_Function_0/NAND4_in[0] ,
         \SB2_1_19/Component_Function_1/NAND4_in[3] ,
         \SB2_1_19/Component_Function_1/NAND4_in[1] ,
         \SB2_1_19/Component_Function_1/NAND4_in[0] ,
         \SB2_1_19/Component_Function_5/NAND4_in[2] ,
         \SB2_1_19/Component_Function_5/NAND4_in[1] ,
         \SB2_1_19/Component_Function_5/NAND4_in[0] ,
         \SB2_1_20/Component_Function_0/NAND4_in[3] ,
         \SB2_1_20/Component_Function_0/NAND4_in[1] ,
         \SB2_1_20/Component_Function_0/NAND4_in[0] ,
         \SB2_1_20/Component_Function_1/NAND4_in[2] ,
         \SB2_1_20/Component_Function_1/NAND4_in[1] ,
         \SB2_1_20/Component_Function_1/NAND4_in[0] ,
         \SB2_1_20/Component_Function_5/NAND4_in[1] ,
         \SB2_1_20/Component_Function_5/NAND4_in[0] ,
         \SB2_1_21/Component_Function_0/NAND4_in[3] ,
         \SB2_1_21/Component_Function_0/NAND4_in[1] ,
         \SB2_1_21/Component_Function_1/NAND4_in[3] ,
         \SB2_1_21/Component_Function_1/NAND4_in[1] ,
         \SB2_1_21/Component_Function_1/NAND4_in[0] ,
         \SB2_1_21/Component_Function_5/NAND4_in[2] ,
         \SB2_1_21/Component_Function_5/NAND4_in[0] ,
         \SB2_1_22/Component_Function_0/NAND4_in[3] ,
         \SB2_1_22/Component_Function_0/NAND4_in[1] ,
         \SB2_1_22/Component_Function_0/NAND4_in[0] ,
         \SB2_1_22/Component_Function_1/NAND4_in[3] ,
         \SB2_1_22/Component_Function_1/NAND4_in[2] ,
         \SB2_1_22/Component_Function_1/NAND4_in[1] ,
         \SB2_1_22/Component_Function_1/NAND4_in[0] ,
         \SB2_1_22/Component_Function_5/NAND4_in[3] ,
         \SB2_1_22/Component_Function_5/NAND4_in[0] ,
         \SB2_1_23/Component_Function_0/NAND4_in[3] ,
         \SB2_1_23/Component_Function_0/NAND4_in[2] ,
         \SB2_1_23/Component_Function_0/NAND4_in[1] ,
         \SB2_1_23/Component_Function_0/NAND4_in[0] ,
         \SB2_1_23/Component_Function_1/NAND4_in[3] ,
         \SB2_1_23/Component_Function_1/NAND4_in[2] ,
         \SB2_1_23/Component_Function_1/NAND4_in[1] ,
         \SB2_1_23/Component_Function_1/NAND4_in[0] ,
         \SB2_1_23/Component_Function_5/NAND4_in[0] ,
         \SB2_1_24/Component_Function_0/NAND4_in[2] ,
         \SB2_1_24/Component_Function_0/NAND4_in[1] ,
         \SB2_1_24/Component_Function_0/NAND4_in[0] ,
         \SB2_1_24/Component_Function_1/NAND4_in[3] ,
         \SB2_1_24/Component_Function_1/NAND4_in[2] ,
         \SB2_1_24/Component_Function_1/NAND4_in[1] ,
         \SB2_1_24/Component_Function_1/NAND4_in[0] ,
         \SB2_1_24/Component_Function_5/NAND4_in[3] ,
         \SB2_1_24/Component_Function_5/NAND4_in[2] ,
         \SB2_1_24/Component_Function_5/NAND4_in[1] ,
         \SB2_1_24/Component_Function_5/NAND4_in[0] ,
         \SB2_1_25/Component_Function_0/NAND4_in[2] ,
         \SB2_1_25/Component_Function_0/NAND4_in[0] ,
         \SB2_1_25/Component_Function_1/NAND4_in[3] ,
         \SB2_1_25/Component_Function_1/NAND4_in[1] ,
         \SB2_1_25/Component_Function_1/NAND4_in[0] ,
         \SB2_1_25/Component_Function_5/NAND4_in[3] ,
         \SB2_1_25/Component_Function_5/NAND4_in[0] ,
         \SB2_1_26/Component_Function_0/NAND4_in[1] ,
         \SB2_1_26/Component_Function_0/NAND4_in[0] ,
         \SB2_1_26/Component_Function_1/NAND4_in[3] ,
         \SB2_1_26/Component_Function_1/NAND4_in[1] ,
         \SB2_1_26/Component_Function_1/NAND4_in[0] ,
         \SB2_1_26/Component_Function_5/NAND4_in[3] ,
         \SB2_1_26/Component_Function_5/NAND4_in[1] ,
         \SB2_1_27/Component_Function_0/NAND4_in[3] ,
         \SB2_1_27/Component_Function_0/NAND4_in[2] ,
         \SB2_1_27/Component_Function_0/NAND4_in[1] ,
         \SB2_1_27/Component_Function_0/NAND4_in[0] ,
         \SB2_1_27/Component_Function_1/NAND4_in[2] ,
         \SB2_1_27/Component_Function_1/NAND4_in[1] ,
         \SB2_1_27/Component_Function_1/NAND4_in[0] ,
         \SB2_1_27/Component_Function_5/NAND4_in[3] ,
         \SB2_1_27/Component_Function_5/NAND4_in[0] ,
         \SB2_1_28/Component_Function_0/NAND4_in[1] ,
         \SB2_1_28/Component_Function_0/NAND4_in[0] ,
         \SB2_1_28/Component_Function_1/NAND4_in[2] ,
         \SB2_1_28/Component_Function_1/NAND4_in[1] ,
         \SB2_1_28/Component_Function_1/NAND4_in[0] ,
         \SB2_1_28/Component_Function_5/NAND4_in[3] ,
         \SB2_1_28/Component_Function_5/NAND4_in[2] ,
         \SB2_1_28/Component_Function_5/NAND4_in[1] ,
         \SB2_1_28/Component_Function_5/NAND4_in[0] ,
         \SB2_1_29/Component_Function_0/NAND4_in[3] ,
         \SB2_1_29/Component_Function_0/NAND4_in[2] ,
         \SB2_1_29/Component_Function_0/NAND4_in[0] ,
         \SB2_1_29/Component_Function_1/NAND4_in[3] ,
         \SB2_1_29/Component_Function_1/NAND4_in[1] ,
         \SB2_1_29/Component_Function_1/NAND4_in[0] ,
         \SB2_1_29/Component_Function_5/NAND4_in[3] ,
         \SB2_1_29/Component_Function_5/NAND4_in[1] ,
         \SB2_1_29/Component_Function_5/NAND4_in[0] ,
         \SB2_1_30/Component_Function_0/NAND4_in[3] ,
         \SB2_1_30/Component_Function_0/NAND4_in[2] ,
         \SB2_1_30/Component_Function_0/NAND4_in[1] ,
         \SB2_1_30/Component_Function_0/NAND4_in[0] ,
         \SB2_1_30/Component_Function_1/NAND4_in[2] ,
         \SB2_1_30/Component_Function_1/NAND4_in[1] ,
         \SB2_1_30/Component_Function_1/NAND4_in[0] ,
         \SB2_1_30/Component_Function_5/NAND4_in[3] ,
         \SB2_1_30/Component_Function_5/NAND4_in[2] ,
         \SB2_1_30/Component_Function_5/NAND4_in[1] ,
         \SB2_1_30/Component_Function_5/NAND4_in[0] ,
         \SB2_1_31/Component_Function_0/NAND4_in[3] ,
         \SB2_1_31/Component_Function_0/NAND4_in[2] ,
         \SB2_1_31/Component_Function_0/NAND4_in[1] ,
         \SB2_1_31/Component_Function_0/NAND4_in[0] ,
         \SB2_1_31/Component_Function_1/NAND4_in[3] ,
         \SB2_1_31/Component_Function_1/NAND4_in[2] ,
         \SB2_1_31/Component_Function_1/NAND4_in[1] ,
         \SB2_1_31/Component_Function_1/NAND4_in[0] ,
         \SB2_1_31/Component_Function_5/NAND4_in[3] ,
         \SB2_1_31/Component_Function_5/NAND4_in[1] ,
         \SB2_1_31/Component_Function_5/NAND4_in[0] ,
         \SB1_2_0/Component_Function_0/NAND4_in[2] ,
         \SB1_2_0/Component_Function_0/NAND4_in[1] ,
         \SB1_2_0/Component_Function_0/NAND4_in[0] ,
         \SB1_2_0/Component_Function_1/NAND4_in[3] ,
         \SB1_2_0/Component_Function_1/NAND4_in[2] ,
         \SB1_2_0/Component_Function_1/NAND4_in[1] ,
         \SB1_2_0/Component_Function_1/NAND4_in[0] ,
         \SB1_2_0/Component_Function_5/NAND4_in[2] ,
         \SB1_2_0/Component_Function_5/NAND4_in[1] ,
         \SB1_2_0/Component_Function_5/NAND4_in[0] ,
         \SB1_2_1/Component_Function_0/NAND4_in[3] ,
         \SB1_2_1/Component_Function_0/NAND4_in[2] ,
         \SB1_2_1/Component_Function_0/NAND4_in[1] ,
         \SB1_2_1/Component_Function_0/NAND4_in[0] ,
         \SB1_2_1/Component_Function_1/NAND4_in[3] ,
         \SB1_2_1/Component_Function_1/NAND4_in[1] ,
         \SB1_2_1/Component_Function_1/NAND4_in[0] ,
         \SB1_2_1/Component_Function_5/NAND4_in[2] ,
         \SB1_2_1/Component_Function_5/NAND4_in[1] ,
         \SB1_2_1/Component_Function_5/NAND4_in[0] ,
         \SB1_2_2/Component_Function_0/NAND4_in[2] ,
         \SB1_2_2/Component_Function_0/NAND4_in[1] ,
         \SB1_2_2/Component_Function_0/NAND4_in[0] ,
         \SB1_2_2/Component_Function_1/NAND4_in[2] ,
         \SB1_2_2/Component_Function_1/NAND4_in[1] ,
         \SB1_2_2/Component_Function_1/NAND4_in[0] ,
         \SB1_2_2/Component_Function_5/NAND4_in[2] ,
         \SB1_2_2/Component_Function_5/NAND4_in[1] ,
         \SB1_2_2/Component_Function_5/NAND4_in[0] ,
         \SB1_2_3/Component_Function_0/NAND4_in[3] ,
         \SB1_2_3/Component_Function_0/NAND4_in[2] ,
         \SB1_2_3/Component_Function_0/NAND4_in[1] ,
         \SB1_2_3/Component_Function_0/NAND4_in[0] ,
         \SB1_2_3/Component_Function_1/NAND4_in[1] ,
         \SB1_2_3/Component_Function_1/NAND4_in[0] ,
         \SB1_2_3/Component_Function_5/NAND4_in[2] ,
         \SB1_2_4/Component_Function_0/NAND4_in[3] ,
         \SB1_2_4/Component_Function_0/NAND4_in[2] ,
         \SB1_2_4/Component_Function_0/NAND4_in[1] ,
         \SB1_2_4/Component_Function_0/NAND4_in[0] ,
         \SB1_2_4/Component_Function_1/NAND4_in[3] ,
         \SB1_2_4/Component_Function_1/NAND4_in[1] ,
         \SB1_2_4/Component_Function_1/NAND4_in[0] ,
         \SB1_2_4/Component_Function_5/NAND4_in[2] ,
         \SB1_2_4/Component_Function_5/NAND4_in[1] ,
         \SB1_2_4/Component_Function_5/NAND4_in[0] ,
         \SB1_2_5/Component_Function_0/NAND4_in[3] ,
         \SB1_2_5/Component_Function_0/NAND4_in[2] ,
         \SB1_2_5/Component_Function_0/NAND4_in[1] ,
         \SB1_2_5/Component_Function_0/NAND4_in[0] ,
         \SB1_2_5/Component_Function_1/NAND4_in[3] ,
         \SB1_2_5/Component_Function_1/NAND4_in[1] ,
         \SB1_2_5/Component_Function_1/NAND4_in[0] ,
         \SB1_2_5/Component_Function_5/NAND4_in[2] ,
         \SB1_2_5/Component_Function_5/NAND4_in[1] ,
         \SB1_2_5/Component_Function_5/NAND4_in[0] ,
         \SB1_2_6/Component_Function_0/NAND4_in[2] ,
         \SB1_2_6/Component_Function_0/NAND4_in[1] ,
         \SB1_2_6/Component_Function_0/NAND4_in[0] ,
         \SB1_2_6/Component_Function_1/NAND4_in[2] ,
         \SB1_2_6/Component_Function_1/NAND4_in[1] ,
         \SB1_2_6/Component_Function_1/NAND4_in[0] ,
         \SB1_2_6/Component_Function_5/NAND4_in[1] ,
         \SB1_2_6/Component_Function_5/NAND4_in[0] ,
         \SB1_2_7/Component_Function_0/NAND4_in[3] ,
         \SB1_2_7/Component_Function_0/NAND4_in[2] ,
         \SB1_2_7/Component_Function_0/NAND4_in[1] ,
         \SB1_2_7/Component_Function_0/NAND4_in[0] ,
         \SB1_2_7/Component_Function_1/NAND4_in[2] ,
         \SB1_2_7/Component_Function_1/NAND4_in[1] ,
         \SB1_2_7/Component_Function_1/NAND4_in[0] ,
         \SB1_2_7/Component_Function_5/NAND4_in[2] ,
         \SB1_2_7/Component_Function_5/NAND4_in[1] ,
         \SB1_2_8/Component_Function_0/NAND4_in[2] ,
         \SB1_2_8/Component_Function_0/NAND4_in[1] ,
         \SB1_2_8/Component_Function_0/NAND4_in[0] ,
         \SB1_2_8/Component_Function_1/NAND4_in[3] ,
         \SB1_2_8/Component_Function_1/NAND4_in[0] ,
         \SB1_2_8/Component_Function_5/NAND4_in[1] ,
         \SB1_2_8/Component_Function_5/NAND4_in[0] ,
         \SB1_2_9/Component_Function_0/NAND4_in[2] ,
         \SB1_2_9/Component_Function_0/NAND4_in[1] ,
         \SB1_2_9/Component_Function_0/NAND4_in[0] ,
         \SB1_2_9/Component_Function_1/NAND4_in[1] ,
         \SB1_2_9/Component_Function_1/NAND4_in[0] ,
         \SB1_2_9/Component_Function_5/NAND4_in[2] ,
         \SB1_2_9/Component_Function_5/NAND4_in[1] ,
         \SB1_2_9/Component_Function_5/NAND4_in[0] ,
         \SB1_2_10/Component_Function_0/NAND4_in[2] ,
         \SB1_2_10/Component_Function_0/NAND4_in[1] ,
         \SB1_2_10/Component_Function_0/NAND4_in[0] ,
         \SB1_2_10/Component_Function_1/NAND4_in[3] ,
         \SB1_2_10/Component_Function_1/NAND4_in[1] ,
         \SB1_2_10/Component_Function_1/NAND4_in[0] ,
         \SB1_2_10/Component_Function_5/NAND4_in[3] ,
         \SB1_2_10/Component_Function_5/NAND4_in[1] ,
         \SB1_2_11/Component_Function_0/NAND4_in[2] ,
         \SB1_2_11/Component_Function_0/NAND4_in[0] ,
         \SB1_2_11/Component_Function_1/NAND4_in[3] ,
         \SB1_2_11/Component_Function_1/NAND4_in[2] ,
         \SB1_2_11/Component_Function_1/NAND4_in[1] ,
         \SB1_2_11/Component_Function_1/NAND4_in[0] ,
         \SB1_2_11/Component_Function_5/NAND4_in[3] ,
         \SB1_2_11/Component_Function_5/NAND4_in[0] ,
         \SB1_2_12/Component_Function_0/NAND4_in[3] ,
         \SB1_2_12/Component_Function_0/NAND4_in[1] ,
         \SB1_2_12/Component_Function_0/NAND4_in[0] ,
         \SB1_2_12/Component_Function_1/NAND4_in[3] ,
         \SB1_2_12/Component_Function_1/NAND4_in[1] ,
         \SB1_2_12/Component_Function_1/NAND4_in[0] ,
         \SB1_2_12/Component_Function_5/NAND4_in[2] ,
         \SB1_2_12/Component_Function_5/NAND4_in[1] ,
         \SB1_2_12/Component_Function_5/NAND4_in[0] ,
         \SB1_2_13/Component_Function_0/NAND4_in[3] ,
         \SB1_2_13/Component_Function_0/NAND4_in[2] ,
         \SB1_2_13/Component_Function_0/NAND4_in[1] ,
         \SB1_2_13/Component_Function_0/NAND4_in[0] ,
         \SB1_2_13/Component_Function_1/NAND4_in[3] ,
         \SB1_2_13/Component_Function_1/NAND4_in[2] ,
         \SB1_2_13/Component_Function_1/NAND4_in[1] ,
         \SB1_2_13/Component_Function_1/NAND4_in[0] ,
         \SB1_2_13/Component_Function_5/NAND4_in[3] ,
         \SB1_2_13/Component_Function_5/NAND4_in[2] ,
         \SB1_2_13/Component_Function_5/NAND4_in[0] ,
         \SB1_2_14/Component_Function_0/NAND4_in[2] ,
         \SB1_2_14/Component_Function_0/NAND4_in[1] ,
         \SB1_2_14/Component_Function_0/NAND4_in[0] ,
         \SB1_2_14/Component_Function_1/NAND4_in[2] ,
         \SB1_2_14/Component_Function_1/NAND4_in[1] ,
         \SB1_2_14/Component_Function_1/NAND4_in[0] ,
         \SB1_2_14/Component_Function_5/NAND4_in[1] ,
         \SB1_2_14/Component_Function_5/NAND4_in[0] ,
         \SB1_2_15/Component_Function_0/NAND4_in[3] ,
         \SB1_2_15/Component_Function_0/NAND4_in[2] ,
         \SB1_2_15/Component_Function_0/NAND4_in[1] ,
         \SB1_2_15/Component_Function_0/NAND4_in[0] ,
         \SB1_2_15/Component_Function_1/NAND4_in[3] ,
         \SB1_2_15/Component_Function_1/NAND4_in[2] ,
         \SB1_2_15/Component_Function_1/NAND4_in[1] ,
         \SB1_2_15/Component_Function_1/NAND4_in[0] ,
         \SB1_2_15/Component_Function_5/NAND4_in[0] ,
         \SB1_2_16/Component_Function_0/NAND4_in[3] ,
         \SB1_2_16/Component_Function_0/NAND4_in[2] ,
         \SB1_2_16/Component_Function_0/NAND4_in[0] ,
         \SB1_2_16/Component_Function_1/NAND4_in[2] ,
         \SB1_2_16/Component_Function_1/NAND4_in[1] ,
         \SB1_2_16/Component_Function_5/NAND4_in[2] ,
         \SB1_2_16/Component_Function_5/NAND4_in[1] ,
         \SB1_2_16/Component_Function_5/NAND4_in[0] ,
         \SB1_2_17/Component_Function_0/NAND4_in[3] ,
         \SB1_2_17/Component_Function_0/NAND4_in[2] ,
         \SB1_2_17/Component_Function_0/NAND4_in[1] ,
         \SB1_2_17/Component_Function_0/NAND4_in[0] ,
         \SB1_2_17/Component_Function_1/NAND4_in[2] ,
         \SB1_2_17/Component_Function_1/NAND4_in[1] ,
         \SB1_2_17/Component_Function_1/NAND4_in[0] ,
         \SB1_2_17/Component_Function_5/NAND4_in[2] ,
         \SB1_2_17/Component_Function_5/NAND4_in[1] ,
         \SB1_2_17/Component_Function_5/NAND4_in[0] ,
         \SB1_2_18/Component_Function_0/NAND4_in[2] ,
         \SB1_2_18/Component_Function_0/NAND4_in[1] ,
         \SB1_2_18/Component_Function_0/NAND4_in[0] ,
         \SB1_2_18/Component_Function_1/NAND4_in[3] ,
         \SB1_2_18/Component_Function_1/NAND4_in[2] ,
         \SB1_2_18/Component_Function_1/NAND4_in[1] ,
         \SB1_2_18/Component_Function_1/NAND4_in[0] ,
         \SB1_2_18/Component_Function_5/NAND4_in[3] ,
         \SB1_2_18/Component_Function_5/NAND4_in[1] ,
         \SB1_2_18/Component_Function_5/NAND4_in[0] ,
         \SB1_2_19/Component_Function_0/NAND4_in[3] ,
         \SB1_2_19/Component_Function_0/NAND4_in[2] ,
         \SB1_2_19/Component_Function_0/NAND4_in[1] ,
         \SB1_2_19/Component_Function_0/NAND4_in[0] ,
         \SB1_2_19/Component_Function_1/NAND4_in[2] ,
         \SB1_2_19/Component_Function_1/NAND4_in[1] ,
         \SB1_2_19/Component_Function_1/NAND4_in[0] ,
         \SB1_2_19/Component_Function_5/NAND4_in[3] ,
         \SB1_2_19/Component_Function_5/NAND4_in[1] ,
         \SB1_2_19/Component_Function_5/NAND4_in[0] ,
         \SB1_2_20/Component_Function_0/NAND4_in[3] ,
         \SB1_2_20/Component_Function_0/NAND4_in[2] ,
         \SB1_2_20/Component_Function_0/NAND4_in[1] ,
         \SB1_2_20/Component_Function_0/NAND4_in[0] ,
         \SB1_2_20/Component_Function_1/NAND4_in[3] ,
         \SB1_2_20/Component_Function_1/NAND4_in[1] ,
         \SB1_2_20/Component_Function_1/NAND4_in[0] ,
         \SB1_2_20/Component_Function_5/NAND4_in[2] ,
         \SB1_2_20/Component_Function_5/NAND4_in[1] ,
         \SB1_2_20/Component_Function_5/NAND4_in[0] ,
         \SB1_2_21/Component_Function_0/NAND4_in[2] ,
         \SB1_2_21/Component_Function_0/NAND4_in[1] ,
         \SB1_2_21/Component_Function_0/NAND4_in[0] ,
         \SB1_2_21/Component_Function_1/NAND4_in[2] ,
         \SB1_2_21/Component_Function_1/NAND4_in[1] ,
         \SB1_2_21/Component_Function_1/NAND4_in[0] ,
         \SB1_2_21/Component_Function_5/NAND4_in[1] ,
         \SB1_2_21/Component_Function_5/NAND4_in[0] ,
         \SB1_2_22/Component_Function_0/NAND4_in[3] ,
         \SB1_2_22/Component_Function_0/NAND4_in[2] ,
         \SB1_2_22/Component_Function_0/NAND4_in[1] ,
         \SB1_2_22/Component_Function_0/NAND4_in[0] ,
         \SB1_2_22/Component_Function_1/NAND4_in[3] ,
         \SB1_2_22/Component_Function_1/NAND4_in[2] ,
         \SB1_2_22/Component_Function_1/NAND4_in[1] ,
         \SB1_2_22/Component_Function_1/NAND4_in[0] ,
         \SB1_2_22/Component_Function_5/NAND4_in[2] ,
         \SB1_2_22/Component_Function_5/NAND4_in[1] ,
         \SB1_2_22/Component_Function_5/NAND4_in[0] ,
         \SB1_2_23/Component_Function_0/NAND4_in[3] ,
         \SB1_2_23/Component_Function_0/NAND4_in[2] ,
         \SB1_2_23/Component_Function_0/NAND4_in[1] ,
         \SB1_2_23/Component_Function_0/NAND4_in[0] ,
         \SB1_2_23/Component_Function_1/NAND4_in[3] ,
         \SB1_2_23/Component_Function_1/NAND4_in[2] ,
         \SB1_2_23/Component_Function_1/NAND4_in[1] ,
         \SB1_2_23/Component_Function_5/NAND4_in[3] ,
         \SB1_2_23/Component_Function_5/NAND4_in[2] ,
         \SB1_2_23/Component_Function_5/NAND4_in[1] ,
         \SB1_2_23/Component_Function_5/NAND4_in[0] ,
         \SB1_2_24/Component_Function_0/NAND4_in[2] ,
         \SB1_2_24/Component_Function_0/NAND4_in[1] ,
         \SB1_2_24/Component_Function_0/NAND4_in[0] ,
         \SB1_2_24/Component_Function_1/NAND4_in[3] ,
         \SB1_2_24/Component_Function_1/NAND4_in[2] ,
         \SB1_2_24/Component_Function_1/NAND4_in[1] ,
         \SB1_2_24/Component_Function_1/NAND4_in[0] ,
         \SB1_2_24/Component_Function_5/NAND4_in[2] ,
         \SB1_2_24/Component_Function_5/NAND4_in[0] ,
         \SB1_2_25/Component_Function_0/NAND4_in[2] ,
         \SB1_2_25/Component_Function_0/NAND4_in[1] ,
         \SB1_2_25/Component_Function_0/NAND4_in[0] ,
         \SB1_2_25/Component_Function_1/NAND4_in[2] ,
         \SB1_2_25/Component_Function_1/NAND4_in[1] ,
         \SB1_2_25/Component_Function_1/NAND4_in[0] ,
         \SB1_2_25/Component_Function_5/NAND4_in[2] ,
         \SB1_2_25/Component_Function_5/NAND4_in[1] ,
         \SB1_2_25/Component_Function_5/NAND4_in[0] ,
         \SB1_2_26/Component_Function_0/NAND4_in[3] ,
         \SB1_2_26/Component_Function_0/NAND4_in[2] ,
         \SB1_2_26/Component_Function_0/NAND4_in[1] ,
         \SB1_2_26/Component_Function_0/NAND4_in[0] ,
         \SB1_2_26/Component_Function_1/NAND4_in[2] ,
         \SB1_2_26/Component_Function_1/NAND4_in[1] ,
         \SB1_2_26/Component_Function_1/NAND4_in[0] ,
         \SB1_2_26/Component_Function_5/NAND4_in[1] ,
         \SB1_2_26/Component_Function_5/NAND4_in[0] ,
         \SB1_2_27/Component_Function_0/NAND4_in[3] ,
         \SB1_2_27/Component_Function_0/NAND4_in[2] ,
         \SB1_2_27/Component_Function_0/NAND4_in[1] ,
         \SB1_2_27/Component_Function_0/NAND4_in[0] ,
         \SB1_2_27/Component_Function_1/NAND4_in[3] ,
         \SB1_2_27/Component_Function_1/NAND4_in[2] ,
         \SB1_2_27/Component_Function_1/NAND4_in[1] ,
         \SB1_2_27/Component_Function_1/NAND4_in[0] ,
         \SB1_2_27/Component_Function_5/NAND4_in[0] ,
         \SB1_2_28/Component_Function_0/NAND4_in[3] ,
         \SB1_2_28/Component_Function_0/NAND4_in[2] ,
         \SB1_2_28/Component_Function_0/NAND4_in[1] ,
         \SB1_2_28/Component_Function_0/NAND4_in[0] ,
         \SB1_2_28/Component_Function_1/NAND4_in[3] ,
         \SB1_2_28/Component_Function_1/NAND4_in[2] ,
         \SB1_2_28/Component_Function_1/NAND4_in[1] ,
         \SB1_2_28/Component_Function_1/NAND4_in[0] ,
         \SB1_2_28/Component_Function_5/NAND4_in[1] ,
         \SB1_2_28/Component_Function_5/NAND4_in[0] ,
         \SB1_2_29/Component_Function_0/NAND4_in[2] ,
         \SB1_2_29/Component_Function_0/NAND4_in[1] ,
         \SB1_2_29/Component_Function_0/NAND4_in[0] ,
         \SB1_2_29/Component_Function_1/NAND4_in[2] ,
         \SB1_2_29/Component_Function_1/NAND4_in[1] ,
         \SB1_2_29/Component_Function_1/NAND4_in[0] ,
         \SB1_2_29/Component_Function_5/NAND4_in[2] ,
         \SB1_2_29/Component_Function_5/NAND4_in[1] ,
         \SB1_2_29/Component_Function_5/NAND4_in[0] ,
         \SB1_2_30/Component_Function_0/NAND4_in[2] ,
         \SB1_2_30/Component_Function_0/NAND4_in[1] ,
         \SB1_2_30/Component_Function_0/NAND4_in[0] ,
         \SB1_2_30/Component_Function_1/NAND4_in[3] ,
         \SB1_2_30/Component_Function_1/NAND4_in[2] ,
         \SB1_2_30/Component_Function_1/NAND4_in[1] ,
         \SB1_2_30/Component_Function_1/NAND4_in[0] ,
         \SB1_2_30/Component_Function_5/NAND4_in[2] ,
         \SB1_2_30/Component_Function_5/NAND4_in[0] ,
         \SB1_2_31/Component_Function_0/NAND4_in[2] ,
         \SB1_2_31/Component_Function_0/NAND4_in[1] ,
         \SB1_2_31/Component_Function_0/NAND4_in[0] ,
         \SB1_2_31/Component_Function_1/NAND4_in[3] ,
         \SB1_2_31/Component_Function_1/NAND4_in[2] ,
         \SB1_2_31/Component_Function_1/NAND4_in[1] ,
         \SB1_2_31/Component_Function_1/NAND4_in[0] ,
         \SB1_2_31/Component_Function_5/NAND4_in[2] ,
         \SB1_2_31/Component_Function_5/NAND4_in[1] ,
         \SB2_2_0/Component_Function_0/NAND4_in[1] ,
         \SB2_2_0/Component_Function_0/NAND4_in[0] ,
         \SB2_2_0/Component_Function_1/NAND4_in[3] ,
         \SB2_2_0/Component_Function_1/NAND4_in[2] ,
         \SB2_2_0/Component_Function_1/NAND4_in[1] ,
         \SB2_2_0/Component_Function_1/NAND4_in[0] ,
         \SB2_2_0/Component_Function_5/NAND4_in[2] ,
         \SB2_2_1/Component_Function_0/NAND4_in[1] ,
         \SB2_2_1/Component_Function_0/NAND4_in[0] ,
         \SB2_2_1/Component_Function_1/NAND4_in[3] ,
         \SB2_2_1/Component_Function_1/NAND4_in[1] ,
         \SB2_2_1/Component_Function_1/NAND4_in[0] ,
         \SB2_2_1/Component_Function_5/NAND4_in[2] ,
         \SB2_2_1/Component_Function_5/NAND4_in[0] ,
         \SB2_2_2/Component_Function_0/NAND4_in[3] ,
         \SB2_2_2/Component_Function_0/NAND4_in[2] ,
         \SB2_2_2/Component_Function_0/NAND4_in[1] ,
         \SB2_2_2/Component_Function_0/NAND4_in[0] ,
         \SB2_2_2/Component_Function_1/NAND4_in[3] ,
         \SB2_2_2/Component_Function_1/NAND4_in[2] ,
         \SB2_2_2/Component_Function_1/NAND4_in[1] ,
         \SB2_2_2/Component_Function_1/NAND4_in[0] ,
         \SB2_2_2/Component_Function_5/NAND4_in[2] ,
         \SB2_2_2/Component_Function_5/NAND4_in[1] ,
         \SB2_2_3/Component_Function_0/NAND4_in[2] ,
         \SB2_2_3/Component_Function_0/NAND4_in[1] ,
         \SB2_2_3/Component_Function_0/NAND4_in[0] ,
         \SB2_2_3/Component_Function_1/NAND4_in[3] ,
         \SB2_2_3/Component_Function_1/NAND4_in[0] ,
         \SB2_2_3/Component_Function_5/NAND4_in[2] ,
         \SB2_2_3/Component_Function_5/NAND4_in[1] ,
         \SB2_2_3/Component_Function_5/NAND4_in[0] ,
         \SB2_2_4/Component_Function_0/NAND4_in[2] ,
         \SB2_2_4/Component_Function_0/NAND4_in[1] ,
         \SB2_2_4/Component_Function_0/NAND4_in[0] ,
         \SB2_2_4/Component_Function_1/NAND4_in[3] ,
         \SB2_2_4/Component_Function_1/NAND4_in[1] ,
         \SB2_2_4/Component_Function_1/NAND4_in[0] ,
         \SB2_2_4/Component_Function_5/NAND4_in[3] ,
         \SB2_2_4/Component_Function_5/NAND4_in[2] ,
         \SB2_2_4/Component_Function_5/NAND4_in[1] ,
         \SB2_2_4/Component_Function_5/NAND4_in[0] ,
         \SB2_2_5/Component_Function_0/NAND4_in[3] ,
         \SB2_2_5/Component_Function_0/NAND4_in[2] ,
         \SB2_2_5/Component_Function_0/NAND4_in[0] ,
         \SB2_2_5/Component_Function_1/NAND4_in[2] ,
         \SB2_2_5/Component_Function_1/NAND4_in[1] ,
         \SB2_2_5/Component_Function_1/NAND4_in[0] ,
         \SB2_2_5/Component_Function_5/NAND4_in[3] ,
         \SB2_2_5/Component_Function_5/NAND4_in[0] ,
         \SB2_2_6/Component_Function_0/NAND4_in[3] ,
         \SB2_2_6/Component_Function_0/NAND4_in[1] ,
         \SB2_2_6/Component_Function_0/NAND4_in[0] ,
         \SB2_2_6/Component_Function_1/NAND4_in[3] ,
         \SB2_2_6/Component_Function_1/NAND4_in[2] ,
         \SB2_2_6/Component_Function_1/NAND4_in[1] ,
         \SB2_2_6/Component_Function_1/NAND4_in[0] ,
         \SB2_2_6/Component_Function_5/NAND4_in[3] ,
         \SB2_2_6/Component_Function_5/NAND4_in[0] ,
         \SB2_2_7/Component_Function_0/NAND4_in[2] ,
         \SB2_2_7/Component_Function_0/NAND4_in[1] ,
         \SB2_2_7/Component_Function_0/NAND4_in[0] ,
         \SB2_2_7/Component_Function_1/NAND4_in[3] ,
         \SB2_2_7/Component_Function_1/NAND4_in[2] ,
         \SB2_2_7/Component_Function_1/NAND4_in[1] ,
         \SB2_2_7/Component_Function_1/NAND4_in[0] ,
         \SB2_2_7/Component_Function_5/NAND4_in[3] ,
         \SB2_2_7/Component_Function_5/NAND4_in[2] ,
         \SB2_2_7/Component_Function_5/NAND4_in[1] ,
         \SB2_2_7/Component_Function_5/NAND4_in[0] ,
         \SB2_2_8/Component_Function_0/NAND4_in[1] ,
         \SB2_2_8/Component_Function_1/NAND4_in[3] ,
         \SB2_2_8/Component_Function_1/NAND4_in[2] ,
         \SB2_2_8/Component_Function_1/NAND4_in[1] ,
         \SB2_2_8/Component_Function_1/NAND4_in[0] ,
         \SB2_2_8/Component_Function_5/NAND4_in[3] ,
         \SB2_2_8/Component_Function_5/NAND4_in[2] ,
         \SB2_2_8/Component_Function_5/NAND4_in[1] ,
         \SB2_2_8/Component_Function_5/NAND4_in[0] ,
         \SB2_2_9/Component_Function_0/NAND4_in[3] ,
         \SB2_2_9/Component_Function_0/NAND4_in[2] ,
         \SB2_2_9/Component_Function_0/NAND4_in[0] ,
         \SB2_2_9/Component_Function_1/NAND4_in[3] ,
         \SB2_2_9/Component_Function_1/NAND4_in[2] ,
         \SB2_2_9/Component_Function_1/NAND4_in[1] ,
         \SB2_2_9/Component_Function_1/NAND4_in[0] ,
         \SB2_2_9/Component_Function_5/NAND4_in[2] ,
         \SB2_2_9/Component_Function_5/NAND4_in[0] ,
         \SB2_2_10/Component_Function_0/NAND4_in[2] ,
         \SB2_2_10/Component_Function_0/NAND4_in[1] ,
         \SB2_2_10/Component_Function_0/NAND4_in[0] ,
         \SB2_2_10/Component_Function_1/NAND4_in[2] ,
         \SB2_2_10/Component_Function_1/NAND4_in[1] ,
         \SB2_2_10/Component_Function_1/NAND4_in[0] ,
         \SB2_2_10/Component_Function_5/NAND4_in[2] ,
         \SB2_2_10/Component_Function_5/NAND4_in[1] ,
         \SB2_2_10/Component_Function_5/NAND4_in[0] ,
         \SB2_2_11/Component_Function_0/NAND4_in[3] ,
         \SB2_2_11/Component_Function_0/NAND4_in[1] ,
         \SB2_2_11/Component_Function_0/NAND4_in[0] ,
         \SB2_2_11/Component_Function_1/NAND4_in[2] ,
         \SB2_2_11/Component_Function_1/NAND4_in[1] ,
         \SB2_2_11/Component_Function_1/NAND4_in[0] ,
         \SB2_2_11/Component_Function_5/NAND4_in[2] ,
         \SB2_2_12/Component_Function_0/NAND4_in[3] ,
         \SB2_2_12/Component_Function_0/NAND4_in[2] ,
         \SB2_2_12/Component_Function_0/NAND4_in[1] ,
         \SB2_2_12/Component_Function_0/NAND4_in[0] ,
         \SB2_2_12/Component_Function_1/NAND4_in[2] ,
         \SB2_2_12/Component_Function_1/NAND4_in[0] ,
         \SB2_2_12/Component_Function_5/NAND4_in[1] ,
         \SB2_2_12/Component_Function_5/NAND4_in[0] ,
         \SB2_2_13/Component_Function_0/NAND4_in[3] ,
         \SB2_2_13/Component_Function_0/NAND4_in[2] ,
         \SB2_2_13/Component_Function_0/NAND4_in[1] ,
         \SB2_2_13/Component_Function_0/NAND4_in[0] ,
         \SB2_2_13/Component_Function_1/NAND4_in[2] ,
         \SB2_2_13/Component_Function_1/NAND4_in[1] ,
         \SB2_2_13/Component_Function_1/NAND4_in[0] ,
         \SB2_2_13/Component_Function_5/NAND4_in[3] ,
         \SB2_2_13/Component_Function_5/NAND4_in[2] ,
         \SB2_2_13/Component_Function_5/NAND4_in[1] ,
         \SB2_2_13/Component_Function_5/NAND4_in[0] ,
         \SB2_2_14/Component_Function_0/NAND4_in[3] ,
         \SB2_2_14/Component_Function_0/NAND4_in[2] ,
         \SB2_2_14/Component_Function_0/NAND4_in[0] ,
         \SB2_2_14/Component_Function_1/NAND4_in[3] ,
         \SB2_2_14/Component_Function_1/NAND4_in[1] ,
         \SB2_2_14/Component_Function_1/NAND4_in[0] ,
         \SB2_2_14/Component_Function_5/NAND4_in[3] ,
         \SB2_2_14/Component_Function_5/NAND4_in[2] ,
         \SB2_2_14/Component_Function_5/NAND4_in[1] ,
         \SB2_2_14/Component_Function_5/NAND4_in[0] ,
         \SB2_2_15/Component_Function_0/NAND4_in[2] ,
         \SB2_2_15/Component_Function_0/NAND4_in[1] ,
         \SB2_2_15/Component_Function_0/NAND4_in[0] ,
         \SB2_2_15/Component_Function_1/NAND4_in[3] ,
         \SB2_2_15/Component_Function_1/NAND4_in[2] ,
         \SB2_2_15/Component_Function_1/NAND4_in[1] ,
         \SB2_2_15/Component_Function_1/NAND4_in[0] ,
         \SB2_2_15/Component_Function_5/NAND4_in[3] ,
         \SB2_2_15/Component_Function_5/NAND4_in[0] ,
         \SB2_2_16/Component_Function_0/NAND4_in[1] ,
         \SB2_2_16/Component_Function_0/NAND4_in[0] ,
         \SB2_2_16/Component_Function_1/NAND4_in[2] ,
         \SB2_2_16/Component_Function_1/NAND4_in[1] ,
         \SB2_2_16/Component_Function_1/NAND4_in[0] ,
         \SB2_2_16/Component_Function_5/NAND4_in[2] ,
         \SB2_2_17/Component_Function_0/NAND4_in[3] ,
         \SB2_2_17/Component_Function_0/NAND4_in[1] ,
         \SB2_2_17/Component_Function_0/NAND4_in[0] ,
         \SB2_2_17/Component_Function_1/NAND4_in[3] ,
         \SB2_2_17/Component_Function_1/NAND4_in[2] ,
         \SB2_2_17/Component_Function_1/NAND4_in[1] ,
         \SB2_2_17/Component_Function_1/NAND4_in[0] ,
         \SB2_2_17/Component_Function_5/NAND4_in[2] ,
         \SB2_2_17/Component_Function_5/NAND4_in[0] ,
         \SB2_2_18/Component_Function_0/NAND4_in[3] ,
         \SB2_2_18/Component_Function_0/NAND4_in[2] ,
         \SB2_2_18/Component_Function_0/NAND4_in[1] ,
         \SB2_2_18/Component_Function_0/NAND4_in[0] ,
         \SB2_2_18/Component_Function_1/NAND4_in[2] ,
         \SB2_2_18/Component_Function_1/NAND4_in[1] ,
         \SB2_2_18/Component_Function_1/NAND4_in[0] ,
         \SB2_2_18/Component_Function_5/NAND4_in[2] ,
         \SB2_2_18/Component_Function_5/NAND4_in[0] ,
         \SB2_2_19/Component_Function_0/NAND4_in[3] ,
         \SB2_2_19/Component_Function_0/NAND4_in[2] ,
         \SB2_2_19/Component_Function_0/NAND4_in[1] ,
         \SB2_2_19/Component_Function_0/NAND4_in[0] ,
         \SB2_2_19/Component_Function_1/NAND4_in[3] ,
         \SB2_2_19/Component_Function_1/NAND4_in[1] ,
         \SB2_2_19/Component_Function_1/NAND4_in[0] ,
         \SB2_2_19/Component_Function_5/NAND4_in[3] ,
         \SB2_2_20/Component_Function_0/NAND4_in[3] ,
         \SB2_2_20/Component_Function_0/NAND4_in[2] ,
         \SB2_2_20/Component_Function_0/NAND4_in[1] ,
         \SB2_2_20/Component_Function_0/NAND4_in[0] ,
         \SB2_2_20/Component_Function_1/NAND4_in[3] ,
         \SB2_2_20/Component_Function_1/NAND4_in[2] ,
         \SB2_2_20/Component_Function_1/NAND4_in[1] ,
         \SB2_2_20/Component_Function_1/NAND4_in[0] ,
         \SB2_2_20/Component_Function_5/NAND4_in[1] ,
         \SB2_2_20/Component_Function_5/NAND4_in[0] ,
         \SB2_2_21/Component_Function_0/NAND4_in[2] ,
         \SB2_2_21/Component_Function_0/NAND4_in[1] ,
         \SB2_2_21/Component_Function_1/NAND4_in[2] ,
         \SB2_2_21/Component_Function_1/NAND4_in[1] ,
         \SB2_2_21/Component_Function_1/NAND4_in[0] ,
         \SB2_2_21/Component_Function_5/NAND4_in[2] ,
         \SB2_2_21/Component_Function_5/NAND4_in[0] ,
         \SB2_2_22/Component_Function_0/NAND4_in[3] ,
         \SB2_2_22/Component_Function_0/NAND4_in[1] ,
         \SB2_2_22/Component_Function_0/NAND4_in[0] ,
         \SB2_2_22/Component_Function_1/NAND4_in[3] ,
         \SB2_2_22/Component_Function_1/NAND4_in[0] ,
         \SB2_2_22/Component_Function_5/NAND4_in[3] ,
         \SB2_2_23/Component_Function_0/NAND4_in[1] ,
         \SB2_2_23/Component_Function_0/NAND4_in[0] ,
         \SB2_2_23/Component_Function_1/NAND4_in[2] ,
         \SB2_2_23/Component_Function_1/NAND4_in[1] ,
         \SB2_2_23/Component_Function_1/NAND4_in[0] ,
         \SB2_2_23/Component_Function_5/NAND4_in[2] ,
         \SB2_2_23/Component_Function_5/NAND4_in[1] ,
         \SB2_2_23/Component_Function_5/NAND4_in[0] ,
         \SB2_2_24/Component_Function_0/NAND4_in[3] ,
         \SB2_2_24/Component_Function_0/NAND4_in[2] ,
         \SB2_2_24/Component_Function_0/NAND4_in[1] ,
         \SB2_2_24/Component_Function_0/NAND4_in[0] ,
         \SB2_2_24/Component_Function_1/NAND4_in[3] ,
         \SB2_2_24/Component_Function_1/NAND4_in[1] ,
         \SB2_2_24/Component_Function_1/NAND4_in[0] ,
         \SB2_2_24/Component_Function_5/NAND4_in[3] ,
         \SB2_2_24/Component_Function_5/NAND4_in[1] ,
         \SB2_2_25/Component_Function_0/NAND4_in[3] ,
         \SB2_2_25/Component_Function_0/NAND4_in[2] ,
         \SB2_2_25/Component_Function_0/NAND4_in[1] ,
         \SB2_2_25/Component_Function_0/NAND4_in[0] ,
         \SB2_2_25/Component_Function_1/NAND4_in[3] ,
         \SB2_2_25/Component_Function_1/NAND4_in[1] ,
         \SB2_2_25/Component_Function_1/NAND4_in[0] ,
         \SB2_2_25/Component_Function_5/NAND4_in[2] ,
         \SB2_2_25/Component_Function_5/NAND4_in[0] ,
         \SB2_2_26/Component_Function_0/NAND4_in[3] ,
         \SB2_2_26/Component_Function_0/NAND4_in[2] ,
         \SB2_2_26/Component_Function_0/NAND4_in[1] ,
         \SB2_2_26/Component_Function_0/NAND4_in[0] ,
         \SB2_2_26/Component_Function_1/NAND4_in[3] ,
         \SB2_2_26/Component_Function_1/NAND4_in[2] ,
         \SB2_2_26/Component_Function_1/NAND4_in[1] ,
         \SB2_2_26/Component_Function_1/NAND4_in[0] ,
         \SB2_2_26/Component_Function_5/NAND4_in[2] ,
         \SB2_2_26/Component_Function_5/NAND4_in[1] ,
         \SB2_2_26/Component_Function_5/NAND4_in[0] ,
         \SB2_2_27/Component_Function_0/NAND4_in[3] ,
         \SB2_2_27/Component_Function_0/NAND4_in[2] ,
         \SB2_2_27/Component_Function_0/NAND4_in[0] ,
         \SB2_2_27/Component_Function_1/NAND4_in[2] ,
         \SB2_2_27/Component_Function_1/NAND4_in[1] ,
         \SB2_2_27/Component_Function_1/NAND4_in[0] ,
         \SB2_2_27/Component_Function_5/NAND4_in[3] ,
         \SB2_2_27/Component_Function_5/NAND4_in[1] ,
         \SB2_2_28/Component_Function_0/NAND4_in[3] ,
         \SB2_2_28/Component_Function_0/NAND4_in[2] ,
         \SB2_2_28/Component_Function_0/NAND4_in[1] ,
         \SB2_2_28/Component_Function_0/NAND4_in[0] ,
         \SB2_2_28/Component_Function_1/NAND4_in[3] ,
         \SB2_2_28/Component_Function_1/NAND4_in[1] ,
         \SB2_2_28/Component_Function_1/NAND4_in[0] ,
         \SB2_2_28/Component_Function_5/NAND4_in[3] ,
         \SB2_2_28/Component_Function_5/NAND4_in[1] ,
         \SB2_2_28/Component_Function_5/NAND4_in[0] ,
         \SB2_2_29/Component_Function_0/NAND4_in[2] ,
         \SB2_2_29/Component_Function_0/NAND4_in[1] ,
         \SB2_2_29/Component_Function_0/NAND4_in[0] ,
         \SB2_2_29/Component_Function_1/NAND4_in[3] ,
         \SB2_2_29/Component_Function_1/NAND4_in[2] ,
         \SB2_2_29/Component_Function_1/NAND4_in[1] ,
         \SB2_2_29/Component_Function_1/NAND4_in[0] ,
         \SB2_2_29/Component_Function_5/NAND4_in[2] ,
         \SB2_2_29/Component_Function_5/NAND4_in[1] ,
         \SB2_2_29/Component_Function_5/NAND4_in[0] ,
         \SB2_2_30/Component_Function_0/NAND4_in[3] ,
         \SB2_2_30/Component_Function_0/NAND4_in[1] ,
         \SB2_2_30/Component_Function_0/NAND4_in[0] ,
         \SB2_2_30/Component_Function_1/NAND4_in[2] ,
         \SB2_2_30/Component_Function_1/NAND4_in[1] ,
         \SB2_2_30/Component_Function_1/NAND4_in[0] ,
         \SB2_2_30/Component_Function_5/NAND4_in[3] ,
         \SB2_2_30/Component_Function_5/NAND4_in[1] ,
         \SB2_2_30/Component_Function_5/NAND4_in[0] ,
         \SB2_2_31/Component_Function_0/NAND4_in[3] ,
         \SB2_2_31/Component_Function_0/NAND4_in[2] ,
         \SB2_2_31/Component_Function_0/NAND4_in[0] ,
         \SB2_2_31/Component_Function_1/NAND4_in[3] ,
         \SB2_2_31/Component_Function_1/NAND4_in[2] ,
         \SB2_2_31/Component_Function_1/NAND4_in[1] ,
         \SB2_2_31/Component_Function_1/NAND4_in[0] ,
         \SB2_2_31/Component_Function_5/NAND4_in[3] ,
         \SB2_2_31/Component_Function_5/NAND4_in[1] ,
         \SB2_2_31/Component_Function_5/NAND4_in[0] ,
         \SB1_3_0/Component_Function_0/NAND4_in[2] ,
         \SB1_3_0/Component_Function_0/NAND4_in[1] ,
         \SB1_3_0/Component_Function_0/NAND4_in[0] ,
         \SB1_3_0/Component_Function_1/NAND4_in[3] ,
         \SB1_3_0/Component_Function_1/NAND4_in[2] ,
         \SB1_3_0/Component_Function_1/NAND4_in[1] ,
         \SB1_3_0/Component_Function_1/NAND4_in[0] ,
         \SB1_3_0/Component_Function_5/NAND4_in[3] ,
         \SB1_3_0/Component_Function_5/NAND4_in[0] ,
         \SB1_3_1/Component_Function_0/NAND4_in[2] ,
         \SB1_3_1/Component_Function_0/NAND4_in[1] ,
         \SB1_3_1/Component_Function_0/NAND4_in[0] ,
         \SB1_3_1/Component_Function_1/NAND4_in[3] ,
         \SB1_3_1/Component_Function_1/NAND4_in[2] ,
         \SB1_3_1/Component_Function_1/NAND4_in[1] ,
         \SB1_3_1/Component_Function_1/NAND4_in[0] ,
         \SB1_3_1/Component_Function_5/NAND4_in[1] ,
         \SB1_3_1/Component_Function_5/NAND4_in[0] ,
         \SB1_3_2/Component_Function_0/NAND4_in[2] ,
         \SB1_3_2/Component_Function_0/NAND4_in[1] ,
         \SB1_3_2/Component_Function_0/NAND4_in[0] ,
         \SB1_3_2/Component_Function_1/NAND4_in[3] ,
         \SB1_3_2/Component_Function_1/NAND4_in[2] ,
         \SB1_3_2/Component_Function_1/NAND4_in[1] ,
         \SB1_3_2/Component_Function_1/NAND4_in[0] ,
         \SB1_3_2/Component_Function_5/NAND4_in[2] ,
         \SB1_3_2/Component_Function_5/NAND4_in[0] ,
         \SB1_3_3/Component_Function_0/NAND4_in[3] ,
         \SB1_3_3/Component_Function_0/NAND4_in[2] ,
         \SB1_3_3/Component_Function_0/NAND4_in[1] ,
         \SB1_3_3/Component_Function_0/NAND4_in[0] ,
         \SB1_3_3/Component_Function_1/NAND4_in[2] ,
         \SB1_3_3/Component_Function_1/NAND4_in[1] ,
         \SB1_3_3/Component_Function_5/NAND4_in[2] ,
         \SB1_3_3/Component_Function_5/NAND4_in[1] ,
         \SB1_3_3/Component_Function_5/NAND4_in[0] ,
         \SB1_3_4/Component_Function_0/NAND4_in[3] ,
         \SB1_3_4/Component_Function_0/NAND4_in[2] ,
         \SB1_3_4/Component_Function_0/NAND4_in[1] ,
         \SB1_3_4/Component_Function_0/NAND4_in[0] ,
         \SB1_3_4/Component_Function_1/NAND4_in[3] ,
         \SB1_3_4/Component_Function_1/NAND4_in[2] ,
         \SB1_3_4/Component_Function_1/NAND4_in[1] ,
         \SB1_3_4/Component_Function_5/NAND4_in[3] ,
         \SB1_3_4/Component_Function_5/NAND4_in[2] ,
         \SB1_3_5/Component_Function_0/NAND4_in[3] ,
         \SB1_3_5/Component_Function_0/NAND4_in[2] ,
         \SB1_3_5/Component_Function_0/NAND4_in[1] ,
         \SB1_3_5/Component_Function_0/NAND4_in[0] ,
         \SB1_3_5/Component_Function_1/NAND4_in[3] ,
         \SB1_3_5/Component_Function_1/NAND4_in[1] ,
         \SB1_3_5/Component_Function_1/NAND4_in[0] ,
         \SB1_3_5/Component_Function_5/NAND4_in[2] ,
         \SB1_3_5/Component_Function_5/NAND4_in[0] ,
         \SB1_3_6/Component_Function_0/NAND4_in[3] ,
         \SB1_3_6/Component_Function_0/NAND4_in[2] ,
         \SB1_3_6/Component_Function_0/NAND4_in[1] ,
         \SB1_3_6/Component_Function_0/NAND4_in[0] ,
         \SB1_3_6/Component_Function_1/NAND4_in[3] ,
         \SB1_3_6/Component_Function_1/NAND4_in[1] ,
         \SB1_3_6/Component_Function_5/NAND4_in[3] ,
         \SB1_3_6/Component_Function_5/NAND4_in[1] ,
         \SB1_3_6/Component_Function_5/NAND4_in[0] ,
         \SB1_3_7/Component_Function_0/NAND4_in[2] ,
         \SB1_3_7/Component_Function_0/NAND4_in[1] ,
         \SB1_3_7/Component_Function_0/NAND4_in[0] ,
         \SB1_3_7/Component_Function_1/NAND4_in[3] ,
         \SB1_3_7/Component_Function_1/NAND4_in[2] ,
         \SB1_3_7/Component_Function_1/NAND4_in[0] ,
         \SB1_3_7/Component_Function_5/NAND4_in[1] ,
         \SB1_3_7/Component_Function_5/NAND4_in[0] ,
         \SB1_3_8/Component_Function_0/NAND4_in[3] ,
         \SB1_3_8/Component_Function_0/NAND4_in[2] ,
         \SB1_3_8/Component_Function_0/NAND4_in[1] ,
         \SB1_3_8/Component_Function_0/NAND4_in[0] ,
         \SB1_3_8/Component_Function_1/NAND4_in[2] ,
         \SB1_3_8/Component_Function_1/NAND4_in[1] ,
         \SB1_3_8/Component_Function_1/NAND4_in[0] ,
         \SB1_3_8/Component_Function_5/NAND4_in[2] ,
         \SB1_3_8/Component_Function_5/NAND4_in[1] ,
         \SB1_3_8/Component_Function_5/NAND4_in[0] ,
         \SB1_3_9/Component_Function_0/NAND4_in[3] ,
         \SB1_3_9/Component_Function_0/NAND4_in[2] ,
         \SB1_3_9/Component_Function_0/NAND4_in[1] ,
         \SB1_3_9/Component_Function_0/NAND4_in[0] ,
         \SB1_3_9/Component_Function_1/NAND4_in[3] ,
         \SB1_3_9/Component_Function_1/NAND4_in[2] ,
         \SB1_3_9/Component_Function_1/NAND4_in[1] ,
         \SB1_3_9/Component_Function_1/NAND4_in[0] ,
         \SB1_3_9/Component_Function_5/NAND4_in[3] ,
         \SB1_3_9/Component_Function_5/NAND4_in[2] ,
         \SB1_3_9/Component_Function_5/NAND4_in[1] ,
         \SB1_3_9/Component_Function_5/NAND4_in[0] ,
         \SB1_3_10/Component_Function_0/NAND4_in[3] ,
         \SB1_3_10/Component_Function_0/NAND4_in[2] ,
         \SB1_3_10/Component_Function_0/NAND4_in[1] ,
         \SB1_3_10/Component_Function_0/NAND4_in[0] ,
         \SB1_3_10/Component_Function_1/NAND4_in[2] ,
         \SB1_3_10/Component_Function_1/NAND4_in[1] ,
         \SB1_3_10/Component_Function_1/NAND4_in[0] ,
         \SB1_3_10/Component_Function_5/NAND4_in[2] ,
         \SB1_3_11/Component_Function_0/NAND4_in[3] ,
         \SB1_3_11/Component_Function_0/NAND4_in[2] ,
         \SB1_3_11/Component_Function_0/NAND4_in[1] ,
         \SB1_3_11/Component_Function_1/NAND4_in[2] ,
         \SB1_3_11/Component_Function_1/NAND4_in[1] ,
         \SB1_3_11/Component_Function_5/NAND4_in[3] ,
         \SB1_3_11/Component_Function_5/NAND4_in[0] ,
         \SB1_3_12/Component_Function_0/NAND4_in[3] ,
         \SB1_3_12/Component_Function_0/NAND4_in[2] ,
         \SB1_3_12/Component_Function_0/NAND4_in[1] ,
         \SB1_3_12/Component_Function_0/NAND4_in[0] ,
         \SB1_3_12/Component_Function_1/NAND4_in[3] ,
         \SB1_3_12/Component_Function_1/NAND4_in[2] ,
         \SB1_3_12/Component_Function_1/NAND4_in[1] ,
         \SB1_3_12/Component_Function_5/NAND4_in[2] ,
         \SB1_3_12/Component_Function_5/NAND4_in[1] ,
         \SB1_3_12/Component_Function_5/NAND4_in[0] ,
         \SB1_3_13/Component_Function_0/NAND4_in[2] ,
         \SB1_3_13/Component_Function_0/NAND4_in[1] ,
         \SB1_3_13/Component_Function_0/NAND4_in[0] ,
         \SB1_3_13/Component_Function_1/NAND4_in[3] ,
         \SB1_3_13/Component_Function_1/NAND4_in[2] ,
         \SB1_3_13/Component_Function_1/NAND4_in[1] ,
         \SB1_3_13/Component_Function_1/NAND4_in[0] ,
         \SB1_3_13/Component_Function_5/NAND4_in[2] ,
         \SB1_3_13/Component_Function_5/NAND4_in[0] ,
         \SB1_3_14/Component_Function_0/NAND4_in[2] ,
         \SB1_3_14/Component_Function_0/NAND4_in[1] ,
         \SB1_3_14/Component_Function_0/NAND4_in[0] ,
         \SB1_3_14/Component_Function_1/NAND4_in[3] ,
         \SB1_3_14/Component_Function_1/NAND4_in[2] ,
         \SB1_3_14/Component_Function_1/NAND4_in[1] ,
         \SB1_3_14/Component_Function_1/NAND4_in[0] ,
         \SB1_3_14/Component_Function_5/NAND4_in[0] ,
         \SB1_3_15/Component_Function_0/NAND4_in[3] ,
         \SB1_3_15/Component_Function_0/NAND4_in[2] ,
         \SB1_3_15/Component_Function_0/NAND4_in[1] ,
         \SB1_3_15/Component_Function_0/NAND4_in[0] ,
         \SB1_3_15/Component_Function_1/NAND4_in[2] ,
         \SB1_3_15/Component_Function_1/NAND4_in[1] ,
         \SB1_3_15/Component_Function_1/NAND4_in[0] ,
         \SB1_3_15/Component_Function_5/NAND4_in[3] ,
         \SB1_3_15/Component_Function_5/NAND4_in[2] ,
         \SB1_3_15/Component_Function_5/NAND4_in[1] ,
         \SB1_3_16/Component_Function_0/NAND4_in[3] ,
         \SB1_3_16/Component_Function_0/NAND4_in[2] ,
         \SB1_3_16/Component_Function_0/NAND4_in[1] ,
         \SB1_3_16/Component_Function_0/NAND4_in[0] ,
         \SB1_3_16/Component_Function_1/NAND4_in[3] ,
         \SB1_3_16/Component_Function_1/NAND4_in[1] ,
         \SB1_3_16/Component_Function_1/NAND4_in[0] ,
         \SB1_3_16/Component_Function_5/NAND4_in[0] ,
         \SB1_3_17/Component_Function_0/NAND4_in[0] ,
         \SB1_3_17/Component_Function_1/NAND4_in[2] ,
         \SB1_3_17/Component_Function_1/NAND4_in[1] ,
         \SB1_3_17/Component_Function_5/NAND4_in[3] ,
         \SB1_3_17/Component_Function_5/NAND4_in[1] ,
         \SB1_3_17/Component_Function_5/NAND4_in[0] ,
         \SB1_3_18/Component_Function_0/NAND4_in[2] ,
         \SB1_3_18/Component_Function_0/NAND4_in[1] ,
         \SB1_3_18/Component_Function_0/NAND4_in[0] ,
         \SB1_3_18/Component_Function_1/NAND4_in[3] ,
         \SB1_3_18/Component_Function_1/NAND4_in[2] ,
         \SB1_3_18/Component_Function_1/NAND4_in[1] ,
         \SB1_3_18/Component_Function_5/NAND4_in[3] ,
         \SB1_3_18/Component_Function_5/NAND4_in[1] ,
         \SB1_3_18/Component_Function_5/NAND4_in[0] ,
         \SB1_3_19/Component_Function_0/NAND4_in[3] ,
         \SB1_3_19/Component_Function_0/NAND4_in[2] ,
         \SB1_3_19/Component_Function_0/NAND4_in[1] ,
         \SB1_3_19/Component_Function_0/NAND4_in[0] ,
         \SB1_3_19/Component_Function_1/NAND4_in[3] ,
         \SB1_3_19/Component_Function_1/NAND4_in[2] ,
         \SB1_3_19/Component_Function_1/NAND4_in[1] ,
         \SB1_3_19/Component_Function_1/NAND4_in[0] ,
         \SB1_3_19/Component_Function_5/NAND4_in[2] ,
         \SB1_3_19/Component_Function_5/NAND4_in[1] ,
         \SB1_3_19/Component_Function_5/NAND4_in[0] ,
         \SB1_3_20/Component_Function_0/NAND4_in[3] ,
         \SB1_3_20/Component_Function_0/NAND4_in[2] ,
         \SB1_3_20/Component_Function_0/NAND4_in[1] ,
         \SB1_3_20/Component_Function_0/NAND4_in[0] ,
         \SB1_3_20/Component_Function_1/NAND4_in[1] ,
         \SB1_3_20/Component_Function_1/NAND4_in[0] ,
         \SB1_3_20/Component_Function_5/NAND4_in[1] ,
         \SB1_3_20/Component_Function_5/NAND4_in[0] ,
         \SB1_3_21/Component_Function_0/NAND4_in[3] ,
         \SB1_3_21/Component_Function_0/NAND4_in[2] ,
         \SB1_3_21/Component_Function_0/NAND4_in[1] ,
         \SB1_3_21/Component_Function_0/NAND4_in[0] ,
         \SB1_3_21/Component_Function_1/NAND4_in[2] ,
         \SB1_3_21/Component_Function_1/NAND4_in[1] ,
         \SB1_3_21/Component_Function_1/NAND4_in[0] ,
         \SB1_3_21/Component_Function_5/NAND4_in[1] ,
         \SB1_3_21/Component_Function_5/NAND4_in[0] ,
         \SB1_3_22/Component_Function_0/NAND4_in[3] ,
         \SB1_3_22/Component_Function_0/NAND4_in[2] ,
         \SB1_3_22/Component_Function_0/NAND4_in[1] ,
         \SB1_3_22/Component_Function_0/NAND4_in[0] ,
         \SB1_3_22/Component_Function_1/NAND4_in[3] ,
         \SB1_3_22/Component_Function_1/NAND4_in[2] ,
         \SB1_3_22/Component_Function_1/NAND4_in[1] ,
         \SB1_3_22/Component_Function_1/NAND4_in[0] ,
         \SB1_3_22/Component_Function_5/NAND4_in[3] ,
         \SB1_3_22/Component_Function_5/NAND4_in[1] ,
         \SB1_3_22/Component_Function_5/NAND4_in[0] ,
         \SB1_3_23/Component_Function_0/NAND4_in[3] ,
         \SB1_3_23/Component_Function_0/NAND4_in[2] ,
         \SB1_3_23/Component_Function_0/NAND4_in[1] ,
         \SB1_3_23/Component_Function_1/NAND4_in[2] ,
         \SB1_3_23/Component_Function_1/NAND4_in[1] ,
         \SB1_3_23/Component_Function_1/NAND4_in[0] ,
         \SB1_3_23/Component_Function_5/NAND4_in[3] ,
         \SB1_3_23/Component_Function_5/NAND4_in[1] ,
         \SB1_3_23/Component_Function_5/NAND4_in[0] ,
         \SB1_3_24/Component_Function_0/NAND4_in[2] ,
         \SB1_3_24/Component_Function_0/NAND4_in[1] ,
         \SB1_3_24/Component_Function_0/NAND4_in[0] ,
         \SB1_3_24/Component_Function_1/NAND4_in[2] ,
         \SB1_3_24/Component_Function_1/NAND4_in[1] ,
         \SB1_3_24/Component_Function_5/NAND4_in[2] ,
         \SB1_3_24/Component_Function_5/NAND4_in[0] ,
         \SB1_3_25/Component_Function_0/NAND4_in[3] ,
         \SB1_3_25/Component_Function_0/NAND4_in[2] ,
         \SB1_3_25/Component_Function_0/NAND4_in[1] ,
         \SB1_3_25/Component_Function_0/NAND4_in[0] ,
         \SB1_3_25/Component_Function_1/NAND4_in[3] ,
         \SB1_3_25/Component_Function_1/NAND4_in[1] ,
         \SB1_3_25/Component_Function_1/NAND4_in[0] ,
         \SB1_3_25/Component_Function_5/NAND4_in[1] ,
         \SB1_3_26/Component_Function_0/NAND4_in[1] ,
         \SB1_3_26/Component_Function_0/NAND4_in[0] ,
         \SB1_3_26/Component_Function_1/NAND4_in[1] ,
         \SB1_3_26/Component_Function_1/NAND4_in[0] ,
         \SB1_3_26/Component_Function_5/NAND4_in[2] ,
         \SB1_3_26/Component_Function_5/NAND4_in[1] ,
         \SB1_3_26/Component_Function_5/NAND4_in[0] ,
         \SB1_3_27/Component_Function_0/NAND4_in[2] ,
         \SB1_3_27/Component_Function_0/NAND4_in[1] ,
         \SB1_3_27/Component_Function_0/NAND4_in[0] ,
         \SB1_3_27/Component_Function_1/NAND4_in[2] ,
         \SB1_3_27/Component_Function_1/NAND4_in[1] ,
         \SB1_3_27/Component_Function_1/NAND4_in[0] ,
         \SB1_3_27/Component_Function_5/NAND4_in[2] ,
         \SB1_3_27/Component_Function_5/NAND4_in[1] ,
         \SB1_3_28/Component_Function_0/NAND4_in[2] ,
         \SB1_3_28/Component_Function_0/NAND4_in[1] ,
         \SB1_3_28/Component_Function_0/NAND4_in[0] ,
         \SB1_3_28/Component_Function_1/NAND4_in[2] ,
         \SB1_3_28/Component_Function_1/NAND4_in[1] ,
         \SB1_3_28/Component_Function_1/NAND4_in[0] ,
         \SB1_3_28/Component_Function_5/NAND4_in[1] ,
         \SB1_3_28/Component_Function_5/NAND4_in[0] ,
         \SB1_3_29/Component_Function_0/NAND4_in[3] ,
         \SB1_3_29/Component_Function_0/NAND4_in[2] ,
         \SB1_3_29/Component_Function_0/NAND4_in[1] ,
         \SB1_3_29/Component_Function_0/NAND4_in[0] ,
         \SB1_3_29/Component_Function_1/NAND4_in[3] ,
         \SB1_3_29/Component_Function_1/NAND4_in[1] ,
         \SB1_3_29/Component_Function_1/NAND4_in[0] ,
         \SB1_3_29/Component_Function_5/NAND4_in[1] ,
         \SB1_3_29/Component_Function_5/NAND4_in[0] ,
         \SB1_3_30/Component_Function_0/NAND4_in[3] ,
         \SB1_3_30/Component_Function_0/NAND4_in[2] ,
         \SB1_3_30/Component_Function_0/NAND4_in[1] ,
         \SB1_3_30/Component_Function_0/NAND4_in[0] ,
         \SB1_3_30/Component_Function_1/NAND4_in[3] ,
         \SB1_3_30/Component_Function_1/NAND4_in[1] ,
         \SB1_3_30/Component_Function_1/NAND4_in[0] ,
         \SB1_3_30/Component_Function_5/NAND4_in[2] ,
         \SB1_3_30/Component_Function_5/NAND4_in[1] ,
         \SB1_3_30/Component_Function_5/NAND4_in[0] ,
         \SB1_3_31/Component_Function_0/NAND4_in[2] ,
         \SB1_3_31/Component_Function_0/NAND4_in[1] ,
         \SB1_3_31/Component_Function_1/NAND4_in[3] ,
         \SB1_3_31/Component_Function_1/NAND4_in[1] ,
         \SB1_3_31/Component_Function_1/NAND4_in[0] ,
         \SB1_3_31/Component_Function_5/NAND4_in[2] ,
         \SB1_3_31/Component_Function_5/NAND4_in[1] ,
         \SB1_3_31/Component_Function_5/NAND4_in[0] ,
         \SB2_3_0/Component_Function_0/NAND4_in[3] ,
         \SB2_3_0/Component_Function_0/NAND4_in[2] ,
         \SB2_3_0/Component_Function_0/NAND4_in[0] ,
         \SB2_3_0/Component_Function_1/NAND4_in[3] ,
         \SB2_3_0/Component_Function_1/NAND4_in[1] ,
         \SB2_3_0/Component_Function_1/NAND4_in[0] ,
         \SB2_3_0/Component_Function_5/NAND4_in[1] ,
         \SB2_3_0/Component_Function_5/NAND4_in[0] ,
         \SB2_3_1/Component_Function_0/NAND4_in[2] ,
         \SB2_3_1/Component_Function_0/NAND4_in[1] ,
         \SB2_3_1/Component_Function_0/NAND4_in[0] ,
         \SB2_3_1/Component_Function_1/NAND4_in[2] ,
         \SB2_3_1/Component_Function_1/NAND4_in[1] ,
         \SB2_3_1/Component_Function_1/NAND4_in[0] ,
         \SB2_3_1/Component_Function_5/NAND4_in[2] ,
         \SB2_3_1/Component_Function_5/NAND4_in[1] ,
         \SB2_3_1/Component_Function_5/NAND4_in[0] ,
         \SB2_3_2/Component_Function_0/NAND4_in[3] ,
         \SB2_3_2/Component_Function_0/NAND4_in[1] ,
         \SB2_3_2/Component_Function_0/NAND4_in[0] ,
         \SB2_3_2/Component_Function_1/NAND4_in[3] ,
         \SB2_3_2/Component_Function_1/NAND4_in[2] ,
         \SB2_3_2/Component_Function_1/NAND4_in[1] ,
         \SB2_3_2/Component_Function_1/NAND4_in[0] ,
         \SB2_3_2/Component_Function_5/NAND4_in[2] ,
         \SB2_3_2/Component_Function_5/NAND4_in[0] ,
         \SB2_3_3/Component_Function_0/NAND4_in[3] ,
         \SB2_3_3/Component_Function_0/NAND4_in[2] ,
         \SB2_3_3/Component_Function_0/NAND4_in[1] ,
         \SB2_3_3/Component_Function_0/NAND4_in[0] ,
         \SB2_3_3/Component_Function_5/NAND4_in[2] ,
         \SB2_3_4/Component_Function_0/NAND4_in[2] ,
         \SB2_3_4/Component_Function_0/NAND4_in[1] ,
         \SB2_3_4/Component_Function_0/NAND4_in[0] ,
         \SB2_3_4/Component_Function_1/NAND4_in[1] ,
         \SB2_3_4/Component_Function_1/NAND4_in[0] ,
         \SB2_3_4/Component_Function_5/NAND4_in[2] ,
         \SB2_3_4/Component_Function_5/NAND4_in[1] ,
         \SB2_3_4/Component_Function_5/NAND4_in[0] ,
         \SB2_3_5/Component_Function_0/NAND4_in[2] ,
         \SB2_3_5/Component_Function_0/NAND4_in[1] ,
         \SB2_3_5/Component_Function_0/NAND4_in[0] ,
         \SB2_3_5/Component_Function_1/NAND4_in[3] ,
         \SB2_3_5/Component_Function_1/NAND4_in[2] ,
         \SB2_3_5/Component_Function_1/NAND4_in[1] ,
         \SB2_3_5/Component_Function_1/NAND4_in[0] ,
         \SB2_3_5/Component_Function_5/NAND4_in[1] ,
         \SB2_3_5/Component_Function_5/NAND4_in[0] ,
         \SB2_3_6/Component_Function_0/NAND4_in[2] ,
         \SB2_3_6/Component_Function_0/NAND4_in[1] ,
         \SB2_3_6/Component_Function_0/NAND4_in[0] ,
         \SB2_3_6/Component_Function_1/NAND4_in[2] ,
         \SB2_3_6/Component_Function_1/NAND4_in[1] ,
         \SB2_3_6/Component_Function_1/NAND4_in[0] ,
         \SB2_3_6/Component_Function_5/NAND4_in[2] ,
         \SB2_3_6/Component_Function_5/NAND4_in[0] ,
         \SB2_3_7/Component_Function_0/NAND4_in[3] ,
         \SB2_3_7/Component_Function_0/NAND4_in[1] ,
         \SB2_3_7/Component_Function_0/NAND4_in[0] ,
         \SB2_3_7/Component_Function_1/NAND4_in[3] ,
         \SB2_3_7/Component_Function_1/NAND4_in[2] ,
         \SB2_3_7/Component_Function_1/NAND4_in[0] ,
         \SB2_3_7/Component_Function_5/NAND4_in[3] ,
         \SB2_3_7/Component_Function_5/NAND4_in[2] ,
         \SB2_3_7/Component_Function_5/NAND4_in[0] ,
         \SB2_3_8/Component_Function_0/NAND4_in[3] ,
         \SB2_3_8/Component_Function_0/NAND4_in[2] ,
         \SB2_3_8/Component_Function_0/NAND4_in[0] ,
         \SB2_3_8/Component_Function_1/NAND4_in[3] ,
         \SB2_3_8/Component_Function_1/NAND4_in[1] ,
         \SB2_3_8/Component_Function_1/NAND4_in[0] ,
         \SB2_3_8/Component_Function_5/NAND4_in[3] ,
         \SB2_3_8/Component_Function_5/NAND4_in[2] ,
         \SB2_3_8/Component_Function_5/NAND4_in[0] ,
         \SB2_3_9/Component_Function_0/NAND4_in[1] ,
         \SB2_3_9/Component_Function_0/NAND4_in[0] ,
         \SB2_3_9/Component_Function_1/NAND4_in[3] ,
         \SB2_3_9/Component_Function_1/NAND4_in[2] ,
         \SB2_3_9/Component_Function_1/NAND4_in[1] ,
         \SB2_3_9/Component_Function_1/NAND4_in[0] ,
         \SB2_3_9/Component_Function_5/NAND4_in[1] ,
         \SB2_3_9/Component_Function_5/NAND4_in[0] ,
         \SB2_3_10/Component_Function_0/NAND4_in[3] ,
         \SB2_3_10/Component_Function_0/NAND4_in[2] ,
         \SB2_3_10/Component_Function_0/NAND4_in[1] ,
         \SB2_3_10/Component_Function_0/NAND4_in[0] ,
         \SB2_3_10/Component_Function_1/NAND4_in[3] ,
         \SB2_3_10/Component_Function_1/NAND4_in[2] ,
         \SB2_3_10/Component_Function_1/NAND4_in[1] ,
         \SB2_3_10/Component_Function_1/NAND4_in[0] ,
         \SB2_3_10/Component_Function_5/NAND4_in[2] ,
         \SB2_3_10/Component_Function_5/NAND4_in[1] ,
         \SB2_3_10/Component_Function_5/NAND4_in[0] ,
         \SB2_3_11/Component_Function_0/NAND4_in[3] ,
         \SB2_3_11/Component_Function_0/NAND4_in[1] ,
         \SB2_3_11/Component_Function_1/NAND4_in[3] ,
         \SB2_3_11/Component_Function_1/NAND4_in[2] ,
         \SB2_3_11/Component_Function_1/NAND4_in[1] ,
         \SB2_3_11/Component_Function_1/NAND4_in[0] ,
         \SB2_3_11/Component_Function_5/NAND4_in[2] ,
         \SB2_3_11/Component_Function_5/NAND4_in[1] ,
         \SB2_3_11/Component_Function_5/NAND4_in[0] ,
         \SB2_3_12/Component_Function_0/NAND4_in[3] ,
         \SB2_3_12/Component_Function_0/NAND4_in[2] ,
         \SB2_3_12/Component_Function_0/NAND4_in[1] ,
         \SB2_3_12/Component_Function_0/NAND4_in[0] ,
         \SB2_3_12/Component_Function_1/NAND4_in[2] ,
         \SB2_3_12/Component_Function_1/NAND4_in[1] ,
         \SB2_3_12/Component_Function_1/NAND4_in[0] ,
         \SB2_3_12/Component_Function_5/NAND4_in[2] ,
         \SB2_3_13/Component_Function_0/NAND4_in[3] ,
         \SB2_3_13/Component_Function_0/NAND4_in[1] ,
         \SB2_3_13/Component_Function_0/NAND4_in[0] ,
         \SB2_3_13/Component_Function_1/NAND4_in[3] ,
         \SB2_3_13/Component_Function_1/NAND4_in[2] ,
         \SB2_3_13/Component_Function_1/NAND4_in[1] ,
         \SB2_3_13/Component_Function_1/NAND4_in[0] ,
         \SB2_3_13/Component_Function_5/NAND4_in[3] ,
         \SB2_3_14/Component_Function_0/NAND4_in[3] ,
         \SB2_3_14/Component_Function_0/NAND4_in[1] ,
         \SB2_3_14/Component_Function_0/NAND4_in[0] ,
         \SB2_3_14/Component_Function_1/NAND4_in[3] ,
         \SB2_3_14/Component_Function_1/NAND4_in[2] ,
         \SB2_3_14/Component_Function_1/NAND4_in[1] ,
         \SB2_3_14/Component_Function_1/NAND4_in[0] ,
         \SB2_3_14/Component_Function_5/NAND4_in[3] ,
         \SB2_3_14/Component_Function_5/NAND4_in[0] ,
         \SB2_3_15/Component_Function_0/NAND4_in[3] ,
         \SB2_3_15/Component_Function_0/NAND4_in[1] ,
         \SB2_3_15/Component_Function_0/NAND4_in[0] ,
         \SB2_3_15/Component_Function_1/NAND4_in[3] ,
         \SB2_3_15/Component_Function_1/NAND4_in[2] ,
         \SB2_3_15/Component_Function_1/NAND4_in[0] ,
         \SB2_3_15/Component_Function_5/NAND4_in[2] ,
         \SB2_3_15/Component_Function_5/NAND4_in[1] ,
         \SB2_3_15/Component_Function_5/NAND4_in[0] ,
         \SB2_3_16/Component_Function_0/NAND4_in[3] ,
         \SB2_3_16/Component_Function_0/NAND4_in[2] ,
         \SB2_3_16/Component_Function_0/NAND4_in[1] ,
         \SB2_3_16/Component_Function_1/NAND4_in[2] ,
         \SB2_3_16/Component_Function_1/NAND4_in[1] ,
         \SB2_3_16/Component_Function_1/NAND4_in[0] ,
         \SB2_3_16/Component_Function_5/NAND4_in[2] ,
         \SB2_3_16/Component_Function_5/NAND4_in[0] ,
         \SB2_3_17/Component_Function_0/NAND4_in[3] ,
         \SB2_3_17/Component_Function_0/NAND4_in[1] ,
         \SB2_3_17/Component_Function_0/NAND4_in[0] ,
         \SB2_3_17/Component_Function_1/NAND4_in[3] ,
         \SB2_3_17/Component_Function_1/NAND4_in[2] ,
         \SB2_3_17/Component_Function_1/NAND4_in[1] ,
         \SB2_3_17/Component_Function_1/NAND4_in[0] ,
         \SB2_3_17/Component_Function_5/NAND4_in[3] ,
         \SB2_3_17/Component_Function_5/NAND4_in[2] ,
         \SB2_3_17/Component_Function_5/NAND4_in[0] ,
         \SB2_3_18/Component_Function_0/NAND4_in[1] ,
         \SB2_3_18/Component_Function_0/NAND4_in[0] ,
         \SB2_3_18/Component_Function_1/NAND4_in[3] ,
         \SB2_3_18/Component_Function_1/NAND4_in[2] ,
         \SB2_3_18/Component_Function_1/NAND4_in[1] ,
         \SB2_3_18/Component_Function_1/NAND4_in[0] ,
         \SB2_3_19/Component_Function_0/NAND4_in[1] ,
         \SB2_3_19/Component_Function_0/NAND4_in[0] ,
         \SB2_3_19/Component_Function_1/NAND4_in[3] ,
         \SB2_3_19/Component_Function_1/NAND4_in[2] ,
         \SB2_3_19/Component_Function_1/NAND4_in[1] ,
         \SB2_3_19/Component_Function_1/NAND4_in[0] ,
         \SB2_3_19/Component_Function_5/NAND4_in[1] ,
         \SB2_3_19/Component_Function_5/NAND4_in[0] ,
         \SB2_3_20/Component_Function_0/NAND4_in[3] ,
         \SB2_3_20/Component_Function_0/NAND4_in[2] ,
         \SB2_3_20/Component_Function_0/NAND4_in[1] ,
         \SB2_3_20/Component_Function_0/NAND4_in[0] ,
         \SB2_3_20/Component_Function_1/NAND4_in[2] ,
         \SB2_3_20/Component_Function_1/NAND4_in[1] ,
         \SB2_3_20/Component_Function_1/NAND4_in[0] ,
         \SB2_3_20/Component_Function_5/NAND4_in[2] ,
         \SB2_3_20/Component_Function_5/NAND4_in[1] ,
         \SB2_3_20/Component_Function_5/NAND4_in[0] ,
         \SB2_3_21/Component_Function_0/NAND4_in[2] ,
         \SB2_3_21/Component_Function_0/NAND4_in[0] ,
         \SB2_3_21/Component_Function_1/NAND4_in[2] ,
         \SB2_3_21/Component_Function_1/NAND4_in[1] ,
         \SB2_3_21/Component_Function_1/NAND4_in[0] ,
         \SB2_3_21/Component_Function_5/NAND4_in[3] ,
         \SB2_3_21/Component_Function_5/NAND4_in[2] ,
         \SB2_3_21/Component_Function_5/NAND4_in[0] ,
         \SB2_3_22/Component_Function_0/NAND4_in[3] ,
         \SB2_3_22/Component_Function_0/NAND4_in[2] ,
         \SB2_3_22/Component_Function_0/NAND4_in[1] ,
         \SB2_3_22/Component_Function_0/NAND4_in[0] ,
         \SB2_3_22/Component_Function_1/NAND4_in[3] ,
         \SB2_3_22/Component_Function_1/NAND4_in[2] ,
         \SB2_3_22/Component_Function_1/NAND4_in[1] ,
         \SB2_3_22/Component_Function_1/NAND4_in[0] ,
         \SB2_3_23/Component_Function_0/NAND4_in[2] ,
         \SB2_3_23/Component_Function_0/NAND4_in[1] ,
         \SB2_3_23/Component_Function_0/NAND4_in[0] ,
         \SB2_3_23/Component_Function_1/NAND4_in[3] ,
         \SB2_3_23/Component_Function_1/NAND4_in[1] ,
         \SB2_3_23/Component_Function_1/NAND4_in[0] ,
         \SB2_3_24/Component_Function_0/NAND4_in[3] ,
         \SB2_3_24/Component_Function_0/NAND4_in[0] ,
         \SB2_3_24/Component_Function_1/NAND4_in[1] ,
         \SB2_3_24/Component_Function_1/NAND4_in[0] ,
         \SB2_3_24/Component_Function_5/NAND4_in[3] ,
         \SB2_3_24/Component_Function_5/NAND4_in[2] ,
         \SB2_3_24/Component_Function_5/NAND4_in[0] ,
         \SB2_3_25/Component_Function_0/NAND4_in[2] ,
         \SB2_3_25/Component_Function_0/NAND4_in[0] ,
         \SB2_3_25/Component_Function_1/NAND4_in[3] ,
         \SB2_3_25/Component_Function_1/NAND4_in[2] ,
         \SB2_3_25/Component_Function_1/NAND4_in[1] ,
         \SB2_3_25/Component_Function_1/NAND4_in[0] ,
         \SB2_3_25/Component_Function_5/NAND4_in[3] ,
         \SB2_3_25/Component_Function_5/NAND4_in[0] ,
         \SB2_3_26/Component_Function_0/NAND4_in[3] ,
         \SB2_3_26/Component_Function_0/NAND4_in[1] ,
         \SB2_3_26/Component_Function_0/NAND4_in[0] ,
         \SB2_3_26/Component_Function_1/NAND4_in[3] ,
         \SB2_3_26/Component_Function_1/NAND4_in[2] ,
         \SB2_3_26/Component_Function_1/NAND4_in[1] ,
         \SB2_3_26/Component_Function_1/NAND4_in[0] ,
         \SB2_3_26/Component_Function_5/NAND4_in[3] ,
         \SB2_3_26/Component_Function_5/NAND4_in[0] ,
         \SB2_3_27/Component_Function_0/NAND4_in[3] ,
         \SB2_3_27/Component_Function_0/NAND4_in[2] ,
         \SB2_3_27/Component_Function_0/NAND4_in[1] ,
         \SB2_3_27/Component_Function_0/NAND4_in[0] ,
         \SB2_3_27/Component_Function_1/NAND4_in[2] ,
         \SB2_3_27/Component_Function_1/NAND4_in[1] ,
         \SB2_3_27/Component_Function_1/NAND4_in[0] ,
         \SB2_3_27/Component_Function_5/NAND4_in[1] ,
         \SB2_3_27/Component_Function_5/NAND4_in[0] ,
         \SB2_3_28/Component_Function_0/NAND4_in[3] ,
         \SB2_3_28/Component_Function_0/NAND4_in[2] ,
         \SB2_3_28/Component_Function_0/NAND4_in[1] ,
         \SB2_3_28/Component_Function_0/NAND4_in[0] ,
         \SB2_3_28/Component_Function_1/NAND4_in[3] ,
         \SB2_3_28/Component_Function_1/NAND4_in[2] ,
         \SB2_3_28/Component_Function_1/NAND4_in[1] ,
         \SB2_3_28/Component_Function_1/NAND4_in[0] ,
         \SB2_3_28/Component_Function_5/NAND4_in[2] ,
         \SB2_3_28/Component_Function_5/NAND4_in[1] ,
         \SB2_3_28/Component_Function_5/NAND4_in[0] ,
         \SB2_3_29/Component_Function_0/NAND4_in[1] ,
         \SB2_3_29/Component_Function_0/NAND4_in[0] ,
         \SB2_3_29/Component_Function_1/NAND4_in[3] ,
         \SB2_3_29/Component_Function_1/NAND4_in[0] ,
         \SB2_3_29/Component_Function_5/NAND4_in[2] ,
         \SB2_3_29/Component_Function_5/NAND4_in[1] ,
         \SB2_3_29/Component_Function_5/NAND4_in[0] ,
         \SB2_3_30/Component_Function_0/NAND4_in[3] ,
         \SB2_3_30/Component_Function_0/NAND4_in[1] ,
         \SB2_3_30/Component_Function_0/NAND4_in[0] ,
         \SB2_3_30/Component_Function_1/NAND4_in[3] ,
         \SB2_3_30/Component_Function_1/NAND4_in[2] ,
         \SB2_3_30/Component_Function_1/NAND4_in[1] ,
         \SB2_3_30/Component_Function_1/NAND4_in[0] ,
         \SB2_3_30/Component_Function_5/NAND4_in[1] ,
         \SB2_3_31/Component_Function_0/NAND4_in[2] ,
         \SB2_3_31/Component_Function_0/NAND4_in[1] ,
         \SB2_3_31/Component_Function_0/NAND4_in[0] ,
         \SB2_3_31/Component_Function_1/NAND4_in[3] ,
         \SB2_3_31/Component_Function_1/NAND4_in[1] ,
         \SB2_3_31/Component_Function_1/NAND4_in[0] ,
         \SB2_3_31/Component_Function_5/NAND4_in[0] ,
         \SB3_0/Component_Function_0/NAND4_in[3] ,
         \SB3_0/Component_Function_0/NAND4_in[2] ,
         \SB3_0/Component_Function_0/NAND4_in[1] ,
         \SB3_0/Component_Function_0/NAND4_in[0] ,
         \SB3_0/Component_Function_1/NAND4_in[2] ,
         \SB3_0/Component_Function_1/NAND4_in[1] ,
         \SB3_0/Component_Function_5/NAND4_in[3] ,
         \SB3_0/Component_Function_5/NAND4_in[1] ,
         \SB3_1/Component_Function_0/NAND4_in[2] ,
         \SB3_1/Component_Function_0/NAND4_in[1] ,
         \SB3_1/Component_Function_0/NAND4_in[0] ,
         \SB3_1/Component_Function_1/NAND4_in[3] ,
         \SB3_1/Component_Function_1/NAND4_in[2] ,
         \SB3_1/Component_Function_1/NAND4_in[0] ,
         \SB3_1/Component_Function_5/NAND4_in[1] ,
         \SB3_1/Component_Function_5/NAND4_in[0] ,
         \SB3_2/Component_Function_0/NAND4_in[2] ,
         \SB3_2/Component_Function_0/NAND4_in[1] ,
         \SB3_2/Component_Function_0/NAND4_in[0] ,
         \SB3_2/Component_Function_1/NAND4_in[1] ,
         \SB3_2/Component_Function_1/NAND4_in[0] ,
         \SB3_2/Component_Function_5/NAND4_in[1] ,
         \SB3_2/Component_Function_5/NAND4_in[0] ,
         \SB3_3/Component_Function_0/NAND4_in[3] ,
         \SB3_3/Component_Function_0/NAND4_in[2] ,
         \SB3_3/Component_Function_0/NAND4_in[1] ,
         \SB3_3/Component_Function_0/NAND4_in[0] ,
         \SB3_3/Component_Function_1/NAND4_in[3] ,
         \SB3_3/Component_Function_1/NAND4_in[1] ,
         \SB3_3/Component_Function_1/NAND4_in[0] ,
         \SB3_3/Component_Function_5/NAND4_in[2] ,
         \SB3_3/Component_Function_5/NAND4_in[1] ,
         \SB3_3/Component_Function_5/NAND4_in[0] ,
         \SB3_4/Component_Function_0/NAND4_in[2] ,
         \SB3_4/Component_Function_0/NAND4_in[1] ,
         \SB3_4/Component_Function_0/NAND4_in[0] ,
         \SB3_4/Component_Function_1/NAND4_in[3] ,
         \SB3_4/Component_Function_1/NAND4_in[1] ,
         \SB3_4/Component_Function_1/NAND4_in[0] ,
         \SB3_4/Component_Function_5/NAND4_in[2] ,
         \SB3_4/Component_Function_5/NAND4_in[1] ,
         \SB3_5/Component_Function_0/NAND4_in[2] ,
         \SB3_5/Component_Function_0/NAND4_in[1] ,
         \SB3_5/Component_Function_0/NAND4_in[0] ,
         \SB3_5/Component_Function_1/NAND4_in[3] ,
         \SB3_5/Component_Function_1/NAND4_in[2] ,
         \SB3_5/Component_Function_1/NAND4_in[1] ,
         \SB3_5/Component_Function_5/NAND4_in[3] ,
         \SB3_6/Component_Function_0/NAND4_in[1] ,
         \SB3_6/Component_Function_0/NAND4_in[0] ,
         \SB3_6/Component_Function_1/NAND4_in[3] ,
         \SB3_6/Component_Function_1/NAND4_in[2] ,
         \SB3_6/Component_Function_1/NAND4_in[1] ,
         \SB3_6/Component_Function_5/NAND4_in[3] ,
         \SB3_6/Component_Function_5/NAND4_in[2] ,
         \SB3_6/Component_Function_5/NAND4_in[1] ,
         \SB3_6/Component_Function_5/NAND4_in[0] ,
         \SB3_7/Component_Function_0/NAND4_in[3] ,
         \SB3_7/Component_Function_0/NAND4_in[1] ,
         \SB3_7/Component_Function_0/NAND4_in[0] ,
         \SB3_7/Component_Function_1/NAND4_in[3] ,
         \SB3_7/Component_Function_1/NAND4_in[2] ,
         \SB3_7/Component_Function_1/NAND4_in[1] ,
         \SB3_7/Component_Function_1/NAND4_in[0] ,
         \SB3_7/Component_Function_5/NAND4_in[2] ,
         \SB3_8/Component_Function_0/NAND4_in[2] ,
         \SB3_8/Component_Function_0/NAND4_in[1] ,
         \SB3_8/Component_Function_0/NAND4_in[0] ,
         \SB3_8/Component_Function_1/NAND4_in[3] ,
         \SB3_8/Component_Function_1/NAND4_in[2] ,
         \SB3_8/Component_Function_1/NAND4_in[1] ,
         \SB3_8/Component_Function_5/NAND4_in[3] ,
         \SB3_8/Component_Function_5/NAND4_in[1] ,
         \SB3_8/Component_Function_5/NAND4_in[0] ,
         \SB3_9/Component_Function_0/NAND4_in[3] ,
         \SB3_9/Component_Function_0/NAND4_in[2] ,
         \SB3_9/Component_Function_0/NAND4_in[1] ,
         \SB3_9/Component_Function_0/NAND4_in[0] ,
         \SB3_9/Component_Function_1/NAND4_in[3] ,
         \SB3_9/Component_Function_1/NAND4_in[1] ,
         \SB3_9/Component_Function_1/NAND4_in[0] ,
         \SB3_9/Component_Function_5/NAND4_in[2] ,
         \SB3_9/Component_Function_5/NAND4_in[0] ,
         \SB3_10/Component_Function_0/NAND4_in[3] ,
         \SB3_10/Component_Function_0/NAND4_in[2] ,
         \SB3_10/Component_Function_0/NAND4_in[1] ,
         \SB3_10/Component_Function_0/NAND4_in[0] ,
         \SB3_10/Component_Function_1/NAND4_in[3] ,
         \SB3_10/Component_Function_1/NAND4_in[0] ,
         \SB3_11/Component_Function_0/NAND4_in[3] ,
         \SB3_11/Component_Function_0/NAND4_in[2] ,
         \SB3_11/Component_Function_0/NAND4_in[1] ,
         \SB3_11/Component_Function_0/NAND4_in[0] ,
         \SB3_11/Component_Function_1/NAND4_in[3] ,
         \SB3_11/Component_Function_1/NAND4_in[2] ,
         \SB3_11/Component_Function_1/NAND4_in[1] ,
         \SB3_11/Component_Function_1/NAND4_in[0] ,
         \SB3_11/Component_Function_5/NAND4_in[2] ,
         \SB3_11/Component_Function_5/NAND4_in[0] ,
         \SB3_12/Component_Function_0/NAND4_in[2] ,
         \SB3_12/Component_Function_0/NAND4_in[1] ,
         \SB3_12/Component_Function_0/NAND4_in[0] ,
         \SB3_12/Component_Function_1/NAND4_in[3] ,
         \SB3_12/Component_Function_1/NAND4_in[1] ,
         \SB3_12/Component_Function_1/NAND4_in[0] ,
         \SB3_12/Component_Function_5/NAND4_in[2] ,
         \SB3_12/Component_Function_5/NAND4_in[1] ,
         \SB3_13/Component_Function_0/NAND4_in[3] ,
         \SB3_13/Component_Function_0/NAND4_in[2] ,
         \SB3_13/Component_Function_0/NAND4_in[1] ,
         \SB3_13/Component_Function_0/NAND4_in[0] ,
         \SB3_13/Component_Function_1/NAND4_in[3] ,
         \SB3_13/Component_Function_1/NAND4_in[2] ,
         \SB3_13/Component_Function_1/NAND4_in[1] ,
         \SB3_13/Component_Function_1/NAND4_in[0] ,
         \SB3_13/Component_Function_5/NAND4_in[2] ,
         \SB3_13/Component_Function_5/NAND4_in[1] ,
         \SB3_14/Component_Function_0/NAND4_in[2] ,
         \SB3_14/Component_Function_0/NAND4_in[1] ,
         \SB3_14/Component_Function_0/NAND4_in[0] ,
         \SB3_14/Component_Function_1/NAND4_in[2] ,
         \SB3_14/Component_Function_1/NAND4_in[1] ,
         \SB3_14/Component_Function_1/NAND4_in[0] ,
         \SB3_14/Component_Function_5/NAND4_in[1] ,
         \SB3_14/Component_Function_5/NAND4_in[0] ,
         \SB3_15/Component_Function_0/NAND4_in[1] ,
         \SB3_15/Component_Function_1/NAND4_in[3] ,
         \SB3_15/Component_Function_1/NAND4_in[2] ,
         \SB3_15/Component_Function_1/NAND4_in[1] ,
         \SB3_15/Component_Function_1/NAND4_in[0] ,
         \SB3_15/Component_Function_5/NAND4_in[3] ,
         \SB3_15/Component_Function_5/NAND4_in[2] ,
         \SB3_15/Component_Function_5/NAND4_in[1] ,
         \SB3_15/Component_Function_5/NAND4_in[0] ,
         \SB3_16/Component_Function_0/NAND4_in[3] ,
         \SB3_16/Component_Function_0/NAND4_in[1] ,
         \SB3_16/Component_Function_0/NAND4_in[0] ,
         \SB3_16/Component_Function_1/NAND4_in[0] ,
         \SB3_16/Component_Function_5/NAND4_in[2] ,
         \SB3_16/Component_Function_5/NAND4_in[1] ,
         \SB3_16/Component_Function_5/NAND4_in[0] ,
         \SB3_17/Component_Function_0/NAND4_in[3] ,
         \SB3_17/Component_Function_0/NAND4_in[2] ,
         \SB3_17/Component_Function_0/NAND4_in[1] ,
         \SB3_17/Component_Function_0/NAND4_in[0] ,
         \SB3_17/Component_Function_1/NAND4_in[3] ,
         \SB3_17/Component_Function_1/NAND4_in[2] ,
         \SB3_17/Component_Function_1/NAND4_in[1] ,
         \SB3_17/Component_Function_1/NAND4_in[0] ,
         \SB3_17/Component_Function_5/NAND4_in[2] ,
         \SB3_17/Component_Function_5/NAND4_in[1] ,
         \SB3_17/Component_Function_5/NAND4_in[0] ,
         \SB3_18/Component_Function_0/NAND4_in[3] ,
         \SB3_18/Component_Function_0/NAND4_in[2] ,
         \SB3_18/Component_Function_0/NAND4_in[1] ,
         \SB3_18/Component_Function_0/NAND4_in[0] ,
         \SB3_18/Component_Function_1/NAND4_in[3] ,
         \SB3_18/Component_Function_1/NAND4_in[1] ,
         \SB3_18/Component_Function_1/NAND4_in[0] ,
         \SB3_18/Component_Function_5/NAND4_in[2] ,
         \SB3_18/Component_Function_5/NAND4_in[0] ,
         \SB3_19/Component_Function_0/NAND4_in[3] ,
         \SB3_19/Component_Function_0/NAND4_in[2] ,
         \SB3_19/Component_Function_0/NAND4_in[1] ,
         \SB3_19/Component_Function_0/NAND4_in[0] ,
         \SB3_19/Component_Function_1/NAND4_in[3] ,
         \SB3_19/Component_Function_1/NAND4_in[2] ,
         \SB3_19/Component_Function_1/NAND4_in[1] ,
         \SB3_19/Component_Function_1/NAND4_in[0] ,
         \SB3_19/Component_Function_5/NAND4_in[3] ,
         \SB3_19/Component_Function_5/NAND4_in[2] ,
         \SB3_19/Component_Function_5/NAND4_in[1] ,
         \SB3_19/Component_Function_5/NAND4_in[0] ,
         \SB3_20/Component_Function_0/NAND4_in[3] ,
         \SB3_20/Component_Function_0/NAND4_in[2] ,
         \SB3_20/Component_Function_0/NAND4_in[1] ,
         \SB3_20/Component_Function_0/NAND4_in[0] ,
         \SB3_20/Component_Function_1/NAND4_in[3] ,
         \SB3_20/Component_Function_1/NAND4_in[2] ,
         \SB3_20/Component_Function_1/NAND4_in[1] ,
         \SB3_20/Component_Function_1/NAND4_in[0] ,
         \SB3_20/Component_Function_5/NAND4_in[1] ,
         \SB3_21/Component_Function_0/NAND4_in[2] ,
         \SB3_21/Component_Function_0/NAND4_in[1] ,
         \SB3_21/Component_Function_0/NAND4_in[0] ,
         \SB3_21/Component_Function_1/NAND4_in[3] ,
         \SB3_21/Component_Function_1/NAND4_in[2] ,
         \SB3_21/Component_Function_1/NAND4_in[1] ,
         \SB3_21/Component_Function_1/NAND4_in[0] ,
         \SB3_21/Component_Function_5/NAND4_in[3] ,
         \SB3_21/Component_Function_5/NAND4_in[1] ,
         \SB3_21/Component_Function_5/NAND4_in[0] ,
         \SB3_22/Component_Function_0/NAND4_in[3] ,
         \SB3_22/Component_Function_0/NAND4_in[2] ,
         \SB3_22/Component_Function_0/NAND4_in[1] ,
         \SB3_22/Component_Function_0/NAND4_in[0] ,
         \SB3_22/Component_Function_1/NAND4_in[2] ,
         \SB3_22/Component_Function_1/NAND4_in[0] ,
         \SB3_22/Component_Function_5/NAND4_in[2] ,
         \SB3_22/Component_Function_5/NAND4_in[1] ,
         \SB3_22/Component_Function_5/NAND4_in[0] ,
         \SB3_23/Component_Function_0/NAND4_in[3] ,
         \SB3_23/Component_Function_0/NAND4_in[2] ,
         \SB3_23/Component_Function_1/NAND4_in[1] ,
         \SB3_23/Component_Function_5/NAND4_in[2] ,
         \SB3_23/Component_Function_5/NAND4_in[1] ,
         \SB3_24/Component_Function_0/NAND4_in[3] ,
         \SB3_24/Component_Function_0/NAND4_in[1] ,
         \SB3_24/Component_Function_0/NAND4_in[0] ,
         \SB3_24/Component_Function_1/NAND4_in[2] ,
         \SB3_24/Component_Function_1/NAND4_in[1] ,
         \SB3_24/Component_Function_1/NAND4_in[0] ,
         \SB3_24/Component_Function_5/NAND4_in[3] ,
         \SB3_25/Component_Function_0/NAND4_in[3] ,
         \SB3_25/Component_Function_0/NAND4_in[2] ,
         \SB3_25/Component_Function_0/NAND4_in[1] ,
         \SB3_25/Component_Function_0/NAND4_in[0] ,
         \SB3_25/Component_Function_1/NAND4_in[2] ,
         \SB3_25/Component_Function_1/NAND4_in[1] ,
         \SB3_25/Component_Function_1/NAND4_in[0] ,
         \SB3_25/Component_Function_5/NAND4_in[3] ,
         \SB3_25/Component_Function_5/NAND4_in[1] ,
         \SB3_25/Component_Function_5/NAND4_in[0] ,
         \SB3_26/Component_Function_0/NAND4_in[3] ,
         \SB3_26/Component_Function_0/NAND4_in[2] ,
         \SB3_26/Component_Function_0/NAND4_in[1] ,
         \SB3_26/Component_Function_0/NAND4_in[0] ,
         \SB3_26/Component_Function_1/NAND4_in[3] ,
         \SB3_26/Component_Function_1/NAND4_in[2] ,
         \SB3_26/Component_Function_1/NAND4_in[1] ,
         \SB3_26/Component_Function_1/NAND4_in[0] ,
         \SB3_26/Component_Function_5/NAND4_in[3] ,
         \SB3_26/Component_Function_5/NAND4_in[1] ,
         \SB3_26/Component_Function_5/NAND4_in[0] ,
         \SB3_27/Component_Function_0/NAND4_in[2] ,
         \SB3_27/Component_Function_0/NAND4_in[1] ,
         \SB3_27/Component_Function_0/NAND4_in[0] ,
         \SB3_27/Component_Function_1/NAND4_in[3] ,
         \SB3_27/Component_Function_1/NAND4_in[2] ,
         \SB3_27/Component_Function_1/NAND4_in[1] ,
         \SB3_27/Component_Function_1/NAND4_in[0] ,
         \SB3_27/Component_Function_5/NAND4_in[3] ,
         \SB3_27/Component_Function_5/NAND4_in[0] ,
         \SB3_28/Component_Function_0/NAND4_in[2] ,
         \SB3_28/Component_Function_0/NAND4_in[1] ,
         \SB3_28/Component_Function_0/NAND4_in[0] ,
         \SB3_28/Component_Function_1/NAND4_in[2] ,
         \SB3_28/Component_Function_1/NAND4_in[1] ,
         \SB3_28/Component_Function_1/NAND4_in[0] ,
         \SB3_28/Component_Function_5/NAND4_in[2] ,
         \SB3_28/Component_Function_5/NAND4_in[1] ,
         \SB3_28/Component_Function_5/NAND4_in[0] ,
         \SB3_29/Component_Function_0/NAND4_in[3] ,
         \SB3_29/Component_Function_0/NAND4_in[2] ,
         \SB3_29/Component_Function_0/NAND4_in[1] ,
         \SB3_29/Component_Function_0/NAND4_in[0] ,
         \SB3_29/Component_Function_1/NAND4_in[2] ,
         \SB3_29/Component_Function_1/NAND4_in[1] ,
         \SB3_29/Component_Function_1/NAND4_in[0] ,
         \SB3_29/Component_Function_5/NAND4_in[0] ,
         \SB3_30/Component_Function_0/NAND4_in[3] ,
         \SB3_30/Component_Function_0/NAND4_in[1] ,
         \SB3_30/Component_Function_0/NAND4_in[0] ,
         \SB3_30/Component_Function_1/NAND4_in[2] ,
         \SB3_30/Component_Function_1/NAND4_in[1] ,
         \SB3_30/Component_Function_1/NAND4_in[0] ,
         \SB3_30/Component_Function_5/NAND4_in[1] ,
         \SB3_30/Component_Function_5/NAND4_in[0] ,
         \SB3_31/Component_Function_0/NAND4_in[2] ,
         \SB3_31/Component_Function_0/NAND4_in[1] ,
         \SB3_31/Component_Function_0/NAND4_in[0] ,
         \SB3_31/Component_Function_1/NAND4_in[3] ,
         \SB3_31/Component_Function_1/NAND4_in[2] ,
         \SB3_31/Component_Function_1/NAND4_in[1] ,
         \SB3_31/Component_Function_1/NAND4_in[0] ,
         \SB3_31/Component_Function_5/NAND4_in[3] ,
         \SB3_31/Component_Function_5/NAND4_in[2] ,
         \SB3_31/Component_Function_5/NAND4_in[1] ,
         \SB3_31/Component_Function_5/NAND4_in[0] ,
         \SB4_0/Component_Function_0/NAND4_in[2] ,
         \SB4_0/Component_Function_0/NAND4_in[1] ,
         \SB4_0/Component_Function_0/NAND4_in[0] ,
         \SB4_0/Component_Function_1/NAND4_in[3] ,
         \SB4_0/Component_Function_1/NAND4_in[2] ,
         \SB4_0/Component_Function_1/NAND4_in[1] ,
         \SB4_0/Component_Function_5/NAND4_in[3] ,
         \SB4_0/Component_Function_5/NAND4_in[2] ,
         \SB4_0/Component_Function_5/NAND4_in[1] ,
         \SB4_0/Component_Function_5/NAND4_in[0] ,
         \SB4_1/Component_Function_0/NAND4_in[3] ,
         \SB4_1/Component_Function_0/NAND4_in[2] ,
         \SB4_1/Component_Function_1/NAND4_in[1] ,
         \SB4_1/Component_Function_1/NAND4_in[0] ,
         \SB4_1/Component_Function_5/NAND4_in[3] ,
         \SB4_1/Component_Function_5/NAND4_in[2] ,
         \SB4_1/Component_Function_5/NAND4_in[0] ,
         \SB4_2/Component_Function_0/NAND4_in[2] ,
         \SB4_2/Component_Function_0/NAND4_in[1] ,
         \SB4_2/Component_Function_0/NAND4_in[0] ,
         \SB4_2/Component_Function_1/NAND4_in[2] ,
         \SB4_2/Component_Function_1/NAND4_in[1] ,
         \SB4_2/Component_Function_1/NAND4_in[0] ,
         \SB4_2/Component_Function_5/NAND4_in[3] ,
         \SB4_2/Component_Function_5/NAND4_in[2] ,
         \SB4_2/Component_Function_5/NAND4_in[0] ,
         \SB4_3/Component_Function_0/NAND4_in[3] ,
         \SB4_3/Component_Function_0/NAND4_in[2] ,
         \SB4_3/Component_Function_0/NAND4_in[1] ,
         \SB4_3/Component_Function_1/NAND4_in[3] ,
         \SB4_3/Component_Function_1/NAND4_in[2] ,
         \SB4_3/Component_Function_1/NAND4_in[1] ,
         \SB4_3/Component_Function_1/NAND4_in[0] ,
         \SB4_3/Component_Function_5/NAND4_in[3] ,
         \SB4_3/Component_Function_5/NAND4_in[2] ,
         \SB4_3/Component_Function_5/NAND4_in[1] ,
         \SB4_3/Component_Function_5/NAND4_in[0] ,
         \SB4_4/Component_Function_0/NAND4_in[3] ,
         \SB4_4/Component_Function_0/NAND4_in[2] ,
         \SB4_4/Component_Function_0/NAND4_in[1] ,
         \SB4_4/Component_Function_0/NAND4_in[0] ,
         \SB4_4/Component_Function_1/NAND4_in[2] ,
         \SB4_4/Component_Function_1/NAND4_in[1] ,
         \SB4_4/Component_Function_1/NAND4_in[0] ,
         \SB4_4/Component_Function_5/NAND4_in[3] ,
         \SB4_4/Component_Function_5/NAND4_in[2] ,
         \SB4_4/Component_Function_5/NAND4_in[1] ,
         \SB4_4/Component_Function_5/NAND4_in[0] ,
         \SB4_5/Component_Function_0/NAND4_in[2] ,
         \SB4_5/Component_Function_0/NAND4_in[1] ,
         \SB4_5/Component_Function_0/NAND4_in[0] ,
         \SB4_5/Component_Function_1/NAND4_in[2] ,
         \SB4_5/Component_Function_1/NAND4_in[1] ,
         \SB4_5/Component_Function_1/NAND4_in[0] ,
         \SB4_5/Component_Function_5/NAND4_in[2] ,
         \SB4_5/Component_Function_5/NAND4_in[1] ,
         \SB4_5/Component_Function_5/NAND4_in[0] ,
         \SB4_6/Component_Function_0/NAND4_in[3] ,
         \SB4_6/Component_Function_0/NAND4_in[1] ,
         \SB4_6/Component_Function_0/NAND4_in[0] ,
         \SB4_6/Component_Function_1/NAND4_in[3] ,
         \SB4_6/Component_Function_1/NAND4_in[2] ,
         \SB4_6/Component_Function_1/NAND4_in[1] ,
         \SB4_6/Component_Function_1/NAND4_in[0] ,
         \SB4_6/Component_Function_5/NAND4_in[3] ,
         \SB4_6/Component_Function_5/NAND4_in[2] ,
         \SB4_6/Component_Function_5/NAND4_in[1] ,
         \SB4_6/Component_Function_5/NAND4_in[0] ,
         \SB4_7/Component_Function_0/NAND4_in[3] ,
         \SB4_7/Component_Function_0/NAND4_in[1] ,
         \SB4_7/Component_Function_0/NAND4_in[0] ,
         \SB4_7/Component_Function_1/NAND4_in[3] ,
         \SB4_7/Component_Function_1/NAND4_in[2] ,
         \SB4_7/Component_Function_1/NAND4_in[1] ,
         \SB4_7/Component_Function_1/NAND4_in[0] ,
         \SB4_7/Component_Function_5/NAND4_in[3] ,
         \SB4_7/Component_Function_5/NAND4_in[1] ,
         \SB4_7/Component_Function_5/NAND4_in[0] ,
         \SB4_8/Component_Function_0/NAND4_in[3] ,
         \SB4_8/Component_Function_0/NAND4_in[2] ,
         \SB4_8/Component_Function_0/NAND4_in[1] ,
         \SB4_8/Component_Function_0/NAND4_in[0] ,
         \SB4_8/Component_Function_1/NAND4_in[3] ,
         \SB4_8/Component_Function_1/NAND4_in[2] ,
         \SB4_8/Component_Function_1/NAND4_in[1] ,
         \SB4_8/Component_Function_5/NAND4_in[2] ,
         \SB4_8/Component_Function_5/NAND4_in[1] ,
         \SB4_8/Component_Function_5/NAND4_in[0] ,
         \SB4_9/Component_Function_0/NAND4_in[3] ,
         \SB4_9/Component_Function_0/NAND4_in[2] ,
         \SB4_9/Component_Function_0/NAND4_in[1] ,
         \SB4_9/Component_Function_1/NAND4_in[1] ,
         \SB4_9/Component_Function_1/NAND4_in[0] ,
         \SB4_9/Component_Function_5/NAND4_in[3] ,
         \SB4_9/Component_Function_5/NAND4_in[2] ,
         \SB4_9/Component_Function_5/NAND4_in[1] ,
         \SB4_9/Component_Function_5/NAND4_in[0] ,
         \SB4_10/Component_Function_0/NAND4_in[2] ,
         \SB4_10/Component_Function_0/NAND4_in[1] ,
         \SB4_10/Component_Function_0/NAND4_in[0] ,
         \SB4_10/Component_Function_1/NAND4_in[3] ,
         \SB4_10/Component_Function_1/NAND4_in[2] ,
         \SB4_10/Component_Function_1/NAND4_in[1] ,
         \SB4_10/Component_Function_5/NAND4_in[2] ,
         \SB4_10/Component_Function_5/NAND4_in[1] ,
         \SB4_10/Component_Function_5/NAND4_in[0] ,
         \SB4_11/Component_Function_0/NAND4_in[3] ,
         \SB4_11/Component_Function_0/NAND4_in[2] ,
         \SB4_11/Component_Function_0/NAND4_in[1] ,
         \SB4_11/Component_Function_1/NAND4_in[3] ,
         \SB4_11/Component_Function_1/NAND4_in[1] ,
         \SB4_11/Component_Function_5/NAND4_in[2] ,
         \SB4_11/Component_Function_5/NAND4_in[1] ,
         \SB4_11/Component_Function_5/NAND4_in[0] ,
         \SB4_12/Component_Function_0/NAND4_in[2] ,
         \SB4_12/Component_Function_0/NAND4_in[1] ,
         \SB4_12/Component_Function_1/NAND4_in[2] ,
         \SB4_12/Component_Function_1/NAND4_in[1] ,
         \SB4_12/Component_Function_1/NAND4_in[0] ,
         \SB4_12/Component_Function_5/NAND4_in[3] ,
         \SB4_12/Component_Function_5/NAND4_in[1] ,
         \SB4_13/Component_Function_0/NAND4_in[2] ,
         \SB4_13/Component_Function_0/NAND4_in[1] ,
         \SB4_13/Component_Function_0/NAND4_in[0] ,
         \SB4_13/Component_Function_1/NAND4_in[2] ,
         \SB4_13/Component_Function_1/NAND4_in[1] ,
         \SB4_13/Component_Function_5/NAND4_in[3] ,
         \SB4_13/Component_Function_5/NAND4_in[2] ,
         \SB4_13/Component_Function_5/NAND4_in[1] ,
         \SB4_13/Component_Function_5/NAND4_in[0] ,
         \SB4_14/Component_Function_0/NAND4_in[3] ,
         \SB4_14/Component_Function_0/NAND4_in[2] ,
         \SB4_14/Component_Function_0/NAND4_in[1] ,
         \SB4_14/Component_Function_1/NAND4_in[3] ,
         \SB4_14/Component_Function_1/NAND4_in[2] ,
         \SB4_14/Component_Function_1/NAND4_in[1] ,
         \SB4_14/Component_Function_1/NAND4_in[0] ,
         \SB4_14/Component_Function_5/NAND4_in[2] ,
         \SB4_14/Component_Function_5/NAND4_in[1] ,
         \SB4_14/Component_Function_5/NAND4_in[0] ,
         \SB4_15/Component_Function_0/NAND4_in[3] ,
         \SB4_15/Component_Function_0/NAND4_in[2] ,
         \SB4_15/Component_Function_0/NAND4_in[1] ,
         \SB4_15/Component_Function_1/NAND4_in[2] ,
         \SB4_15/Component_Function_1/NAND4_in[1] ,
         \SB4_15/Component_Function_1/NAND4_in[0] ,
         \SB4_15/Component_Function_5/NAND4_in[3] ,
         \SB4_15/Component_Function_5/NAND4_in[2] ,
         \SB4_15/Component_Function_5/NAND4_in[1] ,
         \SB4_15/Component_Function_5/NAND4_in[0] ,
         \SB4_16/Component_Function_0/NAND4_in[2] ,
         \SB4_16/Component_Function_0/NAND4_in[1] ,
         \SB4_16/Component_Function_1/NAND4_in[3] ,
         \SB4_16/Component_Function_1/NAND4_in[2] ,
         \SB4_16/Component_Function_1/NAND4_in[1] ,
         \SB4_16/Component_Function_1/NAND4_in[0] ,
         \SB4_16/Component_Function_5/NAND4_in[1] ,
         \SB4_16/Component_Function_5/NAND4_in[0] ,
         \SB4_17/Component_Function_0/NAND4_in[2] ,
         \SB4_17/Component_Function_0/NAND4_in[1] ,
         \SB4_17/Component_Function_0/NAND4_in[0] ,
         \SB4_17/Component_Function_1/NAND4_in[3] ,
         \SB4_17/Component_Function_1/NAND4_in[2] ,
         \SB4_17/Component_Function_1/NAND4_in[1] ,
         \SB4_17/Component_Function_1/NAND4_in[0] ,
         \SB4_17/Component_Function_5/NAND4_in[1] ,
         \SB4_17/Component_Function_5/NAND4_in[0] ,
         \SB4_18/Component_Function_0/NAND4_in[3] ,
         \SB4_18/Component_Function_0/NAND4_in[1] ,
         \SB4_18/Component_Function_0/NAND4_in[0] ,
         \SB4_18/Component_Function_1/NAND4_in[3] ,
         \SB4_18/Component_Function_1/NAND4_in[1] ,
         \SB4_18/Component_Function_1/NAND4_in[0] ,
         \SB4_18/Component_Function_5/NAND4_in[2] ,
         \SB4_19/Component_Function_0/NAND4_in[2] ,
         \SB4_19/Component_Function_0/NAND4_in[1] ,
         \SB4_19/Component_Function_0/NAND4_in[0] ,
         \SB4_19/Component_Function_1/NAND4_in[3] ,
         \SB4_19/Component_Function_1/NAND4_in[2] ,
         \SB4_19/Component_Function_1/NAND4_in[1] ,
         \SB4_19/Component_Function_1/NAND4_in[0] ,
         \SB4_19/Component_Function_5/NAND4_in[3] ,
         \SB4_19/Component_Function_5/NAND4_in[2] ,
         \SB4_19/Component_Function_5/NAND4_in[1] ,
         \SB4_19/Component_Function_5/NAND4_in[0] ,
         \SB4_20/Component_Function_0/NAND4_in[3] ,
         \SB4_20/Component_Function_0/NAND4_in[2] ,
         \SB4_20/Component_Function_0/NAND4_in[1] ,
         \SB4_20/Component_Function_0/NAND4_in[0] ,
         \SB4_20/Component_Function_1/NAND4_in[3] ,
         \SB4_20/Component_Function_1/NAND4_in[2] ,
         \SB4_20/Component_Function_1/NAND4_in[1] ,
         \SB4_20/Component_Function_1/NAND4_in[0] ,
         \SB4_20/Component_Function_5/NAND4_in[3] ,
         \SB4_20/Component_Function_5/NAND4_in[2] ,
         \SB4_20/Component_Function_5/NAND4_in[0] ,
         \SB4_21/Component_Function_0/NAND4_in[3] ,
         \SB4_21/Component_Function_0/NAND4_in[2] ,
         \SB4_21/Component_Function_1/NAND4_in[3] ,
         \SB4_21/Component_Function_1/NAND4_in[2] ,
         \SB4_21/Component_Function_1/NAND4_in[1] ,
         \SB4_21/Component_Function_1/NAND4_in[0] ,
         \SB4_21/Component_Function_5/NAND4_in[3] ,
         \SB4_21/Component_Function_5/NAND4_in[2] ,
         \SB4_21/Component_Function_5/NAND4_in[1] ,
         \SB4_21/Component_Function_5/NAND4_in[0] ,
         \SB4_22/Component_Function_0/NAND4_in[3] ,
         \SB4_22/Component_Function_0/NAND4_in[2] ,
         \SB4_22/Component_Function_0/NAND4_in[1] ,
         \SB4_22/Component_Function_0/NAND4_in[0] ,
         \SB4_22/Component_Function_1/NAND4_in[3] ,
         \SB4_22/Component_Function_1/NAND4_in[1] ,
         \SB4_22/Component_Function_1/NAND4_in[0] ,
         \SB4_22/Component_Function_5/NAND4_in[2] ,
         \SB4_22/Component_Function_5/NAND4_in[1] ,
         \SB4_22/Component_Function_5/NAND4_in[0] ,
         \SB4_23/Component_Function_0/NAND4_in[3] ,
         \SB4_23/Component_Function_0/NAND4_in[2] ,
         \SB4_23/Component_Function_0/NAND4_in[1] ,
         \SB4_23/Component_Function_0/NAND4_in[0] ,
         \SB4_23/Component_Function_1/NAND4_in[2] ,
         \SB4_23/Component_Function_1/NAND4_in[1] ,
         \SB4_23/Component_Function_5/NAND4_in[2] ,
         \SB4_23/Component_Function_5/NAND4_in[1] ,
         \SB4_23/Component_Function_5/NAND4_in[0] ,
         \SB4_24/Component_Function_0/NAND4_in[2] ,
         \SB4_24/Component_Function_0/NAND4_in[1] ,
         \SB4_24/Component_Function_0/NAND4_in[0] ,
         \SB4_24/Component_Function_1/NAND4_in[3] ,
         \SB4_24/Component_Function_1/NAND4_in[2] ,
         \SB4_24/Component_Function_1/NAND4_in[1] ,
         \SB4_24/Component_Function_1/NAND4_in[0] ,
         \SB4_24/Component_Function_5/NAND4_in[2] ,
         \SB4_24/Component_Function_5/NAND4_in[1] ,
         \SB4_24/Component_Function_5/NAND4_in[0] ,
         \SB4_25/Component_Function_0/NAND4_in[3] ,
         \SB4_25/Component_Function_0/NAND4_in[2] ,
         \SB4_25/Component_Function_0/NAND4_in[1] ,
         \SB4_25/Component_Function_1/NAND4_in[3] ,
         \SB4_25/Component_Function_1/NAND4_in[1] ,
         \SB4_25/Component_Function_5/NAND4_in[3] ,
         \SB4_25/Component_Function_5/NAND4_in[2] ,
         \SB4_25/Component_Function_5/NAND4_in[1] ,
         \SB4_25/Component_Function_5/NAND4_in[0] ,
         \SB4_26/Component_Function_0/NAND4_in[3] ,
         \SB4_26/Component_Function_0/NAND4_in[1] ,
         \SB4_26/Component_Function_1/NAND4_in[3] ,
         \SB4_26/Component_Function_1/NAND4_in[2] ,
         \SB4_26/Component_Function_1/NAND4_in[1] ,
         \SB4_26/Component_Function_1/NAND4_in[0] ,
         \SB4_26/Component_Function_5/NAND4_in[2] ,
         \SB4_26/Component_Function_5/NAND4_in[1] ,
         \SB4_26/Component_Function_5/NAND4_in[0] ,
         \SB4_27/Component_Function_0/NAND4_in[2] ,
         \SB4_27/Component_Function_0/NAND4_in[1] ,
         \SB4_27/Component_Function_1/NAND4_in[3] ,
         \SB4_27/Component_Function_1/NAND4_in[2] ,
         \SB4_27/Component_Function_1/NAND4_in[1] ,
         \SB4_27/Component_Function_5/NAND4_in[3] ,
         \SB4_27/Component_Function_5/NAND4_in[1] ,
         \SB4_27/Component_Function_5/NAND4_in[0] ,
         \SB4_28/Component_Function_0/NAND4_in[0] ,
         \SB4_28/Component_Function_1/NAND4_in[3] ,
         \SB4_28/Component_Function_1/NAND4_in[2] ,
         \SB4_28/Component_Function_1/NAND4_in[1] ,
         \SB4_28/Component_Function_5/NAND4_in[2] ,
         \SB4_28/Component_Function_5/NAND4_in[1] ,
         \SB4_28/Component_Function_5/NAND4_in[0] ,
         \SB4_29/Component_Function_1/NAND4_in[1] ,
         \SB4_29/Component_Function_1/NAND4_in[0] ,
         \SB4_29/Component_Function_5/NAND4_in[2] ,
         \SB4_29/Component_Function_5/NAND4_in[0] ,
         \SB4_30/Component_Function_0/NAND4_in[2] ,
         \SB4_30/Component_Function_0/NAND4_in[1] ,
         \SB4_30/Component_Function_1/NAND4_in[3] ,
         \SB4_30/Component_Function_1/NAND4_in[2] ,
         \SB4_30/Component_Function_1/NAND4_in[1] ,
         \SB4_30/Component_Function_1/NAND4_in[0] ,
         \SB4_30/Component_Function_5/NAND4_in[3] ,
         \SB4_30/Component_Function_5/NAND4_in[2] ,
         \SB4_30/Component_Function_5/NAND4_in[0] ,
         \SB4_31/Component_Function_0/NAND4_in[3] ,
         \SB4_31/Component_Function_0/NAND4_in[2] ,
         \SB4_31/Component_Function_0/NAND4_in[1] ,
         \SB4_31/Component_Function_0/NAND4_in[0] ,
         \SB4_31/Component_Function_1/NAND4_in[3] ,
         \SB4_31/Component_Function_1/NAND4_in[2] ,
         \SB4_31/Component_Function_1/NAND4_in[1] ,
         \SB4_31/Component_Function_1/NAND4_in[0] ,
         \SB4_31/Component_Function_5/NAND4_in[2] , n1, n4, n8, n11, n12, n18,
         n19, n22, n23, n35, n37, n41, n43, n44, n49, n54, n62, n69, n77, n78,
         n82, n85, n87, n88, n91, n96, n99, n102, n110, n111, n112, n116, n119,
         n120, n123, n124, n139, n142, n145, n149, n150, n151, n155, n161,
         n164, n167, n168, n171, n174, n175, n179, n2, n3, n5, n6, n7, n9, n10,
         n13, n14, n15, n16, n17, n20, n21, n24, n25, n26, n27, n28, n29, n30,
         n31, n33, n34, n36, n38, n39, n40, n42, n45, n46, n47, n48, n50, n51,
         n52, n53, n55, n56, n57, n58, n59, n60, n61, n63, n64, n65, n66, n67,
         n68, n70, n71, n72, n73, n74, n75, n76, n79, n80, n81, n83, n84, n86,
         n89, n90, n92, n93, n94, n95, n97, n98, n100, n101, n103, n104, n105,
         n106, n107, n108, n109, n113, n114, n115, n117, n118, n121, n122,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n140, n141, n143, n144, n146, n147, n148, n152,
         n153, n154, n156, n158, n159, n160, n162, n163, n165, n166, n169,
         n170, n172, n173, n176, n177, n178, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n569, n570,
         n571, n573, n575, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n590, n593, n597, n599, n606, n607, n611, n612, n613, n616,
         n618, n622, n623, n624, n625, n626, n627, n629, n632, n634, n636,
         n639, n641, n642, n643, n649, n650, n652, n654, n656, n657, n659,
         n660, n661, n667, n669, n670, n671, n672, n673, n674, n675, n679,
         n681, n683, n691, n693, n699, n700, n701, n705, n706, n708, n711,
         n712, n715, n719, n721, n722, n724, n725, n727, n729, n731, n733,
         n735, n737, n739, n740, n741, n744, n747, n756, n757, n759, n760,
         n761, n762, n763, n765, n767, n768, n774, n775, n780, n782, n784,
         n785, n790, n792, n793, n795, n796, n799, n800, n804, n805, n806,
         n807, n809, n817, n820, n821, n822, n823, n826, n827, n828, n832,
         n833, n834, n836, n838, n841, n842, n845, n846, n847, n855, n856,
         n858, n860, n864, n865, n868, n869, n870, n873, n874, n876, n877,
         n878, n880, n882, n884, n885, n886, n887, n890, n893, n894, n899,
         n901, n904, n905, n909, n910, n911, n913, n914, n918, n923, n924,
         n926, n927, n930, n933, n935, n937, n940, n941, n942, n943, n946,
         n947, n949, n950, n951, n952, n953, n954, n957, n959, n960, n962,
         n964, n965, n968, n970, n971, n976, n977, n987, n990, n998, n1001,
         n1002, n1003, n1004, n1006, n1009, n1010, n1013, n1014, n1015, n1016,
         n1017, n1020, n1021, n1023, n1025, n1030, n1031, n1037, n1040, n1042,
         n1043, n1044, n1046, n1048, n1049, n1050, n1052, n1053, n1054, n1058,
         n1059, n1060, n1061, n1062, n1063, n1066, n1071, n1076, n1077, n1078,
         n1079, n1080, n1082, n1086, n1088, n1091, n1092, n1095, n1096, n1097,
         n1099, n1103, n1105, n1106, n1109, n1110, n1114, n1115, n1116, n1117,
         n1120, n1121, n1124, n1125, n1127, n1129, n1130, n1131, n1132, n1133,
         n1138, n1142, n1144, n1146, n1148, n1149, n1151, n1152, n1153, n1156,
         n1157, n1158, n1159, n1161, n1163, n1164, n1167, n1169, n1171, n1174,
         n1176, n1177, n1182, n1183, n1184, n1186, n1189, n1190, n1192, n1195,
         n1196, n1198, n1199, n1201, n1203, n1205, n1206, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1217, n1220, n1221, n1225, n1228, n1230,
         n1232, n1235, n1236, n1238, n1239, n1241, n1245, n1249, n1250, n1251,
         n1255, n1257, n1259, n1260, n1261, n1263, n1264, n1265, n1269, n1270,
         n1271, n1272, n1275, n1277, n1278, n1279, n1280, n1284, n1285, n1286,
         n1287, n1290, n1292, n1293, n1294, n1295, n1297, n1298, n1299, n1302,
         n1303, n1306, n1307, n1310, n1311, n1312, n1313, n1314, n1315, n1317,
         n1318, n1319, n1320, n1321, n1322, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1333, n1334, n1337, n1340, n1341, n1342, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1353, n1354, n1355,
         n1358, n1361, n1362, n1365, n1367, n1370, n1371, n1372, n1373, n1375,
         n1376, n1377, n1379, n1381, n1383, n1384, n1385, n1386, n1388, n1389,
         n1390, n1392, n1393, n1394, n1396, n1400, n1401, n1402, n1403, n1404,
         n1405, n1407, n1408, n1409, n1411, n1412, n1413, n1414, n1416, n1417,
         n1419, n1420, n1421, n1422, n1424, n1425, n1426, n1427, n1429, n1431,
         n1433, n1434, n1436, n1437, n1438, n1439, n1440, n1443, n1444, n1445,
         n1447, n1450, n1451, n1452, n1454, n1457, n1458, n1463, n1464, n1465,
         n1466, n1467, n1469, n1472, n1473, n1477, n1478, n1481, n1482, n1483,
         n1484, n1486, n1488, n1490, n1491, n1493, n1494, n1495, n1496, n1497,
         n1498, n1500, n1501, n1506, n1508, n1511, n1514, n1517, n1518, n1522,
         n1523, n1524, n1527, n1528, n1529, n1531, n1532, n1536, n1537, n1538,
         n1539, n1540, n1541, n1544, n1546, n1547, n1548, n1549, n1550, n1551,
         n1553, n1555, n1556, n1557, n1558, n1560, n1561, n1562, n1563, n1567,
         n1568, n1569, n1570, n1571, n1574, n1575, n1576, n1577, n1578, n1579,
         n1581, n1582, n1584, n1589, n1590, n1593, n1594, n1595, n1597, n1598,
         n1599, n1600, n1601, n1603, n1604, n1608, n1609, n1610, n1613, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1625, n1626, n1627, n1628,
         n1632, n1634, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1678, n1679,
         n1680, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1693, n1694, n1695, n1696, n1697, n1699, n1701, n1702, n1703, n1704,
         n1706, n1707, n1708, n1709, n1710, n1712, n1713, n1715, n1717, n1718,
         n1721, n1724, n1729, n1730, n1733, n1734, n1735, n1736, n1737, n1739,
         n1740, n1741, n1742, n1743, n1745, n1746, n1747, n1748, n1750, n1751,
         n1752, n1754, n1755, n1756, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1773, n1775, n1777, n1783, n1784, n1785,
         n1788, n1789, n1790, n1793, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1804, n1805, n1808, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1819, n1820, n1821, n1822, n1823, n1826, n1827, n1828,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1842, n1844, n1846, n1847, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1860, n1861, n1863, n1864, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1877, n1878, n1880, n1881,
         n1882, n1884, n1885, n1886, n1888, n1890, n1891, n1892, n1894, n1895,
         n1896, n1903, n1905, n1906, n1907, n1908, n1909, n1911, n1912, n1913,
         n1916, n1917, n1918, n1921, n1924, n1925, n1926, n1928, n1931, n1932,
         n1933, n1935, n1936, n1937, n1939, n1940, n1944, n1945, n1946, n1948,
         n1949, n1950, n1951, n1955, n1956, n1958, n1960, n1962, n1964, n1967,
         n1969, n1971, n1976, n1977, n1978, n1979, n1980, n1982, n1984, n1986,
         n1987, n1988, n1989, n1990, n1992, n1993, n1995, n1998, n1999, n2000,
         n2001, n2003, n2004, n2005, n2007, n2008, n2009, n2010, n2011, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2021, n2022, n2023, n2025,
         n2026, n2027, n2028, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2043, n2045, n2046, n2047, n2049, n2050,
         n2051, n2053, n2054, n2055, n2056, n2057, n2060, n2062, n2063, n2067,
         n2069, n2070, n2071, n2072, n2073, n2074, n2076, n2078, n2079, n2080,
         n2081, n2083, n2084, n2086, n2087, n2088, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2106,
         n2108, n2109, n2110, n2112, n2113, n2115, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2125, n2126, n2128, n2131, n2132, n2133, n2134,
         n2135, n2137, n2140, n2142, n2143, n2145, n2149, n2150, n2152, n2153,
         n2154, n2155, n2157, n2158, n2161, n2162, n2164, n2168, n2169, n2170,
         n2171, n2172, n2174, n2176, n2177, n2178, n2179, n2180, n2181, n2184,
         n2185, n2186, n2189, n2190, n2191, n2192, n2193, n2195, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2207, n2208, n2209, n2210,
         n2211, n2212, n2215, n2217, n2218, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2230, n2233, n2234, n2235, n2236, n2237, n2239,
         n2240, n2241, n2243, n2244, n2246, n2248, n2249, n2250, n2251, n2253,
         n2255, n2256, n2257, n2258, n2260, n2261, n2263, n2266, n2267, n2268,
         n2273, n2274, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2291, n2292, n2293, n2294, n2295, n2297, n2298,
         n2299, n2300, n2301, n2303, n2307, n2308, n2309, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2325, n2327, n2329,
         n2330, n2333, n2334, n2338, n2339, n2342, n2343, n2344, n2346, n2348,
         n2351, n2352, n2353, n2355, n2356, n2358, n2359, n2362, n2363, n2364,
         n2366, n2367, n2369, n2371, n2372, n2373, n2375, n2379, n2382, n2383,
         n2385, n2387, n2388, n2389, n2390, n2391, n2392, n2394, n2397, n2401,
         n2402, n2403, n2404, n2405, n2406, n2408, n2409, n2410, n2411, n2412,
         n2414, n2415, n2416, n2417, n2418, n2419, n2421, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2442, n2444, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2459, n2460,
         n2461, n2462, n2463, n2465, n2467, n2469, n2470, n2472, n2473, n2475,
         n2476, n2478, n2480, n2481, n2482, n2483, n2484, n2492, n2493, n2495,
         n2496, n2497, n2498, n2499, n2500, n2502, n2509, n2510, n2511, n2512,
         n2518, n2519, n2520, n2522, n2523, n2524, n2525, n2526, n2527, n2529,
         n2530, n2531, n2534, n2535, n2536, n2539, n2540, n2545, n2546, n2547,
         n2548, n2551, n2553, n2554, n2555, n2556, n2557, n2560, n2561, n2562,
         n2563, n2564, n2565, n2567, n2568, n2569, n2572, n2574, n2575, n2576,
         n2577, n2578, n2581, n2582, n2583, n2584, n2587, n2593, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2605, n2606, n2607, n2609,
         n2610, n2611, n2612, n2613, n2615, n2616, n2617, n2618, n2620, n2621,
         n2622, n2623, n2624, n2626, n2627, n2628, n2629, n2630, n2632, n2633,
         n2634, n2635, n2636, n2637, n2639, n2640, n2644, n2646, n2647, n2650,
         n2651, n2652, n2655, n2657, n2658, n2660, n2661, n2663, n2664, n2665,
         n2666, n2667, n2669, n2670, n2671, n2673, n2675, n2677, n2678, n2679,
         n2680, n2681, n2682, n2686, n2687, n2689, n2690, n2691, n2692, n2693,
         n2695, n2700, n2703, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2715, n2718, n2720, n2723, n2724, n2725, n2726, n2727,
         n2728, n2730, n2735, n2738, n2739, n2742, n2743, n2744, n2745, n2746,
         n2749, n2750, n2751, n2752, n2753, n2756, n2757, n2759, n2761, n2762,
         n2763, n2765, n2766, n2768, n2769, n2773, n2774, n2775, n2776, n2777,
         n2778, n2780, n2781, n2782, n2783, n2784, n2785, n2789, n2790, n2792,
         n2794, n2795, n2796, n2798, n2799, n2801, n2802, n2803, n2805, n2806,
         n2807, n2808, n2809, n2812, n2813, n2815, n2816, n2818, n2819, n2820,
         n2823, n2827, n2828, n2829, n2831, n2833, n2834, n2835, n2837, n2839,
         n2842, n2843, n2844, n2845, n2846, n2847, n2850, n2852, n2853, n2854,
         n2856, n2858, n2862, n2863, n2864, n2865, n2867, n2868, n2870, n2875,
         n2876, n2877, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2889, n2890, n2891, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2901, n2902, n2903, n2904, n2905, n2906, n2908, n2909, n2910, n2911,
         n2913, n2914, n2917, n2920, n2922, n2923, n2924, n2925, n2927, n2930,
         n2931, n2933, n2934, n2935, n2937, n2939, n2940, n2942, n2943, n2945,
         n2947, n2948, n2949, n2951, n2956, n2958, n2960, n2962, n2964, n2965,
         n2967, n2970, n2972, n2973, n2974, n2975, n2976, n2979, n2983, n2984,
         n2985, n2987, n2988, n2989, n2991, n2993, n2994, n2995, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3008, n3009,
         n3010, n3011, n3012, n3015, n3016, n3018, n3023, n3026, n3028, n3029,
         n3031, n3032, n3033, n3034, n3035, n3037, n3039, n3040, n3041, n3042,
         n3049, n3050, n3051, n3052, n3053, n3054, n3057, n3058, n3059, n3065,
         n3066, n3068, n3069, n3070, n3071, n3072, n3073, n3075, n3076, n3077,
         n3079, n3080, n3081, n3089, n3090, n3091, n3092, n3097, n3098, n3099,
         n3100, n3101, n3102, n3105, n3106, n3109, n3110, n3112, n3113, n3114,
         n3118, n3119, n3120, n3122, n3124, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3134, n3137, n3140, n3141, n3143, n3144, n3145, n3147,
         n3148, n3149, n3150, n3152, n3154, n3155, n3156, n3157, n3158, n3161,
         n3162, n3165, n3166, n3168, n3171, n3172, n3173, n3175, n3176, n3177,
         n3178, n3179, n3180, n3183, n3184, n3185, n3189, n3190, n3191, n3192,
         n3195, n3196, n3198, n3201, n3202, n3203, n3207, n3208, n3209, n3211,
         n3212, n3213, n3214, n3215, n3219, n3220, n3222, n3224, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3236, n3239, n3240, n3243,
         n3244, n3247, n3248, n3249, n3251, n3255, n3256, n3258, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3276, n3277, n3278, n3279, n3280, n3282, n3283, n3285, n3286, n3287,
         n3288, n3289, n3291, n3292, n3293, n3294, n3295, n3297, n3300, n3302,
         n3303, n3305, n3306, n3307, n3308, n3309, n3312, n3313, n3314, n3315,
         n3316, n3317, n3320, n3322, n3323, n3327, n3329, n3331, n3332, n3333,
         n3334, n3335, n3338, n3340, n3341, n3342, n3344, n3345, n3347, n3348,
         n3349, n3350, n3353, n3356, n3357, n3360, n3364, n3366, n3367, n3368,
         n3369, n3373, n3374, n3375, n3378, n3381, n3382, n3385, n3386, n3388,
         n3389, n3390, n3392, n3393, n3394, n3395, n3396, n3397, n3399, n3400,
         n3401, n3402, n3404, n3405, n3406, n3407, n3409, n3410, n3411, n3412,
         n3413, n3415, n3416, n3419, n3420, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3430, n3431, n3433, n3434, n3435, n3437, n3439, n3440,
         n3442, n3443, n3445, n3447, n3448, n3450, n3451, n3452, n3454, n3456,
         n3461, n3462, n3463, n3464, n3465, n3466, n3468, n3469, n3471, n3472,
         n3473, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3490, n3492, n3494, n3495, n3496, n3497, n3499,
         n3500, n3501, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3512, n3513, n3514, n3516, n3517, n3520, n3522, n3524, n3525, n3526,
         n3528, n3529, n3531, n3532, n3535, n3536, n3540, n3541, n3543, n3544,
         n3545, n3546, n3547, n3551, n3555, n3556, n3559, n3561, n3564, n3565,
         n3568, n3569, n3572, n3573, n3574, n3575, n3577, n3584, n3585, n3587,
         n3589, n3590, n3591, n3596, n3597, n3602, n3607, n3608, n3610, n3611,
         n3612, n3614, n3615, n3616, n3617, n3618, n3620, n3621, n3622, n3626,
         n3627, n3631, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3650, n3651,
         n3652, n3653, n3654, n3655, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3698, n3699, n3701, n3702, n3704, n3708, n3710, n3711, n3712,
         n3713, n3714, n3715, n3717, n3718, n3723, n3724, n3725, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3756, n3757, n3758, n3759, n3760,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3786, n3787, n3788, n3790, n3791, n3792, n3793,
         n3794, n3796, n3797, n3798, n3799, n3801, n3803, n3805, n3806, n3808,
         n3809, n3810, n3811, n3813, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3825, n3826, n3828, n3829, n3830, n3831, n3833, n3834, n3836,
         n3837, n3838, n3839, n3840, n3842, n3844, n3845, n3846, n3847, n3848,
         n3849, n3852, n3854, n3855, n3856, n3857, n3858, n3860, n3861, n3863,
         n3864, n3865, n3868, n3869, n3870, n3871, n3872, n3874, n3876, n3877,
         n3880, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3908, n3910, n3912, n3913, n3914, n3916, n3917, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3929, n3931,
         n3932, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3952, n3953, n3954,
         n3955, n3956, n3957, n3960, n3961, n3962, n3963, n3964, n3968, n3969,
         n3970, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3984, n3987, n3988, n3990, n3991, n3992, n3993, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4006, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4021, n4022, n4023, n4024, n4026, n4027, n4028, n4029, n4032, n4033,
         n4034, n4035, n4036, n4039, n4041, n4044, n4047, n4048, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4063, n4065, n4066, n4067, n4068, n4070, n4071, n4072, n4073, n4075,
         n4076, n4078, n4079, n4080, n4081, n4083, n4084, n4085, n4086, n4087,
         n4089, n4090, n4091, n4092, n4093, n4095, n4096, n4098, n4101, n4104,
         n4105, n4106, n4107, n4108, n4110, n4111, n4113, n4114, n4115, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4141, n4144, n4145, n4146, n4148, n4149, n4150, n4152, n4154, n4155,
         n4156, n4157, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4169, n4171, n4173, n4174, n4175, n4176, n4177, n4179, n4181, n4182,
         n4183, n4184, n4188, n4189, n4190, n4193, n4195, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4207, n4208, n4210, n4211,
         n4212, n4214, n4216, n4217, n4218, n4221, n4225, n4226, n4227, n4228,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4240, n4241, n4242,
         n4243, n4244, n4246, n4247, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4258, n4259, n4260, n4261, n4263, n4264, n4266, n4268, n4271,
         n4272, n4273, n4274, n4276, n4277, n4279, n4281, n4282, n4283, n4284,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4296, n4298,
         n4299, n4300, n4301, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4311, n4312, n4313, n4314, n4315, n4316, n4318, n4319, n4322, n4323,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4334, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4347, n4348,
         n4349, n4350, n4351, n4352, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4366, n4367, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4381, n4382, n4383, n4384, n4385, n4387, n4388,
         n4389, n4391, n4392, n4393, n4394, n4395, n4396, n4398, n4400, n4401,
         n4402, n4403, n4405, n4406, n4407, n4408, n4409, n4410, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4421, n4422, n4423, n4425,
         n4426, n4427, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4452, n4454, n4455, n4456, n4457, n4459, n4460, n4461, n4462,
         n4463, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4474, n4476,
         n4477, n4480, n4482, n4483, n4485, n4486, n4487, n4488, n4489, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4501, n4504,
         n4506, n4507, n4510, n4511, n4512, n4514, n4515, n4517, n4518, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4575, n4576, n4577, n4578, n4579, n4581, n4582, n4583, n4584, n4585,
         n4586, n4589, n4591, n4592, n4593, n4597, n4598, n4603, n4604, n4605,
         n4607, n4608, n4609, n4610, n4611, n4613, n4614, n4616, n4617, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4635, n4636, n4637, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4650, n4651, n4652, n4654, n4655,
         n4656, n4657, n4658, n4660, n4661, n4662, n4663, n4664, n4665, n4667,
         n4668, n4669, n4670, n4671, n4672, n4674, n4675, n4676, n4679, n4680,
         n4681, n4682, n4683, n4685, n4687, n4688, n4690, n4691, n4692, n4693,
         n4694, n4697, n4698, n4700, n4701, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4722, n4724, n4725, n4726, n4727, n4728, n4730, n4732, n4733,
         n4734, n4736, n4739, n4740, n4742, n4743, n4744, n4745, n4746, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540;

  XOR2_X1 \MC_ARK_ARC_1_0/X7_31_5  ( .A1(\MC_ARK_ARC_1_0/temp5[0] ), .A2(
        \MC_ARK_ARC_1_0/temp6[0] ), .Z(\MC_ARK_ARC_1_0/buf_output[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_31_5  ( .A1(\MC_ARK_ARC_1_0/temp3[0] ), .A2(
        \MC_ARK_ARC_1_0/temp4[0] ), .Z(\MC_ARK_ARC_1_0/temp6[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_31_5  ( .A1(\MC_ARK_ARC_1_0/temp1[0] ), .A2(
        \MC_ARK_ARC_1_0/temp2[0] ), .Z(\MC_ARK_ARC_1_0/temp5[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_31_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[36] ), 
        .A2(n221), .Z(\MC_ARK_ARC_1_0/temp4[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_31_5  ( .A1(\RI5[0][102] ), .A2(\RI5[0][66] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_31_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[138] ), 
        .A2(\RI5[0][162] ), .Z(\MC_ARK_ARC_1_0/temp2[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_31_5  ( .A1(\RI5[0][0] ), .A2(\RI5[0][186] ), .Z(
        \MC_ARK_ARC_1_0/temp1[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_31_4  ( .A1(\MC_ARK_ARC_1_0/temp6[1] ), .A2(
        \MC_ARK_ARC_1_0/temp5[1] ), .Z(\MC_ARK_ARC_1_0/buf_output[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_31_4  ( .A1(\MC_ARK_ARC_1_0/temp3[1] ), .A2(
        \MC_ARK_ARC_1_0/temp4[1] ), .Z(\MC_ARK_ARC_1_0/temp6[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_31_4  ( .A1(\MC_ARK_ARC_1_0/temp1[1] ), .A2(
        \MC_ARK_ARC_1_0/temp2[1] ), .Z(\MC_ARK_ARC_1_0/temp5[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_31_4  ( .A1(\RI5[0][37] ), .A2(n132), .Z(
        \MC_ARK_ARC_1_0/temp4[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_31_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[67] ), 
        .A2(\RI5[0][103] ), .Z(\MC_ARK_ARC_1_0/temp3[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_31_4  ( .A1(\RI5[0][163] ), .A2(\RI5[0][139] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_31_4  ( .A1(\RI5[0][1] ), .A2(\RI5[0][187] ), .Z(
        \MC_ARK_ARC_1_0/temp1[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_31_3  ( .A1(\RI5[0][38] ), .A2(n84), .Z(
        \MC_ARK_ARC_1_0/temp4[2] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_31_3  ( .A1(\RI5[0][104] ), .A2(\RI5[0][68] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[2] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_31_2  ( .A1(\MC_ARK_ARC_1_0/temp3[3] ), .A2(
        \MC_ARK_ARC_1_0/temp4[3] ), .Z(\MC_ARK_ARC_1_0/temp6[3] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_31_2  ( .A1(\RI5[0][39] ), .A2(n162), .Z(
        \MC_ARK_ARC_1_0/temp4[3] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_31_1  ( .A1(\RI5[0][40] ), .A2(n150), .Z(
        \MC_ARK_ARC_1_0/temp4[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_31_1  ( .A1(\RI5[0][106] ), .A2(\RI5[0][70] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_31_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[166] ), 
        .A2(\RI5[0][142] ), .Z(\MC_ARK_ARC_1_0/temp2[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_31_0  ( .A1(\RI5[0][41] ), .A2(n169), .Z(
        \MC_ARK_ARC_1_0/temp4[5] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_31_0  ( .A1(\RI5[0][71] ), .A2(\RI5[0][107] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[5] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_30_5  ( .A1(\MC_ARK_ARC_1_0/temp5[6] ), .A2(
        \MC_ARK_ARC_1_0/temp6[6] ), .Z(\MC_ARK_ARC_1_0/buf_output[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_30_5  ( .A1(\MC_ARK_ARC_1_0/temp3[6] ), .A2(
        \MC_ARK_ARC_1_0/temp4[6] ), .Z(\MC_ARK_ARC_1_0/temp6[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_30_5  ( .A1(\MC_ARK_ARC_1_0/temp2[6] ), .A2(
        \MC_ARK_ARC_1_0/temp1[6] ), .Z(\MC_ARK_ARC_1_0/temp5[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_30_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[42] ), 
        .A2(n537), .Z(\MC_ARK_ARC_1_0/temp4[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_30_5  ( .A1(\RI5[0][108] ), .A2(\RI5[0][72] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_30_5  ( .A1(\RI5[0][168] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[144] ), .Z(\MC_ARK_ARC_1_0/temp2[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_30_5  ( .A1(\RI5[0][6] ), .A2(\RI5[0][0] ), .Z(
        \MC_ARK_ARC_1_0/temp1[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_30_4  ( .A1(\RI5[0][43] ), .A2(n530), .Z(
        \MC_ARK_ARC_1_0/temp4[7] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_30_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[109] ), 
        .A2(\MC_ARK_ARC_1_0/buf_datainput[73] ), .Z(\MC_ARK_ARC_1_0/temp3[7] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_30_4  ( .A1(\SB2_0_7/buf_output[1] ), .A2(
        \RI5[0][145] ), .Z(\MC_ARK_ARC_1_0/temp2[7] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_30_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[7] ), 
        .A2(\RI5[0][1] ), .Z(\MC_ARK_ARC_1_0/temp1[7] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_30_3  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[44] ), 
        .A2(n524), .Z(\MC_ARK_ARC_1_0/temp4[8] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_30_2  ( .A1(\MC_ARK_ARC_1_0/temp5[9] ), .A2(
        \MC_ARK_ARC_1_0/temp6[9] ), .Z(\MC_ARK_ARC_1_0/buf_output[9] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_30_2  ( .A1(\MC_ARK_ARC_1_0/temp3[9] ), .A2(
        \MC_ARK_ARC_1_0/temp4[9] ), .Z(\MC_ARK_ARC_1_0/temp6[9] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_30_2  ( .A1(\RI5[0][45] ), .A2(n125), .Z(
        \MC_ARK_ARC_1_0/temp4[9] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_30_2  ( .A1(\RI5[0][111] ), .A2(\RI5[0][75] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[9] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_30_1  ( .A1(\MC_ARK_ARC_1_0/temp4[10] ), .A2(
        \MC_ARK_ARC_1_0/temp3[10] ), .Z(\MC_ARK_ARC_1_0/temp6[10] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_30_1  ( .A1(\MC_ARK_ARC_1_0/temp1[10] ), .A2(
        \MC_ARK_ARC_1_0/temp2[10] ), .Z(\MC_ARK_ARC_1_0/temp5[10] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_30_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[46] ), 
        .A2(n177), .Z(\MC_ARK_ARC_1_0/temp4[10] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_30_1  ( .A1(\RI5[0][172] ), .A2(\RI5[0][148] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[10] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_30_1  ( .A1(\RI5[0][10] ), .A2(\RI5[0][4] ), .Z(
        \MC_ARK_ARC_1_0/temp1[10] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_30_0  ( .A1(\MC_ARK_ARC_1_0/temp3[11] ), .A2(
        \MC_ARK_ARC_1_0/temp4[11] ), .Z(\MC_ARK_ARC_1_0/temp6[11] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_30_0  ( .A1(\RI5[0][47] ), .A2(n117), .Z(
        \MC_ARK_ARC_1_0/temp4[11] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_30_0  ( .A1(\RI5[0][173] ), .A2(\RI5[0][149] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[11] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_29_5  ( .A1(\MC_ARK_ARC_1_0/temp5[12] ), .A2(
        \MC_ARK_ARC_1_0/temp6[12] ), .Z(\MC_ARK_ARC_1_0/buf_output[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_29_5  ( .A1(\MC_ARK_ARC_1_0/temp3[12] ), .A2(
        \MC_ARK_ARC_1_0/temp4[12] ), .Z(\MC_ARK_ARC_1_0/temp6[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_29_5  ( .A1(\MC_ARK_ARC_1_0/temp1[12] ), .A2(
        \MC_ARK_ARC_1_0/temp2[12] ), .Z(\MC_ARK_ARC_1_0/temp5[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_29_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[48] ), 
        .A2(n507), .Z(\MC_ARK_ARC_1_0/temp4[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_29_5  ( .A1(\RI5[0][174] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[150] ), .Z(\MC_ARK_ARC_1_0/temp2[12] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_29_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[12] ), 
        .A2(\RI5[0][6] ), .Z(\MC_ARK_ARC_1_0/temp1[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_29_4  ( .A1(\MC_ARK_ARC_1_0/temp5[13] ), .A2(
        \MC_ARK_ARC_1_0/temp6[13] ), .Z(\MC_ARK_ARC_1_0/buf_output[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_29_4  ( .A1(\MC_ARK_ARC_1_0/temp1[13] ), .A2(
        \MC_ARK_ARC_1_0/temp2[13] ), .Z(\MC_ARK_ARC_1_0/temp5[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_29_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[49] ), 
        .A2(n91), .Z(\MC_ARK_ARC_1_0/temp4[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_29_4  ( .A1(\RI5[0][175] ), .A2(\RI5[0][151] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_29_3  ( .A1(\MC_ARK_ARC_1_0/temp5[14] ), .A2(
        \MC_ARK_ARC_1_0/temp6[14] ), .Z(\MC_ARK_ARC_1_0/buf_output[14] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_29_3  ( .A1(\MC_ARK_ARC_1_0/temp3[14] ), .A2(
        \MC_ARK_ARC_1_0/temp4[14] ), .Z(\MC_ARK_ARC_1_0/temp6[14] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_29_3  ( .A1(\MC_ARK_ARC_1_0/temp2[14] ), .A2(
        \MC_ARK_ARC_1_0/temp1[14] ), .Z(\MC_ARK_ARC_1_0/temp5[14] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_29_3  ( .A1(\RI5[0][50] ), .A2(n209), .Z(
        \MC_ARK_ARC_1_0/temp4[14] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_29_2  ( .A1(\RI5[0][177] ), .A2(\RI5[0][153] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[15] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_29_1  ( .A1(\RI5[0][52] ), .A2(n488), .Z(
        \MC_ARK_ARC_1_0/temp4[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_29_1  ( .A1(\RI5[0][118] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[82] ), .Z(\MC_ARK_ARC_1_0/temp3[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_29_0  ( .A1(\RI5[0][53] ), .A2(n482), .Z(
        \MC_ARK_ARC_1_0/temp4[17] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_29_0  ( .A1(\RI5[0][83] ), .A2(\RI5[0][119] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[17] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_29_0  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[155] ), 
        .A2(\MC_ARK_ARC_1_0/buf_datainput[179] ), .Z(
        \MC_ARK_ARC_1_0/temp2[17] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_29_0  ( .A1(\RI5[0][11] ), .A2(\RI5[0][17] ), .Z(
        \MC_ARK_ARC_1_0/temp1[17] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_28_5  ( .A1(\MC_ARK_ARC_1_0/temp1[18] ), .A2(
        \MC_ARK_ARC_1_0/temp2[18] ), .Z(\MC_ARK_ARC_1_0/temp5[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_28_5  ( .A1(\RI5[0][54] ), .A2(n477), .Z(
        \MC_ARK_ARC_1_0/temp4[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_28_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[180] ), 
        .A2(\MC_ARK_ARC_1_0/buf_datainput[156] ), .Z(
        \MC_ARK_ARC_1_0/temp2[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_28_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[12] ), 
        .A2(\RI5[0][18] ), .Z(\MC_ARK_ARC_1_0/temp1[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_28_4  ( .A1(\MC_ARK_ARC_1_0/temp5[19] ), .A2(
        \MC_ARK_ARC_1_0/temp6[19] ), .Z(\MC_ARK_ARC_1_0/buf_output[19] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_28_4  ( .A1(\RI5[0][55] ), .A2(n472), .Z(
        \MC_ARK_ARC_1_0/temp4[19] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_28_4  ( .A1(\RI5[0][85] ), .A2(\RI5[0][121] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[19] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_28_4  ( .A1(\RI5[0][181] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[157] ), .Z(\MC_ARK_ARC_1_0/temp2[19] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_28_3  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[56] ), 
        .A2(n467), .Z(\MC_ARK_ARC_1_0/temp4[20] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_28_3  ( .A1(\RI5[0][122] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[86] ), .Z(\MC_ARK_ARC_1_0/temp3[20] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_28_3  ( .A1(\RI5[0][20] ), .A2(\RI5[0][14] ), .Z(
        \MC_ARK_ARC_1_0/temp1[20] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_28_2  ( .A1(\RI5[0][57] ), .A2(n103), .Z(
        \MC_ARK_ARC_1_0/temp4[21] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_28_1  ( .A1(\RI5[0][58] ), .A2(n215), .Z(
        \MC_ARK_ARC_1_0/temp4[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_28_1  ( .A1(\RI5[0][124] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[88] ), .Z(\MC_ARK_ARC_1_0/temp3[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_28_1  ( .A1(\RI5[0][160] ), .A2(\RI5[0][184] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_28_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[22] ), 
        .A2(\RI5[0][16] ), .Z(\MC_ARK_ARC_1_0/temp1[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_28_0  ( .A1(\RI5[0][59] ), .A2(n452), .Z(
        \MC_ARK_ARC_1_0/temp4[23] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_28_0  ( .A1(\RI5[0][185] ), .A2(\RI5[0][161] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[23] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_27_5  ( .A1(\RI5[0][60] ), .A2(n18), .Z(
        \MC_ARK_ARC_1_0/temp4[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_27_5  ( .A1(\RI5[0][126] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[90] ), .Z(\MC_ARK_ARC_1_0/temp3[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_27_5  ( .A1(\RI5[0][162] ), .A2(\RI5[0][186] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_27_4  ( .A1(\MC_ARK_ARC_1_0/temp3[25] ), .A2(
        \MC_ARK_ARC_1_0/temp4[25] ), .Z(\MC_ARK_ARC_1_0/temp6[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_27_4  ( .A1(\MC_ARK_ARC_1_0/temp2[25] ), .A2(
        \MC_ARK_ARC_1_0/temp1[25] ), .Z(\MC_ARK_ARC_1_0/temp5[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_27_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[61] ), 
        .A2(n67), .Z(\MC_ARK_ARC_1_0/temp4[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_27_4  ( .A1(\RI5[0][127] ), .A2(\RI5[0][91] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_27_4  ( .A1(\SB2_0_0/buf_output[1] ), .A2(
        \RI5[0][25] ), .Z(\MC_ARK_ARC_1_0/temp1[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_27_3  ( .A1(\RI5[0][62] ), .A2(n24), .Z(
        \MC_ARK_ARC_1_0/temp4[26] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_27_3  ( .A1(\RI5[0][20] ), .A2(\RI5[0][26] ), .Z(
        \MC_ARK_ARC_1_0/temp1[26] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_27_2  ( .A1(\RI5[0][63] ), .A2(n564), .Z(
        \MC_ARK_ARC_1_0/temp4[27] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_27_1  ( .A1(\RI5[0][64] ), .A2(n196), .Z(
        \MC_ARK_ARC_1_0/temp4[28] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_27_1  ( .A1(\RI5[0][94] ), .A2(\RI5[0][130] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[28] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_27_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[22] ), 
        .A2(\RI5[0][28] ), .Z(\MC_ARK_ARC_1_0/temp1[28] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_27_0  ( .A1(\MC_ARK_ARC_1_0/temp5[29] ), .A2(
        \MC_ARK_ARC_1_0/temp6[29] ), .Z(\MC_ARK_ARC_1_0/buf_output[29] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_27_0  ( .A1(\MC_ARK_ARC_1_0/temp4[29] ), .A2(
        \MC_ARK_ARC_1_0/temp3[29] ), .Z(\MC_ARK_ARC_1_0/temp6[29] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_27_0  ( .A1(\RI5[0][65] ), .A2(n167), .Z(
        \MC_ARK_ARC_1_0/temp4[29] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_27_0  ( .A1(\RI5[0][95] ), .A2(\RI5[0][131] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[29] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_27_0  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[167] ), 
        .A2(\RI5[0][191] ), .Z(\MC_ARK_ARC_1_0/temp2[29] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_26_5  ( .A1(\MC_ARK_ARC_1_0/temp3[30] ), .A2(
        \MC_ARK_ARC_1_0/temp4[30] ), .Z(\MC_ARK_ARC_1_0/temp6[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_26_5  ( .A1(\RI5[0][66] ), .A2(n239), .Z(
        \MC_ARK_ARC_1_0/temp4[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_26_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[132] ), 
        .A2(\MC_ARK_ARC_1_0/buf_datainput[96] ), .Z(\MC_ARK_ARC_1_0/temp3[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_26_5  ( .A1(\RI5[0][168] ), .A2(\RI5[0][0] ), .Z(
        \MC_ARK_ARC_1_0/temp2[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_26_5  ( .A1(\RI5[0][30] ), .A2(\RI5[0][24] ), .Z(
        \MC_ARK_ARC_1_0/temp1[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_26_4  ( .A1(\MC_ARK_ARC_1_0/temp6[31] ), .A2(
        \MC_ARK_ARC_1_0/temp5[31] ), .Z(\MC_ARK_ARC_1_0/buf_output[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_26_4  ( .A1(\MC_ARK_ARC_1_0/temp3[31] ), .A2(
        \MC_ARK_ARC_1_0/temp4[31] ), .Z(\MC_ARK_ARC_1_0/temp6[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_26_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[67] ), 
        .A2(n152), .Z(\MC_ARK_ARC_1_0/temp4[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_26_4  ( .A1(\RI5[0][133] ), .A2(\RI5[0][97] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_26_4  ( .A1(\RI5[0][31] ), .A2(\RI5[0][25] ), .Z(
        \MC_ARK_ARC_1_0/temp1[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_26_3  ( .A1(\RI5[0][68] ), .A2(n40), .Z(
        \MC_ARK_ARC_1_0/temp4[32] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_26_3  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[2] ), 
        .A2(\RI5[0][170] ), .Z(\MC_ARK_ARC_1_0/temp2[32] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_26_3  ( .A1(\RI5[0][32] ), .A2(\RI5[0][26] ), .Z(
        \MC_ARK_ARC_1_0/temp1[32] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_26_2  ( .A1(\MC_ARK_ARC_1_0/temp5[33] ), .A2(
        \MC_ARK_ARC_1_0/temp6[33] ), .Z(\MC_ARK_ARC_1_0/buf_output[33] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_26_2  ( .A1(\MC_ARK_ARC_1_0/temp3[33] ), .A2(
        \MC_ARK_ARC_1_0/temp4[33] ), .Z(\MC_ARK_ARC_1_0/temp6[33] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_26_2  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[69] ), 
        .A2(n539), .Z(\MC_ARK_ARC_1_0/temp4[33] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_26_2  ( .A1(\RI5[0][135] ), .A2(\RI5[0][99] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[33] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_26_1  ( .A1(\RI5[0][70] ), .A2(n199), .Z(
        \MC_ARK_ARC_1_0/temp4[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_26_1  ( .A1(\RI5[0][4] ), .A2(\RI5[0][172] ), .Z(
        \MC_ARK_ARC_1_0/temp2[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_26_1  ( .A1(\RI5[0][34] ), .A2(\RI5[0][28] ), .Z(
        \MC_ARK_ARC_1_0/temp1[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_26_0  ( .A1(\RI5[0][71] ), .A2(n217), .Z(
        \MC_ARK_ARC_1_0/temp4[35] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_25_5  ( .A1(\MC_ARK_ARC_1_0/temp5[36] ), .A2(
        \MC_ARK_ARC_1_0/temp6[36] ), .Z(\MC_ARK_ARC_1_0/buf_output[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_25_5  ( .A1(\MC_ARK_ARC_1_0/temp3[36] ), .A2(
        \MC_ARK_ARC_1_0/temp4[36] ), .Z(\MC_ARK_ARC_1_0/temp6[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_25_5  ( .A1(\RI5[0][72] ), .A2(n156), .Z(
        \MC_ARK_ARC_1_0/temp4[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_25_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[138] ), 
        .A2(\RI5[0][102] ), .Z(\MC_ARK_ARC_1_0/temp3[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_25_5  ( .A1(\RI5[0][174] ), .A2(\RI5[0][6] ), .Z(
        \MC_ARK_ARC_1_0/temp2[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_25_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[36] ), 
        .A2(\RI5[0][30] ), .Z(\MC_ARK_ARC_1_0/temp1[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_25_4  ( .A1(\MC_ARK_ARC_1_0/temp1[37] ), .A2(
        \MC_ARK_ARC_1_0/temp2[37] ), .Z(\MC_ARK_ARC_1_0/temp5[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_25_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[73] ), 
        .A2(n518), .Z(\MC_ARK_ARC_1_0/temp4[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_25_4  ( .A1(\RI5[0][103] ), .A2(\RI5[0][139] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_25_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[7] ), 
        .A2(\RI5[0][175] ), .Z(\MC_ARK_ARC_1_0/temp2[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_25_4  ( .A1(\RI5[0][37] ), .A2(\RI5[0][31] ), .Z(
        \MC_ARK_ARC_1_0/temp1[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_25_3  ( .A1(\MC_ARK_ARC_1_0/temp5[38] ), .A2(
        \MC_ARK_ARC_1_0/temp6[38] ), .Z(\MC_ARK_ARC_1_0/buf_output[38] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_25_3  ( .A1(\RI5[0][8] ), .A2(\RI5[0][176] ), .Z(
        \MC_ARK_ARC_1_0/temp2[38] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_25_3  ( .A1(\RI5[0][38] ), .A2(\RI5[0][32] ), .Z(
        \MC_ARK_ARC_1_0/temp1[38] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_25_2  ( .A1(\RI5[0][75] ), .A2(n126), .Z(
        \MC_ARK_ARC_1_0/temp4[39] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_25_2  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[105] ), 
        .A2(\MC_ARK_ARC_1_0/buf_datainput[141] ), .Z(
        \MC_ARK_ARC_1_0/temp3[39] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_25_1  ( .A1(\MC_ARK_ARC_1_0/temp4[40] ), .A2(
        \MC_ARK_ARC_1_0/temp3[40] ), .Z(\MC_ARK_ARC_1_0/temp6[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_25_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[76] ), 
        .A2(n56), .Z(\MC_ARK_ARC_1_0/temp4[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_25_1  ( .A1(\RI5[0][142] ), .A2(\RI5[0][106] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_25_1  ( .A1(\RI5[0][10] ), .A2(\RI5[0][178] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_25_0  ( .A1(\MC_ARK_ARC_1_0/temp3[41] ), .A2(
        \MC_ARK_ARC_1_0/temp4[41] ), .Z(\MC_ARK_ARC_1_0/temp6[41] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_25_0  ( .A1(\RI5[0][77] ), .A2(n189), .Z(
        \MC_ARK_ARC_1_0/temp4[41] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_25_0  ( .A1(\RI5[0][107] ), .A2(\RI5[0][143] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[41] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_25_0  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[179] ), 
        .A2(\RI5[0][11] ), .Z(\MC_ARK_ARC_1_0/temp2[41] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_24_5  ( .A1(\MC_ARK_ARC_1_0/temp5[42] ), .A2(
        \MC_ARK_ARC_1_0/temp6[42] ), .Z(\MC_ARK_ARC_1_0/buf_output[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_24_5  ( .A1(\MC_ARK_ARC_1_0/temp3[42] ), .A2(
        \MC_ARK_ARC_1_0/temp4[42] ), .Z(\MC_ARK_ARC_1_0/temp6[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_24_5  ( .A1(\MC_ARK_ARC_1_0/temp1[42] ), .A2(
        \MC_ARK_ARC_1_0/temp2[42] ), .Z(\MC_ARK_ARC_1_0/temp5[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_24_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[78] ), 
        .A2(n58), .Z(\MC_ARK_ARC_1_0/temp4[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_24_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[144] ), 
        .A2(\RI5[0][108] ), .Z(\MC_ARK_ARC_1_0/temp3[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_24_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[180] ), 
        .A2(\MC_ARK_ARC_1_0/buf_datainput[12] ), .Z(\MC_ARK_ARC_1_0/temp2[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_24_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[42] ), 
        .A2(\MC_ARK_ARC_1_0/buf_datainput[36] ), .Z(\MC_ARK_ARC_1_0/temp1[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_24_4  ( .A1(\MC_ARK_ARC_1_0/temp3[43] ), .A2(
        \MC_ARK_ARC_1_0/temp4[43] ), .Z(\MC_ARK_ARC_1_0/temp6[43] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_24_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[79] ), 
        .A2(n491), .Z(\MC_ARK_ARC_1_0/temp4[43] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_24_4  ( .A1(\RI5[0][145] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[109] ), .Z(\MC_ARK_ARC_1_0/temp3[43] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_24_4  ( .A1(\RI5[0][13] ), .A2(\RI5[0][181] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[43] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_24_3  ( .A1(\RI5[0][80] ), .A2(n485), .Z(
        \MC_ARK_ARC_1_0/temp4[44] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_24_3  ( .A1(\RI5[0][110] ), .A2(\RI5[0][146] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[44] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_24_3  ( .A1(\RI5[0][182] ), .A2(n5497), .Z(
        \MC_ARK_ARC_1_0/temp2[44] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_24_2  ( .A1(\MC_ARK_ARC_1_0/temp6[45] ), .A2(
        \MC_ARK_ARC_1_0/temp5[45] ), .Z(\MC_ARK_ARC_1_0/buf_output[45] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_24_2  ( .A1(\MC_ARK_ARC_1_0/temp3[45] ), .A2(
        \MC_ARK_ARC_1_0/temp4[45] ), .Z(\MC_ARK_ARC_1_0/temp6[45] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_24_2  ( .A1(\MC_ARK_ARC_1_0/temp2[45] ), .A2(
        \MC_ARK_ARC_1_0/temp1[45] ), .Z(\MC_ARK_ARC_1_0/temp5[45] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_24_2  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[81] ), 
        .A2(n479), .Z(\MC_ARK_ARC_1_0/temp4[45] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_24_2  ( .A1(\RI5[0][39] ), .A2(\RI5[0][45] ), .Z(
        \MC_ARK_ARC_1_0/temp1[45] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_24_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[82] ), 
        .A2(n197), .Z(\MC_ARK_ARC_1_0/temp4[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_24_1  ( .A1(\RI5[0][148] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[112] ), .Z(\MC_ARK_ARC_1_0/temp3[46] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_24_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[46] ), 
        .A2(\RI5[0][40] ), .Z(\MC_ARK_ARC_1_0/temp1[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_24_0  ( .A1(\MC_ARK_ARC_1_0/temp1[47] ), .A2(
        \MC_ARK_ARC_1_0/temp2[47] ), .Z(\MC_ARK_ARC_1_0/temp5[47] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_24_0  ( .A1(\RI5[0][83] ), .A2(n233), .Z(
        \MC_ARK_ARC_1_0/temp4[47] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_24_0  ( .A1(\RI5[0][113] ), .A2(\RI5[0][149] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[47] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_24_0  ( .A1(\RI5[0][17] ), .A2(\RI5[0][185] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[47] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_23_5  ( .A1(\MC_ARK_ARC_1_0/temp5[48] ), .A2(
        \MC_ARK_ARC_1_0/temp6[48] ), .Z(\MC_ARK_ARC_1_0/buf_output[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_23_5  ( .A1(\MC_ARK_ARC_1_0/temp3[48] ), .A2(
        \MC_ARK_ARC_1_0/temp4[48] ), .Z(\MC_ARK_ARC_1_0/temp6[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_23_5  ( .A1(\RI5[0][84] ), .A2(n465), .Z(
        \MC_ARK_ARC_1_0/temp4[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_23_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[48] ), 
        .A2(\MC_ARK_ARC_1_0/buf_datainput[42] ), .Z(\MC_ARK_ARC_1_0/temp1[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_23_4  ( .A1(\MC_ARK_ARC_1_0/temp2[49] ), .A2(
        \MC_ARK_ARC_1_0/temp1[49] ), .Z(\MC_ARK_ARC_1_0/temp5[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_23_4  ( .A1(\RI5[0][85] ), .A2(n133), .Z(
        \MC_ARK_ARC_1_0/temp4[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_23_4  ( .A1(\RI5[0][151] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[115] ), .Z(\MC_ARK_ARC_1_0/temp3[49] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_23_4  ( .A1(\RI5[0][19] ), .A2(\RI5[0][187] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_23_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[49] ), 
        .A2(\RI5[0][43] ), .Z(\MC_ARK_ARC_1_0/temp1[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_23_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[88] ), 
        .A2(n108), .Z(\MC_ARK_ARC_1_0/temp4[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_23_1  ( .A1(\RI5[0][154] ), .A2(\RI5[0][118] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_23_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[46] ), 
        .A2(\RI5[0][52] ), .Z(\MC_ARK_ARC_1_0/temp1[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_23_0  ( .A1(\RI5[0][89] ), .A2(n137), .Z(
        \MC_ARK_ARC_1_0/temp4[53] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_22_5  ( .A1(\MC_ARK_ARC_1_0/temp5[54] ), .A2(
        \MC_ARK_ARC_1_0/temp6[54] ), .Z(\MC_ARK_ARC_1_0/buf_output[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_22_5  ( .A1(\MC_ARK_ARC_1_0/temp4[54] ), .A2(
        \MC_ARK_ARC_1_0/temp3[54] ), .Z(\MC_ARK_ARC_1_0/temp6[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_22_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[90] ), 
        .A2(n241), .Z(\MC_ARK_ARC_1_0/temp4[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_22_5  ( .A1(\RI5[0][120] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[156] ), .Z(\MC_ARK_ARC_1_0/temp3[54] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_22_5  ( .A1(\RI5[0][54] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[48] ), .Z(\MC_ARK_ARC_1_0/temp1[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_22_4  ( .A1(\RI5[0][91] ), .A2(n57), .Z(
        \MC_ARK_ARC_1_0/temp4[55] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_22_4  ( .A1(\RI5[0][1] ), .A2(\RI5[0][25] ), .Z(
        \MC_ARK_ARC_1_0/temp2[55] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_22_3  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[92] ), 
        .A2(n50), .Z(\MC_ARK_ARC_1_0/temp4[56] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_22_2  ( .A1(\RI5[0][93] ), .A2(n136), .Z(
        \MC_ARK_ARC_1_0/temp4[57] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_22_2  ( .A1(\RI5[0][159] ), .A2(\RI5[0][123] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[57] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_22_1  ( .A1(\MC_ARK_ARC_1_0/temp1[58] ), .A2(
        \MC_ARK_ARC_1_0/temp2[58] ), .Z(\MC_ARK_ARC_1_0/temp5[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_22_1  ( .A1(\RI5[0][94] ), .A2(n548), .Z(
        \MC_ARK_ARC_1_0/temp4[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_22_1  ( .A1(\RI5[0][160] ), .A2(\RI5[0][124] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_22_1  ( .A1(\RI5[0][28] ), .A2(\RI5[0][4] ), .Z(
        \MC_ARK_ARC_1_0/temp2[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_22_0  ( .A1(\RI5[0][95] ), .A2(n185), .Z(
        \MC_ARK_ARC_1_0/temp4[59] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_22_0  ( .A1(\RI5[0][161] ), .A2(\RI5[0][125] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[59] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_22_0  ( .A1(\RI5[0][5] ), .A2(\RI5[0][29] ), .Z(
        \MC_ARK_ARC_1_0/temp2[59] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_21_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[96] ), 
        .A2(n107), .Z(\MC_ARK_ARC_1_0/temp4[60] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_21_5  ( .A1(\RI5[0][54] ), .A2(\RI5[0][60] ), .Z(
        \MC_ARK_ARC_1_0/temp1[60] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_21_4  ( .A1(\MC_ARK_ARC_1_0/temp3[61] ), .A2(
        \MC_ARK_ARC_1_0/temp4[61] ), .Z(\MC_ARK_ARC_1_0/temp6[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_21_4  ( .A1(\MC_ARK_ARC_1_0/temp2[61] ), .A2(
        \MC_ARK_ARC_1_0/temp1[61] ), .Z(\MC_ARK_ARC_1_0/temp5[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_21_4  ( .A1(\RI5[0][97] ), .A2(n536), .Z(
        \MC_ARK_ARC_1_0/temp4[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_21_4  ( .A1(\RI5[0][127] ), .A2(\RI5[0][163] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_21_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[7] ), 
        .A2(\RI5[0][31] ), .Z(\MC_ARK_ARC_1_0/temp2[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_21_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[61] ), 
        .A2(\RI5[0][55] ), .Z(\MC_ARK_ARC_1_0/temp1[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_21_3  ( .A1(\MC_ARK_ARC_1_0/temp5[62] ), .A2(
        \MC_ARK_ARC_1_0/temp6[62] ), .Z(\MC_ARK_ARC_1_0/buf_output[62] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_21_3  ( .A1(\MC_ARK_ARC_1_0/temp1[62] ), .A2(
        \MC_ARK_ARC_1_0/temp2[62] ), .Z(\MC_ARK_ARC_1_0/temp5[62] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_21_3  ( .A1(\RI5[0][8] ), .A2(\RI5[0][32] ), .Z(
        \MC_ARK_ARC_1_0/temp2[62] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_21_3  ( .A1(\RI5[0][62] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[56] ), .Z(\MC_ARK_ARC_1_0/temp1[62] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_21_2  ( .A1(\MC_ARK_ARC_1_0/temp3[63] ), .A2(
        \MC_ARK_ARC_1_0/temp4[63] ), .Z(\MC_ARK_ARC_1_0/temp6[63] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_21_2  ( .A1(\RI5[0][99] ), .A2(n124), .Z(
        \MC_ARK_ARC_1_0/temp4[63] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_21_1  ( .A1(\MC_ARK_ARC_1_0/temp5[64] ), .A2(
        \MC_ARK_ARC_1_0/temp6[64] ), .Z(\MC_ARK_ARC_1_0/buf_output[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_21_1  ( .A1(\MC_ARK_ARC_1_0/temp1[64] ), .A2(
        \MC_ARK_ARC_1_0/temp2[64] ), .Z(\MC_ARK_ARC_1_0/temp5[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_21_1  ( .A1(\RI5[0][100] ), .A2(n183), .Z(
        \MC_ARK_ARC_1_0/temp4[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_21_1  ( .A1(\RI5[0][34] ), .A2(\RI5[0][10] ), .Z(
        \MC_ARK_ARC_1_0/temp2[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_21_1  ( .A1(\RI5[0][64] ), .A2(\RI5[0][58] ), .Z(
        \MC_ARK_ARC_1_0/temp1[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_20_5  ( .A1(\RI5[0][102] ), .A2(n511), .Z(
        \MC_ARK_ARC_1_0/temp4[66] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_20_4  ( .A1(\MC_ARK_ARC_1_0/temp5[67] ), .A2(
        \MC_ARK_ARC_1_0/temp6[67] ), .Z(\MC_ARK_ARC_1_0/buf_output[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_20_4  ( .A1(\MC_ARK_ARC_1_0/temp3[67] ), .A2(
        \MC_ARK_ARC_1_0/temp4[67] ), .Z(\MC_ARK_ARC_1_0/temp6[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_20_4  ( .A1(\RI5[0][103] ), .A2(n30), .Z(
        \MC_ARK_ARC_1_0/temp4[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_20_4  ( .A1(\RI5[0][169] ), .A2(\RI5[0][133] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_20_4  ( .A1(\RI5[0][13] ), .A2(\RI5[0][37] ), .Z(
        \MC_ARK_ARC_1_0/temp2[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_20_3  ( .A1(\RI5[0][104] ), .A2(n187), .Z(
        \MC_ARK_ARC_1_0/temp4[68] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_20_3  ( .A1(\RI5[0][14] ), .A2(\RI5[0][38] ), .Z(
        \MC_ARK_ARC_1_0/temp2[68] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_20_2  ( .A1(\RI5[0][171] ), .A2(\RI5[0][135] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[69] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_20_1  ( .A1(\MC_ARK_ARC_1_0/temp2[70] ), .A2(
        \MC_ARK_ARC_1_0/temp1[70] ), .Z(\MC_ARK_ARC_1_0/temp5[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_20_1  ( .A1(\RI5[0][106] ), .A2(n77), .Z(
        \MC_ARK_ARC_1_0/temp4[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_20_1  ( .A1(\RI5[0][172] ), .A2(\RI5[0][136] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_20_1  ( .A1(\RI5[0][16] ), .A2(\RI5[0][40] ), .Z(
        \MC_ARK_ARC_1_0/temp2[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_20_1  ( .A1(\RI5[0][70] ), .A2(\RI5[0][64] ), .Z(
        \MC_ARK_ARC_1_0/temp1[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_19_5  ( .A1(\MC_ARK_ARC_1_0/temp5[72] ), .A2(
        \MC_ARK_ARC_1_0/temp6[72] ), .Z(\MC_ARK_ARC_1_0/buf_output[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_19_5  ( .A1(\MC_ARK_ARC_1_0/temp3[72] ), .A2(
        \MC_ARK_ARC_1_0/temp4[72] ), .Z(\MC_ARK_ARC_1_0/temp6[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_19_5  ( .A1(\RI5[0][108] ), .A2(n481), .Z(
        \MC_ARK_ARC_1_0/temp4[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_19_5  ( .A1(\RI5[0][72] ), .A2(\RI5[0][66] ), .Z(
        \MC_ARK_ARC_1_0/temp1[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_19_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[109] ), 
        .A2(n476), .Z(\MC_ARK_ARC_1_0/temp4[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_19_4  ( .A1(\RI5[0][175] ), .A2(\RI5[0][139] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_19_3  ( .A1(\RI5[0][110] ), .A2(n26), .Z(
        \MC_ARK_ARC_1_0/temp4[74] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_19_2  ( .A1(\RI5[0][111] ), .A2(n100), .Z(
        \MC_ARK_ARC_1_0/temp4[75] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_19_1  ( .A1(\MC_ARK_ARC_1_0/temp2[76] ), .A2(
        \MC_ARK_ARC_1_0/temp1[76] ), .Z(\MC_ARK_ARC_1_0/temp5[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_19_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[112] ), 
        .A2(n462), .Z(\MC_ARK_ARC_1_0/temp4[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_19_0  ( .A1(\MC_ARK_ARC_1_0/temp4[77] ), .A2(
        \MC_ARK_ARC_1_0/temp3[77] ), .Z(\MC_ARK_ARC_1_0/temp6[77] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_19_0  ( .A1(\RI5[0][113] ), .A2(n458), .Z(
        \MC_ARK_ARC_1_0/temp4[77] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_19_0  ( .A1(\RI5[0][23] ), .A2(\RI5[0][47] ), .Z(
        \MC_ARK_ARC_1_0/temp2[77] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_19_0  ( .A1(\RI5[0][77] ), .A2(\RI5[0][71] ), .Z(
        \MC_ARK_ARC_1_0/temp1[77] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_18_5  ( .A1(\MC_ARK_ARC_1_0/temp5[78] ), .A2(
        \MC_ARK_ARC_1_0/temp6[78] ), .Z(\MC_ARK_ARC_1_0/buf_output[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_18_5  ( .A1(\MC_ARK_ARC_1_0/temp3[78] ), .A2(
        \MC_ARK_ARC_1_0/temp4[78] ), .Z(\MC_ARK_ARC_1_0/temp6[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_18_5  ( .A1(\MC_ARK_ARC_1_0/temp1[78] ), .A2(
        \MC_ARK_ARC_1_0/temp2[78] ), .Z(\MC_ARK_ARC_1_0/temp5[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_18_5  ( .A1(n1375), .A2(n451), .Z(
        \MC_ARK_ARC_1_0/temp4[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_18_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[180] ), 
        .A2(\MC_ARK_ARC_1_0/buf_datainput[144] ), .Z(
        \MC_ARK_ARC_1_0/temp3[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_18_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[48] ), 
        .A2(\RI5[0][24] ), .Z(\MC_ARK_ARC_1_0/temp2[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_18_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[78] ), 
        .A2(\RI5[0][72] ), .Z(\MC_ARK_ARC_1_0/temp1[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_18_4  ( .A1(\MC_ARK_ARC_1_0/temp2[79] ), .A2(
        \MC_ARK_ARC_1_0/temp1[79] ), .Z(\MC_ARK_ARC_1_0/temp5[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_18_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[115] ), 
        .A2(n47), .Z(\MC_ARK_ARC_1_0/temp4[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_18_4  ( .A1(\RI5[0][181] ), .A2(\RI5[0][145] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_18_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[49] ), 
        .A2(\RI5[0][25] ), .Z(\MC_ARK_ARC_1_0/temp2[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_18_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[79] ), 
        .A2(\MC_ARK_ARC_1_0/buf_datainput[73] ), .Z(\MC_ARK_ARC_1_0/temp1[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_18_3  ( .A1(\RI5[0][116] ), .A2(n60), .Z(
        \MC_ARK_ARC_1_0/temp4[80] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_18_3  ( .A1(\RI5[0][50] ), .A2(\RI5[0][26] ), .Z(
        \MC_ARK_ARC_1_0/temp2[80] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_18_2  ( .A1(\MC_ARK_ARC_1_0/temp4[81] ), .A2(
        \MC_ARK_ARC_1_0/temp3[81] ), .Z(\MC_ARK_ARC_1_0/temp6[81] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_18_2  ( .A1(\RI5[0][117] ), .A2(n223), .Z(
        \MC_ARK_ARC_1_0/temp4[81] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_18_2  ( .A1(\RI5[0][147] ), .A2(\RI5[0][183] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[81] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_18_1  ( .A1(\MC_ARK_ARC_1_0/temp3[82] ), .A2(
        \MC_ARK_ARC_1_0/temp4[82] ), .Z(\MC_ARK_ARC_1_0/temp6[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_18_1  ( .A1(\RI5[0][118] ), .A2(n219), .Z(
        \MC_ARK_ARC_1_0/temp4[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_18_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[82] ), 
        .A2(\MC_ARK_ARC_1_0/buf_datainput[76] ), .Z(\MC_ARK_ARC_1_0/temp1[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_18_0  ( .A1(\MC_ARK_ARC_1_0/temp5[83] ), .A2(
        \MC_ARK_ARC_1_0/temp6[83] ), .Z(\MC_ARK_ARC_1_0/buf_output[83] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_18_0  ( .A1(\MC_ARK_ARC_1_0/temp3[83] ), .A2(
        \MC_ARK_ARC_1_0/temp4[83] ), .Z(\MC_ARK_ARC_1_0/temp6[83] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_18_0  ( .A1(\RI5[0][119] ), .A2(n170), .Z(
        \MC_ARK_ARC_1_0/temp4[83] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_18_0  ( .A1(\RI5[0][185] ), .A2(\RI5[0][149] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[83] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_18_0  ( .A1(\RI5[0][83] ), .A2(\RI5[0][77] ), .Z(
        \MC_ARK_ARC_1_0/temp1[83] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_17_5  ( .A1(\MC_ARK_ARC_1_0/temp2[84] ), .A2(
        \MC_ARK_ARC_1_0/temp1[84] ), .Z(\MC_ARK_ARC_1_0/temp5[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_17_5  ( .A1(\RI5[0][120] ), .A2(n556), .Z(
        \MC_ARK_ARC_1_0/temp4[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_17_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[150] ), 
        .A2(\RI5[0][186] ), .Z(\MC_ARK_ARC_1_0/temp3[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_17_5  ( .A1(\RI5[0][54] ), .A2(\RI5[0][30] ), .Z(
        \MC_ARK_ARC_1_0/temp2[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_17_5  ( .A1(\RI5[0][84] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[78] ), .Z(\MC_ARK_ARC_1_0/temp1[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_17_4  ( .A1(\RI5[0][121] ), .A2(n551), .Z(
        \MC_ARK_ARC_1_0/temp4[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_17_4  ( .A1(\RI5[0][187] ), .A2(\RI5[0][151] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_17_4  ( .A1(\RI5[0][55] ), .A2(\RI5[0][31] ), .Z(
        \MC_ARK_ARC_1_0/temp2[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_17_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[79] ), 
        .A2(\RI5[0][85] ), .Z(\MC_ARK_ARC_1_0/temp1[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_17_3  ( .A1(\SB2_0_14/buf_output[2] ), .A2(n545), 
        .Z(\MC_ARK_ARC_1_0/temp4[86] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_17_2  ( .A1(\MC_ARK_ARC_1_0/temp6[87] ), .A2(
        \MC_ARK_ARC_1_0/temp5[87] ), .Z(\MC_ARK_ARC_1_0/buf_output[87] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_17_2  ( .A1(\MC_ARK_ARC_1_0/temp3[87] ), .A2(
        \MC_ARK_ARC_1_0/temp4[87] ), .Z(\MC_ARK_ARC_1_0/temp6[87] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_17_2  ( .A1(\RI5[0][123] ), .A2(n166), .Z(
        \MC_ARK_ARC_1_0/temp4[87] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_17_2  ( .A1(\RI5[0][189] ), .A2(\RI5[0][153] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[87] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_17_1  ( .A1(\RI5[0][124] ), .A2(n538), .Z(
        \MC_ARK_ARC_1_0/temp4[88] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_17_1  ( .A1(\RI5[0][190] ), .A2(\RI5[0][154] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[88] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_17_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[88] ), 
        .A2(\MC_ARK_ARC_1_0/buf_datainput[82] ), .Z(\MC_ARK_ARC_1_0/temp1[88] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_17_0  ( .A1(\RI5[0][125] ), .A2(n532), .Z(
        \MC_ARK_ARC_1_0/temp4[89] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_17_0  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[155] ), 
        .A2(\RI5[0][191] ), .Z(\MC_ARK_ARC_1_0/temp3[89] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_17_0  ( .A1(\RI5[0][59] ), .A2(\RI5[0][35] ), .Z(
        \MC_ARK_ARC_1_0/temp2[89] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_17_0  ( .A1(\RI5[0][89] ), .A2(\RI5[0][83] ), .Z(
        \MC_ARK_ARC_1_0/temp1[89] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_16_5  ( .A1(\MC_ARK_ARC_1_0/temp6[90] ), .A2(
        \MC_ARK_ARC_1_0/temp5[90] ), .Z(\MC_ARK_ARC_1_0/buf_output[90] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_16_5  ( .A1(\MC_ARK_ARC_1_0/temp3[90] ), .A2(
        \MC_ARK_ARC_1_0/temp4[90] ), .Z(\MC_ARK_ARC_1_0/temp6[90] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_16_5  ( .A1(\MC_ARK_ARC_1_0/temp1[90] ), .A2(
        \MC_ARK_ARC_1_0/temp2[90] ), .Z(\MC_ARK_ARC_1_0/temp5[90] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_16_5  ( .A1(\RI5[0][126] ), .A2(n200), .Z(
        \MC_ARK_ARC_1_0/temp4[90] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_16_5  ( .A1(\RI5[0][0] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[156] ), .Z(\MC_ARK_ARC_1_0/temp3[90] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_16_5  ( .A1(\RI5[0][60] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[36] ), .Z(\MC_ARK_ARC_1_0/temp2[90] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_16_5  ( .A1(\RI5[0][84] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[90] ), .Z(\MC_ARK_ARC_1_0/temp1[90] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_16_4  ( .A1(\MC_ARK_ARC_1_0/temp6[91] ), .A2(
        \MC_ARK_ARC_1_0/temp5[91] ), .Z(\MC_ARK_ARC_1_0/buf_output[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_16_4  ( .A1(\MC_ARK_ARC_1_0/temp4[91] ), .A2(
        \MC_ARK_ARC_1_0/temp3[91] ), .Z(\MC_ARK_ARC_1_0/temp6[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_16_4  ( .A1(\RI5[0][127] ), .A2(n224), .Z(
        \MC_ARK_ARC_1_0/temp4[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_16_4  ( .A1(\RI5[0][1] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[157] ), .Z(\MC_ARK_ARC_1_0/temp3[91] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_16_4  ( .A1(\RI5[0][37] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[61] ), .Z(\MC_ARK_ARC_1_0/temp2[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_16_3  ( .A1(\RI5[0][62] ), .A2(\RI5[0][38] ), .Z(
        \MC_ARK_ARC_1_0/temp2[92] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_16_2  ( .A1(\RI5[0][129] ), .A2(n193), .Z(
        \MC_ARK_ARC_1_0/temp4[93] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_16_1  ( .A1(\MC_ARK_ARC_1_0/temp6[94] ), .A2(
        \MC_ARK_ARC_1_0/temp5[94] ), .Z(\MC_ARK_ARC_1_0/buf_output[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_16_1  ( .A1(\RI5[0][130] ), .A2(n186), .Z(
        \MC_ARK_ARC_1_0/temp4[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_16_1  ( .A1(\RI5[0][160] ), .A2(\RI5[0][4] ), .Z(
        \MC_ARK_ARC_1_0/temp3[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_16_1  ( .A1(\RI5[0][94] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[88] ), .Z(\MC_ARK_ARC_1_0/temp1[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_16_0  ( .A1(\RI5[0][131] ), .A2(n74), .Z(
        \MC_ARK_ARC_1_0/temp4[95] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_16_0  ( .A1(\RI5[0][161] ), .A2(\RI5[0][5] ), .Z(
        \MC_ARK_ARC_1_0/temp3[95] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_15_5  ( .A1(\MC_ARK_ARC_1_0/temp3[96] ), .A2(
        \MC_ARK_ARC_1_0/temp4[96] ), .Z(\MC_ARK_ARC_1_0/temp6[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_15_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[132] ), 
        .A2(n190), .Z(\MC_ARK_ARC_1_0/temp4[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_15_5  ( .A1(\RI5[0][6] ), .A2(\RI5[0][162] ), .Z(
        \MC_ARK_ARC_1_0/temp3[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_15_5  ( .A1(\RI5[0][66] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[42] ), .Z(\MC_ARK_ARC_1_0/temp2[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_15_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[96] ), 
        .A2(\MC_ARK_ARC_1_0/buf_datainput[90] ), .Z(\MC_ARK_ARC_1_0/temp1[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_15_4  ( .A1(\RI5[0][133] ), .A2(n495), .Z(
        \MC_ARK_ARC_1_0/temp4[97] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_15_4  ( .A1(\SB2_0_2/buf_output[1] ), .A2(
        \RI5[0][163] ), .Z(\MC_ARK_ARC_1_0/temp3[97] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_15_3  ( .A1(\SB2_0_12/buf_output[2] ), .A2(n490), 
        .Z(\MC_ARK_ARC_1_0/temp4[98] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_15_2  ( .A1(\MC_ARK_ARC_1_0/temp3[99] ), .A2(
        \MC_ARK_ARC_1_0/temp4[99] ), .Z(\MC_ARK_ARC_1_0/temp6[99] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_15_2  ( .A1(\RI5[0][135] ), .A2(n484), .Z(
        \MC_ARK_ARC_1_0/temp4[99] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_15_2  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[165] ), 
        .A2(\RI5[0][9] ), .Z(\MC_ARK_ARC_1_0/temp3[99] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_15_2  ( .A1(\RI5[0][93] ), .A2(\RI5[0][99] ), .Z(
        \MC_ARK_ARC_1_0/temp1[99] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_15_1  ( .A1(\RI5[0][136] ), .A2(n76), .Z(
        \MC_ARK_ARC_1_0/temp4[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_15_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[166] ), 
        .A2(\RI5[0][10] ), .Z(\MC_ARK_ARC_1_0/temp3[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_14_5  ( .A1(\MC_ARK_ARC_1_0/temp1[102] ), .A2(
        \MC_ARK_ARC_1_0/temp2[102] ), .Z(\MC_ARK_ARC_1_0/temp5[102] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_14_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[138] ), 
        .A2(n160), .Z(\MC_ARK_ARC_1_0/temp4[102] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_14_5  ( .A1(\RI5[0][168] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[12] ), .Z(\MC_ARK_ARC_1_0/temp3[102] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_14_5  ( .A1(\RI5[0][72] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[48] ), .Z(\MC_ARK_ARC_1_0/temp2[102] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_14_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[96] ), 
        .A2(\RI5[0][102] ), .Z(\MC_ARK_ARC_1_0/temp1[102] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_14_4  ( .A1(\MC_ARK_ARC_1_0/temp6[103] ), .A2(
        \MC_ARK_ARC_1_0/temp5[103] ), .Z(\MC_ARK_ARC_1_0/buf_output[103] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_14_4  ( .A1(\MC_ARK_ARC_1_0/temp3[103] ), .A2(
        \MC_ARK_ARC_1_0/temp4[103] ), .Z(\MC_ARK_ARC_1_0/temp6[103] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_14_4  ( .A1(\RI5[0][139] ), .A2(n131), .Z(
        \MC_ARK_ARC_1_0/temp4[103] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_14_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[73] ), 
        .A2(\MC_ARK_ARC_1_0/buf_datainput[49] ), .Z(
        \MC_ARK_ARC_1_0/temp2[103] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_14_3  ( .A1(\RI5[0][140] ), .A2(n121), .Z(
        \MC_ARK_ARC_1_0/temp4[104] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_14_3  ( .A1(\RI5[0][50] ), .A2(\RI5[0][74] ), .Z(
        \MC_ARK_ARC_1_0/temp2[104] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_14_2  ( .A1(\MC_ARK_ARC_1_0/temp6[105] ), .A2(
        \MC_ARK_ARC_1_0/temp5[105] ), .Z(\MC_ARK_ARC_1_0/buf_output[105] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_14_2  ( .A1(\MC_ARK_ARC_1_0/temp1[105] ), .A2(
        \MC_ARK_ARC_1_0/temp2[105] ), .Z(\MC_ARK_ARC_1_0/temp5[105] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_14_2  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[141] ), 
        .A2(n454), .Z(\MC_ARK_ARC_1_0/temp4[105] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_14_2  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[51] ), 
        .A2(\RI5[0][75] ), .Z(\MC_ARK_ARC_1_0/temp2[105] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_14_1  ( .A1(\MC_ARK_ARC_1_0/temp6[106] ), .A2(
        \MC_ARK_ARC_1_0/temp5[106] ), .Z(\MC_ARK_ARC_1_0/buf_output[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_14_1  ( .A1(\MC_ARK_ARC_1_0/temp3[106] ), .A2(
        \MC_ARK_ARC_1_0/temp4[106] ), .Z(\MC_ARK_ARC_1_0/temp6[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_14_1  ( .A1(\RI5[0][142] ), .A2(n128), .Z(
        \MC_ARK_ARC_1_0/temp4[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_14_1  ( .A1(\RI5[0][16] ), .A2(\RI5[0][172] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_14_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[76] ), 
        .A2(\RI5[0][52] ), .Z(\MC_ARK_ARC_1_0/temp2[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_14_1  ( .A1(\RI5[0][106] ), .A2(\RI5[0][100] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_14_0  ( .A1(\MC_ARK_ARC_1_0/temp1[107] ), .A2(
        \MC_ARK_ARC_1_0/temp2[107] ), .Z(\MC_ARK_ARC_1_0/temp5[107] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_14_0  ( .A1(\RI5[0][143] ), .A2(n444), .Z(
        \MC_ARK_ARC_1_0/temp4[107] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_14_0  ( .A1(\RI5[0][173] ), .A2(\RI5[0][17] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[107] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_14_0  ( .A1(\RI5[0][53] ), .A2(\RI5[0][77] ), .Z(
        \MC_ARK_ARC_1_0/temp2[107] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_14_0  ( .A1(\RI5[0][101] ), .A2(\RI5[0][107] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[107] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_13_5  ( .A1(\MC_ARK_ARC_1_0/temp6[108] ), .A2(
        \MC_ARK_ARC_1_0/temp5[108] ), .Z(\MC_ARK_ARC_1_0/buf_output[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_13_5  ( .A1(\MC_ARK_ARC_1_0/temp3[108] ), .A2(
        \MC_ARK_ARC_1_0/temp4[108] ), .Z(\MC_ARK_ARC_1_0/temp6[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_13_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[144] ), 
        .A2(n191), .Z(\MC_ARK_ARC_1_0/temp4[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_13_5  ( .A1(\RI5[0][54] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[78] ), .Z(\MC_ARK_ARC_1_0/temp2[108] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_13_4  ( .A1(\MC_ARK_ARC_1_0/temp1[109] ), .A2(
        \MC_ARK_ARC_1_0/temp2[109] ), .Z(\MC_ARK_ARC_1_0/temp5[109] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_13_4  ( .A1(\RI5[0][145] ), .A2(n55), .Z(
        \MC_ARK_ARC_1_0/temp4[109] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_13_4  ( .A1(\RI5[0][19] ), .A2(\RI5[0][175] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[109] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_13_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[79] ), 
        .A2(\RI5[0][55] ), .Z(\MC_ARK_ARC_1_0/temp2[109] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_13_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[109] ), 
        .A2(\RI5[0][103] ), .Z(\MC_ARK_ARC_1_0/temp1[109] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_13_3  ( .A1(\SB2_0_10/buf_output[2] ), .A2(n201), 
        .Z(\MC_ARK_ARC_1_0/temp4[110] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_13_2  ( .A1(\RI5[0][147] ), .A2(n557), .Z(
        \MC_ARK_ARC_1_0/temp4[111] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_13_1  ( .A1(\MC_ARK_ARC_1_0/temp4[112] ), .A2(
        \MC_ARK_ARC_1_0/temp3[112] ), .Z(\MC_ARK_ARC_1_0/temp6[112] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_13_1  ( .A1(\RI5[0][148] ), .A2(n553), .Z(
        \MC_ARK_ARC_1_0/temp4[112] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_13_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[22] ), 
        .A2(\RI5[0][178] ), .Z(\MC_ARK_ARC_1_0/temp3[112] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_13_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[82] ), 
        .A2(\RI5[0][58] ), .Z(\MC_ARK_ARC_1_0/temp2[112] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_13_0  ( .A1(\RI5[0][149] ), .A2(n235), .Z(
        \MC_ARK_ARC_1_0/temp4[113] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_12_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[150] ), 
        .A2(n243), .Z(\MC_ARK_ARC_1_0/temp4[114] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_12_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[180] ), 
        .A2(\RI5[0][24] ), .Z(\MC_ARK_ARC_1_0/temp3[114] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_12_5  ( .A1(\RI5[0][60] ), .A2(\RI5[0][84] ), .Z(
        \MC_ARK_ARC_1_0/temp2[114] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_12_5  ( .A1(\RI5[0][114] ), .A2(\RI5[0][108] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[114] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_12_4  ( .A1(\MC_ARK_ARC_1_0/temp4[115] ), .A2(
        \MC_ARK_ARC_1_0/temp3[115] ), .Z(\MC_ARK_ARC_1_0/temp6[115] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_12_4  ( .A1(\RI5[0][151] ), .A2(n540), .Z(
        \MC_ARK_ARC_1_0/temp4[115] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_12_4  ( .A1(\RI5[0][181] ), .A2(\RI5[0][25] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[115] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_12_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[61] ), 
        .A2(\RI5[0][85] ), .Z(\MC_ARK_ARC_1_0/temp2[115] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_12_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[115] ), 
        .A2(\MC_ARK_ARC_1_0/buf_datainput[109] ), .Z(
        \MC_ARK_ARC_1_0/temp1[115] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_12_3  ( .A1(\RI5[0][152] ), .A2(n535), .Z(
        \MC_ARK_ARC_1_0/temp4[116] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_12_3  ( .A1(\RI5[0][110] ), .A2(\RI5[0][116] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[116] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_12_2  ( .A1(\RI5[0][153] ), .A2(n198), .Z(
        \MC_ARK_ARC_1_0/temp4[117] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_12_1  ( .A1(\MC_ARK_ARC_1_0/temp6[118] ), .A2(
        \MC_ARK_ARC_1_0/temp5[118] ), .Z(\MC_ARK_ARC_1_0/buf_output[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_12_1  ( .A1(\MC_ARK_ARC_1_0/temp3[118] ), .A2(
        \MC_ARK_ARC_1_0/temp4[118] ), .Z(\MC_ARK_ARC_1_0/temp6[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_12_1  ( .A1(\MC_ARK_ARC_1_0/temp2[118] ), .A2(
        \MC_ARK_ARC_1_0/temp1[118] ), .Z(\MC_ARK_ARC_1_0/temp5[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_12_1  ( .A1(\RI5[0][154] ), .A2(n212), .Z(
        \MC_ARK_ARC_1_0/temp4[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_12_1  ( .A1(\RI5[0][184] ), .A2(\RI5[0][28] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_12_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[88] ), 
        .A2(\RI5[0][64] ), .Z(\MC_ARK_ARC_1_0/temp2[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_11_5  ( .A1(\MC_ARK_ARC_1_0/temp2[120] ), .A2(
        \MC_ARK_ARC_1_0/temp1[120] ), .Z(\MC_ARK_ARC_1_0/temp5[120] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_11_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[156] ), 
        .A2(n516), .Z(\MC_ARK_ARC_1_0/temp4[120] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_11_5  ( .A1(\RI5[0][186] ), .A2(\RI5[0][30] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[120] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_11_5  ( .A1(\RI5[0][66] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[90] ), .Z(\MC_ARK_ARC_1_0/temp2[120] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_11_5  ( .A1(\RI5[0][120] ), .A2(\RI5[0][114] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[120] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_11_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[157] ), 
        .A2(n510), .Z(\MC_ARK_ARC_1_0/temp4[121] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_11_4  ( .A1(\RI5[0][121] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[115] ), .Z(\MC_ARK_ARC_1_0/temp1[121] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_11_3  ( .A1(\RI5[0][158] ), .A2(n181), .Z(
        \MC_ARK_ARC_1_0/temp4[122] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_11_3  ( .A1(\RI5[0][122] ), .A2(\RI5[0][116] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[122] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_11_2  ( .A1(\RI5[0][159] ), .A2(n154), .Z(
        \MC_ARK_ARC_1_0/temp4[123] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_11_2  ( .A1(\RI5[0][93] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[69] ), .Z(\MC_ARK_ARC_1_0/temp2[123] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_11_2  ( .A1(\RI5[0][117] ), .A2(\RI5[0][123] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[123] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_11_1  ( .A1(\RI5[0][160] ), .A2(n497), .Z(
        \MC_ARK_ARC_1_0/temp4[124] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_11_1  ( .A1(\RI5[0][34] ), .A2(\RI5[0][190] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[124] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_11_1  ( .A1(\RI5[0][94] ), .A2(\RI5[0][70] ), .Z(
        \MC_ARK_ARC_1_0/temp2[124] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_11_0  ( .A1(\RI5[0][161] ), .A2(n148), .Z(
        \MC_ARK_ARC_1_0/temp4[125] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_11_0  ( .A1(\RI5[0][125] ), .A2(\RI5[0][119] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[125] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_10_4  ( .A1(\RI5[0][163] ), .A2(n222), .Z(
        \MC_ARK_ARC_1_0/temp4[127] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_10_4  ( .A1(\RI5[0][37] ), .A2(\RI5[0][1] ), .Z(
        \MC_ARK_ARC_1_0/temp3[127] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_10_4  ( .A1(\RI5[0][97] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[73] ), .Z(\MC_ARK_ARC_1_0/temp2[127] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_10_4  ( .A1(\RI5[0][127] ), .A2(\RI5[0][121] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[127] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_10_3  ( .A1(\MC_ARK_ARC_1_0/temp3[128] ), .A2(
        \MC_ARK_ARC_1_0/temp4[128] ), .Z(\MC_ARK_ARC_1_0/temp6[128] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_10_3  ( .A1(\RI5[0][164] ), .A2(n475), .Z(
        \MC_ARK_ARC_1_0/temp4[128] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_10_3  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[2] ), 
        .A2(\RI5[0][38] ), .Z(\MC_ARK_ARC_1_0/temp3[128] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_10_2  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[165] ), 
        .A2(n470), .Z(\MC_ARK_ARC_1_0/temp4[129] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_10_2  ( .A1(\RI5[0][39] ), .A2(\RI5[0][3] ), .Z(
        \MC_ARK_ARC_1_0/temp3[129] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_10_2  ( .A1(\RI5[0][75] ), .A2(\RI5[0][99] ), .Z(
        \MC_ARK_ARC_1_0/temp2[129] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_10_1  ( .A1(\MC_ARK_ARC_1_0/temp2[130] ), .A2(
        \MC_ARK_ARC_1_0/temp1[130] ), .Z(\MC_ARK_ARC_1_0/temp5[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_10_1  ( .A1(\SB2_0_5/buf_output[4] ), .A2(n216), 
        .Z(\MC_ARK_ARC_1_0/temp4[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_10_1  ( .A1(\SB2_0_11/buf_output[4] ), .A2(
        \RI5[0][124] ), .Z(\MC_ARK_ARC_1_0/temp1[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_10_0  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[167] ), 
        .A2(n236), .Z(\MC_ARK_ARC_1_0/temp4[131] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_10_0  ( .A1(\RI5[0][5] ), .A2(\RI5[0][41] ), .Z(
        \MC_ARK_ARC_1_0/temp3[131] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_10_0  ( .A1(\RI5[0][125] ), .A2(\RI5[0][131] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[131] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_9_5  ( .A1(\RI5[0][168] ), .A2(n457), .Z(
        \MC_ARK_ARC_1_0/temp4[132] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_9_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[42] ), 
        .A2(\RI5[0][6] ), .Z(\MC_ARK_ARC_1_0/temp3[132] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_9_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[132] ), 
        .A2(\RI5[0][126] ), .Z(\MC_ARK_ARC_1_0/temp1[132] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_9_4  ( .A1(\RI5[0][169] ), .A2(n159), .Z(
        \MC_ARK_ARC_1_0/temp4[133] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_9_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[7] ), 
        .A2(\RI5[0][43] ), .Z(\MC_ARK_ARC_1_0/temp3[133] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_9_3  ( .A1(\RI5[0][170] ), .A2(n447), .Z(
        \MC_ARK_ARC_1_0/temp4[134] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_9_2  ( .A1(\RI5[0][171] ), .A2(n442), .Z(
        \MC_ARK_ARC_1_0/temp4[135] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_9_2  ( .A1(\RI5[0][9] ), .A2(\RI5[0][45] ), .Z(
        \MC_ARK_ARC_1_0/temp3[135] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_9_2  ( .A1(\RI5[0][129] ), .A2(\RI5[0][135] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[135] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_9_1  ( .A1(\MC_ARK_ARC_1_0/temp2[136] ), .A2(
        \MC_ARK_ARC_1_0/temp1[136] ), .Z(\MC_ARK_ARC_1_0/temp5[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_9_1  ( .A1(\RI5[0][172] ), .A2(n51), .Z(
        \MC_ARK_ARC_1_0/temp4[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_9_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[46] ), 
        .A2(\RI5[0][10] ), .Z(\MC_ARK_ARC_1_0/temp3[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_9_1  ( .A1(\RI5[0][106] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[82] ), .Z(\MC_ARK_ARC_1_0/temp2[136] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_9_1  ( .A1(\RI5[0][130] ), .A2(\RI5[0][136] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_9_0  ( .A1(\RI5[0][173] ), .A2(n65), .Z(
        \MC_ARK_ARC_1_0/temp4[137] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_8_5  ( .A1(\RI5[0][174] ), .A2(n182), .Z(
        \MC_ARK_ARC_1_0/temp4[138] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_8_4  ( .A1(\MC_ARK_ARC_1_0/temp3[139] ), .A2(
        \MC_ARK_ARC_1_0/temp4[139] ), .Z(\MC_ARK_ARC_1_0/temp6[139] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_8_4  ( .A1(\RI5[0][175] ), .A2(n555), .Z(
        \MC_ARK_ARC_1_0/temp4[139] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_8_4  ( .A1(\RI5[0][13] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[49] ), .Z(\MC_ARK_ARC_1_0/temp3[139] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_8_4  ( .A1(\RI5[0][85] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[109] ), .Z(\MC_ARK_ARC_1_0/temp2[139] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_8_4  ( .A1(\RI5[0][133] ), .A2(\RI5[0][139] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[139] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_8_3  ( .A1(\MC_ARK_ARC_1_0/temp4[140] ), .A2(
        \MC_ARK_ARC_1_0/temp3[140] ), .Z(\MC_ARK_ARC_1_0/temp6[140] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_8_3  ( .A1(\RI5[0][176] ), .A2(n115), .Z(
        \MC_ARK_ARC_1_0/temp4[140] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_8_3  ( .A1(\RI5[0][50] ), .A2(\RI5[0][14] ), .Z(
        \MC_ARK_ARC_1_0/temp3[140] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_8_2  ( .A1(\RI5[0][177] ), .A2(n227), .Z(
        \MC_ARK_ARC_1_0/temp4[141] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_8_2  ( .A1(\RI5[0][135] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[141] ), .Z(\MC_ARK_ARC_1_0/temp1[141] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_8_1  ( .A1(\MC_ARK_ARC_1_0/temp3[142] ), .A2(
        \MC_ARK_ARC_1_0/temp4[142] ), .Z(\MC_ARK_ARC_1_0/temp6[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_8_1  ( .A1(\RI5[0][178] ), .A2(n206), .Z(
        \MC_ARK_ARC_1_0/temp4[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_8_1  ( .A1(\RI5[0][52] ), .A2(\RI5[0][16] ), .Z(
        \MC_ARK_ARC_1_0/temp3[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_8_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[112] ), 
        .A2(\MC_ARK_ARC_1_0/buf_datainput[88] ), .Z(
        \MC_ARK_ARC_1_0/temp2[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_8_1  ( .A1(\RI5[0][142] ), .A2(\RI5[0][136] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_7_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[180] ), 
        .A2(n531), .Z(\MC_ARK_ARC_1_0/temp4[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_7_4  ( .A1(\RI5[0][181] ), .A2(n525), .Z(
        \MC_ARK_ARC_1_0/temp4[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_7_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[115] ), 
        .A2(\RI5[0][91] ), .Z(\MC_ARK_ARC_1_0/temp2[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_7_4  ( .A1(\RI5[0][145] ), .A2(\RI5[0][139] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_7_3  ( .A1(\MC_ARK_ARC_1_0/temp1[146] ), .A2(
        \MC_ARK_ARC_1_0/temp2[146] ), .Z(\MC_ARK_ARC_1_0/temp5[146] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_7_3  ( .A1(\RI5[0][116] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[92] ), .Z(\MC_ARK_ARC_1_0/temp2[146] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_7_3  ( .A1(\RI5[0][146] ), .A2(\RI5[0][140] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[146] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_7_2  ( .A1(\RI5[0][183] ), .A2(n146), .Z(
        \MC_ARK_ARC_1_0/temp4[147] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_7_2  ( .A1(\RI5[0][57] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[21] ), .Z(\MC_ARK_ARC_1_0/temp3[147] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_7_1  ( .A1(\RI5[0][184] ), .A2(n180), .Z(
        \MC_ARK_ARC_1_0/temp4[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_7_1  ( .A1(\RI5[0][94] ), .A2(\RI5[0][118] ), .Z(
        \MC_ARK_ARC_1_0/temp2[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_7_1  ( .A1(\RI5[0][148] ), .A2(\RI5[0][142] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_7_0  ( .A1(\RI5[0][185] ), .A2(n99), .Z(
        \MC_ARK_ARC_1_0/temp4[149] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_6_5  ( .A1(\MC_ARK_ARC_1_0/temp4[150] ), .A2(
        \MC_ARK_ARC_1_0/temp3[150] ), .Z(\MC_ARK_ARC_1_0/temp6[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_6_5  ( .A1(\MC_ARK_ARC_1_0/temp1[150] ), .A2(
        \MC_ARK_ARC_1_0/temp2[150] ), .Z(\MC_ARK_ARC_1_0/temp5[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_6_5  ( .A1(\RI5[0][186] ), .A2(n178), .Z(
        \MC_ARK_ARC_1_0/temp4[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_6_5  ( .A1(\RI5[0][60] ), .A2(\RI5[0][24] ), .Z(
        \MC_ARK_ARC_1_0/temp3[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_6_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[150] ), 
        .A2(\MC_ARK_ARC_1_0/buf_datainput[144] ), .Z(
        \MC_ARK_ARC_1_0/temp1[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_6_4  ( .A1(\MC_ARK_ARC_1_0/temp2[151] ), .A2(
        \MC_ARK_ARC_1_0/temp1[151] ), .Z(\MC_ARK_ARC_1_0/temp5[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_6_4  ( .A1(\RI5[0][187] ), .A2(n499), .Z(
        \MC_ARK_ARC_1_0/temp4[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_6_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[61] ), 
        .A2(\RI5[0][25] ), .Z(\MC_ARK_ARC_1_0/temp3[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_6_4  ( .A1(\RI5[0][121] ), .A2(\RI5[0][97] ), .Z(
        \MC_ARK_ARC_1_0/temp2[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_6_4  ( .A1(\RI5[0][151] ), .A2(\RI5[0][145] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_6_3  ( .A1(\MC_ARK_ARC_1_0/temp5[152] ), .A2(
        \MC_ARK_ARC_1_0/temp6[152] ), .Z(\MC_ARK_ARC_1_0/buf_output[152] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_6_3  ( .A1(\RI5[0][188] ), .A2(n494), .Z(
        \MC_ARK_ARC_1_0/temp4[152] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_6_2  ( .A1(\RI5[0][189] ), .A2(n144), .Z(
        \MC_ARK_ARC_1_0/temp4[153] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_6_2  ( .A1(\RI5[0][123] ), .A2(\RI5[0][99] ), .Z(
        \MC_ARK_ARC_1_0/temp2[153] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_6_1  ( .A1(\MC_ARK_ARC_1_0/temp5[154] ), .A2(
        \MC_ARK_ARC_1_0/temp6[154] ), .Z(\MC_ARK_ARC_1_0/buf_output[154] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_6_1  ( .A1(\MC_ARK_ARC_1_0/temp4[154] ), .A2(
        \MC_ARK_ARC_1_0/temp3[154] ), .Z(\MC_ARK_ARC_1_0/temp6[154] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_6_1  ( .A1(\RI5[0][190] ), .A2(n483), .Z(
        \MC_ARK_ARC_1_0/temp4[154] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_6_1  ( .A1(\RI5[0][64] ), .A2(\RI5[0][28] ), .Z(
        \MC_ARK_ARC_1_0/temp3[154] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_6_1  ( .A1(\RI5[0][124] ), .A2(\RI5[0][100] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[154] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_6_0  ( .A1(\MC_ARK_ARC_1_0/temp3[155] ), .A2(
        \MC_ARK_ARC_1_0/temp4[155] ), .Z(\MC_ARK_ARC_1_0/temp6[155] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_6_0  ( .A1(\RI5[0][191] ), .A2(n202), .Z(
        \MC_ARK_ARC_1_0/temp4[155] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_6_0  ( .A1(\RI5[0][65] ), .A2(\RI5[0][29] ), .Z(
        \MC_ARK_ARC_1_0/temp3[155] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_5_5  ( .A1(\MC_ARK_ARC_1_0/temp3[156] ), .A2(
        \MC_ARK_ARC_1_0/temp4[156] ), .Z(\MC_ARK_ARC_1_0/temp6[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_5_5  ( .A1(\RI5[0][0] ), .A2(n242), .Z(
        \MC_ARK_ARC_1_0/temp4[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_5_5  ( .A1(\RI5[0][66] ), .A2(\RI5[0][30] ), .Z(
        \MC_ARK_ARC_1_0/temp3[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_5_5  ( .A1(\RI5[0][126] ), .A2(\RI5[0][102] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_5_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[156] ), 
        .A2(\MC_ARK_ARC_1_0/buf_datainput[150] ), .Z(
        \MC_ARK_ARC_1_0/temp1[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_5_4  ( .A1(\RI5[0][1] ), .A2(n72), .Z(
        \MC_ARK_ARC_1_0/temp4[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_5_2  ( .A1(\RI5[0][3] ), .A2(n459), .Z(
        \MC_ARK_ARC_1_0/temp4[159] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_5_2  ( .A1(\RI5[0][33] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[69] ), .Z(\MC_ARK_ARC_1_0/temp3[159] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_5_1  ( .A1(\RI5[0][4] ), .A2(n203), .Z(
        \MC_ARK_ARC_1_0/temp4[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_5_1  ( .A1(\RI5[0][34] ), .A2(\RI5[0][70] ), .Z(
        \MC_ARK_ARC_1_0/temp3[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_5_1  ( .A1(\RI5[0][130] ), .A2(\RI5[0][106] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_5_0  ( .A1(\RI5[0][5] ), .A2(n165), .Z(
        \MC_ARK_ARC_1_0/temp4[161] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_5_0  ( .A1(\RI5[0][35] ), .A2(\RI5[0][71] ), .Z(
        \MC_ARK_ARC_1_0/temp3[161] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_5_0  ( .A1(\RI5[0][107] ), .A2(\RI5[0][131] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[161] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_5_0  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[155] ), 
        .A2(\RI5[0][161] ), .Z(\MC_ARK_ARC_1_0/temp1[161] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_4_5  ( .A1(\MC_ARK_ARC_1_0/temp4[162] ), .A2(
        \MC_ARK_ARC_1_0/temp3[162] ), .Z(\MC_ARK_ARC_1_0/temp6[162] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_4_5  ( .A1(\RI5[0][6] ), .A2(n238), .Z(
        \MC_ARK_ARC_1_0/temp4[162] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_4_5  ( .A1(\RI5[0][108] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[132] ), .Z(\MC_ARK_ARC_1_0/temp2[162] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_4_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[156] ), 
        .A2(\RI5[0][162] ), .Z(\MC_ARK_ARC_1_0/temp1[162] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_4_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[7] ), 
        .A2(n440), .Z(\MC_ARK_ARC_1_0/temp4[163] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_4_3  ( .A1(\RI5[0][8] ), .A2(n39), .Z(
        \MC_ARK_ARC_1_0/temp4[164] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_4_2  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[165] ), 
        .A2(\RI5[0][159] ), .Z(\MC_ARK_ARC_1_0/temp1[165] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_4_1  ( .A1(\RI5[0][10] ), .A2(n208), .Z(
        \MC_ARK_ARC_1_0/temp4[166] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_4_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[76] ), 
        .A2(\RI5[0][40] ), .Z(\MC_ARK_ARC_1_0/temp3[166] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_4_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[112] ), 
        .A2(\RI5[0][136] ), .Z(\MC_ARK_ARC_1_0/temp2[166] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_4_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[166] ), 
        .A2(\RI5[0][160] ), .Z(\MC_ARK_ARC_1_0/temp1[166] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_4_0  ( .A1(\RI5[0][11] ), .A2(n161), .Z(
        \MC_ARK_ARC_1_0/temp4[167] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_4_0  ( .A1(\RI5[0][41] ), .A2(\RI5[0][77] ), .Z(
        \MC_ARK_ARC_1_0/temp3[167] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_4_0  ( .A1(\RI5[0][137] ), .A2(\RI5[0][113] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[167] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_3_5  ( .A1(\MC_ARK_ARC_1_0/temp1[168] ), .A2(
        \MC_ARK_ARC_1_0/temp2[168] ), .Z(\MC_ARK_ARC_1_0/temp5[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_3_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[12] ), 
        .A2(n184), .Z(\MC_ARK_ARC_1_0/temp4[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_3_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[78] ), 
        .A2(\MC_ARK_ARC_1_0/buf_datainput[42] ), .Z(
        \MC_ARK_ARC_1_0/temp3[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_3_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[138] ), 
        .A2(\RI5[0][114] ), .Z(\MC_ARK_ARC_1_0/temp2[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_3_5  ( .A1(\RI5[0][168] ), .A2(\RI5[0][162] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_3_4  ( .A1(\MC_ARK_ARC_1_0/temp4[169] ), .A2(
        \MC_ARK_ARC_1_0/temp3[169] ), .Z(\MC_ARK_ARC_1_0/temp6[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_3_4  ( .A1(\MC_ARK_ARC_1_0/temp1[169] ), .A2(
        \MC_ARK_ARC_1_0/temp2[169] ), .Z(\MC_ARK_ARC_1_0/temp5[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_3_4  ( .A1(\RI5[0][13] ), .A2(n544), .Z(
        \MC_ARK_ARC_1_0/temp4[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_3_4  ( .A1(\RI5[0][43] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[79] ), .Z(\MC_ARK_ARC_1_0/temp3[169] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_3_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[115] ), 
        .A2(\RI5[0][139] ), .Z(\MC_ARK_ARC_1_0/temp2[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_3_4  ( .A1(\RI5[0][169] ), .A2(\RI5[0][163] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_3_3  ( .A1(\RI5[0][14] ), .A2(
        \MC_ARK_ARC_1_1/buf_keyinput[51] ), .Z(\MC_ARK_ARC_1_0/temp4[170] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_3_3  ( .A1(\RI5[0][140] ), .A2(\RI5[0][116] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[170] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_3_2  ( .A1(\MC_ARK_ARC_1_0/temp5[171] ), .A2(
        \MC_ARK_ARC_1_0/temp6[171] ), .Z(\MC_ARK_ARC_1_0/buf_output[171] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_3_2  ( .A1(\RI5[0][15] ), .A2(n534), .Z(
        \MC_ARK_ARC_1_0/temp4[171] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_3_1  ( .A1(\MC_ARK_ARC_1_0/temp4[172] ), .A2(
        \MC_ARK_ARC_1_0/temp3[172] ), .Z(\MC_ARK_ARC_1_0/temp6[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_3_1  ( .A1(\RI5[0][16] ), .A2(n122), .Z(
        \MC_ARK_ARC_1_0/temp4[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_3_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[46] ), 
        .A2(\MC_ARK_ARC_1_0/buf_datainput[82] ), .Z(
        \MC_ARK_ARC_1_0/temp3[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_3_1  ( .A1(\RI5[0][142] ), .A2(\RI5[0][118] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_3_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[166] ), 
        .A2(\RI5[0][172] ), .Z(\MC_ARK_ARC_1_0/temp1[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_3_0  ( .A1(\MC_ARK_ARC_1_0/temp3[173] ), .A2(
        \MC_ARK_ARC_1_0/temp4[173] ), .Z(\MC_ARK_ARC_1_0/temp6[173] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_3_0  ( .A1(\MC_ARK_ARC_1_0/temp1[173] ), .A2(
        \MC_ARK_ARC_1_0/temp2[173] ), .Z(\MC_ARK_ARC_1_0/temp5[173] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_3_0  ( .A1(\RI5[0][17] ), .A2(n523), .Z(
        \MC_ARK_ARC_1_0/temp4[173] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_3_0  ( .A1(\RI5[0][83] ), .A2(\RI5[0][47] ), .Z(
        \MC_ARK_ARC_1_0/temp3[173] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_3_0  ( .A1(\RI5[0][143] ), .A2(\RI5[0][119] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[173] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_3_0  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[167] ), 
        .A2(\RI5[0][173] ), .Z(\MC_ARK_ARC_1_0/temp1[173] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_2_5  ( .A1(\RI5[0][18] ), .A2(n519), .Z(
        \MC_ARK_ARC_1_0/temp4[174] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_2_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[144] ), 
        .A2(\RI5[0][120] ), .Z(\MC_ARK_ARC_1_0/temp2[174] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_2_4  ( .A1(\MC_ARK_ARC_1_0/temp4[175] ), .A2(
        \MC_ARK_ARC_1_0/temp3[175] ), .Z(\MC_ARK_ARC_1_0/temp6[175] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_2_4  ( .A1(\RI5[0][19] ), .A2(n83), .Z(
        \MC_ARK_ARC_1_0/temp4[175] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_2_4  ( .A1(\RI5[0][85] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[49] ), .Z(\MC_ARK_ARC_1_0/temp3[175] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_2_4  ( .A1(\RI5[0][145] ), .A2(\RI5[0][121] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[175] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_2_4  ( .A1(\RI5[0][169] ), .A2(\RI5[0][175] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[175] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_2_3  ( .A1(\RI5[0][176] ), .A2(\RI5[0][170] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[176] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_2_2  ( .A1(\MC_ARK_ARC_1_0/temp4[177] ), .A2(
        \MC_ARK_ARC_1_0/temp3[177] ), .Z(\MC_ARK_ARC_1_0/temp6[177] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_2_2  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[21] ), 
        .A2(n505), .Z(\MC_ARK_ARC_1_0/temp4[177] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_2_1  ( .A1(\MC_ARK_ARC_1_0/temp6[178] ), .A2(
        \MC_ARK_ARC_1_0/temp5[178] ), .Z(\MC_ARK_ARC_1_0/buf_output[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_2_1  ( .A1(\MC_ARK_ARC_1_0/temp3[178] ), .A2(
        \MC_ARK_ARC_1_0/temp4[178] ), .Z(\MC_ARK_ARC_1_0/temp6[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_2_1  ( .A1(\MC_ARK_ARC_1_0/temp2[178] ), .A2(
        \MC_ARK_ARC_1_0/temp1[178] ), .Z(\MC_ARK_ARC_1_0/temp5[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_2_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[22] ), 
        .A2(n500), .Z(\MC_ARK_ARC_1_0/temp4[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_2_1  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[88] ), 
        .A2(\RI5[0][52] ), .Z(\MC_ARK_ARC_1_0/temp3[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_2_1  ( .A1(\RI5[0][148] ), .A2(\RI5[0][124] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_2_1  ( .A1(\RI5[0][178] ), .A2(\RI5[0][172] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_2_0  ( .A1(\RI5[0][23] ), .A2(n82), .Z(
        \MC_ARK_ARC_1_0/temp4[179] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_2_0  ( .A1(\RI5[0][173] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[179] ), .Z(\MC_ARK_ARC_1_0/temp1[179] )
         );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_1_5  ( .A1(\RI5[0][24] ), .A2(n492), .Z(
        \MC_ARK_ARC_1_0/temp4[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_1_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[150] ), 
        .A2(\RI5[0][126] ), .Z(\MC_ARK_ARC_1_0/temp2[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X7_1_4  ( .A1(\MC_ARK_ARC_1_0/temp5[181] ), .A2(
        \MC_ARK_ARC_1_0/temp6[181] ), .Z(\MC_ARK_ARC_1_0/buf_output[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_1_4  ( .A1(\MC_ARK_ARC_1_0/temp3[181] ), .A2(
        \MC_ARK_ARC_1_0/temp4[181] ), .Z(\MC_ARK_ARC_1_0/temp6[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_1_4  ( .A1(\MC_ARK_ARC_1_0/temp2[181] ), .A2(
        \MC_ARK_ARC_1_0/temp1[181] ), .Z(\MC_ARK_ARC_1_0/temp5[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_1_4  ( .A1(\RI5[0][25] ), .A2(n486), .Z(
        \MC_ARK_ARC_1_0/temp4[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_1_4  ( .A1(\RI5[0][91] ), .A2(\RI5[0][55] ), .Z(
        \MC_ARK_ARC_1_0/temp3[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_1_4  ( .A1(\RI5[0][127] ), .A2(\RI5[0][151] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_1_4  ( .A1(\RI5[0][181] ), .A2(\RI5[0][175] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_1_3  ( .A1(\MC_ARK_ARC_1_0/temp3[182] ), .A2(
        \MC_ARK_ARC_1_0/temp4[182] ), .Z(\MC_ARK_ARC_1_0/temp6[182] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_1_3  ( .A1(\RI5[0][26] ), .A2(n27), .Z(
        \MC_ARK_ARC_1_0/temp4[182] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_1_2  ( .A1(\MC_ARK_ARC_1_0/temp3[183] ), .A2(
        \MC_ARK_ARC_1_0/temp4[183] ), .Z(\MC_ARK_ARC_1_0/temp6[183] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_1_2  ( .A1(\RI5[0][27] ), .A2(n114), .Z(
        \MC_ARK_ARC_1_0/temp4[183] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_1_1  ( .A1(\RI5[0][28] ), .A2(n226), .Z(
        \MC_ARK_ARC_1_0/temp4[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_1_1  ( .A1(\RI5[0][94] ), .A2(\RI5[0][58] ), .Z(
        \MC_ARK_ARC_1_0/temp3[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_1_1  ( .A1(\RI5[0][184] ), .A2(\RI5[0][178] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X6_1_0  ( .A1(\MC_ARK_ARC_1_0/temp3[185] ), .A2(
        \MC_ARK_ARC_1_0/temp4[185] ), .Z(\MC_ARK_ARC_1_0/temp6[185] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_1_0  ( .A1(\RI5[0][29] ), .A2(n135), .Z(
        \MC_ARK_ARC_1_0/temp4[185] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_1_0  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[155] ), 
        .A2(\RI5[0][131] ), .Z(\MC_ARK_ARC_1_0/temp2[185] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_0_5  ( .A1(\RI5[0][30] ), .A2(n461), .Z(
        \MC_ARK_ARC_1_0/temp4[186] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_0_5  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[96] ), 
        .A2(\RI5[0][60] ), .Z(\MC_ARK_ARC_1_0/temp3[186] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_0_4  ( .A1(\MC_ARK_ARC_1_0/temp1[187] ), .A2(
        \MC_ARK_ARC_1_0/temp2[187] ), .Z(\MC_ARK_ARC_1_0/temp5[187] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_0_4  ( .A1(\RI5[0][31] ), .A2(n143), .Z(
        \MC_ARK_ARC_1_0/temp4[187] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_0_4  ( .A1(\MC_ARK_ARC_1_0/buf_datainput[157] ), 
        .A2(\RI5[0][133] ), .Z(\MC_ARK_ARC_1_0/temp2[187] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_0_3  ( .A1(\SB2_0_29/buf_output[2] ), .A2(n130), 
        .Z(\MC_ARK_ARC_1_0/temp4[188] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_0_2  ( .A1(\RI5[0][33] ), .A2(n446), .Z(
        \MC_ARK_ARC_1_0/temp4[189] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_0_2  ( .A1(\RI5[0][189] ), .A2(\RI5[0][183] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[189] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X5_0_1  ( .A1(\MC_ARK_ARC_1_0/temp1[190] ), .A2(
        \MC_ARK_ARC_1_0/temp2[190] ), .Z(\MC_ARK_ARC_1_0/temp5[190] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_0_1  ( .A1(\RI5[0][34] ), .A2(n225), .Z(
        \MC_ARK_ARC_1_0/temp4[190] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X3_0_1  ( .A1(\RI5[0][64] ), .A2(\RI5[0][100] ), .Z(
        \MC_ARK_ARC_1_0/temp3[190] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X2_0_1  ( .A1(\RI5[0][160] ), .A2(\RI5[0][136] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[190] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X1_0_1  ( .A1(\RI5[0][184] ), .A2(\RI5[0][190] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[190] ) );
  XOR2_X1 \MC_ARK_ARC_1_0/X4_0_0  ( .A1(\RI5[0][35] ), .A2(n80), .Z(
        \MC_ARK_ARC_1_0/temp4[191] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_31_5  ( .A1(\RI5[1][36] ), .A2(n169), .Z(
        \MC_ARK_ARC_1_1/temp4[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_31_5  ( .A1(\RI5[1][102] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[66] ), .Z(\MC_ARK_ARC_1_1/temp3[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_31_4  ( .A1(\MC_ARK_ARC_1_1/temp3[1] ), .A2(
        \MC_ARK_ARC_1_1/temp4[1] ), .Z(\MC_ARK_ARC_1_1/temp6[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_31_4  ( .A1(\RI5[1][37] ), .A2(n36), .Z(
        \MC_ARK_ARC_1_1/temp4[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_31_4  ( .A1(\RI5[1][67] ), .A2(\RI5[1][103] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_31_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[163] ), 
        .A2(\MC_ARK_ARC_1_1/buf_datainput[139] ), .Z(\MC_ARK_ARC_1_1/temp2[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_31_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[1] ), 
        .A2(\MC_ARK_ARC_1_1/buf_datainput[187] ), .Z(\MC_ARK_ARC_1_1/temp1[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_31_3  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[38] ), 
        .A2(n472), .Z(\MC_ARK_ARC_1_1/temp4[2] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_31_2  ( .A1(\RI5[1][39] ), .A2(n439), .Z(
        \MC_ARK_ARC_1_1/temp4[3] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_31_2  ( .A1(\RI5[1][3] ), .A2(\RI5[1][189] ), .Z(
        \MC_ARK_ARC_1_1/temp1[3] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_31_1  ( .A1(\RI5[1][40] ), .A2(n71), .Z(
        \MC_ARK_ARC_1_1/temp4[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_31_1  ( .A1(\RI5[1][166] ), .A2(\RI5[1][142] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_31_1  ( .A1(\RI5[1][4] ), .A2(\RI5[1][190] ), .Z(
        \MC_ARK_ARC_1_1/temp1[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_31_0  ( .A1(\MC_ARK_ARC_1_1/temp3[5] ), .A2(
        \MC_ARK_ARC_1_1/temp4[5] ), .Z(\MC_ARK_ARC_1_1/temp6[5] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_31_0  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[41] ), 
        .A2(n504), .Z(\MC_ARK_ARC_1_1/temp4[5] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_30_5  ( .A1(\MC_ARK_ARC_1_1/temp4[6] ), .A2(
        \MC_ARK_ARC_1_1/temp3[6] ), .Z(\MC_ARK_ARC_1_1/temp6[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_30_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[42] ), 
        .A2(n49), .Z(\MC_ARK_ARC_1_1/temp4[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_30_5  ( .A1(\RI5[1][168] ), .A2(\RI5[1][144] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_30_4  ( .A1(\RI5[1][43] ), .A2(n241), .Z(
        \MC_ARK_ARC_1_1/temp4[7] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_30_4  ( .A1(\RI5[1][7] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[1] ), .Z(\MC_ARK_ARC_1_1/temp1[7] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_30_2  ( .A1(\RI5[1][45] ), .A2(n187), .Z(
        \MC_ARK_ARC_1_1/temp4[9] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_30_2  ( .A1(\RI5[1][75] ), .A2(\RI5[1][111] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[9] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_30_1  ( .A1(\RI5[1][46] ), .A2(n466), .Z(
        \MC_ARK_ARC_1_1/temp4[10] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_30_0  ( .A1(\MC_ARK_ARC_1_1/temp3[11] ), .A2(
        \MC_ARK_ARC_1_1/temp4[11] ), .Z(\MC_ARK_ARC_1_1/temp6[11] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_30_0  ( .A1(\RI5[1][47] ), .A2(n179), .Z(
        \MC_ARK_ARC_1_1/temp4[11] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_30_0  ( .A1(\RI5[1][113] ), .A2(\RI5[1][77] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[11] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_29_5  ( .A1(\RI5[1][48] ), .A2(n218), .Z(
        \MC_ARK_ARC_1_1/temp4[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_29_5  ( .A1(\RI5[1][114] ), .A2(\RI5[1][78] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_29_5  ( .A1(\RI5[1][174] ), .A2(\RI5[1][150] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_29_4  ( .A1(\RI5[1][49] ), .A2(n190), .Z(
        \MC_ARK_ARC_1_1/temp4[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_29_4  ( .A1(\RI5[1][115] ), .A2(\RI5[1][79] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_29_4  ( .A1(\RI5[1][151] ), .A2(\RI5[1][175] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_29_3  ( .A1(\SB2_1_26/buf_output[2] ), .A2(n131), 
        .Z(\MC_ARK_ARC_1_1/temp4[14] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_29_1  ( .A1(\RI5[1][52] ), .A2(n528), .Z(
        \MC_ARK_ARC_1_1/temp4[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_29_1  ( .A1(\RI5[1][82] ), .A2(\RI5[1][118] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_29_1  ( .A1(\RI5[1][16] ), .A2(\RI5[1][10] ), .Z(
        \MC_ARK_ARC_1_1/temp1[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_29_0  ( .A1(\RI5[1][53] ), .A2(n138), .Z(
        \MC_ARK_ARC_1_1/temp4[17] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_28_5  ( .A1(\MC_ARK_ARC_1_1/temp1[18] ), .A2(
        \MC_ARK_ARC_1_1/temp2[18] ), .Z(\MC_ARK_ARC_1_1/temp5[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_28_5  ( .A1(\RI5[1][54] ), .A2(n236), .Z(
        \MC_ARK_ARC_1_1/temp4[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_28_5  ( .A1(\RI5[1][120] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[84] ), .Z(\MC_ARK_ARC_1_1/temp3[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_28_5  ( .A1(\RI5[1][180] ), .A2(\RI5[1][156] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_28_5  ( .A1(\SB2_1_2/buf_output[0] ), .A2(
        \RI5[1][18] ), .Z(\MC_ARK_ARC_1_1/temp1[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_28_4  ( .A1(\MC_ARK_ARC_1_1/temp3[19] ), .A2(
        \MC_ARK_ARC_1_1/temp4[19] ), .Z(\MC_ARK_ARC_1_1/temp6[19] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_28_4  ( .A1(\RI5[1][55] ), .A2(n559), .Z(
        \MC_ARK_ARC_1_1/temp4[19] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_28_3  ( .A1(\RI5[1][56] ), .A2(n53), .Z(
        \MC_ARK_ARC_1_1/temp4[20] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_28_2  ( .A1(\MC_ARK_ARC_1_1/temp3[21] ), .A2(
        \MC_ARK_ARC_1_1/temp4[21] ), .Z(\MC_ARK_ARC_1_1/temp6[21] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_28_2  ( .A1(\RI5[1][57] ), .A2(n494), .Z(
        \MC_ARK_ARC_1_1/temp4[21] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_28_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[123] ), 
        .A2(\RI5[1][87] ), .Z(\MC_ARK_ARC_1_1/temp3[21] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_28_2  ( .A1(\RI5[1][183] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[159] ), .Z(\MC_ARK_ARC_1_1/temp2[21] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_28_2  ( .A1(\RI5[1][21] ), .A2(\RI5[1][15] ), .Z(
        \MC_ARK_ARC_1_1/temp1[21] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_28_1  ( .A1(\MC_ARK_ARC_1_1/temp6[22] ), .A2(
        \MC_ARK_ARC_1_1/temp5[22] ), .Z(\MC_ARK_ARC_1_1/buf_output[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_28_1  ( .A1(\MC_ARK_ARC_1_1/temp1[22] ), .A2(
        \MC_ARK_ARC_1_1/temp2[22] ), .Z(\MC_ARK_ARC_1_1/temp5[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_28_1  ( .A1(\RI5[1][58] ), .A2(n459), .Z(
        \MC_ARK_ARC_1_1/temp4[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_28_1  ( .A1(\RI5[1][184] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[160] ), .Z(\MC_ARK_ARC_1_1/temp2[22] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_28_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[22] ), 
        .A2(\RI5[1][16] ), .Z(\MC_ARK_ARC_1_1/temp1[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_27_5  ( .A1(\MC_ARK_ARC_1_1/temp6[24] ), .A2(
        \MC_ARK_ARC_1_1/temp5[24] ), .Z(\MC_ARK_ARC_1_1/buf_output[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_27_5  ( .A1(\MC_ARK_ARC_1_1/temp3[24] ), .A2(
        \MC_ARK_ARC_1_1/temp4[24] ), .Z(\MC_ARK_ARC_1_1/temp6[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_27_5  ( .A1(\MC_ARK_ARC_1_1/temp1[24] ), .A2(
        \MC_ARK_ARC_1_1/temp2[24] ), .Z(\MC_ARK_ARC_1_1/temp5[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_27_5  ( .A1(\RI5[1][60] ), .A2(n97), .Z(
        \MC_ARK_ARC_1_1/temp4[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_27_5  ( .A1(\RI5[1][90] ), .A2(\RI5[1][126] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_27_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[186] ), 
        .A2(\RI5[1][162] ), .Z(\MC_ARK_ARC_1_1/temp2[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_27_5  ( .A1(\RI5[1][24] ), .A2(\RI5[1][18] ), .Z(
        \MC_ARK_ARC_1_1/temp1[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_27_4  ( .A1(\MC_ARK_ARC_1_1/temp3[25] ), .A2(
        \MC_ARK_ARC_1_1/temp4[25] ), .Z(\MC_ARK_ARC_1_1/temp6[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_27_4  ( .A1(\RI5[1][61] ), .A2(n229), .Z(
        \MC_ARK_ARC_1_1/temp4[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_27_4  ( .A1(\RI5[1][91] ), .A2(\RI5[1][127] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_27_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[163] ), 
        .A2(\MC_ARK_ARC_1_1/buf_datainput[187] ), .Z(
        \MC_ARK_ARC_1_1/temp2[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_27_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[25] ), 
        .A2(\RI5[1][19] ), .Z(\MC_ARK_ARC_1_1/temp1[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_27_3  ( .A1(\RI5[1][62] ), .A2(n456), .Z(
        \MC_ARK_ARC_1_1/temp4[26] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_27_3  ( .A1(\RI5[1][26] ), .A2(\RI5[1][20] ), .Z(
        \MC_ARK_ARC_1_1/temp1[26] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_27_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[63] ), 
        .A2(n84), .Z(\MC_ARK_ARC_1_1/temp4[27] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_27_2  ( .A1(\RI5[1][165] ), .A2(\RI5[1][189] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[27] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_27_1  ( .A1(\MC_ARK_ARC_1_1/temp3[28] ), .A2(
        \MC_ARK_ARC_1_1/temp4[28] ), .Z(\MC_ARK_ARC_1_1/temp6[28] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_27_1  ( .A1(\RI5[1][64] ), .A2(n521), .Z(
        \MC_ARK_ARC_1_1/temp4[28] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_27_1  ( .A1(\RI5[1][130] ), .A2(\RI5[1][94] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[28] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_27_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[28] ), 
        .A2(\MC_ARK_ARC_1_1/buf_datainput[22] ), .Z(\MC_ARK_ARC_1_1/temp1[28] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_27_0  ( .A1(\RI5[1][167] ), .A2(\RI5[1][191] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[29] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_27_0  ( .A1(\RI5[1][23] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[29] ), .Z(\MC_ARK_ARC_1_1/temp1[29] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_26_5  ( .A1(\MC_ARK_ARC_1_1/temp1[30] ), .A2(
        \MC_ARK_ARC_1_1/temp2[30] ), .Z(\MC_ARK_ARC_1_1/temp5[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_26_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[66] ), 
        .A2(n140), .Z(\MC_ARK_ARC_1_1/temp4[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_26_5  ( .A1(\RI5[1][0] ), .A2(\RI5[1][168] ), .Z(
        \MC_ARK_ARC_1_1/temp2[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_26_5  ( .A1(\RI5[1][24] ), .A2(\RI5[1][30] ), .Z(
        \MC_ARK_ARC_1_1/temp1[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_26_4  ( .A1(\MC_ARK_ARC_1_1/temp5[31] ), .A2(
        \MC_ARK_ARC_1_1/temp6[31] ), .Z(\MC_ARK_ARC_1_1/buf_output[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_26_4  ( .A1(\RI5[1][67] ), .A2(n239), .Z(
        \MC_ARK_ARC_1_1/temp4[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_26_4  ( .A1(\RI5[1][133] ), .A2(\RI5[1][97] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_26_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[31] ), 
        .A2(\MC_ARK_ARC_1_1/buf_datainput[25] ), .Z(\MC_ARK_ARC_1_1/temp1[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_26_3  ( .A1(\RI5[1][68] ), .A2(n518), .Z(
        \MC_ARK_ARC_1_1/temp4[32] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_26_3  ( .A1(\RI5[1][134] ), .A2(\RI5[1][98] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[32] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_26_3  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[170] ), 
        .A2(\RI5[1][2] ), .Z(\MC_ARK_ARC_1_1/temp2[32] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_26_2  ( .A1(\RI5[1][69] ), .A2(n485), .Z(
        \MC_ARK_ARC_1_1/temp4[33] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_26_2  ( .A1(n1383), .A2(\RI5[1][27] ), .Z(
        \MC_ARK_ARC_1_1/temp1[33] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_26_1  ( .A1(\MC_ARK_ARC_1_1/temp1[34] ), .A2(
        \MC_ARK_ARC_1_1/temp2[34] ), .Z(\MC_ARK_ARC_1_1/temp5[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_26_1  ( .A1(\RI5[1][70] ), .A2(n450), .Z(
        \MC_ARK_ARC_1_1/temp4[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_26_1  ( .A1(\RI5[1][4] ), .A2(\RI5[1][172] ), .Z(
        \MC_ARK_ARC_1_1/temp2[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_26_1  ( .A1(\RI5[1][34] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[28] ), .Z(\MC_ARK_ARC_1_1/temp1[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_26_0  ( .A1(\RI5[1][71] ), .A2(n548), .Z(
        \MC_ARK_ARC_1_1/temp4[35] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_26_0  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[35] ), 
        .A2(\MC_ARK_ARC_1_1/buf_datainput[29] ), .Z(\MC_ARK_ARC_1_1/temp1[35] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_25_5  ( .A1(\MC_ARK_ARC_1_1/temp3[36] ), .A2(
        \MC_ARK_ARC_1_1/temp4[36] ), .Z(\MC_ARK_ARC_1_1/temp6[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_25_5  ( .A1(\RI5[1][72] ), .A2(n172), .Z(
        \MC_ARK_ARC_1_1/temp4[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_25_5  ( .A1(\RI5[1][138] ), .A2(\RI5[1][102] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_25_4  ( .A1(\MC_ARK_ARC_1_1/temp3[37] ), .A2(
        \MC_ARK_ARC_1_1/temp4[37] ), .Z(\MC_ARK_ARC_1_1/temp6[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_25_4  ( .A1(\MC_ARK_ARC_1_1/temp2[37] ), .A2(
        \MC_ARK_ARC_1_1/temp1[37] ), .Z(\MC_ARK_ARC_1_1/temp5[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_25_4  ( .A1(\RI5[1][73] ), .A2(n59), .Z(
        \MC_ARK_ARC_1_1/temp4[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_25_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[31] ), 
        .A2(\RI5[1][37] ), .Z(\MC_ARK_ARC_1_1/temp1[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_25_3  ( .A1(\MC_ARK_ARC_1_1/temp6[38] ), .A2(
        \MC_ARK_ARC_1_1/temp5[38] ), .Z(\MC_ARK_ARC_1_1/buf_output[38] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_25_3  ( .A1(\MC_ARK_ARC_1_1/temp4[38] ), .A2(
        \MC_ARK_ARC_1_1/temp3[38] ), .Z(\MC_ARK_ARC_1_1/temp6[38] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_25_3  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[74] ), 
        .A2(n448), .Z(\MC_ARK_ARC_1_1/temp4[38] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_25_3  ( .A1(\RI5[1][140] ), .A2(\RI5[1][104] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[38] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_25_2  ( .A1(\MC_ARK_ARC_1_1/temp3[39] ), .A2(
        \MC_ARK_ARC_1_1/temp4[39] ), .Z(\MC_ARK_ARC_1_1/temp6[39] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_25_2  ( .A1(\RI5[1][75] ), .A2(n545), .Z(
        \MC_ARK_ARC_1_1/temp4[39] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_25_2  ( .A1(n1383), .A2(\RI5[1][39] ), .Z(
        \MC_ARK_ARC_1_1/temp1[39] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_25_0  ( .A1(\RI5[1][77] ), .A2(n478), .Z(
        \MC_ARK_ARC_1_1/temp4[41] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_25_0  ( .A1(\RI5[1][11] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[179] ), .Z(\MC_ARK_ARC_1_1/temp2[41] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_24_5  ( .A1(\MC_ARK_ARC_1_1/temp5[42] ), .A2(
        \MC_ARK_ARC_1_1/temp6[42] ), .Z(\MC_ARK_ARC_1_1/buf_output[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_24_5  ( .A1(\MC_ARK_ARC_1_1/temp3[42] ), .A2(
        \MC_ARK_ARC_1_1/temp4[42] ), .Z(\MC_ARK_ARC_1_1/temp6[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_24_5  ( .A1(\RI5[1][78] ), .A2(n444), .Z(
        \MC_ARK_ARC_1_1/temp4[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_24_5  ( .A1(\RI5[1][144] ), .A2(\RI5[1][108] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_24_5  ( .A1(\RI5[1][12] ), .A2(\RI5[1][180] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_24_5  ( .A1(\RI5[1][36] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[42] ), .Z(\MC_ARK_ARC_1_1/temp1[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_24_4  ( .A1(\MC_ARK_ARC_1_1/temp1[43] ), .A2(
        \MC_ARK_ARC_1_1/temp2[43] ), .Z(\MC_ARK_ARC_1_1/temp5[43] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_24_4  ( .A1(\RI5[1][79] ), .A2(n243), .Z(
        \MC_ARK_ARC_1_1/temp4[43] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_24_4  ( .A1(\RI5[1][145] ), .A2(\RI5[1][109] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[43] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_24_4  ( .A1(\RI5[1][181] ), .A2(\RI5[1][13] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[43] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_24_4  ( .A1(\RI5[1][37] ), .A2(\RI5[1][43] ), .Z(
        \MC_ARK_ARC_1_1/temp1[43] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_24_2  ( .A1(\MC_ARK_ARC_1_1/temp4[45] ), .A2(
        \MC_ARK_ARC_1_1/temp3[45] ), .Z(\MC_ARK_ARC_1_1/temp6[45] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_24_2  ( .A1(\RI5[1][81] ), .A2(n475), .Z(
        \MC_ARK_ARC_1_1/temp4[45] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_24_1  ( .A1(\RI5[1][82] ), .A2(n442), .Z(
        \MC_ARK_ARC_1_1/temp4[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_24_1  ( .A1(\RI5[1][148] ), .A2(\RI5[1][112] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_24_1  ( .A1(\RI5[1][46] ), .A2(\RI5[1][40] ), .Z(
        \MC_ARK_ARC_1_1/temp1[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_24_0  ( .A1(\MC_ARK_ARC_1_1/temp3[47] ), .A2(
        \MC_ARK_ARC_1_1/temp4[47] ), .Z(\MC_ARK_ARC_1_1/temp6[47] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_24_0  ( .A1(\RI5[1][83] ), .A2(n206), .Z(
        \MC_ARK_ARC_1_1/temp4[47] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_23_5  ( .A1(\MC_ARK_ARC_1_1/temp3[48] ), .A2(
        \MC_ARK_ARC_1_1/temp4[48] ), .Z(\MC_ARK_ARC_1_1/temp6[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_23_5  ( .A1(\MC_ARK_ARC_1_1/temp1[48] ), .A2(
        \MC_ARK_ARC_1_1/temp2[48] ), .Z(\MC_ARK_ARC_1_1/temp5[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_23_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[84] ), 
        .A2(n163), .Z(\MC_ARK_ARC_1_1/temp4[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_23_5  ( .A1(\RI5[1][150] ), .A2(\RI5[1][114] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_23_5  ( .A1(\RI5[1][18] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[186] ), .Z(\MC_ARK_ARC_1_1/temp2[48] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_23_5  ( .A1(\RI5[1][48] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[42] ), .Z(\MC_ARK_ARC_1_1/temp1[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_23_4  ( .A1(\MC_ARK_ARC_1_1/temp1[49] ), .A2(
        \MC_ARK_ARC_1_1/temp2[49] ), .Z(\MC_ARK_ARC_1_1/temp5[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_23_4  ( .A1(\RI5[1][85] ), .A2(n242), .Z(
        \MC_ARK_ARC_1_1/temp4[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_23_4  ( .A1(\RI5[1][115] ), .A2(\RI5[1][151] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_23_4  ( .A1(\RI5[1][19] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[187] ), .Z(\MC_ARK_ARC_1_1/temp2[49] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_23_4  ( .A1(\RI5[1][49] ), .A2(\RI5[1][43] ), .Z(
        \MC_ARK_ARC_1_1/temp1[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_23_3  ( .A1(\RI5[1][86] ), .A2(n440), .Z(
        \MC_ARK_ARC_1_1/temp4[50] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_23_2  ( .A1(\MC_ARK_ARC_1_1/temp3[51] ), .A2(
        \MC_ARK_ARC_1_1/temp4[51] ), .Z(\MC_ARK_ARC_1_1/temp6[51] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_23_2  ( .A1(\MC_ARK_ARC_1_1/temp2[51] ), .A2(
        \MC_ARK_ARC_1_1/temp1[51] ), .Z(\MC_ARK_ARC_1_1/temp5[51] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_23_2  ( .A1(\RI5[1][87] ), .A2(
        \MC_ARK_ARC_1_1/buf_keyinput[51] ), .Z(\MC_ARK_ARC_1_1/temp4[51] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_23_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[153] ), 
        .A2(\RI5[1][117] ), .Z(\MC_ARK_ARC_1_1/temp3[51] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_23_2  ( .A1(\RI5[1][189] ), .A2(\RI5[1][21] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[51] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_23_1  ( .A1(\RI5[1][88] ), .A2(n505), .Z(
        \MC_ARK_ARC_1_1/temp4[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_23_1  ( .A1(\RI5[1][52] ), .A2(\RI5[1][46] ), .Z(
        \MC_ARK_ARC_1_1/temp1[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_22_5  ( .A1(\MC_ARK_ARC_1_1/temp6[54] ), .A2(
        \MC_ARK_ARC_1_1/temp5[54] ), .Z(\MC_ARK_ARC_1_1/buf_output[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_22_5  ( .A1(\MC_ARK_ARC_1_1/temp3[54] ), .A2(
        \MC_ARK_ARC_1_1/temp4[54] ), .Z(\MC_ARK_ARC_1_1/temp6[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_22_5  ( .A1(\MC_ARK_ARC_1_1/temp2[54] ), .A2(
        \MC_ARK_ARC_1_1/temp1[54] ), .Z(\MC_ARK_ARC_1_1/temp5[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_22_5  ( .A1(\RI5[1][90] ), .A2(n437), .Z(
        \MC_ARK_ARC_1_1/temp4[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_22_5  ( .A1(\RI5[1][156] ), .A2(\RI5[1][120] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_22_5  ( .A1(\RI5[1][24] ), .A2(\RI5[1][0] ), .Z(
        \MC_ARK_ARC_1_1/temp2[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_22_5  ( .A1(\RI5[1][54] ), .A2(\RI5[1][48] ), .Z(
        \MC_ARK_ARC_1_1/temp1[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_22_4  ( .A1(\MC_ARK_ARC_1_1/temp6[55] ), .A2(
        \MC_ARK_ARC_1_1/temp5[55] ), .Z(\MC_ARK_ARC_1_1/buf_output[55] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_22_4  ( .A1(\MC_ARK_ARC_1_1/temp3[55] ), .A2(
        \MC_ARK_ARC_1_1/temp4[55] ), .Z(\MC_ARK_ARC_1_1/temp6[55] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_22_4  ( .A1(\MC_ARK_ARC_1_1/temp2[55] ), .A2(
        \MC_ARK_ARC_1_1/temp1[55] ), .Z(\MC_ARK_ARC_1_1/temp5[55] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_22_4  ( .A1(\RI5[1][91] ), .A2(n244), .Z(
        \MC_ARK_ARC_1_1/temp4[55] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_22_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[25] ), 
        .A2(\MC_ARK_ARC_1_1/buf_datainput[1] ), .Z(\MC_ARK_ARC_1_1/temp2[55] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_22_4  ( .A1(\RI5[1][55] ), .A2(\RI5[1][49] ), .Z(
        \MC_ARK_ARC_1_1/temp1[55] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_22_3  ( .A1(\MC_ARK_ARC_1_1/temp3[56] ), .A2(
        \MC_ARK_ARC_1_1/temp4[56] ), .Z(\MC_ARK_ARC_1_1/temp6[56] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_22_3  ( .A1(\RI5[1][92] ), .A2(n79), .Z(
        \MC_ARK_ARC_1_1/temp4[56] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_22_3  ( .A1(\RI5[1][158] ), .A2(\RI5[1][122] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[56] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_22_2  ( .A1(\MC_ARK_ARC_1_1/temp4[57] ), .A2(
        \MC_ARK_ARC_1_1/temp3[57] ), .Z(\MC_ARK_ARC_1_1/temp6[57] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_22_2  ( .A1(\RI5[1][93] ), .A2(n467), .Z(
        \MC_ARK_ARC_1_1/temp4[57] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_22_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[123] ), 
        .A2(\MC_ARK_ARC_1_1/buf_datainput[159] ), .Z(
        \MC_ARK_ARC_1_1/temp3[57] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_22_1  ( .A1(\MC_ARK_ARC_1_1/temp4[58] ), .A2(
        \MC_ARK_ARC_1_1/temp3[58] ), .Z(\MC_ARK_ARC_1_1/temp6[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_22_1  ( .A1(\RI5[1][94] ), .A2(n564), .Z(
        \MC_ARK_ARC_1_1/temp4[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_22_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[160] ), 
        .A2(\RI5[1][124] ), .Z(\MC_ARK_ARC_1_1/temp3[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_22_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[28] ), 
        .A2(\RI5[1][4] ), .Z(\MC_ARK_ARC_1_1/temp2[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_22_1  ( .A1(\RI5[1][58] ), .A2(\RI5[1][52] ), .Z(
        \MC_ARK_ARC_1_1/temp1[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_21_5  ( .A1(\RI5[1][96] ), .A2(n88), .Z(
        \MC_ARK_ARC_1_1/temp4[60] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_21_5  ( .A1(\RI5[1][126] ), .A2(\RI5[1][162] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[60] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_21_5  ( .A1(\RI5[1][30] ), .A2(\RI5[1][6] ), .Z(
        \MC_ARK_ARC_1_1/temp2[60] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_21_5  ( .A1(\RI5[1][60] ), .A2(\RI5[1][54] ), .Z(
        \MC_ARK_ARC_1_1/temp1[60] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_21_4  ( .A1(\MC_ARK_ARC_1_1/temp5[61] ), .A2(
        \MC_ARK_ARC_1_1/temp6[61] ), .Z(\MC_ARK_ARC_1_1/buf_output[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_21_4  ( .A1(\MC_ARK_ARC_1_1/temp3[61] ), .A2(
        \MC_ARK_ARC_1_1/temp4[61] ), .Z(\MC_ARK_ARC_1_1/temp6[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_21_4  ( .A1(\MC_ARK_ARC_1_1/temp2[61] ), .A2(
        \MC_ARK_ARC_1_1/temp1[61] ), .Z(\MC_ARK_ARC_1_1/temp5[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_21_4  ( .A1(\RI5[1][97] ), .A2(n465), .Z(
        \MC_ARK_ARC_1_1/temp4[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_21_4  ( .A1(\RI5[1][7] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[31] ), .Z(\MC_ARK_ARC_1_1/temp2[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_21_4  ( .A1(\RI5[1][61] ), .A2(\RI5[1][55] ), .Z(
        \MC_ARK_ARC_1_1/temp1[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_21_3  ( .A1(\RI5[1][98] ), .A2(n57), .Z(
        \MC_ARK_ARC_1_1/temp4[62] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_21_3  ( .A1(\RI5[1][164] ), .A2(\RI5[1][128] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[62] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_21_3  ( .A1(\RI5[1][8] ), .A2(\RI5[1][32] ), .Z(
        \MC_ARK_ARC_1_1/temp2[62] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_21_3  ( .A1(\RI5[1][56] ), .A2(\RI5[1][62] ), .Z(
        \MC_ARK_ARC_1_1/temp1[62] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_21_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[99] ), 
        .A2(n529), .Z(\MC_ARK_ARC_1_1/temp4[63] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_21_2  ( .A1(\RI5[1][129] ), .A2(\RI5[1][165] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[63] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_21_2  ( .A1(n1383), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[9] ), .Z(\MC_ARK_ARC_1_1/temp2[63] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_21_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[63] ), 
        .A2(\RI5[1][57] ), .Z(\MC_ARK_ARC_1_1/temp1[63] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_21_1  ( .A1(\MC_ARK_ARC_1_1/temp5[64] ), .A2(
        \MC_ARK_ARC_1_1/temp6[64] ), .Z(\MC_ARK_ARC_1_1/buf_output[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_21_1  ( .A1(\MC_ARK_ARC_1_1/temp3[64] ), .A2(
        \MC_ARK_ARC_1_1/temp4[64] ), .Z(\MC_ARK_ARC_1_1/temp6[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_21_1  ( .A1(\MC_ARK_ARC_1_1/temp2[64] ), .A2(
        \MC_ARK_ARC_1_1/temp1[64] ), .Z(\MC_ARK_ARC_1_1/temp5[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_21_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[100] ), 
        .A2(n498), .Z(\MC_ARK_ARC_1_1/temp4[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_21_1  ( .A1(\RI5[1][130] ), .A2(\RI5[1][166] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_21_1  ( .A1(\RI5[1][34] ), .A2(\RI5[1][10] ), .Z(
        \MC_ARK_ARC_1_1/temp2[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_21_1  ( .A1(\RI5[1][64] ), .A2(\RI5[1][58] ), .Z(
        \MC_ARK_ARC_1_1/temp1[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_21_0  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[101] ), 
        .A2(n462), .Z(\MC_ARK_ARC_1_1/temp4[65] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_20_5  ( .A1(\RI5[1][102] ), .A2(n560), .Z(
        \MC_ARK_ARC_1_1/temp4[66] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_20_5  ( .A1(\RI5[1][168] ), .A2(\RI5[1][132] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[66] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_20_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[66] ), 
        .A2(\RI5[1][60] ), .Z(\MC_ARK_ARC_1_1/temp1[66] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_20_4  ( .A1(\RI5[1][103] ), .A2(n200), .Z(
        \MC_ARK_ARC_1_1/temp4[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_20_3  ( .A1(\RI5[1][104] ), .A2(n495), .Z(
        \MC_ARK_ARC_1_1/temp4[68] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_20_3  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[170] ), 
        .A2(\RI5[1][134] ), .Z(\MC_ARK_ARC_1_1/temp3[68] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_20_3  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[38] ), 
        .A2(\RI5[1][14] ), .Z(\MC_ARK_ARC_1_1/temp2[68] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_20_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[105] ), 
        .A2(n460), .Z(\MC_ARK_ARC_1_1/temp4[69] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_20_2  ( .A1(\RI5[1][15] ), .A2(\RI5[1][39] ), .Z(
        \MC_ARK_ARC_1_1/temp2[69] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_20_1  ( .A1(\RI5[1][106] ), .A2(n557), .Z(
        \MC_ARK_ARC_1_1/temp4[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_20_0  ( .A1(\RI5[1][107] ), .A2(n212), .Z(
        \MC_ARK_ARC_1_1/temp4[71] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_20_0  ( .A1(\RI5[1][137] ), .A2(\RI5[1][173] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[71] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_20_0  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[41] ), 
        .A2(\RI5[1][17] ), .Z(\MC_ARK_ARC_1_1/temp2[71] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_20_0  ( .A1(\RI5[1][65] ), .A2(\RI5[1][71] ), .Z(
        \MC_ARK_ARC_1_1/temp1[71] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_19_5  ( .A1(\MC_ARK_ARC_1_1/temp6[72] ), .A2(
        \MC_ARK_ARC_1_1/temp5[72] ), .Z(\MC_ARK_ARC_1_1/buf_output[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_19_5  ( .A1(\MC_ARK_ARC_1_1/temp3[72] ), .A2(
        \MC_ARK_ARC_1_1/temp4[72] ), .Z(\MC_ARK_ARC_1_1/temp6[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_19_5  ( .A1(\RI5[1][108] ), .A2(n493), .Z(
        \MC_ARK_ARC_1_1/temp4[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_19_5  ( .A1(\RI5[1][138] ), .A2(\RI5[1][174] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_19_5  ( .A1(\RI5[1][72] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[66] ), .Z(\MC_ARK_ARC_1_1/temp1[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_19_4  ( .A1(\MC_ARK_ARC_1_1/temp3[73] ), .A2(
        \MC_ARK_ARC_1_1/temp4[73] ), .Z(\MC_ARK_ARC_1_1/temp6[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_19_4  ( .A1(\RI5[1][109] ), .A2(n457), .Z(
        \MC_ARK_ARC_1_1/temp4[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_19_4  ( .A1(\RI5[1][175] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[139] ), .Z(\MC_ARK_ARC_1_1/temp3[73] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_19_4  ( .A1(\RI5[1][43] ), .A2(\RI5[1][19] ), .Z(
        \MC_ARK_ARC_1_1/temp2[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_19_4  ( .A1(\RI5[1][73] ), .A2(\RI5[1][67] ), .Z(
        \MC_ARK_ARC_1_1/temp1[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_19_3  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[110] ), 
        .A2(n16), .Z(\MC_ARK_ARC_1_1/temp4[74] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_19_2  ( .A1(\RI5[1][75] ), .A2(\RI5[1][69] ), .Z(
        \MC_ARK_ARC_1_1/temp1[75] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_19_1  ( .A1(\RI5[1][112] ), .A2(n489), .Z(
        \MC_ARK_ARC_1_1/temp4[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_19_1  ( .A1(\RI5[1][142] ), .A2(\RI5[1][178] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_19_1  ( .A1(\RI5[1][46] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[22] ), .Z(\MC_ARK_ARC_1_1/temp2[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_19_0  ( .A1(\RI5[1][23] ), .A2(\RI5[1][47] ), .Z(
        \MC_ARK_ARC_1_1/temp2[77] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_18_5  ( .A1(\RI5[1][114] ), .A2(n230), .Z(
        \MC_ARK_ARC_1_1/temp4[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_18_5  ( .A1(\RI5[1][180] ), .A2(\RI5[1][144] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_18_5  ( .A1(\RI5[1][78] ), .A2(\RI5[1][72] ), .Z(
        \MC_ARK_ARC_1_1/temp1[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_18_4  ( .A1(\RI5[1][115] ), .A2(n240), .Z(
        \MC_ARK_ARC_1_1/temp4[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_18_4  ( .A1(\RI5[1][181] ), .A2(\RI5[1][145] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_18_3  ( .A1(\MC_ARK_ARC_1_1/temp3[80] ), .A2(
        \MC_ARK_ARC_1_1/temp4[80] ), .Z(\MC_ARK_ARC_1_1/temp6[80] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_18_3  ( .A1(\RI5[1][116] ), .A2(n38), .Z(
        \MC_ARK_ARC_1_1/temp4[80] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_18_2  ( .A1(\MC_ARK_ARC_1_1/temp3[81] ), .A2(
        \MC_ARK_ARC_1_1/temp4[81] ), .Z(\MC_ARK_ARC_1_1/temp6[81] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_18_2  ( .A1(\RI5[1][117] ), .A2(n130), .Z(
        \MC_ARK_ARC_1_1/temp4[81] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_18_2  ( .A1(\RI5[1][147] ), .A2(\RI5[1][183] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[81] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_18_2  ( .A1(\RI5[1][27] ), .A2(\RI5[1][51] ), .Z(
        \MC_ARK_ARC_1_1/temp2[81] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_18_2  ( .A1(\RI5[1][81] ), .A2(\RI5[1][75] ), .Z(
        \MC_ARK_ARC_1_1/temp1[81] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_18_1  ( .A1(\MC_ARK_ARC_1_1/temp6[82] ), .A2(
        \MC_ARK_ARC_1_1/temp5[82] ), .Z(\MC_ARK_ARC_1_1/buf_output[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_18_1  ( .A1(\MC_ARK_ARC_1_1/temp3[82] ), .A2(
        \MC_ARK_ARC_1_1/temp4[82] ), .Z(\MC_ARK_ARC_1_1/temp6[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_18_1  ( .A1(\MC_ARK_ARC_1_1/temp2[82] ), .A2(
        \MC_ARK_ARC_1_1/temp1[82] ), .Z(\MC_ARK_ARC_1_1/temp5[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_18_1  ( .A1(\RI5[1][118] ), .A2(n162), .Z(
        \MC_ARK_ARC_1_1/temp4[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_18_1  ( .A1(\RI5[1][184] ), .A2(\RI5[1][148] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_18_1  ( .A1(\RI5[1][52] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[28] ), .Z(\MC_ARK_ARC_1_1/temp2[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_18_1  ( .A1(\RI5[1][76] ), .A2(\RI5[1][82] ), .Z(
        \MC_ARK_ARC_1_1/temp1[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_18_0  ( .A1(\RI5[1][77] ), .A2(\RI5[1][83] ), .Z(
        \MC_ARK_ARC_1_1/temp1[83] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_17_5  ( .A1(\RI5[1][120] ), .A2(n482), .Z(
        \MC_ARK_ARC_1_1/temp4[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_17_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[186] ), 
        .A2(\RI5[1][150] ), .Z(\MC_ARK_ARC_1_1/temp3[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_17_4  ( .A1(\SB2_1_15/buf_output[1] ), .A2(n220), 
        .Z(\MC_ARK_ARC_1_1/temp4[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_17_3  ( .A1(\RI5[1][122] ), .A2(n546), .Z(
        \MC_ARK_ARC_1_1/temp4[86] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_17_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[123] ), 
        .A2(n514), .Z(\MC_ARK_ARC_1_1/temp4[87] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_17_1  ( .A1(\RI5[1][124] ), .A2(n95), .Z(
        \MC_ARK_ARC_1_1/temp4[88] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_17_1  ( .A1(\RI5[1][190] ), .A2(\RI5[1][154] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[88] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_17_1  ( .A1(\RI5[1][82] ), .A2(\RI5[1][88] ), .Z(
        \MC_ARK_ARC_1_1/temp1[88] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_17_0  ( .A1(\RI5[1][125] ), .A2(n108), .Z(
        \MC_ARK_ARC_1_1/temp4[89] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_17_0  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[89] ), 
        .A2(\RI5[1][83] ), .Z(\MC_ARK_ARC_1_1/temp1[89] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_16_5  ( .A1(\RI5[1][126] ), .A2(n185), .Z(
        \MC_ARK_ARC_1_1/temp4[90] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_16_5  ( .A1(\RI5[1][90] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[84] ), .Z(\MC_ARK_ARC_1_1/temp1[90] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_16_4  ( .A1(\RI5[1][127] ), .A2(n511), .Z(
        \MC_ARK_ARC_1_1/temp4[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_16_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[1] ), 
        .A2(\RI5[1][157] ), .Z(\MC_ARK_ARC_1_1/temp3[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_16_3  ( .A1(\RI5[1][128] ), .A2(n476), .Z(
        \MC_ARK_ARC_1_1/temp4[92] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_16_2  ( .A1(\RI5[1][129] ), .A2(n443), .Z(
        \MC_ARK_ARC_1_1/temp4[93] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_16_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[63] ), 
        .A2(\RI5[1][39] ), .Z(\MC_ARK_ARC_1_1/temp2[93] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_16_2  ( .A1(\RI5[1][87] ), .A2(\RI5[1][93] ), .Z(
        \MC_ARK_ARC_1_1/temp1[93] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_16_1  ( .A1(\MC_ARK_ARC_1_1/temp6[94] ), .A2(
        \MC_ARK_ARC_1_1/temp5[94] ), .Z(\MC_ARK_ARC_1_1/buf_output[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_16_1  ( .A1(\MC_ARK_ARC_1_1/temp3[94] ), .A2(
        \MC_ARK_ARC_1_1/temp4[94] ), .Z(\MC_ARK_ARC_1_1/temp6[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_16_1  ( .A1(\MC_ARK_ARC_1_1/temp2[94] ), .A2(
        \MC_ARK_ARC_1_1/temp1[94] ), .Z(\MC_ARK_ARC_1_1/temp5[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_16_1  ( .A1(\RI5[1][130] ), .A2(n166), .Z(
        \MC_ARK_ARC_1_1/temp4[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_16_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[160] ), 
        .A2(\RI5[1][4] ), .Z(\MC_ARK_ARC_1_1/temp3[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_16_1  ( .A1(\RI5[1][94] ), .A2(\RI5[1][88] ), .Z(
        \MC_ARK_ARC_1_1/temp1[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_16_0  ( .A1(\MC_ARK_ARC_1_1/temp3[95] ), .A2(
        \MC_ARK_ARC_1_1/temp4[95] ), .Z(\MC_ARK_ARC_1_1/temp6[95] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_16_0  ( .A1(\RI5[1][131] ), .A2(n186), .Z(
        \MC_ARK_ARC_1_1/temp4[95] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_16_0  ( .A1(\RI5[1][65] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[41] ), .Z(\MC_ARK_ARC_1_1/temp2[95] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_15_5  ( .A1(\RI5[1][132] ), .A2(n66), .Z(
        \MC_ARK_ARC_1_1/temp4[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_15_5  ( .A1(\RI5[1][6] ), .A2(\RI5[1][162] ), .Z(
        \MC_ARK_ARC_1_1/temp3[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_15_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[42] ), 
        .A2(\MC_ARK_ARC_1_1/buf_datainput[66] ), .Z(\MC_ARK_ARC_1_1/temp2[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_15_5  ( .A1(\RI5[1][90] ), .A2(\RI5[1][96] ), .Z(
        \MC_ARK_ARC_1_1/temp1[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_15_4  ( .A1(\RI5[1][133] ), .A2(n441), .Z(
        \MC_ARK_ARC_1_1/temp4[97] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_15_4  ( .A1(\RI5[1][67] ), .A2(\RI5[1][43] ), .Z(
        \MC_ARK_ARC_1_1/temp2[97] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_15_3  ( .A1(\RI5[1][134] ), .A2(n540), .Z(
        \MC_ARK_ARC_1_1/temp4[98] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_15_2  ( .A1(\SB2_1_11/buf_output[3] ), .A2(n181), 
        .Z(\MC_ARK_ARC_1_1/temp4[99] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_15_1  ( .A1(\RI5[1][136] ), .A2(n127), .Z(
        \MC_ARK_ARC_1_1/temp4[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_15_1  ( .A1(\RI5[1][70] ), .A2(\RI5[1][46] ), .Z(
        \MC_ARK_ARC_1_1/temp2[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_15_0  ( .A1(\RI5[1][137] ), .A2(n438), .Z(
        \MC_ARK_ARC_1_1/temp4[101] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_14_5  ( .A1(\MC_ARK_ARC_1_1/temp6[102] ), .A2(
        \MC_ARK_ARC_1_1/temp5[102] ), .Z(\MC_ARK_ARC_1_1/buf_output[102] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_14_5  ( .A1(\MC_ARK_ARC_1_1/temp4[102] ), .A2(
        \MC_ARK_ARC_1_1/temp3[102] ), .Z(\MC_ARK_ARC_1_1/temp6[102] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_14_5  ( .A1(\MC_ARK_ARC_1_1/temp1[102] ), .A2(
        \MC_ARK_ARC_1_1/temp2[102] ), .Z(\MC_ARK_ARC_1_1/temp5[102] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_14_5  ( .A1(\RI5[1][138] ), .A2(n139), .Z(
        \MC_ARK_ARC_1_1/temp4[102] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_14_5  ( .A1(\RI5[1][12] ), .A2(\RI5[1][168] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[102] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_14_5  ( .A1(\RI5[1][48] ), .A2(\RI5[1][72] ), .Z(
        \MC_ARK_ARC_1_1/temp2[102] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_14_5  ( .A1(\RI5[1][96] ), .A2(\RI5[1][102] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[102] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_14_4  ( .A1(\MC_ARK_ARC_1_1/temp4[103] ), .A2(
        \MC_ARK_ARC_1_1/temp3[103] ), .Z(\MC_ARK_ARC_1_1/temp6[103] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_14_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[139] ), 
        .A2(n502), .Z(\MC_ARK_ARC_1_1/temp4[103] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_14_4  ( .A1(\RI5[1][13] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[169] ), .Z(\MC_ARK_ARC_1_1/temp3[103] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_14_4  ( .A1(\RI5[1][73] ), .A2(\RI5[1][49] ), .Z(
        \MC_ARK_ARC_1_1/temp2[103] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_14_4  ( .A1(\RI5[1][103] ), .A2(\RI5[1][97] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[103] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_14_3  ( .A1(\MC_ARK_ARC_1_1/temp5[104] ), .A2(
        \MC_ARK_ARC_1_1/temp6[104] ), .Z(\MC_ARK_ARC_1_1/buf_output[104] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_14_3  ( .A1(\MC_ARK_ARC_1_1/temp3[104] ), .A2(
        \MC_ARK_ARC_1_1/temp4[104] ), .Z(\MC_ARK_ARC_1_1/temp6[104] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_14_3  ( .A1(\MC_ARK_ARC_1_1/temp2[104] ), .A2(
        \MC_ARK_ARC_1_1/temp1[104] ), .Z(\MC_ARK_ARC_1_1/temp5[104] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_14_3  ( .A1(\RI5[1][140] ), .A2(n468), .Z(
        \MC_ARK_ARC_1_1/temp4[104] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_14_3  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[74] ), 
        .A2(\RI5[1][50] ), .Z(\MC_ARK_ARC_1_1/temp2[104] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_14_2  ( .A1(\RI5[1][141] ), .A2(n39), .Z(
        \MC_ARK_ARC_1_1/temp4[105] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_14_1  ( .A1(\MC_ARK_ARC_1_1/temp3[106] ), .A2(
        \MC_ARK_ARC_1_1/temp4[106] ), .Z(\MC_ARK_ARC_1_1/temp6[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_14_1  ( .A1(\RI5[1][142] ), .A2(n68), .Z(
        \MC_ARK_ARC_1_1/temp4[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_14_1  ( .A1(\RI5[1][76] ), .A2(\RI5[1][52] ), .Z(
        \MC_ARK_ARC_1_1/temp2[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_14_1  ( .A1(\RI5[1][106] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[100] ), .Z(\MC_ARK_ARC_1_1/temp1[106] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_14_0  ( .A1(\MC_ARK_ARC_1_1/temp5[107] ), .A2(
        \MC_ARK_ARC_1_1/temp6[107] ), .Z(\MC_ARK_ARC_1_1/buf_output[107] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_13_5  ( .A1(\MC_ARK_ARC_1_1/temp3[108] ), .A2(
        \MC_ARK_ARC_1_1/temp4[108] ), .Z(\MC_ARK_ARC_1_1/temp6[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_13_5  ( .A1(\RI5[1][144] ), .A2(n135), .Z(
        \MC_ARK_ARC_1_1/temp4[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_13_5  ( .A1(\RI5[1][78] ), .A2(\RI5[1][54] ), .Z(
        \MC_ARK_ARC_1_1/temp2[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_13_4  ( .A1(\MC_ARK_ARC_1_1/temp3[109] ), .A2(
        \MC_ARK_ARC_1_1/temp4[109] ), .Z(\MC_ARK_ARC_1_1/temp6[109] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_13_4  ( .A1(\RI5[1][145] ), .A2(n562), .Z(
        \MC_ARK_ARC_1_1/temp4[109] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_13_4  ( .A1(\RI5[1][79] ), .A2(\RI5[1][55] ), .Z(
        \MC_ARK_ARC_1_1/temp2[109] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_13_4  ( .A1(\RI5[1][109] ), .A2(\RI5[1][103] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[109] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_13_3  ( .A1(\RI5[1][20] ), .A2(\RI5[1][176] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[110] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_13_2  ( .A1(\RI5[1][21] ), .A2(\RI5[1][177] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[111] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_13_1  ( .A1(\RI5[1][148] ), .A2(n103), .Z(
        \MC_ARK_ARC_1_1/temp4[112] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_13_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[22] ), 
        .A2(\RI5[1][178] ), .Z(\MC_ARK_ARC_1_1/temp3[112] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_13_1  ( .A1(\RI5[1][112] ), .A2(\RI5[1][106] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[112] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_13_0  ( .A1(\RI5[1][149] ), .A2(n196), .Z(
        \MC_ARK_ARC_1_1/temp4[113] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_12_5  ( .A1(\RI5[1][150] ), .A2(n217), .Z(
        \MC_ARK_ARC_1_1/temp4[114] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_12_5  ( .A1(\RI5[1][24] ), .A2(\RI5[1][180] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[114] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_12_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[84] ), 
        .A2(\RI5[1][60] ), .Z(\MC_ARK_ARC_1_1/temp2[114] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_12_5  ( .A1(\RI5[1][114] ), .A2(\RI5[1][108] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[114] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_12_4  ( .A1(\RI5[1][181] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[25] ), .Z(\MC_ARK_ARC_1_1/temp3[115] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_12_3  ( .A1(\RI5[1][86] ), .A2(\RI5[1][62] ), .Z(
        \MC_ARK_ARC_1_1/temp2[116] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_12_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[153] ), 
        .A2(n558), .Z(\MC_ARK_ARC_1_1/temp4[117] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_12_1  ( .A1(\MC_ARK_ARC_1_1/temp4[118] ), .A2(
        \MC_ARK_ARC_1_1/temp3[118] ), .Z(\MC_ARK_ARC_1_1/temp6[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_12_1  ( .A1(\MC_ARK_ARC_1_1/temp2[118] ), .A2(
        \MC_ARK_ARC_1_1/temp1[118] ), .Z(\MC_ARK_ARC_1_1/temp5[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_12_1  ( .A1(\RI5[1][154] ), .A2(n207), .Z(
        \MC_ARK_ARC_1_1/temp4[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_12_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[28] ), 
        .A2(\RI5[1][184] ), .Z(\MC_ARK_ARC_1_1/temp3[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_12_1  ( .A1(\RI5[1][88] ), .A2(\RI5[1][64] ), .Z(
        \MC_ARK_ARC_1_1/temp2[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_12_1  ( .A1(\RI5[1][112] ), .A2(\RI5[1][118] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_12_0  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[155] ), 
        .A2(n204), .Z(\MC_ARK_ARC_1_1/temp4[119] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_11_5  ( .A1(\RI5[1][156] ), .A2(n458), .Z(
        \MC_ARK_ARC_1_1/temp4[120] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_11_5  ( .A1(\RI5[1][30] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[186] ), .Z(\MC_ARK_ARC_1_1/temp3[120] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_11_5  ( .A1(\RI5[1][90] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[66] ), .Z(\MC_ARK_ARC_1_1/temp2[120] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_11_5  ( .A1(\RI5[1][120] ), .A2(\RI5[1][114] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[120] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_11_4  ( .A1(\RI5[1][157] ), .A2(n232), .Z(
        \MC_ARK_ARC_1_1/temp4[121] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_11_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[31] ), 
        .A2(\MC_ARK_ARC_1_1/buf_datainput[187] ), .Z(
        \MC_ARK_ARC_1_1/temp3[121] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_11_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[159] ), 
        .A2(n81), .Z(\MC_ARK_ARC_1_1/temp4[123] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_11_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[123] ), 
        .A2(\RI5[1][117] ), .Z(\MC_ARK_ARC_1_1/temp1[123] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_11_1  ( .A1(\MC_ARK_ARC_1_1/temp6[124] ), .A2(
        \MC_ARK_ARC_1_1/temp5[124] ), .Z(\MC_ARK_ARC_1_1/buf_output[124] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_11_1  ( .A1(\MC_ARK_ARC_1_1/temp3[124] ), .A2(
        \MC_ARK_ARC_1_1/temp4[124] ), .Z(\MC_ARK_ARC_1_1/temp6[124] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_11_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[160] ), 
        .A2(n195), .Z(\MC_ARK_ARC_1_1/temp4[124] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_11_1  ( .A1(\RI5[1][34] ), .A2(\RI5[1][190] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[124] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_11_0  ( .A1(\RI5[1][161] ), .A2(n86), .Z(
        \MC_ARK_ARC_1_1/temp4[125] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_11_0  ( .A1(\RI5[1][119] ), .A2(\RI5[1][125] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[125] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_10_5  ( .A1(\RI5[1][162] ), .A2(n116), .Z(
        \MC_ARK_ARC_1_1/temp4[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_10_5  ( .A1(\RI5[1][72] ), .A2(\RI5[1][96] ), .Z(
        \MC_ARK_ARC_1_1/temp2[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_10_5  ( .A1(\RI5[1][126] ), .A2(\RI5[1][120] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_10_4  ( .A1(\MC_ARK_ARC_1_1/temp6[127] ), .A2(
        \MC_ARK_ARC_1_1/temp5[127] ), .Z(\MC_ARK_ARC_1_1/buf_output[127] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_10_4  ( .A1(\MC_ARK_ARC_1_1/temp3[127] ), .A2(
        \MC_ARK_ARC_1_1/temp4[127] ), .Z(\MC_ARK_ARC_1_1/temp6[127] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_10_4  ( .A1(\MC_ARK_ARC_1_1/temp1[127] ), .A2(
        \MC_ARK_ARC_1_1/temp2[127] ), .Z(\MC_ARK_ARC_1_1/temp5[127] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_10_4  ( .A1(\RI5[1][37] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[1] ), .Z(\MC_ARK_ARC_1_1/temp3[127] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_10_4  ( .A1(\RI5[1][73] ), .A2(\RI5[1][97] ), .Z(
        \MC_ARK_ARC_1_1/temp2[127] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_10_4  ( .A1(\RI5[1][121] ), .A2(\RI5[1][127] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[127] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_10_3  ( .A1(\RI5[1][164] ), .A2(n23), .Z(
        \MC_ARK_ARC_1_1/temp4[128] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_10_2  ( .A1(\RI5[1][165] ), .A2(n115), .Z(
        \MC_ARK_ARC_1_1/temp4[129] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_10_1  ( .A1(\RI5[1][166] ), .A2(n146), .Z(
        \MC_ARK_ARC_1_1/temp4[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_10_1  ( .A1(\RI5[1][76] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[100] ), .Z(\MC_ARK_ARC_1_1/temp2[130] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_10_0  ( .A1(\RI5[1][167] ), .A2(n483), .Z(
        \MC_ARK_ARC_1_1/temp4[131] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_9_5  ( .A1(\RI5[1][168] ), .A2(n165), .Z(
        \MC_ARK_ARC_1_1/temp4[132] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_9_5  ( .A1(\RI5[1][6] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[42] ), .Z(\MC_ARK_ARC_1_1/temp3[132] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_9_4  ( .A1(\MC_ARK_ARC_1_1/temp1[133] ), .A2(
        \MC_ARK_ARC_1_1/temp2[133] ), .Z(\MC_ARK_ARC_1_1/temp5[133] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_9_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[169] ), 
        .A2(n184), .Z(\MC_ARK_ARC_1_1/temp4[133] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_9_4  ( .A1(\RI5[1][7] ), .A2(\RI5[1][43] ), .Z(
        \MC_ARK_ARC_1_1/temp3[133] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_9_3  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[170] ), 
        .A2(n83), .Z(\MC_ARK_ARC_1_1/temp4[134] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_9_3  ( .A1(\RI5[1][44] ), .A2(\RI5[1][8] ), .Z(
        \MC_ARK_ARC_1_1/temp3[134] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_9_1  ( .A1(\RI5[1][172] ), .A2(n52), .Z(
        \MC_ARK_ARC_1_1/temp4[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_9_1  ( .A1(\RI5[1][10] ), .A2(\RI5[1][46] ), .Z(
        \MC_ARK_ARC_1_1/temp3[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_9_1  ( .A1(\RI5[1][82] ), .A2(\RI5[1][106] ), .Z(
        \MC_ARK_ARC_1_1/temp2[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_9_0  ( .A1(\MC_ARK_ARC_1_1/temp4[137] ), .A2(
        \MC_ARK_ARC_1_1/temp3[137] ), .Z(\MC_ARK_ARC_1_1/temp6[137] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_9_0  ( .A1(\RI5[1][173] ), .A2(n194), .Z(
        \MC_ARK_ARC_1_1/temp4[137] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_9_0  ( .A1(\RI5[1][11] ), .A2(\RI5[1][47] ), .Z(
        \MC_ARK_ARC_1_1/temp3[137] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_8_5  ( .A1(\MC_ARK_ARC_1_1/temp1[138] ), .A2(
        \MC_ARK_ARC_1_1/temp2[138] ), .Z(\MC_ARK_ARC_1_1/temp5[138] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_8_5  ( .A1(\RI5[1][174] ), .A2(n512), .Z(
        \MC_ARK_ARC_1_1/temp4[138] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_8_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[84] ), 
        .A2(\RI5[1][108] ), .Z(\MC_ARK_ARC_1_1/temp2[138] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_8_5  ( .A1(\RI5[1][138] ), .A2(\RI5[1][132] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[138] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_8_4  ( .A1(\RI5[1][175] ), .A2(n477), .Z(
        \MC_ARK_ARC_1_1/temp4[139] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_8_4  ( .A1(\RI5[1][85] ), .A2(\RI5[1][109] ), .Z(
        \MC_ARK_ARC_1_1/temp2[139] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_8_4  ( .A1(\RI5[1][133] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[139] ), .Z(\MC_ARK_ARC_1_1/temp1[139] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_8_3  ( .A1(\MC_ARK_ARC_1_1/temp3[140] ), .A2(
        \MC_ARK_ARC_1_1/temp4[140] ), .Z(\MC_ARK_ARC_1_1/temp6[140] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_8_3  ( .A1(\RI5[1][176] ), .A2(n67), .Z(
        \MC_ARK_ARC_1_1/temp4[140] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_8_2  ( .A1(\RI5[1][177] ), .A2(n543), .Z(
        \MC_ARK_ARC_1_1/temp4[141] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_8_1  ( .A1(\MC_ARK_ARC_1_1/temp3[142] ), .A2(
        \MC_ARK_ARC_1_1/temp4[142] ), .Z(\MC_ARK_ARC_1_1/temp6[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_8_1  ( .A1(\RI5[1][178] ), .A2(n509), .Z(
        \MC_ARK_ARC_1_1/temp4[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_8_1  ( .A1(\RI5[1][112] ), .A2(\RI5[1][88] ), .Z(
        \MC_ARK_ARC_1_1/temp2[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_8_0  ( .A1(\MC_ARK_ARC_1_1/temp5[143] ), .A2(
        \MC_ARK_ARC_1_1/temp6[143] ), .Z(\MC_ARK_ARC_1_1/buf_output[143] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_7_5  ( .A1(\MC_ARK_ARC_1_1/temp5[144] ), .A2(
        \MC_ARK_ARC_1_1/temp6[144] ), .Z(\MC_ARK_ARC_1_1/buf_output[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_7_5  ( .A1(\MC_ARK_ARC_1_1/temp3[144] ), .A2(
        \MC_ARK_ARC_1_1/temp4[144] ), .Z(\MC_ARK_ARC_1_1/temp6[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_7_5  ( .A1(\RI5[1][180] ), .A2(n137), .Z(
        \MC_ARK_ARC_1_1/temp4[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_7_5  ( .A1(\RI5[1][54] ), .A2(\RI5[1][18] ), .Z(
        \MC_ARK_ARC_1_1/temp3[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_7_5  ( .A1(\RI5[1][138] ), .A2(\RI5[1][144] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_7_4  ( .A1(\RI5[1][181] ), .A2(n541), .Z(
        \MC_ARK_ARC_1_1/temp4[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_7_3  ( .A1(\RI5[1][182] ), .A2(n506), .Z(
        \MC_ARK_ARC_1_1/temp4[146] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_7_3  ( .A1(\RI5[1][146] ), .A2(\RI5[1][140] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[146] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_7_2  ( .A1(\SB2_1_3/buf_output[3] ), .A2(n471), 
        .Z(\MC_ARK_ARC_1_1/temp4[147] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_7_2  ( .A1(\RI5[1][21] ), .A2(\RI5[1][57] ), .Z(
        \MC_ARK_ARC_1_1/temp3[147] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_7_2  ( .A1(\RI5[1][93] ), .A2(\RI5[1][117] ), .Z(
        \MC_ARK_ARC_1_1/temp2[147] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_7_2  ( .A1(\SB2_1_10/buf_output[3] ), .A2(n5521), 
        .Z(\MC_ARK_ARC_1_1/temp1[147] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_7_1  ( .A1(\MC_ARK_ARC_1_1/temp3[148] ), .A2(
        \MC_ARK_ARC_1_1/temp4[148] ), .Z(\MC_ARK_ARC_1_1/temp6[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_7_1  ( .A1(\RI5[1][184] ), .A2(n223), .Z(
        \MC_ARK_ARC_1_1/temp4[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_7_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[22] ), 
        .A2(\RI5[1][58] ), .Z(\MC_ARK_ARC_1_1/temp3[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_7_1  ( .A1(\RI5[1][118] ), .A2(\RI5[1][94] ), .Z(
        \MC_ARK_ARC_1_1/temp2[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_7_1  ( .A1(\RI5[1][142] ), .A2(\RI5[1][148] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_7_0  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[185] ), 
        .A2(n153), .Z(\MC_ARK_ARC_1_1/temp4[149] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_7_0  ( .A1(\RI5[1][119] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[95] ), .Z(\MC_ARK_ARC_1_1/temp2[149] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_7_0  ( .A1(\RI5[1][149] ), .A2(\RI5[1][143] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[149] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_6_5  ( .A1(\MC_ARK_ARC_1_1/temp3[150] ), .A2(
        \MC_ARK_ARC_1_1/temp4[150] ), .Z(\MC_ARK_ARC_1_1/temp6[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_6_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[186] ), 
        .A2(n503), .Z(\MC_ARK_ARC_1_1/temp4[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_6_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[187] ), 
        .A2(n160), .Z(\MC_ARK_ARC_1_1/temp4[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_6_4  ( .A1(\RI5[1][61] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[25] ), .Z(\MC_ARK_ARC_1_1/temp3[151] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_6_4  ( .A1(\RI5[1][145] ), .A2(\RI5[1][151] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_6_2  ( .A1(\MC_ARK_ARC_1_1/temp1[153] ), .A2(
        \MC_ARK_ARC_1_1/temp2[153] ), .Z(\MC_ARK_ARC_1_1/temp5[153] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_6_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[99] ), 
        .A2(\MC_ARK_ARC_1_1/buf_datainput[123] ), .Z(
        \MC_ARK_ARC_1_1/temp2[153] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_6_1  ( .A1(\RI5[1][190] ), .A2(n501), .Z(
        \MC_ARK_ARC_1_1/temp4[154] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_6_0  ( .A1(\MC_ARK_ARC_1_1/temp3[155] ), .A2(
        \MC_ARK_ARC_1_1/temp4[155] ), .Z(\MC_ARK_ARC_1_1/temp6[155] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_6_0  ( .A1(\RI5[1][191] ), .A2(n44), .Z(
        \MC_ARK_ARC_1_1/temp4[155] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_6_0  ( .A1(\RI5[1][65] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[29] ), .Z(\MC_ARK_ARC_1_1/temp3[155] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_6_0  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[101] ), 
        .A2(\RI5[1][125] ), .Z(\MC_ARK_ARC_1_1/temp2[155] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_5_5  ( .A1(\MC_ARK_ARC_1_1/temp5[156] ), .A2(
        \MC_ARK_ARC_1_1/temp6[156] ), .Z(\MC_ARK_ARC_1_1/buf_output[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_5_5  ( .A1(\MC_ARK_ARC_1_1/temp3[156] ), .A2(
        \MC_ARK_ARC_1_1/temp4[156] ), .Z(\MC_ARK_ARC_1_1/temp6[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_5_5  ( .A1(\RI5[1][0] ), .A2(n65), .Z(
        \MC_ARK_ARC_1_1/temp4[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_5_5  ( .A1(\RI5[1][30] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[66] ), .Z(\MC_ARK_ARC_1_1/temp3[156] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_5_5  ( .A1(\RI5[1][126] ), .A2(\RI5[1][102] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_5_5  ( .A1(\RI5[1][156] ), .A2(\RI5[1][150] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_5_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[1] ), 
        .A2(n531), .Z(\MC_ARK_ARC_1_1/temp4[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_5_3  ( .A1(\MC_ARK_ARC_1_1/temp5[158] ), .A2(
        \MC_ARK_ARC_1_1/temp6[158] ), .Z(\MC_ARK_ARC_1_1/buf_output[158] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_5_3  ( .A1(\RI5[1][2] ), .A2(n499), .Z(
        \MC_ARK_ARC_1_1/temp4[158] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_5_3  ( .A1(\RI5[1][68] ), .A2(\RI5[1][32] ), .Z(
        \MC_ARK_ARC_1_1/temp3[158] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_5_3  ( .A1(\RI5[1][128] ), .A2(\RI5[1][104] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[158] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_5_3  ( .A1(\RI5[1][152] ), .A2(\RI5[1][158] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[158] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_5_2  ( .A1(\MC_ARK_ARC_1_1/temp2[159] ), .A2(
        \MC_ARK_ARC_1_1/temp1[159] ), .Z(\MC_ARK_ARC_1_1/temp5[159] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_5_2  ( .A1(\RI5[1][3] ), .A2(n464), .Z(
        \MC_ARK_ARC_1_1/temp4[159] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_5_1  ( .A1(\MC_ARK_ARC_1_1/temp3[160] ), .A2(
        \MC_ARK_ARC_1_1/temp4[160] ), .Z(\MC_ARK_ARC_1_1/temp6[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_5_1  ( .A1(\MC_ARK_ARC_1_1/temp1[160] ), .A2(
        \MC_ARK_ARC_1_1/temp2[160] ), .Z(\MC_ARK_ARC_1_1/temp5[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_5_1  ( .A1(\RI5[1][4] ), .A2(n214), .Z(
        \MC_ARK_ARC_1_1/temp4[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_5_1  ( .A1(\RI5[1][70] ), .A2(\RI5[1][34] ), .Z(
        \MC_ARK_ARC_1_1/temp3[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_5_1  ( .A1(\RI5[1][106] ), .A2(\RI5[1][130] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_5_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[160] ), 
        .A2(\RI5[1][154] ), .Z(\MC_ARK_ARC_1_1/temp1[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_5_0  ( .A1(\RI5[1][5] ), .A2(n122), .Z(
        \MC_ARK_ARC_1_1/temp4[161] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_5_0  ( .A1(\RI5[1][107] ), .A2(\RI5[1][131] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[161] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_4_5  ( .A1(\RI5[1][6] ), .A2(n188), .Z(
        \MC_ARK_ARC_1_1/temp4[162] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_4_5  ( .A1(\RI5[1][36] ), .A2(\RI5[1][72] ), .Z(
        \MC_ARK_ARC_1_1/temp3[162] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_4_4  ( .A1(\SB2_1_2/buf_output[1] ), .A2(n461), 
        .Z(\MC_ARK_ARC_1_1/temp4[163] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_4_4  ( .A1(\RI5[1][133] ), .A2(\RI5[1][109] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[163] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_4_3  ( .A1(\RI5[1][8] ), .A2(n171), .Z(
        \MC_ARK_ARC_1_1/temp4[164] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_4_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[9] ), 
        .A2(n90), .Z(\MC_ARK_ARC_1_1/temp4[165] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_4_2  ( .A1(\RI5[1][75] ), .A2(\RI5[1][39] ), .Z(
        \MC_ARK_ARC_1_1/temp3[165] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_4_2  ( .A1(\RI5[1][111] ), .A2(\RI5[1][135] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[165] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_4_1  ( .A1(\MC_ARK_ARC_1_1/temp3[166] ), .A2(
        \MC_ARK_ARC_1_1/temp4[166] ), .Z(\MC_ARK_ARC_1_1/temp6[166] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_4_1  ( .A1(\RI5[1][10] ), .A2(n205), .Z(
        \MC_ARK_ARC_1_1/temp4[166] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_4_1  ( .A1(\RI5[1][76] ), .A2(\RI5[1][40] ), .Z(
        \MC_ARK_ARC_1_1/temp3[166] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_3_5  ( .A1(\RI5[1][12] ), .A2(n228), .Z(
        \MC_ARK_ARC_1_1/temp4[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_3_5  ( .A1(\RI5[1][138] ), .A2(\RI5[1][114] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_3_5  ( .A1(\RI5[1][168] ), .A2(\RI5[1][162] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_3_4  ( .A1(\RI5[1][13] ), .A2(n522), .Z(
        \MC_ARK_ARC_1_1/temp4[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_3_3  ( .A1(\RI5[1][14] ), .A2(n45), .Z(
        \MC_ARK_ARC_1_1/temp4[170] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_3_1  ( .A1(\MC_ARK_ARC_1_1/temp5[172] ), .A2(
        \MC_ARK_ARC_1_1/temp6[172] ), .Z(\MC_ARK_ARC_1_1/buf_output[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_3_1  ( .A1(\MC_ARK_ARC_1_1/temp4[172] ), .A2(
        \MC_ARK_ARC_1_1/temp3[172] ), .Z(\MC_ARK_ARC_1_1/temp6[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_3_1  ( .A1(\RI5[1][16] ), .A2(n554), .Z(
        \MC_ARK_ARC_1_1/temp4[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_3_1  ( .A1(\RI5[1][82] ), .A2(\RI5[1][46] ), .Z(
        \MC_ARK_ARC_1_1/temp3[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_3_1  ( .A1(\RI5[1][142] ), .A2(\RI5[1][118] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_3_0  ( .A1(\MC_ARK_ARC_1_1/temp2[173] ), .A2(
        \MC_ARK_ARC_1_1/temp1[173] ), .Z(\MC_ARK_ARC_1_1/temp5[173] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_3_0  ( .A1(\RI5[1][17] ), .A2(n520), .Z(
        \MC_ARK_ARC_1_1/temp4[173] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_3_0  ( .A1(\RI5[1][143] ), .A2(\RI5[1][119] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[173] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_3_0  ( .A1(\RI5[1][167] ), .A2(\RI5[1][173] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[173] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_2_5  ( .A1(\RI5[1][18] ), .A2(n487), .Z(
        \MC_ARK_ARC_1_1/temp4[174] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_2_5  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[84] ), 
        .A2(\RI5[1][48] ), .Z(\MC_ARK_ARC_1_1/temp3[174] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_2_5  ( .A1(\RI5[1][174] ), .A2(\RI5[1][168] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[174] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_2_4  ( .A1(\MC_ARK_ARC_1_1/temp2[175] ), .A2(
        \MC_ARK_ARC_1_1/temp1[175] ), .Z(\MC_ARK_ARC_1_1/temp5[175] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_2_4  ( .A1(\RI5[1][19] ), .A2(n451), .Z(
        \MC_ARK_ARC_1_1/temp4[175] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_2_4  ( .A1(\RI5[1][85] ), .A2(\RI5[1][49] ), .Z(
        \MC_ARK_ARC_1_1/temp3[175] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_2_4  ( .A1(\RI5[1][121] ), .A2(\RI5[1][145] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[175] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_2_4  ( .A1(\RI5[1][175] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[169] ), .Z(\MC_ARK_ARC_1_1/temp1[175] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_2_3  ( .A1(\MC_ARK_ARC_1_1/temp3[176] ), .A2(
        \MC_ARK_ARC_1_1/temp4[176] ), .Z(\MC_ARK_ARC_1_1/temp6[176] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_2_3  ( .A1(\RI5[1][20] ), .A2(n173), .Z(
        \MC_ARK_ARC_1_1/temp4[176] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_2_2  ( .A1(\RI5[1][21] ), .A2(n517), .Z(
        \MC_ARK_ARC_1_1/temp4[177] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_2_1  ( .A1(\MC_ARK_ARC_1_1/temp3[178] ), .A2(
        \MC_ARK_ARC_1_1/temp4[178] ), .Z(\MC_ARK_ARC_1_1/temp6[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_2_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[22] ), 
        .A2(n484), .Z(\MC_ARK_ARC_1_1/temp4[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_2_1  ( .A1(\RI5[1][52] ), .A2(\RI5[1][88] ), .Z(
        \MC_ARK_ARC_1_1/temp3[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_2_1  ( .A1(\RI5[1][148] ), .A2(\RI5[1][124] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_2_1  ( .A1(\RI5[1][178] ), .A2(\RI5[1][172] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_2_0  ( .A1(\RI5[1][23] ), .A2(n449), .Z(
        \MC_ARK_ARC_1_1/temp4[179] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_2_0  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[89] ), 
        .A2(\RI5[1][53] ), .Z(\MC_ARK_ARC_1_1/temp3[179] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_2_0  ( .A1(\RI5[1][125] ), .A2(\RI5[1][149] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[179] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_2_0  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[179] ), 
        .A2(\RI5[1][173] ), .Z(\MC_ARK_ARC_1_1/temp1[179] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_1_5  ( .A1(\MC_ARK_ARC_1_1/temp3[180] ), .A2(
        \MC_ARK_ARC_1_1/temp4[180] ), .Z(\MC_ARK_ARC_1_1/temp6[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_1_5  ( .A1(\RI5[1][24] ), .A2(n235), .Z(
        \MC_ARK_ARC_1_1/temp4[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_1_5  ( .A1(\RI5[1][90] ), .A2(\RI5[1][54] ), .Z(
        \MC_ARK_ARC_1_1/temp3[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_1_5  ( .A1(\RI5[1][126] ), .A2(\RI5[1][150] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_1_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[25] ), 
        .A2(n516), .Z(\MC_ARK_ARC_1_1/temp4[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X7_1_2  ( .A1(\MC_ARK_ARC_1_1/temp5[183] ), .A2(
        \MC_ARK_ARC_1_1/temp6[183] ), .Z(\MC_ARK_ARC_1_1/buf_output[183] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_1_2  ( .A1(\MC_ARK_ARC_1_1/temp3[183] ), .A2(
        \MC_ARK_ARC_1_1/temp4[183] ), .Z(\MC_ARK_ARC_1_1/temp6[183] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_1_2  ( .A1(\RI5[1][27] ), .A2(n9), .Z(
        \MC_ARK_ARC_1_1/temp4[183] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_1_2  ( .A1(\RI5[1][57] ), .A2(\RI5[1][93] ), .Z(
        \MC_ARK_ARC_1_1/temp3[183] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X5_1_1  ( .A1(\MC_ARK_ARC_1_1/temp2[184] ), .A2(
        \MC_ARK_ARC_1_1/temp1[184] ), .Z(\MC_ARK_ARC_1_1/temp5[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_1_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[28] ), 
        .A2(n227), .Z(\MC_ARK_ARC_1_1/temp4[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_1_1  ( .A1(\RI5[1][94] ), .A2(\RI5[1][58] ), .Z(
        \MC_ARK_ARC_1_1/temp3[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_1_1  ( .A1(\RI5[1][130] ), .A2(\RI5[1][154] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_1_1  ( .A1(\RI5[1][178] ), .A2(\RI5[1][184] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_1_0  ( .A1(\MC_ARK_ARC_1_1/temp3[185] ), .A2(
        \MC_ARK_ARC_1_1/temp4[185] ), .Z(\MC_ARK_ARC_1_1/temp6[185] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_1_0  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[29] ), 
        .A2(n180), .Z(\MC_ARK_ARC_1_1/temp4[185] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_0_5  ( .A1(\RI5[1][30] ), .A2(n202), .Z(
        \MC_ARK_ARC_1_1/temp4[186] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_0_5  ( .A1(\RI5[1][60] ), .A2(\RI5[1][96] ), .Z(
        \MC_ARK_ARC_1_1/temp3[186] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_0_5  ( .A1(\RI5[1][132] ), .A2(\RI5[1][156] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[186] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_0_5  ( .A1(\RI5[1][180] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[186] ), .Z(\MC_ARK_ARC_1_1/temp1[186] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_0_4  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[31] ), 
        .A2(n12), .Z(\MC_ARK_ARC_1_1/temp4[187] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_0_3  ( .A1(\RI5[1][32] ), .A2(n3), .Z(
        \MC_ARK_ARC_1_1/temp4[188] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_0_3  ( .A1(\RI5[1][134] ), .A2(\RI5[1][158] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[188] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X6_0_2  ( .A1(\MC_ARK_ARC_1_1/temp3[189] ), .A2(
        \MC_ARK_ARC_1_1/temp4[189] ), .Z(\MC_ARK_ARC_1_1/temp6[189] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_0_2  ( .A1(n1383), .A2(n134), .Z(
        \MC_ARK_ARC_1_1/temp4[189] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_0_2  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[99] ), 
        .A2(\MC_ARK_ARC_1_1/buf_datainput[63] ), .Z(
        \MC_ARK_ARC_1_1/temp3[189] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_0_2  ( .A1(\RI5[1][183] ), .A2(\RI5[1][189] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[189] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X4_0_1  ( .A1(\RI5[1][34] ), .A2(n114), .Z(
        \MC_ARK_ARC_1_1/temp4[190] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X3_0_1  ( .A1(\MC_ARK_ARC_1_1/buf_datainput[100] ), 
        .A2(\RI5[1][64] ), .Z(\MC_ARK_ARC_1_1/temp3[190] ) );
  XOR2_X1 \MC_ARK_ARC_1_1/X2_0_1  ( .A1(\RI5[1][136] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[160] ), .Z(\MC_ARK_ARC_1_1/temp2[190] )
         );
  XOR2_X1 \MC_ARK_ARC_1_1/X1_0_1  ( .A1(\RI5[1][190] ), .A2(\RI5[1][184] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[190] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_185  ( .I(\SB2_1_1/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[185] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_95  ( .I(\SB2_1_16/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[95] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_35  ( .I(\SB2_1_26/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[35] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_31_5  ( .A1(\MC_ARK_ARC_1_2/temp5[0] ), .A2(
        \MC_ARK_ARC_1_2/temp6[0] ), .Z(\MC_ARK_ARC_1_2/buf_output[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_31_5  ( .A1(\MC_ARK_ARC_1_2/temp3[0] ), .A2(
        \MC_ARK_ARC_1_2/temp4[0] ), .Z(\MC_ARK_ARC_1_2/temp6[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_31_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[36] ), 
        .A2(n504), .Z(\MC_ARK_ARC_1_2/temp4[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_31_5  ( .A1(\SB2_2_9/buf_output[0] ), .A2(
        \RI5[2][138] ), .Z(\MC_ARK_ARC_1_2/temp2[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_31_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[0] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[186] ), .Z(\MC_ARK_ARC_1_2/temp1[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_31_4  ( .A1(\RI5[2][37] ), .A2(n532), .Z(
        \MC_ARK_ARC_1_2/temp4[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_31_4  ( .A1(\RI5[2][163] ), .A2(\RI5[2][139] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_31_4  ( .A1(\RI5[2][187] ), .A2(\RI5[2][1] ), .Z(
        \MC_ARK_ARC_1_2/temp1[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_31_3  ( .A1(\MC_ARK_ARC_1_2/temp5[2] ), .A2(
        \MC_ARK_ARC_1_2/temp6[2] ), .Z(\MC_ARK_ARC_1_2/buf_output[2] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_31_3  ( .A1(\MC_ARK_ARC_1_2/temp3[2] ), .A2(
        \MC_ARK_ARC_1_2/temp4[2] ), .Z(\MC_ARK_ARC_1_2/temp6[2] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_31_3  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[38] ), 
        .A2(n182), .Z(\MC_ARK_ARC_1_2/temp4[2] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_31_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[39] ), 
        .A2(n456), .Z(\MC_ARK_ARC_1_2/temp4[3] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_31_2  ( .A1(\RI5[2][69] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[105] ), .Z(\MC_ARK_ARC_1_2/temp3[3] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_31_2  ( .A1(n1390), .A2(\RI5[2][3] ), .Z(
        \MC_ARK_ARC_1_2/temp1[3] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_31_1  ( .A1(\RI5[2][40] ), .A2(n485), .Z(
        \MC_ARK_ARC_1_2/temp4[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_31_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[4] ), 
        .A2(\RI5[2][190] ), .Z(\MC_ARK_ARC_1_2/temp1[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_31_0  ( .A1(\RI5[2][41] ), .A2(n193), .Z(
        \MC_ARK_ARC_1_2/temp4[5] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_30_5  ( .A1(\RI5[2][42] ), .A2(n206), .Z(
        \MC_ARK_ARC_1_2/temp4[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_30_5  ( .A1(\RI5[2][108] ), .A2(\RI5[2][72] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_30_4  ( .A1(\MC_ARK_ARC_1_2/temp3[7] ), .A2(
        \MC_ARK_ARC_1_2/temp4[7] ), .Z(\MC_ARK_ARC_1_2/temp6[7] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_30_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[43] ), 
        .A2(n80), .Z(\MC_ARK_ARC_1_2/temp4[7] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_30_4  ( .A1(\RI5[2][145] ), .A2(\RI5[2][169] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[7] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_30_3  ( .A1(\RI5[2][44] ), .A2(n465), .Z(
        \MC_ARK_ARC_1_2/temp4[8] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_30_3  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[2] ), 
        .A2(\RI5[2][8] ), .Z(\MC_ARK_ARC_1_2/temp1[8] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_30_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[45] ), 
        .A2(n495), .Z(\MC_ARK_ARC_1_2/temp4[9] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_30_1  ( .A1(\RI5[2][46] ), .A2(n211), .Z(
        \MC_ARK_ARC_1_2/temp4[10] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_30_1  ( .A1(\RI5[2][112] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[76] ), .Z(\MC_ARK_ARC_1_2/temp3[10] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_30_1  ( .A1(\RI5[2][10] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[4] ), .Z(\MC_ARK_ARC_1_2/temp1[10] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_30_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[47] ), 
        .A2(n549), .Z(\MC_ARK_ARC_1_2/temp4[11] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_30_0  ( .A1(\RI5[2][77] ), .A2(\RI5[2][113] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[11] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_30_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[149] ), 
        .A2(\RI5[2][173] ), .Z(\MC_ARK_ARC_1_2/temp2[11] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_29_5  ( .A1(\SB2_2_28/buf_output[0] ), .A2(n445), 
        .Z(\MC_ARK_ARC_1_2/temp4[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_29_4  ( .A1(\MC_ARK_ARC_1_2/temp3[13] ), .A2(
        \MC_ARK_ARC_1_2/temp4[13] ), .Z(\MC_ARK_ARC_1_2/temp6[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_29_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[49] ), 
        .A2(n473), .Z(\MC_ARK_ARC_1_2/temp4[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_29_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[115] ), 
        .A2(\RI5[2][79] ), .Z(\MC_ARK_ARC_1_2/temp3[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_29_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[175] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[151] ), .Z(
        \MC_ARK_ARC_1_2/temp2[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_29_4  ( .A1(\RI5[2][13] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[7] ), .Z(\MC_ARK_ARC_1_2/temp1[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_29_3  ( .A1(\RI5[2][8] ), .A2(n570), .Z(
        \MC_ARK_ARC_1_2/temp1[14] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_29_2  ( .A1(\RI5[2][51] ), .A2(n530), .Z(
        \MC_ARK_ARC_1_2/temp4[15] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_29_2  ( .A1(\RI5[2][15] ), .A2(\RI5[2][9] ), .Z(
        \MC_ARK_ARC_1_2/temp1[15] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_29_1  ( .A1(\MC_ARK_ARC_1_2/temp3[16] ), .A2(
        \MC_ARK_ARC_1_2/temp4[16] ), .Z(\MC_ARK_ARC_1_2/temp6[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_29_1  ( .A1(\RI5[2][52] ), .A2(n558), .Z(
        \MC_ARK_ARC_1_2/temp4[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_29_1  ( .A1(\RI5[2][118] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[82] ), .Z(\MC_ARK_ARC_1_2/temp3[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_29_1  ( .A1(\RI5[2][16] ), .A2(\RI5[2][10] ), .Z(
        \MC_ARK_ARC_1_2/temp1[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_29_0  ( .A1(\MC_ARK_ARC_1_2/temp3[17] ), .A2(
        \MC_ARK_ARC_1_2/temp4[17] ), .Z(\MC_ARK_ARC_1_2/temp6[17] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_29_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[53] ), 
        .A2(n195), .Z(\MC_ARK_ARC_1_2/temp4[17] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_28_5  ( .A1(\MC_ARK_ARC_1_2/temp2[18] ), .A2(
        \MC_ARK_ARC_1_2/temp1[18] ), .Z(\MC_ARK_ARC_1_2/temp5[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_28_5  ( .A1(\RI5[2][54] ), .A2(n213), .Z(
        \MC_ARK_ARC_1_2/temp4[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_28_5  ( .A1(\RI5[2][120] ), .A2(\RI5[2][84] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_28_5  ( .A1(\RI5[2][12] ), .A2(\RI5[2][18] ), .Z(
        \MC_ARK_ARC_1_2/temp1[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_28_4  ( .A1(\RI5[2][55] ), .A2(n512), .Z(
        \MC_ARK_ARC_1_2/temp4[19] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_28_4  ( .A1(\RI5[2][157] ), .A2(\RI5[2][181] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[19] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_28_4  ( .A1(\RI5[2][19] ), .A2(\RI5[2][13] ), .Z(
        \MC_ARK_ARC_1_2/temp1[19] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_28_3  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[56] ), 
        .A2(n541), .Z(\MC_ARK_ARC_1_2/temp4[20] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_28_2  ( .A1(\MC_ARK_ARC_1_2/temp5[21] ), .A2(
        \MC_ARK_ARC_1_2/temp6[21] ), .Z(\MC_ARK_ARC_1_2/buf_output[21] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_28_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[58] ), 
        .A2(n464), .Z(\MC_ARK_ARC_1_2/temp4[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_28_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[124] ), 
        .A2(\RI5[2][88] ), .Z(\MC_ARK_ARC_1_2/temp3[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_28_1  ( .A1(\RI5[2][184] ), .A2(\RI5[2][160] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_28_1  ( .A1(\RI5[2][22] ), .A2(\RI5[2][16] ), .Z(
        \MC_ARK_ARC_1_2/temp1[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_28_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[59] ), 
        .A2(n205), .Z(\MC_ARK_ARC_1_2/temp4[23] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_27_5  ( .A1(\MC_ARK_ARC_1_2/temp5[24] ), .A2(
        \MC_ARK_ARC_1_2/temp6[24] ), .Z(\MC_ARK_ARC_1_2/buf_output[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_27_5  ( .A1(\MC_ARK_ARC_1_2/temp3[24] ), .A2(
        \MC_ARK_ARC_1_2/temp4[24] ), .Z(\MC_ARK_ARC_1_2/temp6[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_27_5  ( .A1(\MC_ARK_ARC_1_2/temp2[24] ), .A2(
        \MC_ARK_ARC_1_2/temp1[24] ), .Z(\MC_ARK_ARC_1_2/temp5[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_27_5  ( .A1(\RI5[2][60] ), .A2(n520), .Z(
        \MC_ARK_ARC_1_2/temp4[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_27_5  ( .A1(\RI5[2][126] ), .A2(\RI5[2][90] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_27_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[186] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[162] ), .Z(
        \MC_ARK_ARC_1_2/temp2[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_27_5  ( .A1(\RI5[2][24] ), .A2(\RI5[2][18] ), .Z(
        \MC_ARK_ARC_1_2/temp1[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_27_4  ( .A1(\MC_ARK_ARC_1_2/temp5[25] ), .A2(
        \MC_ARK_ARC_1_2/temp6[25] ), .Z(\MC_ARK_ARC_1_2/buf_output[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_27_4  ( .A1(\MC_ARK_ARC_1_2/temp3[25] ), .A2(
        \MC_ARK_ARC_1_2/temp4[25] ), .Z(\MC_ARK_ARC_1_2/temp6[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_27_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[61] ), 
        .A2(n235), .Z(\MC_ARK_ARC_1_2/temp4[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_27_4  ( .A1(\RI5[2][163] ), .A2(\RI5[2][187] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_27_3  ( .A1(\RI5[2][62] ), .A2(n238), .Z(
        \MC_ARK_ARC_1_2/temp4[26] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_27_2  ( .A1(\RI5[2][63] ), .A2(n472), .Z(
        \MC_ARK_ARC_1_2/temp4[27] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_27_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[129] ), 
        .A2(\RI5[2][93] ), .Z(\MC_ARK_ARC_1_2/temp3[27] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_27_2  ( .A1(\RI5[2][165] ), .A2(\RI5[2][189] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[27] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_27_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[27] ), 
        .A2(\RI5[2][21] ), .Z(\MC_ARK_ARC_1_2/temp1[27] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_27_1  ( .A1(\MC_ARK_ARC_1_2/temp3[28] ), .A2(
        \MC_ARK_ARC_1_2/temp4[28] ), .Z(\MC_ARK_ARC_1_2/temp6[28] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_27_1  ( .A1(\RI5[2][64] ), .A2(n187), .Z(
        \MC_ARK_ARC_1_2/temp4[28] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_27_1  ( .A1(\RI5[2][130] ), .A2(\RI5[2][94] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[28] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_27_1  ( .A1(\RI5[2][190] ), .A2(\RI5[2][166] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[28] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_27_1  ( .A1(\RI5[2][28] ), .A2(\RI5[2][22] ), .Z(
        \MC_ARK_ARC_1_2/temp1[28] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_27_0  ( .A1(\RI5[2][167] ), .A2(\RI5[2][191] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[29] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_26_5  ( .A1(\RI5[2][66] ), .A2(n208), .Z(
        \MC_ARK_ARC_1_2/temp4[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_26_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[132] ), 
        .A2(\RI5[2][96] ), .Z(\MC_ARK_ARC_1_2/temp3[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_26_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[30] ), 
        .A2(\RI5[2][24] ), .Z(\MC_ARK_ARC_1_2/temp1[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_26_4  ( .A1(\RI5[2][67] ), .A2(n452), .Z(
        \MC_ARK_ARC_1_2/temp4[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_26_4  ( .A1(\RI5[2][1] ), .A2(\RI5[2][169] ), .Z(
        \MC_ARK_ARC_1_2/temp2[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_26_2  ( .A1(\RI5[2][69] ), .A2(n31), .Z(
        \MC_ARK_ARC_1_2/temp4[33] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_26_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[99] ), 
        .A2(\RI5[2][135] ), .Z(\MC_ARK_ARC_1_2/temp3[33] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_26_2  ( .A1(\RI5[2][171] ), .A2(\RI5[2][3] ), .Z(
        \MC_ARK_ARC_1_2/temp2[33] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_26_1  ( .A1(\MC_ARK_ARC_1_2/temp1[34] ), .A2(
        \MC_ARK_ARC_1_2/temp2[34] ), .Z(\MC_ARK_ARC_1_2/temp5[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_26_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[70] ), 
        .A2(\MC_ARK_ARC_1_1/buf_keyinput[51] ), .Z(\MC_ARK_ARC_1_2/temp4[34] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_26_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[136] ), 
        .A2(\RI5[2][100] ), .Z(\MC_ARK_ARC_1_2/temp3[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_26_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[4] ), 
        .A2(\RI5[2][172] ), .Z(\MC_ARK_ARC_1_2/temp2[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_26_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[34] ), 
        .A2(\RI5[2][28] ), .Z(\MC_ARK_ARC_1_2/temp1[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_26_0  ( .A1(\RI5[2][71] ), .A2(n564), .Z(
        \MC_ARK_ARC_1_2/temp4[35] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_25_5  ( .A1(\MC_ARK_ARC_1_2/temp6[36] ), .A2(
        \MC_ARK_ARC_1_2/temp5[36] ), .Z(\MC_ARK_ARC_1_2/buf_output[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_25_5  ( .A1(\MC_ARK_ARC_1_2/temp3[36] ), .A2(
        \MC_ARK_ARC_1_2/temp4[36] ), .Z(\MC_ARK_ARC_1_2/temp6[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_25_5  ( .A1(\MC_ARK_ARC_1_2/temp2[36] ), .A2(
        \MC_ARK_ARC_1_2/temp1[36] ), .Z(\MC_ARK_ARC_1_2/temp5[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_25_5  ( .A1(\RI5[2][72] ), .A2(n462), .Z(
        \MC_ARK_ARC_1_2/temp4[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_25_5  ( .A1(\RI5[2][138] ), .A2(\RI5[2][102] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_25_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[6] ), 
        .A2(\RI5[2][174] ), .Z(\MC_ARK_ARC_1_2/temp2[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_25_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[36] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[30] ), .Z(\MC_ARK_ARC_1_2/temp1[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_25_4  ( .A1(\MC_ARK_ARC_1_2/temp1[37] ), .A2(
        \MC_ARK_ARC_1_2/temp2[37] ), .Z(\MC_ARK_ARC_1_2/temp5[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_25_4  ( .A1(\RI5[2][73] ), .A2(n148), .Z(
        \MC_ARK_ARC_1_2/temp4[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_25_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[7] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[175] ), .Z(
        \MC_ARK_ARC_1_2/temp2[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_25_4  ( .A1(\RI5[2][31] ), .A2(\RI5[2][37] ), .Z(
        \MC_ARK_ARC_1_2/temp1[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_25_3  ( .A1(\RI5[2][176] ), .A2(\RI5[2][8] ), .Z(
        \MC_ARK_ARC_1_2/temp2[38] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_25_3  ( .A1(\RI5[2][32] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[38] ), .Z(\MC_ARK_ARC_1_2/temp1[38] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_25_2  ( .A1(\RI5[2][75] ), .A2(n546), .Z(
        \MC_ARK_ARC_1_2/temp4[39] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_25_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[141] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[105] ), .Z(
        \MC_ARK_ARC_1_2/temp3[39] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_25_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[39] ), 
        .A2(\RI5[2][33] ), .Z(\MC_ARK_ARC_1_2/temp1[39] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_25_1  ( .A1(\MC_ARK_ARC_1_2/temp5[40] ), .A2(
        \MC_ARK_ARC_1_2/temp6[40] ), .Z(\MC_ARK_ARC_1_2/buf_output[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_25_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[76] ), 
        .A2(n443), .Z(\MC_ARK_ARC_1_2/temp4[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_25_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[106] ), 
        .A2(\RI5[2][142] ), .Z(\MC_ARK_ARC_1_2/temp3[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_25_1  ( .A1(\RI5[2][178] ), .A2(\RI5[2][10] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_25_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[34] ), 
        .A2(\RI5[2][40] ), .Z(\MC_ARK_ARC_1_2/temp1[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_25_0  ( .A1(\MC_ARK_ARC_1_2/temp3[41] ), .A2(
        \MC_ARK_ARC_1_2/temp4[41] ), .Z(\MC_ARK_ARC_1_2/temp6[41] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_25_0  ( .A1(\RI5[2][77] ), .A2(n127), .Z(
        \MC_ARK_ARC_1_2/temp4[41] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_25_0  ( .A1(\RI5[2][143] ), .A2(\RI5[2][107] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[41] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_25_0  ( .A1(\RI5[2][11] ), .A2(\RI5[2][179] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[41] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_25_0  ( .A1(\RI5[2][41] ), .A2(\RI5[2][35] ), .Z(
        \MC_ARK_ARC_1_2/temp1[41] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_24_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[78] ), 
        .A2(n500), .Z(\MC_ARK_ARC_1_2/temp4[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_24_5  ( .A1(\RI5[2][144] ), .A2(\RI5[2][108] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_24_5  ( .A1(\RI5[2][42] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[36] ), .Z(\MC_ARK_ARC_1_2/temp1[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_24_4  ( .A1(\RI5[2][79] ), .A2(n217), .Z(
        \MC_ARK_ARC_1_2/temp4[43] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_24_4  ( .A1(\RI5[2][109] ), .A2(\RI5[2][145] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[43] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_24_4  ( .A1(\RI5[2][13] ), .A2(\RI5[2][181] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[43] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_24_3  ( .A1(\RI5[2][80] ), .A2(n556), .Z(
        \MC_ARK_ARC_1_2/temp4[44] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_24_3  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[182] ), 
        .A2(n570), .Z(\MC_ARK_ARC_1_2/temp2[44] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_24_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[81] ), 
        .A2(n159), .Z(\MC_ARK_ARC_1_2/temp4[45] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_24_1  ( .A1(\MC_ARK_ARC_1_2/temp3[46] ), .A2(
        \MC_ARK_ARC_1_2/temp4[46] ), .Z(\MC_ARK_ARC_1_2/temp6[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_24_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[82] ), 
        .A2(n480), .Z(\MC_ARK_ARC_1_2/temp4[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_24_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[148] ), 
        .A2(\RI5[2][112] ), .Z(\MC_ARK_ARC_1_2/temp3[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_24_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[83] ), 
        .A2(n509), .Z(\MC_ARK_ARC_1_2/temp4[47] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_23_5  ( .A1(\MC_ARK_ARC_1_2/temp1[48] ), .A2(
        \MC_ARK_ARC_1_2/temp2[48] ), .Z(\MC_ARK_ARC_1_2/temp5[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_23_5  ( .A1(\RI5[2][84] ), .A2(n153), .Z(
        \MC_ARK_ARC_1_2/temp4[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_23_5  ( .A1(\RI5[2][18] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[186] ), .Z(\MC_ARK_ARC_1_2/temp2[48] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_23_4  ( .A1(\RI5[2][85] ), .A2(n563), .Z(
        \MC_ARK_ARC_1_2/temp4[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_23_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[115] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[151] ), .Z(
        \MC_ARK_ARC_1_2/temp3[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_23_4  ( .A1(\RI5[2][19] ), .A2(\RI5[2][187] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_23_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[49] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[43] ), .Z(\MC_ARK_ARC_1_2/temp1[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_23_2  ( .A1(\RI5[2][87] ), .A2(n45), .Z(
        \MC_ARK_ARC_1_2/temp4[51] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_23_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[153] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[117] ), .Z(
        \MC_ARK_ARC_1_2/temp3[51] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_23_1  ( .A1(\MC_ARK_ARC_1_2/temp1[52] ), .A2(
        \MC_ARK_ARC_1_2/temp2[52] ), .Z(\MC_ARK_ARC_1_2/temp5[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_23_1  ( .A1(\RI5[2][22] ), .A2(\RI5[2][190] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_23_1  ( .A1(\RI5[2][52] ), .A2(\RI5[2][46] ), .Z(
        \MC_ARK_ARC_1_2/temp1[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_23_0  ( .A1(\RI5[2][89] ), .A2(n227), .Z(
        \MC_ARK_ARC_1_2/temp4[53] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_23_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[53] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[47] ), .Z(\MC_ARK_ARC_1_2/temp1[53] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_22_5  ( .A1(\MC_ARK_ARC_1_2/temp5[54] ), .A2(
        \MC_ARK_ARC_1_2/temp6[54] ), .Z(\MC_ARK_ARC_1_2/buf_output[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_22_5  ( .A1(\MC_ARK_ARC_1_2/temp3[54] ), .A2(
        \MC_ARK_ARC_1_2/temp4[54] ), .Z(\MC_ARK_ARC_1_2/temp6[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_22_5  ( .A1(\MC_ARK_ARC_1_2/temp1[54] ), .A2(
        \MC_ARK_ARC_1_2/temp2[54] ), .Z(\MC_ARK_ARC_1_2/temp5[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_22_5  ( .A1(\RI5[2][90] ), .A2(
        \MC_ARK_ARC_1_2/buf_keyinput[54] ), .Z(\MC_ARK_ARC_1_2/temp4[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_22_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[156] ), 
        .A2(\RI5[2][120] ), .Z(\MC_ARK_ARC_1_2/temp3[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_22_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[0] ), 
        .A2(\RI5[2][24] ), .Z(\MC_ARK_ARC_1_2/temp2[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_22_4  ( .A1(\MC_ARK_ARC_1_2/temp1[55] ), .A2(
        \MC_ARK_ARC_1_2/temp2[55] ), .Z(\MC_ARK_ARC_1_2/temp5[55] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_22_4  ( .A1(\RI5[2][91] ), .A2(n233), .Z(
        \MC_ARK_ARC_1_2/temp4[55] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_22_4  ( .A1(\SB2_2_3/buf_output[1] ), .A2(
        \RI5[2][25] ), .Z(\MC_ARK_ARC_1_2/temp2[55] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_22_4  ( .A1(\RI5[2][55] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[49] ), .Z(\MC_ARK_ARC_1_2/temp1[55] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_22_3  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[92] ), 
        .A2(n190), .Z(\MC_ARK_ARC_1_2/temp4[56] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_22_2  ( .A1(\RI5[2][93] ), .A2(n525), .Z(
        \MC_ARK_ARC_1_2/temp4[57] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_22_2  ( .A1(\RI5[2][51] ), .A2(\RI5[2][57] ), .Z(
        \MC_ARK_ARC_1_2/temp1[57] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_22_1  ( .A1(\RI5[2][94] ), .A2(n84), .Z(
        \MC_ARK_ARC_1_2/temp4[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_22_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[58] ), 
        .A2(\RI5[2][52] ), .Z(\MC_ARK_ARC_1_2/temp1[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_22_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[95] ), 
        .A2(n129), .Z(\MC_ARK_ARC_1_2/temp4[59] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_22_0  ( .A1(\RI5[2][161] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[125] ), .Z(\MC_ARK_ARC_1_2/temp3[59] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_21_5  ( .A1(\MC_ARK_ARC_1_2/temp3[60] ), .A2(
        \MC_ARK_ARC_1_2/temp4[60] ), .Z(\MC_ARK_ARC_1_2/temp6[60] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_21_5  ( .A1(\RI5[2][96] ), .A2(n478), .Z(
        \MC_ARK_ARC_1_2/temp4[60] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_21_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[162] ), 
        .A2(\RI5[2][126] ), .Z(\MC_ARK_ARC_1_2/temp3[60] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_21_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[30] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[6] ), .Z(\MC_ARK_ARC_1_2/temp2[60] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_21_5  ( .A1(\RI5[2][60] ), .A2(\RI5[2][54] ), .Z(
        \MC_ARK_ARC_1_2/temp1[60] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_21_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[97] ), 
        .A2(n163), .Z(\MC_ARK_ARC_1_2/temp4[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_21_4  ( .A1(\RI5[2][163] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[127] ), .Z(\MC_ARK_ARC_1_2/temp3[61] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_21_4  ( .A1(\RI5[2][31] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[7] ), .Z(\MC_ARK_ARC_1_2/temp2[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_21_4  ( .A1(\RI5[2][55] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[61] ), .Z(\MC_ARK_ARC_1_2/temp1[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_21_3  ( .A1(\RI5[2][98] ), .A2(n244), .Z(
        \MC_ARK_ARC_1_2/temp4[62] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_21_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[99] ), 
        .A2(n561), .Z(\MC_ARK_ARC_1_2/temp4[63] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_21_2  ( .A1(\RI5[2][57] ), .A2(\RI5[2][63] ), .Z(
        \MC_ARK_ARC_1_2/temp1[63] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_21_1  ( .A1(\RI5[2][100] ), .A2(n460), .Z(
        \MC_ARK_ARC_1_2/temp4[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_21_0  ( .A1(\MC_ARK_ARC_1_2/temp3[65] ), .A2(
        \MC_ARK_ARC_1_2/temp4[65] ), .Z(\MC_ARK_ARC_1_2/temp6[65] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_21_0  ( .A1(\RI5[2][101] ), .A2(n489), .Z(
        \MC_ARK_ARC_1_2/temp4[65] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_21_0  ( .A1(\RI5[2][167] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[131] ), .Z(\MC_ARK_ARC_1_2/temp3[65] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_20_5  ( .A1(\MC_ARK_ARC_1_2/temp6[66] ), .A2(
        \MC_ARK_ARC_1_2/temp5[66] ), .Z(\MC_ARK_ARC_1_2/buf_output[66] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_20_5  ( .A1(\MC_ARK_ARC_1_2/temp2[66] ), .A2(
        \MC_ARK_ARC_1_2/temp1[66] ), .Z(\MC_ARK_ARC_1_2/temp5[66] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_20_5  ( .A1(\RI5[2][102] ), .A2(n111), .Z(
        \MC_ARK_ARC_1_2/temp4[66] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_20_5  ( .A1(\RI5[2][168] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[132] ), .Z(\MC_ARK_ARC_1_2/temp3[66] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_20_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[36] ), 
        .A2(\RI5[2][12] ), .Z(\MC_ARK_ARC_1_2/temp2[66] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_20_5  ( .A1(\RI5[2][66] ), .A2(\RI5[2][60] ), .Z(
        \MC_ARK_ARC_1_2/temp1[66] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_20_4  ( .A1(\MC_ARK_ARC_1_2/temp4[67] ), .A2(
        \MC_ARK_ARC_1_2/temp3[67] ), .Z(\MC_ARK_ARC_1_2/temp6[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_20_4  ( .A1(\RI5[2][103] ), .A2(n185), .Z(
        \MC_ARK_ARC_1_2/temp4[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_20_4  ( .A1(\RI5[2][169] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[133] ), .Z(\MC_ARK_ARC_1_2/temp3[67] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_20_4  ( .A1(\RI5[2][13] ), .A2(\RI5[2][37] ), .Z(
        \MC_ARK_ARC_1_2/temp2[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_20_4  ( .A1(\RI5[2][67] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[61] ), .Z(\MC_ARK_ARC_1_2/temp1[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_20_3  ( .A1(\RI5[2][104] ), .A2(n441), .Z(
        \MC_ARK_ARC_1_2/temp4[68] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_20_3  ( .A1(\RI5[2][134] ), .A2(\RI5[2][170] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[68] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_20_3  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[38] ), 
        .A2(n570), .Z(\MC_ARK_ARC_1_2/temp2[68] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_20_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[105] ), 
        .A2(n72), .Z(\MC_ARK_ARC_1_2/temp4[69] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_20_2  ( .A1(\RI5[2][171] ), .A2(\RI5[2][135] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[69] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_20_2  ( .A1(\RI5[2][15] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[39] ), .Z(\MC_ARK_ARC_1_2/temp2[69] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_20_1  ( .A1(\MC_ARK_ARC_1_2/temp3[70] ), .A2(
        \MC_ARK_ARC_1_2/temp4[70] ), .Z(\MC_ARK_ARC_1_2/temp6[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_20_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[106] ), 
        .A2(n209), .Z(\MC_ARK_ARC_1_2/temp4[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_20_1  ( .A1(\RI5[2][40] ), .A2(\RI5[2][16] ), .Z(
        \MC_ARK_ARC_1_2/temp2[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_20_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[70] ), 
        .A2(\RI5[2][64] ), .Z(\MC_ARK_ARC_1_2/temp1[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_20_0  ( .A1(\MC_ARK_ARC_1_2/temp4[71] ), .A2(
        \MC_ARK_ARC_1_2/temp3[71] ), .Z(\MC_ARK_ARC_1_2/temp6[71] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_20_0  ( .A1(\RI5[2][107] ), .A2(n207), .Z(
        \MC_ARK_ARC_1_2/temp4[71] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_20_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[65] ), 
        .A2(\RI5[2][71] ), .Z(\MC_ARK_ARC_1_2/temp1[71] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_19_5  ( .A1(\RI5[2][42] ), .A2(\RI5[2][18] ), .Z(
        \MC_ARK_ARC_1_2/temp2[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_19_4  ( .A1(\RI5[2][109] ), .A2(n165), .Z(
        \MC_ARK_ARC_1_2/temp4[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_19_4  ( .A1(\RI5[2][19] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[43] ), .Z(\MC_ARK_ARC_1_2/temp2[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_19_4  ( .A1(\RI5[2][73] ), .A2(\RI5[2][67] ), .Z(
        \MC_ARK_ARC_1_2/temp1[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_19_3  ( .A1(\RI5[2][110] ), .A2(n94), .Z(
        \MC_ARK_ARC_1_2/temp4[74] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_19_3  ( .A1(\RI5[2][140] ), .A2(\RI5[2][176] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[74] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_19_3  ( .A1(\RI5[2][20] ), .A2(\RI5[2][44] ), .Z(
        \MC_ARK_ARC_1_2/temp2[74] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_19_2  ( .A1(\RI5[2][111] ), .A2(n506), .Z(
        \MC_ARK_ARC_1_2/temp4[75] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_19_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[45] ), 
        .A2(\RI5[2][21] ), .Z(\MC_ARK_ARC_1_2/temp2[75] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_19_1  ( .A1(\RI5[2][112] ), .A2(n70), .Z(
        \MC_ARK_ARC_1_2/temp4[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_19_1  ( .A1(\RI5[2][178] ), .A2(\RI5[2][142] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_19_1  ( .A1(\RI5[2][22] ), .A2(\RI5[2][46] ), .Z(
        \MC_ARK_ARC_1_2/temp2[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_19_0  ( .A1(\MC_ARK_ARC_1_2/temp6[77] ), .A2(
        \MC_ARK_ARC_1_2/temp5[77] ), .Z(\MC_ARK_ARC_1_2/buf_output[77] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_19_0  ( .A1(\MC_ARK_ARC_1_2/temp3[77] ), .A2(
        \MC_ARK_ARC_1_2/temp4[77] ), .Z(\MC_ARK_ARC_1_2/temp6[77] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_19_0  ( .A1(\RI5[2][113] ), .A2(n214), .Z(
        \MC_ARK_ARC_1_2/temp4[77] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_19_0  ( .A1(\RI5[2][143] ), .A2(\RI5[2][179] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[77] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_18_5  ( .A1(\MC_ARK_ARC_1_2/temp5[78] ), .A2(
        \MC_ARK_ARC_1_2/temp6[78] ), .Z(\MC_ARK_ARC_1_2/buf_output[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_18_5  ( .A1(\MC_ARK_ARC_1_2/temp3[78] ), .A2(
        \MC_ARK_ARC_1_2/temp4[78] ), .Z(\MC_ARK_ARC_1_2/temp6[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_18_5  ( .A1(\MC_ARK_ARC_1_2/temp2[78] ), .A2(
        \MC_ARK_ARC_1_2/temp1[78] ), .Z(\MC_ARK_ARC_1_2/temp5[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_18_5  ( .A1(\RI5[2][114] ), .A2(n215), .Z(
        \MC_ARK_ARC_1_2/temp4[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_18_5  ( .A1(\RI5[2][144] ), .A2(\RI5[2][180] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_18_5  ( .A1(\RI5[2][48] ), .A2(\RI5[2][24] ), .Z(
        \MC_ARK_ARC_1_2/temp2[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_18_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[78] ), 
        .A2(\RI5[2][72] ), .Z(\MC_ARK_ARC_1_2/temp1[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_18_4  ( .A1(\MC_ARK_ARC_1_2/temp5[79] ), .A2(
        \MC_ARK_ARC_1_2/temp6[79] ), .Z(\MC_ARK_ARC_1_2/buf_output[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_18_4  ( .A1(\MC_ARK_ARC_1_2/temp3[79] ), .A2(
        \MC_ARK_ARC_1_2/temp4[79] ), .Z(\MC_ARK_ARC_1_2/temp6[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_18_4  ( .A1(\MC_ARK_ARC_1_2/temp1[79] ), .A2(
        \MC_ARK_ARC_1_2/temp2[79] ), .Z(\MC_ARK_ARC_1_2/temp5[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_18_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[115] ), 
        .A2(n64), .Z(\MC_ARK_ARC_1_2/temp4[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_18_4  ( .A1(\RI5[2][145] ), .A2(\RI5[2][181] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_18_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[49] ), 
        .A2(\RI5[2][25] ), .Z(\MC_ARK_ARC_1_2/temp2[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_18_4  ( .A1(\RI5[2][73] ), .A2(\RI5[2][79] ), .Z(
        \MC_ARK_ARC_1_2/temp1[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_18_3  ( .A1(\MC_ARK_ARC_1_2/temp3[80] ), .A2(
        \MC_ARK_ARC_1_2/temp4[80] ), .Z(\MC_ARK_ARC_1_2/temp6[80] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_18_3  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[116] ), 
        .A2(n516), .Z(\MC_ARK_ARC_1_2/temp4[80] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_18_3  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[146] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[182] ), .Z(
        \MC_ARK_ARC_1_2/temp3[80] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_18_2  ( .A1(\MC_ARK_ARC_1_2/temp3[81] ), .A2(
        \MC_ARK_ARC_1_2/temp4[81] ), .Z(\MC_ARK_ARC_1_2/temp6[81] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_18_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[117] ), 
        .A2(n544), .Z(\MC_ARK_ARC_1_2/temp4[81] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_18_2  ( .A1(\RI5[2][147] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[183] ), .Z(\MC_ARK_ARC_1_2/temp3[81] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_18_1  ( .A1(\RI5[2][118] ), .A2(n439), .Z(
        \MC_ARK_ARC_1_2/temp4[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_18_1  ( .A1(\RI5[2][184] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[148] ), .Z(\MC_ARK_ARC_1_2/temp3[82] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_18_1  ( .A1(\RI5[2][28] ), .A2(\RI5[2][52] ), .Z(
        \MC_ARK_ARC_1_2/temp2[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_18_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[82] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[76] ), .Z(\MC_ARK_ARC_1_2/temp1[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_18_0  ( .A1(\RI5[2][119] ), .A2(n100), .Z(
        \MC_ARK_ARC_1_2/temp4[83] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_18_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[29] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[53] ), .Z(\MC_ARK_ARC_1_2/temp2[83] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_17_5  ( .A1(\MC_ARK_ARC_1_2/temp3[84] ), .A2(
        \MC_ARK_ARC_1_2/temp4[84] ), .Z(\MC_ARK_ARC_1_2/temp6[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_17_5  ( .A1(\MC_ARK_ARC_1_2/temp1[84] ), .A2(
        \MC_ARK_ARC_1_2/temp2[84] ), .Z(\MC_ARK_ARC_1_2/temp5[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_17_5  ( .A1(\RI5[2][120] ), .A2(n138), .Z(
        \MC_ARK_ARC_1_2/temp4[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_17_5  ( .A1(\RI5[2][150] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[186] ), .Z(\MC_ARK_ARC_1_2/temp3[84] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_17_5  ( .A1(\RI5[2][54] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[30] ), .Z(\MC_ARK_ARC_1_2/temp2[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_17_5  ( .A1(\RI5[2][84] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[78] ), .Z(\MC_ARK_ARC_1_2/temp1[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_17_4  ( .A1(\MC_ARK_ARC_1_2/temp3[85] ), .A2(
        \MC_ARK_ARC_1_2/temp4[85] ), .Z(\MC_ARK_ARC_1_2/temp6[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_17_4  ( .A1(\RI5[2][121] ), .A2(n97), .Z(
        \MC_ARK_ARC_1_2/temp4[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_17_4  ( .A1(\RI5[2][31] ), .A2(\RI5[2][55] ), .Z(
        \MC_ARK_ARC_1_2/temp2[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_17_3  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[122] ), 
        .A2(n552), .Z(\MC_ARK_ARC_1_2/temp4[86] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_17_2  ( .A1(\RI5[2][123] ), .A2(n47), .Z(
        \MC_ARK_ARC_1_2/temp4[87] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_17_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[124] ), 
        .A2(n475), .Z(\MC_ARK_ARC_1_2/temp4[88] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_17_1  ( .A1(\RI5[2][88] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[82] ), .Z(\MC_ARK_ARC_1_2/temp1[88] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_17_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[125] ), 
        .A2(n63), .Z(\MC_ARK_ARC_1_2/temp4[89] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_16_5  ( .A1(\RI5[2][126] ), .A2(n533), .Z(
        \MC_ARK_ARC_1_2/temp4[90] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_16_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[127] ), 
        .A2(n170), .Z(\MC_ARK_ARC_1_2/temp4[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_16_4  ( .A1(\RI5[2][157] ), .A2(\RI5[2][1] ), .Z(
        \MC_ARK_ARC_1_2/temp3[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_16_4  ( .A1(\RI5[2][91] ), .A2(\RI5[2][85] ), .Z(
        \MC_ARK_ARC_1_2/temp1[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_16_3  ( .A1(\SB2_2_13/buf_output[2] ), .A2(n457), 
        .Z(\MC_ARK_ARC_1_2/temp4[92] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_16_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[129] ), 
        .A2(n486), .Z(\MC_ARK_ARC_1_2/temp4[93] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_16_1  ( .A1(\MC_ARK_ARC_1_2/temp3[94] ), .A2(
        \MC_ARK_ARC_1_2/temp4[94] ), .Z(\MC_ARK_ARC_1_2/temp6[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_16_1  ( .A1(\RI5[2][130] ), .A2(n89), .Z(
        \MC_ARK_ARC_1_2/temp4[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_16_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[4] ), 
        .A2(\RI5[2][160] ), .Z(\MC_ARK_ARC_1_2/temp3[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_16_1  ( .A1(\RI5[2][40] ), .A2(\RI5[2][64] ), .Z(
        \MC_ARK_ARC_1_2/temp2[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_16_1  ( .A1(\RI5[2][94] ), .A2(\RI5[2][88] ), .Z(
        \MC_ARK_ARC_1_2/temp1[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_16_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[131] ), 
        .A2(n542), .Z(\MC_ARK_ARC_1_2/temp4[95] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_16_0  ( .A1(\RI5[2][89] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[95] ), .Z(\MC_ARK_ARC_1_2/temp1[95] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_15_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[132] ), 
        .A2(n438), .Z(\MC_ARK_ARC_1_2/temp4[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_15_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[162] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[6] ), .Z(\MC_ARK_ARC_1_2/temp3[96] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_15_5  ( .A1(\RI5[2][96] ), .A2(\RI5[2][90] ), .Z(
        \MC_ARK_ARC_1_2/temp1[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_15_4  ( .A1(\MC_ARK_ARC_1_2/temp5[97] ), .A2(
        \MC_ARK_ARC_1_2/temp6[97] ), .Z(\MC_ARK_ARC_1_2/buf_output[97] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_15_4  ( .A1(\SB2_2_13/buf_output[1] ), .A2(n135), 
        .Z(\MC_ARK_ARC_1_2/temp4[97] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_15_4  ( .A1(\SB2_2_8/buf_output[1] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[7] ), .Z(\MC_ARK_ARC_1_2/temp3[97] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_15_4  ( .A1(\RI5[2][67] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[43] ), .Z(\MC_ARK_ARC_1_2/temp2[97] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_15_2  ( .A1(\RI5[2][135] ), .A2(n224), .Z(
        \MC_ARK_ARC_1_2/temp4[99] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_15_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[136] ), 
        .A2(n550), .Z(\MC_ARK_ARC_1_2/temp4[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_15_1  ( .A1(\RI5[2][10] ), .A2(\RI5[2][166] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_15_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[70] ), 
        .A2(\RI5[2][46] ), .Z(\MC_ARK_ARC_1_2/temp2[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_14_5  ( .A1(\MC_ARK_ARC_1_2/temp2[102] ), .A2(
        \MC_ARK_ARC_1_2/temp1[102] ), .Z(\MC_ARK_ARC_1_2/temp5[102] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_14_5  ( .A1(\RI5[2][138] ), .A2(n197), .Z(
        \MC_ARK_ARC_1_2/temp4[102] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_14_5  ( .A1(\RI5[2][168] ), .A2(\RI5[2][12] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[102] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_14_5  ( .A1(\RI5[2][102] ), .A2(\RI5[2][96] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[102] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_14_4  ( .A1(\RI5[2][139] ), .A2(n503), .Z(
        \MC_ARK_ARC_1_2/temp4[103] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_14_4  ( .A1(\RI5[2][13] ), .A2(\RI5[2][169] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[103] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_14_4  ( .A1(\RI5[2][73] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[49] ), .Z(\MC_ARK_ARC_1_2/temp2[103] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_14_4  ( .A1(\RI5[2][103] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[97] ), .Z(\MC_ARK_ARC_1_2/temp1[103] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_14_3  ( .A1(\RI5[2][140] ), .A2(n531), .Z(
        \MC_ARK_ARC_1_2/temp4[104] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_14_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[141] ), 
        .A2(n132), .Z(\MC_ARK_ARC_1_2/temp4[105] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_14_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[99] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[105] ), .Z(
        \MC_ARK_ARC_1_2/temp1[105] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_14_1  ( .A1(\MC_ARK_ARC_1_2/temp6[106] ), .A2(
        \MC_ARK_ARC_1_2/temp5[106] ), .Z(\MC_ARK_ARC_1_2/buf_output[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_14_1  ( .A1(\MC_ARK_ARC_1_2/temp3[106] ), .A2(
        \MC_ARK_ARC_1_2/temp4[106] ), .Z(\MC_ARK_ARC_1_2/temp6[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_14_1  ( .A1(\MC_ARK_ARC_1_2/temp1[106] ), .A2(
        \MC_ARK_ARC_1_2/temp2[106] ), .Z(\MC_ARK_ARC_1_2/temp5[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_14_1  ( .A1(\RI5[2][142] ), .A2(n455), .Z(
        \MC_ARK_ARC_1_2/temp4[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_14_1  ( .A1(\RI5[2][16] ), .A2(\RI5[2][172] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_14_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[76] ), 
        .A2(\RI5[2][52] ), .Z(\MC_ARK_ARC_1_2/temp2[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_14_1  ( .A1(\RI5[2][100] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[106] ), .Z(\MC_ARK_ARC_1_2/temp1[106] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_14_0  ( .A1(\RI5[2][143] ), .A2(n106), .Z(
        \MC_ARK_ARC_1_2/temp4[107] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_13_5  ( .A1(\MC_ARK_ARC_1_2/temp3[108] ), .A2(
        \MC_ARK_ARC_1_2/temp4[108] ), .Z(\MC_ARK_ARC_1_2/temp6[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_13_5  ( .A1(\MC_ARK_ARC_1_2/temp1[108] ), .A2(
        \MC_ARK_ARC_1_2/temp2[108] ), .Z(\MC_ARK_ARC_1_2/temp5[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_13_5  ( .A1(\RI5[2][144] ), .A2(n513), .Z(
        \MC_ARK_ARC_1_2/temp4[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_13_5  ( .A1(\RI5[2][18] ), .A2(\RI5[2][174] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_13_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[78] ), 
        .A2(\RI5[2][54] ), .Z(\MC_ARK_ARC_1_2/temp2[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_13_5  ( .A1(\RI5[2][108] ), .A2(\RI5[2][102] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_13_4  ( .A1(\MC_ARK_ARC_1_2/temp3[109] ), .A2(
        \MC_ARK_ARC_1_2/temp4[109] ), .Z(\MC_ARK_ARC_1_2/temp6[109] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_13_4  ( .A1(\RI5[2][145] ), .A2(n169), .Z(
        \MC_ARK_ARC_1_2/temp4[109] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_13_4  ( .A1(\RI5[2][19] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[175] ), .Z(\MC_ARK_ARC_1_2/temp3[109] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_13_3  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[146] ), 
        .A2(n1), .Z(\MC_ARK_ARC_1_2/temp4[110] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_13_3  ( .A1(\RI5[2][176] ), .A2(\RI5[2][20] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[110] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_13_2  ( .A1(\RI5[2][147] ), .A2(n41), .Z(
        \MC_ARK_ARC_1_2/temp4[111] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_13_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[105] ), 
        .A2(\RI5[2][111] ), .Z(\MC_ARK_ARC_1_2/temp1[111] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_13_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[148] ), 
        .A2(n5), .Z(\MC_ARK_ARC_1_2/temp4[112] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_13_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[82] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[58] ), .Z(
        \MC_ARK_ARC_1_2/temp2[112] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_13_1  ( .A1(\RI5[2][112] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[106] ), .Z(\MC_ARK_ARC_1_2/temp1[112] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_13_0  ( .A1(\MC_ARK_ARC_1_2/temp3[113] ), .A2(
        \MC_ARK_ARC_1_2/temp4[113] ), .Z(\MC_ARK_ARC_1_2/temp6[113] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_13_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[149] ), 
        .A2(n125), .Z(\MC_ARK_ARC_1_2/temp4[113] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_13_0  ( .A1(\RI5[2][107] ), .A2(\RI5[2][113] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[113] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_12_5  ( .A1(\MC_ARK_ARC_1_2/temp4[114] ), .A2(
        \MC_ARK_ARC_1_2/temp3[114] ), .Z(\MC_ARK_ARC_1_2/temp6[114] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_12_5  ( .A1(\MC_ARK_ARC_1_2/temp1[114] ), .A2(
        \MC_ARK_ARC_1_2/temp2[114] ), .Z(\MC_ARK_ARC_1_2/temp5[114] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_12_5  ( .A1(\RI5[2][150] ), .A2(n548), .Z(
        \MC_ARK_ARC_1_2/temp4[114] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_12_5  ( .A1(\RI5[2][24] ), .A2(\RI5[2][180] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[114] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_12_5  ( .A1(\RI5[2][84] ), .A2(\RI5[2][60] ), .Z(
        \MC_ARK_ARC_1_2/temp2[114] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_12_4  ( .A1(\MC_ARK_ARC_1_2/temp2[115] ), .A2(
        \MC_ARK_ARC_1_2/temp1[115] ), .Z(\MC_ARK_ARC_1_2/temp5[115] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_12_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[151] ), 
        .A2(n73), .Z(\MC_ARK_ARC_1_2/temp4[115] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_12_4  ( .A1(\RI5[2][25] ), .A2(\RI5[2][181] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[115] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_12_4  ( .A1(\RI5[2][85] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[61] ), .Z(\MC_ARK_ARC_1_2/temp2[115] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_12_4  ( .A1(\RI5[2][109] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[115] ), .Z(\MC_ARK_ARC_1_2/temp1[115] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_12_3  ( .A1(\SB2_2_9/buf_output[2] ), .A2(n242), 
        .Z(\MC_ARK_ARC_1_2/temp4[116] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_12_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[153] ), 
        .A2(n79), .Z(\MC_ARK_ARC_1_2/temp4[117] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_12_1  ( .A1(\SB2_2_7/buf_output[4] ), .A2(n101), 
        .Z(\MC_ARK_ARC_1_2/temp4[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_12_1  ( .A1(\RI5[2][112] ), .A2(\RI5[2][118] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_12_0  ( .A1(\RI5[2][155] ), .A2(n557), .Z(
        \MC_ARK_ARC_1_2/temp4[119] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_12_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[29] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[185] ), .Z(
        \MC_ARK_ARC_1_2/temp3[119] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_12_0  ( .A1(\RI5[2][113] ), .A2(\RI5[2][119] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[119] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_11_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[156] ), 
        .A2(n453), .Z(\MC_ARK_ARC_1_2/temp4[120] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_11_4  ( .A1(\RI5[2][157] ), .A2(n482), .Z(
        \MC_ARK_ARC_1_2/temp4[121] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_11_2  ( .A1(\SB2_2_7/buf_output[3] ), .A2(n540), 
        .Z(\MC_ARK_ARC_1_2/temp4[123] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_11_1  ( .A1(\MC_ARK_ARC_1_2/temp3[124] ), .A2(
        \MC_ARK_ARC_1_2/temp4[124] ), .Z(\MC_ARK_ARC_1_2/temp6[124] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_11_1  ( .A1(\RI5[2][160] ), .A2(n565), .Z(
        \MC_ARK_ARC_1_2/temp4[124] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_11_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[124] ), 
        .A2(\RI5[2][118] ), .Z(\MC_ARK_ARC_1_2/temp1[124] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_10_5  ( .A1(\MC_ARK_ARC_1_2/temp6[126] ), .A2(
        \MC_ARK_ARC_1_2/temp5[126] ), .Z(\MC_ARK_ARC_1_2/buf_output[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_10_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[162] ), 
        .A2(n204), .Z(\MC_ARK_ARC_1_2/temp4[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_10_5  ( .A1(\RI5[2][96] ), .A2(\RI5[2][72] ), .Z(
        \MC_ARK_ARC_1_2/temp2[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_10_5  ( .A1(\RI5[2][126] ), .A2(\RI5[2][120] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_10_4  ( .A1(\RI5[2][163] ), .A2(n210), .Z(
        \MC_ARK_ARC_1_2/temp4[127] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_10_4  ( .A1(\RI5[2][121] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[127] ), .Z(\MC_ARK_ARC_1_2/temp1[127] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_10_3  ( .A1(\RI5[2][164] ), .A2(n547), .Z(
        \MC_ARK_ARC_1_2/temp4[128] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_10_3  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[74] ), 
        .A2(\RI5[2][98] ), .Z(\MC_ARK_ARC_1_2/temp2[128] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_10_2  ( .A1(\RI5[2][165] ), .A2(n67), .Z(
        \MC_ARK_ARC_1_2/temp4[129] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_10_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[39] ), 
        .A2(\RI5[2][3] ), .Z(\MC_ARK_ARC_1_2/temp3[129] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_10_1  ( .A1(\RI5[2][166] ), .A2(n471), .Z(
        \MC_ARK_ARC_1_2/temp4[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_10_1  ( .A1(\RI5[2][40] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[4] ), .Z(\MC_ARK_ARC_1_2/temp3[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_10_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[76] ), 
        .A2(\RI5[2][100] ), .Z(\MC_ARK_ARC_1_2/temp2[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_10_1  ( .A1(\RI5[2][130] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[124] ), .Z(\MC_ARK_ARC_1_2/temp1[130] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_10_0  ( .A1(\MC_ARK_ARC_1_2/temp5[131] ), .A2(
        \MC_ARK_ARC_1_2/temp6[131] ), .Z(\MC_ARK_ARC_1_2/buf_output[131] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_10_0  ( .A1(\SB2_2_4/buf_output[5] ), .A2(n501), 
        .Z(\MC_ARK_ARC_1_2/temp4[131] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_9_5  ( .A1(\RI5[2][168] ), .A2(n527), .Z(
        \MC_ARK_ARC_1_2/temp4[132] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_9_5  ( .A1(\RI5[2][42] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[6] ), .Z(\MC_ARK_ARC_1_2/temp3[132] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_9_4  ( .A1(\RI5[2][169] ), .A2(n228), .Z(
        \MC_ARK_ARC_1_2/temp4[133] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_9_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[133] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[127] ), .Z(
        \MC_ARK_ARC_1_2/temp1[133] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_9_3  ( .A1(\RI5[2][170] ), .A2(n451), .Z(
        \MC_ARK_ARC_1_2/temp4[134] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_9_3  ( .A1(\RI5[2][8] ), .A2(\RI5[2][44] ), .Z(
        \MC_ARK_ARC_1_2/temp3[134] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_9_3  ( .A1(\RI5[2][134] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[128] ), .Z(\MC_ARK_ARC_1_2/temp1[134] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_9_2  ( .A1(\MC_ARK_ARC_1_2/temp4[135] ), .A2(
        \MC_ARK_ARC_1_2/temp3[135] ), .Z(\MC_ARK_ARC_1_2/temp6[135] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_9_2  ( .A1(\RI5[2][171] ), .A2(n62), .Z(
        \MC_ARK_ARC_1_2/temp4[135] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_9_1  ( .A1(\MC_ARK_ARC_1_2/temp6[136] ), .A2(
        \MC_ARK_ARC_1_2/temp5[136] ), .Z(\MC_ARK_ARC_1_2/buf_output[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_9_1  ( .A1(\MC_ARK_ARC_1_2/temp3[136] ), .A2(
        \MC_ARK_ARC_1_2/temp4[136] ), .Z(\MC_ARK_ARC_1_2/temp6[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_9_1  ( .A1(\MC_ARK_ARC_1_2/temp1[136] ), .A2(
        \MC_ARK_ARC_1_2/temp2[136] ), .Z(\MC_ARK_ARC_1_2/temp5[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_9_1  ( .A1(\RI5[2][172] ), .A2(n134), .Z(
        \MC_ARK_ARC_1_2/temp4[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_9_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[136] ), 
        .A2(\RI5[2][130] ), .Z(\MC_ARK_ARC_1_2/temp1[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_9_0  ( .A1(\RI5[2][173] ), .A2(n71), .Z(
        \MC_ARK_ARC_1_2/temp4[137] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_9_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[131] ), 
        .A2(\RI5[2][137] ), .Z(\MC_ARK_ARC_1_2/temp1[137] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_8_5  ( .A1(\MC_ARK_ARC_1_2/temp1[138] ), .A2(
        \MC_ARK_ARC_1_2/temp2[138] ), .Z(\MC_ARK_ARC_1_2/temp5[138] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_8_5  ( .A1(\RI5[2][174] ), .A2(n219), .Z(
        \MC_ARK_ARC_1_2/temp4[138] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_8_5  ( .A1(\RI5[2][48] ), .A2(\RI5[2][12] ), .Z(
        \MC_ARK_ARC_1_2/temp3[138] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_8_5  ( .A1(\RI5[2][108] ), .A2(\RI5[2][84] ), .Z(
        \MC_ARK_ARC_1_2/temp2[138] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_8_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[175] ), 
        .A2(n236), .Z(\MC_ARK_ARC_1_2/temp4[139] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_8_4  ( .A1(\RI5[2][13] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[49] ), .Z(\MC_ARK_ARC_1_2/temp3[139] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_8_4  ( .A1(\RI5[2][109] ), .A2(\RI5[2][85] ), .Z(
        \MC_ARK_ARC_1_2/temp2[139] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_8_3  ( .A1(\MC_ARK_ARC_1_2/temp3[140] ), .A2(
        \MC_ARK_ARC_1_2/temp4[140] ), .Z(\MC_ARK_ARC_1_2/temp6[140] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_8_3  ( .A1(\RI5[2][176] ), .A2(n492), .Z(
        \MC_ARK_ARC_1_2/temp4[140] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_8_3  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[50] ), 
        .A2(n570), .Z(\MC_ARK_ARC_1_2/temp3[140] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_8_2  ( .A1(\MC_ARK_ARC_1_2/temp3[141] ), .A2(
        \MC_ARK_ARC_1_2/temp4[141] ), .Z(\MC_ARK_ARC_1_2/temp6[141] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_8_2  ( .A1(\SB2_2_4/buf_output[3] ), .A2(n29), 
        .Z(\MC_ARK_ARC_1_2/temp4[141] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_8_1  ( .A1(\MC_ARK_ARC_1_2/temp1[142] ), .A2(
        \MC_ARK_ARC_1_2/temp2[142] ), .Z(\MC_ARK_ARC_1_2/temp5[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_8_1  ( .A1(\RI5[2][178] ), .A2(n545), .Z(
        \MC_ARK_ARC_1_2/temp4[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_8_1  ( .A1(\RI5[2][88] ), .A2(\RI5[2][112] ), .Z(
        \MC_ARK_ARC_1_2/temp2[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_8_0  ( .A1(\MC_ARK_ARC_1_2/temp4[143] ), .A2(
        \MC_ARK_ARC_1_2/temp3[143] ), .Z(\MC_ARK_ARC_1_2/temp6[143] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_8_0  ( .A1(\RI5[2][179] ), .A2(n46), .Z(
        \MC_ARK_ARC_1_2/temp4[143] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_8_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[53] ), 
        .A2(\RI5[2][17] ), .Z(\MC_ARK_ARC_1_2/temp3[143] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_7_5  ( .A1(\RI5[2][180] ), .A2(n226), .Z(
        \MC_ARK_ARC_1_2/temp4[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_7_5  ( .A1(\RI5[2][90] ), .A2(\RI5[2][114] ), .Z(
        \MC_ARK_ARC_1_2/temp2[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_7_4  ( .A1(\MC_ARK_ARC_1_2/temp3[145] ), .A2(
        \MC_ARK_ARC_1_2/temp4[145] ), .Z(\MC_ARK_ARC_1_2/temp6[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_7_4  ( .A1(\MC_ARK_ARC_1_2/temp1[145] ), .A2(
        \MC_ARK_ARC_1_2/temp2[145] ), .Z(\MC_ARK_ARC_1_2/temp5[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_7_4  ( .A1(\RI5[2][181] ), .A2(n189), .Z(
        \MC_ARK_ARC_1_2/temp4[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_7_4  ( .A1(\RI5[2][55] ), .A2(\RI5[2][19] ), .Z(
        \MC_ARK_ARC_1_2/temp3[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_7_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[115] ), 
        .A2(\RI5[2][91] ), .Z(\MC_ARK_ARC_1_2/temp2[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_7_3  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[182] ), 
        .A2(n526), .Z(\MC_ARK_ARC_1_2/temp4[146] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_7_2  ( .A1(\SB2_2_3/buf_output[3] ), .A2(n555), 
        .Z(\MC_ARK_ARC_1_2/temp4[147] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_7_2  ( .A1(\RI5[2][93] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[117] ), .Z(\MC_ARK_ARC_1_2/temp2[147] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_7_1  ( .A1(\MC_ARK_ARC_1_2/temp3[148] ), .A2(
        \MC_ARK_ARC_1_2/temp4[148] ), .Z(\MC_ARK_ARC_1_2/temp6[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_7_1  ( .A1(\RI5[2][184] ), .A2(n22), .Z(
        \MC_ARK_ARC_1_2/temp4[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_7_1  ( .A1(\RI5[2][118] ), .A2(\RI5[2][94] ), .Z(
        \MC_ARK_ARC_1_2/temp2[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_7_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[148] ), 
        .A2(\RI5[2][142] ), .Z(\MC_ARK_ARC_1_2/temp1[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_7_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[185] ), 
        .A2(n479), .Z(\MC_ARK_ARC_1_2/temp4[149] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_6_5  ( .A1(\MC_ARK_ARC_1_2/temp6[150] ), .A2(
        \MC_ARK_ARC_1_2/temp5[150] ), .Z(\MC_ARK_ARC_1_2/buf_output[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_6_5  ( .A1(\MC_ARK_ARC_1_2/temp4[150] ), .A2(
        \MC_ARK_ARC_1_2/temp3[150] ), .Z(\MC_ARK_ARC_1_2/temp6[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_6_5  ( .A1(\MC_ARK_ARC_1_2/temp1[150] ), .A2(
        \MC_ARK_ARC_1_2/temp2[150] ), .Z(\MC_ARK_ARC_1_2/temp5[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_6_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[186] ), 
        .A2(n508), .Z(\MC_ARK_ARC_1_2/temp4[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_6_5  ( .A1(\RI5[2][60] ), .A2(\RI5[2][24] ), .Z(
        \MC_ARK_ARC_1_2/temp3[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_6_5  ( .A1(\RI5[2][96] ), .A2(\RI5[2][120] ), .Z(
        \MC_ARK_ARC_1_2/temp2[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_6_5  ( .A1(\RI5[2][144] ), .A2(\RI5[2][150] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_6_4  ( .A1(\MC_ARK_ARC_1_2/temp5[151] ), .A2(
        \MC_ARK_ARC_1_2/temp6[151] ), .Z(\MC_ARK_ARC_1_2/buf_output[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_6_4  ( .A1(\MC_ARK_ARC_1_2/temp3[151] ), .A2(
        \MC_ARK_ARC_1_2/temp4[151] ), .Z(\MC_ARK_ARC_1_2/temp6[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_6_4  ( .A1(\MC_ARK_ARC_1_2/temp2[151] ), .A2(
        \MC_ARK_ARC_1_2/temp1[151] ), .Z(\MC_ARK_ARC_1_2/temp5[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_6_4  ( .A1(\RI5[2][187] ), .A2(n234), .Z(
        \MC_ARK_ARC_1_2/temp4[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_6_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[61] ), 
        .A2(\RI5[2][25] ), .Z(\MC_ARK_ARC_1_2/temp3[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_6_4  ( .A1(\RI5[2][121] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[97] ), .Z(\MC_ARK_ARC_1_2/temp2[151] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_6_4  ( .A1(\RI5[2][145] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[151] ), .Z(\MC_ARK_ARC_1_2/temp1[151] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_6_3  ( .A1(\SB2_2_3/buf_output[2] ), .A2(n562), 
        .Z(\MC_ARK_ARC_1_2/temp4[152] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_6_2  ( .A1(n1390), .A2(n133), .Z(
        \MC_ARK_ARC_1_2/temp4[153] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_6_1  ( .A1(\MC_ARK_ARC_1_2/temp1[154] ), .A2(
        \MC_ARK_ARC_1_2/temp2[154] ), .Z(\MC_ARK_ARC_1_2/temp5[154] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_6_1  ( .A1(\RI5[2][190] ), .A2(n81), .Z(
        \MC_ARK_ARC_1_2/temp4[154] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_6_1  ( .A1(\RI5[2][28] ), .A2(\RI5[2][64] ), .Z(
        \MC_ARK_ARC_1_2/temp3[154] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_6_1  ( .A1(\RI5[2][100] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[124] ), .Z(\MC_ARK_ARC_1_2/temp2[154] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_6_1  ( .A1(\RI5[2][154] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[148] ), .Z(\MC_ARK_ARC_1_2/temp1[154] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_6_0  ( .A1(\RI5[2][191] ), .A2(n112), .Z(
        \MC_ARK_ARC_1_2/temp4[155] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_5_5  ( .A1(\MC_ARK_ARC_1_2/temp3[156] ), .A2(
        \MC_ARK_ARC_1_2/temp4[156] ), .Z(\MC_ARK_ARC_1_2/temp6[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_5_5  ( .A1(\SB2_2_4/buf_output[0] ), .A2(n194), 
        .Z(\MC_ARK_ARC_1_2/temp4[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_5_5  ( .A1(\RI5[2][66] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[30] ), .Z(\MC_ARK_ARC_1_2/temp3[156] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_5_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[156] ), 
        .A2(\RI5[2][150] ), .Z(\MC_ARK_ARC_1_2/temp1[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_5_4  ( .A1(\MC_ARK_ARC_1_2/temp2[157] ), .A2(
        \MC_ARK_ARC_1_2/temp1[157] ), .Z(\MC_ARK_ARC_1_2/temp5[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_5_4  ( .A1(\RI5[2][1] ), .A2(n137), .Z(
        \MC_ARK_ARC_1_2/temp4[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_5_4  ( .A1(\SB2_2_18/buf_output[1] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[127] ), .Z(\MC_ARK_ARC_1_2/temp2[157] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_5_4  ( .A1(\RI5[2][157] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[151] ), .Z(\MC_ARK_ARC_1_2/temp1[157] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_5_3  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[2] ), 
        .A2(n469), .Z(\MC_ARK_ARC_1_2/temp4[158] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_5_3  ( .A1(\RI5[2][32] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[68] ), .Z(\MC_ARK_ARC_1_2/temp3[158] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_5_2  ( .A1(\RI5[2][3] ), .A2(n499), .Z(
        \MC_ARK_ARC_1_2/temp4[159] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_5_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[105] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[129] ), .Z(
        \MC_ARK_ARC_1_2/temp2[159] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_5_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[4] ), 
        .A2(n524), .Z(\MC_ARK_ARC_1_2/temp4[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_5_1  ( .A1(\RI5[2][154] ), .A2(\RI5[2][160] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_5_0  ( .A1(\MC_ARK_ARC_1_2/temp6[161] ), .A2(
        \MC_ARK_ARC_1_2/temp5[161] ), .Z(\MC_ARK_ARC_1_2/buf_output[161] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_5_0  ( .A1(\MC_ARK_ARC_1_2/temp3[161] ), .A2(
        \MC_ARK_ARC_1_2/temp4[161] ), .Z(\MC_ARK_ARC_1_2/temp6[161] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_5_0  ( .A1(\RI5[2][5] ), .A2(n554), .Z(
        \MC_ARK_ARC_1_2/temp4[161] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_4_5  ( .A1(\MC_ARK_ARC_1_2/temp5[162] ), .A2(
        \MC_ARK_ARC_1_2/temp6[162] ), .Z(\MC_ARK_ARC_1_2/buf_output[162] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_4_5  ( .A1(\MC_ARK_ARC_1_2/temp4[162] ), .A2(
        \MC_ARK_ARC_1_2/temp3[162] ), .Z(\MC_ARK_ARC_1_2/temp6[162] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_4_5  ( .A1(\MC_ARK_ARC_1_2/temp2[162] ), .A2(
        \MC_ARK_ARC_1_2/temp1[162] ), .Z(\MC_ARK_ARC_1_2/temp5[162] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_4_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[6] ), 
        .A2(n449), .Z(\MC_ARK_ARC_1_2/temp4[162] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_4_5  ( .A1(\RI5[2][72] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[36] ), .Z(\MC_ARK_ARC_1_2/temp3[162] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_4_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[132] ), 
        .A2(\RI5[2][108] ), .Z(\MC_ARK_ARC_1_2/temp2[162] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_4_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[7] ), 
        .A2(n202), .Z(\MC_ARK_ARC_1_2/temp4[163] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_4_4  ( .A1(\RI5[2][163] ), .A2(\RI5[2][157] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[163] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_4_3  ( .A1(\MC_ARK_ARC_1_2/temp2[164] ), .A2(
        \MC_ARK_ARC_1_2/temp1[164] ), .Z(\MC_ARK_ARC_1_2/temp5[164] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_4_3  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[158] ), 
        .A2(\RI5[2][164] ), .Z(\MC_ARK_ARC_1_2/temp1[164] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_4_2  ( .A1(\RI5[2][9] ), .A2(n536), .Z(
        \MC_ARK_ARC_1_2/temp4[165] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_4_2  ( .A1(\RI5[2][159] ), .A2(\RI5[2][165] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[165] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_4_1  ( .A1(\MC_ARK_ARC_1_2/temp3[166] ), .A2(
        \MC_ARK_ARC_1_2/temp4[166] ), .Z(\MC_ARK_ARC_1_2/temp6[166] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_4_1  ( .A1(\SB2_2_31/buf_output[4] ), .A2(n201), 
        .Z(\MC_ARK_ARC_1_2/temp4[166] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_4_0  ( .A1(\RI5[2][137] ), .A2(\RI5[2][113] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[167] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_4_0  ( .A1(\RI5[2][167] ), .A2(\RI5[2][161] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[167] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_3_5  ( .A1(\MC_ARK_ARC_1_2/temp3[168] ), .A2(
        \MC_ARK_ARC_1_2/temp4[168] ), .Z(\MC_ARK_ARC_1_2/temp6[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_3_5  ( .A1(\RI5[2][12] ), .A2(n488), .Z(
        \MC_ARK_ARC_1_2/temp4[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_3_5  ( .A1(\RI5[2][42] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[78] ), .Z(\MC_ARK_ARC_1_2/temp3[168] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_3_4  ( .A1(\MC_ARK_ARC_1_2/temp3[169] ), .A2(
        \MC_ARK_ARC_1_2/temp4[169] ), .Z(\MC_ARK_ARC_1_2/temp6[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_3_4  ( .A1(\RI5[2][13] ), .A2(n172), .Z(
        \MC_ARK_ARC_1_2/temp4[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_3_4  ( .A1(\RI5[2][79] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[43] ), .Z(\MC_ARK_ARC_1_2/temp3[169] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_3_4  ( .A1(\RI5[2][139] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[115] ), .Z(\MC_ARK_ARC_1_2/temp2[169] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_3_4  ( .A1(\RI5[2][163] ), .A2(\RI5[2][169] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_3_3  ( .A1(\RI5[2][140] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[116] ), .Z(\MC_ARK_ARC_1_2/temp2[170] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_3_2  ( .A1(\RI5[2][15] ), .A2(n440), .Z(
        \MC_ARK_ARC_1_2/temp4[171] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_3_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[81] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[45] ), .Z(
        \MC_ARK_ARC_1_2/temp3[171] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_3_2  ( .A1(\RI5[2][165] ), .A2(\RI5[2][171] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[171] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_3_1  ( .A1(\MC_ARK_ARC_1_2/temp3[172] ), .A2(
        \MC_ARK_ARC_1_2/temp4[172] ), .Z(\MC_ARK_ARC_1_2/temp6[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_3_1  ( .A1(\MC_ARK_ARC_1_2/temp1[172] ), .A2(
        \MC_ARK_ARC_1_2/temp2[172] ), .Z(\MC_ARK_ARC_1_2/temp5[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_3_1  ( .A1(\RI5[2][16] ), .A2(n20), .Z(
        \MC_ARK_ARC_1_2/temp4[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_3_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[82] ), 
        .A2(\RI5[2][46] ), .Z(\MC_ARK_ARC_1_2/temp3[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_3_1  ( .A1(\RI5[2][118] ), .A2(\RI5[2][142] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_3_1  ( .A1(\RI5[2][172] ), .A2(\RI5[2][166] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_3_0  ( .A1(\RI5[2][17] ), .A2(n498), .Z(
        \MC_ARK_ARC_1_2/temp4[173] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_3_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[47] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[83] ), .Z(
        \MC_ARK_ARC_1_2/temp3[173] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_2_5  ( .A1(\MC_ARK_ARC_1_2/temp5[174] ), .A2(
        \MC_ARK_ARC_1_2/temp6[174] ), .Z(\MC_ARK_ARC_1_2/buf_output[174] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_2_5  ( .A1(\MC_ARK_ARC_1_2/temp3[174] ), .A2(
        \MC_ARK_ARC_1_2/temp4[174] ), .Z(\MC_ARK_ARC_1_2/temp6[174] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_2_5  ( .A1(\RI5[2][18] ), .A2(n212), .Z(
        \MC_ARK_ARC_1_2/temp4[174] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_2_4  ( .A1(\RI5[2][19] ), .A2(n230), .Z(
        \MC_ARK_ARC_1_2/temp4[175] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_2_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[49] ), 
        .A2(\RI5[2][85] ), .Z(\MC_ARK_ARC_1_2/temp3[175] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_2_3  ( .A1(\RI5[2][20] ), .A2(n220), .Z(
        \MC_ARK_ARC_1_2/temp4[176] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_2_3  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[146] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[122] ), .Z(
        \MC_ARK_ARC_1_2/temp2[176] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_2_3  ( .A1(\RI5[2][176] ), .A2(\RI5[2][170] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[176] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_2_2  ( .A1(\RI5[2][21] ), .A2(n105), .Z(
        \MC_ARK_ARC_1_2/temp4[177] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_2_2  ( .A1(\RI5[2][51] ), .A2(\RI5[2][87] ), .Z(
        \MC_ARK_ARC_1_2/temp3[177] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_2_1  ( .A1(\MC_ARK_ARC_1_2/temp3[178] ), .A2(
        \MC_ARK_ARC_1_2/temp4[178] ), .Z(\MC_ARK_ARC_1_2/temp6[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_2_1  ( .A1(\MC_ARK_ARC_1_2/temp2[178] ), .A2(
        \MC_ARK_ARC_1_2/temp1[178] ), .Z(\MC_ARK_ARC_1_2/temp5[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_2_1  ( .A1(\RI5[2][22] ), .A2(n96), .Z(
        \MC_ARK_ARC_1_2/temp4[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_2_1  ( .A1(\RI5[2][88] ), .A2(\RI5[2][52] ), .Z(
        \MC_ARK_ARC_1_2/temp3[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_2_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[124] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[148] ), .Z(
        \MC_ARK_ARC_1_2/temp2[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_2_1  ( .A1(\RI5[2][178] ), .A2(\RI5[2][172] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_2_0  ( .A1(\RI5[2][23] ), .A2(n534), .Z(
        \MC_ARK_ARC_1_2/temp4[179] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_2_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[125] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[149] ), .Z(
        \MC_ARK_ARC_1_2/temp2[179] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_1_5  ( .A1(\RI5[2][24] ), .A2(n196), .Z(
        \MC_ARK_ARC_1_2/temp4[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_1_5  ( .A1(\RI5[2][54] ), .A2(\RI5[2][90] ), .Z(
        \MC_ARK_ARC_1_2/temp3[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_1_5  ( .A1(\RI5[2][150] ), .A2(\RI5[2][126] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_1_5  ( .A1(\RI5[2][180] ), .A2(\RI5[2][174] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_1_4  ( .A1(\MC_ARK_ARC_1_2/temp5[181] ), .A2(
        \MC_ARK_ARC_1_2/temp6[181] ), .Z(\MC_ARK_ARC_1_2/buf_output[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_1_4  ( .A1(\MC_ARK_ARC_1_2/temp3[181] ), .A2(
        \MC_ARK_ARC_1_2/temp4[181] ), .Z(\MC_ARK_ARC_1_2/temp6[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_1_4  ( .A1(\MC_ARK_ARC_1_2/temp1[181] ), .A2(
        \MC_ARK_ARC_1_2/temp2[181] ), .Z(\MC_ARK_ARC_1_2/temp5[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_1_4  ( .A1(\RI5[2][25] ), .A2(n458), .Z(
        \MC_ARK_ARC_1_2/temp4[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_1_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[151] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[127] ), .Z(
        \MC_ARK_ARC_1_2/temp2[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_1_4  ( .A1(\RI5[2][181] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[175] ), .Z(\MC_ARK_ARC_1_2/temp1[181] )
         );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_1_3  ( .A1(n3677), .A2(n237), .Z(
        \MC_ARK_ARC_1_2/temp4[182] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_1_3  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[56] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[92] ), .Z(
        \MC_ARK_ARC_1_2/temp3[182] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_1_2  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[27] ), 
        .A2(n515), .Z(\MC_ARK_ARC_1_2/temp4[183] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_1_1  ( .A1(\MC_ARK_ARC_1_2/temp6[184] ), .A2(
        \MC_ARK_ARC_1_2/temp5[184] ), .Z(\MC_ARK_ARC_1_2/buf_output[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_1_1  ( .A1(\MC_ARK_ARC_1_2/temp4[184] ), .A2(
        \MC_ARK_ARC_1_2/temp3[184] ), .Z(\MC_ARK_ARC_1_2/temp6[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_1_1  ( .A1(\RI5[2][28] ), .A2(n40), .Z(
        \MC_ARK_ARC_1_2/temp4[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_1_1  ( .A1(\RI5[2][154] ), .A2(\RI5[2][130] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_1_0  ( .A1(\MC_ARK_ARC_1_2/temp4[185] ), .A2(
        \MC_ARK_ARC_1_2/temp3[185] ), .Z(\MC_ARK_ARC_1_2/temp6[185] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_1_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[29] ), 
        .A2(n223), .Z(\MC_ARK_ARC_1_2/temp4[185] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_0_5  ( .A1(\MC_ARK_ARC_1_2/temp5[186] ), .A2(
        \MC_ARK_ARC_1_2/temp6[186] ), .Z(\MC_ARK_ARC_1_2/buf_output[186] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_0_5  ( .A1(\MC_ARK_ARC_1_2/temp4[186] ), .A2(
        \MC_ARK_ARC_1_2/temp3[186] ), .Z(\MC_ARK_ARC_1_2/temp6[186] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_0_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[30] ), 
        .A2(n216), .Z(\MC_ARK_ARC_1_2/temp4[186] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_0_5  ( .A1(\RI5[2][96] ), .A2(\RI5[2][60] ), .Z(
        \MC_ARK_ARC_1_2/temp3[186] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_0_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[156] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[132] ), .Z(
        \MC_ARK_ARC_1_2/temp2[186] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_0_5  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[186] ), 
        .A2(\RI5[2][180] ), .Z(\MC_ARK_ARC_1_2/temp1[186] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X7_0_4  ( .A1(\MC_ARK_ARC_1_2/temp5[187] ), .A2(
        \MC_ARK_ARC_1_2/temp6[187] ), .Z(\MC_ARK_ARC_1_2/buf_output[187] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_0_4  ( .A1(\MC_ARK_ARC_1_2/temp3[187] ), .A2(
        \MC_ARK_ARC_1_2/temp4[187] ), .Z(\MC_ARK_ARC_1_2/temp6[187] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_0_4  ( .A1(\RI5[2][31] ), .A2(n188), .Z(
        \MC_ARK_ARC_1_2/temp4[187] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_0_4  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[97] ), 
        .A2(\MC_ARK_ARC_1_2/buf_datainput[61] ), .Z(
        \MC_ARK_ARC_1_2/temp3[187] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_0_4  ( .A1(\RI5[2][181] ), .A2(\RI5[2][187] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[187] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_0_3  ( .A1(\RI5[2][32] ), .A2(n156), .Z(
        \MC_ARK_ARC_1_2/temp4[188] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_0_2  ( .A1(\RI5[2][33] ), .A2(n173), .Z(
        \MC_ARK_ARC_1_2/temp4[189] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X5_0_1  ( .A1(\MC_ARK_ARC_1_2/temp2[190] ), .A2(
        \MC_ARK_ARC_1_2/temp1[190] ), .Z(\MC_ARK_ARC_1_2/temp5[190] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_0_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[34] ), 
        .A2(n447), .Z(\MC_ARK_ARC_1_2/temp4[190] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_0_1  ( .A1(\RI5[2][64] ), .A2(\RI5[2][100] ), .Z(
        \MC_ARK_ARC_1_2/temp3[190] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_0_1  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[136] ), 
        .A2(\RI5[2][160] ), .Z(\MC_ARK_ARC_1_2/temp2[190] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X1_0_1  ( .A1(\RI5[2][184] ), .A2(\RI5[2][190] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[190] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X6_0_0  ( .A1(\MC_ARK_ARC_1_2/temp3[191] ), .A2(
        \MC_ARK_ARC_1_2/temp4[191] ), .Z(\MC_ARK_ARC_1_2/temp6[191] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X4_0_0  ( .A1(\RI5[2][35] ), .A2(n474), .Z(
        \MC_ARK_ARC_1_2/temp4[191] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X3_0_0  ( .A1(\MC_ARK_ARC_1_2/buf_datainput[65] ), 
        .A2(\RI5[2][101] ), .Z(\MC_ARK_ARC_1_2/temp3[191] ) );
  XOR2_X1 \MC_ARK_ARC_1_2/X2_0_0  ( .A1(\RI5[2][161] ), .A2(\RI5[2][137] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[191] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_95  ( .I(\SB2_2_16/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[95] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_61  ( .I(\SB2_2_25/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[61] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_53  ( .I(\SB2_2_23/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[53] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_31_5  ( .A1(\MC_ARK_ARC_1_3/temp3[0] ), .A2(
        \MC_ARK_ARC_1_3/temp4[0] ), .Z(\MC_ARK_ARC_1_3/temp6[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_31_5  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[36] ), 
        .A2(n193), .Z(\MC_ARK_ARC_1_3/temp4[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_31_5  ( .A1(\RI5[3][162] ), .A2(\RI5[3][138] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[0] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_31_4  ( .A1(\MC_ARK_ARC_1_3/temp3[1] ), .A2(
        \MC_ARK_ARC_1_3/temp4[1] ), .Z(\MC_ARK_ARC_1_3/temp6[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_31_4  ( .A1(\RI5[3][37] ), .A2(n445), .Z(
        \MC_ARK_ARC_1_3/temp4[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_31_4  ( .A1(\RI5[3][163] ), .A2(\RI5[3][139] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[1] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_31_3  ( .A1(\MC_ARK_ARC_1_3/temp3[2] ), .A2(
        \MC_ARK_ARC_1_3/temp4[2] ), .Z(\MC_ARK_ARC_1_3/temp6[2] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_31_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[38] ), 
        .A2(n512), .Z(\MC_ARK_ARC_1_3/temp4[2] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_31_3  ( .A1(\RI5[3][68] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[104] ), .Z(\MC_ARK_ARC_1_3/temp3[2] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_31_3  ( .A1(\RI5[3][164] ), .A2(\RI5[3][140] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[2] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_31_3  ( .A1(\RI5[3][188] ), .A2(\RI5[3][2] ), .Z(
        \MC_ARK_ARC_1_3/temp1[2] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_31_2  ( .A1(\MC_ARK_ARC_1_3/temp5[3] ), .A2(
        \MC_ARK_ARC_1_3/temp6[3] ), .Z(\MC_ARK_ARC_1_3/buf_output[3] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_31_2  ( .A1(\SB2_3_27/buf_output[3] ), .A2(n238), 
        .Z(\MC_ARK_ARC_1_3/temp4[3] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_31_2  ( .A1(\RI5[3][141] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[165] ), .Z(\MC_ARK_ARC_1_3/temp2[3] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_31_1  ( .A1(\MC_ARK_ARC_1_3/temp5[4] ), .A2(
        \MC_ARK_ARC_1_3/temp6[4] ), .Z(\MC_ARK_ARC_1_3/buf_output[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_31_1  ( .A1(\MC_ARK_ARC_1_3/temp3[4] ), .A2(
        \MC_ARK_ARC_1_3/temp4[4] ), .Z(\MC_ARK_ARC_1_3/temp6[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_31_1  ( .A1(\MC_ARK_ARC_1_3/temp2[4] ), .A2(
        \MC_ARK_ARC_1_3/temp1[4] ), .Z(\MC_ARK_ARC_1_3/temp5[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_31_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[40] ), 
        .A2(n510), .Z(\MC_ARK_ARC_1_3/temp4[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_31_1  ( .A1(\RI5[3][106] ), .A2(\RI5[3][70] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_31_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[166] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[142] ), .Z(\MC_ARK_ARC_1_3/temp2[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_31_1  ( .A1(\RI5[3][4] ), .A2(\RI5[3][190] ), .Z(
        \MC_ARK_ARC_1_3/temp1[4] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_31_0  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[41] ), 
        .A2(n60), .Z(\MC_ARK_ARC_1_3/temp4[5] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_31_0  ( .A1(\RI5[3][107] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[71] ), .Z(\MC_ARK_ARC_1_3/temp3[5] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_30_5  ( .A1(\RI5[3][42] ), .A2(n126), .Z(
        \MC_ARK_ARC_1_3/temp4[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_30_5  ( .A1(\RI5[3][108] ), .A2(\RI5[3][72] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_30_5  ( .A1(\RI5[3][0] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[6] ), .Z(\MC_ARK_ARC_1_3/temp1[6] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_30_4  ( .A1(\RI5[3][43] ), .A2(n8), .Z(
        \MC_ARK_ARC_1_3/temp4[7] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_30_4  ( .A1(\RI5[3][73] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[109] ), .Z(\MC_ARK_ARC_1_3/temp3[7] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_30_4  ( .A1(\RI5[3][7] ), .A2(\RI5[3][1] ), .Z(
        \MC_ARK_ARC_1_3/temp1[7] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_30_3  ( .A1(\SB2_3_27/buf_output[2] ), .A2(n163), 
        .Z(\MC_ARK_ARC_1_3/temp4[8] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_30_2  ( .A1(\MC_ARK_ARC_1_3/temp2[9] ), .A2(
        \MC_ARK_ARC_1_3/temp1[9] ), .Z(\MC_ARK_ARC_1_3/temp5[9] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_30_2  ( .A1(\RI5[3][45] ), .A2(n441), .Z(
        \MC_ARK_ARC_1_3/temp4[9] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_30_2  ( .A1(\RI5[3][75] ), .A2(n1392), .Z(
        \MC_ARK_ARC_1_3/temp3[9] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_30_2  ( .A1(\RI5[3][147] ), .A2(\RI5[3][171] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[9] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_30_2  ( .A1(\RI5[3][3] ), .A2(\RI5[3][9] ), .Z(
        \MC_ARK_ARC_1_3/temp1[9] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_30_1  ( .A1(\RI5[3][46] ), .A2(n506), .Z(
        \MC_ARK_ARC_1_3/temp4[10] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_30_0  ( .A1(\RI5[3][47] ), .A2(n439), .Z(
        \MC_ARK_ARC_1_3/temp4[11] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_29_5  ( .A1(\MC_ARK_ARC_1_3/temp3[12] ), .A2(
        \MC_ARK_ARC_1_3/temp4[12] ), .Z(\MC_ARK_ARC_1_3/temp6[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_29_5  ( .A1(\RI5[3][48] ), .A2(n505), .Z(
        \MC_ARK_ARC_1_3/temp4[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_29_5  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[114] ), 
        .A2(\RI5[3][78] ), .Z(\MC_ARK_ARC_1_3/temp3[12] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_29_5  ( .A1(\RI5[3][150] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[174] ), .Z(\MC_ARK_ARC_1_3/temp2[12] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_29_5  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[12] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[6] ), .Z(\MC_ARK_ARC_1_3/temp1[12] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_29_4  ( .A1(\MC_ARK_ARC_1_3/temp5[13] ), .A2(
        \MC_ARK_ARC_1_3/temp6[13] ), .Z(\MC_ARK_ARC_1_3/buf_output[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_29_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[49] ), 
        .A2(n438), .Z(\MC_ARK_ARC_1_3/temp4[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_29_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[115] ), 
        .A2(\RI5[3][79] ), .Z(\MC_ARK_ARC_1_3/temp3[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_29_4  ( .A1(\RI5[3][175] ), .A2(\RI5[3][151] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_29_4  ( .A1(\RI5[3][13] ), .A2(\RI5[3][7] ), .Z(
        \MC_ARK_ARC_1_3/temp1[13] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_29_3  ( .A1(\RI5[3][50] ), .A2(n503), .Z(
        \MC_ARK_ARC_1_3/temp4[14] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_29_3  ( .A1(\RI5[3][80] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[116] ), .Z(\MC_ARK_ARC_1_3/temp3[14] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_29_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[152] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[176] ), .Z(
        \MC_ARK_ARC_1_3/temp2[14] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_29_2  ( .A1(\MC_ARK_ARC_1_3/temp5[15] ), .A2(
        \MC_ARK_ARC_1_3/temp6[15] ), .Z(\MC_ARK_ARC_1_3/buf_output[15] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_29_2  ( .A1(\MC_ARK_ARC_1_3/temp3[15] ), .A2(
        \MC_ARK_ARC_1_3/temp4[15] ), .Z(\MC_ARK_ARC_1_3/temp6[15] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_29_2  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[51] ), 
        .A2(n241), .Z(\MC_ARK_ARC_1_3/temp4[15] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_29_2  ( .A1(\RI5[3][117] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[81] ), .Z(\MC_ARK_ARC_1_3/temp3[15] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_29_2  ( .A1(\RI5[3][177] ), .A2(\RI5[3][153] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[15] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_29_2  ( .A1(\RI5[3][15] ), .A2(\RI5[3][9] ), .Z(
        \MC_ARK_ARC_1_3/temp1[15] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_29_1  ( .A1(\MC_ARK_ARC_1_3/temp3[16] ), .A2(
        \MC_ARK_ARC_1_3/temp4[16] ), .Z(\MC_ARK_ARC_1_3/temp6[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_29_1  ( .A1(\RI5[3][52] ), .A2(n79), .Z(
        \MC_ARK_ARC_1_3/temp4[16] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_29_0  ( .A1(\MC_ARK_ARC_1_3/temp3[17] ), .A2(
        \MC_ARK_ARC_1_3/temp4[17] ), .Z(\MC_ARK_ARC_1_3/temp6[17] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_29_0  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[53] ), 
        .A2(n565), .Z(\MC_ARK_ARC_1_3/temp4[17] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_29_0  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[119] ), 
        .A2(\RI5[3][83] ), .Z(\MC_ARK_ARC_1_3/temp3[17] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_28_5  ( .A1(\MC_ARK_ARC_1_3/temp5[18] ), .A2(
        \MC_ARK_ARC_1_3/temp6[18] ), .Z(\MC_ARK_ARC_1_3/buf_output[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_28_5  ( .A1(\MC_ARK_ARC_1_3/temp2[18] ), .A2(
        \MC_ARK_ARC_1_3/temp1[18] ), .Z(\MC_ARK_ARC_1_3/temp5[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_28_5  ( .A1(\RI5[3][54] ), .A2(n501), .Z(
        \MC_ARK_ARC_1_3/temp4[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_28_5  ( .A1(\RI5[3][120] ), .A2(\RI5[3][84] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_28_5  ( .A1(\RI5[3][180] ), .A2(\RI5[3][156] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_28_5  ( .A1(\RI5[3][18] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[12] ), .Z(\MC_ARK_ARC_1_3/temp1[18] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_28_4  ( .A1(\MC_ARK_ARC_1_3/temp2[19] ), .A2(
        \MC_ARK_ARC_1_3/temp1[19] ), .Z(\MC_ARK_ARC_1_3/temp5[19] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_28_4  ( .A1(\RI5[3][55] ), .A2(n219), .Z(
        \MC_ARK_ARC_1_3/temp4[19] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_28_4  ( .A1(\RI5[3][121] ), .A2(\RI5[3][85] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[19] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_28_4  ( .A1(\RI5[3][157] ), .A2(\RI5[3][181] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[19] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_28_4  ( .A1(\RI5[3][19] ), .A2(\RI5[3][13] ), .Z(
        \MC_ARK_ARC_1_3/temp1[19] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_28_3  ( .A1(\MC_ARK_ARC_1_3/temp5[20] ), .A2(
        \MC_ARK_ARC_1_3/temp6[20] ), .Z(\MC_ARK_ARC_1_3/buf_output[20] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_28_3  ( .A1(\MC_ARK_ARC_1_3/temp3[20] ), .A2(
        \MC_ARK_ARC_1_3/temp4[20] ), .Z(\MC_ARK_ARC_1_3/temp6[20] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_28_3  ( .A1(\MC_ARK_ARC_1_3/temp1[20] ), .A2(
        \MC_ARK_ARC_1_3/temp2[20] ), .Z(\MC_ARK_ARC_1_3/temp5[20] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_28_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[56] ), 
        .A2(n189), .Z(\MC_ARK_ARC_1_3/temp4[20] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_28_3  ( .A1(\RI5[3][86] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[122] ), .Z(\MC_ARK_ARC_1_3/temp3[20] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_28_3  ( .A1(\RI5[3][20] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[14] ), .Z(\MC_ARK_ARC_1_3/temp1[20] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_28_2  ( .A1(\MC_ARK_ARC_1_3/temp3[21] ), .A2(
        \MC_ARK_ARC_1_3/temp4[21] ), .Z(\MC_ARK_ARC_1_3/temp6[21] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_28_2  ( .A1(\MC_ARK_ARC_1_3/temp2[21] ), .A2(
        \MC_ARK_ARC_1_3/temp1[21] ), .Z(\MC_ARK_ARC_1_3/temp5[21] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_28_2  ( .A1(\RI5[3][57] ), .A2(n562), .Z(
        \MC_ARK_ARC_1_3/temp4[21] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_28_2  ( .A1(\RI5[3][87] ), .A2(n3658), .Z(
        \MC_ARK_ARC_1_3/temp3[21] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_28_2  ( .A1(\RI5[3][159] ), .A2(\RI5[3][183] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[21] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_28_2  ( .A1(\RI5[3][15] ), .A2(\RI5[3][21] ), .Z(
        \MC_ARK_ARC_1_3/temp1[21] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_28_1  ( .A1(\MC_ARK_ARC_1_3/temp2[22] ), .A2(
        \MC_ARK_ARC_1_3/temp1[22] ), .Z(\MC_ARK_ARC_1_3/temp5[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_28_1  ( .A1(\RI5[3][58] ), .A2(n28), .Z(
        \MC_ARK_ARC_1_3/temp4[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_28_1  ( .A1(\RI5[3][124] ), .A2(\RI5[3][88] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_28_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[22] ), 
        .A2(\RI5[3][16] ), .Z(\MC_ARK_ARC_1_3/temp1[22] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_28_0  ( .A1(\RI5[3][59] ), .A2(n201), .Z(
        \MC_ARK_ARC_1_3/temp4[23] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_27_5  ( .A1(\MC_ARK_ARC_1_3/temp5[24] ), .A2(
        \MC_ARK_ARC_1_3/temp6[24] ), .Z(\MC_ARK_ARC_1_3/buf_output[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_27_5  ( .A1(\MC_ARK_ARC_1_3/temp3[24] ), .A2(
        \MC_ARK_ARC_1_3/temp4[24] ), .Z(\MC_ARK_ARC_1_3/temp6[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_27_5  ( .A1(\MC_ARK_ARC_1_3/temp2[24] ), .A2(
        \MC_ARK_ARC_1_3/temp1[24] ), .Z(\MC_ARK_ARC_1_3/temp5[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_27_5  ( .A1(\RI5[3][60] ), .A2(n192), .Z(
        \MC_ARK_ARC_1_3/temp4[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_27_5  ( .A1(n2896), .A2(\RI5[3][126] ), .Z(
        \MC_ARK_ARC_1_3/temp3[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_27_5  ( .A1(\RI5[3][24] ), .A2(\RI5[3][18] ), .Z(
        \MC_ARK_ARC_1_3/temp1[24] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_27_4  ( .A1(\MC_ARK_ARC_1_3/temp2[25] ), .A2(
        \MC_ARK_ARC_1_3/temp1[25] ), .Z(\MC_ARK_ARC_1_3/temp5[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_27_4  ( .A1(\RI5[3][61] ), .A2(n174), .Z(
        \MC_ARK_ARC_1_3/temp4[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_27_4  ( .A1(\RI5[3][187] ), .A2(\RI5[3][163] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_27_4  ( .A1(\RI5[3][19] ), .A2(\RI5[3][25] ), .Z(
        \MC_ARK_ARC_1_3/temp1[25] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_27_2  ( .A1(\MC_ARK_ARC_1_3/temp5[27] ), .A2(
        \MC_ARK_ARC_1_3/temp6[27] ), .Z(\MC_ARK_ARC_1_3/buf_output[27] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_27_2  ( .A1(\RI5[3][63] ), .A2(n559), .Z(
        \MC_ARK_ARC_1_3/temp4[27] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_27_2  ( .A1(\RI5[3][21] ), .A2(\RI5[3][27] ), .Z(
        \MC_ARK_ARC_1_3/temp1[27] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_27_1  ( .A1(\MC_ARK_ARC_1_3/temp2[28] ), .A2(
        \MC_ARK_ARC_1_3/temp1[28] ), .Z(\MC_ARK_ARC_1_3/temp5[28] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_27_1  ( .A1(\RI5[3][64] ), .A2(n6), .Z(
        \MC_ARK_ARC_1_3/temp4[28] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_27_1  ( .A1(\RI5[3][130] ), .A2(\RI5[3][94] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[28] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_27_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[28] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[22] ), .Z(\MC_ARK_ARC_1_3/temp1[28] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_27_0  ( .A1(\RI5[3][65] ), .A2(n558), .Z(
        \MC_ARK_ARC_1_3/temp4[29] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_27_0  ( .A1(\RI5[3][29] ), .A2(\RI5[3][23] ), .Z(
        \MC_ARK_ARC_1_3/temp1[29] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_26_5  ( .A1(\MC_ARK_ARC_1_3/temp5[30] ), .A2(
        \MC_ARK_ARC_1_3/temp6[30] ), .Z(\MC_ARK_ARC_1_3/buf_output[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_26_5  ( .A1(\MC_ARK_ARC_1_3/temp3[30] ), .A2(
        \MC_ARK_ARC_1_3/temp4[30] ), .Z(\MC_ARK_ARC_1_3/temp6[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_26_5  ( .A1(\MC_ARK_ARC_1_3/temp2[30] ), .A2(
        \MC_ARK_ARC_1_3/temp1[30] ), .Z(\MC_ARK_ARC_1_3/temp5[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_26_5  ( .A1(\RI5[3][66] ), .A2(n78), .Z(
        \MC_ARK_ARC_1_3/temp4[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_26_5  ( .A1(\RI5[3][96] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[132] ), .Z(\MC_ARK_ARC_1_3/temp3[30] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_26_5  ( .A1(\RI5[3][0] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[168] ), .Z(\MC_ARK_ARC_1_3/temp2[30] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_26_5  ( .A1(\RI5[3][30] ), .A2(\RI5[3][24] ), .Z(
        \MC_ARK_ARC_1_3/temp1[30] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_26_4  ( .A1(\RI5[3][67] ), .A2(n208), .Z(
        \MC_ARK_ARC_1_3/temp4[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_26_4  ( .A1(\RI5[3][133] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[97] ), .Z(\MC_ARK_ARC_1_3/temp3[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_26_4  ( .A1(\RI5[3][31] ), .A2(\RI5[3][25] ), .Z(
        \MC_ARK_ARC_1_3/temp1[31] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_26_3  ( .A1(\RI5[3][68] ), .A2(n493), .Z(
        \MC_ARK_ARC_1_3/temp4[32] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_26_3  ( .A1(\RI5[3][32] ), .A2(\RI5[3][26] ), .Z(
        \MC_ARK_ARC_1_3/temp1[32] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_26_2  ( .A1(\MC_ARK_ARC_1_3/temp1[33] ), .A2(
        \MC_ARK_ARC_1_3/temp2[33] ), .Z(\MC_ARK_ARC_1_3/temp5[33] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_26_2  ( .A1(\RI5[3][69] ), .A2(n232), .Z(
        \MC_ARK_ARC_1_3/temp4[33] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_26_2  ( .A1(\RI5[3][33] ), .A2(\RI5[3][27] ), .Z(
        \MC_ARK_ARC_1_3/temp1[33] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_26_1  ( .A1(\MC_ARK_ARC_1_3/temp5[34] ), .A2(
        \MC_ARK_ARC_1_3/temp6[34] ), .Z(\MC_ARK_ARC_1_3/buf_output[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_26_1  ( .A1(\MC_ARK_ARC_1_3/temp3[34] ), .A2(
        \MC_ARK_ARC_1_3/temp4[34] ), .Z(\MC_ARK_ARC_1_3/temp6[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_26_1  ( .A1(\MC_ARK_ARC_1_3/temp1[34] ), .A2(
        \MC_ARK_ARC_1_3/temp2[34] ), .Z(\MC_ARK_ARC_1_3/temp5[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_26_1  ( .A1(\RI5[3][70] ), .A2(n491), .Z(
        \MC_ARK_ARC_1_3/temp4[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_26_1  ( .A1(\RI5[3][136] ), .A2(\RI5[3][100] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_26_1  ( .A1(\RI5[3][4] ), .A2(\RI5[3][172] ), .Z(
        \MC_ARK_ARC_1_3/temp2[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_26_1  ( .A1(\RI5[3][34] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[28] ), .Z(\MC_ARK_ARC_1_3/temp1[34] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_26_0  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[71] ), 
        .A2(n164), .Z(\MC_ARK_ARC_1_3/temp4[35] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_26_0  ( .A1(\RI5[3][29] ), .A2(\RI5[3][35] ), .Z(
        \MC_ARK_ARC_1_3/temp1[35] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_25_5  ( .A1(\MC_ARK_ARC_1_3/temp6[36] ), .A2(
        \MC_ARK_ARC_1_3/temp5[36] ), .Z(\MC_ARK_ARC_1_3/buf_output[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_25_5  ( .A1(\MC_ARK_ARC_1_3/temp2[36] ), .A2(
        \MC_ARK_ARC_1_3/temp1[36] ), .Z(\MC_ARK_ARC_1_3/temp5[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_25_5  ( .A1(\RI5[3][72] ), .A2(n144), .Z(
        \MC_ARK_ARC_1_3/temp4[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_25_5  ( .A1(\RI5[3][138] ), .A2(\RI5[3][102] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_25_5  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[174] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[6] ), .Z(\MC_ARK_ARC_1_3/temp2[36] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_25_5  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[36] ), 
        .A2(\RI5[3][30] ), .Z(\MC_ARK_ARC_1_3/temp1[36] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_25_4  ( .A1(\MC_ARK_ARC_1_3/temp2[37] ), .A2(
        \MC_ARK_ARC_1_3/temp1[37] ), .Z(\MC_ARK_ARC_1_3/temp5[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_25_4  ( .A1(\RI5[3][73] ), .A2(n553), .Z(
        \MC_ARK_ARC_1_3/temp4[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_25_4  ( .A1(\RI5[3][139] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[103] ), .Z(\MC_ARK_ARC_1_3/temp3[37] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_25_4  ( .A1(\RI5[3][7] ), .A2(\RI5[3][175] ), .Z(
        \MC_ARK_ARC_1_3/temp2[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_25_4  ( .A1(\RI5[3][31] ), .A2(\RI5[3][37] ), .Z(
        \MC_ARK_ARC_1_3/temp1[37] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_25_3  ( .A1(\MC_ARK_ARC_1_3/temp5[38] ), .A2(
        \MC_ARK_ARC_1_3/temp6[38] ), .Z(\MC_ARK_ARC_1_3/buf_output[38] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_25_3  ( .A1(\MC_ARK_ARC_1_3/temp3[38] ), .A2(
        \MC_ARK_ARC_1_3/temp4[38] ), .Z(\MC_ARK_ARC_1_3/temp6[38] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_25_3  ( .A1(\MC_ARK_ARC_1_3/temp2[38] ), .A2(
        \MC_ARK_ARC_1_3/temp1[38] ), .Z(\MC_ARK_ARC_1_3/temp5[38] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_25_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[74] ), 
        .A2(n487), .Z(\MC_ARK_ARC_1_3/temp4[38] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_25_3  ( .A1(\RI5[3][32] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[38] ), .Z(\MC_ARK_ARC_1_3/temp1[38] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_25_2  ( .A1(\RI5[3][75] ), .A2(n552), .Z(
        \MC_ARK_ARC_1_3/temp4[39] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_25_2  ( .A1(\RI5[3][141] ), .A2(\RI5[3][105] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[39] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_25_2  ( .A1(\RI5[3][177] ), .A2(\RI5[3][9] ), .Z(
        \MC_ARK_ARC_1_3/temp2[39] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_25_1  ( .A1(\MC_ARK_ARC_1_3/temp5[40] ), .A2(
        \MC_ARK_ARC_1_3/temp6[40] ), .Z(\MC_ARK_ARC_1_3/buf_output[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_25_1  ( .A1(\MC_ARK_ARC_1_3/temp3[40] ), .A2(
        \MC_ARK_ARC_1_3/temp4[40] ), .Z(\MC_ARK_ARC_1_3/temp6[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_25_1  ( .A1(\MC_ARK_ARC_1_3/temp2[40] ), .A2(
        \MC_ARK_ARC_1_3/temp1[40] ), .Z(\MC_ARK_ARC_1_3/temp5[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_25_1  ( .A1(\RI5[3][76] ), .A2(n486), .Z(
        \MC_ARK_ARC_1_3/temp4[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_25_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[178] ), 
        .A2(\RI5[3][10] ), .Z(\MC_ARK_ARC_1_3/temp2[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_25_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[40] ), 
        .A2(\RI5[3][34] ), .Z(\MC_ARK_ARC_1_3/temp1[40] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_25_0  ( .A1(\RI5[3][77] ), .A2(n550), .Z(
        \MC_ARK_ARC_1_3/temp4[41] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_25_0  ( .A1(\RI5[3][35] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[41] ), .Z(\MC_ARK_ARC_1_3/temp1[41] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_24_5  ( .A1(\MC_ARK_ARC_1_3/temp6[42] ), .A2(
        \MC_ARK_ARC_1_3/temp5[42] ), .Z(\MC_ARK_ARC_1_3/buf_output[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_24_5  ( .A1(\MC_ARK_ARC_1_3/temp3[42] ), .A2(
        \MC_ARK_ARC_1_3/temp4[42] ), .Z(\MC_ARK_ARC_1_3/temp6[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_24_5  ( .A1(\MC_ARK_ARC_1_3/temp1[42] ), .A2(
        \MC_ARK_ARC_1_3/temp2[42] ), .Z(\MC_ARK_ARC_1_3/temp5[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_24_5  ( .A1(\RI5[3][78] ), .A2(n484), .Z(
        \MC_ARK_ARC_1_3/temp4[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_24_5  ( .A1(\RI5[3][144] ), .A2(\RI5[3][108] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_24_5  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[12] ), 
        .A2(\RI5[3][180] ), .Z(\MC_ARK_ARC_1_3/temp2[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_24_5  ( .A1(\RI5[3][42] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[36] ), .Z(\MC_ARK_ARC_1_3/temp1[42] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_24_4  ( .A1(\RI5[3][79] ), .A2(n548), .Z(
        \MC_ARK_ARC_1_3/temp4[43] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_24_3  ( .A1(\RI5[3][80] ), .A2(n158), .Z(
        \MC_ARK_ARC_1_3/temp4[44] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_24_2  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[81] ), 
        .A2(n547), .Z(\MC_ARK_ARC_1_3/temp4[45] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_24_2  ( .A1(\RI5[3][15] ), .A2(\RI5[3][183] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[45] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_24_1  ( .A1(\MC_ARK_ARC_1_3/temp3[46] ), .A2(
        \MC_ARK_ARC_1_3/temp4[46] ), .Z(\MC_ARK_ARC_1_3/temp6[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_24_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[82] ), 
        .A2(n222), .Z(\MC_ARK_ARC_1_3/temp4[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_24_1  ( .A1(\RI5[3][184] ), .A2(\RI5[3][16] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[46] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_23_5  ( .A1(\RI5[3][84] ), .A2(n479), .Z(
        \MC_ARK_ARC_1_3/temp4[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_23_5  ( .A1(\RI5[3][18] ), .A2(\RI5[3][186] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[48] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_23_4  ( .A1(\MC_ARK_ARC_1_3/temp5[49] ), .A2(
        \MC_ARK_ARC_1_3/temp6[49] ), .Z(\MC_ARK_ARC_1_3/buf_output[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_23_4  ( .A1(\MC_ARK_ARC_1_3/temp4[49] ), .A2(
        \MC_ARK_ARC_1_3/temp3[49] ), .Z(\MC_ARK_ARC_1_3/temp6[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_23_4  ( .A1(\RI5[3][85] ), .A2(n194), .Z(
        \MC_ARK_ARC_1_3/temp4[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_23_4  ( .A1(\RI5[3][151] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[115] ), .Z(\MC_ARK_ARC_1_3/temp3[49] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_23_4  ( .A1(\RI5[3][43] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[49] ), .Z(\MC_ARK_ARC_1_3/temp1[49] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_23_3  ( .A1(\RI5[3][86] ), .A2(n202), .Z(
        \MC_ARK_ARC_1_3/temp4[50] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_23_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[152] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[116] ), .Z(
        \MC_ARK_ARC_1_3/temp3[50] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_23_2  ( .A1(\MC_ARK_ARC_1_3/temp1[51] ), .A2(
        \MC_ARK_ARC_1_3/temp2[51] ), .Z(\MC_ARK_ARC_1_3/temp5[51] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_23_2  ( .A1(\RI5[3][87] ), .A2(n243), .Z(
        \MC_ARK_ARC_1_3/temp4[51] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_23_2  ( .A1(\RI5[3][153] ), .A2(\RI5[3][117] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[51] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_23_2  ( .A1(\RI5[3][189] ), .A2(\RI5[3][21] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[51] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_23_2  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[51] ), 
        .A2(\RI5[3][45] ), .Z(\MC_ARK_ARC_1_3/temp1[51] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_23_1  ( .A1(\MC_ARK_ARC_1_3/temp3[52] ), .A2(
        \MC_ARK_ARC_1_3/temp4[52] ), .Z(\MC_ARK_ARC_1_3/temp6[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_23_1  ( .A1(\RI5[3][88] ), .A2(n105), .Z(
        \MC_ARK_ARC_1_3/temp4[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_23_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[154] ), 
        .A2(\RI5[3][118] ), .Z(\MC_ARK_ARC_1_3/temp3[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_23_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[22] ), 
        .A2(\RI5[3][190] ), .Z(\MC_ARK_ARC_1_3/temp2[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_23_1  ( .A1(\RI5[3][52] ), .A2(\RI5[3][46] ), .Z(
        \MC_ARK_ARC_1_3/temp1[52] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_23_0  ( .A1(\RI5[3][89] ), .A2(n543), .Z(
        \MC_ARK_ARC_1_3/temp4[53] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_22_5  ( .A1(\MC_ARK_ARC_1_3/temp4[54] ), .A2(
        \MC_ARK_ARC_1_3/temp3[54] ), .Z(\MC_ARK_ARC_1_3/temp6[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_22_5  ( .A1(\MC_ARK_ARC_1_3/temp2[54] ), .A2(
        \MC_ARK_ARC_1_3/temp1[54] ), .Z(\MC_ARK_ARC_1_3/temp5[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_22_5  ( .A1(n2896), .A2(n474), .Z(
        \MC_ARK_ARC_1_3/temp4[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_22_5  ( .A1(\RI5[3][156] ), .A2(\RI5[3][120] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_22_5  ( .A1(\RI5[3][48] ), .A2(\RI5[3][54] ), .Z(
        \MC_ARK_ARC_1_3/temp1[54] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_22_4  ( .A1(\MC_ARK_ARC_1_3/temp4[55] ), .A2(
        \MC_ARK_ARC_1_3/temp3[55] ), .Z(\MC_ARK_ARC_1_3/temp6[55] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_22_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[91] ), 
        .A2(n145), .Z(\MC_ARK_ARC_1_3/temp4[55] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_22_4  ( .A1(\RI5[3][121] ), .A2(\RI5[3][157] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[55] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_22_4  ( .A1(\RI5[3][25] ), .A2(\RI5[3][1] ), .Z(
        \MC_ARK_ARC_1_3/temp2[55] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_22_3  ( .A1(\MC_ARK_ARC_1_3/temp4[56] ), .A2(
        \MC_ARK_ARC_1_3/temp3[56] ), .Z(\MC_ARK_ARC_1_3/temp6[56] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_22_3  ( .A1(\RI5[3][92] ), .A2(n66), .Z(
        \MC_ARK_ARC_1_3/temp4[56] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_22_3  ( .A1(\RI5[3][158] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[122] ), .Z(\MC_ARK_ARC_1_3/temp3[56] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_22_2  ( .A1(\RI5[3][93] ), .A2(n107), .Z(
        \MC_ARK_ARC_1_3/temp4[57] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_22_2  ( .A1(\RI5[3][3] ), .A2(\RI5[3][27] ), .Z(
        \MC_ARK_ARC_1_3/temp2[57] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_22_1  ( .A1(\RI5[3][94] ), .A2(n21), .Z(
        \MC_ARK_ARC_1_3/temp4[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_22_1  ( .A1(\RI5[3][4] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[28] ), .Z(\MC_ARK_ARC_1_3/temp2[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_22_1  ( .A1(\RI5[3][58] ), .A2(\RI5[3][52] ), .Z(
        \MC_ARK_ARC_1_3/temp1[58] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_22_0  ( .A1(\RI5[3][95] ), .A2(n142), .Z(
        \MC_ARK_ARC_1_3/temp4[59] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_22_0  ( .A1(\RI5[3][29] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[5] ), .Z(\MC_ARK_ARC_1_3/temp2[59] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_21_5  ( .A1(\MC_ARK_ARC_1_3/temp2[60] ), .A2(
        \MC_ARK_ARC_1_3/temp1[60] ), .Z(\MC_ARK_ARC_1_3/temp5[60] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_21_5  ( .A1(\RI5[3][96] ), .A2(n470), .Z(
        \MC_ARK_ARC_1_3/temp4[60] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_21_5  ( .A1(\RI5[3][162] ), .A2(\RI5[3][126] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[60] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_21_5  ( .A1(\RI5[3][30] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[6] ), .Z(\MC_ARK_ARC_1_3/temp2[60] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_21_5  ( .A1(\RI5[3][60] ), .A2(\RI5[3][54] ), .Z(
        \MC_ARK_ARC_1_3/temp1[60] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_21_4  ( .A1(\MC_ARK_ARC_1_3/temp5[61] ), .A2(
        \MC_ARK_ARC_1_3/temp6[61] ), .Z(\MC_ARK_ARC_1_3/buf_output[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_21_4  ( .A1(\MC_ARK_ARC_1_3/temp3[61] ), .A2(
        \MC_ARK_ARC_1_3/temp4[61] ), .Z(\MC_ARK_ARC_1_3/temp6[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_21_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[97] ), 
        .A2(n538), .Z(\MC_ARK_ARC_1_3/temp4[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_21_4  ( .A1(\RI5[3][163] ), .A2(\RI5[3][127] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_21_4  ( .A1(\RI5[3][31] ), .A2(\RI5[3][7] ), .Z(
        \MC_ARK_ARC_1_3/temp2[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_21_4  ( .A1(\RI5[3][61] ), .A2(\RI5[3][55] ), .Z(
        \MC_ARK_ARC_1_3/temp1[61] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_21_3  ( .A1(\MC_ARK_ARC_1_3/temp2[62] ), .A2(
        \MC_ARK_ARC_1_3/temp1[62] ), .Z(\MC_ARK_ARC_1_3/temp5[62] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_21_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[56] ), 
        .A2(\RI5[3][62] ), .Z(\MC_ARK_ARC_1_3/temp1[62] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_21_2  ( .A1(\MC_ARK_ARC_1_3/temp3[63] ), .A2(
        \MC_ARK_ARC_1_3/temp4[63] ), .Z(\MC_ARK_ARC_1_3/temp6[63] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_21_2  ( .A1(\RI5[3][99] ), .A2(n537), .Z(
        \MC_ARK_ARC_1_3/temp4[63] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_21_2  ( .A1(\RI5[3][129] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[165] ), .Z(\MC_ARK_ARC_1_3/temp3[63] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_21_1  ( .A1(\MC_ARK_ARC_1_3/temp3[64] ), .A2(
        \MC_ARK_ARC_1_3/temp4[64] ), .Z(\MC_ARK_ARC_1_3/temp6[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_21_1  ( .A1(\MC_ARK_ARC_1_3/temp1[64] ), .A2(
        \MC_ARK_ARC_1_3/temp2[64] ), .Z(\MC_ARK_ARC_1_3/temp5[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_21_1  ( .A1(\RI5[3][100] ), .A2(n468), .Z(
        \MC_ARK_ARC_1_3/temp4[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_21_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[166] ), 
        .A2(\RI5[3][130] ), .Z(\MC_ARK_ARC_1_3/temp3[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_21_1  ( .A1(\RI5[3][34] ), .A2(\RI5[3][10] ), .Z(
        \MC_ARK_ARC_1_3/temp2[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_21_1  ( .A1(\RI5[3][64] ), .A2(\RI5[3][58] ), .Z(
        \MC_ARK_ARC_1_3/temp1[64] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_20_5  ( .A1(\RI5[3][102] ), .A2(n466), .Z(
        \MC_ARK_ARC_1_3/temp4[66] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_20_5  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[36] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[12] ), .Z(\MC_ARK_ARC_1_3/temp2[66] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_20_4  ( .A1(\MC_ARK_ARC_1_3/temp3[67] ), .A2(
        \MC_ARK_ARC_1_3/temp4[67] ), .Z(\MC_ARK_ARC_1_3/temp6[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_20_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[103] ), 
        .A2(n199), .Z(\MC_ARK_ARC_1_3/temp4[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_20_4  ( .A1(\RI5[3][169] ), .A2(\RI5[3][133] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_20_4  ( .A1(\RI5[3][37] ), .A2(\RI5[3][13] ), .Z(
        \MC_ARK_ARC_1_3/temp2[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_20_4  ( .A1(\RI5[3][61] ), .A2(\RI5[3][67] ), .Z(
        \MC_ARK_ARC_1_3/temp1[67] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_20_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[104] ), 
        .A2(n43), .Z(\MC_ARK_ARC_1_3/temp4[68] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_20_2  ( .A1(\MC_ARK_ARC_1_3/temp3[69] ), .A2(
        \MC_ARK_ARC_1_3/temp4[69] ), .Z(\MC_ARK_ARC_1_3/temp6[69] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_20_2  ( .A1(\SB2_3_16/buf_output[3] ), .A2(n531), 
        .Z(\MC_ARK_ARC_1_3/temp4[69] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_20_1  ( .A1(\RI5[3][106] ), .A2(n131), .Z(
        \MC_ARK_ARC_1_3/temp4[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_20_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[40] ), 
        .A2(\RI5[3][16] ), .Z(\MC_ARK_ARC_1_3/temp2[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_20_1  ( .A1(\RI5[3][70] ), .A2(\RI5[3][64] ), .Z(
        \MC_ARK_ARC_1_3/temp1[70] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_20_0  ( .A1(\RI5[3][107] ), .A2(n529), .Z(
        \MC_ARK_ARC_1_3/temp4[71] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_20_0  ( .A1(\RI5[3][173] ), .A2(\RI5[3][137] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[71] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_19_5  ( .A1(\MC_ARK_ARC_1_3/temp3[72] ), .A2(
        \MC_ARK_ARC_1_3/temp4[72] ), .Z(\MC_ARK_ARC_1_3/temp6[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_19_5  ( .A1(\RI5[3][108] ), .A2(n463), .Z(
        \MC_ARK_ARC_1_3/temp4[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_19_5  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[174] ), 
        .A2(\RI5[3][138] ), .Z(\MC_ARK_ARC_1_3/temp3[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_19_5  ( .A1(\RI5[3][42] ), .A2(\RI5[3][18] ), .Z(
        \MC_ARK_ARC_1_3/temp2[72] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_19_4  ( .A1(\MC_ARK_ARC_1_3/temp5[73] ), .A2(
        \MC_ARK_ARC_1_3/temp6[73] ), .Z(\MC_ARK_ARC_1_3/buf_output[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_19_4  ( .A1(\MC_ARK_ARC_1_3/temp3[73] ), .A2(
        \MC_ARK_ARC_1_3/temp4[73] ), .Z(\MC_ARK_ARC_1_3/temp6[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_19_4  ( .A1(\MC_ARK_ARC_1_3/temp1[73] ), .A2(
        \MC_ARK_ARC_1_3/temp2[73] ), .Z(\MC_ARK_ARC_1_3/temp5[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_19_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[109] ), 
        .A2(n527), .Z(\MC_ARK_ARC_1_3/temp4[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_19_4  ( .A1(\RI5[3][175] ), .A2(\RI5[3][139] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_19_4  ( .A1(\RI5[3][19] ), .A2(\RI5[3][43] ), .Z(
        \MC_ARK_ARC_1_3/temp2[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_19_4  ( .A1(\RI5[3][67] ), .A2(\RI5[3][73] ), .Z(
        \MC_ARK_ARC_1_3/temp1[73] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_19_3  ( .A1(\MC_ARK_ARC_1_3/temp3[74] ), .A2(
        \MC_ARK_ARC_1_3/temp4[74] ), .Z(\MC_ARK_ARC_1_3/temp6[74] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_19_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[110] ), 
        .A2(n37), .Z(\MC_ARK_ARC_1_3/temp4[74] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_19_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[44] ), 
        .A2(\RI5[3][20] ), .Z(\MC_ARK_ARC_1_3/temp2[74] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_19_2  ( .A1(n1392), .A2(n526), .Z(
        \MC_ARK_ARC_1_3/temp4[75] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_19_2  ( .A1(\RI5[3][141] ), .A2(\RI5[3][177] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[75] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_19_2  ( .A1(\RI5[3][69] ), .A2(\RI5[3][75] ), .Z(
        \MC_ARK_ARC_1_3/temp1[75] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_19_1  ( .A1(\MC_ARK_ARC_1_3/temp1[76] ), .A2(
        \MC_ARK_ARC_1_3/temp2[76] ), .Z(\MC_ARK_ARC_1_3/temp5[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_19_1  ( .A1(\RI5[3][112] ), .A2(n35), .Z(
        \MC_ARK_ARC_1_3/temp4[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_19_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[178] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[142] ), .Z(
        \MC_ARK_ARC_1_3/temp3[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_19_1  ( .A1(\RI5[3][46] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[22] ), .Z(\MC_ARK_ARC_1_3/temp2[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_19_1  ( .A1(\RI5[3][76] ), .A2(\RI5[3][70] ), .Z(
        \MC_ARK_ARC_1_3/temp1[76] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_19_0  ( .A1(\MC_ARK_ARC_1_3/temp3[77] ), .A2(
        \MC_ARK_ARC_1_3/temp4[77] ), .Z(\MC_ARK_ARC_1_3/temp6[77] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_19_0  ( .A1(\RI5[3][113] ), .A2(n90), .Z(
        \MC_ARK_ARC_1_3/temp4[77] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_18_5  ( .A1(\MC_ARK_ARC_1_3/temp5[78] ), .A2(
        \MC_ARK_ARC_1_3/temp6[78] ), .Z(\MC_ARK_ARC_1_3/buf_output[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_18_5  ( .A1(\SB2_3_17/buf_output[0] ), .A2(n459), 
        .Z(\MC_ARK_ARC_1_3/temp4[78] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_18_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[115] ), 
        .A2(n123), .Z(\MC_ARK_ARC_1_3/temp4[79] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_18_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[116] ), 
        .A2(n61), .Z(\MC_ARK_ARC_1_3/temp4[80] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_18_2  ( .A1(\MC_ARK_ARC_1_3/temp3[81] ), .A2(
        \MC_ARK_ARC_1_3/temp4[81] ), .Z(\MC_ARK_ARC_1_3/temp6[81] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_18_2  ( .A1(\RI5[3][117] ), .A2(n522), .Z(
        \MC_ARK_ARC_1_3/temp4[81] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_18_2  ( .A1(\RI5[3][75] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[81] ), .Z(\MC_ARK_ARC_1_3/temp1[81] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_18_1  ( .A1(\RI5[3][118] ), .A2(n143), .Z(
        \MC_ARK_ARC_1_3/temp4[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_18_1  ( .A1(\RI5[3][52] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[28] ), .Z(\MC_ARK_ARC_1_3/temp2[82] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_18_0  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[119] ), 
        .A2(n119), .Z(\MC_ARK_ARC_1_3/temp4[83] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_17_5  ( .A1(\RI5[3][120] ), .A2(n454), .Z(
        \MC_ARK_ARC_1_3/temp4[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_17_5  ( .A1(\RI5[3][150] ), .A2(\RI5[3][186] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_17_5  ( .A1(\RI5[3][84] ), .A2(\RI5[3][78] ), .Z(
        \MC_ARK_ARC_1_3/temp1[84] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_17_4  ( .A1(\RI5[3][121] ), .A2(n183), .Z(
        \MC_ARK_ARC_1_3/temp4[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_17_4  ( .A1(\RI5[3][187] ), .A2(\RI5[3][151] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_17_4  ( .A1(\RI5[3][55] ), .A2(\RI5[3][31] ), .Z(
        \MC_ARK_ARC_1_3/temp2[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_17_4  ( .A1(\RI5[3][85] ), .A2(\RI5[3][79] ), .Z(
        \MC_ARK_ARC_1_3/temp1[85] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_17_3  ( .A1(\MC_ARK_ARC_1_3/temp5[86] ), .A2(
        \MC_ARK_ARC_1_3/temp6[86] ), .Z(\MC_ARK_ARC_1_3/buf_output[86] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_17_3  ( .A1(\MC_ARK_ARC_1_3/temp3[86] ), .A2(
        \MC_ARK_ARC_1_3/temp4[86] ), .Z(\MC_ARK_ARC_1_3/temp6[86] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_17_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[122] ), 
        .A2(n140), .Z(\MC_ARK_ARC_1_3/temp4[86] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_17_2  ( .A1(\RI5[3][123] ), .A2(n240), .Z(
        \MC_ARK_ARC_1_3/temp4[87] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_17_2  ( .A1(\RI5[3][87] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[81] ), .Z(\MC_ARK_ARC_1_3/temp1[87] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_17_1  ( .A1(\MC_ARK_ARC_1_3/temp3[88] ), .A2(
        \MC_ARK_ARC_1_3/temp4[88] ), .Z(\MC_ARK_ARC_1_3/temp6[88] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_17_1  ( .A1(\MC_ARK_ARC_1_3/temp2[88] ), .A2(
        \MC_ARK_ARC_1_3/temp1[88] ), .Z(\MC_ARK_ARC_1_3/temp5[88] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_17_1  ( .A1(\RI5[3][124] ), .A2(n159), .Z(
        \MC_ARK_ARC_1_3/temp4[88] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_17_1  ( .A1(\RI5[3][190] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[154] ), .Z(\MC_ARK_ARC_1_3/temp3[88] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_17_1  ( .A1(\RI5[3][58] ), .A2(\RI5[3][34] ), .Z(
        \MC_ARK_ARC_1_3/temp2[88] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_17_1  ( .A1(\RI5[3][88] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[82] ), .Z(\MC_ARK_ARC_1_3/temp1[88] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_17_0  ( .A1(\RI5[3][125] ), .A2(n48), .Z(
        \MC_ARK_ARC_1_3/temp4[89] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_17_0  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[155] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[191] ), .Z(
        \MC_ARK_ARC_1_3/temp3[89] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_16_5  ( .A1(\RI5[3][126] ), .A2(n129), .Z(
        \MC_ARK_ARC_1_3/temp4[90] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_16_5  ( .A1(\RI5[3][0] ), .A2(\RI5[3][156] ), .Z(
        \MC_ARK_ARC_1_3/temp3[90] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_16_4  ( .A1(\MC_ARK_ARC_1_3/temp6[91] ), .A2(
        \MC_ARK_ARC_1_3/temp5[91] ), .Z(\MC_ARK_ARC_1_3/buf_output[91] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_16_3  ( .A1(\RI5[3][128] ), .A2(n19), .Z(
        \MC_ARK_ARC_1_3/temp4[92] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_16_3  ( .A1(\RI5[3][62] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[38] ), .Z(\MC_ARK_ARC_1_3/temp2[92] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_16_2  ( .A1(\RI5[3][129] ), .A2(n109), .Z(
        \MC_ARK_ARC_1_3/temp4[93] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_16_1  ( .A1(\RI5[3][130] ), .A2(n448), .Z(
        \MC_ARK_ARC_1_3/temp4[94] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_16_0  ( .A1(\RI5[3][131] ), .A2(n514), .Z(
        \MC_ARK_ARC_1_3/temp4[95] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_15_5  ( .A1(\MC_ARK_ARC_1_3/temp3[96] ), .A2(
        \MC_ARK_ARC_1_3/temp4[96] ), .Z(\MC_ARK_ARC_1_3/temp6[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_15_5  ( .A1(\MC_ARK_ARC_1_3/temp1[96] ), .A2(
        \MC_ARK_ARC_1_3/temp2[96] ), .Z(\MC_ARK_ARC_1_3/temp5[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_15_5  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[132] ), 
        .A2(n446), .Z(\MC_ARK_ARC_1_3/temp4[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_15_5  ( .A1(\RI5[3][162] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[6] ), .Z(\MC_ARK_ARC_1_3/temp3[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_15_5  ( .A1(\RI5[3][66] ), .A2(\RI5[3][42] ), .Z(
        \MC_ARK_ARC_1_3/temp2[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_15_5  ( .A1(n2896), .A2(\RI5[3][96] ), .Z(
        \MC_ARK_ARC_1_3/temp1[96] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_15_4  ( .A1(\MC_ARK_ARC_1_3/temp2[97] ), .A2(
        \MC_ARK_ARC_1_3/temp1[97] ), .Z(\MC_ARK_ARC_1_3/temp5[97] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_15_4  ( .A1(\RI5[3][133] ), .A2(n513), .Z(
        \MC_ARK_ARC_1_3/temp4[97] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_15_4  ( .A1(\RI5[3][7] ), .A2(\RI5[3][163] ), .Z(
        \MC_ARK_ARC_1_3/temp3[97] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_15_4  ( .A1(\RI5[3][43] ), .A2(\RI5[3][67] ), .Z(
        \MC_ARK_ARC_1_3/temp2[97] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_15_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[97] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[91] ), .Z(\MC_ARK_ARC_1_3/temp1[97] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_15_3  ( .A1(\MC_ARK_ARC_1_3/temp3[98] ), .A2(
        \MC_ARK_ARC_1_3/temp4[98] ), .Z(\MC_ARK_ARC_1_3/temp6[98] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_15_3  ( .A1(\MC_ARK_ARC_1_3/temp2[98] ), .A2(
        \MC_ARK_ARC_1_3/temp1[98] ), .Z(\MC_ARK_ARC_1_3/temp5[98] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_15_3  ( .A1(\RI5[3][134] ), .A2(n73), .Z(
        \MC_ARK_ARC_1_3/temp4[98] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_15_3  ( .A1(\RI5[3][164] ), .A2(\RI5[3][8] ), .Z(
        \MC_ARK_ARC_1_3/temp3[98] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_15_3  ( .A1(\RI5[3][68] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[44] ), .Z(\MC_ARK_ARC_1_3/temp2[98] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_15_3  ( .A1(\RI5[3][98] ), .A2(\RI5[3][92] ), .Z(
        \MC_ARK_ARC_1_3/temp1[98] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_15_2  ( .A1(\MC_ARK_ARC_1_3/temp6[99] ), .A2(
        \MC_ARK_ARC_1_3/temp5[99] ), .Z(\MC_ARK_ARC_1_3/buf_output[99] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_15_2  ( .A1(\MC_ARK_ARC_1_3/temp2[99] ), .A2(
        \MC_ARK_ARC_1_3/temp1[99] ), .Z(\MC_ARK_ARC_1_3/temp5[99] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_15_2  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[135] ), 
        .A2(n511), .Z(\MC_ARK_ARC_1_3/temp4[99] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_15_2  ( .A1(\RI5[3][69] ), .A2(\RI5[3][45] ), .Z(
        \MC_ARK_ARC_1_3/temp2[99] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_15_1  ( .A1(\MC_ARK_ARC_1_3/temp6[100] ), .A2(
        \MC_ARK_ARC_1_3/temp5[100] ), .Z(\MC_ARK_ARC_1_3/buf_output[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_15_1  ( .A1(\MC_ARK_ARC_1_3/temp3[100] ), .A2(
        \MC_ARK_ARC_1_3/temp4[100] ), .Z(\MC_ARK_ARC_1_3/temp6[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_15_1  ( .A1(\MC_ARK_ARC_1_3/temp1[100] ), .A2(
        \MC_ARK_ARC_1_3/temp2[100] ), .Z(\MC_ARK_ARC_1_3/temp5[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_15_1  ( .A1(\RI5[3][136] ), .A2(n11), .Z(
        \MC_ARK_ARC_1_3/temp4[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_15_1  ( .A1(\RI5[3][10] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[166] ), .Z(\MC_ARK_ARC_1_3/temp3[100] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_15_1  ( .A1(\RI5[3][70] ), .A2(\RI5[3][46] ), .Z(
        \MC_ARK_ARC_1_3/temp2[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_15_1  ( .A1(\RI5[3][100] ), .A2(\RI5[3][94] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[100] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_14_5  ( .A1(\RI5[3][138] ), .A2(n442), .Z(
        \MC_ARK_ARC_1_3/temp4[102] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_14_5  ( .A1(\RI5[3][72] ), .A2(\RI5[3][48] ), .Z(
        \MC_ARK_ARC_1_3/temp2[102] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_14_5  ( .A1(\SB2_3_20/buf_output[0] ), .A2(
        \RI5[3][102] ), .Z(\MC_ARK_ARC_1_3/temp1[102] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_14_4  ( .A1(\MC_ARK_ARC_1_3/temp1[103] ), .A2(
        \MC_ARK_ARC_1_3/temp2[103] ), .Z(\MC_ARK_ARC_1_3/temp5[103] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_14_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[49] ), 
        .A2(\RI5[3][73] ), .Z(\MC_ARK_ARC_1_3/temp2[103] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_14_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[103] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[97] ), .Z(
        \MC_ARK_ARC_1_3/temp1[103] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_14_3  ( .A1(\RI5[3][140] ), .A2(n137), .Z(
        \MC_ARK_ARC_1_3/temp4[104] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_14_2  ( .A1(\RI5[3][141] ), .A2(n507), .Z(
        \MC_ARK_ARC_1_3/temp4[105] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_14_2  ( .A1(\RI5[3][15] ), .A2(\RI5[3][171] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[105] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_14_1  ( .A1(\MC_ARK_ARC_1_3/temp5[106] ), .A2(
        \MC_ARK_ARC_1_3/temp6[106] ), .Z(\MC_ARK_ARC_1_3/buf_output[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_14_1  ( .A1(\MC_ARK_ARC_1_3/temp3[106] ), .A2(
        \MC_ARK_ARC_1_3/temp4[106] ), .Z(\MC_ARK_ARC_1_3/temp6[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_14_1  ( .A1(\MC_ARK_ARC_1_3/temp1[106] ), .A2(
        \MC_ARK_ARC_1_3/temp2[106] ), .Z(\MC_ARK_ARC_1_3/temp5[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_14_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[142] ), 
        .A2(n15), .Z(\MC_ARK_ARC_1_3/temp4[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_14_1  ( .A1(\RI5[3][16] ), .A2(\RI5[3][172] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_14_1  ( .A1(\RI5[3][76] ), .A2(\RI5[3][52] ), .Z(
        \MC_ARK_ARC_1_3/temp2[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_14_1  ( .A1(\RI5[3][106] ), .A2(\RI5[3][100] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[106] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_14_0  ( .A1(\RI5[3][77] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[53] ), .Z(\MC_ARK_ARC_1_3/temp2[107] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_13_5  ( .A1(\MC_ARK_ARC_1_3/temp3[108] ), .A2(
        \MC_ARK_ARC_1_3/temp4[108] ), .Z(\MC_ARK_ARC_1_3/temp6[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_13_5  ( .A1(\RI5[3][144] ), .A2(n4), .Z(
        \MC_ARK_ARC_1_3/temp4[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_13_5  ( .A1(\RI5[3][78] ), .A2(\RI5[3][54] ), .Z(
        \MC_ARK_ARC_1_3/temp2[108] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_13_4  ( .A1(\RI5[3][145] ), .A2(n504), .Z(
        \MC_ARK_ARC_1_3/temp4[109] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_13_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[103] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[109] ), .Z(
        \MC_ARK_ARC_1_3/temp1[109] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_13_3  ( .A1(\RI5[3][146] ), .A2(n437), .Z(
        \MC_ARK_ARC_1_3/temp4[110] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_13_2  ( .A1(\MC_ARK_ARC_1_3/temp3[111] ), .A2(
        \MC_ARK_ARC_1_3/temp4[111] ), .Z(\MC_ARK_ARC_1_3/temp6[111] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_13_2  ( .A1(\RI5[3][147] ), .A2(n178), .Z(
        \MC_ARK_ARC_1_3/temp4[111] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_13_2  ( .A1(\RI5[3][57] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[81] ), .Z(\MC_ARK_ARC_1_3/temp2[111] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_13_2  ( .A1(n1392), .A2(\RI5[3][105] ), .Z(
        \MC_ARK_ARC_1_3/temp1[111] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_13_1  ( .A1(\RI5[3][148] ), .A2(n566), .Z(
        \MC_ARK_ARC_1_3/temp4[112] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_13_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[22] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[178] ), .Z(
        \MC_ARK_ARC_1_3/temp3[112] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_13_0  ( .A1(\RI5[3][149] ), .A2(n187), .Z(
        \MC_ARK_ARC_1_3/temp4[113] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_12_5  ( .A1(\SB2_3_11/buf_output[0] ), .A2(n564), 
        .Z(\MC_ARK_ARC_1_3/temp4[114] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_12_5  ( .A1(\RI5[3][24] ), .A2(\RI5[3][180] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[114] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_12_5  ( .A1(\RI5[3][60] ), .A2(\RI5[3][84] ), .Z(
        \MC_ARK_ARC_1_3/temp2[114] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_12_4  ( .A1(\RI5[3][151] ), .A2(n500), .Z(
        \MC_ARK_ARC_1_3/temp4[115] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_12_4  ( .A1(\RI5[3][25] ), .A2(\RI5[3][181] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[115] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_12_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[115] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[109] ), .Z(
        \MC_ARK_ARC_1_3/temp1[115] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_12_3  ( .A1(\SB2_3_9/buf_output[2] ), .A2(n563), 
        .Z(\MC_ARK_ARC_1_3/temp4[116] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_12_3  ( .A1(\RI5[3][86] ), .A2(\RI5[3][62] ), .Z(
        \MC_ARK_ARC_1_3/temp2[116] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_12_2  ( .A1(\RI5[3][153] ), .A2(n87), .Z(
        \MC_ARK_ARC_1_3/temp4[117] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_12_2  ( .A1(\RI5[3][27] ), .A2(\RI5[3][183] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[117] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_12_1  ( .A1(\MC_ARK_ARC_1_3/temp2[118] ), .A2(
        \MC_ARK_ARC_1_3/temp1[118] ), .Z(\MC_ARK_ARC_1_3/temp5[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_12_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[154] ), 
        .A2(n561), .Z(\MC_ARK_ARC_1_3/temp4[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_12_1  ( .A1(\RI5[3][88] ), .A2(\RI5[3][64] ), .Z(
        \MC_ARK_ARC_1_3/temp2[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_12_1  ( .A1(\RI5[3][118] ), .A2(\RI5[3][112] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[118] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_12_0  ( .A1(\MC_ARK_ARC_1_3/temp5[119] ), .A2(
        \MC_ARK_ARC_1_3/temp6[119] ), .Z(\MC_ARK_ARC_1_3/buf_output[119] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_12_0  ( .A1(\MC_ARK_ARC_1_3/temp3[119] ), .A2(
        \MC_ARK_ARC_1_3/temp4[119] ), .Z(\MC_ARK_ARC_1_3/temp6[119] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_12_0  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[155] ), 
        .A2(n85), .Z(\MC_ARK_ARC_1_3/temp4[119] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_12_0  ( .A1(\RI5[3][29] ), .A2(\RI5[3][185] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[119] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_11_5  ( .A1(\MC_ARK_ARC_1_3/temp6[120] ), .A2(
        \MC_ARK_ARC_1_3/temp5[120] ), .Z(\MC_ARK_ARC_1_3/buf_output[120] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_11_5  ( .A1(\MC_ARK_ARC_1_3/temp4[120] ), .A2(
        \MC_ARK_ARC_1_3/temp3[120] ), .Z(\MC_ARK_ARC_1_3/temp6[120] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_11_5  ( .A1(\RI5[3][156] ), .A2(n175), .Z(
        \MC_ARK_ARC_1_3/temp4[120] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_11_5  ( .A1(\RI5[3][186] ), .A2(\RI5[3][30] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[120] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_11_5  ( .A1(\RI5[3][66] ), .A2(n2895), .Z(
        \MC_ARK_ARC_1_3/temp2[120] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_11_4  ( .A1(\MC_ARK_ARC_1_3/temp4[121] ), .A2(
        \MC_ARK_ARC_1_3/temp3[121] ), .Z(\MC_ARK_ARC_1_3/temp6[121] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_11_4  ( .A1(\RI5[3][157] ), .A2(n497), .Z(
        \MC_ARK_ARC_1_3/temp4[121] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_11_4  ( .A1(\RI5[3][187] ), .A2(\RI5[3][31] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[121] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_11_4  ( .A1(\RI5[3][121] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[115] ), .Z(\MC_ARK_ARC_1_3/temp1[121] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_11_3  ( .A1(\RI5[3][158] ), .A2(n560), .Z(
        \MC_ARK_ARC_1_3/temp4[122] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_11_3  ( .A1(\RI5[3][188] ), .A2(\RI5[3][32] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[122] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_11_3  ( .A1(\RI5[3][68] ), .A2(\RI5[3][92] ), .Z(
        \MC_ARK_ARC_1_3/temp2[122] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_11_2  ( .A1(\RI5[3][159] ), .A2(n496), .Z(
        \MC_ARK_ARC_1_3/temp4[123] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_11_1  ( .A1(\RI5[3][34] ), .A2(\RI5[3][190] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[124] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_11_1  ( .A1(\RI5[3][94] ), .A2(\RI5[3][70] ), .Z(
        \MC_ARK_ARC_1_3/temp2[124] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_11_1  ( .A1(\RI5[3][124] ), .A2(\RI5[3][118] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[124] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_11_0  ( .A1(\RI5[3][161] ), .A2(n494), .Z(
        \MC_ARK_ARC_1_3/temp4[125] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_11_0  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[191] ), 
        .A2(\RI5[3][35] ), .Z(\MC_ARK_ARC_1_3/temp3[125] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_11_0  ( .A1(\RI5[3][95] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[71] ), .Z(\MC_ARK_ARC_1_3/temp2[125] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_10_5  ( .A1(\MC_ARK_ARC_1_3/temp5[126] ), .A2(
        \MC_ARK_ARC_1_3/temp6[126] ), .Z(\MC_ARK_ARC_1_3/buf_output[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_10_5  ( .A1(\MC_ARK_ARC_1_3/temp2[126] ), .A2(
        \MC_ARK_ARC_1_3/temp1[126] ), .Z(\MC_ARK_ARC_1_3/temp5[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_10_5  ( .A1(\RI5[3][162] ), .A2(n147), .Z(
        \MC_ARK_ARC_1_3/temp4[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_10_5  ( .A1(\RI5[3][96] ), .A2(\RI5[3][72] ), .Z(
        \MC_ARK_ARC_1_3/temp2[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_10_5  ( .A1(\RI5[3][126] ), .A2(\RI5[3][120] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[126] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_10_4  ( .A1(\RI5[3][163] ), .A2(n204), .Z(
        \MC_ARK_ARC_1_3/temp4[127] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_10_3  ( .A1(n3679), .A2(n228), .Z(
        \MC_ARK_ARC_1_3/temp4[128] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_10_2  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[165] ), 
        .A2(n229), .Z(\MC_ARK_ARC_1_3/temp4[129] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_10_2  ( .A1(\RI5[3][39] ), .A2(\RI5[3][3] ), .Z(
        \MC_ARK_ARC_1_3/temp3[129] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_10_2  ( .A1(n3658), .A2(\RI5[3][129] ), .Z(
        \MC_ARK_ARC_1_3/temp1[129] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_10_1  ( .A1(\MC_ARK_ARC_1_3/temp5[130] ), .A2(
        \MC_ARK_ARC_1_3/temp6[130] ), .Z(\MC_ARK_ARC_1_3/buf_output[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_10_1  ( .A1(\MC_ARK_ARC_1_3/temp4[130] ), .A2(
        \MC_ARK_ARC_1_3/temp3[130] ), .Z(\MC_ARK_ARC_1_3/temp6[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_10_1  ( .A1(\MC_ARK_ARC_1_3/temp1[130] ), .A2(
        \MC_ARK_ARC_1_3/temp2[130] ), .Z(\MC_ARK_ARC_1_3/temp5[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_10_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[166] ), 
        .A2(n555), .Z(\MC_ARK_ARC_1_3/temp4[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_10_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[40] ), 
        .A2(\RI5[3][4] ), .Z(\MC_ARK_ARC_1_3/temp3[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_10_1  ( .A1(\RI5[3][100] ), .A2(\RI5[3][76] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[130] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_10_0  ( .A1(\MC_ARK_ARC_1_3/temp3[131] ), .A2(
        \MC_ARK_ARC_1_3/temp4[131] ), .Z(\MC_ARK_ARC_1_3/temp6[131] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_10_0  ( .A1(n1365), .A2(n490), .Z(
        \MC_ARK_ARC_1_3/temp4[131] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_9_5  ( .A1(\MC_ARK_ARC_1_3/temp5[132] ), .A2(
        \MC_ARK_ARC_1_3/temp6[132] ), .Z(\MC_ARK_ARC_1_3/buf_output[132] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_9_5  ( .A1(\MC_ARK_ARC_1_3/temp4[132] ), .A2(
        \MC_ARK_ARC_1_3/temp3[132] ), .Z(\MC_ARK_ARC_1_3/temp6[132] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_9_5  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[168] ), 
        .A2(n136), .Z(\MC_ARK_ARC_1_3/temp4[132] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_9_5  ( .A1(\RI5[3][42] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[6] ), .Z(\MC_ARK_ARC_1_3/temp3[132] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_9_5  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[132] ), 
        .A2(\RI5[3][126] ), .Z(\MC_ARK_ARC_1_3/temp1[132] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_9_4  ( .A1(\MC_ARK_ARC_1_3/temp3[133] ), .A2(
        \MC_ARK_ARC_1_3/temp4[133] ), .Z(\MC_ARK_ARC_1_3/temp6[133] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_9_4  ( .A1(\MC_ARK_ARC_1_3/temp1[133] ), .A2(
        \MC_ARK_ARC_1_3/temp2[133] ), .Z(\MC_ARK_ARC_1_3/temp5[133] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_9_4  ( .A1(\RI5[3][169] ), .A2(n488), .Z(
        \MC_ARK_ARC_1_3/temp4[133] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_9_4  ( .A1(\RI5[3][7] ), .A2(\RI5[3][43] ), .Z(
        \MC_ARK_ARC_1_3/temp3[133] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_9_4  ( .A1(\RI5[3][79] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[103] ), .Z(\MC_ARK_ARC_1_3/temp2[133] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_9_4  ( .A1(\RI5[3][133] ), .A2(\RI5[3][127] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[133] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_9_3  ( .A1(\MC_ARK_ARC_1_3/temp6[134] ), .A2(
        \MC_ARK_ARC_1_3/temp5[134] ), .Z(\MC_ARK_ARC_1_3/buf_output[134] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_9_3  ( .A1(\MC_ARK_ARC_1_3/temp2[134] ), .A2(
        \MC_ARK_ARC_1_3/temp1[134] ), .Z(\MC_ARK_ARC_1_3/temp5[134] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_9_3  ( .A1(\RI5[3][170] ), .A2(n230), .Z(
        \MC_ARK_ARC_1_3/temp4[134] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_9_3  ( .A1(\RI5[3][80] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[104] ), .Z(\MC_ARK_ARC_1_3/temp2[134] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_9_3  ( .A1(\RI5[3][134] ), .A2(\RI5[3][128] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[134] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_9_2  ( .A1(\RI5[3][171] ), .A2(n69), .Z(
        \MC_ARK_ARC_1_3/temp4[135] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_9_2  ( .A1(\RI5[3][9] ), .A2(\RI5[3][45] ), .Z(
        \MC_ARK_ARC_1_3/temp3[135] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_9_2  ( .A1(\RI5[3][105] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[81] ), .Z(\MC_ARK_ARC_1_3/temp2[135] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_9_2  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[135] ), 
        .A2(\RI5[3][129] ), .Z(\MC_ARK_ARC_1_3/temp1[135] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_9_1  ( .A1(\MC_ARK_ARC_1_3/temp2[136] ), .A2(
        \MC_ARK_ARC_1_3/temp1[136] ), .Z(\MC_ARK_ARC_1_3/temp5[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_9_1  ( .A1(\RI5[3][172] ), .A2(n551), .Z(
        \MC_ARK_ARC_1_3/temp4[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_9_1  ( .A1(\RI5[3][46] ), .A2(\RI5[3][10] ), .Z(
        \MC_ARK_ARC_1_3/temp3[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_9_1  ( .A1(\RI5[3][106] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[82] ), .Z(\MC_ARK_ARC_1_3/temp2[136] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_9_1  ( .A1(\RI5[3][136] ), .A2(\RI5[3][130] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[136] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_9_0  ( .A1(\MC_ARK_ARC_1_3/temp2[137] ), .A2(
        \MC_ARK_ARC_1_3/temp1[137] ), .Z(\MC_ARK_ARC_1_3/temp5[137] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_9_0  ( .A1(\RI5[3][173] ), .A2(n34), .Z(
        \MC_ARK_ARC_1_3/temp4[137] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_9_0  ( .A1(\RI5[3][11] ), .A2(\RI5[3][47] ), .Z(
        \MC_ARK_ARC_1_3/temp3[137] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_9_0  ( .A1(\RI5[3][107] ), .A2(\RI5[3][83] ), .Z(
        \MC_ARK_ARC_1_3/temp2[137] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_9_0  ( .A1(\RI5[3][131] ), .A2(\RI5[3][137] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[137] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_8_5  ( .A1(\MC_ARK_ARC_1_3/temp4[138] ), .A2(
        \MC_ARK_ARC_1_3/temp3[138] ), .Z(\MC_ARK_ARC_1_3/temp6[138] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_8_5  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[174] ), 
        .A2(n549), .Z(\MC_ARK_ARC_1_3/temp4[138] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_8_5  ( .A1(\RI5[3][48] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[12] ), .Z(\MC_ARK_ARC_1_3/temp3[138] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_8_4  ( .A1(\MC_ARK_ARC_1_3/temp5[139] ), .A2(
        \MC_ARK_ARC_1_3/temp6[139] ), .Z(\MC_ARK_ARC_1_3/buf_output[139] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_8_4  ( .A1(\MC_ARK_ARC_1_3/temp3[139] ), .A2(
        \MC_ARK_ARC_1_3/temp4[139] ), .Z(\MC_ARK_ARC_1_3/temp6[139] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_8_4  ( .A1(\MC_ARK_ARC_1_3/temp1[139] ), .A2(
        \MC_ARK_ARC_1_3/temp2[139] ), .Z(\MC_ARK_ARC_1_3/temp5[139] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_8_4  ( .A1(\RI5[3][175] ), .A2(n213), .Z(
        \MC_ARK_ARC_1_3/temp4[139] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_8_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[49] ), 
        .A2(\RI5[3][13] ), .Z(\MC_ARK_ARC_1_3/temp3[139] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_8_4  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[109] ), 
        .A2(\RI5[3][85] ), .Z(\MC_ARK_ARC_1_3/temp2[139] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_8_4  ( .A1(\RI5[3][139] ), .A2(\RI5[3][133] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[139] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_8_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[176] ), 
        .A2(n155), .Z(\MC_ARK_ARC_1_3/temp4[140] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_8_3  ( .A1(\RI5[3][86] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[110] ), .Z(\MC_ARK_ARC_1_3/temp2[140] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_8_2  ( .A1(\SB2_3_4/buf_output[3] ), .A2(n481), 
        .Z(\MC_ARK_ARC_1_3/temp4[141] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_8_2  ( .A1(\SB2_3_19/buf_output[3] ), .A2(n1392), 
        .Z(\MC_ARK_ARC_1_3/temp2[141] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_8_1  ( .A1(\MC_ARK_ARC_1_3/temp6[142] ), .A2(
        \MC_ARK_ARC_1_3/temp5[142] ), .Z(\MC_ARK_ARC_1_3/buf_output[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_8_1  ( .A1(\MC_ARK_ARC_1_3/temp3[142] ), .A2(
        \MC_ARK_ARC_1_3/temp4[142] ), .Z(\MC_ARK_ARC_1_3/temp6[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_8_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[178] ), 
        .A2(n152), .Z(\MC_ARK_ARC_1_3/temp4[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_8_1  ( .A1(\RI5[3][52] ), .A2(\RI5[3][16] ), .Z(
        \MC_ARK_ARC_1_3/temp3[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_8_1  ( .A1(\RI5[3][112] ), .A2(\RI5[3][88] ), .Z(
        \MC_ARK_ARC_1_3/temp2[142] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_8_0  ( .A1(\MC_ARK_ARC_1_3/temp4[143] ), .A2(
        \MC_ARK_ARC_1_3/temp3[143] ), .Z(\MC_ARK_ARC_1_3/temp6[143] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_8_0  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[179] ), 
        .A2(n480), .Z(\MC_ARK_ARC_1_3/temp4[143] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_8_0  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[17] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[53] ), .Z(
        \MC_ARK_ARC_1_3/temp3[143] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_7_5  ( .A1(\MC_ARK_ARC_1_3/temp5[144] ), .A2(
        \MC_ARK_ARC_1_3/temp6[144] ), .Z(\MC_ARK_ARC_1_3/buf_output[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_7_5  ( .A1(\MC_ARK_ARC_1_3/temp3[144] ), .A2(
        \MC_ARK_ARC_1_3/temp4[144] ), .Z(\MC_ARK_ARC_1_3/temp6[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_7_5  ( .A1(\MC_ARK_ARC_1_3/temp1[144] ), .A2(
        \MC_ARK_ARC_1_3/temp2[144] ), .Z(\MC_ARK_ARC_1_3/temp5[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_7_5  ( .A1(\RI5[3][180] ), .A2(n151), .Z(
        \MC_ARK_ARC_1_3/temp4[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_7_5  ( .A1(\RI5[3][54] ), .A2(\RI5[3][18] ), .Z(
        \MC_ARK_ARC_1_3/temp3[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_7_5  ( .A1(n2896), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[114] ), .Z(\MC_ARK_ARC_1_3/temp2[144] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_7_5  ( .A1(\RI5[3][144] ), .A2(\RI5[3][138] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[144] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_7_4  ( .A1(\MC_ARK_ARC_1_3/temp5[145] ), .A2(
        \MC_ARK_ARC_1_3/temp6[145] ), .Z(\MC_ARK_ARC_1_3/buf_output[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_7_4  ( .A1(\MC_ARK_ARC_1_3/temp4[145] ), .A2(
        \MC_ARK_ARC_1_3/temp3[145] ), .Z(\MC_ARK_ARC_1_3/temp6[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_7_4  ( .A1(\RI5[3][181] ), .A2(n478), .Z(
        \MC_ARK_ARC_1_3/temp4[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_7_4  ( .A1(\RI5[3][19] ), .A2(\RI5[3][55] ), .Z(
        \MC_ARK_ARC_1_3/temp3[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_7_4  ( .A1(\RI5[3][145] ), .A2(\RI5[3][139] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[145] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_7_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[182] ), 
        .A2(n149), .Z(\MC_ARK_ARC_1_3/temp4[146] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_7_3  ( .A1(\RI5[3][92] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[116] ), .Z(\MC_ARK_ARC_1_3/temp2[146] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_7_3  ( .A1(\RI5[3][146] ), .A2(\RI5[3][140] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[146] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_7_2  ( .A1(\RI5[3][183] ), .A2(n477), .Z(
        \MC_ARK_ARC_1_3/temp4[147] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_7_2  ( .A1(\RI5[3][93] ), .A2(\RI5[3][117] ), .Z(
        \MC_ARK_ARC_1_3/temp2[147] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_7_1  ( .A1(\MC_ARK_ARC_1_3/temp3[148] ), .A2(
        \MC_ARK_ARC_1_3/temp4[148] ), .Z(\MC_ARK_ARC_1_3/temp6[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_7_1  ( .A1(\RI5[3][184] ), .A2(n544), .Z(
        \MC_ARK_ARC_1_3/temp4[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_7_1  ( .A1(\RI5[3][58] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[22] ), .Z(\MC_ARK_ARC_1_3/temp3[148] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_7_1  ( .A1(\RI5[3][118] ), .A2(\RI5[3][94] ), .Z(
        \MC_ARK_ARC_1_3/temp2[148] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_7_1  ( .A1(\RI5[3][148] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[142] ), .Z(\MC_ARK_ARC_1_3/temp1[148] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_7_0  ( .A1(\MC_ARK_ARC_1_3/temp3[149] ), .A2(
        \MC_ARK_ARC_1_3/temp4[149] ), .Z(\MC_ARK_ARC_1_3/temp6[149] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_7_0  ( .A1(\RI5[3][185] ), .A2(n2), .Z(
        \MC_ARK_ARC_1_3/temp4[149] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_7_0  ( .A1(\RI5[3][23] ), .A2(\RI5[3][59] ), .Z(
        \MC_ARK_ARC_1_3/temp3[149] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_7_0  ( .A1(\RI5[3][95] ), .A2(n5503), .Z(
        \MC_ARK_ARC_1_3/temp2[149] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_7_0  ( .A1(\RI5[3][143] ), .A2(\RI5[3][149] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[149] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_6_5  ( .A1(\MC_ARK_ARC_1_3/temp5[150] ), .A2(
        \MC_ARK_ARC_1_3/temp6[150] ), .Z(\MC_ARK_ARC_1_3/buf_output[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_6_5  ( .A1(\MC_ARK_ARC_1_3/temp3[150] ), .A2(
        \MC_ARK_ARC_1_3/temp4[150] ), .Z(\MC_ARK_ARC_1_3/temp6[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_6_5  ( .A1(\MC_ARK_ARC_1_3/temp2[150] ), .A2(
        \MC_ARK_ARC_1_3/temp1[150] ), .Z(\MC_ARK_ARC_1_3/temp5[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_6_5  ( .A1(\RI5[3][186] ), .A2(n542), .Z(
        \MC_ARK_ARC_1_3/temp4[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_6_5  ( .A1(\RI5[3][60] ), .A2(\RI5[3][24] ), .Z(
        \MC_ARK_ARC_1_3/temp3[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_6_5  ( .A1(\RI5[3][96] ), .A2(\RI5[3][120] ), .Z(
        \MC_ARK_ARC_1_3/temp2[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_6_5  ( .A1(\RI5[3][150] ), .A2(\RI5[3][144] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[150] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_6_4  ( .A1(\MC_ARK_ARC_1_3/temp5[151] ), .A2(
        \MC_ARK_ARC_1_3/temp6[151] ), .Z(\MC_ARK_ARC_1_3/buf_output[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_6_4  ( .A1(\MC_ARK_ARC_1_3/temp3[151] ), .A2(
        \MC_ARK_ARC_1_3/temp4[151] ), .Z(\MC_ARK_ARC_1_3/temp6[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_6_4  ( .A1(\RI5[3][187] ), .A2(n54), .Z(
        \MC_ARK_ARC_1_3/temp4[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_6_4  ( .A1(\RI5[3][61] ), .A2(\RI5[3][25] ), .Z(
        \MC_ARK_ARC_1_3/temp3[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_6_4  ( .A1(\RI5[3][145] ), .A2(\RI5[3][151] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[151] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_6_3  ( .A1(\RI5[3][188] ), .A2(n169), .Z(
        \MC_ARK_ARC_1_3/temp4[152] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_6_3  ( .A1(\RI5[3][98] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[122] ), .Z(\MC_ARK_ARC_1_3/temp2[152] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_6_2  ( .A1(\MC_ARK_ARC_1_3/temp1[153] ), .A2(
        \MC_ARK_ARC_1_3/temp2[153] ), .Z(\MC_ARK_ARC_1_3/temp5[153] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_6_2  ( .A1(\RI5[3][123] ), .A2(\RI5[3][99] ), .Z(
        \MC_ARK_ARC_1_3/temp2[153] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_6_2  ( .A1(\RI5[3][147] ), .A2(\RI5[3][153] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[153] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_6_1  ( .A1(\RI5[3][190] ), .A2(n13), .Z(
        \MC_ARK_ARC_1_3/temp4[154] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_6_1  ( .A1(\RI5[3][64] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[28] ), .Z(\MC_ARK_ARC_1_3/temp3[154] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_6_1  ( .A1(\RI5[3][124] ), .A2(\RI5[3][100] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[154] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_6_1  ( .A1(\RI5[3][148] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[154] ), .Z(\MC_ARK_ARC_1_3/temp1[154] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_6_0  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[191] ), 
        .A2(n471), .Z(\MC_ARK_ARC_1_3/temp4[155] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_6_0  ( .A1(\RI5[3][125] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[101] ), .Z(\MC_ARK_ARC_1_3/temp2[155] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_5_5  ( .A1(\RI5[3][0] ), .A2(n539), .Z(
        \MC_ARK_ARC_1_3/temp4[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_5_5  ( .A1(\RI5[3][156] ), .A2(\RI5[3][150] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[156] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_5_4  ( .A1(\MC_ARK_ARC_1_3/temp5[157] ), .A2(
        \MC_ARK_ARC_1_3/temp6[157] ), .Z(\MC_ARK_ARC_1_3/buf_output[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_5_4  ( .A1(\RI5[3][1] ), .A2(n226), .Z(
        \MC_ARK_ARC_1_3/temp4[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_5_4  ( .A1(\SB2_3_24/buf_output[1] ), .A2(
        \RI5[3][31] ), .Z(\MC_ARK_ARC_1_3/temp3[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_5_4  ( .A1(\RI5[3][157] ), .A2(\RI5[3][151] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[157] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_5_3  ( .A1(\RI5[3][2] ), .A2(n234), .Z(
        \MC_ARK_ARC_1_3/temp4[158] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_5_2  ( .A1(\RI5[3][3] ), .A2(n469), .Z(
        \MC_ARK_ARC_1_3/temp4[159] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_5_2  ( .A1(\RI5[3][105] ), .A2(\RI5[3][129] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[159] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_5_1  ( .A1(\MC_ARK_ARC_1_3/temp5[160] ), .A2(
        \MC_ARK_ARC_1_3/temp6[160] ), .Z(\MC_ARK_ARC_1_3/buf_output[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_5_1  ( .A1(\MC_ARK_ARC_1_3/temp3[160] ), .A2(
        \MC_ARK_ARC_1_3/temp4[160] ), .Z(\MC_ARK_ARC_1_3/temp6[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_5_1  ( .A1(\RI5[3][4] ), .A2(n98), .Z(
        \MC_ARK_ARC_1_3/temp4[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_5_1  ( .A1(\RI5[3][70] ), .A2(\RI5[3][34] ), .Z(
        \MC_ARK_ARC_1_3/temp3[160] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_5_0  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[5] ), 
        .A2(n467), .Z(\MC_ARK_ARC_1_3/temp4[161] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_4_5  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[6] ), 
        .A2(n534), .Z(\MC_ARK_ARC_1_3/temp4[162] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_4_5  ( .A1(\SB2_3_10/buf_output[0] ), .A2(
        \SB2_3_9/buf_output[0] ), .Z(\MC_ARK_ARC_1_3/temp1[162] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_4_3  ( .A1(\RI5[3][8] ), .A2(n218), .Z(
        \MC_ARK_ARC_1_3/temp4[164] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_4_2  ( .A1(\MC_ARK_ARC_1_3/temp3[165] ), .A2(
        \MC_ARK_ARC_1_3/temp4[165] ), .Z(\MC_ARK_ARC_1_3/temp6[165] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_4_2  ( .A1(\RI5[3][9] ), .A2(n465), .Z(
        \MC_ARK_ARC_1_3/temp4[165] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_4_1  ( .A1(\RI5[3][136] ), .A2(\RI5[3][112] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[166] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_4_0  ( .A1(\RI5[3][11] ), .A2(n464), .Z(
        \MC_ARK_ARC_1_3/temp4[167] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_3_5  ( .A1(\MC_ARK_ARC_1_3/temp5[168] ), .A2(
        \MC_ARK_ARC_1_3/temp6[168] ), .Z(\MC_ARK_ARC_1_3/buf_output[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_3_5  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[12] ), 
        .A2(n528), .Z(\MC_ARK_ARC_1_3/temp4[168] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_3_4  ( .A1(\RI5[3][13] ), .A2(n462), .Z(
        \MC_ARK_ARC_1_3/temp4[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_3_4  ( .A1(\RI5[3][43] ), .A2(\RI5[3][79] ), .Z(
        \MC_ARK_ARC_1_3/temp3[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_3_4  ( .A1(\RI5[3][169] ), .A2(\RI5[3][163] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[169] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_3_3  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[14] ), 
        .A2(n217), .Z(\MC_ARK_ARC_1_3/temp4[170] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_3_2  ( .A1(\RI5[3][15] ), .A2(n461), .Z(
        \MC_ARK_ARC_1_3/temp4[171] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_3_2  ( .A1(\RI5[3][45] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[81] ), .Z(\MC_ARK_ARC_1_3/temp3[171] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_3_1  ( .A1(\RI5[3][16] ), .A2(n53), .Z(
        \MC_ARK_ARC_1_3/temp4[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_3_1  ( .A1(\RI5[3][46] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[82] ), .Z(\MC_ARK_ARC_1_3/temp3[172] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_3_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[142] ), 
        .A2(\RI5[3][118] ), .Z(\MC_ARK_ARC_1_3/temp2[172] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_3_1  ( .A1(\RI5[3][172] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[166] ), .Z(\MC_ARK_ARC_1_3/temp1[172] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_3_0  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[17] ), 
        .A2(n121), .Z(\MC_ARK_ARC_1_3/temp4[173] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_2_5  ( .A1(\RI5[3][18] ), .A2(n207), .Z(
        \MC_ARK_ARC_1_3/temp4[174] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_2_5  ( .A1(\RI5[3][84] ), .A2(\RI5[3][48] ), .Z(
        \MC_ARK_ARC_1_3/temp3[174] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_2_5  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[174] ), 
        .A2(\MC_ARK_ARC_1_3/buf_datainput[168] ), .Z(
        \MC_ARK_ARC_1_3/temp1[174] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_2_4  ( .A1(\RI5[3][19] ), .A2(n215), .Z(
        \MC_ARK_ARC_1_3/temp4[175] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_2_4  ( .A1(\RI5[3][121] ), .A2(\RI5[3][145] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[175] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_2_4  ( .A1(\RI5[3][169] ), .A2(\RI5[3][175] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[175] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_2_3  ( .A1(\MC_ARK_ARC_1_3/temp5[176] ), .A2(
        \MC_ARK_ARC_1_3/temp6[176] ), .Z(\MC_ARK_ARC_1_3/buf_output[176] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_2_3  ( .A1(\RI5[3][146] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[122] ), .Z(\MC_ARK_ARC_1_3/temp2[176] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_2_3  ( .A1(\RI5[3][170] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[176] ), .Z(\MC_ARK_ARC_1_3/temp1[176] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_2_2  ( .A1(\MC_ARK_ARC_1_3/temp3[177] ), .A2(
        \MC_ARK_ARC_1_3/temp4[177] ), .Z(\MC_ARK_ARC_1_3/temp6[177] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_2_2  ( .A1(\RI5[3][21] ), .A2(n118), .Z(
        \MC_ARK_ARC_1_3/temp4[177] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_2_2  ( .A1(\RI5[3][147] ), .A2(n3658), .Z(
        \MC_ARK_ARC_1_3/temp2[177] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_2_2  ( .A1(\RI5[3][177] ), .A2(\RI5[3][171] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[177] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_2_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[22] ), 
        .A2(n224), .Z(\MC_ARK_ARC_1_3/temp4[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_2_1  ( .A1(\RI5[3][88] ), .A2(\RI5[3][52] ), .Z(
        \MC_ARK_ARC_1_3/temp3[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_2_1  ( .A1(\RI5[3][148] ), .A2(\RI5[3][124] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_2_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[178] ), 
        .A2(\RI5[3][172] ), .Z(\MC_ARK_ARC_1_3/temp1[178] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_2_0  ( .A1(\RI5[3][23] ), .A2(n141), .Z(
        \MC_ARK_ARC_1_3/temp4[179] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_1_5  ( .A1(\RI5[3][24] ), .A2(n521), .Z(
        \MC_ARK_ARC_1_3/temp4[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_1_5  ( .A1(n2896), .A2(\RI5[3][54] ), .Z(
        \MC_ARK_ARC_1_3/temp3[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_1_5  ( .A1(\RI5[3][126] ), .A2(\RI5[3][150] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_1_5  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[174] ), 
        .A2(\RI5[3][180] ), .Z(\MC_ARK_ARC_1_3/temp1[180] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_1_4  ( .A1(\MC_ARK_ARC_1_3/temp1[181] ), .A2(
        \MC_ARK_ARC_1_3/temp2[181] ), .Z(\MC_ARK_ARC_1_3/temp5[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_1_4  ( .A1(\RI5[3][25] ), .A2(n453), .Z(
        \MC_ARK_ARC_1_3/temp4[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_1_4  ( .A1(\RI5[3][55] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[91] ), .Z(\MC_ARK_ARC_1_3/temp3[181] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_1_4  ( .A1(\RI5[3][151] ), .A2(\RI5[3][127] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_1_4  ( .A1(\RI5[3][181] ), .A2(\RI5[3][175] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[181] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_1_2  ( .A1(\MC_ARK_ARC_1_3/temp1[183] ), .A2(
        \MC_ARK_ARC_1_3/temp2[183] ), .Z(\MC_ARK_ARC_1_3/temp5[183] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_1_2  ( .A1(\RI5[3][27] ), .A2(n231), .Z(
        \MC_ARK_ARC_1_3/temp4[183] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_1_2  ( .A1(\RI5[3][177] ), .A2(\RI5[3][183] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[183] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X5_1_1  ( .A1(\MC_ARK_ARC_1_3/temp2[184] ), .A2(
        \MC_ARK_ARC_1_3/temp1[184] ), .Z(\MC_ARK_ARC_1_3/temp5[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_1_1  ( .A1(\MC_ARK_ARC_1_3/buf_datainput[28] ), 
        .A2(n518), .Z(\MC_ARK_ARC_1_3/temp4[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_1_1  ( .A1(\RI5[3][58] ), .A2(\RI5[3][94] ), .Z(
        \MC_ARK_ARC_1_3/temp3[184] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_1_1  ( .A1(\RI5[3][184] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[178] ), .Z(\MC_ARK_ARC_1_3/temp1[184] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_0_5  ( .A1(\RI5[3][30] ), .A2(n146), .Z(
        \MC_ARK_ARC_1_3/temp4[186] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_0_5  ( .A1(\RI5[3][156] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[132] ), .Z(\MC_ARK_ARC_1_3/temp2[186] )
         );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_0_5  ( .A1(\RI5[3][186] ), .A2(\RI5[3][180] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[186] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_0_4  ( .A1(\RI5[3][31] ), .A2(n128), .Z(
        \MC_ARK_ARC_1_3/temp4[187] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_0_4  ( .A1(\RI5[3][181] ), .A2(\RI5[3][187] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[187] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X3_0_3  ( .A1(\RI5[3][62] ), .A2(\RI5[3][98] ), .Z(
        \MC_ARK_ARC_1_3/temp3[188] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_0_2  ( .A1(\RI5[3][33] ), .A2(n220), .Z(
        \MC_ARK_ARC_1_3/temp4[189] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X7_0_1  ( .A1(\MC_ARK_ARC_1_3/temp5[190] ), .A2(
        \MC_ARK_ARC_1_3/temp6[190] ), .Z(\MC_ARK_ARC_1_3/buf_output[190] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_0_1  ( .A1(\RI5[3][34] ), .A2(n515), .Z(
        \MC_ARK_ARC_1_3/temp4[190] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X1_0_1  ( .A1(\RI5[3][184] ), .A2(\RI5[3][190] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[190] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X6_0_0  ( .A1(\MC_ARK_ARC_1_3/temp3[191] ), .A2(
        \MC_ARK_ARC_1_3/temp4[191] ), .Z(\MC_ARK_ARC_1_3/temp6[191] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X4_0_0  ( .A1(\RI5[3][35] ), .A2(n447), .Z(
        \MC_ARK_ARC_1_3/temp4[191] ) );
  XOR2_X1 \MC_ARK_ARC_1_3/X2_0_0  ( .A1(\RI5[3][161] ), .A2(\RI5[3][137] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[191] ) );
  INV_X1 \SB1_0_0/INV_5  ( .I(n436), .ZN(\SB1_0_0/i1_5 ) );
  INV_X1 \SB1_0_0/INV_4  ( .I(n404), .ZN(\SB1_0_0/i0[7] ) );
  INV_X1 \SB1_0_0/INV_0  ( .I(n338), .ZN(\SB1_0_0/i3[0] ) );
  INV_X1 \SB1_0_1/INV_5  ( .I(n435), .ZN(\SB1_0_1/i1_5 ) );
  INV_X1 \SB1_0_1/INV_1  ( .I(n336), .ZN(\SB1_0_1/i1_7 ) );
  INV_X1 \SB1_0_1/INV_0  ( .I(n335), .ZN(\SB1_0_1/i3[0] ) );
  INV_X1 \SB1_0_2/INV_5  ( .I(n434), .ZN(\SB1_0_2/i1_5 ) );
  INV_X1 \SB1_0_2/INV_4  ( .I(n400), .ZN(\SB1_0_2/i0[7] ) );
  INV_X1 \SB1_0_2/INV_1  ( .I(n333), .ZN(\SB1_0_2/i1_7 ) );
  INV_X1 \SB1_0_2/INV_0  ( .I(n332), .ZN(\SB1_0_2/i3[0] ) );
  INV_X1 \SB1_0_3/INV_5  ( .I(n433), .ZN(\SB1_0_3/i1_5 ) );
  INV_X1 \SB1_0_3/INV_4  ( .I(n398), .ZN(\SB1_0_3/i0[7] ) );
  INV_X1 \SB1_0_3/INV_1  ( .I(n330), .ZN(\SB1_0_3/i1_7 ) );
  INV_X1 \SB1_0_3/INV_0  ( .I(n329), .ZN(\SB1_0_3/i3[0] ) );
  INV_X1 \SB1_0_4/INV_5  ( .I(n432), .ZN(\SB1_0_4/i1_5 ) );
  INV_X1 \SB1_0_4/INV_4  ( .I(n396), .ZN(\SB1_0_4/i0[7] ) );
  INV_X1 \SB1_0_4/INV_1  ( .I(n327), .ZN(\SB1_0_4/i1_7 ) );
  INV_X1 \SB1_0_4/INV_0  ( .I(n326), .ZN(\SB1_0_4/i3[0] ) );
  INV_X1 \SB1_0_5/INV_5  ( .I(n431), .ZN(\SB1_0_5/i1_5 ) );
  INV_X1 \SB1_0_5/INV_1  ( .I(n324), .ZN(\SB1_0_5/i1_7 ) );
  INV_X1 \SB1_0_7/INV_4  ( .I(n5496), .ZN(\SB1_0_7/i0[7] ) );
  INV_X1 \SB1_0_7/INV_1  ( .I(n318), .ZN(\SB1_0_7/i1_7 ) );
  INV_X1 \SB1_0_7/INV_0  ( .I(n317), .ZN(\SB1_0_7/i3[0] ) );
  INV_X1 \SB1_0_8/INV_1  ( .I(n315), .ZN(\SB1_0_8/i1_7 ) );
  INV_X1 \SB1_0_8/INV_0  ( .I(n314), .ZN(\SB1_0_8/i3[0] ) );
  INV_X1 \SB1_0_9/INV_5  ( .I(n427), .ZN(\SB1_0_9/i1_5 ) );
  INV_X1 \SB1_0_9/INV_1  ( .I(n312), .ZN(\SB1_0_9/i1_7 ) );
  INV_X1 \SB1_0_9/INV_0  ( .I(n311), .ZN(\SB1_0_9/i3[0] ) );
  INV_X1 \SB1_0_10/INV_5  ( .I(n426), .ZN(\SB1_0_10/i1_5 ) );
  INV_X1 \SB1_0_10/INV_1  ( .I(n309), .ZN(\SB1_0_10/i1_7 ) );
  INV_X1 \SB1_0_10/INV_0  ( .I(n308), .ZN(\SB1_0_10/i3[0] ) );
  INV_X1 \SB1_0_11/INV_4  ( .I(n382), .ZN(\SB1_0_11/i0[7] ) );
  INV_X1 \SB1_0_11/INV_1  ( .I(n306), .ZN(\SB1_0_11/i1_7 ) );
  INV_X1 \SB1_0_11/INV_0  ( .I(n305), .ZN(\SB1_0_11/i3[0] ) );
  INV_X1 \SB1_0_12/INV_5  ( .I(n424), .ZN(\SB1_0_12/i1_5 ) );
  INV_X1 \SB1_0_12/INV_4  ( .I(n380), .ZN(\SB1_0_12/i0[7] ) );
  INV_X1 \SB1_0_12/INV_1  ( .I(n303), .ZN(\SB1_0_12/i1_7 ) );
  INV_X1 \SB1_0_12/INV_0  ( .I(n302), .ZN(\SB1_0_12/i3[0] ) );
  INV_X1 \SB1_0_13/INV_4  ( .I(n378), .ZN(\SB1_0_13/i0[7] ) );
  INV_X1 \SB1_0_13/INV_0  ( .I(n299), .ZN(\SB1_0_13/i3[0] ) );
  INV_X1 \SB1_0_14/INV_5  ( .I(n422), .ZN(\SB1_0_14/i1_5 ) );
  INV_X1 \SB1_0_14/INV_4  ( .I(n376), .ZN(\SB1_0_14/i0[7] ) );
  INV_X1 \SB1_0_14/INV_1  ( .I(n297), .ZN(\SB1_0_14/i1_7 ) );
  INV_X1 \SB1_0_15/INV_4  ( .I(n374), .ZN(\SB1_0_15/i0[7] ) );
  INV_X1 \SB1_0_15/INV_1  ( .I(n294), .ZN(\SB1_0_15/i1_7 ) );
  INV_X1 \SB1_0_15/INV_0  ( .I(n293), .ZN(\SB1_0_15/i3[0] ) );
  INV_X1 \SB1_0_16/INV_1  ( .I(n291), .ZN(\SB1_0_16/i1_7 ) );
  INV_X1 \SB1_0_17/INV_5  ( .I(n419), .ZN(\SB1_0_17/i1_5 ) );
  INV_X1 \SB1_0_17/INV_0  ( .I(n287), .ZN(\SB1_0_17/i3[0] ) );
  INV_X1 \SB1_0_18/INV_4  ( .I(n4753), .ZN(\SB1_0_18/i0[7] ) );
  INV_X1 \SB1_0_18/INV_1  ( .I(n285), .ZN(\SB1_0_18/i1_7 ) );
  INV_X1 \SB1_0_18/INV_0  ( .I(n284), .ZN(\SB1_0_18/i3[0] ) );
  INV_X1 \SB1_0_19/INV_5  ( .I(n417), .ZN(\SB1_0_19/i1_5 ) );
  INV_X1 \SB1_0_19/INV_4  ( .I(n366), .ZN(\SB1_0_19/i0[7] ) );
  INV_X1 \SB1_0_19/INV_1  ( .I(n282), .ZN(\SB1_0_19/i1_7 ) );
  INV_X1 \SB1_0_19/INV_0  ( .I(n281), .ZN(\SB1_0_19/i3[0] ) );
  INV_X1 \SB1_0_20/INV_5  ( .I(n416), .ZN(\SB1_0_20/i1_5 ) );
  INV_X1 \SB1_0_20/INV_1  ( .I(n279), .ZN(\SB1_0_20/i1_7 ) );
  INV_X1 \SB1_0_20/INV_0  ( .I(n278), .ZN(\SB1_0_20/i3[0] ) );
  INV_X1 \SB1_0_21/INV_4  ( .I(n362), .ZN(\SB1_0_21/i0[7] ) );
  INV_X1 \SB1_0_21/INV_1  ( .I(n276), .ZN(\SB1_0_21/i1_7 ) );
  INV_X1 \SB1_0_21/INV_0  ( .I(n275), .ZN(\SB1_0_21/i3[0] ) );
  INV_X1 \SB1_0_22/INV_5  ( .I(n414), .ZN(\SB1_0_22/i1_5 ) );
  INV_X1 \SB1_0_22/INV_4  ( .I(n360), .ZN(\SB1_0_22/i0[7] ) );
  INV_X1 \SB1_0_22/INV_1  ( .I(n273), .ZN(\SB1_0_22/i1_7 ) );
  INV_X1 \SB1_0_22/INV_0  ( .I(n272), .ZN(\SB1_0_22/i3[0] ) );
  INV_X1 \SB1_0_23/INV_0  ( .I(n269), .ZN(\SB1_0_23/i3[0] ) );
  INV_X1 \SB1_0_24/INV_5  ( .I(n412), .ZN(\SB1_0_24/i1_5 ) );
  INV_X1 \SB1_0_24/INV_4  ( .I(n356), .ZN(\SB1_0_24/i0[7] ) );
  INV_X1 \SB1_0_24/INV_1  ( .I(n267), .ZN(\SB1_0_24/i1_7 ) );
  INV_X1 \SB1_0_24/INV_0  ( .I(n266), .ZN(\SB1_0_24/i3[0] ) );
  INV_X1 \SB1_0_26/INV_5  ( .I(n410), .ZN(\SB1_0_26/i1_5 ) );
  INV_X1 \SB1_0_26/INV_4  ( .I(n352), .ZN(\SB1_0_26/i0[7] ) );
  INV_X1 \SB1_0_26/INV_1  ( .I(n261), .ZN(\SB1_0_26/i1_7 ) );
  INV_X1 \SB1_0_26/INV_0  ( .I(n260), .ZN(\SB1_0_26/i3[0] ) );
  INV_X1 \SB1_0_27/INV_5  ( .I(n409), .ZN(\SB1_0_27/i1_5 ) );
  INV_X1 \SB1_0_27/INV_4  ( .I(n350), .ZN(\SB1_0_27/i0[7] ) );
  INV_X1 \SB1_0_27/INV_1  ( .I(n258), .ZN(\SB1_0_27/i1_7 ) );
  INV_X1 \SB1_0_27/INV_0  ( .I(n257), .ZN(\SB1_0_27/i3[0] ) );
  INV_X1 \SB1_0_28/INV_4  ( .I(n6314), .ZN(\SB1_0_28/i0[7] ) );
  INV_X1 \SB1_0_28/INV_0  ( .I(n254), .ZN(\SB1_0_28/i3[0] ) );
  INV_X1 \SB1_0_29/INV_4  ( .I(n346), .ZN(\SB1_0_29/i0[7] ) );
  INV_X1 \SB1_0_29/INV_1  ( .I(n252), .ZN(\SB1_0_29/i1_7 ) );
  INV_X1 \SB1_0_30/INV_5  ( .I(n406), .ZN(\SB1_0_30/i1_5 ) );
  INV_X1 \SB1_0_30/INV_1  ( .I(n249), .ZN(\SB1_0_30/i1_7 ) );
  INV_X1 \SB1_0_30/INV_0  ( .I(n248), .ZN(\SB1_0_30/i3[0] ) );
  INV_X1 \SB1_0_31/INV_5  ( .I(n405), .ZN(\SB1_0_31/i1_5 ) );
  INV_X1 \SB1_0_31/INV_4  ( .I(n342), .ZN(\SB1_0_31/i0[7] ) );
  INV_X1 \SB1_0_31/INV_1  ( .I(n246), .ZN(\SB1_0_31/i1_7 ) );
  INV_X1 \SB1_0_31/INV_0  ( .I(n245), .ZN(\SB1_0_31/i3[0] ) );
  INV_X1 \SB2_0_0/INV_4  ( .I(\SB1_0_1/buf_output[4] ), .ZN(\SB2_0_0/i0[7] )
         );
  INV_X1 \SB2_0_0/INV_1  ( .I(\SB1_0_4/buf_output[1] ), .ZN(\SB2_0_0/i1_7 ) );
  INV_X1 \SB2_0_2/INV_1  ( .I(\RI3[0][175] ), .ZN(\SB2_0_2/i1_7 ) );
  INV_X1 \SB2_0_2/INV_0  ( .I(\SB1_0_7/buf_output[0] ), .ZN(\SB2_0_2/i3[0] )
         );
  INV_X1 \SB2_0_4/INV_0  ( .I(\RI3[0][162] ), .ZN(\SB2_0_4/i3[0] ) );
  INV_X1 \SB2_0_5/INV_1  ( .I(\SB1_0_9/buf_output[1] ), .ZN(\SB2_0_5/i1_7 ) );
  INV_X1 \SB2_0_5/INV_0  ( .I(\SB1_0_10/buf_output[0] ), .ZN(\SB2_0_5/i3[0] )
         );
  INV_X1 \SB2_0_6/INV_1  ( .I(\SB1_0_10/buf_output[1] ), .ZN(\SB2_0_6/i1_7 )
         );
  INV_X1 \SB2_0_6/INV_0  ( .I(\SB1_0_11/buf_output[0] ), .ZN(\SB2_0_6/i3[0] )
         );
  INV_X1 \SB2_0_7/INV_1  ( .I(\SB2_0_7/i0[6] ), .ZN(\SB2_0_7/i1_7 ) );
  INV_X1 \SB2_0_7/INV_0  ( .I(\SB1_0_12/buf_output[0] ), .ZN(\SB2_0_7/i3[0] )
         );
  INV_X1 \SB2_0_8/INV_0  ( .I(\SB1_0_13/buf_output[0] ), .ZN(\SB2_0_8/i3[0] )
         );
  INV_X1 \SB2_0_9/INV_0  ( .I(\SB1_0_14/buf_output[0] ), .ZN(\SB2_0_9/i3[0] )
         );
  INV_X1 \SB2_0_11/INV_1  ( .I(\RI3[0][121] ), .ZN(\SB2_0_11/i1_7 ) );
  INV_X1 \SB2_0_12/INV_4  ( .I(\RI3[0][118] ), .ZN(\SB2_0_12/i0[7] ) );
  INV_X1 \SB2_0_12/INV_1  ( .I(\SB1_0_16/buf_output[1] ), .ZN(\SB2_0_12/i1_7 )
         );
  INV_X1 \SB2_0_16/INV_0  ( .I(\SB1_0_21/buf_output[0] ), .ZN(\SB2_0_16/i3[0] ) );
  INV_X1 \SB2_0_17/INV_0  ( .I(\RI3[0][84] ), .ZN(\SB2_0_17/i3[0] ) );
  INV_X1 \SB2_0_18/INV_4  ( .I(\SB1_0_19/buf_output[4] ), .ZN(\SB2_0_18/i0[7] ) );
  INV_X1 \SB2_0_18/INV_1  ( .I(\RI3[0][79] ), .ZN(\SB2_0_18/i1_7 ) );
  INV_X1 \SB2_0_19/INV_0  ( .I(\RI3[0][72] ), .ZN(\SB2_0_19/i3[0] ) );
  INV_X1 \SB2_0_21/INV_4  ( .I(\SB1_0_22/buf_output[4] ), .ZN(\SB2_0_21/i0[7] ) );
  INV_X1 \SB2_0_21/INV_0  ( .I(\SB1_0_26/buf_output[0] ), .ZN(\SB2_0_21/i3[0] ) );
  INV_X1 \SB2_0_22/INV_4  ( .I(\RI3[0][58] ), .ZN(\SB2_0_22/i0[7] ) );
  INV_X2 \SB2_0_22/INV_3  ( .I(\RI3[0][57] ), .ZN(\SB2_0_22/i0[8] ) );
  INV_X1 \SB2_0_23/INV_1  ( .I(\RI3[0][49] ), .ZN(\SB2_0_23/i1_7 ) );
  INV_X1 \SB2_0_24/INV_0  ( .I(\SB1_0_29/buf_output[0] ), .ZN(\SB2_0_24/i3[0] ) );
  INV_X1 \SB2_0_25/INV_4  ( .I(\SB1_0_26/buf_output[4] ), .ZN(\SB2_0_25/i0[7] ) );
  INV_X1 \SB2_0_26/INV_1  ( .I(\SB1_0_30/buf_output[1] ), .ZN(\SB2_0_26/i1_7 )
         );
  INV_X1 \SB2_0_26/INV_0  ( .I(\RI3[0][30] ), .ZN(\SB2_0_26/i3[0] ) );
  INV_X2 \SB2_0_27/INV_3  ( .I(\RI3[0][27] ), .ZN(\SB2_0_27/i0[8] ) );
  INV_X2 \SB2_0_27/INV_2  ( .I(\SB1_0_30/buf_output[2] ), .ZN(\SB2_0_27/i1[9] ) );
  INV_X1 \SB2_0_29/INV_4  ( .I(\SB1_0_30/buf_output[4] ), .ZN(\SB2_0_29/i0[7] ) );
  INV_X1 \SB2_0_29/INV_1  ( .I(\SB1_0_1/buf_output[1] ), .ZN(\SB2_0_29/i1_7 )
         );
  INV_X2 \SB2_0_30/INV_3  ( .I(\RI3[0][9] ), .ZN(\SB2_0_30/i0[8] ) );
  INV_X2 \SB2_0_30/INV_2  ( .I(\RI3[0][8] ), .ZN(\SB2_0_30/i1[9] ) );
  INV_X1 \SB2_0_30/INV_1  ( .I(\RI3[0][7] ), .ZN(\SB2_0_30/i1_7 ) );
  INV_X1 \SB2_0_31/INV_4  ( .I(\SB1_0_0/buf_output[4] ), .ZN(\SB2_0_31/i0[7] )
         );
  INV_X1 \SB2_0_31/INV_1  ( .I(\RI3[0][1] ), .ZN(\SB2_0_31/i1_7 ) );
  INV_X1 \SB2_0_31/INV_0  ( .I(\SB1_0_4/buf_output[0] ), .ZN(\SB2_0_31/i3[0] )
         );
  INV_X1 \SB1_1_0/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[190] ), .ZN(
        \SB1_1_0/i0[7] ) );
  INV_X1 \SB1_1_1/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[184] ), .ZN(
        \SB1_1_1/i0[7] ) );
  INV_X2 \SB1_1_1/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[183] ), .ZN(
        \SB1_1_1/i0[8] ) );
  INV_X1 \SB1_1_2/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[178] ), .ZN(
        \SB1_1_2/i0[7] ) );
  INV_X2 \SB1_1_2/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[177] ), .ZN(
        \SB1_1_2/i0[8] ) );
  INV_X2 \SB1_1_2/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[176] ), .ZN(
        \SB1_1_2/i1[9] ) );
  INV_X1 \SB1_1_3/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[172] ), .ZN(
        \SB1_1_3/i0[7] ) );
  INV_X1 \SB1_1_4/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[166] ), .ZN(
        \SB1_1_4/i0[7] ) );
  INV_X2 \SB1_1_4/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[165] ), .ZN(
        \SB1_1_4/i0[8] ) );
  INV_X1 \SB1_1_5/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[160] ), .ZN(
        \SB1_1_5/i0[7] ) );
  INV_X2 \SB1_1_5/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[159] ), .ZN(
        \SB1_1_5/i0[8] ) );
  INV_X1 \SB1_1_6/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[154] ), .ZN(
        \SB1_1_6/i0[7] ) );
  INV_X2 \SB1_1_6/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[153] ), .ZN(
        \SB1_1_6/i0[8] ) );
  INV_X1 \SB1_1_7/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[148] ), .ZN(
        \SB1_1_7/i0[7] ) );
  INV_X2 \SB1_1_7/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[147] ), .ZN(
        \SB1_1_7/i0[8] ) );
  INV_X1 \SB1_1_7/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[145] ), .ZN(
        \SB1_1_7/i1_7 ) );
  INV_X1 \SB1_1_8/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[142] ), .ZN(
        \SB1_1_8/i0[7] ) );
  INV_X1 \SB1_1_9/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[136] ), .ZN(
        \SB1_1_9/i0[7] ) );
  INV_X2 \SB1_1_9/INV_3  ( .I(n1377), .ZN(\SB1_1_9/i0[8] ) );
  INV_X1 \SB1_1_10/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[130] ), .ZN(
        \SB1_1_10/i0[7] ) );
  INV_X2 \SB1_1_10/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[129] ), .ZN(
        \SB1_1_10/i0[8] ) );
  INV_X2 \SB1_1_10/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[128] ), .ZN(
        \SB1_1_10/i1[9] ) );
  INV_X1 \SB1_1_11/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[124] ), .ZN(
        \SB1_1_11/i0[7] ) );
  INV_X2 \SB1_1_11/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[123] ), .ZN(
        \SB1_1_11/i0[8] ) );
  INV_X1 \SB1_1_11/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[120] ), .ZN(
        \SB1_1_11/i3[0] ) );
  INV_X1 \SB1_1_12/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[118] ), .ZN(
        \SB1_1_12/i0[7] ) );
  INV_X2 \SB1_1_12/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[117] ), .ZN(
        \SB1_1_12/i0[8] ) );
  INV_X2 \SB1_1_12/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[116] ), .ZN(
        \SB1_1_12/i1[9] ) );
  INV_X1 \SB1_1_12/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[115] ), .ZN(
        \SB1_1_12/i1_7 ) );
  INV_X1 \SB1_1_13/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[112] ), .ZN(
        \SB1_1_13/i0[7] ) );
  INV_X2 \SB1_1_13/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[111] ), .ZN(
        \SB1_1_13/i0[8] ) );
  INV_X2 \SB1_1_14/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[105] ), .ZN(
        \SB1_1_14/i0[8] ) );
  INV_X1 \SB1_1_15/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[100] ), .ZN(
        \SB1_1_15/i0[7] ) );
  INV_X1 \SB1_1_15/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[96] ), .ZN(
        \SB1_1_15/i3[0] ) );
  INV_X2 \SB1_1_16/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[93] ), .ZN(
        \SB1_1_16/i0[8] ) );
  INV_X2 \SB1_1_16/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[92] ), .ZN(
        \SB1_1_16/i1[9] ) );
  INV_X1 \SB1_1_17/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[88] ), .ZN(
        \SB1_1_17/i0[7] ) );
  INV_X2 \SB1_1_17/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[87] ), .ZN(
        \SB1_1_17/i0[8] ) );
  INV_X1 \SB1_1_18/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[82] ), .ZN(
        \SB1_1_18/i0[7] ) );
  INV_X1 \SB1_1_18/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[79] ), .ZN(
        \SB1_1_18/i1_7 ) );
  INV_X1 \SB1_1_18/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[78] ), .ZN(
        \SB1_1_18/i3[0] ) );
  INV_X1 \SB1_1_19/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[76] ), .ZN(
        \SB1_1_19/i0[7] ) );
  INV_X2 \SB1_1_19/INV_3  ( .I(n3672), .ZN(\SB1_1_19/i0[8] ) );
  INV_X1 \SB1_1_20/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[70] ), .ZN(
        \SB1_1_20/i0[7] ) );
  INV_X1 \SB1_1_21/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[64] ), .ZN(
        \SB1_1_21/i0[7] ) );
  INV_X2 \SB1_1_21/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[63] ), .ZN(
        \SB1_1_21/i0[8] ) );
  INV_X2 \SB1_1_22/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[57] ), .ZN(
        \SB1_1_22/i0[8] ) );
  INV_X2 \SB1_1_22/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[56] ), .ZN(
        \SB1_1_22/i1[9] ) );
  INV_X1 \SB1_1_23/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[52] ), .ZN(
        \SB1_1_23/i0[7] ) );
  INV_X2 \SB1_1_23/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[51] ), .ZN(
        \SB1_1_23/i0[8] ) );
  INV_X1 \SB1_1_24/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[46] ), .ZN(
        \SB1_1_24/i0[7] ) );
  INV_X1 \SB1_1_24/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[43] ), .ZN(
        \SB1_1_24/i1_7 ) );
  INV_X1 \SB1_1_24/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[42] ), .ZN(
        \SB1_1_24/i3[0] ) );
  INV_X1 \SB1_1_25/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[41] ), .ZN(
        \SB1_1_25/i1_5 ) );
  INV_X1 \SB1_1_25/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[40] ), .ZN(
        \SB1_1_25/i0[7] ) );
  INV_X2 \SB1_1_25/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[39] ), .ZN(
        \SB1_1_25/i0[8] ) );
  INV_X1 \SB1_1_25/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[36] ), .ZN(
        \SB1_1_25/i3[0] ) );
  INV_X1 \SB1_1_26/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[34] ), .ZN(
        \SB1_1_26/i0[7] ) );
  INV_X2 \SB1_1_26/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[32] ), .ZN(
        \SB1_1_26/i1[9] ) );
  INV_X1 \SB1_1_27/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[28] ), .ZN(
        \SB1_1_27/i0[7] ) );
  INV_X1 \SB1_1_28/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[22] ), .ZN(
        \SB1_1_28/i0[7] ) );
  INV_X2 \SB1_1_28/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[21] ), .ZN(
        \SB1_1_28/i0[8] ) );
  INV_X2 \SB1_1_28/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[20] ), .ZN(
        \SB1_1_28/i1[9] ) );
  INV_X1 \SB1_1_29/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[16] ), .ZN(
        \SB1_1_29/i0[7] ) );
  INV_X2 \SB1_1_29/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[15] ), .ZN(
        \SB1_1_29/i0[8] ) );
  INV_X1 \SB1_1_30/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[10] ), .ZN(
        \SB1_1_30/i0[7] ) );
  INV_X2 \SB1_1_30/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[9] ), .ZN(
        \SB1_1_30/i0[8] ) );
  INV_X2 \SB1_1_30/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[8] ), .ZN(
        \SB1_1_30/i1[9] ) );
  INV_X1 \SB1_1_30/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[6] ), .ZN(
        \SB1_1_30/i3[0] ) );
  INV_X1 \SB1_1_31/INV_4  ( .I(\MC_ARK_ARC_1_0/buf_output[4] ), .ZN(
        \SB1_1_31/i0[7] ) );
  INV_X1 \SB1_1_31/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[1] ), .ZN(
        \SB1_1_31/i1_7 ) );
  INV_X1 \SB1_1_31/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[0] ), .ZN(
        \SB1_1_31/i3[0] ) );
  INV_X1 \SB2_1_0/INV_1  ( .I(\SB1_1_4/buf_output[1] ), .ZN(\SB2_1_0/i1_7 ) );
  INV_X1 \SB2_1_0/INV_0  ( .I(\SB1_1_5/buf_output[0] ), .ZN(\SB2_1_0/i3[0] )
         );
  INV_X1 \SB2_1_1/INV_4  ( .I(\SB1_1_2/buf_output[4] ), .ZN(\SB2_1_1/i0[7] )
         );
  INV_X2 \SB2_1_1/INV_3  ( .I(\SB1_1_3/buf_output[3] ), .ZN(\SB2_1_1/i0[8] )
         );
  INV_X1 \SB2_1_2/INV_4  ( .I(\SB1_1_3/buf_output[4] ), .ZN(\SB2_1_2/i0[7] )
         );
  INV_X2 \SB2_1_2/INV_3  ( .I(\SB1_1_4/buf_output[3] ), .ZN(\SB2_1_2/i0[8] )
         );
  INV_X2 \SB2_1_3/INV_3  ( .I(\SB1_1_5/buf_output[3] ), .ZN(\SB2_1_3/i0[8] )
         );
  INV_X2 \SB2_1_4/INV_3  ( .I(\SB1_1_6/buf_output[3] ), .ZN(\SB2_1_4/i0[8] )
         );
  INV_X2 \SB2_1_5/INV_3  ( .I(\SB1_1_7/buf_output[3] ), .ZN(\SB2_1_5/i0[8] )
         );
  INV_X1 \SB2_1_5/INV_0  ( .I(\SB1_1_10/buf_output[0] ), .ZN(\SB2_1_5/i3[0] )
         );
  INV_X1 \SB2_1_6/INV_4  ( .I(\SB1_1_7/buf_output[4] ), .ZN(\SB2_1_6/i0[7] )
         );
  INV_X1 \SB2_1_6/INV_0  ( .I(\SB1_1_11/buf_output[0] ), .ZN(\SB2_1_6/i3[0] )
         );
  INV_X1 \SB2_1_7/INV_0  ( .I(\SB1_1_12/buf_output[0] ), .ZN(\SB2_1_7/i3[0] )
         );
  INV_X1 \SB2_1_8/INV_4  ( .I(\SB1_1_9/buf_output[4] ), .ZN(\SB2_1_8/i0[7] )
         );
  INV_X1 \SB2_1_8/INV_1  ( .I(\SB1_1_12/buf_output[1] ), .ZN(\SB2_1_8/i1_7 )
         );
  INV_X1 \SB2_1_9/INV_4  ( .I(\SB1_1_10/buf_output[4] ), .ZN(\SB2_1_9/i0[7] )
         );
  INV_X1 \SB2_1_9/INV_0  ( .I(\SB1_1_14/buf_output[0] ), .ZN(\SB2_1_9/i3[0] )
         );
  INV_X2 \SB2_1_10/INV_3  ( .I(\SB1_1_12/buf_output[3] ), .ZN(\SB2_1_10/i0[8] ) );
  INV_X1 \SB2_1_10/INV_0  ( .I(\SB1_1_15/buf_output[0] ), .ZN(\SB2_1_10/i3[0] ) );
  INV_X2 \SB2_1_11/INV_3  ( .I(\SB1_1_13/buf_output[3] ), .ZN(\SB2_1_11/i0[8] ) );
  INV_X1 \SB2_1_12/INV_4  ( .I(\SB1_1_13/buf_output[4] ), .ZN(\SB2_1_12/i0[7] ) );
  INV_X2 \SB2_1_12/INV_3  ( .I(\SB1_1_14/buf_output[3] ), .ZN(\SB2_1_12/i0[8] ) );
  INV_X1 \SB2_1_13/INV_4  ( .I(\SB1_1_14/buf_output[4] ), .ZN(\SB2_1_13/i0[7] ) );
  INV_X1 \SB2_1_14/INV_4  ( .I(\SB1_1_15/buf_output[4] ), .ZN(\SB2_1_14/i0[7] ) );
  INV_X1 \SB2_1_14/INV_1  ( .I(\SB1_1_18/buf_output[1] ), .ZN(\SB2_1_14/i1_7 )
         );
  INV_X2 \SB2_1_15/INV_3  ( .I(\SB1_1_17/buf_output[3] ), .ZN(\SB2_1_15/i0[8] ) );
  INV_X1 \SB2_1_15/INV_1  ( .I(\SB1_1_19/buf_output[1] ), .ZN(\SB2_1_15/i1_7 )
         );
  INV_X1 \SB2_1_16/INV_4  ( .I(\SB1_1_17/buf_output[4] ), .ZN(\SB2_1_16/i0[7] ) );
  INV_X1 \SB2_1_16/INV_0  ( .I(\SB1_1_21/buf_output[0] ), .ZN(\SB2_1_16/i3[0] ) );
  INV_X1 \SB2_1_17/INV_4  ( .I(\SB1_1_18/buf_output[4] ), .ZN(\SB2_1_17/i0[7] ) );
  INV_X1 \SB2_1_19/INV_0  ( .I(\SB1_1_24/buf_output[0] ), .ZN(\SB2_1_19/i3[0] ) );
  INV_X1 \SB2_1_20/INV_4  ( .I(\SB1_1_21/buf_output[4] ), .ZN(\SB2_1_20/i0[7] ) );
  INV_X1 \SB2_1_20/INV_0  ( .I(\SB1_1_25/buf_output[0] ), .ZN(\SB2_1_20/i3[0] ) );
  INV_X1 \SB2_1_21/INV_4  ( .I(\SB1_1_22/buf_output[4] ), .ZN(\SB2_1_21/i0[7] ) );
  INV_X1 \SB2_1_22/INV_4  ( .I(\SB1_1_23/buf_output[4] ), .ZN(\SB2_1_22/i0[7] ) );
  INV_X1 \SB2_1_22/INV_0  ( .I(\SB1_1_27/buf_output[0] ), .ZN(\SB2_1_22/i3[0] ) );
  INV_X1 \SB2_1_23/INV_4  ( .I(\SB1_1_24/buf_output[4] ), .ZN(\SB2_1_23/i0[7] ) );
  INV_X2 \SB2_1_23/INV_3  ( .I(\SB1_1_25/buf_output[3] ), .ZN(\SB2_1_23/i0[8] ) );
  INV_X1 \SB2_1_24/INV_4  ( .I(\SB1_1_25/buf_output[4] ), .ZN(\SB2_1_24/i0[7] ) );
  INV_X1 \SB2_1_24/INV_0  ( .I(\SB1_1_29/buf_output[0] ), .ZN(\SB2_1_24/i3[0] ) );
  INV_X1 \SB2_1_25/INV_0  ( .I(\SB1_1_30/buf_output[0] ), .ZN(\SB2_1_25/i3[0] ) );
  INV_X1 \SB2_1_26/INV_4  ( .I(\SB1_1_27/buf_output[4] ), .ZN(\SB2_1_26/i0[7] ) );
  INV_X1 \SB2_1_26/INV_0  ( .I(\SB1_1_31/buf_output[0] ), .ZN(\SB2_1_26/i3[0] ) );
  INV_X1 \SB2_1_27/INV_4  ( .I(\SB1_1_28/buf_output[4] ), .ZN(\SB2_1_27/i0[7] ) );
  INV_X1 \SB2_1_28/INV_4  ( .I(\SB1_1_29/buf_output[4] ), .ZN(\SB2_1_28/i0[7] ) );
  INV_X1 \SB2_1_28/INV_0  ( .I(\SB1_1_1/buf_output[0] ), .ZN(\SB2_1_28/i3[0] )
         );
  INV_X1 \SB2_1_30/INV_1  ( .I(\SB1_1_2/buf_output[1] ), .ZN(\SB2_1_30/i1_7 )
         );
  INV_X1 \SB2_1_30/INV_0  ( .I(\SB1_1_3/buf_output[0] ), .ZN(\SB2_1_30/i3[0] )
         );
  INV_X1 \SB2_1_31/INV_1  ( .I(\SB1_1_3/buf_output[1] ), .ZN(\SB2_1_31/i1_7 )
         );
  INV_X1 \SB1_2_0/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[190] ), .ZN(
        \SB1_2_0/i0[7] ) );
  INV_X2 \SB1_2_0/INV_3  ( .I(n1373), .ZN(\SB1_2_0/i0[8] ) );
  INV_X1 \SB1_2_1/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[184] ), .ZN(
        \SB1_2_1/i0[7] ) );
  INV_X1 \SB1_2_2/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[178] ), .ZN(
        \SB1_2_2/i0[7] ) );
  INV_X2 \SB1_2_2/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[177] ), .ZN(
        \SB1_2_2/i0[8] ) );
  INV_X1 \SB1_2_3/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[172] ), .ZN(
        \SB1_2_3/i0[7] ) );
  INV_X2 \SB1_2_3/INV_2  ( .I(n5487), .ZN(\SB1_2_3/i1[9] ) );
  INV_X1 \SB1_2_4/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[166] ), .ZN(
        \SB1_2_4/i0[7] ) );
  INV_X2 \SB1_2_4/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[165] ), .ZN(
        \SB1_2_4/i0[8] ) );
  INV_X1 \SB1_2_5/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[160] ), .ZN(
        \SB1_2_5/i0[7] ) );
  INV_X1 \SB1_2_6/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[154] ), .ZN(
        \SB1_2_6/i0[7] ) );
  INV_X1 \SB1_2_7/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[148] ), .ZN(
        \SB1_2_7/i0[7] ) );
  INV_X2 \SB1_2_7/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[147] ), .ZN(
        \SB1_2_7/i0[8] ) );
  INV_X2 \SB1_2_8/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[141] ), .ZN(
        \SB1_2_8/i0[8] ) );
  INV_X2 \SB1_2_8/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[140] ), .ZN(
        \SB1_2_8/i1[9] ) );
  INV_X1 \SB1_2_9/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[136] ), .ZN(
        \SB1_2_9/i0[7] ) );
  INV_X2 \SB1_2_9/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[135] ), .ZN(
        \SB1_2_9/i0[8] ) );
  INV_X1 \SB1_2_10/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[130] ), .ZN(
        \SB1_2_10/i0[7] ) );
  INV_X2 \SB1_2_10/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[129] ), .ZN(
        \SB1_2_10/i0[8] ) );
  INV_X1 \SB1_2_11/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[124] ), .ZN(
        \SB1_2_11/i0[7] ) );
  INV_X1 \SB1_2_12/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[118] ), .ZN(
        \SB1_2_12/i0[7] ) );
  INV_X1 \SB1_2_13/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[112] ), .ZN(
        \SB1_2_13/i0[7] ) );
  INV_X2 \SB1_2_13/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[111] ), .ZN(
        \SB1_2_13/i0[8] ) );
  INV_X1 \SB1_2_14/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[106] ), .ZN(
        \SB1_2_14/i0[7] ) );
  INV_X1 \SB1_2_15/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[100] ), .ZN(
        \SB1_2_15/i0[7] ) );
  INV_X2 \SB1_2_15/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[99] ), .ZN(
        \SB1_2_15/i0[8] ) );
  INV_X1 \SB1_2_16/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[94] ), .ZN(
        \SB1_2_16/i0[7] ) );
  INV_X2 \SB1_2_16/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[93] ), .ZN(
        \SB1_2_16/i0[8] ) );
  INV_X2 \SB1_2_16/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[92] ), .ZN(
        \SB1_2_16/i1[9] ) );
  INV_X1 \SB1_2_17/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[88] ), .ZN(
        \SB1_2_17/i0[7] ) );
  INV_X2 \SB1_2_17/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[87] ), .ZN(
        \SB1_2_17/i0[8] ) );
  INV_X1 \SB1_2_18/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[82] ), .ZN(
        \SB1_2_18/i0[7] ) );
  INV_X2 \SB1_2_18/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[80] ), .ZN(
        \SB1_2_18/i1[9] ) );
  INV_X1 \SB1_2_19/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[76] ), .ZN(
        \SB1_2_19/i0[7] ) );
  INV_X2 \SB1_2_19/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[75] ), .ZN(
        \SB1_2_19/i0[8] ) );
  INV_X1 \SB1_2_19/INV_1  ( .I(\MC_ARK_ARC_1_1/buf_output[73] ), .ZN(
        \SB1_2_19/i1_7 ) );
  INV_X1 \SB1_2_19/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[72] ), .ZN(
        \SB1_2_19/i3[0] ) );
  INV_X1 \SB1_2_20/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[70] ), .ZN(
        \SB1_2_20/i0[7] ) );
  INV_X1 \SB1_2_21/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[64] ), .ZN(
        \SB1_2_21/i0[7] ) );
  INV_X1 \SB1_2_22/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[58] ), .ZN(
        \SB1_2_22/i0[7] ) );
  INV_X2 \SB1_2_22/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[57] ), .ZN(
        \SB1_2_22/i0[8] ) );
  INV_X2 \SB1_2_22/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[56] ), .ZN(
        \SB1_2_22/i1[9] ) );
  INV_X1 \SB1_2_22/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[54] ), .ZN(
        \SB1_2_22/i3[0] ) );
  INV_X1 \SB1_2_23/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[52] ), .ZN(
        \SB1_2_23/i0[7] ) );
  INV_X1 \SB1_2_23/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[48] ), .ZN(
        \SB1_2_23/i3[0] ) );
  INV_X1 \SB1_2_24/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[46] ), .ZN(
        \SB1_2_24/i0[7] ) );
  INV_X2 \SB1_2_24/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[45] ), .ZN(
        \SB1_2_24/i0[8] ) );
  INV_X1 \SB1_2_25/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[40] ), .ZN(
        \SB1_2_25/i0[7] ) );
  INV_X2 \SB1_2_25/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[39] ), .ZN(
        \SB1_2_25/i0[8] ) );
  INV_X1 \SB1_2_26/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[34] ), .ZN(
        \SB1_2_26/i0[7] ) );
  INV_X1 \SB1_2_26/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[30] ), .ZN(
        \SB1_2_26/i3[0] ) );
  INV_X1 \SB1_2_27/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[28] ), .ZN(
        \SB1_2_27/i0[7] ) );
  INV_X1 \SB1_2_27/INV_1  ( .I(\MC_ARK_ARC_1_1/buf_output[25] ), .ZN(
        \SB1_2_27/i1_7 ) );
  INV_X1 \SB1_2_27/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[24] ), .ZN(
        \SB1_2_27/i3[0] ) );
  INV_X1 \SB1_2_28/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[22] ), .ZN(
        \SB1_2_28/i0[7] ) );
  INV_X1 \SB1_2_29/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[16] ), .ZN(
        \SB1_2_29/i0[7] ) );
  INV_X1 \SB1_2_29/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[12] ), .ZN(
        \SB1_2_29/i3[0] ) );
  INV_X1 \SB1_2_30/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[10] ), .ZN(
        \SB1_2_30/i0[7] ) );
  INV_X2 \SB1_2_30/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[9] ), .ZN(
        \SB1_2_30/i0[8] ) );
  INV_X2 \SB1_2_30/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[8] ), .ZN(
        \SB1_2_30/i1[9] ) );
  INV_X1 \SB1_2_31/INV_4  ( .I(\MC_ARK_ARC_1_1/buf_output[4] ), .ZN(
        \SB1_2_31/i0[7] ) );
  INV_X2 \SB1_2_31/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[3] ), .ZN(
        \SB1_2_31/i0[8] ) );
  INV_X1 \SB2_2_0/INV_4  ( .I(\SB1_2_1/buf_output[4] ), .ZN(\SB2_2_0/i0[7] )
         );
  INV_X2 \SB2_2_0/INV_3  ( .I(\SB1_2_2/buf_output[3] ), .ZN(\SB2_2_0/i0[8] )
         );
  INV_X1 \SB2_2_0/INV_0  ( .I(\SB1_2_5/buf_output[0] ), .ZN(\SB2_2_0/i3[0] )
         );
  INV_X1 \SB2_2_1/INV_0  ( .I(\SB1_2_6/buf_output[0] ), .ZN(\SB2_2_1/i3[0] )
         );
  INV_X1 \SB2_2_2/INV_4  ( .I(\SB1_2_3/buf_output[4] ), .ZN(\SB2_2_2/i0[7] )
         );
  INV_X1 \SB2_2_2/INV_0  ( .I(\SB1_2_7/buf_output[0] ), .ZN(\SB2_2_2/i3[0] )
         );
  INV_X1 \SB2_2_4/INV_0  ( .I(\SB1_2_9/buf_output[0] ), .ZN(\SB2_2_4/i3[0] )
         );
  INV_X1 \SB2_2_5/INV_0  ( .I(\SB1_2_10/buf_output[0] ), .ZN(\SB2_2_5/i3[0] )
         );
  INV_X1 \SB2_2_6/INV_4  ( .I(\SB1_2_7/buf_output[4] ), .ZN(\SB2_2_6/i0[7] )
         );
  INV_X2 \SB2_2_7/INV_3  ( .I(\SB1_2_9/buf_output[3] ), .ZN(\SB2_2_7/i0[8] )
         );
  INV_X1 \SB2_2_7/INV_0  ( .I(\SB1_2_12/buf_output[0] ), .ZN(\SB2_2_7/i3[0] )
         );
  INV_X1 \SB2_2_9/INV_0  ( .I(\SB1_2_14/buf_output[0] ), .ZN(\SB2_2_9/i3[0] )
         );
  INV_X1 \SB2_2_10/INV_0  ( .I(\SB1_2_15/buf_output[0] ), .ZN(\SB2_2_10/i3[0] ) );
  INV_X1 \SB2_2_11/INV_4  ( .I(\SB1_2_12/buf_output[4] ), .ZN(\SB2_2_11/i0[7] ) );
  INV_X1 \SB2_2_11/INV_0  ( .I(\SB1_2_16/buf_output[0] ), .ZN(\SB2_2_11/i3[0] ) );
  INV_X1 \SB2_2_12/INV_4  ( .I(\SB1_2_13/buf_output[4] ), .ZN(\SB2_2_12/i0[7] ) );
  INV_X1 \SB2_2_12/INV_0  ( .I(\SB1_2_17/buf_output[0] ), .ZN(\SB2_2_12/i3[0] ) );
  INV_X2 \SB2_2_13/INV_3  ( .I(\SB1_2_15/buf_output[3] ), .ZN(\SB2_2_13/i0[8] ) );
  INV_X1 \SB2_2_14/INV_1  ( .I(\SB1_2_18/buf_output[1] ), .ZN(\SB2_2_14/i1_7 )
         );
  INV_X1 \SB2_2_14/INV_0  ( .I(\SB1_2_19/buf_output[0] ), .ZN(\SB2_2_14/i3[0] ) );
  INV_X1 \SB2_2_15/INV_0  ( .I(\SB1_2_20/buf_output[0] ), .ZN(\SB2_2_15/i3[0] ) );
  INV_X1 \SB2_2_16/INV_4  ( .I(\SB1_2_17/buf_output[4] ), .ZN(\SB2_2_16/i0[7] ) );
  INV_X1 \SB2_2_16/INV_0  ( .I(\SB1_2_21/buf_output[0] ), .ZN(\SB2_2_16/i3[0] ) );
  INV_X1 \SB2_2_17/INV_4  ( .I(\SB1_2_18/buf_output[4] ), .ZN(\SB2_2_17/i0[7] ) );
  INV_X1 \SB2_2_17/INV_1  ( .I(\SB1_2_21/buf_output[1] ), .ZN(\SB2_2_17/i1_7 )
         );
  INV_X1 \SB2_2_17/INV_0  ( .I(\SB1_2_22/buf_output[0] ), .ZN(\SB2_2_17/i3[0] ) );
  INV_X1 \SB2_2_18/INV_4  ( .I(\SB1_2_19/buf_output[4] ), .ZN(\SB2_2_18/i0[7] ) );
  INV_X1 \SB2_2_18/INV_0  ( .I(\SB1_2_23/buf_output[0] ), .ZN(\SB2_2_18/i3[0] ) );
  INV_X1 \SB2_2_19/INV_4  ( .I(\SB1_2_20/buf_output[4] ), .ZN(\SB2_2_19/i0[7] ) );
  INV_X2 \SB2_2_19/INV_3  ( .I(\SB1_2_21/buf_output[3] ), .ZN(\SB2_2_19/i0[8] ) );
  INV_X1 \SB2_2_19/INV_0  ( .I(\SB1_2_24/buf_output[0] ), .ZN(\SB2_2_19/i3[0] ) );
  INV_X1 \SB2_2_20/INV_4  ( .I(\SB1_2_21/buf_output[4] ), .ZN(\SB2_2_20/i0[7] ) );
  INV_X2 \SB2_2_20/INV_3  ( .I(\SB1_2_22/buf_output[3] ), .ZN(\SB2_2_20/i0[8] ) );
  INV_X1 \SB2_2_20/INV_0  ( .I(\SB1_2_25/buf_output[0] ), .ZN(\SB2_2_20/i3[0] ) );
  INV_X1 \SB2_2_21/INV_4  ( .I(\SB1_2_22/buf_output[4] ), .ZN(\SB2_2_21/i0[7] ) );
  INV_X1 \SB2_2_22/INV_4  ( .I(\SB1_2_23/buf_output[4] ), .ZN(\SB2_2_22/i0[7] ) );
  INV_X1 \SB2_2_22/INV_0  ( .I(\SB1_2_27/buf_output[0] ), .ZN(\SB2_2_22/i3[0] ) );
  INV_X1 \SB2_2_23/INV_4  ( .I(\SB1_2_24/buf_output[4] ), .ZN(\SB2_2_23/i0[7] ) );
  INV_X2 \SB2_2_23/INV_3  ( .I(\SB1_2_25/buf_output[3] ), .ZN(\SB2_2_23/i0[8] ) );
  INV_X1 \SB2_2_23/INV_0  ( .I(\SB1_2_28/buf_output[0] ), .ZN(\SB2_2_23/i3[0] ) );
  INV_X1 \SB2_2_24/INV_4  ( .I(\SB1_2_25/buf_output[4] ), .ZN(\SB2_2_24/i0[7] ) );
  INV_X1 \SB2_2_24/INV_0  ( .I(\SB1_2_29/buf_output[0] ), .ZN(\SB2_2_24/i3[0] ) );
  INV_X1 \SB2_2_25/INV_4  ( .I(\SB1_2_26/buf_output[4] ), .ZN(\SB2_2_25/i0[7] ) );
  INV_X2 \SB2_2_25/INV_3  ( .I(\SB1_2_27/buf_output[3] ), .ZN(\SB2_2_25/i0[8] ) );
  INV_X1 \SB2_2_25/INV_0  ( .I(\SB1_2_30/buf_output[0] ), .ZN(\SB2_2_25/i3[0] ) );
  INV_X1 \SB2_2_26/INV_4  ( .I(\SB1_2_27/buf_output[4] ), .ZN(\SB2_2_26/i0[7] ) );
  INV_X1 \SB2_2_28/INV_0  ( .I(\SB1_2_1/buf_output[0] ), .ZN(\SB2_2_28/i3[0] )
         );
  INV_X1 \SB2_2_29/INV_0  ( .I(\SB1_2_2/buf_output[0] ), .ZN(\SB2_2_29/i3[0] )
         );
  INV_X1 \SB2_2_30/INV_4  ( .I(\SB2_2_30/i0_4 ), .ZN(\SB2_2_30/i0[7] ) );
  INV_X1 \SB2_2_30/INV_0  ( .I(\SB1_2_3/buf_output[0] ), .ZN(\SB2_2_30/i3[0] )
         );
  INV_X1 \SB1_3_0/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[190] ), .ZN(
        \SB1_3_0/i0[7] ) );
  INV_X1 \SB1_3_0/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[186] ), .ZN(
        \SB1_3_0/i3[0] ) );
  INV_X1 \SB1_3_1/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[184] ), .ZN(
        \SB1_3_1/i0[7] ) );
  INV_X2 \SB1_3_1/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[183] ), .ZN(
        \SB1_3_1/i0[8] ) );
  INV_X1 \SB1_3_2/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[178] ), .ZN(
        \SB1_3_2/i0[7] ) );
  INV_X1 \SB1_3_3/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[172] ), .ZN(
        \SB1_3_3/i0[7] ) );
  INV_X1 \SB1_3_3/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[168] ), .ZN(
        \SB1_3_3/i3[0] ) );
  INV_X1 \SB1_3_4/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[166] ), .ZN(
        \SB1_3_4/i0[7] ) );
  INV_X2 \SB1_3_4/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[165] ), .ZN(
        \SB1_3_4/i0[8] ) );
  INV_X1 \SB1_3_5/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[160] ), .ZN(
        \SB1_3_5/i0[7] ) );
  INV_X1 \SB1_3_6/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[154] ), .ZN(
        \SB1_3_6/i0[7] ) );
  INV_X2 \SB1_3_6/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[153] ), .ZN(
        \SB1_3_6/i0[8] ) );
  INV_X1 \SB1_3_6/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[150] ), .ZN(
        \SB1_3_6/i3[0] ) );
  INV_X1 \SB1_3_7/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[148] ), .ZN(
        \SB1_3_7/i0[7] ) );
  INV_X1 \SB1_3_8/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[142] ), .ZN(
        \SB1_3_8/i0[7] ) );
  INV_X2 \SB1_3_8/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[141] ), .ZN(
        \SB1_3_8/i0[8] ) );
  INV_X2 \SB1_3_8/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[140] ), .ZN(
        \SB1_3_8/i1[9] ) );
  INV_X1 \SB1_3_8/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[138] ), .ZN(
        \SB1_3_8/i3[0] ) );
  INV_X1 \SB1_3_9/INV_5  ( .I(\MC_ARK_ARC_1_2/buf_output[137] ), .ZN(
        \SB1_3_9/i1_5 ) );
  INV_X1 \SB1_3_9/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[136] ), .ZN(
        \SB1_3_9/i0[7] ) );
  INV_X1 \SB1_3_9/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[132] ), .ZN(
        \SB1_3_9/i3[0] ) );
  INV_X1 \SB1_3_10/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[130] ), .ZN(
        \SB1_3_10/i0[7] ) );
  INV_X2 \SB1_3_10/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[129] ), .ZN(
        \SB1_3_10/i0[8] ) );
  INV_X1 \SB1_3_10/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[126] ), .ZN(
        \SB1_3_10/i3[0] ) );
  INV_X1 \SB1_3_12/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[114] ), .ZN(
        \SB1_3_12/i3[0] ) );
  INV_X1 \SB1_3_13/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[112] ), .ZN(
        \SB1_3_13/i0[7] ) );
  INV_X2 \SB1_3_13/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[111] ), .ZN(
        \SB1_3_13/i0[8] ) );
  INV_X2 \SB1_3_13/INV_2  ( .I(n5516), .ZN(\SB1_3_13/i1[9] ) );
  INV_X1 \SB1_3_13/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[108] ), .ZN(
        \SB1_3_13/i3[0] ) );
  INV_X1 \SB1_3_14/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[106] ), .ZN(
        \SB1_3_14/i0[7] ) );
  INV_X1 \SB1_3_15/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[100] ), .ZN(
        \SB1_3_15/i0[7] ) );
  INV_X2 \SB1_3_15/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[99] ), .ZN(
        \SB1_3_15/i0[8] ) );
  INV_X1 \SB1_3_16/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[94] ), .ZN(
        \SB1_3_16/i0[7] ) );
  INV_X1 \SB1_3_16/INV_1  ( .I(\MC_ARK_ARC_1_2/buf_output[91] ), .ZN(
        \SB1_3_16/i1_7 ) );
  INV_X1 \SB1_3_17/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[88] ), .ZN(
        \SB1_3_17/i0[7] ) );
  INV_X2 \SB1_3_17/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[87] ), .ZN(
        \SB1_3_17/i0[8] ) );
  INV_X1 \SB1_3_18/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[82] ), .ZN(
        \SB1_3_18/i0[7] ) );
  INV_X1 \SB1_3_18/INV_1  ( .I(\MC_ARK_ARC_1_2/buf_output[79] ), .ZN(
        \SB1_3_18/i1_7 ) );
  INV_X1 \SB1_3_19/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[76] ), .ZN(
        \SB1_3_19/i0[7] ) );
  INV_X2 \SB1_3_19/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[75] ), .ZN(
        \SB1_3_19/i0[8] ) );
  INV_X1 \SB1_3_19/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[72] ), .ZN(
        \SB1_3_19/i3[0] ) );
  INV_X1 \SB1_3_20/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[70] ), .ZN(
        \SB1_3_20/i0[7] ) );
  INV_X1 \SB1_3_20/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[66] ), .ZN(
        \SB1_3_20/i3[0] ) );
  INV_X2 \SB1_3_21/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[63] ), .ZN(
        \SB1_3_21/i0[8] ) );
  INV_X1 \SB1_3_22/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[58] ), .ZN(
        \SB1_3_22/i0[7] ) );
  INV_X2 \SB1_3_22/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[57] ), .ZN(
        \SB1_3_22/i0[8] ) );
  INV_X2 \SB1_3_22/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[56] ), .ZN(
        \SB1_3_22/i1[9] ) );
  INV_X2 \SB1_3_23/INV_3  ( .I(n5507), .ZN(\SB1_3_23/i0[8] ) );
  INV_X1 \SB1_3_24/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[46] ), .ZN(
        \SB1_3_24/i0[7] ) );
  INV_X2 \SB1_3_24/INV_3  ( .I(n3667), .ZN(\SB1_3_24/i0[8] ) );
  INV_X2 \SB1_3_24/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[44] ), .ZN(
        \SB1_3_24/i1[9] ) );
  INV_X1 \SB1_3_25/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[36] ), .ZN(
        \SB1_3_25/i3[0] ) );
  INV_X1 \SB1_3_26/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[34] ), .ZN(
        \SB1_3_26/i0[7] ) );
  INV_X1 \SB1_3_27/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[28] ), .ZN(
        \SB1_3_27/i0[7] ) );
  INV_X1 \SB1_3_28/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[22] ), .ZN(
        \SB1_3_28/i0[7] ) );
  INV_X1 \SB1_3_29/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[16] ), .ZN(
        \SB1_3_29/i0[7] ) );
  INV_X1 \SB1_3_30/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[10] ), .ZN(
        \SB1_3_30/i0[7] ) );
  INV_X1 \SB1_3_31/INV_4  ( .I(\MC_ARK_ARC_1_2/buf_output[4] ), .ZN(
        \SB1_3_31/i0[7] ) );
  INV_X2 \SB1_3_31/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[3] ), .ZN(
        \SB1_3_31/i0[8] ) );
  INV_X1 \SB2_3_0/INV_0  ( .I(\SB1_3_5/buf_output[0] ), .ZN(\SB2_3_0/i3[0] )
         );
  INV_X1 \SB2_3_1/INV_4  ( .I(\SB1_3_2/buf_output[4] ), .ZN(\SB2_3_1/i0[7] )
         );
  INV_X1 \SB2_3_1/INV_0  ( .I(\SB1_3_6/buf_output[0] ), .ZN(\SB2_3_1/i3[0] )
         );
  INV_X1 \SB2_3_2/INV_4  ( .I(\SB1_3_3/buf_output[4] ), .ZN(\SB2_3_2/i0[7] )
         );
  INV_X1 \SB2_3_2/INV_0  ( .I(\SB1_3_7/buf_output[0] ), .ZN(\SB2_3_2/i3[0] )
         );
  INV_X1 \SB2_3_3/INV_4  ( .I(\SB1_3_4/buf_output[4] ), .ZN(\SB2_3_3/i0[7] )
         );
  INV_X1 \SB2_3_4/INV_4  ( .I(\SB1_3_5/buf_output[4] ), .ZN(\SB2_3_4/i0[7] )
         );
  INV_X1 \SB2_3_5/INV_4  ( .I(\SB1_3_6/buf_output[4] ), .ZN(\SB2_3_5/i0[7] )
         );
  INV_X1 \SB2_3_5/INV_0  ( .I(\SB1_3_10/buf_output[0] ), .ZN(\SB2_3_5/i3[0] )
         );
  INV_X1 \SB2_3_6/INV_4  ( .I(\SB1_3_7/buf_output[4] ), .ZN(\SB2_3_6/i0[7] )
         );
  INV_X1 \SB2_3_6/INV_0  ( .I(\SB1_3_11/buf_output[0] ), .ZN(\SB2_3_6/i3[0] )
         );
  INV_X2 \SB2_3_8/INV_3  ( .I(n3685), .ZN(\SB2_3_8/i0[8] ) );
  INV_X1 \SB2_3_8/INV_0  ( .I(\SB1_3_13/buf_output[0] ), .ZN(\SB2_3_8/i3[0] )
         );
  INV_X1 \SB2_3_9/INV_4  ( .I(\SB1_3_10/buf_output[4] ), .ZN(\SB2_3_9/i0[7] )
         );
  INV_X2 \SB2_3_9/INV_2  ( .I(\SB1_3_12/buf_output[2] ), .ZN(\SB2_3_9/i1[9] )
         );
  INV_X1 \SB2_3_9/INV_0  ( .I(\SB1_3_14/buf_output[0] ), .ZN(\SB2_3_9/i3[0] )
         );
  INV_X1 \SB2_3_10/INV_4  ( .I(\SB1_3_11/buf_output[4] ), .ZN(\SB2_3_10/i0[7] ) );
  INV_X1 \SB2_3_10/INV_1  ( .I(\SB1_3_14/buf_output[1] ), .ZN(\SB2_3_10/i1_7 )
         );
  INV_X1 \SB2_3_10/INV_0  ( .I(\SB1_3_15/buf_output[0] ), .ZN(\SB2_3_10/i3[0] ) );
  INV_X1 \SB2_3_11/INV_0  ( .I(\SB1_3_16/buf_output[0] ), .ZN(\SB2_3_11/i3[0] ) );
  INV_X1 \SB2_3_12/INV_4  ( .I(\SB1_3_13/buf_output[4] ), .ZN(\SB2_3_12/i0[7] ) );
  INV_X1 \SB2_3_13/INV_0  ( .I(\SB1_3_18/buf_output[0] ), .ZN(\SB2_3_13/i3[0] ) );
  INV_X1 \SB2_3_14/INV_4  ( .I(\SB1_3_15/buf_output[4] ), .ZN(\SB2_3_14/i0[7] ) );
  INV_X1 \SB2_3_14/INV_0  ( .I(\SB1_3_19/buf_output[0] ), .ZN(\SB2_3_14/i3[0] ) );
  INV_X1 \SB2_3_15/INV_0  ( .I(\SB1_3_20/buf_output[0] ), .ZN(\SB2_3_15/i3[0] ) );
  INV_X1 \SB2_3_16/INV_4  ( .I(\SB1_3_17/buf_output[4] ), .ZN(\SB2_3_16/i0[7] ) );
  INV_X2 \SB2_3_16/INV_3  ( .I(\SB1_3_18/buf_output[3] ), .ZN(\SB2_3_16/i0[8] ) );
  INV_X1 \SB2_3_17/INV_0  ( .I(\SB1_3_22/buf_output[0] ), .ZN(\SB2_3_17/i3[0] ) );
  INV_X1 \SB2_3_18/INV_4  ( .I(\SB1_3_19/buf_output[4] ), .ZN(\SB2_3_18/i0[7] ) );
  INV_X1 \SB2_3_19/INV_4  ( .I(\SB1_3_20/buf_output[4] ), .ZN(\SB2_3_19/i0[7] ) );
  INV_X1 \SB2_3_19/INV_1  ( .I(\SB1_3_23/buf_output[1] ), .ZN(\SB2_3_19/i1_7 )
         );
  INV_X1 \SB2_3_20/INV_0  ( .I(\SB1_3_25/buf_output[0] ), .ZN(\SB2_3_20/i3[0] ) );
  INV_X1 \SB2_3_21/INV_4  ( .I(\SB1_3_22/buf_output[4] ), .ZN(\SB2_3_21/i0[7] ) );
  INV_X1 \SB2_3_21/INV_1  ( .I(\SB1_3_25/buf_output[1] ), .ZN(\SB2_3_21/i1_7 )
         );
  INV_X1 \SB2_3_21/INV_0  ( .I(\SB1_3_26/buf_output[0] ), .ZN(\SB2_3_21/i3[0] ) );
  INV_X1 \SB2_3_22/INV_4  ( .I(\SB1_3_23/buf_output[4] ), .ZN(\SB2_3_22/i0[7] ) );
  INV_X1 \SB2_3_22/INV_0  ( .I(\SB1_3_27/buf_output[0] ), .ZN(\SB2_3_22/i3[0] ) );
  INV_X1 \SB2_3_23/INV_4  ( .I(\SB1_3_24/buf_output[4] ), .ZN(\SB2_3_23/i0[7] ) );
  INV_X1 \SB2_3_24/INV_0  ( .I(\SB1_3_29/buf_output[0] ), .ZN(\SB2_3_24/i3[0] ) );
  INV_X2 \SB2_3_25/INV_3  ( .I(\SB1_3_27/buf_output[3] ), .ZN(\SB2_3_25/i0[8] ) );
  INV_X1 \SB2_3_27/INV_4  ( .I(\SB1_3_28/buf_output[4] ), .ZN(\SB2_3_27/i0[7] ) );
  INV_X2 \SB2_3_28/INV_3  ( .I(\SB1_3_30/buf_output[3] ), .ZN(\SB2_3_28/i0[8] ) );
  INV_X1 \SB2_3_28/INV_0  ( .I(\SB1_3_1/buf_output[0] ), .ZN(\SB2_3_28/i3[0] )
         );
  INV_X1 \SB2_3_29/INV_0  ( .I(\SB1_3_2/buf_output[0] ), .ZN(\SB2_3_29/i3[0] )
         );
  INV_X1 \SB2_3_30/INV_4  ( .I(\SB1_3_31/buf_output[4] ), .ZN(\SB2_3_30/i0[7] ) );
  INV_X1 \SB2_3_30/INV_0  ( .I(\SB1_3_3/buf_output[0] ), .ZN(\SB2_3_30/i3[0] )
         );
  INV_X1 \SB2_3_31/INV_4  ( .I(\SB1_3_0/buf_output[4] ), .ZN(\SB2_3_31/i0[7] )
         );
  INV_X1 \SB3_1/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[184] ), .ZN(
        \SB3_1/i0[7] ) );
  INV_X1 \SB3_1/INV_1  ( .I(\MC_ARK_ARC_1_3/buf_output[181] ), .ZN(
        \SB3_1/i1_7 ) );
  INV_X1 \SB3_2/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[178] ), .ZN(
        \SB3_2/i0[7] ) );
  INV_X1 \SB3_3/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[172] ), .ZN(
        \SB3_3/i0[7] ) );
  INV_X1 \SB3_3/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[168] ), .ZN(
        \SB3_3/i3[0] ) );
  INV_X1 \SB3_4/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[166] ), .ZN(
        \SB3_4/i0[7] ) );
  INV_X1 \SB3_5/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[160] ), .ZN(
        \SB3_5/i0[7] ) );
  INV_X1 \SB3_5/INV_1  ( .I(\MC_ARK_ARC_1_3/buf_output[157] ), .ZN(
        \SB3_5/i1_7 ) );
  INV_X1 \SB3_5/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[156] ), .ZN(
        \SB3_5/i3[0] ) );
  INV_X1 \SB3_7/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[148] ), .ZN(
        \SB3_7/i0[7] ) );
  INV_X1 \SB3_7/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[144] ), .ZN(
        \SB3_7/i3[0] ) );
  INV_X1 \SB3_8/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[142] ), .ZN(
        \SB3_8/i0[7] ) );
  INV_X1 \SB3_8/INV_1  ( .I(\MC_ARK_ARC_1_3/buf_output[139] ), .ZN(
        \SB3_8/i1_7 ) );
  INV_X1 \SB3_8/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[138] ), .ZN(
        \SB3_8/i3[0] ) );
  INV_X1 \SB3_9/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[136] ), .ZN(
        \SB3_9/i0[7] ) );
  INV_X1 \SB3_9/INV_1  ( .I(\MC_ARK_ARC_1_3/buf_output[133] ), .ZN(
        \SB3_9/i1_7 ) );
  INV_X1 \SB3_9/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[132] ), .ZN(
        \SB3_9/i3[0] ) );
  INV_X1 \SB3_10/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[130] ), .ZN(
        \SB3_10/i0[7] ) );
  INV_X1 \SB3_11/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[124] ), .ZN(
        \SB3_11/i0[7] ) );
  INV_X1 \SB3_11/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[120] ), .ZN(
        \SB3_11/i3[0] ) );
  INV_X1 \SB3_12/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[118] ), .ZN(
        \SB3_12/i0[7] ) );
  INV_X1 \SB3_12/INV_1  ( .I(\MC_ARK_ARC_1_3/buf_output[115] ), .ZN(
        \SB3_12/i1_7 ) );
  INV_X1 \SB3_13/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[112] ), .ZN(
        \SB3_13/i0[7] ) );
  INV_X1 \SB3_14/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[106] ), .ZN(
        \SB3_14/i0[7] ) );
  INV_X1 \SB3_14/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[102] ), .ZN(
        \SB3_14/i3[0] ) );
  INV_X1 \SB3_15/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[100] ), .ZN(
        \SB3_15/i0[7] ) );
  INV_X2 \SB3_15/INV_2  ( .I(\MC_ARK_ARC_1_3/buf_output[98] ), .ZN(
        \SB3_15/i1[9] ) );
  INV_X1 \SB3_15/INV_1  ( .I(\MC_ARK_ARC_1_3/buf_output[97] ), .ZN(
        \SB3_15/i1_7 ) );
  INV_X1 \SB3_15/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[96] ), .ZN(
        \SB3_15/i3[0] ) );
  INV_X1 \SB3_16/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[94] ), .ZN(
        \SB3_16/i0[7] ) );
  INV_X1 \SB3_17/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[88] ), .ZN(
        \SB3_17/i0[7] ) );
  INV_X1 \SB3_17/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[84] ), .ZN(
        \SB3_17/i3[0] ) );
  INV_X1 \SB3_18/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[82] ), .ZN(
        \SB3_18/i0[7] ) );
  INV_X1 \SB3_19/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[76] ), .ZN(
        \SB3_19/i0[7] ) );
  INV_X1 \SB3_19/INV_1  ( .I(\MC_ARK_ARC_1_3/buf_output[73] ), .ZN(
        \SB3_19/i1_7 ) );
  INV_X1 \SB3_20/INV_5  ( .I(\MC_ARK_ARC_1_3/buf_output[71] ), .ZN(
        \SB3_20/i1_5 ) );
  INV_X1 \SB3_20/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[70] ), .ZN(
        \SB3_20/i0[7] ) );
  INV_X1 \SB3_20/INV_1  ( .I(\MC_ARK_ARC_1_3/buf_output[67] ), .ZN(
        \SB3_20/i1_7 ) );
  INV_X1 \SB3_21/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[64] ), .ZN(
        \SB3_21/i0[7] ) );
  INV_X1 \SB3_22/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[58] ), .ZN(
        \SB3_22/i0[7] ) );
  INV_X2 \SB3_22/INV_2  ( .I(\MC_ARK_ARC_1_3/buf_output[56] ), .ZN(
        \SB3_22/i1[9] ) );
  INV_X1 \SB3_22/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[54] ), .ZN(
        \SB3_22/i3[0] ) );
  INV_X1 \SB3_23/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[52] ), .ZN(
        \SB3_23/i0[7] ) );
  INV_X1 \SB3_24/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[46] ), .ZN(
        \SB3_24/i0[7] ) );
  INV_X1 \SB3_24/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[42] ), .ZN(
        \SB3_24/i3[0] ) );
  INV_X1 \SB3_25/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[40] ), .ZN(
        \SB3_25/i0[7] ) );
  INV_X1 \SB3_25/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[36] ), .ZN(
        \SB3_25/i3[0] ) );
  INV_X1 \SB3_26/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[34] ), .ZN(
        \SB3_26/i0[7] ) );
  INV_X1 \SB3_26/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[30] ), .ZN(
        \SB3_26/i3[0] ) );
  INV_X1 \SB3_27/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[28] ), .ZN(
        \SB3_27/i0[7] ) );
  INV_X1 \SB3_27/INV_1  ( .I(\MC_ARK_ARC_1_3/buf_output[25] ), .ZN(
        \SB3_27/i1_7 ) );
  INV_X1 \SB3_27/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[24] ), .ZN(
        \SB3_27/i3[0] ) );
  INV_X1 \SB3_28/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[22] ), .ZN(
        \SB3_28/i0[7] ) );
  INV_X1 \SB3_28/INV_1  ( .I(\MC_ARK_ARC_1_3/buf_output[19] ), .ZN(
        \SB3_28/i1_7 ) );
  INV_X1 \SB3_28/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[18] ), .ZN(
        \SB3_28/i3[0] ) );
  INV_X1 \SB3_29/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[16] ), .ZN(
        \SB3_29/i0[7] ) );
  INV_X1 \SB3_29/INV_1  ( .I(\MC_ARK_ARC_1_3/buf_output[13] ), .ZN(
        \SB3_29/i1_7 ) );
  INV_X1 \SB3_29/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[12] ), .ZN(
        \SB3_29/i3[0] ) );
  INV_X1 \SB3_30/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[10] ), .ZN(
        \SB3_30/i0[7] ) );
  INV_X2 \SB3_30/INV_2  ( .I(\MC_ARK_ARC_1_3/buf_output[8] ), .ZN(
        \SB3_30/i1[9] ) );
  INV_X1 \SB3_31/INV_4  ( .I(\MC_ARK_ARC_1_3/buf_output[4] ), .ZN(
        \SB3_31/i0[7] ) );
  INV_X1 \SB3_31/INV_1  ( .I(\MC_ARK_ARC_1_3/buf_output[1] ), .ZN(
        \SB3_31/i1_7 ) );
  INV_X1 \SB4_0/INV_4  ( .I(\SB3_1/buf_output[4] ), .ZN(\SB4_0/i0[7] ) );
  INV_X2 \SB4_0/INV_3  ( .I(\SB3_2/buf_output[3] ), .ZN(\SB4_0/i0[8] ) );
  INV_X1 \SB4_0/INV_1  ( .I(\SB3_4/buf_output[1] ), .ZN(\SB4_0/i1_7 ) );
  INV_X1 \SB4_0/INV_0  ( .I(\SB3_5/buf_output[0] ), .ZN(\SB4_0/i3[0] ) );
  INV_X1 \SB4_1/INV_4  ( .I(\SB3_2/buf_output[4] ), .ZN(\SB4_1/i0[7] ) );
  INV_X1 \SB4_2/INV_4  ( .I(\SB3_3/buf_output[4] ), .ZN(\SB4_2/i0[7] ) );
  INV_X1 \SB4_3/INV_4  ( .I(\SB3_4/buf_output[4] ), .ZN(\SB4_3/i0[7] ) );
  INV_X1 \SB4_3/INV_1  ( .I(\SB3_7/buf_output[1] ), .ZN(\SB4_3/i1_7 ) );
  INV_X1 \SB4_3/INV_0  ( .I(\SB3_8/buf_output[0] ), .ZN(\SB4_3/i3[0] ) );
  INV_X1 \SB4_4/INV_4  ( .I(\SB3_5/buf_output[4] ), .ZN(\SB4_4/i0[7] ) );
  INV_X1 \SB4_4/INV_0  ( .I(\SB3_9/buf_output[0] ), .ZN(\SB4_4/i3[0] ) );
  INV_X1 \SB4_5/INV_4  ( .I(\SB3_6/buf_output[4] ), .ZN(\SB4_5/i0[7] ) );
  INV_X1 \SB4_5/INV_1  ( .I(\SB3_9/buf_output[1] ), .ZN(\SB4_5/i1_7 ) );
  INV_X1 \SB4_5/INV_0  ( .I(\SB3_10/buf_output[0] ), .ZN(\SB4_5/i3[0] ) );
  INV_X1 \SB4_6/INV_4  ( .I(\SB3_7/buf_output[4] ), .ZN(\SB4_6/i0[7] ) );
  INV_X1 \SB4_6/INV_0  ( .I(\SB3_11/buf_output[0] ), .ZN(\SB4_6/i3[0] ) );
  INV_X1 \SB4_7/INV_4  ( .I(\SB3_8/buf_output[4] ), .ZN(\SB4_7/i0[7] ) );
  INV_X1 \SB4_7/INV_0  ( .I(\SB3_12/buf_output[0] ), .ZN(\SB4_7/i3[0] ) );
  INV_X1 \SB4_8/INV_4  ( .I(\SB3_9/buf_output[4] ), .ZN(\SB4_8/i0[7] ) );
  INV_X1 \SB4_8/INV_0  ( .I(\SB3_13/buf_output[0] ), .ZN(\SB4_8/i3[0] ) );
  INV_X1 \SB4_9/INV_4  ( .I(\SB3_10/buf_output[4] ), .ZN(\SB4_9/i0[7] ) );
  INV_X1 \SB4_9/INV_0  ( .I(\SB3_14/buf_output[0] ), .ZN(\SB4_9/i3[0] ) );
  INV_X1 \SB4_10/INV_4  ( .I(\SB3_11/buf_output[4] ), .ZN(\SB4_10/i0[7] ) );
  INV_X1 \SB4_12/INV_4  ( .I(\SB3_13/buf_output[4] ), .ZN(\SB4_12/i0[7] ) );
  INV_X1 \SB4_13/INV_4  ( .I(\SB3_14/buf_output[4] ), .ZN(\SB4_13/i0[7] ) );
  INV_X1 \SB4_13/INV_0  ( .I(\SB3_18/buf_output[0] ), .ZN(\SB4_13/i3[0] ) );
  INV_X1 \SB4_14/INV_4  ( .I(\SB3_15/buf_output[4] ), .ZN(\SB4_14/i0[7] ) );
  INV_X1 \SB4_15/INV_4  ( .I(\SB3_16/buf_output[4] ), .ZN(\SB4_15/i0[7] ) );
  INV_X1 \SB4_15/INV_0  ( .I(\SB3_20/buf_output[0] ), .ZN(\SB4_15/i3[0] ) );
  INV_X1 \SB4_16/INV_4  ( .I(\SB3_17/buf_output[4] ), .ZN(\SB4_16/i0[7] ) );
  INV_X1 \SB4_17/INV_4  ( .I(\SB3_18/buf_output[4] ), .ZN(\SB4_17/i0[7] ) );
  INV_X1 \SB4_18/INV_4  ( .I(\SB3_19/buf_output[4] ), .ZN(\SB4_18/i0[7] ) );
  INV_X1 \SB4_18/INV_0  ( .I(\SB3_23/buf_output[0] ), .ZN(\SB4_18/i3[0] ) );
  INV_X1 \SB4_19/INV_4  ( .I(\SB3_20/buf_output[4] ), .ZN(\SB4_19/i0[7] ) );
  INV_X1 \SB4_19/INV_0  ( .I(\SB3_24/buf_output[0] ), .ZN(\SB4_19/i3[0] ) );
  INV_X1 \SB4_20/INV_4  ( .I(\SB3_21/buf_output[4] ), .ZN(\SB4_20/i0[7] ) );
  INV_X1 \SB4_20/INV_0  ( .I(\SB3_25/buf_output[0] ), .ZN(\SB4_20/i3[0] ) );
  INV_X1 \SB4_21/INV_4  ( .I(\SB3_22/buf_output[4] ), .ZN(\SB4_21/i0[7] ) );
  INV_X1 \SB4_21/INV_0  ( .I(\SB3_26/buf_output[0] ), .ZN(\SB4_21/i3[0] ) );
  INV_X1 \SB4_22/INV_4  ( .I(\SB3_23/buf_output[4] ), .ZN(\SB4_22/i0[7] ) );
  INV_X1 \SB4_22/INV_0  ( .I(\SB3_27/buf_output[0] ), .ZN(\SB4_22/i3[0] ) );
  INV_X1 \SB4_23/INV_4  ( .I(\SB3_24/buf_output[4] ), .ZN(\SB4_23/i0[7] ) );
  INV_X1 \SB4_23/INV_1  ( .I(\SB3_27/buf_output[1] ), .ZN(\SB4_23/i1_7 ) );
  INV_X1 \SB4_24/INV_4  ( .I(\SB3_25/buf_output[4] ), .ZN(\SB4_24/i0[7] ) );
  INV_X1 \SB4_24/INV_0  ( .I(\SB3_29/buf_output[0] ), .ZN(\SB4_24/i3[0] ) );
  INV_X1 \SB4_25/INV_4  ( .I(\SB3_26/buf_output[4] ), .ZN(\SB4_25/i0[7] ) );
  INV_X1 \SB4_25/INV_0  ( .I(\SB3_30/buf_output[0] ), .ZN(\SB4_25/i3[0] ) );
  INV_X1 \SB4_26/INV_4  ( .I(\SB3_27/buf_output[4] ), .ZN(\SB4_26/i0[7] ) );
  INV_X2 \SB4_26/INV_3  ( .I(\SB3_28/buf_output[3] ), .ZN(\SB4_26/i0[8] ) );
  INV_X1 \SB4_26/INV_1  ( .I(\SB3_30/buf_output[1] ), .ZN(\SB4_26/i1_7 ) );
  INV_X1 \SB4_26/INV_0  ( .I(\SB3_31/buf_output[0] ), .ZN(\SB4_26/i3[0] ) );
  INV_X1 \SB4_27/INV_4  ( .I(\SB3_28/buf_output[4] ), .ZN(\SB4_27/i0[7] ) );
  INV_X1 \SB4_27/INV_0  ( .I(\SB3_0/buf_output[0] ), .ZN(\SB4_27/i3[0] ) );
  INV_X1 \SB4_28/INV_4  ( .I(\SB3_29/buf_output[4] ), .ZN(\SB4_28/i0[7] ) );
  INV_X1 \SB4_28/INV_1  ( .I(\SB3_0/buf_output[1] ), .ZN(\SB4_28/i1_7 ) );
  INV_X1 \SB4_29/INV_5  ( .I(\SB3_29/buf_output[5] ), .ZN(\SB4_29/i1_5 ) );
  INV_X1 \SB4_29/INV_0  ( .I(\SB3_2/buf_output[0] ), .ZN(\SB4_29/i3[0] ) );
  INV_X1 \SB4_30/INV_4  ( .I(\SB3_31/buf_output[4] ), .ZN(\SB4_30/i0[7] ) );
  INV_X1 \SB4_30/INV_0  ( .I(\SB3_3/buf_output[0] ), .ZN(\SB4_30/i3[0] ) );
  INV_X1 \SB4_31/INV_4  ( .I(\SB3_0/buf_output[4] ), .ZN(\SB4_31/i0[7] ) );
  NAND3_X1 \SB1_0_0/Component_Function_2/N1  ( .A1(\SB1_0_0/i1_5 ), .A2(
        \SB1_0_0/i0[10] ), .A3(\SB1_0_0/i1[9] ), .ZN(
        \SB1_0_0/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_0/Component_Function_3/N4  ( .A1(\SB1_0_0/i1_5 ), .A2(
        \SB1_0_0/i0[8] ), .A3(\SB1_0_0/i3[0] ), .ZN(
        \SB1_0_0/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_0/Component_Function_3/N2  ( .A1(\SB1_0_0/i0_0 ), .A2(
        \SB1_0_0/i0_3 ), .A3(\SB1_0_0/i0_4 ), .ZN(
        \SB1_0_0/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_0/Component_Function_4/N4  ( .A1(\SB1_0_0/i1[9] ), .A2(
        \SB1_0_0/i1_5 ), .A3(\SB1_0_0/i0_4 ), .ZN(
        \SB1_0_0/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_0/Component_Function_4/N2  ( .A1(\SB1_0_0/i3[0] ), .A2(
        \SB1_0_0/i0_0 ), .A3(\SB1_0_0/i1_7 ), .ZN(
        \SB1_0_0/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_0/Component_Function_4/N1  ( .A1(\SB1_0_0/i0[9] ), .A2(
        \SB1_0_0/i0_0 ), .A3(\SB1_0_0/i0[8] ), .ZN(
        \SB1_0_0/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_1/Component_Function_2/N4  ( .A1(\SB1_0_1/i1_5 ), .A2(
        \SB1_0_1/i0_0 ), .A3(\SB1_0_1/i0_4 ), .ZN(
        \SB1_0_1/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_1/Component_Function_2/N1  ( .A1(\SB1_0_1/i1_5 ), .A2(
        \SB1_0_1/i0[10] ), .A3(\SB1_0_1/i1[9] ), .ZN(
        \SB1_0_1/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_1/Component_Function_3/N3  ( .A1(\SB1_0_1/i1[9] ), .A2(
        \SB1_0_1/i1_7 ), .A3(\SB1_0_1/i0[10] ), .ZN(
        \SB1_0_1/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_1/Component_Function_4/N4  ( .A1(\SB1_0_1/i1[9] ), .A2(
        \SB1_0_1/i1_5 ), .A3(\SB1_0_1/i0_4 ), .ZN(
        \SB1_0_1/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_1/Component_Function_4/N3  ( .A1(\SB1_0_1/i0[9] ), .A2(
        \SB1_0_1/i0[10] ), .A3(\SB1_0_1/i0_3 ), .ZN(
        \SB1_0_1/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_1/Component_Function_4/N2  ( .A1(\SB1_0_1/i3[0] ), .A2(
        \SB1_0_1/i0_0 ), .A3(\SB1_0_1/i1_7 ), .ZN(
        \SB1_0_1/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_1/Component_Function_4/N1  ( .A1(\SB1_0_1/i0[9] ), .A2(
        \SB1_0_1/i0_0 ), .A3(\SB1_0_1/i0[8] ), .ZN(
        \SB1_0_1/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_2/Component_Function_3/N4  ( .A1(\SB1_0_2/i1_5 ), .A2(
        \SB1_0_2/i0[8] ), .A3(\SB1_0_2/i3[0] ), .ZN(
        \SB1_0_2/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_2/Component_Function_3/N3  ( .A1(\SB1_0_2/i1[9] ), .A2(
        \SB1_0_2/i1_7 ), .A3(\SB1_0_2/i0[10] ), .ZN(
        \SB1_0_2/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_2/Component_Function_4/N3  ( .A1(\SB1_0_2/i0[9] ), .A2(
        \SB1_0_2/i0[10] ), .A3(\SB1_0_2/i0_3 ), .ZN(
        \SB1_0_2/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_3/Component_Function_2/N4  ( .A1(\SB1_0_3/i1_5 ), .A2(
        \SB1_0_3/i0_0 ), .A3(\SB1_0_3/i0_4 ), .ZN(
        \SB1_0_3/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_3/Component_Function_2/N1  ( .A1(\SB1_0_3/i1_5 ), .A2(
        \SB1_0_3/i0[10] ), .A3(\SB1_0_3/i1[9] ), .ZN(
        \SB1_0_3/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_3/Component_Function_3/N4  ( .A1(\SB1_0_3/i1_5 ), .A2(
        \SB1_0_3/i0[8] ), .A3(\SB1_0_3/i3[0] ), .ZN(
        \SB1_0_3/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_3/Component_Function_4/N4  ( .A1(\SB1_0_3/i1[9] ), .A2(
        \SB1_0_3/i1_5 ), .A3(\SB1_0_3/i0_4 ), .ZN(
        \SB1_0_3/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_4/Component_Function_2/N4  ( .A1(\SB1_0_4/i1_5 ), .A2(
        \SB1_0_4/i0_0 ), .A3(\SB1_0_4/i0_4 ), .ZN(
        \SB1_0_4/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_4/Component_Function_2/N3  ( .A1(\SB1_0_4/i0_3 ), .A2(
        \SB1_0_4/i0[8] ), .A3(\SB1_0_4/i0[9] ), .ZN(
        \SB1_0_4/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_4/Component_Function_2/N2  ( .A1(\SB1_0_4/i0_3 ), .A2(
        \SB1_0_4/i0[10] ), .A3(\SB1_0_4/i0[6] ), .ZN(
        \SB1_0_4/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_4/Component_Function_2/N1  ( .A1(\SB1_0_4/i1_5 ), .A2(
        \SB1_0_4/i0[10] ), .A3(\SB1_0_4/i1[9] ), .ZN(
        \SB1_0_4/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_4/Component_Function_4/N4  ( .A1(\SB1_0_4/i1[9] ), .A2(
        \SB1_0_4/i1_5 ), .A3(\SB1_0_4/i0_4 ), .ZN(
        \SB1_0_4/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_4/Component_Function_4/N3  ( .A1(\SB1_0_4/i0[9] ), .A2(
        \SB1_0_4/i0[10] ), .A3(\SB1_0_4/i0_3 ), .ZN(
        \SB1_0_4/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_4/Component_Function_4/N2  ( .A1(\SB1_0_4/i3[0] ), .A2(
        \SB1_0_4/i0_0 ), .A3(\SB1_0_4/i1_7 ), .ZN(
        \SB1_0_4/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_4/Component_Function_4/N1  ( .A1(\SB1_0_4/i0[9] ), .A2(
        \SB1_0_4/i0_0 ), .A3(\SB1_0_4/i0[8] ), .ZN(
        \SB1_0_4/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_5/Component_Function_3/N4  ( .A1(\SB1_0_5/i1_5 ), .A2(
        \SB1_0_5/i0[8] ), .A3(\SB1_0_5/i3[0] ), .ZN(
        \SB1_0_5/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_5/Component_Function_3/N1  ( .A1(\SB1_0_5/i1[9] ), .A2(
        \SB1_0_5/i0_3 ), .A3(\SB1_0_5/i0[6] ), .ZN(
        \SB1_0_5/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_5/Component_Function_4/N4  ( .A1(\SB1_0_5/i1[9] ), .A2(
        \SB1_0_5/i1_5 ), .A3(\SB1_0_5/i0_4 ), .ZN(
        \SB1_0_5/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_6/Component_Function_3/N3  ( .A1(\SB1_0_6/i1[9] ), .A2(
        \SB1_0_6/i1_7 ), .A3(\SB1_0_6/i0[10] ), .ZN(
        \SB1_0_6/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_6/Component_Function_4/N4  ( .A1(\SB1_0_6/i1[9] ), .A2(
        \SB1_0_6/i1_5 ), .A3(\SB1_0_6/i0_4 ), .ZN(
        \SB1_0_6/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_6/Component_Function_4/N1  ( .A1(\SB1_0_6/i0[9] ), .A2(
        \SB1_0_6/i0_0 ), .A3(\SB1_0_6/i0[8] ), .ZN(
        \SB1_0_6/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_7/Component_Function_2/N2  ( .A1(\SB1_0_7/i0_3 ), .A2(
        \SB1_0_7/i0[10] ), .A3(\SB1_0_7/i0[6] ), .ZN(
        \SB1_0_7/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_7/Component_Function_4/N2  ( .A1(\SB1_0_7/i3[0] ), .A2(
        \SB1_0_7/i0_0 ), .A3(\SB1_0_7/i1_7 ), .ZN(
        \SB1_0_7/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_7/Component_Function_4/N1  ( .A1(\SB1_0_7/i0[9] ), .A2(
        \SB1_0_7/i0_0 ), .A3(\SB1_0_7/i0[8] ), .ZN(
        \SB1_0_7/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_8/Component_Function_4/N2  ( .A1(\SB1_0_8/i3[0] ), .A2(
        \SB1_0_8/i0_0 ), .A3(\SB1_0_8/i1_7 ), .ZN(
        \SB1_0_8/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_9/Component_Function_2/N4  ( .A1(\SB1_0_9/i1_5 ), .A2(
        \SB1_0_9/i0_0 ), .A3(\SB1_0_9/i0_4 ), .ZN(
        \SB1_0_9/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_9/Component_Function_2/N1  ( .A1(\SB1_0_9/i1_5 ), .A2(
        \SB1_0_9/i0[10] ), .A3(\SB1_0_9/i1[9] ), .ZN(
        \SB1_0_9/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_9/Component_Function_4/N2  ( .A1(\SB1_0_9/i3[0] ), .A2(
        \SB1_0_9/i0_0 ), .A3(\SB1_0_9/i1_7 ), .ZN(
        \SB1_0_9/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_9/Component_Function_4/N1  ( .A1(\SB1_0_9/i0[9] ), .A2(
        \SB1_0_9/i0_0 ), .A3(\SB1_0_9/i0[8] ), .ZN(
        \SB1_0_9/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_10/Component_Function_2/N3  ( .A1(\SB1_0_10/i0_3 ), .A2(
        \SB1_0_10/i0[8] ), .A3(\SB1_0_10/i0[9] ), .ZN(
        \SB1_0_10/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_10/Component_Function_3/N1  ( .A1(\SB1_0_10/i1[9] ), .A2(
        \SB1_0_10/i0_3 ), .A3(\SB1_0_10/i0[6] ), .ZN(
        \SB1_0_10/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_10/Component_Function_4/N4  ( .A1(\SB1_0_10/i1[9] ), .A2(
        \SB1_0_10/i1_5 ), .A3(\SB1_0_10/i0_4 ), .ZN(
        \SB1_0_10/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_10/Component_Function_4/N3  ( .A1(\SB1_0_10/i0[9] ), .A2(
        \SB1_0_10/i0[10] ), .A3(\SB1_0_10/i0_3 ), .ZN(
        \SB1_0_10/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_11/Component_Function_2/N3  ( .A1(\SB1_0_11/i0_3 ), .A2(
        \SB1_0_11/i0[8] ), .A3(\SB1_0_11/i0[9] ), .ZN(
        \SB1_0_11/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_11/Component_Function_3/N4  ( .A1(\SB1_0_11/i1_5 ), .A2(
        \SB1_0_11/i0[8] ), .A3(\SB1_0_11/i3[0] ), .ZN(
        \SB1_0_11/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_11/Component_Function_4/N1  ( .A1(\SB1_0_11/i0[9] ), .A2(
        \SB1_0_11/i0_0 ), .A3(\SB1_0_11/i0[8] ), .ZN(
        \SB1_0_11/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_12/Component_Function_3/N4  ( .A1(\SB1_0_12/i1_5 ), .A2(
        \SB1_0_12/i0[8] ), .A3(\SB1_0_12/i3[0] ), .ZN(
        \SB1_0_12/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_12/Component_Function_4/N4  ( .A1(\SB1_0_12/i1[9] ), .A2(
        \SB1_0_12/i1_5 ), .A3(\SB1_0_12/i0_4 ), .ZN(
        \SB1_0_12/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_13/Component_Function_2/N1  ( .A1(\SB1_0_13/i1_5 ), .A2(
        \SB1_0_13/i0[10] ), .A3(\SB1_0_13/i1[9] ), .ZN(
        \SB1_0_13/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_13/Component_Function_4/N4  ( .A1(\SB1_0_13/i1[9] ), .A2(
        \SB1_0_13/i1_5 ), .A3(\SB1_0_13/i0_4 ), .ZN(
        \SB1_0_13/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_13/Component_Function_4/N2  ( .A1(\SB1_0_13/i3[0] ), .A2(
        \SB1_0_13/i0_0 ), .A3(\SB1_0_13/i1_7 ), .ZN(
        \SB1_0_13/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_13/Component_Function_4/N1  ( .A1(\SB1_0_13/i0[9] ), .A2(
        \SB1_0_13/i0_0 ), .A3(\SB1_0_13/i0[8] ), .ZN(
        \SB1_0_13/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_14/Component_Function_2/N2  ( .A1(\SB1_0_14/i0_3 ), .A2(
        \SB1_0_14/i0[10] ), .A3(\SB1_0_14/i0[6] ), .ZN(
        \SB1_0_14/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_14/Component_Function_2/N1  ( .A1(\SB1_0_14/i1_5 ), .A2(
        \SB1_0_14/i0[10] ), .A3(\SB1_0_14/i1[9] ), .ZN(
        \SB1_0_14/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_14/Component_Function_3/N3  ( .A1(\SB1_0_14/i1[9] ), .A2(
        \SB1_0_14/i1_7 ), .A3(\SB1_0_14/i0[10] ), .ZN(
        \SB1_0_14/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_14/Component_Function_3/N2  ( .A1(\SB1_0_14/i0_0 ), .A2(
        \SB1_0_14/i0_3 ), .A3(\SB1_0_14/i0_4 ), .ZN(
        \SB1_0_14/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_14/Component_Function_4/N4  ( .A1(\SB1_0_14/i1[9] ), .A2(
        \SB1_0_14/i1_5 ), .A3(\SB1_0_14/i0_4 ), .ZN(
        \SB1_0_14/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_14/Component_Function_4/N2  ( .A1(\SB1_0_14/i3[0] ), .A2(
        \SB1_0_14/i0_0 ), .A3(\SB1_0_14/i1_7 ), .ZN(
        \SB1_0_14/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_15/Component_Function_2/N4  ( .A1(\SB1_0_15/i1_5 ), .A2(
        \SB1_0_15/i0_0 ), .A3(\SB1_0_15/i0_4 ), .ZN(
        \SB1_0_15/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_15/Component_Function_2/N2  ( .A1(\SB1_0_15/i0_3 ), .A2(
        \SB1_0_15/i0[10] ), .A3(\SB1_0_15/i0[6] ), .ZN(
        \SB1_0_15/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_15/Component_Function_3/N4  ( .A1(\SB1_0_15/i1_5 ), .A2(
        \SB1_0_15/i0[8] ), .A3(\SB1_0_15/i3[0] ), .ZN(
        \SB1_0_15/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_15/Component_Function_4/N4  ( .A1(\SB1_0_15/i1[9] ), .A2(
        \SB1_0_15/i1_5 ), .A3(\SB1_0_15/i0_4 ), .ZN(
        \SB1_0_15/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_15/Component_Function_4/N2  ( .A1(\SB1_0_15/i3[0] ), .A2(
        \SB1_0_15/i0_0 ), .A3(\SB1_0_15/i1_7 ), .ZN(
        \SB1_0_15/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_15/Component_Function_4/N1  ( .A1(\SB1_0_15/i0[9] ), .A2(
        \SB1_0_15/i0_0 ), .A3(\SB1_0_15/i0[8] ), .ZN(
        \SB1_0_15/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_16/Component_Function_2/N2  ( .A1(\SB1_0_16/i0_3 ), .A2(
        \SB1_0_16/i0[10] ), .A3(\SB1_0_16/i0[6] ), .ZN(
        \SB1_0_16/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_16/Component_Function_4/N4  ( .A1(\SB1_0_16/i1[9] ), .A2(
        \SB1_0_16/i1_5 ), .A3(n4752), .ZN(
        \SB1_0_16/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_17/Component_Function_3/N4  ( .A1(\SB1_0_17/i1_5 ), .A2(
        \SB1_0_17/i0[8] ), .A3(\SB1_0_17/i3[0] ), .ZN(
        \SB1_0_17/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_17/Component_Function_4/N4  ( .A1(\SB1_0_17/i1[9] ), .A2(
        \SB1_0_17/i1_5 ), .A3(n2899), .ZN(
        \SB1_0_17/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_18/Component_Function_2/N3  ( .A1(\SB1_0_18/i0_3 ), .A2(
        \SB1_0_18/i0[8] ), .A3(\SB1_0_18/i0[9] ), .ZN(
        \SB1_0_18/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_18/Component_Function_3/N4  ( .A1(\SB1_0_18/i1_5 ), .A2(
        \SB1_0_18/i0[8] ), .A3(\SB1_0_18/i3[0] ), .ZN(
        \SB1_0_18/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_19/Component_Function_2/N3  ( .A1(\SB1_0_19/i0_3 ), .A2(
        \SB1_0_19/i0[8] ), .A3(\SB1_0_19/i0[9] ), .ZN(
        \SB1_0_19/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_19/Component_Function_2/N1  ( .A1(\SB1_0_19/i1_5 ), .A2(
        \SB1_0_19/i0[10] ), .A3(\SB1_0_19/i1[9] ), .ZN(
        \SB1_0_19/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_19/Component_Function_3/N2  ( .A1(\SB1_0_19/i0_0 ), .A2(
        \SB1_0_19/i0_3 ), .A3(\SB1_0_19/i0_4 ), .ZN(
        \SB1_0_19/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_19/Component_Function_3/N1  ( .A1(\SB1_0_19/i1[9] ), .A2(
        \SB1_0_19/i0_3 ), .A3(\SB1_0_19/i0[6] ), .ZN(
        \SB1_0_19/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_19/Component_Function_4/N1  ( .A1(\SB1_0_19/i0[9] ), .A2(
        \SB1_0_19/i0_0 ), .A3(\SB1_0_19/i0[8] ), .ZN(
        \SB1_0_19/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_20/Component_Function_2/N4  ( .A1(\SB1_0_20/i1_5 ), .A2(
        \SB1_0_20/i0_0 ), .A3(\SB1_0_20/i0_4 ), .ZN(
        \SB1_0_20/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_20/Component_Function_3/N1  ( .A1(\SB1_0_20/i1[9] ), .A2(
        \SB1_0_20/i0_3 ), .A3(\SB1_0_20/i0[6] ), .ZN(
        \SB1_0_20/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_20/Component_Function_4/N2  ( .A1(\SB1_0_20/i3[0] ), .A2(
        \SB1_0_20/i0_0 ), .A3(\SB1_0_20/i1_7 ), .ZN(
        \SB1_0_20/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_22/Component_Function_2/N3  ( .A1(\SB1_0_22/i0_3 ), .A2(
        \SB1_0_22/i0[8] ), .A3(\SB1_0_22/i0[9] ), .ZN(
        \SB1_0_22/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_22/Component_Function_3/N4  ( .A1(\SB1_0_22/i1_5 ), .A2(
        \SB1_0_22/i0[8] ), .A3(\SB1_0_22/i3[0] ), .ZN(
        \SB1_0_22/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_22/Component_Function_3/N1  ( .A1(\SB1_0_22/i1[9] ), .A2(
        \SB1_0_22/i0_3 ), .A3(\SB1_0_22/i0[6] ), .ZN(
        \SB1_0_22/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_22/Component_Function_4/N4  ( .A1(\SB1_0_22/i1[9] ), .A2(
        \SB1_0_22/i1_5 ), .A3(n360), .ZN(
        \SB1_0_22/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_23/Component_Function_2/N1  ( .A1(\SB1_0_23/i1_5 ), .A2(
        \SB1_0_23/i0[10] ), .A3(\SB1_0_23/i1[9] ), .ZN(
        \SB1_0_23/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_23/Component_Function_4/N2  ( .A1(\SB1_0_23/i3[0] ), .A2(
        \SB1_0_23/i0_0 ), .A3(\SB1_0_23/i1_7 ), .ZN(
        \SB1_0_23/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_23/Component_Function_4/N1  ( .A1(\SB1_0_23/i0[9] ), .A2(
        \SB1_0_23/i0_0 ), .A3(\SB1_0_23/i0[8] ), .ZN(
        \SB1_0_23/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_24/Component_Function_2/N2  ( .A1(\SB1_0_24/i0_3 ), .A2(
        \SB1_0_24/i0[10] ), .A3(\SB1_0_24/i0[6] ), .ZN(
        \SB1_0_24/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_24/Component_Function_2/N1  ( .A1(\SB1_0_24/i1_5 ), .A2(
        \SB1_0_24/i0[10] ), .A3(\SB1_0_24/i1[9] ), .ZN(
        \SB1_0_24/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_24/Component_Function_3/N4  ( .A1(\SB1_0_24/i1_5 ), .A2(
        \SB1_0_24/i0[8] ), .A3(\SB1_0_24/i3[0] ), .ZN(
        \SB1_0_24/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_24/Component_Function_3/N3  ( .A1(\SB1_0_24/i1[9] ), .A2(
        \SB1_0_24/i1_7 ), .A3(\SB1_0_24/i0[10] ), .ZN(
        \SB1_0_24/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_24/Component_Function_3/N2  ( .A1(\SB1_0_24/i0_0 ), .A2(
        \SB1_0_24/i0_3 ), .A3(\SB1_0_24/i0_4 ), .ZN(
        \SB1_0_24/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_24/Component_Function_3/N1  ( .A1(\SB1_0_24/i1[9] ), .A2(
        \SB1_0_24/i0_3 ), .A3(\SB1_0_24/i0[6] ), .ZN(
        \SB1_0_24/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_24/Component_Function_4/N4  ( .A1(\SB1_0_24/i1[9] ), .A2(
        \SB1_0_24/i1_5 ), .A3(\SB1_0_24/i0_4 ), .ZN(
        \SB1_0_24/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_24/Component_Function_4/N3  ( .A1(\SB1_0_24/i0[9] ), .A2(
        \SB1_0_24/i0[10] ), .A3(\SB1_0_24/i0_3 ), .ZN(
        \SB1_0_24/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_24/Component_Function_4/N1  ( .A1(\SB1_0_24/i0[9] ), .A2(
        \SB1_0_24/i0_0 ), .A3(\SB1_0_24/i0[8] ), .ZN(
        \SB1_0_24/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_25/Component_Function_2/N2  ( .A1(\SB1_0_25/i0_3 ), .A2(
        \SB1_0_25/i0[10] ), .A3(\SB1_0_25/i0[6] ), .ZN(
        \SB1_0_25/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_25/Component_Function_4/N2  ( .A1(\SB1_0_25/i3[0] ), .A2(
        \SB1_0_25/i0_0 ), .A3(\SB1_0_25/i1_7 ), .ZN(
        \SB1_0_25/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_26/Component_Function_2/N3  ( .A1(\SB1_0_26/i0_3 ), .A2(
        \SB1_0_26/i0[8] ), .A3(\SB1_0_26/i0[9] ), .ZN(
        \SB1_0_26/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_26/Component_Function_3/N4  ( .A1(\SB1_0_26/i1_5 ), .A2(
        \SB1_0_26/i0[8] ), .A3(\SB1_0_26/i3[0] ), .ZN(
        \SB1_0_26/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_26/Component_Function_3/N1  ( .A1(\SB1_0_26/i1[9] ), .A2(
        \SB1_0_26/i0_3 ), .A3(\SB1_0_26/i0[6] ), .ZN(
        \SB1_0_26/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_26/Component_Function_4/N2  ( .A1(\SB1_0_26/i3[0] ), .A2(
        \SB1_0_26/i0_0 ), .A3(\SB1_0_26/i1_7 ), .ZN(
        \SB1_0_26/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_26/Component_Function_4/N1  ( .A1(\SB1_0_26/i0[9] ), .A2(
        \SB1_0_26/i0_0 ), .A3(\SB1_0_26/i0[8] ), .ZN(
        \SB1_0_26/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_27/Component_Function_2/N4  ( .A1(\SB1_0_27/i1_5 ), .A2(
        \SB1_0_27/i0_0 ), .A3(\SB1_0_27/i0_4 ), .ZN(
        \SB1_0_27/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_27/Component_Function_2/N3  ( .A1(\SB1_0_27/i0_3 ), .A2(
        \SB1_0_27/i0[8] ), .A3(\SB1_0_27/i0[9] ), .ZN(
        \SB1_0_27/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_27/Component_Function_2/N2  ( .A1(\SB1_0_27/i0_3 ), .A2(
        \SB1_0_27/i0[10] ), .A3(\SB1_0_27/i0[6] ), .ZN(
        \SB1_0_27/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_27/Component_Function_2/N1  ( .A1(\SB1_0_27/i1_5 ), .A2(
        \SB1_0_27/i0[10] ), .A3(\SB1_0_27/i1[9] ), .ZN(
        \SB1_0_27/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_27/Component_Function_4/N3  ( .A1(\SB1_0_27/i0[9] ), .A2(
        \SB1_0_27/i0[10] ), .A3(\SB1_0_27/i0_3 ), .ZN(
        \SB1_0_27/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_27/Component_Function_4/N2  ( .A1(\SB1_0_27/i3[0] ), .A2(
        \SB1_0_27/i0_0 ), .A3(\SB1_0_27/i1_7 ), .ZN(
        \SB1_0_27/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_27/Component_Function_4/N1  ( .A1(\SB1_0_27/i0[9] ), .A2(
        \SB1_0_27/i0_0 ), .A3(\SB1_0_27/i0[8] ), .ZN(
        \SB1_0_27/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_28/Component_Function_2/N1  ( .A1(\SB1_0_28/i1_5 ), .A2(
        \SB1_0_28/i0[10] ), .A3(\SB1_0_28/i1[9] ), .ZN(
        \SB1_0_28/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_28/Component_Function_3/N4  ( .A1(\SB1_0_28/i1_5 ), .A2(
        \SB1_0_28/i0[8] ), .A3(\SB1_0_28/i3[0] ), .ZN(
        \SB1_0_28/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_29/Component_Function_4/N4  ( .A1(\SB1_0_29/i1[9] ), .A2(
        \SB1_0_29/i1_5 ), .A3(n346), .ZN(
        \SB1_0_29/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_30/Component_Function_2/N3  ( .A1(\SB1_0_30/i0_3 ), .A2(
        \SB1_0_30/i0[8] ), .A3(\SB1_0_30/i0[9] ), .ZN(
        \SB1_0_30/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_30/Component_Function_2/N2  ( .A1(\SB1_0_30/i0_3 ), .A2(
        \SB1_0_30/i0[10] ), .A3(\SB1_0_30/i0[6] ), .ZN(
        \SB1_0_30/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_30/Component_Function_2/N1  ( .A1(\SB1_0_30/i1_5 ), .A2(
        \SB1_0_30/i0[10] ), .A3(\SB1_0_30/i1[9] ), .ZN(
        \SB1_0_30/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_30/Component_Function_3/N2  ( .A1(\SB1_0_30/i0_0 ), .A2(
        \SB1_0_30/i0_3 ), .A3(\SB1_0_30/i0_4 ), .ZN(
        \SB1_0_30/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_30/Component_Function_3/N1  ( .A1(\SB1_0_30/i1[9] ), .A2(
        \SB1_0_30/i0_3 ), .A3(\SB1_0_30/i0[6] ), .ZN(
        \SB1_0_30/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_30/Component_Function_4/N4  ( .A1(\SB1_0_30/i1[9] ), .A2(
        \SB1_0_30/i1_5 ), .A3(\SB1_0_30/i0_4 ), .ZN(
        \SB1_0_30/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_30/Component_Function_4/N3  ( .A1(\SB1_0_30/i0[9] ), .A2(
        \SB1_0_30/i0[10] ), .A3(\SB1_0_30/i0_3 ), .ZN(
        \SB1_0_30/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_30/Component_Function_4/N2  ( .A1(\SB1_0_30/i3[0] ), .A2(
        \SB1_0_30/i0_0 ), .A3(\SB1_0_30/i1_7 ), .ZN(
        \SB1_0_30/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_30/Component_Function_4/N1  ( .A1(\SB1_0_30/i0[9] ), .A2(
        \SB1_0_30/i0_0 ), .A3(\SB1_0_30/i0[8] ), .ZN(
        \SB1_0_30/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_31/Component_Function_2/N4  ( .A1(\SB1_0_31/i1_5 ), .A2(
        \SB1_0_31/i0_0 ), .A3(\SB1_0_31/i0_4 ), .ZN(
        \SB1_0_31/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_31/Component_Function_2/N1  ( .A1(\SB1_0_31/i1_5 ), .A2(
        \SB1_0_31/i0[10] ), .A3(\SB1_0_31/i1[9] ), .ZN(
        \SB1_0_31/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_31/Component_Function_4/N2  ( .A1(\SB1_0_31/i3[0] ), .A2(
        \SB1_0_31/i0_0 ), .A3(\SB1_0_31/i1_7 ), .ZN(
        \SB1_0_31/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_31/Component_Function_4/N1  ( .A1(\SB1_0_31/i0[9] ), .A2(
        \SB1_0_31/i0_0 ), .A3(\SB1_0_31/i0[8] ), .ZN(
        \SB1_0_31/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_0/Component_Function_4/N4  ( .A1(\SB2_0_0/i1[9] ), .A2(
        \SB2_0_0/i1_5 ), .A3(\RI3[0][190] ), .ZN(
        \SB2_0_0/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_0/Component_Function_4/N1  ( .A1(\SB2_0_0/i0[9] ), .A2(
        \SB2_0_0/i0_0 ), .A3(\SB2_0_0/i0[8] ), .ZN(
        \SB2_0_0/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_1/Component_Function_4/N4  ( .A1(\SB2_0_1/i1[9] ), .A2(
        \SB2_0_1/i1_5 ), .A3(\SB2_0_1/i0_4 ), .ZN(
        \SB2_0_1/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_2/Component_Function_4/N4  ( .A1(\SB2_0_2/i1[9] ), .A2(
        \SB2_0_2/i1_5 ), .A3(\RI3[0][178] ), .ZN(
        \SB2_0_2/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_2/Component_Function_4/N2  ( .A1(\SB2_0_2/i3[0] ), .A2(
        \RI3[0][176] ), .A3(\SB2_0_2/i1_7 ), .ZN(
        \SB2_0_2/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_3/Component_Function_4/N1  ( .A1(\SB2_0_3/i0[9] ), .A2(
        \SB2_0_3/i0_0 ), .A3(\SB2_0_3/i0[8] ), .ZN(
        \SB2_0_3/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_4/Component_Function_4/N2  ( .A1(\SB2_0_4/i3[0] ), .A2(
        \SB2_0_4/i0_0 ), .A3(\SB2_0_4/i1_7 ), .ZN(
        \SB2_0_4/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_4/Component_Function_4/N1  ( .A1(\SB2_0_4/i0[9] ), .A2(
        \SB2_0_4/i0_0 ), .A3(\SB2_0_4/i0[8] ), .ZN(
        \SB2_0_4/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_5/Component_Function_2/N4  ( .A1(\SB2_0_5/i1_5 ), .A2(
        \SB2_0_5/i0_0 ), .A3(\RI3[0][160] ), .ZN(
        \SB2_0_5/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_5/Component_Function_3/N4  ( .A1(\SB2_0_5/i1_5 ), .A2(
        \SB2_0_5/i0[8] ), .A3(\SB2_0_5/i3[0] ), .ZN(
        \SB2_0_5/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_5/Component_Function_4/N2  ( .A1(\SB2_0_5/i3[0] ), .A2(
        \SB2_0_5/i0_0 ), .A3(\SB2_0_5/i1_7 ), .ZN(
        \SB2_0_5/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_5/Component_Function_4/N1  ( .A1(\RI3[0][156] ), .A2(
        \SB2_0_5/i0_0 ), .A3(\SB2_0_5/i0[8] ), .ZN(
        \SB2_0_5/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_6/Component_Function_4/N4  ( .A1(\SB2_0_6/i1[9] ), .A2(
        \SB2_0_6/i1_5 ), .A3(\RI3[0][154] ), .ZN(
        \SB2_0_6/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_6/Component_Function_4/N2  ( .A1(\SB2_0_6/i3[0] ), .A2(
        \SB2_0_6/i0_0 ), .A3(\SB2_0_6/i1_7 ), .ZN(
        \SB2_0_6/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_6/Component_Function_4/N1  ( .A1(\SB2_0_6/i0[9] ), .A2(
        \SB2_0_6/i0_0 ), .A3(\SB2_0_6/i0[8] ), .ZN(
        \SB2_0_6/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_7/Component_Function_4/N4  ( .A1(\SB2_0_7/i1[9] ), .A2(
        \SB2_0_7/i1_5 ), .A3(\SB1_0_8/buf_output[4] ), .ZN(
        \SB2_0_7/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_7/Component_Function_4/N2  ( .A1(\SB2_0_7/i3[0] ), .A2(
        \SB2_0_7/i0_0 ), .A3(\SB2_0_7/i1_7 ), .ZN(
        \SB2_0_7/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_8/Component_Function_4/N2  ( .A1(\SB2_0_8/i3[0] ), .A2(
        \SB2_0_8/i0_0 ), .A3(\SB2_0_8/i1_7 ), .ZN(
        \SB2_0_8/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_8/Component_Function_4/N1  ( .A1(\SB2_0_8/i0[9] ), .A2(
        \SB2_0_8/i0_0 ), .A3(\SB2_0_8/i0[8] ), .ZN(
        \SB2_0_8/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_9/Component_Function_3/N4  ( .A1(n5518), .A2(\SB2_0_9/i0[8] ), .A3(\SB2_0_9/i3[0] ), .ZN(\SB2_0_9/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_9/Component_Function_4/N2  ( .A1(\SB2_0_9/i3[0] ), .A2(
        \RI3[0][134] ), .A3(\SB2_0_9/i1_7 ), .ZN(
        \SB2_0_9/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_9/Component_Function_4/N1  ( .A1(\SB2_0_9/i0[9] ), .A2(
        \RI3[0][134] ), .A3(\SB2_0_9/i0[8] ), .ZN(
        \SB2_0_9/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_10/Component_Function_2/N1  ( .A1(\SB2_0_10/i1_5 ), .A2(
        \SB2_0_10/i0[10] ), .A3(\SB2_0_10/i1[9] ), .ZN(
        \SB2_0_10/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_10/Component_Function_3/N1  ( .A1(\SB2_0_10/i1[9] ), .A2(
        \SB2_0_10/i0_3 ), .A3(\SB2_0_10/i0[6] ), .ZN(
        \SB2_0_10/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_10/Component_Function_4/N2  ( .A1(\SB2_0_10/i3[0] ), .A2(
        \SB2_0_10/i0_0 ), .A3(\SB2_0_10/i1_7 ), .ZN(
        \SB2_0_10/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_11/Component_Function_3/N3  ( .A1(\SB2_0_11/i1[9] ), .A2(
        \SB2_0_11/i1_7 ), .A3(\SB2_0_11/i0[10] ), .ZN(
        \SB2_0_11/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_11/Component_Function_3/N1  ( .A1(\SB2_0_11/i1[9] ), .A2(
        \SB2_0_11/i0_3 ), .A3(\SB2_0_11/i0[6] ), .ZN(
        \SB2_0_11/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_11/Component_Function_4/N1  ( .A1(n1911), .A2(
        \SB2_0_11/i0_0 ), .A3(\SB2_0_11/i0[8] ), .ZN(
        \SB2_0_11/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_12/Component_Function_2/N1  ( .A1(\SB2_0_12/i1_5 ), .A2(
        \SB2_0_12/i0[10] ), .A3(\SB2_0_12/i1[9] ), .ZN(
        \SB2_0_12/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_12/Component_Function_4/N2  ( .A1(\SB2_0_12/i3[0] ), .A2(
        \SB2_0_12/i0_0 ), .A3(\SB2_0_12/i1_7 ), .ZN(
        \SB2_0_12/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_13/Component_Function_4/N1  ( .A1(\SB2_0_13/i0[9] ), .A2(
        \SB2_0_13/i0_0 ), .A3(n1393), .ZN(
        \SB2_0_13/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_14/Component_Function_2/N4  ( .A1(\SB2_0_14/i1_5 ), .A2(
        \RI3[0][104] ), .A3(\RI3[0][106] ), .ZN(
        \SB2_0_14/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_14/Component_Function_4/N2  ( .A1(\SB2_0_14/i3[0] ), .A2(
        \RI3[0][104] ), .A3(\SB2_0_14/i1_7 ), .ZN(
        \SB2_0_14/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_15/Component_Function_4/N2  ( .A1(\SB2_0_15/i3[0] ), .A2(
        \SB2_0_15/i0_0 ), .A3(\SB2_0_15/i1_7 ), .ZN(
        \SB2_0_15/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_15/Component_Function_4/N1  ( .A1(\SB2_0_15/i0[9] ), .A2(
        \SB2_0_15/i0_0 ), .A3(\SB2_0_15/i0[8] ), .ZN(
        \SB2_0_15/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_16/Component_Function_3/N4  ( .A1(\SB2_0_16/i1_5 ), .A2(
        \SB2_0_16/i0[8] ), .A3(\SB2_0_16/i3[0] ), .ZN(
        \SB2_0_16/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_16/Component_Function_4/N2  ( .A1(\SB2_0_16/i3[0] ), .A2(
        \SB2_0_16/i0_0 ), .A3(\SB2_0_16/i1_7 ), .ZN(
        \SB2_0_16/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_16/Component_Function_4/N1  ( .A1(\SB2_0_16/i0[9] ), .A2(
        \SB2_0_16/i0_0 ), .A3(\SB2_0_16/i0[8] ), .ZN(
        \SB2_0_16/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_17/Component_Function_4/N2  ( .A1(\SB2_0_17/i3[0] ), .A2(
        \SB2_0_17/i0_0 ), .A3(\SB2_0_17/i1_7 ), .ZN(
        \SB2_0_17/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_18/Component_Function_4/N2  ( .A1(\SB2_0_18/i3[0] ), .A2(
        \SB2_0_18/i0_0 ), .A3(\SB2_0_18/i1_7 ), .ZN(
        \SB2_0_18/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_19/Component_Function_4/N4  ( .A1(\SB2_0_19/i1[9] ), .A2(
        \SB2_0_19/i1_5 ), .A3(\RI3[0][76] ), .ZN(
        \SB2_0_19/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_19/Component_Function_4/N2  ( .A1(\SB2_0_19/i3[0] ), .A2(
        \SB2_0_19/i0_0 ), .A3(\SB2_0_19/i1_7 ), .ZN(
        \SB2_0_19/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_19/Component_Function_4/N1  ( .A1(\SB2_0_19/i0[9] ), .A2(
        \SB2_0_19/i0_0 ), .A3(\SB2_0_19/i0[8] ), .ZN(
        \SB2_0_19/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_20/Component_Function_3/N1  ( .A1(\SB2_0_20/i1[9] ), .A2(
        \SB2_0_20/i0_3 ), .A3(\SB2_0_20/i0[6] ), .ZN(
        \SB2_0_20/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_20/Component_Function_4/N2  ( .A1(\SB2_0_20/i3[0] ), .A2(
        \SB2_0_20/i0_0 ), .A3(\SB2_0_20/i1_7 ), .ZN(
        \SB2_0_20/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_21/Component_Function_4/N4  ( .A1(\SB2_0_21/i1[9] ), .A2(
        \SB2_0_21/i1_5 ), .A3(\SB1_0_22/buf_output[4] ), .ZN(
        \SB2_0_21/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_21/Component_Function_4/N2  ( .A1(\SB2_0_21/i3[0] ), .A2(
        \SB2_0_21/i0_0 ), .A3(\SB2_0_21/i1_7 ), .ZN(
        \SB2_0_21/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_21/Component_Function_4/N1  ( .A1(\SB2_0_21/i0[9] ), .A2(
        \SB2_0_21/i0_0 ), .A3(\SB2_0_21/i0[8] ), .ZN(
        \SB2_0_21/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_22/Component_Function_4/N1  ( .A1(\RI3[0][54] ), .A2(
        \SB2_0_22/i0_0 ), .A3(\SB2_0_22/i0[8] ), .ZN(
        \SB2_0_22/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_23/Component_Function_4/N2  ( .A1(\SB2_0_23/i3[0] ), .A2(
        \SB2_0_23/i0_0 ), .A3(\SB2_0_23/i1_7 ), .ZN(
        \SB2_0_23/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_23/Component_Function_4/N1  ( .A1(\SB2_0_23/i0[9] ), .A2(
        \SB2_0_23/i0_0 ), .A3(\SB2_0_23/i0[8] ), .ZN(
        \SB2_0_23/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_26/Component_Function_4/N1  ( .A1(\SB2_0_26/i0[9] ), .A2(
        \SB2_0_26/i0_0 ), .A3(\SB2_0_26/i0[8] ), .ZN(
        \SB2_0_26/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_27/Component_Function_4/N2  ( .A1(\SB2_0_27/i3[0] ), .A2(
        \SB2_0_27/i0_0 ), .A3(\SB2_0_27/i1_7 ), .ZN(
        \SB2_0_27/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_28/Component_Function_4/N1  ( .A1(\RI3[0][18] ), .A2(
        \SB2_0_28/i0_0 ), .A3(\SB2_0_28/i0[8] ), .ZN(
        \SB2_0_28/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_29/Component_Function_3/N3  ( .A1(\SB2_0_29/i1[9] ), .A2(
        \SB2_0_29/i1_7 ), .A3(\RI3[0][15] ), .ZN(
        \SB2_0_29/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_29/Component_Function_3/N1  ( .A1(\SB2_0_29/i1[9] ), .A2(
        \SB2_0_29/i0_3 ), .A3(\SB2_0_29/i0[6] ), .ZN(
        \SB2_0_29/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_29/Component_Function_4/N2  ( .A1(\SB2_0_29/i3[0] ), .A2(
        \SB2_0_29/i0_0 ), .A3(\SB2_0_29/i1_7 ), .ZN(
        \SB2_0_29/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_29/Component_Function_4/N1  ( .A1(n2605), .A2(
        \SB2_0_29/i0_0 ), .A3(\SB2_0_29/i0[8] ), .ZN(
        \SB2_0_29/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_30/Component_Function_2/N2  ( .A1(\SB2_0_30/i0_3 ), .A2(
        \SB2_0_30/i0[10] ), .A3(\SB2_0_30/i0[6] ), .ZN(
        \SB2_0_30/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_30/Component_Function_4/N4  ( .A1(\SB2_0_30/i1[9] ), .A2(
        \SB2_0_30/i1_5 ), .A3(\RI3[0][10] ), .ZN(
        \SB2_0_30/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_30/Component_Function_4/N3  ( .A1(\SB2_0_30/i0[9] ), .A2(
        \SB2_0_30/i0[10] ), .A3(\SB2_0_30/i0_3 ), .ZN(
        \SB2_0_30/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_31/Component_Function_2/N1  ( .A1(\SB2_0_31/i1_5 ), .A2(
        \SB2_0_31/i0[10] ), .A3(\SB2_0_31/i1[9] ), .ZN(
        \SB2_0_31/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_31/Component_Function_3/N4  ( .A1(\SB2_0_31/i1_5 ), .A2(
        \SB2_0_31/i0[8] ), .A3(\SB2_0_31/i3[0] ), .ZN(
        \SB2_0_31/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_31/Component_Function_3/N3  ( .A1(\SB2_0_31/i1[9] ), .A2(
        \SB2_0_31/i1_7 ), .A3(\SB2_0_31/i0[10] ), .ZN(
        \SB2_0_31/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_31/Component_Function_3/N1  ( .A1(\SB2_0_31/i1[9] ), .A2(
        \SB2_0_31/i0_3 ), .A3(\SB2_0_31/i0[6] ), .ZN(
        \SB2_0_31/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_31/Component_Function_4/N2  ( .A1(\SB2_0_31/i3[0] ), .A2(
        \SB2_0_31/i0_0 ), .A3(\SB2_0_31/i1_7 ), .ZN(
        \SB2_0_31/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_31/Component_Function_4/N1  ( .A1(\SB2_0_31/i0[9] ), .A2(
        \SB2_0_31/i0_0 ), .A3(\SB2_0_31/i0[8] ), .ZN(
        \SB2_0_31/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_3/Component_Function_4/N1  ( .A1(\SB1_1_3/i0[9] ), .A2(
        \SB1_1_3/i0_0 ), .A3(\SB1_1_3/i0[8] ), .ZN(
        \SB1_1_3/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_4/Component_Function_2/N4  ( .A1(\SB1_1_4/i1_5 ), .A2(
        \SB1_1_4/i0_0 ), .A3(\SB1_1_4/i0_4 ), .ZN(
        \SB1_1_4/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_4/Component_Function_3/N4  ( .A1(\SB1_1_4/i1_5 ), .A2(
        \SB1_1_4/i0[8] ), .A3(\SB1_1_4/i3[0] ), .ZN(
        \SB1_1_4/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_6/Component_Function_4/N3  ( .A1(\SB1_1_6/i0[9] ), .A2(
        \SB1_1_6/i0[10] ), .A3(\SB1_1_6/i0_3 ), .ZN(
        \SB1_1_6/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_8/Component_Function_2/N4  ( .A1(n3647), .A2(\SB1_1_8/i0_0 ), 
        .A3(\SB1_1_8/i0_4 ), .ZN(\SB1_1_8/Component_Function_2/NAND4_in[3] )
         );
  NAND3_X1 \SB1_1_8/Component_Function_3/N3  ( .A1(\SB1_1_8/i1[9] ), .A2(
        \SB1_1_8/i1_7 ), .A3(\SB1_1_8/i0[10] ), .ZN(
        \SB1_1_8/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_9/Component_Function_4/N2  ( .A1(\SB1_1_9/i3[0] ), .A2(
        \SB1_1_9/i0_0 ), .A3(\SB1_1_9/i1_7 ), .ZN(
        \SB1_1_9/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_9/Component_Function_4/N1  ( .A1(\SB1_1_9/i0[9] ), .A2(
        \SB1_1_9/i0_0 ), .A3(\SB1_1_9/i0[8] ), .ZN(
        \SB1_1_9/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_10/Component_Function_2/N1  ( .A1(\SB1_1_10/i1_5 ), .A2(
        \SB1_1_10/i0[10] ), .A3(\SB1_1_10/i1[9] ), .ZN(
        \SB1_1_10/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_10/Component_Function_3/N1  ( .A1(\SB1_1_10/i1[9] ), .A2(
        \SB1_1_10/i0_3 ), .A3(\SB1_1_10/i0[6] ), .ZN(
        \SB1_1_10/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_10/Component_Function_4/N1  ( .A1(\SB1_1_10/i0[9] ), .A2(
        \SB1_1_10/i0_0 ), .A3(\SB1_1_10/i0[8] ), .ZN(
        \SB1_1_10/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_11/Component_Function_2/N3  ( .A1(\SB1_1_11/i0_3 ), .A2(
        \SB1_1_11/i0[8] ), .A3(\SB1_1_11/i0[9] ), .ZN(
        \SB1_1_11/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_11/Component_Function_2/N1  ( .A1(\SB1_1_11/i1_5 ), .A2(
        \SB1_1_11/i0[10] ), .A3(\SB1_1_11/i1[9] ), .ZN(
        \SB1_1_11/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_11/Component_Function_3/N2  ( .A1(\SB1_1_11/i0_0 ), .A2(
        \SB1_1_11/i0_3 ), .A3(\SB1_1_11/i0_4 ), .ZN(
        \SB1_1_11/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_11/Component_Function_4/N1  ( .A1(\SB1_1_11/i0[9] ), .A2(
        \SB1_1_11/i0_0 ), .A3(\SB1_1_11/i0[8] ), .ZN(
        \SB1_1_11/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_12/Component_Function_2/N2  ( .A1(\SB1_1_12/i0_3 ), .A2(
        \SB1_1_12/i0[10] ), .A3(\SB1_1_12/i0[6] ), .ZN(
        \SB1_1_12/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_12/Component_Function_3/N2  ( .A1(\SB1_1_12/i0_0 ), .A2(
        \SB1_1_12/i0_3 ), .A3(\SB1_1_12/i0_4 ), .ZN(
        \SB1_1_12/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_13/Component_Function_4/N1  ( .A1(\SB1_1_13/i0[9] ), .A2(
        \SB1_1_13/i0_0 ), .A3(\SB1_1_13/i0[8] ), .ZN(
        \SB1_1_13/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_14/Component_Function_4/N4  ( .A1(\SB1_1_14/i1[9] ), .A2(
        \SB1_1_14/i1_5 ), .A3(\SB1_1_14/i0_4 ), .ZN(
        \SB1_1_14/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_14/Component_Function_4/N1  ( .A1(\SB1_1_14/i0[9] ), .A2(
        \SB1_1_14/i0_0 ), .A3(\SB1_1_14/i0[8] ), .ZN(
        \SB1_1_14/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_15/Component_Function_3/N1  ( .A1(\SB1_1_15/i1[9] ), .A2(
        \SB1_1_15/i0_3 ), .A3(\SB1_1_15/i0[6] ), .ZN(
        \SB1_1_15/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_15/Component_Function_4/N2  ( .A1(\SB1_1_15/i3[0] ), .A2(
        \SB1_1_15/i0_0 ), .A3(\SB1_1_15/i1_7 ), .ZN(
        \SB1_1_15/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_15/Component_Function_4/N1  ( .A1(\SB1_1_15/i0[9] ), .A2(
        \SB1_1_15/i0_0 ), .A3(\SB1_1_15/i0[8] ), .ZN(
        \SB1_1_15/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_16/Component_Function_2/N2  ( .A1(\SB1_1_16/i0_3 ), .A2(
        \SB1_1_16/i0[10] ), .A3(\SB1_1_16/i0[6] ), .ZN(
        \SB1_1_16/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_17/Component_Function_2/N3  ( .A1(\SB1_1_17/i0_3 ), .A2(
        \SB1_1_17/i0[8] ), .A3(\SB1_1_17/i0[9] ), .ZN(
        \SB1_1_17/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_17/Component_Function_3/N1  ( .A1(\SB1_1_17/i1[9] ), .A2(
        \SB1_1_17/i0_3 ), .A3(\SB1_1_17/i0[6] ), .ZN(
        \SB1_1_17/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_18/Component_Function_2/N3  ( .A1(\SB1_1_18/i0_3 ), .A2(
        \SB1_1_18/i0[8] ), .A3(\SB1_1_18/i0[9] ), .ZN(
        \SB1_1_18/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_18/Component_Function_2/N1  ( .A1(\SB1_1_18/i1_5 ), .A2(
        \SB1_1_18/i0[10] ), .A3(\SB1_1_18/i1[9] ), .ZN(
        \SB1_1_18/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_18/Component_Function_4/N3  ( .A1(\SB1_1_18/i0[9] ), .A2(
        \SB1_1_18/i0[10] ), .A3(\SB1_1_18/i0_3 ), .ZN(
        \SB1_1_18/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_18/Component_Function_4/N2  ( .A1(\SB1_1_18/i3[0] ), .A2(
        \SB1_1_18/i0_0 ), .A3(\SB1_1_18/i1_7 ), .ZN(
        \SB1_1_18/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_18/Component_Function_4/N1  ( .A1(\SB1_1_18/i0[9] ), .A2(
        \SB1_1_18/i0_0 ), .A3(\SB1_1_18/i0[8] ), .ZN(
        \SB1_1_18/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_19/Component_Function_2/N4  ( .A1(\SB1_1_19/i1_5 ), .A2(
        \SB1_1_19/i0_0 ), .A3(\SB1_1_19/i0_4 ), .ZN(
        \SB1_1_19/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_19/Component_Function_3/N1  ( .A1(\SB1_1_19/i1[9] ), .A2(
        \SB1_1_19/i0_3 ), .A3(\SB1_1_19/i0[6] ), .ZN(
        \SB1_1_19/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_20/Component_Function_2/N1  ( .A1(\SB1_1_20/i1_5 ), .A2(
        \SB1_1_20/i0[10] ), .A3(\SB1_1_20/i1[9] ), .ZN(
        \SB1_1_20/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_21/Component_Function_2/N2  ( .A1(\SB1_1_21/i0_3 ), .A2(
        \SB1_1_21/i0[10] ), .A3(\SB1_1_21/i0[6] ), .ZN(
        \SB1_1_21/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_21/Component_Function_4/N2  ( .A1(\SB1_1_21/i3[0] ), .A2(
        \SB1_1_21/i0_0 ), .A3(\SB1_1_21/i1_7 ), .ZN(
        \SB1_1_21/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_21/Component_Function_4/N1  ( .A1(\SB1_1_21/i0[9] ), .A2(
        \SB1_1_21/i0_0 ), .A3(\SB1_1_21/i0[8] ), .ZN(
        \SB1_1_21/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_22/Component_Function_4/N2  ( .A1(\SB1_1_22/i3[0] ), .A2(
        \SB1_1_22/i0_0 ), .A3(\SB1_1_22/i1_7 ), .ZN(
        \SB1_1_22/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_24/Component_Function_4/N2  ( .A1(\SB1_1_24/i3[0] ), .A2(
        \SB1_1_24/i0_0 ), .A3(\SB1_1_24/i1_7 ), .ZN(
        \SB1_1_24/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_24/Component_Function_4/N1  ( .A1(\SB1_1_24/i0[9] ), .A2(
        \SB1_1_24/i0_0 ), .A3(\SB1_1_24/i0[8] ), .ZN(
        \SB1_1_24/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_25/Component_Function_3/N1  ( .A1(\SB1_1_25/i1[9] ), .A2(
        \SB1_1_25/i0_3 ), .A3(\SB1_1_25/i0[6] ), .ZN(
        \SB1_1_25/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_25/Component_Function_4/N3  ( .A1(\SB1_1_25/i0[9] ), .A2(
        \SB1_1_25/i0[10] ), .A3(\SB1_1_25/i0_3 ), .ZN(
        \SB1_1_25/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_25/Component_Function_4/N2  ( .A1(\SB1_1_25/i3[0] ), .A2(
        \SB1_1_25/i0_0 ), .A3(\SB1_1_25/i1_7 ), .ZN(
        \SB1_1_25/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_25/Component_Function_4/N1  ( .A1(\SB1_1_25/i0[9] ), .A2(
        \SB1_1_25/i0_0 ), .A3(\SB1_1_25/i0[8] ), .ZN(
        \SB1_1_25/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_26/Component_Function_2/N3  ( .A1(\SB1_1_26/i0_3 ), .A2(
        \SB1_1_26/i0[8] ), .A3(\SB1_1_26/i0[9] ), .ZN(
        \SB1_1_26/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_26/Component_Function_3/N1  ( .A1(\SB1_1_26/i1[9] ), .A2(
        \SB1_1_26/i0_3 ), .A3(\SB1_1_26/i0[6] ), .ZN(
        \SB1_1_26/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_26/Component_Function_4/N4  ( .A1(\SB1_1_26/i1[9] ), .A2(
        \SB1_1_26/i1_5 ), .A3(\SB1_1_26/i0_4 ), .ZN(
        \SB1_1_26/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_26/Component_Function_4/N1  ( .A1(\SB1_1_26/i0[9] ), .A2(
        \SB1_1_26/i0_0 ), .A3(\SB1_1_26/i0[8] ), .ZN(
        \SB1_1_26/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_29/Component_Function_2/N2  ( .A1(\SB1_1_29/i0_3 ), .A2(
        \SB1_1_29/i0[10] ), .A3(\SB1_1_29/i0[6] ), .ZN(
        \SB1_1_29/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_29/Component_Function_2/N1  ( .A1(\SB1_1_29/i1_5 ), .A2(
        \SB1_1_29/i0[10] ), .A3(\SB1_1_29/i1[9] ), .ZN(
        \SB1_1_29/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_29/Component_Function_3/N1  ( .A1(\SB1_1_29/i1[9] ), .A2(
        \SB1_1_29/i0_3 ), .A3(\SB1_1_29/i0[6] ), .ZN(
        \SB1_1_29/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_29/Component_Function_4/N2  ( .A1(\SB1_1_29/i3[0] ), .A2(
        \SB1_1_29/i0_0 ), .A3(\SB1_1_29/i1_7 ), .ZN(
        \SB1_1_29/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_29/Component_Function_4/N1  ( .A1(\SB1_1_29/i0[9] ), .A2(
        \SB1_1_29/i0_0 ), .A3(\SB1_1_29/i0[8] ), .ZN(
        \SB1_1_29/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_30/Component_Function_2/N3  ( .A1(\SB1_1_30/i0_3 ), .A2(
        \SB1_1_30/i0[8] ), .A3(\SB1_1_30/i0[9] ), .ZN(
        \SB1_1_30/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_30/Component_Function_4/N3  ( .A1(\SB1_1_30/i0[9] ), .A2(
        \SB1_1_30/i0[10] ), .A3(\SB1_1_30/i0_3 ), .ZN(
        \SB1_1_30/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_31/Component_Function_2/N1  ( .A1(\SB1_1_31/i1_5 ), .A2(
        \SB1_1_31/i0[10] ), .A3(\SB1_1_31/i1[9] ), .ZN(
        \SB1_1_31/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_31/Component_Function_3/N3  ( .A1(\SB1_1_31/i1[9] ), .A2(
        \SB1_1_31/i1_7 ), .A3(\SB1_1_31/i0[10] ), .ZN(
        \SB1_1_31/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_0/Component_Function_4/N1  ( .A1(\SB2_1_0/i0[9] ), .A2(
        \SB2_1_0/i0_0 ), .A3(\SB2_1_0/i0[8] ), .ZN(
        \SB2_1_0/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_1/Component_Function_4/N2  ( .A1(\SB2_1_1/i3[0] ), .A2(
        \SB2_1_1/i0_0 ), .A3(\SB2_1_1/i1_7 ), .ZN(
        \SB2_1_1/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_1/Component_Function_4/N1  ( .A1(\SB2_1_1/i0[9] ), .A2(
        \SB2_1_1/i0_0 ), .A3(\SB2_1_1/i0[8] ), .ZN(
        \SB2_1_1/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_2/Component_Function_4/N1  ( .A1(\SB2_1_2/i0[9] ), .A2(
        \SB2_1_2/i0_0 ), .A3(\SB2_1_2/i0[8] ), .ZN(
        \SB2_1_2/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_3/Component_Function_4/N1  ( .A1(\SB2_1_3/i0[9] ), .A2(
        \SB2_1_3/i0_0 ), .A3(\SB2_1_3/i0[8] ), .ZN(
        \SB2_1_3/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_4/Component_Function_2/N4  ( .A1(\SB2_1_4/i1_5 ), .A2(
        \SB1_1_7/buf_output[2] ), .A3(\SB1_1_5/buf_output[4] ), .ZN(
        \SB2_1_4/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_4/Component_Function_4/N2  ( .A1(\SB2_1_4/i3[0] ), .A2(
        \SB1_1_7/buf_output[2] ), .A3(\SB2_1_4/i1_7 ), .ZN(
        \SB2_1_4/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_4/Component_Function_4/N1  ( .A1(\SB2_1_4/i0[9] ), .A2(
        \SB1_1_7/buf_output[2] ), .A3(\SB2_1_4/i0[8] ), .ZN(
        \SB2_1_4/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_5/Component_Function_4/N1  ( .A1(\SB2_1_5/i0[9] ), .A2(
        \SB2_1_5/i0_0 ), .A3(\SB2_1_5/i0[8] ), .ZN(
        \SB2_1_5/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_6/Component_Function_4/N2  ( .A1(\SB2_1_6/i3[0] ), .A2(
        \SB2_1_6/i0_0 ), .A3(\SB2_1_6/i1_7 ), .ZN(
        \SB2_1_6/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_6/Component_Function_4/N1  ( .A1(\SB2_1_6/i0[9] ), .A2(
        \SB2_1_6/i0_0 ), .A3(\SB2_1_6/i0[8] ), .ZN(
        \SB2_1_6/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_7/Component_Function_4/N1  ( .A1(\SB2_1_7/i0[9] ), .A2(
        \SB2_1_7/i0_0 ), .A3(\SB2_1_7/i0[8] ), .ZN(
        \SB2_1_7/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_8/Component_Function_4/N2  ( .A1(\SB2_1_8/i3[0] ), .A2(
        \SB2_1_8/i0_0 ), .A3(\SB2_1_8/i1_7 ), .ZN(
        \SB2_1_8/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_8/Component_Function_4/N1  ( .A1(n2745), .A2(\SB2_1_8/i0_0 ), 
        .A3(\SB2_1_8/i0[8] ), .ZN(\SB2_1_8/Component_Function_4/NAND4_in[0] )
         );
  NAND3_X1 \SB2_1_11/Component_Function_4/N1  ( .A1(\SB2_1_11/i0[9] ), .A2(
        \SB2_1_11/i0_0 ), .A3(\SB2_1_11/i0[8] ), .ZN(
        \SB2_1_11/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_12/Component_Function_4/N2  ( .A1(\SB2_1_12/i3[0] ), .A2(
        \SB2_1_12/i0_0 ), .A3(\SB2_1_12/i1_7 ), .ZN(
        \SB2_1_12/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_12/Component_Function_4/N1  ( .A1(\SB2_1_12/i0[9] ), .A2(
        \SB2_1_12/i0_0 ), .A3(\SB2_1_12/i0[8] ), .ZN(
        \SB2_1_12/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_13/Component_Function_4/N2  ( .A1(n4182), .A2(
        \SB2_1_13/i0_0 ), .A3(\SB2_1_13/i1_7 ), .ZN(
        \SB2_1_13/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_15/Component_Function_4/N2  ( .A1(\SB2_1_15/i3[0] ), .A2(
        \SB2_1_15/i0_0 ), .A3(\SB2_1_15/i1_7 ), .ZN(
        \SB2_1_15/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_15/Component_Function_4/N1  ( .A1(\SB2_1_15/i0[9] ), .A2(
        \SB2_1_15/i0_0 ), .A3(\SB2_1_15/i0[8] ), .ZN(
        \SB2_1_15/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_17/Component_Function_4/N1  ( .A1(\SB2_1_17/i0[9] ), .A2(
        \SB2_1_17/i0_0 ), .A3(\SB2_1_17/i0[8] ), .ZN(
        \SB2_1_17/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_18/Component_Function_4/N1  ( .A1(\SB2_1_18/i0[9] ), .A2(
        \SB2_1_18/i0_0 ), .A3(\SB2_1_18/i0[8] ), .ZN(
        \SB2_1_18/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_20/Component_Function_4/N2  ( .A1(\SB2_1_20/i3[0] ), .A2(
        \SB2_1_20/i0_0 ), .A3(\SB2_1_20/i1_7 ), .ZN(
        \SB2_1_20/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_21/Component_Function_4/N1  ( .A1(\RI3[1][60] ), .A2(
        \SB2_1_21/i0_0 ), .A3(\SB2_1_21/i0[8] ), .ZN(
        \SB2_1_21/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_22/Component_Function_4/N2  ( .A1(\SB2_1_22/i3[0] ), .A2(
        \SB2_1_22/i0_0 ), .A3(\SB2_1_22/i1_7 ), .ZN(
        \SB2_1_22/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_22/Component_Function_4/N1  ( .A1(\SB2_1_22/i0[9] ), .A2(
        \SB2_1_22/i0_0 ), .A3(\SB2_1_22/i0[8] ), .ZN(
        \SB2_1_22/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_23/Component_Function_4/N2  ( .A1(\SB2_1_23/i3[0] ), .A2(
        \SB2_1_23/i0_0 ), .A3(\SB2_1_23/i1_7 ), .ZN(
        \SB2_1_23/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_23/Component_Function_4/N1  ( .A1(\SB2_1_23/i0[9] ), .A2(
        \SB2_1_23/i0_0 ), .A3(\SB2_1_23/i0[8] ), .ZN(
        \SB2_1_23/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_24/Component_Function_4/N2  ( .A1(\SB2_1_24/i3[0] ), .A2(
        \SB2_1_24/i0_0 ), .A3(\SB2_1_24/i1_7 ), .ZN(
        \SB2_1_24/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_25/Component_Function_4/N1  ( .A1(\SB2_1_25/i0[9] ), .A2(
        \SB2_1_25/i0_0 ), .A3(\SB2_1_25/i0[8] ), .ZN(
        \SB2_1_25/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_26/Component_Function_4/N4  ( .A1(\SB2_1_26/i1[9] ), .A2(
        \SB2_1_26/i1_5 ), .A3(\SB1_1_27/buf_output[4] ), .ZN(
        \SB2_1_26/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_26/Component_Function_4/N2  ( .A1(\SB2_1_26/i3[0] ), .A2(
        \SB2_1_26/i0_0 ), .A3(\SB2_1_26/i1_7 ), .ZN(
        \SB2_1_26/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_26/Component_Function_4/N1  ( .A1(\SB2_1_26/i0[9] ), .A2(
        \SB2_1_26/i0_0 ), .A3(\SB2_1_26/i0[8] ), .ZN(
        \SB2_1_26/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_27/Component_Function_4/N2  ( .A1(\SB2_1_27/i3[0] ), .A2(
        \SB2_1_27/i0_0 ), .A3(\SB2_1_27/i1_7 ), .ZN(
        \SB2_1_27/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_28/Component_Function_4/N2  ( .A1(\SB2_1_28/i3[0] ), .A2(
        \SB2_1_28/i0_0 ), .A3(\SB2_1_28/i1_7 ), .ZN(
        \SB2_1_28/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_28/Component_Function_4/N1  ( .A1(\SB2_1_28/i0[9] ), .A2(
        \SB2_1_28/i0_0 ), .A3(\SB2_1_28/i0[8] ), .ZN(
        \SB2_1_28/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_29/Component_Function_4/N4  ( .A1(\SB2_1_29/i1[9] ), .A2(
        \SB2_1_29/i1_5 ), .A3(\SB2_1_29/i0_4 ), .ZN(
        \SB2_1_29/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_29/Component_Function_4/N1  ( .A1(\SB2_1_29/i0[9] ), .A2(
        \SB2_1_29/i0_0 ), .A3(\SB2_1_29/i0[8] ), .ZN(
        \SB2_1_29/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_30/Component_Function_3/N3  ( .A1(\SB2_1_30/i1[9] ), .A2(
        \SB2_1_30/i1_7 ), .A3(\SB1_1_0/buf_output[3] ), .ZN(
        \SB2_1_30/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_30/Component_Function_3/N1  ( .A1(\SB2_1_30/i1[9] ), .A2(
        \SB2_1_30/i0_3 ), .A3(\SB2_1_30/i0[6] ), .ZN(
        \SB2_1_30/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_30/Component_Function_4/N2  ( .A1(\SB2_1_30/i3[0] ), .A2(
        \SB2_1_30/i0_0 ), .A3(\SB2_1_30/i1_7 ), .ZN(
        \SB2_1_30/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_30/Component_Function_4/N1  ( .A1(\SB2_1_30/i0[9] ), .A2(
        \SB2_1_30/i0_0 ), .A3(\SB2_1_30/i0[8] ), .ZN(
        \SB2_1_30/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_31/Component_Function_4/N3  ( .A1(\SB2_1_31/i0[9] ), .A2(
        \SB2_1_31/i0[10] ), .A3(\SB2_1_31/i0_3 ), .ZN(
        \SB2_1_31/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_31/Component_Function_4/N2  ( .A1(\SB2_1_31/i3[0] ), .A2(
        \SB2_1_31/i0_0 ), .A3(\SB2_1_31/i1_7 ), .ZN(
        \SB2_1_31/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_1/Component_Function_2/N1  ( .A1(\SB1_2_1/i1_5 ), .A2(
        \SB1_2_1/i0[10] ), .A3(\SB1_2_1/i1[9] ), .ZN(
        \SB1_2_1/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_1/Component_Function_4/N2  ( .A1(\SB1_2_1/i3[0] ), .A2(
        \SB1_2_1/i0_0 ), .A3(\SB1_2_1/i1_7 ), .ZN(
        \SB1_2_1/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_1/Component_Function_4/N1  ( .A1(\SB1_2_1/i0[9] ), .A2(
        \SB1_2_1/i0_0 ), .A3(\SB1_2_1/i0[8] ), .ZN(
        \SB1_2_1/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_4/Component_Function_4/N3  ( .A1(\SB1_2_4/i0[9] ), .A2(
        \SB1_2_4/i0[10] ), .A3(\SB1_2_4/i0_3 ), .ZN(
        \SB1_2_4/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_5/Component_Function_3/N2  ( .A1(\SB1_2_5/i0_0 ), .A2(
        \SB1_2_5/i0_3 ), .A3(\SB1_2_5/i0_4 ), .ZN(
        \SB1_2_5/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_7/Component_Function_3/N2  ( .A1(\SB1_2_7/i0_0 ), .A2(
        \SB1_2_7/i0_3 ), .A3(\SB1_2_7/i0_4 ), .ZN(
        \SB1_2_7/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_7/Component_Function_4/N2  ( .A1(\SB1_2_7/i3[0] ), .A2(
        \SB1_2_7/i0_0 ), .A3(\SB1_2_7/i1_7 ), .ZN(
        \SB1_2_7/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_7/Component_Function_4/N1  ( .A1(\SB1_2_7/i0[9] ), .A2(
        \SB1_2_7/i0_0 ), .A3(\SB1_2_7/i0[8] ), .ZN(
        \SB1_2_7/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_8/Component_Function_3/N2  ( .A1(\SB1_2_8/i0_0 ), .A2(
        \SB1_2_8/i0_3 ), .A3(\SB1_2_8/i0_4 ), .ZN(
        \SB1_2_8/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_8/Component_Function_4/N1  ( .A1(\SB1_2_8/i0[9] ), .A2(
        \SB1_2_8/i0_0 ), .A3(\SB1_2_8/i0[8] ), .ZN(
        \SB1_2_8/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_10/Component_Function_3/N1  ( .A1(\SB1_2_10/i1[9] ), .A2(
        \SB1_2_10/i0_3 ), .A3(\SB1_2_10/i0[6] ), .ZN(
        \SB1_2_10/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_10/Component_Function_4/N4  ( .A1(\SB1_2_10/i1[9] ), .A2(
        \SB1_2_10/i1_5 ), .A3(\SB1_2_10/i0_4 ), .ZN(
        \SB1_2_10/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_14/Component_Function_4/N1  ( .A1(\SB1_2_14/i0[9] ), .A2(
        \SB1_2_14/i0_0 ), .A3(\SB1_2_14/i0[8] ), .ZN(
        \SB1_2_14/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_15/Component_Function_4/N4  ( .A1(\SB1_2_15/i1[9] ), .A2(
        \SB1_2_15/i1_5 ), .A3(\MC_ARK_ARC_1_1/buf_output[100] ), .ZN(
        \SB1_2_15/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_17/Component_Function_4/N2  ( .A1(\SB1_2_17/i3[0] ), .A2(
        \SB1_2_17/i0_0 ), .A3(\SB1_2_17/i1_7 ), .ZN(
        \SB1_2_17/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_17/Component_Function_4/N1  ( .A1(\SB1_2_17/i0[9] ), .A2(
        \SB1_2_17/i0_0 ), .A3(\SB1_2_17/i0[8] ), .ZN(
        \SB1_2_17/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_18/Component_Function_2/N1  ( .A1(\SB1_2_18/i1_5 ), .A2(
        \SB1_2_18/i0[10] ), .A3(\SB1_2_18/i1[9] ), .ZN(
        \SB1_2_18/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_18/Component_Function_3/N2  ( .A1(\SB1_2_18/i0_0 ), .A2(
        \SB1_2_18/i0_3 ), .A3(\SB1_2_18/i0_4 ), .ZN(
        \SB1_2_18/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_19/Component_Function_2/N1  ( .A1(\SB1_2_19/i1_5 ), .A2(
        \SB1_2_19/i0[10] ), .A3(\SB1_2_19/i1[9] ), .ZN(
        \SB1_2_19/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_19/Component_Function_3/N1  ( .A1(\SB1_2_19/i1[9] ), .A2(
        \SB1_2_19/i0_3 ), .A3(\SB1_2_19/i0[6] ), .ZN(
        \SB1_2_19/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_19/Component_Function_4/N2  ( .A1(\SB1_2_19/i3[0] ), .A2(
        \SB1_2_19/i0_0 ), .A3(\SB1_2_19/i1_7 ), .ZN(
        \SB1_2_19/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_20/Component_Function_4/N2  ( .A1(\SB1_2_20/i3[0] ), .A2(
        \SB1_2_20/i0_0 ), .A3(\SB1_2_20/i1_7 ), .ZN(
        \SB1_2_20/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_20/Component_Function_4/N1  ( .A1(\SB1_2_20/i0[9] ), .A2(
        \SB1_2_20/i0_0 ), .A3(n2893), .ZN(
        \SB1_2_20/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_22/Component_Function_4/N2  ( .A1(\SB1_2_22/i3[0] ), .A2(
        \SB1_2_22/i0_0 ), .A3(\SB1_2_22/i1_7 ), .ZN(
        \SB1_2_22/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_22/Component_Function_4/N1  ( .A1(\SB1_2_22/i0[9] ), .A2(
        \SB1_2_22/i0_0 ), .A3(\SB1_2_22/i0[8] ), .ZN(
        \SB1_2_22/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_23/Component_Function_2/N3  ( .A1(\SB1_2_23/i0_3 ), .A2(
        \SB1_2_23/i0[8] ), .A3(\SB1_2_23/i0[9] ), .ZN(
        \SB1_2_23/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_23/Component_Function_4/N2  ( .A1(\SB1_2_23/i3[0] ), .A2(
        \SB1_2_23/i0_0 ), .A3(\SB1_2_23/i1_7 ), .ZN(
        \SB1_2_23/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_23/Component_Function_4/N1  ( .A1(\SB1_2_23/i0[9] ), .A2(
        \SB1_2_23/i0_0 ), .A3(\SB1_2_23/i0[8] ), .ZN(
        \SB1_2_23/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_24/Component_Function_4/N1  ( .A1(\SB1_2_24/i0[9] ), .A2(
        \SB1_2_24/i0_0 ), .A3(\SB1_2_24/i0[8] ), .ZN(
        \SB1_2_24/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_25/Component_Function_3/N1  ( .A1(\SB1_2_25/i1[9] ), .A2(
        \SB1_2_25/i0_3 ), .A3(\SB1_2_25/i0[6] ), .ZN(
        \SB1_2_25/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_27/Component_Function_2/N3  ( .A1(\SB1_2_27/i0_3 ), .A2(
        \SB1_2_27/i0[8] ), .A3(\SB1_2_27/i0[9] ), .ZN(
        \SB1_2_27/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_27/Component_Function_3/N1  ( .A1(\SB1_2_27/i1[9] ), .A2(
        \SB1_2_27/i0_3 ), .A3(\SB1_2_27/i0[6] ), .ZN(
        \SB1_2_27/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_27/Component_Function_4/N2  ( .A1(\SB1_2_27/i3[0] ), .A2(
        \SB1_2_27/i0_0 ), .A3(\SB1_2_27/i1_7 ), .ZN(
        \SB1_2_27/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_27/Component_Function_4/N1  ( .A1(\SB1_2_27/i0[9] ), .A2(
        \SB1_2_27/i0_0 ), .A3(\SB1_2_27/i0[8] ), .ZN(
        \SB1_2_27/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_28/Component_Function_3/N1  ( .A1(\SB1_2_28/i1[9] ), .A2(
        \SB1_2_28/i0_3 ), .A3(\SB1_2_28/i0[6] ), .ZN(
        \SB1_2_28/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_28/Component_Function_4/N1  ( .A1(\SB1_2_28/i0[9] ), .A2(
        \SB1_2_28/i0_0 ), .A3(\SB1_2_28/i0[8] ), .ZN(
        \SB1_2_28/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_30/Component_Function_2/N2  ( .A1(\SB1_2_30/i0_3 ), .A2(
        \SB1_2_30/i0[10] ), .A3(\SB1_2_30/i0[6] ), .ZN(
        \SB1_2_30/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_30/Component_Function_3/N2  ( .A1(\SB1_2_30/i0_0 ), .A2(
        \SB1_2_30/i0_3 ), .A3(\MC_ARK_ARC_1_1/buf_output[10] ), .ZN(
        \SB1_2_30/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_31/Component_Function_2/N2  ( .A1(\SB1_2_31/i0_3 ), .A2(
        \SB1_2_31/i0[10] ), .A3(\SB1_2_31/i0[6] ), .ZN(
        \SB1_2_31/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_31/Component_Function_4/N4  ( .A1(\SB1_2_31/i1[9] ), .A2(
        \SB1_2_31/i1_5 ), .A3(\SB1_2_31/i0_4 ), .ZN(
        \SB1_2_31/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_0/Component_Function_3/N4  ( .A1(\SB2_2_0/i1_5 ), .A2(
        \SB2_2_0/i0[8] ), .A3(\SB2_2_0/i3[0] ), .ZN(
        \SB2_2_0/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_0/Component_Function_4/N2  ( .A1(\SB2_2_0/i3[0] ), .A2(
        \SB2_2_0/i0_0 ), .A3(\SB2_2_0/i1_7 ), .ZN(
        \SB2_2_0/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_0/Component_Function_4/N1  ( .A1(\SB2_2_0/i0[9] ), .A2(
        \SB2_2_0/i0_0 ), .A3(\SB2_2_0/i0[8] ), .ZN(
        \SB2_2_0/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_2/Component_Function_4/N2  ( .A1(\SB2_2_2/i3[0] ), .A2(
        \SB2_2_2/i0_0 ), .A3(\SB2_2_2/i1_7 ), .ZN(
        \SB2_2_2/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_3/Component_Function_4/N2  ( .A1(\SB2_2_3/i3[0] ), .A2(
        \SB2_2_3/i0_0 ), .A3(\SB2_2_3/i1_7 ), .ZN(
        \SB2_2_3/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_3/Component_Function_4/N1  ( .A1(\SB2_2_3/i0[9] ), .A2(
        \SB2_2_3/i0_0 ), .A3(\SB2_2_3/i0[8] ), .ZN(
        \SB2_2_3/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_4/Component_Function_4/N2  ( .A1(\SB2_2_4/i3[0] ), .A2(
        \SB2_2_4/i0_0 ), .A3(\SB2_2_4/i1_7 ), .ZN(
        \SB2_2_4/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_4/Component_Function_4/N1  ( .A1(\SB2_2_4/i0[9] ), .A2(
        \SB2_2_4/i0_0 ), .A3(\SB2_2_4/i0[8] ), .ZN(
        \SB2_2_4/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_5/Component_Function_4/N2  ( .A1(\SB2_2_5/i3[0] ), .A2(
        \SB2_2_5/i0_0 ), .A3(\SB2_2_5/i1_7 ), .ZN(
        \SB2_2_5/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_7/Component_Function_3/N1  ( .A1(\SB2_2_7/i1[9] ), .A2(
        \SB2_2_7/i0_3 ), .A3(\SB2_2_7/i0[6] ), .ZN(
        \SB2_2_7/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_8/Component_Function_4/N2  ( .A1(\SB2_2_8/i3[0] ), .A2(
        \SB2_2_8/i0_0 ), .A3(\SB2_2_8/i1_7 ), .ZN(
        \SB2_2_8/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_9/Component_Function_4/N2  ( .A1(\SB2_2_9/i3[0] ), .A2(
        \SB2_2_9/i0_0 ), .A3(\SB2_2_9/i1_7 ), .ZN(
        \SB2_2_9/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_11/Component_Function_4/N4  ( .A1(n5515), .A2(
        \SB2_2_11/i1_5 ), .A3(\SB2_2_11/i0_4 ), .ZN(
        \SB2_2_11/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_11/Component_Function_4/N1  ( .A1(\SB2_2_11/i0[9] ), .A2(
        \SB2_2_11/i0_0 ), .A3(\SB2_2_11/i0[8] ), .ZN(
        \SB2_2_11/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_12/Component_Function_4/N2  ( .A1(\SB2_2_12/i3[0] ), .A2(
        \SB2_2_12/i0_0 ), .A3(\SB2_2_12/i1_7 ), .ZN(
        \SB2_2_12/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_12/Component_Function_4/N1  ( .A1(\SB2_2_12/i0[9] ), .A2(
        \SB2_2_12/i0_0 ), .A3(\SB2_2_12/i0[8] ), .ZN(
        \SB2_2_12/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_14/Component_Function_4/N2  ( .A1(\SB2_2_14/i3[0] ), .A2(
        \SB2_2_14/i0_0 ), .A3(\SB2_2_14/i1_7 ), .ZN(
        \SB2_2_14/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_15/Component_Function_3/N3  ( .A1(\SB2_2_15/i1[9] ), .A2(
        \SB2_2_15/i1_7 ), .A3(\SB2_2_15/i0[10] ), .ZN(
        \SB2_2_15/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_15/Component_Function_4/N4  ( .A1(\SB2_2_15/i1[9] ), .A2(
        \SB2_2_15/i1_5 ), .A3(\SB2_2_15/i0_4 ), .ZN(
        \SB2_2_15/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_15/Component_Function_4/N1  ( .A1(\SB2_2_15/i0[9] ), .A2(
        \SB2_2_15/i0_0 ), .A3(\SB2_2_15/i0[8] ), .ZN(
        \SB2_2_15/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_16/Component_Function_4/N4  ( .A1(\SB2_2_16/i1[9] ), .A2(
        \SB2_2_16/i1_5 ), .A3(\SB2_2_16/i0_4 ), .ZN(
        \SB2_2_16/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_16/Component_Function_4/N2  ( .A1(\SB2_2_16/i3[0] ), .A2(
        \SB2_2_16/i0_0 ), .A3(\SB2_2_16/i1_7 ), .ZN(
        \SB2_2_16/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_16/Component_Function_4/N1  ( .A1(\SB2_2_16/i0[9] ), .A2(
        \SB2_2_16/i0_0 ), .A3(\SB2_2_16/i0[8] ), .ZN(
        \SB2_2_16/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_17/Component_Function_4/N2  ( .A1(\SB2_2_17/i3[0] ), .A2(
        \SB2_2_17/i0_0 ), .A3(\SB2_2_17/i1_7 ), .ZN(
        \SB2_2_17/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_17/Component_Function_4/N1  ( .A1(\SB2_2_17/i0[9] ), .A2(
        \SB2_2_17/i0_0 ), .A3(\SB2_2_17/i0[8] ), .ZN(
        \SB2_2_17/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_18/Component_Function_4/N1  ( .A1(\SB2_2_18/i0[9] ), .A2(
        \SB2_2_18/i0_0 ), .A3(\SB2_2_18/i0[8] ), .ZN(
        \SB2_2_18/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_19/Component_Function_4/N1  ( .A1(\SB2_2_19/i0[9] ), .A2(
        \SB2_2_19/i0_0 ), .A3(\SB2_2_19/i0[8] ), .ZN(
        \SB2_2_19/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_20/Component_Function_4/N2  ( .A1(\SB2_2_20/i3[0] ), .A2(
        \SB2_2_20/i0_0 ), .A3(\SB2_2_20/i1_7 ), .ZN(
        \SB2_2_20/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_20/Component_Function_4/N1  ( .A1(\SB2_2_20/i0[9] ), .A2(
        \SB2_2_20/i0_0 ), .A3(\SB2_2_20/i0[8] ), .ZN(
        \SB2_2_20/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_21/Component_Function_4/N4  ( .A1(\SB2_2_21/i1[9] ), .A2(
        \SB2_2_21/i1_5 ), .A3(\SB2_2_21/i0_4 ), .ZN(
        \SB2_2_21/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_22/Component_Function_4/N4  ( .A1(\SB2_2_22/i1[9] ), .A2(
        \SB2_2_22/i1_5 ), .A3(\SB2_2_22/i0_4 ), .ZN(
        \SB2_2_22/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_22/Component_Function_4/N1  ( .A1(\SB2_2_22/i0[9] ), .A2(
        \SB2_2_22/i0_0 ), .A3(\SB2_2_22/i0[8] ), .ZN(
        \SB2_2_22/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_23/Component_Function_4/N1  ( .A1(\SB2_2_23/i0[9] ), .A2(
        \SB2_2_23/i0_0 ), .A3(\SB2_2_23/i0[8] ), .ZN(
        \SB2_2_23/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_24/Component_Function_4/N2  ( .A1(\SB2_2_24/i3[0] ), .A2(
        \SB2_2_24/i0_0 ), .A3(\SB2_2_24/i1_7 ), .ZN(
        \SB2_2_24/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_24/Component_Function_4/N1  ( .A1(\SB2_2_24/i0[9] ), .A2(
        \SB2_2_24/i0_0 ), .A3(\SB2_2_24/i0[8] ), .ZN(
        \SB2_2_24/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_25/Component_Function_4/N2  ( .A1(\SB2_2_25/i3[0] ), .A2(
        \SB2_2_25/i0_0 ), .A3(\SB2_2_25/i1_7 ), .ZN(
        \SB2_2_25/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_25/Component_Function_4/N1  ( .A1(\SB2_2_25/i0[9] ), .A2(
        \SB2_2_25/i0_0 ), .A3(\SB2_2_25/i0[8] ), .ZN(
        \SB2_2_25/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_26/Component_Function_4/N3  ( .A1(\SB2_2_26/i0[9] ), .A2(
        \SB2_2_26/i0[10] ), .A3(\SB2_2_26/i0_3 ), .ZN(
        \SB2_2_26/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_28/Component_Function_4/N4  ( .A1(\SB2_2_28/i1[9] ), .A2(
        \SB2_2_28/i1_5 ), .A3(\SB2_2_28/i0_4 ), .ZN(
        \SB2_2_28/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_28/Component_Function_4/N2  ( .A1(\SB2_2_28/i3[0] ), .A2(
        \SB2_2_28/i0_0 ), .A3(\SB2_2_28/i1_7 ), .ZN(
        \SB2_2_28/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_28/Component_Function_4/N1  ( .A1(\SB2_2_28/i0[9] ), .A2(
        \SB2_2_28/i0_0 ), .A3(\SB2_2_28/i0[8] ), .ZN(
        \SB2_2_28/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_29/Component_Function_2/N1  ( .A1(\SB2_2_29/i1_5 ), .A2(
        \SB2_2_29/i0[10] ), .A3(\SB2_2_29/i1[9] ), .ZN(
        \SB2_2_29/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_29/Component_Function_4/N4  ( .A1(\SB2_2_29/i1[9] ), .A2(
        \SB2_2_29/i1_5 ), .A3(n1837), .ZN(
        \SB2_2_29/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_29/Component_Function_4/N2  ( .A1(\SB2_2_29/i3[0] ), .A2(
        \SB2_2_29/i0_0 ), .A3(\SB2_2_29/i1_7 ), .ZN(
        \SB2_2_29/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_29/Component_Function_4/N1  ( .A1(\SB2_2_29/i0[9] ), .A2(
        \SB2_2_29/i0_0 ), .A3(\SB2_2_29/i0[8] ), .ZN(
        \SB2_2_29/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_30/Component_Function_3/N4  ( .A1(\SB2_2_30/i1_5 ), .A2(
        \SB2_2_30/i0[8] ), .A3(\SB2_2_30/i3[0] ), .ZN(
        \SB2_2_30/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_30/Component_Function_4/N4  ( .A1(\SB2_2_30/i1[9] ), .A2(
        \SB2_2_30/i1_5 ), .A3(n2343), .ZN(
        \SB2_2_30/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_30/Component_Function_4/N1  ( .A1(\SB2_2_30/i0[9] ), .A2(
        \SB2_2_30/i0_0 ), .A3(\SB2_2_30/i0[8] ), .ZN(
        \SB2_2_30/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_31/Component_Function_4/N1  ( .A1(\SB2_2_31/i0[9] ), .A2(
        \SB2_2_31/i0_0 ), .A3(\SB2_2_31/i0[8] ), .ZN(
        \SB2_2_31/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_0/Component_Function_2/N1  ( .A1(\SB1_3_0/i1_5 ), .A2(
        \SB1_3_0/i0[10] ), .A3(\SB1_3_0/i1[9] ), .ZN(
        \SB1_3_0/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_0/Component_Function_4/N4  ( .A1(\SB1_3_0/i1[9] ), .A2(
        \SB1_3_0/i1_5 ), .A3(\SB1_3_0/i0_4 ), .ZN(
        \SB1_3_0/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_0/Component_Function_4/N2  ( .A1(\SB1_3_0/i3[0] ), .A2(
        \SB1_3_0/i0_0 ), .A3(\SB1_3_0/i1_7 ), .ZN(
        \SB1_3_0/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_0/Component_Function_4/N1  ( .A1(\SB1_3_0/i0[9] ), .A2(
        \SB1_3_0/i0_0 ), .A3(\SB1_3_0/i0[8] ), .ZN(
        \SB1_3_0/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_1/Component_Function_2/N1  ( .A1(\SB1_3_1/i1_5 ), .A2(
        \SB1_3_1/i0[10] ), .A3(\SB1_3_1/i1[9] ), .ZN(
        \SB1_3_1/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_1/Component_Function_4/N1  ( .A1(\SB1_3_1/i0[9] ), .A2(
        \SB1_3_1/i0_0 ), .A3(\SB1_3_1/i0[8] ), .ZN(
        \SB1_3_1/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_2/Component_Function_3/N2  ( .A1(\SB1_3_2/i0_0 ), .A2(
        \SB1_3_2/i0_3 ), .A3(\SB1_3_2/i0_4 ), .ZN(
        \SB1_3_2/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_2/Component_Function_4/N2  ( .A1(\SB1_3_2/i3[0] ), .A2(
        \SB1_3_2/i0_0 ), .A3(\SB1_3_2/i1_7 ), .ZN(
        \SB1_3_2/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_3/Component_Function_2/N1  ( .A1(\SB1_3_3/i1_5 ), .A2(
        \SB1_3_3/i0[10] ), .A3(\SB1_3_3/i1[9] ), .ZN(
        \SB1_3_3/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_3/Component_Function_4/N2  ( .A1(\SB1_3_3/i3[0] ), .A2(
        \SB1_3_3/i0_0 ), .A3(\SB1_3_3/i1_7 ), .ZN(
        \SB1_3_3/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_3/Component_Function_4/N1  ( .A1(\SB1_3_3/i0[9] ), .A2(
        \SB1_3_3/i0_0 ), .A3(\SB1_3_3/i0[8] ), .ZN(
        \SB1_3_3/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_5/Component_Function_3/N1  ( .A1(\SB1_3_5/i1[9] ), .A2(
        \SB1_3_5/i0_3 ), .A3(\SB1_3_5/i0[6] ), .ZN(
        \SB1_3_5/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_5/Component_Function_4/N2  ( .A1(\SB1_3_5/i3[0] ), .A2(
        \SB1_3_5/i0_0 ), .A3(\SB1_3_5/i1_7 ), .ZN(
        \SB1_3_5/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_5/Component_Function_4/N1  ( .A1(\SB1_3_5/i0[9] ), .A2(
        \SB1_3_5/i0_0 ), .A3(\SB1_3_5/i0[8] ), .ZN(
        \SB1_3_5/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_6/Component_Function_2/N2  ( .A1(\SB1_3_6/i0_3 ), .A2(
        \SB1_3_6/i0[10] ), .A3(\SB1_3_6/i0[6] ), .ZN(
        \SB1_3_6/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_6/Component_Function_2/N1  ( .A1(\SB1_3_6/i1_5 ), .A2(
        \SB1_3_6/i0[10] ), .A3(\SB1_3_6/i1[9] ), .ZN(
        \SB1_3_6/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_6/Component_Function_4/N2  ( .A1(\SB1_3_6/i3[0] ), .A2(
        \SB1_3_6/i0_0 ), .A3(\SB1_3_6/i1_7 ), .ZN(
        \SB1_3_6/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_6/Component_Function_4/N1  ( .A1(\SB1_3_6/i0[9] ), .A2(
        \SB1_3_6/i0_0 ), .A3(\SB1_3_6/i0[8] ), .ZN(
        \SB1_3_6/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_7/Component_Function_4/N4  ( .A1(\SB1_3_7/i1[9] ), .A2(
        \SB1_3_7/i1_5 ), .A3(\SB1_3_7/i0_4 ), .ZN(
        \SB1_3_7/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_9/Component_Function_4/N2  ( .A1(\SB1_3_9/i3[0] ), .A2(
        \SB1_3_9/i0_0 ), .A3(\SB1_3_9/i1_7 ), .ZN(
        \SB1_3_9/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_10/Component_Function_4/N2  ( .A1(\SB1_3_10/i3[0] ), .A2(
        \SB1_3_10/i0_0 ), .A3(\SB1_3_10/i1_7 ), .ZN(
        \SB1_3_10/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_10/Component_Function_4/N1  ( .A1(\SB1_3_10/i0[9] ), .A2(
        \SB1_3_10/i0_0 ), .A3(\SB1_3_10/i0[8] ), .ZN(
        \SB1_3_10/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_11/Component_Function_4/N2  ( .A1(\SB1_3_11/i3[0] ), .A2(
        \SB1_3_11/i0_0 ), .A3(\SB1_3_11/i1_7 ), .ZN(
        \SB1_3_11/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_11/Component_Function_4/N1  ( .A1(\SB1_3_11/i0[9] ), .A2(
        \SB1_3_11/i0_0 ), .A3(\SB1_3_11/i0[8] ), .ZN(
        \SB1_3_11/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_12/Component_Function_2/N2  ( .A1(\SB1_3_12/i0_3 ), .A2(
        \SB1_3_12/i0[10] ), .A3(\SB1_3_12/i0[6] ), .ZN(
        \SB1_3_12/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_13/Component_Function_2/N1  ( .A1(\SB1_3_13/i1_5 ), .A2(
        \SB1_3_13/i0[10] ), .A3(\SB1_3_13/i1[9] ), .ZN(
        \SB1_3_13/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_13/Component_Function_3/N3  ( .A1(\SB1_3_13/i1[9] ), .A2(
        \SB1_3_13/i1_7 ), .A3(\SB1_3_13/i0[10] ), .ZN(
        \SB1_3_13/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_13/Component_Function_4/N1  ( .A1(\SB1_3_13/i0[9] ), .A2(
        \SB1_3_13/i0_0 ), .A3(\SB1_3_13/i0[8] ), .ZN(
        \SB1_3_13/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_14/Component_Function_3/N2  ( .A1(\SB1_3_14/i0_0 ), .A2(
        \SB1_3_14/i0_3 ), .A3(\SB1_3_14/i0_4 ), .ZN(
        \SB1_3_14/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_14/Component_Function_4/N4  ( .A1(\SB1_3_14/i1[9] ), .A2(
        \SB1_3_14/i1_5 ), .A3(\SB1_3_14/i0_4 ), .ZN(
        \SB1_3_14/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_15/Component_Function_4/N2  ( .A1(\SB1_3_15/i3[0] ), .A2(
        \SB1_3_15/i0_0 ), .A3(\SB1_3_15/i1_7 ), .ZN(
        \SB1_3_15/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_15/Component_Function_4/N1  ( .A1(\SB1_3_15/i0[9] ), .A2(
        \SB1_3_15/i0_0 ), .A3(\SB1_3_15/i0[8] ), .ZN(
        \SB1_3_15/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_16/Component_Function_3/N2  ( .A1(\SB1_3_16/i0_0 ), .A2(
        \SB1_3_16/i0_3 ), .A3(\SB1_3_16/i0_4 ), .ZN(
        \SB1_3_16/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_16/Component_Function_4/N4  ( .A1(\SB1_3_16/i1[9] ), .A2(
        \SB1_3_16/i1_5 ), .A3(\SB1_3_16/i0_4 ), .ZN(
        \SB1_3_16/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_17/Component_Function_2/N3  ( .A1(\SB1_3_17/i0_3 ), .A2(
        \SB1_3_17/i0[8] ), .A3(\SB1_3_17/i0[9] ), .ZN(
        \SB1_3_17/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_18/Component_Function_2/N2  ( .A1(\SB1_3_18/i0_3 ), .A2(
        \SB1_3_18/i0[10] ), .A3(\SB1_3_18/i0[6] ), .ZN(
        \SB1_3_18/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_18/Component_Function_4/N1  ( .A1(\SB1_3_18/i0[9] ), .A2(
        \SB1_3_18/i0_0 ), .A3(\SB1_3_18/i0[8] ), .ZN(
        \SB1_3_18/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_19/Component_Function_4/N2  ( .A1(\SB1_3_19/i3[0] ), .A2(
        \SB1_3_19/i0_0 ), .A3(\SB1_3_19/i1_7 ), .ZN(
        \SB1_3_19/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_20/Component_Function_2/N2  ( .A1(\SB1_3_20/i0_3 ), .A2(
        \SB1_3_20/i0[10] ), .A3(\SB1_3_20/i0[6] ), .ZN(
        \SB1_3_20/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_20/Component_Function_2/N1  ( .A1(\SB1_3_20/i1_5 ), .A2(
        \SB1_3_20/i0[10] ), .A3(\SB1_3_20/i1[9] ), .ZN(
        \SB1_3_20/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_20/Component_Function_3/N1  ( .A1(\SB1_3_20/i1[9] ), .A2(
        \SB1_3_20/i0_3 ), .A3(\SB1_3_20/i0[6] ), .ZN(
        \SB1_3_20/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_20/Component_Function_4/N1  ( .A1(\SB1_3_20/i0[9] ), .A2(
        \SB1_3_20/i0_0 ), .A3(\SB1_3_20/i0[8] ), .ZN(
        \SB1_3_20/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_21/Component_Function_2/N2  ( .A1(\SB1_3_21/i0_3 ), .A2(
        \SB1_3_21/i0[10] ), .A3(\SB1_3_21/i0[6] ), .ZN(
        \SB1_3_21/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_23/Component_Function_4/N1  ( .A1(\SB1_3_23/i0[9] ), .A2(
        \SB1_3_23/i0_0 ), .A3(\SB1_3_23/i0[8] ), .ZN(
        \SB1_3_23/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_24/Component_Function_4/N2  ( .A1(\SB1_3_24/i3[0] ), .A2(
        \SB1_3_24/i0_0 ), .A3(\SB1_3_24/i1_7 ), .ZN(
        \SB1_3_24/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_24/Component_Function_4/N1  ( .A1(\SB1_3_24/i0[9] ), .A2(
        \SB1_3_24/i0_0 ), .A3(\SB1_3_24/i0[8] ), .ZN(
        \SB1_3_24/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_25/Component_Function_2/N3  ( .A1(\SB1_3_25/i0_3 ), .A2(
        \SB1_3_25/i0[8] ), .A3(\SB1_3_25/i0[9] ), .ZN(
        \SB1_3_25/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_25/Component_Function_2/N2  ( .A1(\SB1_3_25/i0_3 ), .A2(
        \SB1_3_25/i0[10] ), .A3(\SB1_3_25/i0[6] ), .ZN(
        \SB1_3_25/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_25/Component_Function_4/N1  ( .A1(\SB1_3_25/i0[9] ), .A2(
        \SB1_3_25/i0_0 ), .A3(\SB1_3_25/i0[8] ), .ZN(
        \SB1_3_25/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_27/Component_Function_2/N2  ( .A1(\SB1_3_27/i0_3 ), .A2(
        \SB1_3_27/i0[10] ), .A3(\SB1_3_27/i0[6] ), .ZN(
        \SB1_3_27/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_27/Component_Function_2/N1  ( .A1(\SB1_3_27/i1_5 ), .A2(
        \SB1_3_27/i0[10] ), .A3(\SB1_3_27/i1[9] ), .ZN(
        \SB1_3_27/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_28/Component_Function_4/N1  ( .A1(\SB1_3_28/i0[9] ), .A2(
        \SB1_3_28/i0_0 ), .A3(\SB1_3_28/i0[8] ), .ZN(
        \SB1_3_28/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_30/Component_Function_4/N2  ( .A1(\SB1_3_30/i3[0] ), .A2(
        \SB1_3_30/i0_0 ), .A3(\SB1_3_30/i1_7 ), .ZN(
        \SB1_3_30/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_30/Component_Function_4/N1  ( .A1(\SB1_3_30/i0[9] ), .A2(
        \SB1_3_30/i0_0 ), .A3(\SB1_3_30/i0[8] ), .ZN(
        \SB1_3_30/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_0/Component_Function_4/N2  ( .A1(\SB2_3_0/i3[0] ), .A2(
        \SB2_3_0/i0_0 ), .A3(\SB2_3_0/i1_7 ), .ZN(
        \SB2_3_0/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_0/Component_Function_4/N1  ( .A1(\SB2_3_0/i0[9] ), .A2(
        \SB2_3_0/i0_0 ), .A3(n5513), .ZN(
        \SB2_3_0/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_1/Component_Function_4/N1  ( .A1(\SB2_3_1/i0[9] ), .A2(
        \SB2_3_1/i0_0 ), .A3(\SB2_3_1/i0[8] ), .ZN(
        \SB2_3_1/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_2/Component_Function_4/N4  ( .A1(\SB2_3_2/i1[9] ), .A2(
        \SB2_3_2/i1_5 ), .A3(\SB2_3_2/i0_4 ), .ZN(
        \SB2_3_2/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_3/Component_Function_4/N1  ( .A1(\SB2_3_3/i0[9] ), .A2(
        \SB2_3_3/i0_0 ), .A3(\SB2_3_3/i0[8] ), .ZN(
        \SB2_3_3/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_4/Component_Function_4/N4  ( .A1(\SB2_3_4/i1[9] ), .A2(n5519), .A3(\SB2_3_4/i0_4 ), .ZN(\SB2_3_4/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_4/Component_Function_4/N2  ( .A1(\SB2_3_4/i3[0] ), .A2(
        \SB2_3_4/i0_0 ), .A3(\SB2_3_4/i1_7 ), .ZN(
        \SB2_3_4/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_4/Component_Function_4/N1  ( .A1(\SB2_3_4/i0[9] ), .A2(
        \SB2_3_4/i0_0 ), .A3(\SB2_3_4/i0[8] ), .ZN(
        \SB2_3_4/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_5/Component_Function_4/N4  ( .A1(n3671), .A2(\SB2_3_5/i1_5 ), 
        .A3(\SB2_3_5/i0_4 ), .ZN(\SB2_3_5/Component_Function_4/NAND4_in[3] )
         );
  NAND3_X1 \SB2_3_5/Component_Function_4/N1  ( .A1(\SB2_3_5/i0[9] ), .A2(
        \SB2_3_5/i0_0 ), .A3(\SB2_3_5/i0[8] ), .ZN(
        \SB2_3_5/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_7/Component_Function_4/N1  ( .A1(\SB2_3_7/i0[9] ), .A2(
        \SB2_3_7/i0_0 ), .A3(\SB2_3_7/i0[8] ), .ZN(
        \SB2_3_7/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_8/Component_Function_2/N3  ( .A1(\SB2_3_8/i0_3 ), .A2(
        \SB2_3_8/i0[8] ), .A3(\SB2_3_8/i0[9] ), .ZN(
        \SB2_3_8/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_8/Component_Function_4/N4  ( .A1(n3669), .A2(\SB2_3_8/i1_5 ), 
        .A3(\SB1_3_9/buf_output[4] ), .ZN(
        \SB2_3_8/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_8/Component_Function_4/N1  ( .A1(\SB2_3_8/i0[9] ), .A2(
        \SB2_3_8/i0_0 ), .A3(\SB2_3_8/i0[8] ), .ZN(
        \SB2_3_8/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_9/Component_Function_2/N3  ( .A1(\SB2_3_9/i0_3 ), .A2(
        \SB2_3_9/i0[8] ), .A3(\SB2_3_9/i0[9] ), .ZN(
        \SB2_3_9/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_9/Component_Function_3/N2  ( .A1(\SB2_3_9/i0_0 ), .A2(
        \SB2_3_9/i0_3 ), .A3(\SB2_3_9/i0_4 ), .ZN(
        \SB2_3_9/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_9/Component_Function_3/N1  ( .A1(\SB2_3_9/i1[9] ), .A2(
        \SB2_3_9/i0_3 ), .A3(\SB2_3_9/i0[6] ), .ZN(
        \SB2_3_9/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_9/Component_Function_4/N2  ( .A1(\SB2_3_9/i3[0] ), .A2(
        \SB2_3_9/i0_0 ), .A3(\SB2_3_9/i1_7 ), .ZN(
        \SB2_3_9/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_10/Component_Function_3/N3  ( .A1(\SB2_3_10/i1[9] ), .A2(
        \SB2_3_10/i1_7 ), .A3(\SB2_3_10/i0[10] ), .ZN(
        \SB2_3_10/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_10/Component_Function_4/N4  ( .A1(\SB2_3_10/i1[9] ), .A2(
        \SB2_3_10/i1_5 ), .A3(\SB2_3_10/i0_4 ), .ZN(
        \SB2_3_10/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_10/Component_Function_4/N2  ( .A1(\SB2_3_10/i3[0] ), .A2(
        \SB2_3_10/i0_0 ), .A3(\SB2_3_10/i1_7 ), .ZN(
        \SB2_3_10/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_10/Component_Function_4/N1  ( .A1(\SB2_3_10/i0[9] ), .A2(
        \SB2_3_10/i0_0 ), .A3(\SB2_3_10/i0[8] ), .ZN(
        \SB2_3_10/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_11/Component_Function_4/N4  ( .A1(\SB2_3_11/i1[9] ), .A2(
        n4768), .A3(n3645), .ZN(\SB2_3_11/Component_Function_4/NAND4_in[3] )
         );
  NAND3_X1 \SB2_3_11/Component_Function_4/N1  ( .A1(\SB2_3_11/i0[9] ), .A2(
        \SB2_3_11/i0_0 ), .A3(\SB2_3_11/i0[8] ), .ZN(
        \SB2_3_11/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_12/Component_Function_4/N4  ( .A1(\SB2_3_12/i1[9] ), .A2(
        \SB2_3_12/i1_5 ), .A3(\SB2_3_12/i0_4 ), .ZN(
        \SB2_3_12/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_12/Component_Function_4/N2  ( .A1(\SB2_3_12/i3[0] ), .A2(
        \SB2_3_12/i0_0 ), .A3(\SB2_3_12/i1_7 ), .ZN(
        \SB2_3_12/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_12/Component_Function_4/N1  ( .A1(n1603), .A2(
        \SB2_3_12/i0_0 ), .A3(n3651), .ZN(
        \SB2_3_12/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_13/Component_Function_4/N2  ( .A1(\SB2_3_13/i3[0] ), .A2(
        \SB2_3_13/i0_0 ), .A3(\SB2_3_13/i1_7 ), .ZN(
        \SB2_3_13/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_13/Component_Function_4/N1  ( .A1(\SB2_3_13/i0[9] ), .A2(
        \SB2_3_13/i0_0 ), .A3(\SB2_3_13/i0[8] ), .ZN(
        \SB2_3_13/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_14/Component_Function_4/N2  ( .A1(\SB2_3_14/i3[0] ), .A2(
        \SB2_3_14/i0_0 ), .A3(\SB2_3_14/i1_7 ), .ZN(
        \SB2_3_14/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_14/Component_Function_4/N1  ( .A1(\SB2_3_14/i0[9] ), .A2(
        \SB2_3_14/i0_0 ), .A3(\SB2_3_14/i0[8] ), .ZN(
        \SB2_3_14/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_15/Component_Function_4/N2  ( .A1(\SB2_3_15/i3[0] ), .A2(
        \SB2_3_15/i0_0 ), .A3(\SB2_3_15/i1_7 ), .ZN(
        \SB2_3_15/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_15/Component_Function_4/N1  ( .A1(\SB2_3_15/i0[9] ), .A2(
        \SB2_3_15/i0_0 ), .A3(n3670), .ZN(
        \SB2_3_15/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_16/Component_Function_4/N2  ( .A1(\SB2_3_16/i3[0] ), .A2(
        \SB2_3_16/i0_0 ), .A3(\SB2_3_16/i1_7 ), .ZN(
        \SB2_3_16/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_18/Component_Function_4/N2  ( .A1(\SB2_3_18/i3[0] ), .A2(
        \SB2_3_18/i0_0 ), .A3(\SB2_3_18/i1_7 ), .ZN(
        \SB2_3_18/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_18/Component_Function_4/N1  ( .A1(\SB2_3_18/i0[9] ), .A2(
        \SB2_3_18/i0_0 ), .A3(\SB2_3_18/i0[8] ), .ZN(
        \SB2_3_18/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_19/Component_Function_4/N4  ( .A1(n5494), .A2(
        \SB2_3_19/i1_5 ), .A3(\SB2_3_19/i0_4 ), .ZN(
        \SB2_3_19/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_19/Component_Function_4/N2  ( .A1(\SB2_3_19/i3[0] ), .A2(
        \SB2_3_19/i0_0 ), .A3(\SB2_3_19/i1_7 ), .ZN(
        \SB2_3_19/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_19/Component_Function_4/N1  ( .A1(\SB2_3_19/i0[9] ), .A2(
        \SB2_3_19/i0_0 ), .A3(\SB2_3_19/i0[8] ), .ZN(
        \SB2_3_19/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_20/Component_Function_3/N2  ( .A1(\SB2_3_20/i0_0 ), .A2(
        \SB2_3_20/i0_3 ), .A3(\SB2_3_20/i0_4 ), .ZN(
        \SB2_3_20/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_20/Component_Function_4/N2  ( .A1(\SB2_3_20/i3[0] ), .A2(
        \SB2_3_20/i0_0 ), .A3(\SB2_3_20/i1_7 ), .ZN(
        \SB2_3_20/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_20/Component_Function_4/N1  ( .A1(\SB2_3_20/i0[9] ), .A2(
        \SB2_3_20/i0_0 ), .A3(\SB2_3_20/i0[8] ), .ZN(
        \SB2_3_20/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_21/Component_Function_2/N1  ( .A1(\SB2_3_21/i1_5 ), .A2(
        \SB2_3_21/i0[10] ), .A3(\SB2_3_21/i1[9] ), .ZN(
        \SB2_3_21/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_21/Component_Function_3/N1  ( .A1(\SB2_3_21/i1[9] ), .A2(
        \SB2_3_21/i0_3 ), .A3(\SB2_3_21/i0[6] ), .ZN(
        \SB2_3_21/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_21/Component_Function_4/N3  ( .A1(\SB2_3_21/i0[9] ), .A2(
        \SB2_3_21/i0[10] ), .A3(\SB2_3_21/i0_3 ), .ZN(
        \SB2_3_21/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_21/Component_Function_4/N2  ( .A1(\SB2_3_21/i3[0] ), .A2(
        \SB2_3_21/i0_0 ), .A3(\SB2_3_21/i1_7 ), .ZN(
        \SB2_3_21/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_21/Component_Function_4/N1  ( .A1(\SB2_3_21/i0[9] ), .A2(
        \SB2_3_21/i0_0 ), .A3(\SB2_3_21/i0[8] ), .ZN(
        \SB2_3_21/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_22/Component_Function_4/N2  ( .A1(\SB2_3_22/i3[0] ), .A2(
        \SB2_3_22/i0_0 ), .A3(\SB2_3_22/i1_7 ), .ZN(
        \SB2_3_22/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_22/Component_Function_4/N1  ( .A1(\SB2_3_22/i0[9] ), .A2(
        \SB2_3_22/i0_0 ), .A3(\SB2_3_22/i0[8] ), .ZN(
        \SB2_3_22/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_23/Component_Function_4/N1  ( .A1(\SB2_3_23/i0[9] ), .A2(
        \SB2_3_23/i0_0 ), .A3(\SB2_3_23/i0[8] ), .ZN(
        \SB2_3_23/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_24/Component_Function_2/N2  ( .A1(\SB2_3_24/i0_3 ), .A2(
        \SB1_3_26/buf_output[3] ), .A3(\SB1_3_28/buf_output[1] ), .ZN(
        \SB2_3_24/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_24/Component_Function_4/N4  ( .A1(\SB2_3_24/i1[9] ), .A2(
        \SB2_3_24/i1_5 ), .A3(\SB2_3_24/i0_4 ), .ZN(
        \SB2_3_24/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_24/Component_Function_4/N2  ( .A1(\SB2_3_24/i3[0] ), .A2(
        \SB2_3_24/i0_0 ), .A3(\SB2_3_24/i1_7 ), .ZN(
        \SB2_3_24/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_24/Component_Function_4/N1  ( .A1(\SB2_3_24/i0[9] ), .A2(
        \SB2_3_24/i0_0 ), .A3(n2906), .ZN(
        \SB2_3_24/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_25/Component_Function_4/N1  ( .A1(\SB2_3_25/i0[9] ), .A2(
        \SB2_3_25/i0_0 ), .A3(\SB2_3_25/i0[8] ), .ZN(
        \SB2_3_25/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_26/Component_Function_4/N2  ( .A1(\SB2_3_26/i3[0] ), .A2(
        \SB2_3_26/i0_0 ), .A3(\SB2_3_26/i1_7 ), .ZN(
        \SB2_3_26/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_26/Component_Function_4/N1  ( .A1(\SB2_3_26/i0[9] ), .A2(
        \SB2_3_26/i0_0 ), .A3(n4750), .ZN(
        \SB2_3_26/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_27/Component_Function_4/N2  ( .A1(\SB2_3_27/i3[0] ), .A2(
        \SB2_3_27/i0_0 ), .A3(\SB2_3_27/i1_7 ), .ZN(
        \SB2_3_27/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_27/Component_Function_4/N1  ( .A1(\RI3[3][24] ), .A2(
        \SB2_3_27/i0_0 ), .A3(\SB2_3_27/i0[8] ), .ZN(
        \SB2_3_27/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_28/Component_Function_4/N2  ( .A1(\SB2_3_28/i3[0] ), .A2(
        \SB2_3_28/i0_0 ), .A3(\SB2_3_28/i1_7 ), .ZN(
        \SB2_3_28/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_28/Component_Function_4/N1  ( .A1(\SB2_3_28/i0[9] ), .A2(
        n5489), .A3(\SB2_3_28/i0[8] ), .ZN(
        \SB2_3_28/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_29/Component_Function_4/N1  ( .A1(\SB2_3_29/i0[9] ), .A2(
        \SB2_3_29/i0_0 ), .A3(\SB2_3_29/i0[8] ), .ZN(
        \SB2_3_29/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_30/Component_Function_4/N2  ( .A1(\SB2_3_30/i3[0] ), .A2(
        \SB2_3_30/i0_0 ), .A3(\SB2_3_30/i1_7 ), .ZN(
        \SB2_3_30/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_30/Component_Function_4/N1  ( .A1(\SB2_3_30/i0[9] ), .A2(
        \SB2_3_30/i0_0 ), .A3(\SB2_3_30/i0[8] ), .ZN(
        \SB2_3_30/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_0/Component_Function_4/N4  ( .A1(\SB3_0/i1[9] ), .A2(
        \SB3_0/i1_5 ), .A3(\SB3_0/i0_4 ), .ZN(
        \SB3_0/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_0/Component_Function_4/N2  ( .A1(\SB3_0/i3[0] ), .A2(
        \SB3_0/i0_0 ), .A3(\SB3_0/i1_7 ), .ZN(
        \SB3_0/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_0/Component_Function_4/N1  ( .A1(\SB3_0/i0[9] ), .A2(
        \SB3_0/i0_0 ), .A3(\SB3_0/i0[8] ), .ZN(
        \SB3_0/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_1/Component_Function_2/N2  ( .A1(\SB3_1/i0_3 ), .A2(
        \SB3_1/i0[10] ), .A3(\SB3_1/i0[6] ), .ZN(
        \SB3_1/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_2/Component_Function_3/N2  ( .A1(\SB3_2/i0_0 ), .A2(
        \SB3_2/i0_3 ), .A3(\SB3_2/i0_4 ), .ZN(
        \SB3_2/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_3/Component_Function_2/N1  ( .A1(\SB3_3/i1_5 ), .A2(
        \SB3_3/i0[10] ), .A3(\SB3_3/i1[9] ), .ZN(
        \SB3_3/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_3/Component_Function_4/N4  ( .A1(\SB3_3/i1[9] ), .A2(
        \SB3_3/i1_5 ), .A3(\SB3_3/i0_4 ), .ZN(
        \SB3_3/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_3/Component_Function_4/N2  ( .A1(\SB3_3/i3[0] ), .A2(
        \SB3_3/i0_0 ), .A3(\SB3_3/i1_7 ), .ZN(
        \SB3_3/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_3/Component_Function_4/N1  ( .A1(\SB3_3/i0[9] ), .A2(
        \SB3_3/i0_0 ), .A3(\SB3_3/i0[8] ), .ZN(
        \SB3_3/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_4/Component_Function_2/N1  ( .A1(n2910), .A2(\SB3_4/i0[10] ), 
        .A3(\SB3_4/i1[9] ), .ZN(\SB3_4/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_4/Component_Function_4/N2  ( .A1(\SB3_4/i3[0] ), .A2(
        \SB3_4/i0_0 ), .A3(\SB3_4/i1_7 ), .ZN(
        \SB3_4/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_4/Component_Function_4/N1  ( .A1(\SB3_4/i0[9] ), .A2(
        \SB3_4/i0_0 ), .A3(\SB3_4/i0[8] ), .ZN(
        \SB3_4/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_5/Component_Function_4/N4  ( .A1(\SB3_5/i1[9] ), .A2(
        \SB3_5/i1_5 ), .A3(\SB3_5/i0_4 ), .ZN(
        \SB3_5/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_6/Component_Function_2/N2  ( .A1(\RI1[4][155] ), .A2(
        \SB3_6/i0[10] ), .A3(\SB3_6/i0[6] ), .ZN(
        \SB3_6/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_6/Component_Function_4/N1  ( .A1(\SB3_6/i0[9] ), .A2(
        \SB3_6/i0_0 ), .A3(\SB3_6/i0[8] ), .ZN(
        \SB3_6/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_7/Component_Function_2/N2  ( .A1(\SB3_7/i0_3 ), .A2(
        \SB3_7/i0[10] ), .A3(\SB3_7/i0[6] ), .ZN(
        \SB3_7/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_7/Component_Function_4/N2  ( .A1(\SB3_7/i3[0] ), .A2(
        \SB3_7/i0_0 ), .A3(\SB3_7/i1_7 ), .ZN(
        \SB3_7/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_7/Component_Function_4/N1  ( .A1(\SB3_7/i0[9] ), .A2(
        \SB3_7/i0_0 ), .A3(\SB3_7/i0[8] ), .ZN(
        \SB3_7/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_8/Component_Function_2/N1  ( .A1(\SB3_8/i1_5 ), .A2(
        \SB3_8/i0[10] ), .A3(\SB3_8/i1[9] ), .ZN(
        \SB3_8/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_8/Component_Function_4/N1  ( .A1(\SB3_8/i0[9] ), .A2(
        \SB3_8/i0_0 ), .A3(\SB3_8/i0[8] ), .ZN(
        \SB3_8/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_9/Component_Function_3/N2  ( .A1(\SB3_9/i0_0 ), .A2(
        \SB3_9/i0_3 ), .A3(\SB3_9/i0_4 ), .ZN(
        \SB3_9/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_9/Component_Function_4/N2  ( .A1(\SB3_9/i3[0] ), .A2(
        \SB3_9/i0_0 ), .A3(\SB3_9/i1_7 ), .ZN(
        \SB3_9/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_9/Component_Function_4/N1  ( .A1(\SB3_9/i0[9] ), .A2(
        \SB3_9/i0_0 ), .A3(\SB3_9/i0[8] ), .ZN(
        \SB3_9/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_10/Component_Function_2/N1  ( .A1(\SB3_10/i1_5 ), .A2(
        \SB3_10/i0[10] ), .A3(\SB3_10/i1[9] ), .ZN(
        \SB3_10/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_10/Component_Function_4/N1  ( .A1(\SB3_10/i0[9] ), .A2(
        \SB3_10/i0_0 ), .A3(\SB3_10/i0[8] ), .ZN(
        \SB3_10/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_11/Component_Function_3/N4  ( .A1(n582), .A2(\SB3_11/i0[8] ), 
        .A3(\SB3_11/i3[0] ), .ZN(\SB3_11/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB3_11/Component_Function_3/N2  ( .A1(\SB3_11/i0_0 ), .A2(
        \SB3_11/i0_3 ), .A3(\SB3_11/i0_4 ), .ZN(
        \SB3_11/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_12/Component_Function_4/N1  ( .A1(\SB3_12/i0[9] ), .A2(
        \SB3_12/i0_0 ), .A3(\SB3_12/i0[8] ), .ZN(
        \SB3_12/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_13/Component_Function_4/N3  ( .A1(\SB3_13/i0[9] ), .A2(
        \SB3_13/i0[10] ), .A3(\SB3_13/i0_3 ), .ZN(
        \SB3_13/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB3_13/Component_Function_4/N2  ( .A1(\SB3_13/i3[0] ), .A2(
        \MC_ARK_ARC_1_3/buf_output[110] ), .A3(\SB3_13/i1_7 ), .ZN(
        \SB3_13/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_14/Component_Function_3/N1  ( .A1(\SB3_14/i1[9] ), .A2(
        \SB3_14/i0_3 ), .A3(\SB3_14/i0[6] ), .ZN(
        \SB3_14/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_14/Component_Function_4/N4  ( .A1(\SB3_14/i1[9] ), .A2(
        \SB3_14/i1_5 ), .A3(\SB3_14/i0_4 ), .ZN(
        \SB3_14/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_14/Component_Function_4/N2  ( .A1(\SB3_14/i3[0] ), .A2(
        \SB3_14/i0_0 ), .A3(\SB3_14/i1_7 ), .ZN(
        \SB3_14/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_15/Component_Function_3/N2  ( .A1(\SB3_15/i0_0 ), .A2(
        \SB3_15/i0_3 ), .A3(\SB3_15/i0_4 ), .ZN(
        \SB3_15/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_15/Component_Function_4/N2  ( .A1(\SB3_15/i3[0] ), .A2(
        \SB3_15/i0_0 ), .A3(\SB3_15/i1_7 ), .ZN(
        \SB3_15/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_15/Component_Function_4/N1  ( .A1(\SB3_15/i0[9] ), .A2(
        \SB3_15/i0_0 ), .A3(\SB3_15/i0[8] ), .ZN(
        \SB3_15/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_16/Component_Function_3/N1  ( .A1(\SB3_16/i1[9] ), .A2(
        \SB3_16/i0_3 ), .A3(\SB3_16/i0[6] ), .ZN(
        \SB3_16/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_16/Component_Function_4/N3  ( .A1(\SB3_16/i0[9] ), .A2(
        \SB3_16/i0[10] ), .A3(\SB3_16/i0_3 ), .ZN(
        \SB3_16/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB3_16/Component_Function_4/N2  ( .A1(\SB3_16/i3[0] ), .A2(
        \SB3_16/i0_0 ), .A3(\SB3_16/i1_7 ), .ZN(
        \SB3_16/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_16/Component_Function_4/N1  ( .A1(\SB3_16/i0[9] ), .A2(
        \SB3_16/i0_0 ), .A3(\SB3_16/i0[8] ), .ZN(
        \SB3_16/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_17/Component_Function_4/N2  ( .A1(\SB3_17/i3[0] ), .A2(
        \SB3_17/i0_0 ), .A3(\SB3_17/i1_7 ), .ZN(
        \SB3_17/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_18/Component_Function_4/N1  ( .A1(\SB3_18/i0[9] ), .A2(
        \SB3_18/i0_0 ), .A3(\SB3_18/i0[8] ), .ZN(
        \SB3_18/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_19/Component_Function_2/N1  ( .A1(\SB3_19/i1_5 ), .A2(
        \SB3_19/i0[10] ), .A3(\SB3_19/i1[9] ), .ZN(
        \SB3_19/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_19/Component_Function_4/N2  ( .A1(\SB3_19/i3[0] ), .A2(
        \SB3_19/i0_0 ), .A3(\SB3_19/i1_7 ), .ZN(
        \SB3_19/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_19/Component_Function_4/N1  ( .A1(\SB3_19/i0[9] ), .A2(
        \SB3_19/i0_0 ), .A3(\SB3_19/i0[8] ), .ZN(
        \SB3_19/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_20/Component_Function_2/N1  ( .A1(\SB3_20/i1_5 ), .A2(
        \SB3_20/i0[10] ), .A3(\SB3_20/i1[9] ), .ZN(
        \SB3_20/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_20/Component_Function_3/N2  ( .A1(\SB3_20/i0_0 ), .A2(
        \SB3_20/i0_3 ), .A3(\SB3_20/i0_4 ), .ZN(
        \SB3_20/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_20/Component_Function_4/N2  ( .A1(\SB3_20/i3[0] ), .A2(
        \SB3_20/i0_0 ), .A3(\SB3_20/i1_7 ), .ZN(
        \SB3_20/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_21/Component_Function_4/N4  ( .A1(\SB3_21/i1[9] ), .A2(
        \SB3_21/i1_5 ), .A3(\SB3_21/i0_4 ), .ZN(
        \SB3_21/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_22/Component_Function_4/N2  ( .A1(\SB3_22/i3[0] ), .A2(
        \SB3_22/i0_0 ), .A3(\SB3_22/i1_7 ), .ZN(
        \SB3_22/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_22/Component_Function_4/N1  ( .A1(\SB3_22/i0[9] ), .A2(
        \SB3_22/i0_0 ), .A3(\SB3_22/i0[8] ), .ZN(
        \SB3_22/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_23/Component_Function_4/N1  ( .A1(\SB3_23/i0[9] ), .A2(
        \SB3_23/i0_0 ), .A3(\SB3_23/i0[8] ), .ZN(
        \SB3_23/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_24/Component_Function_4/N3  ( .A1(\SB3_24/i0[9] ), .A2(
        \SB3_24/i0[10] ), .A3(\SB3_24/i0_3 ), .ZN(
        \SB3_24/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB3_25/Component_Function_2/N3  ( .A1(\SB3_25/i0_3 ), .A2(
        \SB3_25/i0[8] ), .A3(\MC_ARK_ARC_1_3/buf_output[36] ), .ZN(
        \SB3_25/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_25/Component_Function_4/N2  ( .A1(\SB3_25/i3[0] ), .A2(
        \SB3_25/i0_0 ), .A3(\SB3_25/i1_7 ), .ZN(
        \SB3_25/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_25/Component_Function_4/N1  ( .A1(\SB3_25/i0[9] ), .A2(
        \SB3_25/i0_0 ), .A3(\SB3_25/i0[8] ), .ZN(
        \SB3_25/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_26/Component_Function_2/N3  ( .A1(\SB3_26/i0_3 ), .A2(
        \SB3_26/i0[8] ), .A3(\MC_ARK_ARC_1_3/buf_output[30] ), .ZN(
        \SB3_26/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_26/Component_Function_4/N2  ( .A1(\SB3_26/i3[0] ), .A2(
        \SB3_26/i0_0 ), .A3(\SB3_26/i1_7 ), .ZN(
        \SB3_26/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_26/Component_Function_4/N1  ( .A1(\SB3_26/i0[9] ), .A2(
        \SB3_26/i0_0 ), .A3(\SB3_26/i0[8] ), .ZN(
        \SB3_26/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_27/Component_Function_3/N2  ( .A1(\SB3_27/i0_0 ), .A2(
        \SB3_27/i0_3 ), .A3(\SB3_27/i0_4 ), .ZN(
        \SB3_27/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_27/Component_Function_4/N1  ( .A1(\SB3_27/i0[9] ), .A2(
        \SB3_27/i0_0 ), .A3(\SB3_27/i0[8] ), .ZN(
        \SB3_27/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_28/Component_Function_2/N1  ( .A1(\SB3_28/i1_5 ), .A2(
        \SB3_28/i0[10] ), .A3(\SB3_28/i1[9] ), .ZN(
        \SB3_28/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_28/Component_Function_3/N3  ( .A1(\SB3_28/i1[9] ), .A2(
        \SB3_28/i1_7 ), .A3(\SB3_28/i0[10] ), .ZN(
        \SB3_28/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB3_28/Component_Function_4/N2  ( .A1(\SB3_28/i3[0] ), .A2(
        \SB3_28/i0_0 ), .A3(\SB3_28/i1_7 ), .ZN(
        \SB3_28/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_28/Component_Function_4/N1  ( .A1(\SB3_28/i0[9] ), .A2(
        \SB3_28/i0_0 ), .A3(\SB3_28/i0[8] ), .ZN(
        \SB3_28/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_29/Component_Function_3/N4  ( .A1(\SB3_29/i1_5 ), .A2(
        \SB3_29/i0[8] ), .A3(\SB3_29/i3[0] ), .ZN(
        \SB3_29/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB3_29/Component_Function_3/N2  ( .A1(\SB3_29/i0_0 ), .A2(
        \SB3_29/i0_3 ), .A3(\SB3_29/i0_4 ), .ZN(
        \SB3_29/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_29/Component_Function_4/N2  ( .A1(\SB3_29/i3[0] ), .A2(
        \SB3_29/i0_0 ), .A3(\SB3_29/i1_7 ), .ZN(
        \SB3_29/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB3_29/Component_Function_4/N1  ( .A1(\SB3_29/i0[9] ), .A2(
        \SB3_29/i0_0 ), .A3(\SB3_29/i0[8] ), .ZN(
        \SB3_29/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB3_30/Component_Function_2/N3  ( .A1(n5509), .A2(\SB3_30/i0[8] ), 
        .A3(\SB3_30/i0[9] ), .ZN(\SB3_30/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_30/Component_Function_2/N1  ( .A1(\SB3_30/i1_5 ), .A2(
        \SB3_30/i0[10] ), .A3(\SB3_30/i1[9] ), .ZN(
        \SB3_30/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_31/Component_Function_2/N1  ( .A1(\SB3_31/i1_5 ), .A2(
        \SB3_31/i0[10] ), .A3(\SB3_31/i1[9] ), .ZN(
        \SB3_31/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_31/Component_Function_3/N2  ( .A1(\SB3_31/i0_0 ), .A2(
        \SB3_31/i0_3 ), .A3(\SB3_31/i0_4 ), .ZN(
        \SB3_31/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB3_31/Component_Function_4/N4  ( .A1(\SB3_31/i1[9] ), .A2(
        \SB3_31/i1_5 ), .A3(\SB3_31/i0_4 ), .ZN(
        \SB3_31/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB4_0/Component_Function_3/N4  ( .A1(\SB4_0/i1_5 ), .A2(
        \SB4_0/i0[8] ), .A3(\SB4_0/i3[0] ), .ZN(
        \SB4_0/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_2/Component_Function_2/N3  ( .A1(\SB4_2/i0_3 ), .A2(
        \SB4_2/i0[8] ), .A3(\SB4_2/i0[9] ), .ZN(
        \SB4_2/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_3/Component_Function_2/N1  ( .A1(\SB4_3/i1_5 ), .A2(
        \SB3_5/buf_output[3] ), .A3(n1371), .ZN(
        \SB4_3/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB4_3/Component_Function_4/N2  ( .A1(\SB4_3/i3[0] ), .A2(
        \SB3_6/buf_output[2] ), .A3(\SB4_3/i1_7 ), .ZN(
        \SB4_3/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB4_4/Component_Function_3/N4  ( .A1(\SB4_4/i1_5 ), .A2(
        \SB4_4/i0[8] ), .A3(\SB4_4/i3[0] ), .ZN(
        \SB4_4/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_4/Component_Function_4/N1  ( .A1(\SB4_4/i0[9] ), .A2(
        \SB3_7/buf_output[2] ), .A3(\SB4_4/i0[8] ), .ZN(
        \SB4_4/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_5/Component_Function_3/N4  ( .A1(\SB4_5/i1_5 ), .A2(
        \SB4_5/i0[8] ), .A3(\SB4_5/i3[0] ), .ZN(
        \SB4_5/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_6/Component_Function_2/N4  ( .A1(\SB4_6/i1_5 ), .A2(
        \SB4_6/i0_0 ), .A3(\SB4_6/i0_4 ), .ZN(
        \SB4_6/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB4_6/Component_Function_3/N4  ( .A1(\SB4_6/i1_5 ), .A2(n579), 
        .A3(\SB4_6/i3[0] ), .ZN(\SB4_6/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_6/Component_Function_4/N4  ( .A1(\SB4_6/i1[9] ), .A2(
        \SB4_6/i1_5 ), .A3(\SB4_6/i0_4 ), .ZN(
        \SB4_6/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB4_7/Component_Function_2/N1  ( .A1(\SB4_7/i1_5 ), .A2(
        \SB4_7/i0[10] ), .A3(\SB4_7/i1[9] ), .ZN(
        \SB4_7/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB4_7/Component_Function_3/N4  ( .A1(\SB4_7/i1_5 ), .A2(
        \SB4_7/i0[8] ), .A3(\SB4_7/i3[0] ), .ZN(
        \SB4_7/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_7/Component_Function_3/N2  ( .A1(\SB4_7/i0_0 ), .A2(
        \SB4_7/i0_3 ), .A3(\SB4_7/i0_4 ), .ZN(
        \SB4_7/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB4_8/Component_Function_2/N3  ( .A1(\SB4_8/i0_3 ), .A2(
        \SB4_8/i0[8] ), .A3(\SB4_8/i0[9] ), .ZN(
        \SB4_8/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_8/Component_Function_3/N4  ( .A1(\SB4_8/i1_5 ), .A2(
        \SB4_8/i0[8] ), .A3(\SB4_8/i3[0] ), .ZN(
        \SB4_8/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_9/Component_Function_4/N4  ( .A1(\SB4_9/i1[9] ), .A2(
        \SB4_9/i1_5 ), .A3(\SB4_9/i0_4 ), .ZN(
        \SB4_9/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB4_10/Component_Function_2/N1  ( .A1(\SB4_10/i1_5 ), .A2(
        \SB4_10/i0[10] ), .A3(n3653), .ZN(
        \SB4_10/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB4_10/Component_Function_3/N4  ( .A1(\SB4_10/i1_5 ), .A2(
        \SB4_10/i0[8] ), .A3(\SB4_10/i3[0] ), .ZN(
        \SB4_10/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_11/Component_Function_2/N3  ( .A1(\SB4_11/i0_3 ), .A2(
        \SB4_11/i0[8] ), .A3(\SB4_11/i0[9] ), .ZN(
        \SB4_11/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_11/Component_Function_3/N4  ( .A1(n3684), .A2(\SB4_11/i0[8] ), 
        .A3(\SB4_11/i3[0] ), .ZN(\SB4_11/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_11/Component_Function_3/N2  ( .A1(\SB4_11/i0_0 ), .A2(
        \SB4_11/i0_3 ), .A3(\SB4_11/i0_4 ), .ZN(
        \SB4_11/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB4_11/Component_Function_4/N4  ( .A1(\SB4_11/i1[9] ), .A2(n3684), 
        .A3(\SB4_11/i0_4 ), .ZN(\SB4_11/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB4_12/Component_Function_2/N1  ( .A1(\SB4_12/i1_5 ), .A2(
        \SB4_12/i0[10] ), .A3(\SB4_12/i1[9] ), .ZN(
        \SB4_12/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB4_12/Component_Function_3/N4  ( .A1(\SB4_12/i1_5 ), .A2(
        \SB4_12/i0[8] ), .A3(\SB4_12/i3[0] ), .ZN(
        \SB4_12/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_13/Component_Function_2/N2  ( .A1(\SB4_13/i0_3 ), .A2(
        \SB4_13/i0[10] ), .A3(\SB4_13/i0[6] ), .ZN(
        \SB4_13/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_14/Component_Function_2/N3  ( .A1(\SB4_14/i0_3 ), .A2(
        \SB4_14/i0[8] ), .A3(\SB4_14/i0[9] ), .ZN(
        \SB4_14/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_14/Component_Function_3/N4  ( .A1(\SB4_14/i1_5 ), .A2(
        \SB4_14/i0[8] ), .A3(\SB4_14/i3[0] ), .ZN(
        \SB4_14/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_15/Component_Function_3/N4  ( .A1(\SB4_15/i1_5 ), .A2(
        \SB4_15/i0[8] ), .A3(\SB4_15/i3[0] ), .ZN(
        \SB4_15/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_15/Component_Function_4/N4  ( .A1(\SB4_15/i1[9] ), .A2(
        \SB4_15/i1_5 ), .A3(\SB4_15/i0_4 ), .ZN(
        \SB4_15/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB4_18/Component_Function_2/N3  ( .A1(\SB4_18/i0_3 ), .A2(n3662), 
        .A3(\SB4_18/i0[9] ), .ZN(\SB4_18/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_18/Component_Function_4/N4  ( .A1(\SB4_18/i1[9] ), .A2(
        \SB4_18/i1_5 ), .A3(\SB4_18/i0_4 ), .ZN(
        \SB4_18/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB4_19/Component_Function_2/N3  ( .A1(\SB4_19/i0_3 ), .A2(n3668), 
        .A3(\SB4_19/i0[9] ), .ZN(\SB4_19/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_19/Component_Function_3/N4  ( .A1(\SB4_19/i1_5 ), .A2(n3668), 
        .A3(\SB4_19/i3[0] ), .ZN(\SB4_19/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_19/Component_Function_3/N2  ( .A1(\SB4_19/i0_0 ), .A2(
        \SB4_19/i0_3 ), .A3(\SB4_19/i0_4 ), .ZN(
        \SB4_19/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB4_19/Component_Function_4/N4  ( .A1(\SB4_19/i1[9] ), .A2(
        \SB4_19/i1_5 ), .A3(n5486), .ZN(
        \SB4_19/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB4_19/Component_Function_4/N1  ( .A1(\SB4_19/i0[9] ), .A2(
        \SB4_19/i0_0 ), .A3(n3668), .ZN(
        \SB4_19/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_21/Component_Function_2/N3  ( .A1(\SB4_21/i0_3 ), .A2(
        \SB4_21/i0[8] ), .A3(\SB4_21/i0[9] ), .ZN(
        \SB4_21/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_21/Component_Function_3/N4  ( .A1(\SB4_21/i1_5 ), .A2(
        \SB4_21/i0[8] ), .A3(\SB4_21/i3[0] ), .ZN(
        \SB4_21/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_21/Component_Function_4/N4  ( .A1(n3666), .A2(\SB4_21/i1_5 ), 
        .A3(\SB4_21/i0_4 ), .ZN(\SB4_21/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB4_22/Component_Function_4/N4  ( .A1(\SB4_22/i1[9] ), .A2(
        \SB4_22/i1_5 ), .A3(\SB4_22/i0_4 ), .ZN(
        \SB4_22/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB4_23/Component_Function_2/N3  ( .A1(\SB4_23/i0_3 ), .A2(
        \SB4_23/i0[8] ), .A3(\SB4_23/i0[9] ), .ZN(
        \SB4_23/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_23/Component_Function_3/N4  ( .A1(\SB4_23/i1_5 ), .A2(
        \SB4_23/i0[8] ), .A3(\SB4_23/i3[0] ), .ZN(
        \SB4_23/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_24/Component_Function_2/N3  ( .A1(\SB4_24/i0_3 ), .A2(
        \SB4_24/i0[8] ), .A3(\SB4_24/i0[9] ), .ZN(
        \SB4_24/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_24/Component_Function_2/N2  ( .A1(\SB4_24/i0_3 ), .A2(
        \SB4_24/i0[10] ), .A3(\SB4_24/i0[6] ), .ZN(
        \SB4_24/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_24/Component_Function_3/N4  ( .A1(\SB4_24/i1_5 ), .A2(
        \SB4_24/i0[8] ), .A3(\SB4_24/i3[0] ), .ZN(
        \SB4_24/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_24/Component_Function_4/N1  ( .A1(\SB4_24/i0[9] ), .A2(
        \SB4_24/i0_0 ), .A3(\SB4_24/i0[8] ), .ZN(
        \SB4_24/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_25/Component_Function_2/N2  ( .A1(\SB4_25/i0_3 ), .A2(
        \SB4_25/i0[10] ), .A3(\SB4_25/i0[6] ), .ZN(
        \SB4_25/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB4_25/Component_Function_3/N4  ( .A1(\SB4_25/i1_5 ), .A2(
        \SB4_25/i0[8] ), .A3(\SB4_25/i3[0] ), .ZN(
        \SB4_25/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_25/Component_Function_3/N2  ( .A1(\SB4_25/i0_0 ), .A2(
        \SB4_25/i0_3 ), .A3(\SB4_25/i0_4 ), .ZN(
        \SB4_25/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB4_25/Component_Function_4/N4  ( .A1(\SB4_25/i1[9] ), .A2(
        \SB4_25/i1_5 ), .A3(\SB4_25/i0_4 ), .ZN(
        \SB4_25/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB4_25/Component_Function_4/N1  ( .A1(\SB4_25/i0[9] ), .A2(
        \SB4_25/i0_0 ), .A3(\SB4_25/i0[8] ), .ZN(
        \SB4_25/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB4_26/Component_Function_2/N1  ( .A1(\SB4_26/i1_5 ), .A2(
        \SB4_26/i0[10] ), .A3(\SB4_26/i1[9] ), .ZN(
        \SB4_26/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB4_26/Component_Function_3/N4  ( .A1(\SB4_26/i1_5 ), .A2(
        \SB4_26/i0[8] ), .A3(\SB4_26/i3[0] ), .ZN(
        \SB4_26/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_26/Component_Function_3/N2  ( .A1(\SB4_26/i0_0 ), .A2(
        \SB4_26/i0_3 ), .A3(\SB4_26/i0_4 ), .ZN(
        \SB4_26/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB4_26/Component_Function_4/N2  ( .A1(\SB4_26/i3[0] ), .A2(
        \SB4_26/i0_0 ), .A3(\SB4_26/i1_7 ), .ZN(
        \SB4_26/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB4_27/Component_Function_2/N1  ( .A1(\SB4_27/i1_5 ), .A2(
        \SB4_27/i0[10] ), .A3(n1389), .ZN(
        \SB4_27/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB4_27/Component_Function_3/N1  ( .A1(n1389), .A2(\SB4_27/i0_3 ), 
        .A3(\SB4_27/i0[6] ), .ZN(\SB4_27/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB4_27/Component_Function_4/N2  ( .A1(\SB4_27/i3[0] ), .A2(n2897), 
        .A3(\SB4_27/i1_7 ), .ZN(\SB4_27/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB4_28/Component_Function_3/N3  ( .A1(n5514), .A2(\SB4_28/i1_7 ), 
        .A3(\SB4_28/i0[10] ), .ZN(\SB4_28/Component_Function_3/NAND4_in[2] )
         );
  NAND3_X1 \SB4_29/Component_Function_2/N4  ( .A1(\SB4_29/i1_5 ), .A2(
        \SB4_29/i0_0 ), .A3(n1793), .ZN(
        \SB4_29/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB4_29/Component_Function_3/N4  ( .A1(\SB4_29/i1_5 ), .A2(
        \SB4_29/i0[8] ), .A3(\SB4_29/i3[0] ), .ZN(
        \SB4_29/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_30/Component_Function_3/N4  ( .A1(n5525), .A2(\SB4_30/i0[8] ), 
        .A3(\SB4_30/i3[0] ), .ZN(\SB4_30/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB4_31/Component_Function_3/N4  ( .A1(\SB4_31/i1_5 ), .A2(n3652), 
        .A3(\SB4_31/i3[0] ), .ZN(\SB4_31/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_0/Component_Function_0/N3  ( .A1(\SB1_0_0/i0[10] ), .A2(
        \SB1_0_0/i0_4 ), .A3(\SB1_0_0/i0_3 ), .ZN(
        \SB1_0_0/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_0/Component_Function_0/N2  ( .A1(\SB1_0_0/i0[8] ), .A2(
        \SB1_0_0/i0[7] ), .A3(n6028), .ZN(
        \SB1_0_0/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_0/Component_Function_1/N3  ( .A1(\SB1_0_0/i1_5 ), .A2(n1376), 
        .A3(\SB1_0_0/i0[9] ), .ZN(\SB1_0_0/Component_Function_1/NAND4_in[2] )
         );
  NAND2_X1 \SB1_0_0/Component_Function_5/N1  ( .A1(\SB1_0_0/i0_0 ), .A2(
        \SB1_0_0/i3[0] ), .ZN(\SB1_0_0/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_1/Component_Function_0/N2  ( .A1(\SB1_0_1/i0[8] ), .A2(
        \SB1_0_1/i0[7] ), .A3(\SB1_0_1/i0[6] ), .ZN(
        \SB1_0_1/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_1/Component_Function_0/N1  ( .A1(\SB1_0_1/i0[10] ), .A2(
        \SB1_0_1/i0[9] ), .ZN(\SB1_0_1/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_1/Component_Function_1/N3  ( .A1(\SB1_0_1/i1_5 ), .A2(
        \SB1_0_1/i0[6] ), .A3(\SB1_0_1/i0[9] ), .ZN(
        \SB1_0_1/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB1_0_1/Component_Function_1/N1  ( .A1(\SB1_0_1/i0_3 ), .A2(
        \SB1_0_1/i1[9] ), .ZN(\SB1_0_1/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_1/Component_Function_5/N3  ( .A1(\SB1_0_1/i1[9] ), .A2(
        \SB1_0_1/i0_4 ), .A3(\SB1_0_1/i0_3 ), .ZN(
        \SB1_0_1/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_2/Component_Function_0/N2  ( .A1(\SB1_0_2/i0[8] ), .A2(
        \SB1_0_2/i0[7] ), .A3(\SB1_0_2/i0[6] ), .ZN(
        \SB1_0_2/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_2/Component_Function_1/N3  ( .A1(\SB1_0_2/i1_5 ), .A2(
        \SB1_0_2/i0[6] ), .A3(\SB1_0_2/i0[9] ), .ZN(
        \SB1_0_2/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_2/Component_Function_1/N2  ( .A1(\SB1_0_2/i0_3 ), .A2(
        \SB1_0_2/i1_7 ), .A3(\SB1_0_2/i0[8] ), .ZN(
        \SB1_0_2/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_3/Component_Function_0/N2  ( .A1(\SB1_0_3/i0[8] ), .A2(
        \SB1_0_3/i0[7] ), .A3(\SB1_0_3/i0[6] ), .ZN(
        \SB1_0_3/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_3/Component_Function_0/N1  ( .A1(\SB1_0_3/i0[10] ), .A2(
        \SB1_0_3/i0[9] ), .ZN(\SB1_0_3/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_3/Component_Function_1/N3  ( .A1(\SB1_0_3/i1_5 ), .A2(
        \SB1_0_3/i0[6] ), .A3(\SB1_0_3/i0[9] ), .ZN(
        \SB1_0_3/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB1_0_3/Component_Function_1/N1  ( .A1(\SB1_0_3/i0_3 ), .A2(
        \SB1_0_3/i1[9] ), .ZN(\SB1_0_3/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_4/Component_Function_0/N3  ( .A1(\SB1_0_4/i0[10] ), .A2(
        \SB1_0_4/i0_4 ), .A3(\SB1_0_4/i0_3 ), .ZN(
        \SB1_0_4/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_4/Component_Function_0/N2  ( .A1(\SB1_0_4/i0[8] ), .A2(
        \SB1_0_4/i0[7] ), .A3(\SB1_0_4/i0[6] ), .ZN(
        \SB1_0_4/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_4/Component_Function_0/N1  ( .A1(\SB1_0_4/i0[10] ), .A2(
        \SB1_0_4/i0[9] ), .ZN(\SB1_0_4/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_4/Component_Function_1/N4  ( .A1(\SB1_0_4/i1_7 ), .A2(
        \SB1_0_4/i0[8] ), .A3(n396), .ZN(
        \SB1_0_4/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_4/Component_Function_1/N3  ( .A1(\SB1_0_4/i1_5 ), .A2(
        \SB1_0_4/i0[6] ), .A3(\SB1_0_4/i0[9] ), .ZN(
        \SB1_0_4/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_4/Component_Function_1/N2  ( .A1(\SB1_0_4/i0_3 ), .A2(
        \SB1_0_4/i1_7 ), .A3(\SB1_0_4/i0[8] ), .ZN(
        \SB1_0_4/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_4/Component_Function_1/N1  ( .A1(\SB1_0_4/i0_3 ), .A2(
        \SB1_0_4/i1[9] ), .ZN(\SB1_0_4/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_5/Component_Function_0/N3  ( .A1(\SB1_0_5/i0[10] ), .A2(
        \SB1_0_5/i0_4 ), .A3(\SB1_0_5/i0_3 ), .ZN(
        \SB1_0_5/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_0_5/Component_Function_0/N1  ( .A1(\SB1_0_5/i0[10] ), .A2(
        \SB1_0_5/i0[9] ), .ZN(\SB1_0_5/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_5/Component_Function_1/N3  ( .A1(\SB1_0_5/i1_5 ), .A2(
        \SB1_0_5/i0[6] ), .A3(\SB1_0_5/i0[9] ), .ZN(
        \SB1_0_5/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_5/Component_Function_1/N2  ( .A1(\SB1_0_5/i0_3 ), .A2(
        \SB1_0_5/i1_7 ), .A3(\SB1_0_5/i0[8] ), .ZN(
        \SB1_0_5/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_6/Component_Function_0/N4  ( .A1(\SB1_0_6/i0[7] ), .A2(
        \SB1_0_6/i0_3 ), .A3(\SB1_0_6/i0_0 ), .ZN(
        \SB1_0_6/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_6/Component_Function_0/N2  ( .A1(\SB1_0_6/i0[8] ), .A2(
        \SB1_0_6/i0[7] ), .A3(\SB1_0_6/i0[6] ), .ZN(
        \SB1_0_6/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_6/Component_Function_0/N1  ( .A1(\SB1_0_6/i0[10] ), .A2(
        \SB1_0_6/i0[9] ), .ZN(\SB1_0_6/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_6/Component_Function_1/N4  ( .A1(\SB1_0_6/i1_7 ), .A2(
        \SB1_0_6/i0[8] ), .A3(\SB1_0_6/i0_4 ), .ZN(
        \SB1_0_6/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_6/Component_Function_5/N4  ( .A1(n320), .A2(n321), .A3(n392), 
        .ZN(\SB1_0_6/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_7/Component_Function_0/N2  ( .A1(\SB1_0_7/i0[8] ), .A2(
        \SB1_0_7/i0[7] ), .A3(\SB1_0_7/i0[6] ), .ZN(
        \SB1_0_7/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_7/Component_Function_0/N1  ( .A1(\SB1_0_7/i0[10] ), .A2(
        \SB1_0_7/i0[9] ), .ZN(\SB1_0_7/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_7/Component_Function_1/N3  ( .A1(\SB1_0_7/i1_5 ), .A2(
        \SB1_0_7/i0[6] ), .A3(\SB1_0_7/i0[9] ), .ZN(
        \SB1_0_7/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_7/Component_Function_5/N4  ( .A1(\SB1_0_7/i0[9] ), .A2(
        \SB1_0_7/i0[6] ), .A3(n5496), .ZN(
        \SB1_0_7/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_8/Component_Function_0/N2  ( .A1(\SB1_0_8/i0[8] ), .A2(
        \SB1_0_8/i0[7] ), .A3(\SB1_0_8/i0[6] ), .ZN(
        \SB1_0_8/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_8/Component_Function_0/N1  ( .A1(\SB1_0_8/i0[10] ), .A2(
        \SB1_0_8/i0[9] ), .ZN(\SB1_0_8/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_8/Component_Function_1/N4  ( .A1(\SB1_0_8/i1_7 ), .A2(
        \SB1_0_8/i0[8] ), .A3(\SB1_0_8/i0_4 ), .ZN(
        \SB1_0_8/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_8/Component_Function_1/N3  ( .A1(\SB1_0_8/i1_5 ), .A2(
        \SB1_0_8/i0[6] ), .A3(\SB1_0_8/i0[9] ), .ZN(
        \SB1_0_8/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB1_0_8/Component_Function_5/N1  ( .A1(\SB1_0_8/i0_0 ), .A2(
        \SB1_0_8/i3[0] ), .ZN(\SB1_0_8/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_9/Component_Function_0/N4  ( .A1(\SB1_0_9/i0[7] ), .A2(
        \SB1_0_9/i0_3 ), .A3(\SB1_0_9/i0_0 ), .ZN(
        \SB1_0_9/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_9/Component_Function_0/N3  ( .A1(\SB1_0_9/i0[10] ), .A2(
        \SB1_0_9/i0_4 ), .A3(\SB1_0_9/i0_3 ), .ZN(
        \SB1_0_9/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_9/Component_Function_0/N2  ( .A1(\SB1_0_9/i0[8] ), .A2(
        \SB1_0_9/i0[7] ), .A3(\SB1_0_9/i0[6] ), .ZN(
        \SB1_0_9/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_9/Component_Function_0/N1  ( .A1(\SB1_0_9/i0[10] ), .A2(
        \SB1_0_9/i0[9] ), .ZN(\SB1_0_9/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_9/Component_Function_1/N4  ( .A1(\SB1_0_9/i1_7 ), .A2(
        \SB1_0_9/i0[8] ), .A3(\SB1_0_9/i0_4 ), .ZN(
        \SB1_0_9/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_9/Component_Function_1/N2  ( .A1(\SB1_0_9/i0_3 ), .A2(
        \SB1_0_9/i1_7 ), .A3(\SB1_0_9/i0[8] ), .ZN(
        \SB1_0_9/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_9/Component_Function_1/N1  ( .A1(\SB1_0_9/i0_3 ), .A2(
        \SB1_0_9/i1[9] ), .ZN(\SB1_0_9/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_10/Component_Function_0/N3  ( .A1(\SB1_0_10/i0[10] ), .A2(
        \SB1_0_10/i0_4 ), .A3(\SB1_0_10/i0_3 ), .ZN(
        \SB1_0_10/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_10/Component_Function_0/N2  ( .A1(\SB1_0_10/i0[8] ), .A2(
        \SB1_0_10/i0[7] ), .A3(\SB1_0_10/i0[6] ), .ZN(
        \SB1_0_10/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_10/Component_Function_0/N1  ( .A1(\SB1_0_10/i0[10] ), .A2(
        \SB1_0_10/i0[9] ), .ZN(\SB1_0_10/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_10/Component_Function_1/N4  ( .A1(\SB1_0_10/i1_7 ), .A2(
        \SB1_0_10/i0[8] ), .A3(\SB1_0_10/i0_4 ), .ZN(
        \SB1_0_10/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_10/Component_Function_1/N3  ( .A1(\SB1_0_10/i1_5 ), .A2(
        \SB1_0_10/i0[6] ), .A3(\SB1_0_10/i0[9] ), .ZN(
        \SB1_0_10/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_10/Component_Function_1/N2  ( .A1(\SB1_0_10/i0_3 ), .A2(
        \SB1_0_10/i1_7 ), .A3(\SB1_0_10/i0[8] ), .ZN(
        \SB1_0_10/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_10/Component_Function_1/N1  ( .A1(\SB1_0_10/i0_3 ), .A2(
        \SB1_0_10/i1[9] ), .ZN(\SB1_0_10/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_11/Component_Function_0/N3  ( .A1(\SB1_0_11/i0[10] ), .A2(
        \SB1_0_11/i0_4 ), .A3(\SB1_0_11/i0_3 ), .ZN(
        \SB1_0_11/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_11/Component_Function_0/N2  ( .A1(\SB1_0_11/i0[8] ), .A2(
        \SB1_0_11/i0[7] ), .A3(\SB1_0_11/i0[6] ), .ZN(
        \SB1_0_11/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_11/Component_Function_0/N1  ( .A1(\SB1_0_11/i0[10] ), .A2(
        \SB1_0_11/i0[9] ), .ZN(\SB1_0_11/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_11/Component_Function_1/N3  ( .A1(\SB1_0_11/i1_5 ), .A2(
        \SB1_0_11/i0[6] ), .A3(\SB1_0_11/i0[9] ), .ZN(
        \SB1_0_11/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_11/Component_Function_1/N2  ( .A1(\SB1_0_11/i0_3 ), .A2(
        \SB1_0_11/i1_7 ), .A3(\SB1_0_11/i0[8] ), .ZN(
        \SB1_0_11/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_11/Component_Function_1/N1  ( .A1(\SB1_0_11/i0_3 ), .A2(
        \SB1_0_11/i1[9] ), .ZN(\SB1_0_11/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_11/Component_Function_5/N4  ( .A1(\SB1_0_11/i0[9] ), .A2(
        n306), .A3(n382), .ZN(\SB1_0_11/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_12/Component_Function_0/N2  ( .A1(\SB1_0_12/i0[8] ), .A2(
        \SB1_0_12/i0[7] ), .A3(\SB1_0_12/i0[6] ), .ZN(
        \SB1_0_12/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_12/Component_Function_0/N1  ( .A1(\SB1_0_12/i0[10] ), .A2(
        \SB1_0_12/i0[9] ), .ZN(\SB1_0_12/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_12/Component_Function_1/N4  ( .A1(\SB1_0_12/i1_7 ), .A2(
        \SB1_0_12/i0[8] ), .A3(\SB1_0_12/i0_4 ), .ZN(
        \SB1_0_12/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_12/Component_Function_1/N3  ( .A1(\SB1_0_12/i1_5 ), .A2(
        \SB1_0_12/i0[6] ), .A3(\SB1_0_12/i0[9] ), .ZN(
        \SB1_0_12/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_13/Component_Function_0/N2  ( .A1(\SB1_0_13/i0[8] ), .A2(
        \SB1_0_13/i0[7] ), .A3(\SB1_0_13/i0[6] ), .ZN(
        \SB1_0_13/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_13/Component_Function_0/N1  ( .A1(\SB1_0_13/i0[10] ), .A2(
        \SB1_0_13/i0[9] ), .ZN(\SB1_0_13/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_0_13/Component_Function_1/N1  ( .A1(\SB1_0_13/i0_3 ), .A2(
        \SB1_0_13/i1[9] ), .ZN(\SB1_0_13/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_14/Component_Function_0/N3  ( .A1(\SB1_0_14/i0[10] ), .A2(
        \SB1_0_14/i0_4 ), .A3(\SB1_0_14/i0_3 ), .ZN(
        \SB1_0_14/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_14/Component_Function_0/N2  ( .A1(\SB1_0_14/i0[8] ), .A2(
        \SB1_0_14/i0[7] ), .A3(\SB1_0_14/i0[6] ), .ZN(
        \SB1_0_14/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_14/Component_Function_0/N1  ( .A1(\SB1_0_14/i0[10] ), .A2(
        \SB1_0_14/i0[9] ), .ZN(\SB1_0_14/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_14/Component_Function_1/N4  ( .A1(\SB1_0_14/i1_7 ), .A2(
        \SB1_0_14/i0[8] ), .A3(\SB1_0_14/i0_4 ), .ZN(
        \SB1_0_14/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_14/Component_Function_1/N3  ( .A1(\SB1_0_14/i1_5 ), .A2(
        \SB1_0_14/i0[6] ), .A3(\SB1_0_14/i0[9] ), .ZN(
        \SB1_0_14/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB1_0_14/Component_Function_1/N1  ( .A1(\SB1_0_14/i0_3 ), .A2(
        \SB1_0_14/i1[9] ), .ZN(\SB1_0_14/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_14/Component_Function_5/N4  ( .A1(\SB1_0_14/i0[9] ), .A2(
        \SB1_0_14/i0[6] ), .A3(n376), .ZN(
        \SB1_0_14/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_15/Component_Function_0/N3  ( .A1(\SB1_0_15/i0[10] ), .A2(
        \SB1_0_15/i0_4 ), .A3(\SB1_0_15/i0_3 ), .ZN(
        \SB1_0_15/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_15/Component_Function_1/N4  ( .A1(\SB1_0_15/i1_7 ), .A2(
        \SB1_0_15/i0[8] ), .A3(\SB1_0_15/i0_4 ), .ZN(
        \SB1_0_15/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_15/Component_Function_1/N3  ( .A1(\SB1_0_15/i1_5 ), .A2(
        \SB1_0_15/i0[6] ), .A3(\SB1_0_15/i0[9] ), .ZN(
        \SB1_0_15/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_15/Component_Function_1/N2  ( .A1(\SB1_0_15/i0_3 ), .A2(
        \SB1_0_15/i1_7 ), .A3(\SB1_0_15/i0[8] ), .ZN(
        \SB1_0_15/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_15/Component_Function_5/N1  ( .A1(\SB1_0_15/i0_0 ), .A2(
        \SB1_0_15/i3[0] ), .ZN(\SB1_0_15/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_16/Component_Function_0/N2  ( .A1(\SB1_0_16/i0[8] ), .A2(
        \SB1_0_16/i0[7] ), .A3(\SB1_0_16/i0[6] ), .ZN(
        \SB1_0_16/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_16/Component_Function_0/N1  ( .A1(\SB1_0_16/i0[10] ), .A2(
        \SB1_0_16/i0[9] ), .ZN(\SB1_0_16/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_16/Component_Function_1/N3  ( .A1(\SB1_0_16/i1_5 ), .A2(
        \SB1_0_16/i0[6] ), .A3(\SB1_0_16/i0[9] ), .ZN(
        \SB1_0_16/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_17/Component_Function_0/N2  ( .A1(\SB1_0_17/i0[8] ), .A2(
        \SB1_0_17/i0[7] ), .A3(\SB1_0_17/i0[6] ), .ZN(
        \SB1_0_17/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_17/Component_Function_1/N3  ( .A1(\SB1_0_17/i1_5 ), .A2(n288), .A3(\SB1_0_17/i0[9] ), .ZN(\SB1_0_17/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_18/Component_Function_0/N2  ( .A1(\SB1_0_18/i0[8] ), .A2(
        \SB1_0_18/i0[7] ), .A3(\SB1_0_18/i0[6] ), .ZN(
        \SB1_0_18/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_18/Component_Function_0/N1  ( .A1(n1367), .A2(
        \SB1_0_18/i0[9] ), .ZN(\SB1_0_18/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_18/Component_Function_1/N4  ( .A1(\SB1_0_18/i1_7 ), .A2(
        \SB1_0_18/i0[8] ), .A3(n4753), .ZN(
        \SB1_0_18/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_18/Component_Function_1/N3  ( .A1(\SB1_0_18/i1_5 ), .A2(
        \SB1_0_18/i0[6] ), .A3(\SB1_0_18/i0[9] ), .ZN(
        \SB1_0_18/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_19/Component_Function_0/N3  ( .A1(\SB1_0_19/i0[10] ), .A2(
        \SB1_0_19/i0_4 ), .A3(\SB1_0_19/i0_3 ), .ZN(
        \SB1_0_19/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_19/Component_Function_0/N2  ( .A1(\SB1_0_19/i0[8] ), .A2(
        \SB1_0_19/i0[7] ), .A3(\SB1_0_19/i0[6] ), .ZN(
        \SB1_0_19/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_19/Component_Function_1/N4  ( .A1(\SB1_0_19/i1_7 ), .A2(
        \SB1_0_19/i0[8] ), .A3(\SB1_0_19/i0_4 ), .ZN(
        \SB1_0_19/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_19/Component_Function_1/N3  ( .A1(\SB1_0_19/i1_5 ), .A2(
        \SB1_0_19/i0[6] ), .A3(\SB1_0_19/i0[9] ), .ZN(
        \SB1_0_19/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_19/Component_Function_1/N2  ( .A1(\SB1_0_19/i0_3 ), .A2(
        \SB1_0_19/i1_7 ), .A3(\SB1_0_19/i0[8] ), .ZN(
        \SB1_0_19/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_20/Component_Function_0/N1  ( .A1(\SB1_0_20/i0[10] ), .A2(
        \SB1_0_20/i0[9] ), .ZN(\SB1_0_20/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_20/Component_Function_1/N3  ( .A1(\SB1_0_20/i1_5 ), .A2(
        \SB1_0_20/i0[6] ), .A3(\SB1_0_20/i0[9] ), .ZN(
        \SB1_0_20/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB1_0_20/Component_Function_1/N1  ( .A1(\SB1_0_20/i0_3 ), .A2(
        \SB1_0_20/i1[9] ), .ZN(\SB1_0_20/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_0_20/Component_Function_5/N1  ( .A1(\SB1_0_20/i0_0 ), .A2(
        \SB1_0_20/i3[0] ), .ZN(\SB1_0_20/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_21/Component_Function_0/N2  ( .A1(\SB1_0_21/i0[8] ), .A2(
        \SB1_0_21/i0[7] ), .A3(\SB1_0_21/i0[6] ), .ZN(
        \SB1_0_21/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_21/Component_Function_0/N1  ( .A1(\SB1_0_21/i0[10] ), .A2(
        \SB1_0_21/i0[9] ), .ZN(\SB1_0_21/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_21/Component_Function_1/N4  ( .A1(\SB1_0_21/i1_7 ), .A2(
        \SB1_0_21/i0[8] ), .A3(\SB1_0_21/i0_4 ), .ZN(
        \SB1_0_21/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB1_0_21/Component_Function_1/N1  ( .A1(\SB1_0_21/i0_3 ), .A2(
        \SB1_0_21/i1[9] ), .ZN(\SB1_0_21/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_22/Component_Function_0/N2  ( .A1(\SB1_0_22/i0[8] ), .A2(
        \SB1_0_22/i0[7] ), .A3(\SB1_0_22/i0[6] ), .ZN(
        \SB1_0_22/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_22/Component_Function_0/N1  ( .A1(\SB1_0_22/i0[10] ), .A2(
        \SB1_0_22/i0[9] ), .ZN(\SB1_0_22/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_22/Component_Function_1/N3  ( .A1(\SB1_0_22/i1_5 ), .A2(
        \SB1_0_22/i0[6] ), .A3(\SB1_0_22/i0[9] ), .ZN(
        \SB1_0_22/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_22/Component_Function_1/N2  ( .A1(\SB1_0_22/i0_3 ), .A2(
        \SB1_0_22/i1_7 ), .A3(\SB1_0_22/i0[8] ), .ZN(
        \SB1_0_22/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_22/Component_Function_1/N1  ( .A1(\SB1_0_22/i0_3 ), .A2(
        \SB1_0_22/i1[9] ), .ZN(\SB1_0_22/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_23/Component_Function_0/N4  ( .A1(\SB1_0_23/i0[7] ), .A2(
        \SB1_0_23/i0_3 ), .A3(\SB1_0_23/i0_0 ), .ZN(
        \SB1_0_23/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_23/Component_Function_0/N2  ( .A1(\SB1_0_23/i0[8] ), .A2(
        \SB1_0_23/i0[7] ), .A3(\SB1_0_23/i0[6] ), .ZN(
        \SB1_0_23/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_23/Component_Function_1/N2  ( .A1(\SB1_0_23/i0_3 ), .A2(
        \SB1_0_23/i1_7 ), .A3(\SB1_0_23/i0[8] ), .ZN(
        \SB1_0_23/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_23/Component_Function_1/N1  ( .A1(\SB1_0_23/i0_3 ), .A2(
        \SB1_0_23/i1[9] ), .ZN(\SB1_0_23/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_24/Component_Function_0/N4  ( .A1(\SB1_0_24/i0[7] ), .A2(
        \SB1_0_24/i0_3 ), .A3(\SB1_0_24/i0_0 ), .ZN(
        \SB1_0_24/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_24/Component_Function_0/N3  ( .A1(\SB1_0_24/i0[10] ), .A2(
        \SB1_0_24/i0_4 ), .A3(\SB1_0_24/i0_3 ), .ZN(
        \SB1_0_24/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_24/Component_Function_0/N2  ( .A1(\SB1_0_24/i0[8] ), .A2(
        \SB1_0_24/i0[7] ), .A3(\SB1_0_24/i0[6] ), .ZN(
        \SB1_0_24/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_24/Component_Function_0/N1  ( .A1(\SB1_0_24/i0[10] ), .A2(
        \SB1_0_24/i0[9] ), .ZN(\SB1_0_24/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_0_24/Component_Function_1/N1  ( .A1(\SB1_0_24/i0_3 ), .A2(
        \SB1_0_24/i1[9] ), .ZN(\SB1_0_24/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_0_25/Component_Function_0/N1  ( .A1(\SB1_0_25/i0[10] ), .A2(
        \SB1_0_25/i0[9] ), .ZN(\SB1_0_25/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_25/Component_Function_1/N4  ( .A1(\SB1_0_25/i1_7 ), .A2(
        \SB1_0_25/i0[8] ), .A3(\SB1_0_25/i0_4 ), .ZN(
        \SB1_0_25/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_26/Component_Function_0/N2  ( .A1(\SB1_0_26/i0[8] ), .A2(
        \SB1_0_26/i0[7] ), .A3(\SB1_0_26/i0[6] ), .ZN(
        \SB1_0_26/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_26/Component_Function_0/N1  ( .A1(\SB1_0_26/i0[10] ), .A2(
        \SB1_0_26/i0[9] ), .ZN(\SB1_0_26/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_26/Component_Function_1/N4  ( .A1(\SB1_0_26/i1_7 ), .A2(
        \SB1_0_26/i0[8] ), .A3(\SB1_0_26/i0_4 ), .ZN(
        \SB1_0_26/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_26/Component_Function_1/N3  ( .A1(\SB1_0_26/i1_5 ), .A2(
        \SB1_0_26/i0[6] ), .A3(n260), .ZN(
        \SB1_0_26/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB1_0_27/Component_Function_0/N1  ( .A1(\SB1_0_27/i0[10] ), .A2(
        \SB1_0_27/i0[9] ), .ZN(\SB1_0_27/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_27/Component_Function_1/N3  ( .A1(\SB1_0_27/i1_5 ), .A2(
        \SB1_0_27/i0[6] ), .A3(\SB1_0_27/i0[9] ), .ZN(
        \SB1_0_27/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_27/Component_Function_1/N2  ( .A1(\SB1_0_27/i0_3 ), .A2(
        \SB1_0_27/i1_7 ), .A3(\SB1_0_27/i0[8] ), .ZN(
        \SB1_0_27/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_27/Component_Function_1/N1  ( .A1(\SB1_0_27/i0_3 ), .A2(
        \SB1_0_27/i1[9] ), .ZN(\SB1_0_27/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_27/Component_Function_5/N2  ( .A1(\SB1_0_27/i0_0 ), .A2(
        \SB1_0_27/i0[6] ), .A3(\SB1_0_27/i0[10] ), .ZN(
        \SB1_0_27/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_28/Component_Function_0/N3  ( .A1(\SB1_0_28/i0[10] ), .A2(
        \SB1_0_28/i0_4 ), .A3(\SB1_0_28/i0_3 ), .ZN(
        \SB1_0_28/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_29/Component_Function_0/N2  ( .A1(\SB1_0_29/i0[8] ), .A2(
        \SB1_0_29/i0[7] ), .A3(\SB1_0_29/i0[6] ), .ZN(
        \SB1_0_29/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_29/Component_Function_0/N1  ( .A1(\SB1_0_29/i0[10] ), .A2(
        \SB1_0_29/i0[9] ), .ZN(\SB1_0_29/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_29/Component_Function_1/N3  ( .A1(\SB1_0_29/i1_5 ), .A2(
        \SB1_0_29/i0[6] ), .A3(n251), .ZN(
        \SB1_0_29/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB1_0_29/Component_Function_1/N1  ( .A1(\SB1_0_29/i0_3 ), .A2(
        \SB1_0_29/i1[9] ), .ZN(\SB1_0_29/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_30/Component_Function_0/N4  ( .A1(\SB1_0_30/i0[7] ), .A2(
        \SB1_0_30/i0_3 ), .A3(\SB1_0_30/i0_0 ), .ZN(
        \SB1_0_30/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_30/Component_Function_0/N3  ( .A1(\SB1_0_30/i0[10] ), .A2(
        \SB1_0_30/i0_4 ), .A3(\SB1_0_30/i0_3 ), .ZN(
        \SB1_0_30/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_30/Component_Function_0/N2  ( .A1(\SB1_0_30/i0[8] ), .A2(
        \SB1_0_30/i0[7] ), .A3(\SB1_0_30/i0[6] ), .ZN(
        \SB1_0_30/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_30/Component_Function_0/N1  ( .A1(\SB1_0_30/i0[10] ), .A2(
        \SB1_0_30/i0[9] ), .ZN(\SB1_0_30/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_30/Component_Function_1/N4  ( .A1(\SB1_0_30/i1_7 ), .A2(
        \SB1_0_30/i0[8] ), .A3(\SB1_0_30/i0_4 ), .ZN(
        \SB1_0_30/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_30/Component_Function_1/N3  ( .A1(\SB1_0_30/i1_5 ), .A2(
        \SB1_0_30/i0[6] ), .A3(\SB1_0_30/i0[9] ), .ZN(
        \SB1_0_30/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_30/Component_Function_1/N2  ( .A1(\SB1_0_30/i0_3 ), .A2(
        \SB1_0_30/i1_7 ), .A3(\SB1_0_30/i0[8] ), .ZN(
        \SB1_0_30/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_30/Component_Function_1/N1  ( .A1(\SB1_0_30/i0_3 ), .A2(
        \SB1_0_30/i1[9] ), .ZN(\SB1_0_30/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_30/Component_Function_5/N4  ( .A1(\SB1_0_30/i0[9] ), .A2(
        n249), .A3(n344), .ZN(\SB1_0_30/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB1_0_30/Component_Function_5/N1  ( .A1(\SB1_0_30/i0_0 ), .A2(
        \SB1_0_30/i3[0] ), .ZN(\SB1_0_30/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_31/Component_Function_0/N4  ( .A1(\SB1_0_31/i0[7] ), .A2(
        \SB1_0_31/i0_3 ), .A3(\SB1_0_31/i0_0 ), .ZN(
        \SB1_0_31/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_31/Component_Function_0/N3  ( .A1(\SB1_0_31/i0[10] ), .A2(
        \SB1_0_31/i0_4 ), .A3(\SB1_0_31/i0_3 ), .ZN(
        \SB1_0_31/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_31/Component_Function_0/N2  ( .A1(\SB1_0_31/i0[8] ), .A2(
        \SB1_0_31/i0[7] ), .A3(\SB1_0_31/i0[6] ), .ZN(
        \SB1_0_31/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_31/Component_Function_0/N1  ( .A1(\SB1_0_31/i0[10] ), .A2(
        \SB1_0_31/i0[9] ), .ZN(\SB1_0_31/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_31/Component_Function_1/N2  ( .A1(\SB1_0_31/i0_3 ), .A2(
        \SB1_0_31/i1_7 ), .A3(\SB1_0_31/i0[8] ), .ZN(
        \SB1_0_31/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_31/Component_Function_1/N1  ( .A1(\SB1_0_31/i0_3 ), .A2(
        \SB1_0_31/i1[9] ), .ZN(\SB1_0_31/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_31/Component_Function_5/N4  ( .A1(n245), .A2(
        \SB1_0_31/i0[6] ), .A3(n342), .ZN(
        \SB1_0_31/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_0/Component_Function_0/N3  ( .A1(\SB2_0_0/i0[10] ), .A2(
        \RI3[0][190] ), .A3(\RI3[0][191] ), .ZN(
        \SB2_0_0/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_0/Component_Function_0/N2  ( .A1(\SB2_0_0/i0[8] ), .A2(
        \SB2_0_0/i0[7] ), .A3(\SB2_0_0/i0[6] ), .ZN(
        \SB2_0_0/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_0/Component_Function_0/N1  ( .A1(\SB2_0_0/i0[10] ), .A2(
        \SB2_0_0/i0[9] ), .ZN(\SB2_0_0/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_0/Component_Function_1/N4  ( .A1(\SB2_0_0/i1_7 ), .A2(
        \SB2_0_0/i0[8] ), .A3(\RI3[0][190] ), .ZN(
        \SB2_0_0/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB2_0_0/Component_Function_1/N1  ( .A1(\RI3[0][191] ), .A2(
        \SB2_0_0/i1[9] ), .ZN(\SB2_0_0/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_0/Component_Function_5/N1  ( .A1(\SB2_0_0/i0_0 ), .A2(
        \SB2_0_0/i3[0] ), .ZN(\SB2_0_0/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_1/Component_Function_1/N1  ( .A1(\SB2_0_1/i0_3 ), .A2(
        \SB2_0_1/i1[9] ), .ZN(\SB2_0_1/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_2/Component_Function_0/N1  ( .A1(\SB2_0_2/i0[10] ), .A2(
        \SB2_0_2/i0[9] ), .ZN(\SB2_0_2/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_2/Component_Function_5/N1  ( .A1(\RI3[0][176] ), .A2(
        \SB2_0_2/i3[0] ), .ZN(\SB2_0_2/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_3/Component_Function_0/N2  ( .A1(\SB2_0_3/i0[8] ), .A2(
        \SB2_0_3/i0[7] ), .A3(\SB2_0_3/i0[6] ), .ZN(
        \SB2_0_3/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_3/Component_Function_0/N1  ( .A1(\SB2_0_3/i0[10] ), .A2(
        \SB2_0_3/i0[9] ), .ZN(\SB2_0_3/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_3/Component_Function_1/N4  ( .A1(\SB2_0_3/i1_7 ), .A2(
        \SB2_0_3/i0[8] ), .A3(\RI3[0][172] ), .ZN(
        \SB2_0_3/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_3/Component_Function_1/N2  ( .A1(\SB2_0_3/i0_3 ), .A2(
        \SB2_0_3/i1_7 ), .A3(\SB2_0_3/i0[8] ), .ZN(
        \SB2_0_3/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_3/Component_Function_1/N1  ( .A1(\SB2_0_3/i0_3 ), .A2(
        \SB2_0_3/i1[9] ), .ZN(\SB2_0_3/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_4/Component_Function_0/N4  ( .A1(\SB2_0_4/i0[7] ), .A2(
        \SB2_0_4/i0_3 ), .A3(\SB2_0_4/i0_0 ), .ZN(
        \SB2_0_4/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_4/Component_Function_1/N3  ( .A1(\SB2_0_4/i1_5 ), .A2(
        \SB2_0_4/i0[6] ), .A3(\SB2_0_4/i0[9] ), .ZN(
        \SB2_0_4/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_4/Component_Function_1/N2  ( .A1(\SB2_0_4/i0_3 ), .A2(
        \SB2_0_4/i1_7 ), .A3(\SB2_0_4/i0[8] ), .ZN(
        \SB2_0_4/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_4/Component_Function_5/N1  ( .A1(\SB2_0_4/i0_0 ), .A2(
        \SB2_0_4/i3[0] ), .ZN(\SB2_0_4/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_5/Component_Function_0/N1  ( .A1(\SB2_0_5/i0[10] ), .A2(
        \RI3[0][156] ), .ZN(\SB2_0_5/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_5/Component_Function_1/N3  ( .A1(\SB2_0_5/i1_5 ), .A2(
        \SB2_0_5/i0[6] ), .A3(\RI3[0][156] ), .ZN(
        \SB2_0_5/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_0_5/Component_Function_5/N1  ( .A1(\SB2_0_5/i0_0 ), .A2(
        \SB2_0_5/i3[0] ), .ZN(\SB2_0_5/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_6/Component_Function_0/N1  ( .A1(n2765), .A2(\SB2_0_6/i0[9] ), .ZN(\SB2_0_6/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_6/Component_Function_5/N1  ( .A1(\SB2_0_6/i0_0 ), .A2(
        \SB2_0_6/i3[0] ), .ZN(\SB2_0_6/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_7/Component_Function_1/N1  ( .A1(\SB2_0_7/i0_3 ), .A2(
        \SB2_0_7/i1[9] ), .ZN(\SB2_0_7/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_7/Component_Function_5/N1  ( .A1(\SB2_0_7/i0_0 ), .A2(
        \SB2_0_7/i3[0] ), .ZN(\SB2_0_7/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_8/Component_Function_0/N4  ( .A1(\SB2_0_8/i0[7] ), .A2(
        \SB2_0_8/i0_3 ), .A3(\SB2_0_8/i0_0 ), .ZN(
        \SB2_0_8/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_8/Component_Function_0/N2  ( .A1(\SB2_0_8/i0[8] ), .A2(
        \SB2_0_8/i0[7] ), .A3(\SB2_0_8/i0[6] ), .ZN(
        \SB2_0_8/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_8/Component_Function_0/N1  ( .A1(\SB2_0_8/i0[10] ), .A2(
        \SB2_0_8/i0[9] ), .ZN(\SB2_0_8/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_8/Component_Function_1/N4  ( .A1(\SB2_0_8/i1_7 ), .A2(
        \SB2_0_8/i0[8] ), .A3(\RI3[0][142] ), .ZN(
        \SB2_0_8/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB2_0_8/Component_Function_1/N1  ( .A1(\SB2_0_8/i0_3 ), .A2(
        \SB2_0_8/i1[9] ), .ZN(\SB2_0_8/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_9/Component_Function_0/N1  ( .A1(\SB2_0_9/i0[10] ), .A2(
        \SB2_0_9/i0[9] ), .ZN(\SB2_0_9/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_9/Component_Function_1/N3  ( .A1(n5518), .A2(\SB2_0_9/i0[6] ), .A3(\SB2_0_9/i0[9] ), .ZN(\SB2_0_9/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_0_10/Component_Function_0/N1  ( .A1(\SB2_0_10/i0[10] ), .A2(
        n571), .ZN(\SB2_0_10/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_10/Component_Function_1/N1  ( .A1(\SB2_0_10/i0_3 ), .A2(
        \SB2_0_10/i1[9] ), .ZN(\SB2_0_10/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_11/Component_Function_0/N3  ( .A1(\SB2_0_11/i0[10] ), .A2(
        \SB2_0_11/i0_4 ), .A3(\SB2_0_11/i0_3 ), .ZN(
        \SB2_0_11/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB2_0_11/Component_Function_0/N1  ( .A1(\SB2_0_11/i0[10] ), .A2(
        n1911), .ZN(\SB2_0_11/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_11/Component_Function_1/N3  ( .A1(\SB2_0_11/i1_5 ), .A2(
        \SB2_0_11/i0[6] ), .A3(n1911), .ZN(
        \SB2_0_11/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_11/Component_Function_1/N2  ( .A1(\SB2_0_11/i0_3 ), .A2(
        \SB2_0_11/i1_7 ), .A3(\SB2_0_11/i0[8] ), .ZN(
        \SB2_0_11/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_11/Component_Function_1/N1  ( .A1(\SB2_0_11/i0_3 ), .A2(
        \SB2_0_11/i1[9] ), .ZN(\SB2_0_11/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_12/Component_Function_0/N4  ( .A1(\SB2_0_12/i0[7] ), .A2(
        \SB2_0_12/i0_3 ), .A3(\SB2_0_12/i0_0 ), .ZN(
        \SB2_0_12/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_12/Component_Function_0/N3  ( .A1(\SB2_0_12/i0[10] ), .A2(
        \SB2_0_12/i0_4 ), .A3(\SB2_0_12/i0_3 ), .ZN(
        \SB2_0_12/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_12/Component_Function_0/N2  ( .A1(\SB2_0_12/i0[8] ), .A2(
        \SB2_0_12/i0[7] ), .A3(\SB2_0_12/i0[6] ), .ZN(
        \SB2_0_12/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_12/Component_Function_0/N1  ( .A1(\SB2_0_12/i0[10] ), .A2(
        \SB2_0_12/i0[9] ), .ZN(\SB2_0_12/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_12/Component_Function_1/N4  ( .A1(\SB2_0_12/i1_7 ), .A2(
        \SB2_0_12/i0[8] ), .A3(\SB2_0_12/i0_4 ), .ZN(
        \SB2_0_12/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_12/Component_Function_1/N3  ( .A1(\SB2_0_12/i1_5 ), .A2(
        \SB2_0_12/i0[6] ), .A3(\SB2_0_12/i0[9] ), .ZN(
        \SB2_0_12/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_12/Component_Function_1/N2  ( .A1(\SB2_0_12/i0_3 ), .A2(
        \SB2_0_12/i1_7 ), .A3(\SB2_0_12/i0[8] ), .ZN(
        \SB2_0_12/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_12/Component_Function_1/N1  ( .A1(\SB2_0_12/i0_3 ), .A2(
        \SB2_0_12/i1[9] ), .ZN(\SB2_0_12/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_12/Component_Function_5/N1  ( .A1(\SB2_0_12/i0_0 ), .A2(
        \SB2_0_12/i3[0] ), .ZN(\SB2_0_12/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_13/Component_Function_0/N3  ( .A1(\SB2_0_13/i0[10] ), .A2(
        \SB2_0_13/i0_4 ), .A3(\SB2_0_13/i0_3 ), .ZN(
        \SB2_0_13/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_13/Component_Function_0/N2  ( .A1(n1393), .A2(n2711), .A3(
        \SB1_0_17/buf_output[1] ), .ZN(
        \SB2_0_13/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_13/Component_Function_0/N1  ( .A1(\SB2_0_13/i0[10] ), .A2(
        \SB2_0_13/i0[9] ), .ZN(\SB2_0_13/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_13/Component_Function_5/N1  ( .A1(\SB2_0_13/i0_0 ), .A2(
        \SB2_0_13/i3[0] ), .ZN(\SB2_0_13/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_14/Component_Function_0/N4  ( .A1(\SB2_0_14/i0[7] ), .A2(
        \SB2_0_14/i0_3 ), .A3(\RI3[0][104] ), .ZN(
        \SB2_0_14/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB2_0_14/Component_Function_0/N1  ( .A1(\RI3[0][105] ), .A2(
        \SB2_0_14/i0[9] ), .ZN(\SB2_0_14/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_14/Component_Function_5/N1  ( .A1(\RI3[0][104] ), .A2(
        \SB2_0_14/i3[0] ), .ZN(\SB2_0_14/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_15/Component_Function_0/N1  ( .A1(\SB2_0_15/i0[10] ), .A2(
        \SB2_0_15/i0[9] ), .ZN(\SB2_0_15/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_15/Component_Function_1/N3  ( .A1(\SB2_0_15/i1_5 ), .A2(
        \SB2_0_15/i0[6] ), .A3(\RI3[0][96] ), .ZN(
        \SB2_0_15/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_0_15/Component_Function_1/N1  ( .A1(\SB2_0_15/i0_3 ), .A2(
        \SB2_0_15/i1[9] ), .ZN(\SB2_0_15/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_15/Component_Function_5/N1  ( .A1(\SB2_0_15/i0_0 ), .A2(
        \SB2_0_15/i3[0] ), .ZN(\SB2_0_15/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_16/Component_Function_0/N4  ( .A1(n2682), .A2(
        \SB2_0_16/i0_3 ), .A3(\SB2_0_16/i0_0 ), .ZN(
        \SB2_0_16/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_16/Component_Function_0/N2  ( .A1(\SB2_0_16/i0[8] ), .A2(
        n2682), .A3(\SB2_0_16/i0[6] ), .ZN(
        \SB2_0_16/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_16/Component_Function_0/N1  ( .A1(\SB2_0_16/i0[10] ), .A2(
        \SB2_0_16/i0[9] ), .ZN(\SB2_0_16/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_16/Component_Function_1/N1  ( .A1(\SB2_0_16/i0_3 ), .A2(
        \SB2_0_16/i1[9] ), .ZN(\SB2_0_16/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_16/Component_Function_5/N1  ( .A1(\SB2_0_16/i0_0 ), .A2(
        \SB2_0_16/i3[0] ), .ZN(\SB2_0_16/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_17/Component_Function_0/N1  ( .A1(\SB2_0_17/i0[10] ), .A2(
        \RI3[0][84] ), .ZN(\SB2_0_17/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_18/Component_Function_0/N2  ( .A1(\SB2_0_18/i0[8] ), .A2(
        \SB2_0_18/i0[7] ), .A3(\SB2_0_18/i0[6] ), .ZN(
        \SB2_0_18/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_18/Component_Function_1/N2  ( .A1(\SB2_0_18/i0_3 ), .A2(
        \SB2_0_18/i1_7 ), .A3(\SB2_0_18/i0[8] ), .ZN(
        \SB2_0_18/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_18/Component_Function_1/N1  ( .A1(\SB2_0_18/i0_3 ), .A2(
        \SB2_0_18/i1[9] ), .ZN(\SB2_0_18/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_19/Component_Function_0/N4  ( .A1(\SB2_0_19/i0[7] ), .A2(
        \SB2_0_19/i0_3 ), .A3(\SB2_0_19/i0_0 ), .ZN(
        \SB2_0_19/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB2_0_19/Component_Function_0/N1  ( .A1(n2774), .A2(
        \SB2_0_19/i0[9] ), .ZN(\SB2_0_19/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_19/Component_Function_1/N4  ( .A1(\SB2_0_19/i1_7 ), .A2(
        \SB2_0_19/i0[8] ), .A3(\RI3[0][76] ), .ZN(
        \SB2_0_19/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_19/Component_Function_1/N3  ( .A1(\SB2_0_19/i1_5 ), .A2(
        \SB2_0_19/i0[6] ), .A3(\SB2_0_19/i0[9] ), .ZN(
        \SB2_0_19/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_19/Component_Function_1/N2  ( .A1(\SB2_0_19/i0_3 ), .A2(
        \SB2_0_19/i1_7 ), .A3(\SB2_0_19/i0[8] ), .ZN(
        \SB2_0_19/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_19/Component_Function_1/N1  ( .A1(\SB2_0_19/i0_3 ), .A2(
        \SB2_0_19/i1[9] ), .ZN(\SB2_0_19/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_20/Component_Function_0/N1  ( .A1(\SB2_0_20/i0[10] ), .A2(
        \SB2_0_20/i0[9] ), .ZN(\SB2_0_20/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_20/Component_Function_1/N1  ( .A1(\SB2_0_20/i0_3 ), .A2(
        \SB2_0_20/i1[9] ), .ZN(\SB2_0_20/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_20/Component_Function_5/N1  ( .A1(\SB2_0_20/i0_0 ), .A2(
        \SB2_0_20/i3[0] ), .ZN(\SB2_0_20/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_21/Component_Function_0/N4  ( .A1(\SB2_0_21/i0[7] ), .A2(
        \SB2_0_21/i0_3 ), .A3(\SB2_0_21/i0_0 ), .ZN(
        \SB2_0_21/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_21/Component_Function_0/N2  ( .A1(\SB2_0_21/i0[8] ), .A2(
        \SB2_0_21/i0[7] ), .A3(\SB2_0_21/i0[6] ), .ZN(
        \SB2_0_21/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_21/Component_Function_0/N1  ( .A1(\SB2_0_21/i0[10] ), .A2(
        \SB2_0_21/i0[9] ), .ZN(\SB2_0_21/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_21/Component_Function_1/N1  ( .A1(\SB2_0_21/i0_3 ), .A2(
        \SB2_0_21/i1[9] ), .ZN(\SB2_0_21/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_22/Component_Function_0/N2  ( .A1(\SB2_0_22/i0[8] ), .A2(
        \SB2_0_22/i0[7] ), .A3(\SB2_0_22/i0[6] ), .ZN(
        \SB2_0_22/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_22/Component_Function_0/N1  ( .A1(\SB2_0_22/i0[10] ), .A2(
        \RI3[0][54] ), .ZN(\SB2_0_22/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_22/Component_Function_1/N1  ( .A1(\SB2_0_22/i0_3 ), .A2(
        \SB2_0_22/i1[9] ), .ZN(\SB2_0_22/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_22/Component_Function_5/N1  ( .A1(\SB2_0_22/i0_0 ), .A2(
        \SB2_0_22/i3[0] ), .ZN(\SB2_0_22/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_23/Component_Function_0/N4  ( .A1(n2877), .A2(
        \SB2_0_23/i0_3 ), .A3(\SB2_0_23/i0_0 ), .ZN(
        \SB2_0_23/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB2_0_23/Component_Function_0/N1  ( .A1(\SB2_0_23/i0[10] ), .A2(
        \SB2_0_23/i0[9] ), .ZN(\SB2_0_23/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_23/Component_Function_1/N1  ( .A1(\SB2_0_23/i0_3 ), .A2(
        \SB2_0_23/i1[9] ), .ZN(\SB2_0_23/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_24/Component_Function_0/N4  ( .A1(\SB2_0_24/i0[7] ), .A2(
        \SB2_0_24/i0_3 ), .A3(\SB2_0_24/i0_0 ), .ZN(
        \SB2_0_24/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB2_0_24/Component_Function_0/N1  ( .A1(\SB2_0_24/i0[10] ), .A2(
        \SB2_0_24/i0[9] ), .ZN(\SB2_0_24/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_25/Component_Function_0/N2  ( .A1(\SB2_0_25/i0[8] ), .A2(
        \SB2_0_25/i0[7] ), .A3(\RI3[0][37] ), .ZN(
        \SB2_0_25/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_25/Component_Function_1/N4  ( .A1(\SB2_0_25/i1_7 ), .A2(
        \SB2_0_25/i0[8] ), .A3(\SB1_0_26/buf_output[4] ), .ZN(
        \SB2_0_25/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB2_0_25/Component_Function_1/N1  ( .A1(\SB2_0_25/i0_3 ), .A2(
        \SB2_0_25/i1[9] ), .ZN(\SB2_0_25/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_25/Component_Function_5/N1  ( .A1(\SB2_0_25/i0_0 ), .A2(
        \SB2_0_25/i3[0] ), .ZN(\SB2_0_25/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_26/Component_Function_0/N4  ( .A1(\SB2_0_26/i0[7] ), .A2(
        \SB2_0_26/i0_3 ), .A3(\SB2_0_26/i0_0 ), .ZN(
        \SB2_0_26/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_26/Component_Function_0/N2  ( .A1(\SB2_0_26/i0[8] ), .A2(
        \SB2_0_26/i0[7] ), .A3(\SB2_0_26/i0[6] ), .ZN(
        \SB2_0_26/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_26/Component_Function_0/N1  ( .A1(\SB2_0_26/i0[10] ), .A2(
        \SB2_0_26/i0[9] ), .ZN(\SB2_0_26/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_26/Component_Function_1/N3  ( .A1(\SB2_0_26/i1_5 ), .A2(
        \SB2_0_26/i0[6] ), .A3(\SB2_0_26/i0[9] ), .ZN(
        \SB2_0_26/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_0_27/Component_Function_1/N1  ( .A1(\SB2_0_27/i0_3 ), .A2(
        \SB2_0_27/i1[9] ), .ZN(\SB2_0_27/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_28/Component_Function_0/N1  ( .A1(\SB2_0_28/i0[10] ), .A2(
        \RI3[0][18] ), .ZN(\SB2_0_28/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_28/Component_Function_1/N1  ( .A1(\SB2_0_28/i0_3 ), .A2(
        \SB2_0_28/i1[9] ), .ZN(\SB2_0_28/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_29/Component_Function_0/N4  ( .A1(\SB2_0_29/i0[7] ), .A2(
        \SB2_0_29/i0_3 ), .A3(\SB2_0_29/i0_0 ), .ZN(
        \SB2_0_29/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_29/Component_Function_0/N3  ( .A1(\RI3[0][15] ), .A2(
        \SB2_0_29/i0_4 ), .A3(\SB2_0_29/i0_3 ), .ZN(
        \SB2_0_29/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB2_0_29/Component_Function_0/N1  ( .A1(\RI3[0][15] ), .A2(n2605), 
        .ZN(\SB2_0_29/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_29/Component_Function_1/N3  ( .A1(\SB2_0_29/i1_5 ), .A2(
        \SB2_0_29/i0[6] ), .A3(n2605), .ZN(
        \SB2_0_29/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_29/Component_Function_1/N2  ( .A1(\SB2_0_29/i0_3 ), .A2(
        \SB2_0_29/i1_7 ), .A3(\SB2_0_29/i0[8] ), .ZN(
        \SB2_0_29/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_29/Component_Function_1/N1  ( .A1(\SB2_0_29/i0_3 ), .A2(
        \SB2_0_29/i1[9] ), .ZN(\SB2_0_29/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_30/Component_Function_0/N3  ( .A1(\SB2_0_30/i0[10] ), .A2(
        \RI3[0][10] ), .A3(\SB2_0_30/i0_3 ), .ZN(
        \SB2_0_30/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB2_0_30/Component_Function_0/N1  ( .A1(\SB2_0_30/i0[10] ), .A2(
        \SB2_0_30/i0[9] ), .ZN(\SB2_0_30/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_30/Component_Function_1/N1  ( .A1(\SB2_0_30/i0_3 ), .A2(
        \SB2_0_30/i1[9] ), .ZN(\SB2_0_30/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_31/Component_Function_0/N4  ( .A1(\SB2_0_31/i0[7] ), .A2(
        \SB2_0_31/i0_3 ), .A3(\SB2_0_31/i0_0 ), .ZN(
        \SB2_0_31/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_31/Component_Function_0/N3  ( .A1(\SB2_0_31/i0[10] ), .A2(
        \RI3[0][4] ), .A3(\SB2_0_31/i0_3 ), .ZN(
        \SB2_0_31/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_31/Component_Function_0/N2  ( .A1(\SB2_0_31/i0[8] ), .A2(
        \SB2_0_31/i0[7] ), .A3(\SB2_0_31/i0[6] ), .ZN(
        \SB2_0_31/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_31/Component_Function_0/N1  ( .A1(\SB2_0_31/i0[10] ), .A2(
        \SB2_0_31/i0[9] ), .ZN(\SB2_0_31/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_31/Component_Function_1/N3  ( .A1(\SB2_0_31/i1_5 ), .A2(
        \SB2_0_31/i0[6] ), .A3(\SB2_0_31/i0[9] ), .ZN(
        \SB2_0_31/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_31/Component_Function_1/N2  ( .A1(\SB2_0_31/i0_3 ), .A2(
        \SB2_0_31/i1_7 ), .A3(\SB2_0_31/i0[8] ), .ZN(
        \SB2_0_31/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_31/Component_Function_1/N1  ( .A1(\SB2_0_31/i0_3 ), .A2(
        \SB2_0_31/i1[9] ), .ZN(\SB2_0_31/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_0/Component_Function_0/N1  ( .A1(\SB1_1_0/i0[10] ), .A2(
        \SB1_1_0/i0[9] ), .ZN(\SB1_1_0/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_0/Component_Function_1/N4  ( .A1(\SB1_1_0/i1_7 ), .A2(
        \SB1_1_0/i0[8] ), .A3(\SB1_1_0/i0_4 ), .ZN(
        \SB1_1_0/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_1/Component_Function_0/N3  ( .A1(\SB1_1_1/i0[10] ), .A2(
        \SB1_1_1/i0_4 ), .A3(\SB1_1_1/i0_3 ), .ZN(
        \SB1_1_1/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_1/Component_Function_0/N2  ( .A1(\SB1_1_1/i0[8] ), .A2(
        \SB1_1_1/i0[7] ), .A3(\SB1_1_1/i0[6] ), .ZN(
        \SB1_1_1/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_1/Component_Function_0/N1  ( .A1(\SB1_1_1/i0[10] ), .A2(
        \SB1_1_1/i0[9] ), .ZN(\SB1_1_1/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_1/Component_Function_1/N3  ( .A1(\SB1_1_1/i1_5 ), .A2(
        \SB1_1_1/i0[6] ), .A3(\SB1_1_1/i0[9] ), .ZN(
        \SB1_1_1/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_2/Component_Function_0/N3  ( .A1(\SB1_1_2/i0[10] ), .A2(
        \SB1_1_2/i0_4 ), .A3(\SB1_1_2/i0_3 ), .ZN(
        \SB1_1_2/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_1_2/Component_Function_1/N1  ( .A1(\SB1_1_2/i0_3 ), .A2(
        \SB1_1_2/i1[9] ), .ZN(\SB1_1_2/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_3/Component_Function_0/N3  ( .A1(\SB1_1_3/i0[10] ), .A2(
        \SB1_1_3/i0_4 ), .A3(\SB1_1_3/i0_3 ), .ZN(
        \SB1_1_3/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_1_3/Component_Function_0/N1  ( .A1(\SB1_1_3/i0[10] ), .A2(
        \SB1_1_3/i0[9] ), .ZN(\SB1_1_3/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_3/Component_Function_1/N2  ( .A1(\SB1_1_3/i0_3 ), .A2(
        \SB1_1_3/i1_7 ), .A3(\SB1_1_3/i0[8] ), .ZN(
        \SB1_1_3/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_3/Component_Function_1/N1  ( .A1(\SB1_1_3/i0_3 ), .A2(
        \SB1_1_3/i1[9] ), .ZN(\SB1_1_3/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_4/Component_Function_0/N3  ( .A1(\SB1_1_4/i0[10] ), .A2(
        \SB1_1_4/i0_4 ), .A3(\SB1_1_4/i0_3 ), .ZN(
        \SB1_1_4/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_4/Component_Function_0/N2  ( .A1(\SB1_1_4/i0[8] ), .A2(
        \SB1_1_4/i0[7] ), .A3(\SB1_1_4/i0[6] ), .ZN(
        \SB1_1_4/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_4/Component_Function_0/N1  ( .A1(\SB1_1_4/i0[10] ), .A2(
        \SB1_1_4/i0[9] ), .ZN(\SB1_1_4/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_4/Component_Function_1/N1  ( .A1(\SB1_1_4/i0_3 ), .A2(
        \SB1_1_4/i1[9] ), .ZN(\SB1_1_4/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_5/Component_Function_0/N4  ( .A1(\SB1_1_5/i0[7] ), .A2(
        \SB1_1_5/i0_3 ), .A3(\SB1_1_5/i0_0 ), .ZN(
        \SB1_1_5/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_5/Component_Function_0/N3  ( .A1(\SB1_1_5/i0[10] ), .A2(
        \SB1_1_5/i0_4 ), .A3(\SB1_1_5/i0_3 ), .ZN(
        \SB1_1_5/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_1_5/Component_Function_0/N1  ( .A1(\SB1_1_5/i0[10] ), .A2(
        \SB1_1_5/i0[9] ), .ZN(\SB1_1_5/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_5/Component_Function_1/N2  ( .A1(\SB1_1_5/i0_3 ), .A2(
        \SB1_1_5/i1_7 ), .A3(\SB1_1_5/i0[8] ), .ZN(
        \SB1_1_5/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_5/Component_Function_1/N1  ( .A1(\SB1_1_5/i0_3 ), .A2(
        \SB1_1_5/i1[9] ), .ZN(\SB1_1_5/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_6/Component_Function_0/N2  ( .A1(\SB1_1_6/i0[8] ), .A2(
        \SB1_1_6/i0[7] ), .A3(\SB1_1_6/i0[6] ), .ZN(
        \SB1_1_6/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_6/Component_Function_0/N1  ( .A1(\SB1_1_6/i0[10] ), .A2(
        \SB1_1_6/i0[9] ), .ZN(\SB1_1_6/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_7/Component_Function_0/N2  ( .A1(\SB1_1_7/i0[8] ), .A2(
        \SB1_1_7/i0[7] ), .A3(\SB1_1_7/i0[6] ), .ZN(
        \SB1_1_7/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_7/Component_Function_0/N1  ( .A1(\SB1_1_7/i0[10] ), .A2(
        \SB1_1_7/i0[9] ), .ZN(\SB1_1_7/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_7/Component_Function_1/N1  ( .A1(\SB1_1_7/i0_3 ), .A2(
        \SB1_1_7/i1[9] ), .ZN(\SB1_1_7/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_8/Component_Function_0/N1  ( .A1(\SB1_1_8/i0[10] ), .A2(
        \SB1_1_8/i0[9] ), .ZN(\SB1_1_8/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_8/Component_Function_1/N1  ( .A1(\RI1[1][143] ), .A2(
        \SB1_1_8/i1[9] ), .ZN(\SB1_1_8/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_9/Component_Function_0/N3  ( .A1(\SB1_1_9/i0[10] ), .A2(
        \SB1_1_9/i0_4 ), .A3(\SB1_1_9/i0_3 ), .ZN(
        \SB1_1_9/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_1_9/Component_Function_0/N1  ( .A1(\SB1_1_9/i0[10] ), .A2(
        \SB1_1_9/i0[9] ), .ZN(\SB1_1_9/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_9/Component_Function_1/N1  ( .A1(\SB1_1_9/i0_3 ), .A2(
        \SB1_1_9/i1[9] ), .ZN(\SB1_1_9/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_10/Component_Function_0/N3  ( .A1(\SB1_1_10/i0[10] ), .A2(
        \SB1_1_10/i0_4 ), .A3(\SB1_1_10/i0_3 ), .ZN(
        \SB1_1_10/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_10/Component_Function_0/N2  ( .A1(\SB1_1_10/i0[8] ), .A2(
        \SB1_1_10/i0[7] ), .A3(\SB1_1_10/i0[6] ), .ZN(
        \SB1_1_10/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_10/Component_Function_0/N1  ( .A1(\SB1_1_10/i0[10] ), .A2(
        \SB1_1_10/i0[9] ), .ZN(\SB1_1_10/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_10/Component_Function_1/N1  ( .A1(\SB1_1_10/i0_3 ), .A2(
        \SB1_1_10/i1[9] ), .ZN(\SB1_1_10/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_11/Component_Function_0/N2  ( .A1(\SB1_1_11/i0[8] ), .A2(
        \SB1_1_11/i0[7] ), .A3(\SB1_1_11/i0[6] ), .ZN(
        \SB1_1_11/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_11/Component_Function_0/N1  ( .A1(\SB1_1_11/i0[10] ), .A2(
        \SB1_1_11/i0[9] ), .ZN(\SB1_1_11/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_11/Component_Function_1/N3  ( .A1(\SB1_1_11/i1_5 ), .A2(
        \SB1_1_11/i0[6] ), .A3(\SB1_1_11/i0[9] ), .ZN(
        \SB1_1_11/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_12/Component_Function_0/N2  ( .A1(\SB1_1_12/i0[8] ), .A2(
        \SB1_1_12/i0[7] ), .A3(\SB1_1_12/i0[6] ), .ZN(
        \SB1_1_12/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_12/Component_Function_0/N1  ( .A1(\SB1_1_12/i0[10] ), .A2(
        \SB1_1_12/i0[9] ), .ZN(\SB1_1_12/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_12/Component_Function_1/N1  ( .A1(\SB1_1_12/i0_3 ), .A2(
        \SB1_1_12/i1[9] ), .ZN(\SB1_1_12/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_13/Component_Function_0/N3  ( .A1(\SB1_1_13/i0[10] ), .A2(
        \SB1_1_13/i0_4 ), .A3(\SB1_1_13/i0_3 ), .ZN(
        \SB1_1_13/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_14/Component_Function_0/N3  ( .A1(\SB1_1_14/i0[10] ), .A2(
        \SB1_1_14/i0_4 ), .A3(\SB1_1_14/i0_3 ), .ZN(
        \SB1_1_14/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_14/Component_Function_0/N2  ( .A1(\SB1_1_14/i0[8] ), .A2(
        \SB1_1_14/i0[7] ), .A3(\SB1_1_14/i0[6] ), .ZN(
        \SB1_1_14/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_14/Component_Function_0/N1  ( .A1(\SB1_1_14/i0[10] ), .A2(
        \SB1_1_14/i0[9] ), .ZN(\SB1_1_14/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_14/Component_Function_1/N2  ( .A1(\SB1_1_14/i0_3 ), .A2(
        \SB1_1_14/i1_7 ), .A3(\SB1_1_14/i0[8] ), .ZN(
        \SB1_1_14/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_15/Component_Function_0/N1  ( .A1(\SB1_1_15/i0[10] ), .A2(
        \SB1_1_15/i0[9] ), .ZN(\SB1_1_15/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_15/Component_Function_1/N1  ( .A1(\SB1_1_15/i0_3 ), .A2(
        \SB1_1_15/i1[9] ), .ZN(\SB1_1_15/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_17/Component_Function_0/N3  ( .A1(\SB1_1_17/i0[10] ), .A2(
        \SB1_1_17/i0_4 ), .A3(\SB1_1_17/i0_3 ), .ZN(
        \SB1_1_17/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_17/Component_Function_0/N2  ( .A1(\SB1_1_17/i0[8] ), .A2(
        \SB1_1_17/i0[7] ), .A3(\SB1_1_17/i0[6] ), .ZN(
        \SB1_1_17/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_17/Component_Function_0/N1  ( .A1(\SB1_1_17/i0[10] ), .A2(
        \SB1_1_17/i0[9] ), .ZN(\SB1_1_17/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_18/Component_Function_0/N2  ( .A1(\SB1_1_18/i0[8] ), .A2(
        \SB1_1_18/i0[7] ), .A3(\SB1_1_18/i0[6] ), .ZN(
        \SB1_1_18/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_18/Component_Function_0/N1  ( .A1(\SB1_1_18/i0[10] ), .A2(
        \SB1_1_18/i0[9] ), .ZN(\SB1_1_18/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_18/Component_Function_1/N3  ( .A1(\SB1_1_18/i1_5 ), .A2(
        \SB1_1_18/i0[6] ), .A3(\SB1_1_18/i0[9] ), .ZN(
        \SB1_1_18/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_18/Component_Function_1/N2  ( .A1(\SB1_1_18/i0_3 ), .A2(
        \SB1_1_18/i1_7 ), .A3(\SB1_1_18/i0[8] ), .ZN(
        \SB1_1_18/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_18/Component_Function_1/N1  ( .A1(\SB1_1_18/i0_3 ), .A2(
        \SB1_1_18/i1[9] ), .ZN(\SB1_1_18/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_19/Component_Function_0/N2  ( .A1(\SB1_1_19/i0[8] ), .A2(
        \SB1_1_19/i0[7] ), .A3(\SB1_1_19/i0[6] ), .ZN(
        \SB1_1_19/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_19/Component_Function_0/N1  ( .A1(\SB1_1_19/i0[10] ), .A2(
        \SB1_1_19/i0[9] ), .ZN(\SB1_1_19/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_19/Component_Function_1/N1  ( .A1(\SB1_1_19/i0_3 ), .A2(
        \SB1_1_19/i1[9] ), .ZN(\SB1_1_19/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_21/Component_Function_0/N4  ( .A1(\SB1_1_21/i0[7] ), .A2(
        \SB1_1_21/i0_3 ), .A3(\SB1_1_21/i0_0 ), .ZN(
        \SB1_1_21/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB1_1_21/Component_Function_1/N1  ( .A1(\SB1_1_21/i0_3 ), .A2(
        \SB1_1_21/i1[9] ), .ZN(\SB1_1_21/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_22/Component_Function_0/N1  ( .A1(\SB1_1_22/i0[10] ), .A2(
        \SB1_1_22/i0[9] ), .ZN(\SB1_1_22/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_22/Component_Function_1/N1  ( .A1(\RI1[1][59] ), .A2(
        \SB1_1_22/i1[9] ), .ZN(\SB1_1_22/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_23/Component_Function_0/N3  ( .A1(\SB1_1_23/i0[10] ), .A2(
        \SB1_1_23/i0_4 ), .A3(\SB1_1_23/i0_3 ), .ZN(
        \SB1_1_23/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_23/Component_Function_0/N2  ( .A1(\SB1_1_23/i0[8] ), .A2(
        \SB1_1_23/i0[7] ), .A3(\SB1_1_23/i0[6] ), .ZN(
        \SB1_1_23/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_24/Component_Function_0/N2  ( .A1(\SB1_1_24/i0[8] ), .A2(
        \SB1_1_24/i0[7] ), .A3(\SB1_1_24/i0[6] ), .ZN(
        \SB1_1_24/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_25/Component_Function_0/N3  ( .A1(\SB1_1_25/i0[10] ), .A2(
        \SB1_1_25/i0_4 ), .A3(\SB1_1_25/i0_3 ), .ZN(
        \SB1_1_25/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_25/Component_Function_0/N2  ( .A1(\SB1_1_25/i0[8] ), .A2(
        \SB1_1_25/i0[7] ), .A3(\SB1_1_25/i0[6] ), .ZN(
        \SB1_1_25/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_25/Component_Function_0/N1  ( .A1(\SB1_1_25/i0[10] ), .A2(
        \SB1_1_25/i0[9] ), .ZN(\SB1_1_25/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_25/Component_Function_1/N3  ( .A1(\SB1_1_25/i1_5 ), .A2(
        \SB1_1_25/i0[6] ), .A3(\SB1_1_25/i0[9] ), .ZN(
        \SB1_1_25/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_25/Component_Function_5/N2  ( .A1(\SB1_1_25/i0_0 ), .A2(
        \SB1_1_25/i0[6] ), .A3(\SB1_1_25/i0[10] ), .ZN(
        \SB1_1_25/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_26/Component_Function_0/N3  ( .A1(\SB1_1_26/i0[10] ), .A2(
        \SB1_1_26/i0_4 ), .A3(\SB1_1_26/i0_3 ), .ZN(
        \SB1_1_26/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_26/Component_Function_0/N2  ( .A1(\SB1_1_26/i0[8] ), .A2(
        \SB1_1_26/i0[7] ), .A3(\SB1_1_26/i0[6] ), .ZN(
        \SB1_1_26/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_26/Component_Function_0/N1  ( .A1(\SB1_1_26/i0[10] ), .A2(
        \SB1_1_26/i0[9] ), .ZN(\SB1_1_26/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_26/Component_Function_1/N3  ( .A1(\SB1_1_26/i1_5 ), .A2(
        \SB1_1_26/i0[6] ), .A3(\SB1_1_26/i0[9] ), .ZN(
        \SB1_1_26/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_26/Component_Function_1/N2  ( .A1(\SB1_1_26/i0_3 ), .A2(
        \SB1_1_26/i1_7 ), .A3(\SB1_1_26/i0[8] ), .ZN(
        \SB1_1_26/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_27/Component_Function_0/N4  ( .A1(\SB1_1_27/i0[7] ), .A2(
        \SB1_1_27/i0_3 ), .A3(\SB1_1_27/i0_0 ), .ZN(
        \SB1_1_27/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_27/Component_Function_0/N2  ( .A1(\SB1_1_27/i0[8] ), .A2(
        \SB1_1_27/i0[7] ), .A3(\SB1_1_27/i0[6] ), .ZN(
        \SB1_1_27/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_27/Component_Function_0/N1  ( .A1(\SB1_1_27/i0[10] ), .A2(
        \SB1_1_27/i0[9] ), .ZN(\SB1_1_27/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_28/Component_Function_0/N4  ( .A1(\SB1_1_28/i0[7] ), .A2(
        \SB1_1_28/i0_3 ), .A3(\SB1_1_28/i0_0 ), .ZN(
        \SB1_1_28/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB1_1_28/Component_Function_0/N1  ( .A1(\SB1_1_28/i0[10] ), .A2(
        \SB1_1_28/i0[9] ), .ZN(\SB1_1_28/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_29/Component_Function_0/N4  ( .A1(\SB1_1_29/i0[7] ), .A2(
        \SB1_1_29/i0_3 ), .A3(\SB1_1_29/i0_0 ), .ZN(
        \SB1_1_29/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_29/Component_Function_0/N3  ( .A1(\SB1_1_29/i0[10] ), .A2(
        \SB1_1_29/i0_4 ), .A3(\SB1_1_29/i0_3 ), .ZN(
        \SB1_1_29/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_29/Component_Function_0/N2  ( .A1(\SB1_1_29/i0[8] ), .A2(
        \SB1_1_29/i0[7] ), .A3(\SB1_1_29/i0[6] ), .ZN(
        \SB1_1_29/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_29/Component_Function_0/N1  ( .A1(\SB1_1_29/i0[10] ), .A2(
        \SB1_1_29/i0[9] ), .ZN(\SB1_1_29/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_29/Component_Function_1/N1  ( .A1(\SB1_1_29/i0_3 ), .A2(
        \SB1_1_29/i1[9] ), .ZN(\SB1_1_29/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_30/Component_Function_0/N1  ( .A1(\SB1_1_30/i0[10] ), .A2(
        \SB1_1_30/i0[9] ), .ZN(\SB1_1_30/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_31/Component_Function_0/N2  ( .A1(\SB1_1_31/i0[8] ), .A2(
        \SB1_1_31/i0[7] ), .A3(\SB1_1_31/i0[6] ), .ZN(
        \SB1_1_31/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_31/Component_Function_0/N1  ( .A1(\SB1_1_31/i0[10] ), .A2(
        \SB1_1_31/i0[9] ), .ZN(\SB1_1_31/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_31/Component_Function_1/N3  ( .A1(\SB1_1_31/i1_5 ), .A2(
        \SB1_1_31/i0[6] ), .A3(\SB1_1_31/i0[9] ), .ZN(
        \SB1_1_31/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_31/Component_Function_1/N2  ( .A1(\SB1_1_31/i0_3 ), .A2(
        \SB1_1_31/i1_7 ), .A3(\SB1_1_31/i0[8] ), .ZN(
        \SB1_1_31/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_0/Component_Function_0/N1  ( .A1(\SB2_1_0/i0[10] ), .A2(
        \SB2_1_0/i0[9] ), .ZN(\SB2_1_0/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_0/Component_Function_1/N2  ( .A1(\SB2_1_0/i0_3 ), .A2(
        \SB2_1_0/i1_7 ), .A3(\SB2_1_0/i0[8] ), .ZN(
        \SB2_1_0/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_1/Component_Function_0/N4  ( .A1(\SB2_1_1/i0[7] ), .A2(
        \SB2_1_1/i0_3 ), .A3(\SB2_1_1/i0_0 ), .ZN(
        \SB2_1_1/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB2_1_1/Component_Function_1/N1  ( .A1(\SB2_1_1/i0_3 ), .A2(
        \SB2_1_1/i1[9] ), .ZN(\SB2_1_1/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_2/Component_Function_0/N2  ( .A1(\SB2_1_2/i0[8] ), .A2(
        \SB2_1_2/i0[7] ), .A3(\SB2_1_2/i0[6] ), .ZN(
        \SB2_1_2/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_3/Component_Function_0/N3  ( .A1(\SB2_1_3/i0[10] ), .A2(
        n5208), .A3(\SB2_1_3/i0_3 ), .ZN(
        \SB2_1_3/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB2_1_3/Component_Function_0/N1  ( .A1(\SB2_1_3/i0[10] ), .A2(
        \SB2_1_3/i0[9] ), .ZN(\SB2_1_3/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_3/Component_Function_1/N2  ( .A1(\SB2_1_3/i0_3 ), .A2(
        \SB2_1_3/i1_7 ), .A3(\SB2_1_3/i0[8] ), .ZN(
        \SB2_1_3/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_3/Component_Function_1/N1  ( .A1(\SB2_1_3/i0_3 ), .A2(
        \SB2_1_3/i1[9] ), .ZN(\SB2_1_3/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_4/Component_Function_0/N1  ( .A1(\SB2_1_4/i0[10] ), .A2(
        \SB2_1_4/i0[9] ), .ZN(\SB2_1_4/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_4/Component_Function_1/N3  ( .A1(\SB2_1_4/i1_5 ), .A2(
        \SB2_1_4/i0[6] ), .A3(\SB1_1_9/buf_output[0] ), .ZN(
        \SB2_1_4/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_4/Component_Function_1/N2  ( .A1(\SB2_1_4/i0_3 ), .A2(
        \SB2_1_4/i1_7 ), .A3(\SB2_1_4/i0[8] ), .ZN(
        \SB2_1_4/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_5/Component_Function_0/N1  ( .A1(\SB2_1_5/i0[10] ), .A2(
        \SB2_1_5/i0[9] ), .ZN(\SB2_1_5/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_6/Component_Function_0/N2  ( .A1(\SB2_1_6/i0[8] ), .A2(
        \SB2_1_6/i0[7] ), .A3(\SB2_1_6/i0[6] ), .ZN(
        \SB2_1_6/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_6/Component_Function_0/N1  ( .A1(\SB2_1_6/i0[10] ), .A2(
        \SB2_1_6/i0[9] ), .ZN(\SB2_1_6/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_6/Component_Function_1/N4  ( .A1(\SB2_1_6/i1_7 ), .A2(
        \SB2_1_6/i0[8] ), .A3(\SB2_1_6/i0_4 ), .ZN(
        \SB2_1_6/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB2_1_6/Component_Function_1/N1  ( .A1(\SB2_1_6/i0_3 ), .A2(
        \SB2_1_6/i1[9] ), .ZN(\SB2_1_6/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_7/Component_Function_1/N2  ( .A1(\SB2_1_7/i0_3 ), .A2(
        \SB2_1_7/i1_7 ), .A3(\SB2_1_7/i0[8] ), .ZN(
        \SB2_1_7/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_7/Component_Function_5/N1  ( .A1(\SB2_1_7/i0_0 ), .A2(
        \SB2_1_7/i3[0] ), .ZN(\SB2_1_7/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_8/Component_Function_0/N4  ( .A1(\SB2_1_8/i0[7] ), .A2(
        \SB2_1_8/i0_3 ), .A3(\SB2_1_8/i0_0 ), .ZN(
        \SB2_1_8/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_8/Component_Function_0/N2  ( .A1(\SB2_1_8/i0[8] ), .A2(
        \SB2_1_8/i0[7] ), .A3(\SB2_1_8/i0[6] ), .ZN(
        \SB2_1_8/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_9/Component_Function_0/N4  ( .A1(\SB2_1_9/i0[7] ), .A2(
        \SB2_1_9/i0_3 ), .A3(\SB2_1_9/i0_0 ), .ZN(
        \SB2_1_9/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_9/Component_Function_1/N4  ( .A1(\SB2_1_9/i1_7 ), .A2(
        \SB2_1_9/i0[8] ), .A3(\SB1_1_10/buf_output[4] ), .ZN(
        \SB2_1_9/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_10/Component_Function_1/N4  ( .A1(\SB2_1_10/i1_7 ), .A2(
        \SB2_1_10/i0[8] ), .A3(\SB1_1_11/buf_output[4] ), .ZN(
        \SB2_1_10/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_10/Component_Function_1/N2  ( .A1(\SB2_1_10/i0_3 ), .A2(
        \SB2_1_10/i1_7 ), .A3(\SB2_1_10/i0[8] ), .ZN(
        \SB2_1_10/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_11/Component_Function_0/N3  ( .A1(\SB2_1_11/i0[10] ), .A2(
        \SB1_1_12/buf_output[4] ), .A3(\SB2_1_11/i0_3 ), .ZN(
        \SB2_1_11/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_11/Component_Function_1/N3  ( .A1(\SB2_1_11/i1_5 ), .A2(
        \SB2_1_11/i0[6] ), .A3(\SB2_1_11/i0[9] ), .ZN(
        \SB2_1_11/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_1_11/Component_Function_1/N1  ( .A1(\SB2_1_11/i0_3 ), .A2(
        \SB2_1_11/i1[9] ), .ZN(\SB2_1_11/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_11/Component_Function_5/N1  ( .A1(\SB2_1_11/i0_0 ), .A2(
        \SB2_1_11/i3[0] ), .ZN(\SB2_1_11/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_12/Component_Function_0/N2  ( .A1(\SB2_1_12/i0[8] ), .A2(
        \SB2_1_12/i0[7] ), .A3(\SB2_1_12/i0[6] ), .ZN(
        \SB2_1_12/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_12/Component_Function_0/N1  ( .A1(\SB2_1_12/i0[10] ), .A2(
        \SB2_1_12/i0[9] ), .ZN(\SB2_1_12/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_12/Component_Function_1/N1  ( .A1(\SB2_1_12/i0_3 ), .A2(
        \SB2_1_12/i1[9] ), .ZN(\SB2_1_12/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_13/Component_Function_5/N4  ( .A1(\SB1_1_18/buf_output[0] ), 
        .A2(\SB2_1_13/i0[6] ), .A3(\SB2_1_13/i0_4 ), .ZN(
        \SB2_1_13/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB2_1_14/Component_Function_0/N1  ( .A1(\SB2_1_14/i0[10] ), .A2(
        \SB2_1_14/i0[9] ), .ZN(\SB2_1_14/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_14/Component_Function_1/N1  ( .A1(\SB2_1_14/i0_3 ), .A2(
        \SB2_1_14/i1[9] ), .ZN(\SB2_1_14/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_15/Component_Function_1/N2  ( .A1(\SB2_1_15/i0_3 ), .A2(
        \SB2_1_15/i1_7 ), .A3(\SB2_1_15/i0[8] ), .ZN(
        \SB2_1_15/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_15/Component_Function_5/N1  ( .A1(\SB2_1_15/i0_0 ), .A2(
        \SB2_1_15/i3[0] ), .ZN(\SB2_1_15/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_16/Component_Function_0/N4  ( .A1(\SB2_1_16/i0[7] ), .A2(
        \SB2_1_16/i0_3 ), .A3(\SB2_1_16/i0_0 ), .ZN(
        \SB2_1_16/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB2_1_16/Component_Function_0/N1  ( .A1(\SB2_1_16/i0[10] ), .A2(
        \SB2_1_16/i0[9] ), .ZN(\SB2_1_16/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_16/Component_Function_1/N1  ( .A1(\SB2_1_16/i0_3 ), .A2(
        \SB2_1_16/i1[9] ), .ZN(\SB2_1_16/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_17/Component_Function_1/N1  ( .A1(\SB2_1_17/i0_3 ), .A2(
        \SB2_1_17/i1[9] ), .ZN(\SB2_1_17/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_18/Component_Function_0/N3  ( .A1(\SB2_1_18/i0[10] ), .A2(
        \SB2_1_18/i0_4 ), .A3(\SB2_1_18/i0_3 ), .ZN(
        \SB2_1_18/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB2_1_18/Component_Function_0/N1  ( .A1(\SB2_1_18/i0[10] ), .A2(
        \SB2_1_18/i0[9] ), .ZN(\SB2_1_18/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_18/Component_Function_1/N1  ( .A1(\SB2_1_18/i0_3 ), .A2(
        \SB2_1_18/i1[9] ), .ZN(\SB2_1_18/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_19/Component_Function_0/N4  ( .A1(n4149), .A2(
        \SB2_1_19/i0_3 ), .A3(\SB1_1_22/buf_output[2] ), .ZN(
        \SB2_1_19/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_19/Component_Function_1/N2  ( .A1(\SB2_1_19/i0_3 ), .A2(
        \SB2_1_19/i1_7 ), .A3(\SB2_1_19/i0[8] ), .ZN(
        \SB2_1_19/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_20/Component_Function_1/N3  ( .A1(\SB2_1_20/i1_5 ), .A2(
        \SB2_1_20/i0[6] ), .A3(\SB1_1_25/buf_output[0] ), .ZN(
        \SB2_1_20/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_21/Component_Function_0/N2  ( .A1(\SB2_1_21/i0[8] ), .A2(
        \SB2_1_21/i0[7] ), .A3(\SB2_1_21/i0[6] ), .ZN(
        \SB2_1_21/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_22/Component_Function_0/N2  ( .A1(\SB2_1_22/i0[8] ), .A2(
        \SB2_1_22/i0[7] ), .A3(\SB2_1_22/i0[6] ), .ZN(
        \SB2_1_22/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_22/Component_Function_0/N1  ( .A1(\SB2_1_22/i0[10] ), .A2(
        \SB2_1_22/i0[9] ), .ZN(\SB2_1_22/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_22/Component_Function_1/N3  ( .A1(\SB2_1_22/i1_5 ), .A2(
        \SB2_1_22/i0[6] ), .A3(\SB1_1_27/buf_output[0] ), .ZN(
        \SB2_1_22/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_1_22/Component_Function_1/N1  ( .A1(\SB2_1_22/i0_3 ), .A2(
        \SB2_1_22/i1[9] ), .ZN(\SB2_1_22/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_23/Component_Function_0/N2  ( .A1(\SB2_1_23/i0[8] ), .A2(
        \SB2_1_23/i0[7] ), .A3(\SB2_1_23/i0[6] ), .ZN(
        \SB2_1_23/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_23/Component_Function_0/N1  ( .A1(\SB2_1_23/i0[10] ), .A2(
        \SB2_1_23/i0[9] ), .ZN(\SB2_1_23/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_23/Component_Function_1/N1  ( .A1(\SB2_1_23/i0_3 ), .A2(
        \SB2_1_23/i1[9] ), .ZN(\SB2_1_23/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_24/Component_Function_0/N2  ( .A1(\SB2_1_24/i0[8] ), .A2(
        \SB2_1_24/i0[7] ), .A3(\SB2_1_24/i0[6] ), .ZN(
        \SB2_1_24/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_24/Component_Function_1/N4  ( .A1(\SB2_1_24/i1_7 ), .A2(
        \SB2_1_24/i0[8] ), .A3(\SB2_1_24/i0_4 ), .ZN(
        \SB2_1_24/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_24/Component_Function_1/N3  ( .A1(\SB2_1_24/i1_5 ), .A2(
        \SB2_1_24/i0[6] ), .A3(\SB2_1_24/i0[9] ), .ZN(
        \SB2_1_24/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_1_24/Component_Function_1/N1  ( .A1(\SB2_1_24/i0_3 ), .A2(
        \SB2_1_24/i1[9] ), .ZN(\SB2_1_24/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_25/Component_Function_0/N1  ( .A1(\SB2_1_25/i0[10] ), .A2(
        \SB2_1_25/i0[9] ), .ZN(\SB2_1_25/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_25/Component_Function_1/N2  ( .A1(\SB2_1_25/i0_3 ), .A2(
        \SB2_1_25/i1_7 ), .A3(\SB2_1_25/i0[8] ), .ZN(
        \SB2_1_25/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_25/Component_Function_1/N1  ( .A1(\SB2_1_25/i0_3 ), .A2(
        \SB2_1_25/i1[9] ), .ZN(\SB2_1_25/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_26/Component_Function_0/N1  ( .A1(\SB2_1_26/i0[10] ), .A2(
        \SB2_1_26/i0[9] ), .ZN(\SB2_1_26/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_26/Component_Function_1/N1  ( .A1(\SB2_1_26/i0_3 ), .A2(
        \SB2_1_26/i1[9] ), .ZN(\SB2_1_26/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_27/Component_Function_0/N3  ( .A1(\SB2_1_27/i0[10] ), .A2(
        \SB2_1_27/i0_4 ), .A3(\SB2_1_27/i0_3 ), .ZN(
        \SB2_1_27/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_27/Component_Function_0/N2  ( .A1(\SB2_1_27/i0[8] ), .A2(
        \SB2_1_27/i0[7] ), .A3(\SB2_1_27/i0[6] ), .ZN(
        \SB2_1_27/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_27/Component_Function_1/N2  ( .A1(\SB2_1_27/i0_3 ), .A2(
        \SB2_1_27/i1_7 ), .A3(\SB2_1_27/i0[8] ), .ZN(
        \SB2_1_27/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_27/Component_Function_1/N1  ( .A1(\SB2_1_27/i0_3 ), .A2(
        \SB2_1_27/i1[9] ), .ZN(\SB2_1_27/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_27/Component_Function_5/N1  ( .A1(\SB2_1_27/i0_0 ), .A2(
        \SB2_1_27/i3[0] ), .ZN(\SB2_1_27/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_28/Component_Function_0/N1  ( .A1(\SB2_1_28/i0[10] ), .A2(
        \SB2_1_28/i0[9] ), .ZN(\SB2_1_28/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_28/Component_Function_1/N2  ( .A1(\SB2_1_28/i0_3 ), .A2(
        \SB2_1_28/i1_7 ), .A3(\SB2_1_28/i0[8] ), .ZN(
        \SB2_1_28/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_29/Component_Function_0/N1  ( .A1(\SB2_1_29/i0[10] ), .A2(
        \SB2_1_29/i0[9] ), .ZN(\SB2_1_29/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_29/Component_Function_1/N2  ( .A1(\SB2_1_29/i0_3 ), .A2(
        \SB2_1_29/i1_7 ), .A3(\SB2_1_29/i0[8] ), .ZN(
        \SB2_1_29/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_29/Component_Function_1/N1  ( .A1(\SB2_1_29/i0_3 ), .A2(
        \SB2_1_29/i1[9] ), .ZN(\SB2_1_29/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_30/Component_Function_0/N2  ( .A1(\SB2_1_30/i0[8] ), .A2(
        n2828), .A3(\SB2_1_30/i0[6] ), .ZN(
        \SB2_1_30/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_30/Component_Function_0/N1  ( .A1(n3690), .A2(
        \SB2_1_30/i0[9] ), .ZN(\SB2_1_30/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_30/Component_Function_1/N2  ( .A1(\SB2_1_30/i0_3 ), .A2(
        \SB2_1_30/i1_7 ), .A3(\SB2_1_30/i0[8] ), .ZN(
        \SB2_1_30/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_31/Component_Function_0/N4  ( .A1(\SB2_1_31/i0[7] ), .A2(
        \SB2_1_31/i0_3 ), .A3(\SB2_1_31/i0_0 ), .ZN(
        \SB2_1_31/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB2_1_31/Component_Function_0/N1  ( .A1(\SB2_1_31/i0[10] ), .A2(
        \SB2_1_31/i0[9] ), .ZN(\SB2_1_31/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_0/Component_Function_0/N3  ( .A1(\SB1_2_0/i0[10] ), .A2(
        \SB1_2_0/i0_4 ), .A3(\SB1_2_0/i0_3 ), .ZN(
        \SB1_2_0/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_2_0/Component_Function_1/N1  ( .A1(\SB1_2_0/i0_3 ), .A2(
        \SB1_2_0/i1[9] ), .ZN(\SB1_2_0/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_2_1/Component_Function_0/N1  ( .A1(\SB1_2_1/i0[10] ), .A2(
        \SB1_2_1/i0[9] ), .ZN(\SB1_2_1/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_2_1/Component_Function_1/N1  ( .A1(\SB1_2_1/i0_3 ), .A2(
        \SB1_2_1/i1[9] ), .ZN(\SB1_2_1/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_2/Component_Function_0/N3  ( .A1(\SB1_2_2/i0[10] ), .A2(
        \SB1_2_2/i0_4 ), .A3(\SB1_2_2/i0_3 ), .ZN(
        \SB1_2_2/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_2/Component_Function_0/N2  ( .A1(\SB1_2_2/i0[8] ), .A2(
        \SB1_2_2/i0[7] ), .A3(\SB1_2_2/i0[6] ), .ZN(
        \SB1_2_2/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_2/Component_Function_1/N2  ( .A1(\SB1_2_2/i0_3 ), .A2(
        \SB1_2_2/i1_7 ), .A3(\SB1_2_2/i0[8] ), .ZN(
        \SB1_2_2/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_3/Component_Function_0/N1  ( .A1(\SB1_2_3/i0[10] ), .A2(
        \SB1_2_3/i0[9] ), .ZN(\SB1_2_3/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_3/Component_Function_1/N2  ( .A1(\SB1_2_3/i0_3 ), .A2(
        \SB1_2_3/i1_7 ), .A3(\SB1_2_3/i0[8] ), .ZN(
        \SB1_2_3/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_3/Component_Function_1/N1  ( .A1(\SB1_2_3/i0_3 ), .A2(
        \SB1_2_3/i1[9] ), .ZN(\SB1_2_3/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_4/Component_Function_0/N4  ( .A1(\SB1_2_4/i0[7] ), .A2(
        \SB1_2_4/i0_3 ), .A3(\SB1_2_4/i0_0 ), .ZN(
        \SB1_2_4/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_4/Component_Function_0/N3  ( .A1(\SB1_2_4/i0[10] ), .A2(
        \SB1_2_4/i0_4 ), .A3(\SB1_2_4/i0_3 ), .ZN(
        \SB1_2_4/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_2_4/Component_Function_0/N1  ( .A1(\SB1_2_4/i0[10] ), .A2(
        \SB1_2_4/i0[9] ), .ZN(\SB1_2_4/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_5/Component_Function_0/N4  ( .A1(\SB1_2_5/i0[7] ), .A2(
        \SB1_2_5/i0_3 ), .A3(\SB1_2_5/i0_0 ), .ZN(
        \SB1_2_5/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_5/Component_Function_0/N3  ( .A1(\SB1_2_5/i0[10] ), .A2(
        \SB1_2_5/i0_4 ), .A3(\SB1_2_5/i0_3 ), .ZN(
        \SB1_2_5/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_2_5/Component_Function_0/N1  ( .A1(\SB1_2_5/i0[10] ), .A2(
        \SB1_2_5/i0[9] ), .ZN(\SB1_2_5/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_2_5/Component_Function_1/N1  ( .A1(\SB1_2_5/i0_3 ), .A2(
        \SB1_2_5/i1[9] ), .ZN(\SB1_2_5/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_6/Component_Function_0/N3  ( .A1(\SB1_2_6/i0[10] ), .A2(
        \SB1_2_6/i0_4 ), .A3(\SB1_2_6/i0_3 ), .ZN(
        \SB1_2_6/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_2_6/Component_Function_1/N1  ( .A1(\SB1_2_6/i0_3 ), .A2(
        \SB1_2_6/i1[9] ), .ZN(\SB1_2_6/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_7/Component_Function_0/N4  ( .A1(\SB1_2_7/i0[7] ), .A2(
        \SB1_2_7/i0_3 ), .A3(\SB1_2_7/i0_0 ), .ZN(
        \SB1_2_7/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_7/Component_Function_0/N3  ( .A1(\SB1_2_7/i0[10] ), .A2(
        \SB1_2_7/i0_4 ), .A3(\SB1_2_7/i0_3 ), .ZN(
        \SB1_2_7/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_2_7/Component_Function_0/N1  ( .A1(\SB1_2_7/i0[10] ), .A2(
        \SB1_2_7/i0[9] ), .ZN(\SB1_2_7/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_7/Component_Function_1/N3  ( .A1(\SB1_2_7/i1_5 ), .A2(
        \SB1_2_7/i0[6] ), .A3(\SB1_2_7/i0[9] ), .ZN(
        \SB1_2_7/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_8/Component_Function_0/N3  ( .A1(\SB1_2_8/i0[10] ), .A2(
        \SB1_2_8/i0_4 ), .A3(\SB1_2_8/i0_3 ), .ZN(
        \SB1_2_8/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_8/Component_Function_0/N2  ( .A1(\SB1_2_8/i0[8] ), .A2(
        \SB1_2_8/i0[7] ), .A3(\SB1_2_8/i0[6] ), .ZN(
        \SB1_2_8/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_8/Component_Function_0/N1  ( .A1(\SB1_2_8/i0[10] ), .A2(
        \SB1_2_8/i0[9] ), .ZN(\SB1_2_8/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_8/Component_Function_1/N4  ( .A1(\SB1_2_8/i1_7 ), .A2(
        \SB1_2_8/i0[8] ), .A3(\SB1_2_8/i0_4 ), .ZN(
        \SB1_2_8/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB1_2_8/Component_Function_1/N1  ( .A1(\SB1_2_8/i0_3 ), .A2(
        \SB1_2_8/i1[9] ), .ZN(\SB1_2_8/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_9/Component_Function_0/N3  ( .A1(\SB1_2_9/i0[10] ), .A2(
        \SB1_2_9/i0_4 ), .A3(\SB1_2_9/i0_3 ), .ZN(
        \SB1_2_9/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_9/Component_Function_0/N2  ( .A1(\SB1_2_9/i0[8] ), .A2(
        \SB1_2_9/i0[7] ), .A3(\SB1_2_9/i0[6] ), .ZN(
        \SB1_2_9/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_9/Component_Function_0/N1  ( .A1(\SB1_2_9/i0[10] ), .A2(
        \SB1_2_9/i0[9] ), .ZN(\SB1_2_9/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_10/Component_Function_0/N3  ( .A1(\SB1_2_10/i0[10] ), .A2(
        \SB1_2_10/i0_4 ), .A3(\SB1_2_10/i0_3 ), .ZN(
        \SB1_2_10/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_10/Component_Function_0/N2  ( .A1(\SB1_2_10/i0[8] ), .A2(
        \SB1_2_10/i0[7] ), .A3(\SB1_2_10/i0[6] ), .ZN(
        \SB1_2_10/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_10/Component_Function_0/N1  ( .A1(\SB1_2_10/i0[10] ), .A2(
        \SB1_2_10/i0[9] ), .ZN(\SB1_2_10/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_2_10/Component_Function_1/N1  ( .A1(\SB1_2_10/i0_3 ), .A2(
        \SB1_2_10/i1[9] ), .ZN(\SB1_2_10/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_2_11/Component_Function_0/N1  ( .A1(\SB1_2_11/i0[10] ), .A2(
        \SB1_2_11/i0[9] ), .ZN(\SB1_2_11/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_11/Component_Function_1/N4  ( .A1(\SB1_2_11/i1_7 ), .A2(
        \SB1_2_11/i0[8] ), .A3(\SB1_2_11/i0_4 ), .ZN(
        \SB1_2_11/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB1_2_12/Component_Function_0/N1  ( .A1(\SB1_2_12/i0[10] ), .A2(
        \SB1_2_12/i0[9] ), .ZN(\SB1_2_12/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_12/Component_Function_1/N4  ( .A1(\SB1_2_12/i1_7 ), .A2(
        \SB1_2_12/i0[8] ), .A3(\SB1_2_12/i0_4 ), .ZN(
        \SB1_2_12/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_13/Component_Function_0/N3  ( .A1(\SB1_2_13/i0[10] ), .A2(
        \MC_ARK_ARC_1_1/buf_output[112] ), .A3(n5526), .ZN(
        \SB1_2_13/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_13/Component_Function_1/N2  ( .A1(\SB1_2_13/i0_3 ), .A2(
        \SB1_2_13/i1_7 ), .A3(\SB1_2_13/i0[8] ), .ZN(
        \SB1_2_13/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_13/Component_Function_1/N1  ( .A1(\SB1_2_13/i0_3 ), .A2(
        \SB1_2_13/i1[9] ), .ZN(\SB1_2_13/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_14/Component_Function_0/N3  ( .A1(\SB1_2_14/i0[10] ), .A2(
        \SB1_2_14/i0_4 ), .A3(\SB1_2_14/i0_3 ), .ZN(
        \SB1_2_14/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_14/Component_Function_0/N2  ( .A1(\SB1_2_14/i0[8] ), .A2(
        \SB1_2_14/i0[7] ), .A3(\SB1_2_14/i0[6] ), .ZN(
        \SB1_2_14/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_14/Component_Function_1/N1  ( .A1(\SB1_2_14/i0_3 ), .A2(
        \SB1_2_14/i1[9] ), .ZN(\SB1_2_14/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_2_15/Component_Function_0/N1  ( .A1(\SB1_2_15/i0[10] ), .A2(
        \SB1_2_15/i0[9] ), .ZN(\SB1_2_15/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_17/Component_Function_0/N2  ( .A1(\SB1_2_17/i0[8] ), .A2(
        \SB1_2_17/i0[7] ), .A3(\SB1_2_17/i0[6] ), .ZN(
        \SB1_2_17/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_17/Component_Function_0/N1  ( .A1(\SB1_2_17/i0[10] ), .A2(
        \SB1_2_17/i0[9] ), .ZN(\SB1_2_17/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_17/Component_Function_1/N2  ( .A1(\SB1_2_17/i0_3 ), .A2(
        \SB1_2_17/i1_7 ), .A3(\SB1_2_17/i0[8] ), .ZN(
        \SB1_2_17/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_18/Component_Function_0/N2  ( .A1(n4762), .A2(
        \SB1_2_18/i0[7] ), .A3(\SB1_2_18/i0[6] ), .ZN(
        \SB1_2_18/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_18/Component_Function_0/N1  ( .A1(\SB1_2_18/i0[10] ), .A2(
        \SB1_2_18/i0[9] ), .ZN(\SB1_2_18/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_18/Component_Function_1/N2  ( .A1(\SB1_2_18/i0_3 ), .A2(
        \SB1_2_18/i1_7 ), .A3(n4762), .ZN(
        \SB1_2_18/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_18/Component_Function_1/N1  ( .A1(\SB1_2_18/i0_3 ), .A2(
        \SB1_2_18/i1[9] ), .ZN(\SB1_2_18/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_19/Component_Function_0/N4  ( .A1(\SB1_2_19/i0[7] ), .A2(
        \SB1_2_19/i0_3 ), .A3(\SB1_2_19/i0_0 ), .ZN(
        \SB1_2_19/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_19/Component_Function_0/N3  ( .A1(\SB1_2_19/i0[10] ), .A2(
        \MC_ARK_ARC_1_1/buf_output[76] ), .A3(\SB1_2_19/i0_3 ), .ZN(
        \SB1_2_19/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_19/Component_Function_0/N2  ( .A1(\SB1_2_19/i0[8] ), .A2(
        \SB1_2_19/i0[7] ), .A3(\SB1_2_19/i0[6] ), .ZN(
        \SB1_2_19/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_19/Component_Function_0/N1  ( .A1(\SB1_2_19/i0[10] ), .A2(
        \SB1_2_19/i0[9] ), .ZN(\SB1_2_19/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_20/Component_Function_0/N3  ( .A1(\SB1_2_20/i0[10] ), .A2(
        \SB1_2_20/i0_4 ), .A3(\SB1_2_20/i0_3 ), .ZN(
        \SB1_2_20/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_2_20/Component_Function_0/N1  ( .A1(\SB1_2_20/i0[10] ), .A2(
        \SB1_2_20/i0[9] ), .ZN(\SB1_2_20/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_20/Component_Function_1/N4  ( .A1(\SB1_2_20/i1_7 ), .A2(
        n2893), .A3(\SB1_2_20/i0_4 ), .ZN(
        \SB1_2_20/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_20/Component_Function_1/N2  ( .A1(\SB1_2_20/i0_3 ), .A2(
        \SB1_2_20/i1_7 ), .A3(n2893), .ZN(
        \SB1_2_20/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_21/Component_Function_0/N3  ( .A1(\SB1_2_21/i0[10] ), .A2(
        \SB1_2_21/i0_4 ), .A3(\SB1_2_21/i0_3 ), .ZN(
        \SB1_2_21/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_21/Component_Function_0/N2  ( .A1(\SB1_2_21/i0[8] ), .A2(
        \SB1_2_21/i0[7] ), .A3(\SB1_2_21/i0[6] ), .ZN(
        \SB1_2_21/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_21/Component_Function_0/N1  ( .A1(\SB1_2_21/i0[10] ), .A2(
        \SB1_2_21/i0[9] ), .ZN(\SB1_2_21/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_22/Component_Function_0/N4  ( .A1(\SB1_2_22/i0[7] ), .A2(
        \SB1_2_22/i0_3 ), .A3(\SB1_2_22/i0_0 ), .ZN(
        \SB1_2_22/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB1_2_22/Component_Function_0/N1  ( .A1(\SB1_2_22/i0[10] ), .A2(
        \SB1_2_22/i0[9] ), .ZN(\SB1_2_22/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_22/Component_Function_1/N3  ( .A1(\SB1_2_22/i1_5 ), .A2(
        \SB1_2_22/i0[6] ), .A3(\SB1_2_22/i0[9] ), .ZN(
        \SB1_2_22/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_22/Component_Function_1/N2  ( .A1(\SB1_2_22/i0_3 ), .A2(
        \SB1_2_22/i1_7 ), .A3(\SB1_2_22/i0[8] ), .ZN(
        \SB1_2_22/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_23/Component_Function_0/N2  ( .A1(\SB1_2_23/i0[8] ), .A2(
        \SB1_2_23/i0[7] ), .A3(\SB1_2_23/i0[6] ), .ZN(
        \SB1_2_23/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_23/Component_Function_0/N1  ( .A1(\SB1_2_23/i0[10] ), .A2(
        \SB1_2_23/i0[9] ), .ZN(\SB1_2_23/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_23/Component_Function_1/N2  ( .A1(\SB1_2_23/i0_3 ), .A2(
        \SB1_2_23/i1_7 ), .A3(\SB1_2_23/i0[8] ), .ZN(
        \SB1_2_23/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_24/Component_Function_0/N1  ( .A1(\SB1_2_24/i0[10] ), .A2(
        \SB1_2_24/i0[9] ), .ZN(\SB1_2_24/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_24/Component_Function_1/N4  ( .A1(\SB1_2_24/i1_7 ), .A2(
        \SB1_2_24/i0[8] ), .A3(\SB1_2_24/i0_4 ), .ZN(
        \SB1_2_24/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_25/Component_Function_0/N2  ( .A1(\SB1_2_25/i0[8] ), .A2(
        \SB1_2_25/i0[7] ), .A3(\SB1_2_25/i0[6] ), .ZN(
        \SB1_2_25/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_25/Component_Function_0/N1  ( .A1(\SB1_2_25/i0[10] ), .A2(
        \SB1_2_25/i0[9] ), .ZN(\SB1_2_25/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_27/Component_Function_0/N2  ( .A1(\SB1_2_27/i0[8] ), .A2(
        \SB1_2_27/i0[7] ), .A3(\SB1_2_27/i0[6] ), .ZN(
        \SB1_2_27/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_27/Component_Function_0/N1  ( .A1(\SB1_2_27/i0[10] ), .A2(
        \SB1_2_27/i0[9] ), .ZN(\SB1_2_27/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_27/Component_Function_1/N4  ( .A1(\SB1_2_27/i1_7 ), .A2(
        \SB1_2_27/i0[8] ), .A3(\SB1_2_27/i0_4 ), .ZN(
        \SB1_2_27/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_27/Component_Function_1/N2  ( .A1(\SB1_2_27/i0_3 ), .A2(
        \SB1_2_27/i1_7 ), .A3(\SB1_2_27/i0[8] ), .ZN(
        \SB1_2_27/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_27/Component_Function_1/N1  ( .A1(\SB1_2_27/i0_3 ), .A2(
        \SB1_2_27/i1[9] ), .ZN(\SB1_2_27/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_28/Component_Function_0/N4  ( .A1(\SB1_2_28/i0[7] ), .A2(
        \SB1_2_28/i0_3 ), .A3(\SB1_2_28/i0_0 ), .ZN(
        \SB1_2_28/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_28/Component_Function_0/N3  ( .A1(\SB1_2_28/i0[10] ), .A2(
        \SB1_2_28/i0_4 ), .A3(\SB1_2_28/i0_3 ), .ZN(
        \SB1_2_28/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_28/Component_Function_0/N2  ( .A1(\SB1_2_28/i0[8] ), .A2(
        \SB1_2_28/i0[7] ), .A3(\SB1_2_28/i0[6] ), .ZN(
        \SB1_2_28/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_28/Component_Function_0/N1  ( .A1(\SB1_2_28/i0[10] ), .A2(
        \SB1_2_28/i0[9] ), .ZN(\SB1_2_28/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_2_28/Component_Function_1/N1  ( .A1(\SB1_2_28/i0_3 ), .A2(
        \SB1_2_28/i1[9] ), .ZN(\SB1_2_28/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_29/Component_Function_0/N2  ( .A1(\SB1_2_29/i0[8] ), .A2(
        \SB1_2_29/i0[7] ), .A3(\SB1_2_29/i0[6] ), .ZN(
        \SB1_2_29/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_29/Component_Function_0/N1  ( .A1(\SB1_2_29/i0[10] ), .A2(
        \SB1_2_29/i0[9] ), .ZN(\SB1_2_29/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_2_29/Component_Function_1/N1  ( .A1(\RI1[2][17] ), .A2(
        \SB1_2_29/i1[9] ), .ZN(\SB1_2_29/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_30/Component_Function_0/N2  ( .A1(\SB1_2_30/i0[8] ), .A2(
        \SB1_2_30/i0[7] ), .A3(\SB1_2_30/i0[6] ), .ZN(
        \SB1_2_30/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_30/Component_Function_0/N1  ( .A1(\SB1_2_30/i0[10] ), .A2(
        \SB1_2_30/i0[9] ), .ZN(\SB1_2_30/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_2_30/Component_Function_1/N1  ( .A1(\SB1_2_30/i0_3 ), .A2(
        \SB1_2_30/i1[9] ), .ZN(\SB1_2_30/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_31/Component_Function_0/N2  ( .A1(\SB1_2_31/i0[8] ), .A2(
        \SB1_2_31/i0[7] ), .A3(\SB1_2_31/i0[6] ), .ZN(
        \SB1_2_31/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_31/Component_Function_0/N1  ( .A1(\SB1_2_31/i0[10] ), .A2(
        \SB1_2_31/i0[9] ), .ZN(\SB1_2_31/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_31/Component_Function_1/N2  ( .A1(\SB1_2_31/i0_3 ), .A2(
        \SB1_2_31/i1_7 ), .A3(\SB1_2_31/i0[8] ), .ZN(
        \SB1_2_31/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_31/Component_Function_1/N1  ( .A1(\SB1_2_31/i0_3 ), .A2(
        \SB1_2_31/i1[9] ), .ZN(\SB1_2_31/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_0/Component_Function_0/N2  ( .A1(\SB2_2_0/i0[8] ), .A2(
        \SB2_2_0/i0[7] ), .A3(\SB2_2_0/i0[6] ), .ZN(
        \SB2_2_0/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_0/Component_Function_0/N1  ( .A1(\SB2_2_0/i0[10] ), .A2(
        \SB2_2_0/i0[9] ), .ZN(\SB2_2_0/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_0/Component_Function_1/N3  ( .A1(\SB2_2_0/i1_5 ), .A2(
        \SB2_2_0/i0[6] ), .A3(\SB2_2_0/i0[9] ), .ZN(
        \SB2_2_0/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_2_1/Component_Function_0/N1  ( .A1(\SB2_2_1/i0[10] ), .A2(
        \SB2_2_1/i0[9] ), .ZN(\SB2_2_1/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_2/Component_Function_0/N4  ( .A1(\SB2_2_2/i0[7] ), .A2(
        \SB2_2_2/i0_3 ), .A3(\SB2_2_2/i0_0 ), .ZN(
        \SB2_2_2/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB2_2_2/Component_Function_0/N1  ( .A1(\SB2_2_2/i0[10] ), .A2(
        \SB2_2_2/i0[9] ), .ZN(\SB2_2_2/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_2/Component_Function_1/N4  ( .A1(\SB2_2_2/i1_7 ), .A2(
        \SB2_2_2/i0[8] ), .A3(\SB2_2_2/i0_4 ), .ZN(
        \SB2_2_2/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_2/Component_Function_1/N3  ( .A1(\SB2_2_2/i1_5 ), .A2(
        \SB2_2_2/i0[6] ), .A3(\SB2_2_2/i0[9] ), .ZN(
        \SB2_2_2/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_3/Component_Function_0/N2  ( .A1(\SB2_2_3/i0[8] ), .A2(n5886), .A3(\SB2_2_3/i0[6] ), .ZN(\SB2_2_3/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_3/Component_Function_0/N1  ( .A1(\SB2_2_3/i0[10] ), .A2(
        \SB2_2_3/i0[9] ), .ZN(\SB2_2_3/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_3/Component_Function_1/N1  ( .A1(\SB2_2_3/i0_3 ), .A2(
        \SB2_2_3/i1[9] ), .ZN(\SB2_2_3/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_4/Component_Function_0/N1  ( .A1(\SB2_2_4/i0[10] ), .A2(
        \SB2_2_4/i0[9] ), .ZN(\SB2_2_4/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_4/Component_Function_1/N1  ( .A1(\SB2_2_4/i0_3 ), .A2(
        \SB2_2_4/i1[9] ), .ZN(\SB2_2_4/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_4/Component_Function_5/N1  ( .A1(\SB2_2_4/i0_0 ), .A2(
        \SB2_2_4/i3[0] ), .ZN(\SB2_2_4/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_5/Component_Function_0/N1  ( .A1(\SB2_2_5/i0[10] ), .A2(
        \SB2_2_5/i0[9] ), .ZN(\SB2_2_5/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_6/Component_Function_0/N2  ( .A1(\SB2_2_6/i0[8] ), .A2(
        \SB2_2_6/i0[7] ), .A3(\SB2_2_6/i0[6] ), .ZN(
        \SB2_2_6/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_6/Component_Function_0/N1  ( .A1(\SB2_2_6/i0[10] ), .A2(
        \SB2_2_6/i0[9] ), .ZN(\SB2_2_6/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_6/Component_Function_1/N3  ( .A1(\SB2_2_6/i1_5 ), .A2(
        \SB2_2_6/i0[6] ), .A3(\SB2_2_6/i0[9] ), .ZN(
        \SB2_2_6/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_2_6/Component_Function_1/N1  ( .A1(\SB2_2_6/i0_3 ), .A2(
        \SB2_2_6/i1[9] ), .ZN(\SB2_2_6/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_7/Component_Function_0/N3  ( .A1(\SB2_2_7/i0[10] ), .A2(
        \SB1_2_8/buf_output[4] ), .A3(\SB2_2_7/i0_3 ), .ZN(
        \SB2_2_7/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB2_2_7/Component_Function_0/N1  ( .A1(\SB2_2_7/i0[10] ), .A2(
        \SB2_2_7/i0[9] ), .ZN(\SB2_2_7/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_7/Component_Function_1/N4  ( .A1(\SB2_2_7/i1_7 ), .A2(
        \SB2_2_7/i0[8] ), .A3(\SB1_2_8/buf_output[4] ), .ZN(
        \SB2_2_7/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_7/Component_Function_1/N2  ( .A1(\SB2_2_7/i0_3 ), .A2(
        \SB2_2_7/i1_7 ), .A3(\SB2_2_7/i0[8] ), .ZN(
        \SB2_2_7/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_8/Component_Function_1/N1  ( .A1(\SB2_2_8/i0_3 ), .A2(
        \SB2_2_8/i1[9] ), .ZN(\SB2_2_8/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_9/Component_Function_0/N1  ( .A1(\SB2_2_9/i0[10] ), .A2(
        \SB2_2_9/i0[9] ), .ZN(\SB2_2_9/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_10/Component_Function_0/N1  ( .A1(\SB2_2_10/i0[10] ), .A2(
        \SB2_2_10/i0[9] ), .ZN(\SB2_2_10/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_10/Component_Function_1/N3  ( .A1(\SB2_2_10/i1_5 ), .A2(
        \SB2_2_10/i0[6] ), .A3(\SB2_2_10/i0[9] ), .ZN(
        \SB2_2_10/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_10/Component_Function_1/N2  ( .A1(\SB2_2_10/i0_3 ), .A2(
        \SB2_2_10/i1_7 ), .A3(\SB2_2_10/i0[8] ), .ZN(
        \SB2_2_10/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_10/Component_Function_1/N1  ( .A1(\SB2_2_10/i0_3 ), .A2(
        \SB2_2_10/i1[9] ), .ZN(\SB2_2_10/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_11/Component_Function_0/N2  ( .A1(\SB2_2_11/i0[8] ), .A2(
        \SB2_2_11/i0[7] ), .A3(\SB2_2_11/i0[6] ), .ZN(
        \SB2_2_11/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_11/Component_Function_0/N1  ( .A1(n5826), .A2(
        \SB2_2_11/i0[9] ), .ZN(\SB2_2_11/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_11/Component_Function_1/N1  ( .A1(\SB2_2_11/i0_3 ), .A2(
        n5515), .ZN(\SB2_2_11/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_12/Component_Function_0/N4  ( .A1(\SB2_2_12/i0[7] ), .A2(
        \SB2_2_12/i0_3 ), .A3(\SB2_2_12/i0_0 ), .ZN(
        \SB2_2_12/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_12/Component_Function_0/N3  ( .A1(\SB2_2_12/i0[10] ), .A2(
        \SB2_2_12/i0_4 ), .A3(\SB2_2_12/i0_3 ), .ZN(
        \SB2_2_12/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_12/Component_Function_0/N2  ( .A1(\SB2_2_12/i0[8] ), .A2(
        \SB2_2_12/i0[7] ), .A3(\SB2_2_12/i0[6] ), .ZN(
        \SB2_2_12/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_12/Component_Function_0/N1  ( .A1(\SB2_2_12/i0[10] ), .A2(
        \SB2_2_12/i0[9] ), .ZN(\SB2_2_12/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_13/Component_Function_0/N1  ( .A1(\SB2_2_13/i0[10] ), .A2(
        \SB2_2_13/i0[9] ), .ZN(\SB2_2_13/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_13/Component_Function_1/N2  ( .A1(\SB2_2_13/i0_3 ), .A2(
        \SB2_2_13/i1_7 ), .A3(\SB2_2_13/i0[8] ), .ZN(
        \SB2_2_13/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_14/Component_Function_0/N3  ( .A1(\SB2_2_14/i0[10] ), .A2(
        n5932), .A3(\SB2_2_14/i0_3 ), .ZN(
        \SB2_2_14/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB2_2_14/Component_Function_0/N1  ( .A1(\SB2_2_14/i0[10] ), .A2(
        \SB2_2_14/i0[9] ), .ZN(\SB2_2_14/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_14/Component_Function_1/N2  ( .A1(\SB2_2_14/i0_3 ), .A2(
        \SB2_2_14/i1_7 ), .A3(\SB2_2_14/i0[8] ), .ZN(
        \SB2_2_14/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_15/Component_Function_0/N1  ( .A1(\SB2_2_15/i0[10] ), .A2(
        \SB2_2_15/i0[9] ), .ZN(\SB2_2_15/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_15/Component_Function_1/N1  ( .A1(\SB2_2_15/i0_3 ), .A2(
        \SB2_2_15/i1[9] ), .ZN(\SB2_2_15/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_16/Component_Function_0/N2  ( .A1(\SB2_2_16/i0[8] ), .A2(
        \SB2_2_16/i0[7] ), .A3(\SB2_2_16/i0[6] ), .ZN(
        \SB2_2_16/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_16/Component_Function_0/N1  ( .A1(\SB2_2_16/i0[10] ), .A2(
        \SB2_2_16/i0[9] ), .ZN(\SB2_2_16/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_16/Component_Function_1/N3  ( .A1(\SB2_2_16/i1_5 ), .A2(
        \SB2_2_16/i0[6] ), .A3(\SB2_2_16/i0[9] ), .ZN(
        \SB2_2_16/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_17/Component_Function_0/N4  ( .A1(\SB2_2_17/i0[7] ), .A2(
        \SB2_2_17/i0_3 ), .A3(\SB2_2_17/i0_0 ), .ZN(
        \SB2_2_17/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB2_2_17/Component_Function_0/N1  ( .A1(\SB2_2_17/i0[10] ), .A2(
        \SB2_2_17/i0[9] ), .ZN(\SB2_2_17/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_17/Component_Function_1/N2  ( .A1(\SB1_2_17/buf_output[5] ), 
        .A2(\SB2_2_17/i1_7 ), .A3(\SB2_2_17/i0[8] ), .ZN(
        \SB2_2_17/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_18/Component_Function_0/N3  ( .A1(\SB2_2_18/i0[10] ), .A2(
        \SB2_2_18/i0_4 ), .A3(\SB2_2_18/i0_3 ), .ZN(
        \SB2_2_18/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB2_2_18/Component_Function_0/N1  ( .A1(\SB2_2_18/i0[10] ), .A2(
        \SB2_2_18/i0[9] ), .ZN(\SB2_2_18/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_18/Component_Function_1/N1  ( .A1(\SB2_2_18/i0_3 ), .A2(
        \SB2_2_18/i1[9] ), .ZN(\SB2_2_18/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_19/Component_Function_0/N2  ( .A1(\SB2_2_19/i0[8] ), .A2(
        \SB2_2_19/i0[7] ), .A3(\SB2_2_19/i0[6] ), .ZN(
        \SB2_2_19/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_19/Component_Function_1/N2  ( .A1(\SB2_2_19/i0_3 ), .A2(
        \SB2_2_19/i1_7 ), .A3(\SB2_2_19/i0[8] ), .ZN(
        \SB2_2_19/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_20/Component_Function_0/N3  ( .A1(\SB2_2_20/i0[10] ), .A2(
        \SB2_2_20/i0_4 ), .A3(\SB2_2_20/i0_3 ), .ZN(
        \SB2_2_20/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_20/Component_Function_0/N2  ( .A1(\SB2_2_20/i0[8] ), .A2(
        \SB2_2_20/i0[7] ), .A3(\SB2_2_20/i0[6] ), .ZN(
        \SB2_2_20/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_20/Component_Function_0/N1  ( .A1(\SB2_2_20/i0[10] ), .A2(
        \SB2_2_20/i0[9] ), .ZN(\SB2_2_20/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_20/Component_Function_1/N1  ( .A1(\SB2_2_20/i0_3 ), .A2(
        \SB2_2_20/i1[9] ), .ZN(\SB2_2_20/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_21/Component_Function_1/N1  ( .A1(\SB2_2_21/i0_3 ), .A2(
        \SB2_2_21/i1[9] ), .ZN(\SB2_2_21/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_22/Component_Function_0/N2  ( .A1(\SB2_2_22/i0[8] ), .A2(
        \SB2_2_22/i0[7] ), .A3(\SB2_2_22/i0[6] ), .ZN(
        \SB2_2_22/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_23/Component_Function_0/N2  ( .A1(\SB2_2_23/i0[8] ), .A2(
        \SB2_2_23/i0[7] ), .A3(\SB2_2_23/i0[6] ), .ZN(
        \SB2_2_23/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_23/Component_Function_1/N3  ( .A1(\SB2_2_23/i1_5 ), .A2(
        \SB2_2_23/i0[6] ), .A3(\SB2_2_23/i0[9] ), .ZN(
        \SB2_2_23/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_24/Component_Function_0/N2  ( .A1(\SB2_2_24/i0[8] ), .A2(
        \SB2_2_24/i0[7] ), .A3(\SB2_2_24/i0[6] ), .ZN(
        \SB2_2_24/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_24/Component_Function_0/N1  ( .A1(\SB2_2_24/i0[10] ), .A2(
        \SB2_2_24/i0[9] ), .ZN(\SB2_2_24/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_24/Component_Function_1/N1  ( .A1(\SB2_2_24/i0_3 ), .A2(
        \SB2_2_24/i1[9] ), .ZN(\SB2_2_24/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_25/Component_Function_0/N1  ( .A1(\SB2_2_25/i0[10] ), .A2(
        \SB2_2_25/i0[9] ), .ZN(\SB2_2_25/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_25/Component_Function_1/N4  ( .A1(\SB2_2_25/i1_7 ), .A2(
        \SB2_2_25/i0[8] ), .A3(\SB1_2_26/buf_output[4] ), .ZN(
        \SB2_2_25/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB2_2_26/Component_Function_0/N1  ( .A1(\SB2_2_26/i0[10] ), .A2(
        \SB2_2_26/i0[9] ), .ZN(\SB2_2_26/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_26/Component_Function_1/N4  ( .A1(\SB2_2_26/i1_7 ), .A2(
        \SB2_2_26/i0[8] ), .A3(\SB2_2_26/i0_4 ), .ZN(
        \SB2_2_26/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB2_2_26/Component_Function_1/N1  ( .A1(\SB2_2_26/i0_3 ), .A2(
        \SB2_2_26/i1[9] ), .ZN(\SB2_2_26/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_27/Component_Function_0/N4  ( .A1(n6073), .A2(
        \SB2_2_27/i0_3 ), .A3(\SB2_2_27/i0_0 ), .ZN(
        \SB2_2_27/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB2_2_27/Component_Function_0/N1  ( .A1(\SB2_2_27/i0[10] ), .A2(
        \SB1_2_0/buf_output[0] ), .ZN(
        \SB2_2_27/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_27/Component_Function_1/N1  ( .A1(\SB2_2_27/i0_3 ), .A2(
        \SB2_2_27/i1[9] ), .ZN(\SB2_2_27/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_28/Component_Function_0/N4  ( .A1(\SB2_2_28/i0[7] ), .A2(
        \SB2_2_28/i0_3 ), .A3(\SB2_2_28/i0_0 ), .ZN(
        \SB2_2_28/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_28/Component_Function_1/N2  ( .A1(\SB2_2_28/i0_3 ), .A2(
        \SB2_2_28/i1_7 ), .A3(\SB2_2_28/i0[8] ), .ZN(
        \SB2_2_28/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_28/Component_Function_1/N1  ( .A1(\SB2_2_28/i0_3 ), .A2(
        \SB2_2_28/i1[9] ), .ZN(\SB2_2_28/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_28/Component_Function_5/N4  ( .A1(\SB1_2_1/buf_output[0] ), 
        .A2(\SB2_2_28/i0[6] ), .A3(\SB2_2_28/i0_4 ), .ZN(
        \SB2_2_28/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB2_2_29/Component_Function_0/N1  ( .A1(\SB2_2_29/i0[10] ), .A2(
        \SB2_2_29/i0[9] ), .ZN(\SB2_2_29/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_29/Component_Function_1/N1  ( .A1(\SB2_2_29/i0_3 ), .A2(
        \SB2_2_29/i1[9] ), .ZN(\SB2_2_29/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_30/Component_Function_0/N2  ( .A1(\SB2_2_30/i0[8] ), .A2(
        \SB2_2_30/i0[7] ), .A3(\SB2_2_30/i0[6] ), .ZN(
        \SB2_2_30/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_30/Component_Function_0/N1  ( .A1(\SB2_2_30/i0[10] ), .A2(
        \SB2_2_30/i0[9] ), .ZN(\SB2_2_30/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_30/Component_Function_1/N3  ( .A1(\SB2_2_30/i1_5 ), .A2(
        \SB2_2_30/i0[6] ), .A3(\SB2_2_30/i0[9] ), .ZN(
        \SB2_2_30/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_30/Component_Function_1/N2  ( .A1(\SB2_2_30/i0_3 ), .A2(
        \SB2_2_30/i1_7 ), .A3(\SB2_2_30/i0[8] ), .ZN(
        \SB2_2_30/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_31/Component_Function_0/N1  ( .A1(\SB2_2_31/i0[10] ), .A2(
        \SB2_2_31/i0[9] ), .ZN(\SB2_2_31/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_0/Component_Function_0/N3  ( .A1(\SB1_3_0/i0[10] ), .A2(
        \SB1_3_0/i0_4 ), .A3(\SB1_3_0/i0_3 ), .ZN(
        \SB1_3_0/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_0/Component_Function_0/N2  ( .A1(\SB1_3_0/i0[8] ), .A2(
        \SB1_3_0/i0[7] ), .A3(\SB1_3_0/i0[6] ), .ZN(
        \SB1_3_0/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_0/Component_Function_0/N1  ( .A1(\SB1_3_0/i0[10] ), .A2(
        \SB1_3_0/i0[9] ), .ZN(\SB1_3_0/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_0/Component_Function_1/N3  ( .A1(\SB1_3_0/i1_5 ), .A2(
        \SB1_3_0/i0[6] ), .A3(\SB1_3_0/i0[9] ), .ZN(
        \SB1_3_0/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_0/Component_Function_1/N2  ( .A1(\SB1_3_0/i0_3 ), .A2(
        \SB1_3_0/i1_7 ), .A3(\SB1_3_0/i0[8] ), .ZN(
        \SB1_3_0/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_1/Component_Function_0/N2  ( .A1(\SB1_3_1/i0[8] ), .A2(
        \SB1_3_1/i0[7] ), .A3(\SB1_3_1/i0[6] ), .ZN(
        \SB1_3_1/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_1/Component_Function_0/N1  ( .A1(\SB1_3_1/i0[10] ), .A2(
        \SB1_3_1/i0[9] ), .ZN(\SB1_3_1/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_1/Component_Function_1/N2  ( .A1(\SB1_3_1/i0_3 ), .A2(
        \SB1_3_1/i1_7 ), .A3(\SB1_3_1/i0[8] ), .ZN(
        \SB1_3_1/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_1/Component_Function_1/N1  ( .A1(\SB1_3_1/i0_3 ), .A2(
        \SB1_3_1/i1[9] ), .ZN(\SB1_3_1/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_2/Component_Function_0/N3  ( .A1(\SB1_3_2/i0[10] ), .A2(
        \SB1_3_2/i0_4 ), .A3(\SB1_3_2/i0_3 ), .ZN(
        \SB1_3_2/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_3_2/Component_Function_0/N1  ( .A1(\SB1_3_2/i0[10] ), .A2(
        \SB1_3_2/i0[9] ), .ZN(\SB1_3_2/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_3_2/Component_Function_1/N1  ( .A1(\SB1_3_2/i0_3 ), .A2(
        \SB1_3_2/i1[9] ), .ZN(\SB1_3_2/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_3/Component_Function_0/N4  ( .A1(\SB1_3_3/i0[7] ), .A2(
        \SB1_3_3/i0_3 ), .A3(\SB1_3_3/i0_0 ), .ZN(
        \SB1_3_3/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_3/Component_Function_0/N3  ( .A1(\SB1_3_3/i0[10] ), .A2(
        \SB1_3_3/i0_4 ), .A3(\SB1_3_3/i0_3 ), .ZN(
        \SB1_3_3/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_3_3/Component_Function_0/N1  ( .A1(\SB1_3_3/i0[10] ), .A2(
        \SB1_3_3/i0[9] ), .ZN(\SB1_3_3/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_3/Component_Function_1/N2  ( .A1(\SB1_3_3/i0_3 ), .A2(
        \SB1_3_3/i1_7 ), .A3(\SB1_3_3/i0[8] ), .ZN(
        \SB1_3_3/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_4/Component_Function_0/N1  ( .A1(\SB1_3_4/i0[10] ), .A2(
        \SB1_3_4/i0[9] ), .ZN(\SB1_3_4/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_5/Component_Function_0/N4  ( .A1(\SB1_3_5/i0[7] ), .A2(
        \SB1_3_5/i0_3 ), .A3(\SB1_3_5/i0_0 ), .ZN(
        \SB1_3_5/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_5/Component_Function_0/N3  ( .A1(\SB1_3_5/i0[10] ), .A2(
        \SB1_3_5/i0_4 ), .A3(\SB1_3_5/i0_3 ), .ZN(
        \SB1_3_5/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_5/Component_Function_0/N2  ( .A1(\SB1_3_5/i0[8] ), .A2(
        \SB1_3_5/i0[7] ), .A3(\SB1_3_5/i0[6] ), .ZN(
        \SB1_3_5/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_5/Component_Function_0/N1  ( .A1(\SB1_3_5/i0[10] ), .A2(
        \SB1_3_5/i0[9] ), .ZN(\SB1_3_5/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_3_5/Component_Function_1/N1  ( .A1(\SB1_3_5/i0_3 ), .A2(
        \SB1_3_5/i1[9] ), .ZN(\SB1_3_5/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_6/Component_Function_0/N3  ( .A1(\SB1_3_6/i0[10] ), .A2(
        \SB1_3_6/i0_4 ), .A3(\SB1_3_6/i0_3 ), .ZN(
        \SB1_3_6/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_6/Component_Function_0/N2  ( .A1(\SB1_3_6/i0[8] ), .A2(
        \SB1_3_6/i0[7] ), .A3(\SB1_3_6/i0[6] ), .ZN(
        \SB1_3_6/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_6/Component_Function_0/N1  ( .A1(\SB1_3_6/i0[10] ), .A2(
        \SB1_3_6/i0[9] ), .ZN(\SB1_3_6/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_6/Component_Function_1/N4  ( .A1(\SB1_3_6/i1_7 ), .A2(
        \SB1_3_6/i0[8] ), .A3(\SB1_3_6/i0_4 ), .ZN(
        \SB1_3_6/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_6/Component_Function_1/N2  ( .A1(\SB1_3_6/i0_3 ), .A2(
        \SB1_3_6/i1_7 ), .A3(\SB1_3_6/i0[8] ), .ZN(
        \SB1_3_6/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_7/Component_Function_0/N2  ( .A1(\SB1_3_7/i0[8] ), .A2(
        \SB1_3_7/i0[7] ), .A3(\SB1_3_7/i0[6] ), .ZN(
        \SB1_3_7/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_7/Component_Function_0/N1  ( .A1(\SB1_3_7/i0[10] ), .A2(
        \SB1_3_7/i0[9] ), .ZN(\SB1_3_7/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_3_8/Component_Function_0/N1  ( .A1(\SB1_3_8/i0[10] ), .A2(
        \SB1_3_8/i0[9] ), .ZN(\SB1_3_8/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_9/Component_Function_0/N4  ( .A1(\SB1_3_9/i0[7] ), .A2(
        \SB1_3_9/i0_3 ), .A3(\SB1_3_9/i0_0 ), .ZN(
        \SB1_3_9/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB1_3_9/Component_Function_1/N1  ( .A1(\SB1_3_9/i0_3 ), .A2(
        \SB1_3_9/i1[9] ), .ZN(\SB1_3_9/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_10/Component_Function_0/N2  ( .A1(\SB1_3_10/i0[8] ), .A2(
        \SB1_3_10/i0[7] ), .A3(\SB1_3_10/i0[6] ), .ZN(
        \SB1_3_10/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_11/Component_Function_0/N3  ( .A1(\SB1_3_11/i0[10] ), .A2(
        \SB1_3_11/i0_4 ), .A3(\SB1_3_11/i0_3 ), .ZN(
        \SB1_3_11/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_11/Component_Function_0/N2  ( .A1(\SB1_3_11/i0[8] ), .A2(
        n3648), .A3(\SB1_3_11/i0[6] ), .ZN(
        \SB1_3_11/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_13/Component_Function_0/N3  ( .A1(\SB1_3_13/i0[10] ), .A2(
        \SB1_3_13/i0_4 ), .A3(\SB1_3_13/i0_3 ), .ZN(
        \SB1_3_13/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_13/Component_Function_0/N2  ( .A1(\SB1_3_13/i0[8] ), .A2(
        \SB1_3_13/i0[7] ), .A3(\SB1_3_13/i0[6] ), .ZN(
        \SB1_3_13/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_13/Component_Function_0/N1  ( .A1(\SB1_3_13/i0[10] ), .A2(
        \SB1_3_13/i0[9] ), .ZN(\SB1_3_13/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_13/Component_Function_1/N2  ( .A1(\SB1_3_13/i0_3 ), .A2(
        \SB1_3_13/i1_7 ), .A3(\SB1_3_13/i0[8] ), .ZN(
        \SB1_3_13/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_13/Component_Function_1/N1  ( .A1(\SB1_3_13/i0_3 ), .A2(
        \SB1_3_13/i1[9] ), .ZN(\SB1_3_13/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_14/Component_Function_0/N3  ( .A1(\SB1_3_14/i0[10] ), .A2(
        \SB1_3_14/i0_4 ), .A3(\SB1_3_14/i0_3 ), .ZN(
        \SB1_3_14/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_3_14/Component_Function_0/N1  ( .A1(\SB1_3_14/i0[10] ), .A2(
        \SB1_3_14/i0[9] ), .ZN(\SB1_3_14/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_14/Component_Function_1/N4  ( .A1(\SB1_3_14/i1_7 ), .A2(
        \SB1_3_14/i0[8] ), .A3(\SB1_3_14/i0_4 ), .ZN(
        \SB1_3_14/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_14/Component_Function_1/N3  ( .A1(\SB1_3_14/i1_5 ), .A2(
        \SB1_3_14/i0[6] ), .A3(\SB1_3_14/i0[9] ), .ZN(
        \SB1_3_14/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_14/Component_Function_1/N2  ( .A1(\SB1_3_14/i0_3 ), .A2(
        \SB1_3_14/i1_7 ), .A3(\SB1_3_14/i0[8] ), .ZN(
        \SB1_3_14/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_14/Component_Function_1/N1  ( .A1(\SB1_3_14/i0_3 ), .A2(
        \SB1_3_14/i1[9] ), .ZN(\SB1_3_14/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_15/Component_Function_0/N2  ( .A1(\SB1_3_15/i0[8] ), .A2(
        \SB1_3_15/i0[7] ), .A3(\SB1_3_15/i0[6] ), .ZN(
        \SB1_3_15/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_15/Component_Function_0/N1  ( .A1(\SB1_3_15/i0[10] ), .A2(
        \SB1_3_15/i0[9] ), .ZN(\SB1_3_15/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_16/Component_Function_0/N3  ( .A1(\SB1_3_16/i0[10] ), .A2(
        \SB1_3_16/i0_4 ), .A3(\SB1_3_16/i0_3 ), .ZN(
        \SB1_3_16/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_16/Component_Function_0/N2  ( .A1(\SB1_3_16/i0[8] ), .A2(
        \SB1_3_16/i0[7] ), .A3(\SB1_3_16/i0[6] ), .ZN(
        \SB1_3_16/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_16/Component_Function_0/N1  ( .A1(\SB1_3_16/i0[10] ), .A2(
        \SB1_3_16/i0[9] ), .ZN(\SB1_3_16/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_16/Component_Function_1/N4  ( .A1(\SB1_3_16/i1_7 ), .A2(
        \SB1_3_16/i0[8] ), .A3(\SB1_3_16/i0_4 ), .ZN(
        \SB1_3_16/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_16/Component_Function_1/N2  ( .A1(\SB1_3_16/i0_3 ), .A2(
        \SB1_3_16/i1_7 ), .A3(\SB1_3_16/i0[8] ), .ZN(
        \SB1_3_16/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_16/Component_Function_1/N1  ( .A1(\SB1_3_16/i0_3 ), .A2(
        \SB1_3_16/i1[9] ), .ZN(\SB1_3_16/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_3_16/Component_Function_5/N1  ( .A1(\SB1_3_16/i0_0 ), .A2(
        \SB1_3_16/i3[0] ), .ZN(\SB1_3_16/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_18/Component_Function_0/N2  ( .A1(\SB1_3_18/i0[8] ), .A2(
        \SB1_3_18/i0[7] ), .A3(\SB1_3_18/i0[6] ), .ZN(
        \SB1_3_18/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_18/Component_Function_0/N1  ( .A1(\SB1_3_18/i0[10] ), .A2(
        \SB1_3_18/i0[9] ), .ZN(\SB1_3_18/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_18/Component_Function_5/N4  ( .A1(\SB1_3_18/i0[9] ), .A2(
        \SB1_3_18/i0[6] ), .A3(\SB1_3_18/i0_4 ), .ZN(
        \SB1_3_18/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_19/Component_Function_0/N4  ( .A1(\SB1_3_19/i0[7] ), .A2(
        \SB1_3_19/i0_3 ), .A3(\SB1_3_19/i0_0 ), .ZN(
        \SB1_3_19/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_19/Component_Function_0/N2  ( .A1(\SB1_3_19/i0[8] ), .A2(
        \SB1_3_19/i0[7] ), .A3(\SB1_3_19/i0[6] ), .ZN(
        \SB1_3_19/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_19/Component_Function_0/N1  ( .A1(\SB1_3_19/i0[10] ), .A2(
        \SB1_3_19/i0[9] ), .ZN(\SB1_3_19/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_19/Component_Function_1/N4  ( .A1(\SB1_3_19/i1_7 ), .A2(
        \SB1_3_19/i0[8] ), .A3(\SB1_3_19/i0_4 ), .ZN(
        \SB1_3_19/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_19/Component_Function_1/N3  ( .A1(\SB1_3_19/i1_5 ), .A2(
        \SB1_3_19/i0[6] ), .A3(\SB1_3_19/i0[9] ), .ZN(
        \SB1_3_19/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_19/Component_Function_1/N2  ( .A1(\SB1_3_19/i0_3 ), .A2(
        \SB1_3_19/i1_7 ), .A3(\SB1_3_19/i0[8] ), .ZN(
        \SB1_3_19/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_19/Component_Function_1/N1  ( .A1(\SB1_3_19/i0_3 ), .A2(
        \SB1_3_19/i1[9] ), .ZN(\SB1_3_19/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_3_19/Component_Function_5/N1  ( .A1(\SB1_3_19/i0_0 ), .A2(
        \SB1_3_19/i3[0] ), .ZN(\SB1_3_19/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_20/Component_Function_0/N2  ( .A1(\SB1_3_20/i0[8] ), .A2(
        \SB1_3_20/i0[7] ), .A3(\SB1_3_20/i0[6] ), .ZN(
        \SB1_3_20/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_20/Component_Function_0/N1  ( .A1(\SB1_3_20/i0[10] ), .A2(
        \SB1_3_20/i0[9] ), .ZN(\SB1_3_20/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_20/Component_Function_1/N2  ( .A1(\SB1_3_20/i0_3 ), .A2(
        \SB1_3_20/i1_7 ), .A3(\SB1_3_20/i0[8] ), .ZN(
        \SB1_3_20/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_20/Component_Function_1/N1  ( .A1(\SB1_3_20/i0_3 ), .A2(
        \SB1_3_20/i1[9] ), .ZN(\SB1_3_20/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_21/Component_Function_0/N3  ( .A1(\SB1_3_21/i0[10] ), .A2(
        \SB1_3_21/i0_4 ), .A3(\SB1_3_21/i0_3 ), .ZN(
        \SB1_3_21/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_3_21/Component_Function_0/N1  ( .A1(\SB1_3_21/i0[10] ), .A2(
        \SB1_3_21/i0[9] ), .ZN(\SB1_3_21/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_22/Component_Function_0/N4  ( .A1(\SB1_3_22/i0[7] ), .A2(
        \SB1_3_22/i0_3 ), .A3(\SB1_3_22/i0_0 ), .ZN(
        \SB1_3_22/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_22/Component_Function_0/N3  ( .A1(\SB1_3_22/i0[10] ), .A2(
        \SB1_3_22/i0_4 ), .A3(\SB1_3_22/i0_3 ), .ZN(
        \SB1_3_22/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_3_22/Component_Function_0/N1  ( .A1(\SB1_3_22/i0[10] ), .A2(
        \SB1_3_22/i0[9] ), .ZN(\SB1_3_22/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_22/Component_Function_1/N2  ( .A1(\SB1_3_22/i0_3 ), .A2(
        \SB1_3_22/i1_7 ), .A3(\SB1_3_22/i0[8] ), .ZN(
        \SB1_3_22/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_22/Component_Function_1/N1  ( .A1(\SB1_3_22/i0_3 ), .A2(
        \SB1_3_22/i1[9] ), .ZN(\SB1_3_22/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_23/Component_Function_0/N4  ( .A1(\SB1_3_23/i0[7] ), .A2(
        \SB1_3_23/i0_3 ), .A3(\SB1_3_23/i0_0 ), .ZN(
        \SB1_3_23/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_23/Component_Function_0/N3  ( .A1(\SB1_3_23/i0[10] ), .A2(
        \SB1_3_23/i0_4 ), .A3(\SB1_3_23/i0_3 ), .ZN(
        \SB1_3_23/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_23/Component_Function_0/N2  ( .A1(\SB1_3_23/i0[8] ), .A2(
        \SB1_3_23/i0[7] ), .A3(\SB1_3_23/i0[6] ), .ZN(
        \SB1_3_23/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_24/Component_Function_0/N3  ( .A1(\SB1_3_24/i0[10] ), .A2(
        \SB1_3_24/i0_4 ), .A3(\SB1_3_24/i0_3 ), .ZN(
        \SB1_3_24/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_24/Component_Function_0/N2  ( .A1(\SB1_3_24/i0[8] ), .A2(
        \SB1_3_24/i0[7] ), .A3(\SB1_3_24/i0[6] ), .ZN(
        \SB1_3_24/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_24/Component_Function_0/N1  ( .A1(\SB1_3_24/i0[10] ), .A2(
        \SB1_3_24/i0[9] ), .ZN(\SB1_3_24/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_24/Component_Function_1/N3  ( .A1(\SB1_3_24/i1_5 ), .A2(
        \SB1_3_24/i0[6] ), .A3(\SB1_3_24/i0[9] ), .ZN(
        \SB1_3_24/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_24/Component_Function_1/N2  ( .A1(\SB1_3_24/i0_3 ), .A2(
        \SB1_3_24/i1_7 ), .A3(\SB1_3_24/i0[8] ), .ZN(
        \SB1_3_24/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_24/Component_Function_5/N1  ( .A1(\SB1_3_24/i0_0 ), .A2(
        \SB1_3_24/i3[0] ), .ZN(\SB1_3_24/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_25/Component_Function_0/N4  ( .A1(\SB1_3_25/i0[7] ), .A2(
        \SB1_3_25/i0_3 ), .A3(\SB1_3_25/i0_0 ), .ZN(
        \SB1_3_25/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_25/Component_Function_0/N3  ( .A1(\SB1_3_25/i0[10] ), .A2(
        \SB1_3_25/i0_4 ), .A3(\SB1_3_25/i0_3 ), .ZN(
        \SB1_3_25/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_25/Component_Function_0/N2  ( .A1(\SB1_3_25/i0[8] ), .A2(
        \SB1_3_25/i0[7] ), .A3(\SB1_3_25/i0[6] ), .ZN(
        \SB1_3_25/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_25/Component_Function_0/N1  ( .A1(\SB1_3_25/i0[10] ), .A2(
        \SB1_3_25/i0[9] ), .ZN(\SB1_3_25/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_25/Component_Function_1/N4  ( .A1(\SB1_3_25/i1_7 ), .A2(
        \SB1_3_25/i0[8] ), .A3(\SB1_3_25/i0_4 ), .ZN(
        \SB1_3_25/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_25/Component_Function_1/N2  ( .A1(\SB1_3_25/i0_3 ), .A2(
        \SB1_3_25/i1_7 ), .A3(\SB1_3_25/i0[8] ), .ZN(
        \SB1_3_25/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_26/Component_Function_0/N2  ( .A1(\SB1_3_26/i0[8] ), .A2(
        \SB1_3_26/i0[7] ), .A3(\SB1_3_26/i0[6] ), .ZN(
        \SB1_3_26/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_26/Component_Function_0/N1  ( .A1(\SB1_3_26/i0[10] ), .A2(
        \SB1_3_26/i0[9] ), .ZN(\SB1_3_26/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_27/Component_Function_0/N3  ( .A1(\SB1_3_27/i0[10] ), .A2(
        \SB1_3_27/i0_4 ), .A3(\SB1_3_27/i0_3 ), .ZN(
        \SB1_3_27/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_3_27/Component_Function_0/N1  ( .A1(\SB1_3_27/i0[10] ), .A2(
        \SB1_3_27/i0[9] ), .ZN(\SB1_3_27/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_27/Component_Function_1/N2  ( .A1(\SB1_3_27/i0_3 ), .A2(
        \SB1_3_27/i1_7 ), .A3(\SB1_3_27/i0[8] ), .ZN(
        \SB1_3_27/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_27/Component_Function_1/N1  ( .A1(\SB1_3_27/i0_3 ), .A2(
        \SB1_3_27/i1[9] ), .ZN(\SB1_3_27/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_28/Component_Function_1/N3  ( .A1(\SB1_3_28/i1_5 ), .A2(
        \SB1_3_28/i0[6] ), .A3(\SB1_3_28/i0[9] ), .ZN(
        \SB1_3_28/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_28/Component_Function_1/N2  ( .A1(\SB1_3_28/i0_3 ), .A2(
        \SB1_3_28/i1_7 ), .A3(\SB1_3_28/i0[8] ), .ZN(
        \SB1_3_28/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_29/Component_Function_0/N3  ( .A1(\SB1_3_29/i0[10] ), .A2(
        \SB1_3_29/i0_4 ), .A3(\SB1_3_29/i0_3 ), .ZN(
        \SB1_3_29/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_29/Component_Function_1/N2  ( .A1(\SB1_3_29/i0_3 ), .A2(
        \SB1_3_29/i1_7 ), .A3(\SB1_3_29/i0[8] ), .ZN(
        \SB1_3_29/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_30/Component_Function_0/N1  ( .A1(\SB1_3_30/i0[10] ), .A2(
        \SB1_3_30/i0[9] ), .ZN(\SB1_3_30/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_30/Component_Function_1/N2  ( .A1(\SB1_3_30/i0_3 ), .A2(
        \SB1_3_30/i1_7 ), .A3(\SB1_3_30/i0[8] ), .ZN(
        \SB1_3_30/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_30/Component_Function_1/N1  ( .A1(\SB1_3_30/i0_3 ), .A2(
        \SB1_3_30/i1[9] ), .ZN(\SB1_3_30/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_0/Component_Function_0/N4  ( .A1(n2564), .A2(\SB2_3_0/i0_3 ), 
        .A3(\SB2_3_0/i0_0 ), .ZN(\SB2_3_0/Component_Function_0/NAND4_in[3] )
         );
  NAND2_X1 \SB2_3_0/Component_Function_0/N1  ( .A1(\SB2_3_0/i0[10] ), .A2(
        \SB2_3_0/i0[9] ), .ZN(\SB2_3_0/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_0/Component_Function_1/N4  ( .A1(\SB2_3_0/i1_7 ), .A2(n5513), 
        .A3(\SB1_3_1/buf_output[4] ), .ZN(
        \SB2_3_0/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB2_3_0/Component_Function_1/N1  ( .A1(\SB2_3_0/i0_3 ), .A2(
        \SB2_3_0/i1[9] ), .ZN(\SB2_3_0/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_1/Component_Function_0/N2  ( .A1(\SB2_3_1/i0[8] ), .A2(
        \SB2_3_1/i0[7] ), .A3(\SB2_3_1/i0[6] ), .ZN(
        \SB2_3_1/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_1/Component_Function_0/N1  ( .A1(\SB2_3_1/i0[10] ), .A2(
        \SB2_3_1/i0[9] ), .ZN(\SB2_3_1/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_1/Component_Function_1/N3  ( .A1(\SB2_3_1/i1_5 ), .A2(
        \SB2_3_1/i0[6] ), .A3(\SB2_3_1/i0[9] ), .ZN(
        \SB2_3_1/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_3_1/Component_Function_1/N1  ( .A1(\SB2_3_1/i0_3 ), .A2(
        \SB2_3_1/i1[9] ), .ZN(\SB2_3_1/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_2/Component_Function_0/N4  ( .A1(\SB2_3_2/i0[7] ), .A2(
        \SB2_3_2/i0_3 ), .A3(\SB2_3_2/i0_0 ), .ZN(
        \SB2_3_2/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB2_3_2/Component_Function_0/N1  ( .A1(\SB2_3_2/i0[10] ), .A2(
        \SB2_3_2/i0[9] ), .ZN(\SB2_3_2/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_2/Component_Function_1/N4  ( .A1(\SB2_3_2/i1_7 ), .A2(n5491), 
        .A3(\SB1_3_3/buf_output[4] ), .ZN(
        \SB2_3_2/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_3/Component_Function_0/N2  ( .A1(\SB2_3_3/i0[8] ), .A2(
        \SB2_3_3/i0[7] ), .A3(\SB2_3_3/i0[6] ), .ZN(
        \SB2_3_3/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_3/Component_Function_0/N1  ( .A1(\SB2_3_3/i0[10] ), .A2(
        \SB2_3_3/i0[9] ), .ZN(\SB2_3_3/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_4/Component_Function_1/N2  ( .A1(\SB2_3_4/i0_3 ), .A2(
        \SB2_3_4/i1_7 ), .A3(\SB2_3_4/i0[8] ), .ZN(
        \SB2_3_4/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_4/Component_Function_1/N1  ( .A1(\SB2_3_4/i0_3 ), .A2(
        \SB2_3_4/i1[9] ), .ZN(\SB2_3_4/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_5/Component_Function_1/N2  ( .A1(\SB2_3_5/i0_3 ), .A2(
        \SB2_3_5/i1_7 ), .A3(\SB2_3_5/i0[8] ), .ZN(
        \SB2_3_5/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_6/Component_Function_0/N3  ( .A1(\SB2_3_6/i0[10] ), .A2(
        \SB2_3_6/i0_4 ), .A3(\SB2_3_6/i0_3 ), .ZN(
        \SB2_3_6/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_6/Component_Function_0/N2  ( .A1(\SB2_3_6/i0[8] ), .A2(
        \SB2_3_6/i0[7] ), .A3(\SB2_3_6/i0[6] ), .ZN(
        \SB2_3_6/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_6/Component_Function_0/N1  ( .A1(\SB2_3_6/i0[10] ), .A2(
        \SB2_3_6/i0[9] ), .ZN(\SB2_3_6/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_6/Component_Function_1/N3  ( .A1(\SB2_3_6/i1_5 ), .A2(
        \SB2_3_6/i0[6] ), .A3(\SB2_3_6/i0[9] ), .ZN(
        \SB2_3_6/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_3_6/Component_Function_1/N1  ( .A1(\SB2_3_6/i0_3 ), .A2(
        \SB2_3_6/i1[9] ), .ZN(\SB2_3_6/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_6/Component_Function_5/N1  ( .A1(\SB2_3_6/i0_0 ), .A2(
        \SB2_3_6/i3[0] ), .ZN(\SB2_3_6/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_7/Component_Function_0/N1  ( .A1(\SB2_3_7/i0[10] ), .A2(
        \SB2_3_7/i0[9] ), .ZN(\SB2_3_7/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_7/Component_Function_1/N1  ( .A1(\SB2_3_7/i0_3 ), .A2(
        \SB2_3_7/i1[9] ), .ZN(\SB2_3_7/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_8/Component_Function_0/N1  ( .A1(\SB2_3_8/i0[10] ), .A2(
        \SB2_3_8/i0[9] ), .ZN(\SB2_3_8/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_8/Component_Function_1/N1  ( .A1(\SB2_3_8/i0_3 ), .A2(n3669), 
        .ZN(\SB2_3_8/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_9/Component_Function_0/N2  ( .A1(\SB2_3_9/i0[8] ), .A2(
        \SB2_3_9/i0[7] ), .A3(\SB2_3_9/i0[6] ), .ZN(
        \SB2_3_9/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_9/Component_Function_0/N1  ( .A1(\SB2_3_9/i0[10] ), .A2(
        \SB2_3_9/i0[9] ), .ZN(\SB2_3_9/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_9/Component_Function_1/N3  ( .A1(\SB2_3_9/i1_5 ), .A2(
        \SB2_3_9/i0[6] ), .A3(\SB2_3_9/i0[9] ), .ZN(
        \SB2_3_9/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_3_9/Component_Function_1/N1  ( .A1(\SB2_3_9/i0_3 ), .A2(
        \SB2_3_9/i1[9] ), .ZN(\SB2_3_9/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_10/Component_Function_1/N3  ( .A1(\SB2_3_10/i1_5 ), .A2(
        \SB2_3_10/i0[6] ), .A3(\SB2_3_10/i0[9] ), .ZN(
        \SB2_3_10/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_3_10/Component_Function_1/N1  ( .A1(\SB2_3_10/i0_3 ), .A2(
        \SB2_3_10/i1[9] ), .ZN(\SB2_3_10/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_11/Component_Function_1/N1  ( .A1(\SB2_3_11/i0_3 ), .A2(
        \SB2_3_11/i1[9] ), .ZN(\SB2_3_11/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_12/Component_Function_0/N1  ( .A1(\SB2_3_12/i0[10] ), .A2(
        n1603), .ZN(\SB2_3_12/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_12/Component_Function_1/N3  ( .A1(\SB2_3_12/i1_5 ), .A2(
        \SB2_3_12/i0[6] ), .A3(n1603), .ZN(
        \SB2_3_12/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_12/Component_Function_1/N2  ( .A1(\SB2_3_12/i0_3 ), .A2(
        \SB2_3_12/i1_7 ), .A3(n3651), .ZN(
        \SB2_3_12/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_12/Component_Function_1/N1  ( .A1(\SB2_3_12/i0_3 ), .A2(
        \SB2_3_12/i1[9] ), .ZN(\SB2_3_12/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_13/Component_Function_0/N2  ( .A1(\SB2_3_13/i0[8] ), .A2(
        \SB2_3_13/i0[7] ), .A3(\SB2_3_13/i0[6] ), .ZN(
        \SB2_3_13/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_13/Component_Function_0/N1  ( .A1(\SB2_3_13/i0[10] ), .A2(
        \SB2_3_13/i0[9] ), .ZN(\SB2_3_13/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_13/Component_Function_1/N3  ( .A1(\SB2_3_13/i1_5 ), .A2(
        \SB2_3_13/i0[6] ), .A3(\SB2_3_13/i0[9] ), .ZN(
        \SB2_3_13/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_13/Component_Function_1/N2  ( .A1(\SB2_3_13/i0_3 ), .A2(
        \SB2_3_13/i1_7 ), .A3(\SB2_3_13/i0[8] ), .ZN(
        \SB2_3_13/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_13/Component_Function_1/N1  ( .A1(\SB2_3_13/i0_3 ), .A2(
        \SB2_3_13/i1[9] ), .ZN(\SB2_3_13/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_14/Component_Function_0/N2  ( .A1(\SB2_3_14/i0[8] ), .A2(
        \SB2_3_14/i0[7] ), .A3(\SB2_3_14/i0[6] ), .ZN(
        \SB2_3_14/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_14/Component_Function_0/N1  ( .A1(\SB2_3_14/i0[10] ), .A2(
        \SB2_3_14/i0[9] ), .ZN(\SB2_3_14/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_14/Component_Function_1/N4  ( .A1(\SB2_3_14/i1_7 ), .A2(
        \SB2_3_14/i0[8] ), .A3(\SB2_3_14/i0_4 ), .ZN(
        \SB2_3_14/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_14/Component_Function_1/N2  ( .A1(\SB2_3_14/i0_3 ), .A2(
        \SB2_3_14/i1_7 ), .A3(\SB2_3_14/i0[8] ), .ZN(
        \SB2_3_14/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_14/Component_Function_1/N1  ( .A1(\SB2_3_14/i0_3 ), .A2(
        \SB2_3_14/i1[9] ), .ZN(\SB2_3_14/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_14/Component_Function_5/N4  ( .A1(\SB1_3_19/buf_output[0] ), 
        .A2(\SB1_3_18/buf_output[1] ), .A3(\SB1_3_15/buf_output[4] ), .ZN(
        \SB2_3_14/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB2_3_14/Component_Function_5/N1  ( .A1(\SB2_3_14/i0_0 ), .A2(
        \SB2_3_14/i3[0] ), .ZN(\SB2_3_14/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_15/Component_Function_0/N2  ( .A1(n3670), .A2(
        \SB2_3_15/i0[7] ), .A3(\SB2_3_15/i0[6] ), .ZN(
        \SB2_3_15/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_15/Component_Function_1/N1  ( .A1(\SB2_3_15/i0_3 ), .A2(
        \SB2_3_15/i1[9] ), .ZN(\SB2_3_15/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_16/Component_Function_0/N2  ( .A1(\SB2_3_16/i0[8] ), .A2(
        \SB2_3_16/i0[7] ), .A3(\SB2_3_16/i0[6] ), .ZN(
        \SB2_3_16/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_16/Component_Function_1/N2  ( .A1(\SB2_3_16/i0_3 ), .A2(
        \SB2_3_16/i1_7 ), .A3(\SB2_3_16/i0[8] ), .ZN(
        \SB2_3_16/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_17/Component_Function_0/N4  ( .A1(\SB2_3_17/i0[7] ), .A2(
        \SB1_3_17/buf_output[5] ), .A3(\SB2_3_17/i0_0 ), .ZN(
        \SB2_3_17/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_17/Component_Function_0/N2  ( .A1(\SB2_3_17/i0[8] ), .A2(
        \SB2_3_17/i0[7] ), .A3(\SB2_3_17/i0[6] ), .ZN(
        \SB2_3_17/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_17/Component_Function_0/N1  ( .A1(\SB2_3_17/i0[10] ), .A2(
        \SB2_3_17/i0[9] ), .ZN(\SB2_3_17/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_17/Component_Function_1/N1  ( .A1(\SB2_3_17/i0_3 ), .A2(
        \SB2_3_17/i1[9] ), .ZN(\SB2_3_17/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_18/Component_Function_0/N2  ( .A1(\SB2_3_18/i0[8] ), .A2(
        \SB2_3_18/i0[7] ), .A3(\SB2_3_18/i0[6] ), .ZN(
        \SB2_3_18/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_18/Component_Function_0/N1  ( .A1(\SB2_3_18/i0[10] ), .A2(
        \SB2_3_18/i0[9] ), .ZN(\SB2_3_18/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_18/Component_Function_1/N1  ( .A1(\SB2_3_18/i0_3 ), .A2(
        \SB2_3_18/i1[9] ), .ZN(\SB2_3_18/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_19/Component_Function_0/N2  ( .A1(\SB2_3_19/i0[8] ), .A2(
        \SB2_3_19/i0[7] ), .A3(\SB2_3_19/i0[6] ), .ZN(
        \SB2_3_19/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_19/Component_Function_1/N4  ( .A1(\SB2_3_19/i1_7 ), .A2(
        \SB2_3_19/i0[8] ), .A3(\SB2_3_19/i0_4 ), .ZN(
        \SB2_3_19/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_19/Component_Function_1/N3  ( .A1(\SB2_3_19/i1_5 ), .A2(
        \SB2_3_19/i0[6] ), .A3(\SB2_3_19/i0[9] ), .ZN(
        \SB2_3_19/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_19/Component_Function_1/N2  ( .A1(\SB2_3_19/i0_3 ), .A2(
        \SB2_3_19/i1_7 ), .A3(\SB2_3_19/i0[8] ), .ZN(
        \SB2_3_19/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_19/Component_Function_1/N1  ( .A1(\SB2_3_19/i0_3 ), .A2(
        n5494), .ZN(\SB2_3_19/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_20/Component_Function_0/N1  ( .A1(\SB2_3_20/i0[10] ), .A2(
        \SB2_3_20/i0[9] ), .ZN(\SB2_3_20/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_20/Component_Function_1/N2  ( .A1(\SB2_3_20/i0_3 ), .A2(
        \SB2_3_20/i1_7 ), .A3(\SB2_3_20/i0[8] ), .ZN(
        \SB2_3_20/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_20/Component_Function_1/N1  ( .A1(\SB2_3_20/i0_3 ), .A2(
        \SB2_3_20/i1[9] ), .ZN(\SB2_3_20/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_20/Component_Function_5/N1  ( .A1(n1400), .A2(
        \SB2_3_20/i3[0] ), .ZN(\SB2_3_20/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_21/Component_Function_0/N1  ( .A1(\SB2_3_21/i0[10] ), .A2(
        \SB2_3_21/i0[9] ), .ZN(\SB2_3_21/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_21/Component_Function_1/N3  ( .A1(\SB2_3_21/i1_5 ), .A2(
        \SB2_3_21/i0[6] ), .A3(\SB2_3_21/i0[9] ), .ZN(
        \SB2_3_21/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_21/Component_Function_1/N2  ( .A1(\SB2_3_21/i0_3 ), .A2(
        \SB2_3_21/i1_7 ), .A3(\SB2_3_21/i0[8] ), .ZN(
        \SB2_3_21/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_21/Component_Function_1/N1  ( .A1(\SB2_3_21/i0_3 ), .A2(
        \SB2_3_21/i1[9] ), .ZN(\SB2_3_21/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_22/Component_Function_0/N3  ( .A1(\SB2_3_22/i0[10] ), .A2(
        \SB2_3_22/i0_4 ), .A3(\SB2_3_22/i0_3 ), .ZN(
        \SB2_3_22/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_22/Component_Function_1/N2  ( .A1(\SB2_3_22/i0_3 ), .A2(
        \SB2_3_22/i1_7 ), .A3(\SB2_3_22/i0[8] ), .ZN(
        \SB2_3_22/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_22/Component_Function_1/N1  ( .A1(\SB2_3_22/i0_3 ), .A2(
        \SB2_3_22/i1[9] ), .ZN(\SB2_3_22/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_23/Component_Function_0/N2  ( .A1(\SB2_3_23/i0[8] ), .A2(
        \SB2_3_23/i0[7] ), .A3(\SB2_3_23/i0[6] ), .ZN(
        \SB2_3_23/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_23/Component_Function_0/N1  ( .A1(\SB2_3_23/i0[10] ), .A2(
        \SB1_3_28/buf_output[0] ), .ZN(
        \SB2_3_23/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_24/Component_Function_0/N1  ( .A1(\SB1_3_26/buf_output[3] ), 
        .A2(\SB2_3_24/i0[9] ), .ZN(\SB2_3_24/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_24/Component_Function_1/N2  ( .A1(\SB2_3_24/i0_3 ), .A2(
        \SB2_3_24/i1_7 ), .A3(n2906), .ZN(
        \SB2_3_24/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_25/Component_Function_0/N1  ( .A1(\SB2_3_25/i0[10] ), .A2(
        \SB2_3_25/i0[9] ), .ZN(\SB2_3_25/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_25/Component_Function_1/N2  ( .A1(\SB2_3_25/i0_3 ), .A2(
        \SB2_3_25/i1_7 ), .A3(\SB2_3_25/i0[8] ), .ZN(
        \SB2_3_25/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_26/Component_Function_0/N4  ( .A1(\SB2_3_26/i0[7] ), .A2(
        \SB2_3_26/i0_3 ), .A3(\SB2_3_26/i0_0 ), .ZN(
        \SB2_3_26/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB2_3_26/Component_Function_1/N1  ( .A1(\SB2_3_26/i0_3 ), .A2(
        \SB2_3_26/i1[9] ), .ZN(\SB2_3_26/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_27/Component_Function_0/N2  ( .A1(\SB2_3_27/i0[8] ), .A2(
        \SB2_3_27/i0[7] ), .A3(n3680), .ZN(
        \SB2_3_27/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_27/Component_Function_0/N1  ( .A1(\SB2_3_27/i0[10] ), .A2(
        \RI3[3][24] ), .ZN(\SB2_3_27/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_27/Component_Function_1/N1  ( .A1(\SB2_3_27/i0_3 ), .A2(
        \SB2_3_27/i1[9] ), .ZN(\SB2_3_27/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_28/Component_Function_0/N4  ( .A1(\SB2_3_28/i0[7] ), .A2(
        \SB2_3_28/i0_3 ), .A3(n5489), .ZN(
        \SB2_3_28/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB2_3_28/Component_Function_0/N1  ( .A1(n5511), .A2(
        \SB2_3_28/i0[9] ), .ZN(\SB2_3_28/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_28/Component_Function_1/N3  ( .A1(\SB2_3_28/i1_5 ), .A2(
        \SB2_3_28/i0[6] ), .A3(\SB2_3_28/i0[9] ), .ZN(
        \SB2_3_28/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_3_28/Component_Function_1/N1  ( .A1(\SB2_3_28/i0_3 ), .A2(
        n2911), .ZN(\SB2_3_28/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_30/Component_Function_0/N1  ( .A1(\SB2_3_30/i0[10] ), .A2(
        \SB2_3_30/i0[9] ), .ZN(\SB2_3_30/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_31/Component_Function_0/N2  ( .A1(\SB2_3_31/i0[8] ), .A2(
        \SB2_3_31/i0[7] ), .A3(\SB2_3_31/i0[6] ), .ZN(
        \SB2_3_31/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_31/Component_Function_0/N1  ( .A1(\SB2_3_31/i0[10] ), .A2(
        \SB2_3_31/i0[9] ), .ZN(\SB2_3_31/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_31/Component_Function_1/N1  ( .A1(\SB2_3_31/i0_3 ), .A2(
        \SB2_3_31/i1[9] ), .ZN(\SB2_3_31/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_0/Component_Function_0/N3  ( .A1(\SB3_0/i0[10] ), .A2(
        \SB3_0/i0_4 ), .A3(\SB3_0/i0_3 ), .ZN(
        \SB3_0/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB3_0/Component_Function_0/N1  ( .A1(\SB3_0/i0[10] ), .A2(
        \SB3_0/i0[9] ), .ZN(\SB3_0/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_1/Component_Function_0/N2  ( .A1(\SB3_1/i0[8] ), .A2(
        \SB3_1/i0[7] ), .A3(\SB3_1/i0[6] ), .ZN(
        \SB3_1/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_1/Component_Function_1/N1  ( .A1(\SB3_1/i0_3 ), .A2(n4765), 
        .ZN(\SB3_1/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_2/Component_Function_0/N3  ( .A1(\SB3_2/i0[10] ), .A2(
        \SB3_2/i0_4 ), .A3(\SB3_2/i0_3 ), .ZN(
        \SB3_2/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB3_2/Component_Function_0/N1  ( .A1(\SB3_2/i0[10] ), .A2(
        \SB3_2/i0[9] ), .ZN(\SB3_2/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB3_2/Component_Function_1/N1  ( .A1(\SB3_2/i0_3 ), .A2(
        \SB3_2/i1[9] ), .ZN(\SB3_2/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_3/Component_Function_0/N3  ( .A1(\SB3_3/i0[10] ), .A2(
        \SB3_3/i0_4 ), .A3(\SB3_3/i0_3 ), .ZN(
        \SB3_3/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_3/Component_Function_0/N2  ( .A1(\SB3_3/i0[8] ), .A2(
        \SB3_3/i0[7] ), .A3(\SB3_3/i0[6] ), .ZN(
        \SB3_3/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_3/Component_Function_0/N1  ( .A1(\SB3_3/i0[10] ), .A2(
        \SB3_3/i0[9] ), .ZN(\SB3_3/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_3/Component_Function_1/N2  ( .A1(\SB3_3/i0_3 ), .A2(
        \SB3_3/i1_7 ), .A3(\SB3_3/i0[8] ), .ZN(
        \SB3_3/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_3/Component_Function_1/N1  ( .A1(\SB3_3/i0_3 ), .A2(
        \SB3_3/i1[9] ), .ZN(\SB3_3/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_3/Component_Function_5/N2  ( .A1(\SB3_3/i0_0 ), .A2(
        \SB3_3/i0[6] ), .A3(\SB3_3/i0[10] ), .ZN(
        \SB3_3/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB3_4/Component_Function_0/N2  ( .A1(\SB3_4/i0[8] ), .A2(
        \SB3_4/i0[7] ), .A3(\MC_ARK_ARC_1_3/buf_output[163] ), .ZN(
        \SB3_4/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB3_4/Component_Function_1/N4  ( .A1(\SB3_4/i1_7 ), .A2(
        \SB3_4/i0[8] ), .A3(\SB3_4/i0_4 ), .ZN(
        \SB3_4/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_4/Component_Function_1/N2  ( .A1(\SB3_4/i0_3 ), .A2(
        \SB3_4/i1_7 ), .A3(\SB3_4/i0[8] ), .ZN(
        \SB3_4/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_4/Component_Function_1/N1  ( .A1(\SB3_4/i0_3 ), .A2(
        \SB3_4/i1[9] ), .ZN(\SB3_4/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_5/Component_Function_0/N2  ( .A1(\SB3_5/i0[8] ), .A2(
        \SB3_5/i0[7] ), .A3(\SB3_5/i0[6] ), .ZN(
        \SB3_5/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB3_6/Component_Function_0/N2  ( .A1(\SB3_6/i0[8] ), .A2(
        \SB3_6/i0[7] ), .A3(\SB3_6/i0[6] ), .ZN(
        \SB3_6/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_6/Component_Function_0/N1  ( .A1(\SB3_6/i0[10] ), .A2(
        \SB3_6/i0[9] ), .ZN(\SB3_6/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_7/Component_Function_0/N4  ( .A1(\SB3_7/i0[7] ), .A2(
        \SB3_7/i0_3 ), .A3(\SB3_7/i0_0 ), .ZN(
        \SB3_7/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB3_7/Component_Function_0/N1  ( .A1(\SB3_7/i0[10] ), .A2(
        \SB3_7/i0[9] ), .ZN(\SB3_7/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB3_7/Component_Function_1/N1  ( .A1(\SB3_7/i0_3 ), .A2(
        \SB3_7/i1[9] ), .ZN(\SB3_7/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_8/Component_Function_0/N3  ( .A1(\SB3_8/i0[10] ), .A2(
        \SB3_8/i0_4 ), .A3(\SB3_8/i0_3 ), .ZN(
        \SB3_8/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_8/Component_Function_0/N2  ( .A1(\SB3_8/i0[8] ), .A2(
        \SB3_8/i0[7] ), .A3(\SB3_8/i0[6] ), .ZN(
        \SB3_8/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_8/Component_Function_0/N1  ( .A1(\SB3_8/i0[10] ), .A2(
        \SB3_8/i0[9] ), .ZN(\SB3_8/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_8/Component_Function_5/N2  ( .A1(\SB3_8/i0_0 ), .A2(
        \SB3_8/i0[6] ), .A3(\SB3_8/i0[10] ), .ZN(
        \SB3_8/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB3_9/Component_Function_0/N3  ( .A1(\SB3_9/i0[10] ), .A2(
        \SB3_9/i0_4 ), .A3(\SB3_9/i0_3 ), .ZN(
        \SB3_9/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_9/Component_Function_0/N2  ( .A1(\SB3_9/i0[8] ), .A2(
        \SB3_9/i0[7] ), .A3(\SB3_9/i0[6] ), .ZN(
        \SB3_9/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_9/Component_Function_0/N1  ( .A1(\SB3_9/i0[10] ), .A2(
        \SB3_9/i0[9] ), .ZN(\SB3_9/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_9/Component_Function_1/N4  ( .A1(\SB3_9/i1_7 ), .A2(
        \SB3_9/i0[8] ), .A3(\SB3_9/i0_4 ), .ZN(
        \SB3_9/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_9/Component_Function_1/N2  ( .A1(\SB3_9/i0_3 ), .A2(
        \SB3_9/i1_7 ), .A3(\SB3_9/i0[8] ), .ZN(
        \SB3_9/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_9/Component_Function_1/N1  ( .A1(\SB3_9/i0_3 ), .A2(
        \SB3_9/i1[9] ), .ZN(\SB3_9/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB3_9/Component_Function_5/N1  ( .A1(\SB3_9/i0_0 ), .A2(
        \SB3_9/i3[0] ), .ZN(\SB3_9/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_10/Component_Function_0/N4  ( .A1(\SB3_10/i0[7] ), .A2(
        \SB3_10/i0_3 ), .A3(\SB3_10/i0_0 ), .ZN(
        \SB3_10/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB3_10/Component_Function_0/N3  ( .A1(\SB3_10/i0[10] ), .A2(
        \SB3_10/i0_4 ), .A3(\SB3_10/i0_3 ), .ZN(
        \SB3_10/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB3_10/Component_Function_0/N1  ( .A1(\SB3_10/i0[10] ), .A2(
        \SB3_10/i0[9] ), .ZN(\SB3_10/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB3_10/Component_Function_1/N1  ( .A1(\SB3_10/i0_3 ), .A2(
        \SB3_10/i1[9] ), .ZN(\SB3_10/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB3_11/Component_Function_0/N1  ( .A1(\SB3_11/i0[10] ), .A2(
        \SB3_11/i0[9] ), .ZN(\SB3_11/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_11/Component_Function_1/N2  ( .A1(\SB3_11/i0_3 ), .A2(
        \SB3_11/i1_7 ), .A3(\SB3_11/i0[8] ), .ZN(
        \SB3_11/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_11/Component_Function_1/N1  ( .A1(\SB3_11/i0_3 ), .A2(
        \SB3_11/i1[9] ), .ZN(\SB3_11/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_12/Component_Function_0/N3  ( .A1(\SB3_12/i0[10] ), .A2(
        \SB3_12/i0_4 ), .A3(\SB3_12/i0_3 ), .ZN(
        \SB3_12/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_12/Component_Function_0/N2  ( .A1(\SB3_12/i0[8] ), .A2(
        \SB3_12/i0[7] ), .A3(\SB3_12/i0[6] ), .ZN(
        \SB3_12/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_12/Component_Function_0/N1  ( .A1(\SB3_12/i0[10] ), .A2(
        \SB3_12/i0[9] ), .ZN(\SB3_12/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_13/Component_Function_0/N4  ( .A1(\SB3_13/i0[7] ), .A2(
        \SB3_13/i0_3 ), .A3(\MC_ARK_ARC_1_3/buf_output[110] ), .ZN(
        \SB3_13/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB3_13/Component_Function_0/N3  ( .A1(\SB3_13/i0[10] ), .A2(
        \SB3_13/i0_4 ), .A3(\SB3_13/i0_3 ), .ZN(
        \SB3_13/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB3_13/Component_Function_0/N1  ( .A1(\SB3_13/i0[10] ), .A2(
        \SB3_13/i0[9] ), .ZN(\SB3_13/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_13/Component_Function_1/N2  ( .A1(\SB3_13/i0_3 ), .A2(
        \SB3_13/i1_7 ), .A3(\SB3_13/i0[8] ), .ZN(
        \SB3_13/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_13/Component_Function_1/N1  ( .A1(\SB3_13/i0_3 ), .A2(
        \SB3_13/i1[9] ), .ZN(\SB3_13/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_14/Component_Function_0/N3  ( .A1(\SB3_14/i0[10] ), .A2(
        \SB3_14/i0_4 ), .A3(\SB3_14/i0_3 ), .ZN(
        \SB3_14/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_14/Component_Function_0/N2  ( .A1(\SB3_14/i0[8] ), .A2(
        \SB3_14/i0[7] ), .A3(\SB3_14/i0[6] ), .ZN(
        \SB3_14/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_14/Component_Function_0/N1  ( .A1(\SB3_14/i0[10] ), .A2(
        \SB3_14/i0[9] ), .ZN(\SB3_14/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_14/Component_Function_1/N2  ( .A1(\SB3_14/i0_3 ), .A2(
        \SB3_14/i1_7 ), .A3(\SB3_14/i0[8] ), .ZN(
        \SB3_14/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB3_15/Component_Function_0/N2  ( .A1(\SB3_15/i0[8] ), .A2(
        \SB3_15/i0[7] ), .A3(\SB3_15/i0[6] ), .ZN(
        \SB3_15/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_15/Component_Function_1/N1  ( .A1(\SB3_15/i0_3 ), .A2(
        \SB3_15/i1[9] ), .ZN(\SB3_15/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_15/Component_Function_5/N2  ( .A1(\SB3_15/i0_0 ), .A2(
        \SB3_15/i0[6] ), .A3(\SB3_15/i0[10] ), .ZN(
        \SB3_15/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB3_16/Component_Function_0/N2  ( .A1(\SB3_16/i0[8] ), .A2(
        \SB3_16/i0[7] ), .A3(\SB3_16/i0[6] ), .ZN(
        \SB3_16/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_16/Component_Function_1/N1  ( .A1(\SB3_16/i0_3 ), .A2(
        \SB3_16/i1[9] ), .ZN(\SB3_16/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB3_17/Component_Function_0/N1  ( .A1(\SB3_17/i0[10] ), .A2(
        \SB3_17/i0[9] ), .ZN(\SB3_17/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB3_17/Component_Function_1/N1  ( .A1(\SB3_17/i0_3 ), .A2(
        \SB3_17/i1[9] ), .ZN(\SB3_17/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB3_18/Component_Function_0/N1  ( .A1(\SB3_18/i0[10] ), .A2(
        \SB3_18/i0[9] ), .ZN(\SB3_18/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_19/Component_Function_0/N3  ( .A1(\SB3_19/i0[10] ), .A2(
        \SB3_19/i0_4 ), .A3(\SB3_19/i0_3 ), .ZN(
        \SB3_19/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_19/Component_Function_0/N2  ( .A1(\SB3_19/i0[8] ), .A2(
        \SB3_19/i0[7] ), .A3(\SB3_19/i0[6] ), .ZN(
        \SB3_19/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB3_19/Component_Function_1/N4  ( .A1(\SB3_19/i1_7 ), .A2(
        \SB3_19/i0[8] ), .A3(\SB3_19/i0_4 ), .ZN(
        \SB3_19/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_19/Component_Function_1/N2  ( .A1(\SB3_19/i0_3 ), .A2(
        \SB3_19/i1_7 ), .A3(\SB3_19/i0[8] ), .ZN(
        \SB3_19/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_19/Component_Function_1/N1  ( .A1(\SB3_19/i0_3 ), .A2(
        \SB3_19/i1[9] ), .ZN(\SB3_19/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_20/Component_Function_0/N3  ( .A1(\SB3_20/i0[10] ), .A2(
        \SB3_20/i0_4 ), .A3(\SB3_20/i0_3 ), .ZN(
        \SB3_20/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_20/Component_Function_0/N2  ( .A1(\SB3_20/i0[8] ), .A2(
        \SB3_20/i0[7] ), .A3(\SB3_20/i0[6] ), .ZN(
        \SB3_20/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_20/Component_Function_0/N1  ( .A1(\SB3_20/i0[10] ), .A2(
        \SB3_20/i0[9] ), .ZN(\SB3_20/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_20/Component_Function_1/N2  ( .A1(\SB3_20/i0_3 ), .A2(
        \SB3_20/i1_7 ), .A3(\SB3_20/i0[8] ), .ZN(
        \SB3_20/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_20/Component_Function_1/N1  ( .A1(\SB3_20/i0_3 ), .A2(
        \SB3_20/i1[9] ), .ZN(\SB3_20/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_21/Component_Function_0/N2  ( .A1(\SB3_21/i0[8] ), .A2(
        \SB3_21/i0[7] ), .A3(\SB3_21/i0[6] ), .ZN(
        \SB3_21/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB3_21/Component_Function_1/N2  ( .A1(\SB3_21/i0_3 ), .A2(
        \SB3_21/i1_7 ), .A3(\SB3_21/i0[8] ), .ZN(
        \SB3_21/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_21/Component_Function_5/N1  ( .A1(\SB3_21/i0_0 ), .A2(
        \SB3_21/i3[0] ), .ZN(\SB3_21/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_22/Component_Function_0/N3  ( .A1(\SB3_22/i0[10] ), .A2(
        \SB3_22/i0_4 ), .A3(\SB3_22/i0_3 ), .ZN(
        \SB3_22/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB3_22/Component_Function_0/N1  ( .A1(\SB3_22/i0[10] ), .A2(
        \SB3_22/i0[9] ), .ZN(\SB3_22/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_23/Component_Function_0/N4  ( .A1(\SB3_23/i0[7] ), .A2(
        \SB3_23/i0_3 ), .A3(\SB3_23/i0_0 ), .ZN(
        \SB3_23/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB3_23/Component_Function_1/N2  ( .A1(\SB3_23/i0_3 ), .A2(
        \SB3_23/i1_7 ), .A3(\SB3_23/i0[8] ), .ZN(
        \SB3_23/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_24/Component_Function_0/N1  ( .A1(\SB3_24/i0[10] ), .A2(
        \SB3_24/i0[9] ), .ZN(\SB3_24/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_24/Component_Function_1/N2  ( .A1(\SB3_24/i0_3 ), .A2(
        \SB3_24/i1_7 ), .A3(\SB3_24/i0[8] ), .ZN(
        \SB3_24/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_24/Component_Function_1/N1  ( .A1(\SB3_24/i0_3 ), .A2(
        \SB3_24/i1[9] ), .ZN(\SB3_24/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_25/Component_Function_0/N4  ( .A1(\SB3_25/i0[7] ), .A2(
        \SB3_25/i0_3 ), .A3(\SB3_25/i0_0 ), .ZN(
        \SB3_25/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB3_25/Component_Function_0/N3  ( .A1(\SB3_25/i0[10] ), .A2(
        \SB3_25/i0_4 ), .A3(\SB3_25/i0_3 ), .ZN(
        \SB3_25/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB3_25/Component_Function_0/N1  ( .A1(\SB3_25/i0[10] ), .A2(
        \SB3_25/i0[9] ), .ZN(\SB3_25/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_25/Component_Function_1/N3  ( .A1(\SB3_25/i1_5 ), .A2(
        \SB3_25/i0[6] ), .A3(\SB3_25/i0[9] ), .ZN(
        \SB3_25/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_25/Component_Function_1/N2  ( .A1(\SB3_25/i0_3 ), .A2(
        \SB3_25/i1_7 ), .A3(\SB3_25/i0[8] ), .ZN(
        \SB3_25/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_25/Component_Function_1/N1  ( .A1(\SB3_25/i0_3 ), .A2(
        \SB3_25/i1[9] ), .ZN(\SB3_25/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_26/Component_Function_0/N3  ( .A1(\SB3_26/i0[10] ), .A2(
        \SB3_26/i0_4 ), .A3(\SB3_26/i0_3 ), .ZN(
        \SB3_26/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB3_26/Component_Function_0/N1  ( .A1(\SB3_26/i0[10] ), .A2(
        \SB3_26/i0[9] ), .ZN(\SB3_26/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_26/Component_Function_1/N2  ( .A1(\SB3_26/i0_3 ), .A2(
        \SB3_26/i1_7 ), .A3(\SB3_26/i0[8] ), .ZN(
        \SB3_26/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_26/Component_Function_1/N1  ( .A1(\SB3_26/i0_3 ), .A2(
        \SB3_26/i1[9] ), .ZN(\SB3_26/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB3_26/Component_Function_5/N1  ( .A1(\SB3_26/i0_0 ), .A2(
        \SB3_26/i3[0] ), .ZN(\SB3_26/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB3_27/Component_Function_0/N3  ( .A1(\SB3_27/i0[10] ), .A2(
        \SB3_27/i0_4 ), .A3(\SB3_27/i0_3 ), .ZN(
        \SB3_27/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_27/Component_Function_0/N2  ( .A1(\SB3_27/i0[8] ), .A2(
        \SB3_27/i0[7] ), .A3(\SB3_27/i0[6] ), .ZN(
        \SB3_27/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB3_27/Component_Function_1/N4  ( .A1(\SB3_27/i1_7 ), .A2(
        \SB3_27/i0[8] ), .A3(\SB3_27/i0_4 ), .ZN(
        \SB3_27/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_27/Component_Function_1/N2  ( .A1(\SB3_27/i0_3 ), .A2(
        \SB3_27/i1_7 ), .A3(\SB3_27/i0[8] ), .ZN(
        \SB3_27/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_27/Component_Function_1/N1  ( .A1(\SB3_27/i0_3 ), .A2(n4764), 
        .ZN(\SB3_27/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_28/Component_Function_0/N3  ( .A1(\SB3_28/i0[10] ), .A2(
        \SB3_28/i0_4 ), .A3(\SB3_28/i0_3 ), .ZN(
        \SB3_28/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_28/Component_Function_0/N2  ( .A1(\SB3_28/i0[8] ), .A2(
        \SB3_28/i0[7] ), .A3(\SB3_28/i0[6] ), .ZN(
        \SB3_28/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_28/Component_Function_0/N1  ( .A1(\SB3_28/i0[10] ), .A2(
        \SB3_28/i0[9] ), .ZN(\SB3_28/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_28/Component_Function_1/N3  ( .A1(\SB3_28/i1_5 ), .A2(
        \SB3_28/i0[6] ), .A3(\SB3_28/i0[9] ), .ZN(
        \SB3_28/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB3_28/Component_Function_1/N1  ( .A1(\SB3_28/i0_3 ), .A2(
        \SB3_28/i1[9] ), .ZN(\SB3_28/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_29/Component_Function_0/N3  ( .A1(\SB3_29/i0[10] ), .A2(
        \SB3_29/i0_4 ), .A3(\SB3_29/i0_3 ), .ZN(
        \SB3_29/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB3_29/Component_Function_0/N2  ( .A1(\SB3_29/i0[8] ), .A2(
        \SB3_29/i0[7] ), .A3(\SB3_29/i0[6] ), .ZN(
        \SB3_29/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_29/Component_Function_0/N1  ( .A1(\SB3_29/i0[10] ), .A2(
        \SB3_29/i0[9] ), .ZN(\SB3_29/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_29/Component_Function_1/N3  ( .A1(\SB3_29/i1_5 ), .A2(
        \SB3_29/i0[6] ), .A3(\SB3_29/i0[9] ), .ZN(
        \SB3_29/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_29/Component_Function_1/N2  ( .A1(\SB3_29/i0_3 ), .A2(
        \SB3_29/i1_7 ), .A3(\SB3_29/i0[8] ), .ZN(
        \SB3_29/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_29/Component_Function_1/N1  ( .A1(\SB3_29/i0_3 ), .A2(
        \SB3_29/i1[9] ), .ZN(\SB3_29/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB3_30/Component_Function_0/N2  ( .A1(\SB3_30/i0[8] ), .A2(
        \SB3_30/i0[7] ), .A3(\SB3_30/i0[6] ), .ZN(
        \SB3_30/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB3_30/Component_Function_0/N1  ( .A1(\SB3_30/i0[10] ), .A2(
        \SB3_30/i0[9] ), .ZN(\SB3_30/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_30/Component_Function_1/N2  ( .A1(\SB3_30/i0_3 ), .A2(
        \SB3_30/i1_7 ), .A3(\SB3_30/i0[8] ), .ZN(
        \SB3_30/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB3_31/Component_Function_0/N1  ( .A1(\SB3_31/i0[10] ), .A2(
        \SB3_31/i0[9] ), .ZN(\SB3_31/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB3_31/Component_Function_1/N1  ( .A1(\SB3_31/i0_3 ), .A2(
        \SB3_31/i1[9] ), .ZN(\SB3_31/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_0/Component_Function_0/N3  ( .A1(\SB4_0/i0[10] ), .A2(
        \SB4_0/i0_4 ), .A3(\SB4_0/i0_3 ), .ZN(
        \SB4_0/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB4_0/Component_Function_0/N2  ( .A1(\SB4_0/i0[8] ), .A2(
        \SB4_0/i0[7] ), .A3(\SB4_0/i0[6] ), .ZN(
        \SB4_0/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB4_0/Component_Function_1/N4  ( .A1(\SB4_0/i1_7 ), .A2(
        \SB4_0/i0[8] ), .A3(\SB4_0/i0_4 ), .ZN(
        \SB4_0/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_0/Component_Function_1/N3  ( .A1(\SB4_0/i1_5 ), .A2(
        \SB4_0/i0[6] ), .A3(\SB4_0/i0[9] ), .ZN(
        \SB4_0/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_0/Component_Function_1/N2  ( .A1(\SB4_0/i0_3 ), .A2(
        \SB4_0/i1_7 ), .A3(\SB4_0/i0[8] ), .ZN(
        \SB4_0/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB4_0/Component_Function_5/N4  ( .A1(\SB4_0/i0[9] ), .A2(
        \SB4_0/i0[6] ), .A3(\SB4_0/i0_4 ), .ZN(
        \SB4_0/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB4_0/Component_Function_5/N1  ( .A1(\SB3_3/buf_output[2] ), .A2(
        \SB4_0/i3[0] ), .ZN(\SB4_0/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_1/Component_Function_1/N2  ( .A1(\SB4_1/i0_3 ), .A2(
        \SB4_1/i1_7 ), .A3(\SB4_1/i0[8] ), .ZN(
        \SB4_1/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_1/Component_Function_5/N1  ( .A1(\SB4_1/i0_0 ), .A2(
        \SB4_1/i3[0] ), .ZN(\SB4_1/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_2/Component_Function_1/N2  ( .A1(\SB4_2/i0_3 ), .A2(
        \SB4_2/i1_7 ), .A3(\SB4_2/i0[8] ), .ZN(
        \SB4_2/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_2/Component_Function_1/N1  ( .A1(\SB4_2/i0_3 ), .A2(
        \SB4_2/i1[9] ), .ZN(\SB4_2/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_3/Component_Function_1/N3  ( .A1(\SB4_3/i1_5 ), .A2(
        \SB4_3/i0[6] ), .A3(\SB4_3/i0[9] ), .ZN(
        \SB4_3/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB4_3/Component_Function_1/N1  ( .A1(\SB4_3/i0_3 ), .A2(n1371), 
        .ZN(\SB4_3/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_3/Component_Function_5/N4  ( .A1(\SB4_3/i0[9] ), .A2(
        \SB4_3/i0[6] ), .A3(\SB4_3/i0_4 ), .ZN(
        \SB4_3/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB4_3/Component_Function_5/N2  ( .A1(\SB3_6/buf_output[2] ), .A2(
        \SB4_3/i0[6] ), .A3(\SB3_5/buf_output[3] ), .ZN(
        \SB4_3/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB4_4/Component_Function_0/N2  ( .A1(\SB4_4/i0[8] ), .A2(
        \SB4_4/i0[7] ), .A3(\SB4_4/i0[6] ), .ZN(
        \SB4_4/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB4_4/Component_Function_0/N1  ( .A1(\SB4_4/i0[10] ), .A2(
        \SB4_4/i0[9] ), .ZN(\SB4_4/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_4/Component_Function_1/N3  ( .A1(\SB4_4/i1_5 ), .A2(
        \SB4_4/i0[6] ), .A3(\SB4_4/i0[9] ), .ZN(
        \SB4_4/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_4/Component_Function_1/N2  ( .A1(\SB4_4/i0_3 ), .A2(
        \SB4_4/i1_7 ), .A3(\SB4_4/i0[8] ), .ZN(
        \SB4_4/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_4/Component_Function_1/N1  ( .A1(\SB4_4/i0_3 ), .A2(n3655), 
        .ZN(\SB4_4/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_4/Component_Function_5/N3  ( .A1(n3655), .A2(\SB4_4/i0_4 ), 
        .A3(\SB4_4/i0_3 ), .ZN(\SB4_4/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 \SB4_4/Component_Function_5/N1  ( .A1(\SB3_7/buf_output[2] ), .A2(
        \SB4_4/i3[0] ), .ZN(\SB4_4/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_5/Component_Function_1/N3  ( .A1(\SB4_5/i1_5 ), .A2(
        \SB4_5/i0[6] ), .A3(\SB4_5/i0[9] ), .ZN(
        \SB4_5/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_5/Component_Function_1/N2  ( .A1(\SB4_5/i0_3 ), .A2(
        \SB4_5/i1_7 ), .A3(\SB4_5/i0[8] ), .ZN(
        \SB4_5/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_5/Component_Function_1/N1  ( .A1(\SB4_5/i0_3 ), .A2(
        \SB4_5/i1[9] ), .ZN(\SB4_5/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_5/Component_Function_5/N2  ( .A1(\SB4_5/i0_0 ), .A2(
        \SB4_5/i0[6] ), .A3(\SB4_5/i0[10] ), .ZN(
        \SB4_5/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB4_6/Component_Function_0/N4  ( .A1(\SB4_6/i0[7] ), .A2(
        \SB4_6/i0_3 ), .A3(\SB4_6/i0_0 ), .ZN(
        \SB4_6/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB4_6/Component_Function_1/N4  ( .A1(\SB4_6/i1_7 ), .A2(n579), 
        .A3(\SB4_6/i0_4 ), .ZN(\SB4_6/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_6/Component_Function_1/N2  ( .A1(\SB4_6/i0_3 ), .A2(
        \SB4_6/i1_7 ), .A3(n579), .ZN(\SB4_6/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_6/Component_Function_1/N1  ( .A1(\SB4_6/i0_3 ), .A2(
        \SB4_6/i1[9] ), .ZN(\SB4_6/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_6/Component_Function_5/N4  ( .A1(\SB4_6/i0[9] ), .A2(
        \SB4_6/i0[6] ), .A3(\SB4_6/i0_4 ), .ZN(
        \SB4_6/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB4_6/Component_Function_5/N1  ( .A1(\SB4_6/i0_0 ), .A2(
        \SB4_6/i3[0] ), .ZN(\SB4_6/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_7/Component_Function_0/N2  ( .A1(\SB4_7/i0[8] ), .A2(
        \SB4_7/i0[7] ), .A3(\SB4_7/i0[6] ), .ZN(
        \SB4_7/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB4_7/Component_Function_1/N4  ( .A1(\SB4_7/i1_7 ), .A2(
        \SB4_7/i0[8] ), .A3(\SB3_8/buf_output[4] ), .ZN(
        \SB4_7/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_7/Component_Function_1/N3  ( .A1(\SB4_7/i1_5 ), .A2(
        \SB4_7/i0[6] ), .A3(\SB4_7/i0[9] ), .ZN(
        \SB4_7/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_7/Component_Function_1/N2  ( .A1(\SB4_7/i0_3 ), .A2(
        \SB4_7/i1_7 ), .A3(\SB4_7/i0[8] ), .ZN(
        \SB4_7/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB4_7/Component_Function_5/N4  ( .A1(\SB4_7/i0[9] ), .A2(
        \SB4_7/i0[6] ), .A3(\SB4_7/i0_4 ), .ZN(
        \SB4_7/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB4_7/Component_Function_5/N2  ( .A1(\SB4_7/i0_0 ), .A2(
        \SB4_7/i0[6] ), .A3(\SB4_7/i0[10] ), .ZN(
        \SB4_7/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB4_7/Component_Function_5/N1  ( .A1(\SB4_7/i0_0 ), .A2(
        \SB4_7/i3[0] ), .ZN(\SB4_7/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_8/Component_Function_0/N2  ( .A1(\SB4_8/i0[8] ), .A2(
        \SB4_8/i0[7] ), .A3(\SB4_8/i0[6] ), .ZN(
        \SB4_8/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB4_8/Component_Function_1/N3  ( .A1(\SB4_8/i1_5 ), .A2(
        \SB4_8/i0[6] ), .A3(\SB4_8/i0[9] ), .ZN(
        \SB4_8/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_8/Component_Function_5/N3  ( .A1(\SB4_8/i1[9] ), .A2(
        \SB4_8/i0_4 ), .A3(\SB4_8/i0_3 ), .ZN(
        \SB4_8/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB4_9/Component_Function_0/N4  ( .A1(\SB4_9/i0[7] ), .A2(
        \SB4_9/i0_3 ), .A3(\SB4_9/i0_0 ), .ZN(
        \SB4_9/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB4_9/Component_Function_0/N3  ( .A1(\SB4_9/i0[10] ), .A2(
        \SB4_9/i0_4 ), .A3(\SB4_9/i0_3 ), .ZN(
        \SB4_9/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB4_9/Component_Function_0/N2  ( .A1(\SB4_9/i0[8] ), .A2(
        \SB4_9/i0[7] ), .A3(\SB4_9/i0[6] ), .ZN(
        \SB4_9/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB4_9/Component_Function_1/N2  ( .A1(\SB4_9/i0_3 ), .A2(
        \SB4_9/i1_7 ), .A3(\SB4_9/i0[8] ), .ZN(
        \SB4_9/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB4_9/Component_Function_5/N4  ( .A1(\SB4_9/i0[9] ), .A2(
        \SB4_9/i0[6] ), .A3(\SB4_9/i0_4 ), .ZN(
        \SB4_9/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB4_9/Component_Function_5/N3  ( .A1(\SB4_9/i1[9] ), .A2(
        \SB4_9/i0_4 ), .A3(\SB4_9/i0_3 ), .ZN(
        \SB4_9/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 \SB4_9/Component_Function_5/N1  ( .A1(\SB4_9/i0_0 ), .A2(
        \SB4_9/i3[0] ), .ZN(\SB4_9/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_10/Component_Function_1/N4  ( .A1(\SB4_10/i1_7 ), .A2(
        \SB4_10/i0[8] ), .A3(\SB4_10/i0_4 ), .ZN(
        \SB4_10/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_10/Component_Function_1/N3  ( .A1(\SB4_10/i1_5 ), .A2(
        \SB4_10/i0[6] ), .A3(\SB4_10/i0[9] ), .ZN(
        \SB4_10/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_10/Component_Function_1/N2  ( .A1(\SB4_10/i0_3 ), .A2(
        \SB4_10/i1_7 ), .A3(\SB4_10/i0[8] ), .ZN(
        \SB4_10/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_10/Component_Function_5/N1  ( .A1(\SB3_13/buf_output[2] ), 
        .A2(\SB4_10/i3[0] ), .ZN(\SB4_10/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_11/Component_Function_1/N4  ( .A1(\SB4_11/i1_7 ), .A2(
        \SB4_11/i0[8] ), .A3(\SB4_11/i0_4 ), .ZN(
        \SB4_11/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_12/Component_Function_0/N3  ( .A1(\SB4_12/i0[10] ), .A2(
        \SB4_12/i0_4 ), .A3(\SB4_12/i0_3 ), .ZN(
        \SB4_12/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB4_12/Component_Function_0/N2  ( .A1(\SB4_12/i0[8] ), .A2(
        \SB4_12/i0[7] ), .A3(\SB4_12/i0[6] ), .ZN(
        \SB4_12/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB4_12/Component_Function_1/N3  ( .A1(\SB4_12/i1_5 ), .A2(
        \SB4_12/i0[6] ), .A3(\SB4_12/i0[9] ), .ZN(
        \SB4_12/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_12/Component_Function_1/N2  ( .A1(\SB4_12/i0_3 ), .A2(
        \SB4_12/i1_7 ), .A3(\SB4_12/i0[8] ), .ZN(
        \SB4_12/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_12/Component_Function_1/N1  ( .A1(\SB4_12/i0_3 ), .A2(
        \SB4_12/i1[9] ), .ZN(\SB4_12/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_12/Component_Function_5/N4  ( .A1(\SB4_12/i0[9] ), .A2(
        \SB4_12/i0[6] ), .A3(\SB4_12/i0_4 ), .ZN(
        \SB4_12/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB4_12/Component_Function_5/N2  ( .A1(\SB4_12/i0_0 ), .A2(
        \SB4_12/i0[6] ), .A3(\SB4_12/i0[10] ), .ZN(
        \SB4_12/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB4_13/Component_Function_0/N2  ( .A1(n3683), .A2(\SB4_13/i0[7] ), 
        .A3(\SB4_13/i0[6] ), .ZN(\SB4_13/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB4_13/Component_Function_0/N1  ( .A1(\SB4_13/i0[10] ), .A2(
        \SB4_13/i0[9] ), .ZN(\SB4_13/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_13/Component_Function_1/N2  ( .A1(\SB4_13/i0_3 ), .A2(
        \SB4_13/i1_7 ), .A3(n3683), .ZN(
        \SB4_13/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB4_14/Component_Function_1/N2  ( .A1(\SB4_14/i0_3 ), .A2(
        \SB4_14/i1_7 ), .A3(\SB4_14/i0[8] ), .ZN(
        \SB4_14/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB4_14/Component_Function_5/N3  ( .A1(\SB4_14/i1[9] ), .A2(
        \SB4_14/i0_4 ), .A3(\SB4_14/i0_3 ), .ZN(
        \SB4_14/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB4_15/Component_Function_0/N2  ( .A1(\SB4_15/i0[8] ), .A2(
        \SB4_15/i0[7] ), .A3(\SB4_15/i0[6] ), .ZN(
        \SB4_15/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB4_15/Component_Function_1/N3  ( .A1(\SB4_15/i1_5 ), .A2(
        \SB4_15/i0[6] ), .A3(\SB4_15/i0[9] ), .ZN(
        \SB4_15/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_15/Component_Function_1/N2  ( .A1(\SB4_15/i0_3 ), .A2(
        \SB4_15/i1_7 ), .A3(\SB4_15/i0[8] ), .ZN(
        \SB4_15/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_15/Component_Function_1/N1  ( .A1(\SB4_15/i0_3 ), .A2(
        \SB4_15/i1[9] ), .ZN(\SB4_15/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_15/Component_Function_5/N4  ( .A1(\SB4_15/i0[9] ), .A2(
        \SB4_15/i0[6] ), .A3(\SB4_15/i0_4 ), .ZN(
        \SB4_15/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB4_15/Component_Function_5/N3  ( .A1(\SB4_15/i1[9] ), .A2(
        \SB4_15/i0_4 ), .A3(\SB4_15/i0_3 ), .ZN(
        \SB4_15/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB4_15/Component_Function_5/N2  ( .A1(\SB4_15/i0_0 ), .A2(
        \SB4_15/i0[6] ), .A3(\SB4_15/i0[10] ), .ZN(
        \SB4_15/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB4_15/Component_Function_5/N1  ( .A1(\SB4_15/i0_0 ), .A2(
        \SB4_15/i3[0] ), .ZN(\SB4_15/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_16/Component_Function_0/N3  ( .A1(\SB4_16/i0[10] ), .A2(
        \SB4_16/i0_4 ), .A3(\SB4_16/i0_3 ), .ZN(
        \SB4_16/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB4_16/Component_Function_0/N2  ( .A1(\SB4_16/i0[8] ), .A2(
        \SB4_16/i0[7] ), .A3(\SB4_16/i0[6] ), .ZN(
        \SB4_16/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB4_17/Component_Function_0/N3  ( .A1(\SB4_17/i0[10] ), .A2(
        \SB4_17/i0_4 ), .A3(\SB4_17/i0_3 ), .ZN(
        \SB4_17/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB4_17/Component_Function_0/N2  ( .A1(n3661), .A2(\SB4_17/i0[7] ), 
        .A3(\SB4_17/i0[6] ), .ZN(\SB4_17/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB4_17/Component_Function_1/N3  ( .A1(\SB4_17/i1_5 ), .A2(
        \SB4_17/i0[6] ), .A3(\SB4_17/i0[9] ), .ZN(
        \SB4_17/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_17/Component_Function_1/N2  ( .A1(\SB4_17/i0_3 ), .A2(
        \SB4_17/i1_7 ), .A3(n3661), .ZN(
        \SB4_17/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_17/Component_Function_5/N1  ( .A1(\SB4_17/i0_0 ), .A2(
        \SB4_17/i3[0] ), .ZN(\SB4_17/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_18/Component_Function_1/N2  ( .A1(\SB4_18/i0_3 ), .A2(
        \SB4_18/i1_7 ), .A3(n3662), .ZN(
        \SB4_18/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB4_18/Component_Function_5/N3  ( .A1(\SB4_18/i1[9] ), .A2(
        \SB4_18/i0_4 ), .A3(\SB4_18/i0_3 ), .ZN(
        \SB4_18/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB4_19/Component_Function_0/N3  ( .A1(\SB3_21/buf_output[3] ), 
        .A2(\SB4_19/i0_4 ), .A3(\SB4_19/i0_3 ), .ZN(
        \SB4_19/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB4_19/Component_Function_0/N2  ( .A1(n3668), .A2(\SB4_19/i0[7] ), 
        .A3(\SB4_19/i0[6] ), .ZN(\SB4_19/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB4_19/Component_Function_0/N1  ( .A1(\SB3_21/buf_output[3] ), 
        .A2(\SB4_19/i0[9] ), .ZN(\SB4_19/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_19/Component_Function_1/N2  ( .A1(\SB4_19/i0_3 ), .A2(
        \SB4_19/i1_7 ), .A3(n3668), .ZN(
        \SB4_19/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB4_19/Component_Function_5/N2  ( .A1(\SB4_19/i0_0 ), .A2(
        \SB4_19/i0[6] ), .A3(\SB3_21/buf_output[3] ), .ZN(
        \SB4_19/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB4_21/Component_Function_0/N3  ( .A1(\SB4_21/i0[10] ), .A2(
        \SB4_21/i0_4 ), .A3(\SB4_21/i0_3 ), .ZN(
        \SB4_21/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB4_21/Component_Function_1/N4  ( .A1(\SB4_21/i1_7 ), .A2(
        \SB4_21/i0[8] ), .A3(\SB4_21/i0_4 ), .ZN(
        \SB4_21/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_21/Component_Function_1/N3  ( .A1(\SB4_21/i1_5 ), .A2(
        \SB4_21/i0[6] ), .A3(\SB4_21/i0[9] ), .ZN(
        \SB4_21/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_21/Component_Function_1/N2  ( .A1(\SB4_21/i0_3 ), .A2(
        \SB4_21/i1_7 ), .A3(\SB4_21/i0[8] ), .ZN(
        \SB4_21/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_21/Component_Function_1/N1  ( .A1(\SB4_21/i0_3 ), .A2(n3666), 
        .ZN(\SB4_21/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_21/Component_Function_5/N3  ( .A1(n3666), .A2(\SB4_21/i0_4 ), 
        .A3(\SB4_21/i0_3 ), .ZN(\SB4_21/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB4_21/Component_Function_5/N2  ( .A1(\SB3_24/buf_output[2] ), 
        .A2(\SB4_21/i0[6] ), .A3(\SB4_21/i0[10] ), .ZN(
        \SB4_21/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB4_21/Component_Function_5/N1  ( .A1(\SB3_24/buf_output[2] ), 
        .A2(\SB4_21/i3[0] ), .ZN(\SB4_21/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_22/Component_Function_0/N2  ( .A1(\SB4_22/i0[8] ), .A2(
        \SB4_22/i0[7] ), .A3(\SB4_22/i0[6] ), .ZN(
        \SB4_22/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB4_22/Component_Function_1/N2  ( .A1(\SB4_22/i0_3 ), .A2(
        \SB4_22/i1_7 ), .A3(\SB4_22/i0[8] ), .ZN(
        \SB4_22/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB4_23/Component_Function_0/N2  ( .A1(\SB4_23/i0[8] ), .A2(
        \SB4_23/i0[7] ), .A3(\SB4_23/i0[6] ), .ZN(
        \SB4_23/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB4_23/Component_Function_1/N3  ( .A1(\SB4_23/i1_5 ), .A2(
        \SB4_23/i0[6] ), .A3(\SB4_23/i0[9] ), .ZN(
        \SB4_23/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_23/Component_Function_1/N2  ( .A1(\SB4_23/i0_3 ), .A2(
        \SB4_23/i1_7 ), .A3(\SB4_23/i0[8] ), .ZN(
        \SB4_23/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB4_23/Component_Function_5/N2  ( .A1(\SB4_23/i0_0 ), .A2(
        \SB4_23/i0[6] ), .A3(\SB4_23/i0[10] ), .ZN(
        \SB4_23/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB4_23/Component_Function_5/N1  ( .A1(\SB4_23/i0_0 ), .A2(
        \SB4_23/i3[0] ), .ZN(\SB4_23/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_24/Component_Function_0/N2  ( .A1(\SB4_24/i0[8] ), .A2(
        \SB4_24/i0[7] ), .A3(\SB4_24/i0[6] ), .ZN(
        \SB4_24/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB4_24/Component_Function_0/N1  ( .A1(\SB4_24/i0[10] ), .A2(
        \SB4_24/i0[9] ), .ZN(\SB4_24/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB4_24/Component_Function_1/N4  ( .A1(\SB4_24/i1_7 ), .A2(
        \SB4_24/i0[8] ), .A3(\SB4_24/i0_4 ), .ZN(
        \SB4_24/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_24/Component_Function_1/N2  ( .A1(\SB4_24/i0_3 ), .A2(
        \SB4_24/i1_7 ), .A3(\SB4_24/i0[8] ), .ZN(
        \SB4_24/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_24/Component_Function_5/N1  ( .A1(\SB4_24/i0_0 ), .A2(
        \SB4_24/i3[0] ), .ZN(\SB4_24/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_25/Component_Function_0/N3  ( .A1(\SB4_25/i0[10] ), .A2(
        \SB4_25/i0_4 ), .A3(\SB4_25/i0_3 ), .ZN(
        \SB4_25/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB4_25/Component_Function_0/N2  ( .A1(\SB4_25/i0[8] ), .A2(
        \SB4_25/i0[7] ), .A3(\SB4_25/i0[6] ), .ZN(
        \SB4_25/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB4_25/Component_Function_1/N4  ( .A1(\SB4_25/i1_7 ), .A2(
        \SB4_25/i0[8] ), .A3(\SB4_25/i0_4 ), .ZN(
        \SB4_25/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_25/Component_Function_1/N2  ( .A1(\SB4_25/i0_3 ), .A2(
        \SB4_25/i1_7 ), .A3(\SB4_25/i0[8] ), .ZN(
        \SB4_25/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB4_25/Component_Function_5/N4  ( .A1(\SB4_25/i0[9] ), .A2(
        \SB4_25/i0[6] ), .A3(\SB4_25/i0_4 ), .ZN(
        \SB4_25/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB4_25/Component_Function_5/N1  ( .A1(\SB4_25/i0_0 ), .A2(
        \SB4_25/i3[0] ), .ZN(\SB4_25/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_26/Component_Function_0/N2  ( .A1(\SB4_26/i0[8] ), .A2(
        \SB4_26/i0[7] ), .A3(\SB4_26/i0[6] ), .ZN(
        \SB4_26/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB4_26/Component_Function_1/N4  ( .A1(\SB4_26/i1_7 ), .A2(
        \SB4_26/i0[8] ), .A3(\SB4_26/i0_4 ), .ZN(
        \SB4_26/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_26/Component_Function_1/N2  ( .A1(\SB4_26/i0_3 ), .A2(
        \SB4_26/i1_7 ), .A3(\SB4_26/i0[8] ), .ZN(
        \SB4_26/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_26/Component_Function_1/N1  ( .A1(\SB4_26/i0_3 ), .A2(
        \SB4_26/i1[9] ), .ZN(\SB4_26/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_26/Component_Function_5/N3  ( .A1(\SB4_26/i1[9] ), .A2(
        \SB4_26/i0_4 ), .A3(\SB4_26/i0_3 ), .ZN(
        \SB4_26/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 \SB4_26/Component_Function_5/N1  ( .A1(\SB4_26/i0_0 ), .A2(
        \SB4_26/i3[0] ), .ZN(\SB4_26/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_27/Component_Function_0/N2  ( .A1(\SB4_27/i0[8] ), .A2(
        \SB4_27/i0[7] ), .A3(\SB4_27/i0[6] ), .ZN(
        \SB4_27/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB4_27/Component_Function_1/N4  ( .A1(\SB4_27/i1_7 ), .A2(
        \SB4_27/i0[8] ), .A3(\SB4_27/i0_4 ), .ZN(
        \SB4_27/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_27/Component_Function_1/N2  ( .A1(\SB4_27/i0_3 ), .A2(
        \SB4_27/i1_7 ), .A3(\SB4_27/i0[8] ), .ZN(
        \SB4_27/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB4_27/Component_Function_5/N2  ( .A1(n2898), .A2(\SB4_27/i0[6] ), 
        .A3(\SB4_27/i0[10] ), .ZN(\SB4_27/Component_Function_5/NAND4_in[1] )
         );
  NAND2_X1 \SB4_27/Component_Function_5/N1  ( .A1(n2898), .A2(\SB4_27/i3[0] ), 
        .ZN(\SB4_27/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_28/Component_Function_1/N4  ( .A1(\SB4_28/i1_7 ), .A2(
        \SB4_28/i0[8] ), .A3(\SB4_28/i0_4 ), .ZN(
        \SB4_28/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_28/Component_Function_1/N3  ( .A1(\SB4_28/i1_5 ), .A2(
        \SB4_28/i0[6] ), .A3(\SB4_28/i0[9] ), .ZN(
        \SB4_28/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_28/Component_Function_1/N2  ( .A1(\SB4_28/i0_3 ), .A2(
        \SB4_28/i1_7 ), .A3(\SB4_28/i0[8] ), .ZN(
        \SB4_28/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_28/Component_Function_5/N1  ( .A1(\SB4_28/i0_0 ), .A2(
        \SB4_28/i3[0] ), .ZN(\SB4_28/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB4_29/Component_Function_1/N2  ( .A1(\SB4_29/i0_3 ), .A2(
        \SB4_29/i1_7 ), .A3(\SB4_29/i0[8] ), .ZN(
        \SB4_29/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_29/Component_Function_1/N1  ( .A1(\SB4_29/i0_3 ), .A2(
        \SB4_29/i1[9] ), .ZN(\SB4_29/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_31/Component_Function_1/N4  ( .A1(\SB4_31/i1_7 ), .A2(n3652), 
        .A3(\SB4_31/i0_4 ), .ZN(\SB4_31/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB4_31/Component_Function_1/N3  ( .A1(\SB4_31/i1_5 ), .A2(
        \SB4_31/i0[6] ), .A3(\SB4_31/i0[9] ), .ZN(
        \SB4_31/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_31/Component_Function_1/N2  ( .A1(\SB4_31/i0_3 ), .A2(
        \SB4_31/i1_7 ), .A3(n3652), .ZN(
        \SB4_31/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB4_31/Component_Function_1/N1  ( .A1(\SB4_31/i0_3 ), .A2(
        \SB4_31/i1[9] ), .ZN(\SB4_31/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB4_31/Component_Function_5/N3  ( .A1(\SB4_31/i1[9] ), .A2(
        \SB4_31/i0_4 ), .A3(\SB4_31/i0_3 ), .ZN(
        \SB4_31/Component_Function_5/NAND4_in[2] ) );
  BUF_X4 \SB2_0_31/BUF_5  ( .I(\RI3[0][5] ), .Z(\SB2_0_31/i0_3 ) );
  BUF_X4 \SB2_1_22/BUF_5  ( .I(\SB1_1_22/buf_output[5] ), .Z(\SB2_1_22/i0_3 )
         );
  BUF_X4 \SB1_2_0/BUF_5  ( .I(\MC_ARK_ARC_1_1/buf_output[191] ), .Z(
        \SB1_2_0/i0_3 ) );
  BUF_X4 \SB1_2_5/BUF_5  ( .I(\MC_ARK_ARC_1_1/buf_output[161] ), .Z(
        \SB1_2_5/i0_3 ) );
  BUF_X4 \SB1_2_10/BUF_5  ( .I(\MC_ARK_ARC_1_1/buf_output[131] ), .Z(
        \SB1_2_10/i0_3 ) );
  BUF_X4 \SB1_2_12/BUF_5  ( .I(\MC_ARK_ARC_1_1/buf_output[119] ), .Z(
        \SB1_2_12/i0_3 ) );
  BUF_X4 \SB2_2_9/BUF_5  ( .I(\SB1_2_9/buf_output[5] ), .Z(\SB2_2_9/i0_3 ) );
  BUF_X4 \SB1_3_1/BUF_5  ( .I(\MC_ARK_ARC_1_2/buf_output[185] ), .Z(
        \SB1_3_1/i0_3 ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_38  ( .I(\SB2_3_28/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[38] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_74  ( .I(\SB2_2_22/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[74] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_86  ( .I(\SB2_0_20/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[86] ) );
  INV_X2 \SB2_0_12/INV_2  ( .I(\RI3[0][116] ), .ZN(\SB2_0_12/i1[9] ) );
  INV_X2 \SB1_2_22/INV_5  ( .I(\RI1[2][59] ), .ZN(\SB1_2_22/i1_5 ) );
  INV_X2 \SB1_2_20/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[68] ), .ZN(
        \SB1_2_20/i1[9] ) );
  INV_X2 \SB1_2_0/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[188] ), .ZN(
        \SB1_2_0/i1[9] ) );
  INV_X2 \SB1_3_25/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[38] ), .ZN(
        \SB1_3_25/i1[9] ) );
  INV_X2 \SB2_1_18/INV_2  ( .I(\SB1_1_21/buf_output[2] ), .ZN(\SB2_1_18/i1[9] ) );
  INV_X2 \SB1_2_6/INV_3  ( .I(n5522), .ZN(\SB1_2_6/i0[8] ) );
  BUF_X4 \SB1_2_3/BUF_5  ( .I(\MC_ARK_ARC_1_1/buf_output[173] ), .Z(
        \SB1_2_3/i0_3 ) );
  INV_X2 \SB2_0_0/INV_2  ( .I(\RI3[0][188] ), .ZN(\SB2_0_0/i1[9] ) );
  INV_X2 \SB1_1_20/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[68] ), .ZN(
        \SB1_1_20/i1[9] ) );
  INV_X2 \SB1_1_0/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[189] ), .ZN(
        \SB1_1_0/i0[8] ) );
  INV_X2 \SB1_2_25/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[38] ), .ZN(
        \SB1_2_25/i1[9] ) );
  INV_X2 \SB1_3_15/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[98] ), .ZN(
        \SB1_3_15/i1[9] ) );
  INV_X2 \SB3_7/INV_3  ( .I(n3646), .ZN(\SB3_7/i0[8] ) );
  INV_X2 \SB1_1_20/INV_5  ( .I(\RI1[1][71] ), .ZN(\SB1_1_20/i1_5 ) );
  BUF_X4 \SB1_2_23/BUF_5  ( .I(\MC_ARK_ARC_1_1/buf_output[53] ), .Z(
        \SB1_2_23/i0_3 ) );
  BUF_X4 \SB1_3_28/BUF_5  ( .I(\MC_ARK_ARC_1_2/buf_output[23] ), .Z(
        \SB1_3_28/i0_3 ) );
  BUF_X4 \SB1_3_9/BUF_5  ( .I(\MC_ARK_ARC_1_2/buf_output[137] ), .Z(
        \SB1_3_9/i0_3 ) );
  INV_X2 \SB1_2_17/INV_2  ( .I(n5523), .ZN(\SB1_2_17/i1[9] ) );
  INV_X2 \SB1_2_1/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[183] ), .ZN(
        \SB1_2_1/i0[8] ) );
  BUF_X4 \SB2_3_29/BUF_5  ( .I(\SB1_3_29/buf_output[5] ), .Z(\SB2_3_29/i0_3 )
         );
  INV_X2 \SB1_3_10/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[128] ), .ZN(
        \SB1_3_10/i1[9] ) );
  INV_X2 \SB1_3_11/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[123] ), .ZN(
        \SB1_3_11/i0[8] ) );
  INV_X2 \SB1_3_26/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[33] ), .ZN(
        \SB1_3_26/i0[8] ) );
  INV_X2 \SB1_2_24/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[44] ), .ZN(
        \SB1_2_24/i1[9] ) );
  BUF_X2 \SB1_0_20/BUF_1  ( .I(n279), .Z(\SB1_0_20/i0[6] ) );
  INV_X2 \SB1_2_5/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[159] ), .ZN(
        \SB1_2_5/i0[8] ) );
  INV_X2 \SB1_3_31/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[2] ), .ZN(
        \SB1_3_31/i1[9] ) );
  INV_X2 \SB1_2_14/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[105] ), .ZN(
        \SB1_2_14/i0[8] ) );
  INV_X2 \SB2_3_10/INV_2  ( .I(\SB1_3_13/buf_output[2] ), .ZN(\SB2_3_10/i1[9] ) );
  INV_X2 \SB1_3_3/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[170] ), .ZN(
        \SB1_3_3/i1[9] ) );
  INV_X2 \SB3_15/INV_5  ( .I(\MC_ARK_ARC_1_3/buf_output[101] ), .ZN(
        \SB3_15/i1_5 ) );
  INV_X2 \SB2_0_25/INV_2  ( .I(\SB1_0_28/buf_output[2] ), .ZN(\SB2_0_25/i1[9] ) );
  INV_X2 \SB1_2_6/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[152] ), .ZN(
        \SB1_2_6/i1[9] ) );
  INV_X2 \SB1_1_27/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[27] ), .ZN(
        \SB1_1_27/i0[8] ) );
  INV_X2 \SB2_3_0/INV_2  ( .I(\SB1_3_3/buf_output[2] ), .ZN(\SB2_3_0/i1[9] )
         );
  INV_X2 \SB1_0_13/INV_2  ( .I(n301), .ZN(\SB1_0_13/i1[9] ) );
  INV_X2 \SB2_0_21/INV_2  ( .I(\RI3[0][62] ), .ZN(\SB2_0_21/i1[9] ) );
  INV_X2 \SB1_3_7/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[147] ), .ZN(
        \SB1_3_7/i0[8] ) );
  INV_X2 \SB1_1_9/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[134] ), .ZN(
        \SB1_1_9/i1[9] ) );
  BUF_X4 \SB1_1_21/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[65] ), .Z(
        \SB1_1_21/i0_3 ) );
  INV_X2 \SB2_0_22/INV_5  ( .I(\SB1_0_22/buf_output[5] ), .ZN(\SB2_0_22/i1_5 )
         );
  INV_X2 \SB1_3_5/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[158] ), .ZN(
        \SB1_3_5/i1[9] ) );
  INV_X2 \SB3_31/INV_3  ( .I(\MC_ARK_ARC_1_3/buf_output[3] ), .ZN(
        \SB3_31/i0[8] ) );
  NAND3_X1 \SB2_1_12/Component_Function_0/N4  ( .A1(\SB2_1_12/i0[7] ), .A2(
        \SB2_1_12/i0_3 ), .A3(\SB2_1_12/i0_0 ), .ZN(
        \SB2_1_12/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_27/Component_Function_4/N3  ( .A1(\SB1_1_27/i0[9] ), .A2(
        \SB1_1_27/i0[10] ), .A3(\SB1_1_27/i0_3 ), .ZN(
        \SB1_1_27/Component_Function_4/NAND4_in[2] ) );
  NAND4_X2 \SB1_0_15/Component_Function_5/N5  ( .A1(
        \SB1_0_15/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_0_15/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_15/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_0_15/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB1_0_15/buf_output[5] ) );
  NAND4_X2 \SB1_2_22/Component_Function_4/N5  ( .A1(
        \SB1_2_22/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_22/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_22/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_22/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_2_22/buf_output[4] ) );
  INV_X2 \SB1_1_8/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[141] ), .ZN(
        \SB1_1_8/i0[8] ) );
  INV_X2 \SB1_1_25/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[38] ), .ZN(
        \SB1_1_25/i1[9] ) );
  INV_X2 \SB1_1_7/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[146] ), .ZN(
        \SB1_1_7/i1[9] ) );
  BUF_X4 \SB2_3_2/BUF_5  ( .I(\SB1_3_2/buf_output[5] ), .Z(\SB2_3_2/i0_3 ) );
  NAND4_X2 \SB3_3/Component_Function_0/N5  ( .A1(
        \SB3_3/Component_Function_0/NAND4_in[0] ), .A2(
        \SB3_3/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_3/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_3/Component_Function_0/NAND4_in[3] ), .ZN(\SB3_3/buf_output[0] )
         );
  INV_X2 \SB1_2_4/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[164] ), .ZN(
        \SB1_2_4/i1[9] ) );
  INV_X2 \SB2_2_27/INV_2  ( .I(\SB1_2_30/buf_output[2] ), .ZN(\SB2_2_27/i1[9] ) );
  INV_X2 \SB3_7/INV_2  ( .I(\MC_ARK_ARC_1_3/buf_output[146] ), .ZN(
        \SB3_7/i1[9] ) );
  NAND3_X2 \SB1_3_2/Component_Function_5/N3  ( .A1(\SB1_3_2/i1[9] ), .A2(
        \SB1_3_2/i0_4 ), .A3(\SB1_3_2/i0_3 ), .ZN(
        \SB1_3_2/Component_Function_5/NAND4_in[2] ) );
  BUF_X4 \SB2_1_12/BUF_5  ( .I(\SB1_1_12/buf_output[5] ), .Z(\SB2_1_12/i0_3 )
         );
  INV_X2 \SB4_2/INV_5  ( .I(\SB3_2/buf_output[5] ), .ZN(\SB4_2/i1_5 ) );
  INV_X2 \SB1_1_0/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[188] ), .ZN(
        \SB1_1_0/i1[9] ) );
  NAND3_X2 \SB1_0_15/Component_Function_5/N3  ( .A1(\SB1_0_15/i1[9] ), .A2(
        \SB1_0_15/i0_4 ), .A3(\SB1_0_15/i0_3 ), .ZN(
        \SB1_0_15/Component_Function_5/NAND4_in[2] ) );
  INV_X2 \SB1_1_15/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[98] ), .ZN(
        \SB1_1_15/i1[9] ) );
  INV_X2 \SB1_1_13/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[110] ), .ZN(
        \SB1_1_13/i1[9] ) );
  INV_X2 \SB1_3_8/INV_5  ( .I(\RI1[3][143] ), .ZN(\SB1_3_8/i1_5 ) );
  INV_X2 \SB1_3_26/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[32] ), .ZN(
        \SB1_3_26/i1[9] ) );
  BUF_X2 \SB1_0_27/BUF_0  ( .I(n257), .Z(\SB1_0_27/i0[9] ) );
  INV_X2 \SB1_3_16/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[92] ), .ZN(
        \SB1_3_16/i1[9] ) );
  INV_X2 \SB2_1_12/INV_5  ( .I(\SB1_1_12/buf_output[5] ), .ZN(\SB2_1_12/i1_5 )
         );
  INV_X2 \SB1_1_3/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[170] ), .ZN(
        \SB1_1_3/i1[9] ) );
  INV_X2 \SB1_0_15/INV_2  ( .I(n295), .ZN(\SB1_0_15/i1[9] ) );
  BUF_X2 \SB1_0_4/BUF_1  ( .I(n327), .Z(\SB1_0_4/i0[6] ) );
  INV_X2 \SB1_2_29/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[14] ), .ZN(
        \SB1_2_29/i1[9] ) );
  INV_X2 \SB3_30/INV_5  ( .I(n5509), .ZN(\SB3_30/i1_5 ) );
  INV_X2 \SB2_0_3/INV_5  ( .I(\SB1_0_3/buf_output[5] ), .ZN(\SB2_0_3/i1_5 ) );
  INV_X2 \SB1_0_20/INV_2  ( .I(n280), .ZN(\SB1_0_20/i1[9] ) );
  CLKBUF_X8 \SB1_2_4/BUF_5  ( .I(\RI1[2][167] ), .Z(\SB1_2_4/i0_3 ) );
  BUF_X2 \SB1_0_22/BUF_1  ( .I(n273), .Z(\SB1_0_22/i0[6] ) );
  INV_X2 \SB3_16/INV_2  ( .I(\MC_ARK_ARC_1_3/buf_output[92] ), .ZN(
        \SB3_16/i1[9] ) );
  INV_X2 \SB2_2_15/INV_2  ( .I(\SB1_2_18/buf_output[2] ), .ZN(\SB2_2_15/i1[9] ) );
  BUF_X2 \SB1_0_1/BUF_0  ( .I(n335), .Z(\SB1_0_1/i0[9] ) );
  NAND4_X1 \SB2_1_30/Component_Function_3/N5  ( .A1(
        \SB2_1_30/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_30/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_30/Component_Function_3/NAND4_in[3] ), .A4(
        \SB2_1_30/Component_Function_3/NAND4_in[2] ), .ZN(
        \SB2_1_30/buf_output[3] ) );
  INV_X2 \SB1_1_21/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[62] ), .ZN(
        \SB1_1_21/i1[9] ) );
  INV_X2 \SB1_1_23/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[50] ), .ZN(
        \SB1_1_23/i1[9] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_155  ( .I(\SB2_3_6/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[155] ) );
  INV_X2 \SB1_1_31/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[2] ), .ZN(
        \SB1_1_31/i1[9] ) );
  INV_X2 \SB2_1_9/INV_2  ( .I(\SB1_1_12/buf_output[2] ), .ZN(\SB2_1_9/i1[9] )
         );
  BUF_X2 \SB1_0_11/BUF_1  ( .I(n306), .Z(\SB1_0_11/i0[6] ) );
  BUF_X2 \SB1_0_7/BUF_1  ( .I(n318), .Z(\SB1_0_7/i0[6] ) );
  INV_X2 \SB2_2_4/INV_5  ( .I(\SB1_2_4/buf_output[5] ), .ZN(\SB2_2_4/i1_5 ) );
  INV_X2 \SB1_1_19/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[74] ), .ZN(
        \SB1_1_19/i1[9] ) );
  INV_X2 \SB1_0_25/INV_2  ( .I(n265), .ZN(\SB1_0_25/i1[9] ) );
  INV_X2 \SB2_3_3/INV_5  ( .I(\SB1_3_3/buf_output[5] ), .ZN(\SB2_3_3/i1_5 ) );
  INV_X2 \SB1_2_23/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[50] ), .ZN(
        \SB1_2_23/i1[9] ) );
  INV_X2 \SB2_3_4/INV_2  ( .I(\SB1_3_7/buf_output[2] ), .ZN(\SB2_3_4/i1[9] )
         );
  INV_X2 \SB1_1_28/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[23] ), .ZN(
        \SB1_1_28/i1_5 ) );
  INV_X2 \SB1_3_2/INV_5  ( .I(\MC_ARK_ARC_1_2/buf_output[179] ), .ZN(
        \SB1_3_2/i1_5 ) );
  INV_X2 \SB4_11/INV_2  ( .I(\SB3_14/buf_output[2] ), .ZN(\SB4_11/i1[9] ) );
  INV_X2 \SB1_2_26/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[32] ), .ZN(
        \SB1_2_26/i1[9] ) );
  INV_X2 \SB1_1_5/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[158] ), .ZN(
        \SB1_1_5/i1[9] ) );
  INV_X2 \SB1_1_3/INV_5  ( .I(\RI1[1][173] ), .ZN(\SB1_1_3/i1_5 ) );
  INV_X2 \SB3_26/INV_2  ( .I(n1384), .ZN(\SB3_26/i1[9] ) );
  INV_X2 \SB1_2_21/INV_3  ( .I(\MC_ARK_ARC_1_1/buf_output[63] ), .ZN(
        \SB1_2_21/i0[8] ) );
  INV_X2 \SB1_1_4/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[164] ), .ZN(
        \SB1_1_4/i1[9] ) );
  INV_X2 \SB1_2_12/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[116] ), .ZN(
        \SB1_2_12/i1[9] ) );
  INV_X2 \SB1_3_23/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[50] ), .ZN(
        \SB1_3_23/i1[9] ) );
  INV_X2 \SB1_3_11/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[122] ), .ZN(
        \SB1_3_11/i1[9] ) );
  INV_X2 \SB1_3_18/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[80] ), .ZN(
        \SB1_3_18/i1[9] ) );
  NAND4_X2 \SB2_3_3/Component_Function_0/N5  ( .A1(
        \SB2_3_3/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_3_3/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_3/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_3/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB2_3_3/buf_output[0] ) );
  INV_X2 \SB1_1_6/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[152] ), .ZN(
        \SB1_1_6/i1[9] ) );
  INV_X2 \SB2_1_2/INV_5  ( .I(\SB1_1_2/buf_output[5] ), .ZN(\SB2_1_2/i1_5 ) );
  INV_X2 \SB1_1_18/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[80] ), .ZN(
        \SB1_1_18/i1[9] ) );
  INV_X2 \SB1_3_2/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[176] ), .ZN(
        \SB1_3_2/i1[9] ) );
  INV_X2 \SB2_2_29/INV_2  ( .I(\SB1_2_0/buf_output[2] ), .ZN(\SB2_2_29/i1[9] )
         );
  INV_X2 \SB1_3_12/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[116] ), .ZN(
        \SB1_3_12/i1[9] ) );
  NAND3_X1 \SB3_1/Component_Function_4/N3  ( .A1(\SB3_1/i0[9] ), .A2(
        \SB3_1/i0[10] ), .A3(\SB3_1/i0_3 ), .ZN(
        \SB3_1/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB4_6/Component_Function_1/N3  ( .A1(\SB4_6/i1_5 ), .A2(
        \SB4_6/i0[6] ), .A3(\SB4_6/i0[9] ), .ZN(
        \SB4_6/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_22/Component_Function_3/N2  ( .A1(\SB1_2_22/i0_0 ), .A2(
        \SB1_2_22/i0_3 ), .A3(\SB1_2_22/i0_4 ), .ZN(
        \SB1_2_22/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_18/Component_Function_4/N1  ( .A1(\SB2_0_18/i0[9] ), .A2(
        \SB2_0_18/i0_0 ), .A3(\SB2_0_18/i0[8] ), .ZN(
        \SB2_0_18/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_30/Component_Function_2/N4  ( .A1(\SB2_0_30/i1_5 ), .A2(
        \SB2_0_30/i0_0 ), .A3(\RI3[0][10] ), .ZN(
        \SB2_0_30/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_18/Component_Function_2/N4  ( .A1(\SB1_0_18/i1_5 ), .A2(
        \SB1_0_18/i0_0 ), .A3(n4753), .ZN(
        \SB1_0_18/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_15/Component_Function_3/N1  ( .A1(\SB1_0_15/i1[9] ), .A2(
        \SB1_0_15/i0_3 ), .A3(\SB1_0_15/i0[6] ), .ZN(
        \SB1_0_15/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_24/Component_Function_1/N3  ( .A1(\SB1_0_24/i1_5 ), .A2(
        \SB1_0_24/i0[6] ), .A3(\SB1_0_24/i0[9] ), .ZN(
        \SB1_0_24/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB4_0/Component_Function_4/N3  ( .A1(\SB4_0/i0[9] ), .A2(
        \SB4_0/i0[10] ), .A3(\SB4_0/i0_3 ), .ZN(
        \SB4_0/Component_Function_4/NAND4_in[2] ) );
  BUF_X2 \SB1_0_27/BUF_3  ( .I(n349), .Z(\SB1_0_27/i0[10] ) );
  NAND3_X1 \SB1_0_15/Component_Function_3/N2  ( .A1(\SB1_0_15/i0_0 ), .A2(
        \SB1_0_15/i0_3 ), .A3(\SB1_0_15/i0_4 ), .ZN(
        \SB1_0_15/Component_Function_3/NAND4_in[1] ) );
  INV_X2 \SB1_2_31/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[2] ), .ZN(
        \SB1_2_31/i1[9] ) );
  INV_X1 \SB1_0_27/INV_3  ( .I(n349), .ZN(\SB1_0_27/i0[8] ) );
  INV_X2 \SB1_2_10/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[128] ), .ZN(
        \SB1_2_10/i1[9] ) );
  INV_X1 \SB1_0_15/INV_5  ( .I(n421), .ZN(\SB1_0_15/i1_5 ) );
  INV_X2 \SB1_2_21/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[62] ), .ZN(
        \SB1_2_21/i1[9] ) );
  INV_X2 \SB3_13/INV_2  ( .I(n3688), .ZN(\SB3_13/i1[9] ) );
  BUF_X4 \SB2_0_23/BUF_5  ( .I(\SB1_0_23/buf_output[5] ), .Z(\SB2_0_23/i0_3 )
         );
  INV_X2 \SB1_0_25/INV_3  ( .I(n353), .ZN(\SB1_0_25/i0[8] ) );
  INV_X2 \SB2_1_25/INV_5  ( .I(\SB1_1_25/buf_output[5] ), .ZN(\SB2_1_25/i1_5 )
         );
  INV_X2 \SB2_3_12/INV_2  ( .I(\SB1_3_15/buf_output[2] ), .ZN(\SB2_3_12/i1[9] ) );
  INV_X2 \SB2_2_23/INV_5  ( .I(\SB1_2_23/buf_output[5] ), .ZN(\SB2_2_23/i1_5 )
         );
  INV_X2 \SB1_1_26/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[35] ), .ZN(
        \SB1_1_26/i1_5 ) );
  NAND3_X2 \SB1_3_6/Component_Function_5/N4  ( .A1(\SB1_3_6/i0[9] ), .A2(
        \SB1_3_6/i0[6] ), .A3(\SB1_3_6/i0_4 ), .ZN(
        \SB1_3_6/Component_Function_5/NAND4_in[3] ) );
  INV_X2 \SB1_3_17/INV_2  ( .I(n5524), .ZN(\SB1_3_17/i1[9] ) );
  INV_X2 \SB3_21/INV_3  ( .I(n5520), .ZN(\SB3_21/i0[8] ) );
  NAND4_X2 \SB3_29/Component_Function_4/N5  ( .A1(
        \SB3_29/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_29/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_29/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_29/Component_Function_4/NAND4_in[3] ), .ZN(\SB3_29/buf_output[4] ) );
  INV_X2 \SB2_2_20/INV_5  ( .I(\SB1_2_20/buf_output[5] ), .ZN(\SB2_2_20/i1_5 )
         );
  INV_X2 \SB1_1_15/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[101] ), .ZN(
        \SB1_1_15/i1_5 ) );
  INV_X2 \SB2_3_16/INV_5  ( .I(\SB1_3_16/buf_output[5] ), .ZN(\SB2_3_16/i1_5 )
         );
  INV_X2 \SB3_21/INV_2  ( .I(\MC_ARK_ARC_1_3/buf_output[62] ), .ZN(
        \SB3_21/i1[9] ) );
  INV_X2 \SB1_3_31/INV_5  ( .I(\RI1[3][5] ), .ZN(\SB1_3_31/i1_5 ) );
  BUF_X2 \SB1_0_26/BUF_1  ( .I(n261), .Z(\SB1_0_26/i0[6] ) );
  CLKBUF_X4 \SB1_0_1/BUF_4  ( .I(n402), .Z(\SB1_0_1/i0_4 ) );
  BUF_X2 \SB1_0_13/BUF_0  ( .I(n299), .Z(\SB1_0_13/i0[9] ) );
  BUF_X2 \SB1_0_14/BUF_1  ( .I(n297), .Z(\SB1_0_14/i0[6] ) );
  CLKBUF_X4 \SB1_0_8/BUF_2  ( .I(n316), .Z(\SB1_0_8/i0_0 ) );
  BUF_X2 \SB1_0_8/BUF_0  ( .I(n314), .Z(\SB1_0_8/i0[9] ) );
  BUF_X2 \SB1_0_15/BUF_1  ( .I(n294), .Z(\SB1_0_15/i0[6] ) );
  BUF_X2 \SB1_0_15/BUF_0  ( .I(n293), .Z(\SB1_0_15/i0[9] ) );
  BUF_X2 \SB1_0_30/BUF_1  ( .I(n249), .Z(\SB1_0_30/i0[6] ) );
  BUF_X2 \SB1_0_30/BUF_0  ( .I(n248), .Z(\SB1_0_30/i0[9] ) );
  CLKBUF_X4 \SB1_0_15/BUF_2  ( .I(n295), .Z(\SB1_0_15/i0_0 ) );
  CLKBUF_X4 \SB1_0_6/BUF_4  ( .I(n392), .Z(\SB1_0_6/i0_4 ) );
  BUF_X2 \SB1_0_20/BUF_0  ( .I(n278), .Z(\SB1_0_20/i0[9] ) );
  BUF_X2 \SB1_0_24/BUF_1  ( .I(n267), .Z(\SB1_0_24/i0[6] ) );
  BUF_X2 \SB1_0_9/BUF_0  ( .I(n311), .Z(\SB1_0_9/i0[9] ) );
  BUF_X2 \SB1_0_21/BUF_0  ( .I(n275), .Z(\SB1_0_21/i0[9] ) );
  BUF_X2 \SB1_0_24/BUF_0  ( .I(n266), .Z(\SB1_0_24/i0[9] ) );
  BUF_X2 \SB1_0_19/BUF_1  ( .I(n282), .Z(\SB1_0_19/i0[6] ) );
  CLKBUF_X4 \SB1_0_31/BUF_4  ( .I(n342), .Z(\SB1_0_31/i0_4 ) );
  BUF_X2 \SB1_0_10/BUF_0  ( .I(n308), .Z(\SB1_0_10/i0[9] ) );
  CLKBUF_X4 \SB1_0_12/BUF_4  ( .I(n380), .Z(\SB1_0_12/i0_4 ) );
  CLKBUF_X4 \SB1_0_20/BUF_2  ( .I(n280), .Z(\SB1_0_20/i0_0 ) );
  NAND3_X1 \SB1_0_1/Component_Function_5/N4  ( .A1(\SB1_0_1/i0[9] ), .A2(
        \SB1_0_1/i0[6] ), .A3(\SB1_0_1/i0_4 ), .ZN(
        \SB1_0_1/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_9/Component_Function_1/N3  ( .A1(\SB1_0_9/i1_5 ), .A2(
        \SB1_0_9/i0[6] ), .A3(\SB1_0_9/i0[9] ), .ZN(
        \SB1_0_9/Component_Function_1/NAND4_in[2] ) );
  CLKBUF_X4 \SB2_0_10/BUF_2  ( .I(\SB1_0_13/buf_output[2] ), .Z(
        \SB2_0_10/i0_0 ) );
  CLKBUF_X4 \SB2_0_6/BUF_2  ( .I(\RI3[0][152] ), .Z(\SB2_0_6/i0_0 ) );
  CLKBUF_X4 \SB2_0_11/BUF_2  ( .I(\SB1_0_14/buf_output[2] ), .Z(
        \SB2_0_11/i0_0 ) );
  BUF_X4 \SB2_0_22/BUF_5  ( .I(\SB1_0_22/buf_output[5] ), .Z(\SB2_0_22/i0_3 )
         );
  CLKBUF_X4 \SB2_0_15/BUF_2  ( .I(\SB1_0_18/buf_output[2] ), .Z(
        \SB2_0_15/i0_0 ) );
  CLKBUF_X4 \SB2_0_8/BUF_3  ( .I(\SB1_0_10/buf_output[3] ), .Z(
        \SB2_0_8/i0[10] ) );
  CLKBUF_X4 \SB2_0_8/BUF_2  ( .I(\SB1_0_11/buf_output[2] ), .Z(\SB2_0_8/i0_0 )
         );
  CLKBUF_X4 \SB2_0_12/BUF_3  ( .I(\SB1_0_14/buf_output[3] ), .Z(
        \SB2_0_12/i0[10] ) );
  CLKBUF_X4 \SB2_0_4/BUF_2  ( .I(\RI3[0][164] ), .Z(\SB2_0_4/i0_0 ) );
  CLKBUF_X4 \SB2_0_24/BUF_3  ( .I(\RI3[0][45] ), .Z(\SB2_0_24/i0[10] ) );
  CLKBUF_X4 \SB2_0_30/BUF_1  ( .I(\RI3[0][7] ), .Z(\SB2_0_30/i0[6] ) );
  CLKBUF_X4 \SB2_0_19/BUF_2  ( .I(\SB1_0_22/buf_output[2] ), .Z(
        \SB2_0_19/i0_0 ) );
  CLKBUF_X4 \SB2_0_25/BUF_0  ( .I(\SB1_0_30/buf_output[0] ), .Z(
        \SB2_0_25/i0[9] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_82  ( .I(\SB2_0_19/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[82] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_179  ( .I(\SB2_0_2/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[179] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_61  ( .I(\SB2_0_25/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[61] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_155  ( .I(\SB2_0_6/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[155] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_90  ( .I(\SB2_0_21/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[90] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_138  ( .I(\SB2_0_13/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[138] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_42  ( .I(\SB2_0_29/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[42] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_44  ( .I(\SB2_0_27/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[44] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_167  ( .I(\SB2_0_4/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[167] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_48  ( .I(\SB2_0_28/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[48] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_36  ( .I(\SB2_0_30/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[36] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_78  ( .I(\SB2_0_23/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[78] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_144  ( .I(\SB2_0_12/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[144] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_88  ( .I(\SB2_0_18/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[88] ) );
  BUF_X4 \SB1_1_14/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[107] ), .Z(
        \SB1_1_14/i0_3 ) );
  BUF_X4 \SB1_1_28/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[23] ), .Z(
        \SB1_1_28/i0_3 ) );
  CLKBUF_X4 \SB1_1_31/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[0] ), .Z(
        \SB1_1_31/i0[9] ) );
  BUF_X4 \SB1_1_1/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[185] ), .Z(
        \SB1_1_1/i0_3 ) );
  CLKBUF_X4 \SB1_1_25/BUF_2  ( .I(\MC_ARK_ARC_1_0/buf_output[38] ), .Z(
        \SB1_1_25/i0_0 ) );
  CLKBUF_X4 \SB1_1_5/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[156] ), .Z(
        \SB1_1_5/i0[9] ) );
  NAND3_X1 \SB1_1_16/Component_Function_1/N3  ( .A1(\SB1_1_16/i1_5 ), .A2(
        \SB1_1_16/i0[6] ), .A3(\SB1_1_16/i0[9] ), .ZN(
        \SB1_1_16/Component_Function_1/NAND4_in[2] ) );
  CLKBUF_X4 \SB2_1_16/BUF_3  ( .I(\SB1_1_18/buf_output[3] ), .Z(
        \SB2_1_16/i0[10] ) );
  CLKBUF_X4 \SB2_1_25/BUF_2  ( .I(\SB1_1_28/buf_output[2] ), .Z(
        \SB2_1_25/i0_0 ) );
  CLKBUF_X4 \SB2_1_11/BUF_1  ( .I(\SB1_1_15/buf_output[1] ), .Z(
        \SB2_1_11/i0[6] ) );
  CLKBUF_X4 \SB2_1_31/BUF_2  ( .I(\SB1_1_2/buf_output[2] ), .Z(\SB2_1_31/i0_0 ) );
  CLKBUF_X4 \SB2_1_31/BUF_3  ( .I(\SB1_1_1/buf_output[3] ), .Z(
        \SB2_1_31/i0[10] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_25  ( .I(\SB2_1_31/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[25] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_101  ( .I(\SB2_1_15/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[101] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_179  ( .I(\SB2_1_2/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[179] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_38  ( .I(\SB2_1_28/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[38] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_29  ( .I(\SB2_1_27/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[29] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_186  ( .I(\SB2_1_5/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[186] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_169  ( .I(\SB2_1_7/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[169] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_160  ( .I(\SB2_1_6/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[160] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_42  ( .I(\SB2_1_29/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[42] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_84  ( .I(\SB2_1_22/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[84] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_9  ( .I(\SB2_1_0/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[9] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_100  ( .I(\SB2_1_16/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[100] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_28  ( .I(\SB2_1_28/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[28] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_187  ( .I(\SB2_1_4/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[187] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_159  ( .I(\SB2_1_7/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[159] ) );
  CLKBUF_X4 \SB1_2_18/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[79] ), .Z(
        \SB1_2_18/i0[6] ) );
  BUF_X4 \SB1_2_27/BUF_5  ( .I(\MC_ARK_ARC_1_1/buf_output[29] ), .Z(
        \SB1_2_27/i0_3 ) );
  CLKBUF_X4 \SB1_2_8/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[138] ), .Z(
        \SB1_2_8/i0[9] ) );
  NAND3_X1 \SB1_2_23/Component_Function_1/N4  ( .A1(\SB1_2_23/i1_7 ), .A2(
        \SB1_2_23/i0[8] ), .A3(\MC_ARK_ARC_1_1/buf_output[52] ), .ZN(
        \SB1_2_23/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_27/Component_Function_1/N3  ( .A1(\SB1_2_27/i1_5 ), .A2(
        \SB1_2_27/i0[6] ), .A3(\SB1_2_27/i0[9] ), .ZN(
        \SB1_2_27/Component_Function_1/NAND4_in[2] ) );
  CLKBUF_X4 \SB2_2_18/BUF_0  ( .I(\SB1_2_23/buf_output[0] ), .Z(
        \SB2_2_18/i0[9] ) );
  CLKBUF_X4 \SB2_2_31/BUF_2  ( .I(\SB1_2_2/buf_output[2] ), .Z(\SB2_2_31/i0_0 ) );
  CLKBUF_X4 \SB2_2_6/BUF_3  ( .I(\SB1_2_8/buf_output[3] ), .Z(\SB2_2_6/i0[10] ) );
  CLKBUF_X4 \SB2_2_15/BUF_2  ( .I(\SB1_2_18/buf_output[2] ), .Z(
        \SB2_2_15/i0_0 ) );
  NAND3_X1 \SB2_2_7/Component_Function_4/N4  ( .A1(\SB2_2_7/i1[9] ), .A2(
        \SB2_2_7/i1_5 ), .A3(\SB1_2_8/buf_output[4] ), .ZN(
        \SB2_2_7/Component_Function_4/NAND4_in[3] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_106  ( .I(\SB2_2_15/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[106] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_158  ( .I(\SB2_2_8/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[158] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_86  ( .I(\SB2_2_20/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[86] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_132  ( .I(\SB2_2_14/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[132] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_76  ( .I(\SB2_2_20/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[76] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_68  ( .I(\SB2_2_23/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[68] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_30  ( .I(\SB2_2_31/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[30] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_45  ( .I(\SB2_2_26/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[45] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_153  ( .I(\SB2_2_8/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[153] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_38  ( .I(\SB2_2_28/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[38] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_151  ( .I(\SB2_2_10/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[151] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_65  ( .I(\SB2_2_21/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[65] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_124  ( .I(\SB2_2_12/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[124] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_70  ( .I(\SB2_2_21/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[70] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_29  ( .I(\SB2_2_27/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[29] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_175  ( .I(\SB2_2_6/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[175] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_182  ( .I(\SB2_2_4/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[182] ) );
  BUF_X4 \SB1_3_0/BUF_5  ( .I(\MC_ARK_ARC_1_2/buf_output[191] ), .Z(
        \SB1_3_0/i0_3 ) );
  CLKBUF_X4 \SB1_3_3/BUF_2  ( .I(\MC_ARK_ARC_1_2/buf_output[170] ), .Z(
        \SB1_3_3/i0_0 ) );
  CLKBUF_X4 \SB1_3_30/BUF_2  ( .I(\MC_ARK_ARC_1_2/buf_output[8] ), .Z(
        \SB1_3_30/i0_0 ) );
  CLKBUF_X4 \SB2_3_18/BUF_0  ( .I(\SB1_3_23/buf_output[0] ), .Z(
        \SB2_3_18/i0[9] ) );
  CLKBUF_X4 \SB2_3_15/BUF_1  ( .I(\SB1_3_19/buf_output[1] ), .Z(
        \SB2_3_15/i0[6] ) );
  CLKBUF_X4 \SB2_3_29/BUF_0  ( .I(\SB1_3_2/buf_output[0] ), .Z(
        \SB2_3_29/i0[9] ) );
  CLKBUF_X4 \SB2_3_1/BUF_1  ( .I(\SB1_3_5/buf_output[1] ), .Z(\SB2_3_1/i0[6] )
         );
  CLKBUF_X4 \SB2_3_17/BUF_0  ( .I(\SB1_3_22/buf_output[0] ), .Z(
        \SB2_3_17/i0[9] ) );
  CLKBUF_X4 \SB2_3_2/BUF_0  ( .I(\SB1_3_7/buf_output[0] ), .Z(\SB2_3_2/i0[9] )
         );
  CLKBUF_X4 \SB2_3_20/BUF_1  ( .I(\SB1_3_24/buf_output[1] ), .Z(
        \SB2_3_20/i0[6] ) );
  CLKBUF_X4 \SB2_3_22/BUF_2  ( .I(\SB1_3_25/buf_output[2] ), .Z(
        \SB2_3_22/i0_0 ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_5  ( .I(\SB2_3_31/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[5] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_122  ( .I(\SB2_3_14/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[122] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_6  ( .I(\SB2_3_3/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[6] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_12  ( .I(\SB2_3_2/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[12] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_28  ( .I(\SB2_3_28/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[28] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_182  ( .I(\SB2_3_4/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[182] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_40  ( .I(\SB2_3_26/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[40] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_81  ( .I(\SB2_3_20/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[81] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_168  ( .I(\SB2_3_8/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[168] ) );
  CLKBUF_X4 \SB3_31/BUF_0  ( .I(\MC_ARK_ARC_1_3/buf_output[0] ), .Z(
        \SB3_31/i0[9] ) );
  BUF_X2 \SB1_0_7/BUF_0  ( .I(n317), .Z(\SB1_0_7/i0[9] ) );
  BUF_X2 \SB1_0_26/BUF_0  ( .I(n260), .Z(\SB1_0_26/i0[9] ) );
  BUF_X2 \SB1_0_4/BUF_0  ( .I(n326), .Z(\SB1_0_4/i0[9] ) );
  BUF_X2 \SB1_0_18/BUF_0  ( .I(n284), .Z(\SB1_0_18/i0[9] ) );
  BUF_X2 \SB1_0_19/BUF_0  ( .I(n281), .Z(\SB1_0_19/i0[9] ) );
  BUF_X2 \SB1_0_3/BUF_0  ( .I(n329), .Z(\SB1_0_3/i0[9] ) );
  BUF_X2 \SB1_0_31/BUF_0  ( .I(n245), .Z(\SB1_0_31/i0[9] ) );
  BUF_X4 \SB2_0_24/BUF_5  ( .I(\SB1_0_24/buf_output[5] ), .Z(\SB2_0_24/i0_3 )
         );
  BUF_X4 \SB2_0_17/BUF_5  ( .I(\SB1_0_17/buf_output[5] ), .Z(\SB2_0_17/i0_3 )
         );
  BUF_X4 \SB2_0_19/BUF_5  ( .I(\SB1_0_19/buf_output[5] ), .Z(\SB2_0_19/i0_3 )
         );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_157  ( .I(\SB2_0_9/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[157] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_76  ( .I(\SB2_0_20/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[76] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_49  ( .I(\SB2_0_27/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[49] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_96  ( .I(\SB2_0_20/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[96] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_180  ( .I(\SB2_0_6/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[180] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_73  ( .I(\SB2_0_23/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[73] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_69  ( .I(\SB2_0_22/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[69] ) );
  BUF_X4 \SB1_1_10/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[131] ), .Z(
        \SB1_1_10/i0_3 ) );
  BUF_X4 \SB1_1_7/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[148] ), .Z(
        \SB1_1_7/i0_4 ) );
  BUF_X4 \SB1_1_4/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[167] ), .Z(
        \SB1_1_4/i0_3 ) );
  BUF_X4 \SB1_1_23/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[53] ), .Z(
        \SB1_1_23/i0_3 ) );
  BUF_X4 \SB1_1_29/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[17] ), .Z(
        \SB1_1_29/i0_3 ) );
  BUF_X4 \SB1_1_6/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[155] ), .Z(
        \SB1_1_6/i0_3 ) );
  BUF_X4 \SB1_1_2/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[179] ), .Z(
        \SB1_1_2/i0_3 ) );
  BUF_X4 \SB1_1_11/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[125] ), .Z(
        \SB1_1_11/i0_3 ) );
  BUF_X4 \SB1_1_19/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[77] ), .Z(
        \SB1_1_19/i0_3 ) );
  BUF_X4 \SB1_1_27/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[29] ), .Z(
        \SB1_1_27/i0_3 ) );
  BUF_X4 \SB2_1_22/BUF_4  ( .I(\SB1_1_23/buf_output[4] ), .Z(\SB2_1_22/i0_4 )
         );
  BUF_X4 \SB2_1_10/BUF_5  ( .I(\SB1_1_10/buf_output[5] ), .Z(\SB2_1_10/i0_3 )
         );
  BUF_X4 \SB2_1_14/BUF_5  ( .I(\SB1_1_14/buf_output[5] ), .Z(\SB2_1_14/i0_3 )
         );
  BUF_X4 \SB2_1_17/BUF_5  ( .I(\SB1_1_17/buf_output[5] ), .Z(\SB2_1_17/i0_3 )
         );
  BUF_X4 \SB2_1_21/BUF_5  ( .I(\SB1_1_21/buf_output[5] ), .Z(\SB2_1_21/i0_3 )
         );
  BUF_X4 \SB2_1_16/BUF_5  ( .I(\SB1_1_16/buf_output[5] ), .Z(\SB2_1_16/i0_3 )
         );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_1  ( .I(\SB2_1_3/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[1] ) );
  BUF_X4 \SB1_2_24/BUF_3  ( .I(\MC_ARK_ARC_1_1/buf_output[45] ), .Z(
        \SB1_2_24/i0[10] ) );
  BUF_X4 \SB1_2_3/BUF_2  ( .I(\MC_ARK_ARC_1_1/buf_output[170] ), .Z(
        \SB1_2_3/i0_0 ) );
  BUF_X4 \SB1_2_1/BUF_5  ( .I(\MC_ARK_ARC_1_1/buf_output[185] ), .Z(
        \SB1_2_1/i0_3 ) );
  BUF_X4 \SB1_2_15/BUF_5  ( .I(\MC_ARK_ARC_1_1/buf_output[101] ), .Z(
        \SB1_2_15/i0_3 ) );
  BUF_X4 \SB1_2_7/BUF_5  ( .I(\MC_ARK_ARC_1_1/buf_output[149] ), .Z(
        \SB1_2_7/i0_3 ) );
  BUF_X4 \SB1_2_1/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[184] ), .Z(
        \SB1_2_1/i0_4 ) );
  BUF_X4 \SB1_2_13/BUF_5  ( .I(\MC_ARK_ARC_1_1/buf_output[113] ), .Z(
        \SB1_2_13/i0_3 ) );
  BUF_X4 \SB1_2_6/BUF_5  ( .I(\MC_ARK_ARC_1_1/buf_output[155] ), .Z(
        \SB1_2_6/i0_3 ) );
  BUF_X4 \SB1_2_17/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[88] ), .Z(
        \SB1_2_17/i0_4 ) );
  BUF_X4 \SB2_2_27/BUF_5  ( .I(\SB1_2_27/buf_output[5] ), .Z(\SB2_2_27/i0_3 )
         );
  BUF_X4 \SB2_2_21/BUF_5  ( .I(\SB1_2_21/buf_output[5] ), .Z(\SB2_2_21/i0_3 )
         );
  BUF_X4 \SB2_2_21/BUF_4  ( .I(\SB1_2_22/buf_output[4] ), .Z(\SB2_2_21/i0_4 )
         );
  BUF_X4 \SB2_2_13/BUF_5  ( .I(\SB1_2_13/buf_output[5] ), .Z(\SB2_2_13/i0_3 )
         );
  BUF_X4 \SB2_2_18/BUF_5  ( .I(\SB1_2_18/buf_output[5] ), .Z(\SB2_2_18/i0_3 )
         );
  BUF_X4 \SB2_2_5/BUF_5  ( .I(\SB1_2_5/buf_output[5] ), .Z(\SB2_2_5/i0_3 ) );
  BUF_X4 \SB2_2_14/BUF_5  ( .I(\SB1_2_14/buf_output[5] ), .Z(\SB2_2_14/i0_3 )
         );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_7  ( .I(\SB2_2_2/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[7] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_115  ( .I(\SB2_2_16/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[115] ) );
  BUF_X4 \SB1_3_26/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[34] ), .Z(
        \SB1_3_26/i0_4 ) );
  BUF_X4 \SB1_3_11/BUF_5  ( .I(\MC_ARK_ARC_1_2/buf_output[125] ), .Z(
        \SB1_3_11/i0_3 ) );
  BUF_X4 \SB1_3_7/BUF_5  ( .I(\MC_ARK_ARC_1_2/buf_output[149] ), .Z(
        \SB1_3_7/i0_3 ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_91  ( .I(\SB2_3_20/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[91] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_103  ( .I(\SB2_3_18/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[103] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_178  ( .I(\SB2_3_3/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[178] ) );
  INV_X1 \SB1_0_22/INV_3  ( .I(n359), .ZN(\SB1_0_22/i0[8] ) );
  NAND3_X1 \SB1_1_14/Component_Function_3/N2  ( .A1(\SB1_1_14/i0_0 ), .A2(
        \SB1_1_14/i0_3 ), .A3(\SB1_1_14/i0_4 ), .ZN(
        \SB1_1_14/Component_Function_3/NAND4_in[1] ) );
  BUF_X4 \SB1_0_5/BUF_5  ( .I(n431), .Z(\SB1_0_5/i0_3 ) );
  NAND3_X1 \SB2_1_23/Component_Function_1/N4  ( .A1(\SB2_1_23/i1_7 ), .A2(
        \SB2_1_23/i0[8] ), .A3(\SB2_1_23/i0_4 ), .ZN(
        \SB2_1_23/Component_Function_1/NAND4_in[3] ) );
  BUF_X4 \SB1_0_9/BUF_5  ( .I(n427), .Z(\SB1_0_9/i0_3 ) );
  NAND4_X2 \SB2_0_21/Component_Function_4/N5  ( .A1(
        \SB2_0_21/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_21/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_21/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_0_21/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_0_21/buf_output[4] ) );
  NAND4_X2 \SB1_2_18/Component_Function_4/N5  ( .A1(
        \SB1_2_18/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_18/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_18/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_18/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_2_18/buf_output[4] ) );
  BUF_X2 \SB1_0_22/BUF_3  ( .I(n359), .Z(\SB1_0_22/i0[10] ) );
  NAND3_X1 \SB1_0_20/Component_Function_5/N2  ( .A1(\SB1_0_20/i0_0 ), .A2(
        \SB1_0_20/i0[6] ), .A3(\SB1_0_20/i0[10] ), .ZN(
        \SB1_0_20/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 \SB1_0_1/Component_Function_4/N5  ( .A1(
        \SB1_0_1/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_1/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_1/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_1/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_0_1/buf_output[4] ) );
  INV_X1 \SB4_17/INV_0  ( .I(\SB3_22/buf_output[0] ), .ZN(\SB4_17/i3[0] ) );
  NAND3_X2 \SB1_3_8/Component_Function_2/N4  ( .A1(\SB1_3_8/i1_5 ), .A2(
        \SB1_3_8/i0_0 ), .A3(\SB1_3_8/i0_4 ), .ZN(
        \SB1_3_8/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_11/Component_Function_5/N2  ( .A1(\SB2_3_11/i0_0 ), .A2(
        \SB2_3_11/i0[6] ), .A3(\SB1_3_13/buf_output[3] ), .ZN(
        \SB2_3_11/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_11/Component_Function_4/N2  ( .A1(\SB2_3_11/i3[0] ), .A2(
        \SB2_3_11/i0_0 ), .A3(\SB2_3_11/i1_7 ), .ZN(
        \SB2_3_11/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_27/Component_Function_4/N4  ( .A1(\SB1_0_27/i1[9] ), .A2(
        \SB1_0_27/i1_5 ), .A3(\SB1_0_27/i0_4 ), .ZN(
        \SB1_0_27/Component_Function_4/NAND4_in[3] ) );
  BUF_X2 \SB1_0_30/BUF_3  ( .I(n343), .Z(\SB1_0_30/i0[10] ) );
  INV_X1 \SB1_0_30/INV_3  ( .I(n343), .ZN(\SB1_0_30/i0[8] ) );
  NAND4_X2 \SB1_1_15/Component_Function_4/N5  ( .A1(
        \SB1_1_15/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_15/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_15/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_15/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_1_15/buf_output[4] ) );
  NAND4_X2 \SB1_2_23/Component_Function_4/N5  ( .A1(
        \SB1_2_23/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_23/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_23/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_23/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_2_23/buf_output[4] ) );
  NAND3_X1 \SB4_7/Component_Function_0/N4  ( .A1(\SB4_7/i0[7] ), .A2(
        \SB4_7/i0_3 ), .A3(\SB4_7/i0_0 ), .ZN(
        \SB4_7/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB4_17/Component_Function_2/N3  ( .A1(\SB4_17/i0_3 ), .A2(n3661), 
        .A3(\SB4_17/i0[9] ), .ZN(\SB4_17/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB4_19/Component_Function_5/N3  ( .A1(\SB4_19/i1[9] ), .A2(
        \SB4_19/i0_4 ), .A3(\SB4_19/i0_3 ), .ZN(
        \SB4_19/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB4_28/Component_Function_5/N3  ( .A1(n5514), .A2(\SB4_28/i0_4 ), 
        .A3(\SB4_28/i0_3 ), .ZN(\SB4_28/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB4_27/Component_Function_5/N4  ( .A1(\SB4_27/i0[9] ), .A2(
        \SB4_27/i0[6] ), .A3(\SB4_27/i0_4 ), .ZN(
        \SB4_27/Component_Function_5/NAND4_in[3] ) );
  INV_X1 \SB4_23/INV_0  ( .I(\SB3_28/buf_output[0] ), .ZN(\SB4_23/i3[0] ) );
  NAND3_X1 \SB2_3_1/Component_Function_4/N2  ( .A1(\SB2_3_1/i3[0] ), .A2(
        \SB2_3_1/i0_0 ), .A3(\SB2_3_1/i1_7 ), .ZN(
        \SB2_3_1/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_0/Component_Function_5/N4  ( .A1(\SB1_3_0/i0[9] ), .A2(
        \SB1_3_0/i0[6] ), .A3(\SB1_3_0/i0_4 ), .ZN(
        \SB1_3_0/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_13/Component_Function_4/N3  ( .A1(\SB2_0_13/i0[9] ), .A2(
        \SB2_0_13/i0[10] ), .A3(\SB2_0_13/i0_3 ), .ZN(
        \SB2_0_13/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_10/Component_Function_4/N4  ( .A1(\SB2_0_10/i1[9] ), .A2(
        \SB2_0_10/i1_5 ), .A3(\SB2_0_10/i0_4 ), .ZN(
        \SB2_0_10/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_27/Component_Function_1/N4  ( .A1(\SB1_0_27/i1_7 ), .A2(
        \SB1_0_27/i0[8] ), .A3(\SB1_0_27/i0_4 ), .ZN(
        \SB1_0_27/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_26/Component_Function_5/N2  ( .A1(\SB1_0_26/i0_0 ), .A2(
        \SB1_0_26/i0[6] ), .A3(\SB1_0_26/i0[10] ), .ZN(
        \SB1_0_26/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_20/Component_Function_5/N4  ( .A1(\SB1_0_20/i0[9] ), .A2(
        n279), .A3(n364), .ZN(\SB1_0_20/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_9/Component_Function_5/N4  ( .A1(\SB1_0_9/i0[9] ), .A2(
        \SB1_0_9/i0[6] ), .A3(\SB1_0_9/i0_4 ), .ZN(
        \SB1_0_9/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_9/Component_Function_4/N4  ( .A1(\SB1_0_9/i1[9] ), .A2(
        \SB1_0_9/i1_5 ), .A3(\SB1_0_9/i0_4 ), .ZN(
        \SB1_0_9/Component_Function_4/NAND4_in[3] ) );
  NAND4_X2 \SB1_3_20/Component_Function_0/N5  ( .A1(
        \SB1_3_20/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_20/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_20/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_20/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_3_20/buf_output[0] ) );
  NAND4_X2 \SB1_2_27/Component_Function_0/N5  ( .A1(
        \SB1_2_27/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_27/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_27/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_27/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_2_27/buf_output[0] ) );
  NAND4_X2 \SB1_0_13/Component_Function_1/N5  ( .A1(
        \SB1_0_13/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_13/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_13/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_13/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_0_13/buf_output[1] ) );
  BUF_X4 \SB1_0_31/BUF_5  ( .I(n405), .Z(\SB1_0_31/i0_3 ) );
  BUF_X4 \SB1_2_0/BUF_2  ( .I(\MC_ARK_ARC_1_1/buf_output[188] ), .Z(
        \SB1_2_0/i0_0 ) );
  INV_X2 \SB1_0_0/INV_2  ( .I(n340), .ZN(\SB1_0_0/i1[9] ) );
  INV_X2 \SB1_2_21/INV_5  ( .I(n3681), .ZN(\SB1_2_21/i1_5 ) );
  NAND4_X2 \SB1_2_31/Component_Function_1/N5  ( .A1(
        \SB1_2_31/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_31/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_31/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_31/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_2_31/buf_output[1] ) );
  BUF_X4 \SB1_0_19/BUF_5  ( .I(n417), .Z(\SB1_0_19/i0_3 ) );
  INV_X2 \SB2_1_22/INV_5  ( .I(\SB1_1_22/buf_output[5] ), .ZN(\SB2_1_22/i1_5 )
         );
  INV_X2 \SB2_0_16/INV_5  ( .I(\RI3[0][95] ), .ZN(\SB2_0_16/i1_5 ) );
  NAND3_X2 \SB2_1_18/Component_Function_5/N3  ( .A1(\SB2_1_18/i1[9] ), .A2(
        \SB2_1_18/i0_4 ), .A3(\SB2_1_18/i0_3 ), .ZN(
        \SB2_1_18/Component_Function_5/NAND4_in[2] ) );
  INV_X2 \SB2_3_26/INV_5  ( .I(\RI3[3][35] ), .ZN(\SB2_3_26/i1_5 ) );
  INV_X2 \SB1_0_19/INV_2  ( .I(n283), .ZN(\SB1_0_19/i1[9] ) );
  INV_X2 \SB1_0_8/INV_2  ( .I(n316), .ZN(\SB1_0_8/i1[9] ) );
  INV_X2 \SB4_2/INV_3  ( .I(\SB3_4/buf_output[3] ), .ZN(\SB4_2/i0[8] ) );
  NAND4_X2 \SB1_2_18/Component_Function_1/N5  ( .A1(
        \SB1_2_18/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_18/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_18/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_18/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_2_18/buf_output[1] ) );
  BUF_X4 \SB1_0_0/BUF_5  ( .I(n436), .Z(\SB1_0_0/i0_3 ) );
  NAND4_X2 \SB1_3_3/Component_Function_4/N5  ( .A1(
        \SB1_3_3/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_3/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_3/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_3_3/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_3_3/buf_output[4] ) );
  NAND4_X2 \SB2_1_22/Component_Function_1/N5  ( .A1(
        \SB2_1_22/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_22/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_22/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_22/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_1_22/buf_output[1] ) );
  NAND4_X2 \SB1_2_28/Component_Function_0/N5  ( .A1(
        \SB1_2_28/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_28/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_28/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_28/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_2_28/buf_output[0] ) );
  NAND4_X2 \SB2_3_18/Component_Function_1/N5  ( .A1(
        \SB2_3_18/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_18/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_18/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_18/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_3_18/buf_output[1] ) );
  NAND4_X2 \SB1_3_25/Component_Function_0/N5  ( .A1(
        \SB1_3_25/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_25/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_25/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_25/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_3_25/buf_output[0] ) );
  INV_X2 \SB1_0_26/INV_2  ( .I(n262), .ZN(\SB1_0_26/i1[9] ) );
  NAND4_X2 \SB2_0_26/Component_Function_3/N5  ( .A1(
        \SB2_0_26/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_26/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_0_26/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_0_26/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_0_26/buf_output[3] ) );
  NAND3_X1 \SB1_0_26/Component_Function_2/N4  ( .A1(\SB1_0_26/i1_5 ), .A2(
        \SB1_0_26/i0_0 ), .A3(\SB1_0_26/i0_4 ), .ZN(
        \SB1_0_26/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_28/Component_Function_4/N4  ( .A1(\SB1_0_28/i1[9] ), .A2(
        \SB1_0_28/i1_5 ), .A3(\SB1_0_28/i0_4 ), .ZN(
        \SB1_0_28/Component_Function_4/NAND4_in[3] ) );
  INV_X1 \SB3_21/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[60] ), .ZN(
        \SB3_21/i3[0] ) );
  NAND3_X1 \SB1_3_9/Component_Function_4/N4  ( .A1(\SB1_3_9/i1[9] ), .A2(
        \SB1_3_9/i1_5 ), .A3(\SB1_3_9/i0_4 ), .ZN(
        \SB1_3_9/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB4_7/Component_Function_4/N3  ( .A1(\SB4_7/i0[9] ), .A2(
        \SB4_7/i0[10] ), .A3(\SB4_7/i0_3 ), .ZN(
        \SB4_7/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_13/Component_Function_5/N4  ( .A1(\SB2_3_13/i0[9] ), .A2(
        \SB2_3_13/i0[6] ), .A3(\SB1_3_14/buf_output[4] ), .ZN(
        \SB2_3_13/Component_Function_5/NAND4_in[3] ) );
  NAND4_X2 \SB2_1_16/Component_Function_4/N5  ( .A1(
        \SB2_1_16/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_16/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_16/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_1_16/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_1_16/buf_output[4] ) );
  NAND4_X2 \SB1_3_13/Component_Function_2/N5  ( .A1(
        \SB1_3_13/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_13/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_3_13/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_3_13/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB1_3_13/buf_output[2] ) );
  NAND4_X2 \SB1_3_8/Component_Function_2/N5  ( .A1(
        \SB1_3_8/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_8/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_3_8/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_3_8/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB1_3_8/buf_output[2] ) );
  NAND4_X2 \SB1_3_6/Component_Function_4/N5  ( .A1(
        \SB1_3_6/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_6/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_6/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_3_6/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_3_6/buf_output[4] ) );
  NAND4_X2 \SB1_3_22/Component_Function_0/N5  ( .A1(
        \SB1_3_22/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_22/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_22/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_22/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_3_22/buf_output[0] ) );
  NAND3_X2 \SB3_21/Component_Function_5/N2  ( .A1(\SB3_21/i0_0 ), .A2(
        \SB3_21/i0[6] ), .A3(\SB3_21/i0[10] ), .ZN(
        \SB3_21/Component_Function_5/NAND4_in[1] ) );
  INV_X2 \SB3_21/INV_5  ( .I(\RI1[4][65] ), .ZN(\SB3_21/i1_5 ) );
  NAND4_X2 \SB2_2_8/Component_Function_1/N5  ( .A1(
        \SB2_2_8/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_8/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_8/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_8/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_2_8/buf_output[1] ) );
  BUF_X4 \SB1_0_3/BUF_5  ( .I(n433), .Z(\SB1_0_3/i0_3 ) );
  INV_X2 \SB1_0_3/INV_2  ( .I(n331), .ZN(\SB1_0_3/i1[9] ) );
  NAND3_X2 \SB3_21/Component_Function_5/N4  ( .A1(\SB3_21/i0[9] ), .A2(
        \SB3_21/i0[6] ), .A3(\SB3_21/i0_4 ), .ZN(
        \SB3_21/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_19/Component_Function_4/N4  ( .A1(\SB1_0_19/i1[9] ), .A2(
        \SB1_0_19/i1_5 ), .A3(\SB1_0_19/i0_4 ), .ZN(
        \SB1_0_19/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_8/Component_Function_5/N2  ( .A1(\SB1_0_8/i0_0 ), .A2(
        \SB1_0_8/i0[6] ), .A3(\SB1_0_8/i0[10] ), .ZN(
        \SB1_0_8/Component_Function_5/NAND4_in[1] ) );
  INV_X1 \SB2_0_0/INV_0  ( .I(\SB1_0_5/buf_output[0] ), .ZN(\SB2_0_0/i3[0] )
         );
  BUF_X2 \SB2_0_5/BUF_1  ( .I(\SB1_0_9/buf_output[1] ), .Z(\SB2_0_5/i0[6] ) );
  NAND3_X1 \SB2_0_12/Component_Function_4/N4  ( .A1(\SB2_0_12/i1[9] ), .A2(
        \SB2_0_12/i1_5 ), .A3(\SB2_0_12/i0_4 ), .ZN(
        \SB2_0_12/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_25/Component_Function_5/N4  ( .A1(\SB2_0_25/i0[9] ), .A2(
        \RI3[0][37] ), .A3(\RI3[0][40] ), .ZN(
        \SB2_0_25/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_20/Component_Function_5/N3  ( .A1(\SB2_0_20/i1[9] ), .A2(
        \SB2_0_20/i0_4 ), .A3(\SB1_0_20/buf_output[5] ), .ZN(
        \SB2_0_20/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_26/Component_Function_5/N4  ( .A1(\SB2_0_26/i0[9] ), .A2(
        \SB2_0_26/i0[6] ), .A3(\RI3[0][34] ), .ZN(
        \SB2_0_26/Component_Function_5/NAND4_in[3] ) );
  BUF_X2 \SB1_1_12/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[115] ), .Z(
        \SB1_1_12/i0[6] ) );
  BUF_X2 \SB1_1_18/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[79] ), .Z(
        \SB1_1_18/i0[6] ) );
  NAND3_X1 \SB1_1_24/Component_Function_1/N3  ( .A1(\SB1_1_24/i1_5 ), .A2(
        \SB1_1_24/i0[6] ), .A3(\SB1_1_24/i0[9] ), .ZN(
        \SB1_1_24/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_10/Component_Function_2/N2  ( .A1(\SB1_1_10/i0_3 ), .A2(
        \SB1_1_10/i0[10] ), .A3(\SB1_1_10/i0[6] ), .ZN(
        \SB1_1_10/Component_Function_2/NAND4_in[1] ) );
  INV_X2 \SB2_1_0/INV_2  ( .I(\SB1_1_3/buf_output[2] ), .ZN(\SB2_1_0/i1[9] )
         );
  BUF_X4 \SB2_1_2/BUF_5  ( .I(\SB1_1_2/buf_output[5] ), .Z(\SB2_1_2/i0_3 ) );
  INV_X1 \SB2_1_30/INV_5  ( .I(\SB1_1_30/buf_output[5] ), .ZN(\SB2_1_30/i1_5 )
         );
  NAND3_X1 \SB2_1_0/Component_Function_4/N2  ( .A1(\SB2_1_0/i3[0] ), .A2(
        \SB2_1_0/i0_0 ), .A3(\SB2_1_0/i1_7 ), .ZN(
        \SB2_1_0/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_24/Component_Function_4/N4  ( .A1(\SB2_1_24/i1[9] ), .A2(
        \SB2_1_24/i1_5 ), .A3(\SB2_1_24/i0_4 ), .ZN(
        \SB2_1_24/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_25/Component_Function_5/N4  ( .A1(\SB2_1_25/i0[9] ), .A2(
        \SB1_1_29/buf_output[1] ), .A3(\SB1_1_26/buf_output[4] ), .ZN(
        \SB2_1_25/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_3/Component_Function_4/N3  ( .A1(\SB2_1_3/i0[9] ), .A2(
        \SB2_1_3/i0[10] ), .A3(\SB2_1_3/i0_3 ), .ZN(
        \SB2_1_3/Component_Function_4/NAND4_in[2] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_155  ( .I(\SB2_1_6/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[155] ) );
  NAND3_X1 \SB1_2_11/Component_Function_0/N3  ( .A1(\SB1_2_11/i0[10] ), .A2(
        \SB1_2_11/i0_4 ), .A3(\SB1_2_11/i0_3 ), .ZN(
        \SB1_2_11/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_28/Component_Function_4/N3  ( .A1(\SB1_2_28/i0[9] ), .A2(
        \SB1_2_28/i0[10] ), .A3(\SB1_2_28/i0_3 ), .ZN(
        \SB1_2_28/Component_Function_4/NAND4_in[2] ) );
  BUF_X2 \SB2_2_22/BUF_0  ( .I(\SB1_2_27/buf_output[0] ), .Z(\SB2_2_22/i0[9] )
         );
  NAND3_X1 \SB2_2_24/Component_Function_4/N4  ( .A1(\SB2_2_24/i1[9] ), .A2(
        \SB2_2_24/i1_5 ), .A3(\SB2_2_24/i0_4 ), .ZN(
        \SB2_2_24/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_7/Component_Function_2/N4  ( .A1(\SB2_2_7/i1_5 ), .A2(
        \SB2_2_7/i0_0 ), .A3(\SB1_2_8/buf_output[4] ), .ZN(
        \SB2_2_7/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_19/Component_Function_4/N2  ( .A1(\SB2_2_19/i3[0] ), .A2(
        \SB2_2_19/i0_0 ), .A3(\SB2_2_19/i1_7 ), .ZN(
        \SB2_2_19/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_6/Component_Function_5/N4  ( .A1(\SB2_2_6/i0[9] ), .A2(
        \SB1_2_10/buf_output[1] ), .A3(\SB1_2_7/buf_output[4] ), .ZN(
        \SB2_2_6/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_29/Component_Function_5/N3  ( .A1(\SB2_2_29/i1[9] ), .A2(
        \SB2_2_29/i0_4 ), .A3(\SB1_2_29/buf_output[5] ), .ZN(
        \SB2_2_29/Component_Function_5/NAND4_in[2] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_148  ( .I(\SB2_2_8/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[148] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_4  ( .I(\SB2_2_0/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[4] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_149  ( .I(\SB2_2_7/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[149] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_99  ( .I(\SB2_2_17/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[99] ) );
  INV_X1 \SB2_3_11/INV_1  ( .I(\SB1_3_15/buf_output[1] ), .ZN(\SB2_3_11/i1_7 )
         );
  NAND3_X1 \SB2_3_6/Component_Function_4/N4  ( .A1(\SB2_3_6/i1[9] ), .A2(
        \SB2_3_6/i1_5 ), .A3(\SB1_3_7/buf_output[4] ), .ZN(
        \SB2_3_6/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_17/Component_Function_4/N2  ( .A1(\SB2_3_17/i3[0] ), .A2(
        \SB2_3_17/i0_0 ), .A3(\SB2_3_17/i1_7 ), .ZN(
        \SB2_3_17/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_26/Component_Function_4/N4  ( .A1(\SB2_3_26/i1[9] ), .A2(
        \SB2_3_26/i1_5 ), .A3(\SB2_3_26/i0_4 ), .ZN(
        \SB2_3_26/Component_Function_4/NAND4_in[3] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_142  ( .I(\SB2_3_9/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[142] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_71  ( .I(\SB2_3_20/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[71] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_53  ( .I(\SB2_3_23/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[53] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_104  ( .I(\SB2_3_17/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[104] ) );
  BUF_X4 \SB3_4/BUF_5  ( .I(\MC_ARK_ARC_1_3/buf_output[167] ), .Z(\SB3_4/i0_3 ) );
  BUF_X2 \SB3_5/BUF_1  ( .I(\MC_ARK_ARC_1_3/buf_output[157] ), .Z(
        \SB3_5/i0[6] ) );
  BUF_X2 \SB3_15/BUF_1  ( .I(\MC_ARK_ARC_1_3/buf_output[97] ), .Z(
        \SB3_15/i0[6] ) );
  NAND3_X1 \SB3_29/Component_Function_2/N3  ( .A1(\SB3_29/i0_3 ), .A2(
        \SB3_29/i0[8] ), .A3(\SB3_29/i0[9] ), .ZN(
        \SB3_29/Component_Function_2/NAND4_in[2] ) );
  INV_X1 \SB4_1/INV_0  ( .I(\SB3_6/buf_output[0] ), .ZN(\SB4_1/i3[0] ) );
  INV_X1 \SB4_21/INV_1  ( .I(\SB3_25/buf_output[1] ), .ZN(\SB4_21/i1_7 ) );
  NAND3_X1 \SB4_26/Component_Function_0/N4  ( .A1(\SB4_26/i0[7] ), .A2(
        \SB4_26/i0_3 ), .A3(\SB4_26/i0_0 ), .ZN(
        \SB4_26/Component_Function_0/NAND4_in[3] ) );
  BUF_X2 U1 ( .I(Key[94]), .Z(n74) );
  BUF_X2 U13 ( .I(Key[100]), .Z(n189) );
  CLKBUF_X2 U14 ( .I(Key[67]), .Z(n211) );
  CLKBUF_X2 U15 ( .I(Key[66]), .Z(n224) );
  CLKBUF_X2 U16 ( .I(Key[126]), .Z(n222) );
  CLKBUF_X2 U19 ( .I(Key[6]), .Z(n57) );
  CLKBUF_X2 U21 ( .I(Key[37]), .Z(n40) );
  CLKBUF_X2 U22 ( .I(Key[144]), .Z(n72) );
  CLKBUF_X2 U23 ( .I(Key[55]), .Z(n101) );
  CLKBUF_X2 U24 ( .I(Key[34]), .Z(n185) );
  CLKBUF_X2 U27 ( .I(Key[158]), .Z(n10) );
  CLKBUF_X2 U28 ( .I(Key[13]), .Z(n50) );
  CLKBUF_X2 U32 ( .I(Key[27]), .Z(n25) );
  CLKBUF_X2 U35 ( .I(Key[48]), .Z(n98) );
  CLKBUF_X2 U38 ( .I(Key[151]), .Z(n93) );
  CLKBUF_X2 U40 ( .I(Key[41]), .Z(n107) );
  CLKBUF_X2 U44 ( .I(Key[159]), .Z(n215) );
  CLKBUF_X2 U45 ( .I(Key[79]), .Z(n89) );
  CLKBUF_X2 U48 ( .I(Key[145]), .Z(n20) );
  CLKBUF_X2 U50 ( .I(Key[131]), .Z(n94) );
  CLKBUF_X2 U52 ( .I(Key[138]), .Z(n21) );
  BUF_X2 U55 ( .I(Key[16]), .Z(n228) );
  CLKBUF_X2 U60 ( .I(Key[187]), .Z(n24) );
  CLKBUF_X2 U62 ( .I(Key[169]), .Z(n130) );
  CLKBUF_X2 U64 ( .I(Key[117]), .Z(n14) );
  CLKBUF_X2 U67 ( .I(Key[89]), .Z(n36) );
  CLKBUF_X2 U68 ( .I(Key[72]), .Z(n29) );
  CLKBUF_X2 U71 ( .I(Key[93]), .Z(n56) );
  CLKBUF_X2 U72 ( .I(Key[124]), .Z(n158) );
  BUF_X2 U73 ( .I(Key[22]), .Z(n230) );
  CLKBUF_X2 U75 ( .I(Key[103]), .Z(n209) );
  CLKBUF_X2 U79 ( .I(Key[20]), .Z(n136) );
  CLKBUF_X2 U80 ( .I(Key[15]), .Z(n208) );
  CLKBUF_X2 U82 ( .I(Key[118]), .Z(n64) );
  CLKBUF_X2 U83 ( .I(Key[54]), .Z(n113) );
  CLKBUF_X2 U85 ( .I(Key[104]), .Z(n192) );
  CLKBUF_X2 U87 ( .I(Key[83]), .Z(n92) );
  CLKBUF_X2 U89 ( .I(Key[81]), .Z(n180) );
  CLKBUF_X2 U91 ( .I(Key[60]), .Z(n53) );
  CLKBUF_X2 U93 ( .I(Key[153]), .Z(n33) );
  CLKBUF_X2 U97 ( .I(Key[125]), .Z(n59) );
  CLKBUF_X2 U98 ( .I(Key[53]), .Z(n176) );
  CLKBUF_X2 U99 ( .I(Key[33]), .Z(n194) );
  CLKBUF_X2 U100 ( .I(Key[160]), .Z(n61) );
  CLKBUF_X2 U101 ( .I(Key[139]), .Z(n26) );
  CLKBUF_X2 U104 ( .I(Key[171]), .Z(n128) );
  CLKBUF_X2 U108 ( .I(Key[157]), .Z(n121) );
  CLKBUF_X2 U109 ( .I(Key[64]), .Z(n97) );
  CLKBUF_X2 U110 ( .I(Key[161]), .Z(n118) );
  CLKBUF_X2 U111 ( .I(Key[36]), .Z(n3) );
  CLKBUF_X2 U114 ( .I(Key[129]), .Z(n76) );
  CLKBUF_X2 U116 ( .I(Key[150]), .Z(n131) );
  CLKBUF_X2 U119 ( .I(Key[77]), .Z(n109) );
  CLKBUF_X2 U120 ( .I(Key[92]), .Z(n63) );
  CLKBUF_X2 U121 ( .I(Key[115]), .Z(n81) );
  CLKBUF_X2 U122 ( .I(Key[21]), .Z(n86) );
  CLKBUF_X2 U123 ( .I(Key[0]), .Z(n55) );
  CLKBUF_X2 U124 ( .I(Key[127]), .Z(n27) );
  CLKBUF_X2 U125 ( .I(Key[185]), .Z(n191) );
  CLKBUF_X2 U126 ( .I(Key[108]), .Z(n6) );
  CLKBUF_X2 U127 ( .I(Key[42]), .Z(n13) );
  CLKBUF_X2 U128 ( .I(Key[4]), .Z(n65) );
  CLKBUF_X2 U129 ( .I(Key[148]), .Z(n135) );
  CLKBUF_X2 U131 ( .I(Key[19]), .Z(n84) );
  CLKBUF_X2 U132 ( .I(Key[175]), .Z(n9) );
  CLKBUF_X2 U138 ( .I(Key[182]), .Z(n46) );
  CLKBUF_X2 U139 ( .I(Key[122]), .Z(n106) );
  CLKBUF_X2 U142 ( .I(Key[73]), .Z(n48) );
  CLKBUF_X2 U143 ( .I(Key[35]), .Z(n243) );
  BUF_X2 U144 ( .I(Key[70]), .Z(n210) );
  CLKBUF_X2 U145 ( .I(Key[49]), .Z(n70) );
  CLKBUF_X2 U146 ( .I(Key[78]), .Z(n83) );
  CLKBUF_X2 U149 ( .I(Key[101]), .Z(n190) );
  CLKBUF_X2 U150 ( .I(Key[50]), .Z(n68) );
  CLKBUF_X2 U151 ( .I(Key[63]), .Z(n212) );
  CLKBUF_X2 U152 ( .I(Key[176]), .Z(n52) );
  CLKBUF_X2 U154 ( .I(Key[31]), .Z(n17) );
  CLKBUF_X2 U156 ( .I(Key[141]), .Z(n226) );
  CLKBUF_X2 U158 ( .I(Key[52]), .Z(n218) );
  CLKBUF_X2 U159 ( .I(Key[190]), .Z(n80) );
  CLKBUF_X2 U160 ( .I(Key[121]), .Z(n34) );
  CLKBUF_X2 U161 ( .I(Key[17]), .Z(n232) );
  BUF_X2 U162 ( .I(Key[142]), .Z(n233) );
  CLKBUF_X2 U163 ( .I(Key[154]), .Z(n236) );
  CLKBUF_X2 U165 ( .I(Key[128]), .Z(n95) );
  CLKBUF_X2 U166 ( .I(Key[114]), .Z(n45) );
  CLKBUF_X2 U167 ( .I(Key[24]), .Z(n173) );
  CLKBUF_X2 U168 ( .I(Key[107]), .Z(n58) );
  CLKBUF_X2 U169 ( .I(Key[95]), .Z(n178) );
  CLKBUF_X2 U170 ( .I(Key[133]), .Z(n2) );
  CLKBUF_X2 U171 ( .I(Key[116]), .Z(n144) );
  CLKBUF_X2 U172 ( .I(Key[29]), .Z(n184) );
  CLKBUF_X2 U174 ( .I(Key[109]), .Z(n5) );
  CLKBUF_X2 U175 ( .I(Key[140]), .Z(n127) );
  CLKBUF_X2 U176 ( .I(Key[38]), .Z(n166) );
  CLKBUF_X2 U177 ( .I(Key[177]), .Z(n108) );
  BUF_X2 U178 ( .I(Key[130]), .Z(n202) );
  CLKBUF_X2 U185 ( .I(Key[87]), .Z(n186) );
  CLKBUF_X2 U186 ( .I(Key[84]), .Z(n31) );
  CLKBUF_X2 U187 ( .I(Key[99]), .Z(n42) );
  CLKBUF_X2 U189 ( .I(Key[188]), .Z(n223) );
  CLKBUF_X2 U191 ( .I(Key[163]), .Z(n141) );
  CLKBUF_X2 U192 ( .I(Key[174]), .Z(n47) );
  CLKBUF_X2 U193 ( .I(Key[85]), .Z(n134) );
  CLKBUF_X2 U195 ( .I(Key[167]), .Z(n231) );
  CLKBUF_X2 U196 ( .I(Key[149]), .Z(n75) );
  CLKBUF_X2 U197 ( .I(Key[189]), .Z(n51) );
  BUF_X2 U198 ( .I(Key[5]), .Z(n221) );
  BUF_X2 U199 ( .I(Key[2]), .Z(n7) );
  XOR2_X1 U200 ( .A1(Plaintext[180]), .A2(Key[180]), .Z(n335) );
  XOR2_X1 U204 ( .A1(Plaintext[75]), .A2(Key[75]), .Z(n365) );
  XOR2_X1 U205 ( .A1(Plaintext[40]), .A2(Key[40]), .Z(n354) );
  XOR2_X1 U206 ( .A1(Plaintext[76]), .A2(Key[76]), .Z(n366) );
  INV_X1 U207 ( .I(n235), .ZN(n155) );
  INV_X1 U208 ( .I(n225), .ZN(n8) );
  INV_X1 U209 ( .I(n206), .ZN(n145) );
  INV_X1 U210 ( .I(n197), .ZN(n54) );
  INV_X1 U211 ( .I(n212), .ZN(n123) );
  INV_X1 U212 ( .I(n223), .ZN(n4) );
  INV_X1 U213 ( .I(n67), .ZN(n11) );
  INV_X1 U214 ( .I(n133), .ZN(n35) );
  INV_X1 U215 ( .I(n172), .ZN(n110) );
  INV_X1 U216 ( .I(n190), .ZN(n87) );
  INV_X1 U217 ( .I(n214), .ZN(n175) );
  INV_X1 U218 ( .I(n227), .ZN(n151) );
  INV_X1 U219 ( .I(n205), .ZN(n78) );
  INV_X1 U220 ( .I(\MC_ARK_ARC_1_1/buf_keyinput[51] ), .ZN(n142) );
  INV_X1 U221 ( .I(n209), .ZN(n85) );
  INV_X1 U222 ( .I(n165), .ZN(n19) );
  INV_X1 U223 ( .I(n196), .ZN(n174) );
  INV_X1 U224 ( .I(n84), .ZN(n164) );
  INV_X1 U225 ( .I(n211), .ZN(n119) );
  INV_X1 U226 ( .I(n237), .ZN(n69) );
  INV_X1 U227 ( .I(n135), .ZN(n43) );
  INV_X1 U228 ( .I(n185), .ZN(n149) );
  INV_X1 U229 ( .I(n236), .ZN(n37) );
  INV_X1 U230 ( .I(n203), .ZN(n453) );
  INV_X1 U231 ( .I(n115), .ZN(n550) );
  INV_X1 U232 ( .I(n177), .ZN(n111) );
  INV_X1 U233 ( .I(n131), .ZN(n41) );
  INV_X1 U234 ( .I(n180), .ZN(n513) );
  INV_X1 U235 ( .I(n108), .ZN(n445) );
  INV_X1 U236 ( .I(n222), .ZN(n62) );
  INV_X1 U237 ( .I(n186), .ZN(n508) );
  INV_X1 U238 ( .I(n122), .ZN(n527) );
  INV_X1 U239 ( .I(n241), .ZN(n1) );
  INV_X1 U240 ( .I(n65), .ZN(n563) );
  INV_X1 U241 ( .I(n39), .ZN(n565) );
  INV_X1 U242 ( .I(n130), .ZN(n22) );
  INV_X1 U243 ( .I(n55), .ZN(n566) );
  INV_X1 U244 ( .I(n57), .ZN(n561) );
  INV_X1 U245 ( .I(n83), .ZN(n515) );
  INV_X1 U246 ( .I(n181), .ZN(n96) );
  INV_X1 U247 ( .I(n103), .ZN(n463) );
  INV_X1 U248 ( .I(n239), .ZN(n552) );
  INV_X1 U249 ( .I(n162), .ZN(n549) );
  INV_X1 U250 ( .I(n184), .ZN(n547) );
  INV_X1 U251 ( .I(n200), .ZN(n526) );
  INV_X1 U252 ( .I(n146), .ZN(n112) );
  INV_X1 U253 ( .I(n160), .ZN(n469) );
  INV_X1 U254 ( .I(n166), .ZN(n542) );
  INV_X1 U255 ( .I(n114), .ZN(n474) );
  INV_X1 U256 ( .I(n233), .ZN(n49) );
  INV_X1 U257 ( .I(n189), .ZN(n88) );
  INV_X1 U258 ( .I(n210), .ZN(n116) );
  INV_X1 U259 ( .I(n148), .ZN(n493) );
  INV_X1 U260 ( .I(n100), .ZN(n466) );
  INV_X1 U261 ( .I(n117), .ZN(n512) );
  INV_X1 U262 ( .I(n126), .ZN(n509) );
  INV_X1 U263 ( .I(n221), .ZN(n562) );
  INV_X1 U264 ( .I(n74), .ZN(n503) );
  INV_X1 U265 ( .I(n89), .ZN(n514) );
  INV_X1 U266 ( .I(n234), .ZN(n139) );
  INV_X1 U267 ( .I(n27), .ZN(n480) );
  INV_X1 U268 ( .I(n156), .ZN(n522) );
  INV_X1 U270 ( .I(n191), .ZN(n441) );
  INV_X1 U271 ( .I(n170), .ZN(n560) );
  INV_X1 U272 ( .I(n238), .ZN(n12) );
  INV_X1 U273 ( .I(n107), .ZN(n541) );
  INV_X1 U274 ( .I(n64), .ZN(n487) );
  INV_X1 U275 ( .I(n178), .ZN(n502) );
  INV_X1 U276 ( .I(n50), .ZN(n558) );
  INV_X1 U277 ( .I(n80), .ZN(n437) );
  INV_X1 U278 ( .I(n58), .ZN(n496) );
  INV_X1 U279 ( .I(n48), .ZN(n517) );
  INV_X1 U280 ( .I(n182), .ZN(n559) );
  INV_X1 U281 ( .I(n141), .ZN(n455) );
  INV_X1 U282 ( .I(n144), .ZN(n489) );
  INV_X1 U284 ( .I(n40), .ZN(n543) );
  INV_X1 U285 ( .I(n125), .ZN(n521) );
  INV_X1 U286 ( .I(n192), .ZN(n498) );
  INV_X1 U287 ( .I(n60), .ZN(n443) );
  INV_X1 U288 ( .I(n26), .ZN(n471) );
  INV_X1 U290 ( .I(n198), .ZN(n528) );
  INV_X1 U291 ( .I(n136), .ZN(n554) );
  INV_X1 U292 ( .I(n101), .ZN(n529) );
  INV_X1 U293 ( .I(n132), .ZN(n171) );
  INV_X1 U294 ( .I(n152), .ZN(n546) );
  INV_X1 U296 ( .I(n219), .ZN(n179) );
  INV_X1 U297 ( .I(n154), .ZN(n501) );
  INV_X1 U298 ( .I(n121), .ZN(n460) );
  INV_X1 U299 ( .I(n224), .ZN(n120) );
  INV_X1 U300 ( .I(n47), .ZN(n448) );
  INV_X1 U301 ( .I(n93), .ZN(n464) );
  INV_X1 U302 ( .I(n216), .ZN(n44) );
  INV_X1 U303 ( .I(n76), .ZN(n478) );
  INV_X1 U304 ( .I(n183), .ZN(n520) );
  INV_X1 U305 ( .I(n56), .ZN(n504) );
  INV_X1 U306 ( .I(n208), .ZN(n168) );
  INV_X1 U307 ( .I(n72), .ZN(n468) );
  INV_X1 U308 ( .I(n159), .ZN(n23) );
  INV_X1 U309 ( .I(n51), .ZN(n438) );
  INV_X1 U310 ( .I(n128), .ZN(n449) );
  INV_X1 U311 ( .I(n199), .ZN(n533) );
  INV_X1 U312 ( .I(n220), .ZN(n18) );
  INV_X1 U313 ( .I(n204), .ZN(n77) );
  INV_X1 U315 ( .I(n244), .ZN(n537) );
  INV_X1 U316 ( .I(n79), .ZN(n91) );
  INV_X1 U317 ( .I(n31), .ZN(n510) );
  INV_X1 U318 ( .I(n153), .ZN(n538) );
  INV_X1 U319 ( .I(n94), .ZN(n477) );
  INV_X1 U320 ( .I(n42), .ZN(n500) );
  INV_X1 U321 ( .I(n194), .ZN(n150) );
  INV_X1 U322 ( .I(n15), .ZN(n440) );
  INV_X1 U324 ( .I(n134), .ZN(n102) );
  INV_X1 U325 ( .I(n36), .ZN(n507) );
  INV_X1 U326 ( .I(n240), .ZN(n519) );
  INV_X1 U327 ( .I(n232), .ZN(n556) );
  INV_X1 U328 ( .I(n29), .ZN(n518) );
  INV_X1 U329 ( .I(n113), .ZN(n530) );
  INV_X1 U330 ( .I(n109), .ZN(n516) );
  INV_X1 U331 ( .I(n231), .ZN(n451) );
  INV_X1 U332 ( .I(n70), .ZN(n535) );
  INV_X1 U334 ( .I(n59), .ZN(n481) );
  INV_X1 U336 ( .I(n105), .ZN(n476) );
  INV_X1 U337 ( .I(n129), .ZN(n450) );
  INV_X1 U338 ( .I(n46), .ZN(n442) );
  INV_X1 U339 ( .I(n98), .ZN(n536) );
  INV_X1 U340 ( .I(n53), .ZN(n525) );
  INV_X1 U341 ( .I(n86), .ZN(n553) );
  INV_X1 U342 ( .I(n147), .ZN(n557) );
  INV_X1 U343 ( .I(n16), .ZN(n555) );
  INV_X1 U345 ( .I(n229), .ZN(n492) );
  INV_X1 U347 ( .I(n45), .ZN(n491) );
  INV_X1 U348 ( .I(n28), .ZN(n499) );
  INV_X1 U349 ( .I(n228), .ZN(n167) );
  INV_X1 U350 ( .I(n173), .ZN(n551) );
  INV_X1 U351 ( .I(n127), .ZN(n470) );
  INV_X1 U353 ( .I(n90), .ZN(n524) );
  INV_X1 U354 ( .I(n207), .ZN(n124) );
  INV_X1 U355 ( .I(n213), .ZN(n483) );
  INV_X1 U356 ( .I(n138), .ZN(n497) );
  INV_X1 U357 ( .I(n38), .ZN(n486) );
  INV_X1 U358 ( .I(n71), .ZN(n539) );
  INV_X1 U360 ( .I(n230), .ZN(n161) );
  INV_X1 U361 ( .I(n2), .ZN(n475) );
  INV_X1 U362 ( .I(n63), .ZN(n505) );
  INV_X1 U363 ( .I(n81), .ZN(n490) );
  INV_X1 U364 ( .I(n106), .ZN(n484) );
  INV_X1 U365 ( .I(n97), .ZN(n523) );
  INV_X1 U366 ( .I(n66), .ZN(n473) );
  INV_X1 U367 ( .I(n195), .ZN(n454) );
  INV_X1 U368 ( .I(n95), .ZN(n479) );
  INV_X1 U369 ( .I(n188), .ZN(n82) );
  INV_X1 U370 ( .I(n52), .ZN(n446) );
  INV_X1 U372 ( .I(n163), .ZN(n99) );
  INV_X1 U373 ( .I(n140), .ZN(n452) );
  INV_X1 U374 ( .I(n218), .ZN(n532) );
  INV_X1 U375 ( .I(n158), .ZN(n482) );
  INV_X1 U376 ( .I(n73), .ZN(n444) );
  INV_X1 U377 ( .I(n9), .ZN(n447) );
  INV_X1 U378 ( .I(n61), .ZN(n458) );
  XOR2_X1 U379 ( .A1(Key[0]), .A2(Plaintext[0]), .Z(n245) );
  XOR2_X1 U380 ( .A1(Key[1]), .A2(Plaintext[1]), .Z(n246) );
  XOR2_X1 U381 ( .A1(Key[2]), .A2(Plaintext[2]), .Z(n247) );
  XOR2_X1 U382 ( .A1(Key[3]), .A2(Plaintext[3]), .Z(n341) );
  XOR2_X1 U383 ( .A1(Key[4]), .A2(Plaintext[4]), .Z(n342) );
  XOR2_X1 U384 ( .A1(Key[5]), .A2(Plaintext[5]), .Z(n405) );
  XOR2_X1 U385 ( .A1(Key[6]), .A2(Plaintext[6]), .Z(n248) );
  XOR2_X1 U386 ( .A1(Key[7]), .A2(Plaintext[7]), .Z(n249) );
  XOR2_X1 U387 ( .A1(Key[8]), .A2(Plaintext[8]), .Z(n250) );
  XOR2_X1 U388 ( .A1(Key[9]), .A2(Plaintext[9]), .Z(n343) );
  XOR2_X1 U389 ( .A1(Key[10]), .A2(Plaintext[10]), .Z(n344) );
  XOR2_X1 U390 ( .A1(Key[11]), .A2(Plaintext[11]), .Z(n406) );
  XOR2_X1 U391 ( .A1(Key[12]), .A2(Plaintext[12]), .Z(n251) );
  XOR2_X1 U392 ( .A1(Key[13]), .A2(Plaintext[13]), .Z(n252) );
  XOR2_X1 U393 ( .A1(Key[14]), .A2(Plaintext[14]), .Z(n253) );
  XOR2_X1 U394 ( .A1(Key[15]), .A2(Plaintext[15]), .Z(n345) );
  XOR2_X1 U395 ( .A1(Key[16]), .A2(Plaintext[16]), .Z(n346) );
  XOR2_X1 U396 ( .A1(Key[17]), .A2(Plaintext[17]), .Z(n407) );
  XOR2_X1 U397 ( .A1(Key[18]), .A2(Plaintext[18]), .Z(n254) );
  XOR2_X1 U398 ( .A1(Key[19]), .A2(Plaintext[19]), .Z(n255) );
  XOR2_X1 U399 ( .A1(Key[20]), .A2(Plaintext[20]), .Z(n256) );
  XOR2_X1 U400 ( .A1(Key[21]), .A2(Plaintext[21]), .Z(n347) );
  XOR2_X1 U401 ( .A1(Key[22]), .A2(Plaintext[22]), .Z(n348) );
  XOR2_X1 U402 ( .A1(Key[23]), .A2(Plaintext[23]), .Z(n408) );
  XOR2_X1 U403 ( .A1(Key[24]), .A2(Plaintext[24]), .Z(n257) );
  XOR2_X1 U404 ( .A1(Key[25]), .A2(Plaintext[25]), .Z(n258) );
  XOR2_X1 U405 ( .A1(Key[26]), .A2(Plaintext[26]), .Z(n259) );
  XOR2_X1 U406 ( .A1(Key[27]), .A2(Plaintext[27]), .Z(n349) );
  XOR2_X1 U407 ( .A1(Key[28]), .A2(Plaintext[28]), .Z(n350) );
  XOR2_X1 U408 ( .A1(Key[29]), .A2(Plaintext[29]), .Z(n409) );
  XOR2_X1 U409 ( .A1(Key[30]), .A2(Plaintext[30]), .Z(n260) );
  XOR2_X1 U410 ( .A1(Key[31]), .A2(Plaintext[31]), .Z(n261) );
  XOR2_X1 U411 ( .A1(Key[32]), .A2(Plaintext[32]), .Z(n262) );
  XOR2_X1 U412 ( .A1(Key[33]), .A2(Plaintext[33]), .Z(n351) );
  XOR2_X1 U413 ( .A1(Key[34]), .A2(Plaintext[34]), .Z(n352) );
  XOR2_X1 U414 ( .A1(Key[35]), .A2(Plaintext[35]), .Z(n410) );
  XOR2_X1 U415 ( .A1(Key[36]), .A2(Plaintext[36]), .Z(n263) );
  XOR2_X1 U416 ( .A1(Key[37]), .A2(Plaintext[37]), .Z(n264) );
  XOR2_X1 U417 ( .A1(Key[38]), .A2(Plaintext[38]), .Z(n265) );
  XOR2_X1 U418 ( .A1(Key[39]), .A2(Plaintext[39]), .Z(n353) );
  XOR2_X1 U419 ( .A1(Key[41]), .A2(Plaintext[41]), .Z(n411) );
  XOR2_X1 U420 ( .A1(Key[42]), .A2(Plaintext[42]), .Z(n266) );
  XOR2_X1 U421 ( .A1(Key[43]), .A2(Plaintext[43]), .Z(n267) );
  XOR2_X1 U422 ( .A1(Key[44]), .A2(Plaintext[44]), .Z(n268) );
  XOR2_X1 U423 ( .A1(Key[45]), .A2(Plaintext[45]), .Z(n355) );
  XOR2_X1 U424 ( .A1(Key[46]), .A2(Plaintext[46]), .Z(n356) );
  XOR2_X1 U425 ( .A1(Key[47]), .A2(Plaintext[47]), .Z(n412) );
  XOR2_X1 U426 ( .A1(Key[48]), .A2(Plaintext[48]), .Z(n269) );
  XOR2_X1 U427 ( .A1(Key[49]), .A2(Plaintext[49]), .Z(n270) );
  XOR2_X1 U428 ( .A1(Key[50]), .A2(Plaintext[50]), .Z(n271) );
  XOR2_X1 U429 ( .A1(Key[51]), .A2(Plaintext[51]), .Z(n357) );
  XOR2_X1 U430 ( .A1(Key[52]), .A2(Plaintext[52]), .Z(n358) );
  XOR2_X1 U431 ( .A1(Key[53]), .A2(Plaintext[53]), .Z(n413) );
  XOR2_X1 U432 ( .A1(Key[54]), .A2(Plaintext[54]), .Z(n272) );
  XOR2_X1 U433 ( .A1(Key[55]), .A2(Plaintext[55]), .Z(n273) );
  XOR2_X1 U434 ( .A1(Key[56]), .A2(Plaintext[56]), .Z(n274) );
  XOR2_X1 U435 ( .A1(Key[57]), .A2(Plaintext[57]), .Z(n359) );
  XOR2_X1 U436 ( .A1(Key[58]), .A2(Plaintext[58]), .Z(n360) );
  XOR2_X1 U437 ( .A1(Key[59]), .A2(Plaintext[59]), .Z(n414) );
  XOR2_X1 U438 ( .A1(Key[60]), .A2(Plaintext[60]), .Z(n275) );
  XOR2_X1 U439 ( .A1(Key[61]), .A2(Plaintext[61]), .Z(n276) );
  XOR2_X1 U440 ( .A1(Key[62]), .A2(Plaintext[62]), .Z(n277) );
  XOR2_X1 U441 ( .A1(Key[63]), .A2(Plaintext[63]), .Z(n361) );
  XOR2_X1 U442 ( .A1(Key[64]), .A2(Plaintext[64]), .Z(n362) );
  XOR2_X1 U443 ( .A1(Key[65]), .A2(Plaintext[65]), .Z(n415) );
  XOR2_X1 U444 ( .A1(Key[66]), .A2(Plaintext[66]), .Z(n278) );
  XOR2_X1 U445 ( .A1(Key[67]), .A2(Plaintext[67]), .Z(n279) );
  XOR2_X1 U446 ( .A1(Key[68]), .A2(Plaintext[68]), .Z(n280) );
  XOR2_X1 U447 ( .A1(Key[69]), .A2(Plaintext[69]), .Z(n363) );
  XOR2_X1 U448 ( .A1(Key[70]), .A2(Plaintext[70]), .Z(n364) );
  XOR2_X1 U449 ( .A1(Key[71]), .A2(Plaintext[71]), .Z(n416) );
  XOR2_X1 U450 ( .A1(Key[72]), .A2(Plaintext[72]), .Z(n281) );
  XOR2_X1 U451 ( .A1(Key[73]), .A2(Plaintext[73]), .Z(n282) );
  XOR2_X1 U452 ( .A1(Key[74]), .A2(Plaintext[74]), .Z(n283) );
  XOR2_X1 U453 ( .A1(Key[77]), .A2(Plaintext[77]), .Z(n417) );
  XOR2_X1 U454 ( .A1(Key[78]), .A2(Plaintext[78]), .Z(n284) );
  XOR2_X1 U455 ( .A1(Key[79]), .A2(Plaintext[79]), .Z(n285) );
  XOR2_X1 U456 ( .A1(Key[80]), .A2(Plaintext[80]), .Z(n286) );
  XOR2_X1 U457 ( .A1(Key[81]), .A2(Plaintext[81]), .Z(n367) );
  XOR2_X1 U458 ( .A1(Key[82]), .A2(Plaintext[82]), .Z(n368) );
  XOR2_X1 U459 ( .A1(Key[83]), .A2(Plaintext[83]), .Z(n418) );
  XOR2_X1 U460 ( .A1(Key[84]), .A2(Plaintext[84]), .Z(n287) );
  XOR2_X1 U461 ( .A1(Key[85]), .A2(Plaintext[85]), .Z(n288) );
  XOR2_X1 U462 ( .A1(Key[86]), .A2(Plaintext[86]), .Z(n289) );
  XOR2_X1 U463 ( .A1(Key[87]), .A2(Plaintext[87]), .Z(n369) );
  XOR2_X1 U464 ( .A1(Key[88]), .A2(Plaintext[88]), .Z(n370) );
  XOR2_X1 U465 ( .A1(Key[89]), .A2(Plaintext[89]), .Z(n419) );
  XOR2_X1 U466 ( .A1(Key[90]), .A2(Plaintext[90]), .Z(n290) );
  XOR2_X1 U467 ( .A1(Key[91]), .A2(Plaintext[91]), .Z(n291) );
  XOR2_X1 U468 ( .A1(Key[92]), .A2(Plaintext[92]), .Z(n292) );
  XOR2_X1 U469 ( .A1(Key[93]), .A2(Plaintext[93]), .Z(n371) );
  XOR2_X1 U470 ( .A1(Key[94]), .A2(Plaintext[94]), .Z(n372) );
  XOR2_X1 U471 ( .A1(Key[95]), .A2(Plaintext[95]), .Z(n420) );
  XOR2_X1 U472 ( .A1(Key[96]), .A2(Plaintext[96]), .Z(n293) );
  XOR2_X1 U473 ( .A1(Key[97]), .A2(Plaintext[97]), .Z(n294) );
  XOR2_X1 U474 ( .A1(Key[98]), .A2(Plaintext[98]), .Z(n295) );
  XOR2_X1 U475 ( .A1(Key[99]), .A2(Plaintext[99]), .Z(n373) );
  XOR2_X1 U476 ( .A1(Key[100]), .A2(Plaintext[100]), .Z(n374) );
  XOR2_X1 U477 ( .A1(Key[101]), .A2(Plaintext[101]), .Z(n421) );
  XOR2_X1 U478 ( .A1(Key[102]), .A2(Plaintext[102]), .Z(n296) );
  XOR2_X1 U479 ( .A1(Key[103]), .A2(Plaintext[103]), .Z(n297) );
  XOR2_X1 U480 ( .A1(Key[104]), .A2(Plaintext[104]), .Z(n298) );
  XOR2_X1 U481 ( .A1(Key[105]), .A2(Plaintext[105]), .Z(n375) );
  XOR2_X1 U482 ( .A1(Key[106]), .A2(Plaintext[106]), .Z(n376) );
  XOR2_X1 U483 ( .A1(Key[107]), .A2(Plaintext[107]), .Z(n422) );
  XOR2_X1 U484 ( .A1(Key[108]), .A2(Plaintext[108]), .Z(n299) );
  XOR2_X1 U485 ( .A1(Key[109]), .A2(Plaintext[109]), .Z(n300) );
  XOR2_X1 U486 ( .A1(Key[110]), .A2(Plaintext[110]), .Z(n301) );
  XOR2_X1 U487 ( .A1(Key[111]), .A2(Plaintext[111]), .Z(n377) );
  XOR2_X1 U488 ( .A1(Key[112]), .A2(Plaintext[112]), .Z(n378) );
  XOR2_X1 U489 ( .A1(Key[113]), .A2(Plaintext[113]), .Z(n423) );
  XOR2_X1 U490 ( .A1(Key[114]), .A2(Plaintext[114]), .Z(n302) );
  XOR2_X1 U491 ( .A1(Key[115]), .A2(Plaintext[115]), .Z(n303) );
  XOR2_X1 U492 ( .A1(Key[116]), .A2(Plaintext[116]), .Z(n304) );
  XOR2_X1 U493 ( .A1(Key[117]), .A2(Plaintext[117]), .Z(n379) );
  XOR2_X1 U494 ( .A1(Key[118]), .A2(Plaintext[118]), .Z(n380) );
  XOR2_X1 U495 ( .A1(Key[119]), .A2(Plaintext[119]), .Z(n424) );
  XOR2_X1 U496 ( .A1(Key[120]), .A2(Plaintext[120]), .Z(n305) );
  XOR2_X1 U497 ( .A1(Key[121]), .A2(Plaintext[121]), .Z(n306) );
  XOR2_X1 U498 ( .A1(Key[122]), .A2(Plaintext[122]), .Z(n307) );
  XOR2_X1 U499 ( .A1(Key[123]), .A2(Plaintext[123]), .Z(n381) );
  XOR2_X1 U500 ( .A1(Key[124]), .A2(Plaintext[124]), .Z(n382) );
  XOR2_X1 U501 ( .A1(Key[125]), .A2(Plaintext[125]), .Z(n425) );
  XOR2_X1 U502 ( .A1(Key[126]), .A2(Plaintext[126]), .Z(n308) );
  XOR2_X1 U503 ( .A1(Key[127]), .A2(Plaintext[127]), .Z(n309) );
  XOR2_X1 U504 ( .A1(Key[128]), .A2(Plaintext[128]), .Z(n310) );
  XOR2_X1 U505 ( .A1(Key[129]), .A2(Plaintext[129]), .Z(n383) );
  XOR2_X1 U506 ( .A1(Key[130]), .A2(Plaintext[130]), .Z(n384) );
  XOR2_X1 U507 ( .A1(Key[131]), .A2(Plaintext[131]), .Z(n426) );
  XOR2_X1 U508 ( .A1(Key[132]), .A2(Plaintext[132]), .Z(n311) );
  XOR2_X1 U509 ( .A1(Key[133]), .A2(Plaintext[133]), .Z(n312) );
  XOR2_X1 U510 ( .A1(Key[134]), .A2(Plaintext[134]), .Z(n313) );
  XOR2_X1 U511 ( .A1(Key[135]), .A2(Plaintext[135]), .Z(n385) );
  XOR2_X1 U512 ( .A1(Key[136]), .A2(Plaintext[136]), .Z(n386) );
  XOR2_X1 U513 ( .A1(Key[137]), .A2(Plaintext[137]), .Z(n427) );
  XOR2_X1 U514 ( .A1(Key[138]), .A2(Plaintext[138]), .Z(n314) );
  XOR2_X1 U515 ( .A1(Key[139]), .A2(Plaintext[139]), .Z(n315) );
  XOR2_X1 U516 ( .A1(Key[140]), .A2(Plaintext[140]), .Z(n316) );
  XOR2_X1 U517 ( .A1(Key[141]), .A2(Plaintext[141]), .Z(n387) );
  XOR2_X1 U518 ( .A1(Key[142]), .A2(Plaintext[142]), .Z(n388) );
  XOR2_X1 U519 ( .A1(Key[143]), .A2(Plaintext[143]), .Z(n428) );
  XOR2_X1 U520 ( .A1(Key[144]), .A2(Plaintext[144]), .Z(n317) );
  XOR2_X1 U521 ( .A1(Key[145]), .A2(Plaintext[145]), .Z(n318) );
  XOR2_X1 U522 ( .A1(Key[146]), .A2(Plaintext[146]), .Z(n319) );
  XOR2_X1 U523 ( .A1(Key[147]), .A2(Plaintext[147]), .Z(n389) );
  XOR2_X1 U524 ( .A1(Key[148]), .A2(Plaintext[148]), .Z(n390) );
  XOR2_X1 U525 ( .A1(Key[149]), .A2(Plaintext[149]), .Z(n429) );
  XOR2_X1 U526 ( .A1(Key[150]), .A2(Plaintext[150]), .Z(n320) );
  XOR2_X1 U527 ( .A1(Key[151]), .A2(Plaintext[151]), .Z(n321) );
  XOR2_X1 U528 ( .A1(Key[152]), .A2(Plaintext[152]), .Z(n322) );
  XOR2_X1 U529 ( .A1(Key[153]), .A2(Plaintext[153]), .Z(n391) );
  XOR2_X1 U530 ( .A1(Key[154]), .A2(Plaintext[154]), .Z(n392) );
  XOR2_X1 U531 ( .A1(Key[155]), .A2(Plaintext[155]), .Z(n430) );
  XOR2_X1 U532 ( .A1(Key[156]), .A2(Plaintext[156]), .Z(n323) );
  XOR2_X1 U533 ( .A1(Key[157]), .A2(Plaintext[157]), .Z(n324) );
  XOR2_X1 U534 ( .A1(Key[158]), .A2(Plaintext[158]), .Z(n325) );
  XOR2_X1 U535 ( .A1(Key[159]), .A2(Plaintext[159]), .Z(n393) );
  XOR2_X1 U536 ( .A1(Key[160]), .A2(Plaintext[160]), .Z(n394) );
  XOR2_X1 U537 ( .A1(Key[161]), .A2(Plaintext[161]), .Z(n431) );
  XOR2_X1 U538 ( .A1(Key[162]), .A2(Plaintext[162]), .Z(n326) );
  XOR2_X1 U539 ( .A1(Key[163]), .A2(Plaintext[163]), .Z(n327) );
  XOR2_X1 U540 ( .A1(Key[164]), .A2(Plaintext[164]), .Z(n328) );
  XOR2_X1 U541 ( .A1(Key[165]), .A2(Plaintext[165]), .Z(n395) );
  XOR2_X1 U542 ( .A1(Key[166]), .A2(Plaintext[166]), .Z(n396) );
  XOR2_X1 U543 ( .A1(Key[167]), .A2(Plaintext[167]), .Z(n432) );
  XOR2_X1 U544 ( .A1(Key[168]), .A2(Plaintext[168]), .Z(n329) );
  XOR2_X1 U545 ( .A1(Key[169]), .A2(Plaintext[169]), .Z(n330) );
  XOR2_X1 U546 ( .A1(Key[170]), .A2(Plaintext[170]), .Z(n331) );
  XOR2_X1 U547 ( .A1(Key[171]), .A2(Plaintext[171]), .Z(n397) );
  XOR2_X1 U548 ( .A1(Key[172]), .A2(Plaintext[172]), .Z(n398) );
  XOR2_X1 U549 ( .A1(Key[173]), .A2(Plaintext[173]), .Z(n433) );
  XOR2_X1 U550 ( .A1(Key[174]), .A2(Plaintext[174]), .Z(n332) );
  XOR2_X1 U551 ( .A1(Key[175]), .A2(Plaintext[175]), .Z(n333) );
  XOR2_X1 U552 ( .A1(Key[176]), .A2(Plaintext[176]), .Z(n334) );
  XOR2_X1 U553 ( .A1(Key[177]), .A2(Plaintext[177]), .Z(n399) );
  XOR2_X1 U554 ( .A1(Key[178]), .A2(Plaintext[178]), .Z(n400) );
  XOR2_X1 U555 ( .A1(Key[179]), .A2(Plaintext[179]), .Z(n434) );
  XOR2_X1 U556 ( .A1(Key[181]), .A2(Plaintext[181]), .Z(n336) );
  XOR2_X1 U557 ( .A1(Key[182]), .A2(Plaintext[182]), .Z(n337) );
  XOR2_X1 U558 ( .A1(Key[183]), .A2(Plaintext[183]), .Z(n401) );
  XOR2_X1 U559 ( .A1(Key[184]), .A2(Plaintext[184]), .Z(n402) );
  XOR2_X1 U560 ( .A1(Key[185]), .A2(Plaintext[185]), .Z(n435) );
  XOR2_X1 U561 ( .A1(Key[186]), .A2(Plaintext[186]), .Z(n338) );
  XOR2_X1 U562 ( .A1(Key[187]), .A2(Plaintext[187]), .Z(n339) );
  XOR2_X1 U563 ( .A1(Key[188]), .A2(Plaintext[188]), .Z(n340) );
  XOR2_X1 U564 ( .A1(Key[189]), .A2(Plaintext[189]), .Z(n403) );
  XOR2_X1 U565 ( .A1(Key[190]), .A2(Plaintext[190]), .Z(n404) );
  XOR2_X1 U566 ( .A1(Key[191]), .A2(Plaintext[191]), .Z(n436) );
  BUF_X4 \SB2_1_8/BUF_5_0  ( .I(\SB2_1_8/buf_output[5] ), .Z(\RI5[1][143] ) );
  BUF_X4 \SB2_2_25/BUF_5  ( .I(\SB1_2_25/buf_output[5] ), .Z(\SB2_2_25/i0_3 )
         );
  INV_X2 \SB4_14/INV_3  ( .I(\RI3[4][105] ), .ZN(\SB4_14/i0[8] ) );
  NAND4_X2 \SB2_0_20/Component_Function_5/N5  ( .A1(
        \SB2_0_20/Component_Function_5/NAND4_in[0] ), .A2(
        \SB2_0_20/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_0_20/Component_Function_5/NAND4_in[2] ), .A4(
        \SB2_0_20/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB2_0_20/buf_output[5] ) );
  BUF_X4 \SB2_2_20/BUF_5_0  ( .I(\SB2_2_20/buf_output[5] ), .Z(\RI5[2][71] )
         );
  INV_X2 \SB2_0_17/INV_3  ( .I(\SB1_0_19/buf_output[3] ), .ZN(\SB2_0_17/i0[8] ) );
  NAND4_X2 \SB2_1_30/Component_Function_5/N5  ( .A1(
        \SB2_1_30/Component_Function_5/NAND4_in[0] ), .A2(
        \SB2_1_30/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_1_30/Component_Function_5/NAND4_in[2] ), .A4(
        \SB2_1_30/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB2_1_30/buf_output[5] ) );
  NAND4_X2 \SB1_0_19/Component_Function_3/N5  ( .A1(
        \SB1_0_19/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_19/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_19/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_19/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_0_19/buf_output[3] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_41  ( .I(\SB2_1_25/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[41] ) );
  INV_X2 \SB2_0_4/INV_3  ( .I(\RI3[0][165] ), .ZN(\SB2_0_4/i0[8] ) );
  INV_X2 \SB1_0_23/INV_2  ( .I(n271), .ZN(\SB1_0_23/i1[9] ) );
  NAND4_X2 \SB2_2_4/Component_Function_5/N5  ( .A1(
        \SB2_2_4/Component_Function_5/NAND4_in[0] ), .A2(
        \SB2_2_4/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_4/Component_Function_5/NAND4_in[2] ), .A4(
        \SB2_2_4/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB2_2_4/buf_output[5] ) );
  INV_X2 \SB1_1_12/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[119] ), .ZN(
        \SB1_1_12/i1_5 ) );
  INV_X4 \SB3_5/INV_3  ( .I(\SB3_5/i0[10] ), .ZN(\SB3_5/i0[8] ) );
  INV_X2 \SB1_0_9/INV_2  ( .I(n313), .ZN(\SB1_0_9/i1[9] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_191  ( .I(\SB2_3_0/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[191] ) );
  INV_X2 \SB1_3_1/INV_5  ( .I(\MC_ARK_ARC_1_2/buf_output[185] ), .ZN(
        \SB1_3_1/i1_5 ) );
  BUF_X4 \SB1_0_15/BUF_5  ( .I(n421), .Z(\SB1_0_15/i0_3 ) );
  INV_X2 \SB2_1_29/INV_3  ( .I(\SB1_1_31/buf_output[3] ), .ZN(\SB2_1_29/i0[8] ) );
  INV_X2 \SB2_0_12/INV_3  ( .I(\SB1_0_14/buf_output[3] ), .ZN(\SB2_0_12/i0[8] ) );
  INV_X2 \SB1_3_9/INV_3  ( .I(n5502), .ZN(\SB1_3_9/i0[8] ) );
  INV_X2 \SB2_1_13/INV_3  ( .I(\SB1_1_15/buf_output[3] ), .ZN(\SB2_1_13/i0[8] ) );
  INV_X2 \SB2_0_9/INV_3  ( .I(\SB1_0_11/buf_output[3] ), .ZN(\SB2_0_9/i0[8] )
         );
  INV_X2 \SB2_1_20/INV_3  ( .I(\SB1_1_22/buf_output[3] ), .ZN(\SB2_1_20/i0[8] ) );
  INV_X2 \SB1_1_20/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[69] ), .ZN(
        \SB1_1_20/i0[8] ) );
  INV_X2 \SB1_2_30/INV_5  ( .I(\MC_ARK_ARC_1_1/buf_output[11] ), .ZN(
        \SB1_2_30/i1_5 ) );
  NAND4_X2 \SB2_1_6/Component_Function_3/N5  ( .A1(
        \SB2_1_6/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_6/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_6/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_1_6/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_1_6/buf_output[3] ) );
  NAND3_X2 \SB2_2_21/Component_Function_3/N3  ( .A1(\SB2_2_21/i1[9] ), .A2(
        \SB2_2_21/i1_7 ), .A3(\SB2_2_21/i0[10] ), .ZN(
        \SB2_2_21/Component_Function_3/NAND4_in[2] ) );
  BUF_X4 \SB2_1_24/BUF_5  ( .I(\SB1_1_24/buf_output[5] ), .Z(\SB2_1_24/i0_3 )
         );
  NAND3_X2 \SB2_1_6/Component_Function_5/N2  ( .A1(\SB2_1_6/i0_0 ), .A2(
        \SB2_1_6/i0[6] ), .A3(\SB2_1_6/i0[10] ), .ZN(
        \SB2_1_6/Component_Function_5/NAND4_in[1] ) );
  INV_X2 \SB1_2_23/INV_5  ( .I(\MC_ARK_ARC_1_1/buf_output[53] ), .ZN(
        \SB1_2_23/i1_5 ) );
  INV_X2 \SB1_0_15/INV_3  ( .I(n373), .ZN(\SB1_0_15/i0[8] ) );
  BUF_X4 \SB1_0_4/BUF_5  ( .I(n432), .Z(\SB1_0_4/i0_3 ) );
  INV_X2 \SB2_2_28/INV_2  ( .I(\SB1_2_31/buf_output[2] ), .ZN(\SB2_2_28/i1[9] ) );
  BUF_X4 \SB1_0_0/BUF_5_0  ( .I(\SB1_0_0/buf_output[5] ), .Z(\RI3[0][191] ) );
  BUF_X4 \SB2_0_6/BUF_1_0  ( .I(\SB2_0_6/buf_output[1] ), .Z(\RI5[0][175] ) );
  INV_X2 \SB2_1_21/INV_3  ( .I(\SB1_1_23/buf_output[3] ), .ZN(\SB2_1_21/i0[8] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_80  ( .I(\SB2_1_21/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[80] ) );
  BUF_X4 \SB2_2_31/BUF_5_0  ( .I(\SB2_2_31/buf_output[5] ), .Z(\RI5[2][5] ) );
  BUF_X4 \SB2_3_22/BUF_5_0  ( .I(\SB2_3_22/buf_output[5] ), .Z(\RI5[3][59] )
         );
  NAND4_X2 \SB2_1_22/Component_Function_3/N5  ( .A1(
        \SB2_1_22/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_22/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_22/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_1_22/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_1_22/buf_output[3] ) );
  BUF_X4 \SB2_0_20/BUF_1_0  ( .I(\SB2_0_20/buf_output[1] ), .Z(\RI5[0][91] )
         );
  NAND4_X2 \SB2_1_23/Component_Function_4/N5  ( .A1(
        \SB2_1_23/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_23/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_23/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_1_23/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_1_23/buf_output[4] ) );
  INV_X2 \SB2_0_0/INV_3  ( .I(\SB1_0_2/buf_output[3] ), .ZN(\SB2_0_0/i0[8] )
         );
  NAND4_X2 \SB2_3_16/Component_Function_4/N5  ( .A1(
        \SB2_3_16/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_16/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_3_16/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_3_16/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_3_16/buf_output[4] ) );
  INV_X2 \SB1_1_17/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[89] ), .ZN(
        \SB1_1_17/i1_5 ) );
  BUF_X4 \SB1_3_31/BUF_5  ( .I(\RI1[3][5] ), .Z(\SB1_3_31/i0_3 ) );
  INV_X2 \SB2_2_21/INV_5  ( .I(\SB1_2_21/buf_output[5] ), .ZN(\SB2_2_21/i1_5 )
         );
  INV_X2 \SB4_16/INV_2  ( .I(\SB3_19/buf_output[2] ), .ZN(\SB4_16/i1[9] ) );
  INV_X2 \SB2_1_7/INV_2  ( .I(\SB1_1_10/buf_output[2] ), .ZN(\SB2_1_7/i1[9] )
         );
  BUF_X4 \SB2_0_16/BUF_5_0  ( .I(\SB2_0_16/buf_output[5] ), .Z(\RI5[0][95] )
         );
  INV_X2 \SB2_1_6/INV_5  ( .I(\SB1_1_6/buf_output[5] ), .ZN(\SB2_1_6/i1_5 ) );
  BUF_X2 \SB2_3_24/BUF_0  ( .I(\SB1_3_29/buf_output[0] ), .Z(\SB2_3_24/i0[9] )
         );
  INV_X2 \SB2_1_16/INV_3  ( .I(\SB1_1_18/buf_output[3] ), .ZN(\SB2_1_16/i0[8] ) );
  BUF_X4 \SB1_3_2/BUF_5  ( .I(\MC_ARK_ARC_1_2/buf_output[179] ), .Z(
        \SB1_3_2/i0_3 ) );
  INV_X2 \SB1_1_19/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[73] ), .ZN(
        \SB1_1_19/i1_7 ) );
  BUF_X4 \SB2_0_20/BUF_5_0  ( .I(\SB2_0_20/buf_output[5] ), .Z(\RI5[0][71] )
         );
  BUF_X4 \SB1_0_13/BUF_5  ( .I(n423), .Z(\SB1_0_13/i0_3 ) );
  BUF_X4 \SB2_0_24/BUF_5_0  ( .I(\SB2_0_24/buf_output[5] ), .Z(\RI5[0][47] )
         );
  BUF_X4 \SB2_1_19/BUF_5_0  ( .I(\SB2_1_19/buf_output[5] ), .Z(\RI5[1][77] )
         );
  BUF_X4 \SB2_0_14/BUF_5_0  ( .I(\SB2_0_14/buf_output[5] ), .Z(\RI5[0][107] )
         );
  INV_X2 \SB2_2_12/INV_3  ( .I(\SB1_2_14/buf_output[3] ), .ZN(\SB2_2_12/i0[8] ) );
  CLKBUF_X4 \SB1_2_20/BUF_2  ( .I(\MC_ARK_ARC_1_1/buf_output[68] ), .Z(
        \SB1_2_20/i0_0 ) );
  BUF_X4 \SB2_1_15/BUF_3_0  ( .I(\SB2_1_15/buf_output[3] ), .Z(\RI5[1][111] )
         );
  NAND4_X2 \SB2_3_27/Component_Function_3/N5  ( .A1(
        \SB2_3_27/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_27/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_27/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_27/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_3_27/buf_output[3] ) );
  BUF_X2 \SB1_3_0/BUF_0  ( .I(\MC_ARK_ARC_1_2/buf_output[186] ), .Z(
        \SB1_3_0/i0[9] ) );
  BUF_X4 \SB2_0_19/BUF_5_0  ( .I(\SB2_0_19/buf_output[5] ), .Z(\RI5[0][77] )
         );
  INV_X2 \SB1_0_21/INV_2  ( .I(n277), .ZN(\SB1_0_21/i1[9] ) );
  NAND3_X2 \SB1_2_22/Component_Function_2/N3  ( .A1(\SB1_2_22/i0_3 ), .A2(
        \SB1_2_22/i0[8] ), .A3(\SB1_2_22/i0[9] ), .ZN(
        \SB1_2_22/Component_Function_2/NAND4_in[2] ) );
  INV_X4 \SB2_0_29/INV_3  ( .I(\RI3[0][15] ), .ZN(\SB2_0_29/i0[8] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_22  ( .I(\SB2_1_29/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[22] ) );
  BUF_X4 \SB2_0_3/BUF_2_0  ( .I(\SB2_0_3/buf_output[2] ), .Z(\RI5[0][188] ) );
  BUF_X4 \SB1_0_27/BUF_5  ( .I(n409), .Z(\SB1_0_27/i0_3 ) );
  INV_X2 \SB1_0_2/INV_3  ( .I(n399), .ZN(\SB1_0_2/i0[8] ) );
  BUF_X4 \SB2_0_21/BUF_5_0  ( .I(\SB2_0_21/buf_output[5] ), .Z(\RI5[0][65] )
         );
  NAND4_X2 \SB2_0_20/Component_Function_1/N5  ( .A1(
        \SB2_0_20/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_20/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_20/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_20/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_0_20/buf_output[1] ) );
  BUF_X4 \SB2_1_27/BUF_3_0  ( .I(\SB2_1_27/buf_output[3] ), .Z(\RI5[1][39] )
         );
  INV_X2 \SB2_1_29/INV_4  ( .I(\SB2_1_29/i0_4 ), .ZN(\SB2_1_29/i0[7] ) );
  INV_X2 \SB1_2_0/INV_5  ( .I(\MC_ARK_ARC_1_1/buf_output[191] ), .ZN(
        \SB1_2_0/i1_5 ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_2  ( .I(\SB2_2_2/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[2] ) );
  INV_X2 \SB2_3_5/INV_5  ( .I(\SB1_3_5/buf_output[5] ), .ZN(\SB2_3_5/i1_5 ) );
  BUF_X4 \SB2_2_17/BUF_5_0  ( .I(\SB2_2_17/buf_output[5] ), .Z(\RI5[2][89] )
         );
  INV_X2 \SB1_3_16/INV_5  ( .I(\MC_ARK_ARC_1_2/buf_output[95] ), .ZN(
        \SB1_3_16/i1_5 ) );
  NAND4_X2 \SB2_2_29/Component_Function_4/N5  ( .A1(
        \SB2_2_29/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_29/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_2_29/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_2_29/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_2_29/buf_output[4] ) );
  NAND4_X2 \SB2_1_30/Component_Function_4/N5  ( .A1(
        \SB2_1_30/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_30/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_30/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_1_30/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_1_30/buf_output[4] ) );
  BUF_X4 \SB2_1_14/BUF_5_0  ( .I(\SB2_1_14/buf_output[5] ), .Z(\RI5[1][107] )
         );
  NAND4_X2 \SB1_0_4/Component_Function_0/N5  ( .A1(
        \SB1_0_4/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_4/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_4/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_4/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_0_4/buf_output[0] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_41  ( .I(\SB2_3_25/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[41] ) );
  INV_X2 \SB1_3_14/INV_5  ( .I(n3664), .ZN(\SB1_3_14/i1_5 ) );
  NAND3_X2 \SB1_1_22/Component_Function_2/N3  ( .A1(\RI1[1][59] ), .A2(
        \SB1_1_22/i0[8] ), .A3(\SB1_1_22/i0[9] ), .ZN(
        \SB1_1_22/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 \SB1_0_2/BUF_5  ( .I(n434), .Z(\SB1_0_2/i0_3 ) );
  BUF_X4 \SB2_0_17/BUF_5_0  ( .I(\SB2_0_17/buf_output[5] ), .Z(\RI5[0][89] )
         );
  INV_X2 \SB1_0_28/INV_3  ( .I(n347), .ZN(\SB1_0_28/i0[8] ) );
  NAND4_X2 \SB2_1_18/Component_Function_4/N5  ( .A1(
        \SB2_1_18/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_18/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_18/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_1_18/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_1_18/buf_output[4] ) );
  NAND3_X2 \SB1_3_10/Component_Function_3/N4  ( .A1(\SB1_3_10/i1_5 ), .A2(
        \SB1_3_10/i0[8] ), .A3(\SB1_3_10/i3[0] ), .ZN(
        \SB1_3_10/Component_Function_3/NAND4_in[3] ) );
  BUF_X4 \SB2_2_16/BUF_4_0  ( .I(\SB2_2_16/buf_output[4] ), .Z(\RI5[2][100] )
         );
  BUF_X4 \SB1_0_26/BUF_5  ( .I(n410), .Z(\SB1_0_26/i0_3 ) );
  BUF_X4 \SB2_0_23/BUF_5_0  ( .I(\SB2_0_23/buf_output[5] ), .Z(\RI5[0][53] )
         );
  BUF_X4 \SB2_0_1/BUF_4_0  ( .I(\SB2_0_1/buf_output[4] ), .Z(\RI5[0][190] ) );
  INV_X2 \SB1_0_29/INV_2  ( .I(n253), .ZN(\SB1_0_29/i1[9] ) );
  NAND4_X2 \SB1_0_14/Component_Function_0/N5  ( .A1(
        \SB1_0_14/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_14/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_14/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_14/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_0_14/buf_output[0] ) );
  BUF_X4 \SB2_0_13/BUF_5_0  ( .I(\SB2_0_13/buf_output[5] ), .Z(\RI5[0][113] )
         );
  CLKBUF_X4 \SB2_3_10/BUF_3  ( .I(\SB1_3_12/buf_output[3] ), .Z(
        \SB2_3_10/i0[10] ) );
  BUF_X4 \SB2_0_16/BUF_0_0  ( .I(\SB2_0_16/buf_output[0] ), .Z(\RI5[0][120] )
         );
  BUF_X4 \SB2_0_10/BUF_4_0  ( .I(\SB2_0_10/buf_output[4] ), .Z(\RI5[0][136] )
         );
  BUF_X4 \SB2_0_15/BUF_5_0  ( .I(\SB2_0_15/buf_output[5] ), .Z(\RI5[0][101] )
         );
  NAND3_X2 \SB1_1_8/Component_Function_3/N4  ( .A1(n3647), .A2(\SB1_1_8/i0[8] ), .A3(\SB1_1_8/i3[0] ), .ZN(\SB1_1_8/Component_Function_3/NAND4_in[3] ) );
  BUF_X4 \SB2_0_1/BUF_5_0  ( .I(\SB2_0_1/buf_output[5] ), .Z(\RI5[0][185] ) );
  INV_X2 \SB1_0_31/INV_2  ( .I(n247), .ZN(\SB1_0_31/i1[9] ) );
  BUF_X4 \SB2_0_9/BUF_2_0  ( .I(\SB2_0_9/buf_output[2] ), .Z(\RI5[0][152] ) );
  INV_X2 \SB2_2_6/INV_3  ( .I(\SB1_2_8/buf_output[3] ), .ZN(\SB2_2_6/i0[8] )
         );
  INV_X2 \SB1_3_14/INV_2  ( .I(\MC_ARK_ARC_1_2/buf_output[104] ), .ZN(
        \SB1_3_14/i1[9] ) );
  NAND3_X2 \SB1_0_31/Component_Function_3/N2  ( .A1(\SB1_0_31/i0_0 ), .A2(
        \SB1_0_31/i0_3 ), .A3(\SB1_0_31/i0_4 ), .ZN(
        \SB1_0_31/Component_Function_3/NAND4_in[1] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_81  ( .I(\SB2_0_20/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[81] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_36  ( .I(\SB2_3_30/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[36] ) );
  NAND3_X2 \SB2_1_30/Component_Function_5/N4  ( .A1(\SB2_1_30/i0[9] ), .A2(
        \SB2_1_30/i0[6] ), .A3(\SB2_1_30/i0_4 ), .ZN(
        \SB2_1_30/Component_Function_5/NAND4_in[3] ) );
  BUF_X4 \SB2_0_17/BUF_3_0  ( .I(\SB2_0_17/buf_output[3] ), .Z(\RI5[0][99] )
         );
  BUF_X4 \SB2_2_17/BUF_4_0  ( .I(\SB2_2_17/buf_output[4] ), .Z(\RI5[2][94] )
         );
  BUF_X4 \SB2_0_31/BUF_5_0  ( .I(\SB2_0_31/buf_output[5] ), .Z(\RI5[0][5] ) );
  NAND4_X2 \SB2_2_26/Component_Function_0/N5  ( .A1(
        \SB2_2_26/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_26/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_26/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_26/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB2_2_26/buf_output[0] ) );
  BUF_X4 \SB2_0_8/BUF_3_0  ( .I(\SB2_0_8/buf_output[3] ), .Z(\RI5[0][153] ) );
  BUF_X4 \SB2_0_11/BUF_3_0  ( .I(\SB2_0_11/buf_output[3] ), .Z(\RI5[0][135] )
         );
  BUF_X4 \SB2_0_19/BUF_0_0  ( .I(\SB2_0_19/buf_output[0] ), .Z(\RI5[0][102] )
         );
  INV_X2 \SB2_0_29/INV_0  ( .I(n1905), .ZN(\SB2_0_29/i3[0] ) );
  BUF_X4 \SB1_0_31/BUF_3_0  ( .I(\SB1_0_31/buf_output[3] ), .Z(\RI3[0][15] )
         );
  BUF_X4 \SB1_1_3/BUF_5  ( .I(\RI1[1][173] ), .Z(\SB1_1_3/i0_3 ) );
  BUF_X4 \SB1_3_26/BUF_5  ( .I(\MC_ARK_ARC_1_2/buf_output[35] ), .Z(
        \SB1_3_26/i0_3 ) );
  BUF_X4 \SB1_2_11/BUF_5  ( .I(\MC_ARK_ARC_1_1/buf_output[125] ), .Z(
        \SB1_2_11/i0_3 ) );
  BUF_X4 \SB2_0_3/BUF_5_0  ( .I(\SB2_0_3/buf_output[5] ), .Z(\RI5[0][173] ) );
  NAND3_X2 \SB1_2_30/Component_Function_2/N1  ( .A1(\SB1_2_30/i1_5 ), .A2(
        \SB1_2_30/i0[10] ), .A3(\SB1_2_30/i1[9] ), .ZN(
        \SB1_2_30/Component_Function_2/NAND4_in[0] ) );
  CLKBUF_X4 \SB1_3_25/BUF_2  ( .I(\MC_ARK_ARC_1_2/buf_output[38] ), .Z(
        \SB1_3_25/i0_0 ) );
  NAND4_X2 \SB2_0_6/Component_Function_3/N5  ( .A1(
        \SB2_0_6/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_6/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_0_6/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_0_6/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_0_6/buf_output[3] ) );
  BUF_X4 \SB2_0_16/BUF_4_0  ( .I(\SB2_0_16/buf_output[4] ), .Z(\RI5[0][100] )
         );
  BUF_X4 \SB2_0_10/BUF_5_0  ( .I(\SB2_0_10/buf_output[5] ), .Z(\RI5[0][131] )
         );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_56  ( .I(\SB2_3_25/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[56] ) );
  INV_X2 \SB2_1_21/INV_5  ( .I(\SB1_1_21/buf_output[5] ), .ZN(\SB2_1_21/i1_5 )
         );
  NAND4_X2 \SB1_0_9/Component_Function_1/N5  ( .A1(
        \SB1_0_9/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_9/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_9/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_9/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_0_9/buf_output[1] ) );
  BUF_X4 \SB2_0_8/BUF_5_0  ( .I(\SB2_0_8/buf_output[5] ), .Z(\RI5[0][143] ) );
  BUF_X4 \SB2_0_21/BUF_4_0  ( .I(\SB2_0_21/buf_output[4] ), .Z(\RI5[0][70] )
         );
  BUF_X2 \SB1_1_21/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[60] ), .Z(
        \SB1_1_21/i0[9] ) );
  INV_X2 \SB1_0_16/INV_3  ( .I(n371), .ZN(\SB1_0_16/i0[8] ) );
  NAND3_X2 \SB1_0_16/Component_Function_3/N3  ( .A1(\SB1_0_16/i1[9] ), .A2(
        \SB1_0_16/i1_7 ), .A3(\SB1_0_16/i0[10] ), .ZN(
        \SB1_0_16/Component_Function_3/NAND4_in[2] ) );
  BUF_X4 \SB2_0_0/BUF_5_0  ( .I(\SB2_0_0/buf_output[5] ), .Z(\RI5[0][191] ) );
  BUF_X4 \SB2_0_1/BUF_2_0  ( .I(\SB2_0_1/buf_output[2] ), .Z(\RI5[0][8] ) );
  NAND4_X2 \SB2_2_4/Component_Function_4/N5  ( .A1(
        \SB2_2_4/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_4/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_2_4/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_2_4/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_2_4/buf_output[4] ) );
  CLKBUF_X4 \SB2_0_29/BUF_2  ( .I(\SB1_0_0/buf_output[2] ), .Z(\SB2_0_29/i0_0 ) );
  NAND3_X2 \SB1_1_0/Component_Function_3/N1  ( .A1(\SB1_1_0/i1[9] ), .A2(
        \SB1_1_0/i0_3 ), .A3(\SB1_1_0/i0[6] ), .ZN(
        \SB1_1_0/Component_Function_3/NAND4_in[0] ) );
  INV_X2 \SB1_0_7/INV_3  ( .I(n389), .ZN(\SB1_0_7/i0[8] ) );
  NAND3_X2 \SB1_0_4/Component_Function_3/N2  ( .A1(\SB1_0_4/i0_0 ), .A2(
        \SB1_0_4/i0_3 ), .A3(\SB1_0_4/i0_4 ), .ZN(
        \SB1_0_4/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 \SB2_0_28/Component_Function_4/N5  ( .A1(
        \SB2_0_28/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_28/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_28/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_0_28/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_0_28/buf_output[4] ) );
  BUF_X4 \SB2_0_15/BUF_2_0  ( .I(\SB2_0_15/buf_output[2] ), .Z(\RI5[0][116] )
         );
  BUF_X4 \SB2_2_11/BUF_1_0  ( .I(\SB2_2_11/buf_output[1] ), .Z(\RI5[2][145] )
         );
  BUF_X4 \SB1_0_25/BUF_4  ( .I(n354), .Z(\SB1_0_25/i0_4 ) );
  INV_X2 \SB2_2_19/INV_5  ( .I(\SB1_2_19/buf_output[5] ), .ZN(\SB2_2_19/i1_5 )
         );
  INV_X2 \SB1_1_10/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[131] ), .ZN(
        \SB1_1_10/i1_5 ) );
  NAND4_X2 \SB2_2_24/Component_Function_0/N5  ( .A1(
        \SB2_2_24/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_24/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_24/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_24/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB2_2_24/buf_output[0] ) );
  NAND4_X2 \SB2_0_23/Component_Function_1/N5  ( .A1(
        \SB2_0_23/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_23/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_23/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_23/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_0_23/buf_output[1] ) );
  NAND4_X2 \SB1_0_1/Component_Function_1/N5  ( .A1(
        \SB1_0_1/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_1/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_1/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_1/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_0_1/buf_output[1] ) );
  NAND3_X2 \SB2_0_11/Component_Function_4/N2  ( .A1(\SB2_0_11/i3[0] ), .A2(
        \SB2_0_11/i0_0 ), .A3(\SB2_0_11/i1_7 ), .ZN(
        \SB2_0_11/Component_Function_4/NAND4_in[1] ) );
  BUF_X4 \SB2_0_11/BUF_5_0  ( .I(\SB2_0_11/buf_output[5] ), .Z(\RI5[0][125] )
         );
  NAND2_X2 \SB2_0_11/Component_Function_5/N1  ( .A1(\SB2_0_11/i0_0 ), .A2(
        \SB2_0_11/i3[0] ), .ZN(\SB2_0_11/Component_Function_5/NAND4_in[0] ) );
  INV_X2 \SB1_0_14/INV_3  ( .I(n375), .ZN(\SB1_0_14/i0[8] ) );
  BUF_X4 \SB2_0_7/BUF_5_0  ( .I(\SB2_0_7/buf_output[5] ), .Z(\RI5[0][149] ) );
  NAND3_X2 \SB1_0_14/Component_Function_5/N3  ( .A1(\SB1_0_14/i1[9] ), .A2(
        \SB1_0_14/i0_4 ), .A3(\SB1_0_14/i0_3 ), .ZN(
        \SB1_0_14/Component_Function_5/NAND4_in[2] ) );
  BUF_X4 \SB2_2_14/BUF_5_0  ( .I(\SB2_2_14/buf_output[5] ), .Z(\RI5[2][107] )
         );
  NAND4_X2 \SB2_3_26/Component_Function_1/N5  ( .A1(
        \SB2_3_26/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_26/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_26/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_26/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_3_26/buf_output[1] ) );
  BUF_X4 \SB2_0_12/BUF_5_0  ( .I(\SB2_0_12/buf_output[5] ), .Z(\RI5[0][119] )
         );
  NAND3_X2 \SB2_2_23/Component_Function_2/N2  ( .A1(\SB2_2_23/i0_3 ), .A2(
        \SB2_2_23/i0[10] ), .A3(\SB2_2_23/i0[6] ), .ZN(
        \SB2_2_23/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 \SB2_1_17/Component_Function_2/N4  ( .A1(\SB2_1_17/i1_5 ), .A2(
        \SB2_1_17/i0_0 ), .A3(\SB2_1_17/i0_4 ), .ZN(
        \SB2_1_17/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 \SB1_2_23/Component_Function_5/N3  ( .A1(\SB1_2_23/i1[9] ), .A2(
        \SB1_2_23/i0_4 ), .A3(\SB1_2_23/i0_3 ), .ZN(
        \SB1_2_23/Component_Function_5/NAND4_in[2] ) );
  INV_X2 \SB1_1_19/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[77] ), .ZN(
        \SB1_1_19/i1_5 ) );
  BUF_X4 \SB2_0_8/BUF_1_0  ( .I(\SB2_0_8/buf_output[1] ), .Z(\RI5[0][163] ) );
  BUF_X4 \SB2_0_22/BUF_5_0  ( .I(\SB2_0_22/buf_output[5] ), .Z(\RI5[0][59] )
         );
  BUF_X2 U56 ( .I(Key[186]), .Z(n15) );
  BUF_X4 \SB1_0_18/BUF_4_0  ( .I(\SB1_0_18/buf_output[4] ), .Z(\RI3[0][88] )
         );
  INV_X2 \SB1_0_18/INV_2  ( .I(n286), .ZN(\SB1_0_18/i1[9] ) );
  NAND4_X2 \SB2_1_30/Component_Function_0/N5  ( .A1(
        \SB2_1_30/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_30/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_30/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_30/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB2_1_30/buf_output[0] ) );
  BUF_X4 \SB2_2_14/BUF_4_0  ( .I(\SB2_2_14/buf_output[4] ), .Z(\RI5[2][112] )
         );
  NAND4_X2 \SB2_0_15/Component_Function_1/N5  ( .A1(
        \SB2_0_15/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_15/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_15/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_15/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_0_15/buf_output[1] ) );
  NAND3_X2 \SB2_0_15/Component_Function_1/N4  ( .A1(\SB2_0_15/i1_7 ), .A2(
        \SB2_0_15/i0[8] ), .A3(\RI3[0][100] ), .ZN(
        \SB2_0_15/Component_Function_1/NAND4_in[3] ) );
  BUF_X4 \SB2_1_7/BUF_2_0  ( .I(\SB2_1_7/buf_output[2] ), .Z(\RI5[1][164] ) );
  INV_X2 \SB1_2_10/INV_5  ( .I(\MC_ARK_ARC_1_1/buf_output[131] ), .ZN(
        \SB1_2_10/i1_5 ) );
  INV_X2 \SB3_12/INV_5  ( .I(\MC_ARK_ARC_1_3/buf_output[119] ), .ZN(
        \SB3_12/i1_5 ) );
  BUF_X4 \SB2_3_25/BUF_4_0  ( .I(\SB2_3_25/buf_output[4] ), .Z(\RI5[3][46] )
         );
  NAND3_X2 \SB2_2_21/Component_Function_2/N3  ( .A1(\SB2_2_21/i0_3 ), .A2(
        \SB2_2_21/i0[8] ), .A3(\SB2_2_21/i0[9] ), .ZN(
        \SB2_2_21/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 \SB1_0_11/Component_Function_0/N5  ( .A1(
        \SB1_0_11/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_11/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_11/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_11/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_0_11/buf_output[0] ) );
  NAND4_X2 \SB2_2_6/Component_Function_3/N5  ( .A1(
        \SB2_2_6/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_6/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_2_6/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_2_6/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_2_6/buf_output[3] ) );
  NAND3_X2 \SB2_1_12/Component_Function_2/N3  ( .A1(\SB2_1_12/i0_3 ), .A2(
        \SB2_1_12/i0[8] ), .A3(\SB2_1_12/i0[9] ), .ZN(
        \SB2_1_12/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 \SB2_1_21/Component_Function_3/N3  ( .A1(\SB2_1_21/i1[9] ), .A2(
        \SB2_1_21/i1_7 ), .A3(\SB2_1_21/i0[10] ), .ZN(
        \SB2_1_21/Component_Function_3/NAND4_in[2] ) );
  NAND4_X2 \SB2_0_10/Component_Function_1/N5  ( .A1(
        \SB2_0_10/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_10/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_10/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_10/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_0_10/buf_output[1] ) );
  NAND4_X2 \SB2_2_13/Component_Function_0/N5  ( .A1(
        \SB2_2_13/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_2_13/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_13/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_13/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB2_2_13/buf_output[0] ) );
  INV_X2 \SB2_1_19/INV_5  ( .I(\SB1_1_19/buf_output[5] ), .ZN(\SB2_1_19/i1_5 )
         );
  INV_X2 \SB1_0_17/INV_3  ( .I(n369), .ZN(\SB1_0_17/i0[8] ) );
  BUF_X4 \SB2_0_13/BUF_3_0  ( .I(\SB2_0_13/buf_output[3] ), .Z(\RI5[0][123] )
         );
  BUF_X4 \SB2_2_23/BUF_5  ( .I(\SB1_2_23/buf_output[5] ), .Z(\SB2_2_23/i0_3 )
         );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_110  ( .I(\SB2_3_16/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[110] ) );
  BUF_X4 \SB2_0_12/BUF_4_0  ( .I(\SB2_0_12/buf_output[4] ), .Z(\RI5[0][124] )
         );
  BUF_X4 \SB1_0_4/BUF_4_0  ( .I(\SB1_0_4/buf_output[4] ), .Z(\RI3[0][172] ) );
  NAND4_X2 \SB1_0_4/Component_Function_4/N5  ( .A1(
        \SB1_0_4/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_4/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_4/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_4/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_0_4/buf_output[4] ) );
  BUF_X4 \SB2_0_16/BUF_5  ( .I(\RI3[0][95] ), .Z(\SB2_0_16/i0_3 ) );
  NAND3_X2 \SB3_7/Component_Function_1/N4  ( .A1(\SB3_7/i1_7 ), .A2(
        \SB3_7/i0[8] ), .A3(\SB3_7/i0_4 ), .ZN(
        \SB3_7/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 \SB1_2_23/Component_Function_2/N2  ( .A1(\SB1_2_23/i0_3 ), .A2(
        \SB1_2_23/i0[10] ), .A3(\SB1_2_23/i0[6] ), .ZN(
        \SB1_2_23/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 \SB2_0_17/BUF_2_0  ( .I(\SB2_0_17/buf_output[2] ), .Z(\RI5[0][104] )
         );
  INV_X2 \SB1_2_5/INV_5  ( .I(\MC_ARK_ARC_1_1/buf_output[161] ), .ZN(
        \SB1_2_5/i1_5 ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_89  ( .I(\SB2_1_17/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[89] ) );
  CLKBUF_X4 \SB2_0_23/BUF_2  ( .I(\RI3[0][50] ), .Z(\SB2_0_23/i0_0 ) );
  INV_X2 \SB1_0_4/INV_2  ( .I(n328), .ZN(\SB1_0_4/i1[9] ) );
  NAND4_X2 \SB1_0_10/Component_Function_0/N5  ( .A1(
        \SB1_0_10/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_10/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_10/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_10/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_0_10/buf_output[0] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_125  ( .I(\SB2_2_11/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[125] ) );
  INV_X2 \SB2_0_23/INV_5  ( .I(\SB1_0_23/buf_output[5] ), .ZN(\SB2_0_23/i1_5 )
         );
  BUF_X4 \SB2_0_1/BUF_0_0  ( .I(\SB2_0_1/buf_output[0] ), .Z(\RI5[0][18] ) );
  BUF_X4 \SB2_3_23/BUF_5  ( .I(\SB1_3_23/buf_output[5] ), .Z(\SB2_3_23/i0_3 )
         );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_83  ( .I(\SB2_2_18/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[83] ) );
  NAND3_X2 \SB2_2_8/Component_Function_3/N4  ( .A1(\SB2_2_8/i1_5 ), .A2(
        \SB2_2_8/i0[8] ), .A3(\SB2_2_8/i3[0] ), .ZN(
        \SB2_2_8/Component_Function_3/NAND4_in[3] ) );
  NAND4_X2 \SB2_2_20/Component_Function_1/N5  ( .A1(
        \SB2_2_20/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_20/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_20/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_20/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_2_20/buf_output[1] ) );
  NAND4_X2 \SB2_3_26/Component_Function_3/N5  ( .A1(
        \SB2_3_26/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_26/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_26/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_26/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_3_26/buf_output[3] ) );
  CLKBUF_X4 \SB2_0_17/BUF_3  ( .I(\SB1_0_19/buf_output[3] ), .Z(
        \SB2_0_17/i0[10] ) );
  INV_X2 \SB1_0_19/INV_3  ( .I(n365), .ZN(\SB1_0_19/i0[8] ) );
  BUF_X4 \SB2_0_15/BUF_1_0  ( .I(\SB2_0_15/buf_output[1] ), .Z(\RI5[0][121] )
         );
  INV_X2 \SB2_1_17/INV_5  ( .I(\SB1_1_17/buf_output[5] ), .ZN(\SB2_1_17/i1_5 )
         );
  NAND3_X2 \SB2_1_24/Component_Function_5/N2  ( .A1(\SB2_1_24/i0_0 ), .A2(
        \SB2_1_24/i0[6] ), .A3(\SB2_1_24/i0[10] ), .ZN(
        \SB2_1_24/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 \SB2_1_26/Component_Function_3/N2  ( .A1(\SB2_1_26/i0_0 ), .A2(
        \SB2_1_26/i0_3 ), .A3(\SB2_1_26/i0_4 ), .ZN(
        \SB2_1_26/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 \SB2_2_15/Component_Function_1/N5  ( .A1(
        \SB2_2_15/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_15/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_15/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_15/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_2_15/buf_output[1] ) );
  NAND4_X2 \SB2_1_14/Component_Function_1/N5  ( .A1(
        \SB2_1_14/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_14/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_14/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_14/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_1_14/buf_output[1] ) );
  INV_X2 \SB1_2_13/INV_5  ( .I(n5526), .ZN(\SB1_2_13/i1_5 ) );
  CLKBUF_X4 \SB1_0_23/BUF_2  ( .I(n271), .Z(\SB1_0_23/i0_0 ) );
  CLKBUF_X4 \SB1_0_17/BUF_3  ( .I(n369), .Z(\SB1_0_17/i0[10] ) );
  BUF_X4 \SB2_2_24/BUF_4_0  ( .I(\SB2_2_24/buf_output[4] ), .Z(\RI5[2][52] )
         );
  NAND3_X2 \SB2_2_17/Component_Function_2/N3  ( .A1(\SB2_2_17/i0_3 ), .A2(
        \SB2_2_17/i0[8] ), .A3(\SB2_2_17/i0[9] ), .ZN(
        \SB2_2_17/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 \SB1_2_25/BUF_5  ( .I(\MC_ARK_ARC_1_1/buf_output[41] ), .Z(
        \SB1_2_25/i0_3 ) );
  NAND3_X2 \SB2_1_24/Component_Function_2/N2  ( .A1(\SB2_1_24/i0_3 ), .A2(
        \SB2_1_24/i0[10] ), .A3(\SB2_1_24/i0[6] ), .ZN(
        \SB2_1_24/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 \SB1_2_30/Component_Function_2/N3  ( .A1(\SB1_2_30/i0_3 ), .A2(
        \SB1_2_30/i0[8] ), .A3(\SB1_2_30/i0[9] ), .ZN(
        \SB1_2_30/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 \SB1_0_17/Component_Function_2/N2  ( .A1(\SB1_0_17/i0_3 ), .A2(
        \SB1_0_17/i0[10] ), .A3(\SB1_0_17/i0[6] ), .ZN(
        \SB1_0_17/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 \SB1_3_24/Component_Function_2/N3  ( .A1(\SB1_3_24/i0_3 ), .A2(
        \SB1_3_24/i0[8] ), .A3(\SB1_3_24/i0[9] ), .ZN(
        \SB1_3_24/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 \SB2_0_9/Component_Function_3/N1  ( .A1(\SB2_0_9/i1[9] ), .A2(
        \SB2_0_9/i0_3 ), .A3(\SB2_0_9/i0[6] ), .ZN(
        \SB2_0_9/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 \SB2_1_19/BUF_5  ( .I(\SB1_1_19/buf_output[5] ), .Z(\SB2_1_19/i0_3 )
         );
  BUF_X4 \SB1_2_17/BUF_5  ( .I(\MC_ARK_ARC_1_1/buf_output[89] ), .Z(
        \SB1_2_17/i0_3 ) );
  INV_X2 \SB2_1_16/INV_1  ( .I(\SB1_1_20/buf_output[1] ), .ZN(\SB2_1_16/i1_7 )
         );
  NAND2_X2 \SB2_2_8/Component_Function_5/N1  ( .A1(\SB2_2_8/i0_0 ), .A2(
        \SB2_2_8/i3[0] ), .ZN(\SB2_2_8/Component_Function_5/NAND4_in[0] ) );
  NAND4_X2 \SB2_0_11/Component_Function_4/N5  ( .A1(
        \SB2_0_11/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_11/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_11/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_0_11/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_0_11/buf_output[4] ) );
  BUF_X4 \SB2_0_31/BUF_1_0  ( .I(\SB2_0_31/buf_output[1] ), .Z(\RI5[0][25] )
         );
  NAND3_X2 \SB2_2_16/Component_Function_3/N4  ( .A1(\SB2_2_16/i1_5 ), .A2(
        \SB2_2_16/i0[8] ), .A3(\SB2_2_16/i3[0] ), .ZN(
        \SB2_2_16/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 \SB1_2_19/Component_Function_5/N4  ( .A1(\SB1_2_19/i0[9] ), .A2(
        \SB1_2_19/i0[6] ), .A3(\SB1_2_19/i0_4 ), .ZN(
        \SB1_2_19/Component_Function_5/NAND4_in[3] ) );
  INV_X2 \SB1_3_24/INV_5  ( .I(\MC_ARK_ARC_1_2/buf_output[47] ), .ZN(
        \SB1_3_24/i1_5 ) );
  CLKBUF_X4 \SB1_0_9/BUF_2  ( .I(n5517), .Z(\SB1_0_9/i0_0 ) );
  BUF_X2 U115 ( .I(Key[120]), .Z(n38) );
  BUF_X4 \SB2_0_21/BUF_2_0  ( .I(\SB2_0_21/buf_output[2] ), .Z(\RI5[0][80] )
         );
  NAND4_X2 \SB1_0_9/Component_Function_4/N5  ( .A1(
        \SB1_0_9/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_9/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_9/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_9/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_0_9/buf_output[4] ) );
  NAND3_X2 \SB2_2_21/Component_Function_1/N2  ( .A1(\SB2_2_21/i0_3 ), .A2(
        \SB2_2_21/i1_7 ), .A3(\SB2_2_21/i0[8] ), .ZN(
        \SB2_2_21/Component_Function_1/NAND4_in[1] ) );
  BUF_X4 \SB2_0_24/BUF_0_0  ( .I(\SB2_0_24/buf_output[0] ), .Z(\RI5[0][72] )
         );
  NAND3_X2 \SB1_2_13/Component_Function_5/N3  ( .A1(\SB1_2_13/i1[9] ), .A2(
        \SB1_2_13/i0_4 ), .A3(\SB1_2_13/i0_3 ), .ZN(
        \SB1_2_13/Component_Function_5/NAND4_in[2] ) );
  INV_X2 \SB1_3_13/INV_5  ( .I(\MC_ARK_ARC_1_2/buf_output[113] ), .ZN(
        \SB1_3_13/i1_5 ) );
  NAND2_X2 \SB2_3_4/Component_Function_5/N1  ( .A1(\SB2_3_4/i0_0 ), .A2(
        \SB2_3_4/i3[0] ), .ZN(\SB2_3_4/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB2_2_18/Component_Function_3/N3  ( .A1(\SB2_2_18/i1[9] ), .A2(
        \SB2_2_18/i1_7 ), .A3(\SB2_2_18/i0[10] ), .ZN(
        \SB2_2_18/Component_Function_3/NAND4_in[2] ) );
  BUF_X4 \SB2_0_1/BUF_5  ( .I(\SB1_0_1/buf_output[5] ), .Z(\SB2_0_1/i0_3 ) );
  BUF_X4 \SB1_0_17/BUF_2_0  ( .I(\SB1_0_17/buf_output[2] ), .Z(\RI3[0][104] )
         );
  INV_X2 \SB2_2_15/INV_5  ( .I(\SB1_2_15/buf_output[5] ), .ZN(\SB2_2_15/i1_5 )
         );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_110  ( .I(\SB2_1_16/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[110] ) );
  NAND3_X2 \SB1_3_8/Component_Function_2/N2  ( .A1(\SB1_3_8/i0_3 ), .A2(
        \SB1_3_8/i0[10] ), .A3(\SB1_3_8/i0[6] ), .ZN(
        \SB1_3_8/Component_Function_2/NAND4_in[1] ) );
  INV_X2 \SB1_0_12/INV_2  ( .I(n304), .ZN(\SB1_0_12/i1[9] ) );
  NAND4_X2 \SB2_3_10/Component_Function_1/N5  ( .A1(
        \SB2_3_10/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_10/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_10/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_10/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_3_10/buf_output[1] ) );
  BUF_X2 U61 ( .I(Key[178]), .Z(n73) );
  INV_X2 \SB1_0_28/INV_2  ( .I(n256), .ZN(\SB1_0_28/i1[9] ) );
  NAND3_X2 \SB2_1_22/Component_Function_3/N3  ( .A1(\SB2_1_22/i1[9] ), .A2(
        \SB2_1_22/i1_7 ), .A3(\SB2_1_22/i0[10] ), .ZN(
        \SB2_1_22/Component_Function_3/NAND4_in[2] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_131  ( .I(\SB2_2_10/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[131] ) );
  INV_X2 \SB1_0_29/INV_3  ( .I(n345), .ZN(\SB1_0_29/i0[8] ) );
  INV_X2 \SB2_0_28/INV_3  ( .I(\SB1_0_30/buf_output[3] ), .ZN(\SB2_0_28/i0[8] ) );
  BUF_X4 \SB2_0_22/BUF_2_0  ( .I(\SB2_0_22/buf_output[2] ), .Z(\RI5[0][74] )
         );
  NAND2_X2 \SB1_0_19/Component_Function_5/N1  ( .A1(\SB1_0_19/i0_0 ), .A2(
        \SB1_0_19/i3[0] ), .ZN(\SB1_0_19/Component_Function_5/NAND4_in[0] ) );
  NAND2_X2 \SB1_1_13/Component_Function_0/N1  ( .A1(\SB1_1_13/i0[10] ), .A2(
        \SB1_1_13/i0[9] ), .ZN(\SB1_1_13/Component_Function_0/NAND4_in[0] ) );
  BUF_X4 \SB1_0_12/BUF_2_0  ( .I(\SB1_0_12/buf_output[2] ), .Z(\RI3[0][134] )
         );
  NAND4_X2 \SB2_0_28/Component_Function_3/N5  ( .A1(
        \SB2_0_28/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_28/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_0_28/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_0_28/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_0_28/buf_output[3] ) );
  NAND3_X2 \SB1_0_9/Component_Function_3/N2  ( .A1(\SB1_0_9/i0_0 ), .A2(
        \SB1_0_9/i0_3 ), .A3(\SB1_0_9/i0_4 ), .ZN(
        \SB1_0_9/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 \SB1_2_0/Component_Function_5/N3  ( .A1(\SB1_2_0/i1[9] ), .A2(
        \SB1_2_0/i0_4 ), .A3(\SB1_2_0/i0_3 ), .ZN(
        \SB1_2_0/Component_Function_5/NAND4_in[2] ) );
  BUF_X4 \SB2_2_21/BUF_3_0  ( .I(\SB2_2_21/buf_output[3] ), .Z(\RI5[2][75] )
         );
  BUF_X4 \SB2_0_18/BUF_5_0  ( .I(\SB2_0_18/buf_output[5] ), .Z(\RI5[0][83] )
         );
  INV_X2 \SB1_1_29/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[17] ), .ZN(
        \SB1_1_29/i1_5 ) );
  NAND3_X2 \SB1_3_11/Component_Function_4/N4  ( .A1(\SB1_3_11/i1[9] ), .A2(
        n2908), .A3(\SB1_3_11/i0_4 ), .ZN(
        \SB1_3_11/Component_Function_4/NAND4_in[3] ) );
  NAND4_X2 \SB2_3_14/Component_Function_1/N5  ( .A1(
        \SB2_3_14/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_14/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_14/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_14/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_3_14/buf_output[1] ) );
  BUF_X4 \SB2_1_1/BUF_5  ( .I(\SB1_1_1/buf_output[5] ), .Z(\SB2_1_1/i0_3 ) );
  NAND4_X2 \SB2_0_9/Component_Function_1/N5  ( .A1(
        \SB2_0_9/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_9/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_9/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_9/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_0_9/buf_output[1] ) );
  INV_X2 \SB1_2_9/INV_5  ( .I(\MC_ARK_ARC_1_1/buf_output[137] ), .ZN(
        \SB1_2_9/i1_5 ) );
  BUF_X2 \SB2_3_15/BUF_2  ( .I(\SB1_3_18/buf_output[2] ), .Z(\SB2_3_15/i0_0 )
         );
  NAND3_X2 \SB2_2_8/Component_Function_1/N2  ( .A1(\SB2_2_8/i0_3 ), .A2(
        \SB2_2_8/i1_7 ), .A3(\SB2_2_8/i0[8] ), .ZN(
        \SB2_2_8/Component_Function_1/NAND4_in[1] ) );
  NAND4_X2 \SB2_0_19/Component_Function_0/N5  ( .A1(
        \SB2_0_19/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_19/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_19/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_19/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB2_0_19/buf_output[0] ) );
  NAND3_X2 \SB1_2_30/Component_Function_4/N2  ( .A1(\SB1_2_30/i3[0] ), .A2(
        \SB1_2_30/i0_0 ), .A3(\SB1_2_30/i1_7 ), .ZN(
        \SB1_2_30/Component_Function_4/NAND4_in[1] ) );
  NAND4_X2 \SB2_3_12/Component_Function_0/N5  ( .A1(
        \SB2_3_12/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_3_12/Component_Function_0/NAND4_in[0] ), .A3(
        \SB2_3_12/Component_Function_0/NAND4_in[3] ), .A4(
        \SB2_3_12/Component_Function_0/NAND4_in[2] ), .ZN(
        \SB2_3_12/buf_output[0] ) );
  NAND3_X2 \SB1_1_22/Component_Function_2/N4  ( .A1(\SB1_1_22/i1_5 ), .A2(
        \SB1_1_22/i0_0 ), .A3(\SB1_1_22/i0_4 ), .ZN(
        \SB1_1_22/Component_Function_2/NAND4_in[3] ) );
  NAND4_X2 \SB2_2_31/Component_Function_2/N5  ( .A1(
        \SB2_2_31/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_31/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_2_31/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_2_31/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB2_2_31/buf_output[2] ) );
  NAND2_X2 \SB1_2_30/Component_Function_5/N1  ( .A1(\SB1_2_30/i0_0 ), .A2(
        \SB1_2_30/i3[0] ), .ZN(\SB1_2_30/Component_Function_5/NAND4_in[0] ) );
  INV_X2 \SB1_2_30/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[6] ), .ZN(
        \SB1_2_30/i3[0] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_112  ( .I(\SB2_0_14/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[112] ) );
  BUF_X4 \SB2_0_5/BUF_5_0  ( .I(\SB2_0_5/buf_output[5] ), .Z(\RI5[0][161] ) );
  CLKBUF_X4 \SB2_3_5/BUF_2  ( .I(\SB1_3_8/buf_output[2] ), .Z(\SB2_3_5/i0_0 )
         );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_6  ( .I(\SB2_2_3/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[6] ) );
  NAND4_X2 \SB2_2_17/Component_Function_2/N5  ( .A1(
        \SB2_2_17/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_17/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_2_17/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_2_17/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_2_17/buf_output[2] ) );
  INV_X2 \SB1_2_3/INV_5  ( .I(\MC_ARK_ARC_1_1/buf_output[173] ), .ZN(
        \SB1_2_3/i1_5 ) );
  BUF_X4 \SB2_3_18/BUF_5  ( .I(\SB1_3_18/buf_output[5] ), .Z(\SB2_3_18/i0_3 )
         );
  CLKBUF_X4 \SB2_3_20/BUF_3  ( .I(\SB1_3_22/buf_output[3] ), .Z(
        \SB2_3_20/i0[10] ) );
  NAND3_X2 \SB1_1_22/Component_Function_5/N4  ( .A1(\SB1_1_22/i0[9] ), .A2(
        \SB1_1_22/i0[6] ), .A3(\SB1_1_22/i0_4 ), .ZN(
        \SB1_1_22/Component_Function_5/NAND4_in[3] ) );
  INV_X2 \SB2_2_27/INV_5  ( .I(\SB1_2_27/buf_output[5] ), .ZN(\SB2_2_27/i1_5 )
         );
  NAND3_X2 \SB1_1_4/Component_Function_2/N1  ( .A1(\SB1_1_4/i1_5 ), .A2(
        \SB1_1_4/i0[10] ), .A3(\SB1_1_4/i1[9] ), .ZN(
        \SB1_1_4/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB1_0_14/Component_Function_5/N2  ( .A1(\SB1_0_14/i0_0 ), .A2(
        \SB1_0_14/i0[6] ), .A3(\SB1_0_14/i0[10] ), .ZN(
        \SB1_0_14/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 \SB1_2_10/Component_Function_3/N2  ( .A1(\SB1_2_10/i0_0 ), .A2(
        \SB1_2_10/i0_3 ), .A3(\SB1_2_10/i0_4 ), .ZN(
        \SB1_2_10/Component_Function_3/NAND4_in[1] ) );
  BUF_X4 \SB2_0_24/BUF_4_0  ( .I(\SB2_0_24/buf_output[4] ), .Z(\RI5[0][52] )
         );
  NAND3_X2 \SB1_3_10/Component_Function_2/N2  ( .A1(n1388), .A2(
        \SB1_3_10/i0[10] ), .A3(\SB1_3_10/i0[6] ), .ZN(
        \SB1_3_10/Component_Function_2/NAND4_in[1] ) );
  NAND4_X2 \SB2_0_18/Component_Function_4/N5  ( .A1(
        \SB2_0_18/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_18/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_18/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_0_18/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_0_18/buf_output[4] ) );
  NAND3_X2 \SB3_7/Component_Function_4/N4  ( .A1(\SB3_7/i1[9] ), .A2(n4766), 
        .A3(\SB3_7/i0_4 ), .ZN(\SB3_7/Component_Function_4/NAND4_in[3] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_179  ( .I(\SB2_3_2/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[179] ) );
  NAND4_X2 \SB2_0_7/Component_Function_3/N5  ( .A1(
        \SB2_0_7/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_7/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_0_7/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_0_7/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_0_7/buf_output[3] ) );
  INV_X2 \SB1_0_7/INV_2  ( .I(n319), .ZN(\SB1_0_7/i1[9] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_123  ( .I(\SB2_1_13/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[123] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_47  ( .I(\SB2_2_24/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[47] ) );
  BUF_X4 \SB1_1_13/BUF_2  ( .I(\MC_ARK_ARC_1_0/buf_output[110] ), .Z(
        \SB1_1_13/i0_0 ) );
  NAND3_X2 \SB2_3_23/Component_Function_3/N2  ( .A1(\SB2_3_23/i0_0 ), .A2(
        \SB2_3_23/i0_3 ), .A3(\SB2_3_23/i0_4 ), .ZN(
        \SB2_3_23/Component_Function_3/NAND4_in[1] ) );
  INV_X2 \SB2_2_5/INV_5  ( .I(\SB1_2_5/buf_output[5] ), .ZN(\SB2_2_5/i1_5 ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_36  ( .I(\SB2_2_30/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[36] ) );
  NAND3_X2 \SB1_3_10/Component_Function_2/N4  ( .A1(\SB1_3_10/i1_5 ), .A2(
        \SB1_3_10/i0_0 ), .A3(\SB1_3_10/i0_4 ), .ZN(
        \SB1_3_10/Component_Function_2/NAND4_in[3] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_59_1  ( .I(\MC_ARK_ARC_1_0/buf_output[59] ), .Z(
        \RI1[1][59] ) );
  INV_X2 \SB1_0_27/INV_2  ( .I(n259), .ZN(\SB1_0_27/i1[9] ) );
  BUF_X4 \SB2_0_23/BUF_4_0  ( .I(\SB2_0_23/buf_output[4] ), .Z(\RI5[0][58] )
         );
  BUF_X4 \SB2_2_29/BUF_2_0  ( .I(\SB2_2_29/buf_output[2] ), .Z(\RI5[2][32] )
         );
  NAND3_X2 \SB2_1_22/Component_Function_2/N2  ( .A1(\SB2_1_22/i0_3 ), .A2(
        \SB2_1_22/i0[10] ), .A3(\SB2_1_22/i0[6] ), .ZN(
        \SB2_1_22/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 \SB2_0_0/BUF_0_0  ( .I(\SB2_0_0/buf_output[0] ), .Z(\RI5[0][24] ) );
  INV_X2 \SB2_1_14/INV_3  ( .I(\SB1_1_16/buf_output[3] ), .ZN(\SB2_1_14/i0[8] ) );
  NAND3_X2 \SB2_1_13/Component_Function_4/N4  ( .A1(\SB2_1_13/i1[9] ), .A2(
        \SB2_1_13/i1_5 ), .A3(\SB2_1_13/i0_4 ), .ZN(
        \SB2_1_13/Component_Function_4/NAND4_in[3] ) );
  NAND2_X2 \SB1_2_9/Component_Function_5/N1  ( .A1(\SB1_2_9/i0_0 ), .A2(
        \SB1_2_9/i3[0] ), .ZN(\SB1_2_9/Component_Function_5/NAND4_in[0] ) );
  NAND4_X2 \SB2_0_24/Component_Function_4/N5  ( .A1(
        \SB2_0_24/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_24/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_24/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_0_24/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_0_24/buf_output[4] ) );
  NAND3_X2 \SB2_1_21/Component_Function_4/N4  ( .A1(\SB2_1_21/i1[9] ), .A2(
        \SB2_1_21/i1_5 ), .A3(\SB2_1_21/i0_4 ), .ZN(
        \SB2_1_21/Component_Function_4/NAND4_in[3] ) );
  NAND3_X2 \SB1_2_0/Component_Function_1/N3  ( .A1(\SB1_2_0/i1_5 ), .A2(
        \SB1_2_0/i0[6] ), .A3(\SB1_2_0/i0[9] ), .ZN(
        \SB1_2_0/Component_Function_1/NAND4_in[2] ) );
  INV_X2 \SB2_3_29/INV_1  ( .I(\SB1_3_1/buf_output[1] ), .ZN(\SB2_3_29/i1_7 )
         );
  NAND3_X2 \SB1_3_17/Component_Function_5/N2  ( .A1(\SB1_3_17/i0_0 ), .A2(
        \SB1_3_17/i0[6] ), .A3(\SB1_3_17/i0[10] ), .ZN(
        \SB1_3_17/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 \SB2_0_7/BUF_4_0  ( .I(\SB2_0_7/buf_output[4] ), .Z(\RI5[0][154] ) );
  INV_X2 \SB1_1_4/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[167] ), .ZN(
        \SB1_1_4/i1_5 ) );
  INV_X2 \SB2_2_14/INV_5  ( .I(\SB1_2_14/buf_output[5] ), .ZN(\SB2_2_14/i1_5 )
         );
  NAND2_X2 \SB1_0_14/Component_Function_5/N1  ( .A1(\SB1_0_14/i0_0 ), .A2(
        \SB1_0_14/i3[0] ), .ZN(\SB1_0_14/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_122  ( .I(\SB2_2_14/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[122] ) );
  BUF_X2 \SB4_3/BUF_1  ( .I(\SB3_7/buf_output[1] ), .Z(\SB4_3/i0[6] ) );
  INV_X2 \SB1_2_10/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[126] ), .ZN(
        \SB1_2_10/i3[0] ) );
  NAND4_X2 \SB2_3_13/Component_Function_1/N5  ( .A1(
        \SB2_3_13/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_13/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_13/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_13/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_3_13/buf_output[1] ) );
  BUF_X4 \SB2_3_17/BUF_5  ( .I(\SB1_3_17/buf_output[5] ), .Z(\SB2_3_17/i0_3 )
         );
  NAND3_X2 \SB2_1_26/Component_Function_5/N2  ( .A1(\SB2_1_26/i0_0 ), .A2(
        \SB2_1_26/i0[6] ), .A3(\SB2_1_26/i0[10] ), .ZN(
        \SB2_1_26/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 \SB2_3_26/BUF_3_0  ( .I(\SB2_3_26/buf_output[3] ), .Z(\RI5[3][45] )
         );
  NAND3_X2 \SB1_3_31/Component_Function_2/N2  ( .A1(\SB1_3_31/i0_3 ), .A2(
        \SB1_3_31/i0[10] ), .A3(\SB1_3_31/i0[6] ), .ZN(
        \SB1_3_31/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 \SB2_0_21/BUF_3_0  ( .I(\SB2_0_21/buf_output[3] ), .Z(\RI5[0][75] )
         );
  BUF_X4 \SB2_0_7/BUF_2_0  ( .I(\SB2_0_7/buf_output[2] ), .Z(\RI5[0][164] ) );
  NAND3_X2 \SB2_2_17/Component_Function_2/N4  ( .A1(\SB2_2_17/i1_5 ), .A2(
        \SB2_2_17/i0_0 ), .A3(\SB2_2_17/i0_4 ), .ZN(
        \SB2_2_17/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 \SB2_1_27/Component_Function_3/N4  ( .A1(\SB2_1_27/i1_5 ), .A2(
        \SB2_1_27/i0[8] ), .A3(\SB2_1_27/i3[0] ), .ZN(
        \SB2_1_27/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 \SB1_0_31/Component_Function_3/N4  ( .A1(\SB1_0_31/i1_5 ), .A2(
        \SB1_0_31/i0[8] ), .A3(\SB1_0_31/i3[0] ), .ZN(
        \SB1_0_31/Component_Function_3/NAND4_in[3] ) );
  NAND4_X2 \SB2_2_31/Component_Function_3/N5  ( .A1(
        \SB2_2_31/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_31/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_2_31/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_2_31/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_2_31/buf_output[3] ) );
  NAND3_X2 \SB1_2_0/Component_Function_3/N1  ( .A1(\SB1_2_0/i1[9] ), .A2(
        \SB1_2_0/i0_3 ), .A3(\SB1_2_0/i0[6] ), .ZN(
        \SB1_2_0/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 \SB2_3_18/Component_Function_2/N2  ( .A1(\SB2_3_18/i0_3 ), .A2(
        \SB2_3_18/i0[10] ), .A3(\SB2_3_18/i0[6] ), .ZN(
        \SB2_3_18/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 \SB1_0_5/BUF_2_0  ( .I(\SB1_0_5/buf_output[2] ), .Z(\RI3[0][176] ) );
  NAND4_X2 \SB2_0_31/Component_Function_0/N5  ( .A1(
        \SB2_0_31/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_31/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_31/Component_Function_0/NAND4_in[3] ), .A4(
        \SB2_0_31/Component_Function_0/NAND4_in[2] ), .ZN(
        \SB2_0_31/buf_output[0] ) );
  CLKBUF_X4 \SB2_1_29/BUF_1  ( .I(\SB1_1_1/buf_output[1] ), .Z(
        \SB2_1_29/i0[6] ) );
  NAND3_X1 \SB4_1/Component_Function_3/N4  ( .A1(\SB4_1/i1_5 ), .A2(
        \SB4_1/i0[8] ), .A3(\SB4_1/i3[0] ), .ZN(
        \SB4_1/Component_Function_3/NAND4_in[3] ) );
  INV_X2 \SB1_0_13/INV_3  ( .I(n377), .ZN(\SB1_0_13/i0[8] ) );
  BUF_X4 \SB2_0_8/BUF_4_0  ( .I(\SB2_0_8/buf_output[4] ), .Z(\RI5[0][148] ) );
  BUF_X4 \SB2_0_13/BUF_4_0  ( .I(\SB2_0_13/buf_output[4] ), .Z(\RI5[0][118] )
         );
  NAND4_X2 \SB2_0_13/Component_Function_4/N5  ( .A1(
        \SB2_0_13/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_13/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_13/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_0_13/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_0_13/buf_output[4] ) );
  NAND3_X2 \SB2_3_14/Component_Function_3/N4  ( .A1(\SB2_3_14/i1_5 ), .A2(
        \SB2_3_14/i0[8] ), .A3(\SB2_3_14/i3[0] ), .ZN(
        \SB2_3_14/Component_Function_3/NAND4_in[3] ) );
  BUF_X4 \SB2_0_1/BUF_1_0  ( .I(\SB2_0_1/buf_output[1] ), .Z(\RI5[0][13] ) );
  NAND3_X2 \SB2_3_3/Component_Function_3/N4  ( .A1(\SB2_3_3/i1_5 ), .A2(
        \SB2_3_3/i0[8] ), .A3(\SB2_3_3/i3[0] ), .ZN(
        \SB2_3_3/Component_Function_3/NAND4_in[3] ) );
  BUF_X4 \SB2_0_22/BUF_4_0  ( .I(\SB2_0_22/buf_output[4] ), .Z(\RI5[0][64] )
         );
  NAND4_X2 \SB2_0_22/Component_Function_4/N5  ( .A1(
        \SB2_0_22/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_22/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_22/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_0_22/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_0_22/buf_output[4] ) );
  BUF_X4 \SB2_2_29/BUF_5_0  ( .I(\SB2_2_29/buf_output[5] ), .Z(\RI5[2][17] )
         );
  NAND3_X2 \SB1_3_1/Component_Function_2/N3  ( .A1(\SB1_3_1/i0_3 ), .A2(
        \SB1_3_1/i0[8] ), .A3(\SB1_3_1/i0[9] ), .ZN(
        \SB1_3_1/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 \SB1_2_30/Component_Function_1/N3  ( .A1(\SB1_2_30/i1_5 ), .A2(
        \SB1_2_30/i0[6] ), .A3(\SB1_2_30/i0[9] ), .ZN(
        \SB1_2_30/Component_Function_1/NAND4_in[2] ) );
  BUF_X4 \SB2_2_9/BUF_4_0  ( .I(\SB2_2_9/buf_output[4] ), .Z(\RI5[2][142] ) );
  NAND3_X2 \SB2_0_1/Component_Function_2/N1  ( .A1(\SB2_0_1/i1_5 ), .A2(
        \SB2_0_1/i0[10] ), .A3(\SB2_0_1/i1[9] ), .ZN(
        \SB2_0_1/Component_Function_2/NAND4_in[0] ) );
  CLKBUF_X4 \SB2_0_0/BUF_3  ( .I(\SB1_0_2/buf_output[3] ), .Z(\SB2_0_0/i0[10] ) );
  INV_X2 \SB1_0_6/INV_2  ( .I(n322), .ZN(\SB1_0_6/i1[9] ) );
  NAND4_X2 \SB2_0_12/Component_Function_0/N5  ( .A1(
        \SB2_0_12/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_12/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_12/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_12/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB2_0_12/buf_output[0] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_185  ( .I(\SB2_2_1/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[185] ) );
  CLKBUF_X4 \SB2_3_1/BUF_2  ( .I(\SB1_3_4/buf_output[2] ), .Z(\SB2_3_1/i0_0 )
         );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_117  ( .I(\SB2_2_14/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[117] ) );
  BUF_X4 \SB2_0_15/BUF_4_0  ( .I(\SB2_0_15/buf_output[4] ), .Z(\RI5[0][106] )
         );
  BUF_X4 \SB2_0_3/BUF_0_0  ( .I(\SB2_0_3/buf_output[0] ), .Z(\RI5[0][6] ) );
  NAND4_X2 \SB2_0_3/Component_Function_0/N5  ( .A1(
        \SB2_0_3/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_3/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_3/Component_Function_0/NAND4_in[3] ), .A4(
        \SB2_0_3/Component_Function_0/NAND4_in[2] ), .ZN(
        \SB2_0_3/buf_output[0] ) );
  NAND4_X2 \SB1_0_27/Component_Function_4/N5  ( .A1(
        \SB1_0_27/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_27/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_27/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_27/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_0_27/buf_output[4] ) );
  NAND4_X2 \SB2_1_18/Component_Function_1/N5  ( .A1(
        \SB2_1_18/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_18/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_18/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_18/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_1_18/buf_output[1] ) );
  NAND3_X2 \SB2_1_18/Component_Function_1/N4  ( .A1(\SB2_1_18/i1_7 ), .A2(
        \SB2_1_18/i0[8] ), .A3(\SB2_1_18/i0_4 ), .ZN(
        \SB2_1_18/Component_Function_1/NAND4_in[3] ) );
  BUF_X4 \SB1_2_21/BUF_2  ( .I(\MC_ARK_ARC_1_1/buf_output[62] ), .Z(
        \SB1_2_21/i0_0 ) );
  BUF_X4 \SB2_3_8/BUF_4_0  ( .I(\SB2_3_8/buf_output[4] ), .Z(\RI5[3][148] ) );
  NAND4_X2 \SB2_1_24/Component_Function_2/N5  ( .A1(
        \SB2_1_24/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_24/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_1_24/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_1_24/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_1_24/buf_output[2] ) );
  NAND4_X2 \SB2_1_4/Component_Function_4/N5  ( .A1(
        \SB2_1_4/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_4/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_4/Component_Function_4/NAND4_in[3] ), .A4(
        \SB2_1_4/Component_Function_4/NAND4_in[2] ), .ZN(
        \SB2_1_4/buf_output[4] ) );
  NAND3_X2 \SB2_1_20/Component_Function_3/N4  ( .A1(\SB2_1_20/i1_5 ), .A2(
        \SB2_1_20/i0[8] ), .A3(\SB2_1_20/i3[0] ), .ZN(
        \SB2_1_20/Component_Function_3/NAND4_in[3] ) );
  NAND4_X2 \SB2_0_4/Component_Function_2/N5  ( .A1(
        \SB2_0_4/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_4/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_0_4/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_0_4/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB2_0_4/buf_output[2] ) );
  NAND3_X2 \SB2_0_4/Component_Function_2/N3  ( .A1(\SB2_0_4/i0_3 ), .A2(
        \SB2_0_4/i0[8] ), .A3(\SB2_0_4/i0[9] ), .ZN(
        \SB2_0_4/Component_Function_2/NAND4_in[2] ) );
  NAND2_X2 \SB1_0_16/Component_Function_5/N1  ( .A1(\SB1_0_16/i0_0 ), .A2(
        \SB1_0_16/i3[0] ), .ZN(\SB1_0_16/Component_Function_5/NAND4_in[0] ) );
  INV_X2 \SB1_0_23/INV_3  ( .I(n357), .ZN(\SB1_0_23/i0[8] ) );
  BUF_X4 \SB2_0_15/BUF_0_0  ( .I(\SB2_0_15/buf_output[0] ), .Z(\RI5[0][126] )
         );
  CLKBUF_X4 \SB2_3_18/BUF_2  ( .I(\SB1_3_21/buf_output[2] ), .Z(
        \SB2_3_18/i0_0 ) );
  NAND4_X2 \SB1_0_4/Component_Function_1/N5  ( .A1(
        \SB1_0_4/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_4/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_4/Component_Function_1/NAND4_in[3] ), .A4(
        \SB1_0_4/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB1_0_4/buf_output[1] ) );
  NAND3_X2 \SB2_1_31/Component_Function_3/N4  ( .A1(n5510), .A2(
        \SB2_1_31/i0[8] ), .A3(\SB2_1_31/i3[0] ), .ZN(
        \SB2_1_31/Component_Function_3/NAND4_in[3] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_92  ( .I(\SB2_0_19/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[92] ) );
  NAND3_X2 \SB1_2_19/Component_Function_3/N2  ( .A1(\SB1_2_19/i0_0 ), .A2(
        \SB1_2_19/i0_3 ), .A3(\SB1_2_19/i0_4 ), .ZN(
        \SB1_2_19/Component_Function_3/NAND4_in[1] ) );
  BUF_X4 \SB2_0_4/BUF_2_0  ( .I(\SB2_0_4/buf_output[2] ), .Z(\RI5[0][182] ) );
  BUF_X4 \SB1_0_27/BUF_0_0  ( .I(\SB1_0_27/buf_output[0] ), .Z(\RI3[0][54] )
         );
  NAND4_X2 \SB2_2_18/Component_Function_3/N5  ( .A1(
        \SB2_2_18/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_18/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_2_18/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_2_18/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_2_18/buf_output[3] ) );
  BUF_X4 \SB2_0_22/BUF_0_0  ( .I(\SB2_0_22/buf_output[0] ), .Z(\RI5[0][84] )
         );
  INV_X4 \SB2_1_18/INV_1  ( .I(\SB1_1_22/buf_output[1] ), .ZN(\SB2_1_18/i1_7 )
         );
  NAND3_X2 \SB2_0_22/Component_Function_3/N3  ( .A1(\SB2_0_22/i1[9] ), .A2(
        \SB2_0_22/i1_7 ), .A3(\SB2_0_22/i0[10] ), .ZN(
        \SB2_0_22/Component_Function_3/NAND4_in[2] ) );
  CLKBUF_X4 \SB2_3_14/BUF_2  ( .I(\SB1_3_17/buf_output[2] ), .Z(
        \SB2_3_14/i0_0 ) );
  NAND3_X2 \SB2_0_20/Component_Function_3/N4  ( .A1(\SB2_0_20/i1_5 ), .A2(
        \SB2_0_20/i0[8] ), .A3(\SB2_0_20/i3[0] ), .ZN(
        \SB2_0_20/Component_Function_3/NAND4_in[3] ) );
  BUF_X4 \SB2_1_24/BUF_2_0  ( .I(\SB2_1_24/buf_output[2] ), .Z(\RI5[1][62] )
         );
  NAND3_X2 \SB2_1_24/Component_Function_2/N1  ( .A1(\SB2_1_24/i1_5 ), .A2(
        \SB2_1_24/i0[10] ), .A3(\SB2_1_24/i1[9] ), .ZN(
        \SB2_1_24/Component_Function_2/NAND4_in[0] ) );
  NAND2_X2 \SB2_2_14/Component_Function_5/N1  ( .A1(\SB2_2_14/i0_0 ), .A2(
        \SB2_2_14/i3[0] ), .ZN(\SB2_2_14/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 \SB1_0_20/BUF_5  ( .I(n416), .Z(\SB1_0_20/i0_3 ) );
  NAND2_X2 \SB1_2_17/Component_Function_5/N1  ( .A1(\SB1_2_17/i0_0 ), .A2(
        \SB1_2_17/i3[0] ), .ZN(\SB1_2_17/Component_Function_5/NAND4_in[0] ) );
  NAND4_X2 \SB2_0_7/Component_Function_1/N5  ( .A1(
        \SB2_0_7/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_7/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_7/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_0_7/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_0_7/buf_output[1] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_92  ( .I(\SB2_2_19/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[92] ) );
  NAND4_X2 \SB2_0_8/Component_Function_1/N5  ( .A1(
        \SB2_0_8/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_8/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_8/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_8/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_0_8/buf_output[1] ) );
  BUF_X4 \SB2_0_12/BUF_1_0  ( .I(\SB2_0_12/buf_output[1] ), .Z(\RI5[0][139] )
         );
  NAND4_X2 \SB1_0_31/Component_Function_1/N5  ( .A1(
        \SB1_0_31/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_31/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_31/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_31/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_0_31/buf_output[1] ) );
  BUF_X4 \SB2_0_4/BUF_1_0  ( .I(\SB2_0_4/buf_output[1] ), .Z(\RI5[0][187] ) );
  INV_X2 \SB1_0_5/INV_2  ( .I(n3675), .ZN(\SB1_0_5/i1[9] ) );
  BUF_X4 \SB2_0_10/BUF_2_0  ( .I(\SB2_0_10/buf_output[2] ), .Z(\RI5[0][146] )
         );
  NAND3_X2 \SB2_0_15/Component_Function_2/N3  ( .A1(\SB2_0_15/i0_3 ), .A2(
        \SB2_0_15/i0[8] ), .A3(\SB2_0_15/i0[9] ), .ZN(
        \SB2_0_15/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 \SB2_3_5/Component_Function_3/N5  ( .A1(
        \SB2_3_5/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_5/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_5/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_5/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_3_5/buf_output[3] ) );
  NAND3_X2 \SB2_2_18/Component_Function_3/N4  ( .A1(n4769), .A2(
        \SB2_2_18/i0[8] ), .A3(\SB2_2_18/i3[0] ), .ZN(
        \SB2_2_18/Component_Function_3/NAND4_in[3] ) );
  BUF_X4 \SB2_3_12/BUF_2_0  ( .I(\SB2_3_12/buf_output[2] ), .Z(\RI5[3][134] )
         );
  NAND2_X2 \SB1_0_7/Component_Function_5/N1  ( .A1(\SB1_0_7/i0_0 ), .A2(
        \SB1_0_7/i3[0] ), .ZN(\SB1_0_7/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 \SB1_0_1/BUF_5  ( .I(n435), .Z(\SB1_0_1/i0_3 ) );
  NAND3_X2 \SB1_0_24/Component_Function_5/N3  ( .A1(\SB1_0_24/i1[9] ), .A2(
        \SB1_0_24/i0_4 ), .A3(\SB1_0_24/i0_3 ), .ZN(
        \SB1_0_24/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 \SB2_2_29/Component_Function_1/N5  ( .A1(
        \SB2_2_29/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_29/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_29/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_2_29/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_2_29/buf_output[1] ) );
  NAND2_X2 \SB2_1_20/Component_Function_5/N1  ( .A1(\SB2_1_20/i0_0 ), .A2(
        \SB2_1_20/i3[0] ), .ZN(\SB2_1_20/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 \SB2_0_9/BUF_4_0  ( .I(\SB2_0_9/buf_output[4] ), .Z(\RI5[0][142] ) );
  NAND3_X2 \SB2_1_29/Component_Function_0/N4  ( .A1(\SB2_1_29/i0[7] ), .A2(
        \SB2_1_29/i0_3 ), .A3(\SB2_1_29/i0_0 ), .ZN(
        \SB2_1_29/Component_Function_0/NAND4_in[3] ) );
  NAND3_X2 \SB2_2_17/Component_Function_2/N2  ( .A1(\SB2_2_17/i0_3 ), .A2(
        \SB2_2_17/i0[10] ), .A3(\SB2_2_17/i0[6] ), .ZN(
        \SB2_2_17/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 \SB2_3_31/Component_Function_2/N2  ( .A1(\SB2_3_31/i0_3 ), .A2(
        \SB2_3_31/i0[10] ), .A3(\SB2_3_31/i0[6] ), .ZN(
        \SB2_3_31/Component_Function_2/NAND4_in[1] ) );
  NAND2_X2 \SB1_2_22/Component_Function_1/N1  ( .A1(\SB1_2_22/i0_3 ), .A2(
        \SB1_2_22/i1[9] ), .ZN(\SB1_2_22/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 \SB1_2_13/Component_Function_3/N2  ( .A1(\SB1_2_13/i0_0 ), .A2(
        \SB1_2_13/i0_3 ), .A3(\SB1_2_13/i0_4 ), .ZN(
        \SB1_2_13/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 \SB2_2_14/Component_Function_3/N3  ( .A1(\SB2_2_14/i1[9] ), .A2(
        \SB2_2_14/i1_7 ), .A3(\SB2_2_14/i0[10] ), .ZN(
        \SB2_2_14/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 \SB2_1_10/Component_Function_2/N3  ( .A1(\SB2_1_10/i0_3 ), .A2(
        \SB2_1_10/i0[8] ), .A3(\SB2_1_10/i0[9] ), .ZN(
        \SB2_1_10/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 \SB2_0_27/Component_Function_2/N4  ( .A1(\SB2_0_27/i1_5 ), .A2(
        \SB2_0_27/i0_0 ), .A3(\SB2_0_27/i0_4 ), .ZN(
        \SB2_0_27/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 \SB2_2_14/Component_Function_2/N1  ( .A1(\SB2_2_14/i1_5 ), .A2(
        \SB2_2_14/i0[10] ), .A3(\SB2_2_14/i1[9] ), .ZN(
        \SB2_2_14/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 \SB2_3_11/BUF_5_0  ( .I(\SB2_3_11/buf_output[5] ), .Z(\RI5[3][125] )
         );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_132  ( .I(\SB2_0_14/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[132] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_150  ( .I(\SB2_0_11/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[150] ) );
  INV_X2 \SB1_0_12/INV_3  ( .I(n379), .ZN(\SB1_0_12/i0[8] ) );
  BUF_X4 \SB2_2_11/BUF_3_0  ( .I(\SB2_2_11/buf_output[3] ), .Z(\RI5[2][135] )
         );
  NAND3_X2 \SB2_3_10/Component_Function_2/N2  ( .A1(\SB2_3_10/i0_3 ), .A2(
        \SB2_3_10/i0[10] ), .A3(\SB2_3_10/i0[6] ), .ZN(
        \SB2_3_10/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 \SB2_0_31/BUF_0_0  ( .I(\SB2_0_31/buf_output[0] ), .Z(\RI5[0][30] )
         );
  NAND4_X2 \SB2_1_11/Component_Function_3/N5  ( .A1(
        \SB2_1_11/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_11/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_11/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_1_11/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_1_11/buf_output[3] ) );
  INV_X2 \SB1_0_0/INV_3  ( .I(n403), .ZN(\SB1_0_0/i0[8] ) );
  NAND4_X2 \SB2_0_31/Component_Function_1/N5  ( .A1(
        \SB2_0_31/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_31/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_31/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_0_31/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_0_31/buf_output[1] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_31  ( .I(\SB2_1_30/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[31] ) );
  BUF_X4 \SB1_0_24/BUF_5  ( .I(n412), .Z(\SB1_0_24/i0_3 ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_154  ( .I(\SB2_3_7/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[154] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_79  ( .I(\SB2_0_22/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[79] ) );
  NAND4_X2 \SB2_0_22/Component_Function_1/N5  ( .A1(
        \SB2_0_22/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_22/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_22/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_0_22/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_0_22/buf_output[1] ) );
  CLKBUF_X4 \SB1_0_2/BUF_4  ( .I(n400), .Z(\SB1_0_2/i0_4 ) );
  NAND2_X2 \SB1_2_4/Component_Function_5/N1  ( .A1(\SB1_2_4/i0_0 ), .A2(
        \SB1_2_4/i3[0] ), .ZN(\SB1_2_4/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_22  ( .I(\SB2_3_29/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[22] ) );
  INV_X2 \SB3_1/INV_5  ( .I(\MC_ARK_ARC_1_3/buf_output[185] ), .ZN(
        \SB3_1/i1_5 ) );
  NAND3_X2 \SB2_2_18/Component_Function_2/N3  ( .A1(\SB2_2_18/i0_3 ), .A2(
        \SB2_2_18/i0[8] ), .A3(\SB2_2_18/i0[9] ), .ZN(
        \SB2_2_18/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 \SB2_0_8/BUF_2_0  ( .I(\SB2_0_8/buf_output[2] ), .Z(\RI5[0][158] ) );
  BUF_X4 \SB1_0_9/BUF_4_0  ( .I(\SB1_0_9/buf_output[4] ), .Z(\RI3[0][142] ) );
  NAND3_X2 \SB2_2_5/Component_Function_2/N2  ( .A1(\SB2_2_5/i0_3 ), .A2(
        \SB2_2_5/i0[10] ), .A3(\SB2_2_5/i0[6] ), .ZN(
        \SB2_2_5/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 \SB2_1_1/Component_Function_3/N2  ( .A1(\SB2_1_1/i0_0 ), .A2(
        \SB2_1_1/i0_3 ), .A3(\SB2_1_1/i0_4 ), .ZN(
        \SB2_1_1/Component_Function_3/NAND4_in[1] ) );
  BUF_X2 \SB1_1_2/BUF_3  ( .I(\MC_ARK_ARC_1_0/buf_output[177] ), .Z(
        \SB1_1_2/i0[10] ) );
  BUF_X2 \SB1_2_31/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[1] ), .Z(
        \SB1_2_31/i0[6] ) );
  NAND3_X2 \SB2_2_19/Component_Function_2/N3  ( .A1(\SB2_2_19/i0_3 ), .A2(
        \SB2_2_19/i0[8] ), .A3(\SB2_2_19/i0[9] ), .ZN(
        \SB2_2_19/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 \SB2_0_27/Component_Function_1/N5  ( .A1(
        \SB2_0_27/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_27/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_27/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_27/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_0_27/buf_output[1] ) );
  NAND3_X2 \SB1_2_24/Component_Function_2/N4  ( .A1(\SB1_2_24/i1_5 ), .A2(
        \SB1_2_24/i0_0 ), .A3(\SB1_2_24/i0_4 ), .ZN(
        \SB1_2_24/Component_Function_2/NAND4_in[3] ) );
  BUF_X4 \SB2_0_11/BUF_1_0  ( .I(\SB2_0_11/buf_output[1] ), .Z(\RI5[0][145] )
         );
  NAND4_X2 \SB2_3_28/Component_Function_3/N5  ( .A1(
        \SB2_3_28/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_28/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_28/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_28/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_3_28/buf_output[3] ) );
  NAND3_X2 \SB2_1_14/Component_Function_2/N3  ( .A1(\SB2_1_14/i0_3 ), .A2(
        \SB2_1_14/i0[8] ), .A3(\SB2_1_14/i0[9] ), .ZN(
        \SB2_1_14/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 \SB1_3_20/Component_Function_2/N3  ( .A1(\SB1_3_20/i0_3 ), .A2(
        \SB1_3_20/i0[8] ), .A3(\SB1_3_20/i0[9] ), .ZN(
        \SB1_3_20/Component_Function_2/NAND4_in[2] ) );
  CLKBUF_X4 \SB2_1_12/BUF_1  ( .I(\SB1_1_16/buf_output[1] ), .Z(
        \SB2_1_12/i0[6] ) );
  NAND4_X2 \SB2_3_13/Component_Function_3/N5  ( .A1(
        \SB2_3_13/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_13/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_13/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_13/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_3_13/buf_output[3] ) );
  BUF_X2 U77 ( .I(Key[183]), .Z(n225) );
  INV_X2 \SB2_2_23/INV_1  ( .I(\SB1_2_27/buf_output[1] ), .ZN(\SB2_2_23/i1_7 )
         );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_139  ( .I(\SB2_1_12/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[139] ) );
  NAND4_X2 \SB1_0_10/Component_Function_1/N5  ( .A1(
        \SB1_0_10/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_0_10/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_10/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_10/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_0_10/buf_output[1] ) );
  CLKBUF_X4 \SB2_2_27/BUF_0  ( .I(\SB1_2_0/buf_output[0] ), .Z(
        \SB2_2_27/i0[9] ) );
  NAND3_X2 \SB1_2_0/Component_Function_1/N4  ( .A1(\SB1_2_0/i1_7 ), .A2(
        \SB1_2_0/i0[8] ), .A3(\SB1_2_0/i0_4 ), .ZN(
        \SB1_2_0/Component_Function_1/NAND4_in[3] ) );
  BUF_X2 U95 ( .I(Key[74]), .Z(n146) );
  NAND3_X2 \SB2_1_12/Component_Function_2/N2  ( .A1(\SB2_1_12/i0_3 ), .A2(
        \SB2_1_12/i0[10] ), .A3(\SB2_1_12/i0[6] ), .ZN(
        \SB2_1_12/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 \SB2_1_10/Component_Function_2/N2  ( .A1(\SB2_1_10/i0_3 ), .A2(
        \SB2_1_10/i0[10] ), .A3(\SB2_1_10/i0[6] ), .ZN(
        \SB2_1_10/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 \SB2_3_24/BUF_2_0  ( .I(\SB2_3_24/buf_output[2] ), .Z(\RI5[3][62] )
         );
  INV_X2 \SB1_0_21/INV_3  ( .I(n361), .ZN(\SB1_0_21/i0[8] ) );
  NAND3_X2 \SB2_2_21/Component_Function_2/N1  ( .A1(\SB2_2_21/i1_5 ), .A2(
        \SB2_2_21/i0[10] ), .A3(\SB2_2_21/i1[9] ), .ZN(
        \SB2_2_21/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB2_0_3/Component_Function_2/N3  ( .A1(\SB2_0_3/i0_3 ), .A2(
        \SB2_0_3/i0[8] ), .A3(\SB2_0_3/i0[9] ), .ZN(
        \SB2_0_3/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 \SB2_1_2/Component_Function_2/N2  ( .A1(\SB2_1_2/i0_3 ), .A2(
        \SB2_1_2/i0[10] ), .A3(\SB2_1_2/i0[6] ), .ZN(
        \SB2_1_2/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 \SB2_3_12/Component_Function_3/N1  ( .A1(\SB2_3_12/i1[9] ), .A2(
        \SB2_3_12/i0_3 ), .A3(\SB2_3_12/i0[6] ), .ZN(
        \SB2_3_12/Component_Function_3/NAND4_in[0] ) );
  NAND2_X2 \SB2_1_12/Component_Function_5/N1  ( .A1(\SB2_1_12/i0_0 ), .A2(
        \SB2_1_12/i3[0] ), .ZN(\SB2_1_12/Component_Function_5/NAND4_in[0] ) );
  BUF_X2 U92 ( .I(Key[88]), .Z(n163) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_129  ( .I(\SB2_2_12/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[129] ) );
  NAND3_X2 \SB2_2_9/Component_Function_2/N2  ( .A1(\SB2_2_9/i0_3 ), .A2(
        \SB2_2_9/i0[10] ), .A3(\SB2_2_9/i0[6] ), .ZN(
        \SB2_2_9/Component_Function_2/NAND4_in[1] ) );
  BUF_X2 U96 ( .I(Key[132]), .Z(n105) );
  CLKBUF_X2 U33 ( .I(Key[102]), .Z(n28) );
  BUF_X2 U59 ( .I(Key[180]), .Z(n67) );
  CLKBUF_X4 \SB1_0_14/BUF_4  ( .I(n376), .Z(\SB1_0_14/i0_4 ) );
  CLKBUF_X4 \SB1_0_19/BUF_4  ( .I(n366), .Z(\SB1_0_19/i0_4 ) );
  CLKBUF_X4 \SB1_0_14/BUF_3  ( .I(n375), .Z(\SB1_0_14/i0[10] ) );
  INV_X1 U3 ( .I(n7), .ZN(n564) );
  CLKBUF_X4 \SB1_0_21/BUF_3  ( .I(n361), .Z(\SB1_0_21/i0[10] ) );
  CLKBUF_X4 \SB1_0_12/BUF_2  ( .I(n304), .Z(\SB1_0_12/i0_0 ) );
  INV_X1 U10 ( .I(n10), .ZN(n459) );
  CLKBUF_X4 \SB1_0_23/BUF_4  ( .I(n358), .Z(\SB1_0_23/i0_4 ) );
  CLKBUF_X4 \SB1_0_0/BUF_3  ( .I(n403), .Z(\SB1_0_0/i0[10] ) );
  CLKBUF_X4 \SB1_0_3/BUF_1  ( .I(n330), .Z(\SB1_0_3/i0[6] ) );
  CLKBUF_X4 \SB1_0_0/BUF_2  ( .I(n340), .Z(\SB1_0_0/i0_0 ) );
  CLKBUF_X4 \SB1_0_0/BUF_4  ( .I(n404), .Z(\SB1_0_0/i0_4 ) );
  INV_X1 U5 ( .I(n75), .ZN(n465) );
  INV_X1 U11 ( .I(n104), .ZN(n461) );
  CLKBUF_X4 \SB1_0_7/BUF_3  ( .I(n389), .Z(\SB1_0_7/i0[10] ) );
  BUF_X1 \MC_ARK_ARC_1_2/BUF_54_0  ( .I(n225), .Z(
        \MC_ARK_ARC_1_2/buf_keyinput[54] ) );
  CLKBUF_X4 \SB2_0_14/BUF_1  ( .I(\RI3[0][103] ), .Z(\SB2_0_14/i0[6] ) );
  CLKBUF_X4 \SB2_0_16/BUF_2  ( .I(\RI3[0][92] ), .Z(\SB2_0_16/i0_0 ) );
  CLKBUF_X4 \SB1_0_26/BUF_4_0  ( .I(\SB1_0_26/buf_output[4] ), .Z(\RI3[0][40] ) );
  CLKBUF_X4 \SB2_0_10/BUF_3  ( .I(\RI3[0][129] ), .Z(\SB2_0_10/i0[10] ) );
  BUF_X2 \SB1_0_10/BUF_0_0  ( .I(\SB1_0_10/buf_output[0] ), .Z(\RI3[0][156] )
         );
  CLKBUF_X4 \SB2_0_18/BUF_0  ( .I(\SB1_0_23/buf_output[0] ), .Z(
        \SB2_0_18/i0[9] ) );
  CLKBUF_X4 \SB2_0_20/BUF_3  ( .I(\RI3[0][69] ), .Z(\SB2_0_20/i0[10] ) );
  CLKBUF_X4 \SB2_0_12/BUF_4  ( .I(\RI3[0][118] ), .Z(\SB2_0_12/i0_4 ) );
  CLKBUF_X4 \MC_ARK_ARC_1_0/BUF_12  ( .I(\SB2_0_2/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[12] ) );
  CLKBUF_X4 \SB1_1_19/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[73] ), .Z(
        \SB1_1_19/i0[6] ) );
  BUF_X2 \SB1_1_18/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[78] ), .Z(
        \SB1_1_18/i0[9] ) );
  CLKBUF_X4 \SB1_1_18/BUF_2  ( .I(\MC_ARK_ARC_1_0/buf_output[80] ), .Z(
        \SB1_1_18/i0_0 ) );
  CLKBUF_X4 \SB1_1_6/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[154] ), .Z(
        \SB1_1_6/i0_4 ) );
  CLKBUF_X4 \SB1_1_12/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[114] ), .Z(
        \SB1_1_12/i0[9] ) );
  CLKBUF_X4 \SB1_1_18/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[82] ), .Z(
        \SB1_1_18/i0_4 ) );
  CLKBUF_X4 \SB1_1_12/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[118] ), .Z(
        \SB1_1_12/i0_4 ) );
  CLKBUF_X4 \SB1_1_21/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[64] ), .Z(
        \SB1_1_21/i0_4 ) );
  CLKBUF_X4 \SB2_1_10/BUF_3  ( .I(\SB1_1_12/buf_output[3] ), .Z(
        \SB2_1_10/i0[10] ) );
  CLKBUF_X4 \SB2_1_14/BUF_2  ( .I(\SB1_1_17/buf_output[2] ), .Z(
        \SB2_1_14/i0_0 ) );
  CLKBUF_X4 \SB2_1_30/BUF_1  ( .I(\SB1_1_2/buf_output[1] ), .Z(
        \SB2_1_30/i0[6] ) );
  CLKBUF_X4 \SB2_1_31/BUF_1  ( .I(\SB1_1_3/buf_output[1] ), .Z(
        \SB2_1_31/i0[6] ) );
  CLKBUF_X4 \SB2_1_16/BUF_2  ( .I(\SB1_1_19/buf_output[2] ), .Z(
        \SB2_1_16/i0_0 ) );
  CLKBUF_X4 \SB2_1_28/BUF_0  ( .I(\SB1_1_1/buf_output[0] ), .Z(
        \SB2_1_28/i0[9] ) );
  CLKBUF_X4 \SB2_1_18/BUF_2  ( .I(\SB1_1_21/buf_output[2] ), .Z(
        \SB2_1_18/i0_0 ) );
  CLKBUF_X4 \SB2_1_27/BUF_0  ( .I(\SB1_1_0/buf_output[0] ), .Z(
        \SB2_1_27/i0[9] ) );
  CLKBUF_X4 \SB1_2_7/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[145] ), .Z(
        \SB1_2_7/i0[6] ) );
  CLKBUF_X4 \SB1_2_21/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[64] ), .Z(
        \SB1_2_21/i0_4 ) );
  CLKBUF_X4 \SB1_2_19/BUF_3  ( .I(\MC_ARK_ARC_1_1/buf_output[75] ), .Z(
        \SB1_2_19/i0[10] ) );
  CLKBUF_X4 \SB1_2_15/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[96] ), .Z(
        \SB1_2_15/i0[9] ) );
  CLKBUF_X4 \SB1_2_15/BUF_2  ( .I(\MC_ARK_ARC_1_1/buf_output[98] ), .Z(
        \SB1_2_15/i0_0 ) );
  CLKBUF_X4 \SB1_2_20/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[66] ), .Z(
        \SB1_2_20/i0[9] ) );
  CLKBUF_X4 \SB1_2_18/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[82] ), .Z(
        \SB1_2_18/i0_4 ) );
  CLKBUF_X4 \SB1_2_30/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[6] ), .Z(
        \SB1_2_30/i0[9] ) );
  CLKBUF_X4 \SB2_2_17/BUF_1  ( .I(\SB1_2_21/buf_output[1] ), .Z(
        \SB2_2_17/i0[6] ) );
  CLKBUF_X4 \SB2_2_29/BUF_2  ( .I(\SB1_2_0/buf_output[2] ), .Z(\SB2_2_29/i0_0 ) );
  CLKBUF_X4 \SB2_2_24/BUF_4  ( .I(\SB1_2_25/buf_output[4] ), .Z(
        \SB2_2_24/i0_4 ) );
  CLKBUF_X4 \SB2_2_17/BUF_2  ( .I(\SB1_2_20/buf_output[2] ), .Z(
        \SB2_2_17/i0_0 ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_27  ( .I(\SB2_2_29/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[27] ) );
  CLKBUF_X4 \MC_ARK_ARC_1_2/BUF_156  ( .I(\SB2_2_10/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[156] ) );
  CLKBUF_X4 \SB1_3_6/BUF_3  ( .I(\MC_ARK_ARC_1_2/buf_output[153] ), .Z(
        \SB1_3_6/i0[10] ) );
  CLKBUF_X4 \SB1_3_3/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[172] ), .Z(
        \SB1_3_3/i0_4 ) );
  CLKBUF_X4 \SB1_3_1/BUF_3  ( .I(\MC_ARK_ARC_1_2/buf_output[183] ), .Z(
        \SB1_3_1/i0[10] ) );
  CLKBUF_X4 \SB1_3_0/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[190] ), .Z(
        \SB1_3_0/i0_4 ) );
  BUF_X2 \SB1_3_18/BUF_1  ( .I(\MC_ARK_ARC_1_2/buf_output[79] ), .Z(
        \SB1_3_18/i0[6] ) );
  CLKBUF_X4 \SB1_3_19/BUF_3  ( .I(\MC_ARK_ARC_1_2/buf_output[75] ), .Z(
        \SB1_3_19/i0[10] ) );
  CLKBUF_X4 \SB1_3_19/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[76] ), .Z(
        \SB1_3_19/i0_4 ) );
  CLKBUF_X4 \SB2_3_12/BUF_1  ( .I(\SB1_3_16/buf_output[1] ), .Z(
        \SB2_3_12/i0[6] ) );
  CLKBUF_X4 \SB2_3_17/BUF_1  ( .I(\SB1_3_21/buf_output[1] ), .Z(
        \SB2_3_17/i0[6] ) );
  CLKBUF_X4 \SB2_3_23/BUF_0  ( .I(\SB1_3_28/buf_output[0] ), .Z(
        \SB2_3_23/i0[9] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_101  ( .I(\SB2_3_15/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[101] ) );
  CLKBUF_X4 \SB3_7/BUF_2  ( .I(n3654), .Z(\SB3_7/i0_0 ) );
  CLKBUF_X4 \SB3_23/BUF_4  ( .I(\MC_ARK_ARC_1_3/buf_output[52] ), .Z(
        \SB3_23/i0_4 ) );
  CLKBUF_X4 \SB4_7/BUF_0  ( .I(\SB3_12/buf_output[0] ), .Z(\SB4_7/i0[9] ) );
  CLKBUF_X4 \SB4_3/BUF_4  ( .I(\SB3_4/buf_output[4] ), .Z(\SB4_3/i0_4 ) );
  CLKBUF_X4 \SB4_13/BUF_4  ( .I(\SB3_14/buf_output[4] ), .Z(\SB4_13/i0_4 ) );
  NAND3_X2 \SB2_1_4/Component_Function_3/N4  ( .A1(\SB2_1_4/i1_5 ), .A2(
        \SB2_1_4/i0[8] ), .A3(\SB2_1_4/i3[0] ), .ZN(
        \SB2_1_4/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_27/Component_Function_0/N2  ( .A1(\SB1_0_27/i0[8] ), .A2(
        \SB1_0_27/i0[7] ), .A3(\SB1_0_27/i0[6] ), .ZN(
        \SB1_0_27/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_28/Component_Function_4/N1  ( .A1(\SB1_0_28/i0[9] ), .A2(
        \SB1_0_28/i0_0 ), .A3(\SB1_0_28/i0[8] ), .ZN(
        \SB1_0_28/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_27/Component_Function_0/N3  ( .A1(\SB1_0_27/i0[10] ), .A2(
        \SB1_0_27/i0_4 ), .A3(\SB1_0_27/i0_3 ), .ZN(
        \SB1_0_27/Component_Function_0/NAND4_in[2] ) );
  BUF_X2 \SB1_0_12/BUF_0  ( .I(n302), .Z(\SB1_0_12/i0[9] ) );
  NAND3_X1 \SB1_0_31/Component_Function_1/N3  ( .A1(\SB1_0_31/i1_5 ), .A2(
        \SB1_0_31/i0[6] ), .A3(\SB1_0_31/i0[9] ), .ZN(
        \SB1_0_31/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_11/Component_Function_4/N2  ( .A1(\SB1_0_11/i3[0] ), .A2(
        \SB1_0_11/i0_0 ), .A3(\SB1_0_11/i1_7 ), .ZN(
        \SB1_0_11/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_14/Component_Function_4/N3  ( .A1(\SB1_0_14/i0[9] ), .A2(
        \SB1_0_14/i0[10] ), .A3(\SB1_0_14/i0_3 ), .ZN(
        \SB1_0_14/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_7/Component_Function_3/N3  ( .A1(\SB1_0_7/i1[9] ), .A2(
        \SB1_0_7/i1_7 ), .A3(\SB1_0_7/i0[10] ), .ZN(
        \SB1_0_7/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_7/Component_Function_3/N4  ( .A1(\SB1_0_7/i1_5 ), .A2(
        \SB1_0_7/i0[8] ), .A3(\SB1_0_7/i3[0] ), .ZN(
        \SB1_0_7/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_2/Component_Function_0/N4  ( .A1(\SB1_0_2/i0[7] ), .A2(
        \SB1_0_2/i0_3 ), .A3(\SB1_0_2/i0_0 ), .ZN(
        \SB1_0_2/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_27/Component_Function_5/N4  ( .A1(\SB1_0_27/i0[9] ), .A2(
        \SB1_0_27/i0[6] ), .A3(\SB1_0_27/i0_4 ), .ZN(
        \SB1_0_27/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB1_0_2/Component_Function_0/N1  ( .A1(\SB1_0_2/i0[10] ), .A2(
        \SB1_0_2/i0[9] ), .ZN(\SB1_0_2/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_22/Component_Function_4/N1  ( .A1(\SB1_0_22/i0[9] ), .A2(
        \SB1_0_22/i0_0 ), .A3(\SB1_0_22/i0[8] ), .ZN(
        \SB1_0_22/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_30/Component_Function_5/N2  ( .A1(\SB1_0_30/i0_0 ), .A2(
        \SB1_0_30/i0[6] ), .A3(\SB1_0_30/i0[10] ), .ZN(
        \SB1_0_30/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_15/Component_Function_0/N1  ( .A1(\SB1_0_15/i0[10] ), .A2(
        \SB1_0_15/i0[9] ), .ZN(\SB1_0_15/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_7/Component_Function_1/N4  ( .A1(\SB1_0_7/i1_7 ), .A2(
        \SB1_0_7/i0[8] ), .A3(n5496), .ZN(
        \SB1_0_7/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_19/Component_Function_3/N4  ( .A1(\SB1_0_19/i1_5 ), .A2(
        \SB1_0_19/i0[8] ), .A3(\SB1_0_19/i3[0] ), .ZN(
        \SB1_0_19/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_19/Component_Function_4/N2  ( .A1(\SB1_0_19/i3[0] ), .A2(
        \SB1_0_19/i0_0 ), .A3(\SB1_0_19/i1_7 ), .ZN(
        \SB1_0_19/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_13/Component_Function_2/N3  ( .A1(\SB1_0_13/i0_3 ), .A2(
        \SB1_0_13/i0[8] ), .A3(\SB1_0_13/i0[9] ), .ZN(
        \SB1_0_13/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_11/Component_Function_2/N2  ( .A1(\SB1_0_11/i0_3 ), .A2(
        \SB1_0_11/i0[10] ), .A3(\SB1_0_11/i0[6] ), .ZN(
        \SB1_0_11/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_13/Component_Function_2/N2  ( .A1(\SB1_0_13/i0_3 ), .A2(
        \SB1_0_13/i0[10] ), .A3(\SB1_0_13/i0[6] ), .ZN(
        \SB1_0_13/Component_Function_2/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_17/Component_Function_0/N1  ( .A1(\SB1_0_17/i0[10] ), .A2(
        \SB1_0_17/i0[9] ), .ZN(\SB1_0_17/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_20/Component_Function_0/N2  ( .A1(\SB1_0_20/i0[8] ), .A2(
        \SB1_0_20/i0[7] ), .A3(\SB1_0_20/i0[6] ), .ZN(
        \SB1_0_20/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_20/Component_Function_0/N4  ( .A1(\SB1_0_20/i0[7] ), .A2(
        \SB1_0_20/i0_3 ), .A3(\SB1_0_20/i0_0 ), .ZN(
        \SB1_0_20/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_29/Component_Function_1/N2  ( .A1(\SB1_0_29/i0_3 ), .A2(
        \SB1_0_29/i1_7 ), .A3(\SB1_0_29/i0[8] ), .ZN(
        \SB1_0_29/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_26/Component_Function_0/N4  ( .A1(\SB1_0_26/i0[7] ), .A2(
        \SB1_0_26/i0_3 ), .A3(\SB1_0_26/i0_0 ), .ZN(
        \SB1_0_26/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_21/Component_Function_5/N4  ( .A1(\SB1_0_21/i0[9] ), .A2(
        \SB1_0_21/i0[6] ), .A3(\SB1_0_21/i0_4 ), .ZN(
        \SB1_0_21/Component_Function_5/NAND4_in[3] ) );
  BUF_X2 \SB2_0_22/BUF_1  ( .I(\RI3[0][55] ), .Z(\SB2_0_22/i0[6] ) );
  INV_X1 \SB2_0_23/INV_0  ( .I(\RI3[0][48] ), .ZN(\SB2_0_23/i3[0] ) );
  NAND3_X1 \SB2_0_11/Component_Function_5/N4  ( .A1(\SB2_0_11/i0[9] ), .A2(
        \RI3[0][121] ), .A3(\SB2_0_11/i0_4 ), .ZN(
        \SB2_0_11/Component_Function_5/NAND4_in[3] ) );
  INV_X1 \SB2_0_22/INV_1  ( .I(\RI3[0][55] ), .ZN(\SB2_0_22/i1_7 ) );
  BUF_X2 \SB2_0_12/BUF_0  ( .I(\RI3[0][114] ), .Z(\SB2_0_12/i0[9] ) );
  BUF_X2 \SB2_0_26/BUF_0  ( .I(\RI3[0][30] ), .Z(\SB2_0_26/i0[9] ) );
  BUF_X2 \SB2_0_13/BUF_0  ( .I(\SB1_0_18/buf_output[0] ), .Z(\SB2_0_13/i0[9] )
         );
  BUF_X2 \SB2_0_19/BUF_0  ( .I(\RI3[0][72] ), .Z(\SB2_0_19/i0[9] ) );
  BUF_X2 \SB2_0_15/BUF_1  ( .I(\RI3[0][97] ), .Z(\SB2_0_15/i0[6] ) );
  BUF_X2 \SB2_0_21/BUF_0  ( .I(\SB1_0_26/buf_output[0] ), .Z(\SB2_0_21/i0[9] )
         );
  BUF_X2 \SB2_0_20/BUF_0  ( .I(\RI3[0][66] ), .Z(\SB2_0_20/i0[9] ) );
  INV_X1 \SB2_0_15/INV_1  ( .I(\RI3[0][97] ), .ZN(\SB2_0_15/i1_7 ) );
  INV_X1 \SB2_0_3/INV_4  ( .I(\SB1_0_4/buf_output[4] ), .ZN(\SB2_0_3/i0[7] )
         );
  NAND3_X1 \SB2_0_18/Component_Function_3/N2  ( .A1(\SB2_0_18/i0_0 ), .A2(
        \SB2_0_18/i0_3 ), .A3(\RI3[0][82] ), .ZN(
        \SB2_0_18/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_24/Component_Function_3/N4  ( .A1(\SB2_0_24/i1_5 ), .A2(
        \SB2_0_24/i0[8] ), .A3(\SB2_0_24/i3[0] ), .ZN(
        \SB2_0_24/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_16/Component_Function_1/N3  ( .A1(\SB2_0_16/i1_5 ), .A2(
        \SB2_0_16/i0[6] ), .A3(\SB1_0_21/buf_output[0] ), .ZN(
        \SB2_0_16/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_18/Component_Function_1/N3  ( .A1(\SB2_0_18/i1_5 ), .A2(
        \SB2_0_18/i0[6] ), .A3(\SB1_0_23/buf_output[0] ), .ZN(
        \SB2_0_18/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_24/Component_Function_4/N1  ( .A1(\SB2_0_24/i0[9] ), .A2(
        \SB2_0_24/i0_0 ), .A3(\SB2_0_24/i0[8] ), .ZN(
        \SB2_0_24/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_27/Component_Function_1/N2  ( .A1(\SB2_0_27/i0_3 ), .A2(
        \SB2_0_27/i1_7 ), .A3(\SB2_0_27/i0[8] ), .ZN(
        \SB2_0_27/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_26/Component_Function_1/N2  ( .A1(\SB2_0_26/i0_3 ), .A2(
        \SB2_0_26/i1_7 ), .A3(\SB2_0_26/i0[8] ), .ZN(
        \SB2_0_26/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_20/Component_Function_4/N1  ( .A1(\SB2_0_20/i0[9] ), .A2(
        \SB2_0_20/i0_0 ), .A3(\SB2_0_20/i0[8] ), .ZN(
        \SB2_0_20/Component_Function_4/NAND4_in[0] ) );
  INV_X1 \SB2_0_26/INV_4  ( .I(\SB1_0_27/buf_output[4] ), .ZN(\SB2_0_26/i0[7] ) );
  INV_X1 \SB2_0_14/INV_4  ( .I(\SB1_0_15/buf_output[4] ), .ZN(\SB2_0_14/i0[7] ) );
  NAND3_X1 \SB2_0_9/Component_Function_2/N4  ( .A1(n5518), .A2(\RI3[0][134] ), 
        .A3(\SB2_0_9/i0_4 ), .ZN(\SB2_0_9/Component_Function_2/NAND4_in[3] )
         );
  NAND3_X1 \SB2_0_22/Component_Function_4/N2  ( .A1(\SB2_0_22/i3[0] ), .A2(
        \SB2_0_22/i0_0 ), .A3(\SB2_0_22/i1_7 ), .ZN(
        \SB2_0_22/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_15/Component_Function_5/N4  ( .A1(\SB2_0_15/i0[9] ), .A2(
        \SB2_0_15/i0[6] ), .A3(\SB1_0_16/buf_output[4] ), .ZN(
        \SB2_0_15/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_10/Component_Function_0/N3  ( .A1(\SB2_0_10/i0[10] ), .A2(
        \SB2_0_10/i0_4 ), .A3(\SB2_0_10/i0_3 ), .ZN(
        \SB2_0_10/Component_Function_0/NAND4_in[2] ) );
  BUF_X2 \SB1_1_30/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[6] ), .Z(
        \SB1_1_30/i0[9] ) );
  NAND3_X1 \SB1_1_18/Component_Function_0/N4  ( .A1(\SB1_1_18/i0[7] ), .A2(
        \SB1_1_18/i0_3 ), .A3(\SB1_1_18/i0_0 ), .ZN(
        \SB1_1_18/Component_Function_0/NAND4_in[3] ) );
  BUF_X2 \SB1_1_16/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[90] ), .Z(
        \SB1_1_16/i0[9] ) );
  BUF_X2 \SB1_1_31/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[1] ), .Z(
        \SB1_1_31/i0[6] ) );
  BUF_X2 \SB1_1_11/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[120] ), .Z(
        \SB1_1_11/i0[9] ) );
  BUF_X2 \SB1_1_15/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[96] ), .Z(
        \SB1_1_15/i0[9] ) );
  BUF_X2 \SB1_1_6/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[150] ), .Z(
        \SB1_1_6/i0[9] ) );
  BUF_X2 \SB1_1_24/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[42] ), .Z(
        \SB1_1_24/i0[9] ) );
  INV_X2 \SB1_1_30/INV_5  ( .I(\RI1[1][11] ), .ZN(\SB1_1_30/i1_5 ) );
  NAND3_X1 \SB1_1_10/Component_Function_1/N2  ( .A1(\SB1_1_10/i0_3 ), .A2(
        \SB1_1_10/i1_7 ), .A3(\SB1_1_10/i0[8] ), .ZN(
        \SB1_1_10/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_12/Component_Function_4/N3  ( .A1(\SB1_1_12/i0[9] ), .A2(
        \SB1_1_12/i0[10] ), .A3(\SB1_1_12/i0_3 ), .ZN(
        \SB1_1_12/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_17/Component_Function_0/N4  ( .A1(\SB1_1_17/i0[7] ), .A2(
        \SB1_1_17/i0_3 ), .A3(\SB1_1_17/i0_0 ), .ZN(
        \SB1_1_17/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_24/Component_Function_4/N4  ( .A1(\SB1_1_24/i1[9] ), .A2(
        \SB1_1_24/i1_5 ), .A3(\SB1_1_24/i0_4 ), .ZN(
        \SB1_1_24/Component_Function_4/NAND4_in[3] ) );
  INV_X1 \SB1_1_16/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[90] ), .ZN(
        \SB1_1_16/i3[0] ) );
  NAND3_X1 \SB1_1_15/Component_Function_2/N3  ( .A1(\SB1_1_15/i0_3 ), .A2(
        \SB1_1_15/i0[8] ), .A3(\SB1_1_15/i0[9] ), .ZN(
        \SB1_1_15/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_0/Component_Function_2/N4  ( .A1(\SB1_1_0/i1_5 ), .A2(
        \SB1_1_0/i0_0 ), .A3(\SB1_1_0/i0_4 ), .ZN(
        \SB1_1_0/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_5/Component_Function_4/N4  ( .A1(\SB1_1_5/i1[9] ), .A2(
        \SB1_1_5/i1_5 ), .A3(\SB1_1_5/i0_4 ), .ZN(
        \SB1_1_5/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_31/Component_Function_3/N2  ( .A1(\SB1_1_31/i0_0 ), .A2(
        \SB1_1_31/i0_3 ), .A3(\SB1_1_31/i0_4 ), .ZN(
        \SB1_1_31/Component_Function_3/NAND4_in[1] ) );
  BUF_X2 \SB1_1_25/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[36] ), .Z(
        \SB1_1_25/i0[9] ) );
  NAND3_X1 \SB1_1_10/Component_Function_1/N4  ( .A1(\SB1_1_10/i1_7 ), .A2(
        \SB1_1_10/i0[8] ), .A3(\SB1_1_10/i0_4 ), .ZN(
        \SB1_1_10/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_1/Component_Function_3/N2  ( .A1(\SB1_1_1/i0_0 ), .A2(
        \SB1_1_1/i0_3 ), .A3(\SB1_1_1/i0_4 ), .ZN(
        \SB1_1_1/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_8/Component_Function_0/N2  ( .A1(\SB1_1_8/i0[8] ), .A2(
        \SB1_1_8/i0[7] ), .A3(\SB1_1_8/i0[6] ), .ZN(
        \SB1_1_8/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_4/Component_Function_0/N4  ( .A1(\SB1_1_4/i0[7] ), .A2(
        \SB1_1_4/i0_3 ), .A3(\SB1_1_4/i0_0 ), .ZN(
        \SB1_1_4/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_21/Component_Function_1/N3  ( .A1(\SB1_1_21/i1_5 ), .A2(
        \SB1_1_21/i0[6] ), .A3(\SB1_1_21/i0[9] ), .ZN(
        \SB1_1_21/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_24/Component_Function_2/N3  ( .A1(\SB1_1_24/i0_3 ), .A2(
        \SB1_1_24/i0[8] ), .A3(\SB1_1_24/i0[9] ), .ZN(
        \SB1_1_24/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_22/Component_Function_0/N2  ( .A1(\SB1_1_22/i0[8] ), .A2(
        \SB1_1_22/i0[7] ), .A3(\SB1_1_22/i0[6] ), .ZN(
        \SB1_1_22/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_3/Component_Function_2/N3  ( .A1(\SB1_1_3/i0_3 ), .A2(
        \SB1_1_3/i0[8] ), .A3(\SB1_1_3/i0[9] ), .ZN(
        \SB1_1_3/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_0/Component_Function_0/N2  ( .A1(\SB1_1_0/i0[8] ), .A2(
        \SB1_1_0/i0[7] ), .A3(\SB1_1_0/i0[6] ), .ZN(
        \SB1_1_0/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_12/Component_Function_0/N3  ( .A1(\SB1_1_12/i0[10] ), .A2(
        \SB1_1_12/i0_4 ), .A3(\SB1_1_12/i0_3 ), .ZN(
        \SB1_1_12/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_3/Component_Function_3/N2  ( .A1(\SB1_1_3/i0_0 ), .A2(
        \SB1_1_3/i0_3 ), .A3(\SB1_1_3/i0_4 ), .ZN(
        \SB1_1_3/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_7/Component_Function_3/N2  ( .A1(\SB1_1_7/i0_0 ), .A2(
        \SB1_1_7/i0_3 ), .A3(\SB1_1_7/i0_4 ), .ZN(
        \SB1_1_7/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_4/Component_Function_2/N3  ( .A1(\SB1_1_4/i0_3 ), .A2(
        \SB1_1_4/i0[8] ), .A3(\SB1_1_4/i0[9] ), .ZN(
        \SB1_1_4/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_1/Component_Function_3/N3  ( .A1(\SB1_1_1/i1[9] ), .A2(
        \SB1_1_1/i1_7 ), .A3(\SB1_1_1/i0[10] ), .ZN(
        \SB1_1_1/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_6/Component_Function_3/N2  ( .A1(\SB1_1_6/i0_0 ), .A2(
        \SB1_1_6/i0_3 ), .A3(\SB1_1_6/i0_4 ), .ZN(
        \SB1_1_6/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_24/Component_Function_3/N2  ( .A1(\SB1_1_24/i0_0 ), .A2(
        \SB1_1_24/i0_3 ), .A3(\SB1_1_24/i0_4 ), .ZN(
        \SB1_1_24/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_11/Component_Function_1/N2  ( .A1(\SB1_1_11/i0_3 ), .A2(
        \SB1_1_11/i1_7 ), .A3(\SB1_1_11/i0[8] ), .ZN(
        \SB1_1_11/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_30/Component_Function_5/N1  ( .A1(\SB2_1_30/i0_0 ), .A2(
        \SB2_1_30/i3[0] ), .ZN(\SB2_1_30/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_7/Component_Function_4/N3  ( .A1(\SB2_1_7/i0[9] ), .A2(
        \SB2_1_7/i0[10] ), .A3(\SB2_1_7/i0_3 ), .ZN(
        \SB2_1_7/Component_Function_4/NAND4_in[2] ) );
  NAND2_X1 \SB2_1_7/Component_Function_0/N1  ( .A1(\SB2_1_7/i0[10] ), .A2(
        \SB2_1_7/i0[9] ), .ZN(\SB2_1_7/Component_Function_0/NAND4_in[0] ) );
  INV_X1 \SB2_1_29/INV_1  ( .I(\SB1_1_1/buf_output[1] ), .ZN(\SB2_1_29/i1_7 )
         );
  INV_X1 \SB2_1_28/INV_1  ( .I(\SB1_1_0/buf_output[1] ), .ZN(\SB2_1_28/i1_7 )
         );
  NAND3_X1 \SB2_1_1/Component_Function_1/N2  ( .A1(\SB2_1_1/i0_3 ), .A2(
        \SB2_1_1/i1_7 ), .A3(\SB2_1_1/i0[8] ), .ZN(
        \SB2_1_1/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_23/Component_Function_4/N4  ( .A1(\SB2_1_23/i1[9] ), .A2(
        \SB2_1_23/i1_5 ), .A3(\SB2_1_23/i0_4 ), .ZN(
        \SB2_1_23/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_4/Component_Function_4/N4  ( .A1(n3660), .A2(\SB2_1_4/i1_5 ), 
        .A3(\SB1_1_5/buf_output[4] ), .ZN(
        \SB2_1_4/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_14/Component_Function_0/N2  ( .A1(\SB2_1_14/i0[8] ), .A2(
        \SB2_1_14/i0[7] ), .A3(\SB2_1_14/i0[6] ), .ZN(
        \SB2_1_14/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_21/Component_Function_4/N2  ( .A1(n4625), .A2(
        \SB2_1_21/i0_0 ), .A3(\SB2_1_21/i1_7 ), .ZN(
        \SB2_1_21/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_22/Component_Function_2/N1  ( .A1(\SB2_1_22/i1_5 ), .A2(
        \SB2_1_22/i0[10] ), .A3(\SB2_1_22/i1[9] ), .ZN(
        \SB2_1_22/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_1/Component_Function_0/N2  ( .A1(\SB2_1_1/i0[8] ), .A2(
        \SB2_1_1/i0[7] ), .A3(\SB2_1_1/i0[6] ), .ZN(
        \SB2_1_1/Component_Function_0/NAND4_in[1] ) );
  INV_X1 \SB1_2_2/INV_1  ( .I(\MC_ARK_ARC_1_1/buf_output[175] ), .ZN(
        \SB1_2_2/i1_7 ) );
  INV_X1 \SB1_2_14/INV_1  ( .I(\MC_ARK_ARC_1_1/buf_output[103] ), .ZN(
        \SB1_2_14/i1_7 ) );
  INV_X1 \SB1_2_11/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[120] ), .ZN(
        \SB1_2_11/i3[0] ) );
  BUF_X2 \SB1_2_27/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[24] ), .Z(
        \SB1_2_27/i0[9] ) );
  BUF_X2 \SB1_2_19/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[73] ), .Z(
        \SB1_2_19/i0[6] ) );
  INV_X4 \SB1_2_16/INV_5  ( .I(\RI1[2][95] ), .ZN(\SB1_2_16/i1_5 ) );
  INV_X1 \SB1_2_20/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[66] ), .ZN(
        \SB1_2_20/i3[0] ) );
  NAND3_X1 \SB1_2_5/Component_Function_0/N2  ( .A1(\SB1_2_5/i0[8] ), .A2(
        \SB1_2_5/i0[7] ), .A3(\SB1_2_5/i0[6] ), .ZN(
        \SB1_2_5/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_4/Component_Function_4/N4  ( .A1(\SB1_2_4/i1[9] ), .A2(
        \SB1_2_4/i1_5 ), .A3(\SB1_2_4/i0_4 ), .ZN(
        \SB1_2_4/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_17/Component_Function_0/N3  ( .A1(\SB1_2_17/i0[10] ), .A2(
        \SB1_2_17/i0_4 ), .A3(\SB1_2_17/i0_3 ), .ZN(
        \SB1_2_17/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_2_4/Component_Function_1/N1  ( .A1(\SB1_2_4/i0_3 ), .A2(
        \SB1_2_4/i1[9] ), .ZN(\SB1_2_4/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_4/Component_Function_1/N4  ( .A1(\SB1_2_4/i1_7 ), .A2(
        \SB1_2_4/i0[8] ), .A3(\SB1_2_4/i0_4 ), .ZN(
        \SB1_2_4/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_17/Component_Function_0/N4  ( .A1(\SB1_2_17/i0[7] ), .A2(
        \SB1_2_17/i0_3 ), .A3(\SB1_2_17/i0_0 ), .ZN(
        \SB1_2_17/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_21/Component_Function_1/N2  ( .A1(n3682), .A2(
        \SB1_2_21/i1_7 ), .A3(\SB1_2_21/i0[8] ), .ZN(
        \SB1_2_21/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_6/Component_Function_0/N1  ( .A1(\SB1_2_6/i0[10] ), .A2(
        \SB1_2_6/i0[9] ), .ZN(\SB1_2_6/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_20/Component_Function_3/N4  ( .A1(n2909), .A2(n2893), .A3(
        \SB1_2_20/i3[0] ), .ZN(\SB1_2_20/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_16/Component_Function_3/N4  ( .A1(\SB1_2_16/i1_5 ), .A2(
        \SB1_2_16/i0[8] ), .A3(\SB1_2_16/i3[0] ), .ZN(
        \SB1_2_16/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_15/Component_Function_0/N4  ( .A1(\SB1_2_15/i0[7] ), .A2(
        \SB1_2_15/i0_3 ), .A3(\SB1_2_15/i0_0 ), .ZN(
        \SB1_2_15/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_2/Component_Function_2/N1  ( .A1(\SB1_2_2/i1_5 ), .A2(
        \SB1_2_2/i0[10] ), .A3(\SB1_2_2/i1[9] ), .ZN(
        \SB1_2_2/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_11/Component_Function_1/N3  ( .A1(\SB1_2_11/i1_5 ), .A2(
        \SB1_2_11/i0[6] ), .A3(\SB1_2_11/i0[9] ), .ZN(
        \SB1_2_11/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB1_2_12/Component_Function_1/N1  ( .A1(\SB1_2_12/i0_3 ), .A2(
        \SB1_2_12/i1[9] ), .ZN(\SB1_2_12/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB1_2_26/Component_Function_1/N1  ( .A1(\RI1[2][35] ), .A2(
        \SB1_2_26/i1[9] ), .ZN(\SB1_2_26/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_9/Component_Function_3/N1  ( .A1(\SB1_2_9/i1[9] ), .A2(
        \SB1_2_9/i0_3 ), .A3(\SB1_2_9/i0[6] ), .ZN(
        \SB1_2_9/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_12/Component_Function_3/N3  ( .A1(\SB1_2_12/i1[9] ), .A2(
        \SB1_2_12/i1_7 ), .A3(\SB1_2_12/i0[10] ), .ZN(
        \SB1_2_12/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_20/Component_Function_0/N2  ( .A1(n2893), .A2(
        \SB1_2_20/i0[7] ), .A3(\SB1_2_20/i0[6] ), .ZN(
        \SB1_2_20/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_23/Component_Function_3/N1  ( .A1(\SB1_2_23/i1[9] ), .A2(
        \SB1_2_23/i0_3 ), .A3(\SB1_2_23/i0[6] ), .ZN(
        \SB1_2_23/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_22/Component_Function_2/N2  ( .A1(\SB1_2_22/i0_3 ), .A2(
        \SB1_2_22/i0[10] ), .A3(\SB1_2_22/i0[6] ), .ZN(
        \SB1_2_22/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_26/Component_Function_3/N2  ( .A1(\SB2_2_26/i0_0 ), .A2(
        \SB2_2_26/i0_3 ), .A3(\SB2_2_26/i0_4 ), .ZN(
        \SB2_2_26/Component_Function_3/NAND4_in[1] ) );
  BUF_X2 \SB2_2_28/BUF_0  ( .I(\SB1_2_1/buf_output[0] ), .Z(\SB2_2_28/i0[9] )
         );
  NAND3_X1 \SB2_2_22/Component_Function_1/N4  ( .A1(\SB2_2_22/i1_7 ), .A2(
        \SB2_2_22/i0[8] ), .A3(\SB2_2_22/i0_4 ), .ZN(
        \SB2_2_22/Component_Function_1/NAND4_in[3] ) );
  INV_X1 \SB2_2_8/INV_1  ( .I(\SB1_2_12/buf_output[1] ), .ZN(\SB2_2_8/i1_7 )
         );
  NAND2_X1 \SB2_2_23/Component_Function_0/N1  ( .A1(\SB2_2_23/i0[10] ), .A2(
        \SB2_2_23/i0[9] ), .ZN(\SB2_2_23/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_26/Component_Function_1/N2  ( .A1(\SB2_2_26/i0_3 ), .A2(
        \SB2_2_26/i1_7 ), .A3(\SB2_2_26/i0[8] ), .ZN(
        \SB2_2_26/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_17/Component_Function_0/N2  ( .A1(\SB2_2_17/i0[8] ), .A2(
        \SB2_2_17/i0[7] ), .A3(\SB2_2_17/i0[6] ), .ZN(
        \SB2_2_17/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_13/Component_Function_4/N4  ( .A1(\SB2_2_13/i1[9] ), .A2(
        n1394), .A3(n580), .ZN(\SB2_2_13/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_27/Component_Function_5/N4  ( .A1(\SB2_2_27/i0[9] ), .A2(
        \SB2_2_27/i0[6] ), .A3(\SB1_2_28/buf_output[4] ), .ZN(
        \SB2_2_27/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_31/Component_Function_1/N2  ( .A1(\SB2_2_31/i0_3 ), .A2(
        \SB2_2_31/i1_7 ), .A3(\SB2_2_31/i0[8] ), .ZN(
        \SB2_2_31/Component_Function_1/NAND4_in[1] ) );
  INV_X1 \SB1_3_26/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[30] ), .ZN(
        \SB1_3_26/i3[0] ) );
  BUF_X2 \SB1_3_6/BUF_0  ( .I(\MC_ARK_ARC_1_2/buf_output[150] ), .Z(
        \SB1_3_6/i0[9] ) );
  NAND3_X1 \SB1_3_25/Component_Function_4/N3  ( .A1(\SB1_3_25/i0[9] ), .A2(
        \SB1_3_25/i0[10] ), .A3(\SB1_3_25/i0_3 ), .ZN(
        \SB1_3_25/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_29/Component_Function_0/N2  ( .A1(\SB1_3_29/i0[8] ), .A2(
        \SB1_3_29/i0[7] ), .A3(\SB1_3_29/i0[6] ), .ZN(
        \SB1_3_29/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_3_17/Component_Function_0/N1  ( .A1(\SB1_3_17/i0[10] ), .A2(
        \SB1_3_17/i0[9] ), .ZN(\SB1_3_17/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_29/Component_Function_0/N4  ( .A1(\SB1_3_29/i0[7] ), .A2(
        \SB1_3_29/i0_3 ), .A3(\RI1[3][14] ), .ZN(
        \SB1_3_29/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB1_3_29/Component_Function_0/N1  ( .A1(\SB1_3_29/i0[10] ), .A2(
        \SB1_3_29/i0[9] ), .ZN(\SB1_3_29/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_3/Component_Function_3/N2  ( .A1(\SB1_3_3/i0_0 ), .A2(
        \SB1_3_3/i0_3 ), .A3(\SB1_3_3/i0_4 ), .ZN(
        \SB1_3_3/Component_Function_3/NAND4_in[1] ) );
  INV_X1 \SB1_3_17/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[84] ), .ZN(
        \SB1_3_17/i3[0] ) );
  INV_X1 \SB1_3_23/INV_4  ( .I(\SB1_3_23/i0_4 ), .ZN(\SB1_3_23/i0[7] ) );
  NAND3_X1 \SB1_3_5/Component_Function_2/N1  ( .A1(\SB1_3_5/i1_5 ), .A2(
        \SB1_3_5/i0[10] ), .A3(\SB1_3_5/i1[9] ), .ZN(
        \SB1_3_5/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_20/Component_Function_3/N2  ( .A1(\SB1_3_20/i0_0 ), .A2(
        \SB1_3_20/i0_3 ), .A3(\SB1_3_20/i0_4 ), .ZN(
        \SB1_3_20/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_3/Component_Function_4/N4  ( .A1(\SB1_3_3/i1[9] ), .A2(
        \SB1_3_3/i1_5 ), .A3(\SB1_3_3/i0_4 ), .ZN(
        \SB1_3_3/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_16/Component_Function_0/N4  ( .A1(\SB1_3_16/i0[7] ), .A2(
        \SB1_3_16/i0_3 ), .A3(\SB1_3_16/i0_0 ), .ZN(
        \SB1_3_16/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_23/Component_Function_1/N3  ( .A1(\SB1_3_23/i1_5 ), .A2(
        \SB1_3_23/i0[6] ), .A3(\SB1_3_23/i0[9] ), .ZN(
        \SB1_3_23/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_10/Component_Function_1/N3  ( .A1(\SB1_3_10/i1_5 ), .A2(
        \SB1_3_10/i0[6] ), .A3(\SB1_3_10/i0[9] ), .ZN(
        \SB1_3_10/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB1_3_15/Component_Function_1/N1  ( .A1(\SB1_3_15/i0_3 ), .A2(
        \SB1_3_15/i1[9] ), .ZN(\SB1_3_15/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_25/Component_Function_3/N1  ( .A1(\SB1_3_25/i1[9] ), .A2(
        \SB1_3_25/i0_3 ), .A3(\SB1_3_25/i0[6] ), .ZN(
        \SB1_3_25/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_29/Component_Function_3/N3  ( .A1(\SB1_3_29/i1[9] ), .A2(
        \SB1_3_29/i1_7 ), .A3(\SB1_3_29/i0[10] ), .ZN(
        \SB1_3_29/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_27/Component_Function_1/N2  ( .A1(\SB2_3_27/i0_3 ), .A2(
        \SB2_3_27/i1_7 ), .A3(\SB2_3_27/i0[8] ), .ZN(
        \SB2_3_27/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_15/Component_Function_5/N1  ( .A1(n809), .A2(
        \SB2_3_15/i3[0] ), .ZN(\SB2_3_15/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_10/Component_Function_1/N4  ( .A1(\SB2_3_10/i1_7 ), .A2(
        \SB2_3_10/i0[8] ), .A3(\SB1_3_11/buf_output[4] ), .ZN(
        \SB2_3_10/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_31/Component_Function_4/N4  ( .A1(\SB2_3_31/i1[9] ), .A2(
        \SB2_3_31/i1_5 ), .A3(\SB2_3_31/i0_4 ), .ZN(
        \SB2_3_31/Component_Function_4/NAND4_in[3] ) );
  NAND2_X1 \SB2_3_0/Component_Function_5/N1  ( .A1(\SB2_3_0/i0_0 ), .A2(
        \SB2_3_0/i3[0] ), .ZN(\SB2_3_0/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_10/Component_Function_3/N4  ( .A1(\SB2_3_10/i1_5 ), .A2(
        \SB2_3_10/i0[8] ), .A3(\SB2_3_10/i3[0] ), .ZN(
        \SB2_3_10/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_15/Component_Function_4/N4  ( .A1(\SB2_3_15/i1[9] ), .A2(
        \SB2_3_15/i1_5 ), .A3(\SB1_3_16/buf_output[4] ), .ZN(
        \SB2_3_15/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_31/Component_Function_3/N3  ( .A1(\SB2_3_31/i1[9] ), .A2(
        \SB2_3_31/i1_7 ), .A3(\SB2_3_31/i0[10] ), .ZN(
        \SB2_3_31/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_20/Component_Function_1/N3  ( .A1(\SB2_3_20/i1_5 ), .A2(
        \SB2_3_20/i0[6] ), .A3(\SB2_3_20/i0[9] ), .ZN(
        \SB2_3_20/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_8/Component_Function_1/N4  ( .A1(\SB2_3_8/i1_7 ), .A2(
        \SB2_3_8/i0[8] ), .A3(\SB1_3_9/buf_output[4] ), .ZN(
        \SB2_3_8/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_18/Component_Function_1/N3  ( .A1(\SB2_3_18/i1_5 ), .A2(
        \SB2_3_18/i0[6] ), .A3(\SB2_3_18/i0[9] ), .ZN(
        \SB2_3_18/Component_Function_1/NAND4_in[2] ) );
  INV_X1 \SB3_23/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[48] ), .ZN(
        \SB3_23/i3[0] ) );
  INV_X1 \SB3_19/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[72] ), .ZN(
        \SB3_19/i3[0] ) );
  NAND3_X1 \SB3_23/Component_Function_3/N3  ( .A1(\SB3_23/i1[9] ), .A2(
        \SB3_23/i1_7 ), .A3(\SB3_23/i0[10] ), .ZN(
        \SB3_23/Component_Function_3/NAND4_in[2] ) );
  BUF_X2 \SB3_7/BUF_0  ( .I(\MC_ARK_ARC_1_3/buf_output[144] ), .Z(
        \SB3_7/i0[9] ) );
  BUF_X2 \SB3_26/BUF_0  ( .I(\MC_ARK_ARC_1_3/buf_output[30] ), .Z(
        \SB3_26/i0[9] ) );
  NAND3_X1 \SB3_10/Component_Function_1/N4  ( .A1(\SB3_10/i1_7 ), .A2(
        \SB3_10/i0[8] ), .A3(\SB3_10/i0_4 ), .ZN(
        \SB3_10/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_14/Component_Function_1/N3  ( .A1(\SB3_14/i1_5 ), .A2(
        \SB3_14/i0[6] ), .A3(\SB3_14/i0[9] ), .ZN(
        \SB3_14/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_15/Component_Function_5/N4  ( .A1(\SB3_15/i0[9] ), .A2(
        \SB3_15/i0[6] ), .A3(\SB3_15/i0_4 ), .ZN(
        \SB3_15/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB3_28/Component_Function_3/N1  ( .A1(\SB3_28/i1[9] ), .A2(
        \SB3_28/i0_3 ), .A3(\SB3_28/i0[6] ), .ZN(
        \SB3_28/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB3_28/Component_Function_4/N3  ( .A1(\SB3_28/i0[9] ), .A2(
        \SB3_28/i0[10] ), .A3(\SB3_28/i0_3 ), .ZN(
        \SB3_28/Component_Function_4/NAND4_in[2] ) );
  NAND2_X1 \SB3_19/Component_Function_0/N1  ( .A1(\SB3_19/i0[10] ), .A2(
        \SB3_19/i0[9] ), .ZN(\SB3_19/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_21/Component_Function_1/N3  ( .A1(\SB3_21/i1_5 ), .A2(
        \SB3_21/i0[6] ), .A3(\SB3_21/i0[9] ), .ZN(
        \SB3_21/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_16/Component_Function_2/N2  ( .A1(\SB3_16/i0_3 ), .A2(
        \SB3_16/i0[10] ), .A3(\SB3_16/i0[6] ), .ZN(
        \SB3_16/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB3_26/Component_Function_5/N4  ( .A1(\SB3_26/i0[9] ), .A2(
        \SB3_26/i0[6] ), .A3(\SB3_26/i0_4 ), .ZN(
        \SB3_26/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB3_8/Component_Function_1/N3  ( .A1(\SB3_8/i1_5 ), .A2(
        \SB3_8/i0[6] ), .A3(\SB3_8/i0[9] ), .ZN(
        \SB3_8/Component_Function_1/NAND4_in[2] ) );
  INV_X1 \SB4_7/INV_1  ( .I(\SB3_11/buf_output[1] ), .ZN(\SB4_7/i1_7 ) );
  BUF_X2 \SB4_5/BUF_1  ( .I(\SB3_9/buf_output[1] ), .Z(\SB4_5/i0[6] ) );
  INV_X1 \SB4_23/INV_5  ( .I(\SB3_23/buf_output[5] ), .ZN(\SB4_23/i1_5 ) );
  NAND2_X1 \SB4_13/Component_Function_5/N1  ( .A1(\SB4_13/i0_0 ), .A2(
        \SB4_13/i3[0] ), .ZN(\SB4_13/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB4_19/Component_Function_1/N1  ( .A1(\SB4_19/i0_3 ), .A2(
        \SB4_19/i1[9] ), .ZN(\SB4_19/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB4_23/Component_Function_0/N1  ( .A1(\SB4_23/i0[10] ), .A2(
        \SB4_23/i0[9] ), .ZN(\SB4_23/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U180 ( .A1(\SB4_23/i0_4 ), .A2(\SB4_23/i0[6] ), .A3(\SB4_23/i0[9] ), 
        .ZN(n2630) );
  NAND3_X1 U570 ( .A1(\SB4_11/i0[10] ), .A2(\SB4_11/i0[9] ), .A3(\SB4_11/i0_3 ), .ZN(n2636) );
  NAND3_X1 U571 ( .A1(\SB4_25/i0_0 ), .A2(\SB4_25/i0_3 ), .A3(\SB4_25/i0[7] ), 
        .ZN(\SB4_25/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U575 ( .A1(\SB4_2/i0[6] ), .A2(\SB4_2/i0[8] ), .A3(\SB4_2/i0[7] ), 
        .ZN(\SB4_2/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U577 ( .A1(\SB4_19/i0_0 ), .A2(\SB4_19/i3[0] ), .A3(\SB4_19/i1_7 ), 
        .ZN(\SB4_19/Component_Function_4/NAND4_in[1] ) );
  NAND2_X1 U578 ( .A1(\SB4_26/i0[10] ), .A2(\SB4_26/i0[9] ), .ZN(n1709) );
  NAND3_X1 U579 ( .A1(\SB4_12/i0_4 ), .A2(\SB4_12/i1[9] ), .A3(\SB4_12/i0_3 ), 
        .ZN(n2518) );
  BUF_X2 U594 ( .I(\SB3_14/buf_output[1] ), .Z(\SB4_10/i0[6] ) );
  BUF_X2 U597 ( .I(\SB3_19/buf_output[1] ), .Z(\SB4_15/i0[6] ) );
  NAND3_X1 U605 ( .A1(\SB3_3/i0_0 ), .A2(\SB3_3/i1_5 ), .A3(\SB3_3/i0_4 ), 
        .ZN(n2108) );
  NAND3_X1 U607 ( .A1(\SB3_8/i1_7 ), .A2(\SB3_8/i0[8] ), .A3(\SB3_8/i0_4 ), 
        .ZN(\SB3_8/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U609 ( .A1(\SB3_7/i0_4 ), .A2(\SB3_7/i0[9] ), .A3(\SB3_7/i0[6] ), 
        .ZN(n1982) );
  NAND3_X1 U610 ( .A1(\SB3_21/i0_0 ), .A2(\SB3_21/i1_5 ), .A3(\SB3_21/i0_4 ), 
        .ZN(n878) );
  NAND3_X1 U616 ( .A1(\SB3_27/i0_3 ), .A2(n4764), .A3(\SB3_27/i0_4 ), .ZN(
        n2723) );
  NAND3_X1 U618 ( .A1(\SB3_3/i0[6] ), .A2(\SB3_3/i0_4 ), .A3(\SB3_3/i0[9] ), 
        .ZN(n2191) );
  NAND3_X1 U622 ( .A1(\SB3_17/i0_4 ), .A2(\SB3_17/i1[9] ), .A3(\SB3_17/i1_5 ), 
        .ZN(n1600) );
  NAND3_X1 U639 ( .A1(\SB3_18/i0[8] ), .A2(\SB3_18/i3[0] ), .A3(\SB3_18/i1_5 ), 
        .ZN(n2498) );
  NAND3_X1 U640 ( .A1(\SB3_9/i0[8] ), .A2(\SB3_9/i3[0] ), .A3(\SB3_9/i1_5 ), 
        .ZN(n2480) );
  NAND3_X1 U643 ( .A1(\SB3_28/i0_0 ), .A2(\SB3_28/i0[7] ), .A3(\SB3_28/i0_3 ), 
        .ZN(n2484) );
  NAND3_X1 U645 ( .A1(\SB3_8/i3[0] ), .A2(\SB3_8/i0[8] ), .A3(\SB3_8/i1_5 ), 
        .ZN(n2113) );
  BUF_X2 U656 ( .I(\MC_ARK_ARC_1_3/buf_output[115] ), .Z(\SB3_12/i0[6] ) );
  BUF_X2 U659 ( .I(\MC_ARK_ARC_1_3/buf_output[48] ), .Z(\SB3_23/i0[9] ) );
  NAND3_X1 U664 ( .A1(\SB3_23/i0[8] ), .A2(\SB3_23/i1_5 ), .A3(\SB3_23/i3[0] ), 
        .ZN(n2818) );
  INV_X1 U724 ( .I(\SB1_3_18/buf_output[1] ), .ZN(\SB2_3_14/i1_7 ) );
  BUF_X2 U727 ( .I(\SB1_3_18/buf_output[1] ), .Z(\SB2_3_14/i0[6] ) );
  INV_X1 U730 ( .I(\SB1_3_23/buf_output[0] ), .ZN(\SB2_3_18/i3[0] ) );
  NAND3_X1 U755 ( .A1(\SB1_3_19/i0[10] ), .A2(\SB1_3_19/i0_3 ), .A3(
        \SB1_3_19/i0[6] ), .ZN(\SB1_3_19/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U757 ( .A1(\SB1_3_17/i0[8] ), .A2(\SB1_3_17/i3[0] ), .A3(
        \SB1_3_17/i1_5 ), .ZN(\SB1_3_17/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U760 ( .A1(\SB1_3_19/i0_0 ), .A2(\SB1_3_19/i0_3 ), .A3(
        \SB1_3_19/i0_4 ), .ZN(\SB1_3_19/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U776 ( .A1(\SB1_3_20/i3[0] ), .A2(\SB1_3_20/i0_0 ), .A3(
        \SB1_3_20/i1_7 ), .ZN(\SB1_3_20/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U783 ( .A1(\SB1_3_25/i1_5 ), .A2(\SB1_3_25/i3[0] ), .A3(
        \SB1_3_25/i0[8] ), .ZN(n1163) );
  NAND3_X1 U789 ( .A1(\SB1_3_7/i0[8] ), .A2(\SB1_3_7/i1_5 ), .A3(
        \SB1_3_7/i3[0] ), .ZN(\SB1_3_7/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U805 ( .A1(\SB1_3_12/i0_0 ), .A2(\SB1_3_12/i1_7 ), .A3(
        \SB1_3_12/i3[0] ), .ZN(\SB1_3_12/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U806 ( .A1(\SB1_3_16/i0[9] ), .A2(\SB1_3_16/i0[8] ), .A3(
        \SB1_3_16/i0_0 ), .ZN(n1311) );
  NAND3_X1 U813 ( .A1(\SB1_3_9/i0[10] ), .A2(\SB1_3_9/i0_3 ), .A3(
        \SB1_3_9/i0[9] ), .ZN(n2444) );
  NAND3_X1 U830 ( .A1(\SB2_2_23/i3[0] ), .A2(\SB2_2_23/i0_0 ), .A3(
        \SB2_2_23/i1_7 ), .ZN(\SB2_2_23/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U834 ( .A1(\SB2_2_22/i0_3 ), .A2(\SB2_2_22/i0[8] ), .A3(
        \SB2_2_22/i1_7 ), .ZN(n1099) );
  NAND3_X1 U835 ( .A1(n722), .A2(\SB2_2_15/i0[8] ), .A3(\SB2_2_15/i0[6] ), 
        .ZN(\SB2_2_15/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 U857 ( .A1(\SB1_2_13/Component_Function_5/NAND4_in[3] ), .A2(
        \SB1_2_13/Component_Function_5/NAND4_in[0] ), .ZN(n1259) );
  NAND3_X1 U859 ( .A1(\RI1[2][35] ), .A2(\SB1_2_26/i0[7] ), .A3(
        \SB1_2_26/i0_0 ), .ZN(\SB1_2_26/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U866 ( .A1(\RI1[2][47] ), .A2(\SB1_2_24/i0_0 ), .A3(\SB1_2_24/i0_4 ), .ZN(\SB1_2_24/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U868 ( .A1(\SB1_2_8/i0[6] ), .A2(\SB1_2_8/i0_4 ), .A3(
        \SB1_2_8/i0[9] ), .ZN(n2097) );
  NAND3_X1 U869 ( .A1(\SB1_2_3/i0[10] ), .A2(\SB1_2_3/i0_4 ), .A3(
        \SB1_2_3/i0_3 ), .ZN(\SB1_2_3/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 U871 ( .A1(\SB1_2_8/Component_Function_4/NAND4_in[3] ), .A2(n2294), 
        .ZN(n2293) );
  NAND2_X1 U876 ( .A1(\SB1_2_28/Component_Function_4/NAND4_in[3] ), .A2(n2026), 
        .ZN(n2025) );
  NAND3_X1 U879 ( .A1(\SB1_2_4/i0_3 ), .A2(\SB1_2_4/i1[9] ), .A3(
        \SB1_2_4/i0_4 ), .ZN(\SB1_2_4/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U880 ( .A1(\SB1_2_11/i0[9] ), .A2(\SB1_2_11/i0_0 ), .A3(
        \SB1_2_11/i0[8] ), .ZN(n1411) );
  NAND3_X1 U883 ( .A1(\SB1_2_31/i0[9] ), .A2(\SB1_2_31/i1_5 ), .A3(
        \SB1_2_31/i0[6] ), .ZN(\SB1_2_31/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U891 ( .A1(\SB1_2_31/i0_0 ), .A2(\SB1_2_31/i3[0] ), .A3(
        \SB1_2_31/i1_7 ), .ZN(\SB1_2_31/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U900 ( .A1(\SB1_2_9/i0_0 ), .A2(\SB1_2_9/i0_3 ), .A3(
        \SB1_2_9/i0[7] ), .ZN(n1293) );
  NAND3_X1 U904 ( .A1(\SB1_2_6/i0_0 ), .A2(\SB1_2_6/i1_5 ), .A3(\SB1_2_6/i0_4 ), .ZN(\SB1_2_6/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U906 ( .A1(\SB1_2_20/i0[6] ), .A2(\SB1_2_20/i1[9] ), .A3(
        \SB1_2_20/i0_3 ), .ZN(\SB1_2_20/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U907 ( .A1(\SB1_2_16/i1_5 ), .A2(\SB1_2_16/i1[9] ), .A3(
        \SB1_2_16/i0_4 ), .ZN(\SB1_2_16/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U921 ( .A1(\SB1_2_12/i0_0 ), .A2(\SB1_2_12/i1_5 ), .A3(
        \SB1_2_12/i0_4 ), .ZN(n2260) );
  NAND3_X1 U925 ( .A1(\SB1_2_19/i0[10] ), .A2(\SB1_2_19/i1[9] ), .A3(
        \SB1_2_19/i1_7 ), .ZN(n2230) );
  NAND3_X1 U931 ( .A1(\SB1_2_16/i0[8] ), .A2(\SB1_2_16/i1_7 ), .A3(
        \RI1[2][95] ), .ZN(\SB1_2_16/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U944 ( .A1(\SB2_1_6/i0_3 ), .A2(\SB2_1_6/i0_0 ), .A3(
        \SB2_1_6/i0[7] ), .ZN(\SB2_1_6/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U948 ( .A1(\SB2_1_13/i0_3 ), .A2(\SB2_1_13/i1_7 ), .A3(
        \SB2_1_13/i0[8] ), .ZN(\SB2_1_13/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U959 ( .A1(\SB2_1_10/i0_0 ), .A2(\SB2_1_10/i0[9] ), .A3(
        \SB2_1_10/i0[8] ), .ZN(n1344) );
  NAND3_X1 U962 ( .A1(n2535), .A2(\SB2_1_5/i0[8] ), .A3(\SB2_1_5/i0[6] ), .ZN(
        n2078) );
  NAND3_X1 U964 ( .A1(\SB2_1_24/i0_3 ), .A2(\SB2_1_24/i0[8] ), .A3(
        \SB2_1_24/i1_7 ), .ZN(\SB2_1_24/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 U974 ( .A1(\SB2_1_10/i0_0 ), .A2(\SB2_1_10/i3[0] ), .ZN(n977) );
  NAND3_X1 U994 ( .A1(\SB1_1_15/i0[6] ), .A2(\SB1_1_15/i1_5 ), .A3(
        \SB1_1_15/i0[9] ), .ZN(n1445) );
  NAND3_X1 U1000 ( .A1(\SB1_1_20/i0_0 ), .A2(\SB1_1_20/i1_7 ), .A3(
        \SB1_1_20/i3[0] ), .ZN(\SB1_1_20/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U1011 ( .A1(\MC_ARK_ARC_1_0/buf_output[82] ), .A2(\SB1_1_18/i0[8] ), 
        .A3(\SB1_1_18/i1_7 ), .ZN(\SB1_1_18/Component_Function_1/NAND4_in[3] )
         );
  NAND3_X1 U1025 ( .A1(\SB1_1_17/i0_0 ), .A2(\SB1_1_17/i3[0] ), .A3(
        \SB1_1_17/i1_7 ), .ZN(\SB1_1_17/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U1026 ( .A1(\SB1_1_24/i0[8] ), .A2(\SB1_1_24/i3[0] ), .A3(
        \SB1_1_24/i1_5 ), .ZN(n2876) );
  NAND3_X1 U1027 ( .A1(\SB1_1_15/i0_0 ), .A2(\SB1_1_15/i0_3 ), .A3(
        \SB1_1_15/i0[7] ), .ZN(n2835) );
  NAND3_X1 U1038 ( .A1(\SB1_1_30/i0_3 ), .A2(\SB1_1_30/i1[9] ), .A3(
        \SB1_1_30/i0_4 ), .ZN(\SB1_1_30/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1039 ( .A1(\SB1_1_11/i0[10] ), .A2(\SB1_1_11/i0_3 ), .A3(
        \SB1_1_11/i0[9] ), .ZN(\SB1_1_11/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1041 ( .A1(\SB1_1_6/i0[9] ), .A2(\SB1_1_6/i0_4 ), .A3(
        \SB1_1_6/i0[6] ), .ZN(n2095) );
  NAND3_X1 U1042 ( .A1(\SB1_1_11/i0_0 ), .A2(\SB1_1_11/i1_7 ), .A3(
        \SB1_1_11/i3[0] ), .ZN(n1562) );
  NAND3_X1 U1049 ( .A1(\SB1_1_1/i0_4 ), .A2(\SB1_1_1/i0[8] ), .A3(
        \SB1_1_1/i1_7 ), .ZN(n2416) );
  NAND3_X1 U1050 ( .A1(\SB1_1_6/i0[9] ), .A2(\SB1_1_6/i1_5 ), .A3(
        \SB1_1_6/i0[6] ), .ZN(\SB1_1_6/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1051 ( .A1(\SB1_1_19/i0_0 ), .A2(\SB1_1_19/i3[0] ), .A3(
        \SB1_1_19/i1_7 ), .ZN(\SB1_1_19/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U1055 ( .A1(\SB1_1_3/i0_0 ), .A2(\SB1_1_3/i0_3 ), .A3(
        \SB1_1_3/i0[7] ), .ZN(n1133) );
  NAND3_X1 U1056 ( .A1(\SB1_1_13/i0[10] ), .A2(\SB1_1_13/i0[9] ), .A3(
        \SB1_1_13/i0_3 ), .ZN(n1328) );
  INV_X1 U1062 ( .I(\MC_ARK_ARC_1_0/buf_output[108] ), .ZN(\SB1_1_13/i3[0] )
         );
  NAND3_X1 U1070 ( .A1(\SB2_0_24/i0[9] ), .A2(\SB2_0_24/i0_3 ), .A3(
        \SB2_0_24/i0[8] ), .ZN(\SB2_0_24/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1071 ( .A1(n2679), .A2(\SB2_0_27/i0[8] ), .A3(\SB2_0_27/i0_0 ), 
        .ZN(\SB2_0_27/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U1074 ( .A1(\SB2_0_16/i0_0 ), .A2(\SB2_0_16/i1_5 ), .A3(
        \SB2_0_16/i0_4 ), .ZN(\SB2_0_16/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U1078 ( .A1(\SB2_0_25/i1_7 ), .A2(\SB2_0_25/i0_3 ), .A3(
        \SB2_0_25/i0[8] ), .ZN(n1804) );
  NAND3_X1 U1082 ( .A1(\RI3[0][22] ), .A2(\SB1_0_1/buf_output[0] ), .A3(
        \SB1_0_0/buf_output[1] ), .ZN(n2014) );
  NAND3_X1 U1094 ( .A1(\SB1_0_13/buf_output[1] ), .A2(\SB2_0_9/i0[9] ), .A3(
        \SB2_0_9/i0_4 ), .ZN(n1097) );
  INV_X1 U1100 ( .I(\SB1_0_12/buf_output[5] ), .ZN(\SB2_0_12/i1_5 ) );
  INV_X1 U1102 ( .I(\RI3[0][66] ), .ZN(\SB2_0_20/i3[0] ) );
  INV_X1 U1107 ( .I(\RI3[0][126] ), .ZN(\SB2_0_10/i3[0] ) );
  NAND3_X1 U1108 ( .A1(\SB2_0_23/i0[9] ), .A2(\SB2_0_23/i0[6] ), .A3(
        \SB2_0_23/i0_4 ), .ZN(n950) );
  NAND3_X1 U1114 ( .A1(\SB1_0_25/i0_4 ), .A2(n263), .A3(n264), .ZN(n2204) );
  NAND3_X1 U1115 ( .A1(\SB1_0_0/i0_0 ), .A2(\SB1_0_0/i0[10] ), .A3(n1376), 
        .ZN(n1265) );
  NAND3_X1 U1116 ( .A1(\SB1_0_13/i0_3 ), .A2(\SB1_0_13/i0[9] ), .A3(
        \SB1_0_13/i0[10] ), .ZN(n2417) );
  NAND3_X1 U1119 ( .A1(\SB1_0_28/i0_3 ), .A2(\SB1_0_28/i0[6] ), .A3(
        \SB1_0_28/i1[9] ), .ZN(n1990) );
  NAND3_X1 U1121 ( .A1(\SB1_0_17/i0_3 ), .A2(\SB1_0_17/i0_0 ), .A3(
        \SB1_0_17/i0[7] ), .ZN(\SB1_0_17/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U1122 ( .A1(\SB1_0_29/i0[9] ), .A2(\SB1_0_29/i0_3 ), .A3(
        \SB1_0_29/i0[8] ), .ZN(n834) );
  NAND3_X1 U1125 ( .A1(\SB1_0_3/i0_3 ), .A2(\SB1_0_3/i0[6] ), .A3(
        \SB1_0_3/i1[9] ), .ZN(n2253) );
  NAND3_X1 U1127 ( .A1(\SB1_0_28/i0_3 ), .A2(\SB1_0_28/i0[8] ), .A3(
        \SB1_0_28/i1_7 ), .ZN(\SB1_0_28/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U1128 ( .A1(\SB1_0_21/i0_4 ), .A2(\SB1_0_21/i1_5 ), .A3(
        \SB1_0_21/i1[9] ), .ZN(\SB1_0_21/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U1129 ( .A1(\SB1_0_12/i0_0 ), .A2(\SB1_0_12/i0[9] ), .A3(
        \SB1_0_12/i0[8] ), .ZN(\SB1_0_12/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U1132 ( .A1(\SB1_0_28/i0_3 ), .A2(\SB1_0_28/i0_0 ), .A3(
        \SB1_0_28/i0[7] ), .ZN(\SB1_0_28/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U1133 ( .A1(\SB1_0_21/i0_0 ), .A2(\SB1_0_21/i0[9] ), .A3(
        \SB1_0_21/i0[8] ), .ZN(n1214) );
  NAND3_X1 U1134 ( .A1(\SB1_0_14/i0[8] ), .A2(\SB1_0_14/i0[9] ), .A3(
        \SB1_0_14/i0_0 ), .ZN(n2402) );
  NAND3_X1 U1139 ( .A1(\SB1_0_28/i0[10] ), .A2(\SB1_0_28/i0_3 ), .A3(
        \SB1_0_28/i0[9] ), .ZN(n1784) );
  NAND3_X1 U1140 ( .A1(\SB1_0_24/i0_0 ), .A2(\SB1_0_24/i3[0] ), .A3(
        \SB1_0_24/i1_7 ), .ZN(n2424) );
  INV_X1 U1149 ( .I(\SB3_28/buf_output[2] ), .ZN(\SB4_25/i1[9] ) );
  BUF_X2 U1150 ( .I(\SB3_28/buf_output[2] ), .Z(\SB4_25/i0_0 ) );
  INV_X1 U1153 ( .I(\MC_ARK_ARC_1_2/buf_output[37] ), .ZN(\SB1_3_25/i1_7 ) );
  BUF_X2 U1154 ( .I(\MC_ARK_ARC_1_2/buf_output[37] ), .Z(\SB1_3_25/i0[6] ) );
  NAND3_X1 U1155 ( .A1(\SB1_3_3/i0[10] ), .A2(\SB1_3_3/i1[9] ), .A3(
        \SB1_3_3/i1_7 ), .ZN(n1546) );
  NAND3_X1 U1157 ( .A1(\SB1_3_3/i0_3 ), .A2(\SB1_3_3/i0[10] ), .A3(
        \SB1_3_3/i0[6] ), .ZN(\SB1_3_3/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U1167 ( .A1(\SB2_3_8/i0_3 ), .A2(\SB2_3_8/i1_7 ), .A3(
        \SB2_3_8/i0[8] ), .ZN(\SB2_3_8/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U1177 ( .A1(\SB3_19/i1_5 ), .A2(\SB3_19/i0[6] ), .A3(\SB3_19/i0[9] ), .ZN(\SB3_19/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1178 ( .A1(\SB3_19/i0[9] ), .A2(\SB3_19/i0[6] ), .A3(\SB3_19/i0_4 ), .ZN(\SB3_19/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U1182 ( .A1(\SB4_2/i0[6] ), .A2(\SB4_2/i0_3 ), .A3(\SB4_2/i0[10] ), 
        .ZN(n2469) );
  NAND3_X1 U1195 ( .A1(\SB2_0_20/i0[7] ), .A2(\SB2_0_20/i0_3 ), .A3(
        \SB2_0_20/i0_0 ), .ZN(\SB2_0_20/Component_Function_0/NAND4_in[3] ) );
  INV_X1 U1200 ( .I(\MC_ARK_ARC_1_3/buf_output[21] ), .ZN(\SB3_28/i0[8] ) );
  BUF_X2 U1201 ( .I(\MC_ARK_ARC_1_3/buf_output[21] ), .Z(\SB3_28/i0[10] ) );
  NAND3_X1 U1206 ( .A1(\SB1_1_20/i0_3 ), .A2(\SB1_1_20/i0[9] ), .A3(
        \SB1_1_20/i0[10] ), .ZN(n2203) );
  INV_X1 U1209 ( .I(\SB3_18/buf_output[2] ), .ZN(\SB4_15/i1[9] ) );
  BUF_X2 U1210 ( .I(\SB3_18/buf_output[2] ), .Z(\SB4_15/i0_0 ) );
  INV_X1 U1217 ( .I(\MC_ARK_ARC_1_3/buf_output[81] ), .ZN(\SB3_18/i0[8] ) );
  BUF_X2 U1218 ( .I(\MC_ARK_ARC_1_3/buf_output[81] ), .Z(\SB3_18/i0[10] ) );
  INV_X1 U1233 ( .I(\MC_ARK_ARC_1_1/buf_output[1] ), .ZN(\SB1_2_31/i1_7 ) );
  INV_X1 U1246 ( .I(\MC_ARK_ARC_1_0/buf_output[180] ), .ZN(\SB1_1_1/i3[0] ) );
  NAND3_X1 U1253 ( .A1(\SB3_9/i0[7] ), .A2(\SB3_9/i0_3 ), .A3(\SB3_9/i0_0 ), 
        .ZN(\SB3_9/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U1254 ( .A1(\SB3_9/i0_3 ), .A2(\SB3_9/i0[8] ), .A3(\SB3_9/i0[9] ), 
        .ZN(\SB3_9/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1255 ( .A1(\SB1_3_22/i1[9] ), .A2(\SB1_3_22/i0_3 ), .A3(
        \SB1_3_22/i0[6] ), .ZN(\SB1_3_22/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U1257 ( .A1(\SB4_1/i1[9] ), .A2(\SB4_1/i1_5 ), .A3(\SB4_1/i0_4 ), 
        .ZN(\SB4_1/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U1262 ( .A1(\SB4_4/i0[10] ), .A2(n3655), .A3(\SB4_4/i1_7 ), .ZN(
        \SB4_4/Component_Function_3/NAND4_in[2] ) );
  CLKBUF_X4 U1265 ( .I(\MC_ARK_ARC_1_2/buf_output[140] ), .Z(\SB1_3_8/i0_0 )
         );
  NAND2_X1 U1269 ( .A1(\SB4_8/i0[10] ), .A2(\SB4_8/i0[9] ), .ZN(
        \SB4_8/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U1270 ( .A1(\SB4_23/i1[9] ), .A2(\SB4_23/i1_7 ), .A3(
        \SB4_23/i0[10] ), .ZN(\SB4_23/Component_Function_3/NAND4_in[2] ) );
  BUF_X2 U1276 ( .I(\MC_ARK_ARC_1_3/buf_output[181] ), .Z(\SB3_1/i0[6] ) );
  NAND3_X1 U1303 ( .A1(\SB4_23/i0_0 ), .A2(\SB4_23/i0_4 ), .A3(\SB4_23/i1_5 ), 
        .ZN(n2628) );
  INV_X1 U1310 ( .I(\MC_ARK_ARC_1_3/buf_output[78] ), .ZN(\SB3_18/i3[0] ) );
  NAND3_X1 U1311 ( .A1(\SB1_2_25/i1_5 ), .A2(\SB1_2_25/i0[6] ), .A3(
        \SB1_2_25/i0[9] ), .ZN(\SB1_2_25/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1314 ( .A1(\SB1_3_27/i0_3 ), .A2(\SB1_3_27/i0_4 ), .A3(
        \SB1_3_27/i1[9] ), .ZN(\SB1_3_27/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1328 ( .A1(\SB4_25/i3[0] ), .A2(\SB4_25/i0_0 ), .A3(\SB4_25/i1_7 ), 
        .ZN(\SB4_25/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U1329 ( .A1(\SB1_2_14/i0[8] ), .A2(\SB1_2_14/i0[9] ), .A3(
        \MC_ARK_ARC_1_1/buf_output[107] ), .ZN(
        \SB1_2_14/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1333 ( .A1(\SB2_2_5/i0_3 ), .A2(\SB2_2_5/i0_0 ), .A3(
        \SB1_2_6/buf_output[4] ), .ZN(n1661) );
  NAND3_X1 U1336 ( .A1(\SB3_26/i0[10] ), .A2(\SB3_26/i1[9] ), .A3(
        \SB3_26/i1_7 ), .ZN(n2362) );
  NAND3_X1 U1337 ( .A1(\SB3_26/i0[6] ), .A2(\SB3_26/i0[10] ), .A3(
        \SB3_26/i0_3 ), .ZN(n1842) );
  NAND3_X1 U1338 ( .A1(\SB3_26/i0_0 ), .A2(\SB3_26/i0[6] ), .A3(
        \SB3_26/i0[10] ), .ZN(\SB3_26/Component_Function_5/NAND4_in[1] ) );
  INV_X1 U1339 ( .I(\MC_ARK_ARC_1_3/buf_output[99] ), .ZN(\SB3_15/i0[8] ) );
  NAND3_X1 U1342 ( .A1(\SB1_1_31/i1[9] ), .A2(\SB1_1_31/i0_3 ), .A3(
        \SB1_1_31/i0[6] ), .ZN(\SB1_1_31/Component_Function_3/NAND4_in[0] ) );
  NAND2_X1 U1344 ( .A1(\SB1_1_31/i0_3 ), .A2(\SB1_1_31/i1[9] ), .ZN(
        \SB1_1_31/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U1348 ( .A1(\SB2_1_30/i0[8] ), .A2(\SB2_1_30/i1_7 ), .A3(
        \SB2_1_30/i0_4 ), .ZN(n1129) );
  NAND3_X1 U1353 ( .A1(\SB1_0_6/i0_0 ), .A2(\SB1_0_6/i1_5 ), .A3(
        \SB1_0_6/i0_4 ), .ZN(n1279) );
  NAND3_X1 U1354 ( .A1(\SB1_0_6/i0_0 ), .A2(\SB1_0_6/i3[0] ), .A3(
        \SB1_0_6/i1_7 ), .ZN(n1310) );
  NAND2_X1 U1363 ( .A1(\SB4_8/i0_3 ), .A2(\SB4_8/i1[9] ), .ZN(n768) );
  NAND3_X1 U1365 ( .A1(n1389), .A2(\SB4_27/i1_7 ), .A3(\SB4_27/i0[10] ), .ZN(
        \SB4_27/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U1367 ( .A1(\SB2_0_12/i0_4 ), .A2(\SB2_0_12/i0_0 ), .A3(
        \SB2_0_12/i1_5 ), .ZN(n2414) );
  NAND3_X1 U1373 ( .A1(\SB1_2_14/i1_5 ), .A2(\SB1_2_14/i0[10] ), .A3(
        \SB1_2_14/i1[9] ), .ZN(\SB1_2_14/Component_Function_2/NAND4_in[0] ) );
  CLKBUF_X4 U1375 ( .I(\SB1_3_24/buf_output[4] ), .Z(\SB2_3_23/i0_4 ) );
  CLKBUF_X4 U1404 ( .I(\MC_ARK_ARC_1_1/buf_output[104] ), .Z(\SB1_2_14/i0_0 )
         );
  NAND3_X1 U1407 ( .A1(\SB1_0_10/i1[9] ), .A2(\SB1_0_10/i1_7 ), .A3(
        \SB1_0_10/i0[10] ), .ZN(\SB1_0_10/Component_Function_3/NAND4_in[2] )
         );
  NAND3_X1 U1413 ( .A1(\SB2_3_12/i0[6] ), .A2(\SB1_3_13/buf_output[4] ), .A3(
        n1603), .ZN(n2099) );
  BUF_X2 U1419 ( .I(\SB3_10/buf_output[3] ), .Z(\SB4_8/i0[10] ) );
  INV_X1 U1428 ( .I(\SB3_8/buf_output[1] ), .ZN(\SB4_4/i1_7 ) );
  BUF_X2 U1429 ( .I(\SB3_8/buf_output[1] ), .Z(\SB4_4/i0[6] ) );
  BUF_X2 U1430 ( .I(\SB3_6/buf_output[3] ), .Z(\SB4_4/i0[10] ) );
  BUF_X2 U1446 ( .I(\SB1_0_13/buf_output[1] ), .Z(\SB2_0_9/i0[6] ) );
  INV_X1 U1447 ( .I(\SB1_0_13/buf_output[1] ), .ZN(\SB2_0_9/i1_7 ) );
  NAND3_X1 U1448 ( .A1(\SB3_5/i3[0] ), .A2(\SB3_5/i0_0 ), .A3(\SB3_5/i1_7 ), 
        .ZN(\SB3_5/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U1450 ( .A1(\SB1_0_26/buf_output[0] ), .A2(\SB1_0_21/buf_output[5] ), .A3(\SB2_0_21/i0[8] ), .ZN(n1674) );
  NAND3_X1 U1451 ( .A1(\SB2_0_21/i0_3 ), .A2(\SB2_0_21/i1_7 ), .A3(
        \SB2_0_21/i0[8] ), .ZN(\SB2_0_21/Component_Function_1/NAND4_in[1] ) );
  INV_X1 U1458 ( .I(n250), .ZN(\SB1_0_30/i1[9] ) );
  BUF_X2 U1459 ( .I(n250), .Z(\SB1_0_30/i0_0 ) );
  NAND3_X1 U1465 ( .A1(\SB1_3_27/i0[10] ), .A2(\SB1_3_27/i0[9] ), .A3(
        \SB1_3_27/i0_3 ), .ZN(\SB1_3_27/Component_Function_4/NAND4_in[2] ) );
  INV_X1 U1483 ( .I(\MC_ARK_ARC_1_3/buf_output[103] ), .ZN(\SB3_14/i1_7 ) );
  NAND3_X1 U1486 ( .A1(\SB4_26/i0_3 ), .A2(\SB4_26/i0[10] ), .A3(
        \SB4_26/i0[6] ), .ZN(\SB4_26/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U1490 ( .A1(\SB4_6/i0_0 ), .A2(\SB4_6/i0[6] ), .A3(\SB4_6/i0[10] ), 
        .ZN(\SB4_6/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1499 ( .A1(\SB1_1_9/i0[10] ), .A2(\SB1_1_9/i1[9] ), .A3(
        \SB1_1_9/i1_7 ), .ZN(\SB1_1_9/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U1506 ( .A1(\SB1_3_30/i1[9] ), .A2(\SB1_3_30/i1_5 ), .A3(
        \SB1_3_30/i0_4 ), .ZN(\SB1_3_30/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U1513 ( .A1(\SB2_0_12/i0_3 ), .A2(\RI3[0][114] ), .A3(
        \SB2_0_12/i0[8] ), .ZN(\SB2_0_12/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1514 ( .A1(\SB2_0_12/i0[9] ), .A2(\SB2_0_12/i0[10] ), .A3(
        \SB2_0_12/i0_3 ), .ZN(\SB2_0_12/Component_Function_4/NAND4_in[2] ) );
  INV_X1 U1518 ( .I(\SB1_1_10/buf_output[1] ), .ZN(\SB2_1_6/i1_7 ) );
  NAND3_X1 U1521 ( .A1(\SB3_8/i0_3 ), .A2(\SB3_8/i1_7 ), .A3(\SB3_8/i0[8] ), 
        .ZN(\SB3_8/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U1533 ( .A1(\SB1_1_3/i1_7 ), .A2(\SB1_1_3/i0[8] ), .A3(
        \SB1_1_3/i0_4 ), .ZN(\SB1_1_3/Component_Function_1/NAND4_in[3] ) );
  INV_X1 U1537 ( .I(\MC_ARK_ARC_1_3/buf_output[126] ), .ZN(\SB3_10/i3[0] ) );
  INV_X1 U1547 ( .I(\MC_ARK_ARC_1_2/buf_output[48] ), .ZN(\SB1_3_23/i3[0] ) );
  BUF_X2 U1548 ( .I(\MC_ARK_ARC_1_2/buf_output[48] ), .Z(\SB1_3_23/i0[9] ) );
  NAND3_X1 U1552 ( .A1(\SB1_3_4/i0_3 ), .A2(\SB1_3_4/i0[8] ), .A3(
        \SB1_3_4/i0[9] ), .ZN(\SB1_3_4/Component_Function_2/NAND4_in[2] ) );
  BUF_X2 U1568 ( .I(\MC_ARK_ARC_1_3/buf_output[111] ), .Z(\SB3_13/i0[10] ) );
  INV_X1 U1569 ( .I(\MC_ARK_ARC_1_3/buf_output[111] ), .ZN(\SB3_13/i0[8] ) );
  NAND3_X1 U1585 ( .A1(\SB1_2_5/i1[9] ), .A2(\SB1_2_5/i1_5 ), .A3(
        \SB1_2_5/i0_4 ), .ZN(\SB1_2_5/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U1586 ( .A1(\SB1_2_5/i1[9] ), .A2(\SB1_2_5/i0_3 ), .A3(
        \SB1_2_5/i0[6] ), .ZN(\SB1_2_5/Component_Function_3/NAND4_in[0] ) );
  INV_X1 U1609 ( .I(\MC_ARK_ARC_1_2/buf_output[54] ), .ZN(\SB1_3_22/i3[0] ) );
  NAND3_X1 U1610 ( .A1(\SB3_1/i0[10] ), .A2(\SB3_1/i0_4 ), .A3(\SB3_1/i0_3 ), 
        .ZN(\SB3_1/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U1612 ( .A1(\SB3_1/i0[10] ), .A2(n4765), .A3(\SB3_1/i1_7 ), .ZN(
        n1021) );
  NAND3_X1 U1619 ( .A1(\SB4_12/i0_4 ), .A2(\SB4_12/i0_0 ), .A3(\SB4_12/i0_3 ), 
        .ZN(n2465) );
  BUF_X2 U1625 ( .I(\SB1_3_25/buf_output[1] ), .Z(\SB2_3_21/i0[6] ) );
  NAND3_X1 U1627 ( .A1(\SB1_1_6/i0_3 ), .A2(\SB1_1_6/i0[10] ), .A3(
        \SB1_1_6/i0[6] ), .ZN(\SB1_1_6/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U1631 ( .A1(\SB1_2_0/i0_3 ), .A2(\SB1_2_0/i1_7 ), .A3(
        \SB1_2_0/i0[8] ), .ZN(\SB1_2_0/Component_Function_1/NAND4_in[1] ) );
  INV_X1 U1632 ( .I(\MC_ARK_ARC_1_0/buf_output[139] ), .ZN(\SB1_1_8/i1_7 ) );
  CLKBUF_X4 U1646 ( .I(n283), .Z(\SB1_0_19/i0_0 ) );
  INV_X1 U1648 ( .I(\MC_ARK_ARC_1_0/buf_output[151] ), .ZN(\SB1_1_6/i1_7 ) );
  NAND4_X2 U1650 ( .A1(\SB2_1_12/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_12/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_12/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_1_12/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_1_12/buf_output[3] ) );
  INV_X2 U1652 ( .I(\SB1_0_21/buf_output[5] ), .ZN(\SB2_0_21/i1_5 ) );
  NAND3_X1 U1656 ( .A1(\SB3_17/i0[10] ), .A2(\SB3_17/i0_4 ), .A3(\SB3_17/i0_3 ), .ZN(\SB3_17/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U1660 ( .A1(\SB1_0_26/i0[10] ), .A2(\SB1_0_26/i1[9] ), .A3(
        \SB1_0_26/i1_7 ), .ZN(\SB1_0_26/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U1662 ( .A1(\SB1_0_26/i1[9] ), .A2(\SB1_0_26/i1_5 ), .A3(
        \SB1_0_26/i0_4 ), .ZN(\SB1_0_26/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U1666 ( .A1(\SB1_0_13/i1_5 ), .A2(\SB1_0_13/i0[8] ), .A3(
        \SB1_0_13/i3[0] ), .ZN(\SB1_0_13/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U1667 ( .A1(\RI1[1][143] ), .A2(\SB1_1_8/i1_7 ), .A3(
        \SB1_1_8/i0[8] ), .ZN(\SB1_1_8/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U1669 ( .A1(\SB1_1_8/i0[7] ), .A2(\RI1[1][143] ), .A3(
        \SB1_1_8/i0_0 ), .ZN(\SB1_1_8/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U1670 ( .A1(\SB1_1_8/i0[10] ), .A2(\SB1_1_8/i0_4 ), .A3(
        \RI1[1][143] ), .ZN(n1313) );
  INV_X1 U1681 ( .I(\MC_ARK_ARC_1_3/buf_output[31] ), .ZN(\SB3_26/i1_7 ) );
  NAND3_X1 U1682 ( .A1(\SB3_18/i0_3 ), .A2(\SB3_18/i1_7 ), .A3(\SB3_18/i0[8] ), 
        .ZN(\SB3_18/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 U1685 ( .A1(\SB3_18/i0_3 ), .A2(\SB3_18/i1[9] ), .ZN(
        \SB3_18/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U1687 ( .A1(\SB3_18/i0[10] ), .A2(\SB3_18/i0_4 ), .A3(\SB3_18/i0_3 ), .ZN(\SB3_18/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U1688 ( .A1(\SB3_18/i0[9] ), .A2(\SB3_18/i0[10] ), .A3(
        \SB3_18/i0_3 ), .ZN(\SB3_18/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1689 ( .A1(\SB3_18/i0_0 ), .A2(\SB3_18/i0_3 ), .A3(\SB3_18/i0_4 ), 
        .ZN(\SB3_18/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1692 ( .A1(\SB1_3_25/i1[9] ), .A2(\SB1_3_25/i1_5 ), .A3(
        \SB1_3_25/i0_4 ), .ZN(\SB1_3_25/Component_Function_4/NAND4_in[3] ) );
  INV_X1 U1699 ( .I(\MC_ARK_ARC_1_3/buf_output[23] ), .ZN(\SB3_28/i1_5 ) );
  CLKBUF_X4 U1723 ( .I(\MC_ARK_ARC_1_0/buf_output[111] ), .Z(\SB1_1_13/i0[10] ) );
  NAND3_X1 U1740 ( .A1(\SB4_27/i0_4 ), .A2(n2897), .A3(\SB4_27/i1_5 ), .ZN(
        n1156) );
  INV_X1 U1741 ( .I(\MC_ARK_ARC_1_2/buf_output[13] ), .ZN(\SB1_3_29/i1_7 ) );
  INV_X1 U1751 ( .I(\SB3_26/buf_output[3] ), .ZN(\SB4_24/i0[8] ) );
  BUF_X2 U1752 ( .I(\SB3_26/buf_output[3] ), .Z(\SB4_24/i0[10] ) );
  INV_X1 U1755 ( .I(\MC_ARK_ARC_1_0/buf_output[5] ), .ZN(\SB1_1_31/i1_5 ) );
  NOR2_X2 U1758 ( .A1(n1190), .A2(n1189), .ZN(n2535) );
  INV_X1 U1763 ( .I(\MC_ARK_ARC_1_0/buf_output[150] ), .ZN(\SB1_1_6/i3[0] ) );
  NAND3_X1 U1771 ( .A1(\SB1_1_14/i1_5 ), .A2(\SB1_1_14/i0_0 ), .A3(
        \SB1_1_14/i0_4 ), .ZN(\SB1_1_14/Component_Function_2/NAND4_in[3] ) );
  BUF_X2 U1782 ( .I(\SB3_16/buf_output[1] ), .Z(\SB4_12/i0[6] ) );
  BUF_X2 U1793 ( .I(\SB3_20/buf_output[0] ), .Z(\SB4_15/i0[9] ) );
  BUF_X2 U1798 ( .I(\SB3_12/buf_output[2] ), .Z(\SB4_9/i0_0 ) );
  BUF_X2 U1800 ( .I(\SB3_29/buf_output[2] ), .Z(\SB4_26/i0_0 ) );
  BUF_X2 U1806 ( .I(\MC_ARK_ARC_1_3/buf_output[163] ), .Z(\SB3_4/i0[6] ) );
  CLKBUF_X4 U1808 ( .I(\MC_ARK_ARC_1_3/buf_output[61] ), .Z(\SB3_21/i0[6] ) );
  CLKBUF_X4 U1813 ( .I(\SB2_3_10/buf_output[0] ), .Z(\RI5[3][156] ) );
  BUF_X4 U1814 ( .I(\SB2_3_4/buf_output[5] ), .Z(n1365) );
  BUF_X4 U1817 ( .I(\SB2_3_16/buf_output[4] ), .Z(\RI5[3][100] ) );
  CLKBUF_X4 U1818 ( .I(\SB2_3_25/buf_output[1] ), .Z(\RI5[3][61] ) );
  BUF_X4 U1824 ( .I(\SB2_3_19/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[82] ) );
  CLKBUF_X2 U1826 ( .I(\SB1_3_18/buf_output[2] ), .Z(n809) );
  CLKBUF_X4 U1827 ( .I(\SB1_3_29/buf_output[2] ), .Z(\SB2_3_26/i0_0 ) );
  CLKBUF_X4 U1849 ( .I(\SB2_2_15/buf_output[1] ), .Z(\RI5[2][121] ) );
  BUF_X4 U1851 ( .I(\SB2_2_14/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[127] ) );
  BUF_X4 U1853 ( .I(\SB2_2_23/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[58] ) );
  CLKBUF_X4 U1854 ( .I(\SB2_2_20/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[81] ) );
  BUF_X4 U1857 ( .I(\SB2_2_16/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[105] ) );
  BUF_X4 U1860 ( .I(\SB2_2_21/buf_output[1] ), .Z(\RI5[2][85] ) );
  BUF_X4 U1862 ( .I(\SB2_2_19/buf_output[0] ), .Z(\RI5[2][102] ) );
  CLKBUF_X4 U1868 ( .I(\SB1_2_17/buf_output[4] ), .Z(\SB2_2_16/i0_4 ) );
  CLKBUF_X4 U1871 ( .I(\SB1_2_16/buf_output[3] ), .Z(\SB2_2_14/i0[10] ) );
  CLKBUF_X4 U1881 ( .I(\MC_ARK_ARC_1_1/buf_output[126] ), .Z(\SB1_2_10/i0[9] )
         );
  CLKBUF_X4 U1882 ( .I(\MC_ARK_ARC_1_1/buf_output[0] ), .Z(\SB1_2_31/i0[9] )
         );
  BUF_X4 U1891 ( .I(\SB2_1_20/buf_output[0] ), .Z(\RI5[1][96] ) );
  BUF_X4 U1894 ( .I(\SB2_1_31/buf_output[2] ), .Z(\RI5[1][20] ) );
  NAND3_X2 U1896 ( .A1(\SB2_1_16/i0_0 ), .A2(\SB2_1_16/i0[6] ), .A3(
        \SB2_1_16/i0[10] ), .ZN(\SB2_1_16/Component_Function_5/NAND4_in[1] )
         );
  BUF_X2 U1901 ( .I(\SB1_1_27/buf_output[0] ), .Z(\SB2_1_22/i0[9] ) );
  CLKBUF_X4 U1908 ( .I(\MC_ARK_ARC_1_0/buf_output[126] ), .Z(\SB1_1_10/i0[9] )
         );
  BUF_X2 U1909 ( .I(\MC_ARK_ARC_1_0/buf_output[127] ), .Z(\SB1_1_10/i0[6] ) );
  AND2_X1 U1910 ( .A1(\SB1_1_16/i1_7 ), .A2(\SB1_1_16/i3[0] ), .Z(n573) );
  BUF_X4 U1916 ( .I(\SB2_0_17/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[109] ) );
  BUF_X4 U1918 ( .I(\SB2_0_3/buf_output[3] ), .Z(\RI5[0][183] ) );
  CLKBUF_X4 U1922 ( .I(\RI3[0][9] ), .Z(\SB2_0_30/i0[10] ) );
  CLKBUF_X2 U1924 ( .I(\SB2_0_29/i0[9] ), .Z(n1905) );
  NAND2_X1 U1926 ( .A1(\SB1_0_28/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_0_28/Component_Function_4/NAND4_in[0] ), .ZN(n1785) );
  NAND2_X1 U1928 ( .A1(\SB1_0_14/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_0_14/Component_Function_4/NAND4_in[2] ), .ZN(n2403) );
  BUF_X2 U1930 ( .I(n315), .Z(\SB1_0_8/i0[6] ) );
  INV_X1 U1933 ( .I(n386), .ZN(\SB1_0_9/i0[7] ) );
  CLKBUF_X4 U1937 ( .I(n332), .Z(\SB1_0_2/i0[9] ) );
  NAND3_X1 U1938 ( .A1(\SB1_0_10/i0[10] ), .A2(\SB1_0_10/i0_0 ), .A3(
        \SB1_0_10/i0[6] ), .ZN(n2351) );
  NAND3_X1 U1943 ( .A1(\SB1_0_22/i0_4 ), .A2(\SB1_0_22/i1_5 ), .A3(
        \SB1_0_22/i0_0 ), .ZN(\SB1_0_22/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U1945 ( .A1(\SB1_0_29/i0[7] ), .A2(\SB1_0_29/i0_3 ), .A3(
        \SB1_0_29/i0_0 ), .ZN(\SB1_0_29/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U1946 ( .A1(n329), .A2(\SB1_0_3/i0[6] ), .A3(n398), .ZN(
        \SB1_0_3/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U1950 ( .A1(n360), .A2(\SB1_0_22/i0[9] ), .A3(\SB1_0_22/i0[6] ), 
        .ZN(n2773) );
  NAND3_X1 U1952 ( .A1(\SB1_0_22/i0_4 ), .A2(\SB1_0_22/i0[8] ), .A3(
        \SB1_0_22/i1_7 ), .ZN(\SB1_0_22/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U1953 ( .A1(\SB1_0_20/i0[10] ), .A2(\SB1_0_20/i0_4 ), .A3(
        \SB1_0_20/i0_3 ), .ZN(\SB1_0_20/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U1955 ( .A1(\SB1_0_14/i0_3 ), .A2(\SB1_0_14/i1_7 ), .A3(
        \SB1_0_14/i0[8] ), .ZN(\SB1_0_14/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 U1956 ( .A1(\SB1_0_28/i0[10] ), .A2(\SB1_0_28/i0[9] ), .ZN(
        \SB1_0_28/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U1957 ( .A1(\SB1_0_7/i0_3 ), .A2(\SB1_0_7/i0_0 ), .A3(
        \SB1_0_7/i0[7] ), .ZN(n1548) );
  CLKBUF_X4 U1961 ( .I(\SB1_0_22/buf_output[4] ), .Z(\SB2_0_21/i0_4 ) );
  CLKBUF_X4 U1963 ( .I(\SB1_0_14/buf_output[0] ), .Z(\SB2_0_9/i0[9] ) );
  CLKBUF_X4 U1964 ( .I(\SB1_0_4/buf_output[0] ), .Z(\SB2_0_31/i0[9] ) );
  NAND3_X1 U1971 ( .A1(\SB2_0_30/i0_3 ), .A2(\SB2_0_30/i1_7 ), .A3(
        \SB2_0_30/i0[8] ), .ZN(\SB2_0_30/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U1975 ( .A1(\SB2_0_21/i1_5 ), .A2(\SB2_0_21/i0[8] ), .A3(
        \SB2_0_21/i3[0] ), .ZN(\SB2_0_21/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U1980 ( .A1(\SB2_0_11/i1[9] ), .A2(\SB2_0_11/i1_5 ), .A3(
        \SB2_0_11/i0_4 ), .ZN(\SB2_0_11/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U1983 ( .A1(\SB2_0_26/i1[9] ), .A2(\SB2_0_26/i1_5 ), .A3(
        \RI3[0][34] ), .ZN(\SB2_0_26/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U1984 ( .A1(\SB2_0_28/i1[9] ), .A2(\SB2_0_28/i1_5 ), .A3(
        \RI3[0][22] ), .ZN(\SB2_0_28/Component_Function_4/NAND4_in[3] ) );
  CLKBUF_X4 U1992 ( .I(\MC_ARK_ARC_1_0/buf_output[124] ), .Z(\SB1_1_11/i0_4 )
         );
  NAND3_X1 U1994 ( .A1(\SB1_1_2/i1_5 ), .A2(\SB1_1_2/i0[6] ), .A3(
        \SB1_1_2/i0[9] ), .ZN(\SB1_1_2/Component_Function_1/NAND4_in[2] ) );
  CLKBUF_X4 U2000 ( .I(\MC_ARK_ARC_1_0/buf_output[153] ), .Z(\SB1_1_6/i0[10] )
         );
  NAND3_X1 U2001 ( .A1(\SB1_1_28/i1[9] ), .A2(\SB1_1_28/i0_3 ), .A3(
        \SB1_1_28/i0[6] ), .ZN(\SB1_1_28/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2006 ( .A1(\SB1_1_1/i1_5 ), .A2(\SB1_1_1/i0[8] ), .A3(
        \SB1_1_1/i3[0] ), .ZN(\SB1_1_1/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2013 ( .A1(\SB1_1_15/i0[9] ), .A2(\SB1_1_15/i0[10] ), .A3(
        \SB1_1_15/i0_3 ), .ZN(\SB1_1_15/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2014 ( .A1(\SB1_1_18/i0_0 ), .A2(\SB1_1_18/i0_3 ), .A3(
        \SB1_1_18/i0_4 ), .ZN(\SB1_1_18/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2029 ( .A1(\SB2_1_3/i0_0 ), .A2(n5208), .A3(\SB2_1_3/i1_5 ), .ZN(
        n1852) );
  NAND3_X1 U2039 ( .A1(\SB2_1_12/i0[6] ), .A2(\SB2_1_12/i1_5 ), .A3(
        \SB2_1_12/i0[9] ), .ZN(\SB2_1_12/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U2044 ( .A1(\SB2_1_2/i1_7 ), .A2(\SB2_1_2/i0[8] ), .A3(
        \SB1_1_3/buf_output[4] ), .ZN(
        \SB2_1_2/Component_Function_1/NAND4_in[3] ) );
  CLKBUF_X4 U2050 ( .I(\MC_ARK_ARC_1_1/buf_output[55] ), .Z(\SB1_2_22/i0[6] )
         );
  INV_X1 U2054 ( .I(\MC_ARK_ARC_1_1/buf_output[102] ), .ZN(\SB1_2_14/i3[0] )
         );
  NAND3_X1 U2057 ( .A1(\SB1_2_20/i0_3 ), .A2(\SB1_2_20/i0[10] ), .A3(
        \SB1_2_20/i0[6] ), .ZN(\SB1_2_20/Component_Function_2/NAND4_in[1] ) );
  CLKBUF_X4 U2064 ( .I(\MC_ARK_ARC_1_1/buf_output[148] ), .Z(\SB1_2_7/i0_4 )
         );
  NAND3_X1 U2074 ( .A1(\SB1_2_15/i1[9] ), .A2(\SB1_2_15/i0_3 ), .A3(
        \SB1_2_15/i0[6] ), .ZN(\SB1_2_15/Component_Function_3/NAND4_in[0] ) );
  INV_X1 U2080 ( .I(\SB1_2_4/buf_output[1] ), .ZN(\SB2_2_0/i1_7 ) );
  CLKBUF_X4 U2082 ( .I(\SB1_2_21/buf_output[0] ), .Z(\SB2_2_16/i0[9] ) );
  CLKBUF_X4 U2083 ( .I(\SB1_2_11/buf_output[0] ), .Z(\SB2_2_6/i0[9] ) );
  NAND3_X1 U2090 ( .A1(\SB2_2_16/i0_3 ), .A2(\SB2_2_16/i0_0 ), .A3(
        \SB2_2_16/i0[7] ), .ZN(n2650) );
  NAND3_X1 U2102 ( .A1(\SB2_2_23/i0_3 ), .A2(\SB2_2_23/i0[7] ), .A3(
        \SB2_2_23/i0_0 ), .ZN(n2523) );
  INV_X1 U2113 ( .I(\MC_ARK_ARC_1_2/buf_output[162] ), .ZN(\SB1_3_4/i3[0] ) );
  NAND3_X1 U2127 ( .A1(\SB1_3_12/i0[8] ), .A2(\SB1_3_12/i0[7] ), .A3(
        \MC_ARK_ARC_1_2/buf_output[115] ), .ZN(
        \SB1_3_12/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U2144 ( .A1(\SB2_3_30/i0_3 ), .A2(\SB2_3_30/i1_7 ), .A3(
        \SB2_3_30/i0[8] ), .ZN(\SB2_3_30/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U2156 ( .A1(\SB2_3_29/i3[0] ), .A2(\SB2_3_29/i0_0 ), .A3(
        \SB2_3_29/i1_7 ), .ZN(\SB2_3_29/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U2161 ( .A1(\SB2_3_26/i0[6] ), .A2(\SB2_3_26/i0[7] ), .A3(n4750), 
        .ZN(\SB2_3_26/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U2183 ( .A1(\RI1[4][155] ), .A2(\SB3_6/i1[9] ), .A3(\SB3_6/i0[6] ), 
        .ZN(\SB3_6/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2189 ( .A1(\SB3_6/i0[8] ), .A2(\SB3_6/i1_7 ), .A3(\RI1[4][154] ), 
        .ZN(\SB3_6/Component_Function_1/NAND4_in[3] ) );
  BUF_X2 U2193 ( .I(\SB3_0/buf_output[0] ), .Z(\SB4_27/i0[9] ) );
  INV_X1 U2195 ( .I(\SB3_10/buf_output[1] ), .ZN(\SB4_6/i1_7 ) );
  NAND3_X1 U2199 ( .A1(\SB4_25/i0_3 ), .A2(\SB4_25/i0[6] ), .A3(\SB4_25/i1[9] ), .ZN(n2829) );
  NAND3_X1 U2201 ( .A1(\SB4_12/i0_4 ), .A2(\SB4_12/i1_7 ), .A3(\SB4_12/i0[8] ), 
        .ZN(n2032) );
  NAND3_X1 U2205 ( .A1(\SB4_14/i0[6] ), .A2(\SB4_14/i0[8] ), .A3(
        \SB4_14/i0[7] ), .ZN(\SB4_14/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U2207 ( .A1(\SB4_5/i0[10] ), .A2(\SB4_5/i0_3 ), .A3(\SB4_5/i0[6] ), 
        .ZN(n2522) );
  NAND3_X1 U2209 ( .A1(\SB4_0/i0[9] ), .A2(\SB3_3/buf_output[2] ), .A3(
        \SB4_0/i0[8] ), .ZN(\SB4_0/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U2210 ( .A1(\SB3_6/buf_output[2] ), .A2(\SB4_3/i0_4 ), .A3(
        \SB4_3/i1_5 ), .ZN(n2126) );
  NAND2_X1 U2211 ( .A1(\SB4_19/i0_0 ), .A2(\SB4_19/i3[0] ), .ZN(
        \SB4_19/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 U2214 ( .A1(\SB3_6/buf_output[2] ), .A2(\SB4_3/i3[0] ), .ZN(
        \SB4_3/Component_Function_5/NAND4_in[0] ) );
  INV_X1 U2220 ( .I(\SB3_27/buf_output[3] ), .ZN(\SB4_25/i0[8] ) );
  INV_X1 U2221 ( .I(\MC_ARK_ARC_1_3/buf_output[163] ), .ZN(\SB3_4/i1_7 ) );
  XNOR2_X1 U2226 ( .A1(\MC_ARK_ARC_1_3/temp5[125] ), .A2(
        \MC_ARK_ARC_1_3/temp6[125] ), .ZN(n582) );
  NAND4_X2 U2227 ( .A1(\SB1_2_0/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_2_0/Component_Function_2/NAND4_in[0] ), .A3(n2644), .A4(n583), 
        .ZN(\SB1_2_0/buf_output[2] ) );
  NAND3_X2 U2228 ( .A1(\SB1_2_0/i0[9] ), .A2(\SB1_2_0/i0_3 ), .A3(
        \SB1_2_0/i0[8] ), .ZN(n583) );
  XOR2_X1 U2230 ( .A1(\RI5[2][37] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[43] ), 
        .Z(n584) );
  XOR2_X1 U2231 ( .A1(\MC_ARK_ARC_1_2/temp6[85] ), .A2(n585), .Z(
        \MC_ARK_ARC_1_2/buf_output[85] ) );
  NAND4_X2 U2236 ( .A1(\SB2_2_2/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_2_2/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_2_2/Component_Function_0/NAND4_in[1] ), .A4(
        \SB2_2_2/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_2_2/buf_output[0] ) );
  XOR2_X1 U2237 ( .A1(\RI5[1][59] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[95] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[185] ) );
  NAND3_X2 U2254 ( .A1(\SB2_1_16/i0[10] ), .A2(\SB2_1_16/i1_5 ), .A3(
        \SB2_1_16/i1[9] ), .ZN(\SB2_1_16/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U2255 ( .A1(\SB2_2_20/i0_3 ), .A2(\SB2_2_20/i0[9] ), .A3(
        \SB2_2_20/i0[8] ), .ZN(\SB2_2_20/Component_Function_2/NAND4_in[2] ) );
  XOR2_X1 U2258 ( .A1(\RI5[3][65] ), .A2(\RI5[3][29] ), .Z(
        \MC_ARK_ARC_1_3/temp3[155] ) );
  NAND2_X2 U2283 ( .A1(\SB1_0_8/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_0_8/Component_Function_2/NAND4_in[0] ), .ZN(n599) );
  XOR2_X1 U2314 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[123] ), .A2(n5521), .Z(
        n2021) );
  XOR2_X1 U2328 ( .A1(n616), .A2(n1138), .Z(\MC_ARK_ARC_1_1/buf_output[53] )
         );
  XOR2_X1 U2331 ( .A1(\RI5[2][48] ), .A2(\RI5[2][42] ), .Z(
        \MC_ARK_ARC_1_2/temp1[48] ) );
  XOR2_X1 U2332 ( .A1(\RI5[2][48] ), .A2(\RI5[2][54] ), .Z(
        \MC_ARK_ARC_1_2/temp1[54] ) );
  XOR2_X1 U2336 ( .A1(\RI5[0][15] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[51] ), 
        .Z(n618) );
  XOR2_X1 U2346 ( .A1(n623), .A2(n622), .Z(\MC_ARK_ARC_1_1/buf_output[147] )
         );
  XOR2_X1 U2347 ( .A1(\MC_ARK_ARC_1_1/temp2[147] ), .A2(
        \MC_ARK_ARC_1_1/temp4[147] ), .Z(n622) );
  XOR2_X1 U2348 ( .A1(\MC_ARK_ARC_1_1/temp1[147] ), .A2(
        \MC_ARK_ARC_1_1/temp3[147] ), .Z(n623) );
  XOR2_X1 U2351 ( .A1(\RI5[1][5] ), .A2(\RI5[1][173] ), .Z(n624) );
  NAND3_X1 U2354 ( .A1(\SB2_1_31/i0[9] ), .A2(n5510), .A3(\SB2_1_31/i0[6] ), 
        .ZN(\SB2_1_31/Component_Function_1/NAND4_in[2] ) );
  NAND4_X2 U2358 ( .A1(\SB2_1_31/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_1_31/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_31/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_31/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_1_31/buf_output[0] ) );
  XOR2_X1 U2360 ( .A1(\MC_ARK_ARC_1_2/temp5[158] ), .A2(n627), .Z(
        \MC_ARK_ARC_1_2/buf_output[158] ) );
  XOR2_X1 U2361 ( .A1(\MC_ARK_ARC_1_2/temp3[158] ), .A2(
        \MC_ARK_ARC_1_2/temp4[158] ), .Z(n627) );
  INV_X2 U2368 ( .I(\MC_ARK_ARC_1_2/buf_output[53] ), .ZN(\SB1_3_23/i1_5 ) );
  NAND4_X2 U2372 ( .A1(\SB1_1_30/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_1_30/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_1_30/Component_Function_5/NAND4_in[0] ), .A4(n1619), .ZN(
        \SB1_1_30/buf_output[5] ) );
  BUF_X4 U2375 ( .I(\SB1_2_26/buf_output[5] ), .Z(\SB2_2_26/i0_3 ) );
  INV_X2 U2385 ( .I(\RI3[0][33] ), .ZN(\SB2_0_26/i0[8] ) );
  NAND4_X2 U2386 ( .A1(\SB1_0_28/Component_Function_3/NAND4_in[1] ), .A2(n1990), .A3(\SB1_0_28/Component_Function_3/NAND4_in[3] ), .A4(
        \SB1_0_28/Component_Function_3/NAND4_in[2] ), .ZN(\RI3[0][33] ) );
  XOR2_X1 U2387 ( .A1(n634), .A2(\MC_ARK_ARC_1_3/temp4[78] ), .Z(
        \MC_ARK_ARC_1_3/temp6[78] ) );
  XOR2_X1 U2388 ( .A1(\RI5[3][144] ), .A2(\RI5[3][180] ), .Z(n634) );
  XOR2_X1 U2394 ( .A1(\MC_ARK_ARC_1_2/temp1[4] ), .A2(n636), .Z(
        \MC_ARK_ARC_1_2/temp5[4] ) );
  XOR2_X1 U2395 ( .A1(\RI5[2][142] ), .A2(\RI5[2][166] ), .Z(n636) );
  INV_X2 U2397 ( .I(\RI3[0][44] ), .ZN(\SB2_0_24/i1[9] ) );
  NAND4_X2 U2404 ( .A1(\SB2_2_9/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_2_9/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_2_9/Component_Function_4/NAND4_in[3] ), .A4(n639), .ZN(
        \SB2_2_9/buf_output[4] ) );
  XOR2_X1 U2412 ( .A1(n642), .A2(n641), .Z(\MC_ARK_ARC_1_3/temp6[103] ) );
  XOR2_X1 U2413 ( .A1(\RI5[3][13] ), .A2(n508), .Z(n641) );
  XOR2_X1 U2414 ( .A1(\RI5[3][169] ), .A2(\RI5[3][139] ), .Z(n642) );
  NAND4_X2 U2434 ( .A1(\SB2_2_14/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_2_14/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_2_14/Component_Function_0/NAND4_in[0] ), .A4(n649), .ZN(
        \SB2_2_14/buf_output[0] ) );
  XOR2_X1 U2437 ( .A1(\RI5[3][106] ), .A2(\RI5[3][130] ), .Z(n650) );
  INV_X2 U2438 ( .I(\RI3[1][182] ), .ZN(\SB2_1_1/i1[9] ) );
  XOR2_X1 U2451 ( .A1(\MC_ARK_ARC_1_2/temp5[48] ), .A2(n656), .Z(
        \MC_ARK_ARC_1_2/buf_output[48] ) );
  XOR2_X1 U2452 ( .A1(\MC_ARK_ARC_1_2/temp3[48] ), .A2(
        \MC_ARK_ARC_1_2/temp4[48] ), .Z(n656) );
  BUF_X4 U2453 ( .I(\SB2_0_6/buf_output[2] ), .Z(\RI5[0][170] ) );
  NAND3_X1 U2458 ( .A1(\SB1_1_4/i0_3 ), .A2(\SB1_1_4/i0[8] ), .A3(
        \SB1_1_4/i1_7 ), .ZN(\SB1_1_4/Component_Function_1/NAND4_in[1] ) );
  NAND4_X2 U2461 ( .A1(\SB2_2_17/Component_Function_0/NAND4_in[3] ), .A2(n1199), .A3(\SB2_2_17/Component_Function_0/NAND4_in[1] ), .A4(
        \SB2_2_17/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_2_17/buf_output[0] ) );
  NAND4_X2 U2464 ( .A1(\SB2_3_29/Component_Function_0/NAND4_in[1] ), .A2(n659), 
        .A3(n1402), .A4(\SB2_3_29/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_3_29/buf_output[0] ) );
  XOR2_X1 U2467 ( .A1(\MC_ARK_ARC_1_3/temp6[72] ), .A2(n660), .Z(
        \MC_ARK_ARC_1_3/buf_output[72] ) );
  XOR2_X1 U2468 ( .A1(\MC_ARK_ARC_1_3/temp2[72] ), .A2(
        \MC_ARK_ARC_1_3/temp1[72] ), .Z(n660) );
  XOR2_X1 U2469 ( .A1(n661), .A2(\MC_ARK_ARC_1_2/temp2[100] ), .Z(
        \MC_ARK_ARC_1_2/temp5[100] ) );
  XOR2_X1 U2470 ( .A1(\RI5[2][94] ), .A2(\RI5[2][100] ), .Z(n661) );
  NAND3_X2 U2481 ( .A1(\SB2_1_21/i0[10] ), .A2(\SB2_1_21/i1_5 ), .A3(
        \SB2_1_21/i1[9] ), .ZN(\SB2_1_21/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U2490 ( .A1(\MC_ARK_ARC_1_3/temp4[71] ), .A2(
        \MC_ARK_ARC_1_3/temp3[71] ), .Z(\MC_ARK_ARC_1_3/temp6[71] ) );
  NAND4_X2 U2491 ( .A1(\SB1_3_14/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_3_14/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_14/Component_Function_0/NAND4_in[0] ), .A4(n667), .ZN(
        \SB1_3_14/buf_output[0] ) );
  BUF_X4 U2493 ( .I(\SB2_1_19/buf_output[3] ), .Z(\RI5[1][87] ) );
  XOR2_X1 U2498 ( .A1(n671), .A2(n670), .Z(\MC_ARK_ARC_1_2/temp6[101] ) );
  XOR2_X1 U2499 ( .A1(\RI5[2][11] ), .A2(n446), .Z(n670) );
  XOR2_X1 U2500 ( .A1(\RI5[2][167] ), .A2(\RI5[2][137] ), .Z(n671) );
  XOR2_X1 U2501 ( .A1(n672), .A2(\MC_ARK_ARC_1_3/temp2[141] ), .Z(
        \MC_ARK_ARC_1_3/temp5[141] ) );
  XOR2_X1 U2502 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[135] ), .A2(\RI5[3][141] ), 
        .Z(n672) );
  XOR2_X1 U2507 ( .A1(n674), .A2(\MC_ARK_ARC_1_2/temp2[97] ), .Z(
        \MC_ARK_ARC_1_2/temp5[97] ) );
  XOR2_X1 U2508 ( .A1(\RI5[2][91] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[97] ), 
        .Z(n674) );
  NAND4_X2 U2515 ( .A1(\SB1_0_25/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_0_25/Component_Function_1/NAND4_in[0] ), .A3(
        \SB1_0_25/Component_Function_1/NAND4_in[3] ), .A4(
        \SB1_0_25/Component_Function_1/NAND4_in[2] ), .ZN(\RI3[0][61] ) );
  NAND4_X2 U2524 ( .A1(\SB1_0_3/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_3/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_0_3/Component_Function_5/NAND4_in[0] ), .A4(
        \SB1_0_3/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB1_0_3/buf_output[5] ) );
  NAND4_X2 U2528 ( .A1(\SB1_1_10/Component_Function_5/NAND4_in[1] ), .A2(n858), 
        .A3(n1066), .A4(\SB1_1_10/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_10/buf_output[5] ) );
  NAND2_X1 U2541 ( .A1(n2203), .A2(\SB1_1_20/Component_Function_4/NAND4_in[3] ), .ZN(n1040) );
  AND2_X1 U2542 ( .A1(n1967), .A2(n2109), .Z(n2634) );
  NAND3_X1 U2549 ( .A1(n2828), .A2(\SB2_1_30/i0_0 ), .A3(\SB2_1_30/i0_3 ), 
        .ZN(\SB2_1_30/Component_Function_0/NAND4_in[3] ) );
  BUF_X4 U2567 ( .I(\SB2_1_14/buf_output[0] ), .Z(\RI5[1][132] ) );
  XOR2_X1 U2572 ( .A1(n1177), .A2(\MC_ARK_ARC_1_2/temp4[99] ), .Z(n2455) );
  NAND3_X2 U2573 ( .A1(\SB2_3_1/i0[10] ), .A2(\SB2_3_1/i0_0 ), .A3(
        \SB2_3_1/i0[6] ), .ZN(\SB2_3_1/Component_Function_5/NAND4_in[1] ) );
  INV_X2 U2576 ( .I(\SB1_2_17/buf_output[5] ), .ZN(\SB2_2_17/i1_5 ) );
  XOR2_X1 U2578 ( .A1(\RI5[3][189] ), .A2(\RI5[3][183] ), .Z(n693) );
  XOR2_X1 U2583 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[187] ), .A2(\RI5[1][181] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[187] ) );
  NAND2_X1 U2584 ( .A1(\SB2_0_20/i0_4 ), .A2(n1212), .ZN(
        \SB2_0_20/Component_Function_5/NAND4_in[3] ) );
  XOR2_X1 U2588 ( .A1(\RI5[1][191] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[155] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[89] ) );
  NAND3_X2 U2594 ( .A1(\SB2_2_17/i0_3 ), .A2(\SB2_2_17/i0_4 ), .A3(
        \SB2_2_17/i0_0 ), .ZN(\SB2_2_17/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U2602 ( .A1(\SB1_1_6/i0[10] ), .A2(\SB1_1_6/i0[6] ), .A3(
        \SB1_1_6/i0_0 ), .ZN(n699) );
  XOR2_X1 U2605 ( .A1(\MC_ARK_ARC_1_2/temp1[167] ), .A2(
        \MC_ARK_ARC_1_2/temp2[167] ), .Z(n701) );
  BUF_X4 U2611 ( .I(\SB2_1_10/buf_output[5] ), .Z(\RI5[1][131] ) );
  XOR2_X1 U2613 ( .A1(\MC_ARK_ARC_1_0/temp6[140] ), .A2(n706), .Z(
        \MC_ARK_ARC_1_0/buf_output[140] ) );
  XOR2_X1 U2621 ( .A1(n2784), .A2(n708), .Z(\MC_ARK_ARC_1_1/buf_output[16] )
         );
  XOR2_X1 U2622 ( .A1(\MC_ARK_ARC_1_1/temp3[16] ), .A2(
        \MC_ARK_ARC_1_1/temp4[16] ), .Z(n708) );
  XOR2_X1 U2633 ( .A1(\MC_ARK_ARC_1_2/temp5[123] ), .A2(
        \MC_ARK_ARC_1_2/temp6[123] ), .Z(\MC_ARK_ARC_1_2/buf_output[123] ) );
  XOR2_X1 U2637 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[185] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[29] ), .Z(\MC_ARK_ARC_1_1/temp3[119] )
         );
  XOR2_X1 U2641 ( .A1(n712), .A2(\MC_ARK_ARC_1_1/temp6[73] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[73] ) );
  XOR2_X1 U2642 ( .A1(\MC_ARK_ARC_1_1/temp1[73] ), .A2(
        \MC_ARK_ARC_1_1/temp2[73] ), .Z(n712) );
  XOR2_X1 U2644 ( .A1(\RI5[0][110] ), .A2(\RI5[0][134] ), .Z(
        \MC_ARK_ARC_1_0/temp2[164] ) );
  NAND2_X1 U2658 ( .A1(\SB1_1_5/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_1_5/Component_Function_4/NAND4_in[3] ), .ZN(n1157) );
  BUF_X4 U2663 ( .I(\SB2_2_18/buf_output[3] ), .Z(\RI5[2][93] ) );
  NAND3_X1 U2665 ( .A1(\SB1_0_21/i0[10] ), .A2(\SB1_0_21/i1[9] ), .A3(
        \SB1_0_21/i1_7 ), .ZN(n719) );
  XOR2_X1 U2668 ( .A1(n1800), .A2(n721), .Z(n1351) );
  XOR2_X1 U2669 ( .A1(\RI5[3][48] ), .A2(\RI5[3][42] ), .Z(n721) );
  INV_X4 U2670 ( .I(n2369), .ZN(\SB2_0_20/i0_4 ) );
  INV_X2 U2672 ( .I(\SB2_0_6/i0[10] ), .ZN(\SB2_0_6/i0[8] ) );
  XOR2_X1 U2677 ( .A1(n725), .A2(n724), .Z(\MC_ARK_ARC_1_3/temp5[83] ) );
  XOR2_X1 U2678 ( .A1(\RI5[3][29] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[53] ), 
        .Z(n724) );
  XOR2_X1 U2679 ( .A1(\RI5[3][77] ), .A2(\RI5[3][83] ), .Z(n725) );
  XOR2_X1 U2680 ( .A1(\RI5[2][188] ), .A2(\RI5[2][32] ), .Z(n1537) );
  XOR2_X1 U2687 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[152] ), .A2(\RI5[3][188] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[86] ) );
  XOR2_X1 U2690 ( .A1(\RI5[2][110] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[74] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[8] ) );
  XOR2_X1 U2694 ( .A1(\RI5[2][104] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[68] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[2] ) );
  XOR2_X1 U2700 ( .A1(n729), .A2(n185), .Z(Ciphertext[75]) );
  XOR2_X1 U2702 ( .A1(n2799), .A2(\MC_ARK_ARC_1_1/temp6[189] ), .Z(n1373) );
  XOR2_X1 U2704 ( .A1(\RI5[2][137] ), .A2(\RI5[2][173] ), .Z(
        \MC_ARK_ARC_1_2/temp3[71] ) );
  INV_X2 U2705 ( .I(\SB1_2_13/buf_output[2] ), .ZN(\SB2_2_10/i1[9] ) );
  NAND4_X2 U2706 ( .A1(\SB1_2_13/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_13/Component_Function_2/NAND4_in[1] ), .A3(n827), .A4(n2795), 
        .ZN(\SB1_2_13/buf_output[2] ) );
  XOR2_X1 U2712 ( .A1(\MC_ARK_ARC_1_1/temp1[90] ), .A2(n733), .Z(
        \MC_ARK_ARC_1_1/temp5[90] ) );
  XOR2_X1 U2713 ( .A1(\RI5[1][36] ), .A2(\RI5[1][60] ), .Z(n733) );
  NAND4_X2 U2720 ( .A1(\SB2_3_0/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_3_0/Component_Function_0/NAND4_in[0] ), .A3(
        \SB2_3_0/Component_Function_0/NAND4_in[2] ), .A4(n735), .ZN(
        \SB2_3_0/buf_output[0] ) );
  NOR2_X2 U2723 ( .A1(n739), .A2(n737), .ZN(n2564) );
  XOR2_X1 U2728 ( .A1(\MC_ARK_ARC_1_3/temp1[180] ), .A2(
        \MC_ARK_ARC_1_3/temp2[180] ), .Z(n740) );
  INV_X1 U2731 ( .I(\SB1_0_7/buf_output[1] ), .ZN(\SB2_0_3/i1_7 ) );
  NAND4_X2 U2732 ( .A1(\SB1_0_7/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_0_7/Component_Function_1/NAND4_in[0] ), .A3(
        \SB1_0_7/Component_Function_1/NAND4_in[3] ), .A4(
        \SB1_0_7/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB1_0_7/buf_output[1] ) );
  INV_X2 U2734 ( .I(\SB1_2_26/buf_output[3] ), .ZN(\SB2_2_24/i0[8] ) );
  NAND3_X1 U2736 ( .A1(\RI3[1][60] ), .A2(\SB1_1_25/buf_output[1] ), .A3(
        \SB1_1_22/buf_output[4] ), .ZN(n2439) );
  XOR2_X1 U2742 ( .A1(n744), .A2(\MC_ARK_ARC_1_0/temp6[170] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[170] ) );
  NAND2_X1 U2744 ( .A1(\SB1_1_26/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_1_26/Component_Function_0/NAND4_in[1] ), .ZN(n2617) );
  INV_X1 U2745 ( .I(\SB3_21/buf_output[1] ), .ZN(\SB4_17/i1_7 ) );
  NAND4_X2 U2746 ( .A1(\SB3_21/Component_Function_1/NAND4_in[1] ), .A2(
        \SB3_21/Component_Function_1/NAND4_in[3] ), .A3(
        \SB3_21/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_21/Component_Function_1/NAND4_in[0] ), .ZN(\SB3_21/buf_output[1] ) );
  NAND2_X1 U2754 ( .A1(\SB1_0_21/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_0_21/Component_Function_4/NAND4_in[3] ), .ZN(n747) );
  INV_X2 U2757 ( .I(\RI3[0][164] ), .ZN(\SB2_0_4/i1[9] ) );
  NAND4_X2 U2758 ( .A1(\SB1_0_7/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_0_7/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_0_7/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_7/Component_Function_2/NAND4_in[3] ), .ZN(\RI3[0][164] ) );
  XOR2_X1 U2759 ( .A1(n1327), .A2(\MC_ARK_ARC_1_1/temp1[36] ), .Z(
        \MC_ARK_ARC_1_1/temp5[36] ) );
  NAND3_X1 U2774 ( .A1(\SB2_0_6/i0[7] ), .A2(\SB2_0_6/i0[8] ), .A3(
        \SB2_0_6/i0[6] ), .ZN(\SB2_0_6/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U2780 ( .A1(n756), .A2(\MC_ARK_ARC_1_3/temp4[140] ), .Z(n2845) );
  XOR2_X1 U2781 ( .A1(\RI5[3][50] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[14] ), 
        .Z(n756) );
  XOR2_X1 U2782 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[76] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[112] ), .Z(\MC_ARK_ARC_1_0/temp3[10] )
         );
  XOR2_X1 U2783 ( .A1(n757), .A2(\MC_ARK_ARC_1_3/temp5[83] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[83] ) );
  NAND4_X2 U2790 ( .A1(\SB1_0_0/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_0_0/Component_Function_3/NAND4_in[2] ), .A3(
        \SB1_0_0/Component_Function_3/NAND4_in[3] ), .A4(n759), .ZN(
        \RI3[0][9] ) );
  NAND3_X1 U2793 ( .A1(\RI3[0][191] ), .A2(\SB2_0_0/i0_0 ), .A3(
        \SB2_0_0/i0[7] ), .ZN(n760) );
  NAND4_X2 U2794 ( .A1(n842), .A2(\SB1_0_25/Component_Function_0/NAND4_in[1] ), 
        .A3(\SB1_0_25/Component_Function_0/NAND4_in[3] ), .A4(
        \SB1_0_25/Component_Function_0/NAND4_in[0] ), .ZN(\RI3[0][66] ) );
  NAND3_X1 U2795 ( .A1(\SB1_1_20/buf_output[1] ), .A2(\SB2_1_16/i0[8] ), .A3(
        \SB2_1_16/i0[7] ), .ZN(\SB2_1_16/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U2796 ( .A1(\MC_ARK_ARC_1_1/temp3[79] ), .A2(
        \MC_ARK_ARC_1_1/temp4[79] ), .Z(n761) );
  XOR2_X1 U2797 ( .A1(\MC_ARK_ARC_1_0/temp6[10] ), .A2(
        \MC_ARK_ARC_1_0/temp5[10] ), .Z(\MC_ARK_ARC_1_0/buf_output[10] ) );
  XOR2_X1 U2798 ( .A1(n763), .A2(n762), .Z(\MC_ARK_ARC_1_0/buf_output[161] )
         );
  XOR2_X1 U2799 ( .A1(\MC_ARK_ARC_1_0/temp2[161] ), .A2(
        \MC_ARK_ARC_1_0/temp4[161] ), .Z(n762) );
  BUF_X4 U2803 ( .I(\SB2_3_21/buf_output[3] ), .Z(\RI5[3][75] ) );
  XOR2_X1 U2805 ( .A1(n765), .A2(n29), .Z(Ciphertext[53]) );
  NAND4_X2 U2806 ( .A1(\SB4_23/Component_Function_5/NAND4_in[1] ), .A2(
        \SB4_23/Component_Function_5/NAND4_in[2] ), .A3(n2630), .A4(
        \SB4_23/Component_Function_5/NAND4_in[0] ), .ZN(n765) );
  NAND4_X2 U2809 ( .A1(\SB1_2_16/Component_Function_2/NAND4_in[0] ), .A2(n1604), .A3(\SB1_2_16/Component_Function_2/NAND4_in[1] ), .A4(
        \SB1_2_16/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB1_2_16/buf_output[2] ) );
  NAND3_X2 U2812 ( .A1(\SB1_3_24/i0[10] ), .A2(\SB1_3_24/i0_3 ), .A3(
        \SB1_3_24/i0[6] ), .ZN(\SB1_3_24/Component_Function_2/NAND4_in[1] ) );
  XOR2_X1 U2827 ( .A1(\MC_ARK_ARC_1_2/temp5[80] ), .A2(
        \MC_ARK_ARC_1_2/temp6[80] ), .Z(\MC_ARK_ARC_1_2/buf_output[80] ) );
  NAND4_X2 U2828 ( .A1(\SB2_3_12/Component_Function_3/NAND4_in[3] ), .A2(
        \SB2_3_12/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_3_12/Component_Function_3/NAND4_in[0] ), .A4(
        \SB2_3_12/Component_Function_3/NAND4_in[1] ), .ZN(
        \SB2_3_12/buf_output[3] ) );
  NAND4_X2 U2831 ( .A1(n2364), .A2(\SB3_10/Component_Function_1/NAND4_in[3] ), 
        .A3(\SB3_10/Component_Function_1/NAND4_in[0] ), .A4(n1575), .ZN(
        \SB3_10/buf_output[1] ) );
  XOR2_X1 U2835 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[59] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[95] ), .Z(\MC_ARK_ARC_1_2/temp3[185] )
         );
  NAND4_X2 U2838 ( .A1(\SB2_3_25/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_3_25/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_3_25/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_25/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_3_25/buf_output[1] ) );
  NAND3_X1 U2854 ( .A1(\SB1_1_28/i0[10] ), .A2(\SB1_1_28/i0_3 ), .A3(
        \SB1_1_28/i0_4 ), .ZN(\SB1_1_28/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 U2858 ( .A1(\SB2_0_11/i0_3 ), .A2(\SB2_0_11/i1[9] ), .A3(
        \SB2_0_11/i0_4 ), .ZN(n780) );
  NAND4_X2 U2862 ( .A1(\SB2_1_12/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_12/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_12/Component_Function_4/NAND4_in[3] ), .A4(n782), .ZN(
        \SB2_1_12/buf_output[4] ) );
  BUF_X4 U2864 ( .I(\SB2_3_0/buf_output[3] ), .Z(\RI5[3][9] ) );
  NAND4_X2 U2865 ( .A1(\SB2_0_10/Component_Function_0/NAND4_in[1] ), .A2(n1912), .A3(\SB2_0_10/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_10/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_0_10/buf_output[0] ) );
  NAND3_X2 U2878 ( .A1(\SB1_1_4/i0_4 ), .A2(\SB1_1_4/i0_3 ), .A3(
        \SB1_1_4/i1[9] ), .ZN(\SB1_1_4/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U2883 ( .A1(n2083), .A2(\MC_ARK_ARC_1_1/temp6[1] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[1] ) );
  XOR2_X1 U2888 ( .A1(\RI5[0][63] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[69] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[69] ) );
  NAND4_X2 U2889 ( .A1(\SB2_3_17/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_3_17/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_3_17/Component_Function_0/NAND4_in[0] ), .A4(n793), .ZN(
        \SB2_3_17/buf_output[0] ) );
  NAND3_X1 U2894 ( .A1(\SB3_30/i0_3 ), .A2(\SB3_30/i0[10] ), .A3(\SB3_30/i0_4 ), .ZN(n795) );
  NAND4_X2 U2895 ( .A1(n796), .A2(\SB2_2_25/Component_Function_4/NAND4_in[1] ), 
        .A3(\SB2_2_25/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_2_25/Component_Function_4/NAND4_in[2] ), .ZN(
        \SB2_2_25/buf_output[4] ) );
  NAND4_X2 U2905 ( .A1(n1337), .A2(\SB1_1_23/Component_Function_5/NAND4_in[3] ), .A3(\SB1_1_23/Component_Function_5/NAND4_in[0] ), .A4(
        \SB1_1_23/Component_Function_5/NAND4_in[1] ), .ZN(
        \SB1_1_23/buf_output[5] ) );
  NAND3_X2 U2906 ( .A1(\SB2_0_24/i1_7 ), .A2(\SB2_0_24/i0[10] ), .A3(
        \SB2_0_24/i1[9] ), .ZN(n800) );
  NAND3_X1 U2915 ( .A1(\SB1_0_25/i0_3 ), .A2(\SB1_0_25/i1_7 ), .A3(
        \SB1_0_25/i0[8] ), .ZN(\SB1_0_25/Component_Function_1/NAND4_in[1] ) );
  BUF_X4 U2918 ( .I(\SB2_1_31/buf_output[0] ), .Z(\RI5[1][30] ) );
  XOR2_X1 U2920 ( .A1(\RI5[3][66] ), .A2(\RI5[3][30] ), .Z(n805) );
  XOR2_X1 U2922 ( .A1(\SB2_2_27/buf_output[4] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[58] ), .Z(\MC_ARK_ARC_1_2/temp2[88] ) );
  NAND3_X1 U2925 ( .A1(\SB4_30/i0_3 ), .A2(\SB4_30/i0_4 ), .A3(n4751), .ZN(
        \SB4_30/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U2936 ( .A1(\RI5[0][191] ), .A2(\RI5[0][5] ), .Z(
        \MC_ARK_ARC_1_0/temp1[5] ) );
  INV_X2 U2941 ( .I(\MC_ARK_ARC_1_3/buf_output[14] ), .ZN(\SB3_29/i1[9] ) );
  NAND3_X2 U2944 ( .A1(\RI3[0][191] ), .A2(\SB2_0_0/i1[9] ), .A3(\RI3[0][190] ), .ZN(\SB2_0_0/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2948 ( .A1(\SB4_27/i0_4 ), .A2(n2897), .A3(\SB4_27/i0_3 ), .ZN(
        \SB4_27/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2959 ( .A1(\SB3_28/i1_7 ), .A2(\SB3_28/i0_3 ), .A3(\SB3_28/i0[8] ), 
        .ZN(\SB3_28/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U2963 ( .A1(\MC_ARK_ARC_1_3/temp3[75] ), .A2(
        \MC_ARK_ARC_1_3/temp4[75] ), .Z(\MC_ARK_ARC_1_3/temp6[75] ) );
  NAND4_X2 U2968 ( .A1(\SB3_28/Component_Function_4/NAND4_in[1] ), .A2(
        \SB3_28/Component_Function_4/NAND4_in[0] ), .A3(
        \SB3_28/Component_Function_4/NAND4_in[3] ), .A4(
        \SB3_28/Component_Function_4/NAND4_in[2] ), .ZN(\SB3_28/buf_output[4] ) );
  NAND3_X2 U2977 ( .A1(n4763), .A2(\SB2_3_17/i0[8] ), .A3(\SB2_3_17/i3[0] ), 
        .ZN(\SB2_3_17/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U2980 ( .A1(n822), .A2(n1878), .Z(\MC_ARK_ARC_1_1/buf_output[139] )
         );
  XOR2_X1 U2981 ( .A1(\MC_ARK_ARC_1_1/temp1[139] ), .A2(
        \MC_ARK_ARC_1_1/temp3[139] ), .Z(n822) );
  NAND4_X2 U2986 ( .A1(\SB3_23/Component_Function_4/NAND4_in[2] ), .A2(
        \SB3_23/Component_Function_4/NAND4_in[0] ), .A3(
        \SB3_23/Component_Function_4/NAND4_in[1] ), .A4(n823), .ZN(
        \SB3_23/buf_output[4] ) );
  NAND3_X1 U2990 ( .A1(\SB1_0_10/i1_5 ), .A2(\SB1_0_10/i3[0] ), .A3(
        \SB1_0_10/i0[8] ), .ZN(\SB1_0_10/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U2991 ( .A1(\RI5[3][2] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[38] ), 
        .Z(n2311) );
  NAND3_X2 U2992 ( .A1(\SB1_3_31/i0_3 ), .A2(\SB1_3_31/i0[8] ), .A3(
        \SB1_3_31/i0[9] ), .ZN(\SB1_3_31/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 U2993 ( .I(\SB2_1_15/buf_output[0] ), .Z(\RI5[1][126] ) );
  AND2_X1 U2996 ( .A1(\RI3[0][66] ), .A2(\RI3[0][67] ), .Z(n1212) );
  NAND3_X2 U3000 ( .A1(\SB2_2_14/i0_3 ), .A2(\SB2_2_14/i0[8] ), .A3(
        \SB2_2_14/i0[9] ), .ZN(n826) );
  NAND3_X1 U3004 ( .A1(\SB1_3_20/i0_4 ), .A2(\SB1_3_20/i1_7 ), .A3(
        \SB1_3_20/i0[8] ), .ZN(n828) );
  BUF_X4 U3008 ( .I(\SB2_0_18/buf_output[2] ), .Z(\RI5[0][98] ) );
  XOR2_X1 U3016 ( .A1(\RI5[1][50] ), .A2(\RI5[1][56] ), .Z(n1132) );
  XOR2_X1 U3018 ( .A1(\RI5[1][104] ), .A2(\RI5[1][98] ), .Z(
        \MC_ARK_ARC_1_1/temp1[104] ) );
  BUF_X4 U3028 ( .I(\SB2_0_23/buf_output[3] ), .Z(\RI5[0][63] ) );
  INV_X2 U3034 ( .I(\SB1_3_29/buf_output[3] ), .ZN(\SB2_3_27/i0[8] ) );
  NAND3_X1 U3042 ( .A1(\SB1_0_25/i0_3 ), .A2(\SB1_0_25/i0[10] ), .A3(
        \SB1_0_25/i0_4 ), .ZN(n842) );
  XOR2_X1 U3052 ( .A1(n2016), .A2(n847), .Z(n2495) );
  XOR2_X1 U3053 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[186] ), .A2(\RI5[1][0] ), 
        .Z(n847) );
  XOR2_X1 U3073 ( .A1(\MC_ARK_ARC_1_2/temp1[77] ), .A2(n855), .Z(
        \MC_ARK_ARC_1_2/temp5[77] ) );
  XOR2_X1 U3074 ( .A1(\RI5[2][23] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[47] ), 
        .Z(n855) );
  NAND3_X1 U3076 ( .A1(n2774), .A2(\SB2_0_19/i0_3 ), .A3(\SB2_0_19/i0[9] ), 
        .ZN(\SB2_0_19/Component_Function_4/NAND4_in[2] ) );
  XOR2_X1 U3081 ( .A1(\MC_ARK_ARC_1_0/temp1[137] ), .A2(n860), .Z(
        \MC_ARK_ARC_1_0/temp5[137] ) );
  XOR2_X1 U3082 ( .A1(\RI5[0][83] ), .A2(\RI5[0][107] ), .Z(n860) );
  NAND4_X2 U3085 ( .A1(\SB2_1_15/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_1_15/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_1_15/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_15/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_1_15/buf_output[0] ) );
  XOR2_X1 U3102 ( .A1(n868), .A2(\MC_ARK_ARC_1_0/temp6[115] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[115] ) );
  XOR2_X1 U3103 ( .A1(\MC_ARK_ARC_1_0/temp1[115] ), .A2(
        \MC_ARK_ARC_1_0/temp2[115] ), .Z(n868) );
  NAND3_X2 U3107 ( .A1(\SB3_30/i0_3 ), .A2(\SB3_30/i1[9] ), .A3(\SB3_30/i0_4 ), 
        .ZN(n2867) );
  NAND3_X1 U3108 ( .A1(\SB4_20/i0[10] ), .A2(\SB4_20/i1_7 ), .A3(
        \SB4_20/i1[9] ), .ZN(\SB4_20/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U3114 ( .A1(\SB1_1_16/i0_3 ), .A2(\SB1_1_16/i0[8] ), .A3(
        \SB1_1_16/i1_7 ), .ZN(\SB1_1_16/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U3123 ( .A1(\SB4_15/i0_0 ), .A2(\SB4_15/i0[9] ), .A3(\SB4_15/i0[8] ), .ZN(n873) );
  NAND3_X1 U3125 ( .A1(\SB1_2_4/i0_3 ), .A2(\SB1_2_4/i0[8] ), .A3(
        \SB1_2_4/i1_7 ), .ZN(\SB1_2_4/Component_Function_1/NAND4_in[1] ) );
  NAND3_X2 U3126 ( .A1(\SB1_1_0/i0_3 ), .A2(\SB1_1_0/i0_0 ), .A3(
        \SB1_1_0/i0_4 ), .ZN(\SB1_1_0/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3129 ( .A1(\SB1_1_19/i0_3 ), .A2(\SB1_1_19/i0[10] ), .A3(
        \SB1_1_19/i0_4 ), .ZN(\SB1_1_19/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 U3132 ( .A1(\SB2_2_14/i0_3 ), .A2(\SB2_2_14/i1[9] ), .A3(
        \SB2_2_14/i0[6] ), .ZN(\SB2_2_14/Component_Function_3/NAND4_in[0] ) );
  NAND2_X2 U3134 ( .A1(\SB4_18/i0_0 ), .A2(\SB4_18/i3[0] ), .ZN(n876) );
  XOR2_X1 U3136 ( .A1(\RI5[2][123] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[117] ), 
        .Z(n877) );
  XOR2_X1 U3139 ( .A1(\RI5[0][177] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[141] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[75] ) );
  XOR2_X1 U3146 ( .A1(\MC_ARK_ARC_1_1/temp1[171] ), .A2(
        \MC_ARK_ARC_1_1/temp2[171] ), .Z(\MC_ARK_ARC_1_1/temp5[171] ) );
  XOR2_X1 U3156 ( .A1(n884), .A2(\MC_ARK_ARC_1_1/temp2[41] ), .Z(
        \MC_ARK_ARC_1_1/temp5[41] ) );
  XOR2_X1 U3157 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[35] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[41] ), .Z(n884) );
  BUF_X4 U3160 ( .I(\SB2_0_23/buf_output[2] ), .Z(\RI5[0][68] ) );
  NAND3_X1 U3161 ( .A1(\SB1_3_16/i0_0 ), .A2(\SB1_3_16/i1_7 ), .A3(
        \SB1_3_16/i3[0] ), .ZN(n886) );
  NAND4_X2 U3175 ( .A1(\SB2_0_11/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_0_11/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_0_11/Component_Function_1/NAND4_in[2] ), .A4(n1003), .ZN(
        \SB2_0_11/buf_output[1] ) );
  XOR2_X1 U3178 ( .A1(n893), .A2(\MC_ARK_ARC_1_1/temp6[29] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[29] ) );
  XOR2_X1 U3179 ( .A1(\MC_ARK_ARC_1_1/temp2[29] ), .A2(
        \MC_ARK_ARC_1_1/temp1[29] ), .Z(n893) );
  BUF_X4 U3180 ( .I(\SB2_1_29/buf_output[1] ), .Z(\RI5[1][37] ) );
  XOR2_X1 U3183 ( .A1(n894), .A2(\MC_ARK_ARC_1_2/temp6[166] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[166] ) );
  XOR2_X1 U3192 ( .A1(n899), .A2(\MC_ARK_ARC_1_3/temp2[142] ), .Z(
        \MC_ARK_ARC_1_3/temp5[142] ) );
  XOR2_X1 U3193 ( .A1(\RI5[3][136] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[142] ), 
        .Z(n899) );
  NAND4_X2 U3198 ( .A1(\SB2_0_24/Component_Function_1/NAND4_in[3] ), .A2(n1688), .A3(\SB2_0_24/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_24/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_0_24/buf_output[1] ) );
  XOR2_X1 U3203 ( .A1(\MC_ARK_ARC_1_2/temp1[165] ), .A2(
        \MC_ARK_ARC_1_2/temp2[165] ), .Z(\MC_ARK_ARC_1_2/temp5[165] ) );
  NAND4_X2 U3205 ( .A1(\SB2_0_15/Component_Function_0/NAND4_in[3] ), .A2(n2329), .A3(\SB2_0_15/Component_Function_0/NAND4_in[0] ), .A4(n904), .ZN(
        \SB2_0_15/buf_output[0] ) );
  BUF_X4 U3207 ( .I(\SB2_1_25/buf_output[2] ), .Z(\RI5[1][56] ) );
  NAND3_X1 U3208 ( .A1(\SB1_3_16/i0[9] ), .A2(\SB1_3_16/i0_3 ), .A3(
        \SB1_3_16/i0[10] ), .ZN(n905) );
  BUF_X4 U3215 ( .I(\SB2_1_10/buf_output[0] ), .Z(\RI5[1][156] ) );
  NAND3_X2 U3216 ( .A1(\SB2_1_21/i0_3 ), .A2(\RI3[1][60] ), .A3(
        \SB2_1_21/i0[8] ), .ZN(\SB2_1_21/Component_Function_2/NAND4_in[2] ) );
  XOR2_X1 U3221 ( .A1(\MC_ARK_ARC_1_0/temp4[19] ), .A2(
        \MC_ARK_ARC_1_0/temp3[19] ), .Z(\MC_ARK_ARC_1_0/temp6[19] ) );
  NAND4_X2 U3222 ( .A1(\SB1_1_11/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_1_11/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_11/Component_Function_1/NAND4_in[0] ), .A4(n909), .ZN(
        \SB1_1_11/buf_output[1] ) );
  NAND3_X1 U3229 ( .A1(\SB1_1_13/i0[10] ), .A2(\SB1_1_13/i1[9] ), .A3(
        \SB1_1_13/i1_5 ), .ZN(\SB1_1_13/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U3233 ( .A1(\RI5[3][47] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[53] ), 
        .Z(n914) );
  XOR2_X1 U3234 ( .A1(\MC_ARK_ARC_1_3/temp6[118] ), .A2(
        \MC_ARK_ARC_1_3/temp5[118] ), .Z(\MC_ARK_ARC_1_3/buf_output[118] ) );
  XOR2_X1 U3239 ( .A1(\RI5[1][174] ), .A2(\RI5[1][18] ), .Z(
        \MC_ARK_ARC_1_1/temp3[108] ) );
  BUF_X4 U3240 ( .I(\SB2_3_15/buf_output[0] ), .Z(\RI5[3][126] ) );
  NAND4_X2 U3244 ( .A1(\SB2_3_30/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_3_30/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_3_30/Component_Function_3/NAND4_in[3] ), .A4(n918), .ZN(
        \SB2_3_30/buf_output[3] ) );
  XOR2_X1 U3261 ( .A1(\MC_ARK_ARC_1_0/temp2[103] ), .A2(n923), .Z(
        \MC_ARK_ARC_1_0/temp5[103] ) );
  XOR2_X1 U3262 ( .A1(\RI5[0][97] ), .A2(\RI5[0][103] ), .Z(n923) );
  XOR2_X1 U3265 ( .A1(\RI5[1][113] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[89] ), 
        .Z(n926) );
  NAND3_X1 U3266 ( .A1(\SB4_9/i0_4 ), .A2(\SB4_9/i1_5 ), .A3(\SB4_9/i0_0 ), 
        .ZN(n927) );
  INV_X4 U3278 ( .I(n930), .ZN(\RI5[3][8] ) );
  NAND3_X1 U3279 ( .A1(\SB1_0_12/i0[10] ), .A2(\SB1_0_12/i0_0 ), .A3(
        \SB1_0_12/i0[6] ), .ZN(\SB1_0_12/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U3282 ( .A1(\SB2_1_21/i0_4 ), .A2(\SB2_1_21/i0_3 ), .A3(
        \SB2_1_21/i1[9] ), .ZN(\SB2_1_21/Component_Function_5/NAND4_in[2] ) );
  INV_X2 U3286 ( .I(\SB1_1_10/buf_output[3] ), .ZN(\SB2_1_8/i0[8] ) );
  NAND3_X2 U3289 ( .A1(\SB2_1_1/i0_3 ), .A2(\SB2_1_1/i0_4 ), .A3(
        \SB2_1_1/i1[9] ), .ZN(n2449) );
  NAND4_X2 U3290 ( .A1(\SB1_2_0/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_0/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_0/Component_Function_0/NAND4_in[0] ), .A4(n935), .ZN(
        \SB1_2_0/buf_output[0] ) );
  NAND3_X2 U3291 ( .A1(\SB1_2_0/i0_0 ), .A2(\SB1_2_0/i0_3 ), .A3(
        \SB1_2_0/i0[7] ), .ZN(n935) );
  BUF_X4 U3292 ( .I(\SB2_2_19/buf_output[3] ), .Z(\RI5[2][87] ) );
  XOR2_X1 U3295 ( .A1(n937), .A2(\MC_ARK_ARC_1_2/temp3[129] ), .Z(n2761) );
  XOR2_X1 U3296 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[99] ), .A2(\RI5[2][75] ), 
        .Z(n937) );
  BUF_X4 U3299 ( .I(\SB2_3_14/buf_output[3] ), .Z(\RI5[3][117] ) );
  NAND4_X2 U3302 ( .A1(\SB1_2_12/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_2_12/Component_Function_1/NAND4_in[0] ), .A3(
        \SB1_2_12/Component_Function_1/NAND4_in[1] ), .A4(n940), .ZN(
        \SB1_2_12/buf_output[1] ) );
  INV_X2 U3305 ( .I(\SB1_1_30/buf_output[2] ), .ZN(\SB2_1_27/i1[9] ) );
  NAND4_X2 U3310 ( .A1(\SB2_0_27/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_27/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_0_27/Component_Function_4/NAND4_in[1] ), .A4(n943), .ZN(
        \SB2_0_27/buf_output[4] ) );
  NAND3_X1 U3312 ( .A1(\SB2_3_31/i0_3 ), .A2(\SB2_3_31/i0_4 ), .A3(
        \SB2_3_31/i0[10] ), .ZN(\SB2_3_31/Component_Function_0/NAND4_in[2] )
         );
  NAND4_X2 U3315 ( .A1(\SB1_2_8/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_2_8/Component_Function_0/NAND4_in[2] ), .A3(n1813), .A4(
        \SB1_2_8/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_2_8/buf_output[0] ) );
  INV_X4 U3318 ( .I(n1117), .ZN(\SB2_1_13/i1_5 ) );
  NAND3_X1 U3320 ( .A1(\SB3_22/i0_4 ), .A2(\SB3_22/i1_7 ), .A3(\SB3_22/i0[8] ), 
        .ZN(n947) );
  BUF_X4 U3324 ( .I(\SB2_3_31/buf_output[1] ), .Z(\RI5[3][25] ) );
  BUF_X4 U3328 ( .I(\SB2_1_27/buf_output[1] ), .Z(\RI5[1][49] ) );
  NAND3_X2 U3331 ( .A1(\SB2_2_14/i0[10] ), .A2(\SB2_2_14/i0_0 ), .A3(
        \SB2_2_14/i0[6] ), .ZN(\SB2_2_14/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U3332 ( .A1(\MC_ARK_ARC_1_1/temp6[103] ), .A2(n951), .Z(
        \MC_ARK_ARC_1_1/buf_output[103] ) );
  XOR2_X1 U3333 ( .A1(\MC_ARK_ARC_1_1/temp2[103] ), .A2(
        \MC_ARK_ARC_1_1/temp1[103] ), .Z(n951) );
  NAND4_X2 U3334 ( .A1(\SB1_2_20/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_2_20/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_2_20/Component_Function_1/NAND4_in[0] ), .A4(n952), .ZN(
        \SB1_2_20/buf_output[1] ) );
  XOR2_X1 U3339 ( .A1(n1678), .A2(n1116), .Z(\MC_ARK_ARC_1_1/buf_output[187] )
         );
  NAND3_X2 U3349 ( .A1(\SB2_0_13/i0[6] ), .A2(\SB2_0_13/i0[10] ), .A3(
        \SB2_0_13/i0_0 ), .ZN(n957) );
  NAND3_X1 U3355 ( .A1(\SB3_16/i0_3 ), .A2(\SB3_16/i1_7 ), .A3(\SB3_16/i0[8] ), 
        .ZN(n959) );
  XOR2_X1 U3357 ( .A1(\RI5[3][65] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[71] ), 
        .Z(n960) );
  NAND3_X1 U3361 ( .A1(\SB3_0/i1_7 ), .A2(\SB3_0/i0_4 ), .A3(\SB3_0/i0[8] ), 
        .ZN(n962) );
  NAND4_X2 U3364 ( .A1(\SB2_2_23/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_2_23/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_2_23/Component_Function_1/NAND4_in[1] ), .A4(n964), .ZN(
        \SB2_2_23/buf_output[1] ) );
  NAND3_X1 U3366 ( .A1(\SB4_12/i0[6] ), .A2(\SB4_12/i0_3 ), .A3(\SB4_12/i1[9] ), .ZN(n965) );
  INV_X2 U3377 ( .I(\SB1_2_6/buf_output[3] ), .ZN(\SB2_2_4/i0[8] ) );
  INV_X2 U3381 ( .I(n428), .ZN(\SB1_0_8/i1_5 ) );
  XOR2_X1 U3393 ( .A1(n1987), .A2(\MC_ARK_ARC_1_2/temp6[7] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[7] ) );
  BUF_X4 U3400 ( .I(\SB2_3_0/buf_output[0] ), .Z(\RI5[3][24] ) );
  INV_X2 U3411 ( .I(\SB1_2_16/buf_output[2] ), .ZN(\SB2_2_13/i1[9] ) );
  XOR2_X1 U3412 ( .A1(\RI5[3][75] ), .A2(\RI5[3][99] ), .Z(n1693) );
  NAND3_X2 U3422 ( .A1(\SB2_1_17/i0[9] ), .A2(\SB2_1_17/i0_3 ), .A3(
        \SB2_1_17/i0[8] ), .ZN(\SB2_1_17/Component_Function_2/NAND4_in[2] ) );
  XOR2_X1 U3423 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[69] ), .A2(\RI5[0][75] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[75] ) );
  XOR2_X1 U3427 ( .A1(\MC_ARK_ARC_1_2/temp6[38] ), .A2(
        \MC_ARK_ARC_1_2/temp5[38] ), .Z(\MC_ARK_ARC_1_2/buf_output[38] ) );
  NAND3_X2 U3429 ( .A1(\SB2_1_14/i0_0 ), .A2(\SB2_1_14/i0_4 ), .A3(
        \SB2_1_14/i1_5 ), .ZN(n1151) );
  XOR2_X1 U3433 ( .A1(\RI5[1][24] ), .A2(\RI5[1][48] ), .Z(
        \MC_ARK_ARC_1_1/temp2[78] ) );
  BUF_X4 U3434 ( .I(\SB2_2_16/buf_output[0] ), .Z(\RI5[2][120] ) );
  NAND3_X2 U3438 ( .A1(\SB2_2_16/i0_4 ), .A2(\SB2_2_16/i1_7 ), .A3(
        \SB2_2_16/i0[8] ), .ZN(n2299) );
  NAND4_X2 U3444 ( .A1(\SB2_1_13/Component_Function_5/NAND4_in[3] ), .A2(
        \SB2_1_13/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_1_13/Component_Function_5/NAND4_in[0] ), .A4(n990), .ZN(
        \SB2_1_13/buf_output[5] ) );
  NAND4_X2 U3463 ( .A1(\SB2_1_1/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_1/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_1/Component_Function_4/NAND4_in[3] ), .A4(n998), .ZN(
        \SB2_1_1/buf_output[4] ) );
  XOR2_X1 U3472 ( .A1(n1002), .A2(n1001), .Z(\MC_ARK_ARC_1_1/temp6[143] ) );
  XOR2_X1 U3473 ( .A1(\RI5[1][53] ), .A2(n197), .Z(n1001) );
  XOR2_X1 U3474 ( .A1(\RI5[1][17] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[179] ), 
        .Z(n1002) );
  NAND4_X2 U3477 ( .A1(\SB1_2_13/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_2_13/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_2_13/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_2_13/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_2_13/buf_output[0] ) );
  XOR2_X1 U3483 ( .A1(\RI5[0][59] ), .A2(\RI5[0][53] ), .Z(n1869) );
  XOR2_X1 U3489 ( .A1(n2434), .A2(n1006), .Z(\MC_ARK_ARC_1_1/temp5[183] ) );
  XOR2_X1 U3490 ( .A1(\RI5[1][183] ), .A2(\RI5[1][177] ), .Z(n1006) );
  XOR2_X1 U3494 ( .A1(\RI5[2][62] ), .A2(\RI5[2][98] ), .Z(
        \MC_ARK_ARC_1_2/temp3[188] ) );
  XOR2_X1 U3497 ( .A1(\MC_ARK_ARC_1_0/temp6[175] ), .A2(
        \MC_ARK_ARC_1_0/temp5[175] ), .Z(\MC_ARK_ARC_1_0/buf_output[175] ) );
  NAND4_X2 U3498 ( .A1(\SB2_1_12/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_12/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_1_12/Component_Function_2/NAND4_in[2] ), .A4(n1009), .ZN(
        \SB2_1_12/buf_output[2] ) );
  NAND4_X2 U3503 ( .A1(\SB2_1_3/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_1_3/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_1_3/Component_Function_3/NAND4_in[3] ), .A4(n1010), .ZN(
        \SB2_1_3/buf_output[3] ) );
  NAND4_X2 U3512 ( .A1(\SB1_0_22/Component_Function_3/NAND4_in[3] ), .A2(
        \SB1_0_22/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_22/Component_Function_3/NAND4_in[0] ), .A4(n1015), .ZN(
        \RI3[0][69] ) );
  XOR2_X1 U3514 ( .A1(\MC_ARK_ARC_1_3/temp1[23] ), .A2(n1016), .Z(
        \MC_ARK_ARC_1_3/temp5[23] ) );
  XOR2_X1 U3515 ( .A1(\RI5[3][161] ), .A2(\RI5[3][185] ), .Z(n1016) );
  XOR2_X1 U3519 ( .A1(n1017), .A2(\MC_ARK_ARC_1_3/temp1[75] ), .Z(
        \MC_ARK_ARC_1_3/temp5[75] ) );
  XOR2_X1 U3520 ( .A1(\RI5[3][21] ), .A2(\RI5[3][45] ), .Z(n1017) );
  NAND4_X2 U3526 ( .A1(\SB3_29/Component_Function_1/NAND4_in[2] ), .A2(
        \SB3_29/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_29/Component_Function_1/NAND4_in[0] ), .A4(n1020), .ZN(
        \SB3_29/buf_output[1] ) );
  NAND3_X1 U3527 ( .A1(\SB3_29/i0_4 ), .A2(\SB3_29/i1_7 ), .A3(\SB3_29/i0[8] ), 
        .ZN(n1020) );
  XOR2_X1 U3537 ( .A1(\MC_ARK_ARC_1_2/temp2[31] ), .A2(n1466), .Z(n1023) );
  XOR2_X1 U3540 ( .A1(\MC_ARK_ARC_1_2/temp4[127] ), .A2(n1025), .Z(n2623) );
  XOR2_X1 U3541 ( .A1(\RI5[2][37] ), .A2(\RI5[2][1] ), .Z(n1025) );
  BUF_X4 U3542 ( .I(\SB2_0_11/buf_output[2] ), .Z(\RI5[0][140] ) );
  INV_X2 U3548 ( .I(\RI3[0][123] ), .ZN(\SB2_0_11/i0[8] ) );
  XOR2_X1 U3553 ( .A1(\MC_ARK_ARC_1_0/temp1[116] ), .A2(n1030), .Z(
        \MC_ARK_ARC_1_0/temp5[116] ) );
  XOR2_X1 U3554 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[86] ), .A2(\RI5[0][62] ), 
        .Z(n1030) );
  BUF_X4 U3559 ( .I(\SB2_1_1/buf_output[1] ), .Z(\RI5[1][13] ) );
  INV_X1 U3560 ( .I(\SB3_3/buf_output[5] ), .ZN(\SB4_3/i1_5 ) );
  NAND3_X1 U3566 ( .A1(\SB4_28/i0[8] ), .A2(\SB4_28/i1_5 ), .A3(\SB4_28/i3[0] ), .ZN(\SB4_28/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U3567 ( .A1(\MC_ARK_ARC_1_3/temp1[172] ), .A2(
        \MC_ARK_ARC_1_3/temp2[172] ), .Z(\MC_ARK_ARC_1_3/temp5[172] ) );
  INV_X1 U3575 ( .I(\SB1_1_28/buf_output[0] ), .ZN(\SB2_1_23/i3[0] ) );
  NAND4_X2 U3576 ( .A1(\SB1_1_28/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_1_28/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_1_28/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_1_28/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_1_28/buf_output[0] ) );
  NAND4_X2 U3578 ( .A1(\SB2_0_11/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_11/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_0_11/Component_Function_2/NAND4_in[1] ), .A4(
        \SB2_0_11/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_0_11/buf_output[2] ) );
  INV_X1 U3585 ( .I(\SB1_3_28/buf_output[1] ), .ZN(\SB2_3_24/i1_7 ) );
  NAND4_X2 U3586 ( .A1(\SB1_3_28/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_3_28/Component_Function_1/NAND4_in[2] ), .A3(n1295), .A4(
        \SB1_3_28/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_3_28/buf_output[1] ) );
  XOR2_X1 U3588 ( .A1(\MC_ARK_ARC_1_2/temp3[91] ), .A2(
        \MC_ARK_ARC_1_2/temp4[91] ), .Z(n1042) );
  BUF_X4 U3589 ( .I(\SB2_3_12/buf_output[3] ), .Z(\RI5[3][129] ) );
  NAND3_X1 U3590 ( .A1(\SB1_0_29/i0[8] ), .A2(\SB1_0_29/i1_5 ), .A3(
        \SB1_0_29/i3[0] ), .ZN(\SB1_0_29/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 U3592 ( .A1(\SB1_2_10/i0[8] ), .A2(\SB1_2_10/i3[0] ), .A3(
        \SB1_2_10/i1_5 ), .ZN(n1043) );
  NAND4_X2 U3596 ( .A1(\SB2_3_8/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_3_8/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_3_8/Component_Function_0/NAND4_in[0] ), .A4(n1046), .ZN(
        \SB2_3_8/buf_output[0] ) );
  NAND3_X1 U3598 ( .A1(\SB2_0_28/i0[6] ), .A2(\SB2_0_28/i0[7] ), .A3(
        \SB2_0_28/i0[8] ), .ZN(\SB2_0_28/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U3605 ( .A1(\RI5[2][104] ), .A2(\RI5[2][110] ), .Z(n1050) );
  BUF_X4 U3608 ( .I(\SB2_1_4/buf_output[4] ), .Z(\RI5[1][172] ) );
  NAND3_X1 U3609 ( .A1(\SB1_0_11/i0_3 ), .A2(\SB1_0_11/i0[9] ), .A3(
        \SB1_0_11/i0[10] ), .ZN(n1052) );
  INV_X2 U3612 ( .I(\MC_ARK_ARC_1_1/buf_output[182] ), .ZN(\SB1_2_1/i1[9] ) );
  XOR2_X1 U3615 ( .A1(\RI5[1][115] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[139] ), 
        .Z(n1054) );
  INV_X2 U3618 ( .I(\RI3[0][146] ), .ZN(\SB2_0_7/i1[9] ) );
  NAND4_X2 U3619 ( .A1(n2121), .A2(\SB1_0_10/Component_Function_2/NAND4_in[0] ), .A3(\SB1_0_10/Component_Function_2/NAND4_in[2] ), .A4(n2431), .ZN(
        \RI3[0][146] ) );
  XOR2_X1 U3627 ( .A1(\RI5[2][103] ), .A2(\RI5[2][139] ), .Z(n1058) );
  XOR2_X1 U3634 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[182] ), .A2(\RI5[2][176] ), 
        .Z(n1061) );
  XOR2_X1 U3636 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[21] ), .A2(\RI5[0][45] ), 
        .Z(n1062) );
  XOR2_X1 U3640 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[185] ), .A2(\RI5[1][161] ), 
        .Z(n1063) );
  NAND2_X1 U3641 ( .A1(\SB1_1_18/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_1_18/Component_Function_0/NAND4_in[3] ), .ZN(n1756) );
  XOR2_X1 U3652 ( .A1(\MC_ARK_ARC_1_2/temp5[154] ), .A2(n1626), .Z(
        \MC_ARK_ARC_1_2/buf_output[154] ) );
  NAND3_X2 U3668 ( .A1(\SB2_3_18/i0_3 ), .A2(\SB2_3_18/i0[9] ), .A3(
        \SB2_3_18/i0[8] ), .ZN(n1590) );
  XOR2_X1 U3672 ( .A1(\MC_ARK_ARC_1_1/temp5[128] ), .A2(n1078), .Z(
        \MC_ARK_ARC_1_1/buf_output[128] ) );
  XOR2_X1 U3673 ( .A1(n1868), .A2(\MC_ARK_ARC_1_1/temp4[128] ), .Z(n1078) );
  XOR2_X1 U3676 ( .A1(n1080), .A2(n2120), .Z(n1450) );
  XOR2_X1 U3677 ( .A1(\RI5[0][126] ), .A2(\RI5[0][120] ), .Z(n1080) );
  XOR2_X1 U3683 ( .A1(n1088), .A2(\MC_ARK_ARC_1_1/temp3[67] ), .Z(n1286) );
  NAND3_X2 U3684 ( .A1(\SB1_1_11/i0[6] ), .A2(\SB1_1_11/i0_4 ), .A3(
        \SB1_1_11/i0[9] ), .ZN(n2624) );
  NAND3_X2 U3689 ( .A1(\SB1_1_13/i0[10] ), .A2(\SB1_1_13/i0[6] ), .A3(
        \SB1_1_13/i0_3 ), .ZN(\SB1_1_13/Component_Function_2/NAND4_in[1] ) );
  XOR2_X1 U3691 ( .A1(n1622), .A2(n1621), .Z(n2453) );
  XOR2_X1 U3694 ( .A1(\MC_ARK_ARC_1_1/temp3[31] ), .A2(
        \MC_ARK_ARC_1_1/temp4[31] ), .Z(\MC_ARK_ARC_1_1/temp6[31] ) );
  XOR2_X1 U3705 ( .A1(\MC_ARK_ARC_1_2/temp2[95] ), .A2(
        \MC_ARK_ARC_1_2/temp1[95] ), .Z(n2309) );
  XOR2_X1 U3708 ( .A1(\RI5[1][61] ), .A2(\RI5[1][67] ), .Z(n1088) );
  NAND3_X2 U3711 ( .A1(\SB1_2_19/i0_0 ), .A2(\SB1_2_19/i0_4 ), .A3(
        \SB1_2_19/i1_5 ), .ZN(\SB1_2_19/Component_Function_2/NAND4_in[3] ) );
  BUF_X4 U3716 ( .I(\SB1_2_16/buf_output[5] ), .Z(\SB2_2_16/i0_3 ) );
  XOR2_X1 U3722 ( .A1(\RI5[0][113] ), .A2(\RI5[0][107] ), .Z(n1095) );
  XOR2_X1 U3723 ( .A1(\MC_ARK_ARC_1_2/temp1[14] ), .A2(n1096), .Z(
        \MC_ARK_ARC_1_2/temp5[14] ) );
  XOR2_X1 U3724 ( .A1(\RI5[2][152] ), .A2(\RI5[2][176] ), .Z(n1096) );
  XOR2_X1 U3734 ( .A1(n1103), .A2(\MC_ARK_ARC_1_0/temp5[58] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[58] ) );
  XOR2_X1 U3735 ( .A1(\MC_ARK_ARC_1_0/temp4[58] ), .A2(
        \MC_ARK_ARC_1_0/temp3[58] ), .Z(n1103) );
  NAND4_X2 U3739 ( .A1(\SB1_0_13/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_0_13/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_0_13/Component_Function_4/NAND4_in[1] ), .A4(n2417), .ZN(
        \RI3[0][118] ) );
  BUF_X4 U3748 ( .I(\SB2_1_19/buf_output[1] ), .Z(\RI5[1][97] ) );
  XOR2_X1 U3760 ( .A1(\RI5[3][32] ), .A2(\RI5[3][8] ), .Z(
        \MC_ARK_ARC_1_3/temp2[62] ) );
  XOR2_X1 U3763 ( .A1(n1114), .A2(\MC_ARK_ARC_1_0/temp4[56] ), .Z(
        \MC_ARK_ARC_1_0/temp6[56] ) );
  BUF_X4 U3767 ( .I(n407), .Z(\SB1_0_29/i0_3 ) );
  BUF_X4 U3768 ( .I(\SB2_1_21/buf_output[1] ), .Z(\RI5[1][85] ) );
  XOR2_X1 U3770 ( .A1(\MC_ARK_ARC_1_1/temp4[187] ), .A2(
        \MC_ARK_ARC_1_1/temp1[187] ), .Z(n1116) );
  XOR2_X1 U3779 ( .A1(\MC_ARK_ARC_1_0/temp3[13] ), .A2(
        \MC_ARK_ARC_1_0/temp4[13] ), .Z(\MC_ARK_ARC_1_0/temp6[13] ) );
  NAND3_X2 U3780 ( .A1(\SB1_1_12/i0[8] ), .A2(\SB1_1_12/i3[0] ), .A3(
        \SB1_1_12/i1_5 ), .ZN(n1120) );
  INV_X2 U3781 ( .I(\SB1_0_22/buf_output[2] ), .ZN(\SB2_0_19/i1[9] ) );
  NAND2_X1 U3783 ( .A1(\SB1_0_21/Component_Function_4/NAND4_in[1] ), .A2(n1214), .ZN(n1213) );
  NAND4_X2 U3784 ( .A1(\SB1_0_15/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_15/Component_Function_4/NAND4_in[3] ), .A3(
        \SB1_0_15/Component_Function_4/NAND4_in[1] ), .A4(n1121), .ZN(
        \SB1_0_15/buf_output[4] ) );
  XOR2_X1 U3790 ( .A1(\SB2_2_20/buf_output[1] ), .A2(\RI5[2][67] ), .Z(
        \MC_ARK_ARC_1_2/temp2[121] ) );
  NAND4_X2 U3791 ( .A1(\SB1_0_26/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_26/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_0_26/Component_Function_0/NAND4_in[1] ), .A4(n1124), .ZN(
        \SB1_0_26/buf_output[0] ) );
  XOR2_X1 U3794 ( .A1(\MC_ARK_ARC_1_0/temp6[5] ), .A2(n1127), .Z(
        \MC_ARK_ARC_1_0/buf_output[5] ) );
  XOR2_X1 U3795 ( .A1(n2043), .A2(\MC_ARK_ARC_1_0/temp1[5] ), .Z(n1127) );
  XOR2_X1 U3798 ( .A1(\RI5[1][30] ), .A2(\RI5[1][54] ), .Z(
        \MC_ARK_ARC_1_1/temp2[84] ) );
  NAND4_X1 U3799 ( .A1(\SB2_1_30/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_1_30/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_1_30/Component_Function_1/NAND4_in[0] ), .A4(n1129), .ZN(
        \SB2_1_30/buf_output[1] ) );
  NAND3_X2 U3801 ( .A1(\SB1_1_28/i0_0 ), .A2(\SB1_1_28/i1_5 ), .A3(
        \SB1_1_28/i0_4 ), .ZN(n1130) );
  NAND4_X2 U3803 ( .A1(\SB1_0_0/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_0/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_0_0/Component_Function_4/NAND4_in[3] ), .A4(n1131), .ZN(
        \SB1_0_0/buf_output[4] ) );
  NAND4_X2 U3805 ( .A1(\SB1_1_3/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_1_3/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_3/Component_Function_0/NAND4_in[0] ), .A4(n1133), .ZN(
        \SB1_1_3/buf_output[0] ) );
  INV_X2 U3806 ( .I(\SB1_2_16/buf_output[5] ), .ZN(\SB2_2_16/i1_5 ) );
  NAND3_X1 U3807 ( .A1(\SB1_2_31/i0[8] ), .A2(\SB1_2_31/i0_4 ), .A3(
        \SB1_2_31/i1_7 ), .ZN(\SB1_2_31/Component_Function_1/NAND4_in[3] ) );
  XOR2_X1 U3810 ( .A1(\MC_ARK_ARC_1_0/temp3[160] ), .A2(
        \MC_ARK_ARC_1_0/temp4[160] ), .Z(n1255) );
  NAND3_X1 U3817 ( .A1(\SB4_20/i0_0 ), .A2(\SB4_20/i0[8] ), .A3(\SB4_20/i0[9] ), .ZN(\SB4_20/Component_Function_4/NAND4_in[0] ) );
  NAND4_X2 U3827 ( .A1(\SB1_1_18/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_18/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_1_18/Component_Function_5/NAND4_in[3] ), .A4(
        \SB1_1_18/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_18/buf_output[5] ) );
  NAND4_X2 U3833 ( .A1(\SB2_0_30/Component_Function_3/NAND4_in[3] ), .A2(
        \SB2_0_30/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_0_30/Component_Function_3/NAND4_in[0] ), .A4(
        \SB2_0_30/Component_Function_3/NAND4_in[1] ), .ZN(
        \SB2_0_30/buf_output[3] ) );
  NAND3_X1 U3842 ( .A1(\SB1_0_8/i0[8] ), .A2(\SB1_0_8/i1_5 ), .A3(
        \SB1_0_8/i3[0] ), .ZN(n1142) );
  NAND3_X1 U3843 ( .A1(\SB2_0_9/i0_3 ), .A2(\SB2_0_9/i0[7] ), .A3(
        \RI3[0][134] ), .ZN(\SB2_0_9/Component_Function_0/NAND4_in[3] ) );
  XOR2_X1 U3851 ( .A1(\MC_ARK_ARC_1_1/temp3[86] ), .A2(
        \MC_ARK_ARC_1_1/temp4[86] ), .Z(n1146) );
  XOR2_X1 U3856 ( .A1(n1148), .A2(\MC_ARK_ARC_1_0/temp6[41] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[41] ) );
  XOR2_X1 U3857 ( .A1(\MC_ARK_ARC_1_0/temp1[41] ), .A2(
        \MC_ARK_ARC_1_0/temp2[41] ), .Z(n1148) );
  NAND4_X2 U3859 ( .A1(\SB3_30/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_30/Component_Function_2/NAND4_in[2] ), .A3(
        \SB3_30/Component_Function_2/NAND4_in[1] ), .A4(n1669), .ZN(
        \SB3_30/buf_output[2] ) );
  NAND2_X1 U3866 ( .A1(n1713), .A2(n2088), .ZN(n1153) );
  XOR2_X1 U3871 ( .A1(n1768), .A2(n1767), .Z(\MC_ARK_ARC_1_0/buf_output[60] )
         );
  NAND3_X1 U3877 ( .A1(\SB2_1_4/i0[6] ), .A2(\SB2_1_4/i0[8] ), .A3(
        \SB2_1_4/i0[7] ), .ZN(\SB2_1_4/Component_Function_0/NAND4_in[1] ) );
  NOR2_X2 U3878 ( .A1(n1158), .A2(n1157), .ZN(\SB2_1_4/i0[7] ) );
  NAND4_X2 U3882 ( .A1(\SB2_1_12/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_1_12/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_12/Component_Function_0/NAND4_in[0] ), .A4(n1159), .ZN(
        \SB2_1_12/buf_output[0] ) );
  NAND3_X1 U3892 ( .A1(\SB4_18/i0[6] ), .A2(n3662), .A3(\SB4_18/i0[7] ), .ZN(
        \SB4_18/Component_Function_0/NAND4_in[1] ) );
  NAND4_X2 U3902 ( .A1(\SB1_0_26/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_26/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_0_26/Component_Function_5/NAND4_in[3] ), .A4(
        \SB1_0_26/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_0_26/buf_output[5] ) );
  NAND4_X2 U3903 ( .A1(\SB1_0_24/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_24/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_24/Component_Function_2/NAND4_in[2] ), .A4(n1167), .ZN(
        \RI3[0][62] ) );
  NAND4_X2 U3906 ( .A1(\SB1_2_12/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_2_12/Component_Function_0/NAND4_in[0] ), .A3(
        \SB1_2_12/Component_Function_0/NAND4_in[3] ), .A4(n1169), .ZN(
        \SB1_2_12/buf_output[0] ) );
  XOR2_X1 U3908 ( .A1(n1171), .A2(\MC_ARK_ARC_1_2/temp6[147] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[147] ) );
  XOR2_X1 U3909 ( .A1(\MC_ARK_ARC_1_2/temp1[147] ), .A2(
        \MC_ARK_ARC_1_2/temp2[147] ), .Z(n1171) );
  BUF_X4 U3910 ( .I(\SB2_2_12/buf_output[5] ), .Z(\RI5[2][119] ) );
  NAND3_X1 U3914 ( .A1(\SB4_0/i0[10] ), .A2(\SB4_0/i1_5 ), .A3(n1386), .ZN(
        n1174) );
  XOR2_X1 U3920 ( .A1(\RI5[1][130] ), .A2(\RI5[1][136] ), .Z(
        \MC_ARK_ARC_1_1/temp1[136] ) );
  BUF_X4 U3921 ( .I(\SB1_1_28/buf_output[5] ), .Z(\SB2_1_28/i0_3 ) );
  XOR2_X1 U3922 ( .A1(\RI5[3][66] ), .A2(\RI5[3][72] ), .Z(
        \MC_ARK_ARC_1_3/temp1[72] ) );
  XOR2_X1 U3923 ( .A1(n1176), .A2(\MC_ARK_ARC_1_1/temp4[105] ), .Z(
        \MC_ARK_ARC_1_1/temp6[105] ) );
  XOR2_X1 U3924 ( .A1(\RI5[1][171] ), .A2(\RI5[1][15] ), .Z(n1176) );
  XOR2_X1 U3926 ( .A1(\RI5[2][9] ), .A2(\RI5[2][165] ), .Z(n1177) );
  NAND2_X1 U3935 ( .A1(\SB1_2_8/Component_Function_4/NAND4_in[0] ), .A2(n1182), 
        .ZN(n2295) );
  NAND3_X1 U3936 ( .A1(\SB1_2_8/i0_0 ), .A2(\SB1_2_8/i3[0] ), .A3(
        \SB1_2_8/i1_7 ), .ZN(n1182) );
  XOR2_X1 U3939 ( .A1(n1184), .A2(n1183), .Z(n2870) );
  XOR2_X1 U3940 ( .A1(\RI5[0][17] ), .A2(n234), .Z(n1183) );
  NAND2_X1 U3950 ( .A1(\SB1_1_6/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_1_6/Component_Function_4/NAND4_in[3] ), .ZN(n1189) );
  NAND3_X1 U3952 ( .A1(\SB1_0_22/i0_4 ), .A2(\SB1_0_22/i0[10] ), .A3(
        \SB1_0_22/i0_3 ), .ZN(\SB1_0_22/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U3956 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[155] ), .A2(\RI5[3][149] ), 
        .Z(n1192) );
  XOR2_X1 U3961 ( .A1(\MC_ARK_ARC_1_0/temp3[123] ), .A2(
        \MC_ARK_ARC_1_0/temp2[123] ), .Z(n1195) );
  XOR2_X1 U3966 ( .A1(\RI5[3][89] ), .A2(\RI5[3][125] ), .Z(
        \MC_ARK_ARC_1_3/temp3[23] ) );
  NAND3_X1 U3967 ( .A1(\SB1_3_21/i0_3 ), .A2(\SB1_3_21/i0[8] ), .A3(
        \SB1_3_21/i1_7 ), .ZN(\SB1_3_21/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U3969 ( .A1(\SB3_13/i0[8] ), .A2(\SB3_13/i1_5 ), .A3(\SB3_13/i3[0] ), .ZN(n1196) );
  NAND3_X2 U3970 ( .A1(\SB1_0_27/i0_0 ), .A2(\SB1_0_27/i0_3 ), .A3(
        \SB1_0_27/i0_4 ), .ZN(\SB1_0_27/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U3981 ( .A1(\SB2_1_13/Component_Function_0/NAND4_in[1] ), .A2(n2018), .A3(\SB2_1_13/Component_Function_0/NAND4_in[0] ), .A4(n2017), .ZN(
        \SB2_1_13/buf_output[0] ) );
  NAND3_X1 U3983 ( .A1(\SB4_11/i0_3 ), .A2(\SB4_11/i0[6] ), .A3(\SB4_11/i1[9] ), .ZN(\SB4_11/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U3985 ( .A1(\SB1_3_9/i0[8] ), .A2(\SB1_3_9/i0[9] ), .A3(
        \SB1_3_9/i0_0 ), .ZN(n1201) );
  XOR2_X1 U3988 ( .A1(n2495), .A2(\MC_ARK_ARC_1_1/temp6[0] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[0] ) );
  NAND3_X2 U4001 ( .A1(\SB1_0_24/i0_4 ), .A2(\SB1_0_24/i0[9] ), .A3(
        \SB1_0_24/i0[6] ), .ZN(n1205) );
  XOR2_X1 U4003 ( .A1(\MC_ARK_ARC_1_3/temp6[70] ), .A2(n1206), .Z(
        \MC_ARK_ARC_1_3/buf_output[70] ) );
  XOR2_X1 U4004 ( .A1(\MC_ARK_ARC_1_3/temp2[70] ), .A2(
        \MC_ARK_ARC_1_3/temp1[70] ), .Z(n1206) );
  NAND3_X2 U4006 ( .A1(\SB2_1_21/i0[6] ), .A2(\SB2_1_21/i0_3 ), .A3(
        \SB2_1_21/i1[9] ), .ZN(n1208) );
  NAND3_X2 U4009 ( .A1(\SB1_3_6/i0_0 ), .A2(\SB1_3_6/i0_4 ), .A3(
        \SB1_3_6/i1_5 ), .ZN(n1210) );
  XOR2_X1 U4020 ( .A1(\RI5[3][173] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[179] ), 
        .Z(n1217) );
  XOR2_X1 U4021 ( .A1(\RI5[2][147] ), .A2(\RI5[2][123] ), .Z(
        \MC_ARK_ARC_1_2/temp2[177] ) );
  NAND3_X1 U4037 ( .A1(\SB1_2_12/i0_4 ), .A2(\SB1_2_12/i1[9] ), .A3(
        \SB1_2_12/i1_5 ), .ZN(\SB1_2_12/Component_Function_4/NAND4_in[3] ) );
  XOR2_X1 U4042 ( .A1(\MC_ARK_ARC_1_1/temp5[118] ), .A2(
        \MC_ARK_ARC_1_1/temp6[118] ), .Z(\MC_ARK_ARC_1_1/buf_output[118] ) );
  XOR2_X1 U4049 ( .A1(n2497), .A2(\MC_ARK_ARC_1_3/temp6[81] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[81] ) );
  NAND3_X1 U4053 ( .A1(\SB4_15/i0_0 ), .A2(\SB4_15/i1_7 ), .A3(\SB4_15/i3[0] ), 
        .ZN(n1235) );
  XOR2_X1 U4054 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[27] ), .A2(\RI5[2][63] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[153] ) );
  BUF_X4 U4055 ( .I(\SB2_1_29/buf_output[3] ), .Z(\RI5[1][27] ) );
  NAND3_X2 U4057 ( .A1(\SB2_1_20/i0[10] ), .A2(\SB2_1_20/i1_7 ), .A3(
        \SB2_1_20/i1[9] ), .ZN(n1236) );
  NAND3_X1 U4067 ( .A1(n400), .A2(\SB1_0_2/i1_7 ), .A3(\SB1_0_2/i0[8] ), .ZN(
        \SB1_0_2/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U4078 ( .A1(\SB1_0_28/i0[8] ), .A2(\SB1_0_28/i1_7 ), .A3(n6314), 
        .ZN(\SB1_0_28/Component_Function_1/NAND4_in[3] ) );
  BUF_X4 U4088 ( .I(\MC_ARK_ARC_1_2/buf_output[113] ), .Z(\SB1_3_13/i0_3 ) );
  NAND3_X1 U4089 ( .A1(\SB2_1_10/i1[9] ), .A2(\SB1_1_11/buf_output[4] ), .A3(
        \SB2_1_10/i1_5 ), .ZN(\SB2_1_10/Component_Function_4/NAND4_in[3] ) );
  XOR2_X1 U4090 ( .A1(\MC_ARK_ARC_1_0/temp4[94] ), .A2(
        \MC_ARK_ARC_1_0/temp3[94] ), .Z(\MC_ARK_ARC_1_0/temp6[94] ) );
  NAND3_X1 U4094 ( .A1(\SB2_2_9/i0_4 ), .A2(\SB2_2_9/i1_7 ), .A3(
        \SB2_2_9/i0[8] ), .ZN(\SB2_2_9/Component_Function_1/NAND4_in[3] ) );
  XOR2_X1 U4097 ( .A1(\MC_ARK_ARC_1_3/temp3[115] ), .A2(
        \MC_ARK_ARC_1_3/temp4[115] ), .Z(n1257) );
  NAND4_X2 U4098 ( .A1(\SB2_1_16/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_1_16/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_1_16/Component_Function_0/NAND4_in[1] ), .A4(
        \SB2_1_16/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_1_16/buf_output[0] ) );
  NOR2_X2 U4102 ( .A1(n1260), .A2(n1259), .ZN(n1394) );
  NAND2_X1 U4103 ( .A1(n1523), .A2(\SB1_2_13/Component_Function_5/NAND4_in[2] ), .ZN(n1260) );
  XOR2_X1 U4104 ( .A1(\MC_ARK_ARC_1_0/temp2[24] ), .A2(n1261), .Z(
        \MC_ARK_ARC_1_0/temp5[24] ) );
  XOR2_X1 U4105 ( .A1(\RI5[0][18] ), .A2(\RI5[0][24] ), .Z(n1261) );
  NAND3_X1 U4112 ( .A1(\SB3_15/i0_3 ), .A2(\SB3_15/i0[10] ), .A3(\SB3_15/i0_4 ), .ZN(n1264) );
  BUF_X4 U4120 ( .I(\SB1_2_17/buf_output[5] ), .Z(\SB2_2_17/i0_3 ) );
  XOR2_X1 U4124 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[125] ), .A2(\RI5[2][89] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[23] ) );
  XOR2_X1 U4129 ( .A1(\MC_ARK_ARC_1_1/temp6[137] ), .A2(
        \MC_ARK_ARC_1_1/temp5[137] ), .Z(\MC_ARK_ARC_1_1/buf_output[137] ) );
  NAND4_X2 U4132 ( .A1(\SB2_0_20/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_0_20/Component_Function_0/NAND4_in[0] ), .A3(
        \SB2_0_20/Component_Function_0/NAND4_in[2] ), .A4(n1270), .ZN(
        \SB2_0_20/buf_output[0] ) );
  XOR2_X1 U4135 ( .A1(\MC_ARK_ARC_1_2/temp2[68] ), .A2(
        \MC_ARK_ARC_1_2/temp4[68] ), .Z(n1272) );
  XOR2_X1 U4139 ( .A1(n2437), .A2(\MC_ARK_ARC_1_3/temp5[171] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[171] ) );
  XOR2_X1 U4140 ( .A1(\MC_ARK_ARC_1_3/temp4[171] ), .A2(
        \MC_ARK_ARC_1_3/temp3[171] ), .Z(n2437) );
  NAND4_X2 U4141 ( .A1(\SB2_1_20/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_1_20/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_1_20/Component_Function_4/NAND4_in[3] ), .A4(n1275), .ZN(
        \SB2_1_20/buf_output[4] ) );
  NAND3_X1 U4144 ( .A1(\SB4_12/i0[8] ), .A2(\SB4_12/i0_3 ), .A3(\SB4_12/i0[9] ), .ZN(\SB4_12/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 U4145 ( .I(\SB2_2_1/buf_output[1] ), .Z(\RI5[2][13] ) );
  XOR2_X1 U4151 ( .A1(n1280), .A2(\MC_ARK_ARC_1_1/temp6[80] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[80] ) );
  BUF_X4 U4153 ( .I(\SB2_1_18/buf_output[1] ), .Z(\RI5[1][103] ) );
  INV_X2 U4158 ( .I(\SB1_1_29/buf_output[2] ), .ZN(\SB2_1_26/i1[9] ) );
  XOR2_X1 U4161 ( .A1(\MC_ARK_ARC_1_2/temp4[112] ), .A2(
        \MC_ARK_ARC_1_2/temp1[112] ), .Z(n1284) );
  XOR2_X1 U4162 ( .A1(n1885), .A2(\MC_ARK_ARC_1_1/temp6[56] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[56] ) );
  XOR2_X1 U4164 ( .A1(n1286), .A2(n1285), .Z(\MC_ARK_ARC_1_1/buf_output[67] )
         );
  XOR2_X1 U4165 ( .A1(n1314), .A2(\MC_ARK_ARC_1_1/temp4[67] ), .Z(n1285) );
  BUF_X4 U4169 ( .I(\SB2_3_31/buf_output[2] ), .Z(\RI5[3][20] ) );
  BUF_X4 U4172 ( .I(\SB2_0_27/buf_output[3] ), .Z(\RI5[0][39] ) );
  NAND3_X1 U4173 ( .A1(\SB1_0_31/i0[8] ), .A2(\SB1_0_31/i1_7 ), .A3(
        \SB1_0_31/i0_4 ), .ZN(\SB1_0_31/Component_Function_1/NAND4_in[3] ) );
  XOR2_X1 U4176 ( .A1(n1290), .A2(\MC_ARK_ARC_1_1/temp1[66] ), .Z(
        \MC_ARK_ARC_1_1/temp5[66] ) );
  INV_X1 U4178 ( .I(\SB1_3_9/buf_output[0] ), .ZN(\SB2_3_4/i3[0] ) );
  NAND4_X2 U4179 ( .A1(\SB1_3_9/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_3_9/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_9/Component_Function_0/NAND4_in[0] ), .A4(
        \SB1_3_9/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_3_9/buf_output[0] ) );
  XOR2_X1 U4183 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[80] ), .A2(\RI5[1][104] ), 
        .Z(n1292) );
  BUF_X4 U4184 ( .I(n424), .Z(\SB1_0_12/i0_3 ) );
  NAND4_X2 U4185 ( .A1(\SB1_2_9/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_2_9/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_2_9/Component_Function_0/NAND4_in[0] ), .A4(n1293), .ZN(
        \SB1_2_9/buf_output[0] ) );
  BUF_X4 U4186 ( .I(\SB2_2_30/buf_output[4] ), .Z(\RI5[2][16] ) );
  XOR2_X1 U4187 ( .A1(\MC_ARK_ARC_1_1/temp1[10] ), .A2(n1294), .Z(
        \MC_ARK_ARC_1_1/temp5[10] ) );
  XOR2_X1 U4188 ( .A1(\RI5[1][148] ), .A2(\RI5[1][172] ), .Z(n1294) );
  XOR2_X1 U4197 ( .A1(n1298), .A2(\MC_ARK_ARC_1_1/temp5[184] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[184] ) );
  XOR2_X1 U4200 ( .A1(\MC_ARK_ARC_1_1/temp2[25] ), .A2(
        \MC_ARK_ARC_1_1/temp1[25] ), .Z(n1299) );
  NAND3_X1 U4216 ( .A1(\SB4_16/i0[10] ), .A2(\SB4_16/i1_5 ), .A3(
        \SB4_16/i1[9] ), .ZN(\SB4_16/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U4220 ( .A1(\SB2_3_6/Component_Function_2/NAND4_in[0] ), .A2(n2004), 
        .A3(\SB2_3_6/Component_Function_2/NAND4_in[1] ), .A4(
        \SB2_3_6/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB2_3_6/buf_output[2] ) );
  XOR2_X1 U4228 ( .A1(\RI5[0][13] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[7] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[13] ) );
  XOR2_X1 U4231 ( .A1(\MC_ARK_ARC_1_0/temp3[28] ), .A2(
        \MC_ARK_ARC_1_0/temp4[28] ), .Z(n1746) );
  XOR2_X1 U4233 ( .A1(n1307), .A2(\MC_ARK_ARC_1_0/temp2[19] ), .Z(
        \MC_ARK_ARC_1_0/temp5[19] ) );
  XOR2_X1 U4238 ( .A1(\RI5[1][112] ), .A2(\RI5[1][136] ), .Z(
        \MC_ARK_ARC_1_1/temp2[166] ) );
  INV_X1 U4240 ( .I(\SB1_3_16/buf_output[1] ), .ZN(\SB2_3_12/i1_7 ) );
  NAND4_X2 U4242 ( .A1(\SB2_1_29/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_1_29/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_29/Component_Function_1/NAND4_in[0] ), .A4(n1632), .ZN(
        \SB2_1_29/buf_output[1] ) );
  NAND3_X2 U4243 ( .A1(\SB2_3_1/i0_3 ), .A2(\SB2_3_1/i0_4 ), .A3(
        \SB2_3_1/i1[9] ), .ZN(\SB2_3_1/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U4244 ( .A1(\SB2_3_18/i0[10] ), .A2(\SB2_3_18/i0_0 ), .A3(
        \SB2_3_18/i0[6] ), .ZN(n1312) );
  NAND4_X2 U4245 ( .A1(\SB2_2_20/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_2_20/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_2_20/Component_Function_0/NAND4_in[3] ), .A4(
        \SB2_2_20/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_2_20/buf_output[0] ) );
  BUF_X4 U4248 ( .I(\MC_ARK_ARC_1_1/buf_output[128] ), .Z(\SB1_2_10/i0_0 ) );
  XOR2_X1 U4249 ( .A1(\RI5[1][37] ), .A2(\RI5[1][13] ), .Z(n1314) );
  XOR2_X1 U4252 ( .A1(\RI5[0][33] ), .A2(\RI5[0][39] ), .Z(n1315) );
  BUF_X4 U4254 ( .I(\SB2_1_18/buf_output[2] ), .Z(\RI5[1][98] ) );
  XOR2_X1 U4257 ( .A1(\RI5[3][19] ), .A2(\RI5[3][187] ), .Z(
        \MC_ARK_ARC_1_3/temp2[49] ) );
  NAND4_X2 U4259 ( .A1(\SB2_3_28/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_3_28/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_28/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_28/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_3_28/buf_output[0] ) );
  NAND3_X1 U4264 ( .A1(n2911), .A2(n577), .A3(\SB2_3_28/i1_5 ), .ZN(n1320) );
  XOR2_X1 U4265 ( .A1(\MC_ARK_ARC_1_3/temp3[184] ), .A2(
        \MC_ARK_ARC_1_3/temp4[184] ), .Z(n1321) );
  NAND3_X1 U4266 ( .A1(\SB4_0/i0[10] ), .A2(\SB4_0/i1_7 ), .A3(n1386), .ZN(
        n1322) );
  BUF_X4 U4267 ( .I(\SB2_3_28/buf_output[5] ), .Z(\RI5[3][23] ) );
  NAND4_X2 U4270 ( .A1(\SB1_1_25/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_25/Component_Function_5/NAND4_in[3] ), .A3(n2789), .A4(n1324), 
        .ZN(\SB1_1_25/buf_output[5] ) );
  XOR2_X1 U4272 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[42] ), .A2(\RI5[1][78] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[168] ) );
  XOR2_X1 U4279 ( .A1(\RI5[1][174] ), .A2(\RI5[1][6] ), .Z(n1327) );
  BUF_X4 U4284 ( .I(\SB2_1_5/buf_output[4] ), .Z(\RI5[1][166] ) );
  NAND3_X2 U4286 ( .A1(\SB1_0_19/i0_4 ), .A2(\SB1_0_19/i0_3 ), .A3(
        \SB1_0_19/i1[9] ), .ZN(n1330) );
  BUF_X4 U4287 ( .I(\SB2_2_9/buf_output[5] ), .Z(\RI5[2][137] ) );
  BUF_X4 U4288 ( .I(\SB2_1_17/buf_output[1] ), .Z(\RI5[1][109] ) );
  XOR2_X1 U4298 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[110] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[104] ), .Z(\MC_ARK_ARC_1_3/temp1[110] )
         );
  INV_X1 U4300 ( .I(\SB1_0_18/buf_output[0] ), .ZN(\SB2_0_13/i3[0] ) );
  NAND4_X2 U4301 ( .A1(\SB1_0_18/Component_Function_0/NAND4_in[1] ), .A2(n2404), .A3(\SB1_0_18/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_18/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_0_18/buf_output[0] ) );
  BUF_X4 U4302 ( .I(\SB1_1_13/buf_output[5] ), .Z(\SB2_1_13/i0_3 ) );
  XOR2_X1 U4304 ( .A1(\SB2_2_24/buf_output[3] ), .A2(n566), .Z(n1334) );
  NAND2_X1 U4309 ( .A1(\SB1_1_26/Component_Function_0/NAND4_in[0] ), .A2(n2742), .ZN(n2616) );
  NAND3_X1 U4310 ( .A1(\SB1_0_21/i0_0 ), .A2(\SB1_0_21/i3[0] ), .A3(
        \SB1_0_21/i1_7 ), .ZN(\SB1_0_21/Component_Function_4/NAND4_in[1] ) );
  NAND3_X2 U4313 ( .A1(\SB2_1_2/i0[10] ), .A2(\SB2_1_2/i0_0 ), .A3(
        \SB2_1_2/i0[6] ), .ZN(n2583) );
  NAND3_X1 U4314 ( .A1(\SB1_0_28/i0_0 ), .A2(\SB1_0_28/i3[0] ), .A3(
        \SB1_0_28/i1_7 ), .ZN(\SB1_0_28/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U4315 ( .A1(\MC_ARK_ARC_1_1/temp5[152] ), .A2(
        \MC_ARK_ARC_1_1/temp6[152] ), .Z(\MC_ARK_ARC_1_1/buf_output[152] ) );
  XOR2_X1 U4322 ( .A1(\MC_ARK_ARC_1_0/temp5[37] ), .A2(n1340), .Z(
        \MC_ARK_ARC_1_0/buf_output[37] ) );
  XOR2_X1 U4323 ( .A1(\MC_ARK_ARC_1_0/temp3[37] ), .A2(
        \MC_ARK_ARC_1_0/temp4[37] ), .Z(n1340) );
  XOR2_X1 U4324 ( .A1(\RI5[1][81] ), .A2(\RI5[1][117] ), .Z(
        \MC_ARK_ARC_1_1/temp3[15] ) );
  NAND4_X2 U4326 ( .A1(\SB1_1_16/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_16/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_16/Component_Function_3/NAND4_in[2] ), .A4(n1342), .ZN(
        \SB1_1_16/buf_output[3] ) );
  XOR2_X1 U4328 ( .A1(\MC_ARK_ARC_1_0/temp6[129] ), .A2(
        \MC_ARK_ARC_1_0/temp5[129] ), .Z(\MC_ARK_ARC_1_0/buf_output[129] ) );
  BUF_X4 U4330 ( .I(\SB2_3_12/buf_output[1] ), .Z(\RI5[3][139] ) );
  XOR2_X1 U4333 ( .A1(\MC_ARK_ARC_1_2/temp5[109] ), .A2(
        \MC_ARK_ARC_1_2/temp6[109] ), .Z(\MC_ARK_ARC_1_2/buf_output[109] ) );
  INV_X2 U4335 ( .I(\MC_ARK_ARC_1_2/buf_output[1] ), .ZN(\SB1_3_31/i1_7 ) );
  INV_X2 U4337 ( .I(\MC_ARK_ARC_1_0/buf_output[3] ), .ZN(\SB1_1_31/i0[8] ) );
  XOR2_X1 U4341 ( .A1(n1345), .A2(\MC_ARK_ARC_1_0/temp6[185] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[185] ) );
  XOR2_X1 U4345 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[49] ), .A2(\RI5[0][55] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[55] ) );
  NAND3_X1 U4347 ( .A1(\SB2_1_10/i0_0 ), .A2(\SB2_1_10/i3[0] ), .A3(
        \SB2_1_10/i1_7 ), .ZN(n1346) );
  XOR2_X1 U4348 ( .A1(\RI5[1][133] ), .A2(\RI5[1][127] ), .Z(
        \MC_ARK_ARC_1_1/temp1[133] ) );
  XOR2_X1 U4349 ( .A1(n1348), .A2(n1347), .Z(\MC_ARK_ARC_1_1/buf_output[136] )
         );
  XOR2_X1 U4351 ( .A1(\MC_ARK_ARC_1_1/temp3[136] ), .A2(
        \MC_ARK_ARC_1_1/temp1[136] ), .Z(n1348) );
  XOR2_X1 U4353 ( .A1(\MC_ARK_ARC_1_2/temp2[19] ), .A2(
        \MC_ARK_ARC_1_2/temp1[19] ), .Z(n1349) );
  NAND3_X2 U4354 ( .A1(\SB2_2_13/i0_3 ), .A2(n580), .A3(\SB2_2_13/i1[9] ), 
        .ZN(\SB2_2_13/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U4358 ( .A1(\SB3_5/i0[9] ), .A2(\SB3_5/i1_5 ), .A3(\SB3_5/i0[6] ), 
        .ZN(\SB3_5/Component_Function_1/NAND4_in[2] ) );
  XOR2_X1 U4362 ( .A1(n1353), .A2(\MC_ARK_ARC_1_0/temp4[18] ), .Z(
        \MC_ARK_ARC_1_0/temp6[18] ) );
  XOR2_X1 U4363 ( .A1(\RI5[0][84] ), .A2(\RI5[0][120] ), .Z(n1353) );
  XOR2_X1 U4367 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[170] ), .A2(\RI5[1][14] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[104] ) );
  INV_X2 U4368 ( .I(\SB1_3_25/buf_output[2] ), .ZN(\SB2_3_22/i1[9] ) );
  INV_X2 U4370 ( .I(\SB1_2_3/buf_output[5] ), .ZN(\SB2_2_3/i1_5 ) );
  NAND4_X2 U4371 ( .A1(\SB1_0_30/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_0_30/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_30/Component_Function_5/NAND4_in[3] ), .A4(n1355), .ZN(
        \SB1_0_30/buf_output[5] ) );
  NAND3_X2 U4372 ( .A1(\SB1_0_30/i0_3 ), .A2(\SB1_0_30/i0_4 ), .A3(
        \SB1_0_30/i1[9] ), .ZN(n1355) );
  XOR2_X1 U4379 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[56] ), .A2(\RI5[0][80] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[110] ) );
  NAND4_X2 U4381 ( .A1(\SB1_0_23/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_23/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_23/Component_Function_3/NAND4_in[3] ), .A4(n1361), .ZN(
        \RI3[0][63] ) );
  NAND3_X2 U4382 ( .A1(\SB1_0_23/i0[10] ), .A2(\SB1_0_23/i1[9] ), .A3(
        \SB1_0_23/i1_7 ), .ZN(n1361) );
  XOR2_X1 U4384 ( .A1(n1362), .A2(\MC_ARK_ARC_1_0/temp6[172] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[172] ) );
  XOR2_X1 U4385 ( .A1(\MC_ARK_ARC_1_0/temp1[172] ), .A2(
        \MC_ARK_ARC_1_0/temp2[172] ), .Z(n1362) );
  XOR2_X1 U4389 ( .A1(n2143), .A2(\MC_ARK_ARC_1_3/temp5[181] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[181] ) );
  BUF_X4 U4391 ( .I(\SB3_30/buf_output[5] ), .Z(\SB4_30/i0_3 ) );
  BUF_X4 U4399 ( .I(\SB2_1_25/buf_output[1] ), .Z(\RI5[1][61] ) );
  BUF_X4 U4401 ( .I(\SB2_2_13/buf_output[4] ), .Z(\RI5[2][118] ) );
  NAND3_X2 U4402 ( .A1(\SB1_3_11/i0_3 ), .A2(\SB1_3_11/i0_4 ), .A3(
        \SB1_3_11/i1[9] ), .ZN(n2598) );
  BUF_X4 U4404 ( .I(\SB2_3_5/buf_output[3] ), .Z(\RI5[3][171] ) );
  BUF_X4 U4405 ( .I(\SB2_1_9/buf_output[0] ), .Z(\RI5[1][162] ) );
  NAND3_X1 U4413 ( .A1(\SB1_3_26/i0_0 ), .A2(\SB1_3_26/i3[0] ), .A3(
        \SB1_3_26/i1_7 ), .ZN(n2646) );
  NAND3_X1 U4416 ( .A1(\SB3_27/i0[9] ), .A2(\SB3_27/i0[6] ), .A3(\SB3_27/i0_4 ), .ZN(\SB3_27/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U4424 ( .A1(\SB1_3_1/i0[10] ), .A2(\SB1_3_1/i0_0 ), .A3(
        \SB1_3_1/i0[6] ), .ZN(\SB1_3_1/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U4442 ( .A1(\SB2_2_24/i1_7 ), .A2(\SB2_2_24/i0[8] ), .A3(
        \SB2_2_24/i0_4 ), .ZN(\SB2_2_24/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U4443 ( .A1(\SB2_2_24/i1_5 ), .A2(\SB2_2_24/i0[8] ), .A3(
        \SB2_2_24/i3[0] ), .ZN(\SB2_2_24/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U4444 ( .A1(\SB2_2_24/i0_3 ), .A2(\SB2_2_24/i1_7 ), .A3(
        \SB2_2_24/i0[8] ), .ZN(\SB2_2_24/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 U4456 ( .A1(\SB1_1_16/i0_3 ), .A2(\SB1_1_16/i1[9] ), .ZN(
        \SB1_1_16/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U4458 ( .A1(\SB1_1_16/i1[9] ), .A2(\SB1_1_16/i0_3 ), .A3(
        \SB1_1_16/i0[6] ), .ZN(\SB1_1_16/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 U4459 ( .I(\SB2_2_15/buf_output[5] ), .Z(\RI5[2][101] ) );
  NAND3_X1 U4461 ( .A1(\SB1_2_16/i3[0] ), .A2(\SB1_2_16/i0_0 ), .A3(
        \SB1_2_16/i1_7 ), .ZN(\SB1_2_16/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U4463 ( .A1(\SB1_3_12/i1[9] ), .A2(\SB1_3_12/i1_7 ), .A3(
        \SB1_3_12/i0[10] ), .ZN(\SB1_3_12/Component_Function_3/NAND4_in[2] )
         );
  NAND3_X1 U4468 ( .A1(\SB4_11/i0[10] ), .A2(\SB4_11/i0_0 ), .A3(
        \SB4_11/i0[6] ), .ZN(\SB4_11/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U4470 ( .A1(\SB4_11/i0[6] ), .A2(\SB4_11/i0[10] ), .A3(
        \SB4_11/i0_3 ), .ZN(n2635) );
  NAND3_X1 U4471 ( .A1(\SB3_5/i1_5 ), .A2(\SB3_5/i0_0 ), .A3(\SB3_5/i0_4 ), 
        .ZN(\SB3_5/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U4473 ( .A1(n2898), .A2(\SB4_27/i0_3 ), .A3(\SB4_27/i0[7] ), .ZN(
        n2071) );
  NAND2_X1 U4475 ( .A1(\SB4_9/i0[10] ), .A2(\SB4_9/i0[9] ), .ZN(n1913) );
  NAND3_X1 U4483 ( .A1(\SB3_22/i0_0 ), .A2(\SB3_22/i0[6] ), .A3(
        \SB3_22/i0[10] ), .ZN(\SB3_22/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 U4484 ( .I(\SB1_2_6/buf_output[4] ), .Z(\SB2_2_5/i0_4 ) );
  CLKBUF_X4 U4487 ( .I(\MC_ARK_ARC_1_2/buf_output[46] ), .Z(\SB1_3_24/i0_4 )
         );
  CLKBUF_X4 U4488 ( .I(\MC_ARK_ARC_1_3/buf_output[124] ), .Z(\SB3_11/i0_4 ) );
  CLKBUF_X4 U4506 ( .I(\SB1_2_18/buf_output[3] ), .Z(\SB2_2_16/i0[10] ) );
  BUF_X2 U4509 ( .I(\SB3_9/buf_output[2] ), .Z(\SB4_6/i0_0 ) );
  NAND3_X1 U4512 ( .A1(\SB3_7/i1[9] ), .A2(\SB3_7/i0_4 ), .A3(\SB3_7/i0_3 ), 
        .ZN(\SB3_7/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U4525 ( .A1(\SB3_25/i0[9] ), .A2(\SB3_25/i0[6] ), .A3(\SB3_25/i0_4 ), .ZN(\SB3_25/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U4526 ( .A1(\SB3_25/i0[9] ), .A2(\SB3_25/i0[10] ), .A3(
        \SB3_25/i0_3 ), .ZN(\SB3_25/Component_Function_4/NAND4_in[2] ) );
  BUF_X4 U4527 ( .I(\SB2_2_6/buf_output[2] ), .Z(\RI5[2][170] ) );
  INV_X1 U4528 ( .I(\SB3_14/buf_output[1] ), .ZN(\SB4_10/i1_7 ) );
  XOR2_X1 U4529 ( .A1(Key[81]), .A2(Plaintext[81]), .Z(n1367) );
  NAND3_X1 U4535 ( .A1(n2692), .A2(\SB2_3_24/i0_3 ), .A3(\SB2_3_24/i0_0 ), 
        .ZN(\SB2_3_24/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U4541 ( .A1(\SB4_22/i0[10] ), .A2(\SB4_22/i1[9] ), .A3(
        \SB4_22/i1_7 ), .ZN(\SB4_22/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U4542 ( .A1(\SB1_3_22/i0_3 ), .A2(\SB1_3_22/i0_0 ), .A3(
        \SB1_3_22/i0_4 ), .ZN(\SB1_3_22/Component_Function_3/NAND4_in[1] ) );
  CLKBUF_X4 U4543 ( .I(\MC_ARK_ARC_1_2/buf_output[56] ), .Z(\SB1_3_22/i0_0 )
         );
  NAND2_X1 U4548 ( .A1(\SB4_1/i0_3 ), .A2(\SB4_1/i1[9] ), .ZN(
        \SB4_1/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U4549 ( .A1(\SB4_1/i1[9] ), .A2(\SB4_1/i0_4 ), .A3(\SB4_1/i0_3 ), 
        .ZN(\SB4_1/Component_Function_5/NAND4_in[2] ) );
  CLKBUF_X4 U4555 ( .I(\SB3_18/buf_output[3] ), .Z(\SB4_16/i0[10] ) );
  NAND3_X1 U4569 ( .A1(\SB3_24/i0[7] ), .A2(\SB3_24/i0_3 ), .A3(\SB3_24/i0_0 ), 
        .ZN(\SB3_24/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U4573 ( .A1(\SB2_3_6/i0_3 ), .A2(\SB2_3_6/i1_7 ), .A3(
        \SB2_3_6/i0[8] ), .ZN(\SB2_3_6/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U4590 ( .A1(\SB4_26/i0[10] ), .A2(\SB4_26/i0_3 ), .A3(
        \SB4_26/i0[9] ), .ZN(n2372) );
  NAND4_X2 U4592 ( .A1(\SB2_3_19/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_19/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_19/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_19/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_3_19/buf_output[3] ) );
  NAND3_X1 U4596 ( .A1(\SB1_3_23/i0[8] ), .A2(\SB1_3_23/i1_7 ), .A3(
        \SB1_3_23/i0_4 ), .ZN(n2430) );
  NAND3_X1 U4597 ( .A1(\SB3_3/buf_output[2] ), .A2(\SB4_0/i0_3 ), .A3(
        \SB4_0/i0_4 ), .ZN(\SB4_0/Component_Function_3/NAND4_in[1] ) );
  BUF_X2 U4605 ( .I(\MC_ARK_ARC_1_3/buf_output[169] ), .Z(\SB3_3/i0[6] ) );
  INV_X1 U4606 ( .I(\MC_ARK_ARC_1_3/buf_output[169] ), .ZN(\SB3_3/i1_7 ) );
  NAND3_X1 U4610 ( .A1(\SB4_10/i0[10] ), .A2(\SB3_13/buf_output[2] ), .A3(
        \SB4_10/i0[6] ), .ZN(\SB4_10/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U4611 ( .A1(\SB3_13/buf_output[2] ), .A2(\SB4_10/i1_5 ), .A3(
        \SB4_10/i0_4 ), .ZN(n2730) );
  NAND3_X1 U4616 ( .A1(\SB4_16/i0_0 ), .A2(\SB4_16/i0[6] ), .A3(
        \SB4_16/i0[10] ), .ZN(\SB4_16/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 U4620 ( .A1(\SB3_25/i0_0 ), .A2(\SB3_25/i3[0] ), .ZN(
        \SB3_25/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U4621 ( .A1(\SB3_25/i0_0 ), .A2(\SB3_25/i0_3 ), .A3(\SB3_25/i0_4 ), 
        .ZN(\SB3_25/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U4626 ( .A1(\SB3_9/i0[10] ), .A2(\SB3_9/i0_3 ), .A3(\SB3_9/i0[6] ), 
        .ZN(\SB3_9/Component_Function_2/NAND4_in[1] ) );
  NAND4_X2 U4628 ( .A1(n2606), .A2(\SB3_21/Component_Function_5/NAND4_in[0] ), 
        .A3(\SB3_21/Component_Function_5/NAND4_in[1] ), .A4(
        \SB3_21/Component_Function_5/NAND4_in[3] ), .ZN(n1372) );
  NAND3_X1 U4632 ( .A1(\SB4_10/i0_4 ), .A2(n3653), .A3(\SB4_10/i1_5 ), .ZN(
        \SB4_10/Component_Function_4/NAND4_in[3] ) );
  BUF_X4 U4635 ( .I(\SB2_3_17/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[109] ) );
  NAND4_X2 U4636 ( .A1(\SB2_3_17/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_17/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_17/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_3_17/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_3_17/buf_output[1] ) );
  NAND3_X1 U4643 ( .A1(\SB2_3_16/i0[9] ), .A2(\SB2_3_16/i0_0 ), .A3(
        \SB2_3_16/i0[8] ), .ZN(\SB2_3_16/Component_Function_4/NAND4_in[0] ) );
  INV_X1 U4646 ( .I(\SB3_15/buf_output[1] ), .ZN(\SB4_11/i1_7 ) );
  CLKBUF_X4 U4649 ( .I(\MC_ARK_ARC_1_3/buf_output[54] ), .Z(\SB3_22/i0[9] ) );
  CLKBUF_X4 U4650 ( .I(\MC_ARK_ARC_1_3/buf_output[171] ), .Z(\SB3_3/i0[10] )
         );
  NAND3_X1 U4651 ( .A1(\SB1_3_9/i0[10] ), .A2(\SB1_3_9/i0_3 ), .A3(
        \SB1_3_9/i0_4 ), .ZN(\SB1_3_9/Component_Function_0/NAND4_in[2] ) );
  INV_X1 U4663 ( .I(\MC_ARK_ARC_1_2/buf_output[187] ), .ZN(\SB1_3_0/i1_7 ) );
  NAND2_X1 U4665 ( .A1(\SB4_10/i0[10] ), .A2(\SB4_10/i0[9] ), .ZN(
        \SB4_10/Component_Function_0/NAND4_in[0] ) );
  CLKBUF_X4 U4671 ( .I(\SB1_2_12/buf_output[3] ), .Z(\SB2_2_10/i0[10] ) );
  BUF_X4 U4674 ( .I(\MC_ARK_ARC_1_0/buf_output[137] ), .Z(\SB1_1_9/i0_3 ) );
  BUF_X4 U4676 ( .I(\SB2_2_23/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[78] ) );
  NAND3_X1 U4678 ( .A1(\SB4_7/i0_3 ), .A2(\SB4_7/i0[10] ), .A3(\SB4_7/i0[6] ), 
        .ZN(\SB4_7/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U4684 ( .A1(\SB4_19/i0_0 ), .A2(\SB3_20/buf_output[4] ), .A3(
        \SB4_19/i1_5 ), .ZN(n2049) );
  NAND3_X1 U4686 ( .A1(\SB2_1_6/i0_3 ), .A2(\SB2_1_6/i0[8] ), .A3(
        \SB2_1_6/i1_7 ), .ZN(\SB2_1_6/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U4698 ( .A1(Key[187]), .A2(Plaintext[187]), .Z(n1376) );
  INV_X1 U4706 ( .I(\SB3_29/buf_output[1] ), .ZN(\SB4_25/i1_7 ) );
  NAND3_X1 U4713 ( .A1(\SB3_25/i0[10] ), .A2(\SB3_25/i1_5 ), .A3(
        \SB3_25/i1[9] ), .ZN(\SB3_25/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U4714 ( .A1(\SB3_15/i1_7 ), .A2(\SB3_15/i0[8] ), .A3(\SB3_15/i0_4 ), 
        .ZN(\SB3_15/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U4720 ( .A1(\SB2_0_4/i1_5 ), .A2(\SB2_0_4/i0_0 ), .A3(\RI3[0][166] ), .ZN(\SB2_0_4/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U4723 ( .A1(\SB1_0_7/i1_5 ), .A2(\SB1_0_7/i0[10] ), .A3(
        \SB1_0_7/i1[9] ), .ZN(\SB1_0_7/Component_Function_2/NAND4_in[0] ) );
  INV_X1 U4724 ( .I(\MC_ARK_ARC_1_3/buf_output[37] ), .ZN(\SB3_25/i1_7 ) );
  BUF_X2 U4725 ( .I(\SB3_25/buf_output[1] ), .Z(\SB4_21/i0[6] ) );
  CLKBUF_X4 U4728 ( .I(\MC_ARK_ARC_1_3/buf_output[100] ), .Z(\SB3_15/i0_4 ) );
  BUF_X4 U4729 ( .I(\SB2_3_5/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[166] ) );
  NAND3_X1 U4731 ( .A1(\SB1_3_29/i0[9] ), .A2(\SB1_3_29/i0[8] ), .A3(
        \RI1[3][14] ), .ZN(\SB1_3_29/Component_Function_4/NAND4_in[0] ) );
  NAND4_X2 U4739 ( .A1(\SB2_3_16/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_16/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_16/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_16/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_3_16/buf_output[3] ) );
  NAND3_X1 U4741 ( .A1(\SB3_4/i0_0 ), .A2(\SB3_4/i0[6] ), .A3(\SB3_4/i0[10] ), 
        .ZN(\SB3_4/Component_Function_5/NAND4_in[1] ) );
  AND4_X1 U4746 ( .A1(\SB1_1_19/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_19/Component_Function_4/NAND4_in[1] ), .A3(n1495), .A4(n1494), 
        .Z(n1379) );
  NAND4_X2 U4747 ( .A1(\SB2_2_0/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_0/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_2_0/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_2_0/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB2_2_0/buf_output[2] ) );
  NAND3_X1 U4749 ( .A1(\SB2_1_15/i0_3 ), .A2(\SB2_1_15/i0[10] ), .A3(
        \SB2_1_15/i0_4 ), .ZN(\SB2_1_15/Component_Function_0/NAND4_in[2] ) );
  CLKBUF_X4 U4752 ( .I(\MC_ARK_ARC_1_0/buf_output[183] ), .Z(\SB1_1_1/i0[10] )
         );
  NAND2_X1 U4753 ( .A1(\SB4_9/i0_3 ), .A2(\SB4_9/i1[9] ), .ZN(
        \SB4_9/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U4754 ( .A1(\SB3_13/i1_5 ), .A2(\SB3_13/i0_4 ), .A3(\SB3_13/i1[9] ), 
        .ZN(n2600) );
  CLKBUF_X4 U4760 ( .I(\SB1_2_2/buf_output[3] ), .Z(\SB2_2_0/i0[10] ) );
  BUF_X4 U4761 ( .I(\SB2_3_29/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[17] ) );
  BUF_X4 U4768 ( .I(\SB2_3_26/buf_output[5] ), .Z(\RI5[3][35] ) );
  NAND3_X1 U4770 ( .A1(\SB3_20/i0_0 ), .A2(\SB3_20/i1_5 ), .A3(\SB3_20/i0_4 ), 
        .ZN(\SB3_20/Component_Function_2/NAND4_in[3] ) );
  CLKBUF_X4 U4775 ( .I(\SB1_3_20/buf_output[1] ), .Z(\SB2_3_16/i0[6] ) );
  NAND3_X1 U4778 ( .A1(\SB4_22/i0_0 ), .A2(\SB4_22/i0[6] ), .A3(
        \SB4_22/i0[10] ), .ZN(\SB4_22/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 U4783 ( .I(\SB2_3_0/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[14] ) );
  NAND3_X1 U4792 ( .A1(n577), .A2(\SB2_3_28/i1_7 ), .A3(\SB2_3_28/i0[8] ), 
        .ZN(\SB2_3_28/Component_Function_1/NAND4_in[3] ) );
  INV_X1 U4794 ( .I(n358), .ZN(\SB1_0_23/i0[7] ) );
  BUF_X2 U4796 ( .I(\SB3_25/buf_output[3] ), .Z(\SB4_23/i0[10] ) );
  CLKBUF_X4 U4799 ( .I(\MC_ARK_ARC_1_3/buf_output[106] ), .Z(\SB3_14/i0_4 ) );
  NAND3_X1 U4800 ( .A1(\RI1[4][155] ), .A2(\SB3_6/i0[10] ), .A3(\RI1[4][154] ), 
        .ZN(n2527) );
  NAND3_X1 U4802 ( .A1(\SB4_14/i0[9] ), .A2(\SB4_14/i0[10] ), .A3(
        \SB4_14/i0_3 ), .ZN(\SB4_14/Component_Function_4/NAND4_in[2] ) );
  CLKBUF_X4 U4812 ( .I(n1372), .Z(\SB4_21/i0_3 ) );
  NAND3_X1 U4817 ( .A1(\SB4_4/i0[10] ), .A2(\SB4_4/i0_4 ), .A3(\SB4_4/i0_3 ), 
        .ZN(\SB4_4/Component_Function_0/NAND4_in[2] ) );
  CLKBUF_X4 U4818 ( .I(\MC_ARK_ARC_1_0/buf_output[39] ), .Z(\SB1_1_25/i0[10] )
         );
  NAND3_X1 U4819 ( .A1(\SB4_25/i0[10] ), .A2(\SB4_25/i1[9] ), .A3(
        \SB4_25/i1_7 ), .ZN(\SB4_25/Component_Function_3/NAND4_in[2] ) );
  XOR2_X1 U4822 ( .A1(\MC_ARK_ARC_1_3/temp5[171] ), .A2(n2437), .Z(n1385) );
  NAND3_X1 U4827 ( .A1(\SB4_23/i1_5 ), .A2(\SB4_23/i0[10] ), .A3(
        \SB4_23/i1[9] ), .ZN(\SB4_23/Component_Function_2/NAND4_in[0] ) );
  NAND2_X1 U4828 ( .A1(\SB4_23/i0_3 ), .A2(\SB4_23/i1[9] ), .ZN(n1702) );
  CLKBUF_X4 U4835 ( .I(\SB1_0_7/buf_output[3] ), .Z(\SB2_0_5/i0[10] ) );
  NAND3_X1 U4838 ( .A1(\SB2_3_22/i1[9] ), .A2(\SB2_3_22/i1_5 ), .A3(
        \SB2_3_22/i0_4 ), .ZN(\SB2_3_22/Component_Function_4/NAND4_in[3] ) );
  INV_X1 U4846 ( .I(\MC_ARK_ARC_1_3/buf_output[151] ), .ZN(\SB3_6/i1_7 ) );
  NAND3_X1 U4850 ( .A1(\SB2_3_27/i0[10] ), .A2(\SB2_3_27/i0_4 ), .A3(
        \SB2_3_27/i0_3 ), .ZN(\SB2_3_27/Component_Function_0/NAND4_in[2] ) );
  CLKBUF_X4 U4851 ( .I(\MC_ARK_ARC_1_1/buf_output[42] ), .Z(\SB1_2_24/i0[9] )
         );
  NAND3_X2 U4852 ( .A1(\SB1_0_12/i1_5 ), .A2(\SB1_0_12/i0[10] ), .A3(
        \SB1_0_12/i1[9] ), .ZN(\SB1_0_12/Component_Function_2/NAND4_in[0] ) );
  CLKBUF_X4 U4854 ( .I(n259), .Z(\SB1_0_27/i0_0 ) );
  NAND3_X1 U4856 ( .A1(\SB2_0_18/i0_0 ), .A2(\RI3[0][82] ), .A3(
        \SB2_0_18/i1_5 ), .ZN(n1638) );
  NAND3_X1 U4861 ( .A1(\SB1_0_17/i0_0 ), .A2(\SB1_0_17/i0[9] ), .A3(
        \SB1_0_17/i0[8] ), .ZN(n2036) );
  BUF_X2 U4865 ( .I(\SB2_2_2/buf_output[3] ), .Z(n1390) );
  NAND4_X2 U4867 ( .A1(\SB2_2_2/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_2/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_2_2/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_2_2/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_2_2/buf_output[3] ) );
  BUF_X4 U4873 ( .I(\SB2_2_19/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[82] ) );
  AND4_X2 U4874 ( .A1(\SB1_0_15/Component_Function_3/NAND4_in[3] ), .A2(
        \SB1_0_15/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_0_15/Component_Function_3/NAND4_in[1] ), .A4(n2330), .Z(n1393) );
  NAND3_X1 U4877 ( .A1(\SB3_0/i0[9] ), .A2(\SB3_0/i0[6] ), .A3(\SB3_0/i1_5 ), 
        .ZN(\SB3_0/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U4879 ( .A1(\SB3_0/i0[9] ), .A2(\SB3_0/i0_4 ), .A3(\SB3_0/i0[6] ), 
        .ZN(\SB3_0/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U4882 ( .A1(\SB1_1_10/i0[10] ), .A2(\SB1_1_10/i0_0 ), .A3(
        \SB1_1_10/i0[6] ), .ZN(\SB1_1_10/Component_Function_5/NAND4_in[1] ) );
  INV_X1 U4883 ( .I(\MC_ARK_ARC_1_1/buf_output[7] ), .ZN(\SB1_2_30/i1_7 ) );
  BUF_X2 U4884 ( .I(\MC_ARK_ARC_1_1/buf_output[7] ), .Z(\SB1_2_30/i0[6] ) );
  INV_X1 U4885 ( .I(\MC_ARK_ARC_1_0/buf_output[127] ), .ZN(\SB1_1_10/i1_7 ) );
  INV_X1 U4889 ( .I(\RI1[4][41] ), .ZN(\SB3_25/i1_5 ) );
  CLKBUF_X4 U4891 ( .I(\SB3_25/buf_output[5] ), .Z(\SB4_25/i0_3 ) );
  BUF_X4 U4895 ( .I(n415), .Z(\SB1_0_21/i0_3 ) );
  NAND3_X1 U4899 ( .A1(\SB1_0_27/i0_3 ), .A2(\SB1_0_27/i0_0 ), .A3(
        \SB1_0_27/i0[7] ), .ZN(n2273) );
  CLKBUF_X4 U4904 ( .I(\SB1_3_10/buf_output[4] ), .Z(\SB2_3_9/i0_4 ) );
  BUF_X4 U4911 ( .I(\SB2_2_11/buf_output[4] ), .Z(\RI5[2][130] ) );
  CLKBUF_X4 U4914 ( .I(\MC_ARK_ARC_1_0/buf_output[141] ), .Z(\SB1_1_8/i0[10] )
         );
  NAND3_X1 U4923 ( .A1(\SB1_0_14/i0[8] ), .A2(\SB1_0_14/i1_5 ), .A3(
        \SB1_0_14/i3[0] ), .ZN(\SB1_0_14/Component_Function_3/NAND4_in[3] ) );
  CLKBUF_X4 U4926 ( .I(\SB1_1_1/buf_output[2] ), .Z(\SB2_1_30/i0_0 ) );
  NAND3_X1 U4927 ( .A1(\SB2_2_12/i0_3 ), .A2(\SB2_2_12/i0[8] ), .A3(
        \SB2_2_12/i0[9] ), .ZN(\SB2_2_12/Component_Function_2/NAND4_in[2] ) );
  CLKBUF_X4 U4929 ( .I(\MC_ARK_ARC_1_0/buf_output[129] ), .Z(\SB1_1_10/i0[10] ) );
  CLKBUF_X4 U4932 ( .I(\MC_ARK_ARC_1_3/buf_output[32] ), .Z(\SB3_26/i0_0 ) );
  CLKBUF_X4 U4936 ( .I(\MC_ARK_ARC_1_1/buf_output[189] ), .Z(\SB1_2_0/i0[10] )
         );
  BUF_X2 U4937 ( .I(\MC_ARK_ARC_1_3/buf_output[33] ), .Z(\SB3_26/i0[10] ) );
  INV_X1 U4938 ( .I(\MC_ARK_ARC_1_3/buf_output[33] ), .ZN(\SB3_26/i0[8] ) );
  INV_X1 U4939 ( .I(n407), .ZN(\SB1_0_29/i1_5 ) );
  INV_X1 U4944 ( .I(n423), .ZN(\SB1_0_13/i1_5 ) );
  INV_X1 U4945 ( .I(\MC_ARK_ARC_1_3/buf_output[186] ), .ZN(\SB3_0/i3[0] ) );
  INV_X1 U4948 ( .I(\SB1_0_29/buf_output[1] ), .ZN(\SB2_0_25/i1_7 ) );
  BUF_X2 U4949 ( .I(\SB1_0_29/buf_output[1] ), .Z(\RI3[0][37] ) );
  CLKBUF_X4 U4950 ( .I(\RI3[0][116] ), .Z(\SB2_0_12/i0_0 ) );
  OR3_X2 U4951 ( .A1(\SB1_0_27/buf_output[5] ), .A2(\RI3[0][27] ), .A3(
        \SB2_0_27/i0[9] ), .Z(\SB2_0_27/Component_Function_3/NAND4_in[3] ) );
  INV_X1 U4959 ( .I(\MC_ARK_ARC_1_3/buf_output[161] ), .ZN(\SB3_5/i1_5 ) );
  INV_X1 U4961 ( .I(\SB3_10/buf_output[5] ), .ZN(\SB4_10/i1_5 ) );
  INV_X1 U4966 ( .I(\MC_ARK_ARC_1_3/buf_output[173] ), .ZN(\SB3_3/i1_5 ) );
  BUF_X4 U4970 ( .I(\SB2_1_29/buf_output[2] ), .Z(\RI5[1][32] ) );
  XOR2_X1 U4971 ( .A1(\MC_ARK_ARC_1_2/temp4[12] ), .A2(n1404), .Z(n2496) );
  XOR2_X1 U4972 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[78] ), .A2(\RI5[2][114] ), 
        .Z(n1404) );
  XOR2_X1 U4973 ( .A1(n1408), .A2(n1405), .Z(\MC_ARK_ARC_1_1/buf_output[62] )
         );
  XOR2_X1 U4974 ( .A1(\MC_ARK_ARC_1_1/temp2[62] ), .A2(
        \MC_ARK_ARC_1_1/temp1[62] ), .Z(n1405) );
  NAND3_X1 U4975 ( .A1(\SB2_2_15/i0_3 ), .A2(\SB2_2_15/i0[6] ), .A3(
        \SB2_2_15/i1[9] ), .ZN(\SB2_2_15/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U4981 ( .A1(\MC_ARK_ARC_1_1/temp2[72] ), .A2(
        \MC_ARK_ARC_1_1/temp1[72] ), .Z(\MC_ARK_ARC_1_1/temp5[72] ) );
  BUF_X4 U4984 ( .I(\SB2_3_14/buf_output[1] ), .Z(\RI5[3][127] ) );
  NAND3_X1 U4985 ( .A1(\SB1_2_15/i0[6] ), .A2(\SB1_2_15/i0[10] ), .A3(
        \SB1_2_15/i0_3 ), .ZN(\SB1_2_15/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U4986 ( .A1(\SB1_0_7/i0_3 ), .A2(\SB1_0_7/i1[9] ), .A3(
        \SB1_0_7/i0[6] ), .ZN(\SB1_0_7/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U4987 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[34] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[70] ), .Z(\MC_ARK_ARC_1_2/temp3[160] )
         );
  XOR2_X1 U4988 ( .A1(\MC_ARK_ARC_1_1/temp3[62] ), .A2(
        \MC_ARK_ARC_1_1/temp4[62] ), .Z(n1408) );
  XOR2_X1 U4994 ( .A1(n1412), .A2(\MC_ARK_ARC_1_1/temp5[120] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[120] ) );
  XOR2_X1 U4995 ( .A1(\MC_ARK_ARC_1_1/temp3[120] ), .A2(
        \MC_ARK_ARC_1_1/temp4[120] ), .Z(n1412) );
  XOR2_X1 U4996 ( .A1(n1413), .A2(\MC_ARK_ARC_1_1/temp4[27] ), .Z(
        \MC_ARK_ARC_1_1/temp6[27] ) );
  NAND4_X2 U5000 ( .A1(\SB2_1_17/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_1_17/Component_Function_3/NAND4_in[0] ), .A3(n2115), .A4(
        \SB2_1_17/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_1_17/buf_output[3] ) );
  XOR2_X1 U5001 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[79] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[115] ), .Z(\MC_ARK_ARC_1_0/temp3[13] )
         );
  NAND3_X1 U5004 ( .A1(\SB1_0_31/i0_4 ), .A2(\SB1_0_31/i1[9] ), .A3(
        \SB1_0_31/i1_5 ), .ZN(\SB1_0_31/Component_Function_4/NAND4_in[3] ) );
  XOR2_X1 U5005 ( .A1(\RI5[0][63] ), .A2(\RI5[0][27] ), .Z(n1946) );
  XOR2_X1 U5007 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[96] ), .A2(\RI5[0][120] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[150] ) );
  INV_X1 U5008 ( .I(\SB3_19/buf_output[1] ), .ZN(\SB4_15/i1_7 ) );
  NAND4_X2 U5009 ( .A1(\SB3_19/Component_Function_1/NAND4_in[3] ), .A2(
        \SB3_19/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_19/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_19/Component_Function_1/NAND4_in[0] ), .ZN(\SB3_19/buf_output[1] ) );
  XOR2_X1 U5010 ( .A1(\MC_ARK_ARC_1_0/temp5[136] ), .A2(n1417), .Z(
        \MC_ARK_ARC_1_0/buf_output[136] ) );
  XOR2_X1 U5011 ( .A1(\MC_ARK_ARC_1_0/temp4[136] ), .A2(
        \MC_ARK_ARC_1_0/temp3[136] ), .Z(n1417) );
  NAND4_X2 U5016 ( .A1(\SB2_3_5/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_3_5/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_3_5/Component_Function_1/NAND4_in[0] ), .A4(
        \SB2_3_5/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_3_5/buf_output[1] ) );
  BUF_X4 U5017 ( .I(\SB2_3_5/buf_output[1] ), .Z(\RI5[3][181] ) );
  XOR2_X1 U5019 ( .A1(\RI5[1][173] ), .A2(\RI5[1][149] ), .Z(n1419) );
  NAND3_X1 U5021 ( .A1(\SB2_0_5/i0[7] ), .A2(\SB2_0_5/i0[6] ), .A3(
        \SB2_0_5/i0[8] ), .ZN(n1422) );
  XOR2_X1 U5024 ( .A1(\RI5[3][124] ), .A2(\RI5[3][130] ), .Z(
        \MC_ARK_ARC_1_3/temp1[130] ) );
  XOR2_X1 U5026 ( .A1(\MC_ARK_ARC_1_0/temp1[139] ), .A2(
        \MC_ARK_ARC_1_0/temp2[139] ), .Z(n1424) );
  NAND3_X1 U5027 ( .A1(\SB3_27/i0[10] ), .A2(n4764), .A3(\SB3_27/i1_7 ), .ZN(
        \SB3_27/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U5028 ( .A1(\SB4_21/i0[10] ), .A2(\SB4_21/i1_5 ), .A3(n3666), .ZN(
        n1425) );
  NAND4_X2 U5029 ( .A1(\SB1_2_21/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_21/Component_Function_3/NAND4_in[1] ), .A3(n1854), .A4(
        \SB1_2_21/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_2_21/buf_output[3] ) );
  NAND4_X2 U5031 ( .A1(\SB1_2_14/Component_Function_5/NAND4_in[1] ), .A2(n1847), .A3(\SB1_2_14/Component_Function_5/NAND4_in[0] ), .A4(n1427), .ZN(
        \SB1_2_14/buf_output[5] ) );
  XOR2_X1 U5033 ( .A1(\RI5[1][58] ), .A2(\RI5[1][82] ), .Z(
        \MC_ARK_ARC_1_1/temp2[112] ) );
  XOR2_X1 U5038 ( .A1(\RI5[0][74] ), .A2(\RI5[0][80] ), .Z(n1429) );
  BUF_X4 U5041 ( .I(\SB2_1_14/buf_output[4] ), .Z(\RI5[1][112] ) );
  NAND4_X2 U5043 ( .A1(\SB2_2_11/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_2_11/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_2_11/Component_Function_1/NAND4_in[0] ), .A4(n1431), .ZN(
        \SB2_2_11/buf_output[1] ) );
  NAND3_X1 U5044 ( .A1(\SB2_2_4/i0_3 ), .A2(\SB2_2_4/i0[9] ), .A3(
        \SB2_2_4/i0[10] ), .ZN(\SB2_2_4/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U5045 ( .A1(\SB1_2_3/i0[6] ), .A2(\SB1_2_3/i0[8] ), .A3(
        \SB1_2_3/i0[7] ), .ZN(\SB1_2_3/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U5047 ( .A1(\MC_ARK_ARC_1_1/temp4[93] ), .A2(n1433), .Z(n2565) );
  XOR2_X1 U5049 ( .A1(n1434), .A2(n2174), .Z(\MC_ARK_ARC_1_1/buf_output[3] )
         );
  XOR2_X1 U5050 ( .A1(\MC_ARK_ARC_1_1/temp2[3] ), .A2(
        \MC_ARK_ARC_1_1/temp1[3] ), .Z(n1434) );
  XOR2_X1 U5057 ( .A1(\MC_ARK_ARC_1_0/temp6[112] ), .A2(n1437), .Z(
        \MC_ARK_ARC_1_0/buf_output[112] ) );
  XOR2_X1 U5058 ( .A1(\MC_ARK_ARC_1_0/temp2[112] ), .A2(
        \MC_ARK_ARC_1_0/temp1[112] ), .Z(n1437) );
  XOR2_X1 U5060 ( .A1(\RI5[2][168] ), .A2(\RI5[2][174] ), .Z(
        \MC_ARK_ARC_1_2/temp1[174] ) );
  NAND4_X2 U5062 ( .A1(\SB2_0_19/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_0_19/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_0_19/Component_Function_4/NAND4_in[3] ), .A4(
        \SB2_0_19/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB2_0_19/buf_output[4] ) );
  BUF_X4 U5068 ( .I(\SB2_2_0/buf_output[1] ), .Z(\RI5[2][19] ) );
  NAND4_X2 U5071 ( .A1(\SB2_0_28/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_28/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_0_28/Component_Function_2/NAND4_in[2] ), .A4(n1443), .ZN(
        \SB2_0_28/buf_output[2] ) );
  NAND4_X2 U5076 ( .A1(\SB2_0_26/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_26/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_0_26/Component_Function_4/NAND4_in[1] ), .A4(n1447), .ZN(
        \SB2_0_26/buf_output[4] ) );
  NAND3_X2 U5084 ( .A1(\SB2_1_9/i0[10] ), .A2(\SB2_1_9/i0_3 ), .A3(
        \SB2_1_9/i0[6] ), .ZN(n1451) );
  NAND4_X2 U5088 ( .A1(\SB2_0_4/Component_Function_1/NAND4_in[1] ), .A2(n1827), 
        .A3(\SB2_0_4/Component_Function_1/NAND4_in[2] ), .A4(n1454), .ZN(
        \SB2_0_4/buf_output[1] ) );
  XOR2_X1 U5093 ( .A1(\MC_ARK_ARC_1_0/temp2[23] ), .A2(n1458), .Z(
        \MC_ARK_ARC_1_0/temp5[23] ) );
  XOR2_X1 U5094 ( .A1(\RI5[0][17] ), .A2(\RI5[0][23] ), .Z(n1458) );
  NOR2_X2 U5101 ( .A1(n1464), .A2(n1463), .ZN(\SB2_1_10/i0[7] ) );
  XOR2_X1 U5104 ( .A1(n2499), .A2(n2500), .Z(\MC_ARK_ARC_1_0/buf_output[157] )
         );
  XOR2_X1 U5105 ( .A1(\RI5[2][25] ), .A2(\RI5[2][31] ), .Z(n1466) );
  NAND4_X2 U5107 ( .A1(\SB2_3_13/Component_Function_5/NAND4_in[3] ), .A2(n2794), .A3(n2454), .A4(n1467), .ZN(\SB2_3_13/buf_output[5] ) );
  BUF_X4 U5112 ( .I(\SB2_3_2/buf_output[4] ), .Z(\RI5[3][184] ) );
  NAND3_X1 U5114 ( .A1(\SB4_26/i0[10] ), .A2(\SB4_26/i0[6] ), .A3(
        \SB4_26/i0_0 ), .ZN(\SB4_26/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U5118 ( .A1(\SB2_0_2/i0[8] ), .A2(\SB2_0_2/i1_7 ), .A3(
        \SB2_0_2/i0_3 ), .ZN(\SB2_0_2/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U5119 ( .A1(\RI5[3][100] ), .A2(\RI5[3][64] ), .Z(
        \MC_ARK_ARC_1_3/temp3[190] ) );
  NAND4_X2 U5120 ( .A1(\SB2_3_27/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_3_27/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_3_27/Component_Function_0/NAND4_in[3] ), .A4(
        \SB2_3_27/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_3_27/buf_output[0] ) );
  XOR2_X1 U5121 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[70] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[106] ), .Z(\MC_ARK_ARC_1_2/temp3[4] ) );
  XOR2_X1 U5128 ( .A1(n1473), .A2(\MC_ARK_ARC_1_1/temp6[106] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[106] ) );
  XOR2_X1 U5129 ( .A1(\MC_ARK_ARC_1_1/temp2[106] ), .A2(
        \MC_ARK_ARC_1_1/temp1[106] ), .Z(n1473) );
  NAND2_X1 U5137 ( .A1(\SB2_3_26/i0[9] ), .A2(\SB1_3_28/buf_output[3] ), .ZN(
        \SB2_3_26/Component_Function_0/NAND4_in[0] ) );
  XOR2_X1 U5138 ( .A1(\RI5[3][96] ), .A2(\RI5[3][60] ), .Z(
        \MC_ARK_ARC_1_3/temp3[186] ) );
  XOR2_X1 U5139 ( .A1(\MC_ARK_ARC_1_3/temp5[163] ), .A2(n1478), .Z(
        \MC_ARK_ARC_1_3/buf_output[163] ) );
  NAND3_X1 U5141 ( .A1(\SB1_3_31/i0_3 ), .A2(\SB1_3_31/i0[10] ), .A3(
        \SB1_3_31/i0_4 ), .ZN(\SB1_3_31/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 U5145 ( .A1(\SB2_1_2/i0_4 ), .A2(\SB2_1_2/i0_3 ), .A3(
        \SB2_1_2/i0[10] ), .ZN(n1482) );
  INV_X1 U5149 ( .I(\SB3_23/buf_output[1] ), .ZN(\SB4_19/i1_7 ) );
  XOR2_X1 U5153 ( .A1(\MC_ARK_ARC_1_3/temp2[173] ), .A2(n1486), .Z(
        \MC_ARK_ARC_1_3/temp5[173] ) );
  XOR2_X1 U5154 ( .A1(\RI5[3][173] ), .A2(n1365), .Z(n1486) );
  NAND3_X1 U5166 ( .A1(\SB1_3_7/i0[10] ), .A2(\SB1_3_7/i0_3 ), .A3(
        \SB1_3_7/i0_4 ), .ZN(\SB1_3_7/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 U5170 ( .A1(\SB2_1_18/i0_0 ), .A2(\SB2_1_18/i0_4 ), .A3(
        \SB2_1_18/i1_5 ), .ZN(\SB2_1_18/Component_Function_2/NAND4_in[3] ) );
  NAND4_X2 U5171 ( .A1(\SB1_1_19/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_19/Component_Function_4/NAND4_in[1] ), .A3(n1495), .A4(n1494), 
        .ZN(\SB1_1_19/buf_output[4] ) );
  NAND3_X1 U5178 ( .A1(\SB2_2_8/i1[9] ), .A2(\SB2_2_8/i1_5 ), .A3(
        \SB2_2_8/i0_4 ), .ZN(n1831) );
  XOR2_X1 U5179 ( .A1(\MC_ARK_ARC_1_2/temp3[176] ), .A2(
        \MC_ARK_ARC_1_2/temp4[176] ), .Z(n2438) );
  NAND3_X2 U5181 ( .A1(\SB2_1_29/i0[10] ), .A2(\SB2_1_29/i0_0 ), .A3(
        \SB2_1_29/i0[6] ), .ZN(\SB2_1_29/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U5182 ( .A1(n2475), .A2(n1497), .Z(\MC_ARK_ARC_1_3/buf_output[31] )
         );
  XOR2_X1 U5183 ( .A1(\MC_ARK_ARC_1_3/temp4[31] ), .A2(
        \MC_ARK_ARC_1_3/temp3[31] ), .Z(n1497) );
  XOR2_X1 U5189 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[39] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[45] ), .Z(n1500) );
  XOR2_X1 U5190 ( .A1(n1501), .A2(\MC_ARK_ARC_1_3/temp6[8] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[8] ) );
  NAND3_X1 U5199 ( .A1(\SB4_4/i0_4 ), .A2(\SB4_4/i1_7 ), .A3(\SB4_4/i0[8] ), 
        .ZN(n1506) );
  XOR2_X1 U5200 ( .A1(\RI5[3][65] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[101] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[191] ) );
  NAND3_X1 U5210 ( .A1(\SB1_3_25/i0_3 ), .A2(\SB1_3_25/i0_0 ), .A3(
        \SB1_3_25/i0_4 ), .ZN(\SB1_3_25/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U5217 ( .A1(\SB1_1_22/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_22/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_22/Component_Function_3/NAND4_in[3] ), .A4(n1514), .ZN(
        \SB1_1_22/buf_output[3] ) );
  BUF_X4 U5218 ( .I(\SB2_1_20/buf_output[2] ), .Z(\RI5[1][86] ) );
  NAND3_X1 U5223 ( .A1(\SB3_7/i0_0 ), .A2(n4766), .A3(
        \MC_ARK_ARC_1_3/buf_output[148] ), .ZN(
        \SB3_7/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U5225 ( .A1(\SB2_2_7/i0[6] ), .A2(\SB2_2_7/i0[8] ), .A3(
        \SB2_2_7/i0[7] ), .ZN(\SB2_2_7/Component_Function_0/NAND4_in[1] ) );
  NOR2_X2 U5226 ( .A1(n2295), .A2(n2293), .ZN(\SB2_2_7/i0[7] ) );
  NAND3_X1 U5228 ( .A1(\SB4_21/i0[10] ), .A2(\SB4_21/i0[9] ), .A3(
        \SB4_21/i0_3 ), .ZN(n1517) );
  NAND4_X2 U5238 ( .A1(\SB1_0_26/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_0_26/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_0_26/Component_Function_1/NAND4_in[1] ), .A4(
        \SB1_0_26/Component_Function_1/NAND4_in[0] ), .ZN(\RI3[0][55] ) );
  NAND4_X2 U5252 ( .A1(\SB2_1_9/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_1_9/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_9/Component_Function_0/NAND4_in[2] ), .A4(n1528), .ZN(
        \SB2_1_9/buf_output[0] ) );
  XOR2_X1 U5254 ( .A1(\MC_ARK_ARC_1_2/temp2[173] ), .A2(n1529), .Z(
        \MC_ARK_ARC_1_2/temp5[173] ) );
  XOR2_X1 U5255 ( .A1(\RI5[2][167] ), .A2(\RI5[2][173] ), .Z(n1529) );
  NAND4_X2 U5256 ( .A1(\SB1_3_3/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_3_3/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_3_3/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_3_3/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_3_3/buf_output[0] ) );
  XOR2_X1 U5262 ( .A1(\RI5[2][69] ), .A2(\RI5[2][75] ), .Z(n1532) );
  NAND3_X1 U5264 ( .A1(\SB4_6/i0[10] ), .A2(\SB4_6/i1[9] ), .A3(\SB4_6/i1_7 ), 
        .ZN(\SB4_6/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U5265 ( .A1(\RI3[0][37] ), .A2(\SB2_0_25/i0[9] ), .A3(
        \SB2_0_25/i1_5 ), .ZN(\SB2_0_25/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 U5266 ( .A1(\SB1_0_24/Component_Function_4/NAND4_in[2] ), .A2(n2424), .ZN(n2423) );
  XOR2_X1 U5267 ( .A1(\MC_ARK_ARC_1_0/temp6[25] ), .A2(
        \MC_ARK_ARC_1_0/temp5[25] ), .Z(\MC_ARK_ARC_1_0/buf_output[25] ) );
  INV_X2 U5274 ( .I(\RI3[0][67] ), .ZN(\SB2_0_20/i1_7 ) );
  XOR2_X1 U5277 ( .A1(\RI5[1][7] ), .A2(\RI5[1][13] ), .Z(n1536) );
  XOR2_X1 U5279 ( .A1(n1540), .A2(n1539), .Z(n2461) );
  XOR2_X1 U5280 ( .A1(\RI5[3][128] ), .A2(n188), .Z(n1539) );
  XOR2_X1 U5281 ( .A1(\RI5[3][92] ), .A2(\RI5[3][62] ), .Z(n1540) );
  NOR2_X2 U5282 ( .A1(n2123), .A2(n1541), .ZN(n2692) );
  NAND2_X1 U5283 ( .A1(n1704), .A2(\SB1_3_25/Component_Function_4/NAND4_in[3] ), .ZN(n1541) );
  INV_X2 U5286 ( .I(\SB1_1_8/buf_output[3] ), .ZN(\SB2_1_6/i0[8] ) );
  NAND3_X1 U5288 ( .A1(\SB1_0_10/i0_0 ), .A2(\SB1_0_10/i0[9] ), .A3(
        \SB1_0_10/i0[8] ), .ZN(\SB1_0_10/Component_Function_4/NAND4_in[0] ) );
  INV_X2 U5294 ( .I(\SB1_2_24/buf_output[2] ), .ZN(\SB2_2_21/i1[9] ) );
  XOR2_X1 U5303 ( .A1(\RI5[0][113] ), .A2(\RI5[0][77] ), .Z(
        \MC_ARK_ARC_1_0/temp3[11] ) );
  XOR2_X1 U5305 ( .A1(\RI5[1][188] ), .A2(\RI5[1][20] ), .Z(n1551) );
  XOR2_X1 U5307 ( .A1(n1553), .A2(n1595), .Z(\MC_ARK_ARC_1_2/temp5[12] ) );
  XOR2_X1 U5308 ( .A1(\RI5[2][150] ), .A2(\RI5[2][174] ), .Z(n1553) );
  NOR2_X2 U5310 ( .A1(n1557), .A2(n1555), .ZN(n2342) );
  XOR2_X1 U5313 ( .A1(\RI5[0][147] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[141] ), 
        .Z(n2612) );
  INV_X2 U5314 ( .I(\SB1_1_30/buf_output[3] ), .ZN(\SB2_1_28/i0[8] ) );
  NAND4_X2 U5317 ( .A1(\SB1_0_2/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_0_2/Component_Function_3/NAND4_in[2] ), .A3(
        \SB1_0_2/Component_Function_3/NAND4_in[3] ), .A4(
        \SB1_0_2/Component_Function_3/NAND4_in[0] ), .ZN(
        \SB1_0_2/buf_output[3] ) );
  XOR2_X1 U5319 ( .A1(n1383), .A2(\RI5[1][189] ), .Z(
        \MC_ARK_ARC_1_1/temp3[123] ) );
  XOR2_X1 U5325 ( .A1(\RI5[1][117] ), .A2(\RI5[1][111] ), .Z(n1560) );
  NAND4_X2 U5327 ( .A1(\SB2_2_11/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_2_11/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_2_11/Component_Function_4/NAND4_in[1] ), .A4(n1561), .ZN(
        \SB2_2_11/buf_output[4] ) );
  XOR2_X1 U5329 ( .A1(n1563), .A2(\MC_ARK_ARC_1_3/temp2[128] ), .Z(
        \MC_ARK_ARC_1_3/temp5[128] ) );
  XOR2_X1 U5330 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[122] ), .A2(\RI5[3][128] ), 
        .Z(n1563) );
  XOR2_X1 U5343 ( .A1(\RI5[2][171] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[177] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[177] ) );
  XOR2_X1 U5345 ( .A1(\RI5[2][9] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[177] ), 
        .Z(n1571) );
  BUF_X4 U5352 ( .I(\SB2_3_24/buf_output[0] ), .Z(\RI5[3][72] ) );
  NAND3_X2 U5358 ( .A1(\SB2_2_18/i0[6] ), .A2(\SB2_2_18/i1[9] ), .A3(
        \SB2_2_18/i0_3 ), .ZN(\SB2_2_18/Component_Function_3/NAND4_in[0] ) );
  NAND2_X1 U5360 ( .A1(\SB1_1_1/i1[9] ), .A2(\SB1_1_1/i0_3 ), .ZN(
        \SB1_1_1/Component_Function_1/NAND4_in[0] ) );
  NAND4_X2 U5361 ( .A1(\SB3_28/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_28/Component_Function_2/NAND4_in[3] ), .A3(
        \SB3_28/Component_Function_2/NAND4_in[1] ), .A4(
        \SB3_28/Component_Function_2/NAND4_in[2] ), .ZN(\SB3_28/buf_output[2] ) );
  XOR2_X1 U5366 ( .A1(\MC_ARK_ARC_1_3/temp1[168] ), .A2(n1582), .Z(
        \MC_ARK_ARC_1_3/temp5[168] ) );
  XOR2_X1 U5367 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[114] ), .A2(\RI5[3][138] ), 
        .Z(n1582) );
  NAND3_X1 U5373 ( .A1(\SB3_27/i0[8] ), .A2(\SB3_27/i1_5 ), .A3(\SB3_27/i3[0] ), .ZN(n1640) );
  NAND3_X1 U5375 ( .A1(\SB3_10/i0[6] ), .A2(\SB3_10/i0[9] ), .A3(\SB3_10/i1_5 ), .ZN(n2364) );
  NAND3_X1 U5377 ( .A1(\SB2_1_29/i0_0 ), .A2(\SB2_1_29/i3[0] ), .A3(
        \SB2_1_29/i1_7 ), .ZN(\SB2_1_29/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U5383 ( .A1(n1589), .A2(\MC_ARK_ARC_1_2/temp5[52] ), .Z(n2651) );
  XOR2_X1 U5388 ( .A1(n1593), .A2(n70), .Z(Ciphertext[36]) );
  NAND4_X2 U5389 ( .A1(\SB4_25/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_25/Component_Function_0/NAND4_in[1] ), .A3(n2009), .A4(
        \SB4_25/Component_Function_0/NAND4_in[3] ), .ZN(n1593) );
  NAND3_X1 U5391 ( .A1(\SB2_2_3/i0_3 ), .A2(\SB2_2_3/i0[10] ), .A3(
        \SB1_2_4/buf_output[4] ), .ZN(
        \SB2_2_3/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U5392 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[6] ), .A2(\RI5[2][12] ), 
        .Z(n1595) );
  XOR2_X1 U5397 ( .A1(\MC_ARK_ARC_1_2/temp3[40] ), .A2(
        \MC_ARK_ARC_1_2/temp4[40] ), .Z(\MC_ARK_ARC_1_2/temp6[40] ) );
  NAND4_X2 U5398 ( .A1(\SB2_2_20/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_2_20/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_2_20/Component_Function_4/NAND4_in[1] ), .A4(n1598), .ZN(
        \SB2_2_20/buf_output[4] ) );
  NAND4_X2 U5400 ( .A1(\SB2_0_16/Component_Function_3/NAND4_in[3] ), .A2(
        \SB2_0_16/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_0_16/Component_Function_3/NAND4_in[1] ), .A4(n1599), .ZN(
        \SB2_0_16/buf_output[3] ) );
  NAND3_X2 U5401 ( .A1(\SB2_0_16/i0[10] ), .A2(\SB2_0_16/i1[9] ), .A3(
        \SB2_0_16/i1_7 ), .ZN(n1599) );
  INV_X2 U5404 ( .I(\SB1_2_4/buf_output[2] ), .ZN(\SB2_2_1/i1[9] ) );
  XOR2_X1 U5406 ( .A1(\MC_ARK_ARC_1_3/temp6[5] ), .A2(n1601), .Z(\RI1[4][5] )
         );
  NAND3_X2 U5411 ( .A1(\SB1_2_16/i1_5 ), .A2(\SB1_2_16/i0_4 ), .A3(
        \SB1_2_16/i0_0 ), .ZN(n1604) );
  XOR2_X1 U5418 ( .A1(\MC_ARK_ARC_1_3/temp5[169] ), .A2(n1608), .Z(
        \MC_ARK_ARC_1_3/buf_output[169] ) );
  XOR2_X1 U5419 ( .A1(\MC_ARK_ARC_1_3/temp4[169] ), .A2(
        \MC_ARK_ARC_1_3/temp3[169] ), .Z(n1608) );
  NAND4_X2 U5432 ( .A1(n2320), .A2(\SB2_3_27/Component_Function_5/NAND4_in[1] ), .A3(\SB2_3_27/Component_Function_5/NAND4_in[0] ), .A4(n1617), .ZN(
        \SB2_3_27/buf_output[5] ) );
  XOR2_X1 U5433 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[83] ), .A2(\RI5[2][107] ), 
        .Z(n1618) );
  NAND3_X2 U5434 ( .A1(\SB1_1_30/i0[6] ), .A2(\SB1_1_30/i0[9] ), .A3(
        \SB1_1_30/i0_4 ), .ZN(n1619) );
  XOR2_X1 U5437 ( .A1(\RI5[0][187] ), .A2(\RI5[0][31] ), .Z(n1621) );
  XOR2_X1 U5438 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[67] ), .A2(\RI5[0][91] ), 
        .Z(n1622) );
  XOR2_X1 U5444 ( .A1(\MC_ARK_ARC_1_2/temp3[154] ), .A2(
        \MC_ARK_ARC_1_2/temp4[154] ), .Z(n1626) );
  XOR2_X1 U5465 ( .A1(n1636), .A2(\MC_ARK_ARC_1_2/temp1[59] ), .Z(
        \MC_ARK_ARC_1_2/temp5[59] ) );
  XOR2_X1 U5466 ( .A1(\RI5[2][5] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[29] ), 
        .Z(n1636) );
  XOR2_X1 U5467 ( .A1(\MC_ARK_ARC_1_3/temp5[28] ), .A2(n1637), .Z(
        \MC_ARK_ARC_1_3/buf_output[28] ) );
  XOR2_X1 U5468 ( .A1(\MC_ARK_ARC_1_3/temp4[28] ), .A2(
        \MC_ARK_ARC_1_3/temp3[28] ), .Z(n1637) );
  BUF_X4 U5469 ( .I(\SB2_3_22/buf_output[4] ), .Z(\RI5[3][64] ) );
  BUF_X4 U5488 ( .I(\SB2_2_5/buf_output[3] ), .Z(\RI5[2][171] ) );
  XOR2_X1 U5493 ( .A1(\MC_ARK_ARC_1_1/temp4[76] ), .A2(
        \MC_ARK_ARC_1_1/temp3[76] ), .Z(\MC_ARK_ARC_1_1/temp6[76] ) );
  NAND4_X2 U5495 ( .A1(\SB2_1_7/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_1_7/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_1_7/Component_Function_1/NAND4_in[0] ), .A4(n1650), .ZN(
        \SB2_1_7/buf_output[1] ) );
  XOR2_X1 U5497 ( .A1(\MC_ARK_ARC_1_1/temp1[31] ), .A2(n1651), .Z(
        \MC_ARK_ARC_1_1/temp5[31] ) );
  XOR2_X1 U5498 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[169] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[1] ), .Z(n1651) );
  NAND4_X2 U5499 ( .A1(\SB2_3_23/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_3_23/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_3_23/Component_Function_4/NAND4_in[1] ), .A4(n1652), .ZN(
        \SB2_3_23/buf_output[4] ) );
  XOR2_X1 U5502 ( .A1(\MC_ARK_ARC_1_0/temp2[110] ), .A2(
        \MC_ARK_ARC_1_0/temp4[110] ), .Z(n1653) );
  XOR2_X1 U5504 ( .A1(n1656), .A2(n1655), .Z(\MC_ARK_ARC_1_0/buf_output[69] )
         );
  XOR2_X1 U5506 ( .A1(\MC_ARK_ARC_1_0/temp3[69] ), .A2(
        \MC_ARK_ARC_1_0/temp1[69] ), .Z(n1656) );
  NAND3_X1 U5512 ( .A1(\SB4_3/i0[6] ), .A2(n5495), .A3(\SB4_3/i0[7] ), .ZN(
        \SB4_3/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U5515 ( .A1(\RI5[2][42] ), .A2(\RI5[2][66] ), .Z(
        \MC_ARK_ARC_1_2/temp2[96] ) );
  BUF_X4 U5516 ( .I(\SB2_2_5/buf_output[4] ), .Z(\RI5[2][166] ) );
  NAND4_X2 U5517 ( .A1(\SB2_2_29/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_2_29/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_2_29/Component_Function_0/NAND4_in[0] ), .A4(n1662), .ZN(
        \SB2_2_29/buf_output[0] ) );
  XOR2_X1 U5519 ( .A1(\MC_ARK_ARC_1_1/temp2[57] ), .A2(n1664), .Z(
        \MC_ARK_ARC_1_1/temp5[57] ) );
  XOR2_X1 U5520 ( .A1(\RI5[1][51] ), .A2(\RI5[1][57] ), .Z(n1664) );
  BUF_X4 U5530 ( .I(\SB2_0_26/buf_output[1] ), .Z(\RI5[0][55] ) );
  NAND3_X1 U5532 ( .A1(\SB2_0_28/i0_3 ), .A2(\SB2_0_28/i0[10] ), .A3(
        \RI3[0][22] ), .ZN(\SB2_0_28/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U5533 ( .A1(n1673), .A2(n1672), .Z(n1678) );
  XOR2_X1 U5534 ( .A1(\RI5[1][61] ), .A2(\RI5[1][157] ), .Z(n1672) );
  XOR2_X1 U5535 ( .A1(\RI5[1][133] ), .A2(\RI5[1][97] ), .Z(n1673) );
  BUF_X4 U5536 ( .I(\SB2_3_1/buf_output[3] ), .Z(\RI5[3][3] ) );
  XOR2_X1 U5542 ( .A1(\MC_ARK_ARC_1_2/temp6[71] ), .A2(
        \MC_ARK_ARC_1_2/temp5[71] ), .Z(\RI1[3][71] ) );
  XOR2_X1 U5544 ( .A1(\RI5[3][15] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[51] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[141] ) );
  XOR2_X1 U5551 ( .A1(\RI5[2][23] ), .A2(\RI5[2][191] ), .Z(n1743) );
  NAND3_X1 U5552 ( .A1(\SB1_3_21/i0[6] ), .A2(\SB1_3_21/i1[9] ), .A3(
        \SB1_3_21/i0_3 ), .ZN(\SB1_3_21/Component_Function_3/NAND4_in[0] ) );
  NAND4_X2 U5557 ( .A1(\SB2_1_24/Component_Function_5/NAND4_in[1] ), .A2(
        \SB2_1_24/Component_Function_5/NAND4_in[2] ), .A3(
        \SB2_1_24/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_1_24/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_1_24/buf_output[5] ) );
  BUF_X4 U5563 ( .I(\SB2_2_5/buf_output[2] ), .Z(\RI5[2][176] ) );
  NAND4_X2 U5566 ( .A1(\SB2_2_14/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_14/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_14/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_2_14/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_2_14/buf_output[5] ) );
  XOR2_X1 U5568 ( .A1(\RI5[3][129] ), .A2(\RI5[3][153] ), .Z(
        \MC_ARK_ARC_1_3/temp2[183] ) );
  XOR2_X1 U5572 ( .A1(\MC_ARK_ARC_1_0/temp3[35] ), .A2(
        \MC_ARK_ARC_1_0/temp4[35] ), .Z(n1682) );
  XOR2_X1 U5578 ( .A1(n1686), .A2(\MC_ARK_ARC_1_1/temp4[26] ), .Z(n2863) );
  NAND3_X1 U5586 ( .A1(\SB4_23/i0_0 ), .A2(\SB4_23/i0_3 ), .A3(\SB4_23/i0[7] ), 
        .ZN(\SB4_23/Component_Function_0/NAND4_in[3] ) );
  XOR2_X1 U5588 ( .A1(\MC_ARK_ARC_1_3/temp1[129] ), .A2(n1693), .Z(
        \MC_ARK_ARC_1_3/temp5[129] ) );
  INV_X2 U5589 ( .I(\SB1_1_8/buf_output[2] ), .ZN(\SB2_1_5/i1[9] ) );
  XOR2_X1 U5593 ( .A1(\MC_ARK_ARC_1_2/temp3[97] ), .A2(
        \MC_ARK_ARC_1_2/temp4[97] ), .Z(\MC_ARK_ARC_1_2/temp6[97] ) );
  NAND3_X1 U5596 ( .A1(\RI1[2][47] ), .A2(\SB1_2_24/i0[10] ), .A3(
        \SB1_2_24/i0_4 ), .ZN(\SB1_2_24/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U5599 ( .A1(\MC_ARK_ARC_1_3/temp2[113] ), .A2(n4767), .Z(n1699) );
  NAND4_X2 U5601 ( .A1(\SB4_23/Component_Function_1/NAND4_in[2] ), .A2(
        \SB4_23/Component_Function_1/NAND4_in[1] ), .A3(n2632), .A4(n1702), 
        .ZN(n2298) );
  NAND3_X1 U5606 ( .A1(\SB1_2_14/i0_0 ), .A2(\SB1_2_14/i3[0] ), .A3(
        \SB1_2_14/i1_7 ), .ZN(n1706) );
  XOR2_X1 U5612 ( .A1(\MC_ARK_ARC_1_3/temp5[23] ), .A2(n2303), .Z(
        \MC_ARK_ARC_1_3/buf_output[23] ) );
  XOR2_X1 U5615 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[17] ), .A2(\RI5[3][23] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[23] ) );
  NAND4_X2 U5618 ( .A1(\SB2_0_1/Component_Function_5/NAND4_in[1] ), .A2(
        \SB2_0_1/Component_Function_5/NAND4_in[2] ), .A3(
        \SB2_0_1/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_0_1/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_0_1/buf_output[5] ) );
  NAND3_X1 U5621 ( .A1(\SB4_23/i0_4 ), .A2(\SB4_23/i0_3 ), .A3(\SB4_23/i1[9] ), 
        .ZN(\SB4_23/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U5622 ( .A1(\SB2_0_1/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_1/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_0_1/Component_Function_4/NAND4_in[3] ), .A4(
        \SB2_0_1/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB2_0_1/buf_output[4] ) );
  NAND3_X2 U5627 ( .A1(\SB3_15/i0_3 ), .A2(\SB3_15/i1[9] ), .A3(\SB3_15/i0_4 ), 
        .ZN(\SB3_15/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U5634 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[44] ), .A2(\RI5[3][80] ), 
        .Z(n1718) );
  NOR2_X1 U5636 ( .A1(\MC_ARK_ARC_1_1/buf_output[12] ), .A2(
        \MC_ARK_ARC_1_1/buf_output[15] ), .ZN(n1721) );
  NAND3_X1 U5640 ( .A1(\RI3[0][39] ), .A2(\SB2_0_25/i0_3 ), .A3(\RI3[0][40] ), 
        .ZN(n1724) );
  XOR2_X1 U5642 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[46] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[22] ), .Z(\MC_ARK_ARC_1_0/temp2[76] ) );
  NAND3_X2 U5646 ( .A1(\SB2_0_25/i0_0 ), .A2(\RI3[0][39] ), .A3(\RI3[0][37] ), 
        .ZN(\SB2_0_25/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U5648 ( .A1(\MC_ARK_ARC_1_3/temp5[161] ), .A2(n1729), .Z(
        \MC_ARK_ARC_1_3/buf_output[161] ) );
  NAND3_X1 U5658 ( .A1(\SB1_1_25/i0[6] ), .A2(\MC_ARK_ARC_1_0/buf_output[40] ), 
        .A3(\SB1_1_25/i0[9] ), .ZN(\SB1_1_25/Component_Function_5/NAND4_in[3] ) );
  XOR2_X1 U5659 ( .A1(\RI5[1][72] ), .A2(\RI5[1][108] ), .Z(
        \MC_ARK_ARC_1_1/temp3[6] ) );
  NAND3_X1 U5666 ( .A1(\SB1_2_7/i0[8] ), .A2(\SB1_2_7/i0_4 ), .A3(
        \SB1_2_7/i1_7 ), .ZN(n1733) );
  NAND3_X1 U5667 ( .A1(\SB1_3_21/i0[6] ), .A2(\SB1_3_21/i0[9] ), .A3(
        \SB1_3_21/i1_5 ), .ZN(\SB1_3_21/Component_Function_1/NAND4_in[2] ) );
  XOR2_X1 U5670 ( .A1(\MC_ARK_ARC_1_3/temp6[123] ), .A2(
        \MC_ARK_ARC_1_3/temp5[123] ), .Z(\MC_ARK_ARC_1_3/buf_output[123] ) );
  XOR2_X1 U5672 ( .A1(n2087), .A2(n2086), .Z(\MC_ARK_ARC_1_2/buf_output[61] )
         );
  XOR2_X1 U5673 ( .A1(\MC_ARK_ARC_1_1/temp5[6] ), .A2(
        \MC_ARK_ARC_1_1/temp6[6] ), .Z(\MC_ARK_ARC_1_1/buf_output[6] ) );
  XOR2_X1 U5682 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[81] ), .A2(\RI5[2][87] ), 
        .Z(n1736) );
  XOR2_X1 U5683 ( .A1(\MC_ARK_ARC_1_3/temp2[46] ), .A2(n1737), .Z(n2358) );
  XOR2_X1 U5684 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[40] ), .A2(\RI5[3][46] ), 
        .Z(n1737) );
  XOR2_X1 U5685 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[81] ), .A2(\RI5[2][75] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[81] ) );
  NAND3_X1 U5687 ( .A1(\SB4_22/i0[10] ), .A2(\SB4_22/i0_3 ), .A3(
        \SB4_22/i0[6] ), .ZN(\SB4_22/Component_Function_2/NAND4_in[1] ) );
  NAND4_X2 U5689 ( .A1(\SB2_1_28/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_1_28/Component_Function_0/NAND4_in[0] ), .A3(n1740), .A4(n1739), 
        .ZN(\SB2_1_28/buf_output[0] ) );
  NAND4_X2 U5691 ( .A1(\SB1_2_23/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_23/Component_Function_2/NAND4_in[2] ), .A3(
        \SB1_2_23/Component_Function_2/NAND4_in[3] ), .A4(
        \SB1_2_23/Component_Function_2/NAND4_in[1] ), .ZN(
        \SB1_2_23/buf_output[2] ) );
  NAND2_X1 U5692 ( .A1(\SB1_2_28/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_28/Component_Function_4/NAND4_in[2] ), .ZN(n2027) );
  XOR2_X1 U5695 ( .A1(n1743), .A2(\MC_ARK_ARC_1_2/temp1[53] ), .Z(n1834) );
  BUF_X4 U5703 ( .I(\SB2_2_3/buf_output[4] ), .Z(\RI5[2][178] ) );
  NAND3_X2 U5704 ( .A1(\SB2_1_13/i0[10] ), .A2(\SB2_1_13/i1_5 ), .A3(
        \SB2_1_13/i1[9] ), .ZN(\SB2_1_13/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 U5706 ( .I(\SB2_1_8/buf_output[0] ), .Z(\RI5[1][168] ) );
  XOR2_X1 U5709 ( .A1(\RI5[3][33] ), .A2(\RI5[3][57] ), .Z(n1747) );
  NAND3_X1 U5713 ( .A1(\SB2_1_18/i0_3 ), .A2(\SB2_1_18/i0_0 ), .A3(
        \SB2_1_18/i0_4 ), .ZN(\SB2_1_18/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U5715 ( .A1(\SB1_2_21/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_21/Component_Function_4/NAND4_in[3] ), .A3(n1886), .A4(n1751), 
        .ZN(\SB1_2_21/buf_output[4] ) );
  NOR2_X2 U5719 ( .A1(n1756), .A2(n1754), .ZN(n2885) );
  NAND3_X2 U5720 ( .A1(\SB2_2_3/i0[9] ), .A2(\SB1_2_4/buf_output[4] ), .A3(
        \SB2_2_3/i0[6] ), .ZN(n2757) );
  NAND3_X2 U5721 ( .A1(\SB3_17/i0[10] ), .A2(\SB3_17/i0_0 ), .A3(
        \SB3_17/i0[6] ), .ZN(\SB3_17/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U5724 ( .A1(\RI5[0][102] ), .A2(\RI5[0][108] ), .Z(
        \MC_ARK_ARC_1_0/temp1[108] ) );
  NAND4_X2 U5726 ( .A1(n1832), .A2(n1833), .A3(
        \SB1_0_13/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_0_13/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_0_13/buf_output[0] ) );
  NAND3_X1 U5729 ( .A1(\SB2_0_9/i0[7] ), .A2(\SB2_0_9/i0[6] ), .A3(
        \SB2_0_9/i0[8] ), .ZN(\SB2_0_9/Component_Function_0/NAND4_in[1] ) );
  NAND4_X2 U5740 ( .A1(\SB2_3_14/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_3_14/Component_Function_3/NAND4_in[0] ), .A3(n2657), .A4(
        \SB2_3_14/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_3_14/buf_output[3] ) );
  XOR2_X1 U5748 ( .A1(n1764), .A2(n1763), .Z(n2348) );
  XOR2_X1 U5749 ( .A1(\RI5[1][56] ), .A2(n222), .Z(n1763) );
  XOR2_X1 U5750 ( .A1(\SB2_1_30/buf_output[2] ), .A2(\RI5[1][92] ), .Z(n1764)
         );
  INV_X2 U5751 ( .I(\SB1_2_1/buf_output[5] ), .ZN(\SB2_2_1/i1_5 ) );
  XOR2_X1 U5752 ( .A1(\MC_ARK_ARC_1_2/temp1[38] ), .A2(
        \MC_ARK_ARC_1_2/temp2[38] ), .Z(\MC_ARK_ARC_1_2/temp5[38] ) );
  XOR2_X1 U5753 ( .A1(\MC_ARK_ARC_1_3/temp6[103] ), .A2(
        \MC_ARK_ARC_1_3/temp5[103] ), .Z(\MC_ARK_ARC_1_3/buf_output[103] ) );
  NAND3_X1 U5756 ( .A1(n1388), .A2(\SB1_3_10/i0[8] ), .A3(\SB1_3_10/i1_7 ), 
        .ZN(\SB1_3_10/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U5757 ( .A1(\MC_ARK_ARC_1_0/temp2[60] ), .A2(
        \MC_ARK_ARC_1_0/temp4[60] ), .Z(n1767) );
  XOR2_X1 U5758 ( .A1(\MC_ARK_ARC_1_0/temp3[60] ), .A2(
        \MC_ARK_ARC_1_0/temp1[60] ), .Z(n1768) );
  NAND3_X1 U5766 ( .A1(\SB3_14/i0[8] ), .A2(\SB3_14/i3[0] ), .A3(\SB3_14/i1_5 ), .ZN(n1979) );
  NAND3_X1 U5768 ( .A1(\SB3_11/i0_4 ), .A2(\SB3_11/i1[9] ), .A3(n582), .ZN(
        \SB3_11/Component_Function_4/NAND4_in[3] ) );
  INV_X1 U5770 ( .I(\RI3[0][96] ), .ZN(\SB2_0_15/i3[0] ) );
  NAND4_X2 U5771 ( .A1(\SB1_0_20/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_0_20/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_0_20/Component_Function_0/NAND4_in[0] ), .A4(
        \SB1_0_20/Component_Function_0/NAND4_in[2] ), .ZN(\RI3[0][96] ) );
  NAND3_X1 U5774 ( .A1(\SB4_24/i0[6] ), .A2(\SB4_24/i0[10] ), .A3(
        \SB4_24/i0_0 ), .ZN(\SB4_24/Component_Function_5/NAND4_in[1] ) );
  INV_X2 U5782 ( .I(\SB1_3_5/buf_output[3] ), .ZN(\SB2_3_3/i0[8] ) );
  NAND4_X2 U5783 ( .A1(\SB1_3_5/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_5/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_5/Component_Function_3/NAND4_in[2] ), .A4(n2317), .ZN(
        \SB1_3_5/buf_output[3] ) );
  XOR2_X1 U5786 ( .A1(\MC_ARK_ARC_1_2/temp5[13] ), .A2(
        \MC_ARK_ARC_1_2/temp6[13] ), .Z(\MC_ARK_ARC_1_2/buf_output[13] ) );
  BUF_X4 U5794 ( .I(\SB2_3_4/buf_output[1] ), .Z(\RI5[3][187] ) );
  NAND3_X1 U5795 ( .A1(\SB3_24/i0_4 ), .A2(\SB3_24/i0_0 ), .A3(\SB3_24/i0_3 ), 
        .ZN(\SB3_24/Component_Function_3/NAND4_in[1] ) );
  NOR2_X2 U5798 ( .A1(n1785), .A2(n1783), .ZN(n2237) );
  NAND3_X1 U5799 ( .A1(\SB2_0_23/i0[9] ), .A2(\SB2_0_23/i1_5 ), .A3(
        \SB2_0_23/i0[6] ), .ZN(\SB2_0_23/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U5800 ( .A1(\SB2_0_29/i0_3 ), .A2(n2605), .A3(\RI3[0][15] ), .ZN(
        \SB2_0_29/Component_Function_4/NAND4_in[2] ) );
  BUF_X4 U5803 ( .I(\SB2_0_25/buf_output[0] ), .Z(\RI5[0][66] ) );
  XOR2_X1 U5806 ( .A1(\RI5[0][60] ), .A2(\RI5[0][66] ), .Z(
        \MC_ARK_ARC_1_0/temp1[66] ) );
  NAND3_X1 U5807 ( .A1(\SB2_0_25/i0_0 ), .A2(\SB2_0_25/i0_3 ), .A3(
        \SB2_0_25/i0[7] ), .ZN(n1788) );
  BUF_X4 U5813 ( .I(\SB2_3_2/buf_output[3] ), .Z(\RI5[3][189] ) );
  NAND3_X1 U5814 ( .A1(\SB3_26/i0[6] ), .A2(\SB3_26/i0[8] ), .A3(
        \SB3_26/i0[7] ), .ZN(\SB3_26/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U5827 ( .A1(\RI5[2][121] ), .A2(\RI5[2][145] ), .Z(n1797) );
  NAND4_X2 U5828 ( .A1(\SB2_1_22/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_22/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_1_22/Component_Function_2/NAND4_in[1] ), .A4(n1798), .ZN(
        \SB2_1_22/buf_output[2] ) );
  XOR2_X1 U5833 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[114] ), .A2(\RI5[3][150] ), 
        .Z(n1800) );
  NAND3_X1 U5834 ( .A1(\SB3_15/i0_3 ), .A2(\SB3_15/i0[8] ), .A3(\SB3_15/i1_7 ), 
        .ZN(\SB3_15/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U5836 ( .A1(\MC_ARK_ARC_1_3/temp1[32] ), .A2(n1802), .Z(
        \MC_ARK_ARC_1_3/temp5[32] ) );
  XOR2_X1 U5837 ( .A1(\RI5[3][170] ), .A2(\RI5[3][2] ), .Z(n1802) );
  BUF_X4 U5839 ( .I(\SB2_2_22/buf_output[1] ), .Z(\RI5[2][79] ) );
  NAND4_X2 U5841 ( .A1(\SB1_3_24/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_3_24/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_24/Component_Function_0/NAND4_in[0] ), .A4(n1805), .ZN(
        \SB1_3_24/buf_output[0] ) );
  XOR2_X1 U5844 ( .A1(\RI5[0][168] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[132] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[66] ) );
  XOR2_X1 U5847 ( .A1(\RI5[1][146] ), .A2(\RI5[1][152] ), .Z(n1808) );
  NAND3_X2 U5855 ( .A1(\SB1_0_9/i0_3 ), .A2(\SB1_0_9/i0_4 ), .A3(
        \SB1_0_9/i1[9] ), .ZN(n1812) );
  NAND4_X2 U5863 ( .A1(\SB1_3_27/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_3_27/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_3_27/Component_Function_1/NAND4_in[0] ), .A4(n1817), .ZN(
        \SB1_3_27/buf_output[1] ) );
  NAND3_X1 U5864 ( .A1(\SB1_1_1/i0_0 ), .A2(\SB1_1_1/i3[0] ), .A3(
        \SB1_1_1/i1_7 ), .ZN(\SB1_1_1/Component_Function_4/NAND4_in[1] ) );
  NAND3_X2 U5867 ( .A1(\SB1_1_2/i0_4 ), .A2(\SB1_1_2/i1[9] ), .A3(
        \SB1_1_2/i0_3 ), .ZN(n2079) );
  XOR2_X1 U5868 ( .A1(\MC_ARK_ARC_1_3/temp3[37] ), .A2(
        \MC_ARK_ARC_1_3/temp4[37] ), .Z(\MC_ARK_ARC_1_3/temp6[37] ) );
  NAND3_X2 U5869 ( .A1(\SB2_1_18/i1_7 ), .A2(\SB2_1_18/i3[0] ), .A3(
        \SB2_1_18/i0_0 ), .ZN(\SB2_1_18/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U5870 ( .A1(\MC_ARK_ARC_1_0/temp5[167] ), .A2(n1821), .Z(
        \MC_ARK_ARC_1_0/buf_output[167] ) );
  XOR2_X1 U5871 ( .A1(\MC_ARK_ARC_1_0/temp3[167] ), .A2(
        \MC_ARK_ARC_1_0/temp4[167] ), .Z(n1821) );
  XOR2_X1 U5872 ( .A1(n2096), .A2(\MC_ARK_ARC_1_2/temp1[30] ), .Z(
        \MC_ARK_ARC_1_2/temp5[30] ) );
  XOR2_X1 U5873 ( .A1(n1823), .A2(n1822), .Z(\MC_ARK_ARC_1_0/buf_output[85] )
         );
  XOR2_X1 U5874 ( .A1(\MC_ARK_ARC_1_0/temp1[85] ), .A2(
        \MC_ARK_ARC_1_0/temp4[85] ), .Z(n1822) );
  XOR2_X1 U5875 ( .A1(\MC_ARK_ARC_1_0/temp3[85] ), .A2(
        \MC_ARK_ARC_1_0/temp2[85] ), .Z(n1823) );
  XOR2_X1 U5878 ( .A1(n1826), .A2(\MC_ARK_ARC_1_0/temp1[54] ), .Z(
        \MC_ARK_ARC_1_0/temp5[54] ) );
  BUF_X4 U5881 ( .I(\SB2_3_11/buf_output[4] ), .Z(\RI5[3][130] ) );
  NAND3_X1 U5883 ( .A1(\SB2_0_4/i1_7 ), .A2(\RI3[0][166] ), .A3(
        \SB2_0_4/i0[8] ), .ZN(n1827) );
  NAND4_X2 U5884 ( .A1(\SB1_0_15/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_0_15/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_0_15/Component_Function_0/NAND4_in[0] ), .A4(
        \SB1_0_15/Component_Function_0/NAND4_in[1] ), .ZN(\RI3[0][126] ) );
  NAND4_X2 U5885 ( .A1(\SB2_3_16/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_3_16/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_3_16/Component_Function_1/NAND4_in[0] ), .A4(n1828), .ZN(
        \SB2_3_16/buf_output[1] ) );
  NAND4_X2 U5893 ( .A1(\SB2_3_22/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_3_22/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_3_22/Component_Function_4/NAND4_in[3] ), .A4(n2076), .ZN(
        \SB2_3_22/buf_output[4] ) );
  XOR2_X1 U5897 ( .A1(\MC_ARK_ARC_1_3/temp3[33] ), .A2(
        \MC_ARK_ARC_1_3/temp4[33] ), .Z(n2666) );
  XOR2_X1 U5898 ( .A1(\MC_ARK_ARC_1_2/temp5[29] ), .A2(n1908), .Z(
        \MC_ARK_ARC_1_2/buf_output[29] ) );
  XOR2_X1 U5899 ( .A1(n2176), .A2(n2177), .Z(\MC_ARK_ARC_1_0/buf_output[7] )
         );
  NAND3_X1 U5901 ( .A1(\SB4_7/i0[9] ), .A2(\SB4_7/i0_3 ), .A3(\SB4_7/i0[8] ), 
        .ZN(n1830) );
  NAND3_X1 U5903 ( .A1(\SB1_0_13/i0_3 ), .A2(\SB1_0_13/i0_0 ), .A3(
        \SB1_0_13/i0[7] ), .ZN(n1832) );
  NAND3_X1 U5904 ( .A1(\SB1_0_13/i0_3 ), .A2(\SB1_0_13/i0[10] ), .A3(
        \SB1_0_13/i0_4 ), .ZN(n1833) );
  XOR2_X1 U5906 ( .A1(\RI5[1][76] ), .A2(\RI5[1][112] ), .Z(
        \MC_ARK_ARC_1_1/temp3[10] ) );
  NAND3_X1 U5907 ( .A1(\SB2_3_5/i0_0 ), .A2(\SB2_3_5/i3[0] ), .A3(
        \SB2_3_5/i1_7 ), .ZN(\SB2_3_5/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U5908 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[166] ), .A2(\RI5[3][190] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[28] ) );
  BUF_X4 U5911 ( .I(\SB2_1_11/buf_output[1] ), .Z(\RI5[1][145] ) );
  NAND3_X2 U5913 ( .A1(\SB1_3_26/i0[10] ), .A2(\SB1_3_26/i1[9] ), .A3(
        \SB1_3_26/i1_7 ), .ZN(n1838) );
  NAND2_X1 U5915 ( .A1(\SB1_2_2/i1[9] ), .A2(\SB1_2_2/i0_3 ), .ZN(
        \SB1_2_2/Component_Function_1/NAND4_in[0] ) );
  XOR2_X1 U5916 ( .A1(n1839), .A2(n1989), .Z(\MC_ARK_ARC_1_1/buf_output[15] )
         );
  NAND3_X1 U5918 ( .A1(\SB1_3_18/i0_0 ), .A2(\SB1_3_18/i0_3 ), .A3(
        \SB1_3_18/i0[7] ), .ZN(n2546) );
  BUF_X4 U5929 ( .I(\SB2_3_13/buf_output[2] ), .Z(\RI5[3][128] ) );
  XOR2_X1 U5933 ( .A1(n2209), .A2(n1846), .Z(\MC_ARK_ARC_1_0/buf_output[95] )
         );
  XOR2_X1 U5934 ( .A1(\MC_ARK_ARC_1_0/temp3[95] ), .A2(
        \MC_ARK_ARC_1_0/temp4[95] ), .Z(n1846) );
  BUF_X4 U5935 ( .I(\SB2_3_10/buf_output[3] ), .Z(\RI5[3][141] ) );
  XOR2_X1 U5944 ( .A1(\MC_ARK_ARC_1_0/temp3[186] ), .A2(
        \MC_ARK_ARC_1_0/temp4[186] ), .Z(n1850) );
  NAND3_X1 U5949 ( .A1(\SB3_7/i0[8] ), .A2(\SB3_7/i0_3 ), .A3(\SB3_7/i1_7 ), 
        .ZN(\SB3_7/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U5950 ( .A1(\SB1_2_15/i0[6] ), .A2(\SB1_2_15/i0[8] ), .A3(
        \SB1_2_15/i0[7] ), .ZN(\SB1_2_15/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U5954 ( .A1(\MC_ARK_ARC_1_0/buf_output[166] ), .A2(\SB1_1_4/i1_7 ), 
        .A3(\SB1_1_4/i0[8] ), .ZN(\SB1_1_4/Component_Function_1/NAND4_in[3] )
         );
  XOR2_X1 U5961 ( .A1(\MC_ARK_ARC_1_0/temp5[32] ), .A2(n1855), .Z(
        \MC_ARK_ARC_1_0/buf_output[32] ) );
  XOR2_X1 U5962 ( .A1(\MC_ARK_ARC_1_0/temp3[32] ), .A2(
        \MC_ARK_ARC_1_0/temp4[32] ), .Z(n1855) );
  XOR2_X1 U5964 ( .A1(\MC_ARK_ARC_1_0/temp4[153] ), .A2(n1946), .Z(n1856) );
  NAND3_X2 U5972 ( .A1(\SB1_0_7/i0_3 ), .A2(\SB1_0_7/i1[9] ), .A3(n390), .ZN(
        \SB1_0_7/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U5973 ( .A1(\SB2_2_23/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_23/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_2_23/Component_Function_4/NAND4_in[1] ), .A4(n1860), .ZN(
        \SB2_2_23/buf_output[4] ) );
  XOR2_X1 U5977 ( .A1(n1864), .A2(n28), .Z(Ciphertext[167]) );
  NAND4_X2 U5978 ( .A1(\SB4_4/Component_Function_5/NAND4_in[2] ), .A2(
        \SB4_4/Component_Function_5/NAND4_in[1] ), .A3(
        \SB4_4/Component_Function_5/NAND4_in[3] ), .A4(
        \SB4_4/Component_Function_5/NAND4_in[0] ), .ZN(n1864) );
  NAND4_X2 U5979 ( .A1(n2446), .A2(\SB1_2_16/Component_Function_0/NAND4_in[2] ), .A3(\SB1_2_16/Component_Function_0/NAND4_in[3] ), .A4(
        \SB1_2_16/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_2_16/buf_output[0] ) );
  NAND3_X1 U5981 ( .A1(\SB3_24/i0_0 ), .A2(\SB3_24/i1_7 ), .A3(\SB3_24/i3[0] ), 
        .ZN(\SB3_24/Component_Function_4/NAND4_in[1] ) );
  NAND2_X1 U5984 ( .A1(\SB1_0_24/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_0_24/Component_Function_4/NAND4_in[0] ), .ZN(n2425) );
  NAND3_X1 U5985 ( .A1(\SB2_3_20/i0[7] ), .A2(\SB2_3_20/i0_3 ), .A3(
        \SB2_3_20/i0_0 ), .ZN(\SB2_3_20/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U5986 ( .A1(\SB2_2_15/i0_3 ), .A2(\SB2_2_15/i0_4 ), .A3(
        \SB2_2_15/i1[9] ), .ZN(n1866) );
  NAND3_X1 U5987 ( .A1(\SB4_15/i0_0 ), .A2(\SB4_15/i0_4 ), .A3(\SB4_15/i1_5 ), 
        .ZN(n1867) );
  XOR2_X1 U5989 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[38] ), .A2(\RI5[1][2] ), 
        .Z(n1868) );
  XOR2_X1 U5991 ( .A1(n1870), .A2(\MC_ARK_ARC_1_3/temp1[190] ), .Z(
        \MC_ARK_ARC_1_3/temp5[190] ) );
  XOR2_X1 U5992 ( .A1(\RI5[3][160] ), .A2(\RI5[3][136] ), .Z(n1870) );
  NAND4_X2 U5993 ( .A1(\SB2_3_10/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_3_10/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_3_10/Component_Function_4/NAND4_in[1] ), .A4(n1872), .ZN(
        \SB2_3_10/buf_output[4] ) );
  XOR2_X1 U5998 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[27] ), .A2(\RI5[2][33] ), 
        .Z(n1874) );
  NAND3_X2 U5999 ( .A1(\SB2_1_24/i0_3 ), .A2(\SB2_1_24/i1[9] ), .A3(
        \SB2_1_24/i0_4 ), .ZN(\SB2_1_24/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U6001 ( .A1(\RI5[3][131] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[101] ), 
        .Z(n2661) );
  XOR2_X1 U6004 ( .A1(\MC_ARK_ARC_1_0/temp5[137] ), .A2(n1877), .Z(
        \MC_ARK_ARC_1_0/buf_output[137] ) );
  XOR2_X1 U6006 ( .A1(\MC_ARK_ARC_1_1/temp2[139] ), .A2(
        \MC_ARK_ARC_1_1/temp4[139] ), .Z(n1878) );
  NAND4_X2 U6010 ( .A1(\SB1_1_0/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_1_0/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_1_0/Component_Function_0/NAND4_in[0] ), .A4(n1880), .ZN(
        \SB1_1_0/buf_output[0] ) );
  XOR2_X1 U6013 ( .A1(\RI5[3][37] ), .A2(\RI5[3][43] ), .Z(n1882) );
  NAND3_X1 U6015 ( .A1(\SB1_0_28/i0[10] ), .A2(\SB1_0_28/i1[9] ), .A3(
        \SB1_0_28/i1_7 ), .ZN(\SB1_0_28/Component_Function_3/NAND4_in[2] ) );
  NAND4_X2 U6016 ( .A1(\SB1_3_23/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_3_23/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_3_23/Component_Function_0/NAND4_in[2] ), .A4(n2356), .ZN(
        \SB1_3_23/buf_output[0] ) );
  NAND4_X2 U6017 ( .A1(\SB2_3_22/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_3_22/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_3_22/Component_Function_0/NAND4_in[1] ), .A4(
        \SB2_3_22/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_3_22/buf_output[0] ) );
  NAND3_X2 U6018 ( .A1(\SB1_2_21/i0_3 ), .A2(\SB1_2_21/i0[9] ), .A3(
        \SB1_2_21/i0[10] ), .ZN(n1886) );
  NAND3_X1 U6021 ( .A1(\SB4_20/i0[8] ), .A2(\SB4_20/i3[0] ), .A3(n3674), .ZN(
        n1888) );
  XOR2_X1 U6028 ( .A1(n1890), .A2(\MC_ARK_ARC_1_2/temp6[16] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[16] ) );
  XOR2_X1 U6029 ( .A1(\MC_ARK_ARC_1_2/temp1[16] ), .A2(n2092), .Z(n1890) );
  XOR2_X1 U6030 ( .A1(n1891), .A2(\MC_ARK_ARC_1_3/temp5[153] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[153] ) );
  XOR2_X1 U6033 ( .A1(\MC_ARK_ARC_1_3/temp5[173] ), .A2(n1892), .Z(
        \MC_ARK_ARC_1_3/buf_output[173] ) );
  XOR2_X1 U6037 ( .A1(\RI5[0][47] ), .A2(\RI5[0][71] ), .Z(
        \MC_ARK_ARC_1_0/temp2[101] ) );
  NOR2_X2 U6039 ( .A1(n2168), .A2(n1894), .ZN(\SB2_2_1/i0[7] ) );
  BUF_X4 U6041 ( .I(\SB2_2_29/buf_output[0] ), .Z(\RI5[2][42] ) );
  INV_X2 U6042 ( .I(\SB1_3_29/buf_output[5] ), .ZN(\SB2_3_29/i1_5 ) );
  NAND4_X2 U6043 ( .A1(n2227), .A2(\SB2_0_27/Component_Function_5/NAND4_in[2] ), .A3(\SB2_0_27/Component_Function_5/NAND4_in[0] ), .A4(n1895), .ZN(
        \SB2_0_27/buf_output[5] ) );
  NAND3_X2 U6044 ( .A1(\SB2_1_18/i1_7 ), .A2(\SB2_1_18/i0_3 ), .A3(
        \SB2_1_18/i0[8] ), .ZN(\SB2_1_18/Component_Function_1/NAND4_in[1] ) );
  INV_X4 U6054 ( .I(n2563), .ZN(\SB1_3_9/buf_output[4] ) );
  BUF_X4 U6060 ( .I(\SB2_1_6/buf_output[1] ), .Z(\RI5[1][175] ) );
  XOR2_X1 U6062 ( .A1(n1909), .A2(\MC_ARK_ARC_1_0/temp6[182] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[182] ) );
  XOR2_X1 U6067 ( .A1(\SB2_1_4/buf_output[2] ), .A2(\RI5[1][176] ), .Z(
        \MC_ARK_ARC_1_1/temp1[182] ) );
  NAND3_X1 U6068 ( .A1(n2738), .A2(\SB2_0_10/i0_0 ), .A3(\SB2_0_10/i0_3 ), 
        .ZN(n1912) );
  BUF_X4 U6070 ( .I(\SB2_2_30/buf_output[5] ), .Z(\RI5[2][11] ) );
  NAND3_X1 U6078 ( .A1(\SB4_0/i0_3 ), .A2(\SB4_0/i0_4 ), .A3(n1386), .ZN(
        \SB4_0/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U6079 ( .A1(\RI5[1][67] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[31] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[157] ) );
  NAND3_X1 U6080 ( .A1(\SB4_28/i0_3 ), .A2(\SB4_28/i0[10] ), .A3(\SB4_28/i0_4 ), .ZN(n1918) );
  XOR2_X1 U6083 ( .A1(\RI5[3][160] ), .A2(\RI5[3][184] ), .Z(
        \MC_ARK_ARC_1_3/temp2[22] ) );
  NAND2_X1 U6087 ( .A1(\SB4_27/i0_3 ), .A2(n1389), .ZN(n1921) );
  NAND3_X1 U6092 ( .A1(\SB2_1_5/i0_0 ), .A2(\SB2_1_5/i3[0] ), .A3(
        \SB2_1_5/i1_7 ), .ZN(\SB2_1_5/Component_Function_4/NAND4_in[1] ) );
  BUF_X4 U6095 ( .I(\SB2_1_4/buf_output[3] ), .Z(\RI5[1][177] ) );
  XOR2_X1 U6096 ( .A1(\RI5[3][164] ), .A2(\RI5[3][188] ), .Z(n1925) );
  XOR2_X1 U6102 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[105] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[69] ), .Z(\MC_ARK_ARC_1_0/temp3[3] ) );
  BUF_X4 U6105 ( .I(\SB2_2_22/buf_output[0] ), .Z(\RI5[2][84] ) );
  NAND4_X2 U6106 ( .A1(\SB1_0_27/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_0_27/Component_Function_0/NAND4_in[1] ), .A3(n2273), .A4(
        \SB1_0_27/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_0_27/buf_output[0] ) );
  NAND3_X1 U6107 ( .A1(\SB1_2_25/i0[6] ), .A2(\SB1_2_25/i0_3 ), .A3(
        \SB1_2_25/i0[10] ), .ZN(\SB1_2_25/Component_Function_2/NAND4_in[1] )
         );
  XOR2_X1 U6109 ( .A1(n1932), .A2(n1931), .Z(\MC_ARK_ARC_1_3/buf_output[186] )
         );
  XOR2_X1 U6110 ( .A1(\MC_ARK_ARC_1_3/temp2[186] ), .A2(
        \MC_ARK_ARC_1_3/temp4[186] ), .Z(n1931) );
  XOR2_X1 U6111 ( .A1(\MC_ARK_ARC_1_3/temp3[186] ), .A2(
        \MC_ARK_ARC_1_3/temp1[186] ), .Z(n1932) );
  XOR2_X1 U6113 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[104] ), .A2(\RI5[3][128] ), 
        .Z(n1933) );
  XOR2_X1 U6115 ( .A1(n1935), .A2(\MC_ARK_ARC_1_2/temp1[124] ), .Z(
        \MC_ARK_ARC_1_2/temp5[124] ) );
  XOR2_X1 U6116 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[70] ), .A2(\RI5[2][94] ), 
        .Z(n1935) );
  XOR2_X1 U6122 ( .A1(\MC_ARK_ARC_1_2/temp1[183] ), .A2(
        \MC_ARK_ARC_1_2/temp2[183] ), .Z(n1937) );
  BUF_X4 U6132 ( .I(\SB2_2_27/buf_output[2] ), .Z(\RI5[2][44] ) );
  NAND3_X2 U6137 ( .A1(\SB1_1_26/i0_3 ), .A2(\SB1_1_26/i1[9] ), .A3(
        \SB1_1_26/i0_4 ), .ZN(n1940) );
  INV_X2 U6138 ( .I(\SB1_2_1/buf_output[3] ), .ZN(\SB2_2_31/i0[8] ) );
  NAND3_X1 U6144 ( .A1(\SB2_2_30/i0_0 ), .A2(\SB2_2_30/i3[0] ), .A3(
        \SB2_2_30/i1_7 ), .ZN(\SB2_2_30/Component_Function_4/NAND4_in[1] ) );
  INV_X2 U6147 ( .I(\RI3[0][182] ), .ZN(\SB2_0_1/i1[9] ) );
  BUF_X4 U6149 ( .I(\SB2_3_23/buf_output[1] ), .Z(\RI5[3][73] ) );
  BUF_X4 U6151 ( .I(\SB2_2_11/buf_output[0] ), .Z(\RI5[2][150] ) );
  XOR2_X1 U6154 ( .A1(\MC_ARK_ARC_1_0/temp5[151] ), .A2(n1945), .Z(
        \MC_ARK_ARC_1_0/buf_output[151] ) );
  XOR2_X1 U6155 ( .A1(\MC_ARK_ARC_1_0/temp3[151] ), .A2(
        \MC_ARK_ARC_1_0/temp4[151] ), .Z(n1945) );
  NAND4_X2 U6158 ( .A1(\SB3_19/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_19/Component_Function_0/NAND4_in[3] ), .A3(
        \SB3_19/Component_Function_0/NAND4_in[1] ), .A4(
        \SB3_19/Component_Function_0/NAND4_in[0] ), .ZN(\SB3_19/buf_output[0] ) );
  BUF_X4 U6159 ( .I(\SB2_3_2/buf_output[2] ), .Z(\RI5[3][2] ) );
  INV_X2 U6160 ( .I(\SB1_2_11/buf_output[2] ), .ZN(\SB2_2_8/i1[9] ) );
  NAND4_X2 U6161 ( .A1(\SB1_2_11/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_2_11/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_2_11/Component_Function_2/NAND4_in[1] ), .A4(n2843), .ZN(
        \SB1_2_11/buf_output[2] ) );
  NAND3_X1 U6164 ( .A1(\SB4_4/i0[10] ), .A2(\SB3_7/buf_output[2] ), .A3(
        \SB4_4/i0[6] ), .ZN(\SB4_4/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U6166 ( .A1(\MC_ARK_ARC_1_0/temp4[5] ), .A2(
        \MC_ARK_ARC_1_0/temp3[5] ), .Z(\MC_ARK_ARC_1_0/temp6[5] ) );
  XOR2_X1 U6172 ( .A1(\MC_ARK_ARC_1_3/temp3[180] ), .A2(
        \MC_ARK_ARC_1_3/temp4[180] ), .Z(\MC_ARK_ARC_1_3/temp6[180] ) );
  XOR2_X1 U6179 ( .A1(\MC_ARK_ARC_1_2/temp5[180] ), .A2(n1955), .Z(
        \MC_ARK_ARC_1_2/buf_output[180] ) );
  XOR2_X1 U6180 ( .A1(\MC_ARK_ARC_1_2/temp3[180] ), .A2(
        \MC_ARK_ARC_1_2/temp4[180] ), .Z(n1955) );
  BUF_X4 U6181 ( .I(\SB2_2_0/buf_output[0] ), .Z(\RI5[2][24] ) );
  NAND3_X1 U6183 ( .A1(\SB2_3_25/i0[7] ), .A2(\SB2_3_25/i0[6] ), .A3(
        \SB2_3_25/i0[8] ), .ZN(n2134) );
  XOR2_X1 U6187 ( .A1(\MC_ARK_ARC_1_2/temp5[49] ), .A2(n2325), .Z(
        \MC_ARK_ARC_1_2/buf_output[49] ) );
  NAND4_X2 U6188 ( .A1(\SB2_0_5/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_5/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_0_5/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_0_5/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_0_5/buf_output[5] ) );
  XOR2_X1 U6189 ( .A1(\MC_ARK_ARC_1_3/temp6[133] ), .A2(
        \MC_ARK_ARC_1_3/temp5[133] ), .Z(\MC_ARK_ARC_1_3/buf_output[133] ) );
  XOR2_X1 U6201 ( .A1(\MC_ARK_ARC_1_0/temp5[111] ), .A2(n1964), .Z(
        \MC_ARK_ARC_1_0/buf_output[111] ) );
  BUF_X4 U6210 ( .I(\SB2_1_14/buf_output[3] ), .Z(\RI5[1][117] ) );
  BUF_X4 U6218 ( .I(\SB2_0_28/buf_output[2] ), .Z(\RI5[0][38] ) );
  NAND3_X2 U6223 ( .A1(\SB1_0_12/i0_0 ), .A2(\SB1_0_12/i1_5 ), .A3(
        \SB1_0_12/i0_4 ), .ZN(n1978) );
  NAND3_X1 U6225 ( .A1(\SB2_1_27/i0_3 ), .A2(\SB1_1_0/buf_output[0] ), .A3(
        \SB2_1_27/i0[8] ), .ZN(\SB2_1_27/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U6227 ( .A1(\SB4_6/i0_4 ), .A2(\SB4_6/i0_3 ), .A3(\SB4_6/i1[9] ), 
        .ZN(\SB4_6/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U6228 ( .A1(\SB2_1_28/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_28/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_1_28/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_1_28/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_1_28/buf_output[5] ) );
  NAND4_X2 U6229 ( .A1(\SB1_0_19/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_19/Component_Function_4/NAND4_in[2] ), .A3(
        \SB1_0_19/Component_Function_4/NAND4_in[3] ), .A4(
        \SB1_0_19/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB1_0_19/buf_output[4] ) );
  NAND4_X2 U6239 ( .A1(\SB2_2_28/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_2_28/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_28/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_2_28/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_2_28/buf_output[0] ) );
  NAND4_X2 U6243 ( .A1(\SB2_3_29/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_29/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_3_29/Component_Function_4/NAND4_in[1] ), .A4(n1986), .ZN(
        \SB2_3_29/buf_output[4] ) );
  NAND3_X1 U6245 ( .A1(\SB1_2_16/i0_0 ), .A2(\RI1[2][95] ), .A3(
        \SB1_2_16/i0[7] ), .ZN(\SB1_2_16/Component_Function_0/NAND4_in[3] ) );
  NAND3_X2 U6247 ( .A1(\SB2_2_8/i0_3 ), .A2(\SB2_2_8/i0[9] ), .A3(
        \SB2_2_8/i0[8] ), .ZN(\SB2_2_8/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 U6248 ( .I(\SB2_0_28/buf_output[4] ), .Z(\RI5[0][28] ) );
  NAND4_X2 U6249 ( .A1(\SB1_0_19/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_0_19/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_0_19/Component_Function_1/NAND4_in[1] ), .A4(n1988), .ZN(
        \RI3[0][97] ) );
  NAND2_X1 U6250 ( .A1(\SB1_0_19/i1[9] ), .A2(\SB1_0_19/i0_3 ), .ZN(n1988) );
  BUF_X4 U6255 ( .I(\SB2_3_21/buf_output[1] ), .Z(\RI5[3][85] ) );
  BUF_X4 U6256 ( .I(\SB2_3_29/buf_output[3] ), .Z(\RI5[3][27] ) );
  XOR2_X1 U6259 ( .A1(\RI5[2][80] ), .A2(\RI5[2][104] ), .Z(n1993) );
  XOR2_X1 U6271 ( .A1(\MC_ARK_ARC_1_3/temp5[25] ), .A2(n1998), .Z(
        \MC_ARK_ARC_1_3/buf_output[25] ) );
  NAND3_X2 U6274 ( .A1(\SB2_0_9/i1[9] ), .A2(\SB2_0_9/i0[10] ), .A3(n5518), 
        .ZN(\SB2_0_9/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U6275 ( .A1(\SB1_0_12/i0_4 ), .A2(\SB1_0_12/i0[9] ), .A3(
        \SB1_0_12/i0[6] ), .ZN(n2286) );
  NAND3_X2 U6276 ( .A1(\SB2_3_5/i0[10] ), .A2(n3671), .A3(\SB2_3_5/i1_7 ), 
        .ZN(\SB2_3_5/Component_Function_3/NAND4_in[2] ) );
  XOR2_X1 U6277 ( .A1(\RI5[0][38] ), .A2(\RI5[0][74] ), .Z(
        \MC_ARK_ARC_1_0/temp3[164] ) );
  NAND4_X2 U6279 ( .A1(\SB1_1_26/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_26/Component_Function_4/NAND4_in[3] ), .A3(
        \SB1_1_26/Component_Function_4/NAND4_in[1] ), .A4(n1999), .ZN(
        \SB1_1_26/buf_output[4] ) );
  NAND3_X2 U6280 ( .A1(\SB1_1_26/i0[10] ), .A2(\SB1_1_26/i0_3 ), .A3(
        \SB1_1_26/i0[9] ), .ZN(n1999) );
  XOR2_X1 U6282 ( .A1(n2119), .A2(n2000), .Z(\MC_ARK_ARC_1_0/buf_output[180] )
         );
  XOR2_X1 U6283 ( .A1(\MC_ARK_ARC_1_0/temp1[180] ), .A2(n2045), .Z(n2000) );
  BUF_X4 U6284 ( .I(\SB2_1_27/buf_output[0] ), .Z(\RI5[1][54] ) );
  NAND4_X2 U6285 ( .A1(\SB1_2_21/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_2_21/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_21/Component_Function_1/NAND4_in[0] ), .A4(n2001), .ZN(
        \SB1_2_21/buf_output[1] ) );
  NAND3_X1 U6286 ( .A1(\SB1_2_21/i0[8] ), .A2(\SB1_2_21/i0_4 ), .A3(
        \SB1_2_21/i1_7 ), .ZN(n2001) );
  XOR2_X1 U6291 ( .A1(\MC_ARK_ARC_1_3/temp5[32] ), .A2(
        \MC_ARK_ARC_1_3/temp6[32] ), .Z(\MC_ARK_ARC_1_3/buf_output[32] ) );
  XOR2_X1 U6294 ( .A1(n2007), .A2(\MC_ARK_ARC_1_0/temp5[124] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[124] ) );
  XOR2_X1 U6295 ( .A1(\MC_ARK_ARC_1_0/temp3[124] ), .A2(
        \MC_ARK_ARC_1_0/temp4[124] ), .Z(n2007) );
  XOR2_X1 U6296 ( .A1(\MC_ARK_ARC_1_0/temp5[190] ), .A2(n2008), .Z(
        \MC_ARK_ARC_1_0/buf_output[190] ) );
  XOR2_X1 U6297 ( .A1(\MC_ARK_ARC_1_0/temp4[190] ), .A2(
        \MC_ARK_ARC_1_0/temp3[190] ), .Z(n2008) );
  BUF_X4 U6300 ( .I(\SB2_1_14/buf_output[2] ), .Z(\RI5[1][122] ) );
  NAND2_X1 U6302 ( .A1(\SB4_25/i0[9] ), .A2(\SB4_25/i0[10] ), .ZN(n2009) );
  XOR2_X1 U6303 ( .A1(n2010), .A2(n121), .Z(Ciphertext[24]) );
  XOR2_X1 U6305 ( .A1(\RI5[0][34] ), .A2(\RI5[0][58] ), .Z(n2011) );
  NAND4_X2 U6307 ( .A1(\SB3_13/Component_Function_0/NAND4_in[3] ), .A2(
        \SB3_13/Component_Function_0/NAND4_in[2] ), .A3(
        \SB3_13/Component_Function_0/NAND4_in[1] ), .A4(
        \SB3_13/Component_Function_0/NAND4_in[0] ), .ZN(\SB3_13/buf_output[0] ) );
  NAND4_X2 U6308 ( .A1(n2681), .A2(\SB2_0_28/Component_Function_5/NAND4_in[1] ), .A3(\SB2_0_28/Component_Function_5/NAND4_in[0] ), .A4(n2014), .ZN(
        \SB2_0_28/buf_output[5] ) );
  XOR2_X1 U6309 ( .A1(\RI5[1][113] ), .A2(\RI5[1][149] ), .Z(
        \MC_ARK_ARC_1_1/temp3[47] ) );
  XOR2_X1 U6310 ( .A1(\MC_ARK_ARC_1_3/temp2[49] ), .A2(
        \MC_ARK_ARC_1_3/temp1[49] ), .Z(\MC_ARK_ARC_1_3/temp5[49] ) );
  XOR2_X1 U6312 ( .A1(n2831), .A2(\MC_ARK_ARC_1_2/temp5[15] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[15] ) );
  XOR2_X1 U6314 ( .A1(\RI5[1][138] ), .A2(\RI5[1][162] ), .Z(n2016) );
  XOR2_X1 U6318 ( .A1(\MC_ARK_ARC_1_2/temp3[105] ), .A2(
        \MC_ARK_ARC_1_2/temp4[105] ), .Z(n2019) );
  XOR2_X1 U6324 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[69] ), .A2(\RI5[0][45] ), 
        .Z(n2022) );
  NAND3_X1 U6331 ( .A1(\SB1_2_28/i0_0 ), .A2(\SB1_2_28/i3[0] ), .A3(
        \SB1_2_28/i1_7 ), .ZN(n2026) );
  XOR2_X1 U6338 ( .A1(\MC_ARK_ARC_1_3/temp5[141] ), .A2(n2031), .Z(
        \MC_ARK_ARC_1_3/buf_output[141] ) );
  XOR2_X1 U6339 ( .A1(\MC_ARK_ARC_1_3/temp3[141] ), .A2(
        \MC_ARK_ARC_1_3/temp4[141] ), .Z(n2031) );
  NAND2_X2 U6343 ( .A1(\SB1_0_14/Component_Function_4/NAND4_in[1] ), .A2(n2402), .ZN(n2401) );
  INV_X4 U6346 ( .I(n2711), .ZN(\SB2_0_13/i0_4 ) );
  XOR2_X1 U6347 ( .A1(n2034), .A2(\MC_ARK_ARC_1_2/temp6[88] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[88] ) );
  XOR2_X1 U6348 ( .A1(\MC_ARK_ARC_1_2/temp2[88] ), .A2(
        \MC_ARK_ARC_1_2/temp1[88] ), .Z(n2034) );
  XOR2_X1 U6349 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[56] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[92] ), .Z(\MC_ARK_ARC_1_0/temp3[182] )
         );
  NOR2_X2 U6351 ( .A1(n2037), .A2(n2035), .ZN(n2682) );
  NAND2_X1 U6353 ( .A1(\SB4_0/i0_3 ), .A2(n1386), .ZN(n2038) );
  NAND3_X1 U6354 ( .A1(\SB4_15/i0[10] ), .A2(\SB4_15/i0_3 ), .A3(\SB4_15/i0_4 ), .ZN(\SB4_15/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U6359 ( .A1(\SB3_11/i0_0 ), .A2(\SB3_11/i0[8] ), .A3(\SB3_11/i0[9] ), .ZN(n2039) );
  XOR2_X1 U6367 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[167] ), .A2(\RI5[0][143] ), 
        .Z(n2043) );
  XOR2_X1 U6369 ( .A1(\RI5[0][54] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[90] ), 
        .Z(n2045) );
  XOR2_X1 U6372 ( .A1(\RI5[2][130] ), .A2(\RI5[2][166] ), .Z(n2046) );
  XOR2_X1 U6381 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[156] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[162] ), .Z(\MC_ARK_ARC_1_2/temp1[162] )
         );
  BUF_X4 U6382 ( .I(\SB2_2_18/buf_output[0] ), .Z(\RI5[2][108] ) );
  NAND4_X2 U6384 ( .A1(n2128), .A2(\SB2_3_4/Component_Function_3/NAND4_in[2] ), 
        .A3(\SB2_3_4/Component_Function_3/NAND4_in[3] ), .A4(n2053), .ZN(
        \SB2_3_4/buf_output[3] ) );
  XOR2_X1 U6386 ( .A1(\MC_ARK_ARC_1_0/temp3[184] ), .A2(n2055), .Z(n2640) );
  XOR2_X1 U6387 ( .A1(\RI5[0][130] ), .A2(\RI5[0][154] ), .Z(n2055) );
  XOR2_X1 U6388 ( .A1(\RI5[3][189] ), .A2(n242), .Z(n2056) );
  XOR2_X1 U6389 ( .A1(\RI5[3][63] ), .A2(\RI5[3][27] ), .Z(n2057) );
  NAND3_X1 U6394 ( .A1(\SB3_6/i0[8] ), .A2(\SB3_6/i1_7 ), .A3(\RI1[4][155] ), 
        .ZN(\SB3_6/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 U6404 ( .A1(\SB4_25/i0_3 ), .A2(\SB4_25/i1[9] ), .ZN(n2063) );
  NAND3_X1 U6405 ( .A1(\SB2_3_1/i0[10] ), .A2(\SB2_3_1/i0_3 ), .A3(
        \SB2_3_1/i0_4 ), .ZN(\SB2_3_1/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U6408 ( .A1(\SB4_25/i0_0 ), .A2(\SB4_25/i0[10] ), .A3(
        \SB4_25/i0[6] ), .ZN(\SB4_25/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 U6414 ( .I(\SB2_3_1/buf_output[0] ), .Z(\RI5[3][18] ) );
  BUF_X4 U6421 ( .I(\SB2_2_22/buf_output[3] ), .Z(\RI5[2][69] ) );
  XOR2_X1 U6423 ( .A1(\MC_ARK_ARC_1_3/temp2[2] ), .A2(
        \MC_ARK_ARC_1_3/temp1[2] ), .Z(n2069) );
  NAND2_X1 U6425 ( .A1(\SB3_5/i0_3 ), .A2(\SB3_5/i1[9] ), .ZN(n2070) );
  XOR2_X1 U6429 ( .A1(n2073), .A2(\MC_ARK_ARC_1_0/temp1[28] ), .Z(
        \MC_ARK_ARC_1_0/temp5[28] ) );
  BUF_X4 U6431 ( .I(\SB2_3_3/buf_output[3] ), .Z(\RI5[3][183] ) );
  XOR2_X1 U6432 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[176] ), .A2(\RI5[3][8] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[38] ) );
  NAND3_X1 U6433 ( .A1(\SB1_0_19/i0_0 ), .A2(\SB1_0_19/i1_5 ), .A3(
        \SB1_0_19/i0_4 ), .ZN(\SB1_0_19/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U6438 ( .A1(\SB3_25/i0[6] ), .A2(\SB3_25/i0[8] ), .A3(
        \SB3_25/i0[7] ), .ZN(\SB3_25/Component_Function_0/NAND4_in[1] ) );
  NAND3_X2 U6446 ( .A1(\SB1_2_29/i1_5 ), .A2(\SB1_2_29/i1[9] ), .A3(
        \SB1_2_29/i0_4 ), .ZN(\SB1_2_29/Component_Function_4/NAND4_in[3] ) );
  XOR2_X1 U6447 ( .A1(\MC_ARK_ARC_1_0/temp6[150] ), .A2(
        \MC_ARK_ARC_1_0/temp5[150] ), .Z(\MC_ARK_ARC_1_0/buf_output[150] ) );
  XOR2_X1 U6448 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[160] ), .A2(\RI5[1][166] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[166] ) );
  BUF_X4 U6449 ( .I(\SB2_2_17/buf_output[2] ), .Z(\RI5[2][104] ) );
  XOR2_X1 U6450 ( .A1(\MC_ARK_ARC_1_1/temp5[66] ), .A2(n2080), .Z(
        \MC_ARK_ARC_1_1/buf_output[66] ) );
  XOR2_X1 U6451 ( .A1(\MC_ARK_ARC_1_1/temp4[66] ), .A2(
        \MC_ARK_ARC_1_1/temp3[66] ), .Z(n2080) );
  XOR2_X1 U6452 ( .A1(\MC_ARK_ARC_1_1/temp5[119] ), .A2(n2081), .Z(
        \MC_ARK_ARC_1_1/buf_output[119] ) );
  XOR2_X1 U6453 ( .A1(\MC_ARK_ARC_1_1/temp3[119] ), .A2(
        \MC_ARK_ARC_1_1/temp4[119] ), .Z(n2081) );
  NAND4_X2 U6456 ( .A1(\SB2_1_6/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_1_6/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_6/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_1_6/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_1_6/buf_output[4] ) );
  XOR2_X1 U6459 ( .A1(\MC_ARK_ARC_1_1/temp2[1] ), .A2(
        \MC_ARK_ARC_1_1/temp1[1] ), .Z(n2083) );
  XOR2_X1 U6460 ( .A1(\MC_ARK_ARC_1_0/temp4[114] ), .A2(
        \MC_ARK_ARC_1_0/temp2[114] ), .Z(n2448) );
  BUF_X4 U6461 ( .I(\SB2_2_31/buf_output[2] ), .Z(\RI5[2][20] ) );
  BUF_X4 U6462 ( .I(\SB2_3_27/buf_output[0] ), .Z(\RI5[3][54] ) );
  XOR2_X1 U6463 ( .A1(n2084), .A2(\MC_ARK_ARC_1_1/temp2[108] ), .Z(n2418) );
  XOR2_X1 U6464 ( .A1(\RI5[1][102] ), .A2(\RI5[1][108] ), .Z(n2084) );
  XOR2_X1 U6467 ( .A1(\MC_ARK_ARC_1_2/temp1[61] ), .A2(
        \MC_ARK_ARC_1_2/temp2[61] ), .Z(n2086) );
  XOR2_X1 U6468 ( .A1(\MC_ARK_ARC_1_2/temp3[61] ), .A2(
        \MC_ARK_ARC_1_2/temp4[61] ), .Z(n2087) );
  NAND3_X1 U6475 ( .A1(\SB2_1_4/i0[10] ), .A2(\SB2_1_4/i1_5 ), .A3(n3660), 
        .ZN(\SB2_1_4/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U6478 ( .A1(n2091), .A2(n2438), .Z(\MC_ARK_ARC_1_2/buf_output[176] )
         );
  XOR2_X1 U6479 ( .A1(\MC_ARK_ARC_1_2/temp2[176] ), .A2(
        \MC_ARK_ARC_1_2/temp1[176] ), .Z(n2091) );
  XOR2_X1 U6480 ( .A1(\RI5[2][154] ), .A2(\RI5[2][178] ), .Z(n2092) );
  NAND3_X2 U6483 ( .A1(\SB2_0_29/i0[8] ), .A2(\SB2_0_29/i3[0] ), .A3(
        \SB2_0_29/i1_5 ), .ZN(n2093) );
  NAND3_X1 U6484 ( .A1(\SB2_2_1/i0_0 ), .A2(\SB2_2_1/i0[9] ), .A3(
        \SB2_2_1/i0[8] ), .ZN(\SB2_2_1/Component_Function_4/NAND4_in[0] ) );
  INV_X4 U6486 ( .I(\SB2_3_15/i0[7] ), .ZN(\SB1_3_16/buf_output[4] ) );
  NAND3_X1 U6487 ( .A1(\SB2_3_15/i0_0 ), .A2(\SB2_3_15/i0_3 ), .A3(
        \SB2_3_15/i0[7] ), .ZN(\SB2_3_15/Component_Function_0/NAND4_in[3] ) );
  XOR2_X1 U6491 ( .A1(\RI5[2][168] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[0] ), 
        .Z(n2096) );
  NAND3_X1 U6498 ( .A1(\SB1_3_18/i0[9] ), .A2(\SB1_3_18/i1_5 ), .A3(
        \SB1_3_18/i0[6] ), .ZN(\SB1_3_18/Component_Function_1/NAND4_in[2] ) );
  NAND4_X2 U6499 ( .A1(\SB1_1_1/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_1_1/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_1_1/Component_Function_0/NAND4_in[0] ), .A4(n2100), .ZN(
        \SB1_1_1/buf_output[0] ) );
  NAND3_X1 U6501 ( .A1(\SB1_2_9/i0[6] ), .A2(\SB1_2_9/i0_3 ), .A3(
        \SB1_2_9/i0[10] ), .ZN(\SB1_2_9/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U6503 ( .A1(\MC_ARK_ARC_1_3/buf_output[10] ), .A2(\SB3_30/i1_7 ), 
        .A3(\SB3_30/i0[8] ), .ZN(n2101) );
  NAND3_X1 U6505 ( .A1(\SB4_26/i0[6] ), .A2(\SB4_26/i0_4 ), .A3(\SB4_26/i0[9] ), .ZN(n2102) );
  NAND3_X1 U6507 ( .A1(\SB4_26/i0[6] ), .A2(\SB4_26/i0_3 ), .A3(\SB4_26/i1[9] ), .ZN(n2103) );
  XOR2_X1 U6510 ( .A1(n2240), .A2(\MC_ARK_ARC_1_3/temp2[147] ), .Z(
        \MC_ARK_ARC_1_3/temp5[147] ) );
  NAND3_X1 U6519 ( .A1(\SB1_0_29/i0_0 ), .A2(\SB1_0_29/i3[0] ), .A3(
        \SB1_0_29/i1_7 ), .ZN(\SB1_0_29/Component_Function_4/NAND4_in[1] ) );
  BUF_X4 U6520 ( .I(\SB2_0_28/buf_output[1] ), .Z(\RI5[0][43] ) );
  XOR2_X1 U6524 ( .A1(\RI5[3][84] ), .A2(\RI5[3][108] ), .Z(n2110) );
  NAND3_X1 U6527 ( .A1(\SB1_2_2/i0_0 ), .A2(\SB1_2_2/i3[0] ), .A3(
        \SB1_2_2/i1_7 ), .ZN(\SB1_2_2/Component_Function_4/NAND4_in[1] ) );
  INV_X1 U6528 ( .I(\SB3_16/buf_output[1] ), .ZN(\SB4_12/i1_7 ) );
  NAND3_X1 U6533 ( .A1(n2852), .A2(\SB2_1_7/i1_5 ), .A3(\SB2_1_7/i0[9] ), .ZN(
        \SB2_1_7/Component_Function_1/NAND4_in[2] ) );
  XOR2_X1 U6539 ( .A1(\MC_ARK_ARC_1_0/temp2[180] ), .A2(
        \MC_ARK_ARC_1_0/temp4[180] ), .Z(n2119) );
  XOR2_X1 U6540 ( .A1(\RI5[0][72] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[96] ), 
        .Z(n2120) );
  NAND3_X1 U6543 ( .A1(\SB1_0_10/i0_0 ), .A2(\SB1_0_10/i1_5 ), .A3(
        \SB1_0_10/i0_4 ), .ZN(n2121) );
  NAND2_X1 U6545 ( .A1(\SB1_3_25/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_3_25/Component_Function_4/NAND4_in[0] ), .ZN(n2123) );
  NAND4_X2 U6546 ( .A1(\SB1_3_25/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_3_25/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_3_25/Component_Function_1/NAND4_in[0] ), .A4(n2125), .ZN(
        \SB1_3_25/buf_output[1] ) );
  XOR2_X1 U6548 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[82] ), .A2(\RI5[3][118] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[16] ) );
  XOR2_X1 U6552 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[51] ), .A2(\RI5[0][87] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[177] ) );
  XOR2_X1 U6557 ( .A1(\RI5[0][95] ), .A2(\RI5[0][59] ), .Z(
        \MC_ARK_ARC_1_0/temp3[185] ) );
  XOR2_X1 U6558 ( .A1(\RI5[3][177] ), .A2(\RI5[3][21] ), .Z(
        \MC_ARK_ARC_1_3/temp3[111] ) );
  NAND3_X1 U6562 ( .A1(\SB4_6/i0_0 ), .A2(\SB4_6/i0[9] ), .A3(n579), .ZN(
        \SB4_6/Component_Function_4/NAND4_in[0] ) );
  XOR2_X1 U6565 ( .A1(n2132), .A2(\MC_ARK_ARC_1_3/temp4[134] ), .Z(
        \MC_ARK_ARC_1_3/temp6[134] ) );
  XOR2_X1 U6566 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[44] ), .A2(\RI5[3][8] ), 
        .Z(n2132) );
  XOR2_X1 U6571 ( .A1(\MC_ARK_ARC_1_1/temp6[166] ), .A2(n2140), .Z(
        \MC_ARK_ARC_1_1/buf_output[166] ) );
  XOR2_X1 U6572 ( .A1(\MC_ARK_ARC_1_1/temp1[166] ), .A2(
        \MC_ARK_ARC_1_1/temp2[166] ), .Z(n2140) );
  NAND4_X2 U6575 ( .A1(\SB2_2_18/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_2_18/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_2_18/Component_Function_0/NAND4_in[1] ), .A4(
        \SB2_2_18/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_2_18/buf_output[0] ) );
  NAND4_X2 U6576 ( .A1(\SB1_2_18/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_18/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_2_18/Component_Function_5/NAND4_in[0] ), .A4(n2142), .ZN(
        \SB1_2_18/buf_output[5] ) );
  NAND3_X2 U6577 ( .A1(\SB1_2_18/i0_3 ), .A2(\SB1_2_18/i1[9] ), .A3(
        \SB1_2_18/i0_4 ), .ZN(n2142) );
  XOR2_X1 U6578 ( .A1(\MC_ARK_ARC_1_3/temp4[181] ), .A2(
        \MC_ARK_ARC_1_3/temp3[181] ), .Z(n2143) );
  NAND3_X1 U6584 ( .A1(\SB2_3_25/i0[10] ), .A2(\SB2_3_25/i0_3 ), .A3(
        \SB1_3_26/buf_output[4] ), .ZN(
        \SB2_3_25/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U6585 ( .A1(\SB4_12/i0_0 ), .A2(\SB4_12/i0[9] ), .A3(\SB4_12/i0[8] ), .ZN(\SB4_12/Component_Function_4/NAND4_in[0] ) );
  XOR2_X1 U6588 ( .A1(\RI5[0][111] ), .A2(\RI5[0][147] ), .Z(
        \MC_ARK_ARC_1_0/temp3[45] ) );
  NAND4_X2 U6593 ( .A1(\SB1_0_15/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_0_15/Component_Function_2/NAND4_in[3] ), .A3(
        \SB1_0_15/Component_Function_2/NAND4_in[0] ), .A4(n2149), .ZN(
        \RI3[0][116] ) );
  XOR2_X1 U6594 ( .A1(n2150), .A2(\MC_ARK_ARC_1_0/temp4[148] ), .Z(
        \MC_ARK_ARC_1_0/temp6[148] ) );
  XOR2_X1 U6595 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[22] ), .A2(\RI5[0][58] ), 
        .Z(n2150) );
  INV_X2 U6598 ( .I(\SB1_1_1/buf_output[5] ), .ZN(\SB2_1_1/i1_5 ) );
  XOR2_X1 U6599 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[63] ), .A2(\RI5[1][69] ), 
        .Z(n2154) );
  NAND4_X2 U6602 ( .A1(\SB1_3_8/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_3_8/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_3_8/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_3_8/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_3_8/buf_output[0] ) );
  NAND4_X2 U6604 ( .A1(\SB2_0_26/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_0_26/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_0_26/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_26/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_0_26/buf_output[0] ) );
  BUF_X4 U6605 ( .I(\SB2_0_26/buf_output[0] ), .Z(\RI5[0][60] ) );
  INV_X2 U6606 ( .I(\SB1_3_19/buf_output[3] ), .ZN(\SB2_3_17/i0[8] ) );
  XOR2_X1 U6609 ( .A1(\MC_ARK_ARC_1_2/temp5[74] ), .A2(n2157), .Z(
        \MC_ARK_ARC_1_2/buf_output[74] ) );
  XOR2_X1 U6610 ( .A1(\MC_ARK_ARC_1_2/temp3[74] ), .A2(
        \MC_ARK_ARC_1_2/temp4[74] ), .Z(n2157) );
  XOR2_X1 U6613 ( .A1(n2161), .A2(n2162), .Z(\MC_ARK_ARC_1_1/buf_output[126] )
         );
  XOR2_X1 U6615 ( .A1(\MC_ARK_ARC_1_1/temp1[126] ), .A2(
        \MC_ARK_ARC_1_1/temp4[126] ), .Z(n2162) );
  XOR2_X1 U6618 ( .A1(\RI5[1][188] ), .A2(\RI5[1][164] ), .Z(n2164) );
  XOR2_X1 U6624 ( .A1(\RI5[0][34] ), .A2(\RI5[0][40] ), .Z(
        \MC_ARK_ARC_1_0/temp1[40] ) );
  BUF_X4 U6625 ( .I(\SB2_2_25/buf_output[0] ), .Z(\RI5[2][66] ) );
  NAND3_X1 U6626 ( .A1(\SB1_0_7/i0[10] ), .A2(\SB1_0_7/i0_0 ), .A3(
        \SB1_0_7/i0[6] ), .ZN(\SB1_0_7/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U6628 ( .A1(\SB2_2_1/i0[6] ), .A2(\SB2_2_1/i0[7] ), .A3(
        \SB2_2_1/i0[8] ), .ZN(\SB2_2_1/Component_Function_0/NAND4_in[1] ) );
  NAND4_X2 U6629 ( .A1(\SB1_2_10/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_10/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_10/Component_Function_0/NAND4_in[0] ), .A4(n2169), .ZN(
        \SB1_2_10/buf_output[0] ) );
  NAND3_X1 U6633 ( .A1(\SB1_3_27/i0[9] ), .A2(\SB1_3_27/i1_5 ), .A3(
        \SB1_3_27/i0[6] ), .ZN(\SB1_3_27/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U6637 ( .A1(\SB3_16/i0_4 ), .A2(\SB3_16/i1_7 ), .A3(\SB3_16/i0[8] ), 
        .ZN(n2171) );
  XOR2_X1 U6640 ( .A1(\RI5[3][77] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[101] ), 
        .Z(n2172) );
  XOR2_X1 U6642 ( .A1(\MC_ARK_ARC_1_1/temp4[3] ), .A2(
        \MC_ARK_ARC_1_1/temp3[3] ), .Z(n2174) );
  BUF_X4 U6644 ( .I(\SB2_0_27/buf_output[0] ), .Z(\RI5[0][54] ) );
  XOR2_X1 U6646 ( .A1(\MC_ARK_ARC_1_0/temp1[7] ), .A2(
        \MC_ARK_ARC_1_0/temp3[7] ), .Z(n2176) );
  XOR2_X1 U6647 ( .A1(\MC_ARK_ARC_1_0/temp2[7] ), .A2(
        \MC_ARK_ARC_1_0/temp4[7] ), .Z(n2177) );
  INV_X1 U6648 ( .I(\SB1_3_12/buf_output[1] ), .ZN(\SB2_3_8/i1_7 ) );
  BUF_X4 U6651 ( .I(\SB2_1_26/buf_output[1] ), .Z(\RI5[1][55] ) );
  NAND4_X2 U6659 ( .A1(\SB2_2_31/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_2_31/Component_Function_0/NAND4_in[0] ), .A3(
        \SB2_2_31/Component_Function_0/NAND4_in[2] ), .A4(n2181), .ZN(
        \SB2_2_31/buf_output[0] ) );
  XOR2_X1 U6671 ( .A1(n2186), .A2(\MC_ARK_ARC_1_2/temp6[156] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[156] ) );
  NAND4_X2 U6673 ( .A1(n2190), .A2(\SB2_0_17/Component_Function_4/NAND4_in[1] ), .A3(\SB2_0_17/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_0_17/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_0_17/buf_output[4] ) );
  NAND4_X2 U6674 ( .A1(\SB1_1_14/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_1_14/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_1_14/Component_Function_1/NAND4_in[0] ), .A4(n2192), .ZN(
        \SB1_1_14/buf_output[1] ) );
  XOR2_X1 U6675 ( .A1(n2193), .A2(\MC_ARK_ARC_1_3/temp1[169] ), .Z(
        \MC_ARK_ARC_1_3/temp5[169] ) );
  XOR2_X1 U6676 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[115] ), .A2(\RI5[3][139] ), 
        .Z(n2193) );
  INV_X1 U6677 ( .I(\SB1_2_2/buf_output[1] ), .ZN(\SB2_2_30/i1_7 ) );
  XOR2_X1 U6682 ( .A1(\RI5[0][154] ), .A2(\RI5[0][178] ), .Z(n2197) );
  XOR2_X1 U6684 ( .A1(\RI5[0][133] ), .A2(\RI5[0][103] ), .Z(n2198) );
  XOR2_X1 U6685 ( .A1(\RI5[0][127] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[79] ), 
        .Z(n2199) );
  NAND4_X2 U6690 ( .A1(\SB1_0_19/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_0_19/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_19/Component_Function_0/NAND4_in[0] ), .A4(n2201), .ZN(
        \SB1_0_19/buf_output[0] ) );
  XOR2_X1 U6692 ( .A1(\MC_ARK_ARC_1_2/temp2[186] ), .A2(
        \MC_ARK_ARC_1_2/temp1[186] ), .Z(\MC_ARK_ARC_1_2/temp5[186] ) );
  NAND3_X1 U6694 ( .A1(\SB2_3_20/i0[10] ), .A2(\SB2_3_20/i0_3 ), .A3(
        \SB2_3_20/i0[6] ), .ZN(\SB2_3_20/Component_Function_2/NAND4_in[1] ) );
  XOR2_X1 U6696 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[101] ), .A2(\RI5[1][77] ), 
        .Z(n2207) );
  XOR2_X1 U6697 ( .A1(\MC_ARK_ARC_1_0/temp2[108] ), .A2(
        \MC_ARK_ARC_1_0/temp1[108] ), .Z(\MC_ARK_ARC_1_0/temp5[108] ) );
  XOR2_X1 U6698 ( .A1(\MC_ARK_ARC_1_2/temp6[60] ), .A2(n2208), .Z(
        \MC_ARK_ARC_1_2/buf_output[60] ) );
  XOR2_X1 U6699 ( .A1(\MC_ARK_ARC_1_2/temp2[60] ), .A2(
        \MC_ARK_ARC_1_2/temp1[60] ), .Z(n2208) );
  NAND3_X2 U6702 ( .A1(\SB1_1_0/i0[8] ), .A2(\SB1_1_0/i3[0] ), .A3(
        \SB1_1_0/i1_5 ), .ZN(n2211) );
  XOR2_X1 U6703 ( .A1(\MC_ARK_ARC_1_2/temp3[11] ), .A2(
        \MC_ARK_ARC_1_2/temp4[11] ), .Z(n2212) );
  XOR2_X1 U6705 ( .A1(\MC_ARK_ARC_1_0/temp6[163] ), .A2(
        \MC_ARK_ARC_1_0/temp5[163] ), .Z(\MC_ARK_ARC_1_0/buf_output[163] ) );
  NAND3_X2 U6707 ( .A1(\SB1_1_19/i0_4 ), .A2(\SB1_1_19/i1[9] ), .A3(
        \SB1_1_19/i0_3 ), .ZN(\SB1_1_19/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U6709 ( .A1(\SB1_3_27/i0_0 ), .A2(\SB1_3_27/i3[0] ), .A3(
        \SB1_3_27/i1_7 ), .ZN(\SB1_3_27/Component_Function_4/NAND4_in[1] ) );
  NAND3_X2 U6711 ( .A1(\SB2_1_22/i0_3 ), .A2(\SB2_1_22/i0_4 ), .A3(
        \SB2_1_22/i1[9] ), .ZN(n2217) );
  INV_X2 U6715 ( .I(\SB1_1_23/buf_output[5] ), .ZN(\SB2_1_23/i1_5 ) );
  NAND3_X1 U6717 ( .A1(\SB1_3_27/i0_0 ), .A2(\SB1_3_27/i0[9] ), .A3(
        \SB1_3_27/i0[8] ), .ZN(n2221) );
  XOR2_X1 U6721 ( .A1(\MC_ARK_ARC_1_0/temp5[49] ), .A2(n2707), .Z(
        \MC_ARK_ARC_1_0/buf_output[49] ) );
  XOR2_X1 U6722 ( .A1(\MC_ARK_ARC_1_2/temp1[51] ), .A2(n2222), .Z(
        \MC_ARK_ARC_1_2/temp5[51] ) );
  XOR2_X1 U6723 ( .A1(n1390), .A2(\RI5[2][21] ), .Z(n2222) );
  NAND3_X2 U6725 ( .A1(\SB2_1_23/i0_0 ), .A2(\SB2_1_23/i0_4 ), .A3(
        \SB2_1_23/i1_5 ), .ZN(n2223) );
  NAND4_X2 U6727 ( .A1(\SB1_3_10/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_3_10/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_10/Component_Function_0/NAND4_in[3] ), .A4(
        \SB1_3_10/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_3_10/buf_output[0] ) );
  NAND3_X1 U6729 ( .A1(\SB1_1_15/i0[6] ), .A2(\SB1_1_15/i0_3 ), .A3(
        \SB1_1_15/i0[10] ), .ZN(\SB1_1_15/Component_Function_2/NAND4_in[1] )
         );
  XOR2_X1 U6730 ( .A1(\MC_ARK_ARC_1_0/temp1[55] ), .A2(
        \MC_ARK_ARC_1_0/temp2[55] ), .Z(n2409) );
  NAND3_X1 U6731 ( .A1(\SB4_13/i0[10] ), .A2(\SB4_13/i1_7 ), .A3(
        \SB4_13/i1[9] ), .ZN(n2228) );
  NAND3_X1 U6735 ( .A1(\RI1[4][155] ), .A2(\SB3_6/i0_0 ), .A3(\RI1[4][154] ), 
        .ZN(\SB3_6/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U6736 ( .A1(\SB1_1_12/i0[9] ), .A2(\SB1_1_12/i1_5 ), .A3(
        \SB1_1_12/i0[6] ), .ZN(\SB1_1_12/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U6738 ( .A1(\SB4_11/i0[6] ), .A2(\SB4_11/i0[8] ), .A3(
        \SB4_11/i0[7] ), .ZN(\SB4_11/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U6739 ( .A1(\MC_ARK_ARC_1_0/temp2[46] ), .A2(
        \MC_ARK_ARC_1_0/temp1[46] ), .Z(\MC_ARK_ARC_1_0/temp5[46] ) );
  XOR2_X1 U6741 ( .A1(n2460), .A2(n2233), .Z(\MC_ARK_ARC_1_0/buf_output[98] )
         );
  NAND3_X1 U6742 ( .A1(n5493), .A2(\SB2_1_15/i0[8] ), .A3(\SB2_1_15/i0[6] ), 
        .ZN(\SB2_1_15/Component_Function_0/NAND4_in[1] ) );
  BUF_X4 U6743 ( .I(\SB2_2_17/buf_output[0] ), .Z(\RI5[2][114] ) );
  NAND4_X2 U6744 ( .A1(\SB1_0_0/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_0_0/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_0_0/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_0_0/Component_Function_0/NAND4_in[0] ), .ZN(\SB2_0_27/i0[9] ) );
  INV_X1 U6755 ( .I(\SB3_19/buf_output[5] ), .ZN(\SB4_19/i1_5 ) );
  NAND4_X2 U6756 ( .A1(\SB3_19/Component_Function_5/NAND4_in[1] ), .A2(
        \SB3_19/Component_Function_5/NAND4_in[3] ), .A3(
        \SB3_19/Component_Function_5/NAND4_in[2] ), .A4(
        \SB3_19/Component_Function_5/NAND4_in[0] ), .ZN(\SB3_19/buf_output[5] ) );
  NAND3_X1 U6757 ( .A1(\SB4_4/i0_4 ), .A2(\SB4_4/i0[9] ), .A3(\SB4_4/i0[6] ), 
        .ZN(\SB4_4/Component_Function_5/NAND4_in[3] ) );
  BUF_X4 U6758 ( .I(\SB2_3_16/buf_output[0] ), .Z(\RI5[3][120] ) );
  NOR2_X2 U6760 ( .A1(n2244), .A2(n2243), .ZN(\SB2_3_26/i0[7] ) );
  NAND3_X2 U6765 ( .A1(\SB2_2_26/i0_0 ), .A2(\SB2_2_26/i1_5 ), .A3(
        \SB2_2_26/i0_4 ), .ZN(\SB2_2_26/Component_Function_2/NAND4_in[3] ) );
  INV_X2 U6766 ( .I(\RI3[0][129] ), .ZN(\SB2_0_10/i0[8] ) );
  XOR2_X1 U6769 ( .A1(\MC_ARK_ARC_1_0/temp3[44] ), .A2(
        \MC_ARK_ARC_1_0/temp4[44] ), .Z(n2359) );
  XOR2_X1 U6770 ( .A1(n2246), .A2(\MC_ARK_ARC_1_3/temp1[171] ), .Z(
        \MC_ARK_ARC_1_3/temp5[171] ) );
  XOR2_X1 U6771 ( .A1(\RI5[3][141] ), .A2(\RI5[3][117] ), .Z(n2246) );
  NAND3_X1 U6772 ( .A1(\SB1_1_20/i1_5 ), .A2(\SB1_1_20/i0_4 ), .A3(
        \SB1_1_20/i1[9] ), .ZN(\SB1_1_20/Component_Function_4/NAND4_in[3] ) );
  BUF_X4 U6774 ( .I(\SB2_3_10/buf_output[1] ), .Z(\RI5[3][151] ) );
  XOR2_X1 U6775 ( .A1(\MC_ARK_ARC_1_3/temp2[13] ), .A2(
        \MC_ARK_ARC_1_3/temp1[13] ), .Z(\MC_ARK_ARC_1_3/temp5[13] ) );
  NAND4_X2 U6778 ( .A1(\SB2_2_23/Component_Function_0/NAND4_in[1] ), .A2(n2523), .A3(n2524), .A4(\SB2_2_23/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_2_23/buf_output[0] ) );
  NAND4_X2 U6781 ( .A1(\SB2_3_6/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_3_6/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_3_6/Component_Function_0/NAND4_in[0] ), .A4(n2248), .ZN(
        \SB2_3_6/buf_output[0] ) );
  BUF_X4 U6782 ( .I(\SB2_3_5/buf_output[0] ), .Z(\RI5[3][186] ) );
  XOR2_X1 U6786 ( .A1(\MC_ARK_ARC_1_1/temp5[99] ), .A2(n2250), .Z(
        \MC_ARK_ARC_1_1/buf_output[99] ) );
  NAND3_X2 U6789 ( .A1(\SB2_3_10/i0_3 ), .A2(\SB2_3_10/i1[9] ), .A3(
        \SB2_3_10/i0_4 ), .ZN(\SB2_3_10/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U6791 ( .A1(\SB2_3_18/i1_5 ), .A2(\SB2_3_18/i3[0] ), .A3(
        \SB2_3_18/i0[8] ), .ZN(n2251) );
  NAND3_X1 U6795 ( .A1(\SB1_1_1/i0[8] ), .A2(\SB1_1_1/i0_3 ), .A3(
        \SB1_1_1/i1_7 ), .ZN(\SB1_1_1/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U6796 ( .A1(\SB4_31/i0_4 ), .A2(\SB4_31/i1[9] ), .A3(\SB4_31/i1_5 ), 
        .ZN(\SB4_31/Component_Function_4/NAND4_in[3] ) );
  AND2_X1 U6797 ( .A1(\SB1_0_3/Component_Function_3/NAND4_in[1] ), .A2(n2253), 
        .Z(n2710) );
  XOR2_X1 U6801 ( .A1(\RI5[0][189] ), .A2(\RI5[0][3] ), .Z(n2255) );
  NAND3_X2 U6804 ( .A1(\SB2_0_2/i0[8] ), .A2(\SB2_0_2/i3[0] ), .A3(
        \SB2_0_2/i1_5 ), .ZN(\SB2_0_2/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U6807 ( .A1(\SB1_2_29/i0_0 ), .A2(\SB1_2_29/i3[0] ), .A3(
        \SB1_2_29/i1_7 ), .ZN(n2257) );
  NAND3_X2 U6809 ( .A1(\SB1_3_3/i0[6] ), .A2(\SB1_3_3/i0[9] ), .A3(
        \SB1_3_3/i0_4 ), .ZN(n2258) );
  NAND4_X2 U6810 ( .A1(\SB1_1_31/Component_Function_3/NAND4_in[2] ), .A2(
        \SB1_1_31/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_31/Component_Function_3/NAND4_in[0] ), .A4(
        \SB1_1_31/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_1_31/buf_output[3] ) );
  XOR2_X1 U6811 ( .A1(\MC_ARK_ARC_1_3/temp5[98] ), .A2(
        \MC_ARK_ARC_1_3/temp6[98] ), .Z(\MC_ARK_ARC_1_3/buf_output[98] ) );
  NAND3_X1 U6815 ( .A1(\SB4_2/i0_3 ), .A2(\SB4_2/i0[10] ), .A3(\SB4_2/i0_4 ), 
        .ZN(\SB4_2/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U6819 ( .A1(\SB1_0_17/i0[10] ), .A2(\SB1_0_17/i1_5 ), .A3(
        \SB1_0_17/i1[9] ), .ZN(\SB1_0_17/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U6830 ( .A1(\MC_ARK_ARC_1_3/temp3[18] ), .A2(
        \MC_ARK_ARC_1_3/temp4[18] ), .Z(\MC_ARK_ARC_1_3/temp6[18] ) );
  NAND4_X2 U6831 ( .A1(\SB1_3_2/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_3_2/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_2/Component_Function_0/NAND4_in[0] ), .A4(n2263), .ZN(
        \SB1_3_2/buf_output[0] ) );
  NAND3_X1 U6832 ( .A1(\SB1_3_2/i0_0 ), .A2(\SB1_3_2/i0[7] ), .A3(
        \SB1_3_2/i0_3 ), .ZN(n2263) );
  XOR2_X1 U6834 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[86] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[92] ), .Z(n2266) );
  NAND3_X1 U6835 ( .A1(\SB4_14/i0[10] ), .A2(\SB4_14/i1[9] ), .A3(
        \SB4_14/i1_7 ), .ZN(n2267) );
  XOR2_X1 U6836 ( .A1(\MC_ARK_ARC_1_0/temp6[148] ), .A2(n2268), .Z(
        \MC_ARK_ARC_1_0/buf_output[148] ) );
  XOR2_X1 U6837 ( .A1(\MC_ARK_ARC_1_0/temp2[148] ), .A2(
        \MC_ARK_ARC_1_0/temp1[148] ), .Z(n2268) );
  BUF_X4 U6838 ( .I(\SB2_1_16/buf_output[0] ), .Z(\RI5[1][120] ) );
  XOR2_X1 U6841 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[180] ), .A2(\RI5[0][174] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[180] ) );
  XOR2_X1 U6842 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[165] ), .A2(\RI5[3][171] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[171] ) );
  BUF_X4 U6843 ( .I(\SB2_2_1/buf_output[0] ), .Z(\RI5[2][18] ) );
  NAND4_X2 U6847 ( .A1(\SB2_2_25/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_2_25/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_25/Component_Function_0/NAND4_in[3] ), .A4(
        \SB2_2_25/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_2_25/buf_output[0] ) );
  NAND3_X2 U6851 ( .A1(\SB2_0_22/i3[0] ), .A2(\SB2_0_22/i1_5 ), .A3(
        \SB2_0_22/i0[8] ), .ZN(n2274) );
  NAND3_X2 U6852 ( .A1(\SB2_2_23/i0_3 ), .A2(\SB2_2_23/i0[9] ), .A3(
        \SB2_2_23/i0[8] ), .ZN(\SB2_2_23/Component_Function_2/NAND4_in[2] ) );
  XOR2_X1 U6853 ( .A1(\RI5[3][66] ), .A2(\RI5[3][102] ), .Z(
        \MC_ARK_ARC_1_3/temp3[0] ) );
  XOR2_X1 U6854 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[58] ), .A2(\RI5[2][94] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[184] ) );
  BUF_X4 U6856 ( .I(\SB2_1_17/buf_output[0] ), .Z(\RI5[1][114] ) );
  XOR2_X1 U6857 ( .A1(\MC_ARK_ARC_1_1/temp2[168] ), .A2(
        \MC_ARK_ARC_1_1/temp1[168] ), .Z(\MC_ARK_ARC_1_1/temp5[168] ) );
  XOR2_X1 U6858 ( .A1(\MC_ARK_ARC_1_1/temp6[48] ), .A2(
        \MC_ARK_ARC_1_1/temp5[48] ), .Z(\MC_ARK_ARC_1_1/buf_output[48] ) );
  XOR2_X1 U6863 ( .A1(\RI5[0][95] ), .A2(\RI5[0][71] ), .Z(n2278) );
  NAND3_X1 U6864 ( .A1(\SB4_21/i0[10] ), .A2(\SB4_21/i0_3 ), .A3(
        \SB4_21/i0[6] ), .ZN(n2279) );
  NAND3_X1 U6865 ( .A1(\SB4_29/i0_0 ), .A2(\SB4_29/i0[9] ), .A3(\SB4_29/i0[8] ), .ZN(\SB4_29/Component_Function_4/NAND4_in[0] ) );
  BUF_X4 U6866 ( .I(\SB2_3_0/buf_output[1] ), .Z(\RI5[3][19] ) );
  NAND3_X1 U6867 ( .A1(\SB4_10/i0[6] ), .A2(\SB4_10/i0[8] ), .A3(
        \SB4_10/i0[7] ), .ZN(\SB4_10/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U6868 ( .A1(n2280), .A2(n181), .Z(Ciphertext[42]) );
  XOR2_X1 U6872 ( .A1(\MC_ARK_ARC_1_3/temp2[161] ), .A2(n2281), .Z(
        \MC_ARK_ARC_1_3/temp5[161] ) );
  NAND3_X2 U6880 ( .A1(\SB2_0_9/i1[9] ), .A2(\SB2_0_9/i0_3 ), .A3(
        \SB2_0_9/i0_4 ), .ZN(n2287) );
  XOR2_X1 U6881 ( .A1(\RI5[0][159] ), .A2(\RI5[0][3] ), .Z(
        \MC_ARK_ARC_1_0/temp3[93] ) );
  BUF_X4 U6884 ( .I(\SB2_1_9/buf_output[2] ), .Z(\RI5[1][152] ) );
  INV_X2 U6885 ( .I(\RI3[0][99] ), .ZN(\SB2_0_15/i0[8] ) );
  NAND4_X2 U6894 ( .A1(\SB1_1_16/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_1_16/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_1_16/Component_Function_0/NAND4_in[0] ), .A4(
        \SB1_1_16/Component_Function_0/NAND4_in[1] ), .ZN(
        \SB1_1_16/buf_output[0] ) );
  INV_X2 U6895 ( .I(n2291), .ZN(\MC_ARK_ARC_1_3/buf_output[113] ) );
  NAND4_X2 U6900 ( .A1(\SB1_3_27/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_3_27/Component_Function_0/NAND4_in[0] ), .A3(
        \SB1_3_27/Component_Function_0/NAND4_in[1] ), .A4(n2297), .ZN(
        \SB1_3_27/buf_output[0] ) );
  BUF_X4 U6901 ( .I(\SB2_1_0/buf_output[0] ), .Z(\RI5[1][24] ) );
  NAND2_X1 U6902 ( .A1(\SB1_3_23/i1[9] ), .A2(\SB1_3_23/i0_3 ), .ZN(
        \SB1_3_23/Component_Function_1/NAND4_in[0] ) );
  XOR2_X1 U6903 ( .A1(n2298), .A2(n71), .Z(Ciphertext[49]) );
  NAND3_X1 U6904 ( .A1(\SB2_3_0/i0_0 ), .A2(\SB1_3_1/buf_output[4] ), .A3(
        \SB2_3_0/i1_5 ), .ZN(n2300) );
  NAND3_X1 U6906 ( .A1(\SB1_3_19/i0_0 ), .A2(\SB1_3_19/i0_4 ), .A3(
        \SB1_3_19/i1_5 ), .ZN(n2301) );
  BUF_X4 U6909 ( .I(\SB2_2_18/buf_output[4] ), .Z(\RI5[2][88] ) );
  XOR2_X1 U6910 ( .A1(\MC_ARK_ARC_1_3/temp3[23] ), .A2(
        \MC_ARK_ARC_1_3/temp4[23] ), .Z(n2303) );
  XOR2_X1 U6917 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[68] ), .A2(\RI5[2][62] ), 
        .Z(n2308) );
  XOR2_X1 U6922 ( .A1(n2311), .A2(\MC_ARK_ARC_1_3/temp4[128] ), .Z(
        \MC_ARK_ARC_1_3/temp6[128] ) );
  XOR2_X1 U6923 ( .A1(\RI5[1][165] ), .A2(\RI5[1][141] ), .Z(
        \MC_ARK_ARC_1_1/temp2[3] ) );
  BUF_X4 U6924 ( .I(\SB2_3_7/buf_output[5] ), .Z(\RI5[3][149] ) );
  XOR2_X1 U6926 ( .A1(\RI5[0][142] ), .A2(\RI5[0][178] ), .Z(
        \MC_ARK_ARC_1_0/temp3[76] ) );
  NAND2_X1 U6930 ( .A1(\SB1_3_29/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_29/Component_Function_4/NAND4_in[1] ), .ZN(n2334) );
  NAND3_X1 U6933 ( .A1(n4762), .A2(\SB1_2_18/i3[0] ), .A3(\SB1_2_18/i1_5 ), 
        .ZN(n2318) );
  NAND4_X2 U6934 ( .A1(\SB3_28/Component_Function_3/NAND4_in[2] ), .A2(
        \SB3_28/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_28/Component_Function_3/NAND4_in[0] ), .A4(n2319), .ZN(
        \SB3_28/buf_output[3] ) );
  XOR2_X1 U6942 ( .A1(\RI5[2][154] ), .A2(\RI5[2][190] ), .Z(
        \MC_ARK_ARC_1_2/temp3[88] ) );
  NAND3_X1 U6946 ( .A1(\SB2_2_1/i0_0 ), .A2(\SB2_2_1/i3[0] ), .A3(
        \SB2_2_1/i1_7 ), .ZN(\SB2_2_1/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U6947 ( .A1(\MC_ARK_ARC_1_2/temp3[49] ), .A2(
        \MC_ARK_ARC_1_2/temp4[49] ), .Z(n2325) );
  BUF_X4 U6948 ( .I(\SB2_1_31/buf_output[4] ), .Z(\RI5[1][10] ) );
  XOR2_X1 U6951 ( .A1(\RI5[1][13] ), .A2(\RI5[1][49] ), .Z(
        \MC_ARK_ARC_1_1/temp3[139] ) );
  INV_X2 U6952 ( .I(\SB1_0_25/buf_output[2] ), .ZN(\SB2_0_22/i1[9] ) );
  NAND4_X2 U6954 ( .A1(\SB2_3_5/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_3_5/Component_Function_0/NAND4_in[1] ), .A3(n2397), .A4(
        \SB2_3_5/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_3_5/buf_output[0] ) );
  NAND3_X2 U6955 ( .A1(\SB3_30/i0_3 ), .A2(\SB3_30/i0_0 ), .A3(\SB3_30/i0_4 ), 
        .ZN(\SB3_30/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U6956 ( .A1(\SB2_0_6/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_0_6/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_0_6/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_6/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_0_6/buf_output[0] ) );
  NAND3_X2 U6957 ( .A1(\SB2_2_17/i0_3 ), .A2(\SB2_2_17/i1[9] ), .A3(
        \SB2_2_17/i0_4 ), .ZN(\SB2_2_17/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U6958 ( .A1(\SB1_0_16/i0_0 ), .A2(n290), .A3(\SB1_0_16/i0[8] ), 
        .ZN(n2327) );
  XOR2_X1 U6967 ( .A1(\MC_ARK_ARC_1_2/temp2[130] ), .A2(
        \MC_ARK_ARC_1_2/temp1[130] ), .Z(n2333) );
  BUF_X4 U6970 ( .I(\SB2_1_7/buf_output[4] ), .Z(\RI5[1][154] ) );
  XOR2_X1 U6971 ( .A1(\MC_ARK_ARC_1_1/temp6[160] ), .A2(
        \MC_ARK_ARC_1_1/temp5[160] ), .Z(\MC_ARK_ARC_1_1/buf_output[160] ) );
  NAND3_X1 U6972 ( .A1(n3993), .A2(\SB2_3_11/i0[8] ), .A3(\SB2_3_11/i0[6] ), 
        .ZN(\SB2_3_11/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U6977 ( .A1(n2338), .A2(n72), .Z(Ciphertext[173]) );
  NAND4_X2 U6978 ( .A1(\SB4_3/Component_Function_5/NAND4_in[1] ), .A2(
        \SB4_3/Component_Function_5/NAND4_in[2] ), .A3(
        \SB4_3/Component_Function_5/NAND4_in[3] ), .A4(
        \SB4_3/Component_Function_5/NAND4_in[0] ), .ZN(n2338) );
  BUF_X4 U6989 ( .I(\SB2_0_29/buf_output[5] ), .Z(\RI5[0][17] ) );
  XOR2_X1 U6991 ( .A1(\RI5[3][95] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[101] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[101] ) );
  BUF_X4 U6993 ( .I(\SB2_0_28/buf_output[5] ), .Z(\RI5[0][23] ) );
  NAND3_X1 U6995 ( .A1(\SB2_2_11/i0_3 ), .A2(\SB2_2_11/i0_0 ), .A3(
        \SB2_2_11/i0[7] ), .ZN(\SB2_2_11/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U6997 ( .A1(\SB3_5/buf_output[3] ), .A2(\SB4_3/i0_3 ), .A3(
        \SB4_3/i0_4 ), .ZN(\SB4_3/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U6999 ( .A1(\RI5[0][68] ), .A2(\RI5[0][74] ), .Z(n2344) );
  NAND4_X2 U7004 ( .A1(\SB1_1_18/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_1_18/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_1_18/Component_Function_3/NAND4_in[2] ), .A4(n2346), .ZN(
        \SB1_1_18/buf_output[3] ) );
  NAND3_X1 U7005 ( .A1(\SB1_1_18/i0[8] ), .A2(\SB1_1_18/i3[0] ), .A3(
        \SB1_1_18/i1_5 ), .ZN(n2346) );
  XOR2_X1 U7006 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[104] ), .A2(\RI5[3][140] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[38] ) );
  NAND3_X1 U7007 ( .A1(\SB4_27/i0[10] ), .A2(\SB4_27/i0_3 ), .A3(\SB4_27/i0_4 ), .ZN(\SB4_27/Component_Function_0/NAND4_in[2] ) );
  NAND4_X2 U7009 ( .A1(\SB1_2_19/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_2_19/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_2_19/Component_Function_4/NAND4_in[3] ), .A4(
        \SB1_2_19/Component_Function_4/NAND4_in[2] ), .ZN(
        \SB1_2_19/buf_output[4] ) );
  NAND4_X2 U7010 ( .A1(\SB1_2_20/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_20/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_20/Component_Function_4/NAND4_in[3] ), .A4(
        \SB1_2_20/Component_Function_4/NAND4_in[2] ), .ZN(
        \SB1_2_20/buf_output[4] ) );
  XOR2_X1 U7011 ( .A1(\MC_ARK_ARC_1_2/temp6[84] ), .A2(
        \MC_ARK_ARC_1_2/temp5[84] ), .Z(\MC_ARK_ARC_1_2/buf_output[84] ) );
  BUF_X4 U7013 ( .I(\SB2_1_21/buf_output[0] ), .Z(\RI5[1][90] ) );
  XOR2_X1 U7015 ( .A1(\MC_ARK_ARC_1_1/temp4[78] ), .A2(
        \MC_ARK_ARC_1_1/temp3[78] ), .Z(\MC_ARK_ARC_1_1/temp6[78] ) );
  XOR2_X1 U7017 ( .A1(n2776), .A2(\MC_ARK_ARC_1_0/temp6[96] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[96] ) );
  XOR2_X1 U7018 ( .A1(\MC_ARK_ARC_1_0/temp3[97] ), .A2(
        \MC_ARK_ARC_1_0/temp4[97] ), .Z(\MC_ARK_ARC_1_0/temp6[97] ) );
  BUF_X4 U7023 ( .I(\SB2_1_17/buf_output[2] ), .Z(\RI5[1][104] ) );
  XOR2_X1 U7026 ( .A1(n2352), .A2(\MC_ARK_ARC_1_3/temp1[31] ), .Z(n2475) );
  XOR2_X1 U7027 ( .A1(\RI5[3][169] ), .A2(\RI5[3][1] ), .Z(n2352) );
  BUF_X4 U7028 ( .I(\SB2_2_24/buf_output[0] ), .Z(\RI5[2][72] ) );
  XOR2_X1 U7031 ( .A1(\RI5[2][114] ), .A2(\RI5[2][150] ), .Z(
        \MC_ARK_ARC_1_2/temp3[48] ) );
  INV_X2 U7035 ( .I(\SB1_2_31/buf_output[3] ), .ZN(\SB2_2_29/i0[8] ) );
  NAND2_X1 U7037 ( .A1(\SB1_3_23/i0[9] ), .A2(\SB1_3_23/i0[10] ), .ZN(n2356)
         );
  NAND3_X1 U7038 ( .A1(\SB1_2_21/i0[10] ), .A2(\SB1_2_21/i1_5 ), .A3(
        \SB1_2_21/i1[9] ), .ZN(\SB1_2_21/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U7047 ( .A1(\RI5[3][171] ), .A2(\RI5[3][3] ), .Z(
        \MC_ARK_ARC_1_3/temp2[33] ) );
  BUF_X4 U7048 ( .I(\SB2_3_11/buf_output[2] ), .Z(\RI5[3][140] ) );
  NAND3_X1 U7049 ( .A1(\SB4_14/i0_3 ), .A2(\SB4_14/i1[9] ), .A3(\SB4_14/i0[6] ), .ZN(n2363) );
  BUF_X4 U7051 ( .I(\SB2_2_0/buf_output[5] ), .Z(\RI5[2][191] ) );
  XOR2_X1 U7052 ( .A1(\RI5[3][0] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[36] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[126] ) );
  XOR2_X1 U7053 ( .A1(\RI5[1][68] ), .A2(\RI5[1][104] ), .Z(
        \MC_ARK_ARC_1_1/temp3[2] ) );
  XOR2_X1 U7054 ( .A1(\MC_ARK_ARC_1_2/temp6[160] ), .A2(
        \MC_ARK_ARC_1_2/temp5[160] ), .Z(\MC_ARK_ARC_1_2/buf_output[160] ) );
  BUF_X4 U7055 ( .I(\SB2_3_29/buf_output[1] ), .Z(\RI5[3][37] ) );
  BUF_X4 U7056 ( .I(\SB2_1_28/buf_output[0] ), .Z(\RI5[1][48] ) );
  NAND4_X2 U7059 ( .A1(\SB2_0_22/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_0_22/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_0_22/Component_Function_0/NAND4_in[0] ), .A4(n2366), .ZN(
        \SB2_0_22/buf_output[0] ) );
  BUF_X4 U7070 ( .I(\SB2_2_28/buf_output[4] ), .Z(\RI5[2][28] ) );
  NAND3_X1 U7071 ( .A1(\SB2_1_6/i0_3 ), .A2(\SB2_1_6/i0[10] ), .A3(
        \SB2_1_6/i0[9] ), .ZN(\SB2_1_6/Component_Function_4/NAND4_in[2] ) );
  XOR2_X1 U7078 ( .A1(\MC_ARK_ARC_1_0/temp5[166] ), .A2(n2375), .Z(
        \MC_ARK_ARC_1_0/buf_output[166] ) );
  XOR2_X1 U7079 ( .A1(\MC_ARK_ARC_1_0/temp3[166] ), .A2(
        \MC_ARK_ARC_1_0/temp4[166] ), .Z(n2375) );
  BUF_X4 U7083 ( .I(\SB2_1_24/buf_output[0] ), .Z(\RI5[1][72] ) );
  XOR2_X1 U7086 ( .A1(\RI5[0][57] ), .A2(\RI5[0][93] ), .Z(
        \MC_ARK_ARC_1_0/temp3[183] ) );
  NAND4_X2 U7087 ( .A1(\SB2_3_30/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_30/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_3_30/Component_Function_4/NAND4_in[2] ), .A4(n2382), .ZN(
        \SB2_3_30/buf_output[4] ) );
  XOR2_X1 U7089 ( .A1(n2383), .A2(n57), .Z(Ciphertext[71]) );
  NAND4_X2 U7090 ( .A1(\SB4_20/Component_Function_5/NAND4_in[2] ), .A2(
        \SB4_20/Component_Function_5/NAND4_in[3] ), .A3(n2436), .A4(
        \SB4_20/Component_Function_5/NAND4_in[0] ), .ZN(n2383) );
  NAND3_X2 U7092 ( .A1(\SB3_21/i0_3 ), .A2(\SB3_21/i0_0 ), .A3(\SB3_21/i0_4 ), 
        .ZN(\SB3_21/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U7099 ( .A1(\MC_ARK_ARC_1_1/temp4[91] ), .A2(
        \MC_ARK_ARC_1_1/temp3[91] ), .Z(n2388) );
  XOR2_X1 U7102 ( .A1(\MC_ARK_ARC_1_2/temp3[31] ), .A2(
        \MC_ARK_ARC_1_2/temp4[31] ), .Z(n2389) );
  NAND3_X1 U7103 ( .A1(\SB4_6/i0[6] ), .A2(n579), .A3(\SB4_6/i0[7] ), .ZN(
        \SB4_6/Component_Function_0/NAND4_in[1] ) );
  BUF_X4 U7104 ( .I(\SB2_1_19/buf_output[4] ), .Z(\RI5[1][82] ) );
  XOR2_X1 U7106 ( .A1(\MC_ARK_ARC_1_1/temp4[46] ), .A2(
        \MC_ARK_ARC_1_1/temp3[46] ), .Z(n2390) );
  XOR2_X1 U7109 ( .A1(\MC_ARK_ARC_1_0/temp6[15] ), .A2(
        \MC_ARK_ARC_1_0/temp5[15] ), .Z(\MC_ARK_ARC_1_0/buf_output[15] ) );
  NAND3_X1 U7110 ( .A1(\SB4_20/i0[10] ), .A2(\SB4_20/i0_3 ), .A3(
        \SB4_20/i0[6] ), .ZN(\SB4_20/Component_Function_2/NAND4_in[1] ) );
  XOR2_X1 U7115 ( .A1(n2623), .A2(\MC_ARK_ARC_1_2/temp5[127] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[127] ) );
  NAND4_X2 U7117 ( .A1(\SB1_2_23/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_23/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_2_23/Component_Function_5/NAND4_in[3] ), .A4(
        \SB1_2_23/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_2_23/buf_output[5] ) );
  NAND3_X1 U7123 ( .A1(\SB1_1_22/i0[8] ), .A2(\SB1_1_22/i1_7 ), .A3(
        \SB1_1_22/i0_4 ), .ZN(n2728) );
  BUF_X4 U7127 ( .I(\SB2_1_28/buf_output[5] ), .Z(\RI5[1][23] ) );
  BUF_X4 U7130 ( .I(\SB2_1_11/buf_output[5] ), .Z(\RI5[1][125] ) );
  NOR2_X2 U7131 ( .A1(n2403), .A2(n2401), .ZN(n2711) );
  NAND3_X1 U7132 ( .A1(\SB1_0_18/i0_0 ), .A2(\SB1_0_18/i0[7] ), .A3(
        \SB1_0_18/i0_3 ), .ZN(n2404) );
  NAND3_X1 U7133 ( .A1(\SB4_12/i0[10] ), .A2(\SB4_12/i0_3 ), .A3(
        \SB4_12/i0[6] ), .ZN(n2406) );
  XOR2_X1 U7134 ( .A1(\MC_ARK_ARC_1_3/temp3[135] ), .A2(
        \MC_ARK_ARC_1_3/temp4[135] ), .Z(\MC_ARK_ARC_1_3/temp6[135] ) );
  XOR2_X1 U7142 ( .A1(n2410), .A2(\MC_ARK_ARC_1_2/temp5[100] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[100] ) );
  XOR2_X1 U7143 ( .A1(\MC_ARK_ARC_1_2/temp4[100] ), .A2(
        \MC_ARK_ARC_1_2/temp3[100] ), .Z(n2410) );
  BUF_X4 U7145 ( .I(\SB2_1_19/buf_output[0] ), .Z(\RI5[1][102] ) );
  NAND3_X1 U7146 ( .A1(\SB4_23/i0_0 ), .A2(\SB4_23/i1_7 ), .A3(\SB4_23/i3[0] ), 
        .ZN(n2705) );
  XOR2_X1 U7147 ( .A1(\MC_ARK_ARC_1_2/temp5[178] ), .A2(
        \MC_ARK_ARC_1_2/temp6[178] ), .Z(\MC_ARK_ARC_1_2/buf_output[178] ) );
  BUF_X4 U7148 ( .I(\SB2_2_4/buf_output[4] ), .Z(\RI5[2][172] ) );
  NAND3_X2 U7152 ( .A1(\SB2_3_7/i1_7 ), .A2(\SB2_3_7/i0[10] ), .A3(
        \SB2_3_7/i1[9] ), .ZN(\SB2_3_7/Component_Function_3/NAND4_in[2] ) );
  BUF_X4 U7158 ( .I(\SB2_1_20/buf_output[3] ), .Z(\RI5[1][81] ) );
  BUF_X4 U7162 ( .I(\SB2_1_0/buf_output[4] ), .Z(\RI5[1][4] ) );
  NAND4_X2 U7163 ( .A1(\SB1_1_1/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_1_1/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_1/Component_Function_1/NAND4_in[0] ), .A4(n2416), .ZN(
        \SB1_1_1/buf_output[1] ) );
  XOR2_X1 U7164 ( .A1(\MC_ARK_ARC_1_1/temp6[108] ), .A2(n2418), .Z(
        \MC_ARK_ARC_1_1/buf_output[108] ) );
  BUF_X4 U7166 ( .I(\SB2_2_15/buf_output[3] ), .Z(\RI5[2][111] ) );
  NAND3_X1 U7168 ( .A1(\SB1_2_21/i0_3 ), .A2(\SB1_2_21/i1[9] ), .A3(
        \SB1_2_21/i0[6] ), .ZN(\SB1_2_21/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U7169 ( .A1(\SB4_26/i0[10] ), .A2(\SB4_26/i1[9] ), .A3(
        \SB4_26/i1_7 ), .ZN(n2419) );
  XOR2_X1 U7171 ( .A1(\MC_ARK_ARC_1_3/temp4[99] ), .A2(n2421), .Z(
        \MC_ARK_ARC_1_3/temp6[99] ) );
  XOR2_X1 U7172 ( .A1(\RI5[3][9] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[165] ), 
        .Z(n2421) );
  AND3_X1 U7176 ( .A1(\SB1_1_30/i1[9] ), .A2(\SB1_1_30/i1_5 ), .A3(
        \SB1_1_30/i0_4 ), .Z(n2884) );
  NOR2_X2 U7177 ( .A1(n2425), .A2(n2423), .ZN(n2877) );
  INV_X2 U7178 ( .I(n2426), .ZN(\RI1[3][143] ) );
  XNOR2_X1 U7179 ( .A1(\MC_ARK_ARC_1_2/temp6[143] ), .A2(
        \MC_ARK_ARC_1_2/temp5[143] ), .ZN(n2426) );
  XOR2_X1 U7181 ( .A1(\MC_ARK_ARC_1_3/temp3[94] ), .A2(
        \MC_ARK_ARC_1_3/temp4[94] ), .Z(n2427) );
  NAND4_X2 U7186 ( .A1(\SB1_3_23/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_3_23/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_23/Component_Function_1/NAND4_in[0] ), .A4(n2430), .ZN(
        \SB1_3_23/buf_output[1] ) );
  XOR2_X1 U7192 ( .A1(\RI5[0][118] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[112] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[118] ) );
  XOR2_X1 U7194 ( .A1(\RI5[1][129] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[153] ), 
        .Z(n2434) );
  INV_X2 U7200 ( .I(\RI3[0][69] ), .ZN(\SB2_0_20/i0[8] ) );
  NAND4_X2 U7202 ( .A1(\SB2_1_19/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_1_19/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_19/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_19/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_1_19/buf_output[0] ) );
  XOR2_X1 U7203 ( .A1(\RI5[3][131] ), .A2(\RI5[3][125] ), .Z(
        \MC_ARK_ARC_1_3/temp1[131] ) );
  NAND3_X1 U7207 ( .A1(\SB2_1_15/i0_4 ), .A2(\SB2_1_15/i0[8] ), .A3(
        \SB2_1_15/i1_7 ), .ZN(\SB2_1_15/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U7208 ( .A1(\SB1_0_12/i0_0 ), .A2(\SB1_0_12/i3[0] ), .A3(
        \SB1_0_12/i1_7 ), .ZN(\SB1_0_12/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U7211 ( .A1(\SB1_2_16/i0[6] ), .A2(\SB1_2_16/i0[8] ), .A3(
        \SB1_2_16/i0[7] ), .ZN(n2446) );
  XOR2_X1 U7212 ( .A1(n2447), .A2(n2448), .Z(\MC_ARK_ARC_1_0/buf_output[114] )
         );
  XOR2_X1 U7213 ( .A1(\MC_ARK_ARC_1_0/temp3[114] ), .A2(
        \MC_ARK_ARC_1_0/temp1[114] ), .Z(n2447) );
  XOR2_X1 U7214 ( .A1(\RI5[1][91] ), .A2(\RI5[1][85] ), .Z(
        \MC_ARK_ARC_1_1/temp1[91] ) );
  XOR2_X1 U7215 ( .A1(n2450), .A2(n127), .Z(Ciphertext[145]) );
  XOR2_X1 U7218 ( .A1(\MC_ARK_ARC_1_0/temp1[121] ), .A2(
        \MC_ARK_ARC_1_0/temp4[121] ), .Z(n2452) );
  NAND3_X2 U7219 ( .A1(\SB2_3_13/i0[10] ), .A2(\SB2_3_13/i0_0 ), .A3(
        \SB2_3_13/i0[6] ), .ZN(n2454) );
  NAND2_X1 U7220 ( .A1(\SB4_10/i0_3 ), .A2(n3653), .ZN(n2456) );
  NAND4_X2 U7226 ( .A1(\SB1_0_14/Component_Function_3/NAND4_in[2] ), .A2(
        \SB1_0_14/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_14/Component_Function_3/NAND4_in[3] ), .A4(
        \SB1_0_14/Component_Function_3/NAND4_in[0] ), .ZN(
        \SB1_0_14/buf_output[3] ) );
  XOR2_X1 U7227 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[14] ), .A2(\RI5[3][170] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[104] ) );
  NAND3_X2 U7229 ( .A1(\SB1_1_18/i0_4 ), .A2(\SB1_1_18/i1[9] ), .A3(
        \SB1_1_18/i0_3 ), .ZN(\SB1_1_18/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U7239 ( .A1(\MC_ARK_ARC_1_1/temp2[125] ), .A2(
        \MC_ARK_ARC_1_1/temp1[125] ), .Z(n2462) );
  XOR2_X1 U7240 ( .A1(n2463), .A2(n140), .Z(Ciphertext[39]) );
  NAND4_X2 U7241 ( .A1(\SB4_25/Component_Function_3/NAND4_in[3] ), .A2(
        \SB4_25/Component_Function_3/NAND4_in[1] ), .A3(
        \SB4_25/Component_Function_3/NAND4_in[2] ), .A4(n2829), .ZN(n2463) );
  XOR2_X1 U7242 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[56] ), .A2(\RI5[3][32] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[86] ) );
  XOR2_X1 U7246 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[105] ), .A2(\RI5[1][111] ), 
        .Z(n2467) );
  XOR2_X1 U7248 ( .A1(\MC_ARK_ARC_1_2/temp3[188] ), .A2(
        \MC_ARK_ARC_1_2/temp4[188] ), .Z(n2470) );
  BUF_X4 U7249 ( .I(\SB2_1_4/buf_output[5] ), .Z(\RI5[1][167] ) );
  INV_X2 U7250 ( .I(\SB1_1_16/buf_output[5] ), .ZN(\SB2_1_16/i1_5 ) );
  NAND3_X1 U7251 ( .A1(\SB2_2_21/i0_3 ), .A2(\SB2_2_21/i0[10] ), .A3(
        \SB2_2_21/i0[9] ), .ZN(n2473) );
  NAND3_X1 U7253 ( .A1(\SB4_20/i0_0 ), .A2(\SB4_20/i0_3 ), .A3(\SB4_20/i0[7] ), 
        .ZN(\SB4_20/Component_Function_0/NAND4_in[3] ) );
  INV_X1 U7255 ( .I(\SB3_26/buf_output[1] ), .ZN(\SB4_22/i1_7 ) );
  NAND4_X2 U7256 ( .A1(\SB3_26/Component_Function_1/NAND4_in[2] ), .A2(
        \SB3_26/Component_Function_1/NAND4_in[3] ), .A3(
        \SB3_26/Component_Function_1/NAND4_in[0] ), .A4(
        \SB3_26/Component_Function_1/NAND4_in[1] ), .ZN(\SB3_26/buf_output[1] ) );
  XOR2_X1 U7258 ( .A1(\MC_ARK_ARC_1_2/temp2[180] ), .A2(
        \MC_ARK_ARC_1_2/temp1[180] ), .Z(\MC_ARK_ARC_1_2/temp5[180] ) );
  NAND4_X2 U7264 ( .A1(\SB1_0_1/Component_Function_2/NAND4_in[3] ), .A2(
        \SB1_0_1/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_0_1/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_1/Component_Function_2/NAND4_in[1] ), .ZN(\RI3[0][8] ) );
  XOR2_X1 U7265 ( .A1(\MC_ARK_ARC_1_1/temp5[169] ), .A2(n2823), .Z(
        \MC_ARK_ARC_1_1/buf_output[169] ) );
  NOR2_X2 U7268 ( .A1(n2483), .A2(n2481), .ZN(n2753) );
  NAND4_X2 U7271 ( .A1(\SB3_28/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_28/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_28/Component_Function_0/NAND4_in[0] ), .A4(n2484), .ZN(
        \SB3_28/buf_output[0] ) );
  XOR2_X1 U7272 ( .A1(\MC_ARK_ARC_1_0/temp5[4] ), .A2(
        \MC_ARK_ARC_1_0/temp6[4] ), .Z(\MC_ARK_ARC_1_0/buf_output[4] ) );
  XOR2_X1 U7275 ( .A1(\MC_ARK_ARC_1_1/temp3[0] ), .A2(
        \MC_ARK_ARC_1_1/temp4[0] ), .Z(\MC_ARK_ARC_1_1/temp6[0] ) );
  NAND3_X1 U7276 ( .A1(\SB1_0_2/i1_5 ), .A2(\SB1_0_2/i1[9] ), .A3(n400), .ZN(
        \SB1_0_2/Component_Function_4/NAND4_in[3] ) );
  XOR2_X1 U7282 ( .A1(\MC_ARK_ARC_1_3/temp5[69] ), .A2(
        \MC_ARK_ARC_1_3/temp6[69] ), .Z(\MC_ARK_ARC_1_3/buf_output[69] ) );
  NAND4_X2 U7283 ( .A1(\SB1_3_13/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_3_13/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_3_13/Component_Function_0/NAND4_in[0] ), .A4(n2492), .ZN(
        \SB1_3_13/buf_output[0] ) );
  XOR2_X1 U7288 ( .A1(\MC_ARK_ARC_1_1/temp5[51] ), .A2(
        \MC_ARK_ARC_1_1/temp6[51] ), .Z(\MC_ARK_ARC_1_1/buf_output[51] ) );
  XOR2_X1 U7289 ( .A1(\MC_ARK_ARC_1_2/temp5[12] ), .A2(n2496), .Z(
        \MC_ARK_ARC_1_2/buf_output[12] ) );
  XOR2_X1 U7291 ( .A1(\MC_ARK_ARC_1_0/temp2[157] ), .A2(
        \MC_ARK_ARC_1_0/temp4[157] ), .Z(n2500) );
  BUF_X4 U7292 ( .I(\SB2_1_4/buf_output[0] ), .Z(\RI5[1][0] ) );
  XOR2_X1 U7296 ( .A1(\RI5[1][188] ), .A2(n120), .Z(n2502) );
  XOR2_X1 U7304 ( .A1(\MC_ARK_ARC_1_0/temp5[165] ), .A2(n2509), .Z(
        \MC_ARK_ARC_1_0/buf_output[165] ) );
  XOR2_X1 U7308 ( .A1(n2511), .A2(\MC_ARK_ARC_1_0/temp5[168] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[168] ) );
  XOR2_X1 U7309 ( .A1(\MC_ARK_ARC_1_0/temp4[168] ), .A2(
        \MC_ARK_ARC_1_0/temp3[168] ), .Z(n2511) );
  BUF_X4 U7313 ( .I(\SB2_3_23/buf_output[3] ), .Z(\RI5[3][63] ) );
  NAND3_X1 U7322 ( .A1(\SB4_31/i0_0 ), .A2(\SB4_31/i1_5 ), .A3(\SB4_31/i0_4 ), 
        .ZN(n2519) );
  BUF_X4 U7323 ( .I(\SB2_2_13/buf_output[0] ), .Z(\RI5[2][138] ) );
  INV_X2 U7325 ( .I(\SB1_1_29/buf_output[3] ), .ZN(\SB2_1_27/i0[8] ) );
  NAND4_X2 U7326 ( .A1(\SB1_1_29/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_29/Component_Function_3/NAND4_in[2] ), .A3(
        \SB1_1_29/Component_Function_3/NAND4_in[1] ), .A4(
        \SB1_1_29/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_1_29/buf_output[3] ) );
  XOR2_X1 U7327 ( .A1(n2525), .A2(\MC_ARK_ARC_1_2/temp5[102] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[102] ) );
  XOR2_X1 U7328 ( .A1(\MC_ARK_ARC_1_2/temp3[102] ), .A2(
        \MC_ARK_ARC_1_2/temp4[102] ), .Z(n2525) );
  INV_X2 U7329 ( .I(\SB1_2_23/buf_output[2] ), .ZN(\SB2_2_20/i1[9] ) );
  NAND3_X2 U7331 ( .A1(\SB1_2_30/i0[10] ), .A2(\SB1_2_30/i0[9] ), .A3(
        \SB1_2_30/i0_3 ), .ZN(n2526) );
  XOR2_X1 U7335 ( .A1(\SB2_3_19/buf_output[2] ), .A2(n210), .Z(n2530) );
  NAND3_X2 U7345 ( .A1(\SB2_0_2/i1[9] ), .A2(\SB2_0_2/i0_3 ), .A3(
        \RI3[0][178] ), .ZN(\SB2_0_2/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U7349 ( .A1(\MC_ARK_ARC_1_1/temp2[156] ), .A2(
        \MC_ARK_ARC_1_1/temp1[156] ), .Z(\MC_ARK_ARC_1_1/temp5[156] ) );
  NAND4_X2 U7350 ( .A1(\SB1_0_28/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_0_28/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_0_28/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_0_28/Component_Function_0/NAND4_in[0] ), .ZN(\RI3[0][48] ) );
  BUF_X4 U7352 ( .I(\SB2_1_22/buf_output[3] ), .Z(\RI5[1][69] ) );
  NAND4_X2 U7355 ( .A1(\SB2_1_7/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_1_7/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_1_7/Component_Function_4/NAND4_in[1] ), .A4(n2545), .ZN(
        \SB2_1_7/buf_output[4] ) );
  XOR2_X1 U7356 ( .A1(\RI5[3][159] ), .A2(\RI5[3][3] ), .Z(n2547) );
  XOR2_X1 U7357 ( .A1(n2548), .A2(\MC_ARK_ARC_1_3/temp6[16] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[16] ) );
  NAND4_X2 U7362 ( .A1(\SB1_0_3/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_0_3/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_0_3/Component_Function_1/NAND4_in[1] ), .A4(
        \SB1_0_3/Component_Function_1/NAND4_in[0] ), .ZN(\RI3[0][1] ) );
  NAND4_X2 U7365 ( .A1(\SB1_2_8/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_2_8/Component_Function_3/NAND4_in[0] ), .A3(n2796), .A4(
        \SB1_2_8/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_2_8/buf_output[3] ) );
  XOR2_X1 U7369 ( .A1(n2551), .A2(\MC_ARK_ARC_1_3/temp1[115] ), .Z(
        \MC_ARK_ARC_1_3/temp5[115] ) );
  XOR2_X1 U7370 ( .A1(\RI5[3][61] ), .A2(\RI5[3][85] ), .Z(n2551) );
  XOR2_X1 U7371 ( .A1(\MC_ARK_ARC_1_2/temp1[121] ), .A2(
        \MC_ARK_ARC_1_2/temp2[121] ), .Z(\MC_ARK_ARC_1_2/temp5[121] ) );
  XOR2_X1 U7377 ( .A1(\RI5[0][174] ), .A2(\RI5[0][18] ), .Z(
        \MC_ARK_ARC_1_0/temp3[108] ) );
  BUF_X4 U7378 ( .I(\SB2_1_8/buf_output[4] ), .Z(\RI5[1][148] ) );
  BUF_X4 U7379 ( .I(\SB2_3_28/buf_output[0] ), .Z(\RI5[3][48] ) );
  XOR2_X1 U7382 ( .A1(\RI5[2][135] ), .A2(\RI5[2][111] ), .Z(
        \MC_ARK_ARC_1_2/temp2[165] ) );
  BUF_X4 U7384 ( .I(\SB2_2_6/buf_output[5] ), .Z(\RI5[2][155] ) );
  NAND3_X1 U7386 ( .A1(\SB1_1_24/i0_4 ), .A2(\SB1_1_24/i1_7 ), .A3(
        \SB1_1_24/i0[8] ), .ZN(\SB1_1_24/Component_Function_1/NAND4_in[3] ) );
  XOR2_X1 U7387 ( .A1(n2562), .A2(n2561), .Z(\MC_ARK_ARC_1_3/buf_output[170] )
         );
  XOR2_X1 U7388 ( .A1(\MC_ARK_ARC_1_3/temp4[170] ), .A2(
        \MC_ARK_ARC_1_3/temp2[170] ), .Z(n2561) );
  NAND4_X2 U7392 ( .A1(\SB3_3/Component_Function_4/NAND4_in[1] ), .A2(
        \SB3_3/Component_Function_4/NAND4_in[0] ), .A3(
        \SB3_3/Component_Function_4/NAND4_in[3] ), .A4(n2567), .ZN(
        \SB3_3/buf_output[4] ) );
  NAND3_X1 U7393 ( .A1(\SB3_3/i0_3 ), .A2(\SB3_3/i0[10] ), .A3(\SB3_3/i0[9] ), 
        .ZN(n2567) );
  NAND3_X1 U7395 ( .A1(\SB4_19/i0_4 ), .A2(\SB4_19/i0[9] ), .A3(\SB4_19/i0[6] ), .ZN(\SB4_19/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U7396 ( .A1(\SB4_2/i0_4 ), .A2(\SB4_2/i1_7 ), .A3(\SB4_2/i0[8] ), 
        .ZN(n2569) );
  XOR2_X1 U7400 ( .A1(\MC_ARK_ARC_1_1/temp6[19] ), .A2(
        \MC_ARK_ARC_1_1/temp5[19] ), .Z(\MC_ARK_ARC_1_1/buf_output[19] ) );
  XOR2_X1 U7401 ( .A1(\RI5[3][134] ), .A2(\RI5[3][98] ), .Z(
        \MC_ARK_ARC_1_3/temp3[32] ) );
  XOR2_X1 U7404 ( .A1(\RI5[2][155] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[131] ), 
        .Z(n2574) );
  BUF_X4 U7406 ( .I(\SB2_1_30/buf_output[0] ), .Z(\RI5[1][36] ) );
  NAND3_X1 U7407 ( .A1(\SB1_0_15/i0_3 ), .A2(\SB1_0_15/i0[7] ), .A3(
        \SB1_0_15/i0_0 ), .ZN(\SB1_0_15/Component_Function_0/NAND4_in[3] ) );
  XOR2_X1 U7409 ( .A1(\MC_ARK_ARC_1_0/temp3[49] ), .A2(
        \MC_ARK_ARC_1_0/temp4[49] ), .Z(n2707) );
  NAND3_X1 U7410 ( .A1(\SB4_27/i0[9] ), .A2(\SB4_27/i1_5 ), .A3(\SB4_27/i0[6] ), .ZN(\SB4_27/Component_Function_1/NAND4_in[2] ) );
  BUF_X4 U7412 ( .I(\SB2_1_31/buf_output[3] ), .Z(\RI5[1][15] ) );
  NAND3_X1 U7413 ( .A1(\SB4_2/i0[6] ), .A2(\SB4_2/i0_4 ), .A3(\SB4_2/i0[9] ), 
        .ZN(\SB4_2/Component_Function_5/NAND4_in[3] ) );
  BUF_X4 U7417 ( .I(\SB2_1_11/buf_output[0] ), .Z(\RI5[1][150] ) );
  NAND4_X2 U7418 ( .A1(\SB2_2_13/Component_Function_5/NAND4_in[1] ), .A2(
        \SB2_2_13/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_2_13/Component_Function_5/NAND4_in[2] ), .A4(
        \SB2_2_13/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_2_13/buf_output[5] ) );
  NAND3_X1 U7420 ( .A1(\SB1_1_12/i0_4 ), .A2(\SB1_1_12/i1[9] ), .A3(
        \SB1_1_12/i1_5 ), .ZN(n2581) );
  BUF_X4 U7421 ( .I(\SB2_1_20/buf_output[4] ), .Z(\RI5[1][76] ) );
  NAND4_X2 U7422 ( .A1(\SB1_1_23/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_1_23/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_1_23/Component_Function_1/NAND4_in[0] ), .A4(n2582), .ZN(
        \SB1_1_23/buf_output[1] ) );
  XOR2_X1 U7423 ( .A1(\MC_ARK_ARC_1_1/temp6[138] ), .A2(
        \MC_ARK_ARC_1_1/temp5[138] ), .Z(\MC_ARK_ARC_1_1/buf_output[138] ) );
  XOR2_X1 U7430 ( .A1(\MC_ARK_ARC_1_1/temp2[60] ), .A2(
        \MC_ARK_ARC_1_1/temp1[60] ), .Z(n2587) );
  NAND3_X1 U7431 ( .A1(n2899), .A2(\SB1_0_17/i1_7 ), .A3(\SB1_0_17/i0[8] ), 
        .ZN(\SB1_0_17/Component_Function_1/NAND4_in[3] ) );
  BUF_X2 U7437 ( .I(\SB2_0_7/i0[6] ), .Z(n2593) );
  XOR2_X1 U7442 ( .A1(\MC_ARK_ARC_1_1/temp3[63] ), .A2(
        \MC_ARK_ARC_1_1/temp4[63] ), .Z(n2596) );
  XOR2_X1 U7444 ( .A1(\MC_ARK_ARC_1_3/temp2[109] ), .A2(
        \MC_ARK_ARC_1_3/temp1[109] ), .Z(n2597) );
  BUF_X4 U7445 ( .I(\SB2_3_26/buf_output[1] ), .Z(\RI5[3][55] ) );
  INV_X2 U7448 ( .I(\RI3[0][3] ), .ZN(\SB2_0_31/i0[8] ) );
  NAND3_X1 U7452 ( .A1(\SB2_3_13/i0_0 ), .A2(\SB2_3_13/i0_3 ), .A3(
        \SB2_3_13/i0[7] ), .ZN(\SB2_3_13/Component_Function_0/NAND4_in[3] ) );
  NOR2_X2 U7453 ( .A1(n2602), .A2(n2601), .ZN(\SB2_3_13/i0[7] ) );
  XOR2_X1 U7457 ( .A1(\MC_ARK_ARC_1_1/temp3[130] ), .A2(
        \MC_ARK_ARC_1_1/temp4[130] ), .Z(n2603) );
  BUF_X2 U7459 ( .I(\SB2_0_29/i0[9] ), .Z(n2605) );
  NAND3_X2 U7461 ( .A1(\SB3_21/i0_3 ), .A2(\SB3_21/i1[9] ), .A3(\SB3_21/i0_4 ), 
        .ZN(n2606) );
  NAND3_X1 U7463 ( .A1(\SB4_13/i0_4 ), .A2(\SB4_13/i1_7 ), .A3(n3683), .ZN(
        n2607) );
  XOR2_X1 U7465 ( .A1(\MC_ARK_ARC_1_0/temp2[179] ), .A2(
        \MC_ARK_ARC_1_0/temp1[179] ), .Z(\MC_ARK_ARC_1_0/temp5[179] ) );
  BUF_X4 U7466 ( .I(\SB2_2_6/buf_output[4] ), .Z(\RI5[2][160] ) );
  XOR2_X1 U7471 ( .A1(\MC_ARK_ARC_1_3/temp5[182] ), .A2(n2610), .Z(
        \MC_ARK_ARC_1_3/buf_output[182] ) );
  BUF_X4 U7473 ( .I(\SB2_2_21/buf_output[0] ), .Z(\RI5[2][90] ) );
  XOR2_X1 U7475 ( .A1(\MC_ARK_ARC_1_3/temp6[60] ), .A2(
        \MC_ARK_ARC_1_3/temp5[60] ), .Z(\MC_ARK_ARC_1_3/buf_output[60] ) );
  XOR2_X1 U7477 ( .A1(\RI5[2][188] ), .A2(\RI5[2][20] ), .Z(n2611) );
  NAND3_X1 U7480 ( .A1(\SB1_0_20/i1_5 ), .A2(\SB1_0_20/i0_4 ), .A3(
        \SB1_0_20/i1[9] ), .ZN(n2613) );
  NAND3_X2 U7481 ( .A1(\SB2_3_23/i0_3 ), .A2(\SB2_3_23/i1[9] ), .A3(
        \SB2_3_23/i0_4 ), .ZN(n2615) );
  INV_X2 U7482 ( .I(\SB2_1_21/i3[0] ), .ZN(\RI3[1][60] ) );
  NOR2_X2 U7484 ( .A1(n2617), .A2(n2616), .ZN(\SB2_1_21/i3[0] ) );
  NAND4_X2 U7486 ( .A1(\SB1_0_22/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_0_22/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_0_22/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_0_22/Component_Function_0/NAND4_in[0] ), .ZN(\RI3[0][84] ) );
  BUF_X4 U7487 ( .I(\SB2_2_13/buf_output[5] ), .Z(\RI5[2][113] ) );
  XOR2_X1 U7489 ( .A1(\RI5[3][20] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[56] ), 
        .Z(n2620) );
  BUF_X4 U7490 ( .I(\SB2_1_26/buf_output[0] ), .Z(\RI5[1][60] ) );
  XOR2_X1 U7491 ( .A1(\RI5[1][175] ), .A2(\RI5[1][19] ), .Z(
        \MC_ARK_ARC_1_1/temp3[109] ) );
  XOR2_X1 U7494 ( .A1(\MC_ARK_ARC_1_0/temp5[46] ), .A2(n2622), .Z(
        \MC_ARK_ARC_1_0/buf_output[46] ) );
  XOR2_X1 U7495 ( .A1(\MC_ARK_ARC_1_0/temp3[46] ), .A2(
        \MC_ARK_ARC_1_0/temp4[46] ), .Z(n2622) );
  NAND3_X1 U7498 ( .A1(\SB1_0_11/i0_3 ), .A2(\SB1_0_11/i0_0 ), .A3(
        \SB1_0_11/i0[7] ), .ZN(\SB1_0_11/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U7501 ( .A1(\SB2_2_18/i0_0 ), .A2(\SB2_2_18/i3[0] ), .A3(
        \SB2_2_18/i1_7 ), .ZN(\SB2_2_18/Component_Function_4/NAND4_in[1] ) );
  NAND4_X2 U7502 ( .A1(\SB1_0_16/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_0_16/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_16/Component_Function_1/NAND4_in[0] ), .A4(n2626), .ZN(
        \SB1_0_16/buf_output[1] ) );
  NAND3_X1 U7503 ( .A1(n4752), .A2(\SB1_0_16/i1_7 ), .A3(\SB1_0_16/i0[8] ), 
        .ZN(n2626) );
  NAND3_X1 U7504 ( .A1(\SB2_0_8/i0_3 ), .A2(\SB2_0_8/i0[10] ), .A3(
        \RI3[0][142] ), .ZN(\SB2_0_8/Component_Function_0/NAND4_in[2] ) );
  BUF_X4 U7506 ( .I(\SB2_2_18/buf_output[2] ), .Z(\RI5[2][98] ) );
  NAND3_X1 U7513 ( .A1(\SB4_23/i0_4 ), .A2(\SB4_23/i1_7 ), .A3(\SB4_23/i0[8] ), 
        .ZN(n2632) );
  NAND3_X1 U7516 ( .A1(\SB2_0_5/i0[10] ), .A2(\SB2_0_5/i0_0 ), .A3(
        \SB2_0_5/i0[6] ), .ZN(\SB2_0_5/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 U7517 ( .I(\SB2_3_15/buf_output[4] ), .Z(\RI5[3][106] ) );
  NAND4_X2 U7518 ( .A1(\SB1_1_18/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_1_18/Component_Function_4/NAND4_in[2] ), .A3(
        \SB1_1_18/Component_Function_4/NAND4_in[0] ), .A4(n2637), .ZN(
        \SB1_1_18/buf_output[4] ) );
  XOR2_X1 U7523 ( .A1(n2640), .A2(n2639), .Z(\MC_ARK_ARC_1_0/buf_output[184] )
         );
  XOR2_X1 U7524 ( .A1(\MC_ARK_ARC_1_0/temp1[184] ), .A2(
        \MC_ARK_ARC_1_0/temp4[184] ), .Z(n2639) );
  XOR2_X1 U7527 ( .A1(\MC_ARK_ARC_1_3/temp2[178] ), .A2(
        \MC_ARK_ARC_1_3/temp1[178] ), .Z(\MC_ARK_ARC_1_3/temp5[178] ) );
  NAND3_X1 U7528 ( .A1(\SB1_1_7/i0_0 ), .A2(\SB1_1_7/i1_7 ), .A3(
        \SB1_1_7/i3[0] ), .ZN(\SB1_1_7/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U7536 ( .A1(\SB4_24/i0_3 ), .A2(\SB4_24/i1[9] ), .A3(\SB4_24/i0[6] ), .ZN(\SB4_24/Component_Function_3/NAND4_in[0] ) );
  NAND4_X2 U7538 ( .A1(\SB1_2_2/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_2/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_2/Component_Function_0/NAND4_in[0] ), .A4(n2647), .ZN(
        \SB1_2_2/buf_output[0] ) );
  NAND4_X2 U7540 ( .A1(\SB1_0_24/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_0_24/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_0_24/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_0_24/Component_Function_0/NAND4_in[0] ), .ZN(\RI3[0][72] ) );
  NAND3_X1 U7542 ( .A1(\SB1_2_25/i0_0 ), .A2(\SB1_2_25/i3[0] ), .A3(
        \SB1_2_25/i1_7 ), .ZN(\SB1_2_25/Component_Function_4/NAND4_in[1] ) );
  INV_X2 U7543 ( .I(n2651), .ZN(\SB1_3_23/i0_4 ) );
  XOR2_X1 U7544 ( .A1(\MC_ARK_ARC_1_3/temp5[19] ), .A2(n2652), .Z(
        \MC_ARK_ARC_1_3/buf_output[19] ) );
  XOR2_X1 U7545 ( .A1(\MC_ARK_ARC_1_3/temp3[19] ), .A2(
        \MC_ARK_ARC_1_3/temp4[19] ), .Z(n2652) );
  BUF_X4 U7546 ( .I(\SB2_1_14/buf_output[1] ), .Z(\RI5[1][127] ) );
  XOR2_X1 U7551 ( .A1(n1365), .A2(n535), .Z(n2660) );
  NAND3_X1 U7555 ( .A1(\SB4_28/i0_0 ), .A2(\SB4_28/i1_5 ), .A3(\SB4_28/i0_4 ), 
        .ZN(n2663) );
  XOR2_X1 U7556 ( .A1(\RI5[1][113] ), .A2(\RI5[1][137] ), .Z(n2664) );
  NAND4_X2 U7557 ( .A1(\SB2_2_24/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_2_24/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_2_24/Component_Function_4/NAND4_in[1] ), .A4(n2665), .ZN(
        \SB2_2_24/buf_output[4] ) );
  XOR2_X1 U7559 ( .A1(n2666), .A2(\MC_ARK_ARC_1_3/temp5[33] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[33] ) );
  NAND3_X1 U7567 ( .A1(\SB2_0_28/i1[9] ), .A2(\SB2_0_28/i1_5 ), .A3(
        \SB2_0_28/i0[10] ), .ZN(\SB2_0_28/Component_Function_2/NAND4_in[0] )
         );
  NAND3_X1 U7568 ( .A1(\SB4_28/i0_0 ), .A2(\SB4_28/i0[9] ), .A3(\SB4_28/i0[8] ), .ZN(n2671) );
  XOR2_X1 U7571 ( .A1(n2673), .A2(\RI5[0][11] ), .Z(n2709) );
  XOR2_X1 U7573 ( .A1(\MC_ARK_ARC_1_3/temp6[12] ), .A2(n2675), .Z(
        \MC_ARK_ARC_1_3/buf_output[12] ) );
  XOR2_X1 U7574 ( .A1(\MC_ARK_ARC_1_3/temp2[12] ), .A2(
        \MC_ARK_ARC_1_3/temp1[12] ), .Z(n2675) );
  NAND4_X2 U7579 ( .A1(\SB1_0_14/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_0_14/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_14/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_14/Component_Function_1/NAND4_in[0] ), .ZN(\RI3[0][127] ) );
  NAND4_X2 U7580 ( .A1(\SB1_1_13/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_13/Component_Function_3/NAND4_in[2] ), .A3(
        \SB1_1_13/Component_Function_3/NAND4_in[1] ), .A4(n2678), .ZN(
        \SB1_1_13/buf_output[3] ) );
  XOR2_X1 U7581 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[99] ), .A2(\RI5[2][63] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[189] ) );
  BUF_X2 U7582 ( .I(\SB2_0_27/i0[9] ), .Z(n2679) );
  XOR2_X1 U7585 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[179] ), .A2(\RI5[3][143] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[77] ) );
  XOR2_X1 U7598 ( .A1(\MC_ARK_ARC_1_2/temp1[153] ), .A2(
        \MC_ARK_ARC_1_2/temp2[153] ), .Z(n2690) );
  XOR2_X1 U7600 ( .A1(\RI5[1][96] ), .A2(\RI5[1][132] ), .Z(n2691) );
  XOR2_X1 U7601 ( .A1(\RI5[1][135] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[99] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[33] ) );
  NAND3_X1 U7603 ( .A1(\SB4_9/i0_4 ), .A2(\SB4_9/i1_7 ), .A3(\SB4_9/i0[8] ), 
        .ZN(n2693) );
  NAND4_X2 U7604 ( .A1(\SB1_2_22/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_2_22/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_2_22/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_2_22/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_2_22/buf_output[0] ) );
  NAND3_X1 U7606 ( .A1(\SB4_27/i0_3 ), .A2(n1389), .A3(\SB4_27/i0_4 ), .ZN(
        n2695) );
  XOR2_X1 U7614 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[35] ), .A2(\RI5[1][191] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[125] ) );
  XOR2_X1 U7617 ( .A1(\MC_ARK_ARC_1_3/temp4[6] ), .A2(
        \MC_ARK_ARC_1_3/temp3[6] ), .Z(n2881) );
  NAND4_X2 U7624 ( .A1(\SB2_1_13/Component_Function_4/NAND4_in[1] ), .A2(n2703), .A3(\SB2_1_13/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_1_13/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_1_13/buf_output[4] ) );
  INV_X1 U7629 ( .I(\SB3_26/buf_output[5] ), .ZN(\SB4_26/i1_5 ) );
  XOR2_X1 U7631 ( .A1(n2708), .A2(\MC_ARK_ARC_1_0/temp6[11] ), .Z(n2785) );
  XOR2_X1 U7632 ( .A1(n2709), .A2(\MC_ARK_ARC_1_0/temp2[11] ), .Z(n2708) );
  BUF_X4 U7637 ( .I(\SB2_2_26/buf_output[0] ), .Z(\RI5[2][60] ) );
  NAND3_X1 U7639 ( .A1(n388), .A2(\SB1_0_8/i0[9] ), .A3(\SB1_0_8/i0[6] ), .ZN(
        n2715) );
  NAND4_X2 U7640 ( .A1(\SB1_0_22/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_0_22/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_0_22/Component_Function_1/NAND4_in[1] ), .A4(
        \SB1_0_22/Component_Function_1/NAND4_in[0] ), .ZN(\RI3[0][79] ) );
  NAND4_X2 U7641 ( .A1(\SB1_0_15/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_0_15/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_0_15/Component_Function_1/NAND4_in[1] ), .A4(
        \SB1_0_15/Component_Function_1/NAND4_in[0] ), .ZN(\RI3[0][121] ) );
  XOR2_X1 U7642 ( .A1(\RI5[0][87] ), .A2(\RI5[0][63] ), .Z(
        \MC_ARK_ARC_1_0/temp2[117] ) );
  XOR2_X1 U7643 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[177] ), .A2(\RI5[2][21] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[111] ) );
  INV_X4 U7644 ( .I(n2806), .ZN(\SB1_1_22/buf_output[1] ) );
  NAND4_X2 U7648 ( .A1(\SB1_0_24/Component_Function_3/NAND4_in[2] ), .A2(
        \SB1_0_24/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_24/Component_Function_3/NAND4_in[0] ), .A4(
        \SB1_0_24/Component_Function_3/NAND4_in[3] ), .ZN(\RI3[0][57] ) );
  XOR2_X1 U7653 ( .A1(\MC_ARK_ARC_1_2/temp1[126] ), .A2(
        \MC_ARK_ARC_1_2/temp2[126] ), .Z(\MC_ARK_ARC_1_2/temp5[126] ) );
  BUF_X4 U7654 ( .I(\SB2_2_20/buf_output[0] ), .Z(\RI5[2][96] ) );
  BUF_X4 U7657 ( .I(\SB2_1_21/buf_output[3] ), .Z(\RI5[1][75] ) );
  XOR2_X1 U7664 ( .A1(\MC_ARK_ARC_1_2/temp2[80] ), .A2(
        \MC_ARK_ARC_1_2/temp1[80] ), .Z(\MC_ARK_ARC_1_2/temp5[80] ) );
  NAND4_X2 U7665 ( .A1(\SB1_0_31/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_0_31/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_0_31/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_0_31/Component_Function_0/NAND4_in[0] ), .ZN(\RI3[0][30] ) );
  XOR2_X1 U7669 ( .A1(\MC_ARK_ARC_1_1/temp1[120] ), .A2(
        \MC_ARK_ARC_1_1/temp2[120] ), .Z(\MC_ARK_ARC_1_1/temp5[120] ) );
  XOR2_X1 U7675 ( .A1(n2735), .A2(\MC_ARK_ARC_1_0/temp5[79] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[79] ) );
  XOR2_X1 U7676 ( .A1(\MC_ARK_ARC_1_0/temp3[79] ), .A2(
        \MC_ARK_ARC_1_0/temp4[79] ), .Z(n2735) );
  NAND4_X2 U7680 ( .A1(\SB1_0_2/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_0_2/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_0_2/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_0_2/Component_Function_0/NAND4_in[0] ), .ZN(\SB2_0_29/i0[9] ) );
  NAND4_X2 U7681 ( .A1(\SB1_0_14/Component_Function_5/NAND4_in[3] ), .A2(
        \SB1_0_14/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_14/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_0_14/Component_Function_5/NAND4_in[0] ), .ZN(\RI3[0][107] ) );
  NAND4_X2 U7684 ( .A1(\SB1_0_6/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_0_6/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_0_6/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_6/Component_Function_0/NAND4_in[0] ), .ZN(\RI3[0][180] ) );
  BUF_X4 U7685 ( .I(\SB2_2_19/buf_output[5] ), .Z(\RI5[2][77] ) );
  XOR2_X1 U7690 ( .A1(\MC_ARK_ARC_1_0/temp1[165] ), .A2(
        \MC_ARK_ARC_1_0/temp2[165] ), .Z(\MC_ARK_ARC_1_0/temp5[165] ) );
  NAND3_X1 U7693 ( .A1(\SB1_1_26/i0_3 ), .A2(\SB1_1_26/i0[7] ), .A3(
        \SB1_1_26/i0_0 ), .ZN(n2742) );
  BUF_X4 U7697 ( .I(\SB2_2_23/buf_output[1] ), .Z(\RI5[2][73] ) );
  NAND3_X1 U7699 ( .A1(\SB2_1_25/i0_3 ), .A2(\SB2_1_25/i0[10] ), .A3(n1579), 
        .ZN(\SB2_1_25/Component_Function_0/NAND4_in[2] ) );
  BUF_X2 U7700 ( .I(\SB1_1_13/buf_output[0] ), .Z(n2745) );
  NAND3_X1 U7701 ( .A1(\SB4_27/i0_4 ), .A2(n1389), .A3(\SB4_27/i1_5 ), .ZN(
        n2746) );
  XOR2_X1 U7710 ( .A1(\MC_ARK_ARC_1_2/temp3[90] ), .A2(
        \MC_ARK_ARC_1_2/temp4[90] ), .Z(n2751) );
  NAND3_X1 U7718 ( .A1(\SB3_7/buf_output[2] ), .A2(\SB4_4/i3[0] ), .A3(
        \SB4_4/i1_7 ), .ZN(\SB4_4/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U7722 ( .A1(\SB4_13/i0_3 ), .A2(\SB4_13/i0[10] ), .A3(
        \SB4_13/i0[9] ), .ZN(n2759) );
  XOR2_X1 U7725 ( .A1(\RI5[1][103] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[139] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[37] ) );
  NAND3_X1 U7728 ( .A1(\SB4_5/i0_4 ), .A2(\SB4_5/i1[9] ), .A3(\SB4_5/i1_5 ), 
        .ZN(n2766) );
  XOR2_X1 U7731 ( .A1(\MC_ARK_ARC_1_3/temp3[14] ), .A2(
        \MC_ARK_ARC_1_3/temp4[14] ), .Z(n2768) );
  NAND4_X2 U7741 ( .A1(\SB1_0_27/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_0_27/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_0_27/Component_Function_1/NAND4_in[1] ), .A4(
        \SB1_0_27/Component_Function_1/NAND4_in[0] ), .ZN(\RI3[0][49] ) );
  XOR2_X1 U7742 ( .A1(\MC_ARK_ARC_1_0/temp2[38] ), .A2(
        \MC_ARK_ARC_1_0/temp1[38] ), .Z(\MC_ARK_ARC_1_0/temp5[38] ) );
  NAND3_X1 U7743 ( .A1(\SB3_22/i1_5 ), .A2(\SB3_22/i0_4 ), .A3(\SB3_22/i1[9] ), 
        .ZN(\SB3_22/Component_Function_4/NAND4_in[3] ) );
  XOR2_X1 U7746 ( .A1(n2775), .A2(n95), .Z(Ciphertext[61]) );
  XOR2_X1 U7748 ( .A1(\MC_ARK_ARC_1_0/temp2[96] ), .A2(
        \MC_ARK_ARC_1_0/temp1[96] ), .Z(n2776) );
  NAND3_X1 U7749 ( .A1(\SB4_3/i0_3 ), .A2(n1371), .A3(\SB4_3/i0[6] ), .ZN(
        n2777) );
  BUF_X4 U7750 ( .I(\SB2_1_18/buf_output[4] ), .Z(\RI5[1][88] ) );
  BUF_X4 U7751 ( .I(\SB2_1_30/buf_output[4] ), .Z(\RI5[1][16] ) );
  BUF_X4 U7753 ( .I(\SB2_2_29/buf_output[4] ), .Z(\RI5[2][22] ) );
  XOR2_X1 U7758 ( .A1(n2781), .A2(\MC_ARK_ARC_1_2/temp6[94] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[94] ) );
  XOR2_X1 U7759 ( .A1(\MC_ARK_ARC_1_2/temp2[94] ), .A2(
        \MC_ARK_ARC_1_2/temp1[94] ), .Z(n2781) );
  BUF_X4 U7760 ( .I(\SB2_2_22/buf_output[4] ), .Z(\RI5[2][64] ) );
  XOR2_X1 U7761 ( .A1(n2783), .A2(\MC_ARK_ARC_1_1/temp1[44] ), .Z(
        \MC_ARK_ARC_1_1/temp5[44] ) );
  XOR2_X1 U7762 ( .A1(\RI5[1][14] ), .A2(\RI5[1][182] ), .Z(n2783) );
  BUF_X4 U7763 ( .I(\SB2_2_21/buf_output[2] ), .Z(\RI5[2][80] ) );
  INV_X2 U7765 ( .I(n2785), .ZN(\RI1[1][11] ) );
  INV_X2 U7769 ( .I(\SB1_0_1/buf_output[5] ), .ZN(\SB2_0_1/i1_5 ) );
  NAND3_X2 U7771 ( .A1(\SB1_1_25/i0_4 ), .A2(\SB1_1_25/i1[9] ), .A3(
        \SB1_1_25/i0_3 ), .ZN(n2789) );
  XOR2_X1 U7773 ( .A1(\MC_ARK_ARC_1_0/temp6[40] ), .A2(n2790), .Z(
        \MC_ARK_ARC_1_0/buf_output[40] ) );
  XOR2_X1 U7774 ( .A1(\MC_ARK_ARC_1_0/temp2[40] ), .A2(
        \MC_ARK_ARC_1_0/temp1[40] ), .Z(n2790) );
  NAND3_X1 U7775 ( .A1(\SB2_1_29/i1_7 ), .A2(\SB2_1_29/i0_4 ), .A3(
        \SB2_1_29/i0[8] ), .ZN(\SB2_1_29/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U7777 ( .A1(\SB1_1_16/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_1_16/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_16/Component_Function_1/NAND4_in[0] ), .A4(n2792), .ZN(
        \SB1_1_16/buf_output[1] ) );
  NAND3_X2 U7779 ( .A1(\SB1_1_15/i0[10] ), .A2(\SB1_1_15/i0_0 ), .A3(
        \SB1_1_15/i0[6] ), .ZN(\SB1_1_15/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U7784 ( .A1(\SB1_1_13/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_1_13/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_1_13/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_1_13/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_1_13/buf_output[0] ) );
  XOR2_X1 U7785 ( .A1(\MC_ARK_ARC_1_1/temp6[189] ), .A2(n2799), .Z(
        \MC_ARK_ARC_1_1/buf_output[189] ) );
  BUF_X4 U7787 ( .I(\SB2_3_24/buf_output[4] ), .Z(\RI5[3][52] ) );
  XOR2_X1 U7788 ( .A1(\MC_ARK_ARC_1_2/temp6[182] ), .A2(n2801), .Z(
        \MC_ARK_ARC_1_2/buf_output[182] ) );
  INV_X2 U7790 ( .I(n2803), .ZN(\RI1[2][167] ) );
  BUF_X4 U7791 ( .I(\SB2_2_2/buf_output[0] ), .Z(\RI5[2][12] ) );
  XOR2_X1 U7794 ( .A1(\MC_ARK_ARC_1_0/temp3[84] ), .A2(
        \MC_ARK_ARC_1_0/temp4[84] ), .Z(n2805) );
  NAND3_X1 U7795 ( .A1(\SB4_23/i0[10] ), .A2(\SB4_23/i0_3 ), .A3(\SB4_23/i0_4 ), .ZN(\SB4_23/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U7796 ( .A1(\SB4_25/i0_0 ), .A2(\SB4_25/i1_5 ), .A3(\SB4_25/i0_4 ), 
        .ZN(\SB4_25/Component_Function_2/NAND4_in[3] ) );
  NAND4_X2 U7801 ( .A1(\SB1_0_23/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_0_23/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_0_23/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_23/Component_Function_4/NAND4_in[3] ), .ZN(\RI3[0][58] ) );
  NAND3_X1 U7802 ( .A1(\SB1_0_14/i0_3 ), .A2(\SB1_0_14/i0_0 ), .A3(
        \SB1_0_14/i0[7] ), .ZN(\SB1_0_14/Component_Function_0/NAND4_in[3] ) );
  BUF_X4 U7803 ( .I(\SB2_3_22/buf_output[3] ), .Z(\RI5[3][69] ) );
  XOR2_X1 U7804 ( .A1(\MC_ARK_ARC_1_1/temp5[52] ), .A2(n2812), .Z(
        \MC_ARK_ARC_1_1/buf_output[52] ) );
  XOR2_X1 U7806 ( .A1(n2813), .A2(\MC_ARK_ARC_1_2/temp5[37] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[37] ) );
  BUF_X4 U7807 ( .I(\SB2_1_6/buf_output[0] ), .Z(\RI5[1][180] ) );
  NAND3_X1 U7808 ( .A1(\SB2_2_25/i0_3 ), .A2(\SB2_2_25/i0[10] ), .A3(
        \SB2_2_25/i0_4 ), .ZN(\SB2_2_25/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U7812 ( .A1(\MC_ARK_ARC_1_0/temp3[102] ), .A2(
        \MC_ARK_ARC_1_0/temp4[102] ), .Z(n2853) );
  NAND3_X1 U7814 ( .A1(\SB4_8/i0[10] ), .A2(\SB4_8/i1[9] ), .A3(\SB4_8/i1_7 ), 
        .ZN(\SB4_8/Component_Function_3/NAND4_in[2] ) );
  XOR2_X1 U7815 ( .A1(\MC_ARK_ARC_1_2/temp5[14] ), .A2(
        \MC_ARK_ARC_1_2/temp6[14] ), .Z(\MC_ARK_ARC_1_2/buf_output[14] ) );
  BUF_X4 U7817 ( .I(\SB2_2_6/buf_output[0] ), .Z(\RI5[2][180] ) );
  XOR2_X1 U7819 ( .A1(n2816), .A2(\MC_ARK_ARC_1_0/temp5[120] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[120] ) );
  XOR2_X1 U7820 ( .A1(\MC_ARK_ARC_1_0/temp3[120] ), .A2(
        \MC_ARK_ARC_1_0/temp4[120] ), .Z(n2816) );
  NAND4_X2 U7822 ( .A1(\SB1_2_22/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_2_22/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_2_22/Component_Function_1/NAND4_in[3] ), .A4(
        \SB1_2_22/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_2_22/buf_output[1] ) );
  XOR2_X1 U7823 ( .A1(\RI5[3][107] ), .A2(\RI5[3][143] ), .Z(
        \MC_ARK_ARC_1_3/temp3[41] ) );
  XOR2_X1 U7824 ( .A1(\MC_ARK_ARC_1_2/temp6[171] ), .A2(n2819), .Z(
        \MC_ARK_ARC_1_2/buf_output[171] ) );
  XOR2_X1 U7826 ( .A1(n2820), .A2(\MC_ARK_ARC_1_3/temp6[63] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[63] ) );
  XOR2_X1 U7829 ( .A1(\MC_ARK_ARC_1_1/temp3[169] ), .A2(
        \MC_ARK_ARC_1_1/temp4[169] ), .Z(n2823) );
  NAND3_X1 U7831 ( .A1(\SB1_1_10/i0_0 ), .A2(\SB1_1_10/i1_7 ), .A3(
        \SB1_1_10/i3[0] ), .ZN(\SB1_1_10/Component_Function_4/NAND4_in[1] ) );
  BUF_X4 U7832 ( .I(\SB2_1_9/buf_output[4] ), .Z(\RI5[1][142] ) );
  INV_X2 U7834 ( .I(\SB1_3_18/buf_output[5] ), .ZN(\SB2_3_18/i1_5 ) );
  BUF_X4 U7837 ( .I(\SB2_1_23/buf_output[4] ), .Z(\RI5[1][58] ) );
  NAND3_X2 U7838 ( .A1(\SB1_2_0/i0[10] ), .A2(\SB1_2_0/i0[9] ), .A3(
        \SB1_2_0/i0_3 ), .ZN(\SB1_2_0/Component_Function_4/NAND4_in[2] ) );
  XOR2_X1 U7839 ( .A1(n2827), .A2(\MC_ARK_ARC_1_0/temp6[3] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[3] ) );
  NAND3_X1 U7840 ( .A1(\SB1_1_20/i0_3 ), .A2(\SB1_1_20/i0[10] ), .A3(
        \SB1_1_20/i0_4 ), .ZN(\SB1_1_20/Component_Function_0/NAND4_in[2] ) );
  BUF_X4 U7843 ( .I(\SB2_3_20/buf_output[4] ), .Z(\RI5[3][76] ) );
  NAND4_X2 U7848 ( .A1(\SB1_0_9/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_0_9/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_0_9/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_9/Component_Function_0/NAND4_in[0] ), .ZN(\RI3[0][162] ) );
  XOR2_X1 U7850 ( .A1(\MC_ARK_ARC_1_2/temp5[30] ), .A2(n2833), .Z(
        \MC_ARK_ARC_1_2/buf_output[30] ) );
  XOR2_X1 U7851 ( .A1(\MC_ARK_ARC_1_2/temp3[30] ), .A2(
        \MC_ARK_ARC_1_2/temp4[30] ), .Z(n2833) );
  XOR2_X1 U7854 ( .A1(\MC_ARK_ARC_1_0/temp5[162] ), .A2(
        \MC_ARK_ARC_1_0/temp6[162] ), .Z(\MC_ARK_ARC_1_0/buf_output[162] ) );
  NAND3_X2 U7857 ( .A1(\SB2_1_14/i0_4 ), .A2(\SB2_1_14/i0[9] ), .A3(
        \SB2_1_14/i0[6] ), .ZN(n2834) );
  XOR2_X1 U7858 ( .A1(\MC_ARK_ARC_1_3/temp6[21] ), .A2(
        \MC_ARK_ARC_1_3/temp5[21] ), .Z(\MC_ARK_ARC_1_3/buf_output[21] ) );
  NAND3_X1 U7859 ( .A1(\SB1_0_9/i0_3 ), .A2(\SB1_0_9/i0[10] ), .A3(
        \SB1_0_9/i0[9] ), .ZN(\SB1_0_9/Component_Function_4/NAND4_in[2] ) );
  NAND4_X2 U7860 ( .A1(\SB1_1_15/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_1_15/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_15/Component_Function_0/NAND4_in[0] ), .A4(n2835), .ZN(
        \SB1_1_15/buf_output[0] ) );
  XOR2_X1 U7864 ( .A1(n2837), .A2(\MC_ARK_ARC_1_0/temp5[21] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[21] ) );
  NAND3_X1 U7871 ( .A1(\SB4_25/i0[10] ), .A2(\SB4_25/i0_3 ), .A3(
        \SB4_25/i0[9] ), .ZN(n2839) );
  BUF_X4 U7874 ( .I(\SB2_3_23/buf_output[0] ), .Z(\RI5[3][78] ) );
  NAND4_X2 U7880 ( .A1(\SB1_2_24/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_24/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_24/Component_Function_0/NAND4_in[0] ), .A4(n2844), .ZN(
        \SB1_2_24/buf_output[0] ) );
  XOR2_X1 U7882 ( .A1(n2845), .A2(\MC_ARK_ARC_1_3/temp5[140] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[140] ) );
  XOR2_X1 U7883 ( .A1(\MC_ARK_ARC_1_3/temp5[51] ), .A2(n2847), .Z(
        \MC_ARK_ARC_1_3/buf_output[51] ) );
  XOR2_X1 U7884 ( .A1(\MC_ARK_ARC_1_3/temp3[51] ), .A2(
        \MC_ARK_ARC_1_3/temp4[51] ), .Z(n2847) );
  XOR2_X1 U7887 ( .A1(\MC_ARK_ARC_1_0/temp6[56] ), .A2(
        \MC_ARK_ARC_1_0/temp5[56] ), .Z(\MC_ARK_ARC_1_0/buf_output[56] ) );
  XOR2_X1 U7888 ( .A1(\MC_ARK_ARC_1_0/temp2[32] ), .A2(
        \MC_ARK_ARC_1_0/temp1[32] ), .Z(\MC_ARK_ARC_1_0/temp5[32] ) );
  NAND4_X2 U7892 ( .A1(\SB1_3_29/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_3_29/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_3_29/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_3_29/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_3_29/buf_output[0] ) );
  XOR2_X1 U7896 ( .A1(\MC_ARK_ARC_1_1/temp5[177] ), .A2(n2854), .Z(
        \MC_ARK_ARC_1_1/buf_output[177] ) );
  XOR2_X1 U7899 ( .A1(\MC_ARK_ARC_1_2/temp5[168] ), .A2(
        \MC_ARK_ARC_1_2/temp6[168] ), .Z(\MC_ARK_ARC_1_2/buf_output[168] ) );
  NAND3_X1 U7901 ( .A1(\SB3_2/i1_5 ), .A2(\SB3_2/i1[9] ), .A3(\SB3_2/i0_4 ), 
        .ZN(\SB3_2/Component_Function_4/NAND4_in[3] ) );
  NOR2_X2 U7906 ( .A1(n2883), .A2(n2884), .ZN(n2882) );
  NAND3_X1 U7908 ( .A1(\SB1_0_17/i0_0 ), .A2(\SB1_0_17/i3[0] ), .A3(
        \SB1_0_17/i1_7 ), .ZN(\SB1_0_17/Component_Function_4/NAND4_in[1] ) );
  BUF_X4 U7913 ( .I(\SB2_3_23/buf_output[4] ), .Z(\RI5[3][58] ) );
  BUF_X4 U7917 ( .I(\SB2_3_24/buf_output[5] ), .Z(\RI5[3][47] ) );
  INV_X2 U7918 ( .I(n2864), .ZN(\MC_ARK_ARC_1_3/buf_output[101] ) );
  XNOR2_X1 U7919 ( .A1(\MC_ARK_ARC_1_3/temp6[101] ), .A2(
        \MC_ARK_ARC_1_3/temp5[101] ), .ZN(n2864) );
  NAND3_X1 U7920 ( .A1(\SB1_1_25/i0_0 ), .A2(\SB1_1_25/i0_4 ), .A3(
        \SB1_1_25/i1_5 ), .ZN(n2865) );
  XOR2_X1 U7925 ( .A1(\MC_ARK_ARC_1_3/temp3[11] ), .A2(
        \MC_ARK_ARC_1_3/temp4[11] ), .Z(\MC_ARK_ARC_1_3/temp6[11] ) );
  BUF_X4 U7926 ( .I(\SB2_1_13/buf_output[2] ), .Z(\RI5[1][128] ) );
  BUF_X4 U7927 ( .I(\SB2_2_27/buf_output[0] ), .Z(\RI5[2][54] ) );
  XOR2_X1 U7928 ( .A1(\MC_ARK_ARC_1_2/temp5[108] ), .A2(
        \MC_ARK_ARC_1_2/temp6[108] ), .Z(\MC_ARK_ARC_1_2/buf_output[108] ) );
  NAND3_X1 U7930 ( .A1(\SB1_0_17/i0[10] ), .A2(\SB1_0_17/i1[9] ), .A3(
        \SB1_0_17/i1_7 ), .ZN(\SB1_0_17/Component_Function_3/NAND4_in[2] ) );
  XOR2_X1 U7932 ( .A1(\MC_ARK_ARC_1_3/temp5[131] ), .A2(
        \MC_ARK_ARC_1_3/temp6[131] ), .Z(\RI1[4][131] ) );
  NAND3_X2 U7936 ( .A1(\SB1_3_31/i0_3 ), .A2(\SB1_3_31/i1[9] ), .A3(
        \SB1_3_31/i0_4 ), .ZN(\SB1_3_31/Component_Function_5/NAND4_in[2] ) );
  BUF_X4 U7938 ( .I(\SB2_3_31/buf_output[0] ), .Z(\RI5[3][30] ) );
  XOR2_X1 U7942 ( .A1(\MC_ARK_ARC_1_1/temp6[27] ), .A2(
        \MC_ARK_ARC_1_1/temp5[27] ), .Z(\MC_ARK_ARC_1_1/buf_output[27] ) );
  XOR2_X1 U7945 ( .A1(\MC_ARK_ARC_1_0/temp5[76] ), .A2(n2875), .Z(
        \MC_ARK_ARC_1_0/buf_output[76] ) );
  XOR2_X1 U7946 ( .A1(\MC_ARK_ARC_1_0/temp3[76] ), .A2(
        \MC_ARK_ARC_1_0/temp4[76] ), .Z(n2875) );
  NAND3_X1 U7949 ( .A1(\SB4_17/i0[10] ), .A2(\SB4_17/i0_0 ), .A3(
        \SB4_17/i0[6] ), .ZN(\SB4_17/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U7954 ( .A1(\SB4_29/i0[9] ), .A2(n1793), .A3(\SB4_29/i0[6] ), .ZN(
        n2880) );
  BUF_X4 U7955 ( .I(\SB2_3_29/buf_output[0] ), .Z(\RI5[3][42] ) );
  XOR2_X1 U7956 ( .A1(\MC_ARK_ARC_1_3/temp5[6] ), .A2(n2881), .Z(
        \MC_ARK_ARC_1_3/buf_output[6] ) );
  BUF_X4 U7959 ( .I(\SB2_2_25/buf_output[5] ), .Z(\RI5[2][41] ) );
  XOR2_X1 U7960 ( .A1(\MC_ARK_ARC_1_0/temp5[173] ), .A2(
        \MC_ARK_ARC_1_0/temp6[173] ), .Z(\RI1[1][173] ) );
  BUF_X4 U7961 ( .I(\SB2_1_3/buf_output[4] ), .Z(\RI5[1][178] ) );
  BUF_X4 U7962 ( .I(\SB2_1_23/buf_output[1] ), .Z(\RI5[1][73] ) );
  BUF_X4 U7963 ( .I(\SB2_2_7/buf_output[0] ), .Z(\RI5[2][174] ) );
  XOR2_X1 U7965 ( .A1(\MC_ARK_ARC_1_3/temp3[3] ), .A2(
        \MC_ARK_ARC_1_3/temp4[3] ), .Z(\MC_ARK_ARC_1_3/temp6[3] ) );
  XOR2_X1 U7971 ( .A1(\MC_ARK_ARC_1_3/temp4[129] ), .A2(
        \MC_ARK_ARC_1_3/temp3[129] ), .Z(n2886) );
  BUF_X4 U7976 ( .I(\SB2_1_23/buf_output[0] ), .Z(\RI5[1][78] ) );
  BUF_X4 U7977 ( .I(\SB2_2_28/buf_output[5] ), .Z(\RI5[2][23] ) );
  XOR2_X1 U7980 ( .A1(\RI5[1][71] ), .A2(\RI5[1][107] ), .Z(
        \MC_ARK_ARC_1_1/temp3[5] ) );
  NAND3_X2 U7982 ( .A1(\SB1_1_3/i0_3 ), .A2(\SB1_1_3/i1[9] ), .A3(
        \SB1_1_3/i0_4 ), .ZN(\SB1_1_3/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U7983 ( .A1(\MC_ARK_ARC_1_3/temp6[143] ), .A2(
        \MC_ARK_ARC_1_3/temp5[143] ), .Z(\RI1[4][143] ) );
  BUF_X4 U7985 ( .I(\SB2_1_13/buf_output[0] ), .Z(\RI5[1][138] ) );
  BUF_X4 U7987 ( .I(\SB2_1_26/buf_output[4] ), .Z(\RI5[1][40] ) );
  BUF_X4 U7988 ( .I(\SB2_2_25/buf_output[4] ), .Z(\RI5[2][46] ) );
  BUF_X4 U7989 ( .I(\SB2_1_7/buf_output[5] ), .Z(\RI5[1][149] ) );
  BUF_X4 U7990 ( .I(\SB2_3_12/buf_output[4] ), .Z(\RI5[3][124] ) );
  BUF_X4 U7991 ( .I(\SB2_1_22/buf_output[4] ), .Z(\RI5[1][64] ) );
  BUF_X4 U7992 ( .I(\SB2_3_26/buf_output[2] ), .Z(\RI5[3][50] ) );
  BUF_X4 U7993 ( .I(\SB2_2_23/buf_output[3] ), .Z(\RI5[2][63] ) );
  BUF_X4 U7996 ( .I(\SB2_1_13/buf_output[4] ), .Z(\RI5[1][118] ) );
  BUF_X4 U7997 ( .I(\SB2_3_17/buf_output[5] ), .Z(\RI5[3][89] ) );
  BUF_X4 U7998 ( .I(\SB2_1_5/buf_output[5] ), .Z(\RI5[1][161] ) );
  BUF_X4 U8000 ( .I(\SB2_0_27/buf_output[5] ), .Z(\RI5[0][29] ) );
  NAND4_X2 U8001 ( .A1(\SB2_0_27/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_27/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_0_27/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_0_27/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_0_27/buf_output[2] ) );
  NAND4_X2 U8002 ( .A1(\SB1_0_30/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_30/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_30/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_30/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB1_0_30/buf_output[2] ) );
  NAND4_X2 U8004 ( .A1(\SB2_0_29/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_29/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_29/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_29/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB2_0_29/buf_output[0] ) );
  NAND4_X2 U8005 ( .A1(\SB1_0_30/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_30/Component_Function_4/NAND4_in[3] ), .A3(
        \SB1_0_30/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_0_30/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB1_0_30/buf_output[4] ) );
  NAND4_X2 U8006 ( .A1(\SB1_0_30/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_30/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_30/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_30/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_0_30/buf_output[0] ) );
  BUF_X4 U8008 ( .I(\SB2_0_26/buf_output[2] ), .Z(\RI5[0][50] ) );
  BUF_X4 U8009 ( .I(\SB2_0_26/buf_output[3] ), .Z(\RI5[0][45] ) );
  BUF_X4 U8010 ( .I(\SB2_0_26/buf_output[5] ), .Z(\RI5[0][35] ) );
  NAND4_X2 U8016 ( .A1(\SB1_1_18/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_18/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_18/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_18/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_1_18/buf_output[1] ) );
  BUF_X4 U8017 ( .I(\SB2_0_30/buf_output[2] ), .Z(\RI5[0][26] ) );
  NAND4_X2 U8023 ( .A1(\SB1_1_7/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_7/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_7/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_7/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_1_7/buf_output[0] ) );
  NAND4_X2 U8025 ( .A1(\SB1_1_13/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_13/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_13/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_13/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_1_13/buf_output[1] ) );
  NAND4_X2 U8030 ( .A1(\SB1_1_27/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_27/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_27/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_27/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_1_27/buf_output[0] ) );
  NAND4_X2 U8032 ( .A1(\SB1_1_3/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_3/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_3/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_3/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_1_3/buf_output[3] ) );
  NAND4_X2 U8033 ( .A1(\SB1_1_3/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_3/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_3/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_3/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_1_3/buf_output[1] ) );
  NAND4_X2 U8034 ( .A1(\SB1_1_14/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_14/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_14/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_14/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_1_14/buf_output[4] ) );
  NAND4_X2 U8035 ( .A1(\SB1_1_14/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_14/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_14/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_14/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_1_14/buf_output[0] ) );
  NAND4_X2 U8038 ( .A1(\SB1_1_28/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_28/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_28/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_28/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_1_28/buf_output[4] ) );
  NAND4_X2 U8042 ( .A1(\SB1_1_5/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_5/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_5/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_5/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_1_5/buf_output[0] ) );
  NAND4_X2 U8044 ( .A1(\SB1_1_11/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_11/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_11/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_11/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_1_11/buf_output[0] ) );
  NAND4_X2 U8050 ( .A1(\SB1_1_10/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_10/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_10/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_10/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_1_10/buf_output[1] ) );
  BUF_X4 U8057 ( .I(\SB2_1_1/buf_output[4] ), .Z(\RI5[1][190] ) );
  BUF_X4 U8058 ( .I(\SB2_1_1/buf_output[0] ), .Z(\RI5[1][18] ) );
  BUF_X4 U8059 ( .I(\SB2_1_1/buf_output[2] ), .Z(\RI5[1][8] ) );
  BUF_X4 U8060 ( .I(\SB2_1_2/buf_output[2] ), .Z(\RI5[1][2] ) );
  BUF_X4 U8061 ( .I(\SB2_1_2/buf_output[3] ), .Z(\RI5[1][189] ) );
  BUF_X4 U8062 ( .I(\SB2_1_2/buf_output[4] ), .Z(\RI5[1][184] ) );
  BUF_X4 U8065 ( .I(\SB2_1_31/buf_output[5] ), .Z(\RI5[1][5] ) );
  BUF_X4 U8068 ( .I(\SB2_1_0/buf_output[1] ), .Z(\RI5[1][19] ) );
  BUF_X4 U8072 ( .I(\SB2_1_9/buf_output[5] ), .Z(\RI5[1][137] ) );
  NAND4_X2 U8073 ( .A1(\SB1_1_9/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_9/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_9/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_9/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_1_9/buf_output[4] ) );
  NAND4_X2 U8074 ( .A1(\SB1_1_9/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_9/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_9/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_9/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_1_9/buf_output[1] ) );
  BUF_X4 U8075 ( .I(\SB2_1_12/buf_output[0] ), .Z(\RI5[1][144] ) );
  BUF_X4 U8076 ( .I(\SB2_1_12/buf_output[2] ), .Z(\RI5[1][134] ) );
  BUF_X4 U8077 ( .I(\SB2_1_12/buf_output[5] ), .Z(\RI5[1][119] ) );
  BUF_X4 U8078 ( .I(\SB2_1_12/buf_output[4] ), .Z(\RI5[1][124] ) );
  BUF_X4 U8079 ( .I(\SB2_1_13/buf_output[5] ), .Z(\RI5[1][113] ) );
  BUF_X4 U8081 ( .I(\SB2_1_11/buf_output[2] ), .Z(\RI5[1][140] ) );
  BUF_X4 U8082 ( .I(\SB2_1_11/buf_output[4] ), .Z(\RI5[1][130] ) );
  BUF_X4 U8084 ( .I(\SB2_1_15/buf_output[4] ), .Z(\RI5[1][106] ) );
  BUF_X4 U8085 ( .I(\SB2_1_18/buf_output[0] ), .Z(\RI5[1][108] ) );
  BUF_X4 U8086 ( .I(\SB2_1_18/buf_output[5] ), .Z(\RI5[1][83] ) );
  BUF_X4 U8091 ( .I(\SB2_1_17/buf_output[4] ), .Z(\RI5[1][94] ) );
  NAND4_X2 U8092 ( .A1(\SB1_1_21/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_21/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_21/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_21/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_1_21/buf_output[1] ) );
  BUF_X4 U8093 ( .I(\SB2_1_22/buf_output[1] ), .Z(\RI5[1][79] ) );
  BUF_X4 U8094 ( .I(\SB2_1_22/buf_output[5] ), .Z(\RI5[1][59] ) );
  BUF_X4 U8095 ( .I(\SB2_1_23/buf_output[2] ), .Z(\RI5[1][68] ) );
  BUF_X4 U8097 ( .I(\SB2_1_23/buf_output[5] ), .Z(\RI5[1][53] ) );
  NAND4_X2 U8099 ( .A1(\SB1_1_25/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_25/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_25/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_25/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_1_25/buf_output[4] ) );
  BUF_X4 U8101 ( .I(\SB2_1_20/buf_output[5] ), .Z(\RI5[1][71] ) );
  NAND4_X2 U8102 ( .A1(\SB1_1_25/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_25/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_25/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_25/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_1_25/buf_output[0] ) );
  BUF_X4 U8103 ( .I(\SB2_1_21/buf_output[4] ), .Z(\RI5[1][70] ) );
  BUF_X4 U8104 ( .I(\SB2_1_21/buf_output[5] ), .Z(\RI5[1][65] ) );
  NAND4_X2 U8105 ( .A1(\SB1_1_29/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_29/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_1_29/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_1_29/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_1_29/buf_output[4] ) );
  BUF_X4 U8106 ( .I(\SB2_1_24/buf_output[3] ), .Z(\RI5[1][57] ) );
  BUF_X4 U8108 ( .I(\SB2_1_24/buf_output[5] ), .Z(\RI5[1][47] ) );
  BUF_X4 U8109 ( .I(\SB2_1_24/buf_output[4] ), .Z(\RI5[1][52] ) );
  NAND4_X2 U8110 ( .A1(\SB1_1_29/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_1_29/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_29/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_1_29/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_1_29/buf_output[0] ) );
  NAND4_X2 U8113 ( .A1(\SB2_1_28/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_28/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_28/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_1_28/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_1_28/buf_output[4] ) );
  BUF_X4 U8114 ( .I(\SB2_1_29/buf_output[5] ), .Z(\RI5[1][17] ) );
  BUF_X4 U8115 ( .I(\SB2_1_25/buf_output[3] ), .Z(\RI5[1][51] ) );
  BUF_X4 U8119 ( .I(\SB2_0_30/buf_output[5] ), .Z(\RI5[0][11] ) );
  BUF_X4 U8124 ( .I(\SB2_1_3/buf_output[5] ), .Z(\RI5[1][173] ) );
  NAND4_X2 U8130 ( .A1(\SB1_2_20/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_20/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_20/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_20/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_2_20/buf_output[0] ) );
  NAND4_X2 U8134 ( .A1(\SB1_2_28/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_28/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_28/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_28/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_2_28/buf_output[1] ) );
  NAND4_X2 U8139 ( .A1(\SB1_2_1/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_1/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_1/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_1/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_2_1/buf_output[0] ) );
  NAND4_X2 U8145 ( .A1(\SB1_2_5/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_5/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_5/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_5/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_2_5/buf_output[0] ) );
  NAND4_X2 U8146 ( .A1(\SB1_2_30/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_30/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_30/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_30/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_2_30/buf_output[1] ) );
  NAND4_X2 U8147 ( .A1(\SB1_2_0/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_0/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_0/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_0/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_2_0/buf_output[1] ) );
  NAND4_X2 U8148 ( .A1(\SB1_2_6/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_6/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_6/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_6/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_2_6/buf_output[4] ) );
  NAND4_X2 U8155 ( .A1(\SB1_2_23/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_23/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_23/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_23/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_2_23/buf_output[0] ) );
  NAND4_X2 U8157 ( .A1(\SB1_2_3/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_3/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_3/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_3/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_2_3/buf_output[0] ) );
  BUF_X2 U8161 ( .I(\SB2_2_2/buf_output[3] ), .Z(\RI5[2][189] ) );
  BUF_X4 U8162 ( .I(\SB2_2_2/buf_output[5] ), .Z(\RI5[2][179] ) );
  BUF_X4 U8163 ( .I(\SB2_2_2/buf_output[4] ), .Z(\RI5[2][184] ) );
  BUF_X4 U8165 ( .I(\SB2_2_3/buf_output[5] ), .Z(\RI5[2][173] ) );
  NAND4_X2 U8167 ( .A1(\SB2_2_0/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_0/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_2_0/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_2_0/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_2_0/buf_output[4] ) );
  NAND4_X2 U8168 ( .A1(\SB2_2_4/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_4/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_2_4/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_2_4/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_2_4/buf_output[3] ) );
  NAND4_X2 U8173 ( .A1(\SB2_2_8/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_8/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_2_8/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_2_8/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_2_8/buf_output[3] ) );
  BUF_X4 U8174 ( .I(\SB2_2_8/buf_output[0] ), .Z(\RI5[2][168] ) );
  NAND4_X2 U8185 ( .A1(\SB1_2_15/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_15/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_15/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_2_15/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_2_15/buf_output[0] ) );
  BUF_X4 U8188 ( .I(\SB2_2_16/buf_output[2] ), .Z(\RI5[2][110] ) );
  NAND4_X2 U8198 ( .A1(\SB2_2_26/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_26/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_2_26/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_2_26/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_2_26/buf_output[2] ) );
  BUF_X4 U8200 ( .I(\SB2_2_26/buf_output[5] ), .Z(\RI5[2][35] ) );
  NAND4_X2 U8209 ( .A1(\SB1_3_5/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_5/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_5/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_5/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_3_5/buf_output[0] ) );
  NAND4_X2 U8210 ( .A1(\SB1_3_5/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_5/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_5/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_3_5/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_3_5/buf_output[4] ) );
  NAND4_X2 U8211 ( .A1(\SB1_3_10/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_10/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_10/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_3_10/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_3_10/buf_output[4] ) );
  NAND4_X2 U8213 ( .A1(\SB1_3_16/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_16/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_16/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_16/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_3_16/buf_output[0] ) );
  NAND4_X2 U8217 ( .A1(\SB1_3_14/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_14/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_14/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_14/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_3_14/buf_output[1] ) );
  NAND4_X2 U8222 ( .A1(\SB1_3_9/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_9/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_9/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_9/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_3_9/buf_output[1] ) );
  NAND4_X2 U8223 ( .A1(\SB1_3_15/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_15/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_15/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_15/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_3_15/buf_output[0] ) );
  NAND4_X2 U8226 ( .A1(\SB1_3_30/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_30/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_30/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_30/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_3_30/buf_output[0] ) );
  NAND4_X2 U8229 ( .A1(\SB1_3_6/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_3_6/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_6/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_6/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_3_6/buf_output[0] ) );
  BUF_X4 U8233 ( .I(\SB2_3_30/buf_output[4] ), .Z(\RI5[3][16] ) );
  BUF_X4 U8234 ( .I(\SB2_3_30/buf_output[2] ), .Z(\RI5[3][26] ) );
  BUF_X4 U8235 ( .I(\SB2_3_30/buf_output[3] ), .Z(\RI5[3][21] ) );
  BUF_X4 U8236 ( .I(\SB2_3_30/buf_output[5] ), .Z(\RI5[3][11] ) );
  BUF_X4 U8239 ( .I(\SB2_3_1/buf_output[4] ), .Z(\RI5[3][190] ) );
  BUF_X4 U8240 ( .I(\SB2_3_1/buf_output[5] ), .Z(\RI5[3][185] ) );
  NAND4_X2 U8241 ( .A1(\SB1_3_2/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_2/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_2/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_3_2/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_3_2/buf_output[4] ) );
  BUF_X4 U8242 ( .I(\SB2_3_31/buf_output[4] ), .Z(\RI5[3][10] ) );
  BUF_X4 U8245 ( .I(\SB2_3_3/buf_output[2] ), .Z(\RI5[3][188] ) );
  BUF_X4 U8247 ( .I(\SB2_3_3/buf_output[5] ), .Z(\RI5[3][173] ) );
  BUF_X4 U8249 ( .I(\SB2_3_4/buf_output[4] ), .Z(\RI5[3][172] ) );
  BUF_X4 U8251 ( .I(\SB2_3_5/buf_output[5] ), .Z(\RI5[3][161] ) );
  BUF_X4 U8253 ( .I(\SB2_3_6/buf_output[1] ), .Z(\RI5[3][175] ) );
  CLKBUF_X4 U8260 ( .I(\SB2_3_9/buf_output[0] ), .Z(\RI5[3][162] ) );
  BUF_X4 U8262 ( .I(\SB2_3_9/buf_output[5] ), .Z(\RI5[3][137] ) );
  BUF_X4 U8265 ( .I(\SB2_3_10/buf_output[4] ), .Z(\RI5[3][136] ) );
  BUF_X4 U8266 ( .I(\SB2_3_10/buf_output[5] ), .Z(\RI5[3][131] ) );
  BUF_X4 U8267 ( .I(\SB2_3_8/buf_output[2] ), .Z(\RI5[3][158] ) );
  NAND4_X2 U8270 ( .A1(\SB1_3_19/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_3_19/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_19/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_19/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_3_19/buf_output[1] ) );
  BUF_X4 U8272 ( .I(\SB2_3_17/buf_output[4] ), .Z(\RI5[3][94] ) );
  NAND4_X2 U8273 ( .A1(\SB1_3_19/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_19/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_19/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_3_19/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_3_19/buf_output[4] ) );
  BUF_X4 U8275 ( .I(\SB2_3_14/buf_output[4] ), .Z(\RI5[3][112] ) );
  NAND4_X2 U8277 ( .A1(\SB2_3_16/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_3_16/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_16/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_3_16/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_3_16/buf_output[2] ) );
  BUF_X4 U8281 ( .I(\SB2_3_18/buf_output[2] ), .Z(\RI5[3][98] ) );
  BUF_X4 U8282 ( .I(\SB2_3_18/buf_output[0] ), .Z(\RI5[3][108] ) );
  BUF_X4 U8283 ( .I(\SB2_3_18/buf_output[5] ), .Z(\RI5[3][83] ) );
  BUF_X4 U8284 ( .I(\SB2_3_18/buf_output[4] ), .Z(\RI5[3][88] ) );
  CLKBUF_X4 U8285 ( .I(\SB2_3_22/buf_output[0] ), .Z(\RI5[3][84] ) );
  BUF_X4 U8286 ( .I(\SB2_3_27/buf_output[4] ), .Z(\RI5[3][34] ) );
  BUF_X4 U8287 ( .I(\SB2_3_27/buf_output[5] ), .Z(\RI5[3][29] ) );
  BUF_X4 U8289 ( .I(\SB2_3_23/buf_output[2] ), .Z(\RI5[3][68] ) );
  NAND4_X2 U8299 ( .A1(\SB3_7/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_7/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_7/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_7/Component_Function_1/NAND4_in[3] ), .ZN(\SB3_7/buf_output[1] )
         );
  NAND4_X2 U8301 ( .A1(\SB3_0/Component_Function_0/NAND4_in[0] ), .A2(
        \SB3_0/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_0/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_0/Component_Function_0/NAND4_in[3] ), .ZN(\SB3_0/buf_output[0] )
         );
  NAND4_X2 U8302 ( .A1(\SB3_11/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_11/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_11/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_11/Component_Function_1/NAND4_in[3] ), .ZN(\SB3_11/buf_output[1] ) );
  NAND4_X2 U8303 ( .A1(\SB3_11/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_11/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_11/Component_Function_0/NAND4_in[0] ), .A4(
        \SB3_11/Component_Function_0/NAND4_in[3] ), .ZN(\SB3_11/buf_output[0] ) );
  NAND4_X2 U8305 ( .A1(\SB3_17/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_17/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_17/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_17/Component_Function_1/NAND4_in[3] ), .ZN(\SB3_17/buf_output[1] ) );
  NAND4_X2 U8306 ( .A1(\SB3_1/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_1/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_1/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_1/Component_Function_4/NAND4_in[3] ), .ZN(\SB3_1/buf_output[4] )
         );
  NAND4_X2 U8310 ( .A1(\SB3_18/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_18/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_18/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_18/Component_Function_4/NAND4_in[3] ), .ZN(\SB3_18/buf_output[4] ) );
  NAND4_X2 U8311 ( .A1(\SB3_18/Component_Function_0/NAND4_in[0] ), .A2(
        \SB3_18/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_18/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_18/Component_Function_0/NAND4_in[3] ), .ZN(\SB3_18/buf_output[0] ) );
  NAND4_X2 U8314 ( .A1(\SB3_22/Component_Function_0/NAND4_in[0] ), .A2(
        \SB3_22/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_22/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_22/Component_Function_0/NAND4_in[3] ), .ZN(\SB3_22/buf_output[0] ) );
  NAND4_X2 U8317 ( .A1(\SB3_26/Component_Function_0/NAND4_in[0] ), .A2(
        \SB3_26/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_26/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_26/Component_Function_0/NAND4_in[3] ), .ZN(\SB3_26/buf_output[0] ) );
  NAND4_X2 U8318 ( .A1(\SB3_27/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_27/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_27/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_27/Component_Function_4/NAND4_in[3] ), .ZN(\SB3_27/buf_output[4] ) );
  NAND4_X2 U8320 ( .A1(\SB3_27/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_27/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_27/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_27/Component_Function_1/NAND4_in[3] ), .ZN(\SB3_27/buf_output[1] ) );
  NAND4_X2 U8321 ( .A1(\SB3_9/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_9/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_9/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_9/Component_Function_4/NAND4_in[3] ), .ZN(\SB3_9/buf_output[4] )
         );
  NAND4_X2 U8322 ( .A1(\SB3_9/Component_Function_0/NAND4_in[0] ), .A2(
        \SB3_9/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_9/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_9/Component_Function_0/NAND4_in[3] ), .ZN(\SB3_9/buf_output[0] )
         );
  NAND4_X2 U8324 ( .A1(\SB3_15/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_15/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_15/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_15/Component_Function_4/NAND4_in[3] ), .ZN(\SB3_15/buf_output[4] ) );
  NAND4_X2 U8325 ( .A1(\SB3_15/Component_Function_1/NAND4_in[0] ), .A2(
        \SB3_15/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_15/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_15/Component_Function_1/NAND4_in[3] ), .ZN(\SB3_15/buf_output[1] ) );
  NAND4_X2 U8330 ( .A1(\SB3_4/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_4/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_4/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_4/Component_Function_4/NAND4_in[3] ), .ZN(\SB3_4/buf_output[4] )
         );
  NAND4_X2 U8331 ( .A1(\SB3_10/Component_Function_0/NAND4_in[0] ), .A2(
        \SB3_10/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_10/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_10/Component_Function_0/NAND4_in[3] ), .ZN(\SB3_10/buf_output[0] ) );
  NAND4_X2 U8332 ( .A1(\SB3_10/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_10/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_10/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_10/Component_Function_4/NAND4_in[3] ), .ZN(\SB3_10/buf_output[4] ) );
  NAND4_X2 U8335 ( .A1(\SB3_20/Component_Function_0/NAND4_in[0] ), .A2(
        \SB3_20/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_20/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_20/Component_Function_0/NAND4_in[3] ), .ZN(\SB3_20/buf_output[0] ) );
  NAND4_X2 U8338 ( .A1(\SB3_25/Component_Function_0/NAND4_in[0] ), .A2(
        \SB3_25/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_25/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_25/Component_Function_0/NAND4_in[3] ), .ZN(\SB3_25/buf_output[0] ) );
  NAND2_X2 \SB1_0_3/Component_Function_5/N1  ( .A1(\SB1_0_3/i0_0 ), .A2(
        \SB1_0_3/i3[0] ), .ZN(\SB1_0_3/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 \SB2_0_3/BUF_1_0  ( .I(\SB2_0_3/buf_output[1] ), .Z(\RI5[0][1] ) );
  NAND4_X2 \SB2_0_3/Component_Function_1/N5  ( .A1(
        \SB2_0_3/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_3/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_3/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_0_3/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_0_3/buf_output[1] ) );
  NAND3_X2 \SB1_1_7/Component_Function_0/N4  ( .A1(\SB1_1_7/i0[7] ), .A2(
        \SB1_1_7/i0_3 ), .A3(\SB1_1_7/i0_0 ), .ZN(
        \SB1_1_7/Component_Function_0/NAND4_in[3] ) );
  INV_X4 U1728 ( .I(\RI3[0][39] ), .ZN(\SB2_0_25/i0[8] ) );
  NAND3_X2 \SB2_2_3/Component_Function_5/N2  ( .A1(\SB2_2_3/i0_0 ), .A2(
        \SB2_2_3/i0[6] ), .A3(\SB2_2_3/i0[10] ), .ZN(
        \SB2_2_3/Component_Function_5/NAND4_in[1] ) );
  INV_X2 U4934 ( .I(\SB1_3_27/buf_output[5] ), .ZN(\SB2_3_27/i1_5 ) );
  BUF_X4 U4960 ( .I(\SB2_3_8/buf_output[3] ), .Z(\RI5[3][153] ) );
  INV_X2 \SB1_2_15/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[98] ), .ZN(
        \SB1_2_15/i1[9] ) );
  BUF_X2 U1273 ( .I(\MC_ARK_ARC_1_3/buf_output[42] ), .Z(\SB3_24/i0[9] ) );
  NAND3_X2 \SB2_2_29/Component_Function_5/N2  ( .A1(\SB2_2_29/i0_0 ), .A2(
        \SB2_2_29/i0[6] ), .A3(\SB2_2_29/i0[10] ), .ZN(
        \SB2_2_29/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 \SB2_2_0/BUF_3_0  ( .I(\SB2_2_0/buf_output[3] ), .Z(\RI5[2][9] ) );
  INV_X2 \SB1_0_6/INV_3  ( .I(n391), .ZN(\SB1_0_6/i0[8] ) );
  INV_X2 U1773 ( .I(\RI3[0][107] ), .ZN(\SB2_0_14/i1_5 ) );
  BUF_X4 U1355 ( .I(\MC_ARK_ARC_1_1/buf_output[71] ), .Z(\SB1_2_20/i0_3 ) );
  INV_X2 U1744 ( .I(\MC_ARK_ARC_1_1/buf_output[145] ), .ZN(\SB1_2_7/i1_7 ) );
  BUF_X4 \SB1_2_1/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[181] ), .Z(
        \SB1_2_1/i0[6] ) );
  INV_X2 \SB1_2_1/INV_1  ( .I(\MC_ARK_ARC_1_1/buf_output[181] ), .ZN(
        \SB1_2_1/i1_7 ) );
  INV_X2 \SB2_1_14/INV_5  ( .I(\SB1_1_14/buf_output[5] ), .ZN(\SB2_1_14/i1_5 )
         );
  INV_X2 \SB1_3_14/INV_3  ( .I(\MC_ARK_ARC_1_2/buf_output[105] ), .ZN(
        \SB1_3_14/i0[8] ) );
  INV_X2 U1538 ( .I(\MC_ARK_ARC_1_1/buf_output[15] ), .ZN(\SB1_2_29/i0[8] ) );
  BUF_X2 U1188 ( .I(\SB1_3_16/buf_output[0] ), .Z(\SB2_3_11/i0[9] ) );
  NAND4_X2 U4195 ( .A1(\SB2_0_31/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_31/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_31/Component_Function_4/NAND4_in[2] ), .A4(n1297), .ZN(
        \SB2_0_31/buf_output[4] ) );
  NAND4_X2 \SB2_2_25/Component_Function_3/N5  ( .A1(
        \SB2_2_25/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_25/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_2_25/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_2_25/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_2_25/buf_output[3] ) );
  BUF_X4 U1594 ( .I(\MC_ARK_ARC_1_0/buf_output[161] ), .Z(\SB1_1_5/i0_3 ) );
  INV_X2 \SB2_3_19/INV_3  ( .I(\SB1_3_21/buf_output[3] ), .ZN(\SB2_3_19/i0[8] ) );
  NAND3_X2 U2178 ( .A1(\SB3_29/i1_5 ), .A2(\SB3_29/i0_0 ), .A3(\SB3_29/i0_4 ), 
        .ZN(\SB3_29/Component_Function_2/NAND4_in[3] ) );
  INV_X2 \SB1_3_19/INV_5  ( .I(\MC_ARK_ARC_1_2/buf_output[77] ), .ZN(
        \SB1_3_19/i1_5 ) );
  NAND3_X2 U837 ( .A1(\SB2_2_24/i0[10] ), .A2(\SB2_2_24/i0_0 ), .A3(
        \SB2_2_24/i0[6] ), .ZN(\SB2_2_24/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U874 ( .A1(\SB1_2_27/i0_0 ), .A2(\SB1_2_27/i1_5 ), .A3(
        \SB1_2_27/i0_4 ), .ZN(n1801) );
  BUF_X4 \SB1_2_13/BUF_2  ( .I(\MC_ARK_ARC_1_1/buf_output[110] ), .Z(
        \SB1_2_13/i0_0 ) );
  INV_X2 \SB2_2_2/INV_5  ( .I(\SB1_2_2/buf_output[5] ), .ZN(\SB2_2_2/i1_5 ) );
  INV_X2 U1679 ( .I(\MC_ARK_ARC_1_3/buf_output[69] ), .ZN(\SB3_20/i0[8] ) );
  NAND3_X2 \SB3_20/Component_Function_5/N2  ( .A1(\SB3_20/i0_0 ), .A2(
        \SB3_20/i0[6] ), .A3(\SB3_20/i0[10] ), .ZN(
        \SB3_20/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 \SB1_0_31/Component_Function_3/N1  ( .A1(\SB1_0_31/i1[9] ), .A2(
        \SB1_0_31/i0_3 ), .A3(\SB1_0_31/i0[6] ), .ZN(
        \SB1_0_31/Component_Function_3/NAND4_in[0] ) );
  INV_X2 \SB2_3_23/INV_0  ( .I(\SB1_3_28/buf_output[0] ), .ZN(\SB2_3_23/i3[0] ) );
  BUF_X4 U940 ( .I(\SB2_1_10/buf_output[1] ), .Z(\RI5[1][151] ) );
  INV_X2 \SB2_1_24/INV_5  ( .I(\SB1_1_24/buf_output[5] ), .ZN(\SB2_1_24/i1_5 )
         );
  BUF_X4 U669 ( .I(\SB2_3_11/buf_output[0] ), .Z(\RI5[3][150] ) );
  BUF_X4 \SB2_0_5/BUF_1_0  ( .I(\SB2_0_5/buf_output[1] ), .Z(\RI5[0][181] ) );
  INV_X2 \SB1_0_18/INV_3  ( .I(n367), .ZN(\SB1_0_18/i0[8] ) );
  NAND2_X2 \SB1_0_5/Component_Function_5/N1  ( .A1(\SB1_0_5/i0_0 ), .A2(
        \SB1_0_5/i3[0] ), .ZN(\SB1_0_5/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U699 ( .A1(\SB2_3_30/i0_4 ), .A2(\SB2_3_30/i1_5 ), .A3(
        \SB2_3_30/i0_0 ), .ZN(\SB2_3_30/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 \SB2_2_18/Component_Function_5/N3  ( .A1(\SB2_2_18/i1[9] ), .A2(
        \SB2_2_18/i0_4 ), .A3(\SB2_2_18/i0_3 ), .ZN(
        \SB2_2_18/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 \SB1_2_19/Component_Function_4/N4  ( .A1(\SB1_2_19/i1[9] ), .A2(
        \SB1_2_19/i1_5 ), .A3(\SB1_2_19/i0_4 ), .ZN(
        \SB1_2_19/Component_Function_4/NAND4_in[3] ) );
  NAND3_X2 U1517 ( .A1(\SB4_18/i0[10] ), .A2(\SB4_18/i1[9] ), .A3(
        \SB4_18/i1_7 ), .ZN(\SB4_18/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 \SB2_2_18/Component_Function_2/N1  ( .A1(n4769), .A2(
        \SB2_2_18/i0[10] ), .A3(\SB2_2_18/i1[9] ), .ZN(
        \SB2_2_18/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U1701 ( .A1(\SB1_1_7/i0_0 ), .A2(\SB1_1_7/i0_4 ), .A3(
        \SB1_1_7/i1_5 ), .ZN(\SB1_1_7/Component_Function_2/NAND4_in[3] ) );
  BUF_X2 U57 ( .I(Key[47]), .Z(n244) );
  NAND3_X2 U950 ( .A1(\SB2_1_14/i0[10] ), .A2(\SB2_1_14/i0_3 ), .A3(
        \SB2_1_14/i0_4 ), .ZN(\SB2_1_14/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 \SB2_3_5/Component_Function_3/N4  ( .A1(\SB2_3_5/i1_5 ), .A2(
        \SB2_3_5/i0[8] ), .A3(\SB2_3_5/i3[0] ), .ZN(
        \SB2_3_5/Component_Function_3/NAND4_in[3] ) );
  INV_X4 \SB2_3_7/INV_1  ( .I(n1670), .ZN(\SB2_3_7/i1_7 ) );
  NAND4_X2 U1629 ( .A1(\SB2_0_3/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_3/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_3/Component_Function_4/NAND4_in[2] ), .A4(
        \SB2_0_3/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_0_3/buf_output[4] ) );
  NAND3_X2 \SB1_0_9/Component_Function_3/N4  ( .A1(\SB1_0_9/i1_5 ), .A2(
        \SB1_0_9/i0[8] ), .A3(\SB1_0_9/i3[0] ), .ZN(
        \SB1_0_9/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 \SB2_1_26/Component_Function_5/N4  ( .A1(\SB2_1_26/i0[9] ), .A2(
        \SB2_1_26/i0[6] ), .A3(\SB2_1_26/i0_4 ), .ZN(
        \SB2_1_26/Component_Function_5/NAND4_in[3] ) );
  BUF_X4 \SB2_0_21/BUF_1_0  ( .I(\SB2_0_21/buf_output[1] ), .Z(\RI5[0][85] )
         );
  NAND4_X2 \SB2_0_21/Component_Function_1/N5  ( .A1(
        \SB2_0_21/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_0_21/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_0_21/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_0_21/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_0_21/buf_output[1] ) );
  BUF_X4 U666 ( .I(\SB2_3_13/buf_output[0] ), .Z(\RI5[3][138] ) );
  NAND3_X2 \SB2_2_13/Component_Function_5/N2  ( .A1(\SB2_2_13/i0_0 ), .A2(
        \SB2_2_13/i0[6] ), .A3(\SB2_2_13/i0[10] ), .ZN(
        \SB2_2_13/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 U2023 ( .I(\SB1_1_26/buf_output[4] ), .Z(n1579) );
  INV_X2 \SB2_2_28/INV_5  ( .I(\SB1_2_28/buf_output[5] ), .ZN(\SB2_2_28/i1_5 )
         );
  BUF_X4 U4964 ( .I(\MC_ARK_ARC_1_1/buf_output[76] ), .Z(\SB1_2_19/i0_4 ) );
  INV_X2 U1733 ( .I(\MC_ARK_ARC_1_1/buf_output[186] ), .ZN(\SB1_2_0/i3[0] ) );
  BUF_X4 U1064 ( .I(\SB2_0_3/buf_output[4] ), .Z(\RI5[0][178] ) );
  NAND3_X2 \SB2_3_1/Component_Function_3/N1  ( .A1(\SB2_3_1/i1[9] ), .A2(
        \SB2_3_1/i0_3 ), .A3(\SB2_3_1/i0[6] ), .ZN(
        \SB2_3_1/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 \SB1_2_30/Component_Function_1/N4  ( .A1(\SB1_2_30/i1_7 ), .A2(
        \SB1_2_30/i0[8] ), .A3(\SB1_2_30/i0_4 ), .ZN(
        \SB1_2_30/Component_Function_1/NAND4_in[3] ) );
  BUF_X4 U8080 ( .I(\SB2_1_10/buf_output[4] ), .Z(\RI5[1][136] ) );
  BUF_X4 U1747 ( .I(\SB1_1_9/buf_output[5] ), .Z(\SB2_1_9/i0_3 ) );
  INV_X4 \SB2_0_24/INV_1  ( .I(\RI3[0][43] ), .ZN(\SB2_0_24/i1_7 ) );
  NAND3_X2 \SB1_0_5/Component_Function_3/N2  ( .A1(\SB1_0_5/i0_0 ), .A2(
        \SB1_0_5/i0_3 ), .A3(\SB1_0_5/i0_4 ), .ZN(
        \SB1_0_5/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U982 ( .A1(\SB2_1_9/i0[10] ), .A2(\SB2_1_9/i1_5 ), .A3(
        \SB2_1_9/i1[9] ), .ZN(n1538) );
  NAND3_X2 \SB1_2_17/Component_Function_3/N2  ( .A1(\SB1_2_17/i0_0 ), .A2(
        \SB1_2_17/i0_3 ), .A3(\SB1_2_17/i0_4 ), .ZN(
        \SB1_2_17/Component_Function_3/NAND4_in[1] ) );
  INV_X8 \SB1_2_29/INV_5  ( .I(\RI1[2][17] ), .ZN(\SB1_2_29/i1_5 ) );
  BUF_X4 \SB2_2_1/BUF_5  ( .I(\SB1_2_1/buf_output[5] ), .Z(\SB2_2_1/i0_3 ) );
  BUF_X4 \SB1_2_31/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[4] ), .Z(
        \SB1_2_31/i0_4 ) );
  NAND3_X2 \SB2_0_13/Component_Function_1/N2  ( .A1(\SB2_0_13/i0_3 ), .A2(
        \SB2_0_13/i1_7 ), .A3(n1393), .ZN(
        \SB2_0_13/Component_Function_1/NAND4_in[1] ) );
  INV_X2 \SB2_3_6/INV_3  ( .I(\SB1_3_8/buf_output[3] ), .ZN(\SB2_3_6/i0[8] )
         );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_176  ( .I(\SB2_3_5/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[176] ) );
  BUF_X4 U5887 ( .I(\SB2_0_29/buf_output[2] ), .Z(\RI5[0][32] ) );
  NAND4_X2 U5290 ( .A1(\SB2_1_7/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_1_7/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_1_7/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_1_7/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_1_7/buf_output[0] ) );
  INV_X2 \SB2_0_6/INV_5  ( .I(\SB1_0_6/buf_output[5] ), .ZN(\SB2_0_6/i1_5 ) );
  NAND3_X2 \SB3_31/Component_Function_2/N4  ( .A1(\SB3_31/i1_5 ), .A2(
        \SB3_31/i0_0 ), .A3(\SB3_31/i0_4 ), .ZN(
        \SB3_31/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 U1087 ( .A1(n2774), .A2(\SB2_0_19/i0[6] ), .A3(\SB2_0_19/i0_3 ), 
        .ZN(\SB2_0_19/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U5146 ( .A1(\SB2_1_2/i0_3 ), .A2(\SB2_1_2/i0_0 ), .A3(
        \SB2_1_2/i0[7] ), .ZN(n1483) );
  INV_X2 U1470 ( .I(n3657), .ZN(\SB3_24/i1[9] ) );
  BUF_X4 U8107 ( .I(\SB2_1_24/buf_output[1] ), .Z(\RI5[1][67] ) );
  NAND3_X2 \SB2_0_3/Component_Function_3/N3  ( .A1(\SB2_0_3/i1[9] ), .A2(
        \SB2_0_3/i1_7 ), .A3(\SB2_0_3/i0[10] ), .ZN(
        \SB2_0_3/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U1411 ( .A1(\SB1_2_27/i0[10] ), .A2(\SB1_2_27/i0_3 ), .A3(
        \SB1_2_27/i0[6] ), .ZN(\SB1_2_27/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U614 ( .A1(\SB3_13/i0_3 ), .A2(\SB3_13/i1[9] ), .A3(\SB3_13/i0_4 ), 
        .ZN(\SB3_13/Component_Function_5/NAND4_in[2] ) );
  NAND2_X2 \SB1_0_25/Component_Function_5/N1  ( .A1(\SB1_0_25/i0_0 ), .A2(
        \SB1_0_25/i3[0] ), .ZN(\SB1_0_25/Component_Function_5/NAND4_in[0] ) );
  INV_X2 U723 ( .I(\SB1_3_0/buf_output[5] ), .ZN(\SB2_3_0/i1_5 ) );
  BUF_X4 U8268 ( .I(\SB2_3_8/buf_output[1] ), .Z(\RI5[3][163] ) );
  NAND3_X2 \SB1_0_25/Component_Function_2/N3  ( .A1(\SB1_0_25/i0_3 ), .A2(
        \SB1_0_25/i0[8] ), .A3(\SB1_0_25/i0[9] ), .ZN(
        \SB1_0_25/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U1196 ( .A1(\SB2_0_20/i0_3 ), .A2(\SB2_0_20/i0[10] ), .A3(
        \SB2_0_20/i0[6] ), .ZN(\SB2_0_20/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 \SB1_0_24/Component_Function_1/N2  ( .A1(\SB1_0_24/i0_3 ), .A2(
        \SB1_0_24/i1_7 ), .A3(\SB1_0_24/i0[8] ), .ZN(
        \SB1_0_24/Component_Function_1/NAND4_in[1] ) );
  BUF_X4 \SB1_1_26/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[35] ), .Z(
        \SB1_1_26/i0_3 ) );
  NAND4_X2 U6982 ( .A1(\SB2_0_29/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_29/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_29/Component_Function_4/NAND4_in[3] ), .A4(
        \SB2_0_29/Component_Function_4/NAND4_in[2] ), .ZN(
        \SB2_0_29/buf_output[4] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_43  ( .I(\SB2_2_28/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[43] ) );
  BUF_X4 \SB2_0_0/BUF_4_0  ( .I(\SB2_0_0/buf_output[4] ), .Z(\RI5[0][4] ) );
  NAND3_X2 \SB2_0_3/Component_Function_3/N1  ( .A1(\SB2_0_3/i1[9] ), .A2(
        \SB2_0_3/i0_3 ), .A3(\SB2_0_3/i0[6] ), .ZN(
        \SB2_0_3/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 U2035 ( .I(\SB1_1_23/buf_output[5] ), .Z(\SB2_1_23/i0_3 ) );
  NAND3_X2 U4521 ( .A1(\SB1_3_11/i1[9] ), .A2(\SB1_3_11/i0_3 ), .A3(
        \SB1_3_11/i0[6] ), .ZN(\SB1_3_11/Component_Function_3/NAND4_in[0] ) );
  INV_X2 \SB1_3_26/INV_1  ( .I(\MC_ARK_ARC_1_2/buf_output[31] ), .ZN(
        \SB1_3_26/i1_7 ) );
  BUF_X4 U1063 ( .I(\MC_ARK_ARC_1_0/buf_output[83] ), .Z(\SB1_1_18/i0_3 ) );
  NAND3_X2 \SB2_2_31/Component_Function_2/N3  ( .A1(\SB2_2_31/i0_3 ), .A2(
        \SB2_2_31/i0[8] ), .A3(\SB2_2_31/i0[9] ), .ZN(
        \SB2_2_31/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 U1847 ( .I(\MC_ARK_ARC_1_2/buf_output[64] ), .Z(\SB1_3_21/i0_4 ) );
  INV_X2 U734 ( .I(\SB1_3_1/buf_output[5] ), .ZN(\SB2_3_1/i1_5 ) );
  NAND3_X2 U7425 ( .A1(\SB1_1_4/i0_4 ), .A2(\SB1_1_4/i1[9] ), .A3(
        \SB1_1_4/i1_5 ), .ZN(n2584) );
  BUF_X4 U8067 ( .I(\SB2_1_0/buf_output[2] ), .Z(\RI5[1][14] ) );
  INV_X2 U1427 ( .I(\RI3[0][23] ), .ZN(\SB2_0_28/i1_5 ) );
  INV_X4 \SB2_0_11/INV_0  ( .I(n1911), .ZN(\SB2_0_11/i3[0] ) );
  BUF_X4 U1865 ( .I(\SB2_2_0/buf_output[2] ), .Z(n570) );
  NAND3_X2 \SB1_1_28/Component_Function_2/N3  ( .A1(\SB1_1_28/i0_3 ), .A2(
        \SB1_1_28/i0[8] ), .A3(\SB1_1_28/i0[9] ), .ZN(
        \SB1_1_28/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 \SB2_0_28/Component_Function_2/N2  ( .A1(\SB2_0_28/i0_3 ), .A2(
        \SB2_0_28/i0[10] ), .A3(\SB2_0_28/i0[6] ), .ZN(
        \SB2_0_28/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U1066 ( .A1(\SB2_0_28/i0_3 ), .A2(\SB2_0_28/i0_0 ), .A3(
        \RI3[0][22] ), .ZN(\SB2_0_28/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U3504 ( .A1(\SB2_1_3/i0[10] ), .A2(\SB2_1_3/i1[9] ), .A3(
        \SB2_1_3/i1_7 ), .ZN(n1010) );
  BUF_X4 \SB4_18/BUF_3  ( .I(\SB3_20/buf_output[3] ), .Z(\SB4_18/i0[10] ) );
  NAND3_X2 \SB1_2_6/Component_Function_3/N2  ( .A1(\SB1_2_6/i0_0 ), .A2(
        \SB1_2_6/i0_3 ), .A3(\SB1_2_6/i0_4 ), .ZN(
        \SB1_2_6/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U786 ( .A1(\SB1_3_10/i0[10] ), .A2(\SB1_3_10/i1[9] ), .A3(
        \SB1_3_10/i1_7 ), .ZN(n2137) );
  INV_X2 \SB3_24/INV_5  ( .I(\MC_ARK_ARC_1_3/buf_output[47] ), .ZN(
        \SB3_24/i1_5 ) );
  NAND3_X2 \SB2_1_11/Component_Function_3/N4  ( .A1(\SB2_1_11/i1_5 ), .A2(
        \SB2_1_11/i0[8] ), .A3(\SB2_1_11/i3[0] ), .ZN(
        \SB2_1_11/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 \SB1_3_10/Component_Function_4/N4  ( .A1(\SB1_3_10/i1[9] ), .A2(
        \SB1_3_10/i1_5 ), .A3(\SB1_3_10/i0_4 ), .ZN(
        \SB1_3_10/Component_Function_4/NAND4_in[3] ) );
  INV_X2 U1099 ( .I(\SB1_0_17/buf_output[5] ), .ZN(\SB2_0_17/i1_5 ) );
  NAND3_X2 U3976 ( .A1(\SB2_2_8/i0[10] ), .A2(\SB2_2_8/i1_5 ), .A3(
        \SB2_2_8/i1[9] ), .ZN(\SB2_2_8/Component_Function_2/NAND4_in[0] ) );
  INV_X2 U1663 ( .I(\MC_ARK_ARC_1_2/buf_output[74] ), .ZN(\SB1_3_19/i1[9] ) );
  NAND3_X2 \SB2_2_31/Component_Function_2/N4  ( .A1(\SB2_2_31/i1_5 ), .A2(
        \SB2_2_31/i0_0 ), .A3(n569), .ZN(
        \SB2_2_31/Component_Function_2/NAND4_in[3] ) );
  BUF_X4 U8158 ( .I(\SB2_2_1/buf_output[2] ), .Z(\RI5[2][8] ) );
  NAND3_X2 \SB1_0_9/Component_Function_3/N1  ( .A1(\SB1_0_9/i1[9] ), .A2(
        \SB1_0_9/i0_3 ), .A3(\SB1_0_9/i0[6] ), .ZN(
        \SB1_0_9/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 U4703 ( .I(\SB1_2_31/buf_output[5] ), .Z(\SB2_2_31/i0_3 ) );
  NAND3_X2 \SB2_2_7/Component_Function_5/N2  ( .A1(\SB2_2_7/i0_0 ), .A2(
        \SB2_2_7/i0[6] ), .A3(\SB2_2_7/i0[10] ), .ZN(
        \SB2_2_7/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U1607 ( .A1(\SB2_2_7/i0[9] ), .A2(\SB2_2_7/i0[6] ), .A3(
        \SB1_2_8/buf_output[4] ), .ZN(
        \SB2_2_7/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 \SB2_2_0/Component_Function_2/N3  ( .A1(\SB2_2_0/i0_3 ), .A2(
        \SB2_2_0/i0[8] ), .A3(\SB2_2_0/i0[9] ), .ZN(
        \SB2_2_0/Component_Function_2/NAND4_in[2] ) );
  NAND2_X2 \SB1_1_21/Component_Function_5/N1  ( .A1(\SB1_1_21/i0_0 ), .A2(
        \SB1_1_21/i3[0] ), .ZN(\SB1_1_21/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 U1877 ( .I(\SB1_2_3/buf_output[5] ), .Z(\SB2_2_3/i0_3 ) );
  NAND3_X2 \SB1_3_6/Component_Function_5/N2  ( .A1(\SB1_3_6/i0_0 ), .A2(
        \SB1_3_6/i0[6] ), .A3(\SB1_3_6/i0[10] ), .ZN(
        \SB1_3_6/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 U1884 ( .I(\MC_ARK_ARC_1_1/buf_output[171] ), .Z(\SB1_2_3/i0[10] ) );
  NAND2_X1 U3439 ( .A1(\SB1_1_20/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_20/Component_Function_4/NAND4_in[1] ), .ZN(n987) );
  BUF_X4 \SB2_0_19/BUF_3_0  ( .I(\SB2_0_19/buf_output[3] ), .Z(\RI5[0][87] )
         );
  BUF_X4 \SB2_0_4/BUF_4_0  ( .I(\SB2_0_4/buf_output[4] ), .Z(\RI5[0][172] ) );
  BUF_X4 \SB2_0_9/BUF_5  ( .I(\SB1_0_9/buf_output[5] ), .Z(\SB2_0_9/i0_3 ) );
  BUF_X4 \SB2_0_13/BUF_5  ( .I(\RI3[0][113] ), .Z(\SB2_0_13/i0_3 ) );
  BUF_X4 U1929 ( .I(n322), .Z(\SB1_0_6/i0_0 ) );
  BUF_X4 \SB2_2_19/BUF_5  ( .I(\SB1_2_19/buf_output[5] ), .Z(\SB2_2_19/i0_3 )
         );
  NAND3_X2 \SB2_1_31/Component_Function_3/N3  ( .A1(\SB2_1_31/i1[9] ), .A2(
        \SB2_1_31/i1_7 ), .A3(\SB2_1_31/i0[10] ), .ZN(
        \SB2_1_31/Component_Function_3/NAND4_in[2] ) );
  INV_X4 U1104 ( .I(\SB2_0_9/i0[7] ), .ZN(\SB2_0_9/i0_4 ) );
  NAND3_X2 \SB1_2_25/Component_Function_4/N4  ( .A1(\SB1_2_25/i1[9] ), .A2(
        \SB1_2_25/i1_5 ), .A3(\SB1_2_25/i0_4 ), .ZN(
        \SB1_2_25/Component_Function_4/NAND4_in[3] ) );
  INV_X2 U1615 ( .I(\MC_ARK_ARC_1_1/buf_output[23] ), .ZN(\SB1_2_28/i1_5 ) );
  INV_X2 U1313 ( .I(\MC_ARK_ARC_1_1/buf_output[41] ), .ZN(\SB1_2_25/i1_5 ) );
  NAND2_X2 \SB1_2_18/Component_Function_5/N1  ( .A1(\SB1_2_18/i0_0 ), .A2(
        \SB1_2_18/i3[0] ), .ZN(\SB1_2_18/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U2155 ( .A1(\SB2_3_29/i0[10] ), .A2(\SB2_3_29/i0_0 ), .A3(
        \SB2_3_29/i0[6] ), .ZN(\SB2_3_29/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 U1734 ( .I(\SB2_1_15/buf_output[2] ), .Z(\RI5[1][116] ) );
  INV_X2 U1714 ( .I(\MC_ARK_ARC_1_0/buf_output[149] ), .ZN(\SB1_1_7/i1_5 ) );
  NAND2_X2 \SB1_0_21/Component_Function_5/N1  ( .A1(\SB1_0_21/i0_0 ), .A2(
        \SB1_0_21/i3[0] ), .ZN(\SB1_0_21/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 U4803 ( .I(\SB2_2_31/buf_output[1] ), .Z(\RI5[2][25] ) );
  NAND3_X2 U905 ( .A1(\SB1_2_31/i0_3 ), .A2(\SB1_2_31/i1[9] ), .A3(
        \SB1_2_31/i0_4 ), .ZN(\SB1_2_31/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 \SB2_1_28/Component_Function_2/N2  ( .A1(\SB2_1_28/i0_3 ), .A2(
        \SB2_1_28/i0[10] ), .A3(\SB2_1_28/i0[6] ), .ZN(
        \SB2_1_28/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 U1874 ( .I(\SB1_2_30/buf_output[3] ), .Z(\SB2_2_28/i0[10] ) );
  NAND3_X2 \SB1_1_5/Component_Function_2/N3  ( .A1(\SB1_1_5/i0_3 ), .A2(
        \SB1_1_5/i0[8] ), .A3(\SB1_1_5/i0[9] ), .ZN(
        \SB1_1_5/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 \SB2_3_9/Component_Function_5/N2  ( .A1(\SB2_3_9/i0_0 ), .A2(
        \SB2_3_9/i0[6] ), .A3(\SB2_3_9/i0[10] ), .ZN(
        \SB2_3_9/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 \SB3_6/Component_Function_2/N1  ( .A1(\SB3_6/i1_5 ), .A2(
        \SB3_6/i0[10] ), .A3(\SB3_6/i1[9] ), .ZN(
        \SB3_6/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB2_0_3/Component_Function_2/N2  ( .A1(\SB2_0_3/i0_3 ), .A2(
        \SB2_0_3/i0[10] ), .A3(\SB2_0_3/i0[6] ), .ZN(
        \SB2_0_3/Component_Function_2/NAND4_in[1] ) );
  INV_X2 U1267 ( .I(\MC_ARK_ARC_1_3/buf_output[176] ), .ZN(\SB3_2/i1[9] ) );
  BUF_X4 \SB2_1_11/BUF_5  ( .I(\SB1_1_11/buf_output[5] ), .Z(\SB2_1_11/i0_3 )
         );
  NAND2_X2 \SB3_2/Component_Function_5/N1  ( .A1(\SB3_2/i0_0 ), .A2(
        \SB3_2/i3[0] ), .ZN(\SB3_2/Component_Function_5/NAND4_in[0] ) );
  NAND2_X2 \SB2_0_28/Component_Function_5/N1  ( .A1(\SB2_0_28/i0_0 ), .A2(
        \SB2_0_28/i3[0] ), .ZN(\SB2_0_28/Component_Function_5/NAND4_in[0] ) );
  NAND4_X2 U670 ( .A1(\SB2_3_25/Component_Function_0/NAND4_in[2] ), .A2(n2134), 
        .A3(n2133), .A4(\SB2_3_25/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_3_25/buf_output[0] ) );
  NAND2_X2 \SB1_1_20/Component_Function_5/N1  ( .A1(\SB1_1_20/i0_0 ), .A2(
        \SB1_1_20/i3[0] ), .ZN(\SB1_1_20/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U3365 ( .A1(\SB2_2_23/i0_4 ), .A2(\SB2_2_23/i1_7 ), .A3(
        \SB2_2_23/i0[8] ), .ZN(n964) );
  NAND2_X2 \SB3_30/Component_Function_5/N1  ( .A1(\SB3_30/i0_0 ), .A2(
        \SB3_30/i3[0] ), .ZN(\SB3_30/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 U1614 ( .I(\MC_ARK_ARC_1_1/buf_output[23] ), .Z(\SB1_2_28/i0_3 ) );
  BUF_X4 U4935 ( .I(\SB1_3_27/buf_output[5] ), .Z(\SB2_3_27/i0_3 ) );
  BUF_X4 \SB2_0_14/BUF_5  ( .I(\RI3[0][107] ), .Z(\SB2_0_14/i0_3 ) );
  BUF_X4 U1799 ( .I(\SB3_2/buf_output[5] ), .Z(\SB4_2/i0_3 ) );
  NAND3_X2 U3883 ( .A1(\SB2_1_12/i0_3 ), .A2(\SB2_1_12/i0_4 ), .A3(
        \SB2_1_12/i0[10] ), .ZN(n1159) );
  NAND2_X2 \SB1_1_10/Component_Function_5/N1  ( .A1(\SB1_1_10/i0_0 ), .A2(
        \SB1_1_10/i3[0] ), .ZN(\SB1_1_10/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 U8264 ( .I(\SB2_3_10/buf_output[2] ), .Z(\RI5[3][146] ) );
  NAND2_X2 \SB2_1_28/Component_Function_5/N1  ( .A1(\SB2_1_28/i0_0 ), .A2(
        \SB2_1_28/i3[0] ), .ZN(\SB2_1_28/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB1_2_23/Component_Function_4/N4  ( .A1(\SB1_2_23/i1[9] ), .A2(
        \SB1_2_23/i1_5 ), .A3(\SB1_2_23/i0_4 ), .ZN(
        \SB1_2_23/Component_Function_4/NAND4_in[3] ) );
  NAND3_X2 \SB1_2_7/Component_Function_5/N2  ( .A1(\SB1_2_7/i0_0 ), .A2(
        \SB1_2_7/i0[6] ), .A3(\SB1_2_7/i0[10] ), .ZN(
        \SB1_2_7/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U4921 ( .A1(\SB2_3_6/i0[9] ), .A2(\SB2_3_6/i0_3 ), .A3(
        \SB2_3_6/i0[8] ), .ZN(\SB2_3_6/Component_Function_2/NAND4_in[2] ) );
  INV_X4 U1103 ( .I(\SB2_0_28/i0[7] ), .ZN(\RI3[0][22] ) );
  CLKBUF_X4 \SB2_2_30/BUF_2  ( .I(\SB1_2_1/buf_output[2] ), .Z(\SB2_2_30/i0_0 ) );
  BUF_X2 U190 ( .I(Key[105]), .Z(n138) );
  BUF_X4 \SB2_1_15/BUF_5  ( .I(\SB1_1_15/buf_output[5] ), .Z(\SB2_1_15/i0_3 )
         );
  BUF_X4 \SB2_0_7/BUF_5  ( .I(\RI3[0][149] ), .Z(\SB2_0_7/i0_3 ) );
  BUF_X4 \SB2_1_14/BUF_4  ( .I(\SB1_1_15/buf_output[4] ), .Z(\SB2_1_14/i0_4 )
         );
  BUF_X2 U1230 ( .I(\SB3_29/buf_output[3] ), .Z(\SB4_27/i0[10] ) );
  INV_X2 \SB2_2_22/INV_5  ( .I(\SB1_2_22/buf_output[5] ), .ZN(\SB2_2_22/i1_5 )
         );
  INV_X2 \SB1_1_9/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[133] ), .ZN(
        \SB1_1_9/i1_7 ) );
  NAND3_X2 U980 ( .A1(\SB2_1_9/i0_4 ), .A2(\SB2_1_9/i0_3 ), .A3(
        \SB2_1_9/i1[9] ), .ZN(n1436) );
  NAND3_X2 \SB2_2_6/Component_Function_2/N3  ( .A1(\SB2_2_6/i0_3 ), .A2(
        \SB2_2_6/i0[8] ), .A3(\SB2_2_6/i0[9] ), .ZN(
        \SB2_2_6/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 U1713 ( .I(\MC_ARK_ARC_1_0/buf_output[149] ), .Z(\SB1_1_7/i0_3 ) );
  NAND3_X2 \SB2_1_9/Component_Function_2/N3  ( .A1(\SB2_1_9/i0_3 ), .A2(
        \SB2_1_9/i0[8] ), .A3(\SB2_1_9/i0[9] ), .ZN(
        \SB2_1_9/Component_Function_2/NAND4_in[2] ) );
  INV_X2 \SB1_1_9/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[137] ), .ZN(
        \SB1_1_9/i1_5 ) );
  NAND2_X2 U2003 ( .A1(\SB1_1_9/i0_0 ), .A2(\SB1_1_9/i3[0] ), .ZN(
        \SB1_1_9/Component_Function_5/NAND4_in[0] ) );
  NAND2_X2 \SB2_2_13/Component_Function_5/N1  ( .A1(\SB2_2_13/i0_0 ), .A2(
        \SB2_2_13/i3[0] ), .ZN(\SB2_2_13/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_115  ( .I(\SB2_0_16/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[115] ) );
  NAND4_X2 \SB2_0_16/Component_Function_1/N5  ( .A1(
        \SB2_0_16/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_16/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_16/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_16/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_0_16/buf_output[1] ) );
  NAND3_X2 U1037 ( .A1(\SB1_1_12/i0[10] ), .A2(\SB1_1_12/i0_0 ), .A3(
        \SB1_1_12/i0[6] ), .ZN(\SB1_1_12/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 \SB2_1_8/BUF_5  ( .I(\SB1_1_8/buf_output[5] ), .Z(\SB2_1_8/i0_3 ) );
  NAND3_X2 U1043 ( .A1(\SB1_1_18/i0_4 ), .A2(\SB1_1_18/i0[9] ), .A3(
        \SB1_1_18/i0[6] ), .ZN(\SB1_1_18/Component_Function_5/NAND4_in[3] ) );
  NAND2_X2 \SB1_1_6/Component_Function_5/N1  ( .A1(\SB1_1_6/i0_0 ), .A2(
        \SB1_1_6/i3[0] ), .ZN(\SB1_1_6/Component_Function_5/NAND4_in[0] ) );
  BUF_X2 U153 ( .I(Key[165]), .Z(n203) );
  NAND2_X2 \SB2_3_7/Component_Function_5/N1  ( .A1(\SB2_3_7/i0_0 ), .A2(
        \SB2_3_7/i3[0] ), .ZN(\SB2_3_7/Component_Function_5/NAND4_in[0] ) );
  INV_X2 \SB1_1_14/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[104] ), .ZN(
        \SB1_1_14/i1[9] ) );
  INV_X2 U4567 ( .I(\SB1_3_8/buf_output[5] ), .ZN(\SB2_3_8/i1_5 ) );
  NAND3_X2 \SB2_2_13/Component_Function_5/N4  ( .A1(\SB2_2_13/i0[9] ), .A2(
        \SB2_2_13/i0[6] ), .A3(n580), .ZN(
        \SB2_2_13/Component_Function_5/NAND4_in[3] ) );
  BUF_X2 \SB2_1_15/BUF_1  ( .I(\SB1_1_19/buf_output[1] ), .Z(\SB2_1_15/i0[6] )
         );
  BUF_X4 \SB2_0_18/BUF_0_0  ( .I(\SB2_0_18/buf_output[0] ), .Z(\RI5[0][108] )
         );
  NAND3_X2 U942 ( .A1(\SB2_1_12/i0_3 ), .A2(\SB2_1_12/i0_0 ), .A3(
        \SB2_1_12/i0_4 ), .ZN(\SB2_1_12/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U738 ( .A1(\SB1_3_8/i0_3 ), .A2(\SB1_3_8/i1[9] ), .A3(
        \SB1_3_8/i0_4 ), .ZN(\SB1_3_8/Component_Function_5/NAND4_in[2] ) );
  BUF_X4 U4568 ( .I(\SB1_3_8/buf_output[5] ), .Z(\SB2_3_8/i0_3 ) );
  BUF_X2 U105 ( .I(Key[10]), .Z(n170) );
  NAND2_X2 \SB1_2_27/Component_Function_5/N1  ( .A1(\SB1_2_27/i0_0 ), .A2(
        \SB1_2_27/i3[0] ), .ZN(\SB1_2_27/Component_Function_5/NAND4_in[0] ) );
  NAND2_X2 \SB2_1_21/Component_Function_1/N1  ( .A1(\SB2_1_21/i0_3 ), .A2(
        \SB2_1_21/i1[9] ), .ZN(\SB2_1_21/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 U4441 ( .A1(\SB2_0_17/i0[7] ), .A2(\SB2_0_17/i0[8] ), .A3(
        \SB2_0_17/i0[6] ), .ZN(n1697) );
  NAND3_X2 \SB1_1_13/Component_Function_3/N2  ( .A1(\SB1_1_13/i0_0 ), .A2(
        \SB1_1_13/i0_3 ), .A3(\SB1_1_13/i0_4 ), .ZN(
        \SB1_1_13/Component_Function_3/NAND4_in[1] ) );
  CLKBUF_X4 U4433 ( .I(\MC_ARK_ARC_1_3/buf_output[117] ), .Z(\SB3_12/i0[10] )
         );
  NAND3_X2 U3696 ( .A1(\SB2_3_29/i0_3 ), .A2(\SB2_3_29/i0[6] ), .A3(
        \SB2_3_29/i1[9] ), .ZN(\SB2_3_29/Component_Function_3/NAND4_in[0] ) );
  INV_X2 U4432 ( .I(\MC_ARK_ARC_1_3/buf_output[117] ), .ZN(\SB3_12/i0[8] ) );
  NAND3_X2 \SB1_2_10/Component_Function_1/N4  ( .A1(\SB1_2_10/i1_7 ), .A2(
        \SB1_2_10/i0[8] ), .A3(\SB1_2_10/i0_4 ), .ZN(
        \SB1_2_10/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 U2091 ( .A1(\SB2_2_9/i1[9] ), .A2(n3687), .A3(\SB2_2_9/i0_4 ), .ZN(
        \SB2_2_9/Component_Function_4/NAND4_in[3] ) );
  NAND2_X2 \SB1_1_11/Component_Function_5/N1  ( .A1(\SB1_1_11/i0_0 ), .A2(
        \SB1_1_11/i3[0] ), .ZN(\SB1_1_11/Component_Function_5/NAND4_in[0] ) );
  INV_X2 \SB1_1_27/INV_2  ( .I(\MC_ARK_ARC_1_0/buf_output[26] ), .ZN(
        \SB1_1_27/i1[9] ) );
  BUF_X2 U136 ( .I(Key[56]), .Z(n198) );
  BUF_X4 \SB2_0_3/BUF_5  ( .I(\SB1_0_3/buf_output[5] ), .Z(\SB2_0_3/i0_3 ) );
  INV_X2 U2140 ( .I(\SB1_3_22/buf_output[5] ), .ZN(\SB2_3_22/i1_5 ) );
  INV_X2 U1284 ( .I(\MC_ARK_ARC_1_3/buf_output[27] ), .ZN(\SB3_27/i0[8] ) );
  NAND3_X2 \SB1_1_22/Component_Function_3/N4  ( .A1(\SB1_1_22/i1_5 ), .A2(
        \SB1_1_22/i0[8] ), .A3(\SB1_1_22/i3[0] ), .ZN(
        \SB1_1_22/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 \SB1_3_8/Component_Function_5/N2  ( .A1(\SB1_3_8/i0_0 ), .A2(
        \SB1_3_8/i0[6] ), .A3(\SB1_3_8/i0[10] ), .ZN(
        \SB1_3_8/Component_Function_5/NAND4_in[1] ) );
  BUF_X2 U140 ( .I(Key[57]), .Z(n122) );
  BUF_X4 \SB2_2_6/BUF_5  ( .I(\SB1_2_6/buf_output[5] ), .Z(\SB2_2_6/i0_3 ) );
  NAND3_X2 \SB2_2_2/Component_Function_5/N2  ( .A1(\SB2_2_2/i0_0 ), .A2(
        \SB2_2_2/i0[6] ), .A3(\SB2_2_2/i0[10] ), .ZN(
        \SB2_2_2/Component_Function_5/NAND4_in[1] ) );
  INV_X2 U1510 ( .I(\MC_ARK_ARC_1_1/buf_output[27] ), .ZN(\SB1_2_27/i0[8] ) );
  NAND3_X2 \SB2_1_2/Component_Function_3/N3  ( .A1(\SB2_1_2/i1[9] ), .A2(
        \SB2_1_2/i1_7 ), .A3(\SB2_1_2/i0[10] ), .ZN(
        \SB2_1_2/Component_Function_3/NAND4_in[2] ) );
  BUF_X2 U88 ( .I(Key[90]), .Z(n30) );
  INV_X2 \SB2_3_25/INV_5  ( .I(\SB1_3_25/buf_output[5] ), .ZN(\SB2_3_25/i1_5 )
         );
  INV_X2 U1228 ( .I(\MC_ARK_ARC_1_1/buf_output[74] ), .ZN(\SB1_2_19/i1[9] ) );
  INV_X2 \SB1_1_1/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[185] ), .ZN(
        \SB1_1_1/i1_5 ) );
  NAND3_X2 \SB1_1_22/Component_Function_2/N2  ( .A1(\RI1[1][59] ), .A2(
        \SB1_1_22/i0[10] ), .A3(\SB1_1_22/i0[6] ), .ZN(
        \SB1_1_22/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U1137 ( .A1(\SB1_0_27/i0_3 ), .A2(\SB1_0_27/i0_4 ), .A3(
        \SB1_0_27/i1[9] ), .ZN(n2210) );
  BUF_X4 \SB2_0_5/BUF_2_0  ( .I(\SB2_0_5/buf_output[2] ), .Z(\RI5[0][176] ) );
  BUF_X2 \SB2_0_17/BUF_0  ( .I(\RI3[0][84] ), .Z(\SB2_0_17/i0[9] ) );
  CLKBUF_X4 \SB2_1_16/BUF_1  ( .I(\SB1_1_20/buf_output[1] ), .Z(
        \SB2_1_16/i0[6] ) );
  CLKBUF_X4 \SB1_1_27/BUF_2  ( .I(\MC_ARK_ARC_1_0/buf_output[26] ), .Z(
        \SB1_1_27/i0_0 ) );
  NAND3_X2 \SB2_2_12/Component_Function_2/N1  ( .A1(\SB2_2_12/i1_5 ), .A2(
        \SB2_2_12/i0[10] ), .A3(\SB2_2_12/i1[9] ), .ZN(
        \SB2_2_12/Component_Function_2/NAND4_in[0] ) );
  INV_X2 U2271 ( .I(\SB1_2_12/buf_output[5] ), .ZN(\SB2_2_12/i1_5 ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_49  ( .I(\SB2_3_27/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[49] ) );
  NAND3_X2 \SB2_1_24/Component_Function_3/N1  ( .A1(\SB2_1_24/i1[9] ), .A2(
        \SB2_1_24/i0_3 ), .A3(\SB2_1_24/i0[6] ), .ZN(
        \SB2_1_24/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_56  ( .I(\SB2_2_25/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[56] ) );
  NAND3_X2 \SB1_1_7/Component_Function_0/N3  ( .A1(\SB1_1_7/i0[10] ), .A2(
        \SB1_1_7/i0_4 ), .A3(\SB1_1_7/i0_3 ), .ZN(
        \SB1_1_7/Component_Function_0/NAND4_in[2] ) );
  INV_X2 U1466 ( .I(n393), .ZN(\SB1_0_5/i0[8] ) );
  BUF_X4 U1866 ( .I(\SB1_2_12/buf_output[5] ), .Z(\SB2_2_12/i0_3 ) );
  BUF_X2 U179 ( .I(Key[123]), .Z(n213) );
  BUF_X2 U36 ( .I(Key[25]), .Z(n115) );
  NAND3_X2 \SB1_3_23/Component_Function_2/N2  ( .A1(\SB1_3_23/i0_3 ), .A2(
        \SB1_3_23/i0[10] ), .A3(\SB1_3_23/i0[6] ), .ZN(
        \SB1_3_23/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U1193 ( .A1(\SB2_0_20/i0[9] ), .A2(\SB2_0_20/i0_3 ), .A3(
        \SB2_0_20/i0[8] ), .ZN(\SB2_0_20/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U856 ( .A1(\SB2_2_12/i0[10] ), .A2(\SB2_2_12/i1_7 ), .A3(
        \SB2_2_12/i1[9] ), .ZN(\SB2_2_12/Component_Function_3/NAND4_in[2] ) );
  BUF_X4 U1811 ( .I(\SB2_3_7/buf_output[1] ), .Z(\RI5[3][169] ) );
  BUF_X4 U1852 ( .I(\SB2_2_24/buf_output[1] ), .Z(\RI5[2][67] ) );
  INV_X2 U2684 ( .I(\SB1_2_8/buf_output[1] ), .ZN(\SB2_2_4/i1_7 ) );
  NAND3_X2 U7852 ( .A1(\SB2_1_10/i0[9] ), .A2(\SB1_1_11/buf_output[4] ), .A3(
        \SB2_1_10/i0[6] ), .ZN(\SB2_1_10/Component_Function_5/NAND4_in[3] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_66  ( .I(\SB2_1_25/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[66] ) );
  NAND4_X2 U6036 ( .A1(\SB2_1_25/Component_Function_0/NAND4_in[2] ), .A2(n2744), .A3(\SB2_1_25/Component_Function_0/NAND4_in[0] ), .A4(n2743), .ZN(
        \SB2_1_25/buf_output[0] ) );
  NAND3_X2 U1334 ( .A1(\SB2_2_5/i0_0 ), .A2(\SB2_2_5/i1_5 ), .A3(
        \SB2_2_5/i0_4 ), .ZN(n1881) );
  BUF_X4 U1308 ( .I(\MC_ARK_ARC_1_0/buf_output[95] ), .Z(\SB1_1_16/i0_3 ) );
  NAND3_X2 \SB2_2_12/Component_Function_3/N1  ( .A1(\SB2_2_12/i1[9] ), .A2(
        \SB2_2_12/i0_3 ), .A3(\SB2_2_12/i0[6] ), .ZN(
        \SB2_2_12/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U976 ( .A1(\SB2_1_28/i0_3 ), .A2(\SB2_1_28/i0[10] ), .A3(
        \SB2_1_28/i0_4 ), .ZN(n1740) );
  NAND2_X2 \SB1_1_28/Component_Function_5/N1  ( .A1(\SB1_1_28/i0_0 ), .A2(
        \SB1_1_28/i3[0] ), .ZN(\SB1_1_28/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB1_3_23/Component_Function_2/N1  ( .A1(\SB1_3_23/i1_5 ), .A2(
        \SB1_3_23/i0[10] ), .A3(\SB1_3_23/i1[9] ), .ZN(
        \SB1_3_23/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U4657 ( .A1(\SB1_0_6/i0_3 ), .A2(\SB1_0_6/i1_7 ), .A3(
        \SB1_0_6/i0[8] ), .ZN(\SB1_0_6/Component_Function_1/NAND4_in[1] ) );
  NAND3_X2 \SB2_0_8/Component_Function_2/N2  ( .A1(\SB2_0_8/i0_3 ), .A2(
        \SB2_0_8/i0[10] ), .A3(\SB2_0_8/i0[6] ), .ZN(
        \SB2_0_8/Component_Function_2/NAND4_in[1] ) );
  NAND2_X2 U865 ( .A1(\SB1_2_0/Component_Function_4/NAND4_in[2] ), .A2(n1949), 
        .ZN(n1948) );
  BUF_X2 U184 ( .I(Key[113]), .Z(n229) );
  BUF_X4 \SB2_0_9/BUF_0_0  ( .I(\SB2_0_9/buf_output[0] ), .Z(\RI5[0][162] ) );
  INV_X2 U1605 ( .I(\MC_ARK_ARC_1_3/buf_output[75] ), .ZN(\SB3_19/i0[8] ) );
  NAND3_X2 \SB2_0_29/Component_Function_5/N2  ( .A1(\SB2_0_29/i0_0 ), .A2(
        \SB2_0_29/i0[6] ), .A3(\RI3[0][15] ), .ZN(
        \SB2_0_29/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 \SB1_2_18/Component_Function_5/N4  ( .A1(\SB1_2_18/i0[9] ), .A2(
        \SB1_2_18/i0[6] ), .A3(\SB1_2_18/i0_4 ), .ZN(
        \SB1_2_18/Component_Function_5/NAND4_in[3] ) );
  BUF_X4 \SB2_3_15/BUF_5  ( .I(\SB1_3_15/buf_output[5] ), .Z(\SB2_3_15/i0_3 )
         );
  NAND3_X2 \SB2_2_18/Component_Function_0/N2  ( .A1(\SB2_2_18/i0[8] ), .A2(
        \SB2_2_18/i0[7] ), .A3(\SB2_2_18/i0[6] ), .ZN(
        \SB2_2_18/Component_Function_0/NAND4_in[1] ) );
  BUF_X4 U1876 ( .I(\SB1_2_29/buf_output[5] ), .Z(\SB2_2_29/i0_3 ) );
  NAND3_X2 \SB2_3_15/Component_Function_2/N1  ( .A1(\SB2_3_15/i1_5 ), .A2(
        \SB2_3_15/i0[10] ), .A3(\SB2_3_15/i1[9] ), .ZN(
        \SB2_3_15/Component_Function_2/NAND4_in[0] ) );
  INV_X2 U4500 ( .I(\SB1_2_22/buf_output[1] ), .ZN(\SB2_2_18/i1_7 ) );
  BUF_X2 U112 ( .I(Key[164]), .Z(n195) );
  BUF_X2 \SB2_2_2/BUF_3  ( .I(\SB1_2_4/buf_output[3] ), .Z(\SB2_2_2/i0[10] )
         );
  INV_X2 U4435 ( .I(\SB3_31/buf_output[3] ), .ZN(\SB4_29/i0[8] ) );
  BUF_X4 \SB2_0_5/BUF_0_0  ( .I(\SB2_0_5/buf_output[0] ), .Z(\RI5[0][186] ) );
  NAND4_X2 U2958 ( .A1(n1422), .A2(\SB2_0_5/Component_Function_0/NAND4_in[3] ), 
        .A3(\SB2_0_5/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_5/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_0_5/buf_output[0] ) );
  NAND3_X2 \SB1_2_18/Component_Function_2/N3  ( .A1(\SB1_2_18/i0_3 ), .A2(
        n4762), .A3(\SB1_2_18/i0[9] ), .ZN(
        \SB1_2_18/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 \SB1_0_30/BUF_5  ( .I(n406), .Z(\SB1_0_30/i0_3 ) );
  NAND3_X2 U775 ( .A1(\SB1_3_8/i0[10] ), .A2(\SB1_3_8/i1[9] ), .A3(
        \SB1_3_8/i1_7 ), .ZN(\SB1_3_8/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 \SB1_2_21/Component_Function_3/N4  ( .A1(\SB1_2_21/i1_5 ), .A2(
        \SB1_2_21/i0[8] ), .A3(\SB1_2_21/i3[0] ), .ZN(
        \SB1_2_21/Component_Function_3/NAND4_in[3] ) );
  INV_X4 U735 ( .I(n1319), .ZN(\SB1_3_8/buf_output[4] ) );
  NAND3_X2 \SB2_3_3/Component_Function_3/N2  ( .A1(\SB2_3_3/i0_0 ), .A2(
        \SB2_3_3/i0_3 ), .A3(\SB2_3_3/i0_4 ), .ZN(
        \SB2_3_3/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 \SB2_1_31/Component_Function_2/N1  ( .A1(n5510), .A2(
        \SB2_1_31/i0[10] ), .A3(\SB2_1_31/i1[9] ), .ZN(
        \SB2_1_31/Component_Function_2/NAND4_in[0] ) );
  CLKBUF_X2 U34 ( .I(Key[58]), .Z(n217) );
  INV_X2 U3396 ( .I(\SB1_0_19/buf_output[5] ), .ZN(\SB2_0_19/i1_5 ) );
  NAND3_X2 U1013 ( .A1(\SB1_1_10/i0[9] ), .A2(\SB1_1_10/i0_4 ), .A3(
        \SB1_1_10/i0[6] ), .ZN(n1066) );
  BUF_X4 U4600 ( .I(n1381), .Z(\SB3_11/i0_3 ) );
  BUF_X4 U1917 ( .I(\SB2_0_12/buf_output[2] ), .Z(\RI5[0][134] ) );
  CLKBUF_X4 \SB2_2_26/BUF_3  ( .I(\SB1_2_28/buf_output[3] ), .Z(
        \SB2_2_26/i0[10] ) );
  INV_X2 U1572 ( .I(\MC_ARK_ARC_1_1/buf_output[21] ), .ZN(\SB1_2_28/i0[8] ) );
  NAND3_X2 U2040 ( .A1(\SB2_1_3/i1_5 ), .A2(\SB2_1_3/i0[8] ), .A3(
        \SB2_1_3/i3[0] ), .ZN(\SB2_1_3/Component_Function_3/NAND4_in[3] ) );
  NAND2_X2 \SB1_2_0/Component_Function_0/N1  ( .A1(\SB1_2_0/i0[10] ), .A2(
        \SB1_2_0/i0[9] ), .ZN(\SB1_2_0/Component_Function_0/NAND4_in[0] ) );
  NAND3_X2 U1069 ( .A1(\SB2_0_24/i0[10] ), .A2(\SB2_0_24/i1_5 ), .A3(
        \SB2_0_24/i1[9] ), .ZN(n1790) );
  INV_X2 \SB2_3_15/INV_5  ( .I(\SB1_3_15/buf_output[5] ), .ZN(\SB2_3_15/i1_5 )
         );
  BUF_X4 \SB2_0_19/BUF_1_0  ( .I(\SB2_0_19/buf_output[1] ), .Z(\RI5[0][97] )
         );
  NAND4_X2 U3056 ( .A1(\SB2_0_19/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_0_19/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_19/Component_Function_1/NAND4_in[0] ), .A4(
        \SB2_0_19/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_0_19/buf_output[1] ) );
  NAND2_X2 \SB1_3_12/Component_Function_5/N1  ( .A1(\SB1_3_12/i0_0 ), .A2(
        \SB1_3_12/i3[0] ), .ZN(\SB1_3_12/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 U8279 ( .I(\SB2_3_21/buf_output[4] ), .Z(\RI5[3][70] ) );
  INV_X2 U1185 ( .I(\MC_ARK_ARC_1_1/buf_output[26] ), .ZN(\SB1_2_27/i1[9] ) );
  BUF_X4 U4662 ( .I(\SB1_2_31/buf_output[1] ), .Z(\SB2_2_27/i0[6] ) );
  NAND3_X2 U2041 ( .A1(\SB2_1_24/i1_5 ), .A2(\SB2_1_24/i0[8] ), .A3(
        \SB2_1_24/i3[0] ), .ZN(\SB2_1_24/Component_Function_3/NAND4_in[3] ) );
  BUF_X4 \SB2_3_0/BUF_5  ( .I(\SB1_3_0/buf_output[5] ), .Z(\SB2_3_0/i0_3 ) );
  NAND3_X2 \SB2_1_20/Component_Function_2/N3  ( .A1(\SB2_1_20/i0_3 ), .A2(
        \SB2_1_20/i0[8] ), .A3(\SB2_1_20/i0[9] ), .ZN(
        \SB2_1_20/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 \SB1_1_19/Component_Function_2/N1  ( .A1(\SB1_1_19/i1_5 ), .A2(
        \SB1_1_19/i0[10] ), .A3(\SB1_1_19/i1[9] ), .ZN(
        \SB1_1_19/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 U1812 ( .I(\SB2_3_15/buf_output[1] ), .Z(\RI5[3][121] ) );
  NAND3_X2 \SB2_3_15/Component_Function_3/N2  ( .A1(\SB2_3_15/i0_0 ), .A2(
        \SB2_3_15/i0_3 ), .A3(\SB1_3_16/buf_output[4] ), .ZN(
        \SB2_3_15/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_31/Component_Function_3/N4  ( .A1(\SB2_3_31/i1_5 ), .A2(
        \SB2_3_31/i0[8] ), .A3(\SB2_3_31/i3[0] ), .ZN(
        \SB2_3_31/Component_Function_3/NAND4_in[3] ) );
  INV_X4 U3876 ( .I(\SB2_1_4/i0[7] ), .ZN(\SB1_1_5/buf_output[4] ) );
  BUF_X4 U4805 ( .I(\SB2_1_9/buf_output[1] ), .Z(\RI5[1][157] ) );
  NAND3_X2 \SB1_2_8/Component_Function_2/N2  ( .A1(\SB1_2_8/i0_3 ), .A2(
        \SB1_2_8/i0[10] ), .A3(\SB1_2_8/i0[6] ), .ZN(
        \SB1_2_8/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 U6890 ( .I(\SB2_3_22/buf_output[1] ), .Z(\RI5[3][79] ) );
  NAND4_X2 \SB2_3_22/Component_Function_1/N5  ( .A1(
        \SB2_3_22/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_22/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_22/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_22/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_3_22/buf_output[1] ) );
  NAND3_X2 \SB2_1_19/Component_Function_5/N2  ( .A1(\SB1_1_22/buf_output[2] ), 
        .A2(\SB2_1_19/i0[6] ), .A3(\SB2_1_19/i0[10] ), .ZN(
        \SB2_1_19/Component_Function_5/NAND4_in[1] ) );
  INV_X2 U1588 ( .I(\MC_ARK_ARC_1_1/buf_output[158] ), .ZN(\SB1_2_5/i1[9] ) );
  BUF_X2 U63 ( .I(Key[9]), .Z(n196) );
  BUF_X2 U102 ( .I(Key[146]), .Z(n100) );
  BUF_X4 \SB1_2_5/BUF_2  ( .I(\MC_ARK_ARC_1_1/buf_output[158] ), .Z(
        \SB1_2_5/i0_0 ) );
  INV_X2 \SB1_0_9/INV_3  ( .I(n385), .ZN(\SB1_0_9/i0[8] ) );
  BUF_X4 \SB2_0_7/BUF_3  ( .I(\RI3[0][147] ), .Z(\SB2_0_7/i0[10] ) );
  BUF_X4 U8328 ( .I(\SB2_3_28/buf_output[1] ), .Z(\RI5[3][43] ) );
  NAND4_X2 \SB2_3_28/Component_Function_1/N5  ( .A1(
        \SB2_3_28/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_28/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_28/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_28/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_3_28/buf_output[1] ) );
  INV_X2 U6267 ( .I(\SB1_3_9/buf_output[5] ), .ZN(\SB2_3_9/i1_5 ) );
  NAND4_X2 \SB2_3_9/Component_Function_3/N5  ( .A1(
        \SB2_3_9/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_9/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_9/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_9/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_3_9/buf_output[3] ) );
  BUF_X4 U8259 ( .I(\SB2_3_9/buf_output[3] ), .Z(\RI5[3][147] ) );
  NAND2_X2 U1940 ( .A1(\SB1_0_23/i0_0 ), .A2(\SB1_0_23/i3[0] ), .ZN(
        \SB1_0_23/Component_Function_5/NAND4_in[0] ) );
  INV_X2 U1436 ( .I(n292), .ZN(\SB1_0_16/i1[9] ) );
  BUF_X4 \MC_ARK_ARC_1_1/BUF_153  ( .I(\SB2_1_8/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[153] ) );
  INV_X8 \SB2_0_14/INV_3  ( .I(\RI3[0][105] ), .ZN(\SB2_0_14/i0[8] ) );
  INV_X4 U850 ( .I(n722), .ZN(\SB2_2_15/i0_4 ) );
  BUF_X4 U1426 ( .I(\RI3[0][23] ), .Z(\SB2_0_28/i0_3 ) );
  CLKBUF_X4 \SB2_2_15/BUF_1  ( .I(\SB1_2_19/buf_output[1] ), .Z(
        \SB2_2_15/i0[6] ) );
  CLKBUF_X4 \SB1_0_9/BUF_3  ( .I(n385), .Z(\SB1_0_9/i0[10] ) );
  NAND3_X2 U1168 ( .A1(\SB1_3_10/i0_3 ), .A2(\SB1_3_10/i1[9] ), .A3(
        \SB1_3_10/i0[6] ), .ZN(\SB1_3_10/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 \SB2_0_14/Component_Function_3/N1  ( .A1(\SB2_0_14/i1[9] ), .A2(
        \SB2_0_14/i0_3 ), .A3(\SB2_0_14/i0[6] ), .ZN(
        \SB2_0_14/Component_Function_3/NAND4_in[0] ) );
  NAND2_X2 \SB1_2_5/Component_Function_5/N1  ( .A1(\SB1_2_5/i0_0 ), .A2(
        \SB1_2_5/i3[0] ), .ZN(\SB1_2_5/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB1_2_12/Component_Function_2/N3  ( .A1(\SB1_2_12/i0_3 ), .A2(
        \SB1_2_12/i0[8] ), .A3(\SB1_2_12/i0[9] ), .ZN(
        \SB1_2_12/Component_Function_2/NAND4_in[2] ) );
  BUF_X2 U90 ( .I(Key[134]), .Z(n114) );
  NAND3_X2 U6494 ( .A1(\SB2_1_5/i0[9] ), .A2(\SB1_1_6/buf_output[4] ), .A3(
        \SB2_1_5/i0[6] ), .ZN(\SB2_1_5/Component_Function_5/NAND4_in[3] ) );
  INV_X2 U4815 ( .I(\MC_ARK_ARC_1_2/buf_output[21] ), .ZN(\SB1_3_28/i0[8] ) );
  NAND3_X2 U1711 ( .A1(\SB2_0_15/i0_3 ), .A2(\SB2_0_15/i0[10] ), .A3(
        \SB2_0_15/i0[6] ), .ZN(\SB2_0_15/Component_Function_2/NAND4_in[1] ) );
  INV_X2 U1621 ( .I(\SB1_3_7/buf_output[5] ), .ZN(\SB2_3_7/i1_5 ) );
  BUF_X4 U1620 ( .I(\SB1_3_7/buf_output[5] ), .Z(\SB2_3_7/i0_3 ) );
  NAND3_X2 U2947 ( .A1(\SB2_3_15/i0_3 ), .A2(\SB2_3_15/i0[6] ), .A3(
        \SB2_3_15/i1[9] ), .ZN(\SB2_3_15/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 \SB2_0_8/BUF_5  ( .I(\SB1_0_8/buf_output[5] ), .Z(\SB2_0_8/i0_3 ) );
  NAND2_X2 \SB2_1_14/Component_Function_5/N1  ( .A1(\SB2_1_14/i0_0 ), .A2(
        \SB2_1_14/i3[0] ), .ZN(\SB2_1_14/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U5522 ( .A1(\SB2_1_24/i0_3 ), .A2(\SB2_1_24/i0_0 ), .A3(
        \SB2_1_24/i0_4 ), .ZN(\SB2_1_24/Component_Function_3/NAND4_in[1] ) );
  INV_X2 \SB2_0_21/INV_3  ( .I(\RI3[0][63] ), .ZN(\SB2_0_21/i0[8] ) );
  BUF_X4 U8176 ( .I(\SB2_2_5/buf_output[1] ), .Z(\RI5[2][181] ) );
  NAND3_X2 U881 ( .A1(\SB1_2_19/i0[10] ), .A2(\SB1_2_19/i0_0 ), .A3(
        \SB1_2_19/i0[6] ), .ZN(\SB1_2_19/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 \SB1_1_9/Component_Function_3/N2  ( .A1(\SB1_1_9/i0_0 ), .A2(
        \SB1_1_9/i0_3 ), .A3(\SB1_1_9/i0_4 ), .ZN(
        \SB1_1_9/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U965 ( .A1(\SB2_1_12/i0[10] ), .A2(\SB2_1_12/i0_3 ), .A3(
        \SB2_1_12/i0[9] ), .ZN(n782) );
  NAND3_X2 U7782 ( .A1(\SB1_2_13/i0_4 ), .A2(\SB1_2_13/i1_5 ), .A3(
        \SB1_2_13/i0_0 ), .ZN(n2795) );
  BUF_X4 \SB2_0_8/BUF_0_0  ( .I(\SB2_0_8/buf_output[0] ), .Z(\RI5[0][168] ) );
  NAND4_X2 U5243 ( .A1(\SB2_0_8/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_0_8/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_0_8/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_8/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_0_8/buf_output[0] ) );
  INV_X2 U4913 ( .I(\MC_ARK_ARC_1_0/buf_output[83] ), .ZN(\SB1_1_18/i1_5 ) );
  BUF_X4 U1638 ( .I(\MC_ARK_ARC_1_0/buf_output[89] ), .Z(\SB1_1_17/i0_3 ) );
  NAND3_X1 \SB1_3_9/Component_Function_2/N4  ( .A1(\SB1_3_9/i1_5 ), .A2(
        \SB1_3_9/i0_0 ), .A3(\SB1_3_9/i0_4 ), .ZN(
        \SB1_3_9/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 U1072 ( .A1(\SB2_0_15/i0[7] ), .A2(\SB2_0_15/i0[8] ), .A3(
        \SB2_0_15/i0[6] ), .ZN(n2329) );
  BUF_X4 \SB2_2_0/BUF_5  ( .I(\SB1_2_0/buf_output[5] ), .Z(\SB2_2_0/i0_3 ) );
  NAND3_X2 \SB2_0_15/Component_Function_0/N4  ( .A1(\SB2_0_15/i0[7] ), .A2(
        \SB2_0_15/i0_3 ), .A3(\SB2_0_15/i0_0 ), .ZN(
        \SB2_0_15/Component_Function_0/NAND4_in[3] ) );
  NAND3_X2 U1068 ( .A1(\SB2_0_28/i0_3 ), .A2(\SB2_0_28/i1[9] ), .A3(
        \RI3[0][22] ), .ZN(n2681) );
  INV_X2 U1601 ( .I(\SB1_1_29/buf_output[1] ), .ZN(\SB2_1_25/i1_7 ) );
  INV_X4 \SB2_1_25/INV_4  ( .I(n1579), .ZN(\SB2_1_25/i0[7] ) );
  BUF_X4 U1275 ( .I(\SB2_3_20/buf_output[2] ), .Z(\RI5[3][86] ) );
  CLKBUF_X4 \SB2_2_4/BUF_1  ( .I(\SB1_2_8/buf_output[1] ), .Z(\SB2_2_4/i0[6] )
         );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_156  ( .I(\SB2_0_10/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[156] ) );
  CLKBUF_X4 U1602 ( .I(\SB1_1_29/buf_output[1] ), .Z(\SB2_1_25/i0[6] ) );
  BUF_X4 U1919 ( .I(\SB2_0_11/i0[9] ), .Z(n1911) );
  INV_X2 \SB3_3/INV_3  ( .I(n1385), .ZN(\SB3_3/i0[8] ) );
  NAND3_X2 \SB2_2_2/Component_Function_3/N3  ( .A1(\SB2_2_2/i1[9] ), .A2(
        \SB2_2_2/i1_7 ), .A3(\SB2_2_2/i0[10] ), .ZN(
        \SB2_2_2/Component_Function_3/NAND4_in[2] ) );
  BUF_X4 U8172 ( .I(\SB2_2_7/buf_output[2] ), .Z(\RI5[2][164] ) );
  BUF_X2 U113 ( .I(Key[143]), .Z(n160) );
  BUF_X2 U47 ( .I(Key[26]), .Z(n162) );
  NAND3_X2 \SB1_0_5/Component_Function_5/N4  ( .A1(\SB1_0_5/i0[9] ), .A2(
        \SB1_0_5/i0[6] ), .A3(\SB1_0_5/i0_4 ), .ZN(
        \SB1_0_5/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 U3603 ( .A1(\SB2_3_8/i0_0 ), .A2(\SB1_3_9/buf_output[4] ), .A3(
        \SB2_3_8/i1_5 ), .ZN(n1049) );
  NAND3_X2 \SB1_0_5/Component_Function_2/N3  ( .A1(\SB1_0_5/i0_3 ), .A2(
        \SB1_0_5/i0[8] ), .A3(\SB1_0_5/i0[9] ), .ZN(
        \SB1_0_5/Component_Function_2/NAND4_in[2] ) );
  INV_X2 \SB1_1_3/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[169] ), .ZN(
        \SB1_1_3/i1_7 ) );
  INV_X4 U6216 ( .I(n1976), .ZN(\SB2_0_11/i0_4 ) );
  NAND3_X2 U4765 ( .A1(\SB2_0_26/i0[10] ), .A2(\SB2_0_26/i0_3 ), .A3(
        \SB2_0_26/i0[9] ), .ZN(n1447) );
  NAND4_X2 \SB2_0_5/Component_Function_1/N5  ( .A1(
        \SB2_0_5/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_5/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_5/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_0_5/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_0_5/buf_output[1] ) );
  NAND4_X2 \SB2_0_18/Component_Function_1/N5  ( .A1(
        \SB2_0_18/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_18/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_18/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_0_18/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_0_18/buf_output[1] ) );
  BUF_X4 U4517 ( .I(\SB1_2_24/buf_output[5] ), .Z(\SB2_2_24/i0_3 ) );
  NAND3_X2 U4532 ( .A1(\SB2_2_30/i0_0 ), .A2(\SB2_2_30/i0[6] ), .A3(
        \SB2_2_30/i0[10] ), .ZN(\SB2_2_30/Component_Function_5/NAND4_in[1] )
         );
  CLKBUF_X2 U194 ( .I(Key[156]), .Z(n133) );
  NAND3_X2 \SB2_2_31/Component_Function_5/N4  ( .A1(\SB2_2_31/i0[9] ), .A2(
        \SB2_2_31/i0[6] ), .A3(n569), .ZN(
        \SB2_2_31/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 U826 ( .A1(\SB2_2_9/i0[10] ), .A2(\SB2_2_9/i1[9] ), .A3(
        \SB2_2_9/i1_7 ), .ZN(\SB2_2_9/Component_Function_3/NAND4_in[2] ) );
  CLKBUF_X4 U4781 ( .I(\SB2_2_28/buf_output[0] ), .Z(\RI5[2][48] ) );
  BUF_X4 U8121 ( .I(\SB2_1_5/buf_output[1] ), .Z(\RI5[1][181] ) );
  NAND3_X2 \SB2_0_24/Component_Function_5/N4  ( .A1(\SB2_0_24/i0[9] ), .A2(
        \RI3[0][43] ), .A3(\RI3[0][46] ), .ZN(
        \SB2_0_24/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 \SB1_3_22/Component_Function_2/N3  ( .A1(\SB1_3_22/i0_3 ), .A2(
        \SB1_3_22/i0[8] ), .A3(\SB1_3_22/i0[9] ), .ZN(
        \SB1_3_22/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U2709 ( .A1(\SB2_0_23/i0_3 ), .A2(\SB2_0_23/i0[9] ), .A3(
        \SB2_0_23/i0[8] ), .ZN(n731) );
  NAND3_X2 U703 ( .A1(n4763), .A2(\SB2_3_17/i0[6] ), .A3(\SB2_3_17/i0[9] ), 
        .ZN(\SB2_3_17/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 U7478 ( .A1(\SB2_0_3/i0_3 ), .A2(\SB2_0_3/i0[9] ), .A3(
        \SB2_0_3/i0[10] ), .ZN(\SB2_0_3/Component_Function_4/NAND4_in[2] ) );
  BUF_X4 \SB1_3_31/BUF_3  ( .I(\MC_ARK_ARC_1_2/buf_output[3] ), .Z(
        \SB1_3_31/i0[10] ) );
  NAND3_X2 \SB2_1_19/Component_Function_2/N3  ( .A1(\SB2_1_19/i0_3 ), .A2(
        \SB2_1_19/i0[8] ), .A3(\SB2_1_19/i0[9] ), .ZN(
        \SB2_1_19/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 \SB1_1_31/Component_Function_5/N4  ( .A1(\SB1_1_31/i0[9] ), .A2(
        \SB1_1_31/i0[6] ), .A3(\SB1_1_31/i0_4 ), .ZN(
        \SB1_1_31/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 \SB1_1_16/Component_Function_3/N3  ( .A1(\SB1_1_16/i1[9] ), .A2(
        \SB1_1_16/i1_7 ), .A3(\SB1_1_16/i0[10] ), .ZN(
        \SB1_1_16/Component_Function_3/NAND4_in[2] ) );
  INV_X2 U1479 ( .I(\MC_ARK_ARC_1_0/buf_output[85] ), .ZN(\SB1_1_17/i1_7 ) );
  NAND2_X2 \SB1_1_2/Component_Function_5/N1  ( .A1(\SB1_1_2/i0_0 ), .A2(
        \SB1_1_2/i3[0] ), .ZN(\SB1_1_2/Component_Function_5/NAND4_in[0] ) );
  INV_X2 \SB2_0_18/INV_5  ( .I(\SB1_0_18/buf_output[5] ), .ZN(\SB2_0_18/i1_5 )
         );
  CLKBUF_X4 \SB1_1_12/BUF_3  ( .I(\MC_ARK_ARC_1_0/buf_output[117] ), .Z(
        \SB1_1_12/i0[10] ) );
  BUF_X2 U42 ( .I(Key[82]), .Z(n117) );
  NAND3_X1 \SB2_0_6/Component_Function_5/N4  ( .A1(\SB2_0_6/i0[9] ), .A2(
        \SB2_0_6/i0[6] ), .A3(\RI3[0][154] ), .ZN(
        \SB2_0_6/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 \SB1_1_0/Component_Function_5/N1  ( .A1(\SB1_1_0/i0_0 ), .A2(
        \SB1_1_0/i3[0] ), .ZN(\SB1_1_0/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 U4855 ( .I(\SB1_0_18/buf_output[5] ), .Z(\SB2_0_18/i0_3 ) );
  INV_X4 U993 ( .I(n2828), .ZN(\SB2_1_30/i0_4 ) );
  NAND4_X2 U3392 ( .A1(\SB1_0_5/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_0_5/Component_Function_4/NAND4_in[1] ), .A3(n2478), .A4(
        \SB1_0_5/Component_Function_4/NAND4_in[0] ), .ZN(
        \SB1_0_5/buf_output[4] ) );
  BUF_X4 \SB2_0_31/BUF_4_0  ( .I(\SB2_0_31/buf_output[4] ), .Z(\RI5[0][10] )
         );
  INV_X2 \SB4_18/INV_1  ( .I(\SB3_22/buf_output[1] ), .ZN(\SB4_18/i1_7 ) );
  BUF_X4 U1903 ( .I(\SB1_1_18/buf_output[5] ), .Z(\SB2_1_18/i0_3 ) );
  NAND3_X2 \SB2_2_4/Component_Function_2/N1  ( .A1(\SB2_2_4/i1_5 ), .A2(
        \SB2_2_4/i0[10] ), .A3(\SB2_2_4/i1[9] ), .ZN(
        \SB2_2_4/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U870 ( .A1(\SB1_2_24/i0[10] ), .A2(\SB1_2_24/i0_0 ), .A3(
        \SB1_2_24/i0[6] ), .ZN(n887) );
  BUF_X4 \SB2_3_30/BUF_5  ( .I(\SB1_3_30/buf_output[5] ), .Z(\SB2_3_30/i0_3 )
         );
  NAND3_X2 \SB2_3_29/Component_Function_2/N3  ( .A1(\SB2_3_29/i0_3 ), .A2(
        \SB2_3_29/i0[8] ), .A3(\SB2_3_29/i0[9] ), .ZN(
        \SB2_3_29/Component_Function_2/NAND4_in[2] ) );
  INV_X2 U1282 ( .I(\MC_ARK_ARC_1_3/buf_output[164] ), .ZN(\SB3_4/i1[9] ) );
  CLKBUF_X4 \SB2_3_30/BUF_4  ( .I(\SB1_3_31/buf_output[4] ), .Z(
        \SB2_3_30/i0_4 ) );
  NAND3_X2 \SB1_2_0/Component_Function_3/N3  ( .A1(\SB1_2_0/i1[9] ), .A2(
        \SB1_2_0/i1_7 ), .A3(\SB1_2_0/i0[10] ), .ZN(
        \SB1_2_0/Component_Function_3/NAND4_in[2] ) );
  BUF_X4 U3900 ( .I(\SB2_1_7/buf_output[0] ), .Z(\RI5[1][174] ) );
  BUF_X4 U8180 ( .I(\SB2_2_12/buf_output[0] ), .Z(\RI5[2][144] ) );
  NAND3_X2 \SB1_1_26/Component_Function_5/N4  ( .A1(\SB1_1_26/i0[9] ), .A2(
        \SB1_1_26/i0[6] ), .A3(\SB1_1_26/i0_4 ), .ZN(
        \SB1_1_26/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 \SB2_1_18/Component_Function_2/N1  ( .A1(\SB2_1_18/i1_5 ), .A2(
        \SB2_1_18/i0[10] ), .A3(\SB2_1_18/i1[9] ), .ZN(
        \SB2_1_18/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB2_0_18/Component_Function_4/N3  ( .A1(\SB2_0_18/i0[9] ), .A2(
        \SB2_0_18/i0[10] ), .A3(\SB2_0_18/i0_3 ), .ZN(
        \SB2_0_18/Component_Function_4/NAND4_in[2] ) );
  INV_X2 \SB1_1_23/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[53] ), .ZN(
        \SB1_1_23/i1_5 ) );
  CLKBUF_X2 U130 ( .I(Key[28]), .Z(n235) );
  NAND3_X2 \SB2_1_19/Component_Function_2/N2  ( .A1(\SB2_1_19/i0_3 ), .A2(
        \SB2_1_19/i0[10] ), .A3(\SB2_1_19/i0[6] ), .ZN(
        \SB2_1_19/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 \SB2_2_8/Component_Function_5/N2  ( .A1(\SB2_2_8/i0_0 ), .A2(
        \SB2_2_8/i0[6] ), .A3(\SB2_2_8/i0[10] ), .ZN(
        \SB2_2_8/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 \SB1_1_16/BUF_3  ( .I(\MC_ARK_ARC_1_0/buf_output[93] ), .Z(
        \SB1_1_16/i0[10] ) );
  NAND3_X2 U1717 ( .A1(\SB1_3_4/i1[9] ), .A2(\SB1_3_4/i0_4 ), .A3(
        \SB1_3_4/i0_3 ), .ZN(\SB1_3_4/Component_Function_5/NAND4_in[2] ) );
  BUF_X4 \SB2_0_15/BUF_3_0  ( .I(\SB2_0_15/buf_output[3] ), .Z(\RI5[0][111] )
         );
  NAND4_X2 \SB2_0_0/Component_Function_1/N5  ( .A1(
        \SB2_0_0/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_0/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_0/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_0_0/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_0_0/buf_output[1] ) );
  NAND2_X2 \SB1_0_27/Component_Function_5/N1  ( .A1(\SB1_0_27/i0_0 ), .A2(
        \SB1_0_27/i3[0] ), .ZN(\SB1_0_27/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 \SB2_3_15/BUF_3  ( .I(\SB1_3_17/buf_output[3] ), .Z(\SB2_3_15/i0[10] ) );
  BUF_X4 U4967 ( .I(n3659), .Z(\SB1_1_7/i0[10] ) );
  NAND3_X2 U4510 ( .A1(\SB3_7/i0_0 ), .A2(\SB3_7/i0_3 ), .A3(\SB3_7/i0_4 ), 
        .ZN(\SB3_7/Component_Function_3/NAND4_in[1] ) );
  BUF_X4 U8159 ( .I(\SB2_2_1/buf_output[3] ), .Z(\RI5[2][3] ) );
  BUF_X4 \SB1_3_23/BUF_3  ( .I(\MC_ARK_ARC_1_2/buf_output[51] ), .Z(
        \SB1_3_23/i0[10] ) );
  BUF_X4 U8100 ( .I(\SB2_1_20/buf_output[1] ), .Z(\RI5[1][91] ) );
  NAND3_X2 \SB1_2_10/Component_Function_5/N2  ( .A1(\SB1_2_10/i0_0 ), .A2(
        \SB1_2_10/i0[6] ), .A3(\SB1_2_10/i0[10] ), .ZN(
        \SB1_2_10/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 \SB2_2_0/Component_Function_1/N2  ( .A1(\SB2_2_0/i0_3 ), .A2(
        \SB2_2_0/i1_7 ), .A3(\SB2_2_0/i0[8] ), .ZN(
        \SB2_2_0/Component_Function_1/NAND4_in[1] ) );
  NAND3_X2 \SB2_0_21/Component_Function_2/N4  ( .A1(\SB2_0_21/i1_5 ), .A2(
        \SB2_0_21/i0_0 ), .A3(\SB2_0_21/i0_4 ), .ZN(
        \SB2_0_21/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 \SB2_3_5/Component_Function_2/N2  ( .A1(\SB2_3_5/i0_3 ), .A2(
        \SB2_3_5/i0[10] ), .A3(\SB2_3_5/i0[6] ), .ZN(
        \SB2_3_5/Component_Function_2/NAND4_in[1] ) );
  CLKBUF_X4 \SB1_0_25/BUF_1  ( .I(n264), .Z(\SB1_0_25/i0[6] ) );
  BUF_X4 \SB2_2_2/BUF_0  ( .I(\SB1_2_7/buf_output[0] ), .Z(\SB2_2_2/i0[9] ) );
  CLKBUF_X4 U4694 ( .I(\SB1_2_19/buf_output[4] ), .Z(\SB2_2_18/i0_4 ) );
  NAND3_X2 \SB1_2_1/Component_Function_0/N4  ( .A1(\SB1_2_1/i0[7] ), .A2(
        \SB1_2_1/i0_3 ), .A3(\SB1_2_1/i0_0 ), .ZN(
        \SB1_2_1/Component_Function_0/NAND4_in[3] ) );
  NAND3_X2 U5355 ( .A1(\SB2_1_29/i0[6] ), .A2(\SB2_1_29/i0_3 ), .A3(
        \SB2_1_29/i0[10] ), .ZN(\SB2_1_29/Component_Function_2/NAND4_in[1] )
         );
  BUF_X4 U8269 ( .I(\SB2_3_13/buf_output[4] ), .Z(\RI5[3][118] ) );
  BUF_X2 U84 ( .I(Key[30]), .Z(n152) );
  CLKBUF_X4 U1962 ( .I(\RI3[0][44] ), .Z(\SB2_0_24/i0_0 ) );
  NAND3_X2 U933 ( .A1(\SB1_2_12/i0_3 ), .A2(\SB1_2_12/i0_4 ), .A3(
        \SB1_2_12/i1[9] ), .ZN(\SB1_2_12/Component_Function_5/NAND4_in[2] ) );
  BUF_X2 U74 ( .I(Key[68]), .Z(n125) );
  NAND3_X2 U5312 ( .A1(\SB2_2_0/i0[6] ), .A2(\SB2_2_0/i0_3 ), .A3(
        \SB2_2_0/i0[10] ), .ZN(\SB2_2_0/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 \SB2_0_4/BUF_0_0  ( .I(\SB2_0_4/buf_output[0] ), .Z(\RI5[0][0] ) );
  NAND3_X2 U2166 ( .A1(\SB2_3_13/i0[10] ), .A2(\SB2_3_13/i1_7 ), .A3(
        \SB2_3_13/i1[9] ), .ZN(\SB2_3_13/Component_Function_3/NAND4_in[2] ) );
  NAND2_X2 \SB3_21/Component_Function_1/N1  ( .A1(\SB3_21/i0_3 ), .A2(
        \SB3_21/i1[9] ), .ZN(\SB3_21/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 \SB2_0_24/Component_Function_3/N1  ( .A1(\SB2_0_24/i1[9] ), .A2(
        \SB2_0_24/i0_3 ), .A3(\RI3[0][43] ), .ZN(
        \SB2_0_24/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 U1932 ( .I(n255), .Z(\SB1_0_28/i0[6] ) );
  BUF_X4 \SB1_2_28/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[22] ), .Z(
        \SB1_2_28/i0_4 ) );
  BUF_X4 U2114 ( .I(\MC_ARK_ARC_1_2/buf_output[116] ), .Z(\SB1_3_12/i0_0 ) );
  NAND3_X1 \SB1_3_31/Component_Function_0/N2  ( .A1(\SB1_3_31/i0[8] ), .A2(
        \SB1_3_31/i0[7] ), .A3(\SB1_3_31/i0[6] ), .ZN(
        \SB1_3_31/Component_Function_0/NAND4_in[1] ) );
  CLKBUF_X4 \SB2_2_8/BUF_2  ( .I(\SB1_2_11/buf_output[2] ), .Z(\SB2_2_8/i0_0 )
         );
  NAND3_X2 U1089 ( .A1(\SB2_0_25/i0_0 ), .A2(\RI3[0][40] ), .A3(
        \SB2_0_25/i1_5 ), .ZN(n1550) );
  NAND4_X2 U5490 ( .A1(\SB2_2_30/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_30/Component_Function_3/NAND4_in[3] ), .A3(
        \SB2_2_30/Component_Function_3/NAND4_in[1] ), .A4(n1647), .ZN(
        \SB2_2_30/buf_output[3] ) );
  INV_X2 U1469 ( .I(\MC_ARK_ARC_1_2/buf_output[49] ), .ZN(\SB1_3_23/i1_7 ) );
  NAND3_X2 U995 ( .A1(\SB1_1_15/i0_3 ), .A2(\SB1_1_15/i0_4 ), .A3(
        \SB1_1_15/i1[9] ), .ZN(n1696) );
  NAND3_X2 \SB1_0_16/Component_Function_2/N1  ( .A1(\SB1_0_16/i1_5 ), .A2(
        \SB1_0_16/i0[10] ), .A3(\SB1_0_16/i1[9] ), .ZN(
        \SB1_0_16/Component_Function_2/NAND4_in[0] ) );
  INV_X2 U1481 ( .I(\MC_ARK_ARC_1_3/buf_output[122] ), .ZN(\SB3_11/i1[9] ) );
  NAND3_X2 \SB2_3_3/Component_Function_2/N2  ( .A1(\SB2_3_3/i0_3 ), .A2(
        \SB2_3_3/i0[10] ), .A3(\SB2_3_3/i0[6] ), .ZN(
        \SB2_3_3/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U5712 ( .A1(\SB2_2_14/i0_3 ), .A2(n5932), .A3(\SB2_2_14/i1[9] ), 
        .ZN(\SB2_2_14/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 \SB1_0_31/Component_Function_4/N3  ( .A1(\SB1_0_31/i0[9] ), .A2(
        \SB1_0_31/i0[10] ), .A3(\SB1_0_31/i0_3 ), .ZN(
        \SB1_0_31/Component_Function_4/NAND4_in[2] ) );
  BUF_X4 \SB2_0_7/BUF_0_0  ( .I(\SB2_0_7/buf_output[0] ), .Z(\RI5[0][174] ) );
  INV_X2 \SB1_2_3/INV_1  ( .I(\MC_ARK_ARC_1_1/buf_output[169] ), .ZN(
        \SB1_2_3/i1_7 ) );
  BUF_X2 \SB1_1_25/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[37] ), .Z(
        \SB1_1_25/i0[6] ) );
  BUF_X4 \SB1_0_19/BUF_4_0  ( .I(\SB1_0_19/buf_output[4] ), .Z(\RI3[0][82] )
         );
  INV_X2 \SB1_0_31/INV_3  ( .I(n341), .ZN(\SB1_0_31/i0[8] ) );
  INV_X2 \SB1_1_21/INV_0  ( .I(n3131), .ZN(\SB1_1_21/i3[0] ) );
  NAND3_X2 \SB2_1_3/Component_Function_2/N3  ( .A1(\SB2_1_3/i0_3 ), .A2(
        \SB2_1_3/i0[8] ), .A3(\SB2_1_3/i0[9] ), .ZN(
        \SB2_1_3/Component_Function_2/NAND4_in[2] ) );
  BUF_X2 U58 ( .I(Key[65]), .Z(n156) );
  NAND3_X2 \SB2_0_17/Component_Function_3/N4  ( .A1(\SB2_0_17/i1_5 ), .A2(
        \SB2_0_17/i0[8] ), .A3(\SB2_0_17/i3[0] ), .ZN(
        \SB2_0_17/Component_Function_3/NAND4_in[3] ) );
  CLKBUF_X4 U1549 ( .I(\SB1_1_28/buf_output[1] ), .Z(\SB2_1_24/i0[6] ) );
  BUF_X4 U8171 ( .I(\SB2_2_7/buf_output[1] ), .Z(\RI5[2][169] ) );
  NAND3_X2 \SB1_2_17/Component_Function_5/N3  ( .A1(\SB1_2_17/i1[9] ), .A2(
        \SB1_2_17/i0_4 ), .A3(\SB1_2_17/i0_3 ), .ZN(
        \SB1_2_17/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 \SB2_0_4/Component_Function_3/N4  ( .A1(\SB2_0_4/i1_5 ), .A2(
        \SB2_0_4/i0[8] ), .A3(\SB2_0_4/i3[0] ), .ZN(
        \SB2_0_4/Component_Function_3/NAND4_in[3] ) );
  BUF_X4 U8112 ( .I(\SB2_1_27/buf_output[2] ), .Z(\RI5[1][44] ) );
  NAND3_X2 \SB2_3_23/Component_Function_3/N3  ( .A1(\SB2_3_23/i1[9] ), .A2(
        \SB2_3_23/i1_7 ), .A3(\SB2_3_23/i0[10] ), .ZN(
        \SB2_3_23/Component_Function_3/NAND4_in[2] ) );
  BUF_X4 U1841 ( .I(\SB1_3_3/buf_output[5] ), .Z(\SB2_3_3/i0_3 ) );
  INV_X2 U1596 ( .I(\RI1[3][59] ), .ZN(\SB1_3_22/i1_5 ) );
  BUF_X4 U1595 ( .I(\RI1[3][59] ), .Z(\SB1_3_22/i0_3 ) );
  NAND3_X2 U1113 ( .A1(\SB1_0_13/i0[10] ), .A2(\SB1_0_13/i0_0 ), .A3(
        \SB1_0_13/i0[6] ), .ZN(\SB1_0_13/Component_Function_5/NAND4_in[1] ) );
  INV_X2 \SB1_0_6/INV_1  ( .I(n321), .ZN(\SB1_0_6/i1_7 ) );
  BUF_X2 U51 ( .I(Key[152]), .Z(n103) );
  NAND3_X2 \SB2_0_25/Component_Function_2/N3  ( .A1(\SB2_0_25/i0_3 ), .A2(
        \SB2_0_25/i0[8] ), .A3(\SB2_0_25/i0[9] ), .ZN(
        \SB2_0_25/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U4434 ( .A1(\SB3_11/i0[6] ), .A2(\SB3_11/i0[9] ), .A3(\SB3_11/i0_4 ), .ZN(n1490) );
  BUF_X4 U4688 ( .I(\SB1_1_6/buf_output[5] ), .Z(\SB2_1_6/i0_3 ) );
  NAND3_X1 \SB1_0_13/Component_Function_3/N3  ( .A1(\SB1_0_13/i1[9] ), .A2(
        \SB1_0_13/i1_7 ), .A3(\SB1_0_13/i0[10] ), .ZN(
        \SB1_0_13/Component_Function_3/NAND4_in[2] ) );
  INV_X2 U6220 ( .I(n1977), .ZN(\RI1[1][71] ) );
  NAND2_X1 U7270 ( .A1(\SB1_0_2/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_0_2/Component_Function_4/NAND4_in[3] ), .ZN(n2483) );
  BUF_X4 U1170 ( .I(\MC_ARK_ARC_1_2/buf_output[154] ), .Z(\SB1_3_6/i0_4 ) );
  CLKBUF_X2 U134 ( .I(Key[162]), .Z(n143) );
  CLKBUF_X2 U173 ( .I(Key[18]), .Z(n16) );
  CLKBUF_X4 \SB1_0_13/BUF_3  ( .I(n377), .Z(\SB1_0_13/i0[10] ) );
  INV_X1 U333 ( .I(n118), .ZN(n457) );
  CLKBUF_X4 \SB1_0_30/BUF_4  ( .I(n344), .Z(\SB1_0_30/i0_4 ) );
  CLKBUF_X4 U4940 ( .I(n276), .Z(\SB1_0_21/i0[6] ) );
  CLKBUF_X4 U1635 ( .I(n383), .Z(\SB1_0_10/i0[10] ) );
  CLKBUF_X4 \SB1_0_3/BUF_4  ( .I(n398), .Z(\SB1_0_3/i0_4 ) );
  INV_X1 U335 ( .I(n21), .ZN(n472) );
  CLKBUF_X4 \SB1_0_2/BUF_1  ( .I(n333), .Z(\SB1_0_2/i0[6] ) );
  INV_X1 U346 ( .I(n13), .ZN(n540) );
  INV_X1 U352 ( .I(n20), .ZN(n467) );
  CLKBUF_X4 \SB1_0_29/BUF_3  ( .I(n345), .Z(\SB1_0_29/i0[10] ) );
  CLKBUF_X4 \SB1_0_28/BUF_3  ( .I(n347), .Z(\SB1_0_28/i0[10] ) );
  CLKBUF_X4 \SB1_0_26/BUF_2  ( .I(n262), .Z(\SB1_0_26/i0_0 ) );
  CLKBUF_X4 \SB1_0_26/BUF_4  ( .I(n352), .Z(\SB1_0_26/i0_4 ) );
  CLKBUF_X4 \SB1_0_28/BUF_0  ( .I(n254), .Z(\SB1_0_28/i0[9] ) );
  CLKBUF_X4 \SB1_0_6/BUF_3  ( .I(n391), .Z(\SB1_0_6/i0[10] ) );
  INV_X1 U359 ( .I(n34), .ZN(n485) );
  INV_X1 U9 ( .I(n92), .ZN(n511) );
  CLKBUF_X4 \SB1_0_1/BUF_1  ( .I(n336), .Z(\SB1_0_1/i0[6] ) );
  CLKBUF_X4 U1463 ( .I(n401), .Z(\SB1_0_1/i0[10] ) );
  CLKBUF_X4 \SB1_0_11/BUF_3  ( .I(n381), .Z(\SB1_0_11/i0[10] ) );
  CLKBUF_X4 \SB1_0_5/BUF_2  ( .I(n325), .Z(\SB1_0_5/i0_0 ) );
  CLKBUF_X4 U1966 ( .I(\SB1_0_30/buf_output[4] ), .Z(\SB2_0_29/i0_4 ) );
  CLKBUF_X4 U1712 ( .I(\RI3[0][99] ), .Z(\SB2_0_15/i0[10] ) );
  CLKBUF_X4 \SB2_0_10/BUF_1  ( .I(\RI3[0][127] ), .Z(\SB2_0_10/i0[6] ) );
  CLKBUF_X4 \SB2_0_3/BUF_3  ( .I(\SB1_0_5/buf_output[3] ), .Z(\SB2_0_3/i0[10] ) );
  BUF_X2 \SB2_0_8/BUF_0  ( .I(\SB1_0_13/buf_output[0] ), .Z(\SB2_0_8/i0[9] )
         );
  CLKBUF_X4 \SB2_0_26/BUF_3  ( .I(\RI3[0][33] ), .Z(\SB2_0_26/i0[10] ) );
  CLKBUF_X4 \SB2_0_19/BUF_1  ( .I(\SB1_0_23/buf_output[1] ), .Z(
        \SB2_0_19/i0[6] ) );
  BUF_X4 \SB2_0_18/BUF_1_0  ( .I(\SB2_0_18/buf_output[1] ), .Z(\RI5[0][103] )
         );
  CLKBUF_X4 U2817 ( .I(\SB2_0_25/buf_output[5] ), .Z(\RI5[0][41] ) );
  BUF_X4 \SB2_0_1/BUF_3_0  ( .I(\SB2_0_1/buf_output[3] ), .Z(\RI5[0][3] ) );
  CLKBUF_X4 \SB2_0_11/BUF_4_0  ( .I(\SB2_0_11/buf_output[4] ), .Z(
        \RI5[0][130] ) );
  CLKBUF_X4 \SB1_1_23/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[49] ), .Z(
        \SB1_1_23/i0[6] ) );
  CLKBUF_X4 \SB1_1_31/BUF_5  ( .I(\MC_ARK_ARC_1_0/buf_output[5] ), .Z(
        \SB1_1_31/i0_3 ) );
  CLKBUF_X4 U2476 ( .I(\MC_ARK_ARC_1_0/buf_output[170] ), .Z(\SB1_1_3/i0_0 )
         );
  CLKBUF_X4 \SB1_1_26/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[34] ), .Z(
        \SB1_1_26/i0_4 ) );
  CLKBUF_X4 U3428 ( .I(\MC_ARK_ARC_1_0/buf_output[3] ), .Z(\SB1_1_31/i0[10] )
         );
  CLKBUF_X4 \SB1_1_27/BUF_3  ( .I(\MC_ARK_ARC_1_0/buf_output[27] ), .Z(
        \SB1_1_27/i0[10] ) );
  CLKBUF_X4 \SB1_1_0/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[187] ), .Z(
        \SB1_1_0/i0[6] ) );
  CLKBUF_X4 \SB1_1_23/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[48] ), .Z(
        \SB1_1_23/i0[9] ) );
  CLKBUF_X4 \SB1_1_20/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[66] ), .Z(
        \SB1_1_20/i0[9] ) );
  BUF_X2 \SB1_1_6/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[151] ), .Z(
        \SB1_1_6/i0[6] ) );
  CLKBUF_X4 U1058 ( .I(\MC_ARK_ARC_1_0/buf_output[69] ), .Z(\SB1_1_20/i0[10] )
         );
  CLKBUF_X4 \SB1_1_14/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[102] ), .Z(
        \SB1_1_14/i0[9] ) );
  CLKBUF_X4 \SB2_1_1/BUF_2  ( .I(\RI3[1][182] ), .Z(\SB2_1_1/i0_0 ) );
  CLKBUF_X4 \SB2_1_22/BUF_2  ( .I(\SB1_1_25/buf_output[2] ), .Z(
        \SB2_1_22/i0_0 ) );
  CLKBUF_X4 U1695 ( .I(\SB1_1_10/buf_output[3] ), .Z(\SB2_1_8/i0[10] ) );
  CLKBUF_X4 \SB2_1_10/BUF_2  ( .I(\SB1_1_13/buf_output[2] ), .Z(
        \SB2_1_10/i0_0 ) );
  CLKBUF_X4 \SB2_1_24/BUF_4  ( .I(\SB1_1_25/buf_output[4] ), .Z(
        \SB2_1_24/i0_4 ) );
  CLKBUF_X4 \SB2_1_28/BUF_4  ( .I(\SB1_1_29/buf_output[4] ), .Z(
        \SB2_1_28/i0_4 ) );
  CLKBUF_X4 \SB2_1_30/BUF_0  ( .I(\SB1_1_3/buf_output[0] ), .Z(
        \SB2_1_30/i0[9] ) );
  CLKBUF_X4 \SB2_1_2/BUF_3  ( .I(\SB1_1_4/buf_output[3] ), .Z(\SB2_1_2/i0[10] ) );
  CLKBUF_X4 \SB2_1_24/BUF_3  ( .I(\SB1_1_26/buf_output[3] ), .Z(
        \SB2_1_24/i0[10] ) );
  CLKBUF_X4 U4834 ( .I(\SB1_1_6/buf_output[2] ), .Z(\SB2_1_3/i0_0 ) );
  CLKBUF_X4 \SB2_1_2/BUF_2  ( .I(\SB1_1_5/buf_output[2] ), .Z(\SB2_1_2/i0_0 )
         );
  CLKBUF_X4 \SB2_1_23/BUF_3  ( .I(\SB1_1_25/buf_output[3] ), .Z(
        \SB2_1_23/i0[10] ) );
  CLKBUF_X4 U4690 ( .I(\SB1_1_15/buf_output[2] ), .Z(\SB2_1_12/i0_0 ) );
  CLKBUF_X4 \SB2_1_20/BUF_1  ( .I(\SB1_1_24/buf_output[1] ), .Z(
        \SB2_1_20/i0[6] ) );
  CLKBUF_X4 \SB2_1_2/BUF_4  ( .I(\SB1_1_3/buf_output[4] ), .Z(\SB2_1_2/i0_4 )
         );
  CLKBUF_X4 \SB2_1_23/BUF_2  ( .I(\SB1_1_26/buf_output[2] ), .Z(
        \SB2_1_23/i0_0 ) );
  CLKBUF_X4 \SB2_1_21/BUF_1  ( .I(\SB1_1_25/buf_output[1] ), .Z(
        \SB2_1_21/i0[6] ) );
  CLKBUF_X4 \SB2_1_21/BUF_4  ( .I(\SB1_1_22/buf_output[4] ), .Z(
        \SB2_1_21/i0_4 ) );
  CLKBUF_X4 U1893 ( .I(\SB2_1_2/buf_output[0] ), .Z(\RI5[1][12] ) );
  BUF_X4 U6987 ( .I(\SB2_1_18/buf_output[3] ), .Z(\RI5[1][93] ) );
  CLKBUF_X4 U4864 ( .I(\MC_ARK_ARC_1_1/buf_output[105] ), .Z(\SB1_2_14/i0[10] ) );
  CLKBUF_X4 \SB1_2_28/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[18] ), .Z(
        \SB1_2_28/i0[9] ) );
  CLKBUF_X4 U1227 ( .I(\MC_ARK_ARC_1_1/buf_output[74] ), .Z(\SB1_2_19/i0_0 )
         );
  CLKBUF_X4 \SB1_2_17/BUF_2  ( .I(\MC_ARK_ARC_1_1/buf_output[86] ), .Z(
        \SB1_2_17/i0_0 ) );
  CLKBUF_X4 \SB1_2_4/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[166] ), .Z(
        \SB1_2_4/i0_4 ) );
  BUF_X2 \SB1_2_11/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[120] ), .Z(
        \SB1_2_11/i0[9] ) );
  CLKBUF_X4 U1509 ( .I(\MC_ARK_ARC_1_1/buf_output[27] ), .Z(\SB1_2_27/i0[10] )
         );
  CLKBUF_X4 \SB1_2_14/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[102] ), .Z(
        \SB1_2_14/i0[9] ) );
  INV_X4 \SB1_2_26/INV_5  ( .I(\RI1[2][35] ), .ZN(\SB1_2_26/i1_5 ) );
  CLKBUF_X4 \SB1_2_3/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[168] ), .Z(
        \SB1_2_3/i0[9] ) );
  BUF_X2 \SB1_2_14/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[103] ), .Z(
        \SB1_2_14/i0[6] ) );
  CLKBUF_X4 U2060 ( .I(\MC_ARK_ARC_1_1/buf_output[118] ), .Z(\SB1_2_12/i0_4 )
         );
  CLKBUF_X4 \SB2_2_20/BUF_4  ( .I(\SB1_2_21/buf_output[4] ), .Z(
        \SB2_2_20/i0_4 ) );
  CLKBUF_X4 U6434 ( .I(\SB1_2_7/buf_output[4] ), .Z(n2074) );
  CLKBUF_X4 \SB2_2_13/BUF_0  ( .I(\SB1_2_18/buf_output[0] ), .Z(
        \SB2_2_13/i0[9] ) );
  CLKBUF_X4 \SB2_2_2/BUF_4  ( .I(\SB1_2_3/buf_output[4] ), .Z(\SB2_2_2/i0_4 )
         );
  CLKBUF_X4 \SB2_2_23/BUF_2  ( .I(\SB1_2_26/buf_output[2] ), .Z(
        \SB2_2_23/i0_0 ) );
  CLKBUF_X4 \SB2_2_1/BUF_3  ( .I(\SB1_2_3/buf_output[3] ), .Z(\SB2_2_1/i0[10] ) );
  CLKBUF_X4 U1867 ( .I(\SB1_2_12/buf_output[4] ), .Z(\SB2_2_11/i0_4 ) );
  CLKBUF_X4 \SB2_2_19/BUF_0  ( .I(\SB1_2_24/buf_output[0] ), .Z(
        \SB2_2_19/i0[9] ) );
  INV_X2 \SB2_2_5/INV_4  ( .I(\SB2_2_5/i0_4 ), .ZN(\SB2_2_5/i0[7] ) );
  CLKBUF_X4 U4534 ( .I(\SB1_2_2/buf_output[1] ), .Z(\SB2_2_30/i0[6] ) );
  CLKBUF_X4 \SB2_2_14/BUF_2  ( .I(\SB1_2_17/buf_output[2] ), .Z(
        \SB2_2_14/i0_0 ) );
  CLKBUF_X4 U852 ( .I(\SB1_2_31/buf_output[0] ), .Z(\SB2_2_26/i0[9] ) );
  CLKBUF_X4 \SB2_2_9/BUF_0  ( .I(\SB1_2_14/buf_output[0] ), .Z(\SB2_2_9/i0[9] ) );
  BUF_X4 U1858 ( .I(\SB2_2_30/buf_output[1] ), .Z(\RI5[2][31] ) );
  BUF_X4 U8204 ( .I(\SB2_2_30/buf_output[3] ), .Z(\RI5[2][21] ) );
  BUF_X4 U8170 ( .I(\SB2_2_4/buf_output[1] ), .Z(\RI5[2][187] ) );
  CLKBUF_X4 U4912 ( .I(\SB2_2_27/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[34] ) );
  CLKBUF_X4 U7154 ( .I(\SB2_2_20/buf_output[1] ), .Z(\RI5[2][91] ) );
  CLKBUF_X4 U8164 ( .I(\SB2_2_3/buf_output[1] ), .Z(\RI5[2][1] ) );
  CLKBUF_X4 U4601 ( .I(\MC_ARK_ARC_1_2/buf_output[147] ), .Z(\SB1_3_7/i0[10] )
         );
  BUF_X2 \SB1_3_21/BUF_1  ( .I(\MC_ARK_ARC_1_2/buf_output[61] ), .Z(
        \SB1_3_21/i0[6] ) );
  BUF_X4 U4466 ( .I(\MC_ARK_ARC_1_2/buf_output[40] ), .Z(\SB1_3_25/i0_4 ) );
  CLKBUF_X4 \SB1_3_10/BUF_1  ( .I(\MC_ARK_ARC_1_2/buf_output[127] ), .Z(
        \SB1_3_10/i0[6] ) );
  CLKBUF_X4 \SB1_3_14/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[106] ), .Z(
        \SB1_3_14/i0_4 ) );
  CLKBUF_X4 \SB1_3_13/BUF_2  ( .I(\MC_ARK_ARC_1_2/buf_output[110] ), .Z(
        \SB1_3_13/i0_0 ) );
  CLKBUF_X4 \SB1_3_18/BUF_2  ( .I(n5527), .Z(\SB1_3_18/i0_0 ) );
  CLKBUF_X4 \SB1_3_18/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[82] ), .Z(
        \SB1_3_18/i0_4 ) );
  CLKBUF_X4 \SB1_3_14/BUF_2  ( .I(n5506), .Z(\SB1_3_14/i0_0 ) );
  CLKBUF_X4 \SB1_3_4/BUF_3  ( .I(\MC_ARK_ARC_1_2/buf_output[165] ), .Z(
        \SB1_3_4/i0[10] ) );
  CLKBUF_X4 \SB1_3_21/BUF_3  ( .I(\MC_ARK_ARC_1_2/buf_output[63] ), .Z(
        \SB1_3_21/i0[10] ) );
  CLKBUF_X4 U1608 ( .I(\MC_ARK_ARC_1_2/buf_output[54] ), .Z(\SB1_3_22/i0[9] )
         );
  CLKBUF_X4 \SB1_3_26/BUF_3  ( .I(\MC_ARK_ARC_1_2/buf_output[33] ), .Z(
        \SB1_3_26/i0[10] ) );
  CLKBUF_X8 \SB1_3_8/BUF_5  ( .I(\RI1[3][143] ), .Z(\SB1_3_8/i0_3 ) );
  CLKBUF_X4 U1842 ( .I(\SB1_3_11/buf_output[4] ), .Z(\SB2_3_10/i0_4 ) );
  CLKBUF_X4 \SB2_3_1/BUF_4  ( .I(\SB1_3_2/buf_output[4] ), .Z(\SB2_3_1/i0_4 )
         );
  CLKBUF_X4 \SB2_3_22/BUF_4  ( .I(\SB1_3_23/buf_output[4] ), .Z(
        \SB2_3_22/i0_4 ) );
  CLKBUF_X4 \SB2_3_19/BUF_3  ( .I(\SB1_3_21/buf_output[3] ), .Z(
        \SB2_3_19/i0[10] ) );
  CLKBUF_X4 \SB2_3_19/BUF_2  ( .I(\SB1_3_22/buf_output[2] ), .Z(
        \SB2_3_19/i0_0 ) );
  CLKBUF_X4 U2146 ( .I(\SB1_3_20/buf_output[4] ), .Z(\SB2_3_19/i0_4 ) );
  BUF_X4 \SB2_3_5/BUF_5  ( .I(\SB1_3_5/buf_output[5] ), .Z(\SB2_3_5/i0_3 ) );
  CLKBUF_X4 \SB2_3_12/BUF_2  ( .I(\SB1_3_15/buf_output[2] ), .Z(
        \SB2_3_12/i0_0 ) );
  CLKBUF_X4 \SB2_3_16/BUF_4  ( .I(\SB1_3_17/buf_output[4] ), .Z(
        \SB2_3_16/i0_4 ) );
  CLKBUF_X4 \SB2_3_25/BUF_3  ( .I(\SB1_3_27/buf_output[3] ), .Z(
        \SB2_3_25/i0[10] ) );
  BUF_X4 \SB2_3_8/BUF_3  ( .I(\SB1_3_10/buf_output[3] ), .Z(\SB2_3_8/i0[10] )
         );
  CLKBUF_X4 \SB2_3_25/BUF_1  ( .I(\SB1_3_29/buf_output[1] ), .Z(
        \SB2_3_25/i0[6] ) );
  CLKBUF_X4 U1285 ( .I(\MC_ARK_ARC_1_3/buf_output[27] ), .Z(\SB3_27/i0[10] )
         );
  CLKBUF_X4 U1268 ( .I(\MC_ARK_ARC_1_3/buf_output[176] ), .Z(\SB3_2/i0_0 ) );
  CLKBUF_X4 U1536 ( .I(\MC_ARK_ARC_1_3/buf_output[126] ), .Z(\SB3_10/i0[9] )
         );
  CLKBUF_X4 \SB3_31/BUF_4  ( .I(\MC_ARK_ARC_1_3/buf_output[4] ), .Z(
        \SB3_31/i0_4 ) );
  CLKBUF_X4 \SB3_31/BUF_3  ( .I(\MC_ARK_ARC_1_3/buf_output[3] ), .Z(
        \SB3_31/i0[10] ) );
  CLKBUF_X4 \SB3_19/BUF_4  ( .I(\MC_ARK_ARC_1_3/buf_output[76] ), .Z(
        \SB3_19/i0_4 ) );
  BUF_X2 U4844 ( .I(\MC_ARK_ARC_1_3/buf_output[36] ), .Z(\SB3_25/i0[9] ) );
  CLKBUF_X4 \SB3_17/BUF_4  ( .I(\MC_ARK_ARC_1_3/buf_output[88] ), .Z(
        \SB3_17/i0_4 ) );
  CLKBUF_X4 \SB3_20/BUF_1  ( .I(\MC_ARK_ARC_1_3/buf_output[67] ), .Z(
        \SB3_20/i0[6] ) );
  BUF_X2 U1181 ( .I(\MC_ARK_ARC_1_3/buf_output[73] ), .Z(\SB3_19/i0[6] ) );
  CLKBUF_X4 U4575 ( .I(\SB3_15/buf_output[5] ), .Z(\SB4_15/i0_3 ) );
  BUF_X2 \SB4_22/BUF_1  ( .I(\SB3_26/buf_output[1] ), .Z(\SB4_22/i0[6] ) );
  BUF_X2 U4467 ( .I(\SB3_15/buf_output[1] ), .Z(\SB4_11/i0[6] ) );
  BUF_X2 U591 ( .I(\SB3_9/buf_output[3] ), .Z(\SB4_7/i0[10] ) );
  CLKBUF_X4 U1784 ( .I(\SB3_15/buf_output[4] ), .Z(\SB4_14/i0_4 ) );
  NAND3_X2 \SB2_1_12/Component_Function_3/N1  ( .A1(\SB2_1_12/i1[9] ), .A2(
        \SB2_1_12/i0_3 ), .A3(\SB2_1_12/i0[6] ), .ZN(
        \SB2_1_12/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 \SB1_0_16/BUF_4_0  ( .I(\SB1_0_16/buf_output[4] ), .Z(\RI3[0][100] )
         );
  NAND3_X2 \SB1_0_5/Component_Function_5/N2  ( .A1(\SB1_0_5/i0_0 ), .A2(
        \SB1_0_5/i0[6] ), .A3(\SB1_0_5/i0[10] ), .ZN(
        \SB1_0_5/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 \SB2_3_27/Component_Function_4/N4  ( .A1(\SB2_3_27/i1[9] ), .A2(
        \SB2_3_27/i1_5 ), .A3(\SB2_3_27/i0_4 ), .ZN(
        \SB2_3_27/Component_Function_4/NAND4_in[3] ) );
  NAND3_X2 \SB2_0_21/Component_Function_2/N1  ( .A1(\SB2_0_21/i1_5 ), .A2(
        \SB2_0_21/i0[10] ), .A3(\SB2_0_21/i1[9] ), .ZN(
        \SB2_0_21/Component_Function_2/NAND4_in[0] ) );
  INV_X2 U978 ( .I(\SB1_1_18/buf_output[5] ), .ZN(\SB2_1_18/i1_5 ) );
  NAND3_X2 \SB2_0_17/Component_Function_0/N4  ( .A1(\SB2_0_17/i0[7] ), .A2(
        \SB2_0_17/i0_3 ), .A3(\SB2_0_17/i0_0 ), .ZN(
        \SB2_0_17/Component_Function_0/NAND4_in[3] ) );
  NAND3_X2 U1370 ( .A1(\SB1_2_28/i1_5 ), .A2(\SB1_2_28/i0[10] ), .A3(
        \SB1_2_28/i1[9] ), .ZN(\SB1_2_28/Component_Function_2/NAND4_in[0] ) );
  INV_X2 U1675 ( .I(\MC_ARK_ARC_1_1/buf_output[20] ), .ZN(\SB1_2_28/i1[9] ) );
  NAND3_X2 U7584 ( .A1(\SB2_3_11/i0_0 ), .A2(n4768), .A3(n3645), .ZN(
        \SB2_3_11/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 U6415 ( .A1(\SB2_0_29/i0_0 ), .A2(\SB2_0_29/i0_4 ), .A3(
        \SB2_0_29/i1_5 ), .ZN(\SB2_0_29/Component_Function_2/NAND4_in[3] ) );
  INV_X1 \SB1_0_25/INV_1  ( .I(n264), .ZN(\SB1_0_25/i1_7 ) );
  NAND3_X1 \SB1_0_21/Component_Function_1/N2  ( .A1(\SB1_0_21/i0_3 ), .A2(
        \SB1_0_21/i1_7 ), .A3(\SB1_0_21/i0[8] ), .ZN(
        \SB1_0_21/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U7267 ( .A1(\SB1_0_21/i0[6] ), .A2(\SB1_0_21/i0[9] ), .A3(
        \SB1_0_21/i1_5 ), .ZN(\SB1_0_21/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U5759 ( .A1(\SB1_0_27/i0_3 ), .A2(\SB1_0_27/i0[6] ), .A3(
        \SB1_0_27/i1[9] ), .ZN(n1769) );
  NAND3_X1 \SB1_0_3/Component_Function_4/N2  ( .A1(\SB1_0_3/i3[0] ), .A2(
        \SB1_0_3/i0_0 ), .A3(\SB1_0_3/i1_7 ), .ZN(
        \SB1_0_3/Component_Function_4/NAND4_in[1] ) );
  NAND2_X1 \SB1_0_0/Component_Function_0/N1  ( .A1(\SB1_0_0/i0[10] ), .A2(
        \SB1_0_0/i0[9] ), .ZN(\SB1_0_0/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_28/Component_Function_0/N2  ( .A1(\SB1_0_28/i0[8] ), .A2(
        \SB1_0_28/i0[7] ), .A3(\SB1_0_28/i0[6] ), .ZN(
        \SB1_0_28/Component_Function_0/NAND4_in[1] ) );
  INV_X1 \SB1_0_6/INV_0  ( .I(n320), .ZN(\SB1_0_6/i3[0] ) );
  NAND3_X1 \SB1_0_18/Component_Function_4/N2  ( .A1(\SB1_0_18/i3[0] ), .A2(
        \SB1_0_18/i0_0 ), .A3(\SB1_0_18/i1_7 ), .ZN(
        \SB1_0_18/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_13/Component_Function_1/N2  ( .A1(\SB1_0_13/i0_3 ), .A2(
        \SB1_0_13/i1_7 ), .A3(\SB1_0_13/i0[8] ), .ZN(
        \SB1_0_13/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_13/Component_Function_1/N4  ( .A1(\SB1_0_13/i1_7 ), .A2(
        \SB1_0_13/i0[8] ), .A3(\SB1_0_13/i0_4 ), .ZN(
        \SB1_0_13/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U2506 ( .A1(\SB1_0_16/i0_0 ), .A2(\SB1_0_16/i1_5 ), .A3(n4752), 
        .ZN(n673) );
  NAND3_X1 U1110 ( .A1(\SB1_0_13/i0_3 ), .A2(\SB1_0_13/i1[9] ), .A3(
        \SB1_0_13/i0_4 ), .ZN(\SB1_0_13/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_12/Component_Function_1/N2  ( .A1(\SB1_0_12/i0_3 ), .A2(
        \SB1_0_12/i1_7 ), .A3(\SB1_0_12/i0[8] ), .ZN(
        \SB1_0_12/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U4722 ( .A1(\SB1_0_7/i0_3 ), .A2(\SB1_0_7/i0[10] ), .A3(
        \SB1_0_7/i0[9] ), .ZN(n1671) );
  NAND3_X1 \SB1_0_23/Component_Function_4/N3  ( .A1(\SB1_0_23/i0[9] ), .A2(
        \SB1_0_23/i0[10] ), .A3(\SB1_0_23/i0_3 ), .ZN(
        \SB1_0_23/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U7717 ( .A1(\SB1_0_2/i0_0 ), .A2(\SB1_0_2/i3[0] ), .A3(
        \SB1_0_2/i1_7 ), .ZN(\SB1_0_2/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U4117 ( .A1(\SB1_0_28/i0[6] ), .A2(\SB1_0_28/i1_5 ), .A3(
        \SB1_0_28/i0[9] ), .ZN(\SB1_0_28/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1124 ( .A1(\SB1_0_21/i0_3 ), .A2(\SB1_0_21/i0_4 ), .A3(
        \SB1_0_21/i1[9] ), .ZN(\SB1_0_21/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_21/Component_Function_0/N3  ( .A1(\SB1_0_21/i0[10] ), .A2(
        \SB1_0_21/i0_4 ), .A3(\SB1_0_21/i0_3 ), .ZN(
        \SB1_0_21/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_11/Component_Function_5/N2  ( .A1(\SB1_0_11/i0_0 ), .A2(
        \SB1_0_11/i0[6] ), .A3(\SB1_0_11/i0[10] ), .ZN(
        \SB1_0_11/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_25/Component_Function_0/N2  ( .A1(\SB1_0_25/i0[8] ), .A2(
        \SB1_0_25/i0[7] ), .A3(\SB1_0_25/i0[6] ), .ZN(
        \SB1_0_25/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_23/Component_Function_3/N2  ( .A1(\SB1_0_23/i0_0 ), .A2(
        \SB1_0_23/i0_3 ), .A3(\SB1_0_23/i0_4 ), .ZN(
        \SB1_0_23/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_8/Component_Function_4/N1  ( .A1(\SB1_0_8/i0[9] ), .A2(
        \SB1_0_8/i0_0 ), .A3(\SB1_0_8/i0[8] ), .ZN(
        \SB1_0_8/Component_Function_4/NAND4_in[0] ) );
  INV_X1 \SB1_0_17/INV_4  ( .I(n2899), .ZN(\SB1_0_17/i0[7] ) );
  INV_X1 \SB1_0_5/INV_4  ( .I(n394), .ZN(\SB1_0_5/i0[7] ) );
  NAND3_X1 U5945 ( .A1(\SB1_0_13/i0_3 ), .A2(\SB1_0_13/i0[6] ), .A3(
        \SB1_0_13/i1[9] ), .ZN(\SB1_0_13/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_1/Component_Function_2/N3  ( .A1(\SB1_0_1/i0_3 ), .A2(
        \SB1_0_1/i0[8] ), .A3(\SB1_0_1/i0[9] ), .ZN(
        \SB1_0_1/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_10/Component_Function_5/N4  ( .A1(\SB1_0_10/i0[9] ), .A2(
        n309), .A3(n384), .ZN(\SB1_0_10/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U2566 ( .A1(\SB1_0_21/i0_3 ), .A2(\SB1_0_21/i0_0 ), .A3(
        \SB1_0_21/i0_4 ), .ZN(n869) );
  NAND3_X1 \SB1_0_3/Component_Function_0/N3  ( .A1(\SB1_0_3/i0[10] ), .A2(
        \SB1_0_3/i0_4 ), .A3(\SB1_0_3/i0_3 ), .ZN(
        \SB1_0_3/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U1949 ( .A1(\SB1_0_30/i1_5 ), .A2(\SB1_0_30/i0[8] ), .A3(
        \SB1_0_30/i3[0] ), .ZN(\SB1_0_30/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_19/Component_Function_5/N4  ( .A1(\SB1_0_19/i0[9] ), .A2(
        \SB1_0_19/i0[6] ), .A3(\SB1_0_19/i0_4 ), .ZN(
        \SB1_0_19/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U6076 ( .A1(\SB1_0_6/i0[8] ), .A2(\SB1_0_6/i1_5 ), .A3(
        \SB1_0_6/i3[0] ), .ZN(n1916) );
  NAND3_X1 \SB1_0_5/Component_Function_0/N2  ( .A1(\SB1_0_5/i0[8] ), .A2(
        \SB1_0_5/i0[7] ), .A3(\SB1_0_5/i0[6] ), .ZN(
        \SB1_0_5/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_21/Component_Function_2/N3  ( .A1(\SB1_0_21/i0_3 ), .A2(
        \SB1_0_21/i0[8] ), .A3(\SB1_0_21/i0[9] ), .ZN(
        \SB1_0_21/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_26/Component_Function_5/N4  ( .A1(\SB1_0_26/i0[9] ), .A2(
        \SB1_0_26/i0[6] ), .A3(\SB1_0_26/i0_4 ), .ZN(
        \SB1_0_26/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_14/Component_Function_3/N1  ( .A1(\SB1_0_14/i1[9] ), .A2(
        \SB1_0_14/i0_3 ), .A3(\SB1_0_14/i0[6] ), .ZN(
        \SB1_0_14/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U3014 ( .A1(\SB1_0_21/i0_3 ), .A2(\SB1_0_21/i1[9] ), .A3(
        \SB1_0_21/i0[6] ), .ZN(n832) );
  NAND3_X1 \SB1_0_23/Component_Function_1/N3  ( .A1(\SB1_0_23/i1_5 ), .A2(
        \SB1_0_23/i0[6] ), .A3(\SB1_0_23/i0[9] ), .ZN(
        \SB1_0_23/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_28/Component_Function_2/N2  ( .A1(\SB1_0_28/i0_3 ), .A2(
        \SB1_0_28/i0[10] ), .A3(\SB1_0_28/i0[6] ), .ZN(
        \SB1_0_28/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U5546 ( .A1(\SB1_0_28/i0[10] ), .A2(\SB1_0_28/i0_0 ), .A3(
        \SB1_0_28/i0[6] ), .ZN(\SB1_0_28/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_23/Component_Function_1/N4  ( .A1(\SB1_0_23/i1_7 ), .A2(
        \SB1_0_23/i0[8] ), .A3(\SB1_0_23/i0_4 ), .ZN(
        \SB1_0_23/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 U1352 ( .A1(\SB1_0_6/i0_0 ), .A2(\SB1_0_6/i3[0] ), .ZN(
        \SB1_0_6/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_15/Component_Function_5/N4  ( .A1(\SB1_0_15/i0[9] ), .A2(
        n294), .A3(n374), .ZN(\SB1_0_15/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_0_12/Component_Function_3/N2  ( .A1(\SB1_0_12/i0_0 ), .A2(
        \SB1_0_12/i0_3 ), .A3(\SB1_0_12/i0_4 ), .ZN(
        \SB1_0_12/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U7590 ( .A1(\SB1_0_1/i0_3 ), .A2(\SB1_0_1/i0_0 ), .A3(
        \SB1_0_1/i0[7] ), .ZN(\SB1_0_1/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB2_0_23/Component_Function_5/N1  ( .A1(\SB2_0_23/i0_0 ), .A2(
        \SB2_0_23/i3[0] ), .ZN(\SB2_0_23/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_29/Component_Function_5/N1  ( .A1(\SB2_0_29/i0_0 ), .A2(
        \SB2_0_29/i3[0] ), .ZN(\SB2_0_29/Component_Function_5/NAND4_in[0] ) );
  INV_X2 \SB2_0_22/INV_0  ( .I(\RI3[0][54] ), .ZN(\SB2_0_22/i3[0] ) );
  INV_X2 \SB2_0_20/INV_4  ( .I(\SB2_0_20/i0_4 ), .ZN(\SB2_0_20/i0[7] ) );
  INV_X1 \SB2_0_4/INV_1  ( .I(\RI3[0][163] ), .ZN(\SB2_0_4/i1_7 ) );
  INV_X1 \SB2_0_27/INV_1  ( .I(\SB1_0_31/buf_output[1] ), .ZN(\SB2_0_27/i1_7 )
         );
  NAND2_X1 \SB2_0_27/Component_Function_5/N1  ( .A1(\SB2_0_27/i0_0 ), .A2(
        \SB2_0_27/i3[0] ), .ZN(\SB2_0_27/Component_Function_5/NAND4_in[0] ) );
  INV_X1 \SB2_0_12/INV_0  ( .I(\RI3[0][114] ), .ZN(\SB2_0_12/i3[0] ) );
  INV_X1 \SB2_0_25/INV_0  ( .I(\SB1_0_30/buf_output[0] ), .ZN(\SB2_0_25/i3[0] ) );
  NAND3_X1 U1965 ( .A1(\SB2_0_22/i0[10] ), .A2(\SB2_0_22/i0_4 ), .A3(
        \SB2_0_22/i0_3 ), .ZN(\SB2_0_22/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_24/Component_Function_1/N3  ( .A1(\SB2_0_24/i1_5 ), .A2(
        \RI3[0][43] ), .A3(\SB1_0_29/buf_output[0] ), .ZN(
        \SB2_0_24/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_25/Component_Function_3/N3  ( .A1(\SB2_0_25/i1[9] ), .A2(
        \SB2_0_25/i1_7 ), .A3(\RI3[0][39] ), .ZN(
        \SB2_0_25/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_21/Component_Function_1/N4  ( .A1(\SB2_0_21/i1_7 ), .A2(
        \SB2_0_21/i0[8] ), .A3(\SB2_0_21/i0_4 ), .ZN(
        \SB2_0_21/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_31/Component_Function_1/N4  ( .A1(\SB2_0_31/i1_7 ), .A2(
        \SB2_0_31/i0[8] ), .A3(\RI3[0][4] ), .ZN(
        \SB2_0_31/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_6/Component_Function_1/N4  ( .A1(\SB2_0_6/i1_7 ), .A2(
        \SB2_0_6/i0[8] ), .A3(\RI3[0][154] ), .ZN(
        \SB2_0_6/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_13/Component_Function_1/N3  ( .A1(n3663), .A2(
        \SB2_0_13/i0[6] ), .A3(\SB2_0_13/i0[9] ), .ZN(
        \SB2_0_13/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1366 ( .A1(\SB2_0_12/i0[9] ), .A2(\SB2_0_12/i0_4 ), .A3(
        \SB2_0_12/i0[6] ), .ZN(n1701) );
  NAND3_X1 \SB2_0_18/Component_Function_4/N4  ( .A1(\SB2_0_18/i1[9] ), .A2(
        \SB2_0_18/i1_5 ), .A3(\RI3[0][82] ), .ZN(
        \SB2_0_18/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U1098 ( .A1(\SB2_0_11/i0[8] ), .A2(\SB2_0_11/i0_4 ), .A3(
        \SB2_0_11/i1_7 ), .ZN(n1003) );
  NAND3_X1 U4764 ( .A1(\SB2_0_26/i1[9] ), .A2(\SB2_0_26/i0_3 ), .A3(
        \SB2_0_26/i0[6] ), .ZN(\SB2_0_26/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U1979 ( .A1(\SB2_0_8/i1[9] ), .A2(\SB2_0_8/i1_5 ), .A3(
        \RI3[0][142] ), .ZN(\SB2_0_8/Component_Function_4/NAND4_in[3] ) );
  NAND2_X1 \SB2_0_18/Component_Function_5/N1  ( .A1(\SB2_0_18/i0_0 ), .A2(
        \SB2_0_18/i3[0] ), .ZN(\SB2_0_18/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U4992 ( .A1(\SB2_0_4/i0[6] ), .A2(\SB2_0_4/i0[9] ), .A3(
        \RI3[0][166] ), .ZN(n1409) );
  NAND3_X1 \SB2_0_16/Component_Function_4/N4  ( .A1(\SB2_0_16/i1[9] ), .A2(
        \SB2_0_16/i1_5 ), .A3(\SB2_0_16/i0_4 ), .ZN(
        \SB2_0_16/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_18/Component_Function_5/N3  ( .A1(\SB2_0_18/i1[9] ), .A2(
        \RI3[0][82] ), .A3(\SB2_0_18/i0_3 ), .ZN(
        \SB2_0_18/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_23/Component_Function_4/N4  ( .A1(\SB2_0_23/i1[9] ), .A2(
        \SB2_0_23/i1_5 ), .A3(\SB2_0_23/i0_4 ), .ZN(
        \SB2_0_23/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_24/Component_Function_4/N4  ( .A1(\SB2_0_24/i1[9] ), .A2(
        \SB2_0_24/i1_5 ), .A3(\RI3[0][46] ), .ZN(
        \SB2_0_24/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_17/Component_Function_1/N3  ( .A1(\SB2_0_17/i1_5 ), .A2(
        \SB2_0_17/i0[6] ), .A3(\SB2_0_17/i0[9] ), .ZN(
        \SB2_0_17/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U4380 ( .A1(n2774), .A2(\SB2_0_19/i0_3 ), .A3(\RI3[0][76] ), .ZN(
        \SB2_0_19/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_18/Component_Function_0/N3  ( .A1(\SB2_0_18/i0[10] ), .A2(
        \RI3[0][82] ), .A3(\SB2_0_18/i0_3 ), .ZN(
        \SB2_0_18/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U1455 ( .A1(\SB2_0_21/i0_3 ), .A2(\SB2_0_21/i0_4 ), .A3(
        \SB2_0_21/i0_0 ), .ZN(n1995) );
  NAND3_X1 U1978 ( .A1(n2237), .A2(\SB2_0_27/i0[8] ), .A3(\SB2_0_27/i0[6] ), 
        .ZN(n2239) );
  NAND3_X1 \SB2_0_24/Component_Function_1/N4  ( .A1(\SB2_0_24/i1_7 ), .A2(
        \SB2_0_24/i0[8] ), .A3(\RI3[0][46] ), .ZN(
        \SB2_0_24/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_6/Component_Function_5/N2  ( .A1(\SB2_0_6/i0_0 ), .A2(
        \SB2_0_6/i0[6] ), .A3(n2765), .ZN(
        \SB2_0_6/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_5/Component_Function_1/N2  ( .A1(\SB2_0_5/i0_3 ), .A2(
        \SB2_0_5/i1_7 ), .A3(\SB2_0_5/i0[8] ), .ZN(
        \SB2_0_5/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U1967 ( .A1(\SB2_0_22/i0_3 ), .A2(\SB2_0_22/i0[8] ), .A3(
        \SB2_0_22/i1_7 ), .ZN(\SB2_0_22/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U1080 ( .A1(\SB2_0_22/i0_3 ), .A2(\SB2_0_22/i0[10] ), .A3(
        \RI3[0][54] ), .ZN(\SB2_0_22/Component_Function_4/NAND4_in[2] ) );
  NAND2_X1 U2396 ( .A1(n3689), .A2(\SB2_0_5/i0_3 ), .ZN(
        \SB2_0_5/Component_Function_1/NAND4_in[0] ) );
  INV_X1 U7 ( .I(n17), .ZN(n545) );
  INV_X1 U8 ( .I(n33), .ZN(n462) );
  INV_X1 \SB1_1_20/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[66] ), .ZN(
        \SB1_1_20/i3[0] ) );
  BUF_X2 \SB1_1_5/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[160] ), .Z(
        \SB1_1_5/i0_4 ) );
  INV_X1 \SB1_1_5/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[156] ), .ZN(
        \SB1_1_5/i3[0] ) );
  BUF_X2 \SB1_1_1/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[181] ), .Z(
        \SB1_1_1/i0[6] ) );
  INV_X1 \SB1_1_25/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[37] ), .ZN(
        \SB1_1_25/i1_7 ) );
  BUF_X2 U1907 ( .I(\MC_ARK_ARC_1_0/buf_output[108] ), .Z(\SB1_1_13/i0[9] ) );
  BUF_X2 \SB1_1_10/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[130] ), .Z(
        \SB1_1_10/i0_4 ) );
  NAND3_X1 U1991 ( .A1(\SB1_1_18/i0_4 ), .A2(\SB1_1_18/i0[10] ), .A3(
        \SB1_1_18/i0_3 ), .ZN(n1755) );
  NAND3_X1 \SB1_1_5/Component_Function_2/N4  ( .A1(\SB1_1_5/i1_5 ), .A2(
        \SB1_1_5/i0_0 ), .A3(\SB1_1_5/i0_4 ), .ZN(
        \SB1_1_5/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_21/Component_Function_0/N2  ( .A1(\SB1_1_21/i0[8] ), .A2(
        \SB1_1_21/i0[7] ), .A3(\SB1_1_21/i0[6] ), .ZN(
        \SB1_1_21/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_28/Component_Function_1/N1  ( .A1(\SB1_1_28/i0_3 ), .A2(
        \SB1_1_28/i1[9] ), .ZN(\SB1_1_28/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_25/Component_Function_4/N4  ( .A1(\SB1_1_25/i1[9] ), .A2(
        \SB1_1_25/i1_5 ), .A3(\SB1_1_25/i0_4 ), .ZN(
        \SB1_1_25/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_14/Component_Function_0/N4  ( .A1(\SB1_1_14/i0[7] ), .A2(
        \SB1_1_14/i0_3 ), .A3(\SB1_1_14/i0_0 ), .ZN(
        \SB1_1_14/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_28/Component_Function_1/N4  ( .A1(\SB1_1_28/i1_7 ), .A2(
        \SB1_1_28/i0[8] ), .A3(\SB1_1_28/i0_4 ), .ZN(
        \SB1_1_28/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB1_1_4/Component_Function_5/N1  ( .A1(\SB1_1_4/i0_0 ), .A2(
        \SB1_1_4/i3[0] ), .ZN(\SB1_1_4/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_15/Component_Function_0/N2  ( .A1(\SB1_1_15/i0[8] ), .A2(
        \SB1_1_15/i0[7] ), .A3(\SB1_1_15/i0[6] ), .ZN(
        \SB1_1_15/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U999 ( .A1(\SB1_1_11/i1_7 ), .A2(\SB1_1_11/i0_4 ), .A3(
        \SB1_1_11/i0[8] ), .ZN(n909) );
  NAND3_X1 U6905 ( .A1(\SB1_1_0/i0_0 ), .A2(\SB1_1_0/i3[0] ), .A3(
        \SB1_1_0/i1_7 ), .ZN(\SB1_1_0/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_3/Component_Function_4/N2  ( .A1(\SB1_1_3/i3[0] ), .A2(
        \SB1_1_3/i0_0 ), .A3(\SB1_1_3/i1_7 ), .ZN(
        \SB1_1_3/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_15/Component_Function_2/N1  ( .A1(\SB1_1_15/i1_5 ), .A2(
        \SB1_1_15/i0[10] ), .A3(\SB1_1_15/i1[9] ), .ZN(
        \SB1_1_15/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_24/Component_Function_0/N4  ( .A1(\SB1_1_24/i0[7] ), .A2(
        \SB1_1_24/i0_3 ), .A3(\SB1_1_24/i0_0 ), .ZN(
        \SB1_1_24/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_1/Component_Function_4/N4  ( .A1(\SB1_1_1/i1[9] ), .A2(
        \SB1_1_1/i1_5 ), .A3(\SB1_1_1/i0_4 ), .ZN(
        \SB1_1_1/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U1700 ( .A1(\SB1_1_7/i1[9] ), .A2(\SB1_1_7/i1_5 ), .A3(
        \SB1_1_7/i0_4 ), .ZN(\SB1_1_7/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U1052 ( .A1(\SB1_1_12/i0_0 ), .A2(\SB1_1_12/i3[0] ), .A3(
        \SB1_1_12/i1_7 ), .ZN(n1775) );
  NAND3_X1 U1046 ( .A1(\SB1_1_24/i0[10] ), .A2(\SB1_1_24/i0_3 ), .A3(
        \SB1_1_24/i0[9] ), .ZN(\SB1_1_24/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U4206 ( .A1(\SB1_1_20/i0_3 ), .A2(\SB1_1_20/i1[9] ), .A3(
        \SB1_1_20/i0[6] ), .ZN(\SB1_1_20/Component_Function_3/NAND4_in[0] ) );
  NAND2_X1 U2015 ( .A1(\SB1_1_18/Component_Function_0/NAND4_in[0] ), .A2(n1755), .ZN(n1754) );
  NAND3_X1 U5464 ( .A1(\SB1_1_24/i0[10] ), .A2(\SB1_1_24/i0_3 ), .A3(
        \SB1_1_24/i0_4 ), .ZN(\SB1_1_24/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_1_24/Component_Function_0/N1  ( .A1(\SB1_1_24/i0[10] ), .A2(
        \SB1_1_24/i0[9] ), .ZN(\SB1_1_24/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U1005 ( .A1(\SB1_1_24/i0_3 ), .A2(\SB1_1_24/i0[6] ), .A3(
        \SB1_1_24/i0[10] ), .ZN(\SB1_1_24/Component_Function_2/NAND4_in[1] )
         );
  NAND2_X1 U6726 ( .A1(\SB1_1_23/i0[6] ), .A2(n2224), .ZN(
        \SB1_1_23/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_4/Component_Function_3/N1  ( .A1(\SB1_1_4/i1[9] ), .A2(
        \SB1_1_4/i0_3 ), .A3(\SB1_1_4/i0[6] ), .ZN(
        \SB1_1_4/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_12/Component_Function_5/N4  ( .A1(\SB1_1_12/i0[9] ), .A2(
        \SB1_1_12/i0[6] ), .A3(\MC_ARK_ARC_1_0/buf_output[118] ), .ZN(
        \SB1_1_12/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_27/Component_Function_3/N2  ( .A1(\SB1_1_27/i0_0 ), .A2(
        \SB1_1_27/i0_3 ), .A3(\SB1_1_27/i0_4 ), .ZN(
        \SB1_1_27/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U4232 ( .A1(\SB1_1_28/i0[6] ), .A2(\SB1_1_28/i1_5 ), .A3(
        \SB1_1_28/i0[9] ), .ZN(\SB1_1_28/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1995 ( .A1(\SB1_1_26/i0_0 ), .A2(\SB1_1_26/i0_3 ), .A3(
        \SB1_1_26/i0_4 ), .ZN(\SB1_1_26/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U7307 ( .A1(\SB1_1_4/i0_0 ), .A2(\SB1_1_4/i0[9] ), .A3(
        \SB1_1_4/i0[8] ), .ZN(n2510) );
  NAND3_X1 \SB1_1_18/Component_Function_3/N1  ( .A1(\SB1_1_18/i1[9] ), .A2(
        \SB1_1_18/i0_3 ), .A3(\SB1_1_18/i0[6] ), .ZN(
        \SB1_1_18/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U1998 ( .A1(\SB1_1_8/i1_7 ), .A2(\SB1_1_8/i0[8] ), .A3(
        \SB1_1_8/i0_4 ), .ZN(\SB1_1_8/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_4/Component_Function_3/N2  ( .A1(\SB1_1_4/i0_0 ), .A2(
        \SB1_1_4/i0_3 ), .A3(\SB1_1_4/i0_4 ), .ZN(
        \SB1_1_4/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_23/Component_Function_3/N3  ( .A1(\SB1_1_23/i1[9] ), .A2(
        \SB1_1_23/i1_7 ), .A3(\SB1_1_23/i0[10] ), .ZN(
        \SB1_1_23/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U7286 ( .A1(\SB1_1_19/i0_0 ), .A2(\SB1_1_19/i0[7] ), .A3(
        \SB1_1_19/i0_3 ), .ZN(\SB1_1_19/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_29/Component_Function_3/N3  ( .A1(\SB1_1_29/i1[9] ), .A2(
        \SB1_1_29/i1_7 ), .A3(\SB1_1_29/i0[10] ), .ZN(
        \SB1_1_29/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2591 ( .A1(\SB1_1_3/i0_0 ), .A2(\SB1_1_3/i0_4 ), .A3(
        \SB1_1_3/i1_5 ), .ZN(n741) );
  NAND3_X1 \SB1_1_13/Component_Function_0/N2  ( .A1(\SB1_1_13/i0[8] ), .A2(
        \SB1_1_13/i0[7] ), .A3(\SB1_1_13/i0[6] ), .ZN(
        \SB1_1_13/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U2639 ( .A1(\SB1_1_7/i0[8] ), .A2(\SB1_1_7/i0_4 ), .A3(
        \SB1_1_7/i1_7 ), .ZN(\SB1_1_7/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U7204 ( .A1(\SB1_1_0/i0[9] ), .A2(\SB1_1_0/i0[6] ), .A3(
        \SB1_1_0/i1_5 ), .ZN(n2440) );
  NAND3_X1 \SB1_1_5/Component_Function_3/N2  ( .A1(\SB1_1_5/i0_0 ), .A2(
        \SB1_1_5/i0_3 ), .A3(\SB1_1_5/i0_4 ), .ZN(
        \SB1_1_5/Component_Function_3/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_16/Component_Function_0/N1  ( .A1(\SB1_1_16/i0[10] ), .A2(
        \SB1_1_16/i0[9] ), .ZN(\SB1_1_16/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_27/Component_Function_0/N3  ( .A1(\SB1_1_27/i0[10] ), .A2(
        \SB1_1_27/i0_4 ), .A3(\SB1_1_27/i0_3 ), .ZN(
        \SB1_1_27/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_29/Component_Function_4/N4  ( .A1(\SB1_1_29/i1[9] ), .A2(
        \SB1_1_29/i1_5 ), .A3(\SB1_1_29/i0_4 ), .ZN(
        \SB1_1_29/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_19/Component_Function_1/N2  ( .A1(\SB1_1_19/i0_3 ), .A2(
        \SB1_1_19/i1_7 ), .A3(\SB1_1_19/i0[8] ), .ZN(
        \SB1_1_19/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_28/Component_Function_4/N1  ( .A1(\SB1_1_28/i0[9] ), .A2(
        \SB1_1_28/i0_0 ), .A3(\SB1_1_28/i0[8] ), .ZN(
        \SB1_1_28/Component_Function_4/NAND4_in[0] ) );
  INV_X2 U7968 ( .I(n2885), .ZN(\SB1_1_18/buf_output[0] ) );
  INV_X1 \SB2_1_1/INV_0  ( .I(\SB1_1_6/buf_output[0] ), .ZN(\SB2_1_1/i3[0] )
         );
  INV_X1 U1397 ( .I(\SB1_1_4/buf_output[0] ), .ZN(\SB2_1_31/i3[0] ) );
  NAND2_X1 \SB2_1_4/Component_Function_5/N1  ( .A1(\SB1_1_7/buf_output[2] ), 
        .A2(\SB2_1_4/i3[0] ), .ZN(\SB2_1_4/Component_Function_5/NAND4_in[0] )
         );
  INV_X1 U6660 ( .I(\SB1_1_24/buf_output[1] ), .ZN(\SB2_1_20/i1_7 ) );
  INV_X1 \SB2_1_12/INV_1  ( .I(\SB1_1_16/buf_output[1] ), .ZN(\SB2_1_12/i1_7 )
         );
  INV_X1 \SB2_1_7/INV_1  ( .I(\SB1_1_11/buf_output[1] ), .ZN(\SB2_1_7/i1_7 )
         );
  INV_X1 \SB2_1_8/INV_0  ( .I(\SB1_1_13/buf_output[0] ), .ZN(\SB2_1_8/i3[0] )
         );
  NAND2_X1 \SB2_1_13/Component_Function_5/N1  ( .A1(\SB2_1_13/i0_0 ), .A2(
        n4182), .ZN(\SB2_1_13/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 U7483 ( .A1(\SB2_1_21/i0_0 ), .A2(n4625), .ZN(
        \SB2_1_21/Component_Function_5/NAND4_in[0] ) );
  INV_X1 \SB2_1_27/INV_0  ( .I(\SB1_1_0/buf_output[0] ), .ZN(\SB2_1_27/i3[0] )
         );
  NAND3_X1 \SB2_1_14/Component_Function_4/N2  ( .A1(\SB2_1_14/i3[0] ), .A2(
        \SB2_1_14/i0_0 ), .A3(\SB2_1_14/i1_7 ), .ZN(
        \SB2_1_14/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U6443 ( .A1(\SB2_1_29/i0_0 ), .A2(\SB2_1_29/i0_4 ), .A3(
        \SB2_1_29/i0_3 ), .ZN(\SB2_1_29/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_25/Component_Function_1/N4  ( .A1(\SB2_1_25/i1_7 ), .A2(
        \SB2_1_25/i0[8] ), .A3(n1579), .ZN(
        \SB2_1_25/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_1/Component_Function_3/N4  ( .A1(\SB2_1_1/i1_5 ), .A2(
        \SB2_1_1/i0[8] ), .A3(\SB2_1_1/i3[0] ), .ZN(
        \SB2_1_1/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_13/Component_Function_0/N2  ( .A1(\SB2_1_13/i0[8] ), .A2(
        \SB2_1_13/i0[7] ), .A3(\SB2_1_13/i0[6] ), .ZN(
        \SB2_1_13/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_19/Component_Function_4/N2  ( .A1(\SB2_1_19/i3[0] ), .A2(
        \SB1_1_22/buf_output[2] ), .A3(\SB2_1_19/i1_7 ), .ZN(
        \SB2_1_19/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U2042 ( .A1(\SB2_1_17/i0[8] ), .A2(\SB2_1_17/i0[7] ), .A3(
        \SB2_1_17/i0[6] ), .ZN(\SB2_1_17/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_20/Component_Function_0/N2  ( .A1(\SB2_1_20/i0[8] ), .A2(
        \SB2_1_20/i0[7] ), .A3(\SB2_1_20/i0[6] ), .ZN(
        \SB2_1_20/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_2/Component_Function_3/N4  ( .A1(\SB2_1_2/i1_5 ), .A2(
        \SB2_1_2/i0[8] ), .A3(\SB2_1_2/i3[0] ), .ZN(
        \SB2_1_2/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_31/Component_Function_1/N2  ( .A1(\SB2_1_31/i0_3 ), .A2(
        \SB2_1_31/i1_7 ), .A3(\SB2_1_31/i0[8] ), .ZN(
        \SB2_1_31/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_12/Component_Function_3/N4  ( .A1(\SB2_1_12/i1_5 ), .A2(
        \SB2_1_12/i0[8] ), .A3(\SB2_1_12/i3[0] ), .ZN(
        \SB2_1_12/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_16/Component_Function_4/N2  ( .A1(\SB2_1_16/i3[0] ), .A2(
        \SB2_1_16/i0_0 ), .A3(\SB2_1_16/i1_7 ), .ZN(
        \SB2_1_16/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_17/Component_Function_0/N4  ( .A1(\SB2_1_17/i0[7] ), .A2(
        \SB2_1_17/i0_3 ), .A3(\SB2_1_17/i0_0 ), .ZN(
        \SB2_1_17/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U975 ( .A1(n3690), .A2(\SB2_1_30/i0_3 ), .A3(\SB2_1_30/i0[9] ), 
        .ZN(\SB2_1_30/Component_Function_4/NAND4_in[2] ) );
  NAND2_X1 \SB2_1_22/Component_Function_5/N1  ( .A1(\SB2_1_22/i0_0 ), .A2(
        \SB2_1_22/i3[0] ), .ZN(\SB2_1_22/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_17/Component_Function_4/N4  ( .A1(\SB2_1_17/i1[9] ), .A2(
        \SB2_1_17/i1_5 ), .A3(\SB2_1_17/i0_4 ), .ZN(
        \SB2_1_17/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_13/Component_Function_4/N1  ( .A1(\SB1_1_18/buf_output[0] ), 
        .A2(\SB2_1_13/i0_0 ), .A3(\SB2_1_13/i0[8] ), .ZN(
        \SB2_1_13/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_11/Component_Function_4/N4  ( .A1(\SB2_1_11/i1[9] ), .A2(
        \SB2_1_11/i1_5 ), .A3(\SB1_1_12/buf_output[4] ), .ZN(
        \SB2_1_11/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_14/Component_Function_1/N3  ( .A1(\SB2_1_14/i1_5 ), .A2(
        \SB2_1_14/i0[6] ), .A3(\SB2_1_14/i0[9] ), .ZN(
        \SB2_1_14/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_19/Component_Function_4/N1  ( .A1(\SB2_1_19/i0[9] ), .A2(
        \SB1_1_22/buf_output[2] ), .A3(\SB2_1_19/i0[8] ), .ZN(
        \SB2_1_19/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_17/Component_Function_0/N3  ( .A1(\SB2_1_17/i0[10] ), .A2(
        \SB2_1_17/i0_4 ), .A3(\SB2_1_17/i0_3 ), .ZN(
        \SB2_1_17/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB2_1_24/Component_Function_0/N1  ( .A1(\SB2_1_24/i0[10] ), .A2(
        \SB2_1_24/i0[9] ), .ZN(\SB2_1_24/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U4163 ( .A1(n2745), .A2(\SB2_1_8/i0_3 ), .A3(\SB2_1_8/i0[10] ), 
        .ZN(\SB2_1_8/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_18/Component_Function_0/N2  ( .A1(\SB2_1_18/i0[8] ), .A2(
        n1379), .A3(\SB1_1_22/buf_output[1] ), .ZN(
        \SB2_1_18/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_16/Component_Function_4/N1  ( .A1(\SB2_1_16/i0[9] ), .A2(
        \SB2_1_16/i0_0 ), .A3(\SB2_1_16/i0[8] ), .ZN(
        \SB2_1_16/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_26/Component_Function_1/N4  ( .A1(\SB2_1_26/i1_7 ), .A2(
        \SB2_1_26/i0[8] ), .A3(\SB2_1_26/i0_4 ), .ZN(
        \SB2_1_26/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U4700 ( .A1(\SB2_1_28/i0_3 ), .A2(\SB2_1_28/i0_0 ), .A3(
        \SB1_1_29/buf_output[4] ), .ZN(
        \SB2_1_28/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U5655 ( .A1(\SB2_1_24/i0_3 ), .A2(\SB2_1_24/i0[10] ), .A3(
        \SB2_1_24/i0_4 ), .ZN(\SB2_1_24/Component_Function_0/NAND4_in[2] ) );
  INV_X1 \SB1_2_6/INV_1  ( .I(\MC_ARK_ARC_1_1/buf_output[151] ), .ZN(
        \SB1_2_6/i1_7 ) );
  INV_X1 \SB1_2_11/INV_1  ( .I(\MC_ARK_ARC_1_1/buf_output[121] ), .ZN(
        \SB1_2_11/i1_7 ) );
  NAND3_X1 U902 ( .A1(\SB1_2_11/i0[9] ), .A2(\SB1_2_11/i0[10] ), .A3(
        \SB1_2_11/i0_3 ), .ZN(n1569) );
  NAND3_X1 \SB1_2_2/Component_Function_4/N4  ( .A1(\SB1_2_2/i1[9] ), .A2(
        \SB1_2_2/i1_5 ), .A3(\SB1_2_2/i0_4 ), .ZN(
        \SB1_2_2/Component_Function_4/NAND4_in[3] ) );
  BUF_X2 \SB1_2_27/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[25] ), .Z(
        \SB1_2_27/i0[6] ) );
  NAND3_X1 \SB1_2_6/Component_Function_4/N2  ( .A1(\SB1_2_6/i3[0] ), .A2(
        \SB1_2_6/i0_0 ), .A3(\SB1_2_6/i1_7 ), .ZN(
        \SB1_2_6/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_0/Component_Function_4/N1  ( .A1(\SB1_2_0/i0[9] ), .A2(
        \SB1_2_0/i0_0 ), .A3(\SB1_2_0/i0[8] ), .ZN(
        \SB1_2_0/Component_Function_4/NAND4_in[0] ) );
  INV_X1 \SB1_2_15/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[96] ), .ZN(
        \SB1_2_15/i3[0] ) );
  NAND3_X1 \SB1_2_27/Component_Function_0/N4  ( .A1(\SB1_2_27/i0[7] ), .A2(
        \SB1_2_27/i0_3 ), .A3(\SB1_2_27/i0_0 ), .ZN(
        \SB1_2_27/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_10/Component_Function_1/N2  ( .A1(\SB1_2_10/i0_3 ), .A2(
        \SB1_2_10/i1_7 ), .A3(\SB1_2_10/i0[8] ), .ZN(
        \SB1_2_10/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U5960 ( .A1(\SB1_2_21/i0[10] ), .A2(\SB1_2_21/i1[9] ), .A3(
        \SB1_2_21/i1_7 ), .ZN(n1854) );
  NAND3_X1 U932 ( .A1(\SB1_2_12/i0[9] ), .A2(\SB1_2_12/i0[10] ), .A3(
        \SB1_2_12/i0_3 ), .ZN(\SB1_2_12/Component_Function_4/NAND4_in[2] ) );
  NAND2_X1 \SB1_2_15/Component_Function_5/N1  ( .A1(\SB1_2_15/i0_0 ), .A2(
        \SB1_2_15/i3[0] ), .ZN(\SB1_2_15/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_26/Component_Function_4/N2  ( .A1(\SB1_2_26/i3[0] ), .A2(
        \SB1_2_26/i0_0 ), .A3(\SB1_2_26/i1_7 ), .ZN(
        \SB1_2_26/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_22/Component_Function_3/N4  ( .A1(\SB1_2_22/i1_5 ), .A2(
        \SB1_2_22/i0[8] ), .A3(\SB1_2_22/i3[0] ), .ZN(
        \SB1_2_22/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U3335 ( .A1(\SB1_2_20/i0[6] ), .A2(n2909), .A3(\SB1_2_20/i0[9] ), 
        .ZN(n952) );
  NAND3_X1 \SB1_2_7/Component_Function_4/N4  ( .A1(\SB1_2_7/i1[9] ), .A2(
        \SB1_2_7/i1_5 ), .A3(\SB1_2_7/i0_4 ), .ZN(
        \SB1_2_7/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_22/Component_Function_1/N4  ( .A1(\SB1_2_22/i1_7 ), .A2(
        \SB1_2_22/i0[8] ), .A3(\SB1_2_22/i0_4 ), .ZN(
        \SB1_2_22/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB1_2_19/Component_Function_5/N1  ( .A1(\SB1_2_19/i0_0 ), .A2(
        \SB1_2_19/i3[0] ), .ZN(\SB1_2_19/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_19/Component_Function_1/N3  ( .A1(\SB1_2_19/i1_5 ), .A2(
        \SB1_2_19/i0[6] ), .A3(\SB1_2_19/i0[9] ), .ZN(
        \SB1_2_19/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U888 ( .A1(\SB1_2_17/i0_0 ), .A2(\SB1_2_17/i1_5 ), .A3(
        \SB1_2_17/i0_4 ), .ZN(\SB1_2_17/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U7916 ( .A1(\SB1_2_21/i0_3 ), .A2(\SB1_2_21/i1[9] ), .A3(
        \SB1_2_21/i0_4 ), .ZN(n2862) );
  NAND3_X1 \SB1_2_6/Component_Function_3/N1  ( .A1(\SB1_2_6/i1[9] ), .A2(
        \SB1_2_6/i0_3 ), .A3(\SB1_2_6/i0[6] ), .ZN(
        \SB1_2_6/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U862 ( .A1(\SB1_2_11/i0[6] ), .A2(\SB1_2_11/i0[10] ), .A3(
        \SB1_2_11/i0_3 ), .ZN(\SB1_2_11/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_5/Component_Function_1/N4  ( .A1(\SB1_2_5/i1_7 ), .A2(
        \SB1_2_5/i0[8] ), .A3(\SB1_2_5/i0_4 ), .ZN(
        \SB1_2_5/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_22/Component_Function_0/N2  ( .A1(\SB1_2_22/i0[8] ), .A2(
        \SB1_2_22/i0[7] ), .A3(\SB1_2_22/i0[6] ), .ZN(
        \SB1_2_22/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_18/Component_Function_1/N4  ( .A1(\SB1_2_18/i1_7 ), .A2(
        n4762), .A3(\SB1_2_18/i0_4 ), .ZN(
        \SB1_2_18/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_28/Component_Function_1/N3  ( .A1(\SB1_2_28/i1_5 ), .A2(
        \SB1_2_28/i0[6] ), .A3(\SB1_2_28/i0[9] ), .ZN(
        \SB1_2_28/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_0/Component_Function_5/N2  ( .A1(\SB1_2_0/i0_0 ), .A2(
        \SB1_2_0/i0[6] ), .A3(\SB1_2_0/i0[10] ), .ZN(
        \SB1_2_0/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_12/Component_Function_5/N2  ( .A1(\SB1_2_12/i0_0 ), .A2(
        \SB1_2_12/i0[6] ), .A3(\SB1_2_12/i0[10] ), .ZN(
        \SB1_2_12/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U2059 ( .A1(\SB1_2_29/i1_5 ), .A2(\SB1_2_29/i0[6] ), .A3(
        \SB1_2_29/i0[9] ), .ZN(\SB1_2_29/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_3/Component_Function_4/N1  ( .A1(\SB1_2_3/i0[9] ), .A2(
        \SB1_2_3/i0_0 ), .A3(\SB1_2_3/i0[8] ), .ZN(
        \SB1_2_3/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_23/Component_Function_0/N4  ( .A1(\SB1_2_23/i0[7] ), .A2(
        \SB1_2_23/i0_3 ), .A3(\SB1_2_23/i0_0 ), .ZN(
        \SB1_2_23/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_3/Component_Function_0/N4  ( .A1(\SB1_2_3/i0[7] ), .A2(
        \SB1_2_3/i0_3 ), .A3(\SB1_2_3/i0_0 ), .ZN(
        \SB1_2_3/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U6745 ( .A1(\SB1_2_2/i0[10] ), .A2(\SB1_2_2/i1[9] ), .A3(
        \SB1_2_2/i1_7 ), .ZN(\SB1_2_2/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U901 ( .A1(\SB1_2_16/i0_0 ), .A2(\RI1[2][95] ), .A3(\SB1_2_16/i0_4 ), .ZN(\SB1_2_16/Component_Function_3/NAND4_in[1] ) );
  NAND2_X1 \SB1_2_15/Component_Function_1/N1  ( .A1(\SB1_2_15/i0_3 ), .A2(
        \SB1_2_15/i1[9] ), .ZN(\SB1_2_15/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_6/Component_Function_1/N3  ( .A1(\SB1_2_6/i1_5 ), .A2(
        \SB1_2_6/i0[6] ), .A3(\SB1_2_6/i0[9] ), .ZN(
        \SB1_2_6/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U6988 ( .A1(\SB1_2_1/i0[8] ), .A2(\SB1_2_1/i0_4 ), .A3(
        \SB1_2_1/i1_7 ), .ZN(\SB1_2_1/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U4427 ( .A1(\SB1_2_3/i0_3 ), .A2(\SB1_2_3/i0[10] ), .A3(
        \SB1_2_3/i0[6] ), .ZN(\SB1_2_3/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U7596 ( .A1(\SB1_2_21/i0_3 ), .A2(\SB1_2_21/i0_0 ), .A3(
        \SB1_2_21/i0_4 ), .ZN(\SB1_2_21/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U875 ( .A1(\SB1_2_12/i0_3 ), .A2(\SB1_2_12/i0[10] ), .A3(
        \SB1_2_12/i0_4 ), .ZN(n1169) );
  INV_X1 \SB2_2_6/INV_0  ( .I(\SB1_2_11/buf_output[0] ), .ZN(\SB2_2_6/i3[0] )
         );
  INV_X1 \SB2_2_24/INV_1  ( .I(\SB1_2_28/buf_output[1] ), .ZN(\SB2_2_24/i1_7 )
         );
  BUF_X2 \SB2_2_21/BUF_0  ( .I(\SB1_2_26/buf_output[0] ), .Z(\SB2_2_21/i0[9] )
         );
  INV_X1 \SB2_2_28/INV_1  ( .I(\SB1_2_0/buf_output[1] ), .ZN(\SB2_2_28/i1_7 )
         );
  NAND3_X1 \SB2_2_31/Component_Function_0/N4  ( .A1(\SB2_2_31/i0[7] ), .A2(
        \SB2_2_31/i0_3 ), .A3(\SB2_2_31/i0_0 ), .ZN(
        \SB2_2_31/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_20/Component_Function_1/N2  ( .A1(\SB2_2_20/i0_3 ), .A2(
        \SB2_2_20/i1_7 ), .A3(\SB2_2_20/i0[8] ), .ZN(
        \SB2_2_20/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U3417 ( .A1(\SB2_2_4/i0_3 ), .A2(\SB2_2_4/i1_7 ), .A3(
        \SB2_2_4/i0[8] ), .ZN(\SB2_2_4/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U3704 ( .A1(\SB2_2_21/i0_3 ), .A2(\SB2_2_21/i0_0 ), .A3(
        \SB2_2_21/i0[7] ), .ZN(n1086) );
  NAND3_X1 U824 ( .A1(\SB2_2_13/i3[0] ), .A2(\SB2_2_13/i0[8] ), .A3(n1394), 
        .ZN(n2152) );
  NAND2_X1 \SB2_2_18/Component_Function_5/N1  ( .A1(\SB2_2_18/i0_0 ), .A2(
        \SB2_2_18/i3[0] ), .ZN(\SB2_2_18/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_9/Component_Function_5/N1  ( .A1(\SB2_2_9/i0_0 ), .A2(
        \SB2_2_9/i3[0] ), .ZN(\SB2_2_9/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_1/Component_Function_5/N1  ( .A1(\SB2_2_1/i0_0 ), .A2(
        \SB2_2_1/i3[0] ), .ZN(\SB2_2_1/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U1492 ( .A1(\SB2_2_11/i0_3 ), .A2(\SB1_2_12/buf_output[4] ), .A3(
        n5515), .ZN(\SB2_2_11/Component_Function_5/NAND4_in[2] ) );
  INV_X1 \SB2_2_29/INV_4  ( .I(\SB2_2_29/i0_4 ), .ZN(\SB2_2_29/i0[7] ) );
  NAND2_X1 \SB2_2_0/Component_Function_1/N1  ( .A1(\SB2_2_0/i0_3 ), .A2(
        \SB2_2_0/i1[9] ), .ZN(\SB2_2_0/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_9/Component_Function_0/N4  ( .A1(n3333), .A2(\SB2_2_9/i0_3 ), 
        .A3(\SB2_2_9/i0_0 ), .ZN(\SB2_2_9/Component_Function_0/NAND4_in[3] )
         );
  NAND3_X1 U5059 ( .A1(\SB2_2_8/i0[7] ), .A2(\SB2_2_8/i0_0 ), .A3(
        \SB2_2_8/i0_3 ), .ZN(n1438) );
  NAND3_X1 \SB2_2_20/Component_Function_3/N4  ( .A1(\SB2_2_20/i1_5 ), .A2(
        \SB2_2_20/i0[8] ), .A3(\SB2_2_20/i3[0] ), .ZN(
        \SB2_2_20/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_9/Component_Function_4/N1  ( .A1(\SB2_2_9/i0[9] ), .A2(
        \SB2_2_9/i0_0 ), .A3(\SB2_2_9/i0[8] ), .ZN(
        \SB2_2_9/Component_Function_4/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_7/Component_Function_1/N1  ( .A1(\SB2_2_7/i0_3 ), .A2(
        \SB2_2_7/i1[9] ), .ZN(\SB2_2_7/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_13/Component_Function_1/N1  ( .A1(\SB2_2_13/i0_3 ), .A2(
        \SB2_2_13/i1[9] ), .ZN(\SB2_2_13/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_19/Component_Function_0/N1  ( .A1(\SB2_2_19/i0[10] ), .A2(
        \SB2_2_19/i0[9] ), .ZN(\SB2_2_19/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U840 ( .A1(\SB2_2_8/i0[7] ), .A2(\SB2_2_8/i0[8] ), .A3(
        \SB2_2_8/i0[6] ), .ZN(\SB2_2_8/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_24/Component_Function_0/N4  ( .A1(\SB2_2_24/i0[7] ), .A2(
        \SB2_2_24/i0_3 ), .A3(\SB2_2_24/i0_0 ), .ZN(
        \SB2_2_24/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_24/Component_Function_0/N3  ( .A1(\SB2_2_24/i0[10] ), .A2(
        \SB2_2_24/i0_4 ), .A3(\SB2_2_24/i0_3 ), .ZN(
        \SB2_2_24/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U4209 ( .A1(\SB2_2_9/i3[0] ), .A2(n3687), .A3(\SB2_2_9/i0[8] ), 
        .ZN(n1481) );
  INV_X4 \SB1_3_29/INV_2  ( .I(\RI1[3][14] ), .ZN(\SB1_3_29/i1[9] ) );
  BUF_X2 \SB1_3_17/BUF_0  ( .I(\MC_ARK_ARC_1_2/buf_output[84] ), .Z(
        \SB1_3_17/i0[9] ) );
  BUF_X2 \SB1_3_1/BUF_0  ( .I(\MC_ARK_ARC_1_2/buf_output[180] ), .Z(
        \SB1_3_1/i0[9] ) );
  INV_X1 U4807 ( .I(\MC_ARK_ARC_1_2/buf_output[145] ), .ZN(\SB1_3_7/i1_7 ) );
  NAND3_X1 U2111 ( .A1(\SB1_3_8/i0_3 ), .A2(\SB1_3_8/i0[10] ), .A3(
        \SB1_3_8/i0[9] ), .ZN(n606) );
  INV_X1 \SB1_3_21/INV_1  ( .I(\MC_ARK_ARC_1_2/buf_output[61] ), .ZN(
        \SB1_3_21/i1_7 ) );
  INV_X1 U2112 ( .I(\MC_ARK_ARC_1_2/buf_output[127] ), .ZN(\SB1_3_10/i1_7 ) );
  INV_X1 U1647 ( .I(\MC_ARK_ARC_1_2/buf_output[149] ), .ZN(\SB1_3_7/i1_5 ) );
  INV_X1 \SB1_3_30/INV_5  ( .I(\MC_ARK_ARC_1_2/buf_output[11] ), .ZN(
        \SB1_3_30/i1_5 ) );
  NAND2_X1 \SB1_3_28/Component_Function_0/N1  ( .A1(\SB1_3_28/i0[10] ), .A2(
        \SB1_3_28/i0[9] ), .ZN(\SB1_3_28/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U777 ( .A1(\SB1_3_23/i0[8] ), .A2(\SB1_3_23/i3[0] ), .A3(
        \SB1_3_23/i1_5 ), .ZN(n1712) );
  NAND3_X1 U6547 ( .A1(\SB1_3_25/i0[6] ), .A2(\SB1_3_25/i1_5 ), .A3(
        \SB1_3_25/i0[9] ), .ZN(n2125) );
  NAND3_X1 \SB1_3_16/Component_Function_3/N4  ( .A1(\SB1_3_16/i1_5 ), .A2(
        \SB1_3_16/i0[8] ), .A3(\SB1_3_16/i3[0] ), .ZN(
        \SB1_3_16/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U5509 ( .A1(\SB1_3_2/i0[8] ), .A2(\SB1_3_2/i1_5 ), .A3(
        \SB1_3_2/i3[0] ), .ZN(n1658) );
  NAND3_X1 \SB1_3_7/Component_Function_1/N4  ( .A1(\SB1_3_7/i1_7 ), .A2(
        \SB1_3_7/i0[8] ), .A3(\SB1_3_7/i0_4 ), .ZN(
        \SB1_3_7/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U2137 ( .A1(\SB1_3_22/i0_0 ), .A2(\SB1_3_22/i3[0] ), .A3(
        \SB1_3_22/i1_7 ), .ZN(n2118) );
  NAND3_X1 \SB1_3_28/Component_Function_0/N2  ( .A1(\SB1_3_28/i0[8] ), .A2(
        \SB1_3_28/i0[7] ), .A3(\SB1_3_28/i0[6] ), .ZN(
        \SB1_3_28/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_4/Component_Function_0/N4  ( .A1(\SB1_3_4/i0[7] ), .A2(
        \SB1_3_4/i0_3 ), .A3(\SB1_3_4/i0_0 ), .ZN(
        \SB1_3_4/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U1359 ( .A1(\SB1_3_15/i1_5 ), .A2(\SB1_3_15/i0[10] ), .A3(
        \SB1_3_15/i1[9] ), .ZN(\SB1_3_15/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_28/Component_Function_4/N4  ( .A1(\SB1_3_28/i1[9] ), .A2(
        \SB1_3_28/i1_5 ), .A3(\SB1_3_28/i0_4 ), .ZN(
        \SB1_3_28/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U771 ( .A1(\SB1_3_27/i0_0 ), .A2(\SB1_3_27/i0[7] ), .A3(
        \SB1_3_27/i0_3 ), .ZN(n2297) );
  NAND3_X1 \SB1_3_20/Component_Function_4/N4  ( .A1(\SB1_3_20/i1[9] ), .A2(
        \SB1_3_20/i1_5 ), .A3(\SB1_3_20/i0_4 ), .ZN(
        \SB1_3_20/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_1/Component_Function_1/N3  ( .A1(\SB1_3_1/i1_5 ), .A2(
        \SB1_3_1/i0[6] ), .A3(\SB1_3_1/i0[9] ), .ZN(
        \SB1_3_1/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_13/Component_Function_2/N4  ( .A1(\SB1_3_13/i1_5 ), .A2(
        \SB1_3_13/i0_0 ), .A3(\SB1_3_13/i0_4 ), .ZN(
        \SB1_3_13/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U770 ( .A1(\SB1_3_10/i0[6] ), .A2(\SB1_3_10/i0_4 ), .A3(
        \SB1_3_10/i0[9] ), .ZN(n1331) );
  NAND3_X1 \SB1_3_15/Component_Function_2/N2  ( .A1(\SB1_3_15/i0_3 ), .A2(
        \SB1_3_15/i0[10] ), .A3(\SB1_3_15/i0[6] ), .ZN(
        \SB1_3_15/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_19/Component_Function_4/N4  ( .A1(\SB1_3_19/i1[9] ), .A2(
        \SB1_3_19/i1_5 ), .A3(\SB1_3_19/i0_4 ), .ZN(
        \SB1_3_19/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_22/Component_Function_2/N1  ( .A1(\SB1_3_22/i1_5 ), .A2(
        \SB1_3_22/i0[10] ), .A3(\SB1_3_22/i1[9] ), .ZN(
        \SB1_3_22/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U5974 ( .A1(\SB1_3_22/i0[10] ), .A2(\SB1_3_22/i0_3 ), .A3(
        \SB1_3_22/i0[9] ), .ZN(n1861) );
  NAND3_X1 \SB1_3_20/Component_Function_0/N3  ( .A1(\SB1_3_20/i0[10] ), .A2(
        \SB1_3_20/i0_4 ), .A3(\SB1_3_20/i0_3 ), .ZN(
        \SB1_3_20/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_22/Component_Function_4/N4  ( .A1(\SB1_3_22/i1[9] ), .A2(
        \SB1_3_22/i1_5 ), .A3(\SB1_3_22/i0_4 ), .ZN(
        \SB1_3_22/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_2/Component_Function_2/N3  ( .A1(\SB1_3_2/i0_3 ), .A2(
        \SB1_3_2/i0[8] ), .A3(\SB1_3_2/i0[9] ), .ZN(
        \SB1_3_2/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_15/Component_Function_0/N3  ( .A1(\SB1_3_15/i0[10] ), .A2(
        \SB1_3_15/i0_4 ), .A3(\SB1_3_15/i0_3 ), .ZN(
        \SB1_3_15/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_2/Component_Function_1/N4  ( .A1(\SB1_3_2/i1_7 ), .A2(
        \SB1_3_2/i0[8] ), .A3(\SB1_3_2/i0_4 ), .ZN(
        \SB1_3_2/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_23/Component_Function_5/N4  ( .A1(\SB1_3_23/i0[9] ), .A2(
        \SB1_3_23/i0[6] ), .A3(\SB1_3_23/i0_4 ), .ZN(
        \SB1_3_23/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 U750 ( .A1(n905), .A2(n886), .ZN(n2241) );
  NAND3_X1 \SB1_3_28/Component_Function_3/N2  ( .A1(\SB1_3_28/i0_0 ), .A2(
        \SB1_3_28/i0_3 ), .A3(\SB1_3_28/i0_4 ), .ZN(
        \SB1_3_28/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_2/Component_Function_4/N1  ( .A1(\SB1_3_2/i0[9] ), .A2(
        \SB1_3_2/i0_0 ), .A3(\SB1_3_2/i0[8] ), .ZN(
        \SB1_3_2/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U5745 ( .A1(\SB1_3_25/i0[6] ), .A2(\SB1_3_25/i0_4 ), .A3(
        \SB1_3_25/i0[9] ), .ZN(n1761) );
  NAND2_X1 U1693 ( .A1(\SB1_3_25/i0_3 ), .A2(\SB1_3_25/i1[9] ), .ZN(
        \SB1_3_25/Component_Function_1/NAND4_in[0] ) );
  INV_X2 U731 ( .I(\SB2_3_26/i0[7] ), .ZN(\SB2_3_26/i0_4 ) );
  INV_X1 \SB2_3_6/INV_1  ( .I(\SB1_3_10/buf_output[1] ), .ZN(\SB2_3_6/i1_7 )
         );
  NAND3_X1 \SB2_3_13/Component_Function_3/N2  ( .A1(\SB2_3_13/i0_0 ), .A2(
        \SB2_3_13/i0_3 ), .A3(\SB1_3_14/buf_output[4] ), .ZN(
        \SB2_3_13/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_28/Component_Function_3/N3  ( .A1(n2911), .A2(
        \SB2_3_28/i1_7 ), .A3(\SB1_3_30/buf_output[3] ), .ZN(
        \SB2_3_28/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_26/Component_Function_1/N2  ( .A1(\SB2_3_26/i0_3 ), .A2(
        \SB2_3_26/i1_7 ), .A3(n4750), .ZN(
        \SB2_3_26/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_23/Component_Function_4/N2  ( .A1(\SB2_3_23/i3[0] ), .A2(
        \SB2_3_23/i0_0 ), .A3(\SB2_3_23/i1_7 ), .ZN(
        \SB2_3_23/Component_Function_4/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_28/Component_Function_5/N1  ( .A1(\SB2_3_28/i0_0 ), .A2(
        \SB2_3_28/i3[0] ), .ZN(\SB2_3_28/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_1/Component_Function_4/N4  ( .A1(\SB2_3_1/i1[9] ), .A2(
        \SB2_3_1/i1_5 ), .A3(\SB2_3_1/i0_4 ), .ZN(
        \SB2_3_1/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U3267 ( .A1(\SB2_3_18/i0_3 ), .A2(\SB2_3_18/i0[9] ), .A3(
        \SB2_3_18/i0[10] ), .ZN(\SB2_3_18/Component_Function_4/NAND4_in[2] )
         );
  INV_X2 \SB2_3_8/INV_4  ( .I(\SB1_3_9/buf_output[4] ), .ZN(\SB2_3_8/i0[7] )
         );
  INV_X1 \SB2_3_5/INV_1  ( .I(\SB1_3_9/buf_output[1] ), .ZN(\SB2_3_5/i1_7 ) );
  INV_X1 \SB2_3_17/INV_4  ( .I(\SB1_3_18/buf_output[4] ), .ZN(\SB2_3_17/i0[7] ) );
  NAND3_X1 U2141 ( .A1(\SB2_3_26/i1_7 ), .A2(n4750), .A3(\SB2_3_26/i0_4 ), 
        .ZN(\SB2_3_26/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U2912 ( .A1(\SB2_3_25/i0[8] ), .A2(\SB2_3_25/i1_7 ), .A3(
        \SB1_3_26/buf_output[4] ), .ZN(
        \SB2_3_25/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U5861 ( .A1(\SB2_3_29/i0[8] ), .A2(\SB2_3_29/i1_5 ), .A3(
        \SB2_3_29/i3[0] ), .ZN(n1815) );
  NAND3_X1 U2152 ( .A1(\SB2_3_26/i1_5 ), .A2(n4750), .A3(\SB2_3_26/i3[0] ), 
        .ZN(\SB2_3_26/Component_Function_3/NAND4_in[3] ) );
  NAND2_X1 \SB2_3_5/Component_Function_5/N1  ( .A1(\SB2_3_5/i0_0 ), .A2(
        \SB2_3_5/i3[0] ), .ZN(\SB2_3_5/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_8/Component_Function_5/N1  ( .A1(\SB2_3_8/i0_0 ), .A2(
        \SB2_3_8/i3[0] ), .ZN(\SB2_3_8/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U683 ( .A1(\SB2_3_6/i0[10] ), .A2(\SB2_3_6/i1_7 ), .A3(
        \SB2_3_6/i1[9] ), .ZN(n2459) );
  NAND3_X1 \SB2_3_6/Component_Function_3/N1  ( .A1(\SB2_3_6/i1[9] ), .A2(
        \SB2_3_6/i0_3 ), .A3(\SB2_3_6/i0[6] ), .ZN(
        \SB2_3_6/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_27/Component_Function_2/N3  ( .A1(\SB2_3_27/i0_3 ), .A2(
        \SB2_3_27/i0[8] ), .A3(\RI3[3][24] ), .ZN(
        \SB2_3_27/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3680 ( .A1(\SB2_3_18/i0_3 ), .A2(\SB2_3_18/i0_4 ), .A3(
        \SB2_3_18/i0[10] ), .ZN(n1082) );
  NAND3_X1 U4547 ( .A1(\SB2_3_17/i0_3 ), .A2(\SB2_3_17/i1_7 ), .A3(
        \SB2_3_17/i0[8] ), .ZN(\SB2_3_17/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_12/Component_Function_0/N4  ( .A1(\SB2_3_12/i0[7] ), .A2(
        \SB2_3_12/i0_3 ), .A3(\SB2_3_12/i0_0 ), .ZN(
        \SB2_3_12/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U684 ( .A1(\SB2_3_14/i0_0 ), .A2(\SB2_3_14/i0[7] ), .A3(
        \SB2_3_14/i0_3 ), .ZN(\SB2_3_14/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_17/Component_Function_4/N1  ( .A1(\SB2_3_17/i0[9] ), .A2(
        \SB2_3_17/i0_0 ), .A3(\SB2_3_17/i0[8] ), .ZN(
        \SB2_3_17/Component_Function_4/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_19/Component_Function_0/N1  ( .A1(\SB2_3_19/i0[10] ), .A2(
        \SB2_3_19/i0[9] ), .ZN(\SB2_3_19/Component_Function_0/NAND4_in[0] ) );
  INV_X1 \SB3_23/INV_1  ( .I(\MC_ARK_ARC_1_3/buf_output[49] ), .ZN(
        \SB3_23/i1_7 ) );
  BUF_X2 \SB3_28/BUF_0  ( .I(\MC_ARK_ARC_1_3/buf_output[18] ), .Z(
        \SB3_28/i0[9] ) );
  BUF_X2 U1804 ( .I(\MC_ARK_ARC_1_3/buf_output[72] ), .Z(\SB3_19/i0[9] ) );
  BUF_X4 \SB3_13/BUF_5  ( .I(\MC_ARK_ARC_1_3/buf_output[113] ), .Z(
        \SB3_13/i0_3 ) );
  BUF_X2 \SB3_15/BUF_0  ( .I(\MC_ARK_ARC_1_3/buf_output[96] ), .Z(
        \SB3_15/i0[9] ) );
  NAND3_X1 \SB3_13/Component_Function_1/N4  ( .A1(\SB3_13/i1_7 ), .A2(
        \SB3_13/i0[8] ), .A3(\SB3_13/i0_4 ), .ZN(
        \SB3_13/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_18/Component_Function_0/N2  ( .A1(\SB3_18/i0[8] ), .A2(
        \SB3_18/i0[7] ), .A3(\SB3_18/i0[6] ), .ZN(
        \SB3_18/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U5909 ( .A1(\SB3_7/i0[8] ), .A2(\SB3_7/i3[0] ), .A3(n4766), .ZN(
        n1836) );
  NAND3_X1 \SB3_28/Component_Function_5/N3  ( .A1(\SB3_28/i1[9] ), .A2(
        \SB3_28/i0_4 ), .A3(\SB3_28/i0_3 ), .ZN(
        \SB3_28/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB3_24/Component_Function_1/N3  ( .A1(\SB3_24/i1_5 ), .A2(
        \SB3_24/i0[6] ), .A3(\SB3_24/i0[9] ), .ZN(
        \SB3_24/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_21/Component_Function_4/N1  ( .A1(\SB3_21/i0[9] ), .A2(
        \SB3_21/i0_0 ), .A3(\SB3_21/i0[8] ), .ZN(
        \SB3_21/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U1179 ( .A1(\SB3_19/i1[9] ), .A2(\SB3_19/i0_3 ), .A3(\SB3_19/i0[6] ), .ZN(\SB3_19/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U7515 ( .A1(\MC_ARK_ARC_1_3/buf_output[46] ), .A2(\SB3_24/i1[9] ), 
        .A3(\SB3_24/i1_5 ), .ZN(n2633) );
  NAND3_X1 U1654 ( .A1(\SB3_17/i0[9] ), .A2(\SB3_17/i0[10] ), .A3(
        \SB3_17/i0_3 ), .ZN(\SB3_17/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB3_28/Component_Function_2/N2  ( .A1(\SB3_28/i0_3 ), .A2(
        \SB3_28/i0[10] ), .A3(\SB3_28/i0[6] ), .ZN(
        \SB3_28/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U608 ( .A1(\SB3_21/i0_3 ), .A2(\SB3_21/i1[9] ), .A3(\SB3_21/i0[6] ), 
        .ZN(\SB3_21/Component_Function_3/NAND4_in[0] ) );
  NAND4_X2 U3674 ( .A1(\SB3_13/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_13/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_13/Component_Function_2/NAND4_in[3] ), .A4(n1079), .ZN(
        \SB3_13/buf_output[2] ) );
  BUF_X2 \SB4_5/BUF_0  ( .I(\SB3_10/buf_output[0] ), .Z(\SB4_5/i0[9] ) );
  BUF_X2 \SB4_26/BUF_0  ( .I(\SB3_31/buf_output[0] ), .Z(\SB4_26/i0[9] ) );
  INV_X1 \SB4_24/INV_5  ( .I(\SB3_24/buf_output[5] ), .ZN(\SB4_24/i1_5 ) );
  NAND3_X1 \SB4_25/Component_Function_5/N3  ( .A1(\SB4_25/i1[9] ), .A2(
        \SB4_25/i0_4 ), .A3(\SB4_25/i0_3 ), .ZN(
        \SB4_25/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB4_18/Component_Function_3/N2  ( .A1(\SB4_18/i0_0 ), .A2(
        \SB4_18/i0_3 ), .A3(\SB4_18/i0_4 ), .ZN(
        \SB4_18/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3104 ( .A1(\SB4_19/i0_3 ), .A2(\SB3_23/buf_output[1] ), .A3(
        \SB4_19/i1[9] ), .ZN(n870) );
  NAND3_X1 \SB4_16/Component_Function_1/N4  ( .A1(\SB4_16/i1_7 ), .A2(
        \SB4_16/i0[8] ), .A3(\SB4_16/i0_4 ), .ZN(
        \SB4_16/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB4_7/Component_Function_1/N1  ( .A1(\SB4_7/i0_3 ), .A2(
        \SB4_7/i1[9] ), .ZN(\SB4_7/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB4_18/Component_Function_0/N1  ( .A1(\SB4_18/i0[10] ), .A2(
        \SB4_18/i0[9] ), .ZN(\SB4_18/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U43 ( .A1(\SB4_13/i1_5 ), .A2(\SB4_13/i0[6] ), .A3(\SB4_13/i0[9] ), 
        .ZN(\SB4_13/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U155 ( .A1(\SB4_20/i0[6] ), .A2(\SB4_20/i0[8] ), .A3(\SB4_20/i0[7] ), .ZN(\SB4_20/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U371 ( .A1(\SB4_13/i1_5 ), .A2(\SB4_13/i0[10] ), .A3(\SB4_13/i1[9] ), .ZN(\SB4_13/Component_Function_2/NAND4_in[0] ) );
  CLKBUF_X2 U586 ( .I(\SB3_30/buf_output[2] ), .Z(n2898) );
  NAND3_X1 U599 ( .A1(\SB3_20/i0_3 ), .A2(\SB3_20/i0[6] ), .A3(\SB3_20/i1[9] ), 
        .ZN(n3864) );
  NAND3_X1 U600 ( .A1(\SB3_21/i1_5 ), .A2(\SB3_21/i0[8] ), .A3(\SB3_21/i3[0] ), 
        .ZN(n4217) );
  NAND3_X1 U615 ( .A1(\SB3_19/i0[10] ), .A2(\SB3_19/i0_3 ), .A3(\SB3_19/i0[6] ), .ZN(n4065) );
  NAND3_X1 U620 ( .A1(\SB3_10/i0[6] ), .A2(\SB3_10/i1[9] ), .A3(\SB3_10/i0_3 ), 
        .ZN(n4571) );
  NAND3_X1 U623 ( .A1(\SB3_2/i0[10] ), .A2(\SB3_2/i0_3 ), .A3(\SB3_2/i0[9] ), 
        .ZN(n3481) );
  NAND3_X1 U624 ( .A1(\SB3_29/i0_4 ), .A2(\SB3_29/i0[9] ), .A3(\SB3_29/i0[6] ), 
        .ZN(n3406) );
  NAND3_X1 U626 ( .A1(n4766), .A2(\SB3_7/i0[6] ), .A3(\SB3_7/i0[9] ), .ZN(
        \SB3_7/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U628 ( .A1(\SB3_30/i0[9] ), .A2(n5488), .A3(\SB3_30/i0[8] ), .ZN(
        n3891) );
  NAND3_X1 U635 ( .A1(\SB3_30/i0_0 ), .A2(\SB3_30/i1_7 ), .A3(\SB3_30/i3[0] ), 
        .ZN(\SB3_30/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U662 ( .A1(\SB2_3_5/i0_0 ), .A2(\SB1_3_6/buf_output[4] ), .A3(
        \SB2_3_5/i1_5 ), .ZN(n4126) );
  NAND3_X1 U674 ( .A1(\SB2_3_6/i0_4 ), .A2(\SB2_3_6/i1_7 ), .A3(
        \SB2_3_6/i0[8] ), .ZN(n4083) );
  NAND3_X1 U688 ( .A1(\SB2_3_7/i0[8] ), .A2(n3739), .A3(n1670), .ZN(
        \SB2_3_7/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U689 ( .A1(\SB2_3_16/i0[9] ), .A2(\SB2_3_16/i1_5 ), .A3(
        \SB2_3_16/i0[6] ), .ZN(\SB2_3_16/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U691 ( .A1(\SB2_3_9/i0_4 ), .A2(\SB2_3_9/i1[9] ), .A3(
        \SB2_3_9/i1_5 ), .ZN(n4637) );
  NAND3_X1 U715 ( .A1(\SB2_3_31/i0_3 ), .A2(\SB2_3_31/i0[10] ), .A3(
        \SB2_3_31/i0[9] ), .ZN(\SB2_3_31/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U722 ( .A1(\SB2_3_16/i0[9] ), .A2(\SB2_3_16/i0[6] ), .A3(
        \SB1_3_17/buf_output[4] ), .ZN(n4681) );
  NAND3_X1 U737 ( .A1(\SB2_3_30/i0_0 ), .A2(\SB2_3_30/i0[10] ), .A3(
        \SB2_3_30/i0[6] ), .ZN(\SB2_3_30/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U739 ( .A1(\SB2_3_22/i0[6] ), .A2(\SB2_3_22/i1_5 ), .A3(
        \SB2_3_22/i0[9] ), .ZN(\SB2_3_22/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U740 ( .A1(\SB2_3_20/i0_3 ), .A2(\SB2_3_20/i0[9] ), .A3(
        \SB2_3_20/i0[8] ), .ZN(\SB2_3_20/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U746 ( .A1(\SB2_3_28/i0_3 ), .A2(n2911), .A3(n577), .ZN(
        \SB2_3_28/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U748 ( .A1(\SB2_3_22/i0_3 ), .A2(\SB2_3_22/i0[10] ), .A3(
        \SB2_3_22/i0[9] ), .ZN(n2076) );
  NAND3_X1 U785 ( .A1(\SB1_3_28/i0[9] ), .A2(\SB1_3_28/i0_3 ), .A3(
        \SB1_3_28/i0[10] ), .ZN(n4199) );
  NAND3_X1 U787 ( .A1(\SB1_3_22/i0_0 ), .A2(\SB1_3_22/i0[9] ), .A3(
        \SB1_3_22/i0[8] ), .ZN(n3075) );
  NAND3_X1 U788 ( .A1(\SB1_3_13/i0[6] ), .A2(\SB1_3_13/i0[9] ), .A3(
        \SB1_3_13/i0_4 ), .ZN(n4544) );
  NAND3_X1 U791 ( .A1(\SB1_3_28/i0_3 ), .A2(\SB1_3_28/i0_0 ), .A3(
        \SB1_3_28/i0[7] ), .ZN(n3610) );
  NAND3_X1 U792 ( .A1(\SB1_3_29/i0[9] ), .A2(\SB1_3_29/i1_5 ), .A3(
        \SB1_3_29/i0[6] ), .ZN(n1971) );
  NAND3_X1 U793 ( .A1(\SB1_3_30/i0_4 ), .A2(\SB1_3_30/i0_0 ), .A3(
        \SB1_3_30/i1_5 ), .ZN(n3297) );
  NAND3_X1 U811 ( .A1(\SB1_3_2/i0[8] ), .A2(\SB1_3_2/i0_3 ), .A3(
        \SB1_3_2/i1_7 ), .ZN(\SB1_3_2/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U822 ( .A1(\SB1_3_20/i0_3 ), .A2(\SB1_3_20/i1[9] ), .A3(
        \SB1_3_20/i0_4 ), .ZN(n4328) );
  NAND3_X1 U853 ( .A1(\SB1_3_1/i0[6] ), .A2(\SB1_3_1/i0_4 ), .A3(
        \SB1_3_1/i0[9] ), .ZN(n4120) );
  NAND3_X1 U861 ( .A1(\SB1_3_27/i0_3 ), .A2(\SB1_3_27/i0[8] ), .A3(
        \MC_ARK_ARC_1_2/buf_output[24] ), .ZN(n3822) );
  NAND3_X1 U882 ( .A1(\SB1_3_26/i0_4 ), .A2(\SB1_3_26/i0[8] ), .A3(
        \SB1_3_26/i1_7 ), .ZN(n2749) );
  NAND3_X1 U887 ( .A1(\SB1_3_10/i0[8] ), .A2(\SB1_3_10/i1_7 ), .A3(
        \SB1_3_10/i0_4 ), .ZN(n4583) );
  NAND3_X1 U893 ( .A1(\SB1_3_19/i0[8] ), .A2(\SB1_3_19/i3[0] ), .A3(
        \SB1_3_19/i1_5 ), .ZN(n820) );
  NAND3_X1 U894 ( .A1(\SB1_3_27/i0[8] ), .A2(\SB1_3_27/i1_5 ), .A3(
        \SB1_3_27/i3[0] ), .ZN(n4383) );
  NAND3_X1 U915 ( .A1(\SB1_3_21/i0_3 ), .A2(\SB1_3_21/i0[8] ), .A3(
        \SB1_3_21/i0[9] ), .ZN(\SB1_3_21/Component_Function_2/NAND4_in[2] ) );
  BUF_X2 U920 ( .I(\MC_ARK_ARC_1_2/buf_output[108] ), .Z(\SB1_3_13/i0[9] ) );
  NAND3_X1 U941 ( .A1(\SB1_3_1/i0_0 ), .A2(\SB1_3_1/i1_7 ), .A3(
        \SB1_3_1/i3[0] ), .ZN(n4525) );
  NAND3_X1 U945 ( .A1(\SB1_3_29/i1[9] ), .A2(\SB1_3_29/i1_5 ), .A3(
        \SB1_3_29/i0_4 ), .ZN(n953) );
  BUF_X4 U954 ( .I(n6540), .Z(\SB1_3_29/i0_3 ) );
  OAI21_X1 U957 ( .A1(\SB2_2_12/i0_3 ), .A2(\SB2_2_12/i0_4 ), .B(n2901), .ZN(
        n1488) );
  NAND3_X1 U972 ( .A1(\SB1_2_19/buf_output[4] ), .A2(\SB2_2_18/i0[8] ), .A3(
        \SB2_2_18/i1_7 ), .ZN(n4009) );
  NAND3_X1 U979 ( .A1(\SB2_2_27/i0_0 ), .A2(\SB2_2_27/i1_5 ), .A3(
        \SB1_2_28/buf_output[4] ), .ZN(n3198) );
  NAND3_X1 U1001 ( .A1(\SB2_2_28/i0_4 ), .A2(\SB2_2_28/i0[8] ), .A3(
        \SB2_2_28/i1_7 ), .ZN(\SB2_2_28/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U1047 ( .A1(\SB2_2_7/i0[10] ), .A2(\SB2_2_7/i1_7 ), .A3(
        \SB2_2_7/i1[9] ), .ZN(\SB2_2_7/Component_Function_3/NAND4_in[2] ) );
  INV_X1 U1091 ( .I(\SB1_2_6/buf_output[1] ), .ZN(\SB2_2_2/i1_7 ) );
  NAND3_X1 U1105 ( .A1(\SB1_2_1/i0[8] ), .A2(\SB1_2_1/i0[9] ), .A3(
        \SB1_2_1/i0_3 ), .ZN(\SB1_2_1/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1135 ( .A1(\MC_ARK_ARC_1_1/buf_output[130] ), .A2(\SB1_2_10/i0_3 ), 
        .A3(\SB1_2_10/i1[9] ), .ZN(n3591) );
  NAND3_X1 U1141 ( .A1(\SB1_2_21/i0_3 ), .A2(\SB1_2_21/i0[7] ), .A3(
        \SB1_2_21/i0_0 ), .ZN(n4026) );
  NAND3_X1 U1166 ( .A1(\MC_ARK_ARC_1_1/buf_output[70] ), .A2(\SB1_2_20/i0[9] ), 
        .A3(\SB1_2_20/i0[6] ), .ZN(n3338) );
  NAND3_X1 U1180 ( .A1(\RI1[2][35] ), .A2(\SB1_2_26/i1[9] ), .A3(
        \SB1_2_26/i0[6] ), .ZN(\SB1_2_26/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U1187 ( .A1(\SB1_2_29/i0_4 ), .A2(\SB1_2_29/i0_0 ), .A3(
        \RI1[2][17] ), .ZN(n4071) );
  NAND3_X1 U1198 ( .A1(\SB1_2_25/i0_0 ), .A2(\SB1_2_25/i1_5 ), .A3(
        \MC_ARK_ARC_1_1/buf_output[40] ), .ZN(n4444) );
  NAND3_X1 U1203 ( .A1(\SB1_2_15/i0[6] ), .A2(\SB1_2_15/i1_5 ), .A3(
        \SB1_2_15/i0[9] ), .ZN(\SB1_2_15/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1223 ( .A1(\SB1_2_28/i0[8] ), .A2(\SB1_2_28/i3[0] ), .A3(
        \SB1_2_28/i1_5 ), .ZN(\SB1_2_28/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U1224 ( .A1(\SB1_2_11/i0_0 ), .A2(\SB1_2_11/i0_3 ), .A3(
        \SB1_2_11/i0[7] ), .ZN(n4363) );
  NAND3_X1 U1225 ( .A1(\SB1_2_31/i0[10] ), .A2(\SB1_2_31/i1[9] ), .A3(
        \SB1_2_31/i1_7 ), .ZN(\SB1_2_31/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U1226 ( .A1(\SB1_2_2/i0[8] ), .A2(\SB1_2_2/i0_4 ), .A3(
        \SB1_2_2/i1_7 ), .ZN(n4670) );
  NAND3_X1 U1240 ( .A1(\SB1_2_19/i0_0 ), .A2(\SB1_2_19/i0[9] ), .A3(
        \SB1_2_19/i0[8] ), .ZN(\SB1_2_19/Component_Function_4/NAND4_in[0] ) );
  INV_X4 U1248 ( .I(\RI1[2][47] ), .ZN(\SB1_2_24/i1_5 ) );
  NAND3_X1 U1252 ( .A1(\SB2_1_27/i0[9] ), .A2(\SB2_1_27/i1_5 ), .A3(
        \SB2_1_27/i0[6] ), .ZN(\SB2_1_27/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1293 ( .A1(\SB2_1_19/i0[8] ), .A2(n578), .A3(\SB2_1_19/i1_7 ), 
        .ZN(\SB2_1_19/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U1295 ( .A1(n3690), .A2(\SB2_1_30/i0_4 ), .A3(\SB2_1_30/i0_3 ), 
        .ZN(\SB2_1_30/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U1300 ( .A1(\SB1_1_9/buf_output[4] ), .A2(\SB2_1_8/i1_7 ), .A3(
        \SB2_1_8/i0[8] ), .ZN(n3938) );
  NAND3_X1 U1304 ( .A1(\SB2_1_20/i0_0 ), .A2(\SB2_1_20/i0_3 ), .A3(
        \SB2_1_20/i0[7] ), .ZN(\SB2_1_20/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U1312 ( .A1(\SB2_1_9/i0[6] ), .A2(\SB2_1_9/i0[8] ), .A3(
        \SB2_1_9/i0[7] ), .ZN(\SB2_1_9/Component_Function_0/NAND4_in[1] ) );
  INV_X1 U1372 ( .I(\SB1_1_28/buf_output[1] ), .ZN(\SB2_1_24/i1_7 ) );
  INV_X1 U1383 ( .I(\SB1_1_9/buf_output[0] ), .ZN(\SB2_1_4/i3[0] ) );
  NAND3_X1 U1399 ( .A1(\SB1_1_2/i0_0 ), .A2(\SB1_1_2/i0_4 ), .A3(
        \SB1_1_2/i0_3 ), .ZN(\SB1_1_2/Component_Function_3/NAND4_in[1] ) );
  NAND2_X1 U1402 ( .A1(\SB1_1_24/i0_3 ), .A2(\SB1_1_24/i1[9] ), .ZN(n3385) );
  NAND3_X1 U1408 ( .A1(\MC_ARK_ARC_1_0/buf_output[76] ), .A2(\SB1_1_19/i1_7 ), 
        .A3(\SB1_1_19/i0[8] ), .ZN(\SB1_1_19/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U1412 ( .A1(\SB1_1_21/i0_4 ), .A2(\SB1_1_21/i1[9] ), .A3(
        \SB1_1_21/i1_5 ), .ZN(\SB1_1_21/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U1414 ( .A1(\SB1_1_27/i0[8] ), .A2(\SB1_1_27/i0_0 ), .A3(
        \SB1_1_27/i0[9] ), .ZN(\SB1_1_27/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U1437 ( .A1(\SB1_1_10/i0_3 ), .A2(\SB1_1_10/i0_0 ), .A3(
        \SB1_1_10/i0[7] ), .ZN(n4261) );
  NAND3_X1 U1438 ( .A1(\SB1_1_12/i0[9] ), .A2(\SB1_1_12/i0[8] ), .A3(
        \SB1_1_12/i0_0 ), .ZN(n4700) );
  NAND3_X1 U1461 ( .A1(\SB1_1_21/i0_0 ), .A2(\SB1_1_21/i0_4 ), .A3(
        \SB1_1_21/i1_5 ), .ZN(\SB1_1_21/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U1471 ( .A1(\RI1[1][59] ), .A2(\SB1_1_22/i0_0 ), .A3(
        \SB1_1_22/i0[7] ), .ZN(\SB1_1_22/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U1473 ( .A1(\SB1_1_29/i0_3 ), .A2(\SB1_1_29/i0_4 ), .A3(
        \SB1_1_29/i1[9] ), .ZN(\SB1_1_29/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1476 ( .A1(\SB1_1_19/i0_3 ), .A2(\SB1_1_19/i0[9] ), .A3(
        \SB1_1_19/i0[8] ), .ZN(n4101) );
  NAND3_X1 U1477 ( .A1(\SB1_1_13/i0[6] ), .A2(\SB1_1_13/i0[9] ), .A3(
        \SB1_1_13/i1_5 ), .ZN(\SB1_1_13/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 U1478 ( .A1(\SB1_1_22/Component_Function_2/NAND4_in[3] ), .A2(n1493), .ZN(n4174) );
  NAND3_X1 U1484 ( .A1(\SB1_1_21/i0_4 ), .A2(\SB1_1_21/i0[10] ), .A3(
        \SB1_1_21/i0_3 ), .ZN(n4611) );
  NAND3_X1 U1491 ( .A1(\SB1_1_6/i0[10] ), .A2(\SB1_1_6/i1[9] ), .A3(
        \SB1_1_6/i1_7 ), .ZN(n4293) );
  NAND3_X1 U1501 ( .A1(\SB1_1_2/i0[8] ), .A2(\SB1_1_2/i0_4 ), .A3(
        \SB1_1_2/i1_7 ), .ZN(n4138) );
  NAND3_X1 U1502 ( .A1(\SB1_1_26/i0[10] ), .A2(\SB1_1_26/i0_3 ), .A3(
        \SB1_1_26/i0[6] ), .ZN(n4284) );
  NAND3_X1 U1522 ( .A1(\SB2_0_17/i0_3 ), .A2(\SB2_0_17/i0[10] ), .A3(
        \RI3[0][88] ), .ZN(\SB2_0_17/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U1551 ( .A1(\SB2_0_26/i0[10] ), .A2(\SB2_0_26/i0_3 ), .A3(
        \RI3[0][34] ), .ZN(\SB2_0_26/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U1555 ( .A1(\SB2_0_26/i0_3 ), .A2(\SB2_0_26/i1[9] ), .A3(
        \RI3[0][34] ), .ZN(n2015) );
  NAND3_X1 U1556 ( .A1(\RI3[0][4] ), .A2(\SB2_0_31/i1[9] ), .A3(
        \SB2_0_31/i1_5 ), .ZN(n1297) );
  NAND3_X1 U1571 ( .A1(\SB2_0_12/i0[9] ), .A2(\SB2_0_12/i0[8] ), .A3(
        \SB2_0_12/i0_0 ), .ZN(\SB2_0_12/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U1582 ( .A1(\SB2_0_0/i0[10] ), .A2(\SB2_0_0/i1_7 ), .A3(
        \SB2_0_0/i1[9] ), .ZN(n4130) );
  NAND3_X1 U1599 ( .A1(\SB2_0_17/i0_3 ), .A2(\SB2_0_17/i0[10] ), .A3(
        \SB2_0_17/i0[9] ), .ZN(n2190) );
  NAND3_X1 U1616 ( .A1(\RI3[0][58] ), .A2(\RI3[0][55] ), .A3(\RI3[0][54] ), 
        .ZN(n3855) );
  NAND2_X1 U1617 ( .A1(\SB1_0_23/i0[10] ), .A2(\SB1_0_23/i0[9] ), .ZN(
        \SB1_0_23/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U1624 ( .A1(n6314), .A2(\SB1_0_28/i0[6] ), .A3(\SB1_0_28/i0[9] ), 
        .ZN(\SB1_0_28/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 U1626 ( .A1(\SB1_0_8/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_0_8/Component_Function_4/NAND4_in[0] ), .ZN(n3147) );
  NAND3_X1 U1641 ( .A1(\SB1_0_10/i1_5 ), .A2(\SB1_0_10/i0[10] ), .A3(
        \SB1_0_10/i1[9] ), .ZN(\SB1_0_10/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U1649 ( .A1(\SB1_0_2/i0_0 ), .A2(\SB1_0_2/i0[9] ), .A3(
        \SB1_0_2/i0[8] ), .ZN(n2482) );
  NAND2_X1 U1661 ( .A1(\SB1_0_27/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_0_27/Component_Function_3/NAND4_in[3] ), .ZN(n4395) );
  NAND2_X1 U1665 ( .A1(n1769), .A2(n4244), .ZN(n4243) );
  NAND3_X1 U1676 ( .A1(n390), .A2(\SB1_0_7/i1_5 ), .A3(\SB1_0_7/i1[9] ), .ZN(
        n3621) );
  NAND3_X1 U1678 ( .A1(\SB1_0_16/i0[9] ), .A2(n4752), .A3(\SB1_0_16/i0[6] ), 
        .ZN(n4315) );
  NAND3_X1 U1683 ( .A1(\SB1_0_16/i3[0] ), .A2(\SB1_0_16/i1_5 ), .A3(
        \SB1_0_16/i0[8] ), .ZN(n4539) );
  NAND3_X1 U1690 ( .A1(\SB1_0_1/i0[8] ), .A2(\SB1_0_1/i1_5 ), .A3(
        \SB1_0_1/i3[0] ), .ZN(n3419) );
  INV_X1 U1702 ( .I(n290), .ZN(\SB1_0_16/i3[0] ) );
  NAND3_X1 U1703 ( .A1(\SB1_0_25/i0[8] ), .A2(\SB1_0_25/i1_5 ), .A3(
        \SB1_0_25/i3[0] ), .ZN(n3313) );
  NAND3_X1 U1705 ( .A1(\SB1_0_27/i1_5 ), .A2(\SB1_0_27/i3[0] ), .A3(
        \SB1_0_27/i0[8] ), .ZN(\SB1_0_27/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U1706 ( .A1(\SB1_0_12/i0[10] ), .A2(\SB1_0_12/i0_3 ), .A3(
        \SB1_0_12/i0[9] ), .ZN(n3801) );
  NAND3_X1 U1707 ( .A1(\SB1_0_11/i0_3 ), .A2(\SB1_0_11/i0_4 ), .A3(
        \SB1_0_11/i0_0 ), .ZN(\SB1_0_11/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1708 ( .A1(\SB1_0_26/i0[10] ), .A2(\SB1_0_26/i1[9] ), .A3(
        \SB1_0_26/i1_5 ), .ZN(n3463) );
  BUF_X2 U1709 ( .I(n290), .Z(\SB1_0_16/i0[9] ) );
  NAND3_X2 U1725 ( .A1(\SB1_3_13/i0[6] ), .A2(\SB1_3_13/i0_3 ), .A3(
        \SB1_3_13/i1[9] ), .ZN(\SB1_3_13/Component_Function_3/NAND4_in[0] ) );
  INV_X2 U1730 ( .I(\MC_ARK_ARC_1_3/buf_output[74] ), .ZN(\SB3_19/i1[9] ) );
  BUF_X2 U1735 ( .I(\SB2_2_30/buf_output[2] ), .Z(\RI5[2][26] ) );
  BUF_X4 U1753 ( .I(n420), .Z(\SB1_0_16/i0_3 ) );
  NAND3_X2 U1757 ( .A1(\SB1_2_22/i0_3 ), .A2(\SB1_2_22/i1[9] ), .A3(
        \SB1_2_22/i0_4 ), .ZN(\SB1_2_22/Component_Function_5/NAND4_in[2] ) );
  INV_X2 U1766 ( .I(n420), .ZN(\SB1_0_16/i1_5 ) );
  BUF_X4 U1776 ( .I(n413), .Z(\SB1_0_23/i0_3 ) );
  NAND3_X2 U1778 ( .A1(\SB1_0_5/i0[10] ), .A2(\SB1_0_5/i1_7 ), .A3(
        \SB1_0_5/i1[9] ), .ZN(n3627) );
  INV_X4 U1785 ( .I(\SB2_2_1/i0[7] ), .ZN(\SB2_2_1/i0_4 ) );
  INV_X2 U1788 ( .I(n5498), .ZN(\SB1_0_25/i1_5 ) );
  NAND3_X2 U1794 ( .A1(\SB2_2_20/i1_5 ), .A2(\SB2_2_20/i0[10] ), .A3(
        \SB2_2_20/i1[9] ), .ZN(\SB2_2_20/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U1803 ( .A1(\SB2_2_6/i0_3 ), .A2(n2074), .A3(\SB2_2_6/i1[9] ), .ZN(
        n4429) );
  INV_X2 U1816 ( .I(\MC_ARK_ARC_1_2/buf_output[35] ), .ZN(\SB1_3_26/i1_5 ) );
  NAND3_X2 U1819 ( .A1(\SB2_2_6/i0[10] ), .A2(\SB2_2_6/i1_5 ), .A3(
        \SB2_2_6/i1[9] ), .ZN(n4705) );
  BUF_X2 U1820 ( .I(n309), .Z(\SB1_0_10/i0[6] ) );
  BUF_X4 U1828 ( .I(\SB1_1_27/buf_output[5] ), .Z(\SB2_1_27/i0_3 ) );
  NAND3_X2 U1832 ( .A1(\SB3_7/i0[10] ), .A2(\SB3_7/i0[6] ), .A3(\SB3_7/i0_0 ), 
        .ZN(n3445) );
  BUF_X4 U1834 ( .I(\MC_ARK_ARC_1_2/buf_output[2] ), .Z(\SB1_3_31/i0_0 ) );
  INV_X2 U1837 ( .I(\SB1_1_27/buf_output[5] ), .ZN(\SB2_1_27/i1_5 ) );
  NAND3_X1 U1883 ( .A1(\SB2_3_2/i1[9] ), .A2(\SB2_3_2/i0_3 ), .A3(
        \SB2_3_2/i0[6] ), .ZN(\SB2_3_2/Component_Function_3/NAND4_in[0] ) );
  NAND2_X1 U1898 ( .A1(\SB2_2_28/i0_0 ), .A2(\SB2_2_28/i3[0] ), .ZN(
        \SB2_2_28/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U1954 ( .A1(\SB2_3_29/i0[7] ), .A2(\SB2_3_29/i0_3 ), .A3(
        \SB2_3_29/i0_0 ), .ZN(n659) );
  NAND3_X1 U1970 ( .A1(\SB2_3_4/i0_4 ), .A2(\SB2_3_4/i1_7 ), .A3(
        \SB2_3_4/i0[8] ), .ZN(n1484) );
  NAND3_X1 U1988 ( .A1(\SB4_21/i3[0] ), .A2(\SB3_24/buf_output[2] ), .A3(
        \SB4_21/i1_7 ), .ZN(\SB4_21/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U2016 ( .A1(\SB2_3_9/i0_3 ), .A2(\SB1_3_10/buf_output[4] ), .A3(
        \SB2_3_9/i1[9] ), .ZN(n3509) );
  NAND3_X1 U2036 ( .A1(\SB2_3_26/i0_3 ), .A2(\SB2_3_26/i0_4 ), .A3(
        \SB2_3_26/i1[9] ), .ZN(n2050) );
  NAND3_X1 U2037 ( .A1(\SB2_3_26/i1_5 ), .A2(\SB1_3_28/buf_output[3] ), .A3(
        \SB2_3_26/i1[9] ), .ZN(\SB2_3_26/Component_Function_2/NAND4_in[0] ) );
  BUF_X2 U2043 ( .I(\MC_ARK_ARC_1_3/buf_output[141] ), .Z(\SB3_8/i0[10] ) );
  INV_X1 U2047 ( .I(\MC_ARK_ARC_1_3/buf_output[141] ), .ZN(\SB3_8/i0[8] ) );
  NAND3_X1 U2061 ( .A1(\SB2_3_25/i0_0 ), .A2(\SB2_3_25/i0[7] ), .A3(
        \SB2_3_25/i0_3 ), .ZN(n2133) );
  NAND2_X1 U2067 ( .A1(\SB3_15/i0_0 ), .A2(\SB3_15/i3[0] ), .ZN(
        \SB3_15/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U2071 ( .A1(\SB3_15/i0_3 ), .A2(\SB3_15/i0[7] ), .A3(\SB3_15/i0_0 ), 
        .ZN(n1263) );
  NAND3_X1 U2073 ( .A1(\SB4_10/i3[0] ), .A2(\SB3_13/buf_output[2] ), .A3(
        \SB4_10/i1_7 ), .ZN(\SB4_10/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U2084 ( .A1(\SB1_3_30/i0[9] ), .A2(\SB1_3_30/i0[10] ), .A3(
        \SB1_3_30/i0_3 ), .ZN(\SB1_3_30/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2092 ( .A1(\SB1_3_30/i0_3 ), .A2(\SB1_3_30/i0_4 ), .A3(
        \SB1_3_30/i1[9] ), .ZN(\SB1_3_30/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2103 ( .A1(\SB1_3_18/i0_3 ), .A2(\SB1_3_18/i0[8] ), .A3(
        \SB1_3_18/i0[9] ), .ZN(\SB1_3_18/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2104 ( .A1(\SB1_3_18/i0[8] ), .A2(\SB1_3_18/i1_5 ), .A3(
        \SB1_3_18/i3[0] ), .ZN(n3077) );
  CLKBUF_X4 U2106 ( .I(\SB3_19/buf_output[5] ), .Z(\SB4_19/i0_3 ) );
  NAND3_X1 U2124 ( .A1(\SB2_2_6/i1[9] ), .A2(\SB2_2_6/i1_5 ), .A3(n2074), .ZN(
        \SB2_2_6/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U2129 ( .A1(\SB2_2_23/i1[9] ), .A2(\SB2_2_23/i1_5 ), .A3(
        \SB2_2_23/i0_4 ), .ZN(\SB2_2_23/Component_Function_4/NAND4_in[3] ) );
  NAND2_X1 U2130 ( .A1(\SB2_2_23/i0_3 ), .A2(\SB2_2_23/i1[9] ), .ZN(
        \SB2_2_23/Component_Function_1/NAND4_in[0] ) );
  BUF_X2 U2134 ( .I(\SB3_28/buf_output[1] ), .Z(\SB4_24/i0[6] ) );
  INV_X1 U2136 ( .I(\SB3_28/buf_output[1] ), .ZN(\SB4_24/i1_7 ) );
  NAND3_X1 U2139 ( .A1(\SB4_24/i0[10] ), .A2(\SB4_24/i1[9] ), .A3(
        \SB4_24/i1_7 ), .ZN(\SB4_24/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2147 ( .A1(\SB4_24/i1_5 ), .A2(\SB4_24/i0[10] ), .A3(
        \SB4_24/i1[9] ), .ZN(\SB4_24/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U2169 ( .A1(\SB3_22/i0_0 ), .A2(\SB3_22/i0_3 ), .A3(\SB3_22/i0_4 ), 
        .ZN(\SB3_22/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2171 ( .A1(\SB3_22/i0[7] ), .A2(\SB3_22/i0_3 ), .A3(\SB3_22/i0_0 ), 
        .ZN(\SB3_22/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2177 ( .A1(\SB3_22/i0_3 ), .A2(\SB3_22/i0[10] ), .A3(
        \SB3_22/i0[6] ), .ZN(\SB3_22/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U2179 ( .A1(\SB3_22/i0_3 ), .A2(\SB3_22/i0[8] ), .A3(\SB3_22/i0[9] ), .ZN(\SB3_22/Component_Function_2/NAND4_in[2] ) );
  NAND2_X1 U2203 ( .A1(\SB2_3_25/i0_3 ), .A2(\SB2_3_25/i1[9] ), .ZN(
        \SB2_3_25/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U2204 ( .A1(\SB2_3_25/i0_3 ), .A2(\SB1_3_26/buf_output[4] ), .A3(
        \SB2_3_25/i1[9] ), .ZN(n1161) );
  NAND3_X1 U2206 ( .A1(\SB2_3_25/i1_5 ), .A2(\SB2_3_25/i0[10] ), .A3(
        \SB2_3_25/i1[9] ), .ZN(\SB2_3_25/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U2208 ( .A1(\SB2_3_25/i1[9] ), .A2(\SB2_3_25/i0_3 ), .A3(
        \SB2_3_25/i0[6] ), .ZN(\SB2_3_25/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2212 ( .A1(\SB2_3_25/i1[9] ), .A2(\SB1_3_26/buf_output[4] ), .A3(
        \SB2_3_25/i1_5 ), .ZN(n4492) );
  NAND3_X1 U2216 ( .A1(\SB3_13/i0_3 ), .A2(\SB3_13/i0[10] ), .A3(
        \SB3_13/i0[6] ), .ZN(\SB3_13/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U2218 ( .A1(\SB3_13/i1_5 ), .A2(\SB3_13/i0[10] ), .A3(
        \SB3_13/i1[9] ), .ZN(\SB3_13/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U2219 ( .A1(\SB3_13/i0[10] ), .A2(\SB3_13/i1[9] ), .A3(
        \SB3_13/i1_7 ), .ZN(n3617) );
  CLKBUF_X4 U2233 ( .I(\SB2_1_12/buf_output[3] ), .Z(\RI5[1][129] ) );
  INV_X1 U2235 ( .I(\MC_ARK_ARC_1_2/buf_output[24] ), .ZN(\SB1_3_27/i3[0] ) );
  BUF_X2 U2238 ( .I(\MC_ARK_ARC_1_2/buf_output[24] ), .Z(\SB1_3_27/i0[9] ) );
  CLKBUF_X4 U2239 ( .I(\SB3_1/buf_output[4] ), .Z(\SB4_0/i0_4 ) );
  CLKBUF_X4 U2241 ( .I(\SB3_17/buf_output[5] ), .Z(\SB4_17/i0_3 ) );
  NAND3_X1 U2242 ( .A1(\SB4_21/i0[7] ), .A2(\SB4_21/i0_3 ), .A3(
        \SB3_24/buf_output[2] ), .ZN(\SB4_21/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2243 ( .A1(\SB4_17/i0[9] ), .A2(\SB4_17/i0_0 ), .A3(n3661), .ZN(
        \SB4_17/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U2244 ( .A1(\SB4_17/i0_4 ), .A2(\SB4_17/i0_0 ), .A3(\SB4_17/i1_5 ), 
        .ZN(n3564) );
  NAND3_X1 U2247 ( .A1(\SB4_24/i1[9] ), .A2(\SB4_24/i1_5 ), .A3(\SB4_24/i0_4 ), 
        .ZN(\SB4_24/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U2248 ( .A1(\SB4_24/i1_5 ), .A2(\SB4_24/i0_0 ), .A3(\SB4_24/i0_4 ), 
        .ZN(\SB4_24/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U2251 ( .A1(\SB1_2_11/i1_5 ), .A2(\SB1_2_11/i0[10] ), .A3(
        \SB1_2_11/i1[9] ), .ZN(\SB1_2_11/Component_Function_2/NAND4_in[0] ) );
  NAND2_X1 U2252 ( .A1(\SB1_2_11/i0_3 ), .A2(\SB1_2_11/i1[9] ), .ZN(
        \SB1_2_11/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U2253 ( .A1(\SB1_2_11/i1[9] ), .A2(\SB1_2_11/i0_3 ), .A3(
        \SB1_2_11/i0[6] ), .ZN(\SB1_2_11/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2257 ( .A1(\SB1_2_11/i1[9] ), .A2(\SB1_2_11/i1_7 ), .A3(
        \SB1_2_11/i0[10] ), .ZN(\SB1_2_11/Component_Function_3/NAND4_in[2] )
         );
  INV_X1 U2267 ( .I(\RI1[4][29] ), .ZN(\SB3_27/i1_5 ) );
  CLKBUF_X4 U2269 ( .I(\RI1[4][29] ), .Z(\SB3_27/i0_3 ) );
  NAND3_X1 U2270 ( .A1(\SB1_2_9/i1[9] ), .A2(\SB1_2_9/i1_5 ), .A3(
        \MC_ARK_ARC_1_1/buf_output[136] ), .ZN(
        \SB1_2_9/Component_Function_4/NAND4_in[3] ) );
  NAND2_X1 U2273 ( .A1(\SB1_2_9/i0_3 ), .A2(\SB1_2_9/i1[9] ), .ZN(
        \SB1_2_9/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U2279 ( .A1(\SB3_10/i0[6] ), .A2(\SB3_10/i0[10] ), .A3(
        \SB3_10/i0_0 ), .ZN(n4129) );
  NAND3_X1 U2284 ( .A1(\SB3_10/i0_3 ), .A2(\SB3_10/i0[10] ), .A3(
        \SB3_10/i0[6] ), .ZN(\SB3_10/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U2288 ( .A1(\SB2_3_30/i0_3 ), .A2(\SB2_3_30/i0[7] ), .A3(
        \SB2_3_30/i0_0 ), .ZN(\SB2_3_30/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 U2289 ( .A1(\SB2_3_30/i0_3 ), .A2(\SB2_3_30/i1[9] ), .ZN(
        \SB2_3_30/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U2291 ( .A1(\SB2_3_30/i0_3 ), .A2(\SB2_3_30/i0[10] ), .A3(
        \SB2_3_30/i0[9] ), .ZN(\SB2_3_30/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2293 ( .A1(\SB2_3_30/i0_4 ), .A2(\SB2_3_30/i0_3 ), .A3(
        \SB2_3_30/i0[10] ), .ZN(n4540) );
  INV_X1 U2301 ( .I(\MC_ARK_ARC_1_2/buf_output[60] ), .ZN(\SB1_3_21/i3[0] ) );
  BUF_X2 U2318 ( .I(\MC_ARK_ARC_1_3/buf_output[28] ), .Z(\SB3_27/i0_4 ) );
  INV_X1 U2320 ( .I(\MC_ARK_ARC_1_2/buf_output[115] ), .ZN(\SB1_3_12/i1_7 ) );
  NAND3_X1 U2321 ( .A1(\SB4_19/i0[9] ), .A2(\SB3_21/buf_output[3] ), .A3(
        \SB4_19/i0_3 ), .ZN(\SB4_19/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2327 ( .A1(\SB3_1/i1_7 ), .A2(\SB3_1/i0[8] ), .A3(\SB3_1/i0_4 ), 
        .ZN(\SB3_1/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U2344 ( .A1(\SB2_3_16/i0[9] ), .A2(\SB2_3_16/i0[10] ), .A3(
        \SB2_3_16/i0_3 ), .ZN(\SB2_3_16/Component_Function_4/NAND4_in[2] ) );
  CLKBUF_X4 U2353 ( .I(\SB1_2_3/buf_output[1] ), .Z(\SB2_2_31/i0[6] ) );
  INV_X1 U2363 ( .I(\SB3_13/buf_output[3] ), .ZN(\SB4_11/i0[8] ) );
  NAND2_X1 U2367 ( .A1(\SB2_3_11/i0_0 ), .A2(\SB2_3_11/i3[0] ), .ZN(
        \SB2_3_11/Component_Function_5/NAND4_in[0] ) );
  INV_X1 U2374 ( .I(\MC_ARK_ARC_1_2/buf_output[97] ), .ZN(\SB1_3_15/i1_7 ) );
  BUF_X2 U2376 ( .I(\MC_ARK_ARC_1_2/buf_output[97] ), .Z(\SB1_3_15/i0[6] ) );
  CLKBUF_X4 U2378 ( .I(\MC_ARK_ARC_1_3/buf_output[164] ), .Z(\SB3_4/i0_0 ) );
  NAND2_X1 U2391 ( .A1(\SB2_0_17/i0_3 ), .A2(\SB2_0_17/i1[9] ), .ZN(
        \SB2_0_17/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U2416 ( .A1(\SB1_3_15/i0[7] ), .A2(\SB1_3_15/i0_3 ), .A3(
        \SB1_3_15/i0_0 ), .ZN(\SB1_3_15/Component_Function_0/NAND4_in[3] ) );
  INV_X1 U2418 ( .I(\MC_ARK_ARC_1_1/buf_output[31] ), .ZN(\SB1_2_26/i1_7 ) );
  INV_X1 U2428 ( .I(\MC_ARK_ARC_1_0/buf_output[168] ), .ZN(\SB1_1_3/i3[0] ) );
  NAND3_X1 U2432 ( .A1(\SB2_3_19/i0[10] ), .A2(\SB2_3_19/i0_3 ), .A3(
        \SB2_3_19/i0[6] ), .ZN(n1683) );
  NAND3_X1 U2443 ( .A1(\SB3_0/i0[8] ), .A2(\SB3_0/i0[7] ), .A3(\SB3_0/i0[6] ), 
        .ZN(\SB3_0/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U2462 ( .A1(\SB4_28/i0[6] ), .A2(\SB4_28/i0[9] ), .A3(\SB4_28/i0_4 ), .ZN(n2394) );
  NAND3_X1 U2473 ( .A1(\SB3_18/i0_0 ), .A2(\SB3_18/i0[6] ), .A3(
        \SB3_18/i0[10] ), .ZN(n4200) );
  OAI21_X1 U2478 ( .A1(n2902), .A2(n3150), .B(\SB2_3_6/i0_0 ), .ZN(n4016) );
  CLKBUF_X4 U2483 ( .I(\SB1_3_6/buf_output[5] ), .Z(\SB2_3_6/i0_3 ) );
  NAND3_X1 U2489 ( .A1(\SB1_3_18/i0_0 ), .A2(\SB1_3_18/i0_4 ), .A3(
        \SB1_3_18/i0_3 ), .ZN(\SB1_3_18/Component_Function_3/NAND4_in[1] ) );
  BUF_X2 U2509 ( .I(\SB3_15/buf_output[2] ), .Z(\SB4_12/i0_0 ) );
  INV_X1 U2510 ( .I(\SB3_15/buf_output[2] ), .ZN(\SB4_12/i1[9] ) );
  NAND3_X1 U2518 ( .A1(\SB1_1_14/i0[9] ), .A2(\SB1_1_14/i0[10] ), .A3(
        \SB1_1_14/i0_3 ), .ZN(\SB1_1_14/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2526 ( .A1(n1793), .A2(\SB4_29/i1_7 ), .A3(\SB4_29/i0[8] ), .ZN(
        n4096) );
  NAND3_X1 U2530 ( .A1(\SB4_10/i0[10] ), .A2(\SB4_10/i0[6] ), .A3(
        \SB4_10/i0_3 ), .ZN(n1511) );
  NAND3_X1 U2532 ( .A1(\SB4_20/i0[10] ), .A2(\SB4_20/i0_0 ), .A3(
        \SB4_20/i0[6] ), .ZN(n2436) );
  NAND2_X1 U2535 ( .A1(\SB4_20/i0[10] ), .A2(\SB4_20/i0[9] ), .ZN(
        \SB4_20/Component_Function_0/NAND4_in[0] ) );
  INV_X1 U2537 ( .I(\MC_ARK_ARC_1_3/buf_output[55] ), .ZN(\SB3_22/i1_7 ) );
  BUF_X2 U2543 ( .I(\MC_ARK_ARC_1_3/buf_output[55] ), .Z(\SB3_22/i0[6] ) );
  CLKBUF_X4 U2546 ( .I(\MC_ARK_ARC_1_0/buf_output[47] ), .Z(\SB1_1_24/i0_3 )
         );
  NAND3_X1 U2553 ( .A1(\SB4_10/i0[9] ), .A2(\SB3_13/buf_output[2] ), .A3(
        \SB4_10/i0[8] ), .ZN(\SB4_10/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U2555 ( .A1(\SB4_10/i0[9] ), .A2(\SB4_10/i0_3 ), .A3(\SB4_10/i0[8] ), .ZN(n4554) );
  NAND3_X1 U2562 ( .A1(\SB2_3_14/i0_0 ), .A2(\SB2_3_14/i0_3 ), .A3(
        \SB2_3_14/i0_4 ), .ZN(\SB2_3_14/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2563 ( .A1(\SB2_3_14/i0_3 ), .A2(\SB2_3_14/i0_4 ), .A3(
        \SB2_3_14/i1[9] ), .ZN(n4688) );
  INV_X1 U2586 ( .I(\MC_ARK_ARC_1_3/buf_output[145] ), .ZN(\SB3_7/i1_7 ) );
  BUF_X2 U2587 ( .I(\MC_ARK_ARC_1_3/buf_output[145] ), .Z(\SB3_7/i0[6] ) );
  NAND3_X1 U2596 ( .A1(\RI3[0][155] ), .A2(\SB2_0_6/i0[8] ), .A3(
        \SB1_0_11/buf_output[0] ), .ZN(
        \SB2_0_6/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2599 ( .A1(\RI3[0][155] ), .A2(\SB2_0_6/i1_7 ), .A3(
        \SB2_0_6/i0[8] ), .ZN(\SB2_0_6/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U2601 ( .A1(\SB1_3_13/i0_3 ), .A2(\SB1_3_13/i0[10] ), .A3(
        \SB1_3_13/i0[6] ), .ZN(\SB1_3_13/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U2616 ( .A1(\SB4_16/i0_0 ), .A2(\SB4_16/i3[0] ), .A3(\SB4_16/i1_7 ), 
        .ZN(n2680) );
  NAND2_X1 U2617 ( .A1(\SB4_16/i0_0 ), .A2(\SB4_16/i3[0] ), .ZN(
        \SB4_16/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U2618 ( .A1(\SB4_16/i0_0 ), .A2(\SB4_16/i0_3 ), .A3(\SB4_16/i0[7] ), 
        .ZN(n3838) );
  NAND3_X1 U2623 ( .A1(\SB4_16/i0_0 ), .A2(\SB4_16/i0_3 ), .A3(\SB4_16/i0_4 ), 
        .ZN(n3622) );
  NAND3_X1 U2632 ( .A1(\SB2_2_29/i0_3 ), .A2(\SB2_2_29/i0_0 ), .A3(n1837), 
        .ZN(\SB2_2_29/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2646 ( .A1(\SB1_0_26/i0_3 ), .A2(\SB1_0_26/i0[8] ), .A3(
        \SB1_0_26/i1_7 ), .ZN(\SB1_0_26/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U2647 ( .A1(\SB1_0_26/i0_3 ), .A2(\SB1_0_26/i0[10] ), .A3(
        \SB1_0_26/i0[6] ), .ZN(\SB1_0_26/Component_Function_2/NAND4_in[1] ) );
  NAND2_X1 U2648 ( .A1(\SB1_0_26/i0_3 ), .A2(\SB1_0_26/i1[9] ), .ZN(
        \SB1_0_26/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U2649 ( .A1(\SB1_0_26/i0_3 ), .A2(\SB1_0_26/i0_4 ), .A3(
        \SB1_0_26/i1[9] ), .ZN(\SB1_0_26/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2650 ( .A1(\SB1_3_1/i0_4 ), .A2(\SB1_3_1/i1[9] ), .A3(
        \SB1_3_1/i1_5 ), .ZN(\SB1_3_1/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U2653 ( .A1(\SB1_3_1/i0[10] ), .A2(\SB1_3_1/i1[9] ), .A3(
        \SB1_3_1/i1_7 ), .ZN(n3934) );
  NAND3_X1 U2654 ( .A1(\SB1_3_1/i1[9] ), .A2(\SB1_3_1/i0_3 ), .A3(
        \SB1_3_1/i0[6] ), .ZN(\SB1_3_1/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2657 ( .A1(\SB2_1_23/i0_3 ), .A2(\SB2_1_23/i0_4 ), .A3(
        \SB2_1_23/i0[10] ), .ZN(\SB2_1_23/Component_Function_0/NAND4_in[2] )
         );
  NAND3_X1 U2667 ( .A1(\SB2_1_23/i0_3 ), .A2(\SB2_1_23/i0_0 ), .A3(
        \SB2_1_23/i0[7] ), .ZN(\SB2_1_23/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2696 ( .A1(\SB4_9/i0_0 ), .A2(\SB4_9/i0[6] ), .A3(\SB4_9/i0[10] ), 
        .ZN(\SB4_9/Component_Function_5/NAND4_in[1] ) );
  INV_X1 U2701 ( .I(\SB3_3/buf_output[3] ), .ZN(\SB4_1/i0[8] ) );
  NAND3_X1 U2703 ( .A1(\SB3_27/i0_0 ), .A2(\SB3_27/i0_4 ), .A3(\SB3_27/i1_5 ), 
        .ZN(n590) );
  NAND3_X1 U2719 ( .A1(\SB4_9/i0[9] ), .A2(\SB4_9/i0[8] ), .A3(\SB4_9/i0_0 ), 
        .ZN(n3953) );
  NAND3_X1 U2721 ( .A1(\SB4_9/i1_5 ), .A2(\SB4_9/i0[8] ), .A3(\SB4_9/i3[0] ), 
        .ZN(\SB4_9/Component_Function_3/NAND4_in[3] ) );
  INV_X1 U2729 ( .I(\MC_ARK_ARC_1_3/buf_output[174] ), .ZN(\SB3_2/i3[0] ) );
  NAND3_X1 U2735 ( .A1(\SB1_1_1/i1_5 ), .A2(\SB1_1_1/i0[10] ), .A3(
        \SB1_1_1/i1[9] ), .ZN(\SB1_1_1/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U2740 ( .A1(n3653), .A2(\SB4_10/i0_4 ), .A3(\SB4_10/i0_3 ), .ZN(
        \SB4_10/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 U2760 ( .A1(\SB2_2_19/i0_3 ), .A2(\SB2_2_19/i1[9] ), .ZN(
        \SB2_2_19/Component_Function_1/NAND4_in[0] ) );
  INV_X1 U2763 ( .I(\SB3_30/buf_output[3] ), .ZN(\SB4_28/i0[8] ) );
  BUF_X2 U2769 ( .I(n351), .Z(\SB1_0_26/i0[10] ) );
  INV_X1 U2770 ( .I(n351), .ZN(\SB1_0_26/i0[8] ) );
  NAND3_X1 U2771 ( .A1(\SB3_19/i0_3 ), .A2(\SB3_19/i0_4 ), .A3(\SB3_19/i0_0 ), 
        .ZN(n4351) );
  NAND3_X1 U2775 ( .A1(\SB4_17/i0[10] ), .A2(\SB4_17/i0_3 ), .A3(
        \SB4_17/i0[6] ), .ZN(\SB4_17/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U2776 ( .A1(\SB4_17/i0[10] ), .A2(\SB4_17/i0[9] ), .A3(
        \SB4_17/i0_3 ), .ZN(n4156) );
  NAND2_X1 U2779 ( .A1(\SB4_17/i0_3 ), .A2(\SB4_17/i1[9] ), .ZN(
        \SB4_17/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U2785 ( .A1(\SB4_17/i0_0 ), .A2(\SB4_17/i0_3 ), .A3(\SB4_17/i0[7] ), 
        .ZN(n3836) );
  BUF_X2 U2801 ( .I(\MC_ARK_ARC_1_3/buf_output[51] ), .Z(\SB3_23/i0[10] ) );
  INV_X1 U2802 ( .I(\MC_ARK_ARC_1_3/buf_output[51] ), .ZN(\SB3_23/i0[8] ) );
  INV_X1 U2818 ( .I(\MC_ARK_ARC_1_3/buf_output[9] ), .ZN(\SB3_30/i0[8] ) );
  BUF_X2 U2819 ( .I(\MC_ARK_ARC_1_3/buf_output[9] ), .Z(\SB3_30/i0[10] ) );
  NAND3_X1 U2824 ( .A1(\SB3_18/i1[9] ), .A2(\SB3_18/i1_5 ), .A3(\SB3_18/i0_4 ), 
        .ZN(\SB3_18/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U2840 ( .A1(\SB1_3_4/i0_4 ), .A2(\SB1_3_4/i1[9] ), .A3(
        \SB1_3_4/i1_5 ), .ZN(n3450) );
  INV_X1 U2841 ( .I(\MC_ARK_ARC_1_2/buf_output[78] ), .ZN(\SB1_3_18/i3[0] ) );
  INV_X1 U2845 ( .I(\MC_ARK_ARC_1_2/buf_output[85] ), .ZN(\SB1_3_17/i1_7 ) );
  BUF_X2 U2846 ( .I(\MC_ARK_ARC_1_2/buf_output[85] ), .Z(\SB1_3_17/i0[6] ) );
  CLKBUF_X4 U2847 ( .I(\RI1[4][131] ), .Z(\SB3_10/i0_3 ) );
  INV_X1 U2848 ( .I(\RI1[4][131] ), .ZN(\SB3_10/i1_5 ) );
  BUF_X2 U2849 ( .I(\MC_ARK_ARC_1_2/buf_output[181] ), .Z(\SB1_3_1/i0[6] ) );
  INV_X1 U2850 ( .I(\MC_ARK_ARC_1_2/buf_output[181] ), .ZN(\SB1_3_1/i1_7 ) );
  BUF_X2 U2863 ( .I(n288), .Z(\SB1_0_17/i0[6] ) );
  INV_X1 U2866 ( .I(n288), .ZN(\SB1_0_17/i1_7 ) );
  INV_X1 U2874 ( .I(\MC_ARK_ARC_1_2/buf_output[93] ), .ZN(\SB1_3_16/i0[8] ) );
  BUF_X2 U2875 ( .I(\MC_ARK_ARC_1_2/buf_output[93] ), .Z(\SB1_3_16/i0[10] ) );
  NAND3_X1 U2876 ( .A1(\SB3_2/i0_0 ), .A2(\SB3_2/i1_5 ), .A3(\SB3_2/i0_4 ), 
        .ZN(n2313) );
  INV_X1 U2901 ( .I(\SB3_16/buf_output[5] ), .ZN(\SB4_16/i1_5 ) );
  NAND3_X1 U2919 ( .A1(\SB1_3_26/i0[6] ), .A2(\SB1_3_26/i1_5 ), .A3(
        \SB1_3_26/i0[9] ), .ZN(n3011) );
  INV_X1 U2928 ( .I(\SB3_21/buf_output[0] ), .ZN(\SB4_16/i3[0] ) );
  CLKBUF_X4 U2929 ( .I(\SB3_27/buf_output[5] ), .Z(\SB4_27/i0_3 ) );
  NAND3_X1 U2931 ( .A1(\SB4_24/i0_3 ), .A2(\SB4_24/i0[9] ), .A3(
        \SB4_24/i0[10] ), .ZN(n4545) );
  NAND3_X1 U2932 ( .A1(\SB4_24/i0_3 ), .A2(\SB4_24/i0_0 ), .A3(\SB4_24/i0_4 ), 
        .ZN(\SB4_24/Component_Function_3/NAND4_in[1] ) );
  NAND2_X1 U2933 ( .A1(\SB4_24/i0_3 ), .A2(\SB4_24/i1[9] ), .ZN(
        \SB4_24/Component_Function_1/NAND4_in[0] ) );
  INV_X1 U2934 ( .I(\MC_ARK_ARC_1_0/buf_output[140] ), .ZN(\SB1_1_8/i1[9] ) );
  BUF_X2 U2935 ( .I(\MC_ARK_ARC_1_0/buf_output[140] ), .Z(\SB1_1_8/i0_0 ) );
  INV_X1 U2938 ( .I(\MC_ARK_ARC_1_0/buf_output[72] ), .ZN(\SB1_1_19/i3[0] ) );
  NAND3_X1 U2945 ( .A1(\SB1_0_13/i1_5 ), .A2(\SB1_0_13/i0[6] ), .A3(
        \SB1_0_13/i0[9] ), .ZN(\SB1_0_13/Component_Function_1/NAND4_in[2] ) );
  XNOR2_X1 U2952 ( .A1(\MC_ARK_ARC_1_1/temp6[69] ), .A2(
        \MC_ARK_ARC_1_1/temp5[69] ), .ZN(n2893) );
  BUF_X4 U2954 ( .I(\MC_ARK_ARC_1_3/buf_datainput[90] ), .Z(n2896) );
  CLKBUF_X4 U2955 ( .I(\MC_ARK_ARC_1_0/buf_output[184] ), .Z(\SB1_1_1/i0_4 )
         );
  INV_X1 U2960 ( .I(\MC_ARK_ARC_1_0/buf_output[181] ), .ZN(\SB1_1_1/i1_7 ) );
  NAND3_X1 U2965 ( .A1(\SB2_1_15/i0_0 ), .A2(\SB2_1_15/i0_4 ), .A3(
        \SB2_1_15/i1_5 ), .ZN(n2842) );
  NAND3_X2 U2972 ( .A1(\SB2_0_3/i0[10] ), .A2(\RI3[0][172] ), .A3(
        \SB2_0_3/i0_3 ), .ZN(\SB2_0_3/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U2974 ( .A1(\SB1_2_27/i0[10] ), .A2(\SB1_2_27/i0_0 ), .A3(
        \SB1_2_27/i0[6] ), .ZN(n933) );
  NAND3_X1 U2979 ( .A1(\RI1[1][143] ), .A2(\SB1_1_8/i1[9] ), .A3(
        \SB1_1_8/i0[6] ), .ZN(\SB1_1_8/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 U2984 ( .I(\SB1_2_11/buf_output[5] ), .Z(\SB2_2_11/i0_3 ) );
  BUF_X4 U3021 ( .I(\SB1_3_22/buf_output[5] ), .Z(\SB2_3_22/i0_3 ) );
  CLKBUF_X2 U3025 ( .I(\SB1_2_13/buf_output[0] ), .Z(\SB2_2_8/i0[9] ) );
  NAND3_X1 U3030 ( .A1(\SB1_3_13/i1[9] ), .A2(\SB1_3_13/i1_5 ), .A3(
        \SB1_3_13/i0_4 ), .ZN(\SB1_3_13/Component_Function_4/NAND4_in[3] ) );
  CLKBUF_X4 U3031 ( .I(\MC_ARK_ARC_1_2/buf_output[182] ), .Z(\SB1_3_1/i0_0 )
         );
  INV_X1 U3047 ( .I(n408), .ZN(\SB1_0_28/i1_5 ) );
  INV_X1 U3050 ( .I(\MC_ARK_ARC_1_0/buf_output[31] ), .ZN(\SB1_1_26/i1_7 ) );
  BUF_X2 U3051 ( .I(\MC_ARK_ARC_1_0/buf_output[31] ), .Z(\SB1_1_26/i0[6] ) );
  INV_X1 U3055 ( .I(\SB1_3_30/buf_output[1] ), .ZN(\SB2_3_26/i1_7 ) );
  NAND4_X1 U3057 ( .A1(\SB1_0_15/Component_Function_3/NAND4_in[3] ), .A2(
        \SB1_0_15/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_0_15/Component_Function_3/NAND4_in[1] ), .A4(n2330), .ZN(
        \SB1_0_15/buf_output[3] ) );
  BUF_X2 U3058 ( .I(\MC_ARK_ARC_1_3/buf_output[6] ), .Z(\SB3_30/i0[9] ) );
  INV_X1 U3061 ( .I(\MC_ARK_ARC_1_0/buf_output[61] ), .ZN(\SB1_1_21/i1_7 ) );
  BUF_X2 U3062 ( .I(\MC_ARK_ARC_1_0/buf_output[61] ), .Z(\SB1_1_21/i0[6] ) );
  CLKBUF_X4 U3065 ( .I(\MC_ARK_ARC_1_0/buf_output[164] ), .Z(\SB1_1_4/i0_0 )
         );
  NAND3_X1 U3066 ( .A1(\SB1_0_26/i0[10] ), .A2(\SB1_0_26/i0_3 ), .A3(
        \SB1_0_26/i0_4 ), .ZN(n1124) );
  NAND2_X1 U3069 ( .A1(\SB1_1_0/i0_3 ), .A2(\SB1_1_0/i1[9] ), .ZN(n1980) );
  NAND3_X1 U3071 ( .A1(\SB1_1_0/i0[10] ), .A2(\SB1_1_0/i0_4 ), .A3(
        \SB1_1_0/i0_3 ), .ZN(\SB1_1_0/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3072 ( .A1(\SB1_1_0/i0[6] ), .A2(\SB1_1_0/i0_3 ), .A3(
        \SB1_1_0/i0[10] ), .ZN(n1318) );
  BUF_X4 U3079 ( .I(\MC_ARK_ARC_1_2/buf_output[86] ), .Z(\SB1_3_17/i0_0 ) );
  INV_X1 U3080 ( .I(\MC_ARK_ARC_1_2/buf_output[12] ), .ZN(\SB1_3_29/i3[0] ) );
  INV_X1 U3088 ( .I(\SB1_2_15/buf_output[1] ), .ZN(\SB2_2_11/i1_7 ) );
  BUF_X2 U3089 ( .I(\SB1_2_15/buf_output[1] ), .Z(\SB2_2_11/i0[6] ) );
  NAND3_X1 U3091 ( .A1(\MC_ARK_ARC_1_2/buf_output[9] ), .A2(\SB1_3_30/i1[9] ), 
        .A3(\SB1_3_30/i1_7 ), .ZN(n4664) );
  NAND3_X1 U3096 ( .A1(\SB1_3_30/i1_5 ), .A2(\SB1_3_30/i0[10] ), .A3(
        \SB1_3_30/i1[9] ), .ZN(\SB1_3_30/Component_Function_2/NAND4_in[0] ) );
  NAND2_X1 U3099 ( .A1(\SB1_2_20/i0_3 ), .A2(\SB1_2_20/i1[9] ), .ZN(
        \SB1_2_20/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U3101 ( .A1(\SB1_3_21/i0[7] ), .A2(\SB1_3_21/i0_3 ), .A3(
        \SB1_3_21/i0_0 ), .ZN(\SB1_3_21/Component_Function_0/NAND4_in[3] ) );
  NAND3_X2 U3117 ( .A1(\SB2_0_13/i0_4 ), .A2(n1393), .A3(\SB2_0_13/i1_7 ), 
        .ZN(n2040) );
  BUF_X2 U3120 ( .I(\SB1_0_1/buf_output[0] ), .Z(\RI3[0][18] ) );
  INV_X1 U3122 ( .I(\SB1_0_1/buf_output[0] ), .ZN(\SB2_0_28/i3[0] ) );
  INV_X1 U3127 ( .I(\MC_ARK_ARC_1_0/buf_output[58] ), .ZN(\SB1_1_22/i0[7] ) );
  BUF_X4 U3130 ( .I(\SB1_2_16/buf_output[2] ), .Z(\SB2_2_13/i0_0 ) );
  NAND3_X1 U3131 ( .A1(\SB2_2_10/i0[10] ), .A2(\SB2_2_10/i1[9] ), .A3(
        \SB2_2_10/i1_5 ), .ZN(\SB2_2_10/Component_Function_2/NAND4_in[0] ) );
  INV_X1 U3137 ( .I(\MC_ARK_ARC_1_3/buf_output[127] ), .ZN(\SB3_10/i1_7 ) );
  NAND3_X1 U3140 ( .A1(\SB1_2_6/i1[9] ), .A2(\SB1_2_6/i1_5 ), .A3(
        \SB1_2_6/i0_4 ), .ZN(\SB1_2_6/Component_Function_4/NAND4_in[3] ) );
  CLKBUF_X4 U3149 ( .I(\SB3_17/buf_output[4] ), .Z(\SB4_16/i0_4 ) );
  NAND3_X1 U3152 ( .A1(\SB2_2_16/i0[10] ), .A2(\SB2_2_16/i1[9] ), .A3(
        \SB2_2_16/i1_7 ), .ZN(\SB2_2_16/Component_Function_3/NAND4_in[2] ) );
  BUF_X2 U3165 ( .I(n270), .Z(\SB1_0_23/i0[6] ) );
  INV_X1 U3166 ( .I(n270), .ZN(\SB1_0_23/i1_7 ) );
  CLKBUF_X4 U3167 ( .I(\SB1_0_29/buf_output[5] ), .Z(\SB2_0_29/i0_3 ) );
  NAND3_X1 U3170 ( .A1(\SB1_0_23/i1[9] ), .A2(\SB1_0_23/i0_3 ), .A3(
        \SB1_0_23/i0[6] ), .ZN(\SB1_0_23/Component_Function_3/NAND4_in[0] ) );
  CLKBUF_X4 U3184 ( .I(\MC_ARK_ARC_1_1/buf_output[152] ), .Z(\SB1_2_6/i0_0 )
         );
  OR3_X2 U3185 ( .A1(\MC_ARK_ARC_1_0/buf_output[51] ), .A2(
        \MC_ARK_ARC_1_0/buf_output[53] ), .A3(\MC_ARK_ARC_1_0/buf_output[48] ), 
        .Z(n4573) );
  BUF_X2 U3195 ( .I(\SB3_8/buf_output[4] ), .Z(\SB4_7/i0_4 ) );
  BUF_X2 U3199 ( .I(\SB3_14/buf_output[3] ), .Z(\SB4_12/i0[10] ) );
  BUF_X2 U3200 ( .I(\SB3_29/buf_output[1] ), .Z(\SB4_25/i0[6] ) );
  CLKBUF_X4 U3204 ( .I(\MC_ARK_ARC_1_3/buf_output[66] ), .Z(\SB3_20/i0[9] ) );
  BUF_X2 U3209 ( .I(\MC_ARK_ARC_1_3/buf_output[31] ), .Z(\SB3_26/i0[6] ) );
  CLKBUF_X4 U3210 ( .I(\MC_ARK_ARC_1_3/buf_output[44] ), .Z(\SB3_24/i0_0 ) );
  BUF_X2 U3213 ( .I(\MC_ARK_ARC_1_3/buf_output[37] ), .Z(\SB3_25/i0[6] ) );
  CLKBUF_X4 U3214 ( .I(\MC_ARK_ARC_1_3/buf_output[10] ), .Z(\SB3_30/i0_4 ) );
  BUF_X2 U3217 ( .I(\MC_ARK_ARC_1_3/buf_output[139] ), .Z(\SB3_8/i0[6] ) );
  BUF_X4 U3218 ( .I(\SB2_3_16/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[115] ) );
  BUF_X4 U3232 ( .I(\SB2_3_12/buf_output[0] ), .Z(\RI5[3][144] ) );
  AND2_X1 U3235 ( .A1(\SB2_3_6/i3[0] ), .A2(\SB2_3_6/i1_7 ), .Z(n2902) );
  NAND2_X1 U3236 ( .A1(n3680), .A2(n4272), .ZN(n1617) );
  CLKBUF_X4 U3238 ( .I(\SB1_3_13/buf_output[4] ), .Z(\SB2_3_12/i0_4 ) );
  CLKBUF_X4 U3241 ( .I(\SB1_3_28/buf_output[2] ), .Z(\SB2_3_25/i0_0 ) );
  NAND2_X1 U3243 ( .A1(\SB1_3_4/i0[9] ), .A2(n3122), .ZN(
        \SB1_3_4/Component_Function_5/NAND4_in[3] ) );
  BUF_X2 U3245 ( .I(\MC_ARK_ARC_1_2/buf_output[67] ), .Z(\SB1_3_20/i0[6] ) );
  BUF_X4 U3253 ( .I(\SB2_2_5/buf_output[5] ), .Z(\RI5[2][161] ) );
  BUF_X4 U3259 ( .I(\SB1_2_20/buf_output[5] ), .Z(\SB2_2_20/i0_3 ) );
  INV_X4 U3260 ( .I(n3333), .ZN(\SB2_2_9/i0_4 ) );
  CLKBUF_X4 U3272 ( .I(\MC_ARK_ARC_1_1/buf_output[69] ), .Z(\SB1_2_20/i0[10] )
         );
  BUF_X4 U3273 ( .I(n3682), .Z(\SB1_2_21/i0_3 ) );
  BUF_X4 U3274 ( .I(\SB2_1_3/buf_output[0] ), .Z(\RI5[1][6] ) );
  BUF_X4 U3275 ( .I(\SB2_1_5/buf_output[2] ), .Z(\RI5[1][176] ) );
  CLKBUF_X2 U3283 ( .I(\SB2_1_11/i0[7] ), .Z(n3885) );
  CLKBUF_X4 U3287 ( .I(\SB1_1_24/buf_output[3] ), .Z(\SB2_1_22/i0[10] ) );
  BUF_X2 U3293 ( .I(\SB1_1_31/buf_output[0] ), .Z(\SB2_1_26/i0[9] ) );
  NAND2_X1 U3294 ( .A1(\SB1_1_12/Component_Function_4/NAND4_in[2] ), .A2(n2581), .ZN(n4701) );
  NAND2_X1 U3297 ( .A1(\SB1_1_22/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_1_22/Component_Function_1/NAND4_in[0] ), .ZN(n4141) );
  CLKBUF_X4 U3298 ( .I(\MC_ARK_ARC_1_0/buf_output[105] ), .Z(\SB1_1_14/i0[10] ) );
  CLKBUF_X4 U3300 ( .I(\MC_ARK_ARC_1_0/buf_output[174] ), .Z(\SB1_1_2/i0[9] )
         );
  BUF_X4 U3304 ( .I(\SB2_0_31/buf_output[3] ), .Z(\RI5[0][15] ) );
  BUF_X2 U3306 ( .I(\SB1_0_19/buf_output[0] ), .Z(\SB2_0_14/i0[9] ) );
  BUF_X2 U3309 ( .I(n251), .Z(\SB1_0_29/i0[9] ) );
  BUF_X2 U3311 ( .I(n305), .Z(\SB1_0_11/i0[9] ) );
  BUF_X2 U3313 ( .I(n272), .Z(\SB1_0_22/i0[9] ) );
  CLKBUF_X4 U3316 ( .I(n323), .Z(\SB1_0_5/i0[9] ) );
  BUF_X4 U3317 ( .I(n370), .Z(n2899) );
  NAND3_X1 U3319 ( .A1(\SB1_0_21/i0_3 ), .A2(\SB1_0_21/i0[9] ), .A3(
        \SB1_0_21/i0[10] ), .ZN(\SB1_0_21/Component_Function_4/NAND4_in[2] )
         );
  INV_X1 U3322 ( .I(n255), .ZN(\SB1_0_28/i1_7 ) );
  CLKBUF_X4 U3325 ( .I(n350), .Z(\SB1_0_27/i0_4 ) );
  INV_X1 U3329 ( .I(n392), .ZN(\SB1_0_6/i0[7] ) );
  NAND3_X1 U3336 ( .A1(\SB1_0_15/i0_3 ), .A2(\SB1_0_15/i0[9] ), .A3(
        \SB1_0_15/i0[8] ), .ZN(n2149) );
  NAND3_X1 U3337 ( .A1(\SB1_0_8/i0_3 ), .A2(\SB1_0_8/i1_7 ), .A3(
        \SB1_0_8/i0[8] ), .ZN(\SB1_0_8/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U3344 ( .A1(\SB1_0_21/i1_5 ), .A2(\SB1_0_21/i0[8] ), .A3(
        \SB1_0_21/i3[0] ), .ZN(\SB1_0_21/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U3346 ( .A1(\SB1_0_22/i0[10] ), .A2(\SB1_0_22/i1[9] ), .A3(
        \SB1_0_22/i1_7 ), .ZN(n1015) );
  NAND3_X1 U3347 ( .A1(\SB1_0_1/i1_7 ), .A2(\SB1_0_1/i0[8] ), .A3(
        \SB1_0_1/i0_4 ), .ZN(\SB1_0_1/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U3351 ( .A1(\SB1_0_30/i1_5 ), .A2(\SB1_0_30/i0_0 ), .A3(
        \SB1_0_30/i0_4 ), .ZN(\SB1_0_30/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U3352 ( .A1(\SB1_0_12/i0[7] ), .A2(\SB1_0_12/i0_3 ), .A3(
        \SB1_0_12/i0_0 ), .ZN(\SB1_0_12/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U3353 ( .A1(n4753), .A2(\SB1_0_18/i0[9] ), .A3(\SB1_0_18/i0[6] ), 
        .ZN(n1939) );
  NAND3_X1 U3356 ( .A1(\SB1_0_5/i0[7] ), .A2(\SB1_0_5/i0_3 ), .A3(
        \SB1_0_5/i0_0 ), .ZN(\SB1_0_5/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U3358 ( .A1(\SB1_0_2/i1[9] ), .A2(\SB1_0_2/i0_3 ), .A3(
        \SB1_0_2/i0[6] ), .ZN(\SB1_0_2/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U3363 ( .A1(\SB1_0_21/i0_3 ), .A2(\SB1_0_21/i0_0 ), .A3(
        \SB1_0_21/i0[7] ), .ZN(n4669) );
  NAND3_X1 U3367 ( .A1(\SB1_0_1/i0[10] ), .A2(\SB1_0_1/i0_3 ), .A3(
        \SB1_0_1/i0_4 ), .ZN(n3525) );
  NAND3_X1 U3368 ( .A1(\SB1_0_7/i0_3 ), .A2(\SB1_0_7/i0_0 ), .A3(n390), .ZN(
        \SB1_0_7/Component_Function_3/NAND4_in[1] ) );
  CLKBUF_X4 U3370 ( .I(\SB1_0_21/buf_output[1] ), .Z(\SB2_0_17/i0[6] ) );
  CLKBUF_X4 U3371 ( .I(\SB2_0_19/i0[10] ), .Z(n2774) );
  CLKBUF_X4 U3372 ( .I(\SB1_0_1/buf_output[1] ), .Z(\SB2_0_29/i0[6] ) );
  CLKBUF_X4 U3378 ( .I(\RI3[0][2] ), .Z(\SB2_0_31/i0_0 ) );
  NAND3_X1 U3384 ( .A1(\SB2_0_27/i0[8] ), .A2(\SB2_0_27/i1_7 ), .A3(
        \SB2_0_27/i0_4 ), .ZN(\SB2_0_27/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 U3387 ( .A1(\SB2_0_30/i0_0 ), .A2(\SB2_0_30/i3[0] ), .ZN(
        \SB2_0_30/Component_Function_5/NAND4_in[0] ) );
  INV_X1 U3394 ( .I(\SB1_0_19/buf_output[0] ), .ZN(\SB2_0_14/i3[0] ) );
  NAND3_X1 U3397 ( .A1(\SB2_0_16/i0_3 ), .A2(\SB2_0_16/i1_7 ), .A3(
        \SB2_0_16/i0[8] ), .ZN(\SB2_0_16/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U3399 ( .A1(\SB2_0_24/i1_7 ), .A2(\SB2_0_24/i0_0 ), .A3(
        \SB2_0_24/i3[0] ), .ZN(\SB2_0_24/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U3401 ( .A1(\SB2_0_18/i0_0 ), .A2(\SB2_0_18/i0_3 ), .A3(
        \SB2_0_18/i0[7] ), .ZN(n836) );
  NAND2_X1 U3403 ( .A1(\RI3[0][39] ), .A2(\SB2_0_25/i0[9] ), .ZN(
        \SB2_0_25/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U3405 ( .A1(\SB2_0_12/i0_0 ), .A2(\SB2_0_12/i0_3 ), .A3(
        \SB2_0_12/i0_4 ), .ZN(\SB2_0_12/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3407 ( .A1(\SB2_0_26/i1_7 ), .A2(\SB2_0_26/i0[8] ), .A3(
        \RI3[0][34] ), .ZN(\SB2_0_26/Component_Function_1/NAND4_in[3] ) );
  CLKBUF_X4 U3419 ( .I(\SB2_0_5/buf_output[3] ), .Z(\RI5[0][171] ) );
  INV_X1 U3420 ( .I(\MC_ARK_ARC_1_0/buf_output[106] ), .ZN(\SB1_1_14/i0[7] )
         );
  INV_X1 U3421 ( .I(\MC_ARK_ARC_1_0/buf_output[132] ), .ZN(\SB1_1_9/i3[0] ) );
  NAND2_X1 U3426 ( .A1(\SB1_1_22/i1_5 ), .A2(n4522), .ZN(
        \SB1_1_22/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U3432 ( .A1(\SB1_1_24/i0_3 ), .A2(\SB1_1_24/i0_4 ), .A3(
        \SB1_1_24/i1[9] ), .ZN(\SB1_1_24/Component_Function_5/NAND4_in[2] ) );
  INV_X1 U3441 ( .I(\MC_ARK_ARC_1_0/buf_output[162] ), .ZN(\SB1_1_4/i3[0] ) );
  CLKBUF_X4 U3443 ( .I(\MC_ARK_ARC_1_0/buf_output[70] ), .Z(\SB1_1_20/i0_4 )
         );
  CLKBUF_X4 U3445 ( .I(\MC_ARK_ARC_1_0/buf_output[76] ), .Z(\SB1_1_19/i0_4 )
         );
  NAND3_X1 U3448 ( .A1(\SB1_1_14/i0[8] ), .A2(\SB1_1_14/i1_5 ), .A3(
        \SB1_1_14/i3[0] ), .ZN(\SB1_1_14/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U3451 ( .A1(\SB1_1_13/i1_7 ), .A2(\SB1_1_13/i0[8] ), .A3(
        \SB1_1_13/i0_4 ), .ZN(\SB1_1_13/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U3453 ( .A1(\SB1_1_24/i0_3 ), .A2(\SB1_1_24/i1_7 ), .A3(
        \SB1_1_24/i0[8] ), .ZN(n4537) );
  NAND3_X1 U3455 ( .A1(\SB1_1_13/i1[9] ), .A2(\SB1_1_13/i0_3 ), .A3(
        \SB1_1_13/i0[6] ), .ZN(\SB1_1_13/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U3456 ( .A1(\SB1_1_2/i0_0 ), .A2(\SB1_1_2/i1_5 ), .A3(
        \SB1_1_2/i0_4 ), .ZN(\SB1_1_2/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U3460 ( .A1(\SB1_1_30/i1[9] ), .A2(\SB1_1_30/i1_7 ), .A3(
        \SB1_1_30/i0[10] ), .ZN(\SB1_1_30/Component_Function_3/NAND4_in[2] )
         );
  NAND3_X1 U3469 ( .A1(\SB1_1_28/i0[8] ), .A2(\SB1_1_28/i0[7] ), .A3(
        \SB1_1_28/i0[6] ), .ZN(\SB1_1_28/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U3470 ( .A1(\SB1_1_20/i0[8] ), .A2(\SB1_1_20/i0_4 ), .A3(
        \SB1_1_20/i1_7 ), .ZN(\SB1_1_20/Component_Function_1/NAND4_in[3] ) );
  CLKBUF_X4 U3475 ( .I(\SB1_1_13/buf_output[5] ), .Z(n1117) );
  CLKBUF_X2 U3479 ( .I(n2885), .Z(n4182) );
  NAND3_X1 U3482 ( .A1(\SB2_1_30/i1[9] ), .A2(\SB2_1_30/i0_4 ), .A3(
        \SB2_1_30/i1_5 ), .ZN(\SB2_1_30/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U3484 ( .A1(\SB2_1_26/i0_3 ), .A2(\SB2_1_26/i1_7 ), .A3(
        \SB2_1_26/i0[8] ), .ZN(\SB2_1_26/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 U3488 ( .A1(\SB2_1_30/i0_3 ), .A2(\SB2_1_30/i1[9] ), .ZN(
        \SB2_1_30/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U3496 ( .A1(\SB2_1_28/i0[6] ), .A2(\SB2_1_28/i1_5 ), .A3(
        \SB1_1_1/buf_output[0] ), .ZN(
        \SB2_1_28/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U3501 ( .A1(\SB1_1_14/buf_output[4] ), .A2(\SB2_1_13/i1_7 ), .A3(
        \SB2_1_13/i0[8] ), .ZN(n654) );
  NAND3_X1 U3505 ( .A1(\SB2_1_4/i0[7] ), .A2(\SB2_1_4/i0_3 ), .A3(
        \SB1_1_7/buf_output[2] ), .ZN(
        \SB2_1_4/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U3513 ( .A1(\SB2_1_5/i1[9] ), .A2(\SB2_1_5/i1_5 ), .A3(
        \SB1_1_6/buf_output[4] ), .ZN(
        \SB2_1_5/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U3523 ( .A1(\SB2_1_7/i3[0] ), .A2(\SB2_1_7/i0_0 ), .A3(
        \SB2_1_7/i1_7 ), .ZN(\SB2_1_7/Component_Function_4/NAND4_in[1] ) );
  NAND2_X1 U3525 ( .A1(\SB2_1_31/i0_3 ), .A2(\SB2_1_31/i1[9] ), .ZN(
        \SB2_1_31/Component_Function_1/NAND4_in[0] ) );
  INV_X1 U3535 ( .I(\MC_ARK_ARC_1_1/buf_output[0] ), .ZN(\SB1_2_31/i3[0] ) );
  INV_X1 U3543 ( .I(\MC_ARK_ARC_1_1/buf_output[115] ), .ZN(\SB1_2_12/i1_7 ) );
  CLKBUF_X4 U3549 ( .I(\MC_ARK_ARC_1_1/buf_output[178] ), .Z(\SB1_2_2/i0_4 )
         );
  NAND2_X1 U3555 ( .A1(\SB1_2_21/i0_3 ), .A2(\SB1_2_21/i1[9] ), .ZN(
        \SB1_2_21/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U3557 ( .A1(\SB1_2_20/i0_3 ), .A2(\SB1_2_20/i0[9] ), .A3(n2893), 
        .ZN(n4152) );
  NAND3_X1 U3561 ( .A1(\SB1_2_30/i0_0 ), .A2(\SB1_2_30/i0_3 ), .A3(
        \SB1_2_30/i0[7] ), .ZN(n4736) );
  NAND3_X1 U3568 ( .A1(\SB1_2_13/i0[10] ), .A2(\SB1_2_13/i1[9] ), .A3(
        \SB1_2_13/i1_5 ), .ZN(\SB1_2_13/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U3570 ( .A1(\SB1_2_6/i0[9] ), .A2(\SB1_2_6/i0_0 ), .A3(
        \SB1_2_6/i0[8] ), .ZN(\SB1_2_6/Component_Function_4/NAND4_in[0] ) );
  INV_X2 U3573 ( .I(\MC_ARK_ARC_1_1/buf_output[110] ), .ZN(\SB1_2_13/i1[9] )
         );
  NAND3_X1 U3580 ( .A1(\SB1_2_6/i0[8] ), .A2(\SB1_2_6/i0[7] ), .A3(
        \SB1_2_6/i0[6] ), .ZN(\SB1_2_6/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U3582 ( .A1(\SB1_2_29/i0[10] ), .A2(\SB1_2_29/i1[9] ), .A3(
        \SB1_2_29/i1_7 ), .ZN(\SB1_2_29/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U3595 ( .A1(\SB1_2_12/i0[6] ), .A2(\SB1_2_12/i0[8] ), .A3(
        \SB1_2_12/i0[7] ), .ZN(\SB1_2_12/Component_Function_0/NAND4_in[1] ) );
  INV_X1 U3600 ( .I(\SB1_2_20/buf_output[1] ), .ZN(\SB2_2_16/i1_7 ) );
  CLKBUF_X4 U3602 ( .I(\SB1_2_17/buf_output[1] ), .Z(\SB2_2_13/i0[6] ) );
  NAND3_X1 U3604 ( .A1(\SB2_2_6/i3[0] ), .A2(\SB2_2_6/i0_0 ), .A3(
        \SB2_2_6/i1_7 ), .ZN(\SB2_2_6/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U3607 ( .A1(n3333), .A2(\SB2_2_9/i0[6] ), .A3(\SB2_2_9/i0[8] ), 
        .ZN(n1620) );
  NAND3_X1 U3617 ( .A1(\SB2_2_7/i0[9] ), .A2(\SB2_2_7/i1_5 ), .A3(
        \SB2_2_7/i0[6] ), .ZN(\SB2_2_7/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U3623 ( .A1(\SB2_2_24/i1_5 ), .A2(\SB2_2_24/i0[10] ), .A3(
        \SB2_2_24/i1[9] ), .ZN(\SB2_2_24/Component_Function_2/NAND4_in[0] ) );
  CLKBUF_X4 U3626 ( .I(\SB1_2_23/buf_output[4] ), .Z(\SB2_2_22/i0_4 ) );
  CLKBUF_X4 U3628 ( .I(\SB1_2_21/buf_output[2] ), .Z(\SB2_2_18/i0_0 ) );
  NAND3_X1 U3629 ( .A1(\SB2_2_10/i0[8] ), .A2(\SB2_2_10/i0[7] ), .A3(
        \SB2_2_10/i0[6] ), .ZN(\SB2_2_10/Component_Function_0/NAND4_in[1] ) );
  CLKBUF_X4 U3632 ( .I(\SB2_2_7/buf_output[4] ), .Z(\RI5[2][154] ) );
  INV_X1 U3633 ( .I(\MC_ARK_ARC_1_2/buf_output[180] ), .ZN(\SB1_3_1/i3[0] ) );
  NAND3_X1 U3642 ( .A1(\SB1_3_8/i0[9] ), .A2(\SB1_3_8/i0_0 ), .A3(
        \SB1_3_8/i0[8] ), .ZN(\SB1_3_8/Component_Function_4/NAND4_in[0] ) );
  INV_X1 U3645 ( .I(\MC_ARK_ARC_1_2/buf_output[67] ), .ZN(\SB1_3_20/i1_7 ) );
  NAND3_X1 U3649 ( .A1(\SB1_3_19/i0[9] ), .A2(\SB1_3_19/i0_0 ), .A3(
        \SB1_3_19/i0[8] ), .ZN(\SB1_3_19/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U3651 ( .A1(\SB1_3_24/i0[8] ), .A2(\SB1_3_24/i3[0] ), .A3(
        \SB1_3_24/i1_5 ), .ZN(\SB1_3_24/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U3653 ( .A1(n3648), .A2(\SB1_3_11/i0_3 ), .A3(\SB1_3_11/i0_0 ), 
        .ZN(\SB1_3_11/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U3654 ( .A1(\SB1_3_13/i0_3 ), .A2(\SB1_3_13/i0[8] ), .A3(
        \SB1_3_13/i0[9] ), .ZN(\SB1_3_13/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3656 ( .A1(\SB1_3_20/i0[7] ), .A2(\SB1_3_20/i0_3 ), .A3(
        \SB1_3_20/i0_0 ), .ZN(\SB1_3_20/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U3665 ( .A1(\SB1_3_8/i0_4 ), .A2(\SB1_3_8/i0[8] ), .A3(
        \SB1_3_8/i1_7 ), .ZN(n3957) );
  NAND3_X1 U3669 ( .A1(\SB1_3_18/i0_0 ), .A2(\SB1_3_18/i1_7 ), .A3(
        \SB1_3_18/i3[0] ), .ZN(\SB1_3_18/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U3670 ( .A1(\SB1_3_16/i0_3 ), .A2(\SB1_3_16/i0[10] ), .A3(
        \SB1_3_16/i0[6] ), .ZN(\SB1_3_16/Component_Function_2/NAND4_in[1] ) );
  NAND2_X1 U3678 ( .A1(\SB1_3_9/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_3_9/Component_Function_4/NAND4_in[1] ), .ZN(n4698) );
  NAND3_X1 U3679 ( .A1(\SB1_3_24/i0_4 ), .A2(\SB1_3_24/i1[9] ), .A3(
        \SB1_3_24/i1_5 ), .ZN(n4577) );
  NAND3_X1 U3682 ( .A1(\SB1_3_21/i0_4 ), .A2(\SB1_3_21/i0[6] ), .A3(
        \SB1_3_21/i0[9] ), .ZN(n4072) );
  NAND2_X1 U3685 ( .A1(\SB1_3_1/Component_Function_4/NAND4_in[3] ), .A2(n4525), 
        .ZN(n737) );
  NAND2_X1 U3693 ( .A1(\SB2_3_2/i0_3 ), .A2(\SB2_3_2/i1[9] ), .ZN(
        \SB2_3_2/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U3703 ( .A1(n5490), .A2(\SB2_3_28/i1_5 ), .A3(n577), .ZN(n657) );
  NAND3_X1 U3706 ( .A1(n5491), .A2(\SB2_3_2/i0[7] ), .A3(\SB2_3_2/i0[6] ), 
        .ZN(\SB2_3_2/Component_Function_0/NAND4_in[1] ) );
  INV_X1 U3736 ( .I(\MC_ARK_ARC_1_3/buf_output[6] ), .ZN(\SB3_30/i3[0] ) );
  CLKBUF_X4 U3737 ( .I(\MC_ARK_ARC_1_3/buf_output[148] ), .Z(\SB3_7/i0_4 ) );
  BUF_X2 U3741 ( .I(\MC_ARK_ARC_1_3/buf_output[130] ), .Z(\SB3_10/i0_4 ) );
  NAND2_X1 U3747 ( .A1(\SB3_21/i0[10] ), .A2(\SB3_21/i0[9] ), .ZN(
        \SB3_21/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U3752 ( .A1(n4764), .A2(\SB3_27/i1_5 ), .A3(\SB3_27/i0_4 ), .ZN(
        \SB3_27/Component_Function_4/NAND4_in[3] ) );
  INV_X1 U3753 ( .I(\MC_ARK_ARC_1_3/buf_output[79] ), .ZN(\SB3_18/i1_7 ) );
  NAND3_X1 U3758 ( .A1(\SB3_29/i1[9] ), .A2(\SB3_29/i1_5 ), .A3(\SB3_29/i0_4 ), 
        .ZN(\SB3_29/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U3761 ( .A1(\SB3_28/i0_4 ), .A2(\SB3_28/i0[9] ), .A3(\SB3_28/i0[6] ), .ZN(n4511) );
  CLKBUF_X4 U3771 ( .I(\SB3_27/buf_output[2] ), .Z(\SB4_24/i0_0 ) );
  NAND3_X1 U3777 ( .A1(\SB4_1/i0[9] ), .A2(\SB4_1/i0[6] ), .A3(\SB4_1/i0_4 ), 
        .ZN(\SB4_1/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 U3778 ( .A1(\SB4_5/i0[10] ), .A2(\SB4_5/i0[9] ), .ZN(
        \SB4_5/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U3786 ( .A1(\SB4_5/i0[10] ), .A2(\SB4_5/i1[9] ), .A3(\SB4_5/i1_7 ), 
        .ZN(n3424) );
  NAND3_X1 U3789 ( .A1(\SB4_24/i1_5 ), .A2(\SB4_24/i0[6] ), .A3(\SB4_24/i0[9] ), .ZN(\SB4_24/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 U3796 ( .A1(\SB4_16/i0_3 ), .A2(\SB4_16/i1[9] ), .ZN(
        \SB4_16/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U3797 ( .A1(\SB4_17/i0_4 ), .A2(\SB4_17/i0[9] ), .A3(\SB4_17/i0[6] ), .ZN(n1695) );
  NAND3_X1 U3800 ( .A1(\SB4_1/i0_4 ), .A2(\SB4_1/i1_7 ), .A3(\SB4_1/i0[8] ), 
        .ZN(n4391) );
  NAND3_X1 U3802 ( .A1(\SB4_26/i1_5 ), .A2(\SB4_26/i0[6] ), .A3(\SB4_26/i0[9] ), .ZN(\SB4_26/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U3808 ( .A1(\SB4_5/i1_5 ), .A2(\SB4_5/i0[10] ), .A3(\SB4_5/i1[9] ), 
        .ZN(\SB4_5/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U3811 ( .A1(n3674), .A2(\SB4_20/i0[6] ), .A3(\SB4_20/i0[9] ), .ZN(
        \SB4_20/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U3819 ( .A1(\SB4_29/i3[0] ), .A2(\SB4_29/i0_0 ), .A3(\SB4_29/i1_7 ), 
        .ZN(\SB4_29/Component_Function_4/NAND4_in[1] ) );
  NAND2_X1 U3823 ( .A1(\SB4_17/i0[10] ), .A2(\SB4_17/i0[9] ), .ZN(
        \SB4_17/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 U3825 ( .A1(\SB4_22/i0[10] ), .A2(\SB4_22/i0[9] ), .ZN(
        \SB4_22/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U3831 ( .A1(\SB4_14/i1_5 ), .A2(\SB4_14/i0[6] ), .A3(\SB4_14/i0[9] ), .ZN(\SB4_14/Component_Function_1/NAND4_in[2] ) );
  BUF_X2 U3835 ( .I(\SB2_0_17/buf_output[0] ), .Z(n1375) );
  CLKBUF_X4 U3841 ( .I(\SB1_3_1/buf_output[5] ), .Z(\SB2_3_1/i0_3 ) );
  AND2_X1 U3847 ( .A1(\SB2_2_12/i1_7 ), .A2(\SB2_2_12/i0[8] ), .Z(n2901) );
  AND2_X1 U3848 ( .A1(\SB2_3_21/i0_3 ), .A2(\SB2_3_21/i0_0 ), .Z(n2903) );
  AND2_X1 U3849 ( .A1(\SB2_3_3/i1_7 ), .A2(\SB2_3_3/i0[8] ), .Z(n2904) );
  XNOR2_X1 U3850 ( .A1(\SB2_1_10/buf_output[2] ), .A2(n113), .ZN(n2905) );
  AND4_X2 U3852 ( .A1(\SB1_3_26/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_26/Component_Function_3/NAND4_in[1] ), .A3(n1838), .A4(n1760), 
        .Z(n2906) );
  XNOR2_X1 U3862 ( .A1(\MC_ARK_ARC_1_1/temp5[71] ), .A2(n4150), .ZN(n2909) );
  XNOR2_X1 U3863 ( .A1(\MC_ARK_ARC_1_3/temp5[167] ), .A2(
        \MC_ARK_ARC_1_3/temp6[167] ), .ZN(n2910) );
  NAND3_X2 U3868 ( .A1(\SB2_2_5/i0_3 ), .A2(\SB2_2_5/i0[9] ), .A3(
        \SB2_2_5/i0[8] ), .ZN(\SB2_2_5/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 U3869 ( .A1(n1161), .A2(\SB2_3_25/Component_Function_5/NAND4_in[3] ), .A3(n2940), .A4(\SB2_3_25/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_3_25/buf_output[5] ) );
  INV_X2 U3870 ( .I(\MC_ARK_ARC_1_1/buf_output[47] ), .ZN(n2913) );
  XOR2_X1 U3872 ( .A1(n5521), .A2(\RI5[1][111] ), .Z(
        \MC_ARK_ARC_1_1/temp3[45] ) );
  NAND3_X1 U3881 ( .A1(\SB3_10/i0[6] ), .A2(\SB3_10/i0[7] ), .A3(
        \SB3_10/i0[8] ), .ZN(\SB3_10/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U3886 ( .A1(\SB4_5/i0[9] ), .A2(\SB4_5/i0_4 ), .A3(\SB4_5/i0[6] ), 
        .ZN(n2914) );
  XOR2_X1 U3898 ( .A1(n1576), .A2(n2917), .Z(\MC_ARK_ARC_1_3/buf_output[127] )
         );
  XOR2_X1 U3899 ( .A1(\MC_ARK_ARC_1_3/temp3[127] ), .A2(
        \MC_ARK_ARC_1_3/temp4[127] ), .Z(n2917) );
  INV_X2 U3913 ( .I(\RI3[0][149] ), .ZN(\SB2_0_7/i1_5 ) );
  NAND4_X2 U3915 ( .A1(\SB1_0_7/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_7/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_0_7/Component_Function_5/NAND4_in[3] ), .A4(
        \SB1_0_7/Component_Function_5/NAND4_in[0] ), .ZN(\RI3[0][149] ) );
  NAND3_X2 U3928 ( .A1(\RI3[0][4] ), .A2(\SB2_0_31/i0_3 ), .A3(
        \SB2_0_31/i1[9] ), .ZN(n2920) );
  NAND3_X1 U3932 ( .A1(\SB1_0_0/i1_7 ), .A2(n404), .A3(\SB1_0_0/i0[8] ), .ZN(
        \SB1_0_0/Component_Function_1/NAND4_in[3] ) );
  XOR2_X1 U3933 ( .A1(n2924), .A2(\MC_ARK_ARC_1_1/temp2[145] ), .Z(
        \MC_ARK_ARC_1_1/temp5[145] ) );
  XOR2_X1 U3934 ( .A1(\RI5[1][145] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[139] ), 
        .Z(n2924) );
  XOR2_X1 U3937 ( .A1(\MC_ARK_ARC_1_3/temp4[29] ), .A2(n2925), .Z(
        \MC_ARK_ARC_1_3/temp6[29] ) );
  XOR2_X1 U3938 ( .A1(\RI5[3][131] ), .A2(\RI5[3][95] ), .Z(n2925) );
  XOR2_X1 U3943 ( .A1(\RI5[1][129] ), .A2(\RI5[1][135] ), .Z(n2927) );
  XOR2_X1 U3955 ( .A1(\RI5[2][32] ), .A2(\RI5[2][62] ), .Z(n2931) );
  XOR2_X1 U3971 ( .A1(n2935), .A2(n2934), .Z(\MC_ARK_ARC_1_1/temp5[17] ) );
  XOR2_X1 U3975 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[155] ), .A2(\RI5[1][11] ), 
        .Z(n2934) );
  XOR2_X1 U3977 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[179] ), .A2(\RI5[1][17] ), 
        .Z(n2935) );
  NAND3_X2 U3982 ( .A1(\SB2_1_25/i1[9] ), .A2(\SB2_1_25/i0_3 ), .A3(
        \SB2_1_25/i0[6] ), .ZN(\SB2_1_25/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U3987 ( .A1(\SB2_3_20/buf_output[2] ), .A2(n523), .Z(n2937) );
  XOR2_X1 U3990 ( .A1(\RI5[0][128] ), .A2(\RI5[0][104] ), .Z(n2846) );
  XOR2_X1 U3991 ( .A1(\MC_ARK_ARC_1_1/temp6[11] ), .A2(n2939), .Z(
        \MC_ARK_ARC_1_1/buf_output[11] ) );
  NAND4_X2 U3995 ( .A1(n2288), .A2(n2942), .A3(
        \SB2_1_25/Component_Function_5/NAND4_in[0] ), .A4(
        \SB2_1_25/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB2_1_25/buf_output[5] ) );
  NAND3_X2 U3996 ( .A1(\SB2_1_25/i0[6] ), .A2(\SB2_1_25/i0_0 ), .A3(
        \SB2_1_25/i0[10] ), .ZN(n2942) );
  BUF_X2 U3997 ( .I(\SB2_2_30/buf_output[2] ), .Z(n3677) );
  NAND3_X1 U3998 ( .A1(\SB2_0_1/i0_4 ), .A2(\RI3[0][180] ), .A3(
        \SB1_0_5/buf_output[1] ), .ZN(
        \SB2_0_1/Component_Function_5/NAND4_in[3] ) );
  XOR2_X1 U4000 ( .A1(n3741), .A2(n2943), .Z(\MC_ARK_ARC_1_0/buf_output[145] )
         );
  XOR2_X1 U4002 ( .A1(\MC_ARK_ARC_1_0/temp2[145] ), .A2(
        \MC_ARK_ARC_1_0/temp1[145] ), .Z(n2943) );
  NAND3_X2 U4012 ( .A1(\SB2_1_3/i0[6] ), .A2(n5208), .A3(\SB2_1_3/i0[9] ), 
        .ZN(n1421) );
  NAND3_X2 U4015 ( .A1(\SB2_0_28/i0_3 ), .A2(\SB2_0_28/i0[7] ), .A3(
        \SB2_0_28/i0_0 ), .ZN(n3893) );
  NAND3_X2 U4016 ( .A1(\SB1_2_17/i0[6] ), .A2(\SB1_2_17/i0[10] ), .A3(
        \SB1_2_17/i0_0 ), .ZN(\SB1_2_17/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U4017 ( .A1(\SB1_1_5/i0_4 ), .A2(\SB1_1_5/i0[9] ), .A3(
        \MC_ARK_ARC_1_0/buf_output[157] ), .ZN(
        \SB1_1_5/Component_Function_5/NAND4_in[3] ) );
  XOR2_X1 U4024 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[48] ), .A2(\RI5[0][84] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[174] ) );
  XOR2_X1 U4030 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[41] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[5] ), .Z(\MC_ARK_ARC_1_3/temp3[131] ) );
  XOR2_X1 U4031 ( .A1(\MC_ARK_ARC_1_0/temp5[160] ), .A2(n1255), .Z(
        \MC_ARK_ARC_1_0/buf_output[160] ) );
  XOR2_X1 U4032 ( .A1(\MC_ARK_ARC_1_3/temp2[59] ), .A2(n1522), .Z(
        \MC_ARK_ARC_1_3/temp5[59] ) );
  NAND3_X2 U4039 ( .A1(\SB2_1_1/i0[10] ), .A2(\SB2_1_1/i1_5 ), .A3(
        \SB2_1_1/i1[9] ), .ZN(\SB2_1_1/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U4041 ( .A1(n2948), .A2(n2947), .Z(\MC_ARK_ARC_1_3/temp5[95] ) );
  XOR2_X1 U4043 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[41] ), .A2(\RI5[3][95] ), 
        .Z(n2947) );
  XOR2_X1 U4044 ( .A1(\RI5[3][65] ), .A2(\RI5[3][89] ), .Z(n2948) );
  NAND4_X2 U4045 ( .A1(\SB1_0_6/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_0_6/Component_Function_1/NAND4_in[0] ), .A3(
        \SB1_0_6/Component_Function_1/NAND4_in[1] ), .A4(n2949), .ZN(
        \RI3[0][175] ) );
  NAND3_X2 U4046 ( .A1(\SB1_0_6/i0[6] ), .A2(\SB1_0_6/i1_5 ), .A3(
        \SB1_0_6/i0[9] ), .ZN(n2949) );
  INV_X2 U4051 ( .I(\SB1_2_3/buf_output[2] ), .ZN(\SB2_2_0/i1[9] ) );
  XOR2_X1 U4056 ( .A1(\MC_ARK_ARC_1_2/temp2[69] ), .A2(n2951), .Z(
        \MC_ARK_ARC_1_2/temp5[69] ) );
  NAND3_X1 U4071 ( .A1(\SB1_3_7/i0[10] ), .A2(\SB1_3_7/i1[9] ), .A3(
        \SB1_3_7/i1_5 ), .ZN(\SB1_3_7/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U4076 ( .A1(n3894), .A2(n3810), .Z(\MC_ARK_ARC_1_0/temp5[33] ) );
  AND2_X1 U4079 ( .A1(\SB1_1_1/buf_output[2] ), .A2(\SB1_1_0/buf_output[3] ), 
        .Z(n3857) );
  XOR2_X1 U4081 ( .A1(n3821), .A2(n2956), .Z(\MC_ARK_ARC_1_0/buf_output[191] )
         );
  XOR2_X1 U4082 ( .A1(\MC_ARK_ARC_1_0/temp3[191] ), .A2(
        \MC_ARK_ARC_1_0/temp4[191] ), .Z(n2956) );
  XOR2_X1 U4083 ( .A1(n3650), .A2(n215), .Z(n575) );
  BUF_X4 U4084 ( .I(\SB2_1_8/buf_output[2] ), .Z(\RI5[1][158] ) );
  NAND3_X1 U4092 ( .A1(\SB3_1/i0_4 ), .A2(\SB3_1/i0_3 ), .A3(n4765), .ZN(n2958) );
  BUF_X4 U4093 ( .I(\SB2_3_0/buf_output[4] ), .Z(\RI5[3][4] ) );
  INV_X2 U4111 ( .I(\SB3_5/buf_output[2] ), .ZN(\SB4_2/i1[9] ) );
  XOR2_X1 U4121 ( .A1(\MC_ARK_ARC_1_2/temp1[127] ), .A2(n2962), .Z(
        \MC_ARK_ARC_1_2/temp5[127] ) );
  XOR2_X1 U4122 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[97] ), .A2(\RI5[2][73] ), 
        .Z(n2962) );
  NAND4_X2 U4125 ( .A1(\SB3_3/Component_Function_2/NAND4_in[0] ), .A2(n2108), 
        .A3(n1687), .A4(\SB3_3/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB3_3/buf_output[2] ) );
  XOR2_X1 U4128 ( .A1(\RI5[3][162] ), .A2(\RI5[3][186] ), .Z(
        \MC_ARK_ARC_1_3/temp2[24] ) );
  XOR2_X1 U4130 ( .A1(\RI5[3][162] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[168] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[168] ) );
  NAND4_X2 U4136 ( .A1(\SB2_0_2/Component_Function_5/NAND4_in[1] ), .A2(
        \SB2_0_2/Component_Function_5/NAND4_in[2] ), .A3(
        \SB2_0_2/Component_Function_5/NAND4_in[0] ), .A4(n2964), .ZN(
        \SB2_0_2/buf_output[5] ) );
  XOR2_X1 U4138 ( .A1(n2965), .A2(n20), .Z(Ciphertext[132]) );
  NAND4_X2 U4142 ( .A1(\SB4_9/Component_Function_0/NAND4_in[3] ), .A2(
        \SB4_9/Component_Function_0/NAND4_in[2] ), .A3(
        \SB4_9/Component_Function_0/NAND4_in[1] ), .A4(n1913), .ZN(n2965) );
  XOR2_X1 U4156 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[185] ), .A2(\RI5[2][191] ), 
        .Z(n2967) );
  NAND3_X1 U4157 ( .A1(\SB2_2_15/i0_3 ), .A2(\SB2_2_15/i0[10] ), .A3(
        \SB2_2_15/i0_4 ), .ZN(\SB2_2_15/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 U4180 ( .A1(\SB2_2_7/i0[10] ), .A2(\SB2_2_7/i1_5 ), .A3(
        \SB2_2_7/i1[9] ), .ZN(n2970) );
  NAND3_X2 U4192 ( .A1(\SB1_2_1/i0[6] ), .A2(\SB1_2_1/i0[9] ), .A3(
        \SB1_2_1/i0_4 ), .ZN(n2972) );
  NAND4_X2 U4203 ( .A1(\SB1_0_1/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_0_1/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_1/Component_Function_5/NAND4_in[3] ), .A4(n3287), .ZN(
        \SB1_0_1/buf_output[5] ) );
  NAND3_X2 U4207 ( .A1(\SB1_1_17/i0[10] ), .A2(\SB1_1_17/i0_0 ), .A3(
        \SB1_1_17/i0[6] ), .ZN(\SB1_1_17/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U4210 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[67] ), .A2(\RI5[0][43] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[97] ) );
  NAND4_X2 U4212 ( .A1(\SB2_1_17/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_17/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_17/Component_Function_1/NAND4_in[3] ), .A4(n3745), .ZN(
        \SB2_1_17/buf_output[1] ) );
  NAND4_X2 U4213 ( .A1(\SB1_1_16/Component_Function_2/NAND4_in[1] ), .A2(n3860), .A3(n3423), .A4(n2973), .ZN(\RI3[1][110] ) );
  NAND4_X2 U4214 ( .A1(\SB2_3_8/Component_Function_2/NAND4_in[2] ), .A2(n1049), 
        .A3(\SB2_3_8/Component_Function_2/NAND4_in[1] ), .A4(n2974), .ZN(
        \SB2_3_8/buf_output[2] ) );
  NAND3_X2 U4215 ( .A1(n3669), .A2(\SB2_3_8/i0[10] ), .A3(\SB2_3_8/i1_5 ), 
        .ZN(n2974) );
  XOR2_X1 U4221 ( .A1(n2314), .A2(n2975), .Z(n1501) );
  XOR2_X1 U4222 ( .A1(\RI5[3][2] ), .A2(\RI5[3][8] ), .Z(n2975) );
  NAND3_X1 U4239 ( .A1(\SB1_0_6/i0_0 ), .A2(\SB1_0_6/i0[10] ), .A3(n321), .ZN(
        \SB1_0_6/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U4246 ( .A1(\SB4_10/i0[10] ), .A2(\SB4_10/i0[9] ), .A3(
        \SB4_10/i0_3 ), .ZN(\SB4_10/Component_Function_4/NAND4_in[2] ) );
  NAND4_X2 U4262 ( .A1(\SB1_0_16/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_0_16/Component_Function_4/NAND4_in[3] ), .A3(n2327), .A4(
        \SB1_0_16/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB1_0_16/buf_output[4] ) );
  NAND4_X2 U4268 ( .A1(n1815), .A2(\SB2_3_29/Component_Function_3/NAND4_in[2] ), .A3(\SB2_3_29/Component_Function_3/NAND4_in[0] ), .A4(
        \SB2_3_29/Component_Function_3/NAND4_in[1] ), .ZN(
        \SB2_3_29/buf_output[3] ) );
  XOR2_X1 U4277 ( .A1(n2979), .A2(\MC_ARK_ARC_1_3/temp6[108] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[108] ) );
  XOR2_X1 U4280 ( .A1(\MC_ARK_ARC_1_3/temp1[108] ), .A2(
        \MC_ARK_ARC_1_3/temp2[108] ), .Z(n2979) );
  XOR2_X1 U4293 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[122] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[158] ), .Z(n2983) );
  XOR2_X1 U4294 ( .A1(\MC_ARK_ARC_1_0/temp5[70] ), .A2(n2984), .Z(
        \MC_ARK_ARC_1_0/buf_output[70] ) );
  XOR2_X1 U4297 ( .A1(\MC_ARK_ARC_1_0/temp3[70] ), .A2(
        \MC_ARK_ARC_1_0/temp4[70] ), .Z(n2984) );
  INV_X2 U4299 ( .I(\SB1_1_26/buf_output[3] ), .ZN(\SB2_1_24/i0[8] ) );
  NAND4_X2 U4306 ( .A1(\SB1_1_26/Component_Function_3/NAND4_in[0] ), .A2(n4279), .A3(n1407), .A4(\SB1_1_26/Component_Function_3/NAND4_in[1] ), .ZN(
        \SB1_1_26/buf_output[3] ) );
  NAND3_X2 U4320 ( .A1(\SB2_2_27/i0[10] ), .A2(\SB2_2_27/i1_7 ), .A3(
        \SB2_2_27/i1[9] ), .ZN(n2985) );
  INV_X2 U4327 ( .I(\SB1_3_31/buf_output[3] ), .ZN(\SB2_3_29/i0[8] ) );
  XOR2_X1 U4340 ( .A1(n1796), .A2(\MC_ARK_ARC_1_3/temp1[121] ), .Z(n2987) );
  XOR2_X1 U4342 ( .A1(n2989), .A2(n2988), .Z(\MC_ARK_ARC_1_0/temp6[65] ) );
  XOR2_X1 U4343 ( .A1(\RI5[0][131] ), .A2(n172), .Z(n2988) );
  XOR2_X1 U4361 ( .A1(\MC_ARK_ARC_1_3/temp2[122] ), .A2(n2991), .Z(
        \MC_ARK_ARC_1_3/temp5[122] ) );
  XOR2_X1 U4364 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[116] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[122] ), .Z(n2991) );
  NOR2_X2 U4386 ( .A1(n2994), .A2(n4122), .ZN(n930) );
  NAND2_X1 U4387 ( .A1(\SB2_3_1/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_3_1/Component_Function_2/NAND4_in[3] ), .ZN(n2994) );
  XOR2_X1 U4388 ( .A1(\MC_ARK_ARC_1_3/temp2[14] ), .A2(n2995), .Z(
        \MC_ARK_ARC_1_3/temp5[14] ) );
  XOR2_X1 U4390 ( .A1(\RI5[3][8] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[14] ), 
        .Z(n2995) );
  NAND3_X2 U4395 ( .A1(\SB1_1_11/i0[10] ), .A2(\SB1_1_11/i1[9] ), .A3(
        \SB1_1_11/i1_7 ), .ZN(n2200) );
  NAND4_X2 U4398 ( .A1(\SB2_1_22/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_1_22/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_1_22/Component_Function_0/NAND4_in[0] ), .A4(n2997), .ZN(
        \SB2_1_22/buf_output[0] ) );
  NAND3_X2 U4403 ( .A1(\SB2_1_16/i0_3 ), .A2(\SB2_1_16/i0[9] ), .A3(
        \SB2_1_16/i0[8] ), .ZN(n2998) );
  XOR2_X1 U4407 ( .A1(\RI5[1][151] ), .A2(n496), .Z(n2999) );
  XOR2_X1 U4410 ( .A1(\RI5[1][61] ), .A2(\RI5[1][85] ), .Z(n3000) );
  NAND4_X2 U4412 ( .A1(\SB2_0_25/Component_Function_3/NAND4_in[2] ), .A2(n3517), .A3(\SB2_0_25/Component_Function_3/NAND4_in[0] ), .A4(n3001), .ZN(
        \SB2_0_25/buf_output[3] ) );
  NAND3_X2 U4418 ( .A1(\SB2_0_25/i0_0 ), .A2(\RI3[0][40] ), .A3(
        \SB2_0_25/i0_3 ), .ZN(n3001) );
  NAND4_X2 U4419 ( .A1(\SB2_1_25/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_1_25/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_1_25/Component_Function_1/NAND4_in[0] ), .A4(n3002), .ZN(
        \SB2_1_25/buf_output[1] ) );
  NAND4_X2 U4425 ( .A1(n4550), .A2(\SB1_1_21/Component_Function_3/NAND4_in[0] ), .A3(n3229), .A4(n3003), .ZN(\SB1_1_21/buf_output[3] ) );
  NAND3_X2 U4426 ( .A1(\SB1_1_21/i0[10] ), .A2(\SB1_1_21/i1_7 ), .A3(
        \SB1_1_21/i1[9] ), .ZN(n3003) );
  XOR2_X1 U4438 ( .A1(n3006), .A2(n3005), .Z(\MC_ARK_ARC_1_1/temp5[119] ) );
  XOR2_X1 U4446 ( .A1(\RI5[1][65] ), .A2(\RI5[1][119] ), .Z(n3005) );
  XOR2_X1 U4447 ( .A1(\RI5[1][113] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[89] ), 
        .Z(n3006) );
  NAND3_X2 U4454 ( .A1(\SB1_2_29/i0_4 ), .A2(\SB1_2_29/i1[9] ), .A3(
        \RI1[2][17] ), .ZN(\SB1_2_29/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U4457 ( .A1(\SB2_2_14/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_2_14/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_2_14/Component_Function_4/NAND4_in[0] ), .A4(n865), .ZN(
        \SB2_2_14/buf_output[4] ) );
  NAND4_X2 U4462 ( .A1(\SB1_0_28/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_0_28/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_0_28/Component_Function_1/NAND4_in[3] ), .A4(
        \SB1_0_28/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_0_28/buf_output[1] ) );
  XOR2_X1 U4469 ( .A1(n1365), .A2(\MC_ARK_ARC_1_3/buf_datainput[191] ), .Z(
        n3230) );
  XOR2_X1 U4478 ( .A1(n3008), .A2(n209), .Z(Ciphertext[126]) );
  XOR2_X1 U4485 ( .A1(\RI5[1][62] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[38] ), 
        .Z(n3010) );
  XOR2_X1 U4499 ( .A1(\RI5[1][77] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[41] ), 
        .Z(n3012) );
  INV_X2 U4503 ( .I(\SB1_0_6/buf_output[2] ), .ZN(\SB2_0_3/i1[9] ) );
  NAND3_X1 U4531 ( .A1(\SB4_24/i0[9] ), .A2(\SB4_24/i0[6] ), .A3(\SB4_24/i0_4 ), .ZN(n3015) );
  NAND3_X2 U4539 ( .A1(\SB2_0_3/i0_0 ), .A2(\SB2_0_3/i1_5 ), .A3(\RI3[0][172] ), .ZN(n3016) );
  INV_X1 U4540 ( .I(\SB3_29/buf_output[2] ), .ZN(\SB4_26/i1[9] ) );
  XOR2_X1 U4551 ( .A1(\MC_ARK_ARC_1_3/temp2[132] ), .A2(
        \MC_ARK_ARC_1_3/temp1[132] ), .Z(\MC_ARK_ARC_1_3/temp5[132] ) );
  NAND4_X2 U4552 ( .A1(\SB3_29/Component_Function_0/NAND4_in[3] ), .A2(
        \SB3_29/Component_Function_0/NAND4_in[2] ), .A3(
        \SB3_29/Component_Function_0/NAND4_in[1] ), .A4(
        \SB3_29/Component_Function_0/NAND4_in[0] ), .ZN(\SB3_29/buf_output[0] ) );
  NAND3_X2 U4554 ( .A1(\SB2_2_13/i0_0 ), .A2(n580), .A3(n1394), .ZN(n4591) );
  XOR2_X1 U4556 ( .A1(n3018), .A2(\MC_ARK_ARC_1_1/temp6[92] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[92] ) );
  XOR2_X1 U4558 ( .A1(\RI5[3][102] ), .A2(\RI5[3][78] ), .Z(
        \MC_ARK_ARC_1_3/temp2[132] ) );
  INV_X1 U4577 ( .I(\SB3_12/buf_output[4] ), .ZN(\SB4_11/i0[7] ) );
  XOR2_X1 U4580 ( .A1(\RI5[0][57] ), .A2(\RI5[0][63] ), .Z(
        \MC_ARK_ARC_1_0/temp1[63] ) );
  XOR2_X1 U4582 ( .A1(\SB2_1_17/buf_output[3] ), .A2(\RI5[1][93] ), .Z(
        \MC_ARK_ARC_1_1/temp1[99] ) );
  XOR2_X1 U4585 ( .A1(\MC_ARK_ARC_1_2/temp2[93] ), .A2(n3105), .Z(n3023) );
  NAND4_X2 U4604 ( .A1(\SB2_1_4/Component_Function_5/NAND4_in[2] ), .A2(n3512), 
        .A3(\SB2_1_4/Component_Function_5/NAND4_in[0] ), .A4(n3026), .ZN(
        \SB2_1_4/buf_output[5] ) );
  NAND3_X2 U4607 ( .A1(\SB2_1_4/i0[10] ), .A2(\SB2_1_4/i0[6] ), .A3(
        \SB1_1_7/buf_output[2] ), .ZN(n3026) );
  NAND3_X2 U4609 ( .A1(\SB1_1_3/i0[10] ), .A2(\SB1_1_3/i1[9] ), .A3(
        \SB1_1_3/i1_7 ), .ZN(\SB1_1_3/Component_Function_3/NAND4_in[2] ) );
  XOR2_X1 U4617 ( .A1(\MC_ARK_ARC_1_0/temp5[47] ), .A2(n3028), .Z(
        \MC_ARK_ARC_1_0/buf_output[47] ) );
  XOR2_X1 U4618 ( .A1(\MC_ARK_ARC_1_0/temp4[47] ), .A2(
        \MC_ARK_ARC_1_0/temp3[47] ), .Z(n3028) );
  XOR2_X1 U4634 ( .A1(\MC_ARK_ARC_1_1/temp6[134] ), .A2(n4708), .Z(
        \MC_ARK_ARC_1_1/buf_output[134] ) );
  NAND3_X1 U4638 ( .A1(\SB4_18/i0_4 ), .A2(\SB4_18/i1_7 ), .A3(n3662), .ZN(
        \SB4_18/Component_Function_1/NAND4_in[3] ) );
  XOR2_X1 U4642 ( .A1(n2106), .A2(n3742), .Z(\MC_ARK_ARC_1_2/buf_output[128] )
         );
  NAND4_X2 U4644 ( .A1(\SB1_1_17/Component_Function_5/NAND4_in[2] ), .A2(n3302), .A3(\SB1_1_17/Component_Function_5/NAND4_in[1] ), .A4(
        \SB1_1_17/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_17/buf_output[5] ) );
  XOR2_X1 U4645 ( .A1(\MC_ARK_ARC_1_3/temp5[74] ), .A2(
        \MC_ARK_ARC_1_3/temp6[74] ), .Z(\MC_ARK_ARC_1_3/buf_output[74] ) );
  NAND4_X2 U4652 ( .A1(\SB1_0_19/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_19/Component_Function_5/NAND4_in[3] ), .A3(n1330), .A4(
        \SB1_0_19/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_0_19/buf_output[5] ) );
  NAND3_X1 U4654 ( .A1(\SB3_19/i0_4 ), .A2(\SB3_19/i1[9] ), .A3(\SB3_19/i1_5 ), 
        .ZN(n3081) );
  NAND4_X2 U4655 ( .A1(\SB1_1_19/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_19/Component_Function_3/NAND4_in[1] ), .A3(n3702), .A4(
        \SB1_1_19/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_1_19/buf_output[3] ) );
  NAND3_X1 U4670 ( .A1(\SB1_2_14/i0[10] ), .A2(\SB1_2_14/i0_0 ), .A3(
        \SB1_2_14/i0[6] ), .ZN(\SB1_2_14/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U4673 ( .A1(\SB4_17/i0[10] ), .A2(\SB4_17/i1_7 ), .A3(
        \SB4_17/i1[9] ), .ZN(\SB4_17/Component_Function_3/NAND4_in[2] ) );
  NAND4_X1 U4675 ( .A1(n2412), .A2(\SB3_19/Component_Function_3/NAND4_in[0] ), 
        .A3(n4351), .A4(n4159), .ZN(\SB3_19/buf_output[3] ) );
  XOR2_X1 U4685 ( .A1(\MC_ARK_ARC_1_0/temp1[132] ), .A2(n3031), .Z(
        \MC_ARK_ARC_1_0/temp5[132] ) );
  XOR2_X1 U4691 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[78] ), .A2(\RI5[0][102] ), 
        .Z(n3031) );
  NAND3_X2 U4704 ( .A1(\SB2_1_17/i0[10] ), .A2(\SB2_1_17/i0_3 ), .A3(
        \SB2_1_17/i0[9] ), .ZN(n3334) );
  XOR2_X1 U4705 ( .A1(n3033), .A2(\MC_ARK_ARC_1_1/temp6[148] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[148] ) );
  XOR2_X1 U4709 ( .A1(\MC_ARK_ARC_1_1/temp1[148] ), .A2(
        \MC_ARK_ARC_1_1/temp2[148] ), .Z(n3033) );
  NAND4_X2 U4712 ( .A1(\SB2_0_23/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_0_23/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_0_23/Component_Function_0/NAND4_in[0] ), .A4(n3034), .ZN(
        \SB2_0_23/buf_output[0] ) );
  XOR2_X1 U4748 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[74] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[38] ), .Z(n3037) );
  NAND4_X2 U4758 ( .A1(\SB1_0_31/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_0_31/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_0_31/Component_Function_3/NAND4_in[3] ), .A4(n3040), .ZN(
        \SB1_0_31/buf_output[3] ) );
  NAND3_X2 U4759 ( .A1(\SB1_0_31/i0[10] ), .A2(\SB1_0_31/i1[9] ), .A3(
        \SB1_0_31/i1_7 ), .ZN(n3040) );
  NAND3_X2 U4767 ( .A1(\SB2_2_16/i0[10] ), .A2(\SB2_2_16/i0_0 ), .A3(
        \SB2_2_16/i0[6] ), .ZN(n3041) );
  XOR2_X1 U4769 ( .A1(\MC_ARK_ARC_1_0/temp6[183] ), .A2(n3042), .Z(
        \MC_ARK_ARC_1_0/buf_output[183] ) );
  NAND3_X1 U4790 ( .A1(\SB2_3_21/i3[0] ), .A2(\SB2_3_21/i1_5 ), .A3(
        \SB2_3_21/i0[8] ), .ZN(\SB2_3_21/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U4820 ( .A1(\SB1_1_6/i0[10] ), .A2(\SB1_1_6/i1[9] ), .A3(
        \SB1_1_6/i1_5 ), .ZN(\SB1_1_6/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U4825 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[146] ), .A2(\RI5[2][170] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[8] ) );
  INV_X2 U4840 ( .I(\SB3_27/buf_output[2] ), .ZN(\SB4_24/i1[9] ) );
  XOR2_X1 U4842 ( .A1(n1383), .A2(\RI5[1][69] ), .Z(n3050) );
  XOR2_X1 U4849 ( .A1(\RI5[3][20] ), .A2(\RI5[3][26] ), .Z(n3051) );
  NAND3_X1 U4853 ( .A1(\SB1_0_29/i0_4 ), .A2(\SB1_0_29/i0_0 ), .A3(
        \SB1_0_29/i0_3 ), .ZN(\SB1_0_29/Component_Function_3/NAND4_in[1] ) );
  INV_X2 U4858 ( .I(\SB1_0_4/buf_output[5] ), .ZN(\SB2_0_4/i1_5 ) );
  XOR2_X1 U4866 ( .A1(n2568), .A2(n3053), .Z(\RI1[3][89] ) );
  XOR2_X1 U4868 ( .A1(n4360), .A2(\MC_ARK_ARC_1_2/temp4[89] ), .Z(n3053) );
  NAND4_X2 U4871 ( .A1(\SB1_1_15/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_15/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_15/Component_Function_3/NAND4_in[2] ), .A4(n1203), .ZN(
        \SB1_1_15/buf_output[3] ) );
  NAND4_X2 U4876 ( .A1(n3999), .A2(n1490), .A3(
        \SB3_11/Component_Function_5/NAND4_in[0] ), .A4(
        \SB3_11/Component_Function_5/NAND4_in[2] ), .ZN(\SB3_11/buf_output[5] ) );
  NAND3_X1 U4947 ( .A1(\SB1_3_4/i0_0 ), .A2(\SB1_3_4/i1_7 ), .A3(
        \SB1_3_4/i3[0] ), .ZN(n3058) );
  NAND3_X2 U4952 ( .A1(\SB2_2_14/i0[7] ), .A2(\SB2_2_14/i0[6] ), .A3(
        \SB2_2_14/i0[8] ), .ZN(n649) );
  NAND3_X1 U4957 ( .A1(\SB2_3_8/i0[6] ), .A2(\SB2_3_8/i0[9] ), .A3(
        \SB2_3_8/i1_5 ), .ZN(n3059) );
  INV_X1 U4978 ( .I(\SB1_1_23/buf_output[0] ), .ZN(\SB2_1_18/i3[0] ) );
  NAND4_X2 U4979 ( .A1(\SB1_1_23/Component_Function_0/NAND4_in[2] ), .A2(n3124), .A3(\SB1_1_23/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_1_23/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_1_23/buf_output[0] ) );
  XOR2_X1 U4980 ( .A1(\MC_ARK_ARC_1_2/temp3[66] ), .A2(
        \MC_ARK_ARC_1_2/temp4[66] ), .Z(\MC_ARK_ARC_1_2/temp6[66] ) );
  XOR2_X1 U5015 ( .A1(n3065), .A2(n103), .Z(Ciphertext[37]) );
  NAND4_X2 U5018 ( .A1(n3887), .A2(\SB4_25/Component_Function_1/NAND4_in[3] ), 
        .A3(\SB4_25/Component_Function_1/NAND4_in[1] ), .A4(n2063), .ZN(n3065)
         );
  NAND4_X2 U5034 ( .A1(\SB3_12/Component_Function_2/NAND4_in[1] ), .A2(
        \SB3_12/Component_Function_2/NAND4_in[0] ), .A3(
        \SB3_12/Component_Function_2/NAND4_in[2] ), .A4(n3066), .ZN(
        \SB3_12/buf_output[2] ) );
  NAND3_X2 U5035 ( .A1(\SB3_12/i0_0 ), .A2(\SB3_12/i1_5 ), .A3(\SB3_12/i0_4 ), 
        .ZN(n3066) );
  NOR2_X2 U5039 ( .A1(n1117), .A2(\SB1_1_15/buf_output[3] ), .ZN(n1752) );
  INV_X2 U5051 ( .I(\SB1_3_20/buf_output[5] ), .ZN(\SB2_3_20/i1_5 ) );
  XOR2_X1 U5061 ( .A1(n4033), .A2(n3069), .Z(\MC_ARK_ARC_1_2/buf_output[122] )
         );
  NAND4_X2 U5064 ( .A1(\SB2_2_15/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_2_15/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_2_15/Component_Function_4/NAND4_in[1] ), .A4(n3070), .ZN(
        \SB2_2_15/buf_output[4] ) );
  NAND3_X1 U5065 ( .A1(\SB2_2_15/i0_3 ), .A2(\SB2_2_15/i0[9] ), .A3(
        \SB2_2_15/i0[10] ), .ZN(n3070) );
  XOR2_X1 U5066 ( .A1(n3071), .A2(n211), .Z(Ciphertext[66]) );
  NAND4_X2 U5069 ( .A1(\SB4_20/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_20/Component_Function_0/NAND4_in[3] ), .A3(
        \SB4_20/Component_Function_0/NAND4_in[1] ), .A4(
        \SB4_20/Component_Function_0/NAND4_in[0] ), .ZN(n3071) );
  NAND3_X2 U5070 ( .A1(\SB2_2_14/i0[9] ), .A2(\SB2_2_14/i0_4 ), .A3(
        \SB2_2_14/i0[6] ), .ZN(\SB2_2_14/Component_Function_5/NAND4_in[3] ) );
  XOR2_X1 U5073 ( .A1(\MC_ARK_ARC_1_0/temp2[27] ), .A2(n3072), .Z(
        \MC_ARK_ARC_1_0/temp5[27] ) );
  XOR2_X1 U5074 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[21] ), .A2(\RI5[0][27] ), 
        .Z(n3072) );
  XOR2_X1 U5085 ( .A1(\MC_ARK_ARC_1_2/temp5[27] ), .A2(n3073), .Z(
        \MC_ARK_ARC_1_2/buf_output[27] ) );
  XOR2_X1 U5086 ( .A1(\MC_ARK_ARC_1_2/temp4[27] ), .A2(
        \MC_ARK_ARC_1_2/temp3[27] ), .Z(n3073) );
  XOR2_X1 U5098 ( .A1(\RI5[1][177] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[153] ), 
        .Z(n1645) );
  XOR2_X1 U5116 ( .A1(n4504), .A2(n3076), .Z(\MC_ARK_ARC_1_0/temp5[155] ) );
  XOR2_X1 U5117 ( .A1(\RI5[0][101] ), .A2(\RI5[0][125] ), .Z(n3076) );
  NAND3_X1 U5123 ( .A1(\SB1_0_1/i0_3 ), .A2(\SB1_0_1/i0[8] ), .A3(
        \SB1_0_1/i1_7 ), .ZN(\SB1_0_1/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U5136 ( .A1(\SB2_3_26/i0[6] ), .A2(\SB1_3_31/buf_output[0] ), .A3(
        \SB2_3_26/i0_4 ), .ZN(\SB2_3_26/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 U5143 ( .A1(\SB2_1_20/i0_0 ), .A2(\SB2_1_20/i0_3 ), .A3(
        \SB2_1_20/i0_4 ), .ZN(n3079) );
  NAND4_X2 U5147 ( .A1(\SB2_1_14/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_1_14/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_1_14/Component_Function_3/NAND4_in[2] ), .A4(n3080), .ZN(
        \SB2_1_14/buf_output[3] ) );
  NAND4_X2 U5148 ( .A1(\SB3_19/Component_Function_4/NAND4_in[2] ), .A2(
        \SB3_19/Component_Function_4/NAND4_in[0] ), .A3(
        \SB3_19/Component_Function_4/NAND4_in[1] ), .A4(n3081), .ZN(
        \SB3_19/buf_output[4] ) );
  XOR2_X1 U5155 ( .A1(\RI5[0][70] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[76] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[76] ) );
  NAND3_X1 U5169 ( .A1(\SB3_7/i0[6] ), .A2(\SB3_7/i0[7] ), .A3(\SB3_7/i0[8] ), 
        .ZN(\SB3_7/Component_Function_0/NAND4_in[1] ) );
  NAND4_X2 U5176 ( .A1(n1701), .A2(\SB2_0_12/Component_Function_5/NAND4_in[1] ), .A3(\SB2_0_12/Component_Function_5/NAND4_in[0] ), .A4(n3089), .ZN(
        \SB2_0_12/buf_output[5] ) );
  NAND3_X2 U5177 ( .A1(\SB2_2_28/i0[10] ), .A2(\SB2_2_28/i0_3 ), .A3(
        \SB2_2_28/i0_4 ), .ZN(\SB2_2_28/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U5180 ( .A1(\MC_ARK_ARC_1_0/temp2[9] ), .A2(n3090), .Z(
        \MC_ARK_ARC_1_0/temp5[9] ) );
  XOR2_X1 U5187 ( .A1(\RI5[0][9] ), .A2(\RI5[0][3] ), .Z(n3090) );
  NAND3_X1 U5201 ( .A1(\SB1_0_29/i0_0 ), .A2(\SB1_0_29/i0[9] ), .A3(
        \SB1_0_29/i0[8] ), .ZN(n3092) );
  NAND3_X1 U5203 ( .A1(\SB4_4/i0_3 ), .A2(\SB3_7/buf_output[2] ), .A3(
        \SB4_4/i0[7] ), .ZN(\SB4_4/Component_Function_0/NAND4_in[3] ) );
  XOR2_X1 U5216 ( .A1(n838), .A2(\MC_ARK_ARC_1_2/temp3[163] ), .Z(n3097) );
  XOR2_X1 U5221 ( .A1(\RI5[0][35] ), .A2(\RI5[0][11] ), .Z(n3113) );
  NAND3_X2 U5227 ( .A1(\SB2_0_30/i0[10] ), .A2(\SB2_0_30/i1[9] ), .A3(
        \SB2_0_30/i1_5 ), .ZN(n3098) );
  NAND4_X2 U5229 ( .A1(\SB2_3_16/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_3_16/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_3_16/Component_Function_0/NAND4_in[2] ), .A4(n3099), .ZN(
        \SB2_3_16/buf_output[0] ) );
  NAND2_X1 U5230 ( .A1(\SB2_3_16/i0[9] ), .A2(\SB2_3_16/i0[10] ), .ZN(n3099)
         );
  XOR2_X1 U5231 ( .A1(\MC_ARK_ARC_1_2/temp4[107] ), .A2(n3100), .Z(n2609) );
  XOR2_X1 U5232 ( .A1(\RI5[2][173] ), .A2(\RI5[2][17] ), .Z(n3100) );
  NAND3_X2 U5233 ( .A1(\SB2_2_13/i0[10] ), .A2(n1394), .A3(\SB2_2_13/i1[9] ), 
        .ZN(n1610) );
  XOR2_X1 U5234 ( .A1(n3102), .A2(n3101), .Z(n1280) );
  XOR2_X1 U5235 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[80] ), .A2(\RI5[1][26] ), 
        .Z(n3101) );
  NAND3_X2 U5263 ( .A1(\SB2_3_12/i0[10] ), .A2(\SB2_3_12/i1[9] ), .A3(
        \SB2_3_12/i1_7 ), .ZN(\SB2_3_12/Component_Function_3/NAND4_in[2] ) );
  XOR2_X1 U5269 ( .A1(\MC_ARK_ARC_1_2/temp2[25] ), .A2(n3109), .Z(
        \MC_ARK_ARC_1_2/temp5[25] ) );
  XOR2_X1 U5270 ( .A1(\RI5[2][19] ), .A2(\RI5[2][25] ), .Z(n3109) );
  NAND3_X2 U5272 ( .A1(\SB2_2_0/i0_3 ), .A2(\SB2_2_0/i0_0 ), .A3(
        \SB2_2_0/i0_4 ), .ZN(\SB2_2_0/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U5276 ( .A1(n2867), .A2(\SB3_30/Component_Function_5/NAND4_in[1] ), 
        .A3(\SB3_30/Component_Function_5/NAND4_in[0] ), .A4(n3110), .ZN(
        \SB3_30/buf_output[5] ) );
  NAND3_X2 U5278 ( .A1(\SB3_30/i0_4 ), .A2(\SB3_30/i0[9] ), .A3(\SB3_30/i0[6] ), .ZN(n3110) );
  NAND3_X2 U5289 ( .A1(\SB1_0_31/i0_4 ), .A2(\SB1_0_31/i0_3 ), .A3(
        \SB1_0_31/i1[9] ), .ZN(\SB1_0_31/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U5293 ( .A1(\SB2_0_14/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_0_14/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_0_14/Component_Function_2/NAND4_in[1] ), .A4(
        \SB2_0_14/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_0_14/buf_output[2] ) );
  XOR2_X1 U5296 ( .A1(\RI5[3][112] ), .A2(\RI5[3][76] ), .Z(
        \MC_ARK_ARC_1_3/temp3[10] ) );
  NAND4_X2 U5318 ( .A1(\SB1_1_7/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_1_7/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_1_7/Component_Function_5/NAND4_in[3] ), .A4(
        \SB1_1_7/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_7/buf_output[5] ) );
  NAND3_X1 U5321 ( .A1(\SB2_2_28/i0[6] ), .A2(\SB2_2_28/i0[8] ), .A3(
        \SB2_2_28/i0[7] ), .ZN(\SB2_2_28/Component_Function_0/NAND4_in[1] ) );
  NOR2_X2 U5328 ( .A1(n3852), .A2(n1071), .ZN(\SB2_2_28/i0[7] ) );
  XOR2_X1 U5332 ( .A1(n3112), .A2(n201), .Z(Ciphertext[30]) );
  XOR2_X1 U5334 ( .A1(n3113), .A2(n3114), .Z(n3727) );
  XOR2_X1 U5335 ( .A1(\RI5[0][59] ), .A2(\RI5[0][65] ), .Z(n3114) );
  NAND3_X1 U5349 ( .A1(\SB4_11/i0_4 ), .A2(\SB4_11/i0[6] ), .A3(\SB4_11/i0[9] ), .ZN(n3127) );
  NAND3_X2 U5350 ( .A1(\SB1_2_15/i0_4 ), .A2(\SB1_2_15/i0_3 ), .A3(
        \SB1_2_15/i1[9] ), .ZN(n3118) );
  NOR2_X2 U5351 ( .A1(n3120), .A2(n3119), .ZN(n3669) );
  NAND3_X2 U5353 ( .A1(\SB1_3_11/i0[10] ), .A2(n2908), .A3(\SB1_3_11/i1[9] ), 
        .ZN(\SB1_3_11/Component_Function_2/NAND4_in[0] ) );
  NAND2_X1 U5354 ( .A1(\SB1_3_11/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_11/Component_Function_2/NAND4_in[2] ), .ZN(n3120) );
  NAND4_X2 U5363 ( .A1(\SB2_0_25/Component_Function_2/NAND4_in[0] ), .A2(n1550), .A3(n4008), .A4(\SB2_0_25/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB2_0_25/buf_output[2] ) );
  NAND3_X1 U5379 ( .A1(\SB1_1_27/i0_0 ), .A2(\SB1_1_27/i0_4 ), .A3(
        \SB1_1_27/i1_5 ), .ZN(n3128) );
  XOR2_X1 U5380 ( .A1(\RI5[3][33] ), .A2(\RI5[3][9] ), .Z(
        \MC_ARK_ARC_1_3/temp2[63] ) );
  BUF_X2 U5387 ( .I(\MC_ARK_ARC_1_0/buf_output[60] ), .Z(n3131) );
  INV_X2 U5394 ( .I(\SB1_3_22/buf_output[3] ), .ZN(\SB2_3_20/i0[8] ) );
  NAND4_X2 U5395 ( .A1(\SB1_3_22/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_22/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_22/Component_Function_3/NAND4_in[2] ), .A4(n3364), .ZN(
        \SB1_3_22/buf_output[3] ) );
  XOR2_X1 U5402 ( .A1(\RI5[0][126] ), .A2(\RI5[0][162] ), .Z(
        \MC_ARK_ARC_1_0/temp3[60] ) );
  XOR2_X1 U5405 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[124] ), .A2(\RI5[2][160] ), 
        .Z(n3132) );
  XOR2_X1 U5407 ( .A1(\RI5[0][116] ), .A2(\RI5[0][80] ), .Z(
        \MC_ARK_ARC_1_0/temp3[14] ) );
  NAND4_X2 U5410 ( .A1(\SB2_1_17/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_1_17/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_1_17/Component_Function_0/NAND4_in[3] ), .A4(n3134), .ZN(
        \SB2_1_17/buf_output[0] ) );
  NAND2_X1 U5412 ( .A1(\SB2_1_17/i0[10] ), .A2(\SB2_1_17/i0[9] ), .ZN(n3134)
         );
  NAND2_X1 U5417 ( .A1(\SB1_3_27/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_3_27/Component_Function_4/NAND4_in[3] ), .ZN(n2243) );
  NAND3_X1 U5422 ( .A1(\SB4_25/i0[10] ), .A2(\SB4_25/i1_5 ), .A3(
        \SB4_25/i1[9] ), .ZN(n3137) );
  BUF_X4 U5426 ( .I(\SB1_1_25/buf_output[5] ), .Z(\SB2_1_25/i0_3 ) );
  NAND3_X1 U5427 ( .A1(\SB3_19/i0[10] ), .A2(\SB3_19/i1_7 ), .A3(
        \SB3_19/i1[9] ), .ZN(n2412) );
  NAND4_X2 U5430 ( .A1(\SB2_3_27/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_3_27/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_27/Component_Function_1/NAND4_in[0] ), .A4(n3140), .ZN(
        \SB2_3_27/buf_output[1] ) );
  NAND3_X2 U5440 ( .A1(\SB2_0_29/i0[8] ), .A2(\SB2_0_29/i0_3 ), .A3(n2605), 
        .ZN(n3141) );
  NAND3_X1 U5446 ( .A1(\SB4_8/i0_0 ), .A2(\SB4_8/i1_5 ), .A3(\SB4_8/i0_4 ), 
        .ZN(\SB4_8/Component_Function_2/NAND4_in[3] ) );
  XOR2_X1 U5452 ( .A1(n3144), .A2(n3143), .Z(n833) );
  XOR2_X1 U5453 ( .A1(\RI5[0][89] ), .A2(\RI5[0][119] ), .Z(n3143) );
  XOR2_X1 U5454 ( .A1(\RI5[0][65] ), .A2(\RI5[0][113] ), .Z(n3144) );
  AND2_X1 U5457 ( .A1(n3938), .A2(\SB2_1_8/Component_Function_1/NAND4_in[1] ), 
        .Z(n3145) );
  INV_X4 U5461 ( .I(\SB2_0_7/i0[7] ), .ZN(\SB1_0_8/buf_output[4] ) );
  NAND3_X1 U5462 ( .A1(n2593), .A2(\SB2_0_7/i0[8] ), .A3(n6113), .ZN(
        \SB2_0_7/Component_Function_0/NAND4_in[1] ) );
  NOR2_X2 U5463 ( .A1(n3148), .A2(n3147), .ZN(\SB2_0_7/i0[7] ) );
  NAND2_X1 U5471 ( .A1(\SB1_0_8/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_0_8/Component_Function_4/NAND4_in[1] ), .ZN(n3148) );
  XOR2_X1 U5472 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[132] ), .A2(\RI5[2][138] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[138] ) );
  XOR2_X1 U5479 ( .A1(\RI5[1][116] ), .A2(\RI5[1][122] ), .Z(n3149) );
  NAND4_X2 U5489 ( .A1(\SB2_2_7/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_2_7/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_7/Component_Function_0/NAND4_in[0] ), .A4(n3154), .ZN(
        \SB2_2_7/buf_output[0] ) );
  NAND3_X1 U5494 ( .A1(\SB2_2_7/i0_0 ), .A2(\SB2_2_7/i0_3 ), .A3(
        \SB2_2_7/i0[7] ), .ZN(n3154) );
  NAND4_X2 U5501 ( .A1(\SB1_0_12/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_0_12/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_0_12/Component_Function_0/NAND4_in[1] ), .A4(n3155), .ZN(
        \SB1_0_12/buf_output[0] ) );
  NAND4_X2 U5514 ( .A1(\SB3_2/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_2/Component_Function_4/NAND4_in[3] ), .A3(n3481), .A4(n3157), 
        .ZN(\SB3_2/buf_output[4] ) );
  NAND3_X1 U5518 ( .A1(\SB3_2/i0_0 ), .A2(\SB3_2/i1_7 ), .A3(\SB3_2/i3[0] ), 
        .ZN(n3157) );
  NAND3_X1 U5523 ( .A1(\SB4_0/i0_4 ), .A2(\SB4_0/i1_5 ), .A3(
        \SB3_3/buf_output[2] ), .ZN(n3173) );
  XOR2_X1 U5525 ( .A1(n2390), .A2(n3158), .Z(\MC_ARK_ARC_1_1/buf_output[46] )
         );
  NAND2_X2 U5528 ( .A1(n3366), .A2(n2725), .ZN(n2883) );
  NAND3_X2 U5531 ( .A1(\SB2_3_13/i0_3 ), .A2(\SB2_3_13/i1[9] ), .A3(
        \SB1_3_14/buf_output[4] ), .ZN(n2794) );
  XOR2_X1 U5549 ( .A1(\RI5[2][145] ), .A2(\RI5[2][139] ), .Z(
        \MC_ARK_ARC_1_2/temp1[145] ) );
  NAND2_X2 U5550 ( .A1(n2894), .A2(n1488), .ZN(\RI5[2][139] ) );
  NAND3_X1 U5554 ( .A1(\SB2_3_13/i0_3 ), .A2(\SB2_3_13/i0[10] ), .A3(
        \SB1_3_14/buf_output[4] ), .ZN(n3162) );
  NAND4_X2 U5559 ( .A1(\SB1_1_28/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_28/Component_Function_3/NAND4_in[2] ), .A3(n3267), .A4(n846), 
        .ZN(\SB1_1_28/buf_output[3] ) );
  NAND3_X2 U5561 ( .A1(\SB1_2_10/i0[9] ), .A2(\SB1_2_10/i0[8] ), .A3(
        \SB1_2_10/i0_3 ), .ZN(\SB1_2_10/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U5569 ( .A1(\SB2_3_16/i0_3 ), .A2(\SB2_3_16/i0_0 ), .A3(
        \SB2_3_16/i0[7] ), .ZN(\SB2_3_16/Component_Function_0/NAND4_in[3] ) );
  XOR2_X1 U5573 ( .A1(\RI5[0][134] ), .A2(\RI5[0][98] ), .Z(
        \MC_ARK_ARC_1_0/temp3[32] ) );
  XOR2_X1 U5577 ( .A1(\MC_ARK_ARC_1_2/temp3[88] ), .A2(
        \MC_ARK_ARC_1_2/temp4[88] ), .Z(\MC_ARK_ARC_1_2/temp6[88] ) );
  NAND4_X2 U5585 ( .A1(\SB1_0_6/Component_Function_5/NAND4_in[1] ), .A2(n1969), 
        .A3(\SB1_0_6/Component_Function_5/NAND4_in[0] ), .A4(
        \SB1_0_6/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB1_0_6/buf_output[5] ) );
  NAND4_X2 U5590 ( .A1(\SB1_3_26/Component_Function_2/NAND4_in[1] ), .A2(n3931), .A3(n4467), .A4(n3165), .ZN(\SB1_3_26/buf_output[2] ) );
  NAND3_X1 U5592 ( .A1(\SB1_2_13/i0_0 ), .A2(\SB1_2_13/i0[8] ), .A3(
        \SB1_2_13/i0[9] ), .ZN(\SB1_2_13/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U5597 ( .A1(\SB2_3_24/i3[0] ), .A2(n2906), .A3(\SB2_3_24/i1_5 ), 
        .ZN(n1835) );
  XOR2_X1 U5604 ( .A1(\RI5[2][164] ), .A2(\RI5[2][8] ), .Z(n3166) );
  NAND4_X2 U5610 ( .A1(n2712), .A2(\SB1_3_29/Component_Function_5/NAND4_in[1] ), .A3(n4104), .A4(\SB1_3_29/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_29/buf_output[5] ) );
  XOR2_X1 U5623 ( .A1(\RI5[0][188] ), .A2(\RI5[0][164] ), .Z(n3168) );
  XOR2_X1 U5630 ( .A1(\RI5[2][33] ), .A2(\RI5[2][57] ), .Z(n4236) );
  NAND3_X1 U5639 ( .A1(\SB2_0_13/i0_0 ), .A2(\RI3[0][113] ), .A3(n2711), .ZN(
        n3171) );
  XOR2_X1 U5641 ( .A1(n3172), .A2(n64), .Z(Ciphertext[87]) );
  NAND3_X1 U5644 ( .A1(\SB4_9/i0[10] ), .A2(\SB4_9/i1_7 ), .A3(\SB4_9/i1[9] ), 
        .ZN(n3922) );
  INV_X1 U5645 ( .I(\SB1_1_3/buf_output[5] ), .ZN(\SB2_1_3/i1_5 ) );
  NAND4_X2 U5647 ( .A1(\SB1_1_3/Component_Function_5/NAND4_in[1] ), .A2(n1524), 
        .A3(\SB1_1_3/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_1_3/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_3/buf_output[5] ) );
  NAND3_X1 U5656 ( .A1(\SB4_8/i0_0 ), .A2(\SB4_8/i0_3 ), .A3(\SB4_8/i0[7] ), 
        .ZN(\SB4_8/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U5668 ( .A1(\SB4_22/i0_3 ), .A2(\SB4_22/i0[10] ), .A3(\SB4_22/i0_4 ), .ZN(\SB4_22/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U5675 ( .A1(\RI5[3][57] ), .A2(\RI5[3][63] ), .Z(n3177) );
  INV_X1 U5680 ( .I(\SB1_3_13/buf_output[1] ), .ZN(\SB2_3_9/i1_7 ) );
  NAND4_X2 U5681 ( .A1(\SB1_3_13/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_3_13/Component_Function_1/NAND4_in[0] ), .A3(
        \SB1_3_13/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_13/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_3_13/buf_output[1] ) );
  NAND3_X1 U5697 ( .A1(\SB4_22/i0_3 ), .A2(\SB4_22/i0[10] ), .A3(
        \SB4_22/i0[9] ), .ZN(n2808) );
  NAND4_X2 U5698 ( .A1(\SB2_3_20/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_20/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_3_20/Component_Function_5/NAND4_in[0] ), .A4(n3178), .ZN(
        \SB2_3_20/buf_output[5] ) );
  NAND3_X2 U5700 ( .A1(\SB2_3_20/i0[6] ), .A2(\SB2_3_20/i0_4 ), .A3(
        \SB2_3_20/i0[9] ), .ZN(n3178) );
  XOR2_X1 U5702 ( .A1(n3179), .A2(n192), .Z(Ciphertext[85]) );
  NAND3_X1 U5708 ( .A1(\SB3_22/i0[6] ), .A2(\SB3_22/i0[8] ), .A3(
        \SB3_22/i0[7] ), .ZN(\SB3_22/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U5717 ( .A1(\RI5[2][103] ), .A2(\RI5[2][79] ), .Z(
        \MC_ARK_ARC_1_2/temp2[133] ) );
  NAND3_X1 U5722 ( .A1(\SB4_4/i0_3 ), .A2(\SB4_4/i0[10] ), .A3(\SB4_4/i0[9] ), 
        .ZN(n3180) );
  XOR2_X1 U5737 ( .A1(\MC_ARK_ARC_1_1/temp1[141] ), .A2(n3183), .Z(
        \MC_ARK_ARC_1_1/temp5[141] ) );
  XOR2_X1 U5738 ( .A1(\RI5[1][111] ), .A2(\RI5[1][87] ), .Z(n3183) );
  NAND3_X1 U5742 ( .A1(\SB2_3_9/i0_3 ), .A2(\SB2_3_9/i0[10] ), .A3(
        \SB2_3_9/i0_4 ), .ZN(n3184) );
  NAND3_X2 U5747 ( .A1(\SB1_1_0/i1_7 ), .A2(\SB1_1_0/i0[10] ), .A3(
        \SB1_1_0/i1[9] ), .ZN(n2599) );
  XOR2_X1 U5765 ( .A1(\MC_ARK_ARC_1_3/temp3[126] ), .A2(
        \MC_ARK_ARC_1_3/temp4[126] ), .Z(\MC_ARK_ARC_1_3/temp6[126] ) );
  INV_X2 U5769 ( .I(\SB1_0_16/buf_output[2] ), .ZN(\SB2_0_13/i1[9] ) );
  XOR2_X1 U5778 ( .A1(n4119), .A2(\MC_ARK_ARC_1_1/temp2[77] ), .Z(n3189) );
  NAND3_X1 U5781 ( .A1(\SB4_14/i0[10] ), .A2(\SB4_14/i1_5 ), .A3(
        \SB4_14/i1[9] ), .ZN(n3190) );
  XOR2_X1 U5801 ( .A1(n3196), .A2(n3195), .Z(\MC_ARK_ARC_1_2/temp5[5] ) );
  XOR2_X1 U5802 ( .A1(\RI5[2][191] ), .A2(\RI5[2][5] ), .Z(n3195) );
  NAND3_X2 U5815 ( .A1(\SB2_2_0/i0_3 ), .A2(\SB2_2_0/i1[9] ), .A3(
        \SB2_2_0/i0_4 ), .ZN(\SB2_2_0/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U5846 ( .A1(\RI5[1][47] ), .A2(\RI5[1][53] ), .Z(
        \MC_ARK_ARC_1_1/temp1[53] ) );
  XOR2_X1 U5849 ( .A1(\RI5[1][45] ), .A2(\RI5[1][51] ), .Z(
        \MC_ARK_ARC_1_1/temp1[51] ) );
  XOR2_X1 U5850 ( .A1(n3202), .A2(n2255), .Z(n2827) );
  XOR2_X1 U5851 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[165] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[141] ), .Z(n3202) );
  NAND2_X1 U5858 ( .A1(\SB4_12/i0_0 ), .A2(\SB4_12/i3[0] ), .ZN(n3203) );
  XOR2_X1 U5891 ( .A1(\RI5[0][52] ), .A2(\RI5[0][58] ), .Z(
        \MC_ARK_ARC_1_0/temp1[58] ) );
  NAND4_X2 U5905 ( .A1(\SB2_0_6/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_0_6/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_0_6/Component_Function_2/NAND4_in[0] ), .A4(n4079), .ZN(
        \SB2_0_6/buf_output[2] ) );
  XOR2_X1 U5919 ( .A1(\MC_ARK_ARC_1_3/temp4[60] ), .A2(
        \MC_ARK_ARC_1_3/temp3[60] ), .Z(\MC_ARK_ARC_1_3/temp6[60] ) );
  NAND3_X1 U5922 ( .A1(\SB4_30/i0[6] ), .A2(n5525), .A3(\SB4_30/i0[9] ), .ZN(
        \SB4_30/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 U5923 ( .A1(\SB1_2_29/Component_Function_4/NAND4_in[2] ), .A2(n2257), .ZN(n3852) );
  NAND4_X2 U5925 ( .A1(\SB2_2_7/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_7/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_2_7/Component_Function_3/NAND4_in[1] ), .A4(n3207), .ZN(
        \SB2_2_7/buf_output[3] ) );
  XOR2_X1 U5927 ( .A1(n3208), .A2(n25), .Z(Ciphertext[170]) );
  NAND4_X2 U5932 ( .A1(\SB4_3/Component_Function_2/NAND4_in[0] ), .A2(n3228), 
        .A3(n2126), .A4(\SB4_3/Component_Function_2/NAND4_in[2] ), .ZN(n3208)
         );
  NAND4_X2 U5937 ( .A1(\SB2_3_18/Component_Function_2/NAND4_in[0] ), .A2(n1590), .A3(\SB2_3_18/Component_Function_2/NAND4_in[1] ), .A4(n3209), .ZN(
        \SB2_3_18/buf_output[2] ) );
  NAND3_X2 U5939 ( .A1(\SB2_3_18/i0_0 ), .A2(\SB2_3_18/i1_5 ), .A3(
        \SB2_3_18/i0_4 ), .ZN(n3209) );
  XOR2_X1 U5951 ( .A1(n3212), .A2(n3211), .Z(\MC_ARK_ARC_1_3/temp6[91] ) );
  XOR2_X1 U5952 ( .A1(\RI5[3][1] ), .A2(n177), .Z(n3211) );
  XOR2_X1 U5953 ( .A1(\RI5[3][157] ), .A2(\RI5[3][127] ), .Z(n3212) );
  XOR2_X1 U5956 ( .A1(\MC_ARK_ARC_1_0/temp4[174] ), .A2(
        \MC_ARK_ARC_1_0/temp3[174] ), .Z(n3213) );
  BUF_X4 U5957 ( .I(\SB2_3_7/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[174] ) );
  XOR2_X1 U5965 ( .A1(n3215), .A2(n3214), .Z(\MC_ARK_ARC_1_0/buf_output[52] )
         );
  XOR2_X1 U5966 ( .A1(\MC_ARK_ARC_1_0/temp3[52] ), .A2(
        \MC_ARK_ARC_1_0/temp4[52] ), .Z(n3214) );
  NAND3_X2 U5990 ( .A1(\SB2_2_24/i0_4 ), .A2(\SB2_2_24/i0[9] ), .A3(
        \SB2_2_24/i0[6] ), .ZN(\SB2_2_24/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 U6011 ( .A1(\SB2_3_13/i0_3 ), .A2(\SB2_3_13/i0[10] ), .A3(
        \SB2_3_13/i0[6] ), .ZN(n3236) );
  NAND3_X1 U6019 ( .A1(\SB1_2_4/i0_0 ), .A2(\SB1_2_4/i1_7 ), .A3(
        \SB1_2_4/i3[0] ), .ZN(n3219) );
  XOR2_X1 U6023 ( .A1(n3220), .A2(n1284), .Z(\MC_ARK_ARC_1_2/buf_output[112] )
         );
  XOR2_X1 U6024 ( .A1(n4440), .A2(\MC_ARK_ARC_1_2/temp2[112] ), .Z(n3220) );
  INV_X2 U6025 ( .I(\SB1_3_13/buf_output[3] ), .ZN(\SB2_3_11/i0[8] ) );
  NAND4_X2 U6026 ( .A1(\SB1_3_13/Component_Function_3/NAND4_in[2] ), .A2(n841), 
        .A3(\SB1_3_13/Component_Function_3/NAND4_in[0] ), .A4(n1426), .ZN(
        \SB1_3_13/buf_output[3] ) );
  NAND3_X1 U6046 ( .A1(\SB3_19/i0[10] ), .A2(\SB3_19/i0_3 ), .A3(
        \SB3_19/i0[9] ), .ZN(\SB3_19/Component_Function_4/NAND4_in[2] ) );
  NAND4_X2 U6047 ( .A1(\SB2_2_26/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_2_26/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_2_26/Component_Function_4/NAND4_in[1] ), .A4(n3222), .ZN(
        \SB2_2_26/buf_output[4] ) );
  NAND3_X1 U6048 ( .A1(\SB2_2_26/i0_4 ), .A2(\SB2_2_26/i1_5 ), .A3(
        \SB2_2_26/i1[9] ), .ZN(n3222) );
  XOR2_X1 U6053 ( .A1(n4190), .A2(\MC_ARK_ARC_1_2/temp3[111] ), .Z(n4421) );
  NAND3_X1 U6057 ( .A1(\SB4_23/i0_4 ), .A2(\SB4_23/i1_5 ), .A3(\SB4_23/i1[9] ), 
        .ZN(n3224) );
  NAND4_X2 U6064 ( .A1(n4566), .A2(\SB3_26/Component_Function_2/NAND4_in[2] ), 
        .A3(n1842), .A4(\SB3_26/Component_Function_2/NAND4_in[0] ), .ZN(
        \SB3_26/buf_output[2] ) );
  NAND3_X2 U6071 ( .A1(n4625), .A2(\SB2_1_21/i1_5 ), .A3(\SB2_1_21/i0[8] ), 
        .ZN(n3227) );
  INV_X2 U6072 ( .I(\SB1_0_20/buf_output[5] ), .ZN(\SB2_0_20/i1_5 ) );
  NAND4_X2 U6074 ( .A1(\SB1_0_20/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_20/Component_Function_5/NAND4_in[0] ), .A3(n804), .A4(
        \SB1_0_20/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB1_0_20/buf_output[5] ) );
  NAND3_X1 U6081 ( .A1(\SB3_5/buf_output[3] ), .A2(\SB4_3/i0_3 ), .A3(
        \SB4_3/i0[6] ), .ZN(n3228) );
  XOR2_X1 U6088 ( .A1(\MC_ARK_ARC_1_1/temp1[93] ), .A2(
        \MC_ARK_ARC_1_1/temp2[93] ), .Z(n4584) );
  XOR2_X1 U6093 ( .A1(\MC_ARK_ARC_1_3/temp1[92] ), .A2(
        \MC_ARK_ARC_1_3/temp4[92] ), .Z(n4232) );
  XOR2_X1 U6097 ( .A1(n3233), .A2(n3232), .Z(\MC_ARK_ARC_1_2/temp6[170] ) );
  XOR2_X1 U6099 ( .A1(\RI5[2][80] ), .A2(n243), .Z(n3232) );
  XOR2_X1 U6103 ( .A1(\RI5[2][44] ), .A2(n570), .Z(n3233) );
  XOR2_X1 U6104 ( .A1(\MC_ARK_ARC_1_0/temp4[159] ), .A2(
        \MC_ARK_ARC_1_0/temp3[159] ), .Z(n2512) );
  NAND3_X1 U6117 ( .A1(\SB2_0_4/i0[7] ), .A2(\SB2_0_4/i0[6] ), .A3(
        \SB2_0_4/i0[8] ), .ZN(\SB2_0_4/Component_Function_0/NAND4_in[1] ) );
  NAND3_X2 U6118 ( .A1(\SB2_3_0/i1[9] ), .A2(\SB2_3_0/i0_3 ), .A3(
        \SB2_3_0/i0[6] ), .ZN(\SB2_3_0/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 U6124 ( .I(\MC_ARK_ARC_1_1/buf_output[83] ), .Z(\SB1_2_18/i0_3 ) );
  BUF_X2 U6127 ( .I(\SB2_3_13/buf_output[3] ), .Z(\RI5[3][123] ) );
  INV_X2 U6128 ( .I(\SB1_3_14/buf_output[2] ), .ZN(\SB2_3_11/i1[9] ) );
  INV_X2 U6141 ( .I(\MC_ARK_ARC_1_1/buf_output[83] ), .ZN(\SB1_2_18/i1_5 ) );
  XOR2_X1 U6142 ( .A1(n3240), .A2(n3239), .Z(n3350) );
  XOR2_X1 U6143 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[59] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[95] ), .Z(n3239) );
  XOR2_X1 U6145 ( .A1(\RI5[2][143] ), .A2(\RI5[2][23] ), .Z(n3240) );
  XOR2_X1 U6162 ( .A1(\MC_ARK_ARC_1_0/temp4[21] ), .A2(n3243), .Z(n2837) );
  XOR2_X1 U6163 ( .A1(\RI5[0][123] ), .A2(\RI5[0][87] ), .Z(n3243) );
  XOR2_X1 U6176 ( .A1(\MC_ARK_ARC_1_2/temp3[130] ), .A2(
        \MC_ARK_ARC_1_2/temp4[130] ), .Z(n4639) );
  NAND3_X1 U6177 ( .A1(\SB2_2_10/i1[9] ), .A2(n581), .A3(\SB2_2_10/i1_5 ), 
        .ZN(\SB2_2_10/Component_Function_4/NAND4_in[3] ) );
  XOR2_X1 U6178 ( .A1(\MC_ARK_ARC_1_0/temp2[68] ), .A2(n3247), .Z(
        \MC_ARK_ARC_1_0/temp5[68] ) );
  NAND3_X1 U6190 ( .A1(\SB4_15/i0_3 ), .A2(\SB4_15/i0[9] ), .A3(\SB4_15/i0[8] ), .ZN(n3248) );
  XOR2_X1 U6195 ( .A1(n3249), .A2(n128), .Z(Ciphertext[26]) );
  XOR2_X1 U6198 ( .A1(\RI5[1][32] ), .A2(\RI5[1][158] ), .Z(n4111) );
  XOR2_X1 U6199 ( .A1(\MC_ARK_ARC_1_3/temp1[112] ), .A2(n3251), .Z(
        \MC_ARK_ARC_1_3/temp5[112] ) );
  XOR2_X1 U6200 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[82] ), .A2(\RI5[3][58] ), 
        .Z(n3251) );
  XOR2_X1 U6208 ( .A1(n1042), .A2(\MC_ARK_ARC_1_2/temp5[91] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[91] ) );
  NAND4_X2 U6209 ( .A1(\SB1_0_16/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_16/Component_Function_3/NAND4_in[1] ), .A3(n4539), .A4(
        \SB1_0_16/Component_Function_3/NAND4_in[2] ), .ZN(
        \SB1_0_16/buf_output[3] ) );
  XOR2_X1 U6212 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[101] ), .A2(\RI5[1][107] ), 
        .Z(n3903) );
  NAND3_X1 U6213 ( .A1(\SB2_1_3/i0[10] ), .A2(\SB2_1_3/i1_5 ), .A3(
        \SB2_1_3/i1[9] ), .ZN(\SB2_1_3/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U6214 ( .A1(\SB2_3_30/i0[6] ), .A2(\SB2_3_30/i0[7] ), .A3(
        \SB2_3_30/i0[8] ), .ZN(\SB2_3_30/Component_Function_0/NAND4_in[1] ) );
  NAND3_X2 U6217 ( .A1(\SB1_1_23/i0_3 ), .A2(\SB1_1_23/i0[6] ), .A3(
        \SB1_1_23/i1[9] ), .ZN(\SB1_1_23/Component_Function_3/NAND4_in[0] ) );
  INV_X2 U6226 ( .I(\SB1_2_10/buf_output[2] ), .ZN(\SB2_2_7/i1[9] ) );
  XOR2_X1 U6234 ( .A1(n3256), .A2(n3255), .Z(\MC_ARK_ARC_1_3/temp6[101] ) );
  XOR2_X1 U6235 ( .A1(n1365), .A2(n134), .Z(n3255) );
  XOR2_X1 U6236 ( .A1(\RI5[3][11] ), .A2(\RI5[3][137] ), .Z(n3256) );
  NAND4_X2 U6237 ( .A1(\SB1_0_24/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_24/Component_Function_5/NAND4_in[2] ), .A3(n1205), .A4(
        \SB1_0_24/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_0_24/buf_output[5] ) );
  NAND3_X1 U6241 ( .A1(\SB3_18/i0[10] ), .A2(\SB3_18/i1[9] ), .A3(
        \SB3_18/i1_5 ), .ZN(\SB3_18/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U6244 ( .A1(\SB2_2_7/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_7/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_7/Component_Function_5/NAND4_in[0] ), .A4(
        \SB2_2_7/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB2_2_7/buf_output[5] ) );
  XOR2_X1 U6257 ( .A1(\MC_ARK_ARC_1_3/temp5[79] ), .A2(n3258), .Z(
        \MC_ARK_ARC_1_3/buf_output[79] ) );
  XOR2_X1 U6258 ( .A1(\MC_ARK_ARC_1_3/temp3[79] ), .A2(
        \MC_ARK_ARC_1_3/temp4[79] ), .Z(n3258) );
  NAND4_X2 U6263 ( .A1(\SB1_3_5/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_3_5/Component_Function_1/NAND4_in[1] ), .A3(n2185), .A4(
        \SB1_3_5/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_3_5/buf_output[1] ) );
  XOR2_X1 U6264 ( .A1(n2690), .A2(n4569), .Z(\MC_ARK_ARC_1_2/buf_output[153] )
         );
  NAND3_X1 U6266 ( .A1(\SB1_0_16/i0_3 ), .A2(\SB1_0_16/i0[10] ), .A3(n4752), 
        .ZN(\SB1_0_16/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U6269 ( .A1(n3261), .A2(n3260), .Z(\MC_ARK_ARC_1_3/buf_output[45] )
         );
  XOR2_X1 U6270 ( .A1(\MC_ARK_ARC_1_3/temp3[45] ), .A2(
        \MC_ARK_ARC_1_3/temp4[45] ), .Z(n3260) );
  XOR2_X1 U6273 ( .A1(\MC_ARK_ARC_1_3/temp1[45] ), .A2(
        \MC_ARK_ARC_1_3/temp2[45] ), .Z(n3261) );
  NAND3_X2 U6278 ( .A1(\SB2_2_26/i0_4 ), .A2(\SB2_2_26/i0_3 ), .A3(
        \SB2_2_26/i1[9] ), .ZN(\SB2_2_26/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U6289 ( .A1(\SB1_3_6/i0[10] ), .A2(\SB1_3_6/i1[9] ), .A3(
        \SB1_3_6/i1_7 ), .ZN(n3262) );
  XOR2_X1 U6292 ( .A1(\MC_ARK_ARC_1_2/temp1[15] ), .A2(n3263), .Z(
        \MC_ARK_ARC_1_2/temp5[15] ) );
  XOR2_X1 U6293 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[177] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[153] ), .Z(n3263) );
  NAND3_X1 U6311 ( .A1(\SB4_28/i0[6] ), .A2(n5514), .A3(\SB4_28/i0_3 ), .ZN(
        n3266) );
  XOR2_X1 U6313 ( .A1(\SB2_0_9/buf_output[3] ), .A2(\RI5[0][123] ), .Z(
        \MC_ARK_ARC_1_0/temp2[177] ) );
  NAND3_X2 U6319 ( .A1(\SB1_1_28/i0_0 ), .A2(\SB1_1_28/i0_3 ), .A3(
        \SB1_1_28/i0_4 ), .ZN(n3267) );
  NAND3_X2 U6328 ( .A1(\SB2_2_0/i0_3 ), .A2(\SB2_2_0/i0[10] ), .A3(
        \SB2_2_0/i0_4 ), .ZN(n3269) );
  NAND4_X2 U6329 ( .A1(\SB1_2_13/Component_Function_4/NAND4_in[0] ), .A2(n3510), .A3(\SB1_2_13/Component_Function_4/NAND4_in[3] ), .A4(
        \SB1_2_13/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB1_2_13/buf_output[4] ) );
  XOR2_X1 U6332 ( .A1(\RI5[2][37] ), .A2(\RI5[2][73] ), .Z(
        \MC_ARK_ARC_1_2/temp3[163] ) );
  INV_X2 U6340 ( .I(\MC_ARK_ARC_1_0/buf_output[143] ), .ZN(n3270) );
  NAND2_X2 U6341 ( .A1(\SB1_1_16/i0_0 ), .A2(\SB1_1_16/i3[0] ), .ZN(
        \SB1_1_16/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U6342 ( .A1(\SB3_31/i0[9] ), .A2(\SB3_31/i0_4 ), .A3(\SB3_31/i0[6] ), .ZN(\SB3_31/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 U6356 ( .A1(\SB4_27/i0[9] ), .A2(\SB4_27/i0[10] ), .ZN(n3271) );
  INV_X2 U6366 ( .I(\SB1_2_9/buf_output[2] ), .ZN(\SB2_2_6/i1[9] ) );
  NAND4_X2 U6368 ( .A1(\SB1_2_9/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_2_9/Component_Function_2/NAND4_in[2] ), .A3(n3317), .A4(n4108), 
        .ZN(\SB1_2_9/buf_output[2] ) );
  XOR2_X1 U6378 ( .A1(\MC_ARK_ARC_1_3/temp6[67] ), .A2(n4027), .Z(
        \MC_ARK_ARC_1_3/buf_output[67] ) );
  NAND3_X2 U6379 ( .A1(\SB2_2_9/i0[10] ), .A2(n3687), .A3(\SB2_2_9/i1[9] ), 
        .ZN(\SB2_2_9/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U6385 ( .A1(n3276), .A2(n3964), .Z(\MC_ARK_ARC_1_0/buf_output[188] )
         );
  XOR2_X1 U6391 ( .A1(\RI5[0][174] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[138] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[72] ) );
  NAND3_X2 U6396 ( .A1(\SB1_2_19/i0_4 ), .A2(\SB1_2_19/i0_3 ), .A3(
        \SB1_2_19/i1[9] ), .ZN(n3277) );
  NOR2_X2 U6397 ( .A1(n4141), .A2(n3278), .ZN(n2806) );
  XOR2_X1 U6401 ( .A1(\RI5[1][93] ), .A2(\RI5[1][69] ), .Z(
        \MC_ARK_ARC_1_1/temp2[123] ) );
  AOI21_X2 U6402 ( .A1(n3280), .A2(n3279), .B(\SB2_3_1/i1_5 ), .ZN(n4122) );
  NAND4_X2 U6418 ( .A1(\SB1_0_7/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_7/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_7/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_0_7/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_0_7/buf_output[3] ) );
  NAND3_X2 U6420 ( .A1(\SB1_0_23/i0[6] ), .A2(\SB1_0_23/i0[10] ), .A3(
        \SB1_0_23/i0_3 ), .ZN(n3642) );
  NAND3_X2 U6436 ( .A1(\SB2_2_12/i0_4 ), .A2(\SB2_2_12/i0_3 ), .A3(
        \SB2_2_12/i1[9] ), .ZN(n3283) );
  XOR2_X1 U6439 ( .A1(\MC_ARK_ARC_1_2/temp6[53] ), .A2(n1834), .Z(
        \MC_ARK_ARC_1_2/buf_output[53] ) );
  XOR2_X1 U6441 ( .A1(n3744), .A2(\MC_ARK_ARC_1_1/temp3[115] ), .Z(n3285) );
  XOR2_X1 U6442 ( .A1(\SB2_0_6/buf_output[3] ), .A2(\RI5[0][129] ), .Z(
        \MC_ARK_ARC_1_0/temp3[63] ) );
  NAND3_X2 U6444 ( .A1(\SB1_3_31/i0[6] ), .A2(\SB1_3_31/i0_0 ), .A3(
        \SB1_3_31/i0[10] ), .ZN(\SB1_3_31/Component_Function_5/NAND4_in[1] )
         );
  NAND4_X2 U6445 ( .A1(\SB1_3_23/Component_Function_5/NAND4_in[3] ), .A2(
        \SB1_3_23/Component_Function_5/NAND4_in[1] ), .A3(n4398), .A4(
        \SB1_3_23/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_23/buf_output[5] ) );
  NAND4_X2 U6457 ( .A1(\SB1_2_2/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_2/Component_Function_2/NAND4_in[2] ), .A3(n4437), .A4(
        \SB1_2_2/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB1_2_2/buf_output[2] ) );
  XOR2_X1 U6465 ( .A1(\RI5[2][5] ), .A2(\RI5[2][11] ), .Z(
        \MC_ARK_ARC_1_2/temp1[11] ) );
  NAND4_X2 U6469 ( .A1(\SB1_3_0/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_0/Component_Function_2/NAND4_in[2] ), .A3(
        \SB1_3_0/Component_Function_2/NAND4_in[1] ), .A4(n3286), .ZN(
        \SB1_3_0/buf_output[2] ) );
  NAND3_X2 U6470 ( .A1(\SB1_3_0/i0_0 ), .A2(\SB1_3_0/i0_4 ), .A3(
        \SB1_3_0/i1_5 ), .ZN(n3286) );
  NAND4_X2 U6472 ( .A1(\SB1_0_17/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_0_17/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_0_17/Component_Function_0/NAND4_in[0] ), .A4(
        \SB1_0_17/Component_Function_0/NAND4_in[2] ), .ZN(\RI3[0][114] ) );
  XOR2_X1 U6474 ( .A1(\RI5[1][44] ), .A2(\RI5[1][20] ), .Z(n3393) );
  NAND4_X2 U6477 ( .A1(\SB2_1_27/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_27/Component_Function_2/NAND4_in[2] ), .A3(n3840), .A4(n2283), 
        .ZN(\SB2_1_27/buf_output[2] ) );
  NAND3_X2 U6482 ( .A1(\SB2_1_17/i0[6] ), .A2(\SB2_1_17/i0[9] ), .A3(
        \SB2_1_17/i1_5 ), .ZN(n3745) );
  NAND4_X2 U6489 ( .A1(\SB2_0_6/Component_Function_5/NAND4_in[3] ), .A2(
        \SB2_0_6/Component_Function_5/NAND4_in[1] ), .A3(n3883), .A4(
        \SB2_0_6/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_0_6/buf_output[5] ) );
  NAND3_X1 U6492 ( .A1(\SB3_1/i0_0 ), .A2(\SB3_1/i0[9] ), .A3(\SB3_1/i0[8] ), 
        .ZN(\SB3_1/Component_Function_4/NAND4_in[0] ) );
  NAND2_X2 U6493 ( .A1(\SB1_0_1/i0_0 ), .A2(\SB1_0_1/i3[0] ), .ZN(n3287) );
  NAND3_X2 U6495 ( .A1(\SB2_1_27/i0[9] ), .A2(\SB2_1_27/i0_4 ), .A3(
        \SB2_1_27/i0[6] ), .ZN(\SB2_1_27/Component_Function_5/NAND4_in[3] ) );
  XOR2_X1 U6497 ( .A1(n3288), .A2(\MC_ARK_ARC_1_0/temp1[48] ), .Z(
        \MC_ARK_ARC_1_0/temp5[48] ) );
  XOR2_X1 U6504 ( .A1(\RI5[0][18] ), .A2(\RI5[0][186] ), .Z(n3288) );
  NAND4_X2 U6506 ( .A1(\SB2_0_1/Component_Function_0/NAND4_in[0] ), .A2(n2536), 
        .A3(\SB2_0_1/Component_Function_0/NAND4_in[2] ), .A4(n3289), .ZN(
        \SB2_0_1/buf_output[0] ) );
  NAND4_X2 U6511 ( .A1(\SB1_0_4/Component_Function_5/NAND4_in[3] ), .A2(
        \SB1_0_4/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_4/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_0_4/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_0_4/buf_output[5] ) );
  NAND4_X2 U6515 ( .A1(\SB2_3_19/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_3_19/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_3_19/Component_Function_4/NAND4_in[3] ), .A4(n3291), .ZN(
        \SB2_3_19/buf_output[4] ) );
  NAND3_X1 U6517 ( .A1(\SB3_29/i0_0 ), .A2(\SB3_29/i0_3 ), .A3(\SB3_29/i0[7] ), 
        .ZN(\SB3_29/Component_Function_0/NAND4_in[3] ) );
  NAND4_X2 U6518 ( .A1(\SB2_2_6/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_2_6/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_2_6/Component_Function_0/NAND4_in[0] ), .A4(n3292), .ZN(
        \SB2_2_6/buf_output[0] ) );
  XOR2_X1 U6522 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[56] ), .A2(n211), .Z(n3293) );
  XOR2_X1 U6525 ( .A1(\RI5[0][182] ), .A2(\RI5[0][20] ), .Z(n3294) );
  XOR2_X1 U6529 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[186] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[30] ), .Z(\MC_ARK_ARC_1_2/temp3[120] )
         );
  XOR2_X1 U6530 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[152] ), .A2(\RI5[3][146] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[152] ) );
  NAND4_X2 U6532 ( .A1(\SB1_0_25/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_0_25/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_0_25/Component_Function_5/NAND4_in[0] ), .A4(n2204), .ZN(
        \SB1_0_25/buf_output[5] ) );
  NOR2_X2 U6537 ( .A1(n4175), .A2(n4247), .ZN(n1396) );
  NAND4_X2 U6538 ( .A1(\SB3_1/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_1/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_1/Component_Function_0/NAND4_in[0] ), .A4(n3295), .ZN(
        \SB3_1/buf_output[0] ) );
  XOR2_X1 U6563 ( .A1(\RI5[1][5] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[29] ), 
        .Z(n3300) );
  XOR2_X1 U6580 ( .A1(\MC_ARK_ARC_1_2/temp1[10] ), .A2(n3303), .Z(
        \MC_ARK_ARC_1_2/temp5[10] ) );
  XOR2_X1 U6582 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[148] ), .A2(\RI5[2][172] ), 
        .Z(n3303) );
  XOR2_X1 U6607 ( .A1(\MC_ARK_ARC_1_1/temp3[191] ), .A2(n3305), .Z(n3344) );
  XOR2_X1 U6611 ( .A1(\RI5[1][161] ), .A2(\RI5[1][191] ), .Z(n3305) );
  XOR2_X1 U6612 ( .A1(n3306), .A2(\MC_ARK_ARC_1_1/temp4[17] ), .Z(n2391) );
  XOR2_X1 U6616 ( .A1(\RI5[1][83] ), .A2(\RI5[1][119] ), .Z(n3306) );
  NAND4_X2 U6617 ( .A1(n2576), .A2(n1312), .A3(n4692), .A4(n1076), .ZN(
        \SB2_3_18/buf_output[5] ) );
  INV_X1 U6619 ( .I(\RI3[0][5] ), .ZN(\SB2_0_31/i1_5 ) );
  NAND4_X2 U6620 ( .A1(\SB1_0_31/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_31/Component_Function_5/NAND4_in[2] ), .A3(n2180), .A4(
        \SB1_0_31/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[0][5] ) );
  XOR2_X1 U6621 ( .A1(\MC_ARK_ARC_1_1/temp5[87] ), .A2(n3307), .Z(
        \MC_ARK_ARC_1_1/buf_output[87] ) );
  XOR2_X1 U6627 ( .A1(n4210), .A2(\MC_ARK_ARC_1_1/temp4[87] ), .Z(n3307) );
  NAND3_X2 U6636 ( .A1(\SB2_0_0/i0_0 ), .A2(\RI3[0][190] ), .A3(\SB2_0_0/i1_5 ), .ZN(\SB2_0_0/Component_Function_2/NAND4_in[3] ) );
  XOR2_X1 U6639 ( .A1(\RI5[0][170] ), .A2(n5497), .Z(n3309) );
  INV_X2 U6643 ( .I(\SB1_3_13/buf_output[5] ), .ZN(\SB2_3_13/i1_5 ) );
  NAND4_X2 U6654 ( .A1(\SB2_3_31/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_3_31/Component_Function_3/NAND4_in[3] ), .A3(
        \SB2_3_31/Component_Function_3/NAND4_in[0] ), .A4(n3312), .ZN(
        \SB2_3_31/buf_output[3] ) );
  NAND3_X2 U6656 ( .A1(\SB2_3_31/i0_3 ), .A2(\SB2_3_31/i0_4 ), .A3(
        \SB2_3_31/i0_0 ), .ZN(n3312) );
  NAND4_X2 U6658 ( .A1(\SB1_0_22/Component_Function_2/NAND4_in[3] ), .A2(
        \SB1_0_22/Component_Function_2/NAND4_in[2] ), .A3(n3506), .A4(n3314), 
        .ZN(\SB1_0_22/buf_output[2] ) );
  NAND3_X1 U6661 ( .A1(\SB1_0_22/i0[10] ), .A2(\SB1_0_22/i1[9] ), .A3(
        \SB1_0_22/i1_5 ), .ZN(n3314) );
  XOR2_X1 U6662 ( .A1(\MC_ARK_ARC_1_0/temp6[77] ), .A2(n3315), .Z(
        \MC_ARK_ARC_1_0/buf_output[77] ) );
  XOR2_X1 U6663 ( .A1(\MC_ARK_ARC_1_0/temp1[77] ), .A2(
        \MC_ARK_ARC_1_0/temp2[77] ), .Z(n3315) );
  NAND2_X1 U6664 ( .A1(\SB1_3_14/Component_Function_4/NAND4_in[3] ), .A2(n3316), .ZN(n2601) );
  NAND3_X1 U6665 ( .A1(\SB1_3_14/i0_0 ), .A2(\SB1_3_14/i3[0] ), .A3(
        \SB1_3_14/i1_7 ), .ZN(n3316) );
  NAND4_X2 U6679 ( .A1(\SB2_3_13/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_3_13/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_3_13/Component_Function_4/NAND4_in[2] ), .A4(n3320), .ZN(
        \SB2_3_13/buf_output[4] ) );
  NAND4_X2 U6687 ( .A1(\SB2_3_20/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_3_20/Component_Function_2/NAND4_in[2] ), .A3(n3433), .A4(
        \SB2_3_20/Component_Function_2/NAND4_in[0] ), .ZN(
        \SB2_3_20/buf_output[2] ) );
  NAND3_X2 U6701 ( .A1(\SB1_2_19/i0[10] ), .A2(\SB1_2_19/i0_3 ), .A3(
        \SB1_2_19/i0[9] ), .ZN(\SB1_2_19/Component_Function_4/NAND4_in[2] ) );
  XOR2_X1 U6706 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[149] ), .A2(\RI5[2][119] ), 
        .Z(n1491) );
  XOR2_X1 U6713 ( .A1(n4636), .A2(n4635), .Z(\MC_ARK_ARC_1_2/buf_output[134] )
         );
  NAND4_X2 U6719 ( .A1(\SB2_1_23/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_23/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_23/Component_Function_3/NAND4_in[3] ), .A4(
        \SB2_1_23/Component_Function_3/NAND4_in[2] ), .ZN(
        \SB2_1_23/buf_output[3] ) );
  NAND3_X2 U6728 ( .A1(\SB3_21/i0_3 ), .A2(\SB3_21/i0[7] ), .A3(\SB3_21/i0_0 ), 
        .ZN(n2667) );
  NAND3_X2 U6733 ( .A1(\SB2_2_3/i0[10] ), .A2(\SB2_2_3/i1_5 ), .A3(
        \SB2_2_3/i1[9] ), .ZN(n3942) );
  NAND4_X2 U6740 ( .A1(\SB1_0_23/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_23/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_0_23/Component_Function_5/NAND4_in[0] ), .A4(n3322), .ZN(
        \SB1_0_23/buf_output[5] ) );
  NAND3_X1 U6746 ( .A1(\SB1_0_23/i0[9] ), .A2(n358), .A3(n270), .ZN(n3322) );
  NAND4_X2 U6749 ( .A1(n3923), .A2(\SB2_2_24/Component_Function_5/NAND4_in[1] ), .A3(\SB2_2_24/Component_Function_5/NAND4_in[3] ), .A4(n3323), .ZN(
        \SB2_2_24/buf_output[5] ) );
  NAND4_X2 U6759 ( .A1(\SB1_3_17/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_17/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_17/Component_Function_3/NAND4_in[3] ), .A4(n2226), .ZN(
        \SB1_3_17/buf_output[3] ) );
  XOR2_X1 U6767 ( .A1(n3327), .A2(\MC_ARK_ARC_1_2/temp4[137] ), .Z(n3397) );
  XOR2_X1 U6768 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[47] ), .A2(\RI5[2][11] ), 
        .Z(n3327) );
  NAND3_X2 U6785 ( .A1(\SB2_2_0/i0_3 ), .A2(\SB2_2_0/i1[9] ), .A3(
        \SB2_2_0/i0[6] ), .ZN(n1773) );
  NAND3_X2 U6787 ( .A1(\SB2_3_0/i0_3 ), .A2(\SB2_3_0/i1[9] ), .A3(
        \SB1_3_1/buf_output[4] ), .ZN(n3374) );
  AND2_X1 U6793 ( .A1(\SB1_3_22/Component_Function_4/NAND4_in[3] ), .A2(n2118), 
        .Z(n3329) );
  NAND3_X1 U6799 ( .A1(\SB2_2_10/i0[8] ), .A2(\SB2_2_10/i3[0] ), .A3(
        \SB2_2_10/i1_5 ), .ZN(\SB2_2_10/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U6800 ( .A1(n3331), .A2(\MC_ARK_ARC_1_3/temp4[59] ), .Z(
        \MC_ARK_ARC_1_3/temp6[59] ) );
  NAND4_X2 U6805 ( .A1(\SB1_0_22/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_22/Component_Function_4/NAND4_in[3] ), .A3(
        \SB1_0_22/Component_Function_4/NAND4_in[1] ), .A4(n3332), .ZN(
        \SB1_0_22/buf_output[4] ) );
  NAND3_X1 U6806 ( .A1(\SB1_0_22/i0[10] ), .A2(\SB1_0_22/i0_3 ), .A3(
        \SB1_0_22/i0[9] ), .ZN(n3332) );
  NOR2_X2 U6812 ( .A1(n3340), .A2(n3520), .ZN(n3333) );
  XOR2_X1 U6814 ( .A1(\MC_ARK_ARC_1_2/temp5[189] ), .A2(n3335), .Z(
        \MC_ARK_ARC_1_2/buf_output[189] ) );
  XOR2_X1 U6816 ( .A1(\MC_ARK_ARC_1_2/temp3[189] ), .A2(
        \MC_ARK_ARC_1_2/temp4[189] ), .Z(n3335) );
  INV_X2 U6822 ( .I(\SB1_3_0/buf_output[2] ), .ZN(\SB2_3_29/i1[9] ) );
  NAND4_X2 U6823 ( .A1(\SB1_2_20/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_20/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_2_20/Component_Function_5/NAND4_in[0] ), .A4(n3338), .ZN(
        \SB1_2_20/buf_output[5] ) );
  NAND2_X1 U6826 ( .A1(\SB1_1_13/i1[9] ), .A2(\SB1_1_13/i0_3 ), .ZN(
        \SB1_1_13/Component_Function_1/NAND4_in[0] ) );
  NAND4_X2 U6833 ( .A1(\SB2_0_12/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_0_12/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_0_12/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_12/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_0_12/buf_output[1] ) );
  INV_X2 U6844 ( .I(\MC_ARK_ARC_1_1/buf_output[107] ), .ZN(\SB1_2_14/i1_5 ) );
  XOR2_X1 U6845 ( .A1(n1654), .A2(n1653), .Z(\MC_ARK_ARC_1_0/buf_output[110] )
         );
  NAND4_X2 U6855 ( .A1(\SB2_0_14/Component_Function_3/NAND4_in[3] ), .A2(
        \SB2_0_14/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_0_14/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_0_14/Component_Function_3/NAND4_in[1] ), .ZN(
        \SB2_0_14/buf_output[3] ) );
  NAND3_X2 U6859 ( .A1(\SB1_2_28/i0_3 ), .A2(\SB1_2_28/i0_4 ), .A3(
        \SB1_2_28/i1[9] ), .ZN(n4652) );
  NAND2_X2 U6860 ( .A1(n2457), .A2(n4477), .ZN(n3340) );
  XOR2_X1 U6861 ( .A1(n3342), .A2(n3341), .Z(\MC_ARK_ARC_1_0/temp6[15] ) );
  XOR2_X1 U6869 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[81] ), .A2(n205), .Z(n3341) );
  XOR2_X1 U6870 ( .A1(\RI5[0][117] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[51] ), 
        .Z(n3342) );
  INV_X2 U6875 ( .I(\RI3[1][110] ), .ZN(\SB2_1_13/i1[9] ) );
  XOR2_X1 U6879 ( .A1(\RI5[2][160] ), .A2(\RI5[2][166] ), .Z(n3345) );
  NAND3_X2 U6886 ( .A1(\SB1_1_20/i0_3 ), .A2(\SB1_1_20/i0_0 ), .A3(
        \SB1_1_20/i0_4 ), .ZN(\SB1_1_20/Component_Function_3/NAND4_in[1] ) );
  NAND2_X2 U6889 ( .A1(\SB1_2_10/Component_Function_4/NAND4_in[3] ), .A2(n3347), .ZN(n3520) );
  NAND3_X2 U6891 ( .A1(\SB1_2_10/i0[9] ), .A2(\SB1_2_10/i0_3 ), .A3(
        \SB1_2_10/i0[10] ), .ZN(n3347) );
  XOR2_X1 U6896 ( .A1(n3350), .A2(n3349), .Z(\MC_ARK_ARC_1_2/buf_output[149] )
         );
  XOR2_X1 U6897 ( .A1(n1491), .A2(\MC_ARK_ARC_1_2/temp4[149] ), .Z(n3349) );
  XOR2_X1 U6937 ( .A1(\RI5[3][170] ), .A2(\RI5[3][134] ), .Z(n3356) );
  NAND4_X2 U6938 ( .A1(\SB2_1_18/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_1_18/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_1_18/Component_Function_0/NAND4_in[0] ), .A4(n3357), .ZN(
        \SB2_1_18/buf_output[0] ) );
  XOR2_X1 U6943 ( .A1(\MC_ARK_ARC_1_3/temp1[102] ), .A2(
        \MC_ARK_ARC_1_3/temp2[102] ), .Z(n4442) );
  NAND2_X2 U6945 ( .A1(\SB1_3_7/i0_0 ), .A2(\SB1_3_7/i3[0] ), .ZN(
        \SB1_3_7/Component_Function_5/NAND4_in[0] ) );
  NAND4_X2 U6969 ( .A1(\SB1_3_31/Component_Function_1/NAND4_in[1] ), .A2(n3731), .A3(\SB1_3_31/Component_Function_1/NAND4_in[0] ), .A4(
        \SB1_3_31/Component_Function_1/NAND4_in[3] ), .ZN(n3680) );
  XOR2_X1 U6980 ( .A1(n3368), .A2(n3367), .Z(\MC_ARK_ARC_1_1/temp5[86] ) );
  XOR2_X1 U6981 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[80] ), .A2(\RI5[1][56] ), 
        .Z(n3367) );
  XOR2_X1 U6984 ( .A1(\RI5[1][86] ), .A2(\RI5[1][32] ), .Z(n3368) );
  INV_X2 U6994 ( .I(\SB1_1_27/buf_output[3] ), .ZN(\SB2_1_25/i0[8] ) );
  NAND4_X2 U6996 ( .A1(n4376), .A2(\SB1_1_27/Component_Function_3/NAND4_in[1] ), .A3(\SB1_1_27/Component_Function_3/NAND4_in[0] ), .A4(
        \SB1_1_27/Component_Function_3/NAND4_in[2] ), .ZN(
        \SB1_1_27/buf_output[3] ) );
  INV_X2 U6998 ( .I(\SB1_1_9/buf_output[3] ), .ZN(\SB2_1_7/i0[8] ) );
  NAND4_X2 U7012 ( .A1(\SB2_0_8/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_0_8/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_0_8/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_0_8/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB2_0_8/buf_output[4] ) );
  XOR2_X1 U7024 ( .A1(n3373), .A2(\MC_ARK_ARC_1_2/temp6[141] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[141] ) );
  XOR2_X1 U7030 ( .A1(n3735), .A2(n1115), .Z(n3373) );
  NAND4_X2 U7034 ( .A1(\SB2_1_23/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_1_23/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_1_23/Component_Function_1/NAND4_in[1] ), .A4(
        \SB2_1_23/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_1_23/buf_output[1] ) );
  XOR2_X1 U7036 ( .A1(\RI5[0][57] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[81] ), 
        .Z(n3884) );
  XOR2_X1 U7039 ( .A1(n3375), .A2(n2212), .Z(\MC_ARK_ARC_1_2/buf_output[11] )
         );
  XOR2_X1 U7040 ( .A1(\MC_ARK_ARC_1_2/temp2[11] ), .A2(
        \MC_ARK_ARC_1_2/temp1[11] ), .Z(n3375) );
  INV_X2 U7041 ( .I(\MC_ARK_ARC_1_2/buf_output[171] ), .ZN(\SB1_3_3/i0[8] ) );
  NAND4_X2 U7060 ( .A1(\SB1_1_21/Component_Function_0/NAND4_in[3] ), .A2(n4611), .A3(\SB1_1_21/Component_Function_0/NAND4_in[1] ), .A4(n3378), .ZN(
        \SB1_1_21/buf_output[0] ) );
  XOR2_X1 U7063 ( .A1(\RI5[3][137] ), .A2(\RI5[3][143] ), .Z(
        \MC_ARK_ARC_1_3/temp1[143] ) );
  XOR2_X1 U7085 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[74] ), .A2(n507), .Z(n3381) );
  XOR2_X1 U7091 ( .A1(\RI5[2][8] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[38] ), 
        .Z(n3382) );
  NAND3_X2 U7093 ( .A1(\SB2_3_3/i0_4 ), .A2(\SB2_3_3/i1_5 ), .A3(
        \SB2_3_3/i0_0 ), .ZN(\SB2_3_3/Component_Function_2/NAND4_in[3] ) );
  NAND4_X2 U7094 ( .A1(n2060), .A2(\SB2_1_20/Component_Function_1/NAND4_in[1] ), .A3(\SB2_1_20/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_20/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_1_20/buf_output[1] ) );
  NAND3_X2 U7100 ( .A1(\SB2_2_1/i0_3 ), .A2(\SB2_2_1/i0[10] ), .A3(
        \SB2_2_1/i0[6] ), .ZN(\SB2_2_1/Component_Function_2/NAND4_in[1] ) );
  INV_X2 U7101 ( .I(\MC_ARK_ARC_1_2/buf_output[164] ), .ZN(\SB1_3_4/i1[9] ) );
  INV_X1 U7107 ( .I(\SB3_29/buf_output[3] ), .ZN(\SB4_27/i0[8] ) );
  NAND4_X2 U7112 ( .A1(\SB3_29/Component_Function_3/NAND4_in[1] ), .A2(n2023), 
        .A3(\SB3_29/Component_Function_3/NAND4_in[3] ), .A4(
        \SB3_29/Component_Function_3/NAND4_in[0] ), .ZN(\SB3_29/buf_output[3] ) );
  NAND4_X2 U7116 ( .A1(\SB1_1_24/Component_Function_1/NAND4_in[3] ), .A2(n4537), .A3(\SB1_1_24/Component_Function_1/NAND4_in[2] ), .A4(n3385), .ZN(
        \SB1_1_24/buf_output[1] ) );
  NAND2_X1 U7125 ( .A1(\SB4_12/i0[9] ), .A2(\SB4_12/i0[10] ), .ZN(n3388) );
  XOR2_X1 U7126 ( .A1(\MC_ARK_ARC_1_3/temp1[27] ), .A2(n3389), .Z(
        \MC_ARK_ARC_1_3/temp5[27] ) );
  XOR2_X1 U7128 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[165] ), .A2(\RI5[3][189] ), 
        .Z(n3389) );
  XOR2_X1 U7135 ( .A1(n4581), .A2(n3390), .Z(\MC_ARK_ARC_1_2/temp5[21] ) );
  XOR2_X1 U7138 ( .A1(\RI5[2][15] ), .A2(\RI5[2][21] ), .Z(n3390) );
  INV_X2 U7140 ( .I(\SB1_0_8/buf_output[5] ), .ZN(\SB2_0_8/i1_5 ) );
  NAND4_X2 U7149 ( .A1(\SB1_0_8/Component_Function_5/NAND4_in[1] ), .A2(n2539), 
        .A3(\SB1_0_8/Component_Function_5/NAND4_in[0] ), .A4(n2715), .ZN(
        \SB1_0_8/buf_output[5] ) );
  NAND3_X1 U7153 ( .A1(\SB4_0/i1_7 ), .A2(\SB3_3/buf_output[2] ), .A3(
        \SB4_0/i3[0] ), .ZN(n2658) );
  XOR2_X1 U7156 ( .A1(\MC_ARK_ARC_1_1/temp1[74] ), .A2(n3393), .Z(n2062) );
  NAND4_X2 U7170 ( .A1(\SB2_0_8/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_8/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_0_8/Component_Function_3/NAND4_in[3] ), .A4(n3394), .ZN(
        \SB2_0_8/buf_output[3] ) );
  NAND3_X2 U7175 ( .A1(\SB2_0_8/i0_3 ), .A2(\SB2_0_8/i0_0 ), .A3(\RI3[0][142] ), .ZN(n3394) );
  XOR2_X1 U7180 ( .A1(n3395), .A2(n3503), .Z(n2815) );
  XOR2_X1 U7185 ( .A1(\RI5[0][153] ), .A2(\RI5[0][87] ), .Z(n3395) );
  NAND4_X2 U7188 ( .A1(\SB2_1_13/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_1_13/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_1_13/Component_Function_3/NAND4_in[1] ), .A4(n3396), .ZN(
        \SB2_1_13/buf_output[3] ) );
  XOR2_X1 U7190 ( .A1(n3711), .A2(n3397), .Z(\MC_ARK_ARC_1_2/buf_output[137] )
         );
  NAND3_X1 U7199 ( .A1(\SB4_7/i0_3 ), .A2(\SB4_7/i0[6] ), .A3(\SB4_7/i1[9] ), 
        .ZN(n3399) );
  XOR2_X1 U7209 ( .A1(n3400), .A2(n39), .Z(Ciphertext[84]) );
  NAND4_X2 U7210 ( .A1(\SB4_17/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_17/Component_Function_0/NAND4_in[1] ), .A3(n3836), .A4(
        \SB4_17/Component_Function_0/NAND4_in[0] ), .ZN(n3400) );
  NAND3_X1 U7221 ( .A1(\SB1_2_26/i0[8] ), .A2(\SB1_2_26/i0_0 ), .A3(
        \SB1_2_26/i0[9] ), .ZN(\SB1_2_26/Component_Function_4/NAND4_in[0] ) );
  XOR2_X1 U7228 ( .A1(\MC_ARK_ARC_1_2/temp2[170] ), .A2(n3401), .Z(n3825) );
  XOR2_X1 U7230 ( .A1(\RI5[2][170] ), .A2(\RI5[2][164] ), .Z(n3401) );
  XOR2_X1 U7238 ( .A1(n3402), .A2(\MC_ARK_ARC_1_0/temp5[187] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[187] ) );
  XOR2_X1 U7243 ( .A1(\MC_ARK_ARC_1_0/temp3[187] ), .A2(
        \MC_ARK_ARC_1_0/temp4[187] ), .Z(n3402) );
  NAND4_X2 U7269 ( .A1(\SB1_2_1/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_2_1/Component_Function_1/NAND4_in[0] ), .A3(
        \SB1_2_1/Component_Function_1/NAND4_in[3] ), .A4(n3404), .ZN(
        \SB1_2_1/buf_output[1] ) );
  NAND4_X2 U7274 ( .A1(\SB1_1_28/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_28/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_1_28/Component_Function_5/NAND4_in[0] ), .A4(n3405), .ZN(
        \SB1_1_28/buf_output[5] ) );
  XOR2_X1 U7279 ( .A1(n3407), .A2(\MC_ARK_ARC_1_1/temp5[164] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[164] ) );
  XOR2_X1 U7280 ( .A1(\MC_ARK_ARC_1_1/temp4[164] ), .A2(
        \MC_ARK_ARC_1_1/temp3[164] ), .Z(n3407) );
  NAND3_X1 U7290 ( .A1(\SB2_2_22/i0[9] ), .A2(\SB2_2_22/i0[6] ), .A3(
        \SB2_2_22/i1_5 ), .ZN(n3409) );
  NAND3_X2 U7294 ( .A1(\SB2_0_27/i0_3 ), .A2(n2679), .A3(\SB2_0_27/i0[8] ), 
        .ZN(\SB2_0_27/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 U7295 ( .I(\SB1_0_25/buf_output[5] ), .Z(\SB2_0_25/i0_3 ) );
  NAND3_X2 U7297 ( .A1(\SB2_0_31/i0[10] ), .A2(\SB2_0_31/i0_3 ), .A3(
        \SB2_0_31/i0[6] ), .ZN(\SB2_0_31/Component_Function_2/NAND4_in[1] ) );
  XOR2_X1 U7303 ( .A1(n3410), .A2(\MC_ARK_ARC_1_1/temp2[150] ), .Z(
        \MC_ARK_ARC_1_1/temp5[150] ) );
  XOR2_X1 U7310 ( .A1(\RI5[1][144] ), .A2(\RI5[1][150] ), .Z(n3410) );
  NAND4_X2 U7311 ( .A1(\SB2_0_27/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_0_27/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_0_27/Component_Function_3/NAND4_in[1] ), .A4(
        \SB2_0_27/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_0_27/buf_output[3] ) );
  NAND4_X2 U7316 ( .A1(\SB1_2_25/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_2_25/Component_Function_4/NAND4_in[3] ), .A3(
        \SB1_2_25/Component_Function_4/NAND4_in[0] ), .A4(n3411), .ZN(
        \SB1_2_25/buf_output[4] ) );
  NAND3_X2 U7317 ( .A1(\SB1_2_25/i0[10] ), .A2(\SB1_2_25/i0_3 ), .A3(
        \SB1_2_25/i0[9] ), .ZN(n3411) );
  NOR2_X2 U7318 ( .A1(n3413), .A2(n3412), .ZN(n3671) );
  NAND3_X1 U7338 ( .A1(\SB1_3_14/i0[6] ), .A2(\SB1_3_14/i0_3 ), .A3(
        \SB1_3_14/i0[10] ), .ZN(\SB1_3_14/Component_Function_2/NAND4_in[1] )
         );
  XOR2_X1 U7341 ( .A1(\MC_ARK_ARC_1_0/temp3[80] ), .A2(
        \MC_ARK_ARC_1_0/temp4[80] ), .Z(n3416) );
  XOR2_X1 U7347 ( .A1(\MC_ARK_ARC_1_1/temp5[83] ), .A2(n1527), .Z(
        \MC_ARK_ARC_1_1/buf_output[83] ) );
  NAND4_X2 U7353 ( .A1(\SB1_0_1/Component_Function_3/NAND4_in[2] ), .A2(
        \SB1_0_1/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_1/Component_Function_3/NAND4_in[0] ), .A4(n3419), .ZN(
        \RI3[0][3] ) );
  XOR2_X1 U7360 ( .A1(n2154), .A2(\MC_ARK_ARC_1_1/temp2[69] ), .Z(
        \MC_ARK_ARC_1_1/temp5[69] ) );
  XOR2_X1 U7367 ( .A1(n2292), .A2(n3422), .Z(n3937) );
  XOR2_X1 U7376 ( .A1(n3426), .A2(n3425), .Z(\MC_ARK_ARC_1_3/temp5[44] ) );
  XOR2_X1 U7380 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[182] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[38] ), .Z(n3425) );
  XOR2_X1 U7381 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[44] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[14] ), .Z(n3426) );
  XOR2_X1 U7391 ( .A1(n3427), .A2(n3428), .Z(n625) );
  XOR2_X1 U7394 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[25] ), .A2(\RI5[1][79] ), 
        .Z(n3427) );
  XOR2_X1 U7397 ( .A1(\RI5[1][73] ), .A2(\RI5[1][49] ), .Z(n3428) );
  NAND4_X2 U7402 ( .A1(\SB2_3_28/Component_Function_5/NAND4_in[1] ), .A2(
        \SB2_3_28/Component_Function_5/NAND4_in[2] ), .A3(
        \SB2_3_28/Component_Function_5/NAND4_in[0] ), .A4(n3430), .ZN(
        \SB2_3_28/buf_output[5] ) );
  INV_X2 U7403 ( .I(\SB1_3_17/buf_output[2] ), .ZN(\SB2_3_14/i1[9] ) );
  XOR2_X1 U7408 ( .A1(n3431), .A2(\MC_ARK_ARC_1_3/temp5[76] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[76] ) );
  XOR2_X1 U7411 ( .A1(\MC_ARK_ARC_1_3/temp4[76] ), .A2(
        \MC_ARK_ARC_1_3/temp3[76] ), .Z(n3431) );
  NAND3_X1 U7424 ( .A1(\SB1_3_29/i1_7 ), .A2(\RI1[3][14] ), .A3(
        \SB1_3_29/i3[0] ), .ZN(\SB1_3_29/Component_Function_4/NAND4_in[1] ) );
  INV_X2 U7426 ( .I(\SB1_0_7/buf_output[3] ), .ZN(\SB2_0_5/i0[8] ) );
  INV_X2 U7428 ( .I(\SB1_3_26/buf_output[2] ), .ZN(\SB2_3_23/i1[9] ) );
  NAND4_X2 U7436 ( .A1(n1835), .A2(\SB2_3_24/Component_Function_3/NAND4_in[0] ), .A3(\SB2_3_24/Component_Function_3/NAND4_in[1] ), .A4(n3435), .ZN(
        \SB2_3_24/buf_output[3] ) );
  INV_X2 U7447 ( .I(\MC_ARK_ARC_1_1/buf_output[79] ), .ZN(\SB1_2_18/i1_7 ) );
  NAND4_X2 U7458 ( .A1(\SB2_2_1/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_1/Component_Function_3/NAND4_in[3] ), .A3(
        \SB2_2_1/Component_Function_3/NAND4_in[2] ), .A4(n3437), .ZN(
        \SB2_2_1/buf_output[3] ) );
  NAND4_X2 U7468 ( .A1(\SB1_3_23/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_3_23/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_3_23/Component_Function_3/NAND4_in[2] ), .A4(n1712), .ZN(
        \SB1_3_23/buf_output[3] ) );
  XOR2_X1 U7470 ( .A1(\RI5[2][119] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[83] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[17] ) );
  NAND4_X2 U7474 ( .A1(\SB2_0_18/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_18/Component_Function_5/NAND4_in[1] ), .A3(n3633), .A4(
        \SB2_0_18/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_0_18/buf_output[5] ) );
  NAND3_X1 U7476 ( .A1(\SB3_19/i0[10] ), .A2(\SB3_19/i0_0 ), .A3(
        \SB3_19/i0[6] ), .ZN(\SB3_19/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U7485 ( .A1(\RI5[0][59] ), .A2(\RI5[0][83] ), .Z(
        \MC_ARK_ARC_1_0/temp2[113] ) );
  NAND4_X2 U7505 ( .A1(\SB2_0_29/Component_Function_5/NAND4_in[0] ), .A2(n4610), .A3(\SB2_0_29/Component_Function_5/NAND4_in[1] ), .A4(n3439), .ZN(
        \SB2_0_29/buf_output[5] ) );
  NAND3_X2 U7511 ( .A1(\SB1_0_20/i0[10] ), .A2(\SB1_0_20/i0[6] ), .A3(
        \SB1_0_20/i0_3 ), .ZN(n3442) );
  XOR2_X1 U7519 ( .A1(\RI5[1][125] ), .A2(\RI5[1][131] ), .Z(n3443) );
  NAND3_X2 U7520 ( .A1(\SB2_0_14/i1[9] ), .A2(\SB2_0_14/i1_7 ), .A3(
        \RI3[0][105] ), .ZN(\SB2_0_14/Component_Function_3/NAND4_in[2] ) );
  NAND4_X2 U7535 ( .A1(\SB3_7/Component_Function_5/NAND4_in[2] ), .A2(n1982), 
        .A3(n1680), .A4(n3445), .ZN(\SB3_7/buf_output[5] ) );
  XOR2_X1 U7548 ( .A1(\MC_ARK_ARC_1_3/temp6[147] ), .A2(
        \MC_ARK_ARC_1_3/temp5[147] ), .Z(\MC_ARK_ARC_1_3/buf_output[147] ) );
  XOR2_X1 U7549 ( .A1(\MC_ARK_ARC_1_3/temp3[147] ), .A2(
        \MC_ARK_ARC_1_3/temp4[147] ), .Z(\MC_ARK_ARC_1_3/temp6[147] ) );
  NAND4_X2 U7550 ( .A1(\SB2_2_5/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_2_5/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_2_5/Component_Function_4/NAND4_in[3] ), .A4(n3447), .ZN(
        \SB2_2_5/buf_output[4] ) );
  NAND3_X2 U7560 ( .A1(\SB2_2_5/i0[10] ), .A2(\SB2_2_5/i0_3 ), .A3(
        \SB2_2_5/i0[9] ), .ZN(n3447) );
  BUF_X4 U7561 ( .I(\MC_ARK_ARC_1_0/buf_output[75] ), .Z(\SB1_1_19/i0[10] ) );
  NAND4_X2 U7562 ( .A1(\SB1_2_5/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_5/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_2_5/Component_Function_5/NAND4_in[0] ), .A4(n3448), .ZN(
        \SB1_2_5/buf_output[5] ) );
  NAND3_X2 U7563 ( .A1(\SB1_2_5/i0[9] ), .A2(\SB1_2_5/i0[6] ), .A3(
        \SB1_2_5/i0_4 ), .ZN(n3448) );
  BUF_X4 U7575 ( .I(\SB2_3_17/buf_output[3] ), .Z(\RI5[3][99] ) );
  NAND4_X2 U7576 ( .A1(\SB1_3_23/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_23/Component_Function_4/NAND4_in[3] ), .A3(n3479), .A4(n3452), 
        .ZN(\SB1_3_23/buf_output[4] ) );
  XOR2_X1 U7589 ( .A1(\MC_ARK_ARC_1_0/temp3[68] ), .A2(
        \MC_ARK_ARC_1_0/temp4[68] ), .Z(n3454) );
  NAND3_X1 U7594 ( .A1(\SB4_27/i0[9] ), .A2(n2898), .A3(\SB4_27/i0[8] ), .ZN(
        n3456) );
  NAND3_X1 U7605 ( .A1(\SB1_0_17/i0[6] ), .A2(\SB1_0_17/i0_3 ), .A3(
        \SB1_0_17/i1[9] ), .ZN(\SB1_0_17/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U7613 ( .A1(\RI5[3][145] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[109] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[43] ) );
  XOR2_X1 U7622 ( .A1(\RI5[3][26] ), .A2(\RI5[3][62] ), .Z(
        \MC_ARK_ARC_1_3/temp3[152] ) );
  BUF_X2 U7625 ( .I(\SB2_1_30/buf_output[5] ), .Z(n3650) );
  NAND4_X2 U7626 ( .A1(\SB1_0_26/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_0_26/Component_Function_2/NAND4_in[3] ), .A3(
        \SB1_0_26/Component_Function_2/NAND4_in[1] ), .A4(n3463), .ZN(
        \RI3[0][50] ) );
  INV_X1 U7630 ( .I(\SB3_12/buf_output[2] ), .ZN(\SB4_9/i1[9] ) );
  NAND4_X2 U7634 ( .A1(\SB2_3_4/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_4/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_3_4/Component_Function_4/NAND4_in[3] ), .A4(n3464), .ZN(
        \SB2_3_4/buf_output[4] ) );
  XOR2_X1 U7650 ( .A1(n2661), .A2(n2660), .Z(\MC_ARK_ARC_1_3/temp6[65] ) );
  NAND3_X1 U7652 ( .A1(n1793), .A2(\SB4_29/i0_3 ), .A3(\SB4_29/i1[9] ), .ZN(
        \SB4_29/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U7655 ( .A1(\SB1_1_4/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_4/Component_Function_3/NAND4_in[1] ), .A3(n4734), .A4(
        \SB1_1_4/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_1_4/buf_output[3] ) );
  NAND3_X1 U7659 ( .A1(\SB4_29/i0_0 ), .A2(\SB4_29/i0_3 ), .A3(\SB4_29/i0[7] ), 
        .ZN(n4225) );
  NAND4_X2 U7660 ( .A1(n3561), .A2(n2178), .A3(
        \SB2_0_24/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_0_24/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_0_24/buf_output[5] ) );
  NAND3_X2 U7667 ( .A1(\SB2_1_22/i0_4 ), .A2(\SB2_1_22/i0[6] ), .A3(
        \SB2_1_22/i0[9] ), .ZN(\SB2_1_22/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 U7668 ( .A1(\SB2_1_20/i1[9] ), .A2(\SB2_1_20/i0_3 ), .A3(
        \SB2_1_20/i0[6] ), .ZN(\SB2_1_20/Component_Function_3/NAND4_in[0] ) );
  NAND4_X2 U7673 ( .A1(\SB1_2_26/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_26/Component_Function_2/NAND4_in[1] ), .A3(n4704), .A4(
        \SB1_2_26/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB1_2_26/buf_output[2] ) );
  NAND4_X2 U7678 ( .A1(\SB1_2_29/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_2_29/Component_Function_0/NAND4_in[0] ), .A3(
        \SB1_2_29/Component_Function_0/NAND4_in[2] ), .A4(n3466), .ZN(
        \SB1_2_29/buf_output[0] ) );
  NAND3_X1 U7682 ( .A1(\SB1_2_29/i0_0 ), .A2(\RI1[2][17] ), .A3(
        \SB1_2_29/i0[7] ), .ZN(n3466) );
  NAND3_X2 U7687 ( .A1(\SB2_2_23/i0_3 ), .A2(\SB2_2_23/i0[8] ), .A3(
        \SB2_2_23/i1_7 ), .ZN(\SB2_2_23/Component_Function_1/NAND4_in[1] ) );
  NAND3_X2 U7692 ( .A1(\SB4_18/i0[6] ), .A2(\SB4_18/i0[10] ), .A3(
        \SB4_18/i0_3 ), .ZN(n3468) );
  NAND3_X1 U7707 ( .A1(\SB4_4/i0_4 ), .A2(n3655), .A3(\SB4_4/i1_5 ), .ZN(n3471) );
  XOR2_X1 U7709 ( .A1(n3472), .A2(\MC_ARK_ARC_1_0/temp1[31] ), .Z(
        \MC_ARK_ARC_1_0/temp5[31] ) );
  XOR2_X1 U7713 ( .A1(\RI5[0][169] ), .A2(\RI5[0][1] ), .Z(n3472) );
  XOR2_X1 U7714 ( .A1(\MC_ARK_ARC_1_3/temp1[164] ), .A2(n3473), .Z(
        \MC_ARK_ARC_1_3/temp5[164] ) );
  XOR2_X1 U7715 ( .A1(\RI5[3][134] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[110] ), 
        .Z(n3473) );
  XOR2_X1 U7729 ( .A1(\MC_ARK_ARC_1_0/temp5[27] ), .A2(n3476), .Z(
        \MC_ARK_ARC_1_0/buf_output[27] ) );
  XOR2_X1 U7730 ( .A1(\MC_ARK_ARC_1_0/temp3[27] ), .A2(
        \MC_ARK_ARC_1_0/temp4[27] ), .Z(n3476) );
  INV_X2 U7732 ( .I(\RI3[0][50] ), .ZN(\SB2_0_23/i1[9] ) );
  XOR2_X1 U7735 ( .A1(n3477), .A2(n3478), .Z(\MC_ARK_ARC_1_1/temp5[110] ) );
  XOR2_X1 U7739 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[80] ), .A2(\RI5[1][56] ), 
        .Z(n3477) );
  XOR2_X1 U7740 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[110] ), .A2(\RI5[1][104] ), 
        .Z(n3478) );
  NAND3_X2 U7744 ( .A1(\SB2_0_21/i0[10] ), .A2(\SB2_0_21/i1_7 ), .A3(
        \SB2_0_21/i1[9] ), .ZN(n3797) );
  NAND3_X2 U7752 ( .A1(\SB1_3_23/i0[10] ), .A2(\SB1_3_23/i0_3 ), .A3(
        \SB1_3_23/i0[9] ), .ZN(n3479) );
  NAND3_X2 U7764 ( .A1(\SB2_0_14/i1[9] ), .A2(\SB2_0_14/i1_5 ), .A3(
        \RI3[0][105] ), .ZN(\SB2_0_14/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U7767 ( .A1(\SB2_0_17/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_0_17/Component_Function_0/NAND4_in[2] ), .A3(n1697), .A4(
        \SB2_0_17/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_0_17/buf_output[0] ) );
  NAND4_X2 U7776 ( .A1(n4163), .A2(\SB1_0_17/Component_Function_5/NAND4_in[2] ), .A3(\SB1_0_17/Component_Function_5/NAND4_in[0] ), .A4(n3482), .ZN(
        \SB1_0_17/buf_output[5] ) );
  NAND3_X2 U7778 ( .A1(\SB1_0_17/i0[6] ), .A2(n2899), .A3(\SB1_0_17/i0[9] ), 
        .ZN(n3482) );
  NAND3_X2 U7786 ( .A1(\SB2_2_3/i0_3 ), .A2(\SB2_2_3/i1[9] ), .A3(
        \SB2_2_3/i0[6] ), .ZN(\SB2_2_3/Component_Function_3/NAND4_in[0] ) );
  NAND4_X2 U7793 ( .A1(\SB1_2_27/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_27/Component_Function_3/NAND4_in[1] ), .A3(n3522), .A4(
        \SB1_2_27/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_2_27/buf_output[3] ) );
  XOR2_X1 U7798 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[177] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[183] ), .Z(\MC_ARK_ARC_1_2/temp1[183] )
         );
  XOR2_X1 U7813 ( .A1(n3484), .A2(n3483), .Z(\MC_ARK_ARC_1_2/temp5[132] ) );
  XOR2_X1 U7818 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[132] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[78] ), .Z(n3484) );
  NAND3_X2 U7830 ( .A1(\SB2_2_30/i0_3 ), .A2(\SB2_2_30/i1[9] ), .A3(n2343), 
        .ZN(n3485) );
  BUF_X4 U7861 ( .I(\SB1_0_15/buf_output[5] ), .Z(\SB2_0_15/i0_3 ) );
  NAND4_X2 U7865 ( .A1(\SB2_2_11/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_2_11/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_11/Component_Function_0/NAND4_in[0] ), .A4(n3490), .ZN(
        \SB2_2_11/buf_output[0] ) );
  XOR2_X1 U7870 ( .A1(n3492), .A2(\MC_ARK_ARC_1_1/temp5[123] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[123] ) );
  XOR2_X1 U7872 ( .A1(\MC_ARK_ARC_1_1/temp4[123] ), .A2(
        \MC_ARK_ARC_1_1/temp3[123] ), .Z(n3492) );
  XOR2_X1 U7876 ( .A1(\RI5[1][14] ), .A2(\RI5[1][8] ), .Z(
        \MC_ARK_ARC_1_1/temp1[14] ) );
  INV_X2 U7877 ( .I(\SB1_3_6/buf_output[3] ), .ZN(\SB2_3_4/i0[8] ) );
  XOR2_X1 U7900 ( .A1(\MC_ARK_ARC_1_2/temp5[92] ), .A2(n3496), .Z(
        \MC_ARK_ARC_1_2/buf_output[92] ) );
  BUF_X4 U7903 ( .I(\SB2_3_29/buf_output[2] ), .Z(\RI5[3][32] ) );
  XOR2_X1 U7904 ( .A1(\MC_ARK_ARC_1_2/temp5[3] ), .A2(n3497), .Z(
        \MC_ARK_ARC_1_2/buf_output[3] ) );
  XOR2_X1 U7909 ( .A1(\MC_ARK_ARC_1_2/temp3[3] ), .A2(
        \MC_ARK_ARC_1_2/temp4[3] ), .Z(n3497) );
  XOR2_X1 U7914 ( .A1(\MC_ARK_ARC_1_1/temp4[35] ), .A2(n3499), .Z(n2433) );
  XOR2_X1 U7915 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[101] ), .A2(\RI5[1][137] ), 
        .Z(n3499) );
  XOR2_X1 U7922 ( .A1(\MC_ARK_ARC_1_0/temp5[24] ), .A2(n3500), .Z(
        \MC_ARK_ARC_1_0/buf_output[24] ) );
  XOR2_X1 U7933 ( .A1(\MC_ARK_ARC_1_0/temp3[24] ), .A2(
        \MC_ARK_ARC_1_0/temp4[24] ), .Z(n3500) );
  NAND4_X2 U7943 ( .A1(\SB2_0_15/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_15/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_0_15/Component_Function_4/NAND4_in[1] ), .A4(n3501), .ZN(
        \SB2_0_15/buf_output[4] ) );
  INV_X2 U7944 ( .I(\SB1_0_15/buf_output[5] ), .ZN(\SB2_0_15/i1_5 ) );
  XOR2_X1 U7947 ( .A1(\SB2_0_14/buf_output[3] ), .A2(n450), .Z(n3503) );
  NAND3_X2 U7948 ( .A1(\SB1_0_16/i0_0 ), .A2(\SB1_0_16/i0[10] ), .A3(
        \SB1_0_16/i0[6] ), .ZN(n3505) );
  NAND3_X1 U7950 ( .A1(\SB1_0_22/i0[10] ), .A2(\SB1_0_22/i0_3 ), .A3(
        \SB1_0_22/i0[6] ), .ZN(n3506) );
  NAND4_X2 U7951 ( .A1(\SB2_0_17/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_0_17/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_17/Component_Function_1/NAND4_in[0] ), .A4(n3507), .ZN(
        \SB2_0_17/buf_output[1] ) );
  NAND4_X2 U7952 ( .A1(\SB1_1_19/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_19/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_19/Component_Function_1/NAND4_in[3] ), .A4(n3508), .ZN(
        \SB1_1_19/buf_output[1] ) );
  XOR2_X1 U7957 ( .A1(\RI5[1][147] ), .A2(n209), .Z(
        \MC_ARK_ARC_1_1/temp4[111] ) );
  NAND4_X2 U7981 ( .A1(\SB1_1_2/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_1_2/Component_Function_0/NAND4_in[0] ), .A3(
        \SB1_1_2/Component_Function_0/NAND4_in[3] ), .A4(
        \SB1_1_2/Component_Function_0/NAND4_in[1] ), .ZN(
        \SB1_1_2/buf_output[0] ) );
  NAND4_X2 U8011 ( .A1(\SB2_3_24/Component_Function_2/NAND4_in[3] ), .A2(
        \SB2_3_24/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_24/Component_Function_2/NAND4_in[0] ), .A4(n3833), .ZN(
        \SB2_3_24/buf_output[2] ) );
  XOR2_X1 U8015 ( .A1(\MC_ARK_ARC_1_0/temp6[74] ), .A2(n3513), .Z(
        \MC_ARK_ARC_1_0/buf_output[74] ) );
  NAND3_X2 U8021 ( .A1(\SB2_1_9/i0_0 ), .A2(\SB2_1_9/i0_4 ), .A3(
        \SB2_1_9/i1_5 ), .ZN(n3514) );
  XOR2_X1 U8027 ( .A1(\MC_ARK_ARC_1_1/temp1[28] ), .A2(n3516), .Z(
        \MC_ARK_ARC_1_1/temp5[28] ) );
  XOR2_X1 U8028 ( .A1(\RI5[1][166] ), .A2(\RI5[1][190] ), .Z(n3516) );
  NAND3_X2 U8037 ( .A1(\SB2_0_25/i0[8] ), .A2(\SB2_0_25/i3[0] ), .A3(
        \SB2_0_25/i1_5 ), .ZN(n3517) );
  NAND3_X2 U8041 ( .A1(\SB1_0_23/i0[9] ), .A2(\SB1_0_23/i0_3 ), .A3(
        \SB1_0_23/i0[8] ), .ZN(n3574) );
  INV_X1 U8043 ( .I(\SB1_1_19/buf_output[0] ), .ZN(\SB2_1_14/i3[0] ) );
  NAND4_X2 U8047 ( .A1(\SB1_1_19/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_1_19/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_1_19/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_1_19/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_1_19/buf_output[0] ) );
  BUF_X4 U8053 ( .I(\RI1[3][71] ), .Z(\SB1_3_20/i0_3 ) );
  XOR2_X1 U8071 ( .A1(\MC_ARK_ARC_1_2/temp1[71] ), .A2(n3524), .Z(
        \MC_ARK_ARC_1_2/temp5[71] ) );
  XOR2_X1 U8087 ( .A1(\RI5[2][41] ), .A2(\RI5[2][17] ), .Z(n3524) );
  INV_X2 U8096 ( .I(\RI1[3][71] ), .ZN(\SB1_3_20/i1_5 ) );
  NAND3_X1 U8098 ( .A1(\SB1_2_29/i0[8] ), .A2(\RI1[2][17] ), .A3(
        \SB1_2_29/i1_7 ), .ZN(\SB1_2_29/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 U8120 ( .A1(n2442), .A2(n3760), .ZN(n607) );
  NAND4_X2 U8125 ( .A1(\SB1_0_1/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_0_1/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_0_1/Component_Function_0/NAND4_in[0] ), .A4(n3525), .ZN(
        \SB1_0_1/buf_output[0] ) );
  NAND4_X2 U8126 ( .A1(\SB2_0_23/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_0_23/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_0_23/Component_Function_4/NAND4_in[1] ), .A4(n3526), .ZN(
        \SB2_0_23/buf_output[4] ) );
  NAND3_X2 U8132 ( .A1(\SB1_0_5/i0_3 ), .A2(\SB1_0_5/i0_4 ), .A3(
        \SB1_0_5/i1[9] ), .ZN(\SB1_0_5/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U8135 ( .A1(n3529), .A2(n3528), .Z(n4110) );
  XOR2_X1 U8136 ( .A1(\RI5[0][113] ), .A2(\RI5[0][89] ), .Z(n3528) );
  XOR2_X1 U8137 ( .A1(\RI5[0][137] ), .A2(\RI5[0][143] ), .Z(n3529) );
  NAND3_X1 U8142 ( .A1(\SB1_1_24/i0[10] ), .A2(\SB1_1_24/i1_5 ), .A3(
        \SB1_1_24/i1[9] ), .ZN(\SB1_1_24/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 U8143 ( .I(\SB1_3_4/buf_output[5] ), .Z(\SB2_3_4/i0_3 ) );
  XOR2_X1 U8150 ( .A1(\RI5[3][57] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[51] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[57] ) );
  XOR2_X1 U8154 ( .A1(\MC_ARK_ARC_1_2/temp2[49] ), .A2(
        \MC_ARK_ARC_1_2/temp1[49] ), .Z(\MC_ARK_ARC_1_2/temp5[49] ) );
  XOR2_X1 U8186 ( .A1(n3535), .A2(\MC_ARK_ARC_1_1/temp2[188] ), .Z(n3540) );
  XOR2_X1 U8187 ( .A1(\RI5[1][182] ), .A2(\RI5[1][188] ), .Z(n3535) );
  NAND4_X2 U8189 ( .A1(\SB1_1_4/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_1_4/Component_Function_2/NAND4_in[3] ), .A3(
        \SB1_1_4/Component_Function_2/NAND4_in[0] ), .A4(n3536), .ZN(
        \RI3[1][182] ) );
  NAND3_X2 U8192 ( .A1(\SB1_1_4/i0[10] ), .A2(\SB1_1_4/i0[6] ), .A3(
        \SB1_1_4/i0_3 ), .ZN(n3536) );
  XOR2_X1 U8194 ( .A1(\MC_ARK_ARC_1_0/temp4[129] ), .A2(
        \MC_ARK_ARC_1_0/temp3[129] ), .Z(\MC_ARK_ARC_1_0/temp6[129] ) );
  XOR2_X1 U8206 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[165] ), .A2(\RI5[0][189] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[27] ) );
  NAND3_X2 U8212 ( .A1(\SB2_0_30/i0_0 ), .A2(\RI3[0][10] ), .A3(
        \SB2_0_30/i0_3 ), .ZN(\SB2_0_30/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U8216 ( .A1(\SB2_1_24/i0_0 ), .A2(\SB2_1_24/i1_5 ), .A3(
        \SB2_1_24/i0_4 ), .ZN(\SB2_1_24/Component_Function_2/NAND4_in[3] ) );
  XOR2_X1 U8221 ( .A1(\MC_ARK_ARC_1_1/temp4[190] ), .A2(
        \MC_ARK_ARC_1_1/temp3[190] ), .Z(n3541) );
  NAND4_X2 U8237 ( .A1(\SB1_0_27/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_27/Component_Function_5/NAND4_in[3] ), .A3(n2210), .A4(
        \SB1_0_27/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_0_27/buf_output[5] ) );
  XOR2_X1 U8243 ( .A1(\RI5[1][124] ), .A2(\RI5[1][130] ), .Z(n3543) );
  NAND3_X2 U8246 ( .A1(\SB2_3_6/i0[10] ), .A2(\SB2_3_6/i0_3 ), .A3(
        \SB2_3_6/i0[9] ), .ZN(\SB2_3_6/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U8250 ( .A1(\SB4_22/i0_3 ), .A2(\SB4_22/i1[9] ), .A3(\SB4_22/i0[6] ), .ZN(\SB4_22/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U8258 ( .A1(\SB3_31/i0_3 ), .A2(\SB3_31/i0[8] ), .A3(\SB3_31/i0[9] ), .ZN(\SB3_31/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 U8263 ( .A1(\SB2_3_8/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_8/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_3_8/Component_Function_5/NAND4_in[0] ), .A4(n3544), .ZN(
        \SB2_3_8/buf_output[5] ) );
  XOR2_X1 U8274 ( .A1(\MC_ARK_ARC_1_1/temp5[151] ), .A2(n3545), .Z(
        \MC_ARK_ARC_1_1/buf_output[151] ) );
  XOR2_X1 U8278 ( .A1(\MC_ARK_ARC_1_1/temp3[151] ), .A2(
        \MC_ARK_ARC_1_1/temp4[151] ), .Z(n3545) );
  INV_X2 U8288 ( .I(\RI3[0][80] ), .ZN(\SB2_0_18/i1[9] ) );
  NAND4_X2 U8290 ( .A1(\SB1_0_21/Component_Function_2/NAND4_in[0] ), .A2(n4650), .A3(\SB1_0_21/Component_Function_2/NAND4_in[2] ), .A4(n4651), .ZN(
        \RI3[0][80] ) );
  NAND4_X2 U8291 ( .A1(\SB1_2_7/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_7/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_7/Component_Function_4/NAND4_in[3] ), .A4(n3546), .ZN(
        \SB1_2_7/buf_output[4] ) );
  XOR2_X1 U8292 ( .A1(\RI5[2][159] ), .A2(\RI5[2][3] ), .Z(
        \MC_ARK_ARC_1_2/temp3[93] ) );
  XOR2_X1 U8297 ( .A1(n237), .A2(\MC_ARK_ARC_1_0/buf_datainput[36] ), .Z(n3547) );
  NAND4_X2 U8327 ( .A1(\SB2_0_4/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_0_4/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_0_4/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_4/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_0_4/buf_output[0] ) );
  NAND3_X2 U8336 ( .A1(\SB1_2_22/i0[10] ), .A2(\SB1_2_22/i1[9] ), .A3(
        \SB1_2_22/i1_7 ), .ZN(n1496) );
  NAND3_X1 U8339 ( .A1(\SB1_1_27/i0[8] ), .A2(\SB1_1_27/i0_4 ), .A3(
        \SB1_1_27/i1_7 ), .ZN(n3551) );
  NAND4_X2 U8340 ( .A1(\SB2_0_9/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_0_9/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_9/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_0_9/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_0_9/buf_output[0] ) );
  INV_X2 U8343 ( .I(\MC_ARK_ARC_1_0/buf_output[122] ), .ZN(\SB1_1_11/i1[9] )
         );
  INV_X2 U8351 ( .I(\SB1_3_16/buf_output[2] ), .ZN(\SB2_3_13/i1[9] ) );
  XOR2_X1 U8357 ( .A1(\MC_ARK_ARC_1_3/temp1[125] ), .A2(
        \MC_ARK_ARC_1_3/temp2[125] ), .Z(\MC_ARK_ARC_1_3/temp5[125] ) );
  NAND4_X2 U8358 ( .A1(\SB3_11/Component_Function_4/NAND4_in[3] ), .A2(n2039), 
        .A3(\SB3_11/Component_Function_4/NAND4_in[1] ), .A4(n3556), .ZN(
        \SB3_11/buf_output[4] ) );
  XOR2_X1 U8360 ( .A1(\RI5[3][37] ), .A2(\RI5[3][1] ), .Z(
        \MC_ARK_ARC_1_3/temp3[127] ) );
  XOR2_X1 U8365 ( .A1(\RI5[3][169] ), .A2(\RI5[3][145] ), .Z(
        \MC_ARK_ARC_1_3/temp2[7] ) );
  XOR2_X1 U8368 ( .A1(\MC_ARK_ARC_1_0/temp3[93] ), .A2(
        \MC_ARK_ARC_1_0/temp4[93] ), .Z(n3559) );
  XOR2_X1 U8371 ( .A1(\RI5[0][8] ), .A2(n5497), .Z(\MC_ARK_ARC_1_0/temp1[14] )
         );
  NAND3_X1 U8372 ( .A1(\SB2_1_29/i0[10] ), .A2(\SB2_1_29/i0_3 ), .A3(
        \SB2_1_29/i0_4 ), .ZN(\SB2_1_29/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U8375 ( .A1(\SB2_3_28/i0[6] ), .A2(\SB2_3_28/i0[8] ), .A3(
        \SB2_3_28/i0[7] ), .ZN(\SB2_3_28/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U8379 ( .A1(\SB2_0_12/i0[10] ), .A2(\SB2_0_12/i1_7 ), .A3(
        \SB2_0_12/i1[9] ), .ZN(\SB2_0_12/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U8380 ( .A1(\SB2_1_28/i0[10] ), .A2(\SB2_1_28/i0_0 ), .A3(
        \SB2_1_28/i0[6] ), .ZN(\SB2_1_28/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U8381 ( .A1(\MC_ARK_ARC_1_3/temp6[54] ), .A2(
        \MC_ARK_ARC_1_3/temp5[54] ), .Z(\MC_ARK_ARC_1_3/buf_output[54] ) );
  NAND4_X2 U8382 ( .A1(\SB1_2_7/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_2_7/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_2_7/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_2_7/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_2_7/buf_output[0] ) );
  NAND3_X2 U8386 ( .A1(\SB2_0_24/i0_3 ), .A2(\RI3[0][46] ), .A3(
        \SB2_0_24/i1[9] ), .ZN(n3561) );
  XOR2_X1 U8392 ( .A1(\MC_ARK_ARC_1_0/temp1[16] ), .A2(n2197), .Z(
        \MC_ARK_ARC_1_0/temp5[16] ) );
  NAND4_X2 U8393 ( .A1(\SB2_3_10/Component_Function_2/NAND4_in[2] ), .A2(n2677), .A3(\SB2_3_10/Component_Function_2/NAND4_in[1] ), .A4(n3565), .ZN(
        \SB2_3_10/buf_output[2] ) );
  NAND3_X1 U8395 ( .A1(\SB3_18/i0_0 ), .A2(\SB3_18/i3[0] ), .A3(\SB3_18/i1_7 ), 
        .ZN(\SB3_18/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U8399 ( .A1(n3569), .A2(n3568), .Z(\RI1[4][87] ) );
  XOR2_X1 U8400 ( .A1(n3699), .A2(\MC_ARK_ARC_1_3/temp4[87] ), .Z(n3568) );
  XOR2_X1 U8401 ( .A1(n1747), .A2(\MC_ARK_ARC_1_3/temp1[87] ), .Z(n3569) );
  NAND3_X1 U8410 ( .A1(\SB2_1_28/i0_4 ), .A2(\SB2_1_28/i1_7 ), .A3(
        \SB2_1_28/i0[8] ), .ZN(n3573) );
  NAND4_X2 U8411 ( .A1(\SB1_0_23/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_23/Component_Function_2/NAND4_in[3] ), .A3(n3642), .A4(n3574), 
        .ZN(\RI3[0][68] ) );
  XOR2_X1 U8413 ( .A1(\RI5[2][123] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[99] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[153] ) );
  NAND3_X1 U8414 ( .A1(\SB1_1_19/buf_output[1] ), .A2(\SB2_1_15/i1_5 ), .A3(
        \SB1_1_20/buf_output[0] ), .ZN(
        \SB2_1_15/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 U8417 ( .A1(\SB1_2_29/i0[8] ), .A2(\SB1_2_29/i0[9] ), .A3(
        \RI1[2][17] ), .ZN(n3575) );
  XOR2_X1 U8420 ( .A1(\RI5[3][106] ), .A2(\RI5[3][112] ), .Z(
        \MC_ARK_ARC_1_3/temp1[112] ) );
  XOR2_X1 U8421 ( .A1(\RI5[2][152] ), .A2(\RI5[2][188] ), .Z(
        \MC_ARK_ARC_1_2/temp3[86] ) );
  NAND3_X1 U8422 ( .A1(\SB1_2_8/i0_4 ), .A2(\SB1_2_8/i1[9] ), .A3(
        \SB1_2_8/i1_5 ), .ZN(\SB1_2_8/Component_Function_4/NAND4_in[3] ) );
  XOR2_X1 U8424 ( .A1(\MC_ARK_ARC_1_2/temp1[159] ), .A2(
        \MC_ARK_ARC_1_2/temp2[159] ), .Z(n3577) );
  BUF_X4 U8425 ( .I(\SB2_2_29/buf_output[1] ), .Z(\RI5[2][37] ) );
  BUF_X4 U8426 ( .I(\MC_ARK_ARC_1_0/buf_output[74] ), .Z(\SB1_1_19/i0_0 ) );
  XOR2_X1 U8427 ( .A1(n3772), .A2(\MC_ARK_ARC_1_1/temp1[151] ), .Z(
        \MC_ARK_ARC_1_1/temp5[151] ) );
  XOR2_X1 U8433 ( .A1(\MC_ARK_ARC_1_3/temp1[7] ), .A2(
        \MC_ARK_ARC_1_3/temp2[7] ), .Z(\MC_ARK_ARC_1_3/temp5[7] ) );
  NAND3_X2 U8436 ( .A1(\SB1_2_8/i0_3 ), .A2(\SB1_2_8/i1[9] ), .A3(
        \SB1_2_8/i0_4 ), .ZN(n976) );
  NAND3_X2 U8440 ( .A1(\SB2_3_15/i0[10] ), .A2(\SB2_3_15/i0_3 ), .A3(
        \SB2_3_15/i0[6] ), .ZN(\SB2_3_15/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U8443 ( .A1(\SB2_3_17/i0[6] ), .A2(\SB2_3_17/i0[10] ), .A3(
        \SB2_3_17/i0_0 ), .ZN(n3584) );
  NAND4_X2 U8444 ( .A1(\SB3_26/Component_Function_5/NAND4_in[1] ), .A2(
        \SB3_26/Component_Function_5/NAND4_in[3] ), .A3(
        \SB3_26/Component_Function_5/NAND4_in[0] ), .A4(n3585), .ZN(
        \SB3_26/buf_output[5] ) );
  NAND3_X1 U8449 ( .A1(\SB2_2_29/i0[7] ), .A2(\SB2_2_29/i0[8] ), .A3(
        \SB2_2_29/i0[6] ), .ZN(\SB2_2_29/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U8450 ( .A1(\MC_ARK_ARC_1_2/temp6[72] ), .A2(n4512), .Z(
        \MC_ARK_ARC_1_2/buf_output[72] ) );
  XOR2_X1 U8451 ( .A1(n3587), .A2(n21), .Z(Ciphertext[35]) );
  NAND4_X2 U8452 ( .A1(\SB4_26/Component_Function_5/NAND4_in[1] ), .A2(
        \SB4_26/Component_Function_5/NAND4_in[2] ), .A3(n2102), .A4(
        \SB4_26/Component_Function_5/NAND4_in[0] ), .ZN(n3587) );
  BUF_X4 U8455 ( .I(\MC_ARK_ARC_1_3/buf_output[71] ), .Z(\SB3_20/i0_3 ) );
  NAND3_X2 U8458 ( .A1(\SB1_3_16/i0_3 ), .A2(\SB1_3_16/i0[6] ), .A3(
        \SB1_3_16/i1[9] ), .ZN(n4616) );
  NAND3_X2 U8460 ( .A1(\SB2_2_13/i0[10] ), .A2(\SB2_2_13/i1[9] ), .A3(
        \SB2_2_13/i1_7 ), .ZN(\SB2_2_13/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U8461 ( .A1(\SB1_0_5/i0_0 ), .A2(\SB1_0_5/i1_5 ), .A3(
        \SB1_0_5/i0_4 ), .ZN(n4716) );
  NAND3_X1 U8462 ( .A1(\SB4_27/i1_5 ), .A2(\SB4_27/i3[0] ), .A3(\SB4_27/i0[8] ), .ZN(\SB4_27/Component_Function_3/NAND4_in[3] ) );
  NAND4_X2 U8467 ( .A1(\SB2_2_6/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_6/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_2_6/Component_Function_1/NAND4_in[1] ), .A4(
        \SB2_2_6/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_2_6/buf_output[1] ) );
  NAND4_X2 U8468 ( .A1(\SB1_0_26/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_0_26/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_0_26/Component_Function_4/NAND4_in[3] ), .A4(
        \SB1_0_26/Component_Function_4/NAND4_in[2] ), .ZN(
        \SB1_0_26/buf_output[4] ) );
  NAND3_X1 U8469 ( .A1(\SB2_1_24/i0_0 ), .A2(\SB2_1_24/i0[9] ), .A3(
        \SB2_1_24/i0[8] ), .ZN(\SB2_1_24/Component_Function_4/NAND4_in[0] ) );
  XOR2_X1 U8471 ( .A1(\MC_ARK_ARC_1_2/temp5[139] ), .A2(n3589), .Z(
        \MC_ARK_ARC_1_2/buf_output[139] ) );
  XOR2_X1 U8472 ( .A1(\MC_ARK_ARC_1_2/temp3[139] ), .A2(
        \MC_ARK_ARC_1_2/temp4[139] ), .Z(n3589) );
  XOR2_X1 U8473 ( .A1(\RI5[1][52] ), .A2(\RI5[1][16] ), .Z(
        \MC_ARK_ARC_1_1/temp3[142] ) );
  NAND3_X2 U8474 ( .A1(\SB3_11/i0_3 ), .A2(\SB3_11/i1[9] ), .A3(\SB3_11/i0_4 ), 
        .ZN(\SB3_11/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U8476 ( .A1(n3590), .A2(n73), .Z(Ciphertext[123]) );
  NAND4_X2 U8477 ( .A1(\SB4_11/Component_Function_3/NAND4_in[1] ), .A2(
        \SB4_11/Component_Function_3/NAND4_in[0] ), .A3(
        \SB4_11/Component_Function_3/NAND4_in[2] ), .A4(
        \SB4_11/Component_Function_3/NAND4_in[3] ), .ZN(n3590) );
  NAND3_X1 U8480 ( .A1(\SB1_2_6/i0_3 ), .A2(\SB1_2_6/i0[8] ), .A3(
        \SB1_2_6/i1_7 ), .ZN(\SB1_2_6/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U8484 ( .A1(\MC_ARK_ARC_1_2/temp5[157] ), .A2(n683), .Z(
        \MC_ARK_ARC_1_2/buf_output[157] ) );
  XOR2_X1 U8486 ( .A1(\MC_ARK_ARC_1_0/temp3[4] ), .A2(
        \MC_ARK_ARC_1_0/temp4[4] ), .Z(\MC_ARK_ARC_1_0/temp6[4] ) );
  XOR2_X1 U8500 ( .A1(n3596), .A2(n799), .Z(\MC_ARK_ARC_1_1/buf_output[84] )
         );
  XOR2_X1 U8501 ( .A1(\MC_ARK_ARC_1_1/temp3[84] ), .A2(
        \MC_ARK_ARC_1_1/temp4[84] ), .Z(n3596) );
  NAND3_X1 U8503 ( .A1(\SB4_7/i0_3 ), .A2(\SB4_7/i0_4 ), .A3(\SB4_7/i0[10] ), 
        .ZN(n3597) );
  NAND4_X2 U8512 ( .A1(\SB2_0_26/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_0_26/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_0_26/Component_Function_1/NAND4_in[3] ), .A4(n3602), .ZN(
        \SB2_0_26/buf_output[1] ) );
  NAND2_X1 U8513 ( .A1(\SB2_0_26/i0_3 ), .A2(\SB2_0_26/i1[9] ), .ZN(n3602) );
  NAND3_X1 U8515 ( .A1(\SB4_16/i3[0] ), .A2(\SB4_16/i0[8] ), .A3(\SB4_16/i1_5 ), .ZN(\SB4_16/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U8521 ( .A1(n3607), .A2(n4107), .Z(\MC_ARK_ARC_1_3/temp5[47] ) );
  XOR2_X1 U8522 ( .A1(\RI5[3][185] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[17] ), 
        .Z(n3607) );
  XOR2_X1 U8523 ( .A1(n3608), .A2(\MC_ARK_ARC_1_1/temp5[129] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[129] ) );
  XOR2_X1 U8524 ( .A1(\MC_ARK_ARC_1_1/temp4[129] ), .A2(
        \MC_ARK_ARC_1_1/temp3[129] ), .Z(n3608) );
  NAND4_X2 U8527 ( .A1(\SB1_3_28/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_3_28/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_28/Component_Function_0/NAND4_in[0] ), .A4(n3610), .ZN(
        \SB1_3_28/buf_output[0] ) );
  XOR2_X1 U8528 ( .A1(\MC_ARK_ARC_1_3/temp1[127] ), .A2(n3611), .Z(n1576) );
  XOR2_X1 U8529 ( .A1(\RI5[3][73] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[97] ), 
        .Z(n3611) );
  NAND3_X2 U8530 ( .A1(\SB1_2_19/i0_3 ), .A2(\SB1_2_19/i0[9] ), .A3(
        \SB1_2_19/i0[8] ), .ZN(n4499) );
  NAND4_X2 U8531 ( .A1(\SB2_1_25/Component_Function_2/NAND4_in[1] ), .A2(n4517), .A3(n4724), .A4(n3612), .ZN(\SB2_1_25/buf_output[2] ) );
  NAND3_X2 U8535 ( .A1(\SB2_3_31/i0_3 ), .A2(\SB2_3_31/i0[6] ), .A3(
        \SB2_3_31/i1[9] ), .ZN(\SB2_3_31/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U8537 ( .A1(\SB1_2_6/i0_3 ), .A2(\SB1_2_6/i0_4 ), .A3(
        \SB1_2_6/i1[9] ), .ZN(n3614) );
  NAND3_X2 U8538 ( .A1(\SB2_1_7/i0_3 ), .A2(\SB2_1_7/i1[9] ), .A3(n5790), .ZN(
        \SB2_1_7/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U8540 ( .A1(\SB2_2_18/i0_4 ), .A2(n4769), .A3(\SB2_2_18/i0_0 ), 
        .ZN(n3616) );
  NAND3_X1 U8541 ( .A1(\SB1_2_11/i0_0 ), .A2(\SB1_2_11/i1_7 ), .A3(
        \SB1_2_11/i3[0] ), .ZN(n2088) );
  BUF_X4 U8542 ( .I(\SB1_3_10/buf_output[5] ), .Z(\SB2_3_10/i0_3 ) );
  INV_X2 U8543 ( .I(\SB1_1_7/buf_output[5] ), .ZN(\SB2_1_7/i1_5 ) );
  INV_X2 U8546 ( .I(\MC_ARK_ARC_1_3/buf_output[105] ), .ZN(\SB3_14/i0[8] ) );
  NAND4_X2 U8549 ( .A1(n1420), .A2(n1196), .A3(
        \SB3_13/Component_Function_3/NAND4_in[0] ), .A4(n3617), .ZN(
        \SB3_13/buf_output[3] ) );
  INV_X2 U8552 ( .I(\SB1_3_10/buf_output[5] ), .ZN(\SB2_3_10/i1_5 ) );
  NAND2_X1 U8554 ( .A1(\SB4_11/i0[10] ), .A2(\SB4_11/i0[9] ), .ZN(n4216) );
  XOR2_X1 U8556 ( .A1(n3620), .A2(n1962), .Z(\MC_ARK_ARC_1_1/buf_output[8] )
         );
  XOR2_X1 U8557 ( .A1(n2739), .A2(n3990), .Z(n3620) );
  XOR2_X1 U8558 ( .A1(n4739), .A2(n4740), .Z(n3688) );
  XOR2_X1 U8559 ( .A1(\MC_ARK_ARC_1_3/temp2[110] ), .A2(
        \MC_ARK_ARC_1_3/temp4[110] ), .Z(n4739) );
  XOR2_X1 U8561 ( .A1(\RI5[0][122] ), .A2(\RI5[0][146] ), .Z(
        \MC_ARK_ARC_1_0/temp2[176] ) );
  XOR2_X1 U8564 ( .A1(\RI5[2][23] ), .A2(\RI5[2][179] ), .Z(
        \MC_ARK_ARC_1_2/temp3[113] ) );
  NAND4_X2 U8569 ( .A1(\SB2_0_21/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_0_21/Component_Function_0/NAND4_in[1] ), .A3(n1077), .A4(
        \SB2_0_21/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_0_21/buf_output[0] ) );
  NAND2_X2 U8570 ( .A1(\SB1_3_31/i0_0 ), .A2(\SB1_3_31/i3[0] ), .ZN(
        \SB1_3_31/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 U8571 ( .I(\SB1_3_31/buf_output[5] ), .Z(\SB2_3_31/i0_3 ) );
  NAND3_X1 U8580 ( .A1(\SB4_11/i0_0 ), .A2(\SB4_11/i0[9] ), .A3(\SB4_11/i0[8] ), .ZN(n3626) );
  INV_X2 U8582 ( .I(\SB1_3_31/buf_output[5] ), .ZN(\SB2_3_31/i1_5 ) );
  NAND3_X2 U8584 ( .A1(\SB2_0_3/i0[10] ), .A2(\SB2_0_3/i0_0 ), .A3(
        \SB2_0_3/i0[6] ), .ZN(\SB2_0_3/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U8585 ( .A1(\SB1_0_5/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_5/Component_Function_3/NAND4_in[3] ), .A3(
        \SB1_0_5/Component_Function_3/NAND4_in[1] ), .A4(n3627), .ZN(
        \SB1_0_5/buf_output[3] ) );
  INV_X2 U8589 ( .I(\SB1_2_11/buf_output[3] ), .ZN(\SB2_2_9/i0[8] ) );
  BUF_X4 U8592 ( .I(\MC_ARK_ARC_1_0/buf_output[191] ), .Z(\SB1_1_0/i0_3 ) );
  INV_X2 U8595 ( .I(\MC_ARK_ARC_1_0/buf_output[191] ), .ZN(\SB1_1_0/i1_5 ) );
  NAND3_X2 U8598 ( .A1(\SB2_1_17/i0[6] ), .A2(\SB2_1_17/i0[9] ), .A3(
        \SB2_1_17/i0_4 ), .ZN(n3631) );
  NAND4_X2 U8602 ( .A1(\SB1_1_24/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_1_24/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_1_24/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_1_24/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_1_24/buf_output[0] ) );
  XOR2_X1 U8603 ( .A1(n1642), .A2(n1641), .Z(\MC_ARK_ARC_1_1/buf_output[157] )
         );
  XOR2_X1 U8605 ( .A1(n1584), .A2(n4339), .Z(n3634) );
  XOR2_X1 U8606 ( .A1(\MC_ARK_ARC_1_2/temp2[26] ), .A2(
        \MC_ARK_ARC_1_2/temp4[26] ), .Z(n3635) );
  XOR2_X1 U8611 ( .A1(n3639), .A2(n3638), .Z(n1908) );
  XOR2_X1 U8612 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[131] ), .A2(n198), .Z(
        n3638) );
  XOR2_X1 U8613 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[65] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[95] ), .Z(n3639) );
  XOR2_X1 U8614 ( .A1(\MC_ARK_ARC_1_0/temp5[8] ), .A2(n3640), .Z(
        \MC_ARK_ARC_1_0/buf_output[8] ) );
  XOR2_X1 U8615 ( .A1(n3766), .A2(\MC_ARK_ARC_1_0/temp4[8] ), .Z(n3640) );
  NAND4_X2 U8616 ( .A1(\SB1_1_30/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_1_30/Component_Function_2/NAND4_in[1] ), .A3(n1414), .A4(n3641), 
        .ZN(\SB1_1_30/buf_output[2] ) );
  NAND3_X2 U8617 ( .A1(\SB1_1_30/i0[10] ), .A2(\SB1_1_30/i1[9] ), .A3(
        \SB1_1_30/i1_5 ), .ZN(n3641) );
  NAND4_X2 U8619 ( .A1(\SB2_0_20/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_20/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_0_20/Component_Function_2/NAND4_in[1] ), .A4(n3643), .ZN(
        \SB2_0_20/buf_output[2] ) );
  NAND3_X2 U8620 ( .A1(\SB2_0_20/i0_0 ), .A2(\SB2_0_20/i1_5 ), .A3(
        \SB2_0_20/i0_4 ), .ZN(n3643) );
  XOR2_X1 U8621 ( .A1(\MC_ARK_ARC_1_0/temp6[82] ), .A2(n3644), .Z(
        \MC_ARK_ARC_1_0/buf_output[82] ) );
  XOR2_X1 U8622 ( .A1(n4575), .A2(\MC_ARK_ARC_1_0/temp1[82] ), .Z(n3644) );
  BUF_X2 U8623 ( .I(\SB2_1_30/buf_output[5] ), .Z(\RI5[1][11] ) );
  BUF_X4 U8628 ( .I(n411), .Z(\SB1_0_25/i0_3 ) );
  BUF_X4 U8630 ( .I(\MC_ARK_ARC_1_1/buf_output[11] ), .Z(\SB1_2_30/i0_3 ) );
  BUF_X4 U8631 ( .I(\SB2_3_1/buf_output[1] ), .Z(\RI5[3][13] ) );
  BUF_X4 U8632 ( .I(\SB2_3_6/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[165] ) );
  NAND3_X1 U8634 ( .A1(\SB4_20/i0_3 ), .A2(\SB4_20/i1_7 ), .A3(\SB4_20/i0[8] ), 
        .ZN(\SB4_20/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 U8635 ( .A1(\SB4_20/i0_3 ), .A2(\SB4_20/i1[9] ), .ZN(
        \SB4_20/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U8636 ( .A1(\SB4_20/i0_3 ), .A2(\SB4_20/i0[9] ), .A3(\SB4_20/i0[8] ), .ZN(\SB4_20/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U8637 ( .A1(\SB4_20/i0_3 ), .A2(\SB4_20/i0[6] ), .A3(\SB4_20/i1[9] ), .ZN(\SB4_20/Component_Function_3/NAND4_in[0] ) );
  NAND2_X1 U8642 ( .A1(\SB3_14/i0_3 ), .A2(\SB3_14/i1[9] ), .ZN(
        \SB3_14/Component_Function_1/NAND4_in[0] ) );
  INV_X2 U8647 ( .I(\MC_ARK_ARC_1_2/buf_output[159] ), .ZN(\SB1_3_5/i0[8] ) );
  CLKBUF_X4 U8649 ( .I(\MC_ARK_ARC_1_3/buf_output[46] ), .Z(\SB3_24/i0_4 ) );
  NAND2_X1 U8650 ( .A1(\SB4_21/i0[10] ), .A2(\SB4_21/i0[9] ), .ZN(n4402) );
  NAND3_X1 U8653 ( .A1(\SB3_3/i1[9] ), .A2(\SB3_3/i0_4 ), .A3(\SB3_3/i0_3 ), 
        .ZN(\SB3_3/Component_Function_5/NAND4_in[2] ) );
  CLKBUF_X4 U8654 ( .I(\SB1_2_28/buf_output[0] ), .Z(\SB2_2_23/i0[9] ) );
  XOR2_X1 U8656 ( .A1(\MC_ARK_ARC_1_3/temp6[147] ), .A2(
        \MC_ARK_ARC_1_3/temp5[147] ), .Z(n3646) );
  NAND3_X1 U8658 ( .A1(\SB1_2_26/i0[10] ), .A2(\SB1_2_26/i1_5 ), .A3(
        \SB1_2_26/i1[9] ), .ZN(\SB1_2_26/Component_Function_2/NAND4_in[0] ) );
  BUF_X2 U8661 ( .I(\SB3_3/buf_output[3] ), .Z(\SB4_1/i0[10] ) );
  CLKBUF_X4 U8664 ( .I(\SB1_2_27/buf_output[2] ), .Z(\SB2_2_24/i0_0 ) );
  CLKBUF_X4 U8665 ( .I(\MC_ARK_ARC_1_3/buf_output[64] ), .Z(\SB3_21/i0_4 ) );
  NAND3_X1 U8673 ( .A1(\SB3_3/i0[8] ), .A2(\SB3_3/i1_5 ), .A3(\SB3_3/i3[0] ), 
        .ZN(n1799) );
  CLKBUF_X4 U8677 ( .I(\SB2_2_13/buf_output[3] ), .Z(\RI5[2][123] ) );
  BUF_X2 U8679 ( .I(\MC_ARK_ARC_1_3/buf_output[49] ), .Z(\SB3_23/i0[6] ) );
  NAND3_X1 U8680 ( .A1(\SB3_23/i0[10] ), .A2(\SB3_23/i0_0 ), .A3(
        \SB3_23/i0[6] ), .ZN(\SB3_23/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U8681 ( .A1(\SB3_23/i0[6] ), .A2(\SB3_23/i0[8] ), .A3(
        \SB3_23/i0[7] ), .ZN(n946) );
  NAND3_X1 U8682 ( .A1(\SB4_31/i0[10] ), .A2(\SB4_31/i1[9] ), .A3(
        \SB4_31/i1_7 ), .ZN(\SB4_31/Component_Function_3/NAND4_in[2] ) );
  INV_X1 U8685 ( .I(\MC_ARK_ARC_1_2/buf_output[124] ), .ZN(n3648) );
  CLKBUF_X4 U8686 ( .I(\MC_ARK_ARC_1_3/buf_output[112] ), .Z(\SB3_13/i0_4 ) );
  BUF_X4 U8687 ( .I(\SB2_2_19/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[97] ) );
  NAND3_X1 U8689 ( .A1(\SB2_3_0/i1[9] ), .A2(\SB2_3_0/i1_5 ), .A3(
        \SB1_3_1/buf_output[4] ), .ZN(
        \SB2_3_0/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U8693 ( .A1(\SB2_3_26/i1[9] ), .A2(\SB2_3_26/i0_3 ), .A3(
        \SB2_3_26/i0[6] ), .ZN(\SB2_3_26/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U8694 ( .A1(\SB2_3_26/i0_3 ), .A2(\SB2_3_26/i0_0 ), .A3(
        \SB2_3_26/i0_4 ), .ZN(\SB2_3_26/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U8697 ( .A1(\SB1_2_3/i0_4 ), .A2(\SB1_2_3/i1[9] ), .A3(
        \SB1_2_3/i0_3 ), .ZN(\SB1_2_3/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U8700 ( .A1(\SB4_13/i0_4 ), .A2(\SB4_13/i1[9] ), .A3(\SB4_13/i1_5 ), 
        .ZN(n901) );
  BUF_X2 U8701 ( .I(\MC_ARK_ARC_1_1/buf_output[187] ), .Z(\SB1_2_0/i0[6] ) );
  INV_X1 U8702 ( .I(\MC_ARK_ARC_1_1/buf_output[187] ), .ZN(\SB1_2_0/i1_7 ) );
  INV_X1 U8706 ( .I(\MC_ARK_ARC_1_3/buf_output[83] ), .ZN(\SB3_18/i1_5 ) );
  NAND3_X1 U8708 ( .A1(\SB3_17/i0[7] ), .A2(\SB3_17/i0_3 ), .A3(\SB3_17/i0_0 ), 
        .ZN(\SB3_17/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U8712 ( .A1(\SB1_1_13/i0_3 ), .A2(\SB1_1_13/i1_7 ), .A3(
        \SB1_1_13/i0[8] ), .ZN(\SB1_1_13/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U8713 ( .A1(\SB3_10/i0_3 ), .A2(\SB3_10/i1[9] ), .A3(\SB3_10/i0_4 ), 
        .ZN(n2367) );
  BUF_X4 U8714 ( .I(\MC_ARK_ARC_1_3/buf_output[149] ), .Z(\SB3_7/i0_3 ) );
  INV_X1 U8715 ( .I(\MC_ARK_ARC_1_3/buf_output[66] ), .ZN(\SB3_20/i3[0] ) );
  NAND3_X1 U8717 ( .A1(\SB1_3_17/i1_5 ), .A2(\SB1_3_17/i0[10] ), .A3(
        \SB1_3_17/i1[9] ), .ZN(\SB1_3_17/Component_Function_2/NAND4_in[0] ) );
  INV_X1 U8719 ( .I(\MC_ARK_ARC_1_0/buf_output[94] ), .ZN(\SB1_1_16/i0[7] ) );
  BUF_X4 U8722 ( .I(\MC_ARK_ARC_1_2/buf_output[47] ), .Z(\SB1_3_24/i0_3 ) );
  NAND3_X1 U8727 ( .A1(\SB3_15/i0_3 ), .A2(\SB3_15/i0[8] ), .A3(\SB3_15/i0[9] ), .ZN(\SB3_15/Component_Function_2/NAND4_in[2] ) );
  CLKBUF_X8 U8728 ( .I(\MC_ARK_ARC_1_3/buf_output[101] ), .Z(\SB3_15/i0_3 ) );
  NAND2_X1 U8729 ( .A1(\SB1_2_26/i0[10] ), .A2(\SB1_2_26/i0[9] ), .ZN(
        \SB1_2_26/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U8730 ( .A1(\SB1_2_26/i0[10] ), .A2(\RI1[2][35] ), .A3(
        \SB1_2_26/i0[6] ), .ZN(\SB1_2_26/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U8731 ( .A1(\SB1_2_26/i0[10] ), .A2(\RI1[2][35] ), .A3(
        \SB1_2_26/i0[9] ), .ZN(n1717) );
  NAND3_X1 U8732 ( .A1(\SB1_2_26/i0[10] ), .A2(\SB1_2_26/i1[9] ), .A3(
        \SB1_2_26/i1_7 ), .ZN(n1574) );
  NAND3_X1 U8734 ( .A1(\SB4_11/i0[10] ), .A2(\SB4_11/i1[9] ), .A3(
        \SB4_11/i1_7 ), .ZN(\SB4_11/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U8735 ( .A1(\SB4_11/i0[10] ), .A2(n3684), .A3(\SB4_11/i1[9] ), .ZN(
        n2686) );
  CLKBUF_X2 U8737 ( .I(Key[119]), .Z(n237) );
  NAND3_X1 U8739 ( .A1(\SB1_2_11/i0_3 ), .A2(\SB1_2_11/i1_7 ), .A3(
        \SB1_2_11/i0[8] ), .ZN(\SB1_2_11/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U8741 ( .A1(\SB3_26/i1_5 ), .A2(\SB3_26/i0[8] ), .A3(\SB3_26/i3[0] ), .ZN(\SB3_26/Component_Function_3/NAND4_in[3] ) );
  BUF_X2 U8743 ( .I(\SB3_19/buf_output[3] ), .Z(\SB4_17/i0[10] ) );
  NAND3_X1 U8745 ( .A1(\SB4_13/i0_3 ), .A2(\SB4_13/i0[6] ), .A3(\SB4_13/i1[9] ), .ZN(\SB4_13/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U8746 ( .A1(\SB4_13/i0_3 ), .A2(\SB4_13/i0_0 ), .A3(\SB4_13/i0[7] ), 
        .ZN(n4746) );
  NAND3_X1 U8749 ( .A1(\SB2_1_5/i0_3 ), .A2(\SB2_1_5/i1_7 ), .A3(
        \SB2_1_5/i0[8] ), .ZN(\SB2_1_5/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U8750 ( .A1(n2535), .A2(\SB2_1_5/i0_0 ), .A3(\SB2_1_5/i0_3 ), .ZN(
        \SB2_1_5/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 U8755 ( .A1(\SB4_20/i0_0 ), .A2(\SB4_20/i3[0] ), .ZN(
        \SB4_20/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U8756 ( .A1(\SB4_20/i3[0] ), .A2(\SB4_20/i0_0 ), .A3(\SB4_20/i1_7 ), 
        .ZN(\SB4_20/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U8758 ( .A1(\SB4_19/i1_5 ), .A2(\SB4_19/i0[6] ), .A3(\SB4_19/i0[9] ), .ZN(\SB4_19/Component_Function_1/NAND4_in[2] ) );
  INV_X1 U8759 ( .I(\SB3_1/buf_output[1] ), .ZN(\SB4_29/i1_7 ) );
  CLKBUF_X12 U8760 ( .I(Key[155]), .Z(n104) );
  BUF_X2 U8763 ( .I(\MC_ARK_ARC_1_3/buf_output[109] ), .Z(\SB3_13/i0[6] ) );
  INV_X1 U8764 ( .I(\MC_ARK_ARC_1_3/buf_output[109] ), .ZN(\SB3_13/i1_7 ) );
  NAND2_X1 U8767 ( .A1(\SB4_11/i0_0 ), .A2(\SB4_11/i3[0] ), .ZN(
        \SB4_11/Component_Function_5/NAND4_in[0] ) );
  CLKBUF_X12 U8772 ( .I(Key[14]), .Z(n147) );
  CLKBUF_X4 U8773 ( .I(\SB3_21/buf_output[4] ), .Z(\SB4_20/i0_4 ) );
  NAND2_X1 U8775 ( .A1(\SB3_27/i0_0 ), .A2(\SB3_27/i3[0] ), .ZN(
        \SB3_27/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U8778 ( .A1(\SB2_2_29/i0_0 ), .A2(\SB2_2_29/i1_5 ), .A3(n1837), 
        .ZN(n4501) );
  NAND3_X1 U8780 ( .A1(\SB3_21/buf_output[3] ), .A2(\SB4_19/i1[9] ), .A3(
        \SB4_19/i1_7 ), .ZN(n1228) );
  BUF_X2 U8782 ( .I(\SB3_19/buf_output[0] ), .Z(\SB4_14/i0[9] ) );
  INV_X1 U8783 ( .I(\SB3_19/buf_output[0] ), .ZN(\SB4_14/i3[0] ) );
  NAND3_X1 U8784 ( .A1(\SB1_1_27/i0[8] ), .A2(\SB1_1_27/i1_5 ), .A3(
        \SB1_1_27/i3[0] ), .ZN(n4376) );
  NAND3_X1 U8789 ( .A1(\SB4_28/i0[10] ), .A2(\SB4_28/i1_5 ), .A3(n5514), .ZN(
        \SB4_28/Component_Function_2/NAND4_in[0] ) );
  NAND2_X1 U8790 ( .A1(\SB4_28/i0[10] ), .A2(\SB4_28/i0[9] ), .ZN(
        \SB4_28/Component_Function_0/NAND4_in[0] ) );
  CLKBUF_X4 U8791 ( .I(\MC_ARK_ARC_1_3/buf_output[70] ), .Z(\SB3_20/i0_4 ) );
  NAND2_X1 U8794 ( .A1(\SB4_8/i0_0 ), .A2(\SB4_8/i3[0] ), .ZN(
        \SB4_8/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U8800 ( .A1(\SB1_1_16/i0_4 ), .A2(\SB1_1_16/i0_0 ), .A3(
        \SB1_1_16/i1_5 ), .ZN(n3860) );
  NAND3_X1 U8801 ( .A1(\SB1_1_16/i0[7] ), .A2(\SB1_1_16/i0_3 ), .A3(
        \SB1_1_16/i0_0 ), .ZN(\SB1_1_16/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U8804 ( .A1(\SB3_5/buf_output[3] ), .A2(\SB4_3/i0_3 ), .A3(
        \SB4_3/i0[9] ), .ZN(n3926) );
  NAND3_X1 U8811 ( .A1(\SB3_28/i0_3 ), .A2(\SB3_28/i0[8] ), .A3(\SB3_28/i0[9] ), .ZN(\SB3_28/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U8813 ( .A1(\SB1_1_3/i1_5 ), .A2(\SB1_1_3/i0[10] ), .A3(
        \SB1_1_3/i1[9] ), .ZN(\SB1_1_3/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U8818 ( .A1(\SB3_26/i1[9] ), .A2(\SB3_26/i0_3 ), .A3(\SB3_26/i0[6] ), .ZN(\SB3_26/Component_Function_3/NAND4_in[0] ) );
  INV_X2 U8820 ( .I(\MC_ARK_ARC_1_1/buf_output[139] ), .ZN(\SB1_2_8/i1_7 ) );
  CLKBUF_X4 U8821 ( .I(\SB3_27/buf_output[4] ), .Z(\SB4_26/i0_4 ) );
  AND4_X2 U8823 ( .A1(\SB3_1/Component_Function_3/NAND4_in[1] ), .A2(
        \SB3_1/Component_Function_3/NAND4_in[0] ), .A3(n1021), .A4(n4668), .Z(
        n3652) );
  NAND2_X1 U8827 ( .A1(\SB4_14/i0_3 ), .A2(\SB4_14/i1[9] ), .ZN(
        \SB4_14/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U8828 ( .A1(\SB4_14/i0_3 ), .A2(\SB4_14/i0[10] ), .A3(
        \SB4_14/i0[6] ), .ZN(\SB4_14/Component_Function_2/NAND4_in[1] ) );
  CLKBUF_X4 U8834 ( .I(\RI3[4][105] ), .Z(\SB4_14/i0[10] ) );
  NAND3_X1 U8837 ( .A1(\SB3_30/i0_3 ), .A2(\SB3_30/i0[7] ), .A3(\SB3_30/i0_0 ), 
        .ZN(\SB3_30/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 U8839 ( .A1(\SB4_30/i0_0 ), .A2(\SB4_30/i3[0] ), .ZN(
        \SB4_30/Component_Function_5/NAND4_in[0] ) );
  BUF_X2 U8843 ( .I(\MC_ARK_ARC_1_2/buf_output[102] ), .Z(\SB1_3_14/i0[9] ) );
  INV_X1 U8844 ( .I(\MC_ARK_ARC_1_2/buf_output[102] ), .ZN(\SB1_3_14/i3[0] )
         );
  INV_X1 U8847 ( .I(\SB1_3_24/buf_output[0] ), .ZN(\SB2_3_19/i3[0] ) );
  CLKBUF_X4 U8848 ( .I(\SB1_3_24/buf_output[0] ), .Z(\SB2_3_19/i0[9] ) );
  NAND3_X1 U8850 ( .A1(\SB3_8/i1[9] ), .A2(\SB3_8/i1_5 ), .A3(\SB3_8/i0_4 ), 
        .ZN(\SB3_8/Component_Function_4/NAND4_in[3] ) );
  AND4_X2 U8852 ( .A1(\SB3_7/Component_Function_2/NAND4_in[1] ), .A2(
        \SB3_7/Component_Function_2/NAND4_in[3] ), .A3(
        \SB3_7/Component_Function_2/NAND4_in[0] ), .A4(n4727), .Z(n3655) );
  INV_X1 U8856 ( .I(\MC_ARK_ARC_1_3/buf_output[35] ), .ZN(\SB3_26/i1_5 ) );
  NAND3_X1 U8858 ( .A1(\SB1_1_5/i0[9] ), .A2(\SB1_1_5/i0[10] ), .A3(
        \SB1_1_5/i0_3 ), .ZN(\SB1_1_5/Component_Function_4/NAND4_in[2] ) );
  CLKBUF_X4 U8859 ( .I(\MC_ARK_ARC_1_0/buf_output[159] ), .Z(\SB1_1_5/i0[10] )
         );
  CLKBUF_X4 U8862 ( .I(\SB3_14/buf_output[2] ), .Z(\SB4_11/i0_0 ) );
  NAND3_X1 U8863 ( .A1(\SB1_3_28/i0[10] ), .A2(\SB1_3_28/i0_3 ), .A3(
        \SB1_3_28/i0_4 ), .ZN(\SB1_3_28/Component_Function_0/NAND4_in[2] ) );
  INV_X1 U8867 ( .I(\MC_ARK_ARC_1_1/buf_output[67] ), .ZN(\SB1_2_20/i1_7 ) );
  CLKBUF_X4 U8868 ( .I(\MC_ARK_ARC_1_3/buf_output[56] ), .Z(\SB3_22/i0_0 ) );
  INV_X1 U8871 ( .I(\SB3_16/buf_output[0] ), .ZN(\SB4_11/i3[0] ) );
  NAND3_X1 U8872 ( .A1(\SB3_10/i1_7 ), .A2(\SB3_10/i0_0 ), .A3(\SB3_10/i3[0] ), 
        .ZN(\SB3_10/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U8873 ( .A1(\SB3_10/i1_5 ), .A2(\SB3_10/i0_0 ), .A3(\SB3_10/i0_4 ), 
        .ZN(\SB3_10/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U8874 ( .A1(\SB3_10/i0_0 ), .A2(\SB3_10/i0_3 ), .A3(\SB3_10/i0_4 ), 
        .ZN(\SB3_10/Component_Function_3/NAND4_in[1] ) );
  AND4_X2 U8881 ( .A1(\SB3_19/Component_Function_3/NAND4_in[0] ), .A2(n2412), 
        .A3(n4351), .A4(n4159), .Z(n3661) );
  INV_X1 U8882 ( .I(\SB1_1_9/buf_output[1] ), .ZN(\SB2_1_5/i1_7 ) );
  NAND3_X1 U8884 ( .A1(\SB3_30/i1_5 ), .A2(\SB3_30/i0[6] ), .A3(\SB3_30/i0[9] ), .ZN(\SB3_30/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U8885 ( .A1(\SB3_30/i0_3 ), .A2(\SB3_30/i0[10] ), .A3(
        \SB3_30/i0[9] ), .ZN(\SB3_30/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U8886 ( .A1(\SB2_3_11/i3[0] ), .A2(\SB2_3_11/i0[8] ), .A3(n4768), 
        .ZN(\SB2_3_11/Component_Function_3/NAND4_in[3] ) );
  INV_X1 U8892 ( .I(\MC_ARK_ARC_1_3/buf_output[7] ), .ZN(\SB3_30/i1_7 ) );
  NAND3_X1 U8894 ( .A1(\SB3_28/i0_0 ), .A2(\SB3_28/i1_5 ), .A3(\SB3_28/i0_4 ), 
        .ZN(\SB3_28/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U8895 ( .A1(\SB3_28/i0_0 ), .A2(\SB3_28/i0[6] ), .A3(
        \SB3_28/i0[10] ), .ZN(\SB3_28/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 U8896 ( .A1(\SB3_28/i0_0 ), .A2(\SB3_28/i3[0] ), .ZN(
        \SB3_28/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U8899 ( .A1(n1793), .A2(\SB4_29/i1[9] ), .A3(\SB4_29/i1_5 ), .ZN(
        \SB4_29/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U8901 ( .A1(\SB1_3_8/i1_5 ), .A2(\SB1_3_8/i1[9] ), .A3(
        \MC_ARK_ARC_1_2/buf_output[142] ), .ZN(n2442) );
  NAND3_X1 U8903 ( .A1(\SB3_19/i0[8] ), .A2(\SB3_19/i3[0] ), .A3(\SB3_19/i1_5 ), .ZN(n4159) );
  NAND3_X1 U8905 ( .A1(\SB1_1_14/i0[8] ), .A2(\SB1_1_14/i0[9] ), .A3(
        \SB1_1_14/i0_3 ), .ZN(\SB1_1_14/Component_Function_2/NAND4_in[2] ) );
  INV_X1 U8906 ( .I(\MC_ARK_ARC_1_2/buf_output[73] ), .ZN(\SB1_3_19/i1_7 ) );
  INV_X1 U8908 ( .I(\MC_ARK_ARC_1_3/buf_output[90] ), .ZN(\SB3_16/i3[0] ) );
  CLKBUF_X4 U8910 ( .I(\SB3_19/buf_output[2] ), .Z(\SB4_16/i0_0 ) );
  NAND3_X1 U8916 ( .A1(\SB3_17/i0_0 ), .A2(\SB3_17/i0_4 ), .A3(\SB3_17/i1_5 ), 
        .ZN(\SB3_17/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U8919 ( .A1(\SB4_14/i0[9] ), .A2(\SB4_14/i0_0 ), .A3(\SB4_14/i0[8] ), .ZN(\SB4_14/Component_Function_4/NAND4_in[0] ) );
  NAND2_X1 U8920 ( .A1(\SB4_14/i0_0 ), .A2(\SB4_14/i3[0] ), .ZN(
        \SB4_14/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U8924 ( .A1(\SB4_20/i0[10] ), .A2(\SB4_20/i0_4 ), .A3(\SB4_20/i0_3 ), .ZN(\SB4_20/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U8925 ( .A1(n3674), .A2(\SB4_20/i0[10] ), .A3(\SB4_20/i1[9] ), .ZN(
        \SB4_20/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U8926 ( .A1(\SB2_3_16/i1[9] ), .A2(\SB2_3_16/i1_5 ), .A3(
        \SB2_3_16/i0_4 ), .ZN(\SB2_3_16/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U8927 ( .A1(\SB2_3_16/i0_3 ), .A2(\SB2_3_16/i1[9] ), .A3(
        \SB2_3_16/i0[6] ), .ZN(\SB2_3_16/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U8928 ( .A1(\SB2_3_16/i0[10] ), .A2(\SB2_3_16/i1_5 ), .A3(
        \SB2_3_16/i1[9] ), .ZN(\SB2_3_16/Component_Function_2/NAND4_in[0] ) );
  NAND2_X1 U8929 ( .A1(\SB2_3_16/i0_3 ), .A2(\SB2_3_16/i1[9] ), .ZN(
        \SB2_3_16/Component_Function_1/NAND4_in[0] ) );
  CLKBUF_X4 U8934 ( .I(\SB1_3_1/buf_output[3] ), .Z(\SB2_3_31/i0[10] ) );
  AND4_X2 U8937 ( .A1(\SB3_20/Component_Function_3/NAND4_in[1] ), .A2(n2577), 
        .A3(n612), .A4(n3864), .Z(n3662) );
  NAND3_X1 U8938 ( .A1(\SB3_20/i0[8] ), .A2(\SB3_20/i3[0] ), .A3(\SB3_20/i1_5 ), .ZN(n612) );
  BUF_X2 U8939 ( .I(\SB1_1_16/buf_output[0] ), .Z(\SB2_1_11/i0[9] ) );
  INV_X1 U8940 ( .I(\SB1_1_16/buf_output[0] ), .ZN(\SB2_1_11/i3[0] ) );
  NAND2_X1 U8943 ( .A1(\SB1_1_11/i0_3 ), .A2(\SB1_1_11/i1[9] ), .ZN(
        \SB1_1_11/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U8944 ( .A1(\SB1_1_11/i1[9] ), .A2(\SB1_1_11/i1_5 ), .A3(
        \SB1_1_11/i0_4 ), .ZN(\SB1_1_11/Component_Function_4/NAND4_in[3] ) );
  BUF_X4 U8949 ( .I(\SB1_0_28/buf_output[1] ), .Z(\RI3[0][43] ) );
  AND4_X2 U8950 ( .A1(\SB1_0_13/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_13/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_0_13/Component_Function_5/NAND4_in[0] ), .A4(n4259), .Z(n3663) );
  NAND3_X1 U8953 ( .A1(\SB2_3_28/i0_3 ), .A2(\SB2_3_28/i1_7 ), .A3(
        \SB2_3_28/i0[8] ), .ZN(\SB2_3_28/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U8956 ( .A1(\SB4_17/i1_5 ), .A2(n3661), .A3(\SB4_17/i3[0] ), .ZN(
        \SB4_17/Component_Function_3/NAND4_in[3] ) );
  AND4_X2 U8959 ( .A1(\SB3_24/Component_Function_2/NAND4_in[1] ), .A2(n3888), 
        .A3(\SB3_24/Component_Function_2/NAND4_in[3] ), .A4(n3759), .Z(n3666)
         );
  XOR2_X1 U8961 ( .A1(\MC_ARK_ARC_1_2/temp6[45] ), .A2(
        \MC_ARK_ARC_1_2/temp5[45] ), .Z(n3667) );
  NAND3_X1 U8962 ( .A1(\SB2_1_22/i0_3 ), .A2(\SB2_1_22/i0[10] ), .A3(
        \SB2_1_22/i0[9] ), .ZN(n4690) );
  BUF_X2 U8964 ( .I(\MC_ARK_ARC_1_2/buf_output[78] ), .Z(\SB1_3_18/i0[9] ) );
  AND4_X2 U8965 ( .A1(\SB3_21/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_21/Component_Function_3/NAND4_in[1] ), .A3(n4217), .A4(n2005), 
        .Z(n3668) );
  BUF_X2 U8967 ( .I(\MC_ARK_ARC_1_3/buf_output[187] ), .Z(\SB3_0/i0[6] ) );
  INV_X1 U8968 ( .I(\MC_ARK_ARC_1_3/buf_output[187] ), .ZN(\SB3_0/i1_7 ) );
  BUF_X2 U8969 ( .I(\MC_ARK_ARC_1_3/buf_output[12] ), .Z(\SB3_29/i0[9] ) );
  AND4_X2 U8975 ( .A1(\SB1_3_17/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_3_17/Component_Function_3/NAND4_in[0] ), .A3(n2226), .A4(
        \SB1_3_17/Component_Function_3/NAND4_in[3] ), .Z(n3670) );
  NAND3_X1 U8976 ( .A1(\SB1_2_31/i1[9] ), .A2(\SB1_2_31/i0_3 ), .A3(
        \SB1_2_31/i0[6] ), .ZN(\SB1_2_31/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U8980 ( .A1(\MC_ARK_ARC_1_0/temp6[75] ), .A2(n1198), .Z(n3672) );
  XOR2_X1 U8981 ( .A1(\MC_ARK_ARC_1_2/temp6[177] ), .A2(n3730), .Z(n3673) );
  INV_X1 U8982 ( .I(\MC_ARK_ARC_1_3/buf_output[20] ), .ZN(\SB3_28/i1[9] ) );
  BUF_X2 U8983 ( .I(\MC_ARK_ARC_1_3/buf_output[20] ), .Z(\SB3_28/i0_0 ) );
  INV_X1 U8984 ( .I(\RI3[4][23] ), .ZN(\SB4_28/i1_5 ) );
  BUF_X2 U8985 ( .I(\SB1_2_0/buf_output[3] ), .Z(\SB2_2_30/i0[10] ) );
  INV_X1 U8986 ( .I(\SB1_2_0/buf_output[3] ), .ZN(\SB2_2_30/i0[8] ) );
  NAND3_X1 U8987 ( .A1(\SB3_17/i1[9] ), .A2(\SB3_17/i0_4 ), .A3(\SB3_17/i0_3 ), 
        .ZN(\SB3_17/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U8990 ( .A1(Key[158]), .A2(Plaintext[158]), .Z(n3675) );
  NAND4_X2 U8994 ( .A1(\SB2_2_30/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_30/Component_Function_2/NAND4_in[3] ), .A3(
        \SB2_2_30/Component_Function_2/NAND4_in[2] ), .A4(n4556), .ZN(
        \SB2_2_30/buf_output[2] ) );
  NAND4_X2 U8995 ( .A1(n3776), .A2(\SB1_3_10/Component_Function_2/NAND4_in[1] ), .A3(\SB1_3_10/Component_Function_2/NAND4_in[3] ), .A4(n4541), .ZN(n3678) );
  NAND4_X1 U8996 ( .A1(n3882), .A2(\SB2_3_7/Component_Function_2/NAND4_in[0] ), 
        .A3(n1059), .A4(n3765), .ZN(n3679) );
  CLKBUF_X4 U8997 ( .I(\SB1_3_0/buf_output[2] ), .Z(\SB2_3_29/i0_0 ) );
  INV_X1 U9001 ( .I(\SB4_29/i0_4 ), .ZN(\SB4_29/i0[7] ) );
  NAND3_X1 U9002 ( .A1(\SB3_30/i0_4 ), .A2(\SB3_30/i1[9] ), .A3(\SB3_30/i1_5 ), 
        .ZN(\SB3_30/Component_Function_4/NAND4_in[3] ) );
  XOR2_X1 U9004 ( .A1(\MC_ARK_ARC_1_1/temp6[65] ), .A2(n2807), .Z(n3682) );
  CLKBUF_X4 U9005 ( .I(\MC_ARK_ARC_1_1/buf_output[63] ), .Z(\SB1_2_21/i0[10] )
         );
  NAND3_X1 U9008 ( .A1(\RI1[1][59] ), .A2(\SB1_1_22/i0[8] ), .A3(
        \SB1_1_22/i1_7 ), .ZN(\SB1_1_22/Component_Function_1/NAND4_in[1] ) );
  INV_X4 U9009 ( .I(\RI1[1][59] ), .ZN(\SB1_1_22/i1_5 ) );
  BUF_X2 U9011 ( .I(\SB3_15/buf_output[3] ), .Z(\SB4_13/i0[10] ) );
  AND4_X2 U9015 ( .A1(\SB3_15/Component_Function_3/NAND4_in[1] ), .A2(n4423), 
        .A3(\SB3_15/Component_Function_3/NAND4_in[0] ), .A4(n4137), .Z(n3683)
         );
  NAND3_X1 U9016 ( .A1(\SB3_17/i0[9] ), .A2(\SB3_17/i0_0 ), .A3(\SB3_17/i0[8] ), .ZN(\SB3_17/Component_Function_4/NAND4_in[0] ) );
  INV_X1 U9018 ( .I(\SB1_0_25/buf_output[5] ), .ZN(\SB2_0_25/i1_5 ) );
  INV_X1 U9020 ( .I(\MC_ARK_ARC_1_3/buf_output[108] ), .ZN(\SB3_13/i3[0] ) );
  NAND2_X1 U9021 ( .A1(\SB4_29/i0_0 ), .A2(\SB4_29/i3[0] ), .ZN(
        \SB4_29/Component_Function_5/NAND4_in[0] ) );
  BUF_X2 U9026 ( .I(n300), .Z(\SB1_0_13/i0[6] ) );
  INV_X1 U9027 ( .I(n300), .ZN(\SB1_0_13/i1_7 ) );
  CLKBUF_X4 U9028 ( .I(\MC_ARK_ARC_1_0/buf_output[158] ), .Z(\SB1_1_5/i0_0 )
         );
  NAND3_X1 U9031 ( .A1(\SB1_2_0/i0_3 ), .A2(\SB1_2_0/i0[10] ), .A3(
        \SB1_2_0/i0[6] ), .ZN(\SB1_2_0/Component_Function_2/NAND4_in[1] ) );
  CLKBUF_X4 U9032 ( .I(\MC_ARK_ARC_1_0/buf_output[33] ), .Z(\SB1_1_26/i0[10] )
         );
  INV_X1 U9033 ( .I(\MC_ARK_ARC_1_3/buf_output[61] ), .ZN(\SB3_21/i1_7 ) );
  INV_X1 U9034 ( .I(n251), .ZN(\SB1_0_29/i3[0] ) );
  INV_X1 U9035 ( .I(n415), .ZN(\SB1_0_21/i1_5 ) );
  INV_X1 U9036 ( .I(n323), .ZN(\SB1_0_5/i3[0] ) );
  NAND4_X2 U9040 ( .A1(\SB1_3_10/Component_Function_3/NAND4_in[3] ), .A2(
        \SB1_3_10/Component_Function_3/NAND4_in[0] ), .A3(n2137), .A4(n4264), 
        .ZN(n3685) );
  AND4_X2 U9049 ( .A1(\SB1_2_9/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_2_9/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_2_9/Component_Function_5/NAND4_in[0] ), .A4(n3886), .Z(n3687) );
  CLKBUF_X4 U9051 ( .I(\SB1_2_6/buf_output[1] ), .Z(\SB2_2_2/i0[6] ) );
  NAND4_X2 U9054 ( .A1(\SB1_1_0/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_0/Component_Function_3/NAND4_in[1] ), .A3(n2599), .A4(n2211), 
        .ZN(n3690) );
  NAND3_X2 U9056 ( .A1(\SB2_0_17/i0[6] ), .A2(\SB2_0_17/i0[9] ), .A3(
        \RI3[0][88] ), .ZN(n2618) );
  XOR2_X1 U9057 ( .A1(\MC_ARK_ARC_1_0/temp1[128] ), .A2(n3691), .Z(
        \MC_ARK_ARC_1_0/temp5[128] ) );
  XOR2_X1 U9058 ( .A1(\RI5[0][98] ), .A2(\RI5[0][74] ), .Z(n3691) );
  XOR2_X1 U9060 ( .A1(n3692), .A2(n50), .Z(Ciphertext[168]) );
  NAND3_X1 U9062 ( .A1(\SB1_3_14/i0[6] ), .A2(\SB1_3_14/i0[8] ), .A3(
        \SB1_3_14/i0[7] ), .ZN(\SB1_3_14/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U9063 ( .A1(\SB2_3_0/i0_3 ), .A2(\SB2_3_0/i0[9] ), .A3(n5513), .ZN(
        \SB2_3_0/Component_Function_2/NAND4_in[2] ) );
  XOR2_X1 U9065 ( .A1(\RI5[3][35] ), .A2(\RI5[3][11] ), .Z(n4629) );
  NAND3_X2 U9066 ( .A1(\SB2_2_9/i0_3 ), .A2(\SB2_2_9/i0[6] ), .A3(
        \SB2_2_9/i1[9] ), .ZN(\SB2_2_9/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U9068 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[63] ), .A2(\RI5[1][87] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[117] ) );
  NAND3_X2 U9069 ( .A1(\SB2_0_11/i3[0] ), .A2(\SB2_0_11/i1_5 ), .A3(
        \SB2_0_11/i0[8] ), .ZN(n3693) );
  XOR2_X1 U9070 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[41] ), .A2(\RI5[1][5] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[131] ) );
  XOR2_X1 U9075 ( .A1(\RI5[3][61] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[97] ), 
        .Z(n3694) );
  NAND3_X2 U9077 ( .A1(\SB2_1_31/i0_3 ), .A2(\SB2_1_31/i0_4 ), .A3(
        \SB2_1_31/i1[9] ), .ZN(n3695) );
  XOR2_X1 U9078 ( .A1(\RI5[1][18] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[42] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[72] ) );
  NAND3_X2 U9088 ( .A1(\SB2_2_9/i0_3 ), .A2(\SB2_2_9/i0_4 ), .A3(
        \SB2_2_9/i1[9] ), .ZN(\SB2_2_9/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U9089 ( .A1(\RI5[3][189] ), .A2(\RI5[3][153] ), .Z(n3699) );
  NAND4_X2 U9092 ( .A1(\SB2_2_19/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_2_19/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_2_19/Component_Function_1/NAND4_in[3] ), .A4(n3701), .ZN(
        \SB2_2_19/buf_output[1] ) );
  NAND3_X2 U9093 ( .A1(\SB1_1_19/i0[10] ), .A2(\SB1_1_19/i1[9] ), .A3(
        \SB1_1_19/i1_7 ), .ZN(n3702) );
  NAND4_X2 U9094 ( .A1(\SB1_3_11/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_11/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_3_11/Component_Function_2/NAND4_in[2] ), .A4(n3949), .ZN(
        \SB1_3_11/buf_output[2] ) );
  NAND3_X2 U9095 ( .A1(\SB1_2_23/i0_4 ), .A2(\SB1_2_23/i0[9] ), .A3(
        \SB1_2_23/i0[6] ), .ZN(\SB1_2_23/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U9099 ( .A1(\SB1_1_11/i0[8] ), .A2(\SB1_1_11/i1_5 ), .A3(
        \SB1_1_11/i3[0] ), .ZN(n3704) );
  NAND4_X2 U9103 ( .A1(\SB2_3_20/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_3_20/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_3_20/Component_Function_4/NAND4_in[0] ), .A4(n3708), .ZN(
        \SB2_3_20/buf_output[4] ) );
  XOR2_X1 U9108 ( .A1(\MC_ARK_ARC_1_1/temp5[140] ), .A2(
        \MC_ARK_ARC_1_1/temp6[140] ), .Z(\MC_ARK_ARC_1_1/buf_output[140] ) );
  NAND4_X2 U9109 ( .A1(\SB2_0_12/Component_Function_2/NAND4_in[0] ), .A2(n2414), .A3(\SB2_0_12/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_0_12/Component_Function_2/NAND4_in[1] ), .ZN(
        \SB2_0_12/buf_output[2] ) );
  NAND3_X2 U9111 ( .A1(\SB2_0_27/i0[10] ), .A2(\SB2_0_27/i0_3 ), .A3(
        \SB2_0_27/i0[6] ), .ZN(\SB2_0_27/Component_Function_2/NAND4_in[1] ) );
  NAND4_X2 U9114 ( .A1(\SB1_0_30/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_0_30/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_0_30/Component_Function_1/NAND4_in[1] ), .A4(
        \SB1_0_30/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_0_30/buf_output[1] ) );
  NAND2_X2 U9116 ( .A1(\SB2_1_2/i0_3 ), .A2(\SB2_1_2/i1[9] ), .ZN(n3710) );
  XOR2_X1 U9117 ( .A1(n1618), .A2(\MC_ARK_ARC_1_2/temp1[137] ), .Z(n3711) );
  XOR2_X1 U9118 ( .A1(n3713), .A2(n3712), .Z(n4553) );
  XOR2_X1 U9119 ( .A1(\RI5[1][27] ), .A2(n70), .Z(n3712) );
  XOR2_X1 U9120 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[63] ), .A2(\RI5[1][189] ), 
        .Z(n3713) );
  NAND3_X2 U9121 ( .A1(\SB2_1_2/i0_3 ), .A2(\SB2_1_2/i1[9] ), .A3(
        \SB2_1_2/i0[6] ), .ZN(n1317) );
  XOR2_X1 U9122 ( .A1(\MC_ARK_ARC_1_3/temp2[16] ), .A2(n3714), .Z(n2548) );
  XOR2_X1 U9123 ( .A1(\RI5[3][10] ), .A2(\RI5[3][16] ), .Z(n3714) );
  XOR2_X1 U9124 ( .A1(n3715), .A2(\MC_ARK_ARC_1_3/temp5[136] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[136] ) );
  XOR2_X1 U9125 ( .A1(\MC_ARK_ARC_1_3/temp4[136] ), .A2(
        \MC_ARK_ARC_1_3/temp3[136] ), .Z(n3715) );
  INV_X2 U9126 ( .I(\SB1_1_19/buf_output[3] ), .ZN(\SB2_1_17/i0[8] ) );
  XOR2_X1 U9134 ( .A1(n1321), .A2(\MC_ARK_ARC_1_3/temp5[184] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[184] ) );
  NAND3_X2 U9139 ( .A1(\SB2_1_29/i0[7] ), .A2(\SB2_1_29/i0[6] ), .A3(
        \SB2_1_29/i0[8] ), .ZN(n4496) );
  NAND3_X1 U9142 ( .A1(\SB4_20/i0[6] ), .A2(\SB4_20/i0_4 ), .A3(\SB4_20/i0[9] ), .ZN(\SB4_20/Component_Function_5/NAND4_in[3] ) );
  NAND4_X2 U9143 ( .A1(\SB2_1_5/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_1_5/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_5/Component_Function_1/NAND4_in[2] ), .A4(n3724), .ZN(
        \SB2_1_5/buf_output[1] ) );
  XOR2_X1 U9144 ( .A1(\RI5[0][110] ), .A2(\RI5[0][74] ), .Z(n3766) );
  XOR2_X1 U9145 ( .A1(\RI5[1][27] ), .A2(\RI5[1][183] ), .Z(
        \MC_ARK_ARC_1_1/temp3[117] ) );
  NAND3_X2 U9146 ( .A1(\SB2_2_11/i0[6] ), .A2(\SB2_2_11/i0_0 ), .A3(n5826), 
        .ZN(n3725) );
  XOR2_X1 U9147 ( .A1(\RI5[3][157] ), .A2(\RI5[3][133] ), .Z(
        \MC_ARK_ARC_1_3/temp2[187] ) );
  XOR2_X1 U9150 ( .A1(\MC_ARK_ARC_1_3/temp5[35] ), .A2(n3728), .Z(
        \MC_ARK_ARC_1_3/buf_output[35] ) );
  NAND4_X2 U9152 ( .A1(\SB2_0_6/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_6/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_0_6/Component_Function_4/NAND4_in[1] ), .A4(n3729), .ZN(
        \SB2_0_6/buf_output[4] ) );
  NAND3_X2 U9156 ( .A1(\SB1_3_31/i0[6] ), .A2(\SB1_3_31/i0[9] ), .A3(
        \SB1_3_31/i1_5 ), .ZN(n3731) );
  NAND4_X2 U9157 ( .A1(\SB2_2_9/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_9/Component_Function_3/NAND4_in[2] ), .A3(n1481), .A4(n3732), 
        .ZN(\SB2_2_9/buf_output[3] ) );
  NAND3_X2 U9158 ( .A1(\SB2_2_9/i0_3 ), .A2(\SB2_2_9/i0_0 ), .A3(
        \SB2_2_9/i0_4 ), .ZN(n3732) );
  NAND3_X1 U9160 ( .A1(\SB4_29/i0[10] ), .A2(\SB4_29/i1_5 ), .A3(
        \SB4_29/i1[9] ), .ZN(\SB4_29/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U9161 ( .A1(\SB1_0_12/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_0_12/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_12/Component_Function_1/NAND4_in[3] ), .A4(n3733), .ZN(
        \RI3[0][139] ) );
  NAND4_X2 U9163 ( .A1(\SB2_2_17/Component_Function_5/NAND4_in[2] ), .A2(n4661), .A3(n4307), .A4(\SB2_2_17/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_2_17/buf_output[5] ) );
  XOR2_X1 U9166 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[141] ), .A2(\RI5[2][135] ), 
        .Z(n3735) );
  NAND3_X2 U9168 ( .A1(\SB2_2_26/i0[10] ), .A2(\SB2_2_26/i0[6] ), .A3(
        \SB2_2_26/i0_0 ), .ZN(\SB2_2_26/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U9169 ( .A1(\RI5[0][171] ), .A2(\RI5[0][147] ), .Z(
        \MC_ARK_ARC_1_0/temp2[9] ) );
  NAND4_X2 U9171 ( .A1(n3776), .A2(\SB1_3_10/Component_Function_2/NAND4_in[1] ), .A3(\SB1_3_10/Component_Function_2/NAND4_in[3] ), .A4(n4541), .ZN(
        \SB1_3_10/buf_output[2] ) );
  NAND4_X2 U9172 ( .A1(\SB1_0_5/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_0_5/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_0_5/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_0_5/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_0_5/buf_output[0] ) );
  NAND3_X1 U9174 ( .A1(\SB2_0_0/i0[9] ), .A2(\RI3[0][191] ), .A3(
        \SB2_0_0/i0[10] ), .ZN(n3736) );
  INV_X1 U9175 ( .I(\SB1_3_2/buf_output[1] ), .ZN(\SB2_3_30/i1_7 ) );
  NAND4_X2 U9176 ( .A1(\SB1_3_2/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_3_2/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_2/Component_Function_1/NAND4_in[0] ), .A4(
        \SB1_3_2/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB1_3_2/buf_output[1] ) );
  XOR2_X1 U9179 ( .A1(n4415), .A2(n3738), .Z(\MC_ARK_ARC_1_0/buf_output[22] )
         );
  XOR2_X1 U9180 ( .A1(\MC_ARK_ARC_1_0/temp4[22] ), .A2(
        \MC_ARK_ARC_1_0/temp3[22] ), .Z(n3738) );
  INV_X2 U9182 ( .I(\SB1_0_5/buf_output[3] ), .ZN(\SB2_0_3/i0[8] ) );
  XOR2_X1 U9183 ( .A1(\SB2_2_25/buf_output[3] ), .A2(\SB2_2_31/buf_output[3] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[141] ) );
  BUF_X2 U9184 ( .I(n1319), .Z(n3739) );
  NOR2_X2 U9185 ( .A1(n607), .A2(n3740), .ZN(n1319) );
  NAND3_X2 U9186 ( .A1(\SB2_0_0/i0[9] ), .A2(\RI3[0][191] ), .A3(
        \SB2_0_0/i0[8] ), .ZN(\SB2_0_0/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U9187 ( .A1(\SB2_0_0/i0[9] ), .A2(\SB2_0_0/i1_5 ), .A3(
        \SB2_0_0/i0[6] ), .ZN(\SB2_0_0/Component_Function_1/NAND4_in[2] ) );
  XOR2_X1 U9188 ( .A1(\MC_ARK_ARC_1_0/temp3[145] ), .A2(
        \MC_ARK_ARC_1_0/temp4[145] ), .Z(n3741) );
  XOR2_X1 U9189 ( .A1(n4060), .A2(\MC_ARK_ARC_1_2/temp4[128] ), .Z(n3742) );
  NAND3_X1 U9191 ( .A1(\SB2_0_1/i0_3 ), .A2(\SB2_0_1/i0[6] ), .A3(
        \SB2_0_1/i1[9] ), .ZN(\SB2_0_1/Component_Function_3/NAND4_in[0] ) );
  NAND4_X2 U9192 ( .A1(\SB1_1_24/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_1_24/Component_Function_4/NAND4_in[2] ), .A3(
        \SB1_1_24/Component_Function_4/NAND4_in[0] ), .A4(
        \SB1_1_24/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_1_24/buf_output[4] ) );
  NAND4_X2 U9195 ( .A1(\SB2_1_19/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_1_19/Component_Function_2/NAND4_in[2] ), .A3(n4381), .A4(n3743), 
        .ZN(\SB2_1_19/buf_output[2] ) );
  NAND3_X2 U9196 ( .A1(\SB1_1_22/buf_output[2] ), .A2(n578), .A3(
        \SB2_1_19/i1_5 ), .ZN(n3743) );
  NAND3_X2 U9197 ( .A1(\SB1_3_14/i0[9] ), .A2(\SB1_3_14/i0_4 ), .A3(
        \SB1_3_14/i0[6] ), .ZN(n3746) );
  XOR2_X1 U9199 ( .A1(n3747), .A2(n238), .Z(Ciphertext[82]) );
  NAND3_X1 U9202 ( .A1(\SB3_20/i0_4 ), .A2(\SB3_20/i1_5 ), .A3(\SB3_20/i1[9] ), 
        .ZN(n3748) );
  XOR2_X1 U9203 ( .A1(\RI5[2][134] ), .A2(\RI5[2][110] ), .Z(
        \MC_ARK_ARC_1_2/temp2[164] ) );
  XOR2_X1 U9204 ( .A1(\SB2_1_16/buf_output[3] ), .A2(\RI5[1][69] ), .Z(
        \MC_ARK_ARC_1_1/temp3[3] ) );
  NAND3_X2 U9205 ( .A1(\SB2_2_18/i0_4 ), .A2(\SB2_2_18/i1[9] ), .A3(n4769), 
        .ZN(n4135) );
  XOR2_X1 U9206 ( .A1(n3751), .A2(n3750), .Z(n1589) );
  XOR2_X1 U9207 ( .A1(\RI5[2][118] ), .A2(n48), .Z(n3750) );
  XOR2_X1 U9208 ( .A1(\RI5[2][154] ), .A2(\RI5[2][88] ), .Z(n3751) );
  NAND3_X2 U9209 ( .A1(\SB1_2_10/i0_0 ), .A2(\SB1_2_10/i0_4 ), .A3(
        \SB1_2_10/i1_5 ), .ZN(n611) );
  NAND4_X2 U9214 ( .A1(\SB1_3_18/Component_Function_5/NAND4_in[3] ), .A2(
        \SB1_3_18/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_3_18/Component_Function_5/NAND4_in[0] ), .A4(n3754), .ZN(
        \SB1_3_18/buf_output[5] ) );
  XOR2_X1 U9220 ( .A1(\RI5[0][137] ), .A2(\RI5[0][161] ), .Z(
        \MC_ARK_ARC_1_0/temp2[191] ) );
  NAND4_X2 U9223 ( .A1(\SB2_1_26/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_26/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_26/Component_Function_4/NAND4_in[3] ), .A4(n3757), .ZN(
        \SB2_1_26/buf_output[4] ) );
  NAND4_X2 U9225 ( .A1(\SB2_0_9/Component_Function_4/NAND4_in[3] ), .A2(n4319), 
        .A3(\SB2_0_9/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_0_9/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB2_0_9/buf_output[4] ) );
  XOR2_X1 U9227 ( .A1(n2409), .A2(n3758), .Z(\MC_ARK_ARC_1_0/buf_output[55] )
         );
  XOR2_X1 U9228 ( .A1(n4343), .A2(\MC_ARK_ARC_1_0/temp4[55] ), .Z(n3758) );
  NAND4_X2 U9229 ( .A1(\SB3_24/Component_Function_2/NAND4_in[1] ), .A2(n3888), 
        .A3(\SB3_24/Component_Function_2/NAND4_in[3] ), .A4(n3759), .ZN(
        \SB3_24/buf_output[2] ) );
  NAND3_X2 U9230 ( .A1(\SB2_1_22/i0[8] ), .A2(\SB2_1_22/i1_5 ), .A3(
        \SB2_1_22/i3[0] ), .ZN(\SB2_1_22/Component_Function_3/NAND4_in[3] ) );
  INV_X2 U9231 ( .I(\SB1_3_19/buf_output[5] ), .ZN(\SB2_3_19/i1_5 ) );
  NAND3_X1 U9232 ( .A1(\SB1_3_8/i0_0 ), .A2(\SB1_3_8/i1_7 ), .A3(
        \SB1_3_8/i3[0] ), .ZN(n3760) );
  XOR2_X1 U9235 ( .A1(\RI5[2][159] ), .A2(\RI5[2][135] ), .Z(n3762) );
  XOR2_X1 U9236 ( .A1(n3764), .A2(n3763), .Z(\MC_ARK_ARC_1_1/buf_output[132] )
         );
  XOR2_X1 U9237 ( .A1(\MC_ARK_ARC_1_1/temp1[132] ), .A2(
        \MC_ARK_ARC_1_1/temp4[132] ), .Z(n3763) );
  XOR2_X1 U9240 ( .A1(\MC_ARK_ARC_1_2/temp5[173] ), .A2(n3767), .Z(
        \MC_ARK_ARC_1_2/buf_output[173] ) );
  XOR2_X1 U9241 ( .A1(\MC_ARK_ARC_1_2/temp3[173] ), .A2(
        \MC_ARK_ARC_1_2/temp4[173] ), .Z(n3767) );
  XOR2_X1 U9242 ( .A1(n3769), .A2(n3768), .Z(n2209) );
  XOR2_X1 U9243 ( .A1(\RI5[0][95] ), .A2(\RI5[0][65] ), .Z(n3768) );
  XOR2_X1 U9244 ( .A1(\RI5[0][41] ), .A2(\RI5[0][89] ), .Z(n3769) );
  NAND3_X2 U9245 ( .A1(\SB2_1_13/i0[6] ), .A2(\SB2_1_13/i0_3 ), .A3(
        \SB2_1_13/i1[9] ), .ZN(\SB2_1_13/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U9247 ( .A1(\SB1_3_8/i0_3 ), .A2(\SB1_3_8/i0_4 ), .A3(
        \SB1_3_8/i0_0 ), .ZN(\SB1_3_8/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U9251 ( .A1(\SB2_2_2/i0_4 ), .A2(\SB2_2_2/i0_3 ), .A3(
        \SB2_2_2/i1[9] ), .ZN(\SB2_2_2/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U9252 ( .A1(\SB2_2_3/i0_3 ), .A2(\SB2_2_3/i0[10] ), .A3(
        \SB2_2_3/i0[6] ), .ZN(n1149) );
  NAND3_X2 U9253 ( .A1(\SB2_1_1/i0[10] ), .A2(\SB2_1_1/i0_0 ), .A3(
        \SB2_1_1/i0[6] ), .ZN(\SB2_1_1/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U9255 ( .A1(\SB2_0_5/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_5/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_0_5/Component_Function_2/NAND4_in[3] ), .A4(n3770), .ZN(
        \SB2_0_5/buf_output[2] ) );
  NAND3_X2 U9257 ( .A1(\SB2_2_2/i0_4 ), .A2(\SB2_2_2/i0_0 ), .A3(
        \SB2_2_2/i1_5 ), .ZN(n3771) );
  XOR2_X1 U9259 ( .A1(\RI5[1][97] ), .A2(\RI5[1][121] ), .Z(n3772) );
  NOR2_X2 U9260 ( .A1(n4227), .A2(n3773), .ZN(n1976) );
  NAND2_X1 U9261 ( .A1(\SB1_0_12/Component_Function_4/NAND4_in[0] ), .A2(n3801), .ZN(n3773) );
  NAND4_X2 U9262 ( .A1(\SB2_1_4/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_1_4/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_1_4/Component_Function_1/NAND4_in[0] ), .A4(n3774), .ZN(
        \SB2_1_4/buf_output[1] ) );
  NAND3_X1 U9263 ( .A1(\SB1_1_5/buf_output[4] ), .A2(\SB2_1_4/i1_7 ), .A3(
        \SB2_1_4/i0[8] ), .ZN(n3774) );
  NAND3_X2 U9264 ( .A1(\SB1_3_10/i0[10] ), .A2(\SB1_3_10/i1[9] ), .A3(
        \SB1_3_10/i1_5 ), .ZN(n3776) );
  XOR2_X1 U9267 ( .A1(\RI5[1][118] ), .A2(\RI5[1][154] ), .Z(n3777) );
  NAND3_X2 U9270 ( .A1(\SB2_1_26/i0_0 ), .A2(\SB2_1_26/i0_4 ), .A3(
        \SB2_1_26/i1_5 ), .ZN(n3778) );
  NAND3_X2 U9271 ( .A1(\SB2_0_14/i0[8] ), .A2(\SB2_0_14/i3[0] ), .A3(
        \SB2_0_14/i1_5 ), .ZN(\SB2_0_14/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U9272 ( .A1(n3779), .A2(\MC_ARK_ARC_1_1/buf_keyinput[51] ), .Z(
        Ciphertext[90]) );
  NAND3_X2 U9274 ( .A1(\SB2_0_26/i0[10] ), .A2(\SB2_0_26/i1[9] ), .A3(
        \SB2_0_26/i1_7 ), .ZN(\SB2_0_26/Component_Function_3/NAND4_in[2] ) );
  XOR2_X1 U9275 ( .A1(n3781), .A2(n3780), .Z(\MC_ARK_ARC_1_3/temp5[69] ) );
  XOR2_X1 U9277 ( .A1(\RI5[3][15] ), .A2(\RI5[3][69] ), .Z(n3781) );
  XOR2_X1 U9280 ( .A1(\MC_ARK_ARC_1_2/temp2[33] ), .A2(n1874), .Z(n3782) );
  NAND3_X1 U9282 ( .A1(\SB3_17/i0[6] ), .A2(\SB3_17/i0_3 ), .A3(\SB3_17/i1[9] ), .ZN(\SB3_17/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U9284 ( .A1(\RI5[1][73] ), .A2(\RI5[1][109] ), .Z(
        \MC_ARK_ARC_1_1/temp3[7] ) );
  XOR2_X1 U9288 ( .A1(\MC_ARK_ARC_1_0/temp2[176] ), .A2(n4144), .Z(n3784) );
  XOR2_X1 U9289 ( .A1(n3787), .A2(n3786), .Z(\MC_ARK_ARC_1_2/buf_output[32] )
         );
  NAND3_X1 U9292 ( .A1(\SB1_3_6/i1[9] ), .A2(\SB1_3_6/i0_4 ), .A3(
        \SB1_3_6/i1_5 ), .ZN(\SB1_3_6/Component_Function_4/NAND4_in[3] ) );
  XOR2_X1 U9293 ( .A1(n3788), .A2(\MC_ARK_ARC_1_0/temp2[163] ), .Z(
        \MC_ARK_ARC_1_0/temp5[163] ) );
  XOR2_X1 U9294 ( .A1(\RI5[0][163] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[157] ), 
        .Z(n3788) );
  XOR2_X1 U9297 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[146] ), .A2(\RI5[2][152] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[152] ) );
  NAND4_X2 U9298 ( .A1(\SB1_0_25/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_0_25/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_0_25/Component_Function_2/NAND4_in[2] ), .A4(n2629), .ZN(
        \SB1_0_25/buf_output[2] ) );
  NAND3_X2 U9300 ( .A1(\SB1_1_7/i0[9] ), .A2(\SB1_1_7/i0_3 ), .A3(
        \SB1_1_7/i0[8] ), .ZN(\SB1_1_7/Component_Function_2/NAND4_in[2] ) );
  XOR2_X1 U9302 ( .A1(\RI5[0][59] ), .A2(\RI5[0][23] ), .Z(
        \MC_ARK_ARC_1_0/temp3[149] ) );
  NAND4_X2 U9305 ( .A1(\SB1_1_9/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_1_9/Component_Function_0/NAND4_in[1] ), .A3(n3920), .A4(
        \SB1_1_9/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_1_9/buf_output[0] ) );
  NAND3_X2 U9307 ( .A1(\SB1_0_12/i0_3 ), .A2(\SB1_0_12/i0[6] ), .A3(
        \SB1_0_12/i1[9] ), .ZN(n3790) );
  NAND3_X1 U9308 ( .A1(\SB4_28/i0[9] ), .A2(\SB4_28/i0_3 ), .A3(\SB4_28/i0[8] ), .ZN(\SB4_28/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 U9311 ( .A1(n4308), .A2(\SB1_3_28/Component_Function_5/NAND4_in[1] ), .A3(n4179), .A4(\SB1_3_28/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_28/buf_output[5] ) );
  XOR2_X1 U9318 ( .A1(\MC_ARK_ARC_1_1/temp1[99] ), .A2(n3794), .Z(
        \MC_ARK_ARC_1_1/temp5[99] ) );
  XOR2_X1 U9319 ( .A1(\RI5[1][45] ), .A2(\RI5[1][69] ), .Z(n3794) );
  NAND2_X1 U9322 ( .A1(\SB4_11/i0_3 ), .A2(\SB4_11/i1[9] ), .ZN(n3796) );
  NAND4_X2 U9323 ( .A1(\SB2_0_21/Component_Function_3/NAND4_in[3] ), .A2(n1995), .A3(n4076), .A4(n3797), .ZN(\SB2_0_21/buf_output[3] ) );
  XOR2_X1 U9325 ( .A1(\MC_ARK_ARC_1_1/temp2[128] ), .A2(n3798), .Z(
        \MC_ARK_ARC_1_1/temp5[128] ) );
  XOR2_X1 U9326 ( .A1(\RI5[1][128] ), .A2(\RI5[1][122] ), .Z(n3798) );
  XOR2_X1 U9328 ( .A1(\RI5[2][64] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[58] ), 
        .Z(n3799) );
  NAND3_X2 U9331 ( .A1(\SB2_3_20/i0[10] ), .A2(\SB2_3_20/i0_0 ), .A3(
        \SB2_3_20/i0[6] ), .ZN(\SB2_3_20/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U9335 ( .A1(\SB1_3_22/i0[10] ), .A2(\SB1_3_22/i1[9] ), .A3(
        \SB1_3_22/i1_7 ), .ZN(\SB1_3_22/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U9336 ( .A1(\SB3_26/i0_3 ), .A2(\SB3_26/i0[9] ), .A3(
        \SB3_26/i0[10] ), .ZN(\SB3_26/Component_Function_4/NAND4_in[2] ) );
  XOR2_X1 U9337 ( .A1(n3803), .A2(\MC_ARK_ARC_1_3/temp5[9] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[9] ) );
  XOR2_X1 U9338 ( .A1(\MC_ARK_ARC_1_3/temp3[9] ), .A2(
        \MC_ARK_ARC_1_3/temp4[9] ), .Z(n3803) );
  INV_X1 U9339 ( .I(\SB3_10/buf_output[3] ), .ZN(\SB4_8/i0[8] ) );
  NAND4_X2 U9340 ( .A1(\SB3_10/Component_Function_3/NAND4_in[1] ), .A2(n4013), 
        .A3(n4571), .A4(n2879), .ZN(\SB3_10/buf_output[3] ) );
  NAND3_X1 U9343 ( .A1(\SB4_16/i0[6] ), .A2(\SB4_16/i0_3 ), .A3(\SB4_16/i1[9] ), .ZN(n2411) );
  NAND3_X2 U9345 ( .A1(\SB1_0_12/i0_3 ), .A2(\SB1_0_12/i0_4 ), .A3(
        \SB1_0_12/i1[9] ), .ZN(\SB1_0_12/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U9348 ( .A1(\SB1_3_7/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_3_7/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_7/Component_Function_0/NAND4_in[0] ), .A4(n3805), .ZN(
        \SB1_3_7/buf_output[0] ) );
  XOR2_X1 U9350 ( .A1(\MC_ARK_ARC_1_3/temp2[177] ), .A2(
        \MC_ARK_ARC_1_3/temp1[177] ), .Z(n3806) );
  NAND3_X2 U9353 ( .A1(\SB2_1_25/i0[6] ), .A2(\SB2_1_25/i0[7] ), .A3(
        \SB2_1_25/i0[8] ), .ZN(n2743) );
  NAND3_X1 U9354 ( .A1(\SB2_3_23/i0_0 ), .A2(\SB1_3_24/buf_output[4] ), .A3(
        \SB2_3_23/i1_5 ), .ZN(n4576) );
  XOR2_X1 U9363 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[185] ), .A2(\RI5[2][17] ), 
        .Z(n2235) );
  NAND4_X2 U9365 ( .A1(n4199), .A2(\SB1_3_28/Component_Function_4/NAND4_in[0] ), .A3(\SB1_3_28/Component_Function_4/NAND4_in[1] ), .A4(
        \SB1_3_28/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_3_28/buf_output[4] ) );
  XOR2_X1 U9366 ( .A1(\RI5[0][33] ), .A2(\RI5[0][27] ), .Z(n3810) );
  XOR2_X1 U9367 ( .A1(\SB2_2_26/buf_output[4] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[76] ), .Z(\MC_ARK_ARC_1_2/temp3[166] )
         );
  XOR2_X1 U9368 ( .A1(\MC_ARK_ARC_1_2/temp6[67] ), .A2(n3811), .Z(
        \MC_ARK_ARC_1_2/buf_output[67] ) );
  XOR2_X1 U9369 ( .A1(\MC_ARK_ARC_1_2/temp1[67] ), .A2(
        \MC_ARK_ARC_1_2/temp2[67] ), .Z(n3811) );
  XOR2_X1 U9371 ( .A1(\MC_ARK_ARC_1_1/temp1[16] ), .A2(n3813), .Z(n2784) );
  XOR2_X1 U9372 ( .A1(\RI5[1][154] ), .A2(\RI5[1][178] ), .Z(n3813) );
  XOR2_X1 U9377 ( .A1(n3816), .A2(\MC_ARK_ARC_1_2/temp6[169] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[169] ) );
  XOR2_X1 U9378 ( .A1(\MC_ARK_ARC_1_2/temp1[169] ), .A2(
        \MC_ARK_ARC_1_2/temp2[169] ), .Z(n3816) );
  XOR2_X1 U9379 ( .A1(n3818), .A2(n3817), .Z(\MC_ARK_ARC_1_1/temp5[105] ) );
  XOR2_X1 U9380 ( .A1(\RI5[1][75] ), .A2(\RI5[1][51] ), .Z(n3817) );
  XOR2_X1 U9381 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[105] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[99] ), .Z(n3818) );
  NAND3_X1 U9382 ( .A1(\SB2_1_29/i0[6] ), .A2(\SB2_1_29/i0_4 ), .A3(
        \SB1_1_2/buf_output[0] ), .ZN(
        \SB2_1_29/Component_Function_5/NAND4_in[3] ) );
  NAND2_X2 U9383 ( .A1(n2882), .A2(\SB1_1_30/Component_Function_4/NAND4_in[2] ), .ZN(\SB2_1_29/i0_4 ) );
  NAND4_X2 U9390 ( .A1(\SB1_3_27/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_27/Component_Function_2/NAND4_in[0] ), .A3(n1152), .A4(n3822), 
        .ZN(\SB1_3_27/buf_output[2] ) );
  XOR2_X1 U9393 ( .A1(\MC_ARK_ARC_1_2/temp6[170] ), .A2(n3825), .Z(
        \MC_ARK_ARC_1_2/buf_output[170] ) );
  NAND4_X2 U9395 ( .A1(\SB1_2_0/Component_Function_5/NAND4_in[1] ), .A2(n4425), 
        .A3(\SB1_2_0/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_2_0/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_2_0/buf_output[5] ) );
  NAND4_X2 U9400 ( .A1(\SB1_2_6/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_6/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_6/Component_Function_0/NAND4_in[0] ), .A4(n3829), .ZN(
        \SB1_2_6/buf_output[0] ) );
  NAND3_X1 U9401 ( .A1(\SB1_2_6/i0_0 ), .A2(\SB1_2_6/i0_3 ), .A3(
        \SB1_2_6/i0[7] ), .ZN(n3829) );
  NAND3_X2 U9402 ( .A1(\SB3_20/i0[9] ), .A2(\SB3_20/i0[8] ), .A3(\SB3_20/i0_3 ), .ZN(n3830) );
  OR2_X1 U9403 ( .A1(n4273), .A2(\SB1_1_24/buf_output[0] ), .Z(
        \SB2_1_19/Component_Function_5/NAND4_in[0] ) );
  XOR2_X1 U9404 ( .A1(n4004), .A2(n3831), .Z(n2807) );
  XOR2_X1 U9405 ( .A1(\RI5[1][59] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[35] ), 
        .Z(n3831) );
  XOR2_X1 U9406 ( .A1(\RI5[2][40] ), .A2(\RI5[2][46] ), .Z(
        \MC_ARK_ARC_1_2/temp1[46] ) );
  NAND2_X2 U9407 ( .A1(\SB1_1_22/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_1_22/Component_Function_2/NAND4_in[1] ), .ZN(n4175) );
  NAND3_X2 U9410 ( .A1(\SB2_3_24/i0[9] ), .A2(\SB2_3_24/i0_3 ), .A3(n2906), 
        .ZN(n3833) );
  XOR2_X1 U9411 ( .A1(\RI5[0][27] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[51] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[81] ) );
  XOR2_X1 U9413 ( .A1(\MC_ARK_ARC_1_0/temp2[59] ), .A2(
        \MC_ARK_ARC_1_0/temp4[59] ), .Z(n3834) );
  XOR2_X1 U9416 ( .A1(n3837), .A2(\MC_ARK_ARC_1_2/temp6[50] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[50] ) );
  NAND3_X1 U9417 ( .A1(\SB1_1_2/i0[8] ), .A2(\SB1_1_2/i0[6] ), .A3(
        \SB1_1_2/i0[7] ), .ZN(\SB1_1_2/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U9418 ( .A1(n3839), .A2(\MC_ARK_ARC_1_3/temp2[86] ), .Z(
        \MC_ARK_ARC_1_3/temp5[86] ) );
  XOR2_X1 U9419 ( .A1(\RI5[3][80] ), .A2(\RI5[3][86] ), .Z(n3839) );
  XOR2_X1 U9423 ( .A1(n4713), .A2(n3842), .Z(\MC_ARK_ARC_1_0/buf_output[39] )
         );
  XOR2_X1 U9424 ( .A1(n1315), .A2(\MC_ARK_ARC_1_0/temp4[39] ), .Z(n3842) );
  XOR2_X1 U9427 ( .A1(\MC_ARK_ARC_1_2/temp5[57] ), .A2(n3844), .Z(
        \MC_ARK_ARC_1_2/buf_output[57] ) );
  XOR2_X1 U9428 ( .A1(\MC_ARK_ARC_1_2/temp3[57] ), .A2(
        \MC_ARK_ARC_1_2/temp4[57] ), .Z(n3844) );
  XOR2_X1 U9430 ( .A1(n3845), .A2(n1195), .Z(\MC_ARK_ARC_1_0/buf_output[123] )
         );
  XOR2_X1 U9431 ( .A1(\MC_ARK_ARC_1_0/temp1[123] ), .A2(
        \MC_ARK_ARC_1_0/temp4[123] ), .Z(n3845) );
  XOR2_X1 U9434 ( .A1(\MC_ARK_ARC_1_0/temp2[21] ), .A2(n3846), .Z(
        \MC_ARK_ARC_1_0/temp5[21] ) );
  XOR2_X1 U9435 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[21] ), .A2(\RI5[0][15] ), 
        .Z(n3846) );
  NAND4_X2 U9437 ( .A1(\SB2_1_24/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_1_24/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_1_24/Component_Function_0/NAND4_in[0] ), .A4(n3847), .ZN(
        \SB2_1_24/buf_output[0] ) );
  NAND3_X1 U9439 ( .A1(\SB4_15/i0_3 ), .A2(\SB4_15/i0_4 ), .A3(\SB4_15/i0_0 ), 
        .ZN(n3848) );
  NAND4_X2 U9440 ( .A1(\SB1_3_15/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_3_15/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_3_15/Component_Function_1/NAND4_in[0] ), .A4(n3849), .ZN(
        \SB1_3_15/buf_output[1] ) );
  NAND3_X1 U9441 ( .A1(\SB2_2_13/i0[6] ), .A2(\SB2_2_13/i0[8] ), .A3(n5779), 
        .ZN(\SB2_2_13/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 U9450 ( .A1(\SB4_15/i0[10] ), .A2(\SB4_15/i0[9] ), .ZN(n3854) );
  NAND4_X2 U9451 ( .A1(\SB1_1_17/Component_Function_1/NAND4_in[3] ), .A2(n3872), .A3(\SB1_1_17/Component_Function_1/NAND4_in[0] ), .A4(n3941), .ZN(
        \SB1_1_17/buf_output[1] ) );
  XOR2_X1 U9457 ( .A1(\MC_ARK_ARC_1_0/temp2[44] ), .A2(n3856), .Z(n4274) );
  XOR2_X1 U9458 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[44] ), .A2(\RI5[0][38] ), 
        .Z(n3856) );
  NAND2_X1 U9459 ( .A1(\SB2_1_30/i0[6] ), .A2(n3857), .ZN(
        \SB2_1_30/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U9463 ( .A1(\SB1_1_12/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_1_12/Component_Function_2/NAND4_in[0] ), .A3(n1627), .A4(n3858), 
        .ZN(\SB1_1_12/buf_output[2] ) );
  NAND3_X2 U9464 ( .A1(\SB1_1_12/i0_0 ), .A2(\SB1_1_12/i0_4 ), .A3(
        \SB1_1_12/i1_5 ), .ZN(n3858) );
  XOR2_X1 U9465 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[34] ), .A2(\RI5[2][190] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[124] ) );
  NAND4_X2 U9470 ( .A1(\SB3_19/Component_Function_2/NAND4_in[0] ), .A2(n4065), 
        .A3(\SB3_19/Component_Function_2/NAND4_in[2] ), .A4(n3863), .ZN(
        \SB3_19/buf_output[2] ) );
  NAND4_X2 U9471 ( .A1(\SB3_20/Component_Function_3/NAND4_in[1] ), .A2(n2577), 
        .A3(n612), .A4(n3864), .ZN(\SB3_20/buf_output[3] ) );
  XOR2_X1 U9472 ( .A1(n3865), .A2(n4084), .Z(\MC_ARK_ARC_1_2/buf_output[73] )
         );
  XOR2_X1 U9478 ( .A1(\RI5[3][161] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[5] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[95] ) );
  XOR2_X1 U9481 ( .A1(n4385), .A2(\MC_ARK_ARC_1_2/temp1[113] ), .Z(n3991) );
  NAND3_X1 U9484 ( .A1(\SB4_0/i0_3 ), .A2(\SB3_3/buf_output[2] ), .A3(
        \SB4_0/i0[7] ), .ZN(n3868) );
  XOR2_X1 U9486 ( .A1(n3870), .A2(n3869), .Z(\MC_ARK_ARC_1_1/buf_output[33] )
         );
  XOR2_X1 U9487 ( .A1(\MC_ARK_ARC_1_1/temp1[33] ), .A2(
        \MC_ARK_ARC_1_1/temp4[33] ), .Z(n3869) );
  NAND3_X1 U9489 ( .A1(\SB4_9/i0[9] ), .A2(\SB4_9/i0[6] ), .A3(\SB4_9/i1_5 ), 
        .ZN(n3871) );
  XOR2_X1 U9493 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[65] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[59] ), .Z(n3874) );
  XOR2_X1 U9495 ( .A1(\RI5[1][119] ), .A2(n226), .Z(n3876) );
  XOR2_X1 U9496 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[89] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[155] ), .Z(n3877) );
  XOR2_X1 U9503 ( .A1(\RI5[2][147] ), .A2(\RI5[2][111] ), .Z(n3880) );
  XOR2_X1 U9506 ( .A1(\MC_ARK_ARC_1_3/temp3[43] ), .A2(
        \MC_ARK_ARC_1_3/temp4[43] ), .Z(n2033) );
  XOR2_X1 U9507 ( .A1(\RI5[2][91] ), .A2(\RI5[2][55] ), .Z(
        \MC_ARK_ARC_1_2/temp3[181] ) );
  NAND4_X2 U9509 ( .A1(\SB3_30/Component_Function_4/NAND4_in[2] ), .A2(
        \SB3_30/Component_Function_4/NAND4_in[3] ), .A3(n3891), .A4(
        \SB3_30/Component_Function_4/NAND4_in[1] ), .ZN(\SB4_29/i0_4 ) );
  XOR2_X1 U9510 ( .A1(n3884), .A2(n1924), .Z(\MC_ARK_ARC_1_0/temp5[111] ) );
  NAND3_X1 U9511 ( .A1(n5493), .A2(\SB2_1_15/i0_0 ), .A3(\SB2_1_15/i0_3 ), 
        .ZN(\SB2_1_15/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U9521 ( .A1(\SB4_25/i0[9] ), .A2(\SB4_25/i1_5 ), .A3(\SB4_25/i0[6] ), .ZN(n3887) );
  NAND4_X2 U9522 ( .A1(n795), .A2(\SB3_30/Component_Function_0/NAND4_in[3] ), 
        .A3(\SB3_30/Component_Function_0/NAND4_in[0] ), .A4(
        \SB3_30/Component_Function_0/NAND4_in[1] ), .ZN(\SB3_30/buf_output[0] ) );
  NAND4_X2 U9523 ( .A1(\SB2_3_15/Component_Function_5/NAND4_in[2] ), .A2(n4485), .A3(\SB2_3_15/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_3_15/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_3_15/buf_output[5] ) );
  XOR2_X1 U9524 ( .A1(n4456), .A2(\MC_ARK_ARC_1_1/temp6[5] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[5] ) );
  NAND4_X2 U9530 ( .A1(\SB2_2_5/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_2_5/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_2_5/Component_Function_1/NAND4_in[0] ), .A4(n3916), .ZN(
        \SB2_2_5/buf_output[1] ) );
  NAND3_X2 U9531 ( .A1(\SB2_2_12/i0[10] ), .A2(\SB2_2_12/i0_3 ), .A3(
        \SB2_2_12/i0[6] ), .ZN(n3892) );
  NAND4_X2 U9532 ( .A1(\SB2_0_28/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_0_28/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_0_28/Component_Function_0/NAND4_in[0] ), .A4(n3893), .ZN(
        \SB2_0_28/buf_output[0] ) );
  XOR2_X1 U9533 ( .A1(\RI5[0][171] ), .A2(\RI5[0][3] ), .Z(n3894) );
  XOR2_X1 U9535 ( .A1(\RI5[2][87] ), .A2(\RI5[2][111] ), .Z(n1115) );
  NAND3_X2 U9537 ( .A1(\SB2_0_14/i0[6] ), .A2(\SB2_0_14/i0_3 ), .A3(
        \RI3[0][105] ), .ZN(\SB2_0_14/Component_Function_2/NAND4_in[1] ) );
  INV_X2 U9540 ( .I(\RI3[0][20] ), .ZN(\SB2_0_28/i1[9] ) );
  NAND4_X2 U9541 ( .A1(\SB1_0_31/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_31/Component_Function_2/NAND4_in[3] ), .A3(
        \SB1_0_31/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_31/Component_Function_2/NAND4_in[1] ), .ZN(\RI3[0][20] ) );
  NAND4_X2 U9543 ( .A1(\SB1_1_25/Component_Function_1/NAND4_in[2] ), .A2(n1625), .A3(n4468), .A4(n3895), .ZN(\SB1_1_25/buf_output[1] ) );
  NAND4_X2 U9544 ( .A1(\SB3_21/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_21/Component_Function_0/NAND4_in[1] ), .A3(n2667), .A4(
        \SB3_21/Component_Function_0/NAND4_in[0] ), .ZN(\SB3_21/buf_output[0] ) );
  NAND3_X1 U9546 ( .A1(\SB3_23/i0_4 ), .A2(\SB3_23/i0[8] ), .A3(\SB3_23/i1_7 ), 
        .ZN(n3896) );
  INV_X2 U9547 ( .I(\SB1_3_28/buf_output[2] ), .ZN(\SB2_3_25/i1[9] ) );
  XOR2_X1 U9550 ( .A1(\RI5[3][20] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[176] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[110] ) );
  XOR2_X1 U9552 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[105] ), .A2(\RI5[0][111] ), 
        .Z(n1924) );
  NAND3_X2 U9553 ( .A1(\SB1_0_9/i0[10] ), .A2(\SB1_0_9/i1[9] ), .A3(
        \SB1_0_9/i1_7 ), .ZN(n3897) );
  NAND3_X2 U9558 ( .A1(\SB1_2_28/i0[10] ), .A2(\SB1_2_28/i1[9] ), .A3(
        \SB1_2_28/i1_7 ), .ZN(n3899) );
  NAND3_X2 U9561 ( .A1(\SB2_3_23/i0[9] ), .A2(\SB2_3_23/i0[8] ), .A3(
        \SB2_3_23/i0_3 ), .ZN(n3900) );
  XOR2_X1 U9562 ( .A1(\RI5[3][173] ), .A2(\RI5[3][149] ), .Z(n3901) );
  XOR2_X1 U9563 ( .A1(n1808), .A2(n3902), .Z(\MC_ARK_ARC_1_1/temp5[152] ) );
  XOR2_X1 U9564 ( .A1(\RI5[1][122] ), .A2(\RI5[1][98] ), .Z(n3902) );
  NAND3_X1 U9566 ( .A1(\SB2_0_9/i0_3 ), .A2(\SB2_0_9/i0[10] ), .A3(
        \SB2_0_9/i0[9] ), .ZN(n4319) );
  NAND3_X2 U9568 ( .A1(\SB2_0_8/i0_3 ), .A2(\SB2_0_8/i0[9] ), .A3(
        \SB2_0_8/i0[8] ), .ZN(\SB2_0_8/Component_Function_2/NAND4_in[2] ) );
  XOR2_X1 U9569 ( .A1(\MC_ARK_ARC_1_0/temp3[164] ), .A2(n3904), .Z(n3921) );
  XOR2_X1 U9570 ( .A1(\RI5[0][158] ), .A2(\RI5[0][164] ), .Z(n3904) );
  XOR2_X1 U9571 ( .A1(\RI5[1][21] ), .A2(\RI5[1][45] ), .Z(
        \MC_ARK_ARC_1_1/temp2[75] ) );
  XOR2_X1 U9572 ( .A1(\RI5[0][39] ), .A2(\RI5[0][63] ), .Z(n3905) );
  NAND3_X1 U9573 ( .A1(\SB3_1/i0_0 ), .A2(\SB3_1/i3[0] ), .A3(\SB3_1/i1_7 ), 
        .ZN(\SB3_1/Component_Function_4/NAND4_in[1] ) );
  NAND4_X2 U9575 ( .A1(n4226), .A2(n4439), .A3(
        \SB3_20/Component_Function_5/NAND4_in[1] ), .A4(n3908), .ZN(
        \SB3_20/buf_output[5] ) );
  NAND4_X2 U9576 ( .A1(\SB3_21/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_21/Component_Function_3/NAND4_in[1] ), .A3(n4217), .A4(n2005), 
        .ZN(\SB3_21/buf_output[3] ) );
  XOR2_X1 U9579 ( .A1(n3910), .A2(\MC_ARK_ARC_1_2/temp6[70] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[70] ) );
  XOR2_X1 U9580 ( .A1(\MC_ARK_ARC_1_2/temp2[70] ), .A2(
        \MC_ARK_ARC_1_2/temp1[70] ), .Z(n3910) );
  XOR2_X1 U9581 ( .A1(\MC_ARK_ARC_1_2/temp1[40] ), .A2(
        \MC_ARK_ARC_1_2/temp2[40] ), .Z(\MC_ARK_ARC_1_2/temp5[40] ) );
  XOR2_X1 U9588 ( .A1(n1634), .A2(n3914), .Z(\MC_ARK_ARC_1_0/buf_output[134] )
         );
  XOR2_X1 U9589 ( .A1(\MC_ARK_ARC_1_0/temp4[134] ), .A2(
        \MC_ARK_ARC_1_0/temp2[134] ), .Z(n3914) );
  NAND3_X2 U9592 ( .A1(\SB2_2_5/i0_4 ), .A2(\SB2_2_5/i1_7 ), .A3(
        \SB2_2_5/i0[8] ), .ZN(n3916) );
  NAND4_X2 U9595 ( .A1(\SB2_2_27/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_2_27/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_2_27/Component_Function_1/NAND4_in[2] ), .A4(n3917), .ZN(
        \SB2_2_27/buf_output[1] ) );
  XOR2_X1 U9599 ( .A1(n2011), .A2(\MC_ARK_ARC_1_0/temp1[88] ), .Z(n3919) );
  NAND3_X2 U9602 ( .A1(\SB1_2_9/i0[10] ), .A2(\SB1_2_9/i0_0 ), .A3(
        \SB1_2_9/i0[6] ), .ZN(\SB1_2_9/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U9603 ( .A1(\SB1_1_9/i0[8] ), .A2(\SB1_1_9/i1_7 ), .A3(
        \SB1_1_9/i0_4 ), .ZN(\SB1_1_9/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 U9604 ( .A1(\SB2_2_24/i0_4 ), .A2(\SB2_2_24/i1[9] ), .A3(
        \SB2_2_24/i0_3 ), .ZN(n3923) );
  XOR2_X1 U9606 ( .A1(\RI5[0][158] ), .A2(n48), .Z(n3924) );
  XOR2_X1 U9607 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[2] ), .A2(\RI5[0][128] ), 
        .Z(n3925) );
  XOR2_X1 U9608 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[105] ), .A2(\RI5[1][141] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[39] ) );
  NAND3_X1 U9609 ( .A1(\SB4_3/i0_3 ), .A2(n1371), .A3(\SB4_3/i0_4 ), .ZN(
        \SB4_3/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U9610 ( .A1(n3927), .A2(\MC_ARK_ARC_1_2/temp4[147] ), .Z(
        \MC_ARK_ARC_1_2/temp6[147] ) );
  XOR2_X1 U9611 ( .A1(\RI5[2][57] ), .A2(\RI5[2][21] ), .Z(n3927) );
  NAND3_X1 U9614 ( .A1(\SB3_9/i0[10] ), .A2(\SB3_9/i1[9] ), .A3(\SB3_9/i1_7 ), 
        .ZN(\SB3_9/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U9615 ( .A1(\SB4_7/i0[10] ), .A2(\SB4_7/i1[9] ), .A3(\SB4_7/i1_7 ), 
        .ZN(n3929) );
  INV_X2 U9616 ( .I(\SB1_1_26/buf_output[2] ), .ZN(\SB2_1_23/i1[9] ) );
  XOR2_X1 U9618 ( .A1(\RI5[1][164] ), .A2(\RI5[1][8] ), .Z(
        \MC_ARK_ARC_1_1/temp3[98] ) );
  OAI21_X2 U9620 ( .A1(n3992), .A2(\SB2_3_11/i0[9] ), .B(\SB2_3_11/i0[10] ), 
        .ZN(n3932) );
  XOR2_X1 U9623 ( .A1(n767), .A2(\MC_ARK_ARC_1_1/temp6[95] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[95] ) );
  XOR2_X1 U9625 ( .A1(\MC_ARK_ARC_1_0/temp3[17] ), .A2(
        \MC_ARK_ARC_1_0/temp4[17] ), .Z(n2051) );
  XOR2_X1 U9628 ( .A1(\MC_ARK_ARC_1_3/temp6[77] ), .A2(n3937), .Z(\RI1[4][77] ) );
  XOR2_X1 U9631 ( .A1(\MC_ARK_ARC_1_2/temp3[119] ), .A2(
        \MC_ARK_ARC_1_2/temp4[119] ), .Z(n3939) );
  NAND4_X2 U9632 ( .A1(\SB1_1_22/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_1_22/Component_Function_4/NAND4_in[1] ), .A3(n4356), .A4(n3940), 
        .ZN(\SB1_1_22/buf_output[4] ) );
  NAND3_X1 U9635 ( .A1(\SB2_2_4/i0_4 ), .A2(\SB1_2_9/buf_output[0] ), .A3(
        \SB1_2_8/buf_output[1] ), .ZN(
        \SB2_2_4/Component_Function_5/NAND4_in[3] ) );
  XOR2_X1 U9637 ( .A1(\MC_ARK_ARC_1_0/temp1[89] ), .A2(
        \MC_ARK_ARC_1_0/temp2[89] ), .Z(\MC_ARK_ARC_1_0/temp5[89] ) );
  NAND4_X2 U9643 ( .A1(\SB1_2_11/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_2_11/Component_Function_1/NAND4_in[0] ), .A3(
        \SB1_2_11/Component_Function_1/NAND4_in[1] ), .A4(
        \SB1_2_11/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_2_11/buf_output[1] ) );
  XOR2_X1 U9646 ( .A1(\MC_ARK_ARC_1_3/temp2[43] ), .A2(n1882), .Z(n3943) );
  XOR2_X1 U9648 ( .A1(\MC_ARK_ARC_1_1/temp2[158] ), .A2(
        \MC_ARK_ARC_1_1/temp1[158] ), .Z(\MC_ARK_ARC_1_1/temp5[158] ) );
  NAND4_X2 U9650 ( .A1(\SB2_3_25/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_25/Component_Function_3/NAND4_in[1] ), .A3(n4207), .A4(
        \SB2_3_25/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_3_25/buf_output[3] ) );
  XOR2_X1 U9651 ( .A1(\RI5[1][136] ), .A2(\RI5[1][172] ), .Z(
        \MC_ARK_ARC_1_1/temp3[70] ) );
  XOR2_X1 U9652 ( .A1(\RI5[0][117] ), .A2(\RI5[0][111] ), .Z(n3944) );
  NAND4_X2 U9653 ( .A1(\SB1_3_0/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_3_0/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_3_0/Component_Function_4/NAND4_in[3] ), .A4(n3945), .ZN(
        \SB1_3_0/buf_output[4] ) );
  NAND4_X2 U9655 ( .A1(n1344), .A2(\SB2_1_10/Component_Function_4/NAND4_in[3] ), .A3(n1346), .A4(n3946), .ZN(\SB2_1_10/buf_output[4] ) );
  NAND3_X2 U9657 ( .A1(\SB2_2_27/i0_0 ), .A2(\SB2_2_27/i0_3 ), .A3(
        \SB1_2_28/buf_output[4] ), .ZN(n3947) );
  NAND3_X2 U9658 ( .A1(\SB2_0_14/i0_3 ), .A2(\RI3[0][104] ), .A3(\RI3[0][106] ), .ZN(\SB2_0_14/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U9659 ( .A1(\SB4_18/i0[10] ), .A2(\SB4_18/i1_5 ), .A3(
        \SB4_18/i1[9] ), .ZN(n3948) );
  NAND3_X2 U9660 ( .A1(\SB1_3_11/i0_4 ), .A2(\SB1_3_11/i0[8] ), .A3(
        \SB1_3_11/i1_7 ), .ZN(n775) );
  XOR2_X1 U9667 ( .A1(\RI5[0][137] ), .A2(\RI5[0][101] ), .Z(
        \MC_ARK_ARC_1_0/temp3[35] ) );
  XOR2_X1 U9668 ( .A1(\MC_ARK_ARC_1_1/temp5[154] ), .A2(n3952), .Z(
        \MC_ARK_ARC_1_1/buf_output[154] ) );
  XOR2_X1 U9669 ( .A1(\MC_ARK_ARC_1_1/temp3[154] ), .A2(
        \MC_ARK_ARC_1_1/temp4[154] ), .Z(n3952) );
  NAND4_X2 U9670 ( .A1(\SB2_1_4/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_4/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_1_4/Component_Function_3/NAND4_in[3] ), .A4(n790), .ZN(
        \SB2_1_4/buf_output[3] ) );
  NAND3_X2 U9671 ( .A1(\SB2_3_22/i0_4 ), .A2(\SB2_3_22/i0_3 ), .A3(
        \SB2_3_22/i1[9] ), .ZN(n3954) );
  NAND3_X1 U9672 ( .A1(\SB1_2_11/i0_3 ), .A2(\SB1_2_11/i0[9] ), .A3(
        \SB1_2_11/i0[8] ), .ZN(\SB1_2_11/Component_Function_2/NAND4_in[2] ) );
  XOR2_X1 U9675 ( .A1(\RI5[1][125] ), .A2(n533), .Z(n3955) );
  NAND3_X2 U9677 ( .A1(\SB1_1_7/i0_3 ), .A2(\SB1_1_7/i1[9] ), .A3(
        \SB1_1_7/i0[6] ), .ZN(\SB1_1_7/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U9679 ( .A1(\SB1_1_16/i0[10] ), .A2(\SB1_1_16/i0_0 ), .A3(
        \SB1_1_16/i0[6] ), .ZN(\SB1_1_16/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U9680 ( .A1(\SB1_1_2/i0[9] ), .A2(\SB1_1_2/i0_3 ), .A3(
        \MC_ARK_ARC_1_0/buf_output[177] ), .ZN(
        \SB1_1_2/Component_Function_4/NAND4_in[2] ) );
  XOR2_X1 U9681 ( .A1(\RI5[2][101] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[95] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[101] ) );
  NAND4_X2 U9682 ( .A1(\SB1_1_8/Component_Function_2/NAND4_in[3] ), .A2(n911), 
        .A3(\SB1_1_8/Component_Function_2/NAND4_in[2] ), .A4(n910), .ZN(
        \SB1_1_8/buf_output[2] ) );
  XOR2_X1 U9683 ( .A1(\RI5[0][149] ), .A2(\RI5[0][125] ), .Z(
        \MC_ARK_ARC_1_0/temp2[179] ) );
  NAND3_X2 U9684 ( .A1(\SB2_1_13/i1_5 ), .A2(\SB2_1_13/i0_0 ), .A3(
        \SB2_1_13/i0_4 ), .ZN(n4493) );
  NAND4_X2 U9686 ( .A1(\SB1_0_27/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_27/Component_Function_2/NAND4_in[3] ), .A3(
        \SB1_0_27/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_0_27/Component_Function_2/NAND4_in[1] ), .ZN(\RI3[0][44] ) );
  NAND3_X2 U9687 ( .A1(\SB2_1_12/i0[10] ), .A2(\SB2_1_12/i0[6] ), .A3(
        \SB2_1_12/i0_0 ), .ZN(\SB2_1_12/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U9691 ( .A1(n2172), .A2(\MC_ARK_ARC_1_3/temp1[131] ), .Z(
        \MC_ARK_ARC_1_3/temp5[131] ) );
  XOR2_X1 U9692 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[185] ), .A2(\RI5[2][161] ), 
        .Z(n3961) );
  NAND4_X2 U9693 ( .A1(\SB1_1_26/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_1_26/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_1_26/Component_Function_1/NAND4_in[0] ), .A4(n3962), .ZN(
        \SB1_1_26/buf_output[1] ) );
  NAND3_X1 U9694 ( .A1(\SB1_1_26/i0[8] ), .A2(\SB1_1_26/i0_4 ), .A3(
        \SB1_1_26/i1_7 ), .ZN(n3962) );
  NAND3_X1 U9700 ( .A1(\SB3_0/i0[6] ), .A2(\SB3_0/i0[10] ), .A3(\SB3_0/i0_3 ), 
        .ZN(n3968) );
  NAND4_X2 U9701 ( .A1(\SB1_1_12/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_1_12/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_12/Component_Function_0/NAND4_in[0] ), .A4(n3969), .ZN(
        \SB1_1_12/buf_output[0] ) );
  NAND3_X1 U9702 ( .A1(\SB1_1_12/i0_0 ), .A2(\SB1_1_12/i0_3 ), .A3(
        \SB1_1_12/i0[7] ), .ZN(n3969) );
  XOR2_X1 U9703 ( .A1(n3970), .A2(\MC_ARK_ARC_1_3/temp6[187] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[187] ) );
  XOR2_X1 U9704 ( .A1(\MC_ARK_ARC_1_3/temp2[187] ), .A2(
        \MC_ARK_ARC_1_3/temp1[187] ), .Z(n3970) );
  XOR2_X1 U9706 ( .A1(n2453), .A2(n2452), .Z(\MC_ARK_ARC_1_0/buf_output[121] )
         );
  NAND3_X1 U9707 ( .A1(\SB1_3_7/i0[10] ), .A2(\SB1_3_7/i1_7 ), .A3(
        \SB1_3_7/i1[9] ), .ZN(n3972) );
  XOR2_X1 U9708 ( .A1(\SB2_0_2/buf_output[3] ), .A2(\SB2_0_30/buf_output[3] ), 
        .Z(n3977) );
  XOR2_X1 U9709 ( .A1(n1375), .A2(\MC_ARK_ARC_1_0/buf_datainput[150] ), .Z(
        \MC_ARK_ARC_1_0/temp3[48] ) );
  XOR2_X1 U9711 ( .A1(n4073), .A2(n3974), .Z(\MC_ARK_ARC_1_2/buf_output[64] )
         );
  INV_X1 U9713 ( .I(\SB1_2_16/buf_output[1] ), .ZN(\SB2_2_12/i1_7 ) );
  NAND4_X2 U9715 ( .A1(n3975), .A2(\SB2_3_4/Component_Function_5/NAND4_in[2] ), 
        .A3(\SB2_3_4/Component_Function_5/NAND4_in[0] ), .A4(
        \SB2_3_4/Component_Function_5/NAND4_in[1] ), .ZN(
        \SB2_3_4/buf_output[5] ) );
  NAND3_X2 U9716 ( .A1(\SB2_3_4/i0[6] ), .A2(\SB2_3_4/i0_4 ), .A3(
        \SB2_3_4/i0[9] ), .ZN(n3975) );
  XOR2_X1 U9718 ( .A1(\MC_ARK_ARC_1_3/temp3[50] ), .A2(
        \MC_ARK_ARC_1_3/temp4[50] ), .Z(n2809) );
  NAND3_X1 U9719 ( .A1(\SB3_24/i0[6] ), .A2(\SB3_24/i0_4 ), .A3(\SB3_24/i0[9] ), .ZN(\SB3_24/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 U9721 ( .A1(\SB1_3_17/i0_4 ), .A2(\SB1_3_17/i1[9] ), .A3(
        \SB1_3_17/i0_3 ), .ZN(n3976) );
  XOR2_X1 U9722 ( .A1(n3978), .A2(n3977), .Z(n4656) );
  XOR2_X1 U9725 ( .A1(n3980), .A2(n2051), .Z(\MC_ARK_ARC_1_0/buf_output[17] )
         );
  XOR2_X1 U9726 ( .A1(\MC_ARK_ARC_1_0/temp2[17] ), .A2(
        \MC_ARK_ARC_1_0/temp1[17] ), .Z(n3980) );
  NAND4_X2 U9729 ( .A1(\SB1_3_1/Component_Function_5/NAND4_in[1] ), .A2(n4120), 
        .A3(n1106), .A4(\SB1_3_1/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_1/buf_output[5] ) );
  INV_X2 U9730 ( .I(\RI3[0][152] ), .ZN(\SB2_0_6/i1[9] ) );
  NAND4_X2 U9731 ( .A1(\SB1_0_9/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_9/Component_Function_2/NAND4_in[3] ), .A3(n4028), .A4(
        \SB1_0_9/Component_Function_2/NAND4_in[2] ), .ZN(\RI3[0][152] ) );
  XOR2_X1 U9732 ( .A1(\MC_ARK_ARC_1_3/temp5[47] ), .A2(
        \MC_ARK_ARC_1_3/temp6[47] ), .Z(\MC_ARK_ARC_1_3/buf_output[47] ) );
  XOR2_X1 U9733 ( .A1(\MC_ARK_ARC_1_1/temp3[186] ), .A2(
        \MC_ARK_ARC_1_1/temp4[186] ), .Z(n1325) );
  NAND4_X2 U9734 ( .A1(\SB2_0_12/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_0_12/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_0_12/Component_Function_4/NAND4_in[3] ), .A4(
        \SB2_0_12/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB2_0_12/buf_output[4] ) );
  NAND2_X1 U9741 ( .A1(\SB1_3_1/Component_Function_4/NAND4_in[0] ), .A2(n3984), 
        .ZN(n739) );
  XOR2_X1 U9745 ( .A1(\RI5[1][96] ), .A2(\RI5[1][120] ), .Z(
        \MC_ARK_ARC_1_1/temp2[150] ) );
  XOR2_X1 U9747 ( .A1(n3988), .A2(n224), .Z(Ciphertext[107]) );
  NAND3_X1 U9753 ( .A1(\SB2_2_27/i0_0 ), .A2(\SB2_2_27/i3[0] ), .A3(
        \SB2_2_27/i1_7 ), .ZN(\SB2_2_27/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U9754 ( .A1(\RI5[1][2] ), .A2(\RI5[1][8] ), .Z(n3990) );
  NAND3_X1 U9760 ( .A1(\SB1_3_23/i0_3 ), .A2(\SB1_3_23/i0[8] ), .A3(
        \SB1_3_23/i1_7 ), .ZN(\SB1_3_23/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U9762 ( .A1(\RI5[0][18] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[42] ), 
        .Z(n3996) );
  NAND2_X1 U9763 ( .A1(\SB3_16/i0[9] ), .A2(\SB3_16/i0[10] ), .ZN(
        \SB3_16/Component_Function_0/NAND4_in[0] ) );
  XOR2_X1 U9764 ( .A1(n3997), .A2(n4536), .Z(\MC_ARK_ARC_1_3/buf_output[66] )
         );
  XOR2_X1 U9765 ( .A1(\MC_ARK_ARC_1_3/temp4[66] ), .A2(
        \MC_ARK_ARC_1_3/temp3[66] ), .Z(n3997) );
  AND2_X1 U9766 ( .A1(\SB2_3_19/Component_Function_0/NAND4_in[1] ), .A2(n2112), 
        .Z(n2285) );
  XOR2_X1 U9767 ( .A1(n3998), .A2(\MC_ARK_ARC_1_3/temp4[58] ), .Z(
        \MC_ARK_ARC_1_3/temp6[58] ) );
  XOR2_X1 U9768 ( .A1(\RI5[3][160] ), .A2(\RI5[3][124] ), .Z(n3998) );
  NAND3_X1 U9770 ( .A1(\SB2_3_12/i0[10] ), .A2(\SB2_3_12/i0_3 ), .A3(n1603), 
        .ZN(n4000) );
  XOR2_X1 U9772 ( .A1(\RI5[3][181] ), .A2(\RI5[3][13] ), .Z(
        \MC_ARK_ARC_1_3/temp2[43] ) );
  NAND4_X2 U9773 ( .A1(\SB1_1_20/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_1_20/Component_Function_0/NAND4_in[1] ), .A3(n1110), .A4(n4001), 
        .ZN(\SB1_1_20/buf_output[0] ) );
  XOR2_X1 U9775 ( .A1(n3650), .A2(\RI5[1][65] ), .Z(n4004) );
  INV_X1 U9778 ( .I(\SB3_17/buf_output[0] ), .ZN(\SB4_12/i3[0] ) );
  NAND4_X2 U9779 ( .A1(\SB3_17/Component_Function_0/NAND4_in[3] ), .A2(
        \SB3_17/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_17/Component_Function_0/NAND4_in[2] ), .A4(
        \SB3_17/Component_Function_0/NAND4_in[0] ), .ZN(\SB3_17/buf_output[0] ) );
  XOR2_X1 U9780 ( .A1(n4006), .A2(n144), .Z(Ciphertext[169]) );
  NAND3_X1 U9785 ( .A1(\SB4_13/i0_3 ), .A2(\SB4_13/i0_4 ), .A3(\SB4_13/i1[9] ), 
        .ZN(\SB4_13/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U9786 ( .A1(\SB2_0_25/i0_3 ), .A2(\SB1_0_29/buf_output[1] ), .A3(
        \RI3[0][39] ), .ZN(n4008) );
  NAND3_X2 U9787 ( .A1(\SB1_3_28/i0[6] ), .A2(\SB1_3_28/i0_4 ), .A3(
        \SB1_3_28/i0[9] ), .ZN(n4179) );
  NAND4_X2 U9788 ( .A1(\SB2_2_18/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_18/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_2_18/Component_Function_1/NAND4_in[1] ), .A4(n4009), .ZN(
        \SB2_2_18/buf_output[1] ) );
  XOR2_X1 U9790 ( .A1(\MC_ARK_ARC_1_2/temp5[138] ), .A2(n4010), .Z(
        \MC_ARK_ARC_1_2/buf_output[138] ) );
  XOR2_X1 U9791 ( .A1(\MC_ARK_ARC_1_2/temp3[138] ), .A2(
        \MC_ARK_ARC_1_2/temp4[138] ), .Z(n4010) );
  INV_X4 U9792 ( .I(\SB2_2_4/i0[7] ), .ZN(\SB2_2_4/i0_4 ) );
  NOR2_X2 U9794 ( .A1(n4012), .A2(n4011), .ZN(\SB2_2_4/i0[7] ) );
  XOR2_X1 U9797 ( .A1(\MC_ARK_ARC_1_1/temp3[158] ), .A2(
        \MC_ARK_ARC_1_1/temp4[158] ), .Z(\MC_ARK_ARC_1_1/temp6[158] ) );
  NAND4_X2 U9799 ( .A1(n4230), .A2(\SB3_16/Component_Function_0/NAND4_in[3] ), 
        .A3(\SB3_16/Component_Function_0/NAND4_in[0] ), .A4(
        \SB3_16/Component_Function_0/NAND4_in[1] ), .ZN(\SB3_16/buf_output[0] ) );
  NAND3_X1 U9800 ( .A1(\SB3_10/i0[10] ), .A2(\SB3_10/i1[9] ), .A3(
        \SB3_10/i1_7 ), .ZN(n4013) );
  NAND4_X2 U9803 ( .A1(\SB1_0_9/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_9/Component_Function_5/NAND4_in[3] ), .A3(n1812), .A4(
        \SB1_0_9/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_0_9/buf_output[5] ) );
  XOR2_X1 U9804 ( .A1(\RI5[2][77] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[53] ), 
        .Z(n1232) );
  XOR2_X1 U9805 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[116] ), .A2(\RI5[3][140] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[170] ) );
  NAND4_X2 U9808 ( .A1(\SB2_1_8/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_1_8/Component_Function_0/NAND4_in[1] ), .A3(n4529), .A4(n4014), 
        .ZN(\SB2_1_8/buf_output[0] ) );
  NAND3_X1 U9810 ( .A1(\SB1_0_4/i0_4 ), .A2(\SB1_0_4/i0[9] ), .A3(
        \SB1_0_4/i0[6] ), .ZN(\SB1_0_4/Component_Function_5/NAND4_in[3] ) );
  XOR2_X1 U9811 ( .A1(\RI5[3][160] ), .A2(n132), .Z(
        \MC_ARK_ARC_1_3/temp4[124] ) );
  AND2_X1 U9812 ( .A1(\SB2_3_6/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_3_6/Component_Function_4/NAND4_in[3] ), .Z(n4017) );
  NAND3_X1 U9814 ( .A1(\SB4_8/i0_0 ), .A2(\SB4_8/i0[9] ), .A3(\SB4_8/i0[8] ), 
        .ZN(n4018) );
  INV_X2 U9820 ( .I(\SB1_1_21/buf_output[3] ), .ZN(\SB2_1_19/i0[8] ) );
  NAND4_X2 U9822 ( .A1(\SB2_3_17/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_3_17/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_3_17/Component_Function_4/NAND4_in[3] ), .A4(n4021), .ZN(
        \SB2_3_17/buf_output[4] ) );
  XOR2_X1 U9823 ( .A1(\RI5[2][120] ), .A2(\RI5[2][144] ), .Z(
        \MC_ARK_ARC_1_2/temp2[174] ) );
  NAND4_X2 U9827 ( .A1(\SB1_1_5/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_1_5/Component_Function_1/NAND4_in[0] ), .A3(
        \SB1_1_5/Component_Function_1/NAND4_in[3] ), .A4(
        \SB1_1_5/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB1_1_5/buf_output[1] ) );
  NAND3_X1 U9828 ( .A1(\SB1_1_5/i0_0 ), .A2(\SB1_1_5/i0[8] ), .A3(
        \SB1_1_5/i0[9] ), .ZN(n4023) );
  NAND4_X2 U9829 ( .A1(\SB2_2_12/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_2_12/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_2_12/Component_Function_0/NAND4_in[1] ), .A4(
        \SB2_2_12/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_2_12/buf_output[0] ) );
  NAND3_X1 U9830 ( .A1(\SB1_2_16/i1_7 ), .A2(\SB1_2_16/i0_4 ), .A3(
        \SB1_2_16/i0[8] ), .ZN(n4024) );
  NAND4_X2 U9834 ( .A1(\SB1_2_21/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_21/Component_Function_0/NAND4_in[0] ), .A3(
        \SB1_2_21/Component_Function_0/NAND4_in[1] ), .A4(n4026), .ZN(
        \SB1_2_21/buf_output[0] ) );
  NAND4_X2 U9835 ( .A1(\SB1_1_27/Component_Function_5/NAND4_in[1] ), .A2(n1745), .A3(n4087), .A4(\SB1_1_27/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_27/buf_output[5] ) );
  XOR2_X1 U9837 ( .A1(\MC_ARK_ARC_1_3/temp1[67] ), .A2(
        \MC_ARK_ARC_1_3/temp2[67] ), .Z(n4027) );
  XOR2_X1 U9839 ( .A1(\MC_ARK_ARC_1_3/temp6[0] ), .A2(n4029), .Z(
        \MC_ARK_ARC_1_3/buf_output[0] ) );
  XOR2_X1 U9840 ( .A1(\MC_ARK_ARC_1_3/temp2[0] ), .A2(
        \MC_ARK_ARC_1_3/temp1[0] ), .Z(n4029) );
  INV_X1 U9841 ( .I(\SB3_5/buf_output[5] ), .ZN(\SB4_5/i1_5 ) );
  INV_X2 U9847 ( .I(\SB1_0_10/buf_output[3] ), .ZN(\SB2_0_8/i0[8] ) );
  NAND4_X2 U9848 ( .A1(\SB1_0_10/Component_Function_3/NAND4_in[2] ), .A2(
        \SB1_0_10/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_0_10/Component_Function_3/NAND4_in[1] ), .A4(
        \SB1_0_10/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_0_10/buf_output[3] ) );
  NAND4_X2 U9849 ( .A1(\SB2_0_9/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_9/Component_Function_3/NAND4_in[3] ), .A3(
        \SB2_0_9/Component_Function_3/NAND4_in[1] ), .A4(n4032), .ZN(
        \SB2_0_9/buf_output[3] ) );
  NAND3_X2 U9850 ( .A1(\SB2_0_9/i1[9] ), .A2(\SB2_0_9/i0[10] ), .A3(
        \SB2_0_9/i1_7 ), .ZN(n4032) );
  XOR2_X1 U9852 ( .A1(n1537), .A2(\MC_ARK_ARC_1_2/temp2[122] ), .Z(n4033) );
  INV_X2 U9856 ( .I(n4034), .ZN(\RI1[2][59] ) );
  XNOR2_X1 U9857 ( .A1(\MC_ARK_ARC_1_1/temp6[59] ), .A2(n4133), .ZN(n4034) );
  INV_X2 U9858 ( .I(\RI3[0][2] ), .ZN(\SB2_0_31/i1[9] ) );
  NAND4_X2 U9860 ( .A1(\SB1_3_13/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_13/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_13/Component_Function_4/NAND4_in[3] ), .A4(n4035), .ZN(
        \SB1_3_13/buf_output[4] ) );
  XOR2_X1 U9863 ( .A1(\MC_ARK_ARC_1_3/temp3[104] ), .A2(
        \MC_ARK_ARC_1_3/temp4[104] ), .Z(\MC_ARK_ARC_1_3/temp6[104] ) );
  NAND3_X2 U9864 ( .A1(\SB2_2_18/i0_4 ), .A2(\SB2_2_18/i0[6] ), .A3(
        \SB2_2_18/i0[9] ), .ZN(n4039) );
  XOR2_X1 U9865 ( .A1(\MC_ARK_ARC_1_0/temp2[106] ), .A2(
        \MC_ARK_ARC_1_0/temp1[106] ), .Z(\MC_ARK_ARC_1_0/temp5[106] ) );
  XOR2_X1 U9868 ( .A1(\MC_ARK_ARC_1_3/temp3[85] ), .A2(
        \MC_ARK_ARC_1_3/temp4[85] ), .Z(n4041) );
  XOR2_X1 U9871 ( .A1(n1058), .A2(\MC_ARK_ARC_1_2/temp4[37] ), .Z(n2813) );
  NAND3_X1 U9872 ( .A1(\SB3_24/i0[6] ), .A2(\SB3_24/i0_3 ), .A3(
        \SB3_24/i0[10] ), .ZN(\SB3_24/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U9873 ( .A1(\SB3_24/i0[6] ), .A2(\SB3_24/i0[8] ), .A3(
        \SB3_24/i0[7] ), .ZN(\SB3_24/Component_Function_0/NAND4_in[1] ) );
  INV_X2 U9874 ( .I(\SB1_3_25/buf_output[3] ), .ZN(\SB2_3_23/i0[8] ) );
  NAND4_X2 U9875 ( .A1(\SB1_3_25/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_25/Component_Function_3/NAND4_in[1] ), .A3(n1163), .A4(
        \SB1_3_25/Component_Function_3/NAND4_in[2] ), .ZN(
        \SB1_3_25/buf_output[3] ) );
  XOR2_X1 U9878 ( .A1(n681), .A2(n2597), .Z(\MC_ARK_ARC_1_3/buf_output[109] )
         );
  XOR2_X1 U9880 ( .A1(\RI5[3][107] ), .A2(\RI5[3][143] ), .Z(n4348) );
  XOR2_X1 U9882 ( .A1(\MC_ARK_ARC_1_3/temp5[7] ), .A2(n4044), .Z(
        \MC_ARK_ARC_1_3/buf_output[7] ) );
  XOR2_X1 U9883 ( .A1(\MC_ARK_ARC_1_3/temp3[7] ), .A2(
        \MC_ARK_ARC_1_3/temp4[7] ), .Z(n4044) );
  NAND4_X2 U9884 ( .A1(\SB2_2_30/Component_Function_4/NAND4_in[3] ), .A2(n1694), .A3(\SB2_2_30/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_2_30/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB2_2_30/buf_output[4] ) );
  NAND4_X2 U9885 ( .A1(\SB2_3_6/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_3_6/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_3_6/Component_Function_1/NAND4_in[0] ), .A4(n4083), .ZN(
        \SB2_3_6/buf_output[1] ) );
  NAND3_X2 U9887 ( .A1(\SB1_2_15/i3[0] ), .A2(\SB1_2_15/i0[8] ), .A3(
        \SB1_2_15/i1_5 ), .ZN(n4085) );
  INV_X2 U9888 ( .I(\SB1_1_14/buf_output[2] ), .ZN(\SB2_1_11/i1[9] ) );
  XOR2_X1 U9894 ( .A1(\RI5[2][48] ), .A2(\RI5[2][84] ), .Z(
        \MC_ARK_ARC_1_2/temp3[174] ) );
  INV_X2 U9895 ( .I(\SB1_1_2/buf_output[3] ), .ZN(\SB2_1_0/i0[8] ) );
  XOR2_X1 U9897 ( .A1(n4047), .A2(n4048), .Z(\MC_ARK_ARC_1_2/buf_output[22] )
         );
  XOR2_X1 U9898 ( .A1(\MC_ARK_ARC_1_2/temp1[22] ), .A2(
        \MC_ARK_ARC_1_2/temp2[22] ), .Z(n4047) );
  XOR2_X1 U9899 ( .A1(\MC_ARK_ARC_1_2/temp4[22] ), .A2(
        \MC_ARK_ARC_1_2/temp3[22] ), .Z(n4048) );
  XOR2_X1 U9900 ( .A1(\MC_ARK_ARC_1_3/temp5[56] ), .A2(
        \MC_ARK_ARC_1_3/temp6[56] ), .Z(\MC_ARK_ARC_1_3/buf_output[56] ) );
  NAND3_X1 U9901 ( .A1(\SB3_5/buf_output[3] ), .A2(\SB4_3/i1_7 ), .A3(n1371), 
        .ZN(\SB4_3/Component_Function_3/NAND4_in[2] ) );
  NAND4_X2 U9903 ( .A1(\SB1_3_0/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_3_0/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_3_0/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_0/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_3_0/buf_output[1] ) );
  NAND3_X1 U9904 ( .A1(\SB4_9/i0[6] ), .A2(\SB4_9/i0_3 ), .A3(\SB4_9/i1[9] ), 
        .ZN(n4051) );
  NAND3_X1 U9908 ( .A1(\SB3_13/i0[6] ), .A2(\SB3_13/i0[9] ), .A3(\SB3_13/i1_5 ), .ZN(\SB3_13/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U9909 ( .A1(\SB3_13/i0[6] ), .A2(\SB3_13/i0[8] ), .A3(
        \SB3_13/i0[7] ), .ZN(\SB3_13/Component_Function_0/NAND4_in[1] ) );
  NAND4_X2 U9910 ( .A1(\SB3_8/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_8/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_8/Component_Function_0/NAND4_in[0] ), .A4(n4052), .ZN(
        \SB3_8/buf_output[0] ) );
  XOR2_X1 U9911 ( .A1(n4055), .A2(n4054), .Z(n4204) );
  XOR2_X1 U9913 ( .A1(\RI5[3][39] ), .A2(\RI5[3][87] ), .Z(n4055) );
  NAND3_X2 U9915 ( .A1(\SB2_0_3/i0_3 ), .A2(\RI3[0][172] ), .A3(
        \SB2_0_3/i1[9] ), .ZN(n4056) );
  NAND4_X2 U9916 ( .A1(\SB3_18/Component_Function_1/NAND4_in[1] ), .A2(
        \SB3_18/Component_Function_1/NAND4_in[3] ), .A3(
        \SB3_18/Component_Function_1/NAND4_in[0] ), .A4(n4057), .ZN(
        \SB3_18/buf_output[1] ) );
  NAND3_X1 U9917 ( .A1(\SB3_18/i0[6] ), .A2(\SB3_18/i0_3 ), .A3(
        \SB3_18/i0[10] ), .ZN(n4058) );
  XOR2_X1 U9919 ( .A1(\RI5[3][121] ), .A2(\RI5[3][127] ), .Z(
        \MC_ARK_ARC_1_3/temp1[127] ) );
  NAND3_X2 U9920 ( .A1(\SB2_1_24/i0_3 ), .A2(\SB2_1_24/i0[9] ), .A3(
        \SB2_1_24/i0[8] ), .ZN(\SB2_1_24/Component_Function_2/NAND4_in[2] ) );
  INV_X4 U9921 ( .I(n4231), .ZN(\RI3[0][39] ) );
  XOR2_X1 U9923 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[40] ), .A2(\RI5[3][64] ), 
        .Z(n4059) );
  NAND3_X2 U9924 ( .A1(\SB2_3_29/i0_3 ), .A2(\RI3[3][16] ), .A3(
        \SB2_3_29/i1[9] ), .ZN(\SB2_3_29/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U9926 ( .A1(\SB1_1_15/i0_3 ), .A2(\SB1_1_15/i0[8] ), .A3(
        \SB1_1_15/i1_7 ), .ZN(\SB1_1_15/Component_Function_1/NAND4_in[1] ) );
  NAND4_X2 U9927 ( .A1(\SB2_1_15/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_1_15/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_1_15/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_15/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_1_15/buf_output[1] ) );
  NAND3_X2 U9928 ( .A1(\SB2_1_12/i0[10] ), .A2(\SB2_1_12/i1[9] ), .A3(
        \SB2_1_12/i1_7 ), .ZN(\SB2_1_12/Component_Function_3/NAND4_in[2] ) );
  INV_X2 U9929 ( .I(\SB1_1_28/buf_output[3] ), .ZN(\SB2_1_26/i0[8] ) );
  XOR2_X1 U9931 ( .A1(\RI5[1][145] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[169] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[7] ) );
  XOR2_X1 U9932 ( .A1(n4061), .A2(\MC_ARK_ARC_1_0/temp6[97] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[97] ) );
  XOR2_X1 U9933 ( .A1(\MC_ARK_ARC_1_0/temp2[97] ), .A2(
        \MC_ARK_ARC_1_0/temp1[97] ), .Z(n4061) );
  INV_X2 U9935 ( .I(\SB1_1_15/buf_output[5] ), .ZN(\SB2_1_15/i1_5 ) );
  XOR2_X1 U9937 ( .A1(\RI5[3][77] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[71] ), 
        .Z(n2292) );
  XOR2_X1 U9939 ( .A1(\RI5[2][18] ), .A2(\RI5[2][54] ), .Z(n4063) );
  NAND3_X1 U9941 ( .A1(\SB4_14/i0[9] ), .A2(\SB4_14/i0[6] ), .A3(\SB4_14/i0_4 ), .ZN(n2572) );
  NAND4_X2 U9942 ( .A1(\SB1_2_19/Component_Function_3/NAND4_in[0] ), .A2(n2230), .A3(\SB1_2_19/Component_Function_3/NAND4_in[3] ), .A4(
        \SB1_2_19/Component_Function_3/NAND4_in[1] ), .ZN(
        \SB1_2_19/buf_output[3] ) );
  NAND3_X2 U9943 ( .A1(\SB1_0_14/i0_0 ), .A2(\SB1_0_14/i0_4 ), .A3(
        \SB1_0_14/i1_5 ), .ZN(\SB1_0_14/Component_Function_2/NAND4_in[3] ) );
  XOR2_X1 U9944 ( .A1(\MC_ARK_ARC_1_1/temp5[171] ), .A2(n4066), .Z(
        \MC_ARK_ARC_1_1/buf_output[171] ) );
  NAND3_X1 U9949 ( .A1(\SB1_1_2/i0[8] ), .A2(\SB1_1_2/i0_3 ), .A3(
        \SB1_1_2/i1_7 ), .ZN(\SB1_1_2/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U9950 ( .A1(\MC_ARK_ARC_1_3/temp4[109] ), .A2(n4068), .Z(n681) );
  XOR2_X1 U9951 ( .A1(\RI5[3][19] ), .A2(\RI5[3][175] ), .Z(n4068) );
  XOR2_X1 U9955 ( .A1(n2761), .A2(n4070), .Z(\MC_ARK_ARC_1_2/buf_output[129] )
         );
  XOR2_X1 U9956 ( .A1(\MC_ARK_ARC_1_2/temp4[129] ), .A2(
        \MC_ARK_ARC_1_2/temp1[129] ), .Z(n4070) );
  NAND3_X2 U9961 ( .A1(\SB2_0_21/i0_3 ), .A2(\SB2_0_21/i1[9] ), .A3(
        \SB2_0_21/i0[6] ), .ZN(n4076) );
  XOR2_X1 U9968 ( .A1(n4081), .A2(n4080), .Z(\MC_ARK_ARC_1_0/temp6[62] ) );
  XOR2_X1 U9969 ( .A1(\RI5[0][164] ), .A2(n101), .Z(n4080) );
  NAND3_X2 U9972 ( .A1(\SB2_0_21/i0_3 ), .A2(\SB2_0_21/i0_4 ), .A3(
        \SB2_0_21/i0[10] ), .ZN(n1077) );
  XOR2_X1 U9973 ( .A1(\MC_ARK_ARC_1_2/temp2[73] ), .A2(
        \MC_ARK_ARC_1_2/temp1[73] ), .Z(n4084) );
  NAND4_X2 U9974 ( .A1(n4093), .A2(\SB2_2_24/Component_Function_1/NAND4_in[3] ), .A3(\SB2_2_24/Component_Function_1/NAND4_in[1] ), .A4(
        \SB2_2_24/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_2_24/buf_output[1] ) );
  XOR2_X1 U9975 ( .A1(\MC_ARK_ARC_1_1/temp5[21] ), .A2(
        \MC_ARK_ARC_1_1/temp6[21] ), .Z(\MC_ARK_ARC_1_1/buf_output[21] ) );
  NAND4_X2 U9976 ( .A1(\SB2_1_24/Component_Function_3/NAND4_in[0] ), .A2(n4234), .A3(\SB2_1_24/Component_Function_3/NAND4_in[1] ), .A4(
        \SB2_1_24/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_1_24/buf_output[3] ) );
  NAND3_X1 U9977 ( .A1(\SB4_14/i0_3 ), .A2(\SB4_14/i0_4 ), .A3(\SB4_14/i0[10] ), .ZN(\SB4_14/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U9978 ( .A1(\SB4_10/i0[10] ), .A2(\SB4_10/i0_3 ), .A3(\SB4_10/i0_4 ), .ZN(\SB4_10/Component_Function_0/NAND4_in[2] ) );
  INV_X2 U9979 ( .I(\SB1_1_27/buf_output[2] ), .ZN(\SB2_1_24/i1[9] ) );
  NAND4_X2 U9982 ( .A1(\SB1_1_27/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_1_27/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_1_27/Component_Function_4/NAND4_in[1] ), .A4(
        \SB1_1_27/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_1_27/buf_output[4] ) );
  XOR2_X1 U9983 ( .A1(n4235), .A2(n4086), .Z(\MC_ARK_ARC_1_1/buf_output[96] )
         );
  XOR2_X1 U9984 ( .A1(\MC_ARK_ARC_1_1/temp3[96] ), .A2(
        \MC_ARK_ARC_1_1/temp4[96] ), .Z(n4086) );
  NAND2_X2 U9985 ( .A1(n2261), .A2(\SB2_3_4/i0_0 ), .ZN(
        \SB2_3_4/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U9986 ( .A1(\RI5[3][55] ), .A2(\RI5[3][79] ), .Z(
        \MC_ARK_ARC_1_3/temp2[109] ) );
  NAND3_X1 U9989 ( .A1(\SB2_3_21/i0[10] ), .A2(\SB2_3_21/i1[9] ), .A3(
        \SB2_3_21/i1_7 ), .ZN(n4089) );
  XOR2_X1 U9990 ( .A1(n4090), .A2(\MC_ARK_ARC_1_3/temp1[104] ), .Z(n4091) );
  XOR2_X1 U9991 ( .A1(\RI5[3][50] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[74] ), 
        .Z(n4090) );
  NAND3_X2 U9992 ( .A1(\SB1_0_5/i0[10] ), .A2(\SB1_0_5/i0_3 ), .A3(
        \SB1_0_5/i0[6] ), .ZN(n4241) );
  XOR2_X1 U9993 ( .A1(\MC_ARK_ARC_1_3/temp6[104] ), .A2(n4091), .Z(
        \MC_ARK_ARC_1_3/buf_output[104] ) );
  NAND3_X1 U9995 ( .A1(\SB2_2_24/i0[6] ), .A2(\SB2_2_24/i0[9] ), .A3(
        \SB2_2_24/i1_5 ), .ZN(n4093) );
  NAND3_X1 U9999 ( .A1(\SB1_0_29/i0[10] ), .A2(\SB1_0_29/i1_5 ), .A3(
        \SB1_0_29/i1[9] ), .ZN(n4095) );
  NAND3_X1 U10000 ( .A1(\SB1_2_28/i0_3 ), .A2(\SB1_2_28/i0[8] ), .A3(
        \SB1_2_28/i1_7 ), .ZN(\SB1_2_28/Component_Function_1/NAND4_in[1] ) );
  NAND3_X2 U10002 ( .A1(\SB2_1_11/i0[9] ), .A2(\SB2_1_11/i0[8] ), .A3(
        \SB2_1_11/i0_3 ), .ZN(\SB2_1_11/Component_Function_2/NAND4_in[2] ) );
  XOR2_X1 U10009 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[133] ), .A2(\RI5[2][139] ), .Z(\MC_ARK_ARC_1_2/temp1[139] ) );
  NAND3_X2 U10012 ( .A1(\SB1_3_29/i0[9] ), .A2(\SB1_3_29/i0_4 ), .A3(
        \SB1_3_29/i0[6] ), .ZN(n4104) );
  NAND4_X2 U10014 ( .A1(\SB4_14/Component_Function_0/NAND4_in[3] ), .A2(
        \SB4_14/Component_Function_0/NAND4_in[2] ), .A3(
        \SB4_14/Component_Function_0/NAND4_in[1] ), .A4(n784), .ZN(n4123) );
  NAND3_X1 U10015 ( .A1(\SB1_1_23/i0_0 ), .A2(\SB1_1_23/i0[9] ), .A3(
        \SB1_1_23/i0[8] ), .ZN(\SB1_1_23/Component_Function_4/NAND4_in[0] ) );
  XOR2_X1 U10018 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[41] ), .A2(\RI5[3][47] ), 
        .Z(n4107) );
  XOR2_X1 U10019 ( .A1(\MC_ARK_ARC_1_3/temp5[14] ), .A2(n2768), .Z(
        \MC_ARK_ARC_1_3/buf_output[14] ) );
  NAND3_X1 U10020 ( .A1(\SB1_3_26/i0_0 ), .A2(\SB1_3_26/i0[8] ), .A3(
        \SB1_3_26/i0[9] ), .ZN(\SB1_3_26/Component_Function_4/NAND4_in[0] ) );
  NAND4_X2 U10021 ( .A1(\SB2_0_31/Component_Function_2/NAND4_in[0] ), .A2(
        n4546), .A3(\SB2_0_31/Component_Function_2/NAND4_in[1] ), .A4(
        \SB2_0_31/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB2_0_31/buf_output[2] ) );
  XOR2_X1 U10023 ( .A1(\RI5[2][77] ), .A2(\RI5[2][71] ), .Z(
        \MC_ARK_ARC_1_2/temp1[77] ) );
  NAND4_X2 U10028 ( .A1(\SB2_3_26/Component_Function_0/NAND4_in[3] ), .A2(
        n1936), .A3(\SB2_3_26/Component_Function_0/NAND4_in[0] ), .A4(
        \SB2_3_26/Component_Function_0/NAND4_in[1] ), .ZN(
        \SB2_3_26/buf_output[0] ) );
  NAND3_X1 U10029 ( .A1(\SB1_1_2/i0_0 ), .A2(\SB1_1_2/i0_3 ), .A3(
        \SB1_1_2/i0[7] ), .ZN(\SB1_1_2/Component_Function_0/NAND4_in[3] ) );
  XOR2_X1 U10030 ( .A1(n4110), .A2(n2870), .Z(\MC_ARK_ARC_1_0/buf_output[143] ) );
  XOR2_X1 U10034 ( .A1(n4114), .A2(n4115), .Z(\MC_ARK_ARC_1_2/buf_output[104] ) );
  XOR2_X1 U10035 ( .A1(\MC_ARK_ARC_1_2/temp2[104] ), .A2(n4687), .Z(n4114) );
  XOR2_X1 U10036 ( .A1(n4221), .A2(\MC_ARK_ARC_1_2/temp4[104] ), .Z(n4115) );
  NAND3_X2 U10037 ( .A1(\SB2_1_29/i0[9] ), .A2(\SB2_1_29/i0_3 ), .A3(
        \SB2_1_29/i0[8] ), .ZN(\SB2_1_29/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U10042 ( .A1(\SB1_2_6/i0[10] ), .A2(\SB1_2_6/i0_0 ), .A3(
        \SB1_2_6/i0[6] ), .ZN(\SB1_2_6/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U10043 ( .A1(\RI1[1][59] ), .A2(\SB1_1_22/i0[10] ), .A3(
        \SB1_1_22/i0_4 ), .ZN(\SB1_1_22/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U10044 ( .A1(\MC_ARK_ARC_1_3/temp5[64] ), .A2(
        \MC_ARK_ARC_1_3/temp6[64] ), .Z(\MC_ARK_ARC_1_3/buf_output[64] ) );
  INV_X4 U10045 ( .I(n4273), .ZN(\SB1_1_22/buf_output[2] ) );
  XOR2_X1 U10046 ( .A1(\RI5[1][77] ), .A2(n203), .Z(n4118) );
  XOR2_X1 U10047 ( .A1(\RI5[1][113] ), .A2(\RI5[1][71] ), .Z(n4119) );
  NAND2_X2 U10049 ( .A1(\SB2_2_0/i0_0 ), .A2(\SB2_2_0/i3[0] ), .ZN(n4121) );
  XOR2_X1 U10050 ( .A1(n4123), .A2(n27), .Z(Ciphertext[102]) );
  XOR2_X1 U10051 ( .A1(\MC_ARK_ARC_1_1/temp5[110] ), .A2(n4124), .Z(n4557) );
  XOR2_X1 U10052 ( .A1(\MC_ARK_ARC_1_1/temp3[110] ), .A2(n2905), .Z(n4124) );
  XOR2_X1 U10054 ( .A1(\RI5[3][159] ), .A2(\RI5[3][153] ), .Z(n4125) );
  NAND3_X1 U10055 ( .A1(\SB4_11/i0_3 ), .A2(\SB4_11/i0[8] ), .A3(\SB4_11/i1_7 ), .ZN(\SB4_11/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U10056 ( .A1(n3683), .A2(\SB4_13/i3[0] ), .A3(\SB4_13/i1_5 ), .ZN(
        \SB4_13/Component_Function_3/NAND4_in[3] ) );
  NAND4_X2 U10057 ( .A1(\SB2_3_5/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_3_5/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_3_5/Component_Function_2/NAND4_in[1] ), .A4(n4126), .ZN(
        \SB2_3_5/buf_output[2] ) );
  XOR2_X1 U10059 ( .A1(\MC_ARK_ARC_1_3/temp3[155] ), .A2(
        \MC_ARK_ARC_1_3/temp4[155] ), .Z(n4127) );
  XOR2_X1 U10063 ( .A1(\MC_ARK_ARC_1_0/temp3[66] ), .A2(n4128), .Z(n4162) );
  XOR2_X1 U10064 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[12] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[36] ), .Z(n4128) );
  XOR2_X1 U10066 ( .A1(n4132), .A2(\MC_ARK_ARC_1_0/temp3[39] ), .Z(n4713) );
  XOR2_X1 U10067 ( .A1(\RI5[0][9] ), .A2(\RI5[0][177] ), .Z(n4132) );
  XOR2_X1 U10069 ( .A1(\MC_ARK_ARC_1_3/temp2[156] ), .A2(
        \MC_ARK_ARC_1_3/temp1[156] ), .Z(n4134) );
  NAND4_X2 U10070 ( .A1(\SB2_2_18/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_18/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_2_18/Component_Function_4/NAND4_in[2] ), .A4(n4135), .ZN(
        \SB2_2_18/buf_output[4] ) );
  NAND3_X1 U10071 ( .A1(\SB3_15/i1[9] ), .A2(\SB3_15/i0[10] ), .A3(
        \SB3_15/i1_7 ), .ZN(n4137) );
  NAND4_X2 U10072 ( .A1(\SB1_1_2/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_1_2/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_1_2/Component_Function_1/NAND4_in[0] ), .A4(n4138), .ZN(
        \SB1_1_2/buf_output[1] ) );
  NAND4_X2 U10073 ( .A1(\SB2_3_4/Component_Function_1/NAND4_in[1] ), .A2(n1484), .A3(\SB2_3_4/Component_Function_1/NAND4_in[0] ), .A4(n4139), .ZN(
        \SB2_3_4/buf_output[1] ) );
  XOR2_X1 U10074 ( .A1(\RI5[3][106] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[142] ), .Z(\MC_ARK_ARC_1_3/temp3[40] ) );
  XOR2_X1 U10075 ( .A1(\RI5[1][3] ), .A2(\RI5[1][27] ), .Z(
        \MC_ARK_ARC_1_1/temp2[57] ) );
  XOR2_X1 U10078 ( .A1(\MC_ARK_ARC_1_2/temp3[171] ), .A2(
        \MC_ARK_ARC_1_2/temp4[171] ), .Z(\MC_ARK_ARC_1_2/temp6[171] ) );
  XOR2_X1 U10079 ( .A1(\RI5[0][20] ), .A2(n102), .Z(n4144) );
  NAND3_X1 U10080 ( .A1(\SB2_1_9/i0_0 ), .A2(\SB2_1_9/i3[0] ), .A3(
        \SB2_1_9/i1_7 ), .ZN(\SB2_1_9/Component_Function_4/NAND4_in[1] ) );
  NAND3_X2 U10081 ( .A1(\SB2_1_2/i0_4 ), .A2(\SB2_1_2/i0_3 ), .A3(
        \SB2_1_2/i1[9] ), .ZN(\SB2_1_2/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U10087 ( .A1(\MC_ARK_ARC_1_1/temp5[12] ), .A2(n4148), .Z(
        \MC_ARK_ARC_1_1/buf_output[12] ) );
  XOR2_X1 U10088 ( .A1(\MC_ARK_ARC_1_1/temp3[12] ), .A2(
        \MC_ARK_ARC_1_1/temp4[12] ), .Z(n4148) );
  NAND3_X2 U10089 ( .A1(\SB2_1_14/i0[10] ), .A2(\SB2_1_14/i0_0 ), .A3(
        \SB2_1_14/i0[6] ), .ZN(\SB2_1_14/Component_Function_5/NAND4_in[1] ) );
  NOR2_X2 U10091 ( .A1(n1040), .A2(n987), .ZN(n4149) );
  XOR2_X1 U10093 ( .A1(\MC_ARK_ARC_1_1/temp3[71] ), .A2(
        \MC_ARK_ARC_1_1/temp4[71] ), .Z(n4150) );
  NAND3_X1 U10094 ( .A1(\SB2_2_19/i0_3 ), .A2(\SB2_2_19/i0[10] ), .A3(
        \SB2_2_19/i0_4 ), .ZN(\SB2_2_19/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U10097 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[97] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[133] ), .Z(\MC_ARK_ARC_1_2/temp3[31] )
         );
  NAND3_X1 U10100 ( .A1(\SB1_3_15/i0_3 ), .A2(\SB1_3_15/i0[8] ), .A3(
        \SB1_3_15/i1_7 ), .ZN(\SB1_3_15/Component_Function_1/NAND4_in[1] ) );
  INV_X2 U10104 ( .I(\RI3[0][68] ), .ZN(\SB2_0_20/i1[9] ) );
  NAND3_X2 U10105 ( .A1(\SB2_1_1/i0[10] ), .A2(\SB2_1_1/i1[9] ), .A3(
        \SB2_1_1/i1_7 ), .ZN(n4155) );
  NAND4_X2 U10106 ( .A1(\SB2_0_16/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_0_16/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_0_16/Component_Function_4/NAND4_in[1] ), .A4(n4157), .ZN(
        \SB2_0_16/buf_output[4] ) );
  INV_X2 U10112 ( .I(\SB1_3_20/buf_output[3] ), .ZN(\SB2_3_18/i0[8] ) );
  NAND4_X2 U10113 ( .A1(\SB1_3_20/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_3_20/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_3_20/Component_Function_3/NAND4_in[2] ), .A4(n1186), .ZN(
        \SB1_3_20/buf_output[3] ) );
  XOR2_X1 U10115 ( .A1(\RI5[1][0] ), .A2(\RI5[1][6] ), .Z(n4160) );
  XOR2_X1 U10116 ( .A1(\MC_ARK_ARC_1_0/temp1[162] ), .A2(
        \MC_ARK_ARC_1_0/temp2[162] ), .Z(\MC_ARK_ARC_1_0/temp5[162] ) );
  XOR2_X1 U10117 ( .A1(n4162), .A2(n4161), .Z(\MC_ARK_ARC_1_0/buf_output[66] )
         );
  XOR2_X1 U10118 ( .A1(\MC_ARK_ARC_1_0/temp4[66] ), .A2(
        \MC_ARK_ARC_1_0/temp1[66] ), .Z(n4161) );
  NAND3_X1 U10119 ( .A1(\SB1_0_17/i0_0 ), .A2(\SB1_0_17/i0[10] ), .A3(
        \SB1_0_17/i0[6] ), .ZN(n4163) );
  NAND4_X2 U10120 ( .A1(\SB2_0_30/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_0_30/Component_Function_0/NAND4_in[0] ), .A3(
        \SB2_0_30/Component_Function_0/NAND4_in[2] ), .A4(n4164), .ZN(
        \SB2_0_30/buf_output[0] ) );
  NAND3_X1 U10122 ( .A1(\SB1_0_11/i0[10] ), .A2(\SB1_0_11/i1[9] ), .A3(
        \SB1_0_11/i1_5 ), .ZN(n652) );
  XOR2_X1 U10124 ( .A1(n4165), .A2(\MC_ARK_ARC_1_0/temp6[30] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[30] ) );
  XOR2_X1 U10125 ( .A1(\MC_ARK_ARC_1_0/temp2[30] ), .A2(
        \MC_ARK_ARC_1_0/temp1[30] ), .Z(n4165) );
  XOR2_X1 U10127 ( .A1(\MC_ARK_ARC_1_1/temp5[173] ), .A2(n4166), .Z(
        \MC_ARK_ARC_1_1/buf_output[173] ) );
  XOR2_X1 U10128 ( .A1(\MC_ARK_ARC_1_1/temp4[173] ), .A2(n4393), .Z(n4166) );
  XOR2_X1 U10130 ( .A1(n2805), .A2(\MC_ARK_ARC_1_0/temp5[84] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[84] ) );
  NAND3_X2 U10132 ( .A1(\SB2_0_9/i0[10] ), .A2(\RI3[0][134] ), .A3(
        \SB2_0_9/i0[6] ), .ZN(n4318) );
  XOR2_X1 U10134 ( .A1(\MC_ARK_ARC_1_1/temp5[14] ), .A2(
        \MC_ARK_ARC_1_1/temp6[14] ), .Z(\MC_ARK_ARC_1_1/buf_output[14] ) );
  NAND3_X1 U10135 ( .A1(\SB4_15/i0[10] ), .A2(\SB4_15/i0_3 ), .A3(
        \SB4_15/i0[6] ), .ZN(\SB4_15/Component_Function_2/NAND4_in[1] ) );
  NAND4_X2 U10138 ( .A1(\SB1_2_29/Component_Function_5/NAND4_in[1] ), .A2(
        n4288), .A3(\SB1_2_29/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_2_29/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_2_29/buf_output[5] ) );
  NAND4_X2 U10141 ( .A1(\SB2_1_2/Component_Function_0/NAND4_in[1] ), .A2(n1482), .A3(n1483), .A4(\SB2_1_2/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_1_2/buf_output[0] ) );
  NAND3_X1 U10142 ( .A1(\SB3_19/i0_3 ), .A2(\SB3_19/i0_0 ), .A3(\SB3_19/i0[7] ), .ZN(\SB3_19/Component_Function_0/NAND4_in[3] ) );
  XOR2_X1 U10148 ( .A1(\RI5[3][88] ), .A2(\RI5[3][94] ), .Z(
        \MC_ARK_ARC_1_3/temp1[94] ) );
  NAND4_X2 U10149 ( .A1(\SB2_2_19/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_2_19/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_2_19/Component_Function_4/NAND4_in[3] ), .A4(n4169), .ZN(
        \SB2_2_19/buf_output[4] ) );
  NAND4_X2 U10150 ( .A1(\SB2_3_17/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_3_17/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_17/Component_Function_2/NAND4_in[3] ), .A4(n4171), .ZN(
        \SB2_3_17/buf_output[2] ) );
  NAND3_X2 U10151 ( .A1(\SB2_3_17/i0[10] ), .A2(n4763), .A3(\SB2_3_17/i1[9] ), 
        .ZN(n4171) );
  NOR2_X2 U10155 ( .A1(n4175), .A2(n4174), .ZN(n4273) );
  NAND3_X2 U10156 ( .A1(\SB1_1_22/i1_5 ), .A2(\SB1_1_22/i0[10] ), .A3(
        \SB1_1_22/i1[9] ), .ZN(n1493) );
  XOR2_X1 U10157 ( .A1(n4177), .A2(n4176), .Z(n1989) );
  XOR2_X1 U10158 ( .A1(\RI5[1][51] ), .A2(n201), .Z(n4176) );
  NAND4_X2 U10164 ( .A1(\SB2_1_6/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_1_6/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_1_6/Component_Function_1/NAND4_in[0] ), .A4(n4181), .ZN(
        \SB2_1_6/buf_output[1] ) );
  NAND3_X1 U10165 ( .A1(\SB2_1_6/i0[6] ), .A2(\SB2_1_6/i1_5 ), .A3(
        \SB1_1_11/buf_output[0] ), .ZN(n4181) );
  XOR2_X1 U10166 ( .A1(n2455), .A2(n4183), .Z(\MC_ARK_ARC_1_2/buf_output[99] )
         );
  XOR2_X1 U10168 ( .A1(n2427), .A2(n4184), .Z(\MC_ARK_ARC_1_3/buf_output[94] )
         );
  NAND3_X2 U10169 ( .A1(\SB1_3_23/i0_0 ), .A2(\SB1_3_23/i0[10] ), .A3(
        \SB1_3_23/i0[6] ), .ZN(\SB1_3_23/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U10175 ( .A1(\SB3_18/buf_output[4] ), .A2(\SB4_17/i1_5 ), .A3(
        \SB4_17/i1[9] ), .ZN(n4188) );
  INV_X2 U10176 ( .I(\SB1_2_29/buf_output[5] ), .ZN(\SB2_2_29/i1_5 ) );
  NAND3_X1 U10177 ( .A1(\SB3_15/i0[10] ), .A2(\MC_ARK_ARC_1_3/buf_output[97] ), 
        .A3(\MC_ARK_ARC_1_3/buf_output[101] ), .ZN(
        \SB3_15/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U10190 ( .A1(\SB2_1_27/i0_3 ), .A2(\SB2_1_27/i0_4 ), .A3(
        \SB2_1_27/i1[9] ), .ZN(n4195) );
  XOR2_X1 U10193 ( .A1(\RI5[0][68] ), .A2(n93), .Z(n4197) );
  XOR2_X1 U10194 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[2] ), .A2(\RI5[0][32] ), 
        .Z(n4198) );
  NAND3_X1 U10196 ( .A1(\SB1_2_19/i0[8] ), .A2(\SB1_2_19/i1_5 ), .A3(
        \SB1_2_19/i3[0] ), .ZN(\SB1_2_19/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U10197 ( .A1(\SB2_2_22/i0[6] ), .A2(\SB1_2_27/buf_output[0] ), .A3(
        \SB2_2_22/i0_4 ), .ZN(\SB2_2_22/Component_Function_5/NAND4_in[3] ) );
  XOR2_X1 U10199 ( .A1(\RI5[3][69] ), .A2(\RI5[3][105] ), .Z(
        \MC_ARK_ARC_1_3/temp3[3] ) );
  NAND4_X2 U10202 ( .A1(n2782), .A2(n1333), .A3(
        \SB1_3_16/Component_Function_5/NAND4_in[0] ), .A4(n4203), .ZN(
        \SB1_3_16/buf_output[5] ) );
  XOR2_X1 U10203 ( .A1(\MC_ARK_ARC_1_2/temp3[93] ), .A2(
        \MC_ARK_ARC_1_2/temp4[93] ), .Z(\MC_ARK_ARC_1_2/temp6[93] ) );
  XOR2_X1 U10204 ( .A1(n4205), .A2(\MC_ARK_ARC_1_3/temp1[81] ), .Z(n2497) );
  XOR2_X1 U10205 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[51] ), .A2(\RI5[3][27] ), 
        .Z(n4205) );
  XOR2_X1 U10206 ( .A1(\RI5[3][183] ), .A2(\RI5[3][147] ), .Z(
        \MC_ARK_ARC_1_3/temp3[81] ) );
  XOR2_X1 U10208 ( .A1(\SB2_0_25/buf_output[5] ), .A2(\RI5[0][17] ), .Z(
        \MC_ARK_ARC_1_0/temp2[71] ) );
  NAND4_X2 U10209 ( .A1(\SB3_26/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_26/Component_Function_3/NAND4_in[3] ), .A3(n2362), .A4(n4208), 
        .ZN(\SB3_26/buf_output[3] ) );
  XOR2_X1 U10210 ( .A1(\RI5[1][189] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[153] ), .Z(n4210) );
  XOR2_X1 U10212 ( .A1(\RI5[3][146] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[110] ), .Z(n4211) );
  NAND3_X1 U10213 ( .A1(\SB3_14/i0_0 ), .A2(\SB3_14/i0[8] ), .A3(
        \SB3_14/i0[9] ), .ZN(n4212) );
  XOR2_X1 U10214 ( .A1(\RI5[0][93] ), .A2(\RI5[0][129] ), .Z(
        \MC_ARK_ARC_1_0/temp3[27] ) );
  XOR2_X1 U10215 ( .A1(\MC_ARK_ARC_1_2/temp1[174] ), .A2(
        \MC_ARK_ARC_1_2/temp2[174] ), .Z(\MC_ARK_ARC_1_2/temp5[174] ) );
  XOR2_X1 U10219 ( .A1(\MC_ARK_ARC_1_3/temp3[105] ), .A2(
        \MC_ARK_ARC_1_3/temp4[105] ), .Z(n4214) );
  XOR2_X1 U10220 ( .A1(\MC_ARK_ARC_1_3/temp4[190] ), .A2(
        \MC_ARK_ARC_1_3/temp3[190] ), .Z(\MC_ARK_ARC_1_3/temp6[190] ) );
  NAND4_X2 U10224 ( .A1(\SB1_1_30/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_1_30/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_1_30/Component_Function_1/NAND4_in[0] ), .A4(n4218), .ZN(
        \SB1_1_30/buf_output[1] ) );
  XOR2_X1 U10225 ( .A1(\RI5[1][50] ), .A2(\RI5[1][86] ), .Z(
        \MC_ARK_ARC_1_1/temp3[176] ) );
  NAND3_X2 U10226 ( .A1(\SB2_1_24/i0[6] ), .A2(\SB2_1_24/i0_4 ), .A3(
        \SB2_1_24/i0[9] ), .ZN(\SB2_1_24/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U10227 ( .A1(\SB1_1_28/i0_3 ), .A2(\SB1_1_28/i0[8] ), .A3(
        \SB1_1_28/i1_7 ), .ZN(\SB1_1_28/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U10230 ( .A1(\RI5[2][98] ), .A2(\RI5[2][104] ), .Z(n4221) );
  NAND3_X1 U10232 ( .A1(\SB4_25/i0[9] ), .A2(\SB4_25/i0_3 ), .A3(
        \SB4_25/i0[8] ), .ZN(\SB4_25/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U10234 ( .A1(\SB2_1_24/i0[10] ), .A2(\SB2_1_24/i1_7 ), .A3(
        \SB2_1_24/i1[9] ), .ZN(n4234) );
  XOR2_X1 U10235 ( .A1(\RI5[1][15] ), .A2(\RI5[1][51] ), .Z(
        \MC_ARK_ARC_1_1/temp3[141] ) );
  XOR2_X1 U10238 ( .A1(\RI5[1][7] ), .A2(\RI5[1][175] ), .Z(
        \MC_ARK_ARC_1_1/temp2[37] ) );
  XOR2_X1 U10239 ( .A1(\MC_ARK_ARC_1_1/temp1[7] ), .A2(
        \MC_ARK_ARC_1_1/temp2[7] ), .Z(n4287) );
  NAND4_X2 U10242 ( .A1(\SB2_1_31/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_1_31/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_31/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_31/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_1_31/buf_output[1] ) );
  XOR2_X1 U10244 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[154] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[178] ), .Z(\MC_ARK_ARC_1_3/temp2[16] )
         );
  NAND3_X2 U10245 ( .A1(\SB1_3_16/i0[10] ), .A2(\SB1_3_16/i1[9] ), .A3(
        \SB1_3_16/i1_5 ), .ZN(\SB1_3_16/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U10246 ( .A1(\SB2_3_17/i0_3 ), .A2(\SB2_3_17/i1[9] ), .A3(
        \SB2_3_17/i0_4 ), .ZN(\SB2_3_17/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U10247 ( .A1(\RI5[2][17] ), .A2(\RI5[2][23] ), .Z(n882) );
  NAND2_X1 U10248 ( .A1(\SB1_0_12/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_0_12/Component_Function_4/NAND4_in[1] ), .ZN(n4227) );
  NAND3_X1 U10251 ( .A1(\SB3_16/i0_3 ), .A2(\SB3_16/i0[10] ), .A3(
        \SB3_16/i0_4 ), .ZN(n4230) );
  NOR2_X2 U10252 ( .A1(n4243), .A2(n4395), .ZN(n4231) );
  XOR2_X1 U10253 ( .A1(n4232), .A2(n4233), .Z(\MC_ARK_ARC_1_3/buf_output[92] )
         );
  XOR2_X1 U10254 ( .A1(\MC_ARK_ARC_1_3/temp3[92] ), .A2(
        \MC_ARK_ARC_1_3/temp2[92] ), .Z(n4233) );
  NAND3_X1 U10256 ( .A1(\RI3[0][160] ), .A2(\SB2_0_5/i1_7 ), .A3(
        \SB2_0_5/i0[8] ), .ZN(\SB2_0_5/Component_Function_1/NAND4_in[3] ) );
  XOR2_X1 U10257 ( .A1(\MC_ARK_ARC_1_1/temp1[96] ), .A2(
        \MC_ARK_ARC_1_1/temp2[96] ), .Z(n4235) );
  XOR2_X1 U10260 ( .A1(n2809), .A2(\MC_ARK_ARC_1_3/temp5[50] ), .Z(n1401) );
  XOR2_X1 U10261 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[182] ), .A2(\RI5[3][158] ), .Z(\MC_ARK_ARC_1_3/temp2[20] ) );
  NAND3_X2 U10263 ( .A1(\SB2_1_13/i0[10] ), .A2(\SB1_1_18/buf_output[0] ), 
        .A3(\SB2_1_13/i0_3 ), .ZN(n2703) );
  NAND3_X1 U10270 ( .A1(\SB3_21/buf_output[3] ), .A2(\SB4_19/i1[9] ), .A3(
        \SB4_19/i1_5 ), .ZN(\SB4_19/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U10272 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[176] ), .A2(\RI5[3][140] ), .Z(\MC_ARK_ARC_1_3/temp3[74] ) );
  XOR2_X1 U10273 ( .A1(\MC_ARK_ARC_1_2/temp1[139] ), .A2(
        \MC_ARK_ARC_1_2/temp2[139] ), .Z(\MC_ARK_ARC_1_2/temp5[139] ) );
  XOR2_X1 U10274 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[68] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[92] ), .Z(\MC_ARK_ARC_1_2/temp2[122] )
         );
  NAND3_X2 U10275 ( .A1(\SB2_1_16/i0[6] ), .A2(\SB2_1_16/i0_3 ), .A3(
        \SB2_1_16/i0[10] ), .ZN(\SB2_1_16/Component_Function_2/NAND4_in[1] )
         );
  NAND3_X1 U10276 ( .A1(\SB1_0_5/i0_0 ), .A2(\SB1_0_5/i3[0] ), .A3(
        \SB1_0_5/i1_7 ), .ZN(\SB1_0_5/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U10277 ( .A1(\SB2_3_8/i0_3 ), .A2(\SB2_3_8/i0[10] ), .A3(
        \SB1_3_9/buf_output[4] ), .ZN(
        \SB2_3_8/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U10278 ( .A1(\SB3_20/i0[9] ), .A2(\SB3_20/i0[10] ), .A3(
        \SB3_20/i0_3 ), .ZN(\SB3_20/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U10281 ( .A1(\SB1_1_27/i0[10] ), .A2(\SB1_1_27/i0[6] ), .A3(
        \SB1_1_27/i0_3 ), .ZN(\SB1_1_27/Component_Function_2/NAND4_in[1] ) );
  XOR2_X1 U10283 ( .A1(\RI5[0][135] ), .A2(\RI5[0][111] ), .Z(
        \MC_ARK_ARC_1_0/temp2[165] ) );
  NAND3_X1 U10284 ( .A1(\SB1_3_29/i1[9] ), .A2(\SB1_3_29/i1_5 ), .A3(
        \SB1_3_29/i0[10] ), .ZN(\SB1_3_29/Component_Function_2/NAND4_in[0] )
         );
  NAND3_X2 U10285 ( .A1(\SB2_2_3/i0_3 ), .A2(\SB1_2_4/buf_output[4] ), .A3(
        \SB2_2_3/i1[9] ), .ZN(\SB2_2_3/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U10287 ( .A1(n4246), .A2(\MC_ARK_ARC_1_1/temp2[5] ), .Z(n4456) );
  XOR2_X1 U10288 ( .A1(\RI5[1][5] ), .A2(\RI5[1][191] ), .Z(n4246) );
  NAND4_X2 U10291 ( .A1(\SB2_2_31/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_2_31/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_2_31/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_31/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_2_31/buf_output[1] ) );
  NAND4_X2 U10294 ( .A1(\SB2_2_19/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_2_19/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_2_19/Component_Function_0/NAND4_in[3] ), .A4(
        \SB2_2_19/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_2_19/buf_output[0] ) );
  NAND3_X2 U10297 ( .A1(\SB4_18/i0_0 ), .A2(\SB4_18/i0[6] ), .A3(
        \SB4_18/i0[10] ), .ZN(n4251) );
  XOR2_X1 U10299 ( .A1(\RI5[1][171] ), .A2(\RI5[1][3] ), .Z(
        \MC_ARK_ARC_1_1/temp2[33] ) );
  XOR2_X1 U10301 ( .A1(\MC_ARK_ARC_1_2/temp3[183] ), .A2(
        \MC_ARK_ARC_1_2/temp4[183] ), .Z(n4253) );
  XOR2_X1 U10302 ( .A1(\MC_ARK_ARC_1_1/temp5[34] ), .A2(n4254), .Z(
        \MC_ARK_ARC_1_1/buf_output[34] ) );
  XOR2_X1 U10304 ( .A1(\MC_ARK_ARC_1_1/temp6[180] ), .A2(n4255), .Z(
        \MC_ARK_ARC_1_1/buf_output[180] ) );
  XOR2_X1 U10305 ( .A1(n4586), .A2(\MC_ARK_ARC_1_1/temp2[180] ), .Z(n4255) );
  XOR2_X1 U10306 ( .A1(\SB2_2_12/buf_output[2] ), .A2(n481), .Z(n4256) );
  NAND3_X2 U10310 ( .A1(\SB4_18/i0_0 ), .A2(\SB4_18/i3[0] ), .A3(\SB4_18/i1_7 ), .ZN(n2627) );
  NAND3_X1 U10313 ( .A1(\SB1_0_22/i0_0 ), .A2(\SB1_0_22/i0[7] ), .A3(
        \SB1_0_22/i0_3 ), .ZN(\SB1_0_22/Component_Function_0/NAND4_in[3] ) );
  NAND4_X2 U10314 ( .A1(\SB2_0_10/Component_Function_5/NAND4_in[1] ), .A2(
        \SB2_0_10/Component_Function_5/NAND4_in[2] ), .A3(
        \SB2_0_10/Component_Function_5/NAND4_in[3] ), .A4(n4258), .ZN(
        \SB2_0_10/buf_output[5] ) );
  NAND4_X2 U10315 ( .A1(\SB1_0_13/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_13/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_0_13/Component_Function_5/NAND4_in[0] ), .A4(n4259), .ZN(
        \RI3[0][113] ) );
  NAND3_X1 U10316 ( .A1(\SB2_0_27/i0[6] ), .A2(n2679), .A3(\SB2_0_27/i1_5 ), 
        .ZN(\SB2_0_27/Component_Function_1/NAND4_in[2] ) );
  NAND4_X2 U10322 ( .A1(\SB1_1_10/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_1_10/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_10/Component_Function_0/NAND4_in[0] ), .A4(n4261), .ZN(
        \SB1_1_10/buf_output[0] ) );
  INV_X2 U10323 ( .I(\SB1_2_27/buf_output[2] ), .ZN(\SB2_2_24/i1[9] ) );
  NAND4_X2 U10324 ( .A1(\SB1_2_27/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_27/Component_Function_2/NAND4_in[2] ), .A3(
        \SB1_2_27/Component_Function_2/NAND4_in[1] ), .A4(n1801), .ZN(
        \SB1_2_27/buf_output[2] ) );
  NAND3_X1 U10325 ( .A1(\SB2_1_22/i0_3 ), .A2(\SB2_1_22/i0_0 ), .A3(
        \SB2_1_22/i0[7] ), .ZN(\SB2_1_22/Component_Function_0/NAND4_in[3] ) );
  NAND4_X2 U10326 ( .A1(\SB1_2_17/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_2_17/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_2_17/Component_Function_0/NAND4_in[3] ), .A4(
        \SB1_2_17/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_2_17/buf_output[0] ) );
  NAND4_X2 U10327 ( .A1(\SB2_2_3/Component_Function_4/NAND4_in[1] ), .A2(n4263), .A3(\SB2_2_3/Component_Function_4/NAND4_in[0] ), .A4(n2802), .ZN(
        \SB2_2_3/buf_output[4] ) );
  INV_X2 U10330 ( .I(\SB1_2_19/buf_output[3] ), .ZN(\SB2_2_17/i0[8] ) );
  NAND3_X1 U10332 ( .A1(\SB2_2_3/i0_3 ), .A2(\SB2_2_3/i0[10] ), .A3(
        \SB2_2_3/i0[9] ), .ZN(n4263) );
  NAND3_X1 U10334 ( .A1(\SB1_1_5/i0[10] ), .A2(\SB1_1_5/i1_5 ), .A3(
        \SB1_1_5/i1[9] ), .ZN(\SB1_1_5/Component_Function_2/NAND4_in[0] ) );
  INV_X2 U10337 ( .I(\SB3_21/buf_output[2] ), .ZN(\SB4_18/i1[9] ) );
  XOR2_X1 U10341 ( .A1(n4266), .A2(n1272), .Z(\MC_ARK_ARC_1_2/buf_output[68] )
         );
  XOR2_X1 U10342 ( .A1(\MC_ARK_ARC_1_2/temp3[68] ), .A2(n2308), .Z(n4266) );
  XOR2_X1 U10346 ( .A1(\RI5[1][125] ), .A2(n168), .Z(n4268) );
  NAND4_X2 U10348 ( .A1(\SB1_3_29/Component_Function_3/NAND4_in[2] ), .A2(
        \SB1_3_29/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_3_29/Component_Function_3/NAND4_in[1] ), .A4(
        \SB1_3_29/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_3_29/buf_output[3] ) );
  XOR2_X1 U10350 ( .A1(\RI5[2][15] ), .A2(\RI5[2][171] ), .Z(
        \MC_ARK_ARC_1_2/temp3[105] ) );
  NAND2_X2 U10352 ( .A1(\SB1_2_31/i0_0 ), .A2(\SB1_2_31/i3[0] ), .ZN(n4271) );
  XOR2_X1 U10354 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[119] ), .A2(\RI5[3][125] ), .Z(\MC_ARK_ARC_1_3/temp1[125] ) );
  XOR2_X1 U10356 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[74] ), .A2(\RI5[1][98] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[128] ) );
  NAND3_X2 U10357 ( .A1(\SB3_20/i0[9] ), .A2(\SB3_20/i0_4 ), .A3(
        \SB3_20/i0[6] ), .ZN(n4439) );
  NAND3_X1 U10358 ( .A1(\SB4_20/i0_3 ), .A2(\SB4_20/i0_4 ), .A3(\SB4_20/i1[9] ), .ZN(\SB4_20/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U10359 ( .A1(\SB3_20/i0[9] ), .A2(\SB3_20/i1_5 ), .A3(
        \SB3_20/i0[6] ), .ZN(\SB3_20/Component_Function_1/NAND4_in[2] ) );
  XOR2_X1 U10360 ( .A1(n2359), .A2(n4274), .Z(\MC_ARK_ARC_1_0/buf_output[44] )
         );
  XOR2_X1 U10363 ( .A1(n4276), .A2(n4277), .Z(\MC_ARK_ARC_1_1/temp5[87] ) );
  XOR2_X1 U10364 ( .A1(n1383), .A2(\RI5[1][87] ), .Z(n4276) );
  XOR2_X1 U10365 ( .A1(\RI5[1][81] ), .A2(\RI5[1][57] ), .Z(n4277) );
  NAND3_X1 U10368 ( .A1(\SB1_1_26/i3[0] ), .A2(\SB1_1_26/i0[8] ), .A3(
        \SB1_1_26/i1_5 ), .ZN(n4279) );
  XOR2_X1 U10370 ( .A1(\MC_ARK_ARC_1_3/temp5[117] ), .A2(n4281), .Z(
        \MC_ARK_ARC_1_3/buf_output[117] ) );
  XOR2_X1 U10371 ( .A1(\MC_ARK_ARC_1_3/temp3[117] ), .A2(
        \MC_ARK_ARC_1_3/temp4[117] ), .Z(n4281) );
  XOR2_X1 U10373 ( .A1(\RI5[0][41] ), .A2(\RI5[0][47] ), .Z(
        \MC_ARK_ARC_1_0/temp1[47] ) );
  NAND2_X2 U10374 ( .A1(\SB2_1_11/i0[9] ), .A2(\SB2_1_11/i0[10] ), .ZN(
        \SB2_1_11/Component_Function_0/NAND4_in[0] ) );
  NAND4_X2 U10380 ( .A1(\SB2_1_11/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_1_11/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_11/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_1_11/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_1_11/buf_output[1] ) );
  XOR2_X1 U10382 ( .A1(n4290), .A2(\MC_ARK_ARC_1_3/temp4[8] ), .Z(
        \MC_ARK_ARC_1_3/temp6[8] ) );
  XOR2_X1 U10383 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[74] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[110] ), .Z(n4290) );
  NAND2_X1 U10384 ( .A1(\SB4_28/i0_3 ), .A2(n5514), .ZN(n4291) );
  NAND3_X2 U10385 ( .A1(\SB2_1_18/i0[9] ), .A2(\SB2_1_18/i0_3 ), .A3(
        \SB2_1_18/i0[8] ), .ZN(\SB2_1_18/Component_Function_2/NAND4_in[2] ) );
  XOR2_X1 U10386 ( .A1(\MC_ARK_ARC_1_0/temp6[81] ), .A2(n2170), .Z(
        \MC_ARK_ARC_1_0/buf_output[81] ) );
  NAND4_X2 U10387 ( .A1(\SB2_3_29/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_29/Component_Function_5/NAND4_in[1] ), .A3(n1734), .A4(
        \SB2_3_29/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_3_29/buf_output[5] ) );
  XOR2_X1 U10388 ( .A1(\MC_ARK_ARC_1_3/temp6[17] ), .A2(
        \MC_ARK_ARC_1_3/temp5[17] ), .Z(\MC_ARK_ARC_1_3/buf_output[17] ) );
  NAND4_X2 U10389 ( .A1(\SB3_28/Component_Function_5/NAND4_in[1] ), .A2(
        \SB3_28/Component_Function_5/NAND4_in[2] ), .A3(n4511), .A4(
        \SB3_28/Component_Function_5/NAND4_in[0] ), .ZN(\RI3[4][23] ) );
  XOR2_X1 U10393 ( .A1(\MC_ARK_ARC_1_3/temp6[22] ), .A2(
        \MC_ARK_ARC_1_3/temp5[22] ), .Z(\MC_ARK_ARC_1_3/buf_output[22] ) );
  NAND4_X2 U10395 ( .A1(\SB1_3_1/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_3_1/Component_Function_1/NAND4_in[0] ), .A3(
        \SB1_3_1/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_1/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_3_1/buf_output[1] ) );
  XOR2_X1 U10396 ( .A1(n1856), .A2(\MC_ARK_ARC_1_0/temp5[153] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[153] ) );
  XOR2_X1 U10404 ( .A1(\MC_ARK_ARC_1_0/temp4[131] ), .A2(
        \MC_ARK_ARC_1_0/temp2[131] ), .Z(n4299) );
  XOR2_X1 U10405 ( .A1(\MC_ARK_ARC_1_0/temp3[131] ), .A2(
        \MC_ARK_ARC_1_0/temp1[131] ), .Z(n4300) );
  XOR2_X1 U10407 ( .A1(\MC_ARK_ARC_1_3/temp2[55] ), .A2(
        \MC_ARK_ARC_1_3/temp1[55] ), .Z(n4303) );
  NAND3_X1 U10408 ( .A1(\SB4_22/i0_3 ), .A2(\SB4_22/i0_4 ), .A3(\SB4_22/i1[9] ), .ZN(\SB4_22/Component_Function_5/NAND4_in[2] ) );
  NAND2_X2 U10409 ( .A1(n4305), .A2(n4304), .ZN(\RI5[3][1] ) );
  XOR2_X1 U10411 ( .A1(\MC_ARK_ARC_1_2/temp6[42] ), .A2(n4306), .Z(
        \MC_ARK_ARC_1_2/buf_output[42] ) );
  XOR2_X1 U10413 ( .A1(\RI5[2][48] ), .A2(\RI5[2][72] ), .Z(
        \MC_ARK_ARC_1_2/temp2[102] ) );
  XOR2_X1 U10414 ( .A1(\RI5[0][41] ), .A2(\RI5[0][35] ), .Z(
        \MC_ARK_ARC_1_0/temp1[41] ) );
  NAND3_X2 U10415 ( .A1(\SB2_2_17/i0_4 ), .A2(\SB2_2_17/i0[9] ), .A3(
        \SB2_2_17/i0[6] ), .ZN(n4307) );
  NAND3_X2 U10418 ( .A1(\SB1_2_26/i0_4 ), .A2(\SB1_2_26/i1[9] ), .A3(
        \RI1[2][35] ), .ZN(n4311) );
  NAND3_X2 U10419 ( .A1(\SB2_3_29/i0_3 ), .A2(\RI3[3][16] ), .A3(
        \SB2_3_29/i0_0 ), .ZN(\SB2_3_29/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U10420 ( .A1(n4313), .A2(n4312), .Z(\MC_ARK_ARC_1_3/temp5[117] ) );
  XOR2_X1 U10421 ( .A1(\RI5[3][63] ), .A2(\RI5[3][117] ), .Z(n4312) );
  XOR2_X1 U10423 ( .A1(\MC_ARK_ARC_1_0/temp2[164] ), .A2(
        \MC_ARK_ARC_1_0/temp4[164] ), .Z(n4314) );
  XOR2_X1 U10425 ( .A1(\MC_ARK_ARC_1_2/temp2[13] ), .A2(
        \MC_ARK_ARC_1_2/temp1[13] ), .Z(\MC_ARK_ARC_1_2/temp5[13] ) );
  XOR2_X1 U10426 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[109] ), .A2(\RI5[0][133] ), .Z(\MC_ARK_ARC_1_0/temp2[163] ) );
  NAND4_X2 U10429 ( .A1(\SB1_0_5/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_5/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_0_5/Component_Function_5/NAND4_in[0] ), .A4(
        \SB1_0_5/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[0][161] ) );
  NAND4_X2 U10431 ( .A1(\SB1_2_17/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_2_17/Component_Function_5/NAND4_in[1] ), .A3(n4316), .A4(
        \SB1_2_17/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_2_17/buf_output[5] ) );
  XOR2_X1 U10433 ( .A1(\RI5[1][4] ), .A2(\RI5[1][10] ), .Z(
        \MC_ARK_ARC_1_1/temp1[10] ) );
  XOR2_X1 U10434 ( .A1(\RI5[1][24] ), .A2(\RI5[1][60] ), .Z(
        \MC_ARK_ARC_1_1/temp3[150] ) );
  XOR2_X1 U10435 ( .A1(\MC_ARK_ARC_1_2/temp4[53] ), .A2(
        \MC_ARK_ARC_1_2/temp3[53] ), .Z(\MC_ARK_ARC_1_2/temp6[53] ) );
  XOR2_X1 U10436 ( .A1(\MC_ARK_ARC_1_1/temp6[150] ), .A2(
        \MC_ARK_ARC_1_1/temp5[150] ), .Z(\MC_ARK_ARC_1_1/buf_output[150] ) );
  NAND3_X2 U10437 ( .A1(\SB2_2_27/i0[10] ), .A2(\SB2_2_27/i0_0 ), .A3(
        \SB2_2_27/i0[6] ), .ZN(\SB2_2_27/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U10440 ( .A1(\RI5[0][186] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[156] ), .Z(n1690) );
  OR3_X1 U10442 ( .A1(\SB2_0_5/i0_0 ), .A2(\SB2_0_5/i0[8] ), .A3(\RI3[0][161] ), .Z(\SB2_0_5/Component_Function_2/NAND4_in[0] ) );
  INV_X2 U10443 ( .I(\SB1_2_24/buf_output[3] ), .ZN(\SB2_2_22/i0[8] ) );
  XOR2_X1 U10445 ( .A1(\RI5[1][157] ), .A2(\RI5[1][181] ), .Z(
        \MC_ARK_ARC_1_1/temp2[19] ) );
  XOR2_X1 U10449 ( .A1(\RI5[1][12] ), .A2(\RI5[1][6] ), .Z(
        \MC_ARK_ARC_1_1/temp1[12] ) );
  NAND4_X2 U10452 ( .A1(\SB2_1_1/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_1_1/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_1_1/Component_Function_1/NAND4_in[2] ), .A4(n4322), .ZN(
        \SB2_1_1/buf_output[1] ) );
  NAND4_X2 U10454 ( .A1(\SB2_1_2/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_1_2/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_1_2/Component_Function_4/NAND4_in[1] ), .A4(n4323), .ZN(
        \SB2_1_2/buf_output[4] ) );
  NAND3_X2 U10458 ( .A1(\SB1_2_4/i0_0 ), .A2(\SB1_2_4/i1_5 ), .A3(
        \SB1_2_4/i0_4 ), .ZN(n4326) );
  XOR2_X1 U10459 ( .A1(n4327), .A2(n2863), .Z(\MC_ARK_ARC_1_1/buf_output[26] )
         );
  XOR2_X1 U10460 ( .A1(n2164), .A2(\MC_ARK_ARC_1_1/temp1[26] ), .Z(n4327) );
  NAND3_X1 U10462 ( .A1(\SB4_7/i0_0 ), .A2(\SB4_7/i1_7 ), .A3(\SB4_7/i3[0] ), 
        .ZN(n4329) );
  NAND4_X2 U10464 ( .A1(\SB2_3_20/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_3_20/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_20/Component_Function_0/NAND4_in[2] ), .A4(
        \SB2_3_20/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_3_20/buf_output[0] ) );
  XOR2_X1 U10465 ( .A1(\RI5[3][148] ), .A2(\RI5[3][112] ), .Z(
        \MC_ARK_ARC_1_3/temp3[46] ) );
  NAND3_X1 U10466 ( .A1(\SB4_15/i0_3 ), .A2(\SB4_15/i0[7] ), .A3(\SB4_15/i0_0 ), .ZN(\SB4_15/Component_Function_0/NAND4_in[3] ) );
  NAND4_X2 U10467 ( .A1(n1264), .A2(\SB3_15/Component_Function_0/NAND4_in[1] ), 
        .A3(n1263), .A4(n4330), .ZN(\SB3_15/buf_output[0] ) );
  NAND2_X1 U10468 ( .A1(\SB3_15/i0[9] ), .A2(\SB3_15/i0[10] ), .ZN(n4330) );
  XOR2_X1 U10469 ( .A1(\MC_ARK_ARC_1_3/temp5[128] ), .A2(
        \MC_ARK_ARC_1_3/temp6[128] ), .Z(\MC_ARK_ARC_1_3/buf_output[128] ) );
  XOR2_X1 U10470 ( .A1(\MC_ARK_ARC_1_3/temp5[96] ), .A2(
        \MC_ARK_ARC_1_3/temp6[96] ), .Z(\MC_ARK_ARC_1_3/buf_output[96] ) );
  NAND4_X2 U10471 ( .A1(\SB3_24/Component_Function_0/NAND4_in[3] ), .A2(
        \SB3_24/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_24/Component_Function_0/NAND4_in[0] ), .A4(n4331), .ZN(
        \SB3_24/buf_output[0] ) );
  INV_X1 U10474 ( .I(\SB3_15/buf_output[5] ), .ZN(\SB4_15/i1_5 ) );
  NAND4_X2 U10475 ( .A1(\SB3_15/Component_Function_5/NAND4_in[1] ), .A2(
        \SB3_15/Component_Function_5/NAND4_in[3] ), .A3(
        \SB3_15/Component_Function_5/NAND4_in[2] ), .A4(
        \SB3_15/Component_Function_5/NAND4_in[0] ), .ZN(\SB3_15/buf_output[5] ) );
  XOR2_X1 U10476 ( .A1(n2358), .A2(\MC_ARK_ARC_1_3/temp6[46] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[46] ) );
  NAND4_X2 U10477 ( .A1(\SB3_28/Component_Function_1/NAND4_in[2] ), .A2(
        \SB3_28/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_28/Component_Function_1/NAND4_in[0] ), .A4(n4332), .ZN(
        \SB3_28/buf_output[1] ) );
  NAND3_X1 U10478 ( .A1(\SB3_28/i0_4 ), .A2(\SB3_28/i0[8] ), .A3(\SB3_28/i1_7 ), .ZN(n4332) );
  NAND3_X2 U10481 ( .A1(\SB2_0_4/i0[10] ), .A2(\SB2_0_4/i1[9] ), .A3(
        \SB2_0_4/i1_7 ), .ZN(\SB2_0_4/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U10483 ( .A1(\SB1_2_17/i0[6] ), .A2(\SB1_2_17/i0[9] ), .A3(
        \SB1_2_17/i1_5 ), .ZN(\SB1_2_17/Component_Function_1/NAND4_in[2] ) );
  XOR2_X1 U10487 ( .A1(\RI5[0][99] ), .A2(\RI5[0][63] ), .Z(n4337) );
  NAND4_X2 U10488 ( .A1(n4585), .A2(
        \SB1_3_24/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_3_24/Component_Function_2/NAND4_in[2] ), .A4(n4338), .ZN(
        \SB1_3_24/buf_output[2] ) );
  XOR2_X1 U10489 ( .A1(\RI5[2][26] ), .A2(\RI5[2][20] ), .Z(n4339) );
  NAND3_X1 U10490 ( .A1(\SB2_0_11/i0_4 ), .A2(\SB1_0_14/buf_output[2] ), .A3(
        \SB2_0_11/i1_5 ), .ZN(\SB2_0_11/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 U10491 ( .A1(\SB1_1_30/i0[10] ), .A2(\SB1_1_30/i0_0 ), .A3(
        \SB1_1_30/i0[6] ), .ZN(\SB1_1_30/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U10495 ( .A1(\RI5[1][151] ), .A2(\RI5[1][127] ), .Z(n4342) );
  NAND3_X1 U10497 ( .A1(\SB4_14/i0_0 ), .A2(\SB4_14/i0_3 ), .A3(\SB4_14/i0[7] ), .ZN(\SB4_14/Component_Function_0/NAND4_in[3] ) );
  NAND3_X2 U10498 ( .A1(\SB2_3_7/i1_7 ), .A2(\SB2_3_7/i0_0 ), .A3(
        \SB2_3_7/i3[0] ), .ZN(\SB2_3_7/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U10499 ( .A1(\RI5[0][121] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[157] ), .Z(n4343) );
  NAND3_X1 U10500 ( .A1(\SB4_17/i0_4 ), .A2(\SB4_17/i0_3 ), .A3(\SB4_17/i1[9] ), .ZN(n4344) );
  NAND4_X2 U10501 ( .A1(\SB2_2_16/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_2_16/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_2_16/Component_Function_1/NAND4_in[0] ), .A4(n2299), .ZN(
        \SB2_2_16/buf_output[1] ) );
  XOR2_X1 U10503 ( .A1(\RI5[1][92] ), .A2(\RI5[1][68] ), .Z(n4345) );
  XOR2_X1 U10505 ( .A1(n4348), .A2(n4347), .Z(n4401) );
  XOR2_X1 U10506 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[101] ), .A2(n181), .Z(
        n4347) );
  XOR2_X1 U10508 ( .A1(\RI5[2][102] ), .A2(\RI5[2][66] ), .Z(
        \MC_ARK_ARC_1_2/temp3[0] ) );
  NAND3_X1 U10511 ( .A1(\SB4_17/i0[10] ), .A2(\SB4_17/i1_5 ), .A3(
        \SB4_17/i1[9] ), .ZN(n4352) );
  INV_X1 U10518 ( .I(n4355), .ZN(n4354) );
  NAND2_X1 U10519 ( .A1(\SB1_3_9/buf_output[3] ), .A2(\SB1_3_11/buf_output[1] ), .ZN(n4355) );
  XOR2_X1 U10520 ( .A1(\MC_ARK_ARC_1_1/temp3[117] ), .A2(
        \MC_ARK_ARC_1_1/temp4[117] ), .Z(n4357) );
  NAND4_X2 U10521 ( .A1(\SB1_2_1/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_2_1/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_2_1/Component_Function_3/NAND4_in[3] ), .A4(n4358), .ZN(
        \SB1_2_1/buf_output[3] ) );
  NAND3_X2 U10522 ( .A1(\SB1_2_1/i0[10] ), .A2(\SB1_2_1/i1[9] ), .A3(
        \SB1_2_1/i1_7 ), .ZN(n4358) );
  XOR2_X1 U10523 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[105] ), .A2(\RI5[0][99] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[105] ) );
  NAND4_X2 U10526 ( .A1(\SB1_3_26/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_3_26/Component_Function_3/NAND4_in[0] ), .A3(n1838), .A4(n1760), 
        .ZN(\SB1_3_26/buf_output[3] ) );
  XOR2_X1 U10527 ( .A1(n4359), .A2(n1061), .Z(n2801) );
  XOR2_X1 U10528 ( .A1(\RI5[2][152] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[128] ), .Z(n4359) );
  XOR2_X1 U10530 ( .A1(\RI5[2][155] ), .A2(\RI5[2][191] ), .Z(n4360) );
  XOR2_X1 U10531 ( .A1(n2462), .A2(n4361), .Z(\MC_ARK_ARC_1_1/buf_output[125] ) );
  XOR2_X1 U10532 ( .A1(\MC_ARK_ARC_1_1/temp3[125] ), .A2(
        \MC_ARK_ARC_1_1/temp4[125] ), .Z(n4361) );
  NAND4_X2 U10533 ( .A1(\SB1_2_11/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_11/Component_Function_0/NAND4_in[0] ), .A3(n4363), .A4(n4362), 
        .ZN(\SB1_2_11/buf_output[0] ) );
  NAND3_X1 U10534 ( .A1(\SB1_2_11/i0[6] ), .A2(\SB1_2_11/i0[7] ), .A3(
        \SB1_2_11/i0[8] ), .ZN(n4362) );
  XOR2_X1 U10537 ( .A1(\MC_ARK_ARC_1_1/temp3[121] ), .A2(
        \MC_ARK_ARC_1_1/temp4[121] ), .Z(n4654) );
  NAND4_X2 U10538 ( .A1(\SB3_17/Component_Function_4/NAND4_in[1] ), .A2(
        \SB3_17/Component_Function_4/NAND4_in[0] ), .A3(
        \SB3_17/Component_Function_4/NAND4_in[2] ), .A4(n1600), .ZN(
        \SB3_17/buf_output[4] ) );
  XOR2_X1 U10539 ( .A1(\MC_ARK_ARC_1_3/temp6[88] ), .A2(
        \MC_ARK_ARC_1_3/temp5[88] ), .Z(\MC_ARK_ARC_1_3/buf_output[88] ) );
  XOR2_X1 U10540 ( .A1(\RI5[3][93] ), .A2(\RI5[3][99] ), .Z(
        \MC_ARK_ARC_1_3/temp1[99] ) );
  NAND3_X1 U10541 ( .A1(\SB3_9/i0_4 ), .A2(\SB3_9/i0[6] ), .A3(
        \MC_ARK_ARC_1_3/buf_output[132] ), .ZN(n4366) );
  XOR2_X1 U10543 ( .A1(n4367), .A2(\MC_ARK_ARC_1_3/temp6[111] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[111] ) );
  XOR2_X1 U10544 ( .A1(\MC_ARK_ARC_1_3/temp1[111] ), .A2(
        \MC_ARK_ARC_1_3/temp2[111] ), .Z(n4367) );
  NAND3_X1 U10547 ( .A1(\SB1_0_11/i0_3 ), .A2(\SB1_0_11/i1[9] ), .A3(
        \SB1_0_11/i0[6] ), .ZN(\SB1_0_11/Component_Function_3/NAND4_in[0] ) );
  NAND4_X2 U10550 ( .A1(\SB1_2_27/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_2_27/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_27/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_27/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_2_27/buf_output[1] ) );
  XOR2_X1 U10551 ( .A1(\MC_ARK_ARC_1_2/temp4[182] ), .A2(
        \MC_ARK_ARC_1_2/temp3[182] ), .Z(\MC_ARK_ARC_1_2/temp6[182] ) );
  NAND4_X2 U10552 ( .A1(\SB2_3_0/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_0/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_3_0/Component_Function_1/NAND4_in[1] ), .A4(n4371), .ZN(
        \SB2_3_0/buf_output[1] ) );
  NOR2_X2 U10556 ( .A1(n4701), .A2(n4427), .ZN(\SB2_1_11/i0[7] ) );
  XOR2_X1 U10558 ( .A1(\MC_ARK_ARC_1_2/temp2[105] ), .A2(
        \MC_ARK_ARC_1_2/temp1[105] ), .Z(n4374) );
  XOR2_X1 U10559 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[132] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[168] ), .Z(\MC_ARK_ARC_1_3/temp3[66] )
         );
  INV_X2 U10560 ( .I(\SB1_1_20/buf_output[2] ), .ZN(\SB2_1_17/i1[9] ) );
  NAND4_X2 U10561 ( .A1(\SB1_1_20/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_1_20/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_1_20/Component_Function_2/NAND4_in[3] ), .A4(
        \SB1_1_20/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB1_1_20/buf_output[2] ) );
  XOR2_X1 U10562 ( .A1(\RI5[2][41] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[47] ), 
        .Z(n4375) );
  NAND4_X2 U10571 ( .A1(\SB2_1_25/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_25/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_25/Component_Function_4/NAND4_in[2] ), .A4(n4382), .ZN(
        \SB2_1_25/buf_output[4] ) );
  XOR2_X1 U10573 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[83] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[59] ), .Z(n4385) );
  NAND3_X1 U10574 ( .A1(\SB2_3_30/i0[8] ), .A2(\SB2_3_30/i1_7 ), .A3(
        \SB1_3_31/buf_output[4] ), .ZN(
        \SB2_3_30/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U10576 ( .A1(\SB1_2_31/i0[10] ), .A2(\SB1_2_31/i0_3 ), .A3(
        \SB1_2_31/i0_4 ), .ZN(\SB1_2_31/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U10577 ( .A1(n4622), .A2(n2348), .Z(\MC_ARK_ARC_1_1/buf_output[182] ) );
  NAND3_X1 U10579 ( .A1(\SB1_3_19/i0[10] ), .A2(\SB1_3_19/i0[6] ), .A3(
        \SB1_3_19/i0_0 ), .ZN(\SB1_3_19/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U10587 ( .A1(\SB2_1_25/i0_0 ), .A2(\SB2_1_25/i1_5 ), .A3(n1579), 
        .ZN(n4724) );
  XOR2_X1 U10590 ( .A1(\MC_ARK_ARC_1_1/temp5[145] ), .A2(n4389), .Z(
        \MC_ARK_ARC_1_1/buf_output[145] ) );
  XOR2_X1 U10591 ( .A1(\MC_ARK_ARC_1_1/temp3[145] ), .A2(
        \MC_ARK_ARC_1_1/temp4[145] ), .Z(n4389) );
  NAND4_X2 U10592 ( .A1(\SB3_15/Component_Function_2/NAND4_in[2] ), .A2(
        \SB3_15/Component_Function_2/NAND4_in[0] ), .A3(
        \SB3_15/Component_Function_2/NAND4_in[1] ), .A4(
        \SB3_15/Component_Function_2/NAND4_in[3] ), .ZN(\SB3_15/buf_output[2] ) );
  NAND4_X2 U10593 ( .A1(\SB1_3_24/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_24/Component_Function_4/NAND4_in[1] ), .A3(n4577), .A4(
        \SB1_3_24/Component_Function_4/NAND4_in[2] ), .ZN(
        \SB1_3_24/buf_output[4] ) );
  XOR2_X1 U10594 ( .A1(n2853), .A2(\MC_ARK_ARC_1_0/temp5[102] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[102] ) );
  NAND3_X1 U10595 ( .A1(\SB1_2_7/i0[6] ), .A2(\SB1_2_7/i0[8] ), .A3(
        \SB1_2_7/i0[7] ), .ZN(\SB1_2_7/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U10596 ( .A1(\SB1_0_29/i0[9] ), .A2(\SB1_0_29/i0[10] ), .A3(
        \SB1_0_29/i0_3 ), .ZN(n2225) );
  NAND3_X1 U10598 ( .A1(\SB1_1_20/i0[8] ), .A2(\SB1_1_20/i0_0 ), .A3(
        \SB1_1_20/i0[9] ), .ZN(\SB1_1_20/Component_Function_4/NAND4_in[0] ) );
  XOR2_X1 U10600 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[51] ), .A2(\RI5[3][75] ), 
        .Z(n4392) );
  XOR2_X1 U10601 ( .A1(\RI5[1][47] ), .A2(\RI5[1][83] ), .Z(n4393) );
  NAND4_X2 U10602 ( .A1(\SB1_3_4/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_3_4/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_3_4/Component_Function_1/NAND4_in[1] ), .A4(n4394), .ZN(
        \SB1_3_4/buf_output[1] ) );
  XOR2_X1 U10605 ( .A1(n4396), .A2(\MC_ARK_ARC_1_3/temp4[53] ), .Z(n1518) );
  XOR2_X1 U10606 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[119] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[155] ), .Z(n4396) );
  NAND3_X2 U10609 ( .A1(\SB1_3_23/i0_3 ), .A2(\SB1_3_23/i1[9] ), .A3(
        \SB1_3_23/i0_4 ), .ZN(n4398) );
  XOR2_X1 U10610 ( .A1(n4400), .A2(n4401), .Z(\MC_ARK_ARC_1_3/buf_output[107] ) );
  XOR2_X1 U10611 ( .A1(\MC_ARK_ARC_1_3/temp2[107] ), .A2(n4486), .Z(n4400) );
  INV_X2 U10613 ( .I(n1400), .ZN(\SB2_3_20/i1[9] ) );
  NAND4_X2 U10614 ( .A1(\SB1_3_23/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_23/Component_Function_2/NAND4_in[0] ), .A3(n2778), .A4(n2493), 
        .ZN(n1400) );
  NAND3_X2 U10615 ( .A1(\SB2_1_11/i0_0 ), .A2(\SB2_1_11/i1_5 ), .A3(
        \SB1_1_12/buf_output[4] ), .ZN(
        \SB2_1_11/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U10619 ( .A1(n6230), .A2(\SB2_2_4/i0[6] ), .A3(\SB2_2_4/i0[8] ), 
        .ZN(\SB2_2_4/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U10620 ( .A1(\MC_ARK_ARC_1_2/temp2[184] ), .A2(n4405), .Z(
        \MC_ARK_ARC_1_2/temp5[184] ) );
  XOR2_X1 U10621 ( .A1(\RI5[2][178] ), .A2(\RI5[2][184] ), .Z(n4405) );
  XOR2_X1 U10622 ( .A1(n4406), .A2(\MC_ARK_ARC_1_2/temp4[126] ), .Z(
        \MC_ARK_ARC_1_2/temp6[126] ) );
  XOR2_X1 U10623 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[0] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[36] ), .Z(n4406) );
  XOR2_X1 U10624 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[36] ), .A2(\RI5[0][72] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[162] ) );
  XOR2_X1 U10625 ( .A1(n4407), .A2(n2195), .Z(\MC_ARK_ARC_1_2/buf_output[87] )
         );
  XOR2_X1 U10626 ( .A1(n1736), .A2(\MC_ARK_ARC_1_2/temp4[87] ), .Z(n4407) );
  XOR2_X1 U10627 ( .A1(n4409), .A2(\MC_ARK_ARC_1_0/temp2[129] ), .Z(
        \MC_ARK_ARC_1_0/temp5[129] ) );
  XOR2_X1 U10628 ( .A1(\RI5[0][129] ), .A2(\RI5[0][123] ), .Z(n4409) );
  XOR2_X1 U10629 ( .A1(\MC_ARK_ARC_1_3/temp1[6] ), .A2(n4410), .Z(
        \MC_ARK_ARC_1_3/temp5[6] ) );
  XOR2_X1 U10630 ( .A1(\RI5[3][144] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[168] ), .Z(n4410) );
  NAND3_X2 U10634 ( .A1(\SB1_3_3/i0[9] ), .A2(\SB1_3_3/i0[8] ), .A3(
        \SB1_3_3/i0_3 ), .ZN(n4412) );
  XOR2_X1 U10636 ( .A1(\MC_ARK_ARC_1_2/temp1[168] ), .A2(n4414), .Z(
        \MC_ARK_ARC_1_2/temp5[168] ) );
  XOR2_X1 U10637 ( .A1(\RI5[2][114] ), .A2(\RI5[2][138] ), .Z(n4414) );
  NAND3_X1 U10638 ( .A1(\SB1_2_27/i0[10] ), .A2(\SB1_2_27/i1_5 ), .A3(
        \SB1_2_27/i1[9] ), .ZN(\SB1_2_27/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U10639 ( .A1(\RI5[0][122] ), .A2(\RI5[0][158] ), .Z(n1114) );
  XOR2_X1 U10640 ( .A1(\MC_ARK_ARC_1_0/temp1[22] ), .A2(
        \MC_ARK_ARC_1_0/temp2[22] ), .Z(n4415) );
  XOR2_X1 U10645 ( .A1(\RI5[2][77] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[131] ), 
        .Z(n4416) );
  XOR2_X1 U10646 ( .A1(n4418), .A2(n4417), .Z(\MC_ARK_ARC_1_3/temp6[47] ) );
  XOR2_X1 U10647 ( .A1(\RI5[3][149] ), .A2(n545), .Z(n4417) );
  XOR2_X1 U10648 ( .A1(\RI5[3][113] ), .A2(\RI5[3][83] ), .Z(n4418) );
  NAND3_X1 U10651 ( .A1(\SB1_1_22/i1_5 ), .A2(\SB1_1_22/i1[9] ), .A3(
        \SB1_1_22/i0_4 ), .ZN(\SB1_1_22/Component_Function_4/NAND4_in[3] ) );
  NAND4_X2 U10652 ( .A1(\SB2_0_16/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_0_16/Component_Function_2/NAND4_in[0] ), .A3(n4621), .A4(
        \SB2_0_16/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_0_16/buf_output[2] ) );
  XOR2_X1 U10653 ( .A1(\RI5[3][60] ), .A2(\RI5[3][66] ), .Z(
        \MC_ARK_ARC_1_3/temp1[66] ) );
  NAND4_X2 U10654 ( .A1(\SB3_14/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_14/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_14/Component_Function_0/NAND4_in[0] ), .A4(n4419), .ZN(
        \SB3_14/buf_output[0] ) );
  NAND3_X1 U10655 ( .A1(\SB3_14/i0_3 ), .A2(\SB3_14/i0_0 ), .A3(\SB3_14/i0[7] ), .ZN(n4419) );
  NAND4_X2 U10657 ( .A1(\SB1_0_21/Component_Function_0/NAND4_in[2] ), .A2(
        n4669), .A3(\SB1_0_21/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_0_21/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_0_21/buf_output[0] ) );
  NAND4_X2 U10660 ( .A1(\SB2_1_0/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_1_0/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_1_0/Component_Function_4/NAND4_in[1] ), .A4(n4422), .ZN(
        \SB2_1_0/buf_output[4] ) );
  NAND3_X1 U10662 ( .A1(\SB3_15/i1_5 ), .A2(\SB3_15/i0[8] ), .A3(
        \SB3_15/i3[0] ), .ZN(n4423) );
  XOR2_X1 U10664 ( .A1(\RI5[2][103] ), .A2(\RI5[2][67] ), .Z(
        \MC_ARK_ARC_1_2/temp3[1] ) );
  NAND3_X1 U10665 ( .A1(\SB3_6/i1[9] ), .A2(\RI1[4][154] ), .A3(\RI1[4][155] ), 
        .ZN(\SB3_6/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U10666 ( .A1(\SB1_2_0/i0[6] ), .A2(\SB1_2_0/i0[9] ), .A3(
        \SB1_2_0/i0_4 ), .ZN(n4425) );
  XOR2_X1 U10668 ( .A1(\RI5[2][91] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[127] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[25] ) );
  XOR2_X1 U10670 ( .A1(\RI5[2][71] ), .A2(\RI5[2][107] ), .Z(
        \MC_ARK_ARC_1_2/temp3[5] ) );
  INV_X4 U10671 ( .I(\SB2_2_31/i0[7] ), .ZN(n569) );
  NAND3_X1 U10672 ( .A1(\SB2_2_31/i0[6] ), .A2(\SB2_2_31/i0[8] ), .A3(
        \SB2_2_31/i0[7] ), .ZN(n2181) );
  NOR2_X2 U10673 ( .A1(n1950), .A2(n1948), .ZN(\SB2_2_31/i0[7] ) );
  NAND4_X2 U10674 ( .A1(\SB1_1_30/Component_Function_3/NAND4_in[2] ), .A2(
        \SB1_1_30/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_30/Component_Function_3/NAND4_in[0] ), .A4(n4430), .ZN(
        \SB1_1_30/buf_output[3] ) );
  NAND4_X2 U10675 ( .A1(\SB3_2/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_2/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_2/Component_Function_0/NAND4_in[0] ), .A4(n4431), .ZN(
        \SB3_2/buf_output[0] ) );
  XOR2_X1 U10678 ( .A1(n4433), .A2(n4434), .Z(\MC_ARK_ARC_1_2/buf_output[1] )
         );
  XOR2_X1 U10679 ( .A1(\MC_ARK_ARC_1_2/temp2[1] ), .A2(
        \MC_ARK_ARC_1_2/temp3[1] ), .Z(n4433) );
  XOR2_X1 U10680 ( .A1(\MC_ARK_ARC_1_2/temp1[1] ), .A2(
        \MC_ARK_ARC_1_2/temp4[1] ), .Z(n4434) );
  XOR2_X1 U10681 ( .A1(\MC_ARK_ARC_1_2/temp4[4] ), .A2(
        \MC_ARK_ARC_1_2/temp3[4] ), .Z(n4435) );
  XOR2_X1 U10682 ( .A1(n4436), .A2(\MC_ARK_ARC_1_1/temp1[189] ), .Z(n2799) );
  XOR2_X1 U10683 ( .A1(\RI5[1][135] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[159] ), .Z(n4436) );
  NAND3_X2 U10684 ( .A1(\SB1_2_2/i0[10] ), .A2(\SB1_2_2/i0_3 ), .A3(
        \SB1_2_2/i0[6] ), .ZN(n4437) );
  XOR2_X1 U10685 ( .A1(\RI5[2][178] ), .A2(\RI5[2][22] ), .Z(n4440) );
  NAND3_X1 U10686 ( .A1(\SB1_1_6/buf_output[4] ), .A2(\SB2_1_5/i1_7 ), .A3(
        \SB2_1_5/i0[8] ), .ZN(\SB2_1_5/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U10688 ( .A1(\SB2_1_6/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_1_6/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_6/Component_Function_0/NAND4_in[0] ), .A4(n4441), .ZN(
        \SB2_1_6/buf_output[0] ) );
  NAND3_X1 U10689 ( .A1(\SB1_1_6/i0_0 ), .A2(\SB1_1_6/i3[0] ), .A3(
        \SB1_1_6/i1_7 ), .ZN(\SB1_1_6/Component_Function_4/NAND4_in[1] ) );
  INV_X1 U10692 ( .I(\SB3_31/buf_output[5] ), .ZN(\SB4_31/i1_5 ) );
  XOR2_X1 U10694 ( .A1(n4442), .A2(\MC_ARK_ARC_1_3/temp6[102] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[102] ) );
  XOR2_X1 U10695 ( .A1(\MC_ARK_ARC_1_1/temp2[19] ), .A2(n4443), .Z(
        \MC_ARK_ARC_1_1/temp5[19] ) );
  XOR2_X1 U10696 ( .A1(\RI5[1][19] ), .A2(\RI5[1][13] ), .Z(n4443) );
  XOR2_X1 U10698 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[74] ), .A2(\RI5[3][98] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[128] ) );
  NAND4_X2 U10699 ( .A1(\SB2_0_11/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_0_11/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_0_11/Component_Function_0/NAND4_in[0] ), .A4(n4445), .ZN(
        \SB2_0_11/buf_output[0] ) );
  XOR2_X1 U10702 ( .A1(n4446), .A2(n4447), .Z(\MC_ARK_ARC_1_1/temp5[121] ) );
  XOR2_X1 U10703 ( .A1(\RI5[1][91] ), .A2(\RI5[1][121] ), .Z(n4446) );
  XOR2_X1 U10704 ( .A1(\RI5[1][115] ), .A2(\RI5[1][67] ), .Z(n4447) );
  NAND4_X2 U10710 ( .A1(\SB1_2_19/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_19/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_2_19/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_2_19/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_2_19/buf_output[0] ) );
  NAND4_X2 U10711 ( .A1(\SB2_2_14/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_2_14/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_2_14/Component_Function_1/NAND4_in[0] ), .A4(n4452), .ZN(
        \SB2_2_14/buf_output[1] ) );
  INV_X2 U10712 ( .I(\RI3[0][45] ), .ZN(\SB2_0_24/i0[8] ) );
  NAND4_X2 U10713 ( .A1(\SB1_0_26/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_26/Component_Function_3/NAND4_in[2] ), .A3(
        \SB1_0_26/Component_Function_3/NAND4_in[3] ), .A4(
        \SB1_0_26/Component_Function_3/NAND4_in[1] ), .ZN(\RI3[0][45] ) );
  NAND3_X2 U10715 ( .A1(\SB2_2_27/i0[10] ), .A2(\SB2_2_27/i0_3 ), .A3(
        \SB2_2_27/i0[6] ), .ZN(n4455) );
  NAND2_X1 U10716 ( .A1(n2225), .A2(
        \SB1_0_29/Component_Function_4/NAND4_in[3] ), .ZN(n1048) );
  XOR2_X1 U10718 ( .A1(\RI5[3][60] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[36] ), 
        .Z(n4457) );
  NAND3_X1 U10720 ( .A1(\SB4_0/i0[10] ), .A2(\SB3_3/buf_output[2] ), .A3(
        \SB4_0/i0[6] ), .ZN(\SB4_0/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U10721 ( .A1(n4461), .A2(n4460), .Z(\MC_ARK_ARC_1_3/buf_output[68] )
         );
  XOR2_X1 U10722 ( .A1(n4645), .A2(\MC_ARK_ARC_1_3/temp4[68] ), .Z(n4460) );
  XOR2_X1 U10724 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[167] ), .A2(n473), .Z(
        n4462) );
  XOR2_X1 U10725 ( .A1(\RI5[0][137] ), .A2(\RI5[0][11] ), .Z(n4463) );
  XOR2_X1 U10727 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[44] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[92] ), .Z(n4465) );
  NAND3_X1 U10728 ( .A1(\SB2_1_31/i0[8] ), .A2(\SB2_1_31/i1_7 ), .A3(
        \SB2_1_31/i0_4 ), .ZN(\SB2_1_31/Component_Function_1/NAND4_in[3] ) );
  XOR2_X1 U10730 ( .A1(\SB2_0_17/buf_output[4] ), .A2(\RI5[0][100] ), .Z(n4466) );
  NAND2_X1 U10731 ( .A1(\SB1_1_25/i1[9] ), .A2(\SB1_1_25/i0_3 ), .ZN(n4468) );
  INV_X2 U10732 ( .I(\SB1_2_8/buf_output[5] ), .ZN(\SB2_2_8/i1_5 ) );
  XOR2_X1 U10734 ( .A1(n4469), .A2(\MC_ARK_ARC_1_2/temp1[3] ), .Z(
        \MC_ARK_ARC_1_2/temp5[3] ) );
  XOR2_X1 U10736 ( .A1(\RI5[1][133] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[169] ), .Z(\MC_ARK_ARC_1_1/temp3[67] ) );
  XOR2_X1 U10737 ( .A1(n2057), .A2(n2056), .Z(n1891) );
  NAND3_X1 U10738 ( .A1(\SB3_21/i0_0 ), .A2(\SB3_21/i3[0] ), .A3(\SB3_21/i1_7 ), .ZN(\SB3_21/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U10739 ( .A1(\SB2_2_15/buf_output[1] ), .A2(\RI5[2][85] ), .Z(n4470)
         );
  NAND3_X1 U10740 ( .A1(\SB1_3_27/i0[6] ), .A2(\SB1_3_27/i0_3 ), .A3(
        \SB1_3_27/i1[9] ), .ZN(n4471) );
  NAND3_X1 U10742 ( .A1(\SB3_6/i0[10] ), .A2(\SB3_6/i1[9] ), .A3(\SB3_6/i1_7 ), 
        .ZN(\SB3_6/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U10743 ( .A1(\SB1_1_14/i1_7 ), .A2(\SB1_1_14/i0_0 ), .A3(
        \SB1_1_14/i3[0] ), .ZN(\SB1_1_14/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U10747 ( .A1(\RI5[1][71] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[95] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[125] ) );
  NAND4_X2 U10748 ( .A1(\SB1_2_31/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_2_31/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_31/Component_Function_4/NAND4_in[2] ), .A4(n4474), .ZN(
        \SB2_2_30/i0_4 ) );
  NAND3_X1 U10750 ( .A1(\SB4_12/i0_0 ), .A2(\SB4_12/i1_7 ), .A3(\SB4_12/i3[0] ), .ZN(n4476) );
  INV_X2 U10754 ( .I(\SB1_2_7/buf_output[3] ), .ZN(\SB2_2_5/i0[8] ) );
  NAND4_X2 U10755 ( .A1(\SB1_2_7/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_2_7/Component_Function_3/NAND4_in[0] ), .A3(n2856), .A4(n1819), 
        .ZN(\SB1_2_7/buf_output[3] ) );
  XOR2_X1 U10756 ( .A1(n4480), .A2(\MC_ARK_ARC_1_3/temp4[57] ), .Z(
        \MC_ARK_ARC_1_3/temp6[57] ) );
  XOR2_X1 U10757 ( .A1(\RI5[3][159] ), .A2(n3658), .Z(n4480) );
  NAND3_X1 U10760 ( .A1(\SB4_28/i0_4 ), .A2(n5514), .A3(\SB4_28/i1_5 ), .ZN(
        n4482) );
  NAND4_X2 U10761 ( .A1(\SB1_0_24/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_0_24/Component_Function_1/NAND4_in[0] ), .A3(
        \SB1_0_24/Component_Function_1/NAND4_in[1] ), .A4(n4483), .ZN(
        \RI3[0][67] ) );
  NAND3_X1 U10762 ( .A1(\SB1_0_24/i0[8] ), .A2(\SB1_0_24/i1_7 ), .A3(n356), 
        .ZN(n4483) );
  NOR2_X2 U10763 ( .A1(n747), .A2(n1213), .ZN(n2369) );
  NAND3_X1 U10765 ( .A1(\SB2_3_26/i0_3 ), .A2(\SB2_3_26/i0_4 ), .A3(
        \SB1_3_28/buf_output[3] ), .ZN(n1936) );
  XOR2_X1 U10767 ( .A1(\RI5[3][173] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[17] ), 
        .Z(n4486) );
  XOR2_X1 U10768 ( .A1(\MC_ARK_ARC_1_1/temp5[10] ), .A2(n4487), .Z(
        \MC_ARK_ARC_1_1/buf_output[10] ) );
  XOR2_X1 U10769 ( .A1(\MC_ARK_ARC_1_1/temp3[10] ), .A2(
        \MC_ARK_ARC_1_1/temp4[10] ), .Z(n4487) );
  NAND4_X2 U10770 ( .A1(\SB1_2_26/Component_Function_3/NAND4_in[3] ), .A2(
        n1574), .A3(\SB1_2_26/Component_Function_3/NAND4_in[0] ), .A4(n4488), 
        .ZN(\SB1_2_26/buf_output[3] ) );
  NAND3_X2 U10771 ( .A1(\SB2_1_20/i0[10] ), .A2(\SB2_1_20/i0_0 ), .A3(
        \SB2_1_20/i0[6] ), .ZN(\SB2_1_20/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U10772 ( .A1(\RI5[3][98] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[104] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[104] ) );
  NAND3_X1 U10773 ( .A1(n1793), .A2(\SB4_29/i0_3 ), .A3(\SB4_29/i0[10] ), .ZN(
        n4489) );
  XOR2_X1 U10774 ( .A1(\RI5[3][80] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[56] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[110] ) );
  NAND4_X2 U10778 ( .A1(\SB2_1_13/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_13/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_1_13/Component_Function_2/NAND4_in[2] ), .A4(n4493), .ZN(
        \SB2_1_13/buf_output[2] ) );
  NAND4_X2 U10779 ( .A1(\SB2_2_3/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_2_3/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_3/Component_Function_0/NAND4_in[0] ), .A4(n4494), .ZN(
        \SB2_2_3/buf_output[0] ) );
  XOR2_X1 U10781 ( .A1(\MC_ARK_ARC_1_1/temp4[41] ), .A2(n4495), .Z(
        \MC_ARK_ARC_1_1/temp6[41] ) );
  NAND4_X2 U10783 ( .A1(\SB2_1_29/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_1_29/Component_Function_0/NAND4_in[0] ), .A3(
        \SB2_1_29/Component_Function_0/NAND4_in[2] ), .A4(n4496), .ZN(
        \SB2_1_29/buf_output[0] ) );
  NAND3_X2 U10785 ( .A1(\SB2_2_26/i0[10] ), .A2(\SB2_2_26/i1[9] ), .A3(
        \SB2_2_26/i1_7 ), .ZN(n4497) );
  INV_X2 U10786 ( .I(\SB1_2_20/buf_output[2] ), .ZN(\SB2_2_17/i1[9] ) );
  XOR2_X1 U10794 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[155] ), .A2(\RI5[0][149] ), .Z(n4504) );
  XOR2_X1 U10795 ( .A1(\RI5[1][36] ), .A2(\RI5[1][12] ), .Z(n1290) );
  NAND4_X2 U10797 ( .A1(\SB2_1_11/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_1_11/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_11/Component_Function_0/NAND4_in[0] ), .A4(n4506), .ZN(
        \SB2_1_11/buf_output[0] ) );
  XOR2_X1 U10798 ( .A1(n2476), .A2(n4507), .Z(\MC_ARK_ARC_1_1/buf_output[20] )
         );
  XOR2_X1 U10799 ( .A1(\MC_ARK_ARC_1_1/temp3[20] ), .A2(
        \MC_ARK_ARC_1_1/temp4[20] ), .Z(n4507) );
  XOR2_X1 U10800 ( .A1(\MC_ARK_ARC_1_3/temp3[5] ), .A2(
        \MC_ARK_ARC_1_3/temp4[5] ), .Z(\MC_ARK_ARC_1_3/temp6[5] ) );
  XOR2_X1 U10801 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[177] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[141] ), .Z(\MC_ARK_ARC_1_2/temp3[75] )
         );
  XOR2_X1 U10802 ( .A1(\RI5[3][146] ), .A2(\RI5[3][170] ), .Z(n2314) );
  NAND4_X2 U10805 ( .A1(\SB2_0_16/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_0_16/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_0_16/Component_Function_0/NAND4_in[0] ), .A4(n4510), .ZN(
        \SB2_0_16/buf_output[0] ) );
  XOR2_X1 U10807 ( .A1(\MC_ARK_ARC_1_3/temp4[13] ), .A2(
        \MC_ARK_ARC_1_3/temp3[13] ), .Z(\MC_ARK_ARC_1_3/temp6[13] ) );
  XOR2_X1 U10808 ( .A1(\MC_ARK_ARC_1_2/temp1[72] ), .A2(
        \MC_ARK_ARC_1_2/temp2[72] ), .Z(n4512) );
  XOR2_X1 U10811 ( .A1(\MC_ARK_ARC_1_0/temp5[16] ), .A2(n4514), .Z(
        \MC_ARK_ARC_1_0/buf_output[16] ) );
  XOR2_X1 U10812 ( .A1(\MC_ARK_ARC_1_0/temp4[16] ), .A2(
        \MC_ARK_ARC_1_0/temp3[16] ), .Z(n4514) );
  NAND3_X1 U10813 ( .A1(\SB4_12/i0_0 ), .A2(\SB4_12/i0_3 ), .A3(\SB4_12/i0[7] ), .ZN(n4515) );
  NAND4_X2 U10814 ( .A1(\SB2_3_30/Component_Function_0/NAND4_in[1] ), .A2(
        n4540), .A3(\SB2_3_30/Component_Function_0/NAND4_in[3] ), .A4(
        \SB2_3_30/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_3_30/buf_output[0] ) );
  NAND4_X2 U10818 ( .A1(\SB1_3_1/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_3_1/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_3_1/Component_Function_0/NAND4_in[0] ), .A4(n4518), .ZN(
        \SB1_3_1/buf_output[0] ) );
  NAND3_X2 U10819 ( .A1(\SB2_0_3/i0[10] ), .A2(\SB2_0_3/i1_5 ), .A3(
        \SB2_0_3/i1[9] ), .ZN(\SB2_0_3/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U10820 ( .A1(\SB4_24/i0_3 ), .A2(\SB4_24/i0[10] ), .A3(
        \SB4_24/i0_4 ), .ZN(\SB4_24/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 U10822 ( .A1(\SB2_1_21/i0[10] ), .A2(\SB2_1_21/i0_3 ), .A3(
        \RI3[1][60] ), .ZN(n4542) );
  NAND4_X2 U10826 ( .A1(\SB2_2_21/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_21/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_21/Component_Function_1/NAND4_in[2] ), .A4(n4520), .ZN(
        \SB2_2_21/buf_output[1] ) );
  NAND3_X2 U10827 ( .A1(\SB2_2_21/i0_4 ), .A2(\SB2_2_21/i1_7 ), .A3(
        \SB2_2_21/i0[8] ), .ZN(n4520) );
  NAND4_X2 U10828 ( .A1(\SB1_2_30/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_2_30/Component_Function_2/NAND4_in[2] ), .A3(
        \SB1_2_30/Component_Function_2/NAND4_in[0] ), .A4(n4521), .ZN(
        \SB1_2_30/buf_output[2] ) );
  XOR2_X1 U10832 ( .A1(\RI5[0][188] ), .A2(\RI5[0][152] ), .Z(n4523) );
  NAND3_X2 U10834 ( .A1(\SB2_3_0/i0[10] ), .A2(\SB2_3_0/i1[9] ), .A3(
        \SB2_3_0/i1_7 ), .ZN(n4680) );
  NAND3_X2 U10837 ( .A1(\SB2_1_0/i0[10] ), .A2(\SB2_1_0/i0_0 ), .A3(
        \SB2_1_0/i0[6] ), .ZN(n968) );
  XOR2_X1 U10838 ( .A1(\MC_ARK_ARC_1_0/temp6[156] ), .A2(n4526), .Z(
        \MC_ARK_ARC_1_0/buf_output[156] ) );
  XOR2_X1 U10839 ( .A1(\MC_ARK_ARC_1_0/temp1[156] ), .A2(
        \MC_ARK_ARC_1_0/temp2[156] ), .Z(n4526) );
  XOR2_X1 U10840 ( .A1(\MC_ARK_ARC_1_2/temp5[190] ), .A2(n4527), .Z(
        \MC_ARK_ARC_1_2/buf_output[190] ) );
  XOR2_X1 U10841 ( .A1(\MC_ARK_ARC_1_2/temp4[190] ), .A2(
        \MC_ARK_ARC_1_2/temp3[190] ), .Z(n4527) );
  XOR2_X1 U10842 ( .A1(\RI5[1][129] ), .A2(\RI5[1][93] ), .Z(n1413) );
  XOR2_X1 U10843 ( .A1(\SB2_2_13/buf_output[3] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[129] ), .Z(\MC_ARK_ARC_1_2/temp1[129] )
         );
  NAND3_X1 U10844 ( .A1(\SB2_3_20/i1[9] ), .A2(\SB2_3_20/i0_4 ), .A3(
        \SB2_3_20/i1_5 ), .ZN(\SB2_3_20/Component_Function_4/NAND4_in[3] ) );
  NAND3_X2 U10845 ( .A1(\SB1_2_13/i0_3 ), .A2(\SB1_2_13/i0[8] ), .A3(
        \SB1_2_13/i0[9] ), .ZN(n827) );
  NAND3_X1 U10848 ( .A1(\SB2_1_10/i0_3 ), .A2(\SB2_1_10/i0[10] ), .A3(
        \SB1_1_11/buf_output[4] ), .ZN(n4528) );
  INV_X1 U10851 ( .I(\SB3_15/buf_output[0] ), .ZN(\SB4_10/i3[0] ) );
  NAND4_X2 U10852 ( .A1(\SB1_2_26/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_2_26/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_26/Component_Function_1/NAND4_in[0] ), .A4(n4531), .ZN(
        \SB1_2_26/buf_output[1] ) );
  XOR2_X1 U10854 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[179] ), .A2(\RI5[3][23] ), 
        .Z(n4532) );
  NAND4_X2 U10855 ( .A1(\SB2_0_6/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_0_6/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_0_6/Component_Function_1/NAND4_in[0] ), .A4(n4533), .ZN(
        \SB2_0_6/buf_output[1] ) );
  NAND2_X2 U10858 ( .A1(n4640), .A2(n970), .ZN(
        \MC_ARK_ARC_1_3/buf_datainput[90] ) );
  NAND4_X2 U10862 ( .A1(\SB2_1_0/Component_Function_0/NAND4_in[1] ), .A2(n1708), .A3(\SB2_1_0/Component_Function_0/NAND4_in[0] ), .A4(n4535), .ZN(
        \SB2_1_0/buf_output[0] ) );
  XOR2_X1 U10864 ( .A1(\MC_ARK_ARC_1_3/temp2[66] ), .A2(
        \MC_ARK_ARC_1_3/temp1[66] ), .Z(n4536) );
  NAND3_X1 U10865 ( .A1(\SB2_1_20/i0_4 ), .A2(\SB2_1_20/i1_7 ), .A3(
        \SB2_1_20/i0[8] ), .ZN(n2060) );
  XOR2_X1 U10866 ( .A1(\MC_ARK_ARC_1_2/temp2[85] ), .A2(n4538), .Z(n585) );
  XOR2_X1 U10867 ( .A1(\RI5[2][79] ), .A2(\RI5[2][85] ), .Z(n4538) );
  NAND3_X2 U10869 ( .A1(\SB1_3_10/i0_3 ), .A2(\SB1_3_10/i0[8] ), .A3(
        \SB1_3_10/i0[9] ), .ZN(n4541) );
  INV_X2 U10870 ( .I(\SB1_2_10/buf_output[3] ), .ZN(\SB2_2_8/i0[8] ) );
  NAND4_X2 U10871 ( .A1(\SB1_2_10/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_10/Component_Function_3/NAND4_in[2] ), .A3(
        \SB1_2_10/Component_Function_3/NAND4_in[1] ), .A4(n1043), .ZN(
        \SB1_2_10/buf_output[3] ) );
  NAND4_X2 U10872 ( .A1(\SB2_1_21/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_21/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_21/Component_Function_4/NAND4_in[3] ), .A4(n4542), .ZN(
        \SB2_1_21/buf_output[4] ) );
  NAND4_X2 U10873 ( .A1(\SB2_1_24/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_1_24/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_24/Component_Function_4/NAND4_in[0] ), .A4(n4543), .ZN(
        \SB2_1_24/buf_output[4] ) );
  NAND3_X1 U10875 ( .A1(\SB2_0_31/i0_0 ), .A2(\SB1_0_0/buf_output[4] ), .A3(
        \SB2_0_31/i1_5 ), .ZN(n4546) );
  NAND4_X2 U10876 ( .A1(\SB1_2_29/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_2_29/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_29/Component_Function_1/NAND4_in[0] ), .A4(n4548), .ZN(
        \SB1_2_29/buf_output[1] ) );
  NAND4_X2 U10877 ( .A1(\SB2_1_19/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_19/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_19/Component_Function_3/NAND4_in[2] ), .A4(n4549), .ZN(
        \SB2_1_19/buf_output[3] ) );
  NAND3_X1 U10878 ( .A1(\SB1_1_21/i0_0 ), .A2(\SB1_1_21/i0_4 ), .A3(
        \SB1_1_21/i0_3 ), .ZN(n4550) );
  NAND3_X1 U10879 ( .A1(\SB3_17/i3[0] ), .A2(\SB3_17/i0[8] ), .A3(
        \SB3_17/i1_5 ), .ZN(n4551) );
  XOR2_X1 U10881 ( .A1(n4553), .A2(\MC_ARK_ARC_1_1/temp5[153] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[153] ) );
  INV_X2 U10883 ( .I(\SB1_1_1/buf_output[3] ), .ZN(\SB2_1_31/i0[8] ) );
  NAND4_X2 U10884 ( .A1(\SB1_1_1/Component_Function_3/NAND4_in[2] ), .A2(
        \SB1_1_1/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_1/Component_Function_3/NAND4_in[0] ), .A4(
        \SB1_1_1/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_1_1/buf_output[3] ) );
  NAND3_X1 U10886 ( .A1(\SB3_17/i0[10] ), .A2(\SB3_17/i1[9] ), .A3(
        \SB3_17/i1_5 ), .ZN(\SB3_17/Component_Function_2/NAND4_in[0] ) );
  INV_X2 U10887 ( .I(n4557), .ZN(\MC_ARK_ARC_1_1/buf_output[110] ) );
  NAND3_X1 U10889 ( .A1(\SB4_9/i0_0 ), .A2(\SB4_9/i3[0] ), .A3(\SB4_9/i1_7 ), 
        .ZN(n4558) );
  NAND3_X1 U10890 ( .A1(\SB4_24/i0_3 ), .A2(\SB4_24/i1[9] ), .A3(\SB4_24/i0_4 ), .ZN(\SB4_24/Component_Function_5/NAND4_in[2] ) );
  NAND2_X2 U10892 ( .A1(\SB2_3_22/i0_0 ), .A2(\SB2_3_22/i3[0] ), .ZN(n4560) );
  NAND3_X1 U10893 ( .A1(\SB3_5/i0[8] ), .A2(\SB3_5/i0_3 ), .A3(\SB3_5/i1_7 ), 
        .ZN(\SB3_5/Component_Function_1/NAND4_in[1] ) );
  INV_X2 U10896 ( .I(\SB3_2/buf_output[2] ), .ZN(\SB4_31/i1[9] ) );
  NAND3_X2 U10899 ( .A1(\SB2_1_17/i0_3 ), .A2(\SB2_1_17/i0_4 ), .A3(
        \SB2_1_17/i1[9] ), .ZN(n1211) );
  NAND3_X1 U10900 ( .A1(\SB4_7/i0_0 ), .A2(\SB4_7/i0[9] ), .A3(\SB4_7/i0[8] ), 
        .ZN(n4567) );
  XOR2_X1 U10902 ( .A1(\MC_ARK_ARC_1_2/temp3[153] ), .A2(
        \MC_ARK_ARC_1_2/temp4[153] ), .Z(n4569) );
  XOR2_X1 U10903 ( .A1(n4570), .A2(\MC_ARK_ARC_1_0/temp4[34] ), .Z(n2669) );
  XOR2_X1 U10904 ( .A1(\RI5[0][100] ), .A2(\RI5[0][136] ), .Z(n4570) );
  XOR2_X1 U10905 ( .A1(\MC_ARK_ARC_1_2/temp1[128] ), .A2(
        \MC_ARK_ARC_1_2/temp2[128] ), .Z(n2106) );
  XOR2_X1 U10906 ( .A1(n1544), .A2(n4572), .Z(\MC_ARK_ARC_1_1/buf_output[13] )
         );
  XOR2_X1 U10907 ( .A1(\MC_ARK_ARC_1_1/temp3[13] ), .A2(
        \MC_ARK_ARC_1_1/temp2[13] ), .Z(n4572) );
  NAND4_X2 U10908 ( .A1(\SB1_1_23/Component_Function_3/NAND4_in[2] ), .A2(
        \SB1_1_23/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_23/Component_Function_3/NAND4_in[0] ), .A4(n4573), .ZN(
        \SB1_1_23/buf_output[3] ) );
  NAND3_X1 U10909 ( .A1(\SB1_2_26/i1_5 ), .A2(\SB1_2_26/i0[9] ), .A3(
        \SB1_2_26/i0[6] ), .ZN(\SB1_2_26/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 U10910 ( .A1(\SB2_1_17/i0[10] ), .A2(\SB2_1_17/i1_7 ), .A3(
        \SB2_1_17/i1[9] ), .ZN(n2115) );
  XOR2_X1 U10912 ( .A1(\RI5[0][28] ), .A2(\RI5[0][52] ), .Z(n4575) );
  XOR2_X1 U10913 ( .A1(\MC_ARK_ARC_1_1/temp3[162] ), .A2(
        \MC_ARK_ARC_1_1/temp4[162] ), .Z(\MC_ARK_ARC_1_1/temp6[162] ) );
  NAND2_X1 U10914 ( .A1(\SB2_1_15/i0[9] ), .A2(\SB2_1_15/i0[10] ), .ZN(
        \SB2_1_15/Component_Function_0/NAND4_in[0] ) );
  XOR2_X1 U10917 ( .A1(\MC_ARK_ARC_1_1/temp3[184] ), .A2(
        \MC_ARK_ARC_1_1/temp4[184] ), .Z(n1298) );
  NAND3_X1 U10918 ( .A1(\SB4_22/i0[8] ), .A2(\SB4_22/i3[0] ), .A3(
        \SB4_22/i1_5 ), .ZN(n4579) );
  XOR2_X1 U10919 ( .A1(\RI5[2][159] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[183] ), .Z(n4581) );
  XOR2_X1 U10921 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[105] ), .A2(\RI5[1][129] ), .Z(\MC_ARK_ARC_1_1/temp2[159] ) );
  NAND4_X2 U10922 ( .A1(\SB1_3_10/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_3_10/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_3_10/Component_Function_1/NAND4_in[0] ), .A4(n4583), .ZN(
        \SB1_3_10/buf_output[1] ) );
  XOR2_X1 U10923 ( .A1(n2565), .A2(n4584), .Z(\MC_ARK_ARC_1_1/buf_output[93] )
         );
  NAND3_X1 U10927 ( .A1(\SB4_13/i0[10] ), .A2(\SB4_13/i0_0 ), .A3(
        \SB4_13/i0[6] ), .ZN(\SB4_13/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U10929 ( .A1(\RI5[1][174] ), .A2(\RI5[1][180] ), .Z(n4586) );
  XOR2_X1 U10930 ( .A1(\RI5[0][159] ), .A2(\RI5[0][183] ), .Z(
        \MC_ARK_ARC_1_0/temp2[21] ) );
  NAND3_X1 U10932 ( .A1(\SB1_3_13/i0_0 ), .A2(\SB1_3_13/i3[0] ), .A3(
        \SB1_3_13/i1_7 ), .ZN(\SB1_3_13/Component_Function_4/NAND4_in[1] ) );
  NAND4_X2 U10934 ( .A1(\SB1_2_8/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_2_8/Component_Function_1/NAND4_in[0] ), .A3(n4674), .A4(n4589), 
        .ZN(\SB1_2_8/buf_output[1] ) );
  NAND4_X2 U10935 ( .A1(\SB1_0_11/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_0_11/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_0_11/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_0_11/Component_Function_1/NAND4_in[0] ), .ZN(\SB2_0_7/i0[6] ) );
  INV_X1 U10936 ( .I(\SB1_1_8/buf_output[0] ), .ZN(\SB2_1_3/i3[0] ) );
  NAND4_X2 U10937 ( .A1(\SB1_1_8/Component_Function_0/NAND4_in[3] ), .A2(n1313), .A3(\SB1_1_8/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_1_8/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_1_8/buf_output[0] ) );
  XOR2_X1 U10941 ( .A1(\MC_ARK_ARC_1_3/temp5[159] ), .A2(n4593), .Z(
        \MC_ARK_ARC_1_3/buf_output[159] ) );
  XOR2_X1 U10942 ( .A1(\MC_ARK_ARC_1_3/temp4[159] ), .A2(
        \MC_ARK_ARC_1_3/temp3[159] ), .Z(n4593) );
  NAND3_X2 U10950 ( .A1(\SB2_1_10/i0_3 ), .A2(\SB1_1_11/buf_output[4] ), .A3(
        \SB2_1_10/i1[9] ), .ZN(n4720) );
  XOR2_X1 U10951 ( .A1(\RI5[2][111] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[117] ), .Z(n1230) );
  XOR2_X1 U10958 ( .A1(\MC_ARK_ARC_1_3/temp2[120] ), .A2(n4603), .Z(
        \MC_ARK_ARC_1_3/temp5[120] ) );
  XOR2_X1 U10959 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[114] ), .A2(\RI5[3][120] ), .Z(n4603) );
  NAND3_X1 U10960 ( .A1(\SB4_10/i0[9] ), .A2(\SB4_10/i0_4 ), .A3(
        \SB4_10/i0[6] ), .ZN(n4604) );
  NAND3_X1 U10961 ( .A1(\SB4_15/i0_3 ), .A2(\SB4_15/i0[6] ), .A3(
        \SB4_15/i1[9] ), .ZN(n4605) );
  XOR2_X1 U10964 ( .A1(n4607), .A2(n173), .Z(Ciphertext[101]) );
  NAND4_X2 U10965 ( .A1(\SB4_15/Component_Function_5/NAND4_in[1] ), .A2(
        \SB4_15/Component_Function_5/NAND4_in[2] ), .A3(
        \SB4_15/Component_Function_5/NAND4_in[3] ), .A4(
        \SB4_15/Component_Function_5/NAND4_in[0] ), .ZN(n4607) );
  NAND4_X2 U10967 ( .A1(n1724), .A2(
        \SB2_0_25/Component_Function_0/NAND4_in[1] ), .A3(n1788), .A4(
        \SB2_0_25/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_0_25/buf_output[0] ) );
  NAND4_X2 U10970 ( .A1(\SB1_0_29/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_0_29/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_0_29/Component_Function_1/NAND4_in[0] ), .A4(n4608), .ZN(
        \SB1_0_29/buf_output[1] ) );
  NAND3_X1 U10971 ( .A1(\SB1_0_29/i1_7 ), .A2(\SB1_0_29/i0[8] ), .A3(n346), 
        .ZN(n4608) );
  XOR2_X1 U10972 ( .A1(n4609), .A2(n1690), .Z(\MC_ARK_ARC_1_0/temp5[186] ) );
  XOR2_X1 U10973 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[180] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[132] ), .Z(n4609) );
  INV_X2 U10976 ( .I(\SB1_1_18/buf_output[2] ), .ZN(\SB2_1_15/i1[9] ) );
  INV_X2 U10978 ( .I(\RI3[0][81] ), .ZN(\SB2_0_18/i0[8] ) );
  XOR2_X1 U10981 ( .A1(\MC_ARK_ARC_1_3/temp1[145] ), .A2(n4613), .Z(
        \MC_ARK_ARC_1_3/temp5[145] ) );
  XOR2_X1 U10982 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[115] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[91] ), .Z(n4613) );
  INV_X1 U10983 ( .I(\SB3_7/buf_output[5] ), .ZN(\SB4_7/i1_5 ) );
  NAND3_X1 U10985 ( .A1(\SB1_3_19/buf_output[1] ), .A2(n809), .A3(
        \SB1_3_17/buf_output[3] ), .ZN(
        \SB2_3_15/Component_Function_5/NAND4_in[1] ) );
  AND2_X1 U10987 ( .A1(\SB2_3_21/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_3_21/Component_Function_0/NAND4_in[0] ), .Z(n4640) );
  XOR2_X1 U10989 ( .A1(\RI5[0][3] ), .A2(\RI5[0][27] ), .Z(n4619) );
  XOR2_X1 U10990 ( .A1(n4620), .A2(n223), .Z(Ciphertext[97]) );
  XOR2_X1 U10992 ( .A1(\RI5[1][152] ), .A2(\RI5[1][188] ), .Z(
        \MC_ARK_ARC_1_1/temp3[86] ) );
  XOR2_X1 U10994 ( .A1(\MC_ARK_ARC_1_1/temp2[182] ), .A2(
        \MC_ARK_ARC_1_1/temp1[182] ), .Z(n4622) );
  XOR2_X1 U10995 ( .A1(n4623), .A2(\MC_ARK_ARC_1_2/temp5[34] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[34] ) );
  XOR2_X1 U10996 ( .A1(\MC_ARK_ARC_1_2/temp3[34] ), .A2(
        \MC_ARK_ARC_1_2/temp4[34] ), .Z(n4623) );
  NAND3_X1 U10997 ( .A1(\SB2_0_2/i0[8] ), .A2(\RI3[0][178] ), .A3(
        \SB2_0_2/i1_7 ), .ZN(\SB2_0_2/Component_Function_1/NAND4_in[3] ) );
  XOR2_X1 U10998 ( .A1(\RI5[0][173] ), .A2(\RI5[0][5] ), .Z(n4624) );
  XOR2_X1 U11003 ( .A1(\MC_ARK_ARC_1_0/temp3[89] ), .A2(
        \MC_ARK_ARC_1_0/temp4[89] ), .Z(n4627) );
  XOR2_X1 U11005 ( .A1(\MC_ARK_ARC_1_0/temp2[160] ), .A2(n4630), .Z(
        \MC_ARK_ARC_1_0/temp5[160] ) );
  XOR2_X1 U11006 ( .A1(\RI5[0][160] ), .A2(\RI5[0][154] ), .Z(n4630) );
  NAND3_X2 U11010 ( .A1(\SB2_1_21/i0_4 ), .A2(\SB2_1_21/i1_5 ), .A3(
        \SB2_1_21/i0_0 ), .ZN(n711) );
  NAND4_X2 U11013 ( .A1(\SB1_1_28/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_1_28/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_1_28/Component_Function_1/NAND4_in[3] ), .A4(
        \SB1_1_28/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_1_28/buf_output[1] ) );
  NAND3_X2 U11014 ( .A1(\SB1_2_13/i0_0 ), .A2(\SB1_2_13/i0[10] ), .A3(
        \SB1_2_13/i0[6] ), .ZN(n1523) );
  NAND3_X1 U11015 ( .A1(\SB3_2/i0[9] ), .A2(\SB3_2/i0[8] ), .A3(\SB3_2/i0_0 ), 
        .ZN(\SB3_2/Component_Function_4/NAND4_in[0] ) );
  NAND3_X2 U11017 ( .A1(\SB1_1_15/i0[10] ), .A2(\SB1_1_15/i1[9] ), .A3(
        \SB1_1_15/i1_7 ), .ZN(\SB1_1_15/Component_Function_3/NAND4_in[2] ) );
  INV_X2 U11020 ( .I(\SB1_2_22/buf_output[2] ), .ZN(\SB2_2_19/i1[9] ) );
  NAND3_X1 U11022 ( .A1(\SB2_2_26/i0_0 ), .A2(\SB2_2_26/i0[9] ), .A3(
        \SB2_2_26/i0[8] ), .ZN(\SB2_2_26/Component_Function_4/NAND4_in[0] ) );
  XOR2_X1 U11023 ( .A1(\MC_ARK_ARC_1_2/temp1[134] ), .A2(
        \MC_ARK_ARC_1_2/temp4[134] ), .Z(n4635) );
  XOR2_X1 U11024 ( .A1(\MC_ARK_ARC_1_2/temp3[134] ), .A2(n1993), .Z(n4636) );
  NAND4_X2 U11026 ( .A1(\SB2_3_9/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_3_9/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_3_9/Component_Function_4/NAND4_in[0] ), .A4(n4637), .ZN(
        \SB2_3_9/buf_output[4] ) );
  NAND3_X1 U11028 ( .A1(\SB2_3_10/i0_3 ), .A2(\SB2_3_10/i0[10] ), .A3(
        \SB2_3_10/i0_4 ), .ZN(\SB2_3_10/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 U11029 ( .A1(\SB2_1_21/i0_4 ), .A2(\SB2_1_21/i0[10] ), .A3(
        \SB2_1_21/i0_3 ), .ZN(n4697) );
  XOR2_X1 U11030 ( .A1(n4639), .A2(n2333), .Z(\MC_ARK_ARC_1_2/buf_output[130] ) );
  NOR2_X2 U11032 ( .A1(n1144), .A2(n4641), .ZN(\SB2_0_9/i0[7] ) );
  NAND4_X2 U11033 ( .A1(\SB4_24/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_24/Component_Function_0/NAND4_in[1] ), .A3(
        \SB4_24/Component_Function_0/NAND4_in[0] ), .A4(n4642), .ZN(n2280) );
  NAND3_X1 U11034 ( .A1(\SB3_24/buf_output[2] ), .A2(\SB4_21/i0[8] ), .A3(
        \SB4_21/i0[9] ), .ZN(n4643) );
  XOR2_X1 U11036 ( .A1(\RI5[3][68] ), .A2(\RI5[3][62] ), .Z(n4645) );
  NAND3_X1 U11037 ( .A1(\SB2_1_13/i0_0 ), .A2(\SB2_1_13/i0_3 ), .A3(
        \SB2_1_13/i0[7] ), .ZN(n2017) );
  NAND3_X2 U11039 ( .A1(\SB1_1_10/i0_3 ), .A2(\SB1_1_10/i1[9] ), .A3(
        \SB1_1_10/i0_4 ), .ZN(n858) );
  XOR2_X1 U11040 ( .A1(n4647), .A2(n4648), .Z(\MC_ARK_ARC_1_1/temp5[154] ) );
  XOR2_X1 U11041 ( .A1(\RI5[1][148] ), .A2(\RI5[1][154] ), .Z(n4647) );
  XOR2_X1 U11042 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[100] ), .A2(\RI5[1][124] ), .Z(n4648) );
  NAND3_X2 U11043 ( .A1(\SB2_0_2/i1[9] ), .A2(\SB2_0_2/i1_7 ), .A3(
        \SB2_0_2/i0[10] ), .ZN(n4655) );
  NAND3_X1 U11045 ( .A1(\SB1_0_21/i0_0 ), .A2(\SB1_0_21/i0_4 ), .A3(
        \SB1_0_21/i1_5 ), .ZN(n4650) );
  NAND3_X2 U11046 ( .A1(\SB2_1_31/i0[9] ), .A2(\SB2_1_31/i0[6] ), .A3(
        \SB2_1_31/i0_4 ), .ZN(\SB2_1_31/Component_Function_5/NAND4_in[3] ) );
  INV_X1 U11047 ( .I(\SB3_8/buf_output[5] ), .ZN(\SB4_8/i1_5 ) );
  NAND4_X2 U11048 ( .A1(\SB3_8/Component_Function_5/NAND4_in[1] ), .A2(n2889), 
        .A3(\SB3_8/Component_Function_5/NAND4_in[3] ), .A4(
        \SB3_8/Component_Function_5/NAND4_in[0] ), .ZN(\SB3_8/buf_output[5] )
         );
  NAND4_X2 U11049 ( .A1(\SB1_1_4/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_1_4/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_1_4/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_1_4/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_1_4/buf_output[0] ) );
  INV_X1 U11050 ( .I(\SB1_2_11/buf_output[1] ), .ZN(\SB2_2_7/i1_7 ) );
  XOR2_X1 U11053 ( .A1(n4654), .A2(\MC_ARK_ARC_1_1/temp5[121] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[121] ) );
  XOR2_X1 U11056 ( .A1(n2815), .A2(n4656), .Z(\MC_ARK_ARC_1_0/buf_output[51] )
         );
  XOR2_X1 U11059 ( .A1(n4658), .A2(\MC_ARK_ARC_1_3/temp6[138] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[138] ) );
  NAND4_X2 U11064 ( .A1(\SB3_7/Component_Function_3/NAND4_in[1] ), .A2(
        \SB3_7/Component_Function_3/NAND4_in[0] ), .A3(n1836), .A4(n4660), 
        .ZN(\SB3_7/buf_output[3] ) );
  NAND3_X2 U11065 ( .A1(\SB2_2_17/i0[10] ), .A2(\SB2_2_17/i0[6] ), .A3(
        \SB2_2_17/i0_0 ), .ZN(n4661) );
  NAND4_X2 U11067 ( .A1(\SB2_0_18/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_0_18/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_0_18/Component_Function_3/NAND4_in[3] ), .A4(n4663), .ZN(
        \SB2_0_18/buf_output[3] ) );
  XOR2_X1 U11068 ( .A1(\MC_ARK_ARC_1_3/temp2[61] ), .A2(
        \MC_ARK_ARC_1_3/temp1[61] ), .Z(\MC_ARK_ARC_1_3/temp5[61] ) );
  XOR2_X1 U11070 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[92] ), .A2(\RI5[0][68] ), 
        .Z(n4665) );
  INV_X2 U11071 ( .I(\SB1_0_11/buf_output[2] ), .ZN(\SB2_0_8/i1[9] ) );
  NAND3_X2 U11074 ( .A1(\SB2_3_8/i3[0] ), .A2(\SB2_3_8/i0[8] ), .A3(
        \SB2_3_8/i1_5 ), .ZN(n4728) );
  NAND4_X2 U11079 ( .A1(\SB1_2_2/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_2_2/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_2_2/Component_Function_1/NAND4_in[0] ), .A4(n4670), .ZN(
        \SB1_2_2/buf_output[1] ) );
  NAND3_X1 U11080 ( .A1(\SB3_27/i0_0 ), .A2(\SB3_27/i3[0] ), .A3(\SB3_27/i1_7 ), .ZN(\SB3_27/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U11083 ( .A1(\SB1_3_17/i0[6] ), .A2(\SB1_3_17/i0[9] ), .A3(
        \SB1_3_17/i1_5 ), .ZN(\SB1_3_17/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 U11085 ( .A1(\SB2_0_13/i0_0 ), .A2(n3663), .A3(\SB2_0_13/i0_4 ), 
        .ZN(n4672) );
  XOR2_X1 U11088 ( .A1(\RI5[2][66] ), .A2(\RI5[2][72] ), .Z(
        \MC_ARK_ARC_1_2/temp1[72] ) );
  NOR2_X2 U11089 ( .A1(n1053), .A2(n4675), .ZN(n2738) );
  NAND4_X2 U11090 ( .A1(\SB2_2_10/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_2_10/Component_Function_0/NAND4_in[0] ), .A3(
        \SB2_2_10/Component_Function_0/NAND4_in[2] ), .A4(n4676), .ZN(
        \SB2_2_10/buf_output[0] ) );
  NAND3_X1 U11091 ( .A1(n3680), .A2(\RI3[3][24] ), .A3(\SB2_3_27/i1_5 ), .ZN(
        \SB2_3_27/Component_Function_1/NAND4_in[2] ) );
  XOR2_X1 U11095 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[58] ), .A2(\RI5[2][22] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[148] ) );
  NAND4_X2 U11096 ( .A1(\SB2_3_0/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_3_0/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_3_0/Component_Function_3/NAND4_in[3] ), .A4(n4680), .ZN(
        \SB2_3_0/buf_output[3] ) );
  NAND3_X1 U11097 ( .A1(\SB2_2_26/i0[8] ), .A2(\SB2_2_26/i3[0] ), .A3(
        \SB2_2_26/i1_5 ), .ZN(\SB2_2_26/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U11100 ( .A1(n4683), .A2(\MC_ARK_ARC_1_1/temp5[168] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[168] ) );
  XOR2_X1 U11101 ( .A1(\MC_ARK_ARC_1_1/temp4[168] ), .A2(
        \MC_ARK_ARC_1_1/temp3[168] ), .Z(n4683) );
  NAND4_X2 U11103 ( .A1(\SB1_0_17/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_17/Component_Function_3/NAND4_in[2] ), .A3(
        \SB1_0_17/Component_Function_3/NAND4_in[3] ), .A4(n4685), .ZN(
        \RI3[0][99] ) );
  NAND3_X1 U11105 ( .A1(\SB4_28/i0[10] ), .A2(\SB4_28/i0_0 ), .A3(
        \SB4_28/i0[6] ), .ZN(\SB4_28/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U11106 ( .A1(n570), .A2(\RI5[2][170] ), .Z(n4687) );
  XOR2_X1 U11109 ( .A1(\RI5[1][64] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[28] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[154] ) );
  XOR2_X1 U11116 ( .A1(n4693), .A2(n7), .Z(Ciphertext[43]) );
  NAND4_X2 U11117 ( .A1(\SB4_24/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_24/Component_Function_1/NAND4_in[3] ), .A3(
        \SB4_24/Component_Function_1/NAND4_in[0] ), .A4(
        \SB4_24/Component_Function_1/NAND4_in[2] ), .ZN(n4693) );
  NAND3_X1 U11118 ( .A1(\SB2_1_2/i0_3 ), .A2(\SB2_1_2/i0[10] ), .A3(
        \SB2_1_2/i0[9] ), .ZN(\SB2_1_2/Component_Function_4/NAND4_in[2] ) );
  XOR2_X1 U11119 ( .A1(\MC_ARK_ARC_1_1/temp2[42] ), .A2(
        \MC_ARK_ARC_1_1/temp1[42] ), .Z(\MC_ARK_ARC_1_1/temp5[42] ) );
  NAND4_X2 U11120 ( .A1(\SB2_3_18/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_18/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_3_18/Component_Function_4/NAND4_in[2] ), .A4(n4694), .ZN(
        \SB2_3_18/buf_output[4] ) );
  INV_X2 U11122 ( .I(\SB1_3_27/buf_output[2] ), .ZN(\SB2_3_24/i1[9] ) );
  NAND4_X2 U11123 ( .A1(\SB1_0_8/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_0_8/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_0_8/Component_Function_1/NAND4_in[0] ), .A4(
        \SB1_0_8/Component_Function_1/NAND4_in[2] ), .ZN(\RI3[0][163] ) );
  NAND3_X2 U11124 ( .A1(\SB2_1_21/i0_4 ), .A2(\SB2_1_21/i0_3 ), .A3(
        \SB2_1_21/i0_0 ), .ZN(n4748) );
  XOR2_X1 U11125 ( .A1(\MC_ARK_ARC_1_0/temp1[161] ), .A2(
        \MC_ARK_ARC_1_0/temp3[161] ), .Z(n763) );
  NOR2_X2 U11128 ( .A1(n1014), .A2(n4698), .ZN(n2563) );
  XOR2_X1 U11131 ( .A1(n1536), .A2(\MC_ARK_ARC_1_1/temp4[13] ), .Z(n1544) );
  XOR2_X1 U11134 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[50] ), .A2(n3677), .Z(
        \MC_ARK_ARC_1_2/temp2[80] ) );
  NAND3_X2 U11137 ( .A1(\SB1_2_26/i1_5 ), .A2(\SB1_2_26/i0_4 ), .A3(
        \SB1_2_26/i0_0 ), .ZN(n4704) );
  NAND4_X2 U11138 ( .A1(n2858), .A2(n1616), .A3(
        \SB2_2_6/Component_Function_2/NAND4_in[2] ), .A4(n4705), .ZN(
        \SB2_2_6/buf_output[2] ) );
  XOR2_X1 U11139 ( .A1(n4706), .A2(n6), .Z(Ciphertext[113]) );
  NAND4_X2 U11140 ( .A1(\SB4_13/Component_Function_5/NAND4_in[2] ), .A2(
        \SB4_13/Component_Function_5/NAND4_in[1] ), .A3(
        \SB4_13/Component_Function_5/NAND4_in[0] ), .A4(
        \SB4_13/Component_Function_5/NAND4_in[3] ), .ZN(n4706) );
  XOR2_X1 U11141 ( .A1(n4707), .A2(n141), .Z(Ciphertext[162]) );
  NAND4_X2 U11142 ( .A1(\SB4_4/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_4/Component_Function_0/NAND4_in[1] ), .A3(
        \SB4_4/Component_Function_0/NAND4_in[3] ), .A4(
        \SB4_4/Component_Function_0/NAND4_in[0] ), .ZN(n4707) );
  NAND4_X2 U11143 ( .A1(\SB2_1_21/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_1_21/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_21/Component_Function_1/NAND4_in[0] ), .A4(n4709), .ZN(
        \SB2_1_21/buf_output[1] ) );
  XOR2_X1 U11144 ( .A1(\MC_ARK_ARC_1_0/temp5[186] ), .A2(n1850), .Z(
        \MC_ARK_ARC_1_0/buf_output[186] ) );
  NAND3_X1 U11145 ( .A1(\SB1_2_9/i0_4 ), .A2(\SB1_2_9/i1_7 ), .A3(
        \SB1_2_9/i0[8] ), .ZN(n4710) );
  NAND4_X2 U11147 ( .A1(\SB2_1_2/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_1_2/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_1_2/Component_Function_3/NAND4_in[3] ), .A4(n1317), .ZN(
        \SB2_1_2/buf_output[3] ) );
  NAND4_X2 U11152 ( .A1(\SB1_1_5/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_5/Component_Function_5/NAND4_in[3] ), .A3(n4745), .A4(
        \SB1_1_5/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_5/buf_output[5] ) );
  NAND3_X1 U11154 ( .A1(\SB1_2_26/i0[8] ), .A2(\RI1[2][35] ), .A3(
        \SB1_2_26/i1_7 ), .ZN(\SB1_2_26/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U11156 ( .A1(\RI5[1][131] ), .A2(\RI5[1][167] ), .Z(
        \MC_ARK_ARC_1_1/temp3[65] ) );
  NAND4_X2 U11157 ( .A1(\SB1_2_26/Component_Function_4/NAND4_in[0] ), .A2(
        n1717), .A3(\SB1_2_26/Component_Function_4/NAND4_in[1] ), .A4(n4714), 
        .ZN(\SB1_2_26/buf_output[4] ) );
  NAND3_X2 U11159 ( .A1(\SB2_3_22/i0[10] ), .A2(\SB2_3_22/i0_0 ), .A3(
        \SB2_3_22/i0[6] ), .ZN(n4715) );
  NAND3_X1 U11160 ( .A1(\SB1_3_28/i1[9] ), .A2(\SB1_3_28/i0[10] ), .A3(
        \SB1_3_28/i1_5 ), .ZN(\SB1_3_28/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U11161 ( .A1(\SB2_3_7/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_7/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_3_7/Component_Function_5/NAND4_in[0] ), .A4(n4717), .ZN(
        \SB2_3_7/buf_output[5] ) );
  NAND4_X2 U11162 ( .A1(\SB1_1_7/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_1_7/Component_Function_3/NAND4_in[2] ), .A3(
        \SB1_1_7/Component_Function_3/NAND4_in[0] ), .A4(n4718), .ZN(
        \SB1_1_7/buf_output[3] ) );
  AND2_X1 U11163 ( .A1(n2510), .A2(n4719), .Z(n2282) );
  NAND3_X2 U11166 ( .A1(\SB1_1_13/i0[10] ), .A2(\SB1_1_13/i0_0 ), .A3(
        \SB1_1_13/i0[6] ), .ZN(\SB1_1_13/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U11168 ( .A1(n4722), .A2(n2021), .Z(\MC_ARK_ARC_1_1/temp5[177] ) );
  XOR2_X1 U11169 ( .A1(\RI5[1][171] ), .A2(\RI5[1][177] ), .Z(n4722) );
  INV_X2 U11170 ( .I(\SB1_2_2/buf_output[2] ), .ZN(\SB2_2_31/i1[9] ) );
  NAND3_X2 U11174 ( .A1(\SB2_3_23/i0[9] ), .A2(\SB2_3_23/i0_4 ), .A3(
        \SB2_3_23/i0[6] ), .ZN(n4725) );
  XOR2_X1 U11175 ( .A1(\MC_ARK_ARC_1_1/temp6[185] ), .A2(
        \MC_ARK_ARC_1_1/temp5[185] ), .Z(\MC_ARK_ARC_1_1/buf_output[185] ) );
  XOR2_X1 U11177 ( .A1(\MC_ARK_ARC_1_2/temp3[117] ), .A2(
        \MC_ARK_ARC_1_2/temp4[117] ), .Z(n4726) );
  XOR2_X1 U11191 ( .A1(\RI5[2][184] ), .A2(\RI5[2][16] ), .Z(n4733) );
  NAND3_X2 U11192 ( .A1(\SB1_1_4/i0[10] ), .A2(\SB1_1_4/i1[9] ), .A3(
        \SB1_1_4/i1_7 ), .ZN(n4734) );
  NAND4_X2 U11195 ( .A1(\SB1_2_30/Component_Function_0/NAND4_in[0] ), .A2(
        \SB1_2_30/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_2_30/Component_Function_0/NAND4_in[1] ), .A4(n4736), .ZN(
        \SB1_2_30/buf_output[0] ) );
  NAND3_X2 U11196 ( .A1(\SB2_1_2/i0_3 ), .A2(\SB2_1_2/i1_7 ), .A3(
        \SB2_1_2/i0[8] ), .ZN(n1851) );
  XOR2_X1 U11201 ( .A1(\MC_ARK_ARC_1_3/temp3[110] ), .A2(
        \MC_ARK_ARC_1_3/temp1[110] ), .Z(n4740) );
  NAND3_X1 U11202 ( .A1(\SB1_1_20/i0_3 ), .A2(\SB1_1_20/i0[6] ), .A3(
        \SB1_1_20/i0[10] ), .ZN(\SB1_1_20/Component_Function_2/NAND4_in[1] )
         );
  NAND3_X1 U11205 ( .A1(\SB4_26/i0_4 ), .A2(\SB4_26/i1[9] ), .A3(\SB4_26/i1_5 ), .ZN(n4742) );
  XOR2_X1 U11206 ( .A1(\MC_ARK_ARC_1_2/temp3[159] ), .A2(
        \MC_ARK_ARC_1_2/temp4[159] ), .Z(n4743) );
  NAND3_X2 U11208 ( .A1(\SB1_1_1/i0[6] ), .A2(\SB1_1_1/i0[9] ), .A3(
        \SB1_1_1/i0_4 ), .ZN(n4744) );
  NAND3_X2 U11209 ( .A1(\SB2_0_11/i0_0 ), .A2(\SB2_0_11/i0[10] ), .A3(
        \SB2_0_11/i0[6] ), .ZN(\SB2_0_11/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U11210 ( .A1(\SB1_1_5/i0_3 ), .A2(\SB1_1_5/i1[9] ), .A3(
        \SB1_1_5/i0_4 ), .ZN(n4745) );
  NAND4_X2 U11213 ( .A1(\SB1_2_13/Component_Function_3/NAND4_in[1] ), .A2(
        n2122), .A3(n2763), .A4(\SB1_2_13/Component_Function_3/NAND4_in[3] ), 
        .ZN(n4749) );
  AND4_X2 U11215 ( .A1(\SB1_3_28/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_3_28/Component_Function_3/NAND4_in[0] ), .A3(n2316), .A4(
        \SB1_3_28/Component_Function_3/NAND4_in[3] ), .Z(n4750) );
  BUF_X4 \SB2_0_31/BUF_3  ( .I(\RI3[0][3] ), .Z(\SB2_0_31/i0[10] ) );
  NAND3_X2 U4329 ( .A1(\SB2_1_25/i0_3 ), .A2(\SB2_1_25/i0_0 ), .A3(n1579), 
        .ZN(n2067) );
  INV_X2 \SB3_23/INV_2  ( .I(n1401), .ZN(\SB3_23/i1[9] ) );
  NAND3_X2 \SB1_1_28/Component_Function_2/N2  ( .A1(\SB1_1_28/i0_3 ), .A2(
        \SB1_1_28/i0[10] ), .A3(\SB1_1_28/i0[6] ), .ZN(
        \SB1_1_28/Component_Function_2/NAND4_in[1] ) );
  INV_X2 U952 ( .I(\MC_ARK_ARC_1_2/buf_output[26] ), .ZN(\SB1_3_27/i1[9] ) );
  INV_X2 U2715 ( .I(\MC_ARK_ARC_1_2/buf_output[65] ), .ZN(\SB1_3_21/i1_5 ) );
  BUF_X4 \SB2_2_15/BUF_0  ( .I(\SB1_2_20/buf_output[0] ), .Z(\SB2_2_15/i0[9] )
         );
  INV_X2 U8494 ( .I(\SB1_2_30/buf_output[5] ), .ZN(\SB2_2_30/i1_5 ) );
  INV_X2 U647 ( .I(\MC_ARK_ARC_1_3/buf_output[17] ), .ZN(\SB3_29/i1_5 ) );
  NAND3_X2 U2545 ( .A1(\SB1_3_9/i0[8] ), .A2(\SB1_3_9/i0[9] ), .A3(
        \SB1_3_9/i0_3 ), .ZN(n4106) );
  NAND4_X2 U5492 ( .A1(\SB2_2_1/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_2_1/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_1/Component_Function_1/NAND4_in[0] ), .A4(n1649), .ZN(
        \SB2_2_1/buf_output[1] ) );
  NAND2_X2 \SB1_2_1/Component_Function_5/N1  ( .A1(\SB1_2_1/i0_0 ), .A2(
        \SB1_2_1/i3[0] ), .ZN(\SB1_2_1/Component_Function_5/NAND4_in[0] ) );
  NAND4_X1 \SB2_0_29/Component_Function_1/N5  ( .A1(
        \SB2_0_29/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_0_29/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_29/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_29/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_0_29/buf_output[1] ) );
  NAND3_X2 U927 ( .A1(\SB1_3_9/i0_0 ), .A2(\SB1_3_9/i0_3 ), .A3(\SB1_3_9/i0_4 ), .ZN(\SB1_3_9/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 \SB3_29/Component_Function_3/N1  ( .A1(\SB3_29/i1[9] ), .A2(
        \SB3_29/i0_3 ), .A3(\SB3_29/i0[6] ), .ZN(
        \SB3_29/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U1302 ( .A1(\SB2_1_14/i0[10] ), .A2(\SB2_1_14/i1_7 ), .A3(
        \SB2_1_14/i1[9] ), .ZN(\SB2_1_14/Component_Function_3/NAND4_in[2] ) );
  BUF_X4 \SB1_3_29/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[16] ), .Z(
        \SB1_3_29/i0_4 ) );
  NAND3_X2 U6583 ( .A1(\SB2_2_25/i0_4 ), .A2(\SB2_2_25/i0[9] ), .A3(
        \SB2_2_25/i0[6] ), .ZN(n2145) );
  INV_X2 U2355 ( .I(\MC_ARK_ARC_1_0/buf_output[86] ), .ZN(\SB1_1_17/i1[9] ) );
  BUF_X2 U2120 ( .I(\MC_ARK_ARC_1_2/buf_output[12] ), .Z(\SB1_3_29/i0[9] ) );
  NAND3_X2 U1444 ( .A1(\SB1_1_7/i0_3 ), .A2(\SB1_1_7/i0_4 ), .A3(
        \SB1_1_7/i1[9] ), .ZN(\SB1_1_7/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 \SB2_1_7/Component_Function_2/N3  ( .A1(\SB2_1_7/i0_3 ), .A2(
        \SB2_1_7/i0[8] ), .A3(\SB2_1_7/i0[9] ), .ZN(
        \SB2_1_7/Component_Function_2/NAND4_in[2] ) );
  INV_X4 U5099 ( .I(\SB2_1_10/i0[7] ), .ZN(\SB1_1_11/buf_output[4] ) );
  NAND2_X2 U1008 ( .A1(\SB1_1_11/Component_Function_4/NAND4_in[3] ), .A2(n1562), .ZN(n1463) );
  INV_X2 U1634 ( .I(n383), .ZN(\SB1_0_10/i0[8] ) );
  BUF_X4 U1664 ( .I(\MC_ARK_ARC_1_2/buf_output[74] ), .Z(\SB1_3_19/i0_0 ) );
  NAND3_X2 \SB1_2_17/Component_Function_4/N4  ( .A1(\SB1_2_17/i1[9] ), .A2(
        \SB1_2_17/i1_5 ), .A3(\SB1_2_17/i0_4 ), .ZN(
        \SB1_2_17/Component_Function_4/NAND4_in[3] ) );
  BUF_X4 \SB1_3_30/BUF_5  ( .I(\MC_ARK_ARC_1_2/buf_output[11] ), .Z(
        \SB1_3_30/i0_3 ) );
  INV_X2 U651 ( .I(\MC_ARK_ARC_1_3/buf_output[95] ), .ZN(\SB3_16/i1_5 ) );
  NAND3_X2 U3745 ( .A1(\SB3_6/i1_5 ), .A2(\SB3_6/i1[9] ), .A3(\RI1[4][154] ), 
        .ZN(n785) );
  NAND2_X2 U1190 ( .A1(\SB1_2_17/i0_3 ), .A2(\SB1_2_17/i1[9] ), .ZN(
        \SB1_2_17/Component_Function_1/NAND4_in[0] ) );
  INV_X2 U956 ( .I(\MC_ARK_ARC_1_2/buf_output[182] ), .ZN(\SB1_3_1/i1[9] ) );
  NAND3_X2 U2733 ( .A1(\SB1_1_1/i0_0 ), .A2(\SB1_1_1/i0[6] ), .A3(
        \SB1_1_1/i0[10] ), .ZN(\SB1_1_1/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 \SB1_0_4/Component_Function_5/N3  ( .A1(\SB1_0_4/i1[9] ), .A2(
        \SB1_0_4/i0_4 ), .A3(\SB1_0_4/i0_3 ), .ZN(
        \SB1_0_4/Component_Function_5/NAND4_in[2] ) );
  BUF_X4 \MC_ARK_ARC_1_3/BUF_154_1  ( .I(\MC_ARK_ARC_1_3/buf_output[154] ), 
        .Z(\RI1[4][154] ) );
  NAND3_X2 U3019 ( .A1(\SB2_1_29/i1_5 ), .A2(\SB2_1_29/i0[8] ), .A3(
        \SB2_1_29/i3[0] ), .ZN(\SB2_1_29/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 U685 ( .A1(\SB2_3_10/i0[10] ), .A2(\SB2_3_10/i1_5 ), .A3(
        \SB2_3_10/i1[9] ), .ZN(n3565) );
  NAND3_X2 U997 ( .A1(\SB1_1_17/i0_4 ), .A2(\SB1_1_17/i1_5 ), .A3(
        \SB1_1_17/i0_0 ), .ZN(n2013) );
  NAND2_X2 \SB1_0_4/Component_Function_5/N1  ( .A1(\SB1_0_4/i0_0 ), .A2(
        \SB1_0_4/i3[0] ), .ZN(\SB1_0_4/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U2738 ( .A1(\SB1_1_1/i0[10] ), .A2(\SB1_1_1/i0[9] ), .A3(
        \SB1_1_1/i0_3 ), .ZN(\SB1_1_1/Component_Function_4/NAND4_in[2] ) );
  NAND3_X2 \SB2_3_17/Component_Function_2/N4  ( .A1(n4763), .A2(
        \SB2_3_17/i0_0 ), .A3(\SB2_3_17/i0_4 ), .ZN(
        \SB2_3_17/Component_Function_2/NAND4_in[3] ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_49  ( .I(\SB2_2_27/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[49] ) );
  INV_X2 U1566 ( .I(n5504), .ZN(\SB3_17/i0[8] ) );
  BUF_X4 \SB2_0_4/BUF_3_0  ( .I(\SB2_0_4/buf_output[3] ), .Z(\RI5[0][177] ) );
  NAND3_X2 U2884 ( .A1(n3669), .A2(\SB2_3_8/i0_3 ), .A3(\SB2_3_8/i0[6] ), .ZN(
        \SB2_3_8/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 \SB2_2_14/Component_Function_4/N1  ( .A1(\SB2_2_14/i0[9] ), .A2(
        \SB2_2_14/i0_0 ), .A3(\SB2_2_14/i0[8] ), .ZN(
        \SB2_2_14/Component_Function_4/NAND4_in[0] ) );
  NAND3_X2 U2276 ( .A1(\SB2_2_14/i0_3 ), .A2(\SB2_2_14/i0[10] ), .A3(
        \SB2_2_14/i0[9] ), .ZN(n865) );
  NAND3_X2 U5396 ( .A1(\SB2_2_14/i0_3 ), .A2(\SB2_2_14/i0_0 ), .A3(n5932), 
        .ZN(n1597) );
  NAND3_X2 U1495 ( .A1(\SB1_1_16/i0[10] ), .A2(\SB1_1_16/i1[9] ), .A3(
        \SB1_1_16/i1_5 ), .ZN(n2973) );
  INV_X2 \SB1_2_14/INV_2  ( .I(\MC_ARK_ARC_1_1/buf_output[104] ), .ZN(
        \SB1_2_14/i1[9] ) );
  NAND3_X2 U3007 ( .A1(\SB2_1_22/i0_3 ), .A2(\SB2_1_22/i0[8] ), .A3(
        \SB2_1_22/i0[9] ), .ZN(\SB2_1_22/Component_Function_2/NAND4_in[2] ) );
  BUF_X2 U568 ( .I(\SB3_24/buf_output[0] ), .Z(\SB4_19/i0[9] ) );
  NAND3_X2 U7173 ( .A1(\SB2_0_31/i0[9] ), .A2(\SB2_0_31/i0_3 ), .A3(
        \SB2_0_31/i0[8] ), .ZN(\SB2_0_31/Component_Function_2/NAND4_in[2] ) );
  INV_X2 U936 ( .I(\MC_ARK_ARC_1_2/buf_output[161] ), .ZN(\SB1_3_5/i1_5 ) );
  INV_X2 U2548 ( .I(\MC_ARK_ARC_1_0/buf_output[47] ), .ZN(\SB1_1_24/i1_5 ) );
  NAND3_X2 \SB1_1_25/Component_Function_2/N1  ( .A1(\SB1_1_25/i1_5 ), .A2(
        \SB1_1_25/i0[10] ), .A3(\SB1_1_25/i1[9] ), .ZN(
        \SB1_1_25/Component_Function_2/NAND4_in[0] ) );
  NAND2_X2 \SB2_2_17/Component_Function_1/N1  ( .A1(\SB2_2_17/i0_3 ), .A2(
        \SB2_2_17/i1[9] ), .ZN(\SB2_2_17/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 U1274 ( .A1(\SB2_1_13/i0[10] ), .A2(\SB2_1_13/i1[9] ), .A3(
        \SB2_1_13/i1_7 ), .ZN(\SB2_1_13/Component_Function_3/NAND4_in[2] ) );
  INV_X4 U9756 ( .I(n3645), .ZN(n3993) );
  NAND3_X2 \SB1_2_5/Component_Function_2/N4  ( .A1(\SB1_2_5/i1_5 ), .A2(
        \SB1_2_5/i0_0 ), .A3(\SB1_2_5/i0_4 ), .ZN(
        \SB1_2_5/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 \SB2_2_2/Component_Function_3/N1  ( .A1(\SB2_2_2/i1[9] ), .A2(
        \SB2_2_2/i0_3 ), .A3(\SB2_2_2/i0[6] ), .ZN(
        \SB2_2_2/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 U1802 ( .I(\MC_ARK_ARC_1_3/buf_output[62] ), .Z(\SB3_21/i0_0 ) );
  BUF_X4 \SB1_2_24/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[43] ), .Z(
        \SB1_2_24/i0[6] ) );
  NAND3_X2 \SB2_2_7/Component_Function_3/N2  ( .A1(\SB2_2_7/i0_0 ), .A2(
        \SB2_2_7/i0_3 ), .A3(\SB1_2_8/buf_output[4] ), .ZN(
        \SB2_2_7/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U696 ( .A1(\RI3[3][16] ), .A2(\SB2_3_29/i1[9] ), .A3(
        \SB2_3_29/i1_5 ), .ZN(n1986) );
  NAND3_X2 U2342 ( .A1(\SB2_3_16/i0_3 ), .A2(\SB2_3_16/i0_0 ), .A3(
        \SB2_3_16/i0_4 ), .ZN(\SB2_3_16/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U4897 ( .A1(\SB2_2_8/i1_5 ), .A2(\SB2_2_8/i0_0 ), .A3(
        \SB2_2_8/i0_4 ), .ZN(\SB2_2_8/Component_Function_2/NAND4_in[3] ) );
  NAND2_X2 \SB1_2_8/Component_Function_5/N1  ( .A1(\SB1_2_8/i0_0 ), .A2(
        \SB1_2_8/i3[0] ), .ZN(\SB1_2_8/Component_Function_5/NAND4_in[0] ) );
  BUF_X2 \SB2_0_16/BUF_0  ( .I(\SB1_0_21/buf_output[0] ), .Z(\SB2_0_16/i0[9] )
         );
  INV_X2 U2527 ( .I(\SB1_1_10/buf_output[5] ), .ZN(\SB2_1_10/i1_5 ) );
  INV_X2 U4557 ( .I(\RI1[4][5] ), .ZN(\SB3_31/i1_5 ) );
  NAND3_X2 U2882 ( .A1(\SB2_3_8/i0_3 ), .A2(n3669), .A3(
        \SB1_3_9/buf_output[4] ), .ZN(
        \SB2_3_8/Component_Function_5/NAND4_in[2] ) );
  INV_X2 U1508 ( .I(\MC_ARK_ARC_1_2/buf_output[8] ), .ZN(\SB1_3_30/i1[9] ) );
  BUF_X4 \SB1_1_0/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[190] ), .Z(
        \SB1_1_0/i0_4 ) );
  INV_X2 \SB2_0_13/INV_1  ( .I(\SB1_0_17/buf_output[1] ), .ZN(\SB2_0_13/i1_7 )
         );
  NAND2_X2 \SB1_2_28/Component_Function_5/N1  ( .A1(\SB1_2_28/i0_0 ), .A2(
        \SB1_2_28/i3[0] ), .ZN(\SB1_2_28/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U7195 ( .A1(\SB2_0_14/i1[9] ), .A2(\SB2_0_14/i1_5 ), .A3(
        \RI3[0][106] ), .ZN(\SB2_0_14/Component_Function_4/NAND4_in[3] ) );
  NAND3_X2 U4137 ( .A1(\SB2_0_2/i0[6] ), .A2(\SB2_0_2/i0[9] ), .A3(
        \RI3[0][178] ), .ZN(n2964) );
  BUF_X4 U1997 ( .I(\MC_ARK_ARC_1_0/buf_output[41] ), .Z(\SB1_1_25/i0_3 ) );
  NAND3_X2 U660 ( .A1(\SB2_3_7/i0_0 ), .A2(\SB1_3_8/buf_output[4] ), .A3(
        \SB2_3_7/i1_5 ), .ZN(n3765) );
  NAND3_X2 U5744 ( .A1(\SB2_2_21/i0_3 ), .A2(\SB2_2_21/i0[10] ), .A3(
        \SB2_2_21/i0_4 ), .ZN(\SB2_2_21/Component_Function_0/NAND4_in[2] ) );
  INV_X2 \SB2_3_7/INV_0  ( .I(\SB1_3_12/buf_output[0] ), .ZN(\SB2_3_7/i3[0] )
         );
  NAND2_X2 \SB2_1_1/Component_Function_5/N1  ( .A1(\SB2_1_1/i0_0 ), .A2(
        \SB2_1_1/i3[0] ), .ZN(\SB2_1_1/Component_Function_5/NAND4_in[0] ) );
  NAND4_X2 U2429 ( .A1(\SB2_3_2/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_3_2/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_2/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_2/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_3_2/buf_output[1] ) );
  NAND2_X2 \SB1_1_5/Component_Function_5/N1  ( .A1(\SB1_1_5/i0_0 ), .A2(
        \SB1_1_5/i3[0] ), .ZN(\SB1_1_5/Component_Function_5/NAND4_in[0] ) );
  NAND2_X2 U2077 ( .A1(\SB1_2_19/i0_3 ), .A2(\SB1_2_19/i1[9] ), .ZN(
        \SB1_2_19/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 U3719 ( .A1(\SB1_0_28/Component_Function_4/NAND4_in[3] ), .A2(n1784), .ZN(n1783) );
  NAND3_X2 \SB1_0_5/Component_Function_2/N1  ( .A1(\SB1_0_5/i1_5 ), .A2(
        \SB1_0_5/i0[10] ), .A3(\SB1_0_5/i1[9] ), .ZN(
        \SB1_0_5/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 U1467 ( .I(n393), .Z(\SB1_0_5/i0[10] ) );
  NAND3_X2 U4448 ( .A1(\SB3_11/i1_7 ), .A2(\SB3_11/i0[8] ), .A3(\SB3_11/i0_4 ), 
        .ZN(\SB3_11/Component_Function_1/NAND4_in[3] ) );
  BUF_X4 U2869 ( .I(\MC_ARK_ARC_1_2/buf_output[188] ), .Z(\SB1_3_0/i0_0 ) );
  NAND3_X2 U3009 ( .A1(\SB2_1_22/i1[9] ), .A2(\SB2_1_22/i0_3 ), .A3(
        \SB2_1_22/i0[6] ), .ZN(\SB2_1_22/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 \SB2_3_17/Component_Function_4/N4  ( .A1(\SB2_3_17/i1[9] ), .A2(
        n4763), .A3(\SB2_3_17/i0_4 ), .ZN(
        \SB2_3_17/Component_Function_4/NAND4_in[3] ) );
  NAND3_X2 U3597 ( .A1(\SB2_3_8/i0[7] ), .A2(\SB2_3_8/i0[8] ), .A3(
        \SB2_3_8/i0[6] ), .ZN(n1046) );
  NAND2_X2 \SB2_1_0/Component_Function_5/N1  ( .A1(\SB2_1_0/i0_0 ), .A2(
        \SB2_1_0/i3[0] ), .ZN(\SB2_1_0/Component_Function_5/NAND4_in[0] ) );
  INV_X2 U2870 ( .I(\MC_ARK_ARC_1_2/buf_output[188] ), .ZN(\SB1_3_0/i1[9] ) );
  BUF_X4 U667 ( .I(\SB2_3_30/buf_output[1] ), .Z(\RI5[3][31] ) );
  NAND2_X2 \SB2_3_1/Component_Function_5/N1  ( .A1(\SB2_3_1/i0_0 ), .A2(
        \SB2_3_1/i3[0] ), .ZN(\SB2_3_1/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U1358 ( .A1(\SB1_3_15/i0[8] ), .A2(\SB1_3_15/i1_5 ), .A3(
        \SB1_3_15/i3[0] ), .ZN(n1037) );
  BUF_X4 U8923 ( .I(\RI1[4][5] ), .Z(\SB3_31/i0_3 ) );
  INV_X2 \SB1_2_10/INV_1  ( .I(\MC_ARK_ARC_1_1/buf_output[127] ), .ZN(
        \SB1_2_10/i1_7 ) );
  NAND3_X2 U3667 ( .A1(\SB1_3_26/i0_4 ), .A2(\SB1_3_26/i0_0 ), .A3(
        \SB1_3_26/i1_5 ), .ZN(n3165) );
  NAND3_X2 \SB1_2_14/Component_Function_2/N2  ( .A1(\SB1_2_14/i0_3 ), .A2(
        \SB1_2_14/i0[10] ), .A3(\SB1_2_14/i0[6] ), .ZN(
        \SB1_2_14/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 \SB2_0_20/Component_Function_5/N2  ( .A1(\SB2_0_20/i0_0 ), .A2(
        \SB2_0_20/i0[6] ), .A3(\SB2_0_20/i0[10] ), .ZN(
        \SB2_0_20/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U3414 ( .A1(\SB2_0_22/i1[9] ), .A2(\SB2_0_22/i1_5 ), .A3(
        \SB2_0_22/i0_4 ), .ZN(\SB2_0_22/Component_Function_4/NAND4_in[3] ) );
  NAND3_X2 U9656 ( .A1(\SB2_1_10/i0[10] ), .A2(\SB2_1_10/i0_3 ), .A3(
        \SB2_1_10/i0[9] ), .ZN(n3946) );
  NAND3_X2 U9455 ( .A1(\SB1_1_9/i0_0 ), .A2(\SB1_1_9/i1_5 ), .A3(
        \SB1_1_9/i0_4 ), .ZN(n1221) );
  NAND3_X2 U1432 ( .A1(\SB1_1_29/i0[8] ), .A2(\SB1_1_29/i1_5 ), .A3(
        \SB1_1_29/i3[0] ), .ZN(\SB1_1_29/Component_Function_3/NAND4_in[3] ) );
  OAI21_X2 U6466 ( .A1(n4758), .A2(n573), .B(\SB1_1_16/i0_0 ), .ZN(n2256) );
  NAND3_X2 U678 ( .A1(\SB2_3_5/i0_3 ), .A2(\SB2_3_5/i0[9] ), .A3(
        \SB2_3_5/i0[8] ), .ZN(\SB2_3_5/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U807 ( .A1(\SB1_3_23/i0[10] ), .A2(\SB1_3_23/i1[9] ), .A3(
        \SB1_3_23/i1_7 ), .ZN(\SB1_3_23/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U2899 ( .A1(\SB2_3_31/i0_3 ), .A2(\SB2_3_31/i0_0 ), .A3(
        \SB2_3_31/i0[7] ), .ZN(n924) );
  NAND3_X2 U966 ( .A1(\SB2_1_26/i0[10] ), .A2(\SB2_1_26/i1[9] ), .A3(
        \SB2_1_26/i1_7 ), .ZN(\SB2_1_26/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 \SB1_0_31/Component_Function_2/N2  ( .A1(\SB1_0_31/i0_3 ), .A2(
        \SB1_0_31/i0[10] ), .A3(\SB1_0_31/i0[6] ), .ZN(
        \SB1_0_31/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U1382 ( .A1(\SB2_1_25/i0_3 ), .A2(\SB2_1_25/i1[9] ), .A3(n1579), 
        .ZN(n2288) );
  INV_X2 U3100 ( .I(\MC_ARK_ARC_1_1/buf_output[85] ), .ZN(\SB1_2_17/i1_7 ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_22  ( .I(\SB2_0_29/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[22] ) );
  NAND3_X2 \SB1_0_31/Component_Function_5/N2  ( .A1(\SB1_0_31/i0_0 ), .A2(
        \SB1_0_31/i0[6] ), .A3(\SB1_0_31/i0[10] ), .ZN(
        \SB1_0_31/Component_Function_5/NAND4_in[1] ) );
  INV_X2 U2463 ( .I(\MC_ARK_ARC_1_2/buf_output[9] ), .ZN(\SB1_3_30/i0[8] ) );
  NAND3_X2 U1263 ( .A1(\SB2_1_1/i0_3 ), .A2(\SB2_1_1/i0[10] ), .A3(
        \SB2_1_1/i0[9] ), .ZN(n998) );
  BUF_X2 U2999 ( .I(Key[110]), .Z(n205) );
  BUF_X4 U2151 ( .I(\SB3_31/buf_output[5] ), .Z(\SB4_31/i0_3 ) );
  INV_X2 U752 ( .I(\SB1_3_2/buf_output[5] ), .ZN(\SB2_3_2/i1_5 ) );
  NAND3_X2 \SB2_0_19/Component_Function_2/N4  ( .A1(\SB2_0_19/i1_5 ), .A2(
        \SB2_0_19/i0_0 ), .A3(\RI3[0][76] ), .ZN(
        \SB2_0_19/Component_Function_2/NAND4_in[3] ) );
  NAND2_X2 \SB1_3_2/Component_Function_5/N1  ( .A1(\SB1_3_2/i0_0 ), .A2(
        \SB1_3_2/i3[0] ), .ZN(\SB1_3_2/Component_Function_5/NAND4_in[0] ) );
  INV_X2 U2402 ( .I(\SB1_1_20/buf_output[5] ), .ZN(\SB2_1_20/i1_5 ) );
  NAND3_X2 U842 ( .A1(\SB2_2_4/i0[10] ), .A2(\SB2_2_4/i1[9] ), .A3(
        \SB2_2_4/i1_7 ), .ZN(\SB2_2_4/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U1606 ( .A1(\SB2_0_14/i0[6] ), .A2(\RI3[0][105] ), .A3(
        \RI3[0][104] ), .ZN(\SB2_0_14/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U1456 ( .A1(\SB2_0_21/i0_3 ), .A2(\SB2_0_21/i0_4 ), .A3(
        \SB2_0_21/i1[9] ), .ZN(n2353) );
  INV_X2 \SB1_0_3/INV_3  ( .I(n397), .ZN(\SB1_0_3/i0[8] ) );
  NAND3_X2 U990 ( .A1(\SB2_2_24/i0[10] ), .A2(\SB2_2_24/i1_7 ), .A3(
        \SB2_2_24/i1[9] ), .ZN(n4408) );
  NAND2_X2 U5445 ( .A1(\SB1_1_31/Component_Function_4/NAND4_in[1] ), .A2(n2557), .ZN(n2556) );
  NAND3_X2 U2433 ( .A1(\SB3_17/i0_3 ), .A2(\SB3_17/i0[8] ), .A3(\SB3_17/i0[9] ), .ZN(\SB3_17/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 \SB2_1_27/Component_Function_3/N1  ( .A1(\SB2_1_27/i1[9] ), .A2(
        \SB2_1_27/i0_3 ), .A3(\SB2_1_27/i0[6] ), .ZN(
        \SB2_1_27/Component_Function_3/NAND4_in[0] ) );
  INV_X2 \SB2_0_26/INV_5  ( .I(\SB1_0_26/buf_output[5] ), .ZN(\SB2_0_26/i1_5 )
         );
  BUF_X2 \SB2_0_3/BUF_1  ( .I(\SB1_0_7/buf_output[1] ), .Z(\SB2_0_3/i0[6] ) );
  NAND2_X2 \SB1_1_23/Component_Function_1/N1  ( .A1(\SB1_1_23/i0_3 ), .A2(
        \SB1_1_23/i1[9] ), .ZN(\SB1_1_23/Component_Function_1/NAND4_in[0] ) );
  NAND2_X2 U3508 ( .A1(\SB2_1_31/i0_0 ), .A2(\SB2_1_31/i3[0] ), .ZN(
        \SB2_1_31/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U3098 ( .A1(\SB1_2_20/i1[9] ), .A2(\SB1_2_20/i0_4 ), .A3(
        \SB1_2_20/i0_3 ), .ZN(\SB1_2_20/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 \SB1_3_22/Component_Function_1/N4  ( .A1(\SB1_3_22/i1_7 ), .A2(
        \SB1_3_22/i0[8] ), .A3(\SB1_3_22/i0_4 ), .ZN(
        \SB1_3_22/Component_Function_1/NAND4_in[3] ) );
  NAND4_X1 \SB2_3_11/Component_Function_1/N5  ( .A1(
        \SB2_3_11/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_11/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_11/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_3_11/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_3_11/buf_output[1] ) );
  NAND3_X2 \SB2_1_28/Component_Function_2/N1  ( .A1(\SB2_1_28/i1_5 ), .A2(
        \SB2_1_28/i0[10] ), .A3(\SB2_1_28/i1[9] ), .ZN(
        \SB2_1_28/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB1_2_21/Component_Function_5/N2  ( .A1(\SB1_2_21/i0_0 ), .A2(
        \SB1_2_21/i0[6] ), .A3(\SB1_2_21/i0[10] ), .ZN(
        \SB1_2_21/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 U4804 ( .I(\SB2_1_28/buf_output[3] ), .Z(n1383) );
  INV_X2 \SB2_1_28/INV_5  ( .I(\SB1_1_28/buf_output[5] ), .ZN(\SB2_1_28/i1_5 )
         );
  NAND2_X2 U3348 ( .A1(\SB1_0_31/i0_0 ), .A2(\SB1_0_31/i3[0] ), .ZN(n2180) );
  INV_X2 U8861 ( .I(\MC_ARK_ARC_1_2/buf_output[119] ), .ZN(\SB1_3_12/i1_5 ) );
  NAND3_X2 U1969 ( .A1(\SB2_0_4/i1[9] ), .A2(\RI3[0][166] ), .A3(
        \SB2_0_4/i0_3 ), .ZN(\SB2_0_4/Component_Function_5/NAND4_in[2] ) );
  INV_X2 U2627 ( .I(\MC_ARK_ARC_1_3/buf_output[2] ), .ZN(\SB3_31/i1[9] ) );
  BUF_X4 U2628 ( .I(\MC_ARK_ARC_1_3/buf_output[2] ), .Z(\SB3_31/i0_0 ) );
  NAND3_X2 U3006 ( .A1(\SB2_1_22/i0_3 ), .A2(\SB2_1_22/i0[10] ), .A3(
        \SB2_1_22/i0_4 ), .ZN(n2997) );
  NAND3_X2 \SB2_2_8/Component_Function_3/N1  ( .A1(\SB2_2_8/i1[9] ), .A2(
        \SB2_2_8/i0_3 ), .A3(\SB2_2_8/i0[6] ), .ZN(
        \SB2_2_8/Component_Function_3/NAND4_in[0] ) );
  INV_X2 \SB1_1_20/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[67] ), .ZN(
        \SB1_1_20/i1_7 ) );
  NAND3_X2 U1307 ( .A1(\SB2_1_17/i3[0] ), .A2(\SB2_1_17/i1_5 ), .A3(
        \SB2_1_17/i0[8] ), .ZN(\SB2_1_17/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 U3764 ( .A1(\SB3_31/i0[10] ), .A2(\SB3_31/i1[9] ), .A3(
        \SB3_31/i1_7 ), .ZN(n2072) );
  BUF_X4 \SB2_0_28/BUF_3  ( .I(\SB1_0_30/buf_output[3] ), .Z(\SB2_0_28/i0[10] ) );
  NAND3_X2 U7809 ( .A1(\SB2_0_13/i0_0 ), .A2(\SB2_0_13/i0_4 ), .A3(
        \SB2_0_13/i0_3 ), .ZN(\SB2_0_13/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U1148 ( .A1(\SB1_2_26/i0[9] ), .A2(\SB1_2_26/i0[6] ), .A3(
        \SB1_2_26/i0_4 ), .ZN(n2575) );
  NAND3_X2 \SB2_1_26/Component_Function_3/N1  ( .A1(\SB2_1_26/i1[9] ), .A2(
        \SB2_1_26/i0_3 ), .A3(\SB2_1_26/i0[6] ), .ZN(
        \SB2_1_26/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U3963 ( .A1(\SB2_2_17/i0_3 ), .A2(\SB2_2_17/i1[9] ), .A3(
        \SB2_2_17/i0[6] ), .ZN(\SB2_2_17/Component_Function_3/NAND4_in[0] ) );
  CLKBUF_X4 U3360 ( .I(n321), .Z(\SB1_0_6/i0[6] ) );
  BUF_X4 \SB1_1_9/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[133] ), .Z(
        \SB1_1_9/i0[6] ) );
  INV_X2 U2826 ( .I(\MC_ARK_ARC_1_1/buf_output[109] ), .ZN(\SB1_2_13/i1_7 ) );
  NAND3_X2 U6327 ( .A1(\SB1_3_2/i0[10] ), .A2(\SB1_3_2/i1[9] ), .A3(
        \SB1_3_2/i1_5 ), .ZN(\SB1_3_2/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 \SB2_3_16/BUF_5  ( .I(\SB1_3_16/buf_output[5] ), .Z(\SB2_3_16/i0_3 )
         );
  INV_X2 \SB2_2_13/INV_1  ( .I(\SB1_2_17/buf_output[1] ), .ZN(\SB2_2_13/i1_7 )
         );
  BUF_X4 U8998 ( .I(\RI3[0][183] ), .Z(\SB2_0_1/i0[10] ) );
  INV_X2 U1400 ( .I(\SB1_3_28/buf_output[5] ), .ZN(\SB2_3_28/i1_5 ) );
  NAND2_X2 \SB1_3_28/Component_Function_5/N1  ( .A1(\SB1_3_28/i0_0 ), .A2(
        \SB1_3_28/i3[0] ), .ZN(\SB1_3_28/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U1245 ( .A1(\SB1_3_22/i0[9] ), .A2(\SB1_3_22/i0[6] ), .A3(
        \SB1_3_22/i0_4 ), .ZN(\SB1_3_22/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 \SB2_2_21/Component_Function_0/N2  ( .A1(\SB2_2_21/i0[8] ), .A2(
        \SB2_2_21/i0[7] ), .A3(\SB2_2_21/i0[6] ), .ZN(
        \SB2_2_21/Component_Function_0/NAND4_in[1] ) );
  NAND3_X2 \SB2_0_3/Component_Function_3/N2  ( .A1(\SB2_0_3/i0_0 ), .A2(
        \SB2_0_3/i0_3 ), .A3(\RI3[0][172] ), .ZN(
        \SB2_0_3/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U3622 ( .A1(\SB2_2_30/i0[10] ), .A2(\SB2_2_30/i1_7 ), .A3(
        \SB2_2_30/i1[9] ), .ZN(n1647) );
  NAND3_X2 U2890 ( .A1(\SB2_3_8/i0_3 ), .A2(\SB2_3_8/i0[6] ), .A3(
        \SB2_3_8/i0[10] ), .ZN(\SB2_3_8/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U590 ( .A1(\SB3_7/i0_3 ), .A2(\SB3_7/i0[8] ), .A3(\SB3_7/i0[9] ), 
        .ZN(n4727) );
  NAND3_X2 \SB1_2_16/Component_Function_1/N3  ( .A1(\SB1_2_16/i1_5 ), .A2(
        \SB1_2_16/i0[6] ), .A3(\SB1_2_16/i0[9] ), .ZN(
        \SB1_2_16/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 \SB2_3_10/Component_Function_5/N2  ( .A1(\SB2_3_10/i0_0 ), .A2(
        \SB2_3_10/i0[6] ), .A3(\SB2_3_10/i0[10] ), .ZN(
        \SB2_3_10/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 U3147 ( .I(\MC_ARK_ARC_1_1/buf_output[95] ), .Z(\RI1[2][95] ) );
  NAND3_X2 U1472 ( .A1(\SB1_3_4/i0_0 ), .A2(\SB1_3_4/i0_4 ), .A3(
        \SB1_3_4/i1_5 ), .ZN(n2670) );
  NAND3_X2 U2885 ( .A1(\SB2_3_8/i0_3 ), .A2(\SB2_3_8/i0[10] ), .A3(
        \SB2_3_8/i0[9] ), .ZN(n4282) );
  NAND2_X2 U1281 ( .A1(n1752), .A2(n4182), .ZN(n3396) );
  NAND3_X2 \SB2_2_27/Component_Function_0/N3  ( .A1(\SB2_2_27/i0[10] ), .A2(
        \SB1_2_28/buf_output[4] ), .A3(\SB2_2_27/i0_3 ), .ZN(
        \SB2_2_27/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 U2655 ( .A1(\SB2_1_23/i0_3 ), .A2(\SB2_1_23/i0_4 ), .A3(
        \SB2_1_23/i1[9] ), .ZN(n1992) );
  INV_X8 \SB2_0_14/INV_2  ( .I(\RI3[0][104] ), .ZN(\SB2_0_14/i1[9] ) );
  BUF_X4 U8191 ( .I(\SB2_2_17/buf_output[1] ), .Z(\RI5[2][109] ) );
  NAND4_X2 \SB2_2_17/Component_Function_1/N5  ( .A1(
        \SB2_2_17/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_17/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_17/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_2_17/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_2_17/buf_output[1] ) );
  INV_X2 \SB2_3_15/INV_1  ( .I(\SB1_3_19/buf_output[1] ), .ZN(\SB2_3_15/i1_7 )
         );
  NAND3_X2 \SB1_2_10/Component_Function_2/N2  ( .A1(\SB1_2_10/i0_3 ), .A2(
        \SB1_2_10/i0[10] ), .A3(\SB1_2_10/i0[6] ), .ZN(
        \SB1_2_10/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U873 ( .A1(\SB1_3_26/i0[10] ), .A2(\SB1_3_26/i1[9] ), .A3(
        \SB1_3_26/i1_5 ), .ZN(n4467) );
  NAND3_X2 U3440 ( .A1(\SB1_3_24/i0[10] ), .A2(\SB1_3_24/i1[9] ), .A3(
        \SB1_3_24/i1_7 ), .ZN(\SB1_3_24/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U2128 ( .A1(\SB2_2_23/i1[9] ), .A2(\SB2_2_23/i1_7 ), .A3(
        \SB2_2_23/i0[10] ), .ZN(\SB2_2_23/Component_Function_3/NAND4_in[2] )
         );
  NAND3_X2 \SB1_2_25/Component_Function_3/N2  ( .A1(\SB1_2_25/i0_0 ), .A2(
        \SB1_2_25/i0_3 ), .A3(\SB1_2_25/i0_4 ), .ZN(
        \SB1_2_25/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 \SB1_0_4/Component_Function_5/N2  ( .A1(\SB1_0_4/i0_0 ), .A2(
        \SB1_0_4/i0[6] ), .A3(\SB1_0_4/i0[10] ), .ZN(
        \SB1_0_4/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 \SB1_2_25/BUF_3  ( .I(\MC_ARK_ARC_1_1/buf_output[39] ), .Z(
        \SB1_2_25/i0[10] ) );
  INV_X2 U1067 ( .I(\SB1_2_26/buf_output[2] ), .ZN(\SB2_2_23/i1[9] ) );
  NAND3_X2 U4595 ( .A1(\SB1_3_23/i0_0 ), .A2(\SB1_3_23/i1_5 ), .A3(
        \SB1_3_23/i0_4 ), .ZN(n2778) );
  INV_X2 U3845 ( .I(\MC_ARK_ARC_1_1/buf_output[33] ), .ZN(\SB1_2_26/i0[8] ) );
  BUF_X4 \SB2_3_13/BUF_5  ( .I(\SB1_3_13/buf_output[5] ), .Z(\SB2_3_13/i0_3 )
         );
  NAND3_X2 U2272 ( .A1(\SB1_2_9/i0[10] ), .A2(\SB1_2_9/i1_5 ), .A3(
        \SB1_2_9/i1[9] ), .ZN(n3317) );
  NAND3_X2 U3671 ( .A1(\SB1_3_16/i0_3 ), .A2(\SB1_3_16/i0_4 ), .A3(
        \SB1_3_16/i1[9] ), .ZN(n1333) );
  INV_X2 U1244 ( .I(\MC_ARK_ARC_1_1/buf_output[134] ), .ZN(\SB1_2_9/i1[9] ) );
  INV_X2 U4495 ( .I(\MC_ARK_ARC_1_2/buf_output[103] ), .ZN(\SB1_3_14/i1_7 ) );
  NAND3_X2 U2589 ( .A1(\RI3[0][155] ), .A2(\SB2_0_6/i1[9] ), .A3(\RI3[0][154] ), .ZN(n3883) );
  NAND3_X2 U2756 ( .A1(\SB2_2_19/i0[10] ), .A2(\SB2_2_19/i1_5 ), .A3(
        \SB2_2_19/i1[9] ), .ZN(\SB2_2_19/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U8726 ( .A1(n3647), .A2(\SB1_1_8/i1[9] ), .A3(\SB1_1_8/i0[10] ), 
        .ZN(n911) );
  NAND3_X2 U765 ( .A1(\SB1_3_26/i0[6] ), .A2(\SB1_3_26/i0[9] ), .A3(
        \SB1_3_26/i0_4 ), .ZN(n1871) );
  NAND3_X2 \SB1_3_27/Component_Function_4/N4  ( .A1(\SB1_3_27/i1[9] ), .A2(
        \SB1_3_27/i1_5 ), .A3(\SB1_3_27/i0_4 ), .ZN(
        \SB1_3_27/Component_Function_4/NAND4_in[3] ) );
  INV_X2 U3690 ( .I(\SB1_3_23/buf_output[5] ), .ZN(\SB2_3_23/i1_5 ) );
  INV_X2 U1379 ( .I(\MC_ARK_ARC_1_3/buf_output[191] ), .ZN(\SB3_0/i1_5 ) );
  INV_X2 U2275 ( .I(\MC_ARK_ARC_1_2/buf_output[101] ), .ZN(\SB1_3_15/i1_5 ) );
  BUF_X4 \SB1_0_20/BUF_4  ( .I(n364), .Z(\SB1_0_20/i0_4 ) );
  BUF_X4 \SB2_1_27/BUF_1  ( .I(\SB1_1_31/buf_output[1] ), .Z(\SB2_1_27/i0[6] )
         );
  BUF_X4 U1921 ( .I(\SB1_0_12/buf_output[0] ), .Z(\SB2_0_7/i0[9] ) );
  NAND3_X2 U8666 ( .A1(\SB1_1_14/i0[8] ), .A2(\SB1_1_14/i0_4 ), .A3(
        \SB1_1_14/i1_7 ), .ZN(n2192) );
  NAND3_X2 U3020 ( .A1(\SB2_1_29/i1_5 ), .A2(\SB2_1_29/i0[10] ), .A3(
        \SB2_1_29/i1[9] ), .ZN(\SB2_1_29/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U3917 ( .A1(\SB1_0_12/i0[10] ), .A2(\SB1_0_12/i1[9] ), .A3(
        \SB1_0_12/i1_7 ), .ZN(n2655) );
  NAND3_X2 U1368 ( .A1(\SB2_1_4/i0_3 ), .A2(\SB1_1_5/buf_output[4] ), .A3(
        \SB1_1_7/buf_output[2] ), .ZN(n790) );
  INV_X2 \SB1_3_9/INV_1  ( .I(\MC_ARK_ARC_1_2/buf_output[133] ), .ZN(
        \SB1_3_9/i1_7 ) );
  BUF_X2 U1658 ( .I(Key[170]), .Z(n129) );
  NAND3_X2 \SB2_2_2/Component_Function_3/N4  ( .A1(\SB2_2_2/i1_5 ), .A2(
        \SB2_2_2/i0[8] ), .A3(\SB2_2_2/i3[0] ), .ZN(
        \SB2_2_2/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 \SB1_0_20/Component_Function_2/N1  ( .A1(\SB1_0_20/i1_5 ), .A2(
        \SB1_0_20/i0[10] ), .A3(\SB1_0_20/i1[9] ), .ZN(
        \SB1_0_20/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U2165 ( .A1(\SB3_22/i0_0 ), .A2(\SB3_22/i1_5 ), .A3(\SB3_22/i0_4 ), 
        .ZN(n3494) );
  NAND3_X2 U3530 ( .A1(\SB2_1_20/i0[10] ), .A2(\SB2_1_20/i0_3 ), .A3(
        \SB2_1_20/i0[9] ), .ZN(n1275) );
  NAND3_X2 U9224 ( .A1(\SB2_1_26/i0_3 ), .A2(\SB2_1_26/i0[10] ), .A3(
        \SB2_1_26/i0[9] ), .ZN(n3757) );
  NAND2_X2 \SB2_1_15/Component_Function_1/N1  ( .A1(\SB2_1_15/i0_3 ), .A2(
        \SB2_1_15/i1[9] ), .ZN(\SB2_1_15/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 U1387 ( .A1(\SB1_1_27/i0_4 ), .A2(\SB1_1_27/i1[9] ), .A3(
        \SB1_1_27/i0_3 ), .ZN(n4087) );
  NAND3_X2 U947 ( .A1(\SB2_1_8/i0_3 ), .A2(n2745), .A3(\SB2_1_8/i0[8] ), .ZN(
        \SB2_1_8/Component_Function_2/NAND4_in[2] ) );
  NAND2_X2 U2162 ( .A1(\SB3_22/i0_0 ), .A2(\SB3_22/i3[0] ), .ZN(
        \SB3_22/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB1_2_6/Component_Function_4/N3  ( .A1(\SB1_2_6/i0[9] ), .A2(
        \SB1_2_6/i0[10] ), .A3(\SB1_2_6/i0_3 ), .ZN(
        \SB1_2_6/Component_Function_4/NAND4_in[2] ) );
  NAND3_X2 U1558 ( .A1(\RI3[0][88] ), .A2(\SB2_0_17/i1_7 ), .A3(
        \SB2_0_17/i0[8] ), .ZN(n3507) );
  NAND4_X2 U4954 ( .A1(\SB2_2_7/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_2_7/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_2_7/Component_Function_1/NAND4_in[0] ), .A4(
        \SB2_2_7/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_2_7/buf_output[1] ) );
  NAND3_X2 \SB2_1_14/Component_Function_3/N2  ( .A1(\SB2_1_14/i0_0 ), .A2(
        \SB2_1_14/i0_3 ), .A3(\SB2_1_14/i0_4 ), .ZN(
        \SB2_1_14/Component_Function_3/NAND4_in[1] ) );
  INV_X2 U2249 ( .I(\MC_ARK_ARC_1_1/buf_output[123] ), .ZN(\SB1_2_11/i0[8] )
         );
  NAND3_X2 \SB2_3_7/Component_Function_3/N4  ( .A1(\SB2_3_7/i1_5 ), .A2(
        \SB2_3_7/i0[8] ), .A3(\SB2_3_7/i3[0] ), .ZN(
        \SB2_3_7/Component_Function_3/NAND4_in[3] ) );
  INV_X2 U3087 ( .I(\MC_ARK_ARC_1_1/buf_output[119] ), .ZN(\SB1_2_12/i1_5 ) );
  BUF_X4 \SB1_0_18/BUF_1  ( .I(n285), .Z(\SB1_0_18/i0[6] ) );
  CLKBUF_X8 U1805 ( .I(\RI1[1][71] ), .Z(\SB1_1_20/i0_3 ) );
  NAND3_X2 \SB1_1_6/Component_Function_1/N4  ( .A1(\SB1_1_6/i1_7 ), .A2(
        \SB1_1_6/i0[8] ), .A3(\SB1_1_6/i0_4 ), .ZN(
        \SB1_1_6/Component_Function_1/NAND4_in[3] ) );
  INV_X2 \SB2_0_1/INV_1  ( .I(\SB1_0_5/buf_output[1] ), .ZN(\SB2_0_1/i1_7 ) );
  NAND3_X2 U913 ( .A1(\SB1_3_19/i0_3 ), .A2(\SB1_3_19/i1[9] ), .A3(
        \SB1_3_19/i0_4 ), .ZN(\SB1_3_19/Component_Function_5/NAND4_in[2] ) );
  BUF_X4 U2407 ( .I(\SB1_1_20/buf_output[5] ), .Z(\SB2_1_20/i0_3 ) );
  NAND3_X2 U2761 ( .A1(\SB2_2_19/i0_3 ), .A2(\SB2_2_19/i0_4 ), .A3(
        \SB2_2_19/i1[9] ), .ZN(n4561) );
  NAND3_X2 \SB2_0_4/Component_Function_0/N3  ( .A1(\SB2_0_4/i0[10] ), .A2(
        \RI3[0][166] ), .A3(\SB2_0_4/i0_3 ), .ZN(
        \SB2_0_4/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 \SB1_2_22/Component_Function_2/N1  ( .A1(\SB1_2_22/i1_5 ), .A2(
        \SB1_2_22/i0[10] ), .A3(\SB1_2_22/i1[9] ), .ZN(
        \SB1_2_22/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U8921 ( .A1(\SB4_14/i0_0 ), .A2(\SB4_14/i0[6] ), .A3(
        \SB4_14/i0[10] ), .ZN(\SB4_14/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 U3577 ( .I(\MC_ARK_ARC_1_3/buf_output[185] ), .Z(\SB3_1/i0_3 ) );
  BUF_X4 U4566 ( .I(\SB1_0_4/buf_output[5] ), .Z(\SB2_0_4/i0_3 ) );
  NAND3_X2 \SB2_2_4/Component_Function_2/N4  ( .A1(\SB2_2_4/i1_5 ), .A2(
        \SB2_2_4/i0_0 ), .A3(\SB2_2_4/i0_4 ), .ZN(
        \SB2_2_4/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 \SB2_3_5/Component_Function_5/N2  ( .A1(\SB2_3_5/i0_0 ), .A2(
        \SB2_3_5/i0[6] ), .A3(\SB2_3_5/i0[10] ), .ZN(
        \SB2_3_5/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 \SB2_1_10/Component_Function_3/N4  ( .A1(\SB2_1_10/i1_5 ), .A2(
        \SB2_1_10/i0[8] ), .A3(\SB2_1_10/i3[0] ), .ZN(
        \SB2_1_10/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 \SB2_2_4/Component_Function_3/N4  ( .A1(\SB2_2_4/i1_5 ), .A2(
        \SB2_2_4/i0[8] ), .A3(\SB2_2_4/i3[0] ), .ZN(
        \SB2_2_4/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 \SB2_0_28/Component_Function_5/N2  ( .A1(\SB2_0_28/i0_0 ), .A2(
        \SB2_0_28/i0[6] ), .A3(\SB2_0_28/i0[10] ), .ZN(
        \SB2_0_28/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 \SB1_0_25/Component_Function_3/N1  ( .A1(\SB1_0_25/i1[9] ), .A2(
        \SB1_0_25/i0_3 ), .A3(\SB1_0_25/i0[6] ), .ZN(
        \SB1_0_25/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 \SB1_2_3/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[172] ), .Z(
        \SB1_2_3/i0_4 ) );
  NAND3_X2 U10564 ( .A1(\SB2_2_14/i1[9] ), .A2(n5932), .A3(\SB2_2_14/i1_5 ), 
        .ZN(\SB2_2_14/Component_Function_4/NAND4_in[3] ) );
  AND4_X2 U2196 ( .A1(\SB3_8/Component_Function_3/NAND4_in[1] ), .A2(
        \SB3_8/Component_Function_3/NAND4_in[0] ), .A3(
        \SB3_8/Component_Function_3/NAND4_in[2] ), .A4(n2113), .Z(n579) );
  NAND3_X2 \SB2_0_12/Component_Function_5/N2  ( .A1(\SB2_0_12/i0_0 ), .A2(
        \SB2_0_12/i0[6] ), .A3(\SB2_0_12/i0[10] ), .ZN(
        \SB2_0_12/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 \SB1_3_19/BUF_5  ( .I(\MC_ARK_ARC_1_2/buf_output[77] ), .Z(
        \SB1_3_19/i0_3 ) );
  NAND2_X2 \SB2_1_24/Component_Function_5/N1  ( .A1(\SB2_1_24/i0_0 ), .A2(
        \SB2_1_24/i3[0] ), .ZN(\SB2_1_24/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U4627 ( .A1(\SB3_9/i1_5 ), .A2(\SB3_9/i0[10] ), .A3(\SB3_9/i1[9] ), 
        .ZN(\SB3_9/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 U2837 ( .I(\SB1_1_12/buf_output[1] ), .Z(\SB2_1_8/i0[6] ) );
  NAND2_X2 \SB1_1_23/Component_Function_5/N1  ( .A1(\SB1_1_23/i0_0 ), .A2(
        \SB1_1_23/i3[0] ), .ZN(\SB1_1_23/Component_Function_5/NAND4_in[0] ) );
  INV_X2 U1759 ( .I(\MC_ARK_ARC_1_2/buf_output[29] ), .ZN(\SB1_3_27/i1_5 ) );
  NAND2_X2 \SB2_2_12/Component_Function_1/N1  ( .A1(\SB2_2_12/i0_3 ), .A2(
        \SB2_2_12/i1[9] ), .ZN(\SB2_2_12/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 \SB2_0_18/Component_Function_5/N2  ( .A1(\SB2_0_18/i0_0 ), .A2(
        \SB2_0_18/i0[6] ), .A3(\SB2_0_18/i0[10] ), .ZN(
        \SB2_0_18/Component_Function_5/NAND4_in[1] ) );
  INV_X2 U8973 ( .I(\SB1_3_24/buf_output[2] ), .ZN(\SB2_3_21/i1[9] ) );
  INV_X2 U3186 ( .I(\SB1_2_0/buf_output[5] ), .ZN(\SB2_2_0/i1_5 ) );
  NAND2_X2 \SB2_3_10/Component_Function_5/N1  ( .A1(\SB2_3_10/i0_0 ), .A2(
        \SB2_3_10/i3[0] ), .ZN(\SB2_3_10/Component_Function_5/NAND4_in[0] ) );
  NAND2_X2 \SB1_2_24/Component_Function_5/N1  ( .A1(\SB1_2_24/i0_0 ), .A2(
        \SB1_2_24/i3[0] ), .ZN(\SB1_2_24/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U2682 ( .A1(\SB1_3_4/i0[6] ), .A2(\SB1_3_4/i0[10] ), .A3(
        \SB1_3_4/i0_0 ), .ZN(n2284) );
  NAND3_X2 U687 ( .A1(\SB2_3_12/i0[10] ), .A2(\SB2_3_12/i0_3 ), .A3(
        \SB2_3_12/i0[6] ), .ZN(n4113) );
  INV_X2 \SB4_2/INV_1  ( .I(\SB3_6/buf_output[1] ), .ZN(\SB4_2/i1_7 ) );
  NAND3_X2 U1189 ( .A1(\SB4_31/i0_0 ), .A2(\SB4_31/i0_3 ), .A3(\SB4_31/i0_4 ), 
        .ZN(\SB4_31/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U2125 ( .A1(\SB4_2/i0_4 ), .A2(\SB4_2/i1_5 ), .A3(\SB4_2/i1[9] ), 
        .ZN(n4592) );
  NAND3_X2 U1374 ( .A1(\SB2_1_4/i0_3 ), .A2(\SB1_1_5/buf_output[4] ), .A3(
        n3660), .ZN(\SB2_1_4/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U854 ( .A1(\SB2_2_0/i0[10] ), .A2(\SB2_2_0/i1[9] ), .A3(
        \SB2_2_0/i1_7 ), .ZN(n2553) );
  NAND3_X2 U2581 ( .A1(\SB1_0_19/i0[10] ), .A2(\SB1_0_19/i1[9] ), .A3(
        \SB1_0_19/i1_7 ), .ZN(\SB1_0_19/Component_Function_3/NAND4_in[2] ) );
  BUF_X4 U3142 ( .I(\SB2_1_3/buf_output[2] ), .Z(\RI5[1][188] ) );
  NAND2_X2 \SB1_3_31/Component_Function_1/N1  ( .A1(\SB1_3_31/i0_3 ), .A2(
        \SB1_3_31/i1[9] ), .ZN(\SB1_3_31/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 \SB1_1_23/Component_Function_5/N4  ( .A1(\SB1_1_23/i0[9] ), .A2(
        \SB1_1_23/i0[6] ), .A3(\SB1_1_23/i0_4 ), .ZN(
        \SB1_1_23/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 U1390 ( .A1(\SB1_1_18/i0[10] ), .A2(\SB1_1_18/i0_3 ), .A3(
        \SB1_1_18/i0[6] ), .ZN(\SB1_1_18/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 U2568 ( .I(\SB1_3_12/buf_output[5] ), .Z(\SB2_3_12/i0_3 ) );
  NAND3_X2 U7905 ( .A1(\SB2_2_6/i0_0 ), .A2(\SB2_2_6/i1_5 ), .A3(n2074), .ZN(
        n2858) );
  BUF_X4 \SB1_0_5/BUF_4_0  ( .I(\SB1_0_5/buf_output[4] ), .Z(\RI3[0][166] ) );
  INV_X2 \SB2_2_6/INV_5  ( .I(\SB1_2_6/buf_output[5] ), .ZN(\SB2_2_6/i1_5 ) );
  NAND3_X2 \SB1_3_31/Component_Function_1/N4  ( .A1(\SB1_3_31/i1_7 ), .A2(
        \SB1_3_31/i0[8] ), .A3(\SB1_3_31/i0_4 ), .ZN(
        \SB1_3_31/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 \SB1_2_19/Component_Function_2/N2  ( .A1(\SB1_2_19/i0_3 ), .A2(
        \SB1_2_19/i0[10] ), .A3(\SB1_2_19/i0[6] ), .ZN(
        \SB1_2_19/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U4660 ( .A1(\SB1_0_6/i0_3 ), .A2(\SB1_0_6/i0_4 ), .A3(
        \SB1_0_6/i1[9] ), .ZN(n1969) );
  NAND3_X2 U1152 ( .A1(\SB1_2_9/i0_0 ), .A2(\SB1_2_9/i0_4 ), .A3(
        \SB1_2_9/i1_5 ), .ZN(n4108) );
  NAND3_X2 U7627 ( .A1(\SB1_1_19/i0_4 ), .A2(\SB1_1_19/i0[6] ), .A3(
        \SB1_1_19/i0[9] ), .ZN(n2706) );
  INV_X2 U3174 ( .I(\MC_ARK_ARC_1_2/buf_output[155] ), .ZN(\SB1_3_6/i1_5 ) );
  BUF_X4 U2558 ( .I(\SB1_0_6/buf_output[5] ), .Z(\RI3[0][155] ) );
  NAND2_X2 \SB2_0_3/Component_Function_5/N1  ( .A1(\SB2_0_3/i0_0 ), .A2(
        \SB2_0_3/i3[0] ), .ZN(\SB2_0_3/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U9665 ( .A1(\SB2_3_17/i0_3 ), .A2(\SB2_3_17/i0[10] ), .A3(
        \SB2_3_17/i0_4 ), .ZN(n793) );
  NAND3_X2 U2681 ( .A1(\SB2_2_15/i0[6] ), .A2(\SB2_2_15/i0_3 ), .A3(
        \SB2_2_15/i0[10] ), .ZN(n3152) );
  NAND3_X2 \SB2_2_16/Component_Function_2/N2  ( .A1(\SB2_2_16/i0_3 ), .A2(
        \SB2_2_16/i0[10] ), .A3(\SB2_2_16/i0[6] ), .ZN(
        \SB2_2_16/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 \SB2_1_9/Component_Function_4/N3  ( .A1(\SB2_1_9/i0[9] ), .A2(
        \SB2_1_9/i0[10] ), .A3(\SB2_1_9/i0_3 ), .ZN(
        \SB2_1_9/Component_Function_4/NAND4_in[2] ) );
  INV_X2 U3516 ( .I(\SB1_2_13/buf_output[3] ), .ZN(\SB2_2_11/i0[8] ) );
  NAND3_X2 \SB1_1_31/Component_Function_0/N3  ( .A1(\SB1_1_31/i0[10] ), .A2(
        \SB1_1_31/i0_4 ), .A3(\SB1_1_31/i0_3 ), .ZN(
        \SB1_1_31/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 \SB2_0_3/Component_Function_0/N4  ( .A1(\SB2_0_3/i0[7] ), .A2(
        \SB2_0_3/i0_3 ), .A3(\SB2_0_3/i0_0 ), .ZN(
        \SB2_0_3/Component_Function_0/NAND4_in[3] ) );
  NAND3_X2 U2390 ( .A1(\SB2_0_17/i1[9] ), .A2(\SB2_0_17/i1_7 ), .A3(
        \SB2_0_17/i0[10] ), .ZN(\SB2_0_17/Component_Function_3/NAND4_in[2] )
         );
  NAND3_X2 U961 ( .A1(\SB2_1_8/i0_0 ), .A2(\SB2_1_8/i1_5 ), .A3(\SB2_1_8/i0_4 ), .ZN(n2379) );
  BUF_X4 U1385 ( .I(\SB1_1_15/buf_output[0] ), .Z(\SB2_1_10/i0[9] ) );
  BUF_X4 U1899 ( .I(\SB1_1_13/buf_output[4] ), .Z(\SB2_1_12/i0_4 ) );
  NAND3_X2 \SB1_3_6/Component_Function_3/N2  ( .A1(\SB1_3_6/i0_0 ), .A2(
        \SB1_3_6/i0_3 ), .A3(\SB1_3_6/i0_4 ), .ZN(
        \SB1_3_6/Component_Function_3/NAND4_in[1] ) );
  INV_X2 U2791 ( .I(\MC_ARK_ARC_1_3/buf_output[188] ), .ZN(\SB3_0/i1[9] ) );
  NAND3_X2 U5688 ( .A1(\SB2_2_3/i0_3 ), .A2(\SB2_2_3/i0_0 ), .A3(
        \SB1_2_4/buf_output[4] ), .ZN(
        \SB2_2_3/Component_Function_3/NAND4_in[1] ) );
  BUF_X4 U2325 ( .I(\MC_ARK_ARC_1_2/buf_output[155] ), .Z(\SB1_3_6/i0_3 ) );
  BUF_X4 U2872 ( .I(\SB1_1_4/buf_output[5] ), .Z(\SB2_1_4/i0_3 ) );
  CLKBUF_X4 U8972 ( .I(\SB1_3_24/buf_output[2] ), .Z(\SB2_3_21/i0_0 ) );
  BUF_X4 \SB1_2_3/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[169] ), .Z(
        \SB1_2_3/i0[6] ) );
  NAND3_X2 U1191 ( .A1(\SB1_2_6/i0[10] ), .A2(\SB1_2_6/i0_3 ), .A3(
        \SB1_2_6/i0[6] ), .ZN(n4438) );
  NAND3_X2 U1453 ( .A1(\SB1_1_9/i0_3 ), .A2(\SB1_1_9/i1[9] ), .A3(
        \SB1_1_9/i0_4 ), .ZN(n3936) );
  BUF_X4 \SB2_0_13/BUF_1_0  ( .I(\SB2_0_13/buf_output[1] ), .Z(\RI5[0][133] )
         );
  NAND4_X2 U1515 ( .A1(\SB2_0_13/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_0_13/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_0_13/Component_Function_1/NAND4_in[0] ), .A4(n2040), .ZN(
        \SB2_0_13/buf_output[1] ) );
  BUF_X4 U8257 ( .I(\SB2_3_2/buf_output[1] ), .Z(\RI5[3][7] ) );
  NAND3_X2 U7124 ( .A1(\SB2_3_5/i0_3 ), .A2(\SB2_3_5/i0_0 ), .A3(
        \SB2_3_5/i0[7] ), .ZN(n2397) );
  NAND2_X2 \SB1_0_28/Component_Function_5/N1  ( .A1(\SB1_0_28/i0_0 ), .A2(
        \SB1_0_28/i3[0] ), .ZN(\SB1_0_28/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB2_3_18/Component_Function_1/N4  ( .A1(\SB2_3_18/i1_7 ), .A2(
        \SB2_3_18/i0[8] ), .A3(\SB2_3_18/i0_4 ), .ZN(
        \SB2_3_18/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 U773 ( .A1(\SB1_3_20/i3[0] ), .A2(\SB1_3_20/i1_5 ), .A3(
        \SB1_3_20/i0[8] ), .ZN(n1186) );
  NAND3_X2 U1973 ( .A1(\SB2_3_4/i0_3 ), .A2(\SB2_3_4/i0[9] ), .A3(
        \SB2_3_4/i0[8] ), .ZN(n3465) );
  NAND3_X2 U1516 ( .A1(\SB2_0_7/i0_3 ), .A2(\SB2_0_7/i0_0 ), .A3(
        \SB1_0_8/buf_output[4] ), .ZN(
        \SB2_0_7/Component_Function_3/NAND4_in[1] ) );
  INV_X2 \SB1_2_6/INV_5  ( .I(\MC_ARK_ARC_1_1/buf_output[155] ), .ZN(
        \SB1_2_6/i1_5 ) );
  NAND3_X2 \SB2_3_5/Component_Function_0/N2  ( .A1(\SB2_3_5/i0[8] ), .A2(
        \SB2_3_5/i0[7] ), .A3(\SB2_3_5/i0[6] ), .ZN(
        \SB2_3_5/Component_Function_0/NAND4_in[1] ) );
  NAND3_X2 U1968 ( .A1(\SB2_0_7/i0_3 ), .A2(\SB2_0_7/i1[9] ), .A3(
        \SB1_0_8/buf_output[4] ), .ZN(n1440) );
  NAND3_X2 U794 ( .A1(\SB1_3_5/i0_0 ), .A2(\SB1_3_5/i0_4 ), .A3(\SB1_3_5/i0_3 ), .ZN(\SB1_3_5/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U831 ( .A1(\SB1_3_1/i0_0 ), .A2(\SB1_3_1/i1_5 ), .A3(\SB1_3_1/i0_4 ), .ZN(n4286) );
  NAND3_X2 \SB4_2/Component_Function_3/N1  ( .A1(\SB4_2/i1[9] ), .A2(
        \SB4_2/i0_3 ), .A3(\SB4_2/i0[6] ), .ZN(
        \SB4_2/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 \SB1_1_22/BUF_3  ( .I(\MC_ARK_ARC_1_0/buf_output[57] ), .Z(
        \SB1_1_22/i0[10] ) );
  CLKBUF_X4 U9037 ( .I(\SB1_1_5/buf_output[3] ), .Z(\SB2_1_3/i0[10] ) );
  BUF_X2 U31 ( .I(Key[172]), .Z(n165) );
  NAND3_X2 U3409 ( .A1(\SB2_0_19/i1[9] ), .A2(\SB2_0_19/i0_3 ), .A3(
        \SB2_0_19/i0[6] ), .ZN(\SB2_0_19/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U3354 ( .A1(\SB1_0_21/i0_3 ), .A2(\SB1_0_21/i0[10] ), .A3(
        \SB1_0_21/i0[6] ), .ZN(n4651) );
  NAND2_X2 \SB2_2_23/Component_Function_5/N1  ( .A1(\SB2_2_23/i0_0 ), .A2(
        \SB2_2_23/i3[0] ), .ZN(\SB2_2_23/Component_Function_5/NAND4_in[0] ) );
  INV_X2 U1845 ( .I(\MC_ARK_ARC_1_2/buf_output[134] ), .ZN(\SB1_3_9/i1[9] ) );
  NAND4_X2 U5743 ( .A1(n2546), .A2(\SB1_3_18/Component_Function_0/NAND4_in[0] ), .A3(\SB1_3_18/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_18/Component_Function_0/NAND4_in[1] ), .ZN(
        \SB1_3_18/buf_output[0] ) );
  INV_X2 U2471 ( .I(\MC_ARK_ARC_1_2/buf_output[81] ), .ZN(\SB1_3_18/i0[8] ) );
  INV_X2 U3350 ( .I(\SB1_2_31/buf_output[5] ), .ZN(\SB2_2_31/i1_5 ) );
  NAND3_X2 U1360 ( .A1(\SB1_3_15/i1[9] ), .A2(\SB1_3_15/i1_5 ), .A3(
        \SB1_3_15/i0_4 ), .ZN(\SB1_3_15/Component_Function_4/NAND4_in[3] ) );
  BUF_X4 \SB2_2_8/BUF_5  ( .I(\SB1_2_8/buf_output[5] ), .Z(\SB2_2_8/i0_3 ) );
  CLKBUF_X4 U8684 ( .I(\MC_ARK_ARC_1_3/buf_output[156] ), .Z(\SB3_5/i0[9] ) );
  BUF_X2 U86 ( .I(Key[23]), .Z(n239) );
  BUF_X4 \SB1_1_9/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[132] ), .Z(
        \SB1_1_9/i0[9] ) );
  INV_X2 \SB1_0_11/INV_3  ( .I(n381), .ZN(\SB1_0_11/i0[8] ) );
  INV_X2 U1762 ( .I(\MC_ARK_ARC_1_0/buf_output[157] ), .ZN(\SB1_1_5/i1_7 ) );
  NAND3_X2 U9221 ( .A1(\SB2_1_31/i1[9] ), .A2(\SB2_1_31/i0_4 ), .A3(n5510), 
        .ZN(n3792) );
  NAND3_X2 \SB1_1_0/Component_Function_4/N4  ( .A1(\SB1_1_0/i1[9] ), .A2(
        \SB1_1_0/i1_5 ), .A3(\SB1_1_0/i0_4 ), .ZN(
        \SB1_1_0/Component_Function_4/NAND4_in[3] ) );
  NAND3_X2 U5425 ( .A1(\SB2_3_27/i0_4 ), .A2(\SB2_3_27/i0_3 ), .A3(
        \SB2_3_27/i1[9] ), .ZN(n2320) );
  NAND3_X2 \SB2_1_5/Component_Function_2/N3  ( .A1(\SB2_1_5/i0_3 ), .A2(
        \SB2_1_5/i0[8] ), .A3(\SB2_1_5/i0[9] ), .ZN(
        \SB2_1_5/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U3044 ( .A1(\SB2_3_4/i0_3 ), .A2(\SB2_3_4/i1[9] ), .A3(
        \SB2_3_4/i0_4 ), .ZN(\SB2_3_4/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U3828 ( .A1(\SB3_15/i0_3 ), .A2(\SB3_15/i0[9] ), .A3(
        \SB3_15/i0[10] ), .ZN(\SB3_15/Component_Function_4/NAND4_in[2] ) );
  NAND3_X2 \SB2_2_30/Component_Function_2/N3  ( .A1(\SB2_2_30/i0_3 ), .A2(
        \SB2_2_30/i0[8] ), .A3(\SB2_2_30/i0[9] ), .ZN(
        \SB2_2_30/Component_Function_2/NAND4_in[2] ) );
  NAND2_X2 \SB1_3_21/Component_Function_5/N1  ( .A1(\SB1_3_21/i0_0 ), .A2(
        \SB1_3_21/i3[0] ), .ZN(\SB1_3_21/Component_Function_5/NAND4_in[0] ) );
  NAND2_X2 \SB2_3_5/Component_Function_1/N1  ( .A1(\SB2_3_5/i0_3 ), .A2(n3671), 
        .ZN(\SB2_3_5/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 U3224 ( .A1(\SB1_1_8/i0[10] ), .A2(\SB1_1_8/i0[6] ), .A3(
        \RI1[1][143] ), .ZN(n910) );
  NAND3_X2 U2100 ( .A1(\SB2_2_17/i1_5 ), .A2(\SB2_2_17/i0[10] ), .A3(
        \SB2_2_17/i1[9] ), .ZN(\SB2_2_17/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U3606 ( .A1(\SB2_2_0/i0_3 ), .A2(\SB2_2_0/i0[10] ), .A3(
        \SB2_2_0/i0[9] ), .ZN(\SB2_2_0/Component_Function_4/NAND4_in[2] ) );
  BUF_X4 U3046 ( .I(n408), .Z(\SB1_0_28/i0_3 ) );
  NAND3_X2 \SB1_1_27/Component_Function_5/N2  ( .A1(\SB1_1_27/i0_0 ), .A2(
        \SB1_1_27/i0[6] ), .A3(\SB1_1_27/i0[10] ), .ZN(
        \SB1_1_27/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U714 ( .A1(\SB2_3_16/i0[8] ), .A2(\SB2_3_16/i3[0] ), .A3(
        \SB2_3_16/i1_5 ), .ZN(\SB2_3_16/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 \SB2_2_5/Component_Function_4/N1  ( .A1(\SB2_2_5/i0[9] ), .A2(
        \SB2_2_5/i0_0 ), .A3(\SB2_2_5/i0[8] ), .ZN(
        \SB2_2_5/Component_Function_4/NAND4_in[0] ) );
  NAND3_X2 \SB1_2_18/Component_Function_4/N3  ( .A1(\SB1_2_18/i0[9] ), .A2(
        \SB1_2_18/i0[10] ), .A3(\SB1_2_18/i0_3 ), .ZN(
        \SB1_2_18/Component_Function_4/NAND4_in[2] ) );
  NAND3_X2 U6135 ( .A1(\SB1_3_21/i0[7] ), .A2(\SB1_3_21/i0[8] ), .A3(
        \SB1_3_21/i0[6] ), .ZN(\SB1_3_21/Component_Function_0/NAND4_in[1] ) );
  NAND3_X2 U790 ( .A1(\SB1_3_23/i0_3 ), .A2(\SB1_3_23/i0[6] ), .A3(
        \SB1_3_23/i1[9] ), .ZN(\SB1_3_23/Component_Function_3/NAND4_in[0] ) );
  BUF_X4 U8989 ( .I(\MC_ARK_ARC_1_2/buf_output[177] ), .Z(\SB1_3_2/i0[10] ) );
  BUF_X4 U8705 ( .I(\MC_ARK_ARC_1_3/buf_output[83] ), .Z(\SB3_18/i0_3 ) );
  NAND3_X1 \SB2_0_8/Component_Function_3/N4  ( .A1(\SB2_0_8/i1_5 ), .A2(
        \SB2_0_8/i0[8] ), .A3(\SB2_0_8/i3[0] ), .ZN(
        \SB2_0_8/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 U2131 ( .A1(\SB2_2_23/i0_3 ), .A2(\SB2_2_23/i0_4 ), .A3(
        \SB2_2_23/i1[9] ), .ZN(\SB2_2_23/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U11171 ( .A1(\SB2_3_25/i0_0 ), .A2(\SB2_3_25/i0_3 ), .A3(
        \SB1_3_26/buf_output[4] ), .ZN(
        \SB2_3_25/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U2579 ( .A1(\SB1_0_19/i0[10] ), .A2(\SB1_0_19/i0[6] ), .A3(
        \SB1_0_19/i0_3 ), .ZN(n1287) );
  INV_X2 \SB1_2_24/INV_1  ( .I(\MC_ARK_ARC_1_1/buf_output[43] ), .ZN(
        \SB1_2_24/i1_7 ) );
  NAND3_X2 \SB1_3_0/Component_Function_3/N2  ( .A1(\SB1_3_0/i0_0 ), .A2(
        \SB1_3_0/i0_3 ), .A3(\SB1_3_0/i0_4 ), .ZN(
        \SB1_3_0/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 \SB2_0_26/Component_Function_2/N3  ( .A1(\SB2_0_26/i0_3 ), .A2(
        \SB2_0_26/i0[8] ), .A3(\SB2_0_26/i0[9] ), .ZN(
        \SB2_0_26/Component_Function_2/NAND4_in[2] ) );
  NAND2_X2 \SB1_3_30/Component_Function_5/N1  ( .A1(\SB1_3_30/i0_0 ), .A2(
        \SB1_3_30/i3[0] ), .ZN(\SB1_3_30/Component_Function_5/NAND4_in[0] ) );
  INV_X2 U1511 ( .I(\MC_ARK_ARC_1_0/buf_output[33] ), .ZN(\SB1_1_26/i0[8] ) );
  INV_X2 U1677 ( .I(\SB1_1_26/buf_output[1] ), .ZN(\SB2_1_22/i1_7 ) );
  NAND3_X2 \SB1_2_23/Component_Function_4/N3  ( .A1(\SB1_2_23/i0[9] ), .A2(
        \SB1_2_23/i0[10] ), .A3(\SB1_2_23/i0_3 ), .ZN(
        \SB1_2_23/Component_Function_4/NAND4_in[2] ) );
  NAND2_X2 \SB2_0_1/Component_Function_5/N1  ( .A1(\SB2_0_1/i0_0 ), .A2(
        \SB2_0_1/i3[0] ), .ZN(\SB2_0_1/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U567 ( .A1(\SB4_2/i0[6] ), .A2(\SB4_2/i1_5 ), .A3(\SB4_2/i0[9] ), 
        .ZN(\SB4_2/Component_Function_1/NAND4_in[2] ) );
  BUF_X2 \MC_ARK_ARC_1_1/BUF_51_0  ( .I(Key[43]), .Z(
        \MC_ARK_ARC_1_1/buf_keyinput[51] ) );
  BUF_X4 \SB1_2_24/BUF_2  ( .I(\MC_ARK_ARC_1_1/buf_output[44] ), .Z(
        \SB1_2_24/i0_0 ) );
  BUF_X4 U8833 ( .I(\MC_ARK_ARC_1_2/buf_output[161] ), .Z(\SB1_3_5/i0_3 ) );
  BUF_X2 U20 ( .I(Key[51]), .Z(n199) );
  BUF_X4 \SB2_2_0/BUF_4  ( .I(\SB1_2_1/buf_output[4] ), .Z(\SB2_2_0/i0_4 ) );
  BUF_X4 \SB2_1_28/BUF_1  ( .I(\SB1_1_0/buf_output[1] ), .Z(\SB2_1_28/i0[6] )
         );
  NAND3_X2 \SB1_2_10/Component_Function_3/N3  ( .A1(\SB1_2_10/i1[9] ), .A2(
        \SB1_2_10/i1_7 ), .A3(\SB1_2_10/i0[10] ), .ZN(
        \SB1_2_10/Component_Function_3/NAND4_in[2] ) );
  BUF_X4 \SB2_1_25/BUF_0  ( .I(\SB1_1_30/buf_output[0] ), .Z(\SB2_1_25/i0[9] )
         );
  NAND3_X2 U9030 ( .A1(\SB1_1_17/i0[10] ), .A2(\SB1_1_17/i1[9] ), .A3(
        \SB1_1_17/i1_7 ), .ZN(\SB1_1_17/Component_Function_3/NAND4_in[2] ) );
  NAND2_X2 \SB2_3_31/Component_Function_5/N1  ( .A1(\SB2_3_31/i0_0 ), .A2(
        \SB2_3_31/i3[0] ), .ZN(\SB2_3_31/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U7521 ( .A1(\SB1_3_31/i0_3 ), .A2(\SB1_3_31/i0[8] ), .A3(
        \SB1_3_31/i1_7 ), .ZN(\SB1_3_31/Component_Function_1/NAND4_in[1] ) );
  AND4_X2 U569 ( .A1(n4226), .A2(n4439), .A3(
        \SB3_20/Component_Function_5/NAND4_in[1] ), .A4(n3908), .Z(n3674) );
  BUF_X4 \SB1_1_9/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[136] ), .Z(
        \SB1_1_9/i0_4 ) );
  NAND3_X2 U2099 ( .A1(\SB2_2_6/i0[10] ), .A2(\SB2_2_6/i0[6] ), .A3(
        \SB2_2_6/i0_3 ), .ZN(n1616) );
  INV_X8 \SB2_0_9/INV_2  ( .I(\RI3[0][134] ), .ZN(\SB2_0_9/i1[9] ) );
  BUF_X2 \SB2_0_24/BUF_0  ( .I(\SB1_0_29/buf_output[0] ), .Z(\SB2_0_24/i0[9] )
         );
  INV_X2 U2975 ( .I(\SB1_2_7/buf_output[5] ), .ZN(\SB2_2_7/i1_5 ) );
  NAND3_X2 U4439 ( .A1(\SB1_3_10/i0_3 ), .A2(\SB1_3_10/i1[9] ), .A3(
        \SB1_3_10/i0_4 ), .ZN(\SB1_3_10/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U3754 ( .A1(\SB1_1_20/i0_3 ), .A2(\SB1_1_20/i0[7] ), .A3(
        \SB1_1_20/i0_0 ), .ZN(n1110) );
  NAND3_X2 \SB3_20/Component_Function_4/N1  ( .A1(\SB3_20/i0[9] ), .A2(
        \SB3_20/i0_0 ), .A3(\SB3_20/i0[8] ), .ZN(
        \SB3_20/Component_Function_4/NAND4_in[0] ) );
  BUF_X4 U2714 ( .I(\MC_ARK_ARC_1_2/buf_output[65] ), .Z(\SB1_3_21/i0_3 ) );
  NAND3_X2 \SB2_0_3/Component_Function_1/N3  ( .A1(\SB2_0_3/i1_5 ), .A2(
        \SB2_0_3/i0[6] ), .A3(\SB2_0_3/i0[9] ), .ZN(
        \SB2_0_3/Component_Function_1/NAND4_in[2] ) );
  BUF_X4 \SB1_1_23/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[52] ), .Z(
        \SB1_1_23/i0_4 ) );
  NAND3_X2 U2717 ( .A1(\SB2_3_16/i0[10] ), .A2(\SB2_3_16/i1[9] ), .A3(
        \SB2_3_16/i1_7 ), .ZN(\SB2_3_16/Component_Function_3/NAND4_in[2] ) );
  BUF_X4 U3135 ( .I(\SB1_1_29/buf_output[5] ), .Z(\SB2_1_29/i0_3 ) );
  NAND3_X2 U631 ( .A1(\SB3_5/i0[8] ), .A2(\SB3_5/i1_7 ), .A3(\SB3_5/i0_4 ), 
        .ZN(\SB3_5/Component_Function_1/NAND4_in[3] ) );
  CLKBUF_X4 U1531 ( .I(\RI3[0][180] ), .Z(\SB2_0_1/i0[9] ) );
  BUF_X2 U3840 ( .I(\SB3_23/buf_output[3] ), .Z(\SB4_21/i0[10] ) );
  NAND3_X2 \SB2_1_14/Component_Function_1/N2  ( .A1(\SB2_1_14/i0_3 ), .A2(
        \SB2_1_14/i1_7 ), .A3(\SB2_1_14/i0[8] ), .ZN(
        \SB2_1_14/Component_Function_1/NAND4_in[1] ) );
  NAND3_X2 \SB2_0_10/Component_Function_1/N4  ( .A1(\SB2_0_10/i1_7 ), .A2(
        \SB2_0_10/i0[8] ), .A3(\SB2_0_10/i0_4 ), .ZN(
        \SB2_0_10/Component_Function_1/NAND4_in[3] ) );
  NAND2_X2 \SB1_1_1/Component_Function_5/N1  ( .A1(\SB1_1_1/i0_0 ), .A2(
        \SB1_1_1/i3[0] ), .ZN(\SB1_1_1/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB3_20/Component_Function_0/N4  ( .A1(\SB3_20/i0[7] ), .A2(
        \SB3_20/i0_3 ), .A3(\SB3_20/i0_0 ), .ZN(
        \SB3_20/Component_Function_0/NAND4_in[3] ) );
  NAND2_X2 \SB2_2_7/Component_Function_5/N1  ( .A1(\SB2_2_7/i0_0 ), .A2(
        \SB2_2_7/i3[0] ), .ZN(\SB2_2_7/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U2287 ( .A1(\SB2_3_30/i1[9] ), .A2(\SB2_3_30/i0_3 ), .A3(
        \SB2_3_30/i0[6] ), .ZN(\SB2_3_30/Component_Function_3/NAND4_in[0] ) );
  NAND2_X2 \SB2_2_10/Component_Function_5/N1  ( .A1(\SB2_2_10/i0_0 ), .A2(
        \SB2_2_10/i3[0] ), .ZN(\SB2_2_10/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U3616 ( .A1(\SB2_2_10/i1[9] ), .A2(\SB2_2_10/i1_7 ), .A3(
        \SB2_2_10/i0[10] ), .ZN(\SB2_2_10/Component_Function_3/NAND4_in[2] )
         );
  NAND2_X2 \SB1_2_21/Component_Function_5/N1  ( .A1(\SB1_2_21/i0_0 ), .A2(
        \SB1_2_21/i3[0] ), .ZN(\SB1_2_21/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 U951 ( .I(\MC_ARK_ARC_1_2/buf_output[141] ), .Z(\SB1_3_8/i0[10] ) );
  NAND3_X2 U1032 ( .A1(\SB2_2_15/i0_0 ), .A2(\SB2_2_15/i0_4 ), .A3(
        \SB2_2_15/i1_5 ), .ZN(\SB2_2_15/Component_Function_2/NAND4_in[3] ) );
  NAND2_X2 \SB2_3_24/Component_Function_5/N1  ( .A1(\SB2_3_24/i0_0 ), .A2(
        \SB2_3_24/i3[0] ), .ZN(\SB2_3_24/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 U2399 ( .I(\SB3_18/buf_output[5] ), .Z(\SB4_18/i0_3 ) );
  NAND3_X2 U9385 ( .A1(\SB2_3_24/i0_3 ), .A2(\SB2_3_24/i0_0 ), .A3(
        \SB2_3_24/i0_4 ), .ZN(\SB2_3_24/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U1497 ( .A1(\SB1_1_13/i0_3 ), .A2(\SB1_1_13/i0[9] ), .A3(
        \SB1_1_13/i0[8] ), .ZN(n4240) );
  NAND2_X2 U884 ( .A1(\SB1_2_16/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_2_16/Component_Function_4/NAND4_in[0] ), .ZN(n1660) );
  NAND3_X2 U1305 ( .A1(\SB2_1_24/i0_0 ), .A2(\SB2_1_24/i0_3 ), .A3(
        \SB2_1_24/i0[7] ), .ZN(n3847) );
  INV_X4 U2107 ( .I(\SB1_3_21/i0_4 ), .ZN(\SB1_3_21/i0[7] ) );
  NAND3_X2 \SB2_0_10/Component_Function_3/N4  ( .A1(\SB2_0_10/i1_5 ), .A2(
        \SB2_0_10/i0[8] ), .A3(\SB2_0_10/i3[0] ), .ZN(
        \SB2_0_10/Component_Function_3/NAND4_in[3] ) );
  BUF_X4 \SB1_3_15/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[100] ), .Z(
        \SB1_3_15/i0_4 ) );
  NAND3_X2 U1007 ( .A1(\SB1_1_24/i0_4 ), .A2(\SB1_1_24/i0[9] ), .A3(
        \SB1_1_24/i0[6] ), .ZN(\SB1_1_24/Component_Function_5/NAND4_in[3] ) );
  BUF_X4 \SB2_2_5/BUF_2  ( .I(\SB1_2_8/buf_output[2] ), .Z(\SB2_2_5/i0_0 ) );
  BUF_X4 \MC_ARK_ARC_1_2/BUF_131_1  ( .I(\MC_ARK_ARC_1_2/buf_output[131] ), 
        .Z(\RI1[3][131] ) );
  BUF_X2 U39 ( .I(Key[11]), .Z(n182) );
  BUF_X4 \SB2_1_14/BUF_1  ( .I(\SB1_1_18/buf_output[1] ), .Z(\SB2_1_14/i0[6] )
         );
  CLKBUF_X2 U30 ( .I(Key[137]), .Z(n242) );
  INV_X4 U2949 ( .I(\RI1[1][143] ), .ZN(n3647) );
  BUF_X2 \SB1_1_24/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[43] ), .Z(
        \SB1_1_24/i0[6] ) );
  BUF_X4 U3338 ( .I(n341), .Z(\SB1_0_31/i0[10] ) );
  NAND2_X2 \SB2_3_5/Component_Function_0/N1  ( .A1(\SB2_3_5/i0[10] ), .A2(
        \SB2_3_5/i0[9] ), .ZN(\SB2_3_5/Component_Function_0/NAND4_in[0] ) );
  NAND2_X2 U2377 ( .A1(\SB3_4/i0_0 ), .A2(\SB3_4/i3[0] ), .ZN(n3475) );
  INV_X4 U756 ( .I(\SB2_3_25/i0[7] ), .ZN(\SB1_3_26/buf_output[4] ) );
  NAND3_X2 U2917 ( .A1(\SB1_3_26/i1_5 ), .A2(\SB1_3_26/i1[9] ), .A3(
        \SB1_3_26/i0_4 ), .ZN(\SB1_3_26/Component_Function_4/NAND4_in[3] ) );
  BUF_X4 \SB2_2_2/BUF_5  ( .I(\SB1_2_2/buf_output[5] ), .Z(\SB2_2_2/i0_3 ) );
  NAND3_X2 \SB2_1_17/Component_Function_1/N4  ( .A1(\SB2_1_17/i1_7 ), .A2(
        \SB2_1_17/i0[8] ), .A3(\SB2_1_17/i0_4 ), .ZN(
        \SB2_1_17/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 \SB1_3_9/Component_Function_5/N4  ( .A1(\SB1_3_9/i0[9] ), .A2(
        \SB1_3_9/i0[6] ), .A3(\SB1_3_9/i0_4 ), .ZN(
        \SB1_3_9/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 U7964 ( .A1(\SB3_15/i1_5 ), .A2(\SB3_15/i1[9] ), .A3(\SB3_15/i0_4 ), 
        .ZN(\SB3_15/Component_Function_4/NAND4_in[3] ) );
  INV_X2 U1512 ( .I(\MC_ARK_ARC_1_0/buf_output[125] ), .ZN(\SB1_1_11/i1_5 ) );
  INV_X2 \SB1_0_10/INV_4  ( .I(\SB1_0_10/i0_4 ), .ZN(\SB1_0_10/i0[7] ) );
  NAND3_X2 U2022 ( .A1(\SB3_16/i0_0 ), .A2(\SB3_16/i0[6] ), .A3(
        \SB3_16/i0[10] ), .ZN(\SB3_16/Component_Function_5/NAND4_in[1] ) );
  CLKBUF_X4 U754 ( .I(\SB1_3_13/buf_output[3] ), .Z(\SB2_3_11/i0[10] ) );
  NAND3_X1 U10201 ( .A1(\SB2_2_20/i0_0 ), .A2(\SB2_2_20/i0_4 ), .A3(
        \SB2_2_20/i1_5 ), .ZN(n4202) );
  NAND4_X2 U11184 ( .A1(\SB2_0_10/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_10/Component_Function_3/NAND4_in[3] ), .A3(n4730), .A4(
        \SB2_0_10/Component_Function_3/NAND4_in[1] ), .ZN(
        \SB2_0_10/buf_output[3] ) );
  BUF_X2 U668 ( .I(\SB2_3_11/buf_output[1] ), .Z(\RI5[3][145] ) );
  NAND2_X2 U2021 ( .A1(\SB3_16/i0_0 ), .A2(\SB3_16/i3[0] ), .ZN(
        \SB3_16/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB1_1_17/Component_Function_4/N3  ( .A1(\SB1_1_17/i0[9] ), .A2(
        \SB1_1_17/i0[10] ), .A3(\SB1_1_17/i0_3 ), .ZN(
        \SB1_1_17/Component_Function_4/NAND4_in[2] ) );
  BUF_X4 U1335 ( .I(\MC_ARK_ARC_1_1/buf_output[141] ), .Z(\SB1_2_8/i0[10] ) );
  INV_X2 \SB2_1_11/INV_1  ( .I(\SB1_1_15/buf_output[1] ), .ZN(\SB2_1_11/i1_7 )
         );
  NAND2_X2 U3846 ( .A1(\SB1_0_10/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_0_10/Component_Function_4/NAND4_in[3] ), .ZN(n1144) );
  NAND3_X2 \SB2_3_25/Component_Function_3/N4  ( .A1(\SB2_3_25/i1_5 ), .A2(
        \SB2_3_25/i0[8] ), .A3(\SB2_3_25/i3[0] ), .ZN(
        \SB2_3_25/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 U3151 ( .A1(\SB2_2_16/i0[10] ), .A2(\SB2_2_16/i1_5 ), .A3(
        \SB2_2_16/i1[9] ), .ZN(\SB2_2_16/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB2_0_30/Component_Function_3/N1  ( .A1(\SB2_0_30/i1[9] ), .A2(
        \SB2_0_30/i0_3 ), .A3(\SB2_0_30/i0[6] ), .ZN(
        \SB2_0_30/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U3675 ( .A1(\SB1_3_24/i0_0 ), .A2(\SB1_3_24/i0[7] ), .A3(
        \SB1_3_24/i0_3 ), .ZN(n1805) );
  BUF_X4 \SB1_1_17/BUF_3  ( .I(\MC_ARK_ARC_1_0/buf_output[87] ), .Z(
        \SB1_1_17/i0[10] ) );
  NAND3_X2 \SB4_11/Component_Function_5/N3  ( .A1(\SB4_11/i1[9] ), .A2(
        \SB4_11/i0_4 ), .A3(\SB4_11/i0_3 ), .ZN(
        \SB4_11/Component_Function_5/NAND4_in[2] ) );
  BUF_X4 U2274 ( .I(\MC_ARK_ARC_1_2/buf_output[101] ), .Z(\SB1_3_15/i0_3 ) );
  NAND3_X2 U5173 ( .A1(\SB1_1_19/i0_4 ), .A2(\SB1_1_19/i1_5 ), .A3(
        \SB1_1_19/i1[9] ), .ZN(n1495) );
  NAND3_X2 U704 ( .A1(\SB2_3_4/i0_0 ), .A2(\SB2_3_4/i0_4 ), .A3(n5519), .ZN(
        n1896) );
  NAND3_X2 \SB2_0_0/Component_Function_2/N1  ( .A1(\SB2_0_0/i1_5 ), .A2(
        \SB2_0_0/i0[10] ), .A3(\SB2_0_0/i1[9] ), .ZN(
        \SB2_0_0/Component_Function_2/NAND4_in[0] ) );
  INV_X4 U5320 ( .I(\SB2_2_28/i0[7] ), .ZN(\SB2_2_28/i0_4 ) );
  NAND3_X2 U943 ( .A1(\SB2_1_28/i0[10] ), .A2(\SB2_1_28/i0[9] ), .A3(
        \SB2_1_28/i0_3 ), .ZN(\SB2_1_28/Component_Function_4/NAND4_in[2] ) );
  NAND3_X2 \SB1_3_11/Component_Function_3/N3  ( .A1(\SB1_3_11/i1[9] ), .A2(
        \SB1_3_11/i1_7 ), .A3(\SB1_3_11/i0[10] ), .ZN(
        \SB1_3_11/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_12/Component_Function_1/N2  ( .A1(\SB1_3_12/i0_3 ), .A2(
        \SB1_3_12/i1_7 ), .A3(\SB1_3_12/i0[8] ), .ZN(
        \SB1_3_12/Component_Function_1/NAND4_in[1] ) );
  BUF_X4 U2978 ( .I(\SB1_2_7/buf_output[5] ), .Z(\SB2_2_7/i0_3 ) );
  BUF_X4 U3078 ( .I(\MC_ARK_ARC_1_1/buf_output[50] ), .Z(\SB1_2_23/i0_0 ) );
  BUF_X4 U1815 ( .I(\SB2_3_25/buf_output[0] ), .Z(\RI5[3][66] ) );
  NAND3_X2 \SB2_0_7/Component_Function_0/N4  ( .A1(n6113), .A2(\SB2_0_7/i0_3 ), 
        .A3(\SB2_0_7/i0_0 ), .ZN(\SB2_0_7/Component_Function_0/NAND4_in[3] )
         );
  NAND3_X2 \SB2_1_13/Component_Function_3/N2  ( .A1(\SB2_1_13/i0_0 ), .A2(
        \SB2_1_13/i0_3 ), .A3(\SB2_1_13/i0_4 ), .ZN(
        \SB2_1_13/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 \SB2_0_10/Component_Function_5/N3  ( .A1(\SB2_0_10/i1[9] ), .A2(
        \SB2_0_10/i0_4 ), .A3(\SB2_0_10/i0_3 ), .ZN(
        \SB2_0_10/Component_Function_5/NAND4_in[2] ) );
  NAND2_X2 \SB2_0_14/Component_Function_1/N1  ( .A1(\SB2_0_14/i0_3 ), .A2(
        \SB2_0_14/i1[9] ), .ZN(\SB2_0_14/Component_Function_1/NAND4_in[0] ) );
  BUF_X4 U8643 ( .I(\MC_ARK_ARC_1_2/buf_output[123] ), .Z(\SB1_3_11/i0[10] )
         );
  NAND3_X2 U8845 ( .A1(\SB2_3_4/i0_3 ), .A2(\SB2_3_4/i0[10] ), .A3(
        \SB2_3_4/i0[6] ), .ZN(\SB2_3_4/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 U8913 ( .I(\RI1[4][53] ), .Z(\SB3_23/i0_3 ) );
  CLKBUF_X4 \SB2_0_13/BUF_1  ( .I(\SB1_0_17/buf_output[1] ), .Z(
        \SB2_0_13/i0[6] ) );
  BUF_X2 U1904 ( .I(\SB1_1_11/buf_output[0] ), .Z(\SB2_1_6/i0[9] ) );
  NAND3_X2 \SB1_3_11/Component_Function_3/N2  ( .A1(\SB1_3_11/i0_0 ), .A2(
        \SB1_3_11/i0_3 ), .A3(\SB1_3_11/i0_4 ), .ZN(
        \SB1_3_11/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U851 ( .A1(\SB1_3_16/i0[10] ), .A2(\SB1_3_16/i0[6] ), .A3(
        \SB1_3_16/i0_0 ), .ZN(n4203) );
  NAND3_X2 U2340 ( .A1(\SB2_3_16/i0_3 ), .A2(\SB2_3_16/i0[8] ), .A3(
        \SB2_3_16/i0[9] ), .ZN(\SB2_3_16/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U2486 ( .A1(\SB1_3_18/i0_0 ), .A2(\SB1_3_18/i0[10] ), .A3(
        \SB1_3_18/i0[6] ), .ZN(\SB1_3_18/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 U9050 ( .I(\MC_ARK_ARC_1_1/buf_output[153] ), .Z(\SB1_2_6/i0[10] ) );
  BUF_X4 U8199 ( .I(\SB2_2_26/buf_output[1] ), .Z(\RI5[2][55] ) );
  NAND4_X2 U9314 ( .A1(\SB2_2_26/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_2_26/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_2_26/Component_Function_1/NAND4_in[1] ), .A4(
        \SB2_2_26/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_2_26/buf_output[1] ) );
  INV_X2 \SB2_3_18/INV_1  ( .I(\SB1_3_22/buf_output[1] ), .ZN(\SB2_3_18/i1_7 )
         );
  INV_X2 U2921 ( .I(\MC_ARK_ARC_1_2/buf_output[62] ), .ZN(\SB1_3_21/i1[9] ) );
  NAND3_X2 U2213 ( .A1(\SB2_3_25/i0[10] ), .A2(\SB2_3_25/i1_7 ), .A3(
        \SB2_3_25/i1[9] ), .ZN(n4207) );
  NAND2_X2 U8888 ( .A1(\SB3_12/i0_0 ), .A2(\SB3_12/i3[0] ), .ZN(n1613) );
  NAND3_X2 U2025 ( .A1(\SB2_1_7/i0_3 ), .A2(\SB2_1_7/i0[10] ), .A3(n2852), 
        .ZN(\SB2_1_7/Component_Function_2/NAND4_in[1] ) );
  INV_X2 \SB1_1_27/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[25] ), .ZN(
        \SB1_1_27/i1_7 ) );
  BUF_X4 \MC_ARK_ARC_1_0/BUF_141  ( .I(\SB2_0_10/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[141] ) );
  NAND3_X2 U1739 ( .A1(\SB1_1_27/i1_5 ), .A2(\SB1_1_27/i0[6] ), .A3(
        \SB1_1_27/i0[9] ), .ZN(\SB1_1_27/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 U9250 ( .A1(\SB1_3_15/i0[8] ), .A2(\SB1_3_15/i0_4 ), .A3(
        \SB1_3_15/i1_7 ), .ZN(n3849) );
  NAND3_X2 U9619 ( .A1(n3932), .A2(\SB2_3_11/Component_Function_0/NAND4_in[1] ), .A3(\SB2_3_11/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB2_3_11/buf_output[0] ) );
  NAND2_X2 \SB1_1_7/Component_Function_5/N1  ( .A1(\SB1_1_7/i0_0 ), .A2(
        \SB1_1_7/i3[0] ), .ZN(\SB1_1_7/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB1_2_2/Component_Function_4/N3  ( .A1(\SB1_2_2/i0[9] ), .A2(
        \SB1_2_2/i0[10] ), .A3(\SB1_2_2/i0_3 ), .ZN(
        \SB1_2_2/Component_Function_4/NAND4_in[2] ) );
  NAND3_X2 \SB2_1_11/Component_Function_5/N3  ( .A1(\SB2_1_11/i1[9] ), .A2(
        \SB1_1_12/buf_output[4] ), .A3(\SB2_1_11/i0_3 ), .ZN(
        \SB2_1_11/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U1600 ( .A1(\SB2_0_9/i0_3 ), .A2(\SB2_0_9/i0[10] ), .A3(
        \SB2_0_9/i0[6] ), .ZN(n4373) );
  NAND2_X2 \SB1_0_13/Component_Function_5/N1  ( .A1(\SB1_0_13/i0_0 ), .A2(
        \SB1_0_13/i3[0] ), .ZN(\SB1_0_13/Component_Function_5/NAND4_in[0] ) );
  BUF_X2 U2365 ( .I(\SB3_13/buf_output[3] ), .Z(\SB4_11/i0[10] ) );
  NAND3_X2 U8889 ( .A1(\SB3_12/i0_0 ), .A2(\SB3_12/i0[6] ), .A3(
        \SB3_12/i0[10] ), .ZN(\SB3_12/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U11018 ( .A1(\SB1_1_27/i0_3 ), .A2(\SB1_1_27/i0[6] ), .A3(
        \SB1_1_27/i1[9] ), .ZN(\SB1_1_27/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U1266 ( .A1(\SB2_1_14/i3[0] ), .A2(\SB2_1_14/i0[8] ), .A3(
        \SB2_1_14/i1_5 ), .ZN(n3080) );
  INV_X2 U10888 ( .I(\SB1_2_26/buf_output[5] ), .ZN(\SB2_2_26/i1_5 ) );
  NAND3_X2 U1035 ( .A1(\SB2_2_17/i0[6] ), .A2(\SB2_2_17/i0[9] ), .A3(
        \SB2_2_17/i1_5 ), .ZN(\SB2_2_17/Component_Function_1/NAND4_in[2] ) );
  BUF_X4 \SB2_2_22/BUF_3  ( .I(\SB1_2_24/buf_output[3] ), .Z(\SB2_2_22/i0[10] ) );
  NAND3_X2 U2737 ( .A1(\SB1_1_1/i0[10] ), .A2(\SB1_1_1/i0[6] ), .A3(
        \SB1_1_1/i0_3 ), .ZN(n3386) );
  BUF_X4 \SB1_2_4/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[163] ), .Z(
        \SB1_2_4/i0[6] ) );
  NAND3_X2 U1445 ( .A1(\SB1_1_2/i0[10] ), .A2(\SB1_1_2/i0[6] ), .A3(
        \SB1_1_2/i0_0 ), .ZN(n1742) );
  BUF_X4 U8931 ( .I(\SB1_1_7/buf_output[5] ), .Z(\SB2_1_7/i0_3 ) );
  BUF_X4 U4832 ( .I(\MC_ARK_ARC_1_0/buf_output[152] ), .Z(\SB1_1_6/i0_0 ) );
  CLKBUF_X4 U5275 ( .I(\SB2_3_7/buf_output[2] ), .Z(\RI5[3][164] ) );
  BUF_X4 \SB2_0_4/BUF_3  ( .I(\RI3[0][165] ), .Z(\SB2_0_4/i0[10] ) );
  BUF_X4 \SB2_1_20/BUF_4  ( .I(\SB1_1_21/buf_output[4] ), .Z(\SB2_1_20/i0_4 )
         );
  CLKBUF_X4 U758 ( .I(\SB1_3_9/buf_output[3] ), .Z(\SB2_3_7/i0[10] ) );
  BUF_X2 U135 ( .I(Key[136]), .Z(n66) );
  NAND3_X2 U10295 ( .A1(\SB1_1_6/i0[8] ), .A2(\SB1_1_6/i1_5 ), .A3(
        \SB1_1_6/i3[0] ), .ZN(n2700) );
  NAND2_X2 \SB1_2_24/Component_Function_1/N1  ( .A1(\RI1[2][47] ), .A2(
        \SB1_2_24/i1[9] ), .ZN(\SB1_2_24/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 U1474 ( .A1(\SB1_1_1/i0_0 ), .A2(\SB1_1_1/i0_4 ), .A3(
        \SB1_1_1/i1_5 ), .ZN(n1906) );
  NAND3_X2 \SB2_2_22/Component_Function_2/N1  ( .A1(\SB2_2_22/i1_5 ), .A2(
        \SB2_2_22/i0[10] ), .A3(\SB2_2_22/i1[9] ), .ZN(
        \SB2_2_22/Component_Function_2/NAND4_in[0] ) );
  NAND2_X2 \SB1_1_14/Component_Function_5/N1  ( .A1(\SB1_1_14/i0_0 ), .A2(
        \SB1_1_14/i3[0] ), .ZN(\SB1_1_14/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U8930 ( .A1(\SB2_3_16/i0_3 ), .A2(\SB2_3_16/i1[9] ), .A3(
        \SB2_3_16/i0_4 ), .ZN(\SB2_3_16/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U10635 ( .A1(\SB1_2_24/i0[10] ), .A2(\SB1_2_24/i1[9] ), .A3(
        \SB1_2_24/i1_7 ), .ZN(n4413) );
  NAND3_X2 U672 ( .A1(\SB2_3_25/i0_0 ), .A2(\SB2_3_25/i0[10] ), .A3(
        \SB2_3_25/i0[6] ), .ZN(n2940) );
  BUF_X4 U1863 ( .I(\SB2_2_24/buf_output[2] ), .Z(\RI5[2][62] ) );
  NAND2_X2 \SB2_2_15/Component_Function_5/N1  ( .A1(\SB2_2_15/i0_0 ), .A2(
        \SB2_2_15/i3[0] ), .ZN(\SB2_2_15/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB1_1_1/Component_Function_2/N3  ( .A1(\SB1_1_1/i0_3 ), .A2(
        \SB1_1_1/i0[8] ), .A3(\SB1_1_1/i0[9] ), .ZN(
        \SB1_1_1/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U955 ( .A1(\SB2_1_31/i0[9] ), .A2(\SB2_1_31/i0_3 ), .A3(
        \SB2_1_31/i0[8] ), .ZN(n597) );
  BUF_X4 \SB2_1_23/BUF_4  ( .I(\SB1_1_24/buf_output[4] ), .Z(\SB2_1_23/i0_4 )
         );
  NAND3_X2 U1280 ( .A1(\SB2_1_27/i0[10] ), .A2(\SB2_1_27/i0_3 ), .A3(
        \SB2_1_27/i0[6] ), .ZN(n3840) );
  NAND3_X2 U1452 ( .A1(\SB1_1_17/i0[9] ), .A2(\SB1_1_17/i1_5 ), .A3(
        \SB1_1_17/i0[6] ), .ZN(n3941) );
  NAND3_X2 U2511 ( .A1(\SB2_2_12/i0[10] ), .A2(\SB2_2_12/i0_0 ), .A3(
        \SB2_2_12/i0[6] ), .ZN(\SB2_2_12/Component_Function_5/NAND4_in[1] ) );
  INV_X4 U7658 ( .I(\RI3[0][147] ), .ZN(\SB2_0_7/i0[8] ) );
  BUF_X4 U1237 ( .I(\MC_ARK_ARC_1_1/buf_output[107] ), .Z(\SB1_2_14/i0_3 ) );
  NAND2_X2 \SB2_1_16/Component_Function_5/N1  ( .A1(\SB2_1_16/i0_0 ), .A2(
        \SB2_1_16/i3[0] ), .ZN(\SB2_1_16/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB1_1_2/Component_Function_5/N4  ( .A1(\SB1_1_2/i0[9] ), .A2(
        \SB1_1_2/i0[6] ), .A3(\SB1_1_2/i0_4 ), .ZN(
        \SB1_1_2/Component_Function_5/NAND4_in[3] ) );
  CLKBUF_X4 \SB1_3_15/BUF_3  ( .I(\MC_ARK_ARC_1_2/buf_output[99] ), .Z(
        \SB1_3_15/i0[10] ) );
  CLKBUF_X4 U4928 ( .I(\MC_ARK_ARC_1_2/buf_output[111] ), .Z(\SB1_3_13/i0[10] ) );
  NAND3_X2 U2685 ( .A1(\SB2_3_19/i0[10] ), .A2(\SB2_3_19/i0_0 ), .A3(
        \SB2_3_19/i0[6] ), .ZN(\SB2_3_19/Component_Function_5/NAND4_in[1] ) );
  BUF_X4 U7833 ( .I(\SB2_0_29/buf_output[3] ), .Z(\RI5[0][27] ) );
  INV_X2 U8793 ( .I(\MC_ARK_ARC_1_2/buf_output[117] ), .ZN(\SB1_3_12/i0[8] )
         );
  NAND3_X2 U3853 ( .A1(\SB1_2_31/i0[6] ), .A2(\SB1_2_31/i0[9] ), .A3(
        \SB1_2_31/i0_4 ), .ZN(n1444) );
  NAND3_X2 \SB3_4/Component_Function_3/N2  ( .A1(\SB3_4/i0_0 ), .A2(
        \SB3_4/i0_3 ), .A3(\SB3_4/i0_4 ), .ZN(
        \SB3_4/Component_Function_3/NAND4_in[1] ) );
  NAND2_X2 \SB2_1_2/Component_Function_0/N1  ( .A1(\SB2_1_2/i0[10] ), .A2(
        \SB2_1_2/i0[9] ), .ZN(\SB2_1_2/Component_Function_0/NAND4_in[0] ) );
  NAND3_X2 \SB1_2_11/Component_Function_3/N2  ( .A1(\SB1_2_11/i0_0 ), .A2(
        \SB1_2_11/i0_3 ), .A3(\SB1_2_11/i0_4 ), .ZN(
        \SB1_2_11/Component_Function_3/NAND4_in[1] ) );
  INV_X2 U4715 ( .I(n334), .ZN(\SB1_0_2/i1[9] ) );
  BUF_X4 \SB4_20/BUF_5  ( .I(\SB3_20/buf_output[5] ), .Z(\SB4_20/i0_3 ) );
  INV_X2 \SB2_2_10/INV_1  ( .I(\SB1_2_14/buf_output[1] ), .ZN(\SB2_2_10/i1_7 )
         );
  INV_X2 \SB2_2_31/INV_0  ( .I(\SB1_2_4/buf_output[0] ), .ZN(\SB2_2_31/i3[0] )
         );
  NAND2_X2 U1117 ( .A1(\SB1_0_2/i0_0 ), .A2(\SB1_0_2/i3[0] ), .ZN(n1715) );
  BUF_X4 U4445 ( .I(\SB1_1_22/buf_output[3] ), .Z(\SB2_1_20/i0[10] ) );
  INV_X2 \SB2_2_31/INV_1  ( .I(\SB1_2_3/buf_output[1] ), .ZN(\SB2_2_31/i1_7 )
         );
  NAND3_X2 U3594 ( .A1(\SB2_2_12/i1_5 ), .A2(\SB2_2_12/i0[6] ), .A3(
        \SB2_2_12/i0[9] ), .ZN(\SB2_2_12/Component_Function_1/NAND4_in[2] ) );
  INV_X4 U7389 ( .I(n2564), .ZN(\SB1_3_1/buf_output[4] ) );
  NAND3_X2 \SB2_1_27/Component_Function_3/N2  ( .A1(\SB2_1_27/i0_0 ), .A2(
        \SB2_1_27/i0_3 ), .A3(\SB2_1_27/i0_4 ), .ZN(
        \SB2_1_27/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U1272 ( .A1(\SB2_1_4/i0_3 ), .A2(\SB2_1_4/i0[10] ), .A3(
        \SB2_1_4/i0[9] ), .ZN(\SB2_1_4/Component_Function_4/NAND4_in[2] ) );
  NAND3_X2 U3574 ( .A1(n2593), .A2(\SB2_0_7/i0_3 ), .A3(\SB2_0_7/i0[10] ), 
        .ZN(\SB2_0_7/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U4455 ( .A1(\SB1_1_16/i0[9] ), .A2(\SB1_1_16/i0_3 ), .A3(
        \SB1_1_16/i0[10] ), .ZN(n1956) );
  NAND2_X2 \SB2_2_26/Component_Function_5/N1  ( .A1(\SB2_2_26/i0_0 ), .A2(
        \SB2_2_26/i3[0] ), .ZN(\SB2_2_26/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB2_2_26/Component_Function_0/N4  ( .A1(\SB2_2_26/i0[7] ), .A2(
        \SB2_2_26/i0_3 ), .A3(\SB2_2_26/i0_0 ), .ZN(
        \SB2_2_26/Component_Function_0/NAND4_in[3] ) );
  BUF_X4 U8644 ( .I(\SB1_3_11/buf_output[1] ), .Z(n1670) );
  BUF_X4 U3418 ( .I(\SB1_1_4/buf_output[1] ), .Z(\SB2_1_0/i0[6] ) );
  NAND3_X2 \SB2_2_5/Component_Function_1/N2  ( .A1(\SB2_2_5/i0_3 ), .A2(
        \SB2_2_5/i1_7 ), .A3(\SB2_2_5/i0[8] ), .ZN(
        \SB2_2_5/Component_Function_1/NAND4_in[1] ) );
  NAND3_X2 \SB2_0_22/Component_Function_1/N4  ( .A1(\SB2_0_22/i1_7 ), .A2(
        \SB2_0_22/i0[8] ), .A3(\SB2_0_22/i0_4 ), .ZN(
        \SB2_0_22/Component_Function_1/NAND4_in[3] ) );
  NAND2_X2 \SB1_1_18/Component_Function_5/N1  ( .A1(\SB1_1_18/i0_0 ), .A2(
        \SB1_1_18/i3[0] ), .ZN(\SB1_1_18/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U2032 ( .A1(\SB2_1_18/i0[10] ), .A2(\SB2_1_18/i0[9] ), .A3(
        \SB2_1_18/i0_3 ), .ZN(\SB2_1_18/Component_Function_4/NAND4_in[2] ) );
  NAND3_X2 U2523 ( .A1(\SB2_3_2/i0[10] ), .A2(\SB2_3_2/i0_3 ), .A3(
        \SB2_3_2/i0[9] ), .ZN(n679) );
  NAND3_X2 U9317 ( .A1(\SB2_2_5/i0[6] ), .A2(\SB2_2_5/i0_3 ), .A3(
        \SB2_2_5/i1[9] ), .ZN(n3793) );
  BUF_X4 \SB1_1_27/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[25] ), .Z(
        \SB1_1_27/i0[6] ) );
  BUF_X2 \SB4_17/BUF_1  ( .I(\SB3_21/buf_output[1] ), .Z(\SB4_17/i0[6] ) );
  CLKBUF_X4 U3231 ( .I(\SB2_3_21/buf_output[5] ), .Z(\RI5[3][65] ) );
  BUF_X2 U117 ( .I(Key[98]), .Z(n154) );
  BUF_X4 U3599 ( .I(\SB1_2_26/buf_output[1] ), .Z(\SB2_2_22/i0[6] ) );
  NAND2_X2 U1287 ( .A1(\SB1_3_22/i0_0 ), .A2(\SB1_3_22/i3[0] ), .ZN(
        \SB1_3_22/Component_Function_5/NAND4_in[0] ) );
  NAND4_X2 U2245 ( .A1(\SB4_17/Component_Function_1/NAND4_in[2] ), .A2(
        \SB4_17/Component_Function_1/NAND4_in[1] ), .A3(
        \SB4_17/Component_Function_1/NAND4_in[0] ), .A4(
        \SB4_17/Component_Function_1/NAND4_in[3] ), .ZN(n3179) );
  NAND4_X2 \SB2_3_30/Component_Function_1/N5  ( .A1(
        \SB2_3_30/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_30/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_30/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_3_30/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_3_30/buf_output[1] ) );
  NAND3_X2 \SB3_26/Component_Function_0/N4  ( .A1(\SB3_26/i0[7] ), .A2(
        \SB3_26/i0_3 ), .A3(\SB3_26/i0_0 ), .ZN(
        \SB3_26/Component_Function_0/NAND4_in[3] ) );
  NAND3_X2 \SB2_0_13/Component_Function_2/N3  ( .A1(\SB2_0_13/i0_3 ), .A2(
        n1393), .A3(\SB1_0_18/buf_output[0] ), .ZN(
        \SB2_0_13/Component_Function_2/NAND4_in[2] ) );
  NAND2_X2 \SB1_3_14/Component_Function_5/N1  ( .A1(\SB1_3_14/i0_0 ), .A2(
        \SB1_3_14/i3[0] ), .ZN(\SB1_3_14/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB2_0_13/Component_Function_3/N4  ( .A1(n3663), .A2(n1393), .A3(
        \SB2_0_13/i3[0] ), .ZN(\SB2_0_13/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 U3534 ( .A1(\SB1_2_16/i0[9] ), .A2(\SB1_2_16/i0_0 ), .A3(
        \SB1_2_16/i0[8] ), .ZN(\SB1_2_16/Component_Function_4/NAND4_in[0] ) );
  NAND3_X2 U1951 ( .A1(\SB1_0_25/i1_5 ), .A2(\SB1_0_25/i0[10] ), .A3(
        \SB1_0_25/i1[9] ), .ZN(\SB1_0_25/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB1_3_28/Component_Function_5/N2  ( .A1(\SB1_3_28/i0_0 ), .A2(
        \SB1_3_28/i0[6] ), .A3(\SB1_3_28/i0[10] ), .ZN(
        \SB1_3_28/Component_Function_5/NAND4_in[1] ) );
  NAND2_X2 U1418 ( .A1(n1493), .A2(\SB1_1_22/Component_Function_2/NAND4_in[3] ), .ZN(n4247) );
  NAND3_X2 U2645 ( .A1(\SB1_0_26/i0[9] ), .A2(\SB1_0_26/i0[10] ), .A3(
        \SB1_0_26/i0_3 ), .ZN(\SB1_0_26/Component_Function_4/NAND4_in[2] ) );
  INV_X2 \SB2_0_2/INV_5  ( .I(\RI3[0][179] ), .ZN(\SB2_0_2/i1_5 ) );
  INV_X4 U2739 ( .I(\SB2_3_28/i0[7] ), .ZN(n577) );
  BUF_X2 U49 ( .I(Key[166]), .Z(n140) );
  NAND4_X1 \SB2_3_19/Component_Function_1/N5  ( .A1(
        \SB2_3_19/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_19/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_19/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_3_19/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_3_19/buf_output[1] ) );
  INV_X2 \SB4_1/INV_2  ( .I(\SB3_4/buf_output[2] ), .ZN(\SB4_1/i1[9] ) );
  NAND2_X2 \SB2_1_13/Component_Function_0/N1  ( .A1(\SB2_1_13/i0[10] ), .A2(
        \SB1_1_18/buf_output[0] ), .ZN(
        \SB2_1_13/Component_Function_0/NAND4_in[0] ) );
  NAND3_X2 \SB2_0_17/Component_Function_2/N2  ( .A1(\SB2_0_17/i0_3 ), .A2(
        \SB2_0_17/i0[10] ), .A3(\SB2_0_17/i0[6] ), .ZN(
        \SB2_0_17/Component_Function_2/NAND4_in[1] ) );
  INV_X2 U1323 ( .I(\MC_ARK_ARC_1_3/buf_output[135] ), .ZN(\SB3_9/i0[8] ) );
  INV_X2 U3164 ( .I(\RI3[0][139] ), .ZN(\SB2_0_8/i1_7 ) );
  NAND3_X2 \SB2_1_4/Component_Function_3/N1  ( .A1(n3660), .A2(\SB2_1_4/i0_3 ), 
        .A3(\SB2_1_4/i0[6] ), .ZN(\SB2_1_4/Component_Function_3/NAND4_in[0] )
         );
  NAND3_X2 U6876 ( .A1(\SB2_1_27/i0_0 ), .A2(\SB2_1_27/i1_5 ), .A3(
        \SB2_1_27/i0_4 ), .ZN(n2283) );
  NAND3_X2 U996 ( .A1(\SB1_1_28/i0[10] ), .A2(\SB1_1_28/i0_3 ), .A3(
        \SB1_1_28/i0[9] ), .ZN(\SB1_1_28/Component_Function_4/NAND4_in[2] ) );
  NAND3_X2 U2126 ( .A1(\SB2_2_23/i0[10] ), .A2(\SB2_2_23/i1_5 ), .A3(
        \SB2_2_23/i1[9] ), .ZN(\SB2_2_23/Component_Function_2/NAND4_in[0] ) );
  BUF_X2 U41 ( .I(Key[86]), .Z(n126) );
  NAND3_X2 \SB1_1_26/Component_Function_5/N2  ( .A1(\SB1_1_26/i0_0 ), .A2(
        \SB1_1_26/i0[6] ), .A3(\SB1_1_26/i0[10] ), .ZN(
        \SB1_1_26/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U1364 ( .A1(\SB2_1_23/i0[10] ), .A2(\SB2_1_23/i1[9] ), .A3(
        \SB2_1_23/i1_7 ), .ZN(\SB2_1_23/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U2909 ( .A1(\SB1_1_26/i0[10] ), .A2(\SB1_1_26/i1[9] ), .A3(
        \SB1_1_26/i1_5 ), .ZN(n2405) );
  NAND2_X2 \SB2_3_23/Component_Function_1/N1  ( .A1(\SB2_3_23/i0_3 ), .A2(
        \SB2_3_23/i1[9] ), .ZN(\SB2_3_23/Component_Function_1/NAND4_in[0] ) );
  BUF_X4 U8646 ( .I(\SB1_3_18/buf_output[4] ), .Z(\SB2_3_17/i0_4 ) );
  BUF_X2 U103 ( .I(Key[32]), .Z(n227) );
  INV_X2 U4872 ( .I(\SB3_8/buf_output[2] ), .ZN(\SB4_5/i1[9] ) );
  NAND3_X2 U576 ( .A1(\SB4_31/i0_0 ), .A2(\SB4_31/i1_7 ), .A3(\SB4_31/i3[0] ), 
        .ZN(n2428) );
  NAND2_X2 \SB2_1_8/Component_Function_5/N1  ( .A1(\SB2_1_8/i0_0 ), .A2(
        \SB2_1_8/i3[0] ), .ZN(\SB2_1_8/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB1_3_0/Component_Function_3/N1  ( .A1(\SB1_3_0/i1[9] ), .A2(
        \SB1_3_0/i0_3 ), .A3(\SB1_3_0/i0[6] ), .ZN(
        \SB1_3_0/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 \SB2_2_28/Component_Function_3/N1  ( .A1(\SB2_2_28/i1[9] ), .A2(
        \SB2_2_28/i0_3 ), .A3(\SB2_2_28/i0[6] ), .ZN(
        \SB2_2_28/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U6365 ( .A1(\SB2_3_30/i0_3 ), .A2(\SB2_3_30/i0[6] ), .A3(
        \SB2_3_30/i0[10] ), .ZN(\SB2_3_30/Component_Function_2/NAND4_in[1] )
         );
  NAND3_X2 U6251 ( .A1(\SB2_1_28/i0[6] ), .A2(\SB2_1_28/i0_4 ), .A3(
        \SB2_1_28/i0[9] ), .ZN(\SB2_1_28/Component_Function_5/NAND4_in[3] ) );
  INV_X2 U4452 ( .I(n5499), .ZN(\SB3_9/i1[9] ) );
  NAND2_X2 \SB1_2_23/Component_Function_5/N1  ( .A1(\SB1_2_23/i0_0 ), .A2(
        \SB1_2_23/i3[0] ), .ZN(\SB1_2_23/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U2631 ( .A1(\SB2_2_29/i0_3 ), .A2(\SB2_2_29/i0_0 ), .A3(
        \SB2_2_29/i0[7] ), .ZN(n1662) );
  NAND3_X2 U1096 ( .A1(\SB1_2_29/i0[9] ), .A2(\SB1_2_29/i0[6] ), .A3(
        \SB1_2_29/i0_4 ), .ZN(n4288) );
  INV_X2 U4507 ( .I(\MC_ARK_ARC_1_3/buf_output[137] ), .ZN(\SB3_9/i1_5 ) );
  NAND3_X2 U5056 ( .A1(\SB1_3_0/i0[8] ), .A2(\SB1_3_0/i3[0] ), .A3(
        \SB1_3_0/i1_5 ), .ZN(\SB1_3_0/Component_Function_3/NAND4_in[3] ) );
  NAND4_X2 U6383 ( .A1(\SB4_7/Component_Function_1/NAND4_in[2] ), .A2(
        \SB4_7/Component_Function_1/NAND4_in[1] ), .A3(
        \SB4_7/Component_Function_1/NAND4_in[3] ), .A4(
        \SB4_7/Component_Function_1/NAND4_in[0] ), .ZN(n2450) );
  NAND3_X2 U1388 ( .A1(\SB1_1_11/i1[9] ), .A2(\SB1_1_11/i0_4 ), .A3(
        \SB1_1_11/i0_3 ), .ZN(\SB1_1_11/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U2822 ( .A1(\SB3_18/i0_4 ), .A2(\SB3_18/i1[9] ), .A3(\SB3_18/i0_3 ), 
        .ZN(\SB3_18/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U1532 ( .A1(\SB2_0_24/i0[10] ), .A2(\SB2_0_24/i0_0 ), .A3(
        \RI3[0][43] ), .ZN(n2178) );
  BUF_X4 \SB1_3_27/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[28] ), .Z(
        \SB1_3_27/i0_4 ) );
  BUF_X4 \SB1_1_31/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[4] ), .Z(
        \SB1_1_31/i0_4 ) );
  BUF_X2 U106 ( .I(Key[112]), .Z(n148) );
  NAND3_X1 U5127 ( .A1(\SB2_3_20/i0_4 ), .A2(\SB2_3_20/i1_5 ), .A3(
        \SB2_3_20/i0_0 ), .ZN(n3433) );
  NAND3_X2 U1130 ( .A1(\SB1_0_29/i0[10] ), .A2(\SB1_0_29/i1[9] ), .A3(
        \SB1_0_29/i1_7 ), .ZN(n1277) );
  NAND3_X2 U2577 ( .A1(\SB1_0_19/i0_0 ), .A2(\SB1_0_19/i0[6] ), .A3(
        \SB1_0_19/i0[10] ), .ZN(\SB1_0_19/Component_Function_5/NAND4_in[1] )
         );
  INV_X2 U1565 ( .I(\MC_ARK_ARC_1_3/buf_output[123] ), .ZN(\SB3_11/i0[8] ) );
  NAND3_X1 U800 ( .A1(\SB1_3_30/i0_0 ), .A2(\SB1_3_30/i0[6] ), .A3(
        \SB1_3_30/i0[10] ), .ZN(\SB1_3_30/Component_Function_5/NAND4_in[1] )
         );
  NAND3_X2 U3485 ( .A1(\SB2_1_7/i1[9] ), .A2(\SB2_1_7/i1_7 ), .A3(
        \SB2_1_7/i0[10] ), .ZN(\SB2_1_7/Component_Function_3/NAND4_in[2] ) );
  NAND2_X2 \SB2_1_20/Component_Function_0/N1  ( .A1(\SB2_1_20/i0[10] ), .A2(
        \SB2_1_20/i0[9] ), .ZN(\SB2_1_20/Component_Function_0/NAND4_in[0] ) );
  NAND3_X2 U2334 ( .A1(\SB1_3_21/i0[10] ), .A2(\SB1_3_21/i1[9] ), .A3(
        \SB1_3_21/i1_7 ), .ZN(n1663) );
  NAND3_X2 \SB2_1_7/Component_Function_2/N1  ( .A1(\SB2_1_7/i1_5 ), .A2(
        \SB2_1_7/i0[10] ), .A3(\SB2_1_7/i1[9] ), .ZN(
        \SB2_1_7/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB2_1_7/Component_Function_3/N1  ( .A1(\SB2_1_7/i1[9] ), .A2(
        \SB2_1_7/i0_3 ), .A3(n2852), .ZN(
        \SB2_1_7/Component_Function_3/NAND4_in[0] ) );
  INV_X2 U2550 ( .I(\MC_ARK_ARC_1_3/buf_output[158] ), .ZN(\SB3_5/i1[9] ) );
  NAND3_X2 \SB2_2_18/Component_Function_1/N3  ( .A1(n4769), .A2(
        \SB2_2_18/i0[6] ), .A3(\SB2_2_18/i0[9] ), .ZN(
        \SB2_2_18/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 \SB1_2_8/Component_Function_3/N1  ( .A1(\SB1_2_8/i1[9] ), .A2(
        \SB1_2_8/i0_3 ), .A3(\SB1_2_8/i0[6] ), .ZN(
        \SB1_2_8/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 \SB2_2_6/Component_Function_3/N4  ( .A1(\SB2_2_6/i1_5 ), .A2(
        \SB2_2_6/i0[8] ), .A3(\SB2_2_6/i3[0] ), .ZN(
        \SB2_2_6/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 U6045 ( .A1(\SB2_2_24/i0_3 ), .A2(\SB2_2_24/i0[6] ), .A3(
        \SB2_2_24/i1[9] ), .ZN(\SB2_2_24/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U6219 ( .A1(\SB1_3_11/i0[8] ), .A2(n2908), .A3(\SB1_3_11/i3[0] ), 
        .ZN(n4377) );
  NAND3_X2 \SB2_1_17/Component_Function_3/N2  ( .A1(\SB2_1_17/i0_0 ), .A2(
        \SB2_1_17/i0_3 ), .A3(\SB2_1_17/i0_4 ), .ZN(
        \SB2_1_17/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 \SB2_2_2/Component_Function_3/N2  ( .A1(\SB2_2_2/i0_0 ), .A2(
        \SB2_2_2/i0_3 ), .A3(\SB2_2_2/i0_4 ), .ZN(
        \SB2_2_2/Component_Function_3/NAND4_in[1] ) );
  INV_X2 U9012 ( .I(\MC_ARK_ARC_1_2/buf_output[152] ), .ZN(\SB1_3_6/i1[9] ) );
  NAND3_X2 \SB1_2_14/Component_Function_1/N3  ( .A1(\SB1_2_14/i1_5 ), .A2(
        \SB1_2_14/i0[6] ), .A3(\SB1_2_14/i0[9] ), .ZN(
        \SB1_2_14/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 U3115 ( .A1(\SB1_3_21/i0_0 ), .A2(\SB1_3_21/i0[6] ), .A3(
        \SB1_3_21/i0[10] ), .ZN(\SB1_3_21/Component_Function_5/NAND4_in[1] )
         );
  NAND2_X2 U2580 ( .A1(\SB1_0_19/i0[10] ), .A2(\SB1_0_19/i0[9] ), .ZN(
        \SB1_0_19/Component_Function_0/NAND4_in[0] ) );
  CLKBUF_X4 \SB4_0/BUF_3  ( .I(\SB3_2/buf_output[3] ), .Z(\SB4_0/i0[10] ) );
  NAND3_X2 \SB2_2_2/Component_Function_1/N2  ( .A1(\SB2_2_2/i0_3 ), .A2(
        \SB2_2_2/i1_7 ), .A3(\SB2_2_2/i0[8] ), .ZN(
        \SB2_2_2/Component_Function_1/NAND4_in[1] ) );
  BUF_X4 U3254 ( .I(\SB2_2_10/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[146] ) );
  NAND2_X2 U849 ( .A1(\SB1_3_27/i0_0 ), .A2(\SB1_3_27/i3[0] ), .ZN(n4459) );
  CLKBUF_X4 U4451 ( .I(\SB3_31/buf_output[2] ), .Z(\SB4_28/i0_0 ) );
  NAND2_X2 U572 ( .A1(\SB4_31/i0_0 ), .A2(\SB4_31/i3[0] ), .ZN(n2179) );
  BUF_X4 U8945 ( .I(\SB2_3_27/buf_output[3] ), .Z(\RI5[3][39] ) );
  BUF_X4 U2764 ( .I(\MC_ARK_ARC_1_3/buf_output[47] ), .Z(\SB3_24/i0_3 ) );
  NAND3_X2 U4696 ( .A1(\SB1_3_5/i0_4 ), .A2(\SB1_3_5/i0_0 ), .A3(
        \SB1_3_5/i1_5 ), .ZN(n2003) );
  BUF_X4 U8825 ( .I(\SB2_3_15/buf_output[3] ), .Z(n1392) );
  NAND3_X2 U1993 ( .A1(\SB1_1_20/i0[10] ), .A2(\SB1_1_20/i1[9] ), .A3(
        \SB1_1_20/i1_7 ), .ZN(\SB1_1_20/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 \SB2_2_30/Component_Function_2/N1  ( .A1(\SB2_2_30/i1_5 ), .A2(
        \SB2_2_30/i0[10] ), .A3(\SB2_2_30/i1[9] ), .ZN(
        \SB2_2_30/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 U1960 ( .I(\SB1_0_31/buf_output[1] ), .Z(\SB2_0_27/i0[6] ) );
  NAND3_X2 U1350 ( .A1(\SB2_1_28/i0_3 ), .A2(\SB2_1_28/i0_0 ), .A3(
        \SB2_1_28/i0[7] ), .ZN(n1739) );
  BUF_X4 U6496 ( .I(\SB2_1_28/buf_output[1] ), .Z(\RI5[1][43] ) );
  NAND4_X2 U8409 ( .A1(\SB2_1_28/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_1_28/Component_Function_1/NAND4_in[0] ), .A3(n3573), .A4(
        \SB2_1_28/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_1_28/buf_output[1] ) );
  NAND3_X2 U2505 ( .A1(\SB3_5/i0_3 ), .A2(\SB3_5/i1[9] ), .A3(\SB3_5/i0[6] ), 
        .ZN(n2249) );
  NAND3_X2 U686 ( .A1(\SB2_3_6/i0_0 ), .A2(\SB2_3_6/i1_5 ), .A3(\SB2_3_6/i0_4 ), .ZN(n2004) );
  NAND3_X2 U5273 ( .A1(\SB2_1_9/i0[10] ), .A2(\SB2_1_9/i0_0 ), .A3(
        \SB2_1_9/i0[6] ), .ZN(\SB2_1_9/Component_Function_5/NAND4_in[1] ) );
  INV_X2 U3027 ( .I(\SB1_1_5/buf_output[5] ), .ZN(\SB2_1_5/i1_5 ) );
  BUF_X4 U3026 ( .I(\SB1_1_5/buf_output[5] ), .Z(\SB2_1_5/i0_3 ) );
  NAND3_X2 U8979 ( .A1(\SB2_1_20/i1[9] ), .A2(\SB2_1_20/i1_5 ), .A3(
        \SB2_1_20/i0_4 ), .ZN(\SB2_1_20/Component_Function_4/NAND4_in[3] ) );
  NAND3_X2 U4278 ( .A1(\SB1_0_2/i0_4 ), .A2(\SB1_0_2/i1_5 ), .A3(
        \SB1_0_2/i0_0 ), .ZN(n1326) );
  NAND3_X2 U953 ( .A1(\SB2_1_27/i0[10] ), .A2(\SB2_1_27/i1_5 ), .A3(
        \SB2_1_27/i1[9] ), .ZN(\SB2_1_27/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB2_3_13/Component_Function_2/N1  ( .A1(\SB2_3_13/i1_5 ), .A2(
        \SB2_3_13/i0[10] ), .A3(\SB2_3_13/i1[9] ), .ZN(
        \SB2_3_13/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB1_3_15/Component_Function_3/N1  ( .A1(\SB1_3_15/i1[9] ), .A2(
        \SB1_3_15/i0_3 ), .A3(\SB1_3_15/i0[6] ), .ZN(
        \SB1_3_15/Component_Function_3/NAND4_in[0] ) );
  INV_X4 U1384 ( .I(n2535), .ZN(\SB1_1_6/buf_output[4] ) );
  INV_X2 U2614 ( .I(\MC_ARK_ARC_1_3/buf_output[152] ), .ZN(\SB3_6/i1[9] ) );
  NAND3_X2 U1160 ( .A1(\SB1_2_26/i0[10] ), .A2(\SB1_2_26/i0_0 ), .A3(
        \SB1_2_26/i0[6] ), .ZN(\SB1_2_26/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U986 ( .A1(\SB2_2_19/i0_3 ), .A2(\SB2_2_19/i0[10] ), .A3(
        \SB2_2_19/i0[9] ), .ZN(n4169) );
  NAND2_X2 \SB2_1_7/Component_Function_1/N1  ( .A1(\SB2_1_7/i0_3 ), .A2(
        \SB2_1_7/i1[9] ), .ZN(\SB2_1_7/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 \SB1_1_10/Component_Function_2/N4  ( .A1(\SB1_1_10/i1_5 ), .A2(
        \SB1_1_10/i0_0 ), .A3(\SB1_1_10/i0_4 ), .ZN(
        \SB1_1_10/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 U8738 ( .A1(\SB2_3_12/i1_5 ), .A2(\SB2_3_12/i0[10] ), .A3(
        \SB2_3_12/i1[9] ), .ZN(\SB2_3_12/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 U1889 ( .I(\MC_ARK_ARC_1_1/buf_output[182] ), .Z(\SB1_2_1/i0_0 ) );
  CLKBUF_X4 U4894 ( .I(\SB1_3_9/buf_output[2] ), .Z(\SB2_3_6/i0_0 ) );
  BUF_X2 \SB2_0_2/BUF_0  ( .I(\SB1_0_7/buf_output[0] ), .Z(\SB2_0_2/i0[9] ) );
  BUF_X2 U201 ( .I(Key[184]), .Z(n137) );
  NAND3_X2 U867 ( .A1(\SB1_3_27/i0_0 ), .A2(\SB1_3_27/i1_5 ), .A3(
        \SB1_3_27/i0_4 ), .ZN(n1152) );
  NAND2_X2 \SB2_1_9/Component_Function_5/N1  ( .A1(\SB2_1_9/i0_0 ), .A2(
        \SB2_1_9/i3[0] ), .ZN(\SB2_1_9/Component_Function_5/NAND4_in[0] ) );
  CLKBUF_X4 \SB2_3_6/BUF_0  ( .I(\SB1_3_11/buf_output[0] ), .Z(\SB2_3_6/i0[9] ) );
  INV_X2 \SB2_1_9/INV_1  ( .I(\SB1_1_13/buf_output[1] ), .ZN(\SB2_1_9/i1_7 )
         );
  BUF_X4 \SB2_2_16/BUF_1  ( .I(\SB1_2_20/buf_output[1] ), .Z(\SB2_2_16/i0[6] )
         );
  NAND3_X2 \SB1_1_7/Component_Function_2/N1  ( .A1(\SB1_1_7/i1_5 ), .A2(
        \SB1_1_7/i0[10] ), .A3(\SB1_1_7/i1[9] ), .ZN(
        \SB1_1_7/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U701 ( .A1(\SB2_3_2/i0[10] ), .A2(\SB2_3_2/i0_3 ), .A3(
        \SB2_3_2/i0[6] ), .ZN(\SB2_3_2/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 \SB1_3_2/BUF_1  ( .I(\MC_ARK_ARC_1_2/buf_output[175] ), .Z(
        \SB1_3_2/i0[6] ) );
  NAND3_X1 U926 ( .A1(\SB1_2_7/i0[8] ), .A2(\SB1_2_7/i1_5 ), .A3(
        \SB1_2_7/i3[0] ), .ZN(n1819) );
  NAND2_X2 \SB4_2/Component_Function_5/N1  ( .A1(\SB4_2/i0_0 ), .A2(
        \SB4_2/i3[0] ), .ZN(\SB4_2/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U8935 ( .A1(\SB3_5/i0[8] ), .A2(\SB3_5/i0_3 ), .A3(\SB3_5/i0[9] ), 
        .ZN(\SB3_5/Component_Function_2/NAND4_in[2] ) );
  NAND2_X1 U4680 ( .A1(\SB3_5/i0_0 ), .A2(\SB3_5/i3[0] ), .ZN(n2135) );
  NAND3_X2 \SB2_0_4/Component_Function_2/N1  ( .A1(\SB2_0_4/i1_5 ), .A2(
        \SB2_0_4/i0[10] ), .A3(\SB2_0_4/i1[9] ), .ZN(
        \SB2_0_4/Component_Function_2/NAND4_in[0] ) );
  INV_X2 U2698 ( .I(n289), .ZN(\SB1_0_17/i1[9] ) );
  BUF_X2 U53 ( .I(Key[61]), .Z(n90) );
  NAND3_X2 U11025 ( .A1(\SB2_0_10/i0_4 ), .A2(n571), .A3(\SB2_0_10/i0[6] ), 
        .ZN(\SB2_0_10/Component_Function_5/NAND4_in[3] ) );
  NAND2_X2 \SB1_2_12/Component_Function_5/N1  ( .A1(\SB1_2_12/i0_0 ), .A2(
        \SB1_2_12/i3[0] ), .ZN(\SB1_2_12/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB2_0_29/Component_Function_0/N2  ( .A1(\SB2_0_29/i0[8] ), .A2(
        \SB2_0_29/i0[7] ), .A3(\SB2_0_29/i0[6] ), .ZN(
        \SB2_0_29/Component_Function_0/NAND4_in[1] ) );
  NAND3_X2 \SB2_3_27/Component_Function_2/N1  ( .A1(\SB2_3_27/i1_5 ), .A2(
        \SB2_3_27/i0[10] ), .A3(\SB2_3_27/i1[9] ), .ZN(
        \SB2_3_27/Component_Function_2/NAND4_in[0] ) );
  INV_X2 U1981 ( .I(\SB3_7/buf_output[3] ), .ZN(\SB4_5/i0[8] ) );
  BUF_X2 U147 ( .I(Key[59]), .Z(n200) );
  NAND3_X2 \SB1_3_0/Component_Function_2/N2  ( .A1(\SB1_3_0/i0_3 ), .A2(
        \SB1_3_0/i0[10] ), .A3(\SB1_3_0/i0[6] ), .ZN(
        \SB1_3_0/Component_Function_2/NAND4_in[1] ) );
  NAND2_X2 \SB1_3_13/Component_Function_5/N1  ( .A1(\SB1_3_13/i0_0 ), .A2(
        \SB1_3_13/i3[0] ), .ZN(\SB1_3_13/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 \SB2_3_8/BUF_2  ( .I(\SB1_3_11/buf_output[2] ), .Z(\SB2_3_8/i0_0 ) );
  NAND3_X2 U10824 ( .A1(\RI3[0][166] ), .A2(\SB2_0_4/i1_5 ), .A3(
        \SB2_0_4/i1[9] ), .ZN(\SB2_0_4/Component_Function_4/NAND4_in[3] ) );
  NAND2_X2 \SB4_5/Component_Function_5/N1  ( .A1(\SB4_5/i0_0 ), .A2(
        \SB4_5/i3[0] ), .ZN(\SB4_5/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 U3017 ( .I(\SB1_0_11/buf_output[5] ), .Z(\SB2_0_11/i0_3 ) );
  NAND4_X2 U5030 ( .A1(\SB2_0_2/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_0_2/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_0_2/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_0_2/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_0_2/buf_output[1] ) );
  BUF_X4 \SB2_0_2/BUF_5  ( .I(\RI3[0][179] ), .Z(\SB2_0_2/i0_3 ) );
  NAND3_X2 \SB1_2_3/Component_Function_3/N3  ( .A1(\SB1_2_3/i1[9] ), .A2(
        \SB1_2_3/i1_7 ), .A3(\SB1_2_3/i0[10] ), .ZN(
        \SB1_2_3/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U2132 ( .A1(\SB2_2_23/i0_3 ), .A2(\SB2_2_23/i0[6] ), .A3(
        \SB2_2_23/i1[9] ), .ZN(\SB2_2_23/Component_Function_3/NAND4_in[0] ) );
  NAND2_X2 U2184 ( .A1(\SB1_3_8/i0_0 ), .A2(\SB1_3_8/i3[0] ), .ZN(
        \SB1_3_8/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U4194 ( .A1(\SB2_0_20/i0[10] ), .A2(\SB2_0_20/i1_5 ), .A3(
        \SB2_0_20/i1[9] ), .ZN(\SB2_0_20/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U3468 ( .A1(\SB1_1_2/i1[9] ), .A2(\SB1_1_2/i1_5 ), .A3(
        \SB1_1_2/i0_4 ), .ZN(\SB1_1_2/Component_Function_4/NAND4_in[3] ) );
  NAND3_X2 \SB1_0_22/Component_Function_3/N2  ( .A1(\SB1_0_22/i0_0 ), .A2(
        \SB1_0_22/i0_3 ), .A3(\SB1_0_22/i0_4 ), .ZN(
        \SB1_0_22/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U10268 ( .A1(\SB2_0_2/i1[9] ), .A2(\SB2_0_2/i0[10] ), .A3(
        \SB2_0_2/i1_5 ), .ZN(\SB2_0_2/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U5196 ( .A1(\SB2_1_8/i0[10] ), .A2(\SB2_1_8/i0[6] ), .A3(
        \SB2_1_8/i0_3 ), .ZN(n3091) );
  BUF_X2 \MC_ARK_ARC_1_0/BUF_46  ( .I(\SB2_0_25/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[46] ) );
  BUF_X4 U8855 ( .I(\MC_ARK_ARC_1_3/buf_output[35] ), .Z(\SB3_26/i0_3 ) );
  NAND3_X2 \SB2_2_5/Component_Function_4/N4  ( .A1(\SB2_2_5/i1[9] ), .A2(
        \SB2_2_5/i1_5 ), .A3(\SB2_2_5/i0_4 ), .ZN(
        \SB2_2_5/Component_Function_4/NAND4_in[3] ) );
  INV_X2 U8993 ( .I(n274), .ZN(\SB1_0_22/i1[9] ) );
  NAND3_X2 U3398 ( .A1(\SB2_0_19/i1_5 ), .A2(n2774), .A3(\SB2_0_19/i1[9] ), 
        .ZN(\SB2_0_19/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U1256 ( .A1(\SB2_1_4/i0_3 ), .A2(\SB1_1_5/buf_output[4] ), .A3(
        \SB2_1_4/i0[10] ), .ZN(n845) );
  NAND2_X2 \SB1_0_22/Component_Function_5/N1  ( .A1(\SB1_0_22/i0_0 ), .A2(
        \SB1_0_22/i3[0] ), .ZN(\SB1_0_22/Component_Function_5/NAND4_in[0] ) );
  BUF_X4 \SB1_0_22/BUF_5  ( .I(n414), .Z(\SB1_0_22/i0_3 ) );
  NAND3_X2 U5822 ( .A1(\SB2_3_2/i0_0 ), .A2(\SB2_3_2/i0_4 ), .A3(
        \SB2_3_2/i1_5 ), .ZN(\SB2_3_2/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 \SB2_0_19/Component_Function_3/N3  ( .A1(\SB2_0_19/i1[9] ), .A2(
        \SB2_0_19/i1_7 ), .A3(n2774), .ZN(
        \SB2_0_19/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U8655 ( .A1(\SB2_3_23/i1_5 ), .A2(\SB2_3_23/i0[10] ), .A3(
        \SB2_3_23/i1[9] ), .ZN(\SB2_3_23/Component_Function_2/NAND4_in[0] ) );
  BUF_X2 U183 ( .I(Key[45]), .Z(n153) );
  NAND3_X2 \SB2_0_28/Component_Function_2/N3  ( .A1(\SB2_0_28/i0_3 ), .A2(
        \SB2_0_28/i0[8] ), .A3(\RI3[0][18] ), .ZN(
        \SB2_0_28/Component_Function_2/NAND4_in[2] ) );
  NAND2_X2 U4697 ( .A1(\SB1_3_5/i0_0 ), .A2(\SB1_3_5/i3[0] ), .ZN(
        \SB1_3_5/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U9219 ( .A1(n2687), .A2(\SB2_1_0/i0[9] ), .A3(\SB2_1_0/i0[6] ), 
        .ZN(n3756) );
  NAND3_X2 U2927 ( .A1(\SB3_30/i1_5 ), .A2(\SB3_30/i0[8] ), .A3(\SB3_30/i3[0] ), .ZN(n807) );
  INV_X2 U2115 ( .I(\MC_ARK_ARC_1_1/buf_output[51] ), .ZN(\SB1_2_23/i0[8] ) );
  NAND3_X2 \SB2_1_26/Component_Function_3/N4  ( .A1(\SB2_1_26/i1_5 ), .A2(
        \SB2_1_26/i0[8] ), .A3(\SB2_1_26/i3[0] ), .ZN(
        \SB2_1_26/Component_Function_3/NAND4_in[3] ) );
  BUF_X2 U141 ( .I(Key[71]), .Z(n240) );
  NAND3_X2 U1562 ( .A1(\SB2_0_7/i0_0 ), .A2(\SB2_0_7/i1_5 ), .A3(
        \SB1_0_8/buf_output[4] ), .ZN(n4292) );
  NAND3_X2 U2590 ( .A1(\RI3[0][155] ), .A2(n2765), .A3(\SB2_0_6/i0[6] ), .ZN(
        \SB2_0_6/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U2398 ( .A1(\SB2_0_17/i0_3 ), .A2(\SB2_0_17/i0[6] ), .A3(
        \SB2_0_17/i1[9] ), .ZN(n705) );
  NAND3_X2 U2122 ( .A1(\SB1_3_1/i0_0 ), .A2(\SB1_3_1/i0_3 ), .A3(
        \SB1_3_1/i0_4 ), .ZN(\SB1_3_1/Component_Function_3/NAND4_in[1] ) );
  NAND2_X2 \SB1_0_17/Component_Function_5/N1  ( .A1(\SB1_0_17/i0_0 ), .A2(
        \SB1_0_17/i3[0] ), .ZN(\SB1_0_17/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB2_2_5/Component_Function_0/N4  ( .A1(\SB2_2_5/i0[7] ), .A2(
        \SB2_2_5/i0_3 ), .A3(\SB2_2_5/i0_0 ), .ZN(
        \SB2_2_5/Component_Function_0/NAND4_in[3] ) );
  NAND2_X2 U10231 ( .A1(\SB1_1_11/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_1_11/Component_Function_4/NAND4_in[0] ), .ZN(n1464) );
  NAND3_X2 U1016 ( .A1(\SB2_2_19/i0_0 ), .A2(\SB2_2_19/i0_3 ), .A3(
        \SB2_2_19/i0[7] ), .ZN(\SB2_2_19/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U4533 ( .A1(\SB2_2_30/i0[9] ), .A2(\SB2_2_30/i0[6] ), .A3(
        \SB2_2_30/i0_4 ), .ZN(\SB2_2_30/Component_Function_5/NAND4_in[3] ) );
  CLKBUF_X2 U188 ( .I(Key[168]), .Z(n159) );
  NAND2_X2 U695 ( .A1(\SB2_3_25/i0_0 ), .A2(\SB2_3_25/i3[0] ), .ZN(
        \SB2_3_25/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U6965 ( .A1(\SB1_3_22/i0[8] ), .A2(\SB1_3_22/i3[0] ), .A3(
        \SB1_3_22/i1_5 ), .ZN(n3364) );
  NAND3_X2 U3894 ( .A1(\SB2_3_8/i0[9] ), .A2(\SB1_3_9/buf_output[4] ), .A3(
        \SB2_3_8/i0[6] ), .ZN(\SB2_3_8/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 U1423 ( .A1(\SB1_1_30/i0[8] ), .A2(\SB1_1_30/i1_5 ), .A3(
        \SB1_1_30/i3[0] ), .ZN(n4430) );
  BUF_X2 U2 ( .I(Key[3]), .Z(n219) );
  NAND3_X1 U2821 ( .A1(\SB3_18/i0_3 ), .A2(\SB3_18/i0[6] ), .A3(\SB3_18/i1[9] ), .ZN(\SB3_18/Component_Function_3/NAND4_in[0] ) );
  CLKBUF_X4 U8669 ( .I(\SB2_3_14/buf_output[5] ), .Z(\RI5[3][107] ) );
  INV_X2 \SB2_3_25/INV_0  ( .I(\SB1_3_30/buf_output[0] ), .ZN(\SB2_3_25/i3[0] ) );
  NAND3_X2 \SB1_3_30/Component_Function_3/N2  ( .A1(\SB1_3_30/i0_0 ), .A2(
        \SB1_3_30/i0_3 ), .A3(\SB1_3_30/i0_4 ), .ZN(
        \SB1_3_30/Component_Function_3/NAND4_in[1] ) );
  BUF_X4 U4843 ( .I(\MC_ARK_ARC_1_0/buf_output[145] ), .Z(\SB1_1_7/i0[6] ) );
  NAND3_X2 U1079 ( .A1(n571), .A2(\SB2_0_10/i1_5 ), .A3(\SB2_0_10/i0[6] ), 
        .ZN(\SB2_0_10/Component_Function_1/NAND4_in[2] ) );
  NAND2_X2 U761 ( .A1(\SB1_3_10/i3[0] ), .A2(\SB1_3_10/i0_0 ), .ZN(n1329) );
  BUF_X4 U8966 ( .I(\MC_ARK_ARC_1_2/buf_output[128] ), .Z(\SB1_3_10/i0_0 ) );
  NAND3_X2 \SB2_2_28/Component_Function_2/N4  ( .A1(\SB2_2_28/i1_5 ), .A2(
        \SB2_2_28/i0_0 ), .A3(\SB2_2_28/i0_4 ), .ZN(
        \SB2_2_28/Component_Function_2/NAND4_in[3] ) );
  NAND2_X2 U10293 ( .A1(\SB2_2_19/i0_0 ), .A2(\SB2_2_19/i3[0] ), .ZN(n4250) );
  NAND3_X2 U596 ( .A1(\SB3_7/i0_4 ), .A2(\SB3_7/i0[10] ), .A3(\SB3_7/i0_3 ), 
        .ZN(n4289) );
  BUF_X2 \SB4_19/BUF_1  ( .I(\SB3_23/buf_output[1] ), .Z(\SB4_19/i0[6] ) );
  NAND3_X2 U1084 ( .A1(\SB2_0_19/i0[8] ), .A2(\SB2_0_19/i3[0] ), .A3(
        \SB2_0_19/i1_5 ), .ZN(n1239) );
  INV_X2 U1746 ( .I(\SB1_1_9/buf_output[5] ), .ZN(\SB2_1_9/i1_5 ) );
  NAND3_X2 U2556 ( .A1(\SB2_0_6/i1_5 ), .A2(n2765), .A3(\SB2_0_6/i1[9] ), .ZN(
        \SB2_0_6/Component_Function_2/NAND4_in[0] ) );
  NAND2_X2 \SB1_0_18/Component_Function_5/N1  ( .A1(\SB1_0_18/i0_0 ), .A2(
        \SB1_0_18/i3[0] ), .ZN(\SB1_0_18/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U7696 ( .A1(\SB2_1_25/i0[7] ), .A2(\SB2_1_25/i0_0 ), .A3(
        \SB2_1_25/i0_3 ), .ZN(n2744) );
  NAND2_X2 \SB3_31/Component_Function_5/N1  ( .A1(\SB3_31/i0_0 ), .A2(
        \SB3_31/i3[0] ), .ZN(\SB3_31/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U3951 ( .A1(\SB2_0_27/i0_3 ), .A2(\SB2_0_27/i1[9] ), .A3(
        \SB2_0_27/i0_4 ), .ZN(\SB2_0_27/Component_Function_5/NAND4_in[2] ) );
  BUF_X4 U3644 ( .I(\MC_ARK_ARC_1_2/buf_output[184] ), .Z(\SB1_3_1/i0_4 ) );
  NAND3_X2 \SB1_2_31/Component_Function_2/N1  ( .A1(\SB1_2_31/i1_5 ), .A2(
        \SB1_2_31/i0[10] ), .A3(\SB1_2_31/i1[9] ), .ZN(
        \SB1_2_31/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 \SB2_3_9/Component_Function_1/N5  ( .A1(
        \SB2_3_9/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_3_9/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_3_9/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_3_9/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_3_9/buf_output[1] ) );
  NAND3_X2 U2317 ( .A1(\SB3_7/i0[10] ), .A2(\SB3_7/i1[9] ), .A3(\SB3_7/i1_7 ), 
        .ZN(n4660) );
  NAND3_X2 \SB2_2_28/Component_Function_2/N1  ( .A1(\SB2_2_28/i1_5 ), .A2(
        \SB2_2_28/i0[10] ), .A3(\SB2_2_28/i1[9] ), .ZN(
        \SB2_2_28/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 U4892 ( .I(\SB2_0_2/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[7] ) );
  NAND3_X2 U3471 ( .A1(\SB1_3_19/i0[10] ), .A2(\SB1_3_19/i1[9] ), .A3(
        \SB1_3_19/i1_5 ), .ZN(\SB1_3_19/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB2_3_22/Component_Function_3/N2  ( .A1(\SB2_3_22/i0_0 ), .A2(
        \SB2_3_22/i0_3 ), .A3(\SB2_3_22/i0_4 ), .ZN(
        \SB2_3_22/Component_Function_3/NAND4_in[1] ) );
  INV_X2 U2297 ( .I(\SB1_3_8/buf_output[0] ), .ZN(\SB2_3_3/i3[0] ) );
  NAND3_X1 U1597 ( .A1(n2765), .A2(\SB2_0_6/i1_7 ), .A3(\SB2_0_6/i1[9] ), .ZN(
        \SB2_0_6/Component_Function_3/NAND4_in[2] ) );
  BUF_X4 U8663 ( .I(\SB1_2_14/buf_output[2] ), .Z(\SB2_2_11/i0_0 ) );
  NAND2_X2 \SB1_1_26/Component_Function_5/N1  ( .A1(\SB1_1_26/i0_0 ), .A2(
        \SB1_1_26/i3[0] ), .ZN(\SB1_1_26/Component_Function_5/NAND4_in[0] ) );
  NAND2_X2 \SB2_3_2/Component_Function_5/N1  ( .A1(\SB2_3_2/i0_0 ), .A2(
        \SB2_3_2/i3[0] ), .ZN(\SB2_3_2/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U7075 ( .A1(\SB1_3_19/i0[10] ), .A2(\SB1_3_19/i1[9] ), .A3(
        \SB1_3_19/i1_7 ), .ZN(n2373) );
  NAND3_X2 \SB1_2_18/Component_Function_0/N3  ( .A1(\SB1_2_18/i0[10] ), .A2(
        \SB1_2_18/i0_4 ), .A3(\SB1_2_18/i0_3 ), .ZN(
        \SB1_2_18/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 U5376 ( .A1(\SB2_3_23/i0[8] ), .A2(\SB2_3_23/i1_7 ), .A3(
        \SB2_3_23/i0_4 ), .ZN(\SB2_3_23/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 U5892 ( .A1(\SB1_3_24/i0[10] ), .A2(\SB1_3_24/i0[9] ), .A3(
        \SB1_3_24/i0_3 ), .ZN(\SB1_3_24/Component_Function_4/NAND4_in[2] ) );
  NAND3_X2 U2197 ( .A1(\SB1_3_8/i1_5 ), .A2(\SB1_3_8/i0[8] ), .A3(
        \SB1_3_8/i3[0] ), .ZN(n4296) );
  NAND3_X2 U3655 ( .A1(\SB1_3_3/i0[8] ), .A2(\SB1_3_3/i0_4 ), .A3(
        \SB1_3_3/i1_7 ), .ZN(n1684) );
  INV_X4 U6337 ( .I(n3270), .ZN(\RI1[1][143] ) );
  NAND3_X2 \SB2_2_2/Component_Function_0/N3  ( .A1(\SB2_2_2/i0[10] ), .A2(
        \SB2_2_2/i0_4 ), .A3(\SB2_2_2/i0_3 ), .ZN(
        \SB2_2_2/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 \SB2_1_17/Component_Function_1/N2  ( .A1(\SB2_1_17/i0_3 ), .A2(
        \SB2_1_17/i1_7 ), .A3(\SB2_1_17/i0[8] ), .ZN(
        \SB2_1_17/Component_Function_1/NAND4_in[1] ) );
  NAND3_X2 U2834 ( .A1(\SB2_3_4/i0[10] ), .A2(\SB2_3_4/i1[9] ), .A3(
        \SB2_3_4/i1_7 ), .ZN(\SB2_3_4/Component_Function_3/NAND4_in[2] ) );
  CLKBUF_X4 \SB3_3/BUF_0  ( .I(\MC_ARK_ARC_1_3/buf_output[168] ), .Z(
        \SB3_3/i0[9] ) );
  INV_X1 U283 ( .I(n30), .ZN(n506) );
  CLKBUF_X4 U1580 ( .I(\SB3_4/buf_output[0] ), .Z(\SB4_31/i0[9] ) );
  BUF_X2 U70 ( .I(Key[1]), .Z(n39) );
  BUF_X4 \SB2_2_24/BUF_1  ( .I(\SB1_2_28/buf_output[1] ), .Z(\SB2_2_24/i0[6] )
         );
  CLKBUF_X2 U78 ( .I(Key[179]), .Z(n238) );
  INV_X2 U2907 ( .I(\MC_ARK_ARC_1_2/buf_output[189] ), .ZN(\SB1_3_0/i0[8] ) );
  INV_X2 U2302 ( .I(\MC_ARK_ARC_1_3/buf_output[45] ), .ZN(\SB3_24/i0[8] ) );
  NAND3_X2 U2916 ( .A1(\SB1_3_26/i0[8] ), .A2(\SB1_3_26/i1_5 ), .A3(
        \SB1_3_26/i3[0] ), .ZN(n1760) );
  BUF_X4 \SB2_3_3/BUF_3  ( .I(\SB1_3_5/buf_output[3] ), .Z(\SB2_3_3/i0[10] )
         );
  NAND3_X2 U9965 ( .A1(\SB2_0_6/i0_0 ), .A2(\SB2_0_6/i1_5 ), .A3(\RI3[0][154] ), .ZN(n4079) );
  NAND3_X2 U798 ( .A1(\SB1_3_31/i0[6] ), .A2(\SB1_3_31/i0_4 ), .A3(
        \SB1_3_31/i0[9] ), .ZN(n1251) );
  CLKBUF_X2 U137 ( .I(Key[106]), .Z(n188) );
  BUF_X4 U3442 ( .I(\MC_ARK_ARC_1_0/buf_output[21] ), .Z(\SB1_1_28/i0[10] ) );
  BUF_X4 U9052 ( .I(\MC_ARK_ARC_1_1/buf_output[16] ), .Z(\SB1_2_29/i0_4 ) );
  NAND3_X2 U7002 ( .A1(\SB3_5/i0_3 ), .A2(\SB3_5/i0_0 ), .A3(\SB3_5/i0_4 ), 
        .ZN(\SB3_5/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 \SB1_3_18/Component_Function_2/N1  ( .A1(\SB1_3_18/i1_5 ), .A2(
        \SB1_3_18/i0[10] ), .A3(\SB1_3_18/i1[9] ), .ZN(
        \SB1_3_18/Component_Function_2/NAND4_in[0] ) );
  NAND2_X2 \SB2_0_4/Component_Function_0/N1  ( .A1(\SB2_0_4/i0[10] ), .A2(
        \SB2_0_4/i0[9] ), .ZN(\SB2_0_4/Component_Function_0/NAND4_in[0] ) );
  INV_X2 U2492 ( .I(\MC_ARK_ARC_1_3/buf_output[116] ), .ZN(\SB3_12/i1[9] ) );
  NAND3_X2 \SB2_2_31/Component_Function_2/N2  ( .A1(\SB2_2_31/i0_3 ), .A2(
        \SB2_2_31/i0[10] ), .A3(\SB2_2_31/i0[6] ), .ZN(
        \SB2_2_31/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 U8826 ( .I(\MC_ARK_ARC_1_2/buf_output[83] ), .Z(\SB1_3_18/i0_3 ) );
  NAND3_X2 \SB1_0_12/Component_Function_2/N3  ( .A1(\SB1_0_12/i0_3 ), .A2(
        \SB1_0_12/i0[8] ), .A3(\SB1_0_12/i0[9] ), .ZN(
        \SB1_0_12/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U2174 ( .A1(\SB3_5/i0_3 ), .A2(\SB3_5/i1[9] ), .A3(\SB3_5/i0_4 ), 
        .ZN(n2158) );
  NAND3_X2 \SB2_0_30/Component_Function_5/N3  ( .A1(\SB2_0_30/i1[9] ), .A2(
        \RI3[0][10] ), .A3(\SB2_0_30/i0_3 ), .ZN(
        \SB2_0_30/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U1315 ( .A1(\SB2_1_6/i0_3 ), .A2(\SB2_1_6/i0[10] ), .A3(
        \SB2_1_6/i0_4 ), .ZN(n4441) );
  INV_X2 \SB1_0_14/INV_0  ( .I(n296), .ZN(\SB1_0_14/i3[0] ) );
  NAND3_X2 U8641 ( .A1(\SB1_3_19/i0[10] ), .A2(\SB1_3_19/i0[9] ), .A3(
        \SB1_3_19/i0_3 ), .ZN(\SB1_3_19/Component_Function_4/NAND4_in[2] ) );
  NAND3_X2 U1559 ( .A1(\SB3_31/i0_0 ), .A2(\SB3_31/i0[6] ), .A3(
        \SB3_31/i0[10] ), .ZN(\SB3_31/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 \SB1_0_18/Component_Function_5/N2  ( .A1(\SB1_0_18/i0_0 ), .A2(
        \SB1_0_18/i0[6] ), .A3(n367), .ZN(
        \SB1_0_18/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 \SB2_2_31/Component_Function_3/N1  ( .A1(\SB2_2_31/i1[9] ), .A2(
        \SB2_2_31/i0_3 ), .A3(\SB2_2_31/i0[6] ), .ZN(
        \SB2_2_31/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 \SB2_2_31/Component_Function_1/N3  ( .A1(\SB2_2_31/i1_5 ), .A2(
        \SB2_2_31/i0[6] ), .A3(\SB2_2_31/i0[9] ), .ZN(
        \SB2_2_31/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 U5754 ( .A1(\SB1_2_11/i0[6] ), .A2(\SB1_2_11/i0[9] ), .A3(
        \SB1_2_11/i0_4 ), .ZN(\SB1_2_11/Component_Function_5/NAND4_in[3] ) );
  BUF_X2 U81 ( .I(Key[111]), .Z(n204) );
  BUF_X4 U3547 ( .I(\MC_ARK_ARC_1_1/buf_output[3] ), .Z(\SB1_2_31/i0[10] ) );
  BUF_X4 \SB4_18/BUF_0  ( .I(\SB3_23/buf_output[0] ), .Z(\SB4_18/i0[9] ) );
  BUF_X2 U107 ( .I(Key[181]), .Z(n60) );
  BUF_X4 \SB2_2_31/BUF_3  ( .I(\SB1_2_1/buf_output[3] ), .Z(\SB2_2_31/i0[10] )
         );
  NAND4_X2 U4888 ( .A1(\SB2_3_20/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_3_20/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_3_20/Component_Function_1/NAND4_in[0] ), .A4(n3054), .ZN(
        \SB2_3_20/buf_output[1] ) );
  INV_X2 U6608 ( .I(\SB2_0_11/i0_4 ), .ZN(\SB2_0_11/i0[7] ) );
  NAND2_X2 \SB2_2_17/Component_Function_5/N1  ( .A1(\SB2_2_17/i0_0 ), .A2(
        \SB2_2_17/i3[0] ), .ZN(\SB2_2_17/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB1_0_2/Component_Function_0/N3  ( .A1(\SB1_0_2/i0[10] ), .A2(
        \SB1_0_2/i0_4 ), .A3(\SB1_0_2/i0_3 ), .ZN(
        \SB1_0_2/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 \SB3_5/Component_Function_5/N4  ( .A1(\SB3_5/i0[9] ), .A2(
        \SB3_5/i0[6] ), .A3(\SB3_5/i0_4 ), .ZN(
        \SB3_5/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 U8711 ( .A1(\SB1_1_13/i0[8] ), .A2(\SB1_1_13/i1_5 ), .A3(
        \SB1_1_13/i3[0] ), .ZN(n2678) );
  NAND2_X2 \SB2_2_5/Component_Function_1/N1  ( .A1(\SB2_2_5/i0_3 ), .A2(
        \SB2_2_5/i1[9] ), .ZN(\SB2_2_5/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 \SB1_2_21/Component_Function_2/N3  ( .A1(\SB1_2_21/i0_3 ), .A2(
        \SB1_2_21/i0[8] ), .A3(\SB1_2_21/i0[9] ), .ZN(
        \SB1_2_21/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U2786 ( .A1(\SB2_2_29/i0_3 ), .A2(\SB2_2_29/i1[9] ), .A3(
        \SB2_2_29/i0[6] ), .ZN(\SB2_2_29/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 \SB1_0_18/Component_Function_3/N2  ( .A1(\SB1_0_18/i0_0 ), .A2(
        \SB1_0_18/i0_3 ), .A3(n4753), .ZN(
        \SB1_0_18/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_29/Component_Function_1/N4  ( .A1(\SB1_1_29/i1_7 ), .A2(
        \SB1_1_29/i0[8] ), .A3(\SB1_1_29/i0_4 ), .ZN(
        \SB1_1_29/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 U5500 ( .A1(\SB2_3_23/i0_4 ), .A2(\SB2_3_23/i1[9] ), .A3(
        \SB2_3_23/i1_5 ), .ZN(n1652) );
  BUF_X2 U133 ( .I(Key[7]), .Z(n201) );
  BUF_X4 \SB4_2/BUF_4  ( .I(\SB3_3/buf_output[4] ), .Z(\SB4_2/i0_4 ) );
  NAND3_X2 \SB2_0_0/Component_Function_2/N2  ( .A1(\RI3[0][191] ), .A2(
        \SB2_0_0/i0[10] ), .A3(\SB2_0_0/i0[6] ), .ZN(
        \SB2_0_0/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 \SB3_27/Component_Function_4/N3  ( .A1(\SB3_27/i0[9] ), .A2(
        \SB3_27/i0[10] ), .A3(\SB3_27/i0_3 ), .ZN(
        \SB3_27/Component_Function_4/NAND4_in[2] ) );
  NAND3_X2 \SB2_2_0/Component_Function_1/N4  ( .A1(\SB2_2_0/i1_7 ), .A2(
        \SB2_2_0/i0[8] ), .A3(\SB2_2_0/i0_4 ), .ZN(
        \SB2_2_0/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 \SB1_0_2/Component_Function_2/N1  ( .A1(\SB1_0_2/i1_5 ), .A2(
        \SB1_0_2/i0[10] ), .A3(\SB1_0_2/i1[9] ), .ZN(
        \SB1_0_2/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U692 ( .A1(\SB1_3_14/buf_output[4] ), .A2(\SB2_3_13/i1[9] ), .A3(
        \SB2_3_13/i1_5 ), .ZN(n3320) );
  BUF_X4 U1496 ( .I(\MC_ARK_ARC_1_1/buf_output[106] ), .Z(\SB1_2_14/i0_4 ) );
  NAND3_X2 \SB2_3_13/Component_Function_2/N3  ( .A1(\SB2_3_13/i0_3 ), .A2(
        \SB2_3_13/i0[8] ), .A3(\SB2_3_13/i0[9] ), .ZN(
        \SB2_3_13/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 U1077 ( .I(\SB1_2_11/buf_output[1] ), .Z(\SB2_2_7/i0[6] ) );
  NAND2_X1 U1318 ( .A1(\SB3_14/i0_0 ), .A2(\SB3_14/i3[0] ), .ZN(
        \SB3_14/Component_Function_5/NAND4_in[0] ) );
  NAND2_X2 \SB2_1_10/Component_Function_1/N1  ( .A1(\SB2_1_10/i0_3 ), .A2(
        \SB2_1_10/i1[9] ), .ZN(\SB2_1_10/Component_Function_1/NAND4_in[0] ) );
  BUF_X4 U4845 ( .I(\MC_ARK_ARC_1_0/buf_output[135] ), .Z(\SB1_1_9/i0[10] ) );
  CLKBUF_X4 U8117 ( .I(\SB2_1_26/buf_output[2] ), .Z(\RI5[1][50] ) );
  NAND2_X2 \SB2_2_28/Component_Function_0/N1  ( .A1(\SB2_2_28/i0[10] ), .A2(
        \SB2_2_28/i0[9] ), .ZN(\SB2_2_28/Component_Function_0/NAND4_in[0] ) );
  NAND3_X2 \SB2_0_7/Component_Function_2/N1  ( .A1(\SB2_0_7/i1_5 ), .A2(
        \RI3[0][147] ), .A3(\SB2_0_7/i1[9] ), .ZN(
        \SB2_0_7/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 U1598 ( .I(\MC_ARK_ARC_1_1/buf_output[52] ), .Z(\SB1_2_23/i0_4 ) );
  BUF_X4 U8261 ( .I(\SB2_3_9/buf_output[1] ), .Z(\RI5[3][157] ) );
  NAND2_X2 \SB2_2_2/Component_Function_1/N1  ( .A1(\SB2_2_2/i0_3 ), .A2(
        \SB2_2_2/i1[9] ), .ZN(\SB2_2_2/Component_Function_1/NAND4_in[0] ) );
  NAND4_X2 U2448 ( .A1(\SB2_1_13/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_1_13/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_1_13/Component_Function_1/NAND4_in[2] ), .A4(n654), .ZN(
        \SB2_1_13/buf_output[1] ) );
  NAND3_X2 \SB2_1_13/Component_Function_1/N3  ( .A1(\SB2_1_13/i1_5 ), .A2(
        \SB1_1_17/buf_output[1] ), .A3(\SB1_1_18/buf_output[0] ), .ZN(
        \SB2_1_13/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 \SB2_0_24/Component_Function_2/N4  ( .A1(\SB2_0_24/i1_5 ), .A2(
        \SB2_0_24/i0_0 ), .A3(\RI3[0][46] ), .ZN(
        \SB2_0_24/Component_Function_2/NAND4_in[3] ) );
  NAND2_X2 U1475 ( .A1(\SB1_1_17/i0_3 ), .A2(\SB1_1_17/i1[9] ), .ZN(
        \SB1_1_17/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 U6829 ( .A1(\SB1_0_25/i0[6] ), .A2(\SB1_0_25/i1_5 ), .A3(
        \SB1_0_25/i0[9] ), .ZN(\SB1_0_25/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 U10427 ( .A1(\SB2_3_22/i0[10] ), .A2(\SB2_3_22/i1_5 ), .A3(
        \SB2_3_22/i1[9] ), .ZN(\SB2_3_22/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 \SB1_0_31/Component_Function_2/N3  ( .A1(\SB1_0_31/i0_3 ), .A2(
        \SB1_0_31/i0[8] ), .A3(\SB1_0_31/i0[9] ), .ZN(
        \SB1_0_31/Component_Function_2/NAND4_in[2] ) );
  BUF_X2 U2946 ( .I(\SB1_0_15/buf_output[3] ), .Z(\SB2_0_13/i0[10] ) );
  NAND3_X2 U6412 ( .A1(\SB2_1_7/i0[7] ), .A2(\SB2_1_7/i0[8] ), .A3(n2852), 
        .ZN(\SB2_1_7/Component_Function_0/NAND4_in[1] ) );
  NAND3_X2 U3658 ( .A1(\SB1_3_9/i0[8] ), .A2(\SB1_3_9/i1_7 ), .A3(
        \SB1_3_9/i0_4 ), .ZN(\SB1_3_9/Component_Function_1/NAND4_in[3] ) );
  INV_X4 \SB2_2_14/INV_4  ( .I(n5932), .ZN(\SB2_2_14/i0[7] ) );
  NAND3_X2 \SB1_0_11/Component_Function_1/N4  ( .A1(\SB1_0_11/i1_7 ), .A2(
        \SB1_0_11/i0[8] ), .A3(\SB1_0_11/i0_4 ), .ZN(
        \SB1_0_11/Component_Function_1/NAND4_in[3] ) );
  INV_X2 \SB1_1_14/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[107] ), .ZN(
        \SB1_1_14/i1_5 ) );
  NAND3_X2 \SB1_1_14/Component_Function_5/N3  ( .A1(\SB1_1_14/i1[9] ), .A2(
        \SB1_1_14/i0_4 ), .A3(\SB1_1_14/i0_3 ), .ZN(
        \SB1_1_14/Component_Function_5/NAND4_in[2] ) );
  BUF_X2 U94 ( .I(Key[44]), .Z(n71) );
  BUF_X4 U3688 ( .I(\SB2_1_11/buf_output[3] ), .Z(\RI5[1][135] ) );
  BUF_X2 U2142 ( .I(\SB1_3_7/buf_output[1] ), .Z(\SB2_3_3/i0[6] ) );
  NAND3_X2 U9578 ( .A1(\SB3_1/i0_0 ), .A2(\SB3_1/i0[10] ), .A3(\SB3_1/i0[6] ), 
        .ZN(\SB3_1/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 \SB2_0_7/Component_Function_1/N3  ( .A1(\SB2_0_7/i1_5 ), .A2(n2593), 
        .A3(\SB2_0_7/i0[9] ), .ZN(\SB2_0_7/Component_Function_1/NAND4_in[2] )
         );
  NAND3_X2 U1587 ( .A1(\SB2_0_21/i0_3 ), .A2(\SB2_0_21/i0[9] ), .A3(
        \SB2_0_21/i0[10] ), .ZN(\SB2_0_21/Component_Function_4/NAND4_in[2] )
         );
  INV_X2 U8970 ( .I(\MC_ARK_ARC_1_1/buf_output[125] ), .ZN(\SB1_2_11/i1_5 ) );
  NAND3_X2 U1292 ( .A1(\SB2_1_11/i0[6] ), .A2(\SB1_1_16/buf_output[0] ), .A3(
        \SB1_1_12/buf_output[4] ), .ZN(n3987) );
  NAND2_X2 \SB2_1_20/Component_Function_1/N1  ( .A1(\SB2_1_20/i0_3 ), .A2(
        \SB2_1_20/i1[9] ), .ZN(\SB2_1_20/Component_Function_1/NAND4_in[0] ) );
  INV_X2 \SB1_1_27/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[29] ), .ZN(
        \SB1_1_27/i1_5 ) );
  NAND3_X2 \SB1_1_2/Component_Function_4/N1  ( .A1(\SB1_1_2/i0[9] ), .A2(
        \SB1_1_2/i0_0 ), .A3(\SB1_1_2/i0[8] ), .ZN(
        \SB1_1_2/Component_Function_4/NAND4_in[0] ) );
  NAND3_X2 \SB1_2_5/Component_Function_2/N2  ( .A1(\SB1_2_5/i0_3 ), .A2(
        \SB1_2_5/i0[10] ), .A3(\SB1_2_5/i0[6] ), .ZN(
        \SB1_2_5/Component_Function_2/NAND4_in[1] ) );
  INV_X4 U3895 ( .I(n5790), .ZN(\SB2_1_7/i0[7] ) );
  BUF_X4 \SB2_2_2/BUF_2  ( .I(\SB1_2_5/buf_output[2] ), .Z(\SB2_2_2/i0_0 ) );
  NAND3_X1 U6471 ( .A1(\SB1_2_13/i0[6] ), .A2(\SB1_2_13/i0[8] ), .A3(
        \SB1_2_13/i0[7] ), .ZN(\SB1_2_13/Component_Function_0/NAND4_in[1] ) );
  CLKBUF_X2 U164 ( .I(Key[135]), .Z(n197) );
  NAND2_X2 U1540 ( .A1(\SB2_0_10/i0_0 ), .A2(\SB2_0_10/i3[0] ), .ZN(n4258) );
  NAND3_X2 U8951 ( .A1(\SB1_0_13/i0[6] ), .A2(\SB1_0_13/i0_4 ), .A3(
        \SB1_0_13/i0[9] ), .ZN(n4259) );
  NAND3_X2 U8668 ( .A1(\SB3_12/i1[9] ), .A2(\SB3_12/i1_7 ), .A3(
        \SB3_12/i0[10] ), .ZN(\SB3_12/Component_Function_3/NAND4_in[2] ) );
  OAI21_X2 U3380 ( .A1(n2903), .A2(n971), .B(\SB2_3_21/i0[7] ), .ZN(n970) );
  BUF_X4 U2724 ( .I(\SB1_2_7/buf_output[3] ), .Z(\SB2_2_5/i0[10] ) );
  NAND2_X2 \SB2_0_24/Component_Function_5/N1  ( .A1(\SB2_0_24/i0_0 ), .A2(
        \SB2_0_24/i3[0] ), .ZN(\SB2_0_24/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 \SB1_2_18/Component_Function_4/N4  ( .A1(\SB1_2_18/i1[9] ), .A2(
        \SB1_2_18/i1_5 ), .A3(\SB1_2_18/i0_4 ), .ZN(
        \SB1_2_18/Component_Function_4/NAND4_in[3] ) );
  NAND3_X2 \SB3_7/Component_Function_3/N1  ( .A1(\SB3_7/i1[9] ), .A2(
        \SB3_7/i0_3 ), .A3(\SB3_7/i0[6] ), .ZN(
        \SB3_7/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U2930 ( .A1(\SB4_24/i0_3 ), .A2(\SB4_24/i0_0 ), .A3(\SB4_24/i0[7] ), 
        .ZN(n4642) );
  BUF_X4 \SB2_0_21/BUF_2  ( .I(\RI3[0][62] ), .Z(\SB2_0_21/i0_0 ) );
  CLKBUF_X2 U202 ( .I(Key[91]), .Z(n181) );
  NAND3_X2 \SB2_3_6/Component_Function_3/N4  ( .A1(\SB2_3_6/i1_5 ), .A2(
        \SB2_3_6/i0[8] ), .A3(\SB2_3_6/i3[0] ), .ZN(
        \SB2_3_6/Component_Function_3/NAND4_in[3] ) );
  BUF_X2 U2465 ( .I(\MC_ARK_ARC_1_2/buf_output[9] ), .Z(\SB1_3_30/i0[10] ) );
  CLKBUF_X4 \SB1_3_24/BUF_0  ( .I(\MC_ARK_ARC_1_2/buf_output[42] ), .Z(
        \SB1_3_24/i0[9] ) );
  NAND2_X1 U3968 ( .A1(\SB1_2_3/i0_0 ), .A2(\SB1_2_3/i3[0] ), .ZN(n2933) );
  BUF_X4 U8988 ( .I(\SB2_0_9/buf_output[3] ), .Z(\RI5[0][147] ) );
  NAND3_X2 U7636 ( .A1(\SB1_1_16/i0[6] ), .A2(\SB1_1_16/i0[9] ), .A3(
        \SB1_1_16/i0_4 ), .ZN(n2713) );
  NAND4_X2 U4641 ( .A1(\SB1_2_14/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_14/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_2_14/Component_Function_2/NAND4_in[2] ), .A4(n1225), .ZN(
        \SB1_2_14/buf_output[2] ) );
  NAND3_X2 \SB2_1_29/Component_Function_3/N1  ( .A1(\SB2_1_29/i1[9] ), .A2(
        \SB2_1_29/i0_3 ), .A3(\SB2_1_29/i0[6] ), .ZN(
        \SB2_1_29/Component_Function_3/NAND4_in[0] ) );
  BUF_X2 U25 ( .I(Key[76]), .Z(n172) );
  BUF_X4 U1892 ( .I(\SB2_1_26/buf_output[3] ), .Z(\RI5[1][45] ) );
  CLKBUF_X4 \MC_ARK_ARC_1_0/BUF_2  ( .I(\SB2_0_2/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[2] ) );
  INV_X2 U4625 ( .I(\MC_ARK_ARC_1_2/buf_output[173] ), .ZN(\SB1_3_3/i1_5 ) );
  BUF_X4 U4624 ( .I(\MC_ARK_ARC_1_2/buf_output[173] ), .Z(\SB1_3_3/i0_3 ) );
  NAND3_X2 \SB2_1_27/Component_Function_4/N1  ( .A1(\SB2_1_27/i0[9] ), .A2(
        \SB2_1_27/i0_0 ), .A3(\SB2_1_27/i0[8] ), .ZN(
        \SB2_1_27/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U2277 ( .A1(\SB4_29/i0_3 ), .A2(\SB4_29/i0[8] ), .A3(\SB4_29/i0[9] ), .ZN(\SB4_29/Component_Function_2/NAND4_in[2] ) );
  CLKBUF_X4 \SB2_2_10/BUF_1  ( .I(\SB1_2_14/buf_output[1] ), .Z(
        \SB2_2_10/i0[6] ) );
  BUF_X4 U8992 ( .I(\SB3_31/buf_output[3] ), .Z(\SB4_29/i0[10] ) );
  CLKBUF_X2 U157 ( .I(Key[147]), .Z(n216) );
  BUF_X4 \SB1_3_9/BUF_1  ( .I(\MC_ARK_ARC_1_2/buf_output[133] ), .Z(
        \SB1_3_9/i0[6] ) );
  NAND3_X2 \SB2_2_30/Component_Function_3/N1  ( .A1(\SB2_2_30/i1[9] ), .A2(
        \SB2_2_30/i0_3 ), .A3(\SB2_2_30/i0[6] ), .ZN(
        \SB2_2_30/Component_Function_3/NAND4_in[0] ) );
  NAND2_X2 \SB1_3_8/Component_Function_1/N1  ( .A1(\SB1_3_8/i0_3 ), .A2(
        \SB1_3_8/i1[9] ), .ZN(\SB1_3_8/Component_Function_1/NAND4_in[0] ) );
  NAND4_X2 U5357 ( .A1(\SB2_0_30/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_0_30/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_0_30/Component_Function_4/NAND4_in[1] ), .A4(
        \SB2_0_30/Component_Function_4/NAND4_in[0] ), .ZN(
        \SB2_0_30/buf_output[4] ) );
  NAND3_X2 U3465 ( .A1(\SB1_1_0/i0[9] ), .A2(\SB1_1_0/i0_3 ), .A3(
        \SB1_1_0/i0[8] ), .ZN(n1577) );
  NAND3_X2 U4766 ( .A1(\SB2_0_26/i0_3 ), .A2(\SB2_0_26/i0[10] ), .A3(
        \SB2_0_26/i0[6] ), .ZN(\SB2_0_26/Component_Function_2/NAND4_in[1] ) );
  BUF_X2 U148 ( .I(Key[80]), .Z(n193) );
  BUF_X2 U17 ( .I(Key[69]), .Z(n183) );
  NAND3_X2 U5072 ( .A1(\SB2_0_28/i0_0 ), .A2(\RI3[0][22] ), .A3(
        \SB2_0_28/i1_5 ), .ZN(n1443) );
  NAND3_X2 U8695 ( .A1(\SB1_3_26/i0[9] ), .A2(\SB1_3_26/i0[10] ), .A3(
        \SB1_3_26/i0_3 ), .ZN(\SB1_3_26/Component_Function_4/NAND4_in[2] ) );
  NAND2_X1 U4990 ( .A1(\SB1_2_0/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_0/Component_Function_4/NAND4_in[1] ), .ZN(n1950) );
  NAND3_X2 U2893 ( .A1(\SB1_3_29/i1[9] ), .A2(\SB1_3_29/i0_3 ), .A3(
        \SB1_3_29/i0_4 ), .ZN(n2712) );
  CLKBUF_X4 U7569 ( .I(\MC_ARK_ARC_1_2/buf_output[14] ), .Z(\RI1[3][14] ) );
  INV_X2 \SB2_2_29/INV_1  ( .I(\SB1_2_1/buf_output[1] ), .ZN(\SB2_2_29/i1_7 )
         );
  NAND3_X2 \SB2_0_1/Component_Function_3/N3  ( .A1(\SB2_0_1/i1[9] ), .A2(
        \SB2_0_1/i1_7 ), .A3(\SB2_0_1/i0[10] ), .ZN(
        \SB2_0_1/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U1697 ( .A1(\SB1_0_3/i0_3 ), .A2(\SB1_0_3/i0_4 ), .A3(
        \SB1_0_3/i1[9] ), .ZN(\SB1_0_3/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 \SB1_1_17/Component_Function_4/N1  ( .A1(\SB1_1_17/i0[9] ), .A2(
        \SB1_1_17/i0_0 ), .A3(\SB1_1_17/i0[8] ), .ZN(
        \SB1_1_17/Component_Function_4/NAND4_in[0] ) );
  BUF_X4 \SB1_2_10/BUF_3  ( .I(\MC_ARK_ARC_1_1/buf_output[129] ), .Z(
        \SB1_2_10/i0[10] ) );
  CLKBUF_X4 \SB2_3_4/BUF_3  ( .I(\SB1_3_6/buf_output[3] ), .Z(\SB2_3_4/i0[10] ) );
  INV_X2 \SB2_1_17/INV_1  ( .I(\SB1_1_21/buf_output[1] ), .ZN(\SB2_1_17/i1_7 )
         );
  INV_X2 \SB1_1_2/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[175] ), .ZN(
        \SB1_1_2/i1_7 ) );
  NAND3_X2 U2392 ( .A1(\SB2_0_17/i0_3 ), .A2(\SB2_0_17/i1[9] ), .A3(
        \RI3[0][88] ), .ZN(\SB2_0_17/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3521 ( .A1(\SB2_1_26/i0[10] ), .A2(\SB2_1_26/i0_3 ), .A3(
        \SB2_1_26/i0_4 ), .ZN(n4075) );
  NAND3_X2 \SB2_3_29/Component_Function_1/N4  ( .A1(\SB2_3_29/i1_7 ), .A2(
        \SB2_3_29/i0[8] ), .A3(\RI3[3][16] ), .ZN(
        \SB2_3_29/Component_Function_1/NAND4_in[3] ) );
  BUF_X4 U2194 ( .I(\SB3_4/buf_output[1] ), .Z(\SB4_0/i0[6] ) );
  BUF_X4 \SB1_2_11/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[124] ), .Z(
        \SB1_2_11/i0_4 ) );
  NAND3_X2 \SB1_3_8/Component_Function_2/N1  ( .A1(\SB1_3_8/i1_5 ), .A2(
        \SB1_3_8/i0[10] ), .A3(\SB1_3_8/i1[9] ), .ZN(
        \SB1_3_8/Component_Function_2/NAND4_in[0] ) );
  BUF_X4 U11078 ( .I(\MC_ARK_ARC_1_1/buf_output[35] ), .Z(\RI1[2][35] ) );
  NAND3_X2 U832 ( .A1(\SB2_2_23/i0_3 ), .A2(\SB2_2_23/i0[10] ), .A3(
        \SB2_2_23/i0[9] ), .ZN(n1860) );
  CLKBUF_X4 U3467 ( .I(\SB2_2_8/buf_output[1] ), .Z(\RI5[2][163] ) );
  NAND3_X1 U10554 ( .A1(\SB1_1_12/i0_4 ), .A2(\SB1_1_12/i1_7 ), .A3(
        \SB1_1_12/i0[8] ), .ZN(\SB1_1_12/Component_Function_1/NAND4_in[3] ) );
  BUF_X2 U37 ( .I(Key[62]), .Z(n207) );
  BUF_X4 \SB2_1_1/BUF_3  ( .I(\SB1_1_3/buf_output[3] ), .Z(\SB2_1_1/i0[10] )
         );
  CLKBUF_X4 \SB2_3_25/BUF_0  ( .I(\SB1_3_30/buf_output[0] ), .Z(
        \SB2_3_25/i0[9] ) );
  BUF_X4 U3045 ( .I(\MC_ARK_ARC_1_0/buf_output[68] ), .Z(\SB1_1_20/i0_0 ) );
  BUF_X4 U3457 ( .I(\MC_ARK_ARC_1_0/buf_output[146] ), .Z(\SB1_1_7/i0_0 ) );
  BUF_X4 \SB3_4/BUF_4  ( .I(\MC_ARK_ARC_1_3/buf_output[166] ), .Z(\SB3_4/i0_4 ) );
  BUF_X4 \SB2_1_18/BUF_3  ( .I(\SB1_1_20/buf_output[3] ), .Z(\SB2_1_18/i0[10] ) );
  CLKBUF_X4 U652 ( .I(\MC_ARK_ARC_1_3/buf_output[136] ), .Z(\SB3_9/i0_4 ) );
  BUF_X2 U76 ( .I(Key[40]), .Z(n169) );
  CLKBUF_X4 \SB4_2/BUF_1  ( .I(\SB3_6/buf_output[1] ), .Z(\SB4_2/i0[6] ) );
  BUF_X2 U54 ( .I(Key[173]), .Z(n220) );
  CLKBUF_X4 U2307 ( .I(\MC_ARK_ARC_1_3/buf_output[45] ), .Z(\SB3_24/i0[10] )
         );
  BUF_X4 \SB1_0_21/BUF_2  ( .I(n277), .Z(\SB1_0_21/i0_0 ) );
  CLKBUF_X4 \SB1_2_29/BUF_2  ( .I(\MC_ARK_ARC_1_1/buf_output[14] ), .Z(
        \SB1_2_29/i0_0 ) );
  CLKBUF_X4 U7216 ( .I(\SB2_3_24/buf_output[3] ), .Z(\RI5[3][57] ) );
  CLKBUF_X2 U18 ( .I(Key[39]), .Z(n206) );
  NAND2_X2 \SB1_2_29/Component_Function_5/N1  ( .A1(\SB1_2_29/i0_0 ), .A2(
        \SB1_2_29/i3[0] ), .ZN(\SB1_2_29/Component_Function_5/NAND4_in[0] ) );
  INV_X2 \SB2_3_23/INV_1  ( .I(\SB1_3_27/buf_output[1] ), .ZN(\SB2_3_23/i1_7 )
         );
  INV_X1 U289 ( .I(n143), .ZN(n456) );
  BUF_X4 U4623 ( .I(\SB2_1_16/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[105] ) );
  NAND3_X2 \SB2_1_26/Component_Function_2/N1  ( .A1(\SB2_1_26/i1_5 ), .A2(
        \SB2_1_26/i0[10] ), .A3(\SB2_1_26/i1[9] ), .ZN(
        \SB2_1_26/Component_Function_2/NAND4_in[0] ) );
  CLKBUF_X2 U69 ( .I(Key[8]), .Z(n214) );
  BUF_X4 \SB3_5/BUF_3  ( .I(\MC_ARK_ARC_1_3/buf_output[159] ), .Z(
        \SB3_5/i0[10] ) );
  INV_X4 \SB1_2_4/INV_5  ( .I(\RI1[2][167] ), .ZN(\SB1_2_4/i1_5 ) );
  NAND3_X2 U2093 ( .A1(n3687), .A2(\SB2_2_9/i0_0 ), .A3(\SB2_2_9/i0_4 ), .ZN(
        \SB2_2_9/Component_Function_2/NAND4_in[3] ) );
  NAND2_X2 U768 ( .A1(\SB1_3_8/Component_Function_2/NAND4_in[3] ), .A2(
        \SB1_3_8/Component_Function_2/NAND4_in[2] ), .ZN(n3412) );
  NAND2_X2 U3242 ( .A1(n606), .A2(\SB1_3_8/Component_Function_4/NAND4_in[0] ), 
        .ZN(n3740) );
  BUF_X4 U4653 ( .I(\MC_ARK_ARC_1_3/buf_output[147] ), .Z(\SB3_7/i0[10] ) );
  NAND3_X1 U716 ( .A1(\SB2_3_26/i0_3 ), .A2(\SB1_3_28/buf_output[3] ), .A3(
        \SB2_3_26/i0[6] ), .ZN(\SB2_3_26/Component_Function_2/NAND4_in[1] ) );
  CLKBUF_X2 U29 ( .I(Key[46]), .Z(n234) );
  NAND3_X2 \SB1_0_22/Component_Function_5/N3  ( .A1(\SB1_0_22/i1[9] ), .A2(
        \SB1_0_22/i0_4 ), .A3(\SB1_0_22/i0_3 ), .ZN(
        \SB1_0_22/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 \SB2_0_17/Component_Function_2/N1  ( .A1(\SB2_0_17/i1_5 ), .A2(
        \SB2_0_17/i0[10] ), .A3(\SB2_0_17/i1[9] ), .ZN(
        \SB2_0_17/Component_Function_2/NAND4_in[0] ) );
  NAND2_X2 \SB2_0_31/Component_Function_5/N1  ( .A1(\SB2_0_31/i0_0 ), .A2(
        \SB2_0_31/i3[0] ), .ZN(\SB2_0_31/Component_Function_5/NAND4_in[0] ) );
  NAND2_X2 U2772 ( .A1(\SB3_19/i0_0 ), .A2(\SB3_19/i3[0] ), .ZN(
        \SB3_19/Component_Function_5/NAND4_in[0] ) );
  NAND2_X2 \SB2_2_25/Component_Function_5/N1  ( .A1(\SB2_2_25/i0_0 ), .A2(
        \SB2_2_25/i3[0] ), .ZN(\SB2_2_25/Component_Function_5/NAND4_in[0] ) );
  NAND3_X2 U5821 ( .A1(\SB2_0_29/i0_3 ), .A2(\SB2_0_29/i0[6] ), .A3(
        \RI3[0][15] ), .ZN(n1903) );
  CLKBUF_X4 \SB2_2_9/BUF_2  ( .I(\SB1_2_12/buf_output[2] ), .Z(\SB2_2_9/i0_0 )
         );
  CLKBUF_X4 U8819 ( .I(\SB1_3_16/buf_output[3] ), .Z(\SB2_3_14/i0[10] ) );
  CLKBUF_X4 U3341 ( .I(n371), .Z(\SB1_0_16/i0[10] ) );
  CLKBUF_X4 \SB1_0_23/BUF_3  ( .I(n357), .Z(\SB1_0_23/i0[10] ) );
  CLKBUF_X4 U1696 ( .I(n253), .Z(\SB1_0_29/i0_0 ) );
  CLKBUF_X4 \SB1_0_2/BUF_3  ( .I(n399), .Z(\SB1_0_2/i0[10] ) );
  CLKBUF_X4 U2699 ( .I(n289), .Z(\SB1_0_17/i0_0 ) );
  CLKBUF_X4 \SB1_0_12/BUF_3  ( .I(n379), .Z(\SB1_0_12/i0[10] ) );
  CLKBUF_X4 U1931 ( .I(n356), .Z(\SB1_0_24/i0_4 ) );
  CLKBUF_X4 U4716 ( .I(n334), .Z(\SB1_0_2/i0_0 ) );
  CLKBUF_X4 U8122 ( .I(n274), .Z(\SB1_0_22/i0_0 ) );
  CLKBUF_X4 \SB1_0_28/BUF_2  ( .I(n256), .Z(\SB1_0_28/i0_0 ) );
  CLKBUF_X4 \SB1_0_18/BUF_2  ( .I(n286), .Z(\SB1_0_18/i0_0 ) );
  CLKBUF_X4 \SB1_0_22/BUF_4  ( .I(n360), .Z(\SB1_0_22/i0_4 ) );
  CLKBUF_X4 \SB1_0_11/BUF_5  ( .I(n425), .Z(\SB1_0_11/i0_3 ) );
  CLKBUF_X4 \SB1_0_7/BUF_2  ( .I(n319), .Z(\SB1_0_7/i0_0 ) );
  CLKBUF_X4 \SB1_0_31/BUF_1  ( .I(n246), .Z(\SB1_0_31/i0[6] ) );
  CLKBUF_X4 \SB1_0_9/BUF_1  ( .I(n312), .Z(\SB1_0_9/i0[6] ) );
  CLKBUF_X4 \SB1_0_11/BUF_4  ( .I(n382), .Z(\SB1_0_11/i0_4 ) );
  CLKBUF_X4 \SB1_0_16/BUF_1  ( .I(n291), .Z(\SB1_0_16/i0[6] ) );
  INV_X1 U344 ( .I(n68), .ZN(n534) );
  CLKBUF_X4 \SB1_0_8/BUF_3  ( .I(n387), .Z(\SB1_0_8/i0[10] ) );
  CLKBUF_X4 U3326 ( .I(n353), .Z(\SB1_0_25/i0[10] ) );
  CLKBUF_X4 U3064 ( .I(n301), .Z(\SB1_0_13/i0_0 ) );
  INV_X1 U4 ( .I(n176), .ZN(n531) );
  INV_X1 U269 ( .I(n24), .ZN(n439) );
  CLKBUF_X4 \SB1_0_5/BUF_1  ( .I(n324), .Z(\SB1_0_5/i0[6] ) );
  CLKBUF_X4 \SB1_0_3/BUF_3  ( .I(n397), .Z(\SB1_0_3/i0[10] ) );
  CLKBUF_X4 \SB1_0_5/BUF_4  ( .I(n394), .Z(\SB1_0_5/i0_4 ) );
  CLKBUF_X4 \SB1_0_3/BUF_2  ( .I(n331), .Z(\SB1_0_3/i0_0 ) );
  CLKBUF_X4 U1936 ( .I(n378), .Z(\SB1_0_13/i0_4 ) );
  CLKBUF_X4 \SB1_0_14/BUF_0  ( .I(n296), .Z(\SB1_0_14/i0[9] ) );
  CLKBUF_X4 \SB1_0_15/BUF_3  ( .I(n373), .Z(\SB1_0_15/i0[10] ) );
  INV_X1 U3731 ( .I(n5), .ZN(n494) );
  NAND2_X1 U5707 ( .A1(\SB1_0_2/Component_Function_4/NAND4_in[1] ), .A2(n2482), 
        .ZN(n2481) );
  CLKBUF_X4 \SB2_0_22/BUF_4  ( .I(\RI3[0][58] ), .Z(\SB2_0_22/i0_4 ) );
  BUF_X2 \SB2_0_6/BUF_0  ( .I(\SB1_0_11/buf_output[0] ), .Z(\SB2_0_6/i0[9] )
         );
  CLKBUF_X4 \SB2_0_0/BUF_2  ( .I(\RI3[0][188] ), .Z(\SB2_0_0/i0_0 ) );
  CLKBUF_X4 \SB2_0_25/BUF_2  ( .I(\SB1_0_28/buf_output[2] ), .Z(
        \SB2_0_25/i0_0 ) );
  CLKBUF_X4 U1920 ( .I(\SB1_0_1/buf_output[4] ), .Z(\RI3[0][190] ) );
  CLKBUF_X4 U1923 ( .I(\SB2_0_6/i0[10] ), .Z(n2765) );
  CLKBUF_X4 \SB2_0_18/BUF_1  ( .I(\RI3[0][79] ), .Z(\SB2_0_18/i0[6] ) );
  CLKBUF_X2 U1925 ( .I(\SB2_0_27/i0[9] ), .Z(n1091) );
  CLKBUF_X4 U1927 ( .I(\RI3[0][126] ), .Z(n571) );
  CLKBUF_X4 \SB2_0_7/BUF_2  ( .I(\RI3[0][146] ), .Z(\SB2_0_7/i0_0 ) );
  CLKBUF_X4 \SB2_0_22/BUF_2  ( .I(\SB1_0_25/buf_output[2] ), .Z(
        \SB2_0_22/i0_0 ) );
  BUF_X2 \SB2_0_26/BUF_1  ( .I(\SB1_0_30/buf_output[1] ), .Z(\SB2_0_26/i0[6] )
         );
  CLKBUF_X4 \SB2_0_18/BUF_3  ( .I(\RI3[0][81] ), .Z(\SB2_0_18/i0[10] ) );
  CLKBUF_X4 \SB2_0_3/BUF_2  ( .I(\SB1_0_6/buf_output[2] ), .Z(\SB2_0_3/i0_0 )
         );
  CLKBUF_X4 \SB2_0_23/BUF_3  ( .I(\SB1_0_25/buf_output[3] ), .Z(
        \SB2_0_23/i0[10] ) );
  CLKBUF_X4 \SB2_0_27/BUF_3  ( .I(\RI3[0][27] ), .Z(\SB2_0_27/i0[10] ) );
  BUF_X2 U1623 ( .I(\RI3[0][49] ), .Z(\SB2_0_23/i0[6] ) );
  CLKBUF_X4 \SB2_0_11/BUF_3  ( .I(\RI3[0][123] ), .Z(\SB2_0_11/i0[10] ) );
  CLKBUF_X4 \SB2_0_21/BUF_3  ( .I(\RI3[0][63] ), .Z(\SB2_0_21/i0[10] ) );
  CLKBUF_X4 U1653 ( .I(\SB1_0_21/buf_output[5] ), .Z(\SB2_0_21/i0_3 ) );
  CLKBUF_X4 \SB2_0_9/BUF_3  ( .I(\SB1_0_11/buf_output[3] ), .Z(
        \SB2_0_9/i0[10] ) );
  CLKBUF_X4 \SB2_0_16/BUF_3  ( .I(\RI3[0][93] ), .Z(\SB2_0_16/i0[10] ) );
  CLKBUF_X4 U1628 ( .I(\SB1_0_30/buf_output[2] ), .Z(\SB2_0_27/i0_0 ) );
  CLKBUF_X4 \SB2_0_28/BUF_2  ( .I(\RI3[0][20] ), .Z(\SB2_0_28/i0_0 ) );
  CLKBUF_X4 \SB2_0_8/BUF_1  ( .I(\RI3[0][139] ), .Z(\SB2_0_8/i0[6] ) );
  CLKBUF_X4 \SB2_0_16/BUF_1  ( .I(\RI3[0][91] ), .Z(\SB2_0_16/i0[6] ) );
  CLKBUF_X4 \SB2_0_1/BUF_1  ( .I(\SB1_0_5/buf_output[1] ), .Z(\SB2_0_1/i0[6] )
         );
  CLKBUF_X4 U4763 ( .I(\SB1_0_26/buf_output[5] ), .Z(\SB2_0_26/i0_3 ) );
  CLKBUF_X4 \SB2_0_20/BUF_1  ( .I(\RI3[0][67] ), .Z(\SB2_0_20/i0[6] ) );
  CLKBUF_X4 \SB2_0_20/BUF_5  ( .I(\SB1_0_20/buf_output[5] ), .Z(
        \SB2_0_20/i0_3 ) );
  CLKBUF_X4 \SB2_0_3/BUF_0  ( .I(\SB1_0_8/buf_output[0] ), .Z(\SB2_0_3/i0[9] )
         );
  CLKBUF_X4 U4836 ( .I(\RI3[0][161] ), .Z(\SB2_0_5/i0_3 ) );
  CLKBUF_X4 \SB2_0_21/BUF_1  ( .I(\RI3[0][61] ), .Z(\SB2_0_21/i0[6] ) );
  CLKBUF_X4 \SB2_0_30/BUF_2  ( .I(\RI3[0][8] ), .Z(\SB2_0_30/i0_0 ) );
  CLKBUF_X4 U1756 ( .I(\SB2_0_18/buf_output[3] ), .Z(\RI5[0][93] ) );
  CLKBUF_X4 \SB2_0_31/BUF_2_0  ( .I(\SB2_0_31/buf_output[2] ), .Z(\RI5[0][20] ) );
  CLKBUF_X4 \MC_ARK_ARC_1_0/BUF_166  ( .I(\SB2_0_5/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[166] ) );
  CLKBUF_X4 U1915 ( .I(\SB2_0_28/buf_output[3] ), .Z(\RI5[0][33] ) );
  CLKBUF_X4 \SB2_0_9/BUF_5_0  ( .I(\SB2_0_9/buf_output[5] ), .Z(\RI5[0][137] )
         );
  CLKBUF_X4 \SB2_0_12/BUF_3_0  ( .I(\SB2_0_12/buf_output[3] ), .Z(
        \RI5[0][129] ) );
  CLKBUF_X4 U7999 ( .I(\SB2_0_27/buf_output[4] ), .Z(\RI5[0][34] ) );
  BUF_X2 U3838 ( .I(\SB2_0_17/buf_output[0] ), .Z(\RI5[0][114] ) );
  CLKBUF_X4 \SB2_0_14/BUF_1_0  ( .I(\SB2_0_14/buf_output[1] ), .Z(
        \RI5[0][127] ) );
  CLKBUF_X4 U2629 ( .I(\SB2_0_13/buf_output[2] ), .Z(\RI5[0][128] ) );
  CLKBUF_X4 \SB2_0_10/BUF_1_0  ( .I(\SB2_0_10/buf_output[1] ), .Z(
        \RI5[0][151] ) );
  CLKBUF_X4 U3415 ( .I(\SB2_0_6/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[165] ) );
  BUF_X4 \SB2_0_2/BUF_4_0  ( .I(\SB2_0_2/buf_output[4] ), .Z(\RI5[0][184] ) );
  CLKBUF_X4 \SB2_0_7/BUF_3_0  ( .I(\SB2_0_7/buf_output[3] ), .Z(\RI5[0][159] )
         );
  CLKBUF_X4 U1911 ( .I(\SB2_0_25/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[56] ) );
  CLKBUF_X4 \SB2_0_2/BUF_3_0  ( .I(\SB2_0_2/buf_output[3] ), .Z(\RI5[0][189] )
         );
  CLKBUF_X4 \MC_ARK_ARC_1_0/BUF_51  ( .I(\SB2_0_25/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[51] ) );
  CLKBUF_X4 U8740 ( .I(\SB2_0_7/buf_output[1] ), .Z(\RI5[0][169] ) );
  CLKBUF_X4 U1504 ( .I(\MC_ARK_ARC_1_0/buf_output[58] ), .Z(\SB1_1_22/i0_4 )
         );
  CLKBUF_X4 \SB1_1_28/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[19] ), .Z(
        \SB1_1_28/i0[6] ) );
  CLKBUF_X4 \SB1_1_5/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[157] ), .Z(
        \SB1_1_5/i0[6] ) );
  CLKBUF_X4 \SB1_1_24/BUF_3  ( .I(\MC_ARK_ARC_1_0/buf_output[45] ), .Z(
        \SB1_1_24/i0[10] ) );
  CLKBUF_X4 \SB1_1_8/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[142] ), .Z(
        \SB1_1_8/i0_4 ) );
  CLKBUF_X4 U1633 ( .I(\MC_ARK_ARC_1_0/buf_output[139] ), .Z(\SB1_1_8/i0[6] )
         );
  CLKBUF_X4 U1645 ( .I(\MC_ARK_ARC_1_0/buf_output[9] ), .Z(\SB1_1_30/i0[10] )
         );
  CLKBUF_X4 \SB1_1_13/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[112] ), .Z(
        \SB1_1_13/i0_4 ) );
  CLKBUF_X4 U4809 ( .I(\MC_ARK_ARC_1_0/buf_output[122] ), .Z(\SB1_1_11/i0_0 )
         );
  CLKBUF_X4 \SB1_1_4/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[166] ), .Z(
        \SB1_1_4/i0_4 ) );
  CLKBUF_X4 U1060 ( .I(\MC_ARK_ARC_1_0/buf_output[121] ), .Z(\SB1_1_11/i0[6] )
         );
  CLKBUF_X4 U1480 ( .I(\MC_ARK_ARC_1_0/buf_output[85] ), .Z(\SB1_1_17/i0[6] )
         );
  CLKBUF_X4 U8812 ( .I(\MC_ARK_ARC_1_0/buf_output[171] ), .Z(\SB1_1_3/i0[10] )
         );
  CLKBUF_X4 \SB1_1_2/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[178] ), .Z(
        \SB1_1_2/i0_4 ) );
  CLKBUF_X4 U8802 ( .I(\MC_ARK_ARC_1_0/buf_output[92] ), .Z(\SB1_1_16/i0_0 )
         );
  CLKBUF_X4 \SB1_1_29/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[16] ), .Z(
        \SB1_1_29/i0_4 ) );
  CLKBUF_X4 \SB1_1_0/BUF_3  ( .I(\MC_ARK_ARC_1_0/buf_output[189] ), .Z(
        \SB1_1_0/i0[10] ) );
  CLKBUF_X4 \SB1_1_3/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[172] ), .Z(
        \SB1_1_3/i0_4 ) );
  CLKBUF_X4 \SB1_1_26/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[30] ), .Z(
        \SB1_1_26/i0[9] ) );
  CLKBUF_X4 U3301 ( .I(\MC_ARK_ARC_1_0/buf_output[175] ), .Z(\SB1_1_2/i0[6] )
         );
  CLKBUF_X4 U4773 ( .I(\MC_ARK_ARC_1_0/buf_output[98] ), .Z(\SB1_1_15/i0_0 )
         );
  CLKBUF_X4 U4963 ( .I(\MC_ARK_ARC_1_0/buf_output[32] ), .Z(\SB1_1_26/i0_0 )
         );
  CLKBUF_X4 \SB1_1_20/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[67] ), .Z(
        \SB1_1_20/i0[6] ) );
  CLKBUF_X4 U2427 ( .I(\MC_ARK_ARC_1_0/buf_output[168] ), .Z(\SB1_1_3/i0[9] )
         );
  CLKBUF_X4 \SB1_1_15/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[100] ), .Z(
        \SB1_1_15/i0_4 ) );
  CLKBUF_X4 \SB1_1_27/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[28] ), .Z(
        \SB1_1_27/i0_4 ) );
  CLKBUF_X4 U8879 ( .I(\MC_ARK_ARC_1_0/buf_output[84] ), .Z(\SB1_1_17/i0[9] )
         );
  CLKBUF_X4 U4699 ( .I(\MC_ARK_ARC_1_0/buf_output[123] ), .Z(\SB1_1_11/i0[10] ) );
  CLKBUF_X4 \SB1_1_21/BUF_2  ( .I(\MC_ARK_ARC_1_0/buf_output[62] ), .Z(
        \SB1_1_21/i0_0 ) );
  CLKBUF_X4 \SB1_1_29/BUF_3  ( .I(\MC_ARK_ARC_1_0/buf_output[15] ), .Z(
        \SB1_1_29/i0[10] ) );
  CLKBUF_X4 U1503 ( .I(\MC_ARK_ARC_1_0/buf_output[12] ), .Z(\SB1_1_29/i0[9] )
         );
  CLKBUF_X4 U3015 ( .I(\MC_ARK_ARC_1_0/buf_output[20] ), .Z(\SB1_1_28/i0_0 )
         );
  CLKBUF_X4 U2356 ( .I(\MC_ARK_ARC_1_0/buf_output[86] ), .Z(\SB1_1_17/i0_0 )
         );
  CLKBUF_X4 \SB1_1_14/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[103] ), .Z(
        \SB1_1_14/i0[6] ) );
  CLKBUF_X4 \SB1_1_30/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[10] ), .Z(
        \SB1_1_30/i0_4 ) );
  CLKBUF_X4 \SB1_1_3/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[169] ), .Z(
        \SB1_1_3/i0[6] ) );
  CLKBUF_X4 U2937 ( .I(\MC_ARK_ARC_1_0/buf_output[72] ), .Z(\SB1_1_19/i0[9] )
         );
  CLKBUF_X4 \SB1_1_4/BUF_3  ( .I(\MC_ARK_ARC_1_0/buf_output[165] ), .Z(
        \SB1_1_4/i0[10] ) );
  CLKBUF_X4 \SB1_1_16/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[91] ), .Z(
        \SB1_1_16/i0[6] ) );
  CLKBUF_X4 \SB1_1_8/BUF_0  ( .I(\MC_ARK_ARC_1_0/buf_output[138] ), .Z(
        \SB1_1_8/i0[9] ) );
  NAND2_X1 U10509 ( .A1(n4700), .A2(n1775), .ZN(n4427) );
  CLKBUF_X4 U2722 ( .I(\SB1_1_28/buf_output[3] ), .Z(\SB2_1_26/i0[10] ) );
  CLKBUF_X4 U3285 ( .I(\SB1_1_23/buf_output[1] ), .Z(\SB2_1_19/i0[6] ) );
  CLKBUF_X4 \SB2_1_26/BUF_2  ( .I(\SB1_1_29/buf_output[2] ), .Z(
        \SB2_1_26/i0_0 ) );
  CLKBUF_X4 \SB2_1_21/BUF_2  ( .I(\SB1_1_24/buf_output[2] ), .Z(
        \SB2_1_21/i0_0 ) );
  CLKBUF_X4 \SB2_1_20/BUF_0  ( .I(\SB1_1_25/buf_output[0] ), .Z(
        \SB2_1_20/i0[9] ) );
  CLKBUF_X4 \SB2_1_26/BUF_4  ( .I(\SB1_1_27/buf_output[4] ), .Z(
        \SB2_1_26/i0_4 ) );
  CLKBUF_X4 \SB2_1_27/BUF_3  ( .I(\SB1_1_29/buf_output[3] ), .Z(
        \SB2_1_27/i0[10] ) );
  CLKBUF_X4 U9046 ( .I(\SB1_1_0/buf_output[2] ), .Z(\SB2_1_29/i0_0 ) );
  CLKBUF_X4 \SB2_1_9/BUF_4  ( .I(\SB1_1_10/buf_output[4] ), .Z(\SB2_1_9/i0_4 )
         );
  CLKBUF_X4 \SB2_1_9/BUF_0  ( .I(\SB1_1_14/buf_output[0] ), .Z(\SB2_1_9/i0[9] ) );
  NAND2_X1 U5924 ( .A1(n2728), .A2(\SB1_1_22/Component_Function_1/NAND4_in[2] ), .ZN(n3278) );
  CLKBUF_X4 \SB2_1_13/BUF_3  ( .I(\SB1_1_15/buf_output[3] ), .Z(
        \SB2_1_13/i0[10] ) );
  CLKBUF_X4 \SB2_1_10/BUF_1  ( .I(\SB1_1_14/buf_output[1] ), .Z(
        \SB2_1_10/i0[6] ) );
  CLKBUF_X4 \SB2_1_29/BUF_3  ( .I(\SB1_1_31/buf_output[3] ), .Z(
        \SB2_1_29/i0[10] ) );
  CLKBUF_X4 U2017 ( .I(\SB1_1_9/buf_output[3] ), .Z(\SB2_1_7/i0[10] ) );
  BUF_X2 \SB2_1_31/BUF_0  ( .I(\SB1_1_4/buf_output[0] ), .Z(\SB2_1_31/i0[9] )
         );
  CLKBUF_X4 \SB2_1_1/BUF_0  ( .I(\SB1_1_6/buf_output[0] ), .Z(\SB2_1_1/i0[9] )
         );
  CLKBUF_X4 \SB2_1_12/BUF_3  ( .I(\SB1_1_14/buf_output[3] ), .Z(
        \SB2_1_12/i0[10] ) );
  CLKBUF_X4 \SB2_1_2/BUF_1  ( .I(\SB1_1_6/buf_output[1] ), .Z(\SB2_1_2/i0[6] )
         );
  CLKBUF_X4 \SB2_1_2/BUF_0  ( .I(\SB1_1_7/buf_output[0] ), .Z(\SB2_1_2/i0[9] )
         );
  CLKBUF_X4 \SB2_1_4/BUF_3  ( .I(\SB1_1_6/buf_output[3] ), .Z(\SB2_1_4/i0[10] ) );
  CLKBUF_X4 \SB2_1_13/BUF_4  ( .I(\SB1_1_14/buf_output[4] ), .Z(
        \SB2_1_13/i0_4 ) );
  CLKBUF_X4 \SB2_1_12/BUF_0  ( .I(\SB1_1_17/buf_output[0] ), .Z(
        \SB2_1_12/i0[9] ) );
  CLKBUF_X4 \SB2_1_0/BUF_0  ( .I(\SB1_1_5/buf_output[0] ), .Z(\SB2_1_0/i0[9] )
         );
  CLKBUF_X4 \SB2_1_11/BUF_2  ( .I(\SB1_1_14/buf_output[2] ), .Z(
        \SB2_1_11/i0_0 ) );
  CLKBUF_X4 \SB2_1_20/BUF_2  ( .I(\SB1_1_23/buf_output[2] ), .Z(
        \SB2_1_20/i0_0 ) );
  CLKBUF_X4 U8774 ( .I(\SB1_1_3/buf_output[2] ), .Z(\SB2_1_0/i0_0 ) );
  CLKBUF_X4 \SB2_1_17/BUF_1  ( .I(\SB1_1_21/buf_output[1] ), .Z(
        \SB2_1_17/i0[6] ) );
  CLKBUF_X4 U8720 ( .I(\SB1_1_16/buf_output[3] ), .Z(\SB2_1_14/i0[10] ) );
  CLKBUF_X4 \SB2_1_17/BUF_4  ( .I(\SB1_1_18/buf_output[4] ), .Z(
        \SB2_1_17/i0_4 ) );
  CLKBUF_X4 \SB2_1_28/BUF_2  ( .I(\SB1_1_31/buf_output[2] ), .Z(
        \SB2_1_28/i0_0 ) );
  CLKBUF_X4 U3284 ( .I(\SB1_1_27/buf_output[2] ), .Z(\SB2_1_24/i0_0 ) );
  CLKBUF_X4 \SB2_1_23/BUF_1  ( .I(\SB1_1_27/buf_output[1] ), .Z(
        \SB2_1_23/i0[6] ) );
  CLKBUF_X4 U3507 ( .I(\SB1_1_19/buf_output[3] ), .Z(\SB2_1_17/i0[10] ) );
  CLKBUF_X4 U992 ( .I(\SB1_1_11/buf_output[1] ), .Z(n2852) );
  CLKBUF_X4 \SB2_1_6/BUF_2  ( .I(\SB1_1_9/buf_output[2] ), .Z(\SB2_1_6/i0_0 )
         );
  BUF_X2 \SB2_1_3/BUF_0  ( .I(\SB1_1_8/buf_output[0] ), .Z(\SB2_1_3/i0[9] ) );
  CLKBUF_X4 \SB2_1_25/BUF_3  ( .I(\SB1_1_27/buf_output[3] ), .Z(
        \SB2_1_25/i0[10] ) );
  CLKBUF_X4 \SB2_1_15/BUF_3  ( .I(\SB1_1_17/buf_output[3] ), .Z(
        \SB2_1_15/i0[10] ) );
  CLKBUF_X4 U2019 ( .I(\SB1_1_7/buf_output[4] ), .Z(\SB2_1_6/i0_4 ) );
  CLKBUF_X4 \SB2_1_3/BUF_1  ( .I(\SB1_1_7/buf_output[1] ), .Z(\SB2_1_3/i0[6] )
         );
  CLKBUF_X4 U8842 ( .I(\SB1_1_24/buf_output[0] ), .Z(\SB2_1_19/i0[9] ) );
  BUF_X4 U2031 ( .I(\SB1_1_3/buf_output[5] ), .Z(\SB2_1_3/i0_3 ) );
  CLKBUF_X4 U8883 ( .I(\SB1_1_9/buf_output[1] ), .Z(\SB2_1_5/i0[6] ) );
  CLKBUF_X4 \SB2_1_8/BUF_4  ( .I(\SB1_1_9/buf_output[4] ), .Z(\SB2_1_8/i0_4 )
         );
  CLKBUF_X4 U4860 ( .I(\SB1_1_7/buf_output[3] ), .Z(\SB2_1_5/i0[10] ) );
  CLKBUF_X4 \SB2_1_5/BUF_0  ( .I(\SB1_1_10/buf_output[0] ), .Z(\SB2_1_5/i0[9] ) );
  CLKBUF_X4 U4693 ( .I(\SB1_1_23/buf_output[0] ), .Z(\SB2_1_18/i0[9] ) );
  CLKBUF_X4 \SB2_1_14/BUF_0  ( .I(\SB1_1_19/buf_output[0] ), .Z(
        \SB2_1_14/i0[9] ) );
  BUF_X4 U3814 ( .I(\SB1_1_19/buf_output[4] ), .Z(\SB2_1_18/i0_4 ) );
  CLKBUF_X4 \SB2_1_7/BUF_2  ( .I(\SB1_1_10/buf_output[2] ), .Z(\SB2_1_7/i0_0 )
         );
  CLKBUF_X4 \SB2_1_27/BUF_2  ( .I(\SB1_1_30/buf_output[2] ), .Z(
        \SB2_1_27/i0_0 ) );
  CLKBUF_X2 U10999 ( .I(\SB2_1_21/i3[0] ), .Z(n4625) );
  CLKBUF_X4 \SB2_1_19/BUF_3  ( .I(\SB1_1_21/buf_output[3] ), .Z(
        \SB2_1_19/i0[10] ) );
  CLKBUF_X4 U4915 ( .I(\SB1_1_8/buf_output[3] ), .Z(\SB2_1_6/i0[10] ) );
  CLKBUF_X4 U1895 ( .I(\SB2_1_2/buf_output[1] ), .Z(\RI5[1][7] ) );
  CLKBUF_X4 U8610 ( .I(\SB2_1_17/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[99] ) );
  CLKBUF_X4 \SB2_1_6/BUF_3_0  ( .I(\SB2_1_6/buf_output[3] ), .Z(\RI5[1][165] )
         );
  CLKBUF_X4 U5456 ( .I(\SB2_1_30/buf_output[3] ), .Z(\RI5[1][21] ) );
  CLKBUF_X4 U3276 ( .I(\SB2_1_6/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[170] ) );
  CLKBUF_X4 U7811 ( .I(\SB2_1_4/buf_output[2] ), .Z(\RI5[1][182] ) );
  CLKBUF_X4 U3277 ( .I(\SB2_1_27/buf_output[4] ), .Z(\RI5[1][34] ) );
  BUF_X4 U3533 ( .I(\SB2_1_13/buf_output[1] ), .Z(\RI5[1][133] ) );
  CLKBUF_X4 U7986 ( .I(\SB2_1_3/buf_output[3] ), .Z(\RI5[1][183] ) );
  CLKBUF_X4 U3551 ( .I(\MC_ARK_ARC_1_1/buf_output[159] ), .Z(\SB1_2_5/i0[10] )
         );
  CLKBUF_X4 \SB1_2_8/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[139] ), .Z(
        \SB1_2_8/i0[6] ) );
  CLKBUF_X4 U4953 ( .I(\MC_ARK_ARC_1_1/buf_output[165] ), .Z(\SB1_2_4/i0[10] )
         );
  CLKBUF_X4 \SB1_2_18/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[78] ), .Z(
        \SB1_2_18/i0[9] ) );
  CLKBUF_X4 \SB1_2_22/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[58] ), .Z(
        \SB1_2_22/i0_4 ) );
  CLKBUF_X4 \SB1_2_15/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[100] ), .Z(
        \SB1_2_15/i0_4 ) );
  CLKBUF_X4 U1539 ( .I(\MC_ARK_ARC_1_1/buf_output[15] ), .Z(\SB1_2_29/i0[10] )
         );
  CLKBUF_X4 \SB1_2_5/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[160] ), .Z(
        \SB1_2_5/i0_4 ) );
  CLKBUF_X4 \SB1_2_23/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[49] ), .Z(
        \SB1_2_23/i0[6] ) );
  CLKBUF_X4 \SB1_2_25/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[40] ), .Z(
        \SB1_2_25/i0_4 ) );
  CLKBUF_X4 U2053 ( .I(\MC_ARK_ARC_1_1/buf_output[38] ), .Z(\SB1_2_25/i0_0 )
         );
  CLKBUF_X4 \SB1_2_31/BUF_2  ( .I(\MC_ARK_ARC_1_1/buf_output[2] ), .Z(
        \SB1_2_31/i0_0 ) );
  CLKBUF_X4 \SB1_2_30/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[10] ), .Z(
        \SB1_2_30/i0_4 ) );
  CLKBUF_X4 \SB1_2_10/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[127] ), .Z(
        \SB1_2_10/i0[6] ) );
  CLKBUF_X4 U1161 ( .I(\MC_ARK_ARC_1_1/buf_output[61] ), .Z(\SB1_2_21/i0[6] )
         );
  CLKBUF_X4 \SB1_2_11/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[121] ), .Z(
        \SB1_2_11/i0[6] ) );
  CLKBUF_X4 \SB1_2_0/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[186] ), .Z(
        \SB1_2_0/i0[9] ) );
  CLKBUF_X4 U2973 ( .I(\MC_ARK_ARC_1_1/buf_output[8] ), .Z(\SB1_2_30/i0_0 ) );
  CLKBUF_X4 U4147 ( .I(\MC_ARK_ARC_1_1/buf_output[164] ), .Z(\SB1_2_4/i0_0 )
         );
  CLKBUF_X4 \SB1_2_16/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[90] ), .Z(
        \SB1_2_16/i0[9] ) );
  CLKBUF_X4 U2052 ( .I(\MC_ARK_ARC_1_1/buf_output[130] ), .Z(\SB1_2_10/i0_4 )
         );
  CLKBUF_X4 \SB1_2_27/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[28] ), .Z(
        \SB1_2_27/i0_4 ) );
  CLKBUF_X4 U1674 ( .I(\MC_ARK_ARC_1_1/buf_output[20] ), .Z(\SB1_2_28/i0_0 )
         );
  CLKBUF_X4 U2058 ( .I(\MC_ARK_ARC_1_1/buf_output[34] ), .Z(\SB1_2_26/i0_4 )
         );
  CLKBUF_X4 U3518 ( .I(\MC_ARK_ARC_1_1/buf_output[177] ), .Z(\SB1_2_2/i0[10] )
         );
  CLKBUF_X4 U9041 ( .I(\MC_ARK_ARC_1_1/buf_output[156] ), .Z(\SB1_2_5/i0[9] )
         );
  CLKBUF_X4 U8877 ( .I(\MC_ARK_ARC_1_1/buf_output[21] ), .Z(\SB1_2_28/i0[10] )
         );
  CLKBUF_X4 U1888 ( .I(\MC_ARK_ARC_1_1/buf_output[92] ), .Z(\SB1_2_16/i0_0 )
         );
  CLKBUF_X4 U3844 ( .I(\MC_ARK_ARC_1_1/buf_output[33] ), .Z(\SB1_2_26/i0[10] )
         );
  CLKBUF_X4 U6526 ( .I(\MC_ARK_ARC_1_1/buf_output[26] ), .Z(\SB1_2_27/i0_0 )
         );
  CLKBUF_X8 U8716 ( .I(\RI1[2][59] ), .Z(\SB1_2_22/i0_3 ) );
  CLKBUF_X4 \SB1_2_24/BUF_4  ( .I(\MC_ARK_ARC_1_1/buf_output[46] ), .Z(
        \SB1_2_24/i0_4 ) );
  CLKBUF_X4 U2880 ( .I(\MC_ARK_ARC_1_1/buf_output[108] ), .Z(\SB1_2_13/i0[9] )
         );
  CLKBUF_X4 \SB1_2_12/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[114] ), .Z(
        \SB1_2_12/i0[9] ) );
  CLKBUF_X4 \SB1_2_25/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[36] ), .Z(
        \SB1_2_25/i0[9] ) );
  CLKBUF_X4 U1761 ( .I(\MC_ARK_ARC_1_1/buf_output[32] ), .Z(\SB1_2_26/i0_0 )
         );
  CLKBUF_X4 \SB1_2_22/BUF_3  ( .I(\MC_ARK_ARC_1_1/buf_output[57] ), .Z(
        \SB1_2_22/i0[10] ) );
  CLKBUF_X4 \SB1_2_15/BUF_3  ( .I(\MC_ARK_ARC_1_1/buf_output[99] ), .Z(
        \SB1_2_15/i0[10] ) );
  CLKBUF_X4 U8769 ( .I(\MC_ARK_ARC_1_1/buf_output[94] ), .Z(\SB1_2_16/i0_4 )
         );
  CLKBUF_X4 \SB1_2_7/BUF_3  ( .I(\MC_ARK_ARC_1_1/buf_output[147] ), .Z(
        \SB1_2_7/i0[10] ) );
  CLKBUF_X4 U2829 ( .I(\MC_ARK_ARC_1_1/buf_output[109] ), .Z(\SB1_2_13/i0[6] )
         );
  CLKBUF_X4 \SB2_2_19/BUF_3  ( .I(\SB1_2_21/buf_output[3] ), .Z(
        \SB2_2_19/i0[10] ) );
  CLKBUF_X4 \SB2_2_0/BUF_2  ( .I(\SB1_2_3/buf_output[2] ), .Z(\SB2_2_0/i0_0 )
         );
  CLKBUF_X4 \SB2_2_5/BUF_0  ( .I(\SB1_2_10/buf_output[0] ), .Z(\SB2_2_5/i0[9] ) );
  CLKBUF_X4 \SB2_2_16/BUF_2  ( .I(\SB1_2_19/buf_output[2] ), .Z(
        \SB2_2_16/i0_0 ) );
  CLKBUF_X4 \SB2_2_14/BUF_1  ( .I(\SB1_2_18/buf_output[1] ), .Z(
        \SB2_2_14/i0[6] ) );
  CLKBUF_X4 \SB2_2_7/BUF_2  ( .I(\SB1_2_10/buf_output[2] ), .Z(\SB2_2_7/i0_0 )
         );
  CLKBUF_X4 \SB2_2_26/BUF_1  ( .I(\SB1_2_30/buf_output[1] ), .Z(
        \SB2_2_26/i0[6] ) );
  CLKBUF_X4 U3264 ( .I(\SB1_2_19/buf_output[0] ), .Z(\SB2_2_14/i0[9] ) );
  NAND2_X1 U6012 ( .A1(\SB1_2_4/Component_Function_4/NAND4_in[2] ), .A2(n3219), 
        .ZN(n1557) );
  CLKBUF_X4 \SB2_2_3/BUF_2  ( .I(\SB1_2_6/buf_output[2] ), .Z(\SB2_2_3/i0_0 )
         );
  CLKBUF_X4 U2551 ( .I(\SB1_2_26/buf_output[4] ), .Z(\SB2_2_25/i0_4 ) );
  CLKBUF_X4 U1875 ( .I(\SB1_2_6/buf_output[3] ), .Z(\SB2_2_4/i0[10] ) );
  CLKBUF_X4 \SB2_2_27/BUF_2  ( .I(\SB1_2_30/buf_output[2] ), .Z(
        \SB2_2_27/i0_0 ) );
  CLKBUF_X4 \SB2_2_1/BUF_0  ( .I(\SB1_2_6/buf_output[0] ), .Z(\SB2_2_1/i0[9] )
         );
  CLKBUF_X4 \SB2_2_28/BUF_1  ( .I(\SB1_2_0/buf_output[1] ), .Z(
        \SB2_2_28/i0[6] ) );
  CLKBUF_X4 \SB2_2_1/BUF_2  ( .I(\SB1_2_4/buf_output[2] ), .Z(\SB2_2_1/i0_0 )
         );
  CLKBUF_X4 U1872 ( .I(\SB1_2_31/buf_output[3] ), .Z(\SB2_2_29/i0[10] ) );
  CLKBUF_X4 \SB2_2_1/BUF_1  ( .I(\SB1_2_5/buf_output[1] ), .Z(\SB2_2_1/i0[6] )
         );
  CLKBUF_X4 U1870 ( .I(\SB2_2_30/i0_4 ), .Z(n2343) );
  CLKBUF_X4 \SB2_2_7/BUF_3  ( .I(\SB1_2_9/buf_output[3] ), .Z(\SB2_2_7/i0[10] ) );
  CLKBUF_X4 \SB2_2_17/BUF_0  ( .I(\SB1_2_22/buf_output[0] ), .Z(
        \SB2_2_17/i0[9] ) );
  CLKBUF_X4 \SB2_2_20/BUF_0  ( .I(\SB1_2_25/buf_output[0] ), .Z(
        \SB2_2_20/i0[9] ) );
  CLKBUF_X4 \SB2_2_15/BUF_5  ( .I(\SB1_2_15/buf_output[5] ), .Z(
        \SB2_2_15/i0_3 ) );
  CLKBUF_X4 \SB2_2_15/BUF_3  ( .I(\SB1_2_17/buf_output[3] ), .Z(
        \SB2_2_15/i0[10] ) );
  CLKBUF_X4 \SB2_2_24/BUF_0  ( .I(\SB1_2_29/buf_output[0] ), .Z(
        \SB2_2_24/i0[9] ) );
  CLKBUF_X4 \SB2_2_25/BUF_3  ( .I(\SB1_2_27/buf_output[3] ), .Z(
        \SB2_2_25/i0[10] ) );
  CLKBUF_X4 \SB2_2_9/BUF_3  ( .I(\SB1_2_11/buf_output[3] ), .Z(
        \SB2_2_9/i0[10] ) );
  CLKBUF_X4 \SB2_2_9/BUF_1  ( .I(\SB1_2_13/buf_output[1] ), .Z(\SB2_2_9/i0[6] ) );
  CLKBUF_X4 U3601 ( .I(\SB1_2_4/buf_output[1] ), .Z(\SB2_2_0/i0[6] ) );
  CLKBUF_X4 U4677 ( .I(\SB1_2_25/buf_output[3] ), .Z(\SB2_2_23/i0[10] ) );
  CLKBUF_X4 U3063 ( .I(\SB1_2_4/buf_output[5] ), .Z(\SB2_2_4/i0_3 ) );
  CLKBUF_X4 U1878 ( .I(\SB1_2_7/buf_output[2] ), .Z(\SB2_2_4/i0_0 ) );
  CLKBUF_X4 \SB2_2_13/BUF_3  ( .I(\SB1_2_15/buf_output[3] ), .Z(
        \SB2_2_13/i0[10] ) );
  CLKBUF_X4 \SB2_2_10/BUF_0  ( .I(\SB1_2_15/buf_output[0] ), .Z(
        \SB2_2_10/i0[9] ) );
  CLKBUF_X4 \SB2_2_21/BUF_3  ( .I(\SB1_2_23/buf_output[3] ), .Z(
        \SB2_2_21/i0[10] ) );
  CLKBUF_X4 U1083 ( .I(\SB1_2_16/buf_output[1] ), .Z(\SB2_2_12/i0[6] ) );
  CLKBUF_X4 \SB2_2_21/BUF_1  ( .I(\SB1_2_25/buf_output[1] ), .Z(
        \SB2_2_21/i0[6] ) );
  CLKBUF_X4 \SB2_2_7/BUF_0  ( .I(\SB1_2_12/buf_output[0] ), .Z(\SB2_2_7/i0[9] ) );
  CLKBUF_X4 U2087 ( .I(\SB1_2_20/buf_output[4] ), .Z(\SB2_2_19/i0_4 ) );
  CLKBUF_X4 \SB2_2_19/BUF_2  ( .I(\SB1_2_22/buf_output[2] ), .Z(
        \SB2_2_19/i0_0 ) );
  CLKBUF_X4 \SB2_2_31/BUF_0  ( .I(\SB1_2_4/buf_output[0] ), .Z(
        \SB2_2_31/i0[9] ) );
  CLKBUF_X4 \SB2_2_5/BUF_1  ( .I(\SB1_2_9/buf_output[1] ), .Z(\SB2_2_5/i0[6] )
         );
  CLKBUF_X4 U4146 ( .I(\SB1_2_22/buf_output[1] ), .Z(\SB2_2_18/i0[6] ) );
  CLKBUF_X4 \SB2_2_23/BUF_1  ( .I(\SB1_2_27/buf_output[1] ), .Z(
        \SB2_2_23/i0[6] ) );
  CLKBUF_X4 \SB2_2_26/BUF_2  ( .I(\SB1_2_29/buf_output[2] ), .Z(
        \SB2_2_26/i0_0 ) );
  CLKBUF_X4 \SB2_2_21/BUF_2  ( .I(\SB1_2_24/buf_output[2] ), .Z(
        \SB2_2_21/i0_0 ) );
  CLKBUF_X4 U3269 ( .I(\SB1_2_29/buf_output[3] ), .Z(\SB2_2_27/i0[10] ) );
  CLKBUF_X4 U4109 ( .I(\SB2_2_18/buf_output[1] ), .Z(\RI5[2][103] ) );
  CLKBUF_X4 \MC_ARK_ARC_1_2/BUF_133  ( .I(\SB2_2_13/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[133] ) );
  CLKBUF_X4 \SB2_2_26/BUF_4_0  ( .I(\SB2_2_26/buf_output[4] ), .Z(\RI5[2][40] ) );
  CLKBUF_X4 U3138 ( .I(\SB2_2_13/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[128] ) );
  CLKBUF_X4 U3255 ( .I(\SB2_2_26/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[50] ) );
  CLKBUF_X4 \MC_ARK_ARC_1_2/BUF_136  ( .I(\SB2_2_10/buf_output[4] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[136] ) );
  CLKBUF_X4 U6918 ( .I(\SB2_2_15/buf_output[0] ), .Z(\RI5[2][126] ) );
  CLKBUF_X4 U7995 ( .I(\SB2_2_4/buf_output[5] ), .Z(\RI5[2][167] ) );
  CLKBUF_X4 U8196 ( .I(\SB2_2_28/buf_output[3] ), .Z(\RI5[2][33] ) );
  CLKBUF_X4 U2472 ( .I(\MC_ARK_ARC_1_2/buf_output[81] ), .Z(\SB1_3_18/i0[10] )
         );
  CLKBUF_X4 \SB1_3_6/BUF_1  ( .I(\MC_ARK_ARC_1_2/buf_output[151] ), .Z(
        \SB1_3_6/i0[6] ) );
  CLKBUF_X4 U8709 ( .I(\MC_ARK_ARC_1_2/buf_output[130] ), .Z(\SB1_3_10/i0_4 )
         );
  CLKBUF_X4 \SB1_3_2/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[178] ), .Z(
        \SB1_3_2/i0_4 ) );
  CLKBUF_X4 U2995 ( .I(\MC_ARK_ARC_1_2/buf_output[88] ), .Z(\SB1_3_17/i0_4 )
         );
  CLKBUF_X4 U2110 ( .I(\MC_ARK_ARC_1_2/buf_output[105] ), .Z(\SB1_3_14/i0[10] ) );
  CLKBUF_X4 \SB1_3_31/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[4] ), .Z(
        \SB1_3_31/i0_4 ) );
  CLKBUF_X4 \SB1_3_20/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[70] ), .Z(
        \SB1_3_20/i0_4 ) );
  CLKBUF_X4 U4396 ( .I(\MC_ARK_ARC_1_2/buf_output[1] ), .Z(\SB1_3_31/i0[6] )
         );
  CLKBUF_X4 U4494 ( .I(\MC_ARK_ARC_1_2/buf_output[103] ), .Z(\SB1_3_14/i0[6] )
         );
  CLKBUF_X4 \SB1_3_9/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[136] ), .Z(
        \SB1_3_9/i0_4 ) );
  CLKBUF_X4 \SB1_3_7/BUF_0  ( .I(\MC_ARK_ARC_1_2/buf_output[144] ), .Z(
        \SB1_3_7/i0[9] ) );
  CLKBUF_X4 U4968 ( .I(\MC_ARK_ARC_1_2/buf_output[158] ), .Z(\SB1_3_5/i0_0 )
         );
  CLKBUF_X4 \SB1_3_5/BUF_0  ( .I(\MC_ARK_ARC_1_2/buf_output[156] ), .Z(
        \SB1_3_5/i0[9] ) );
  CLKBUF_X4 U4431 ( .I(\MC_ARK_ARC_1_2/buf_output[160] ), .Z(\SB1_3_5/i0_4 )
         );
  CLKBUF_X4 \SB1_3_16/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[94] ), .Z(
        \SB1_3_16/i0_4 ) );
  CLKBUF_X4 U4397 ( .I(\MC_ARK_ARC_1_2/buf_output[124] ), .Z(\SB1_3_11/i0_4 )
         );
  CLKBUF_X4 U917 ( .I(\MC_ARK_ARC_1_2/buf_output[148] ), .Z(\SB1_3_7/i0_4 ) );
  CLKBUF_X4 \SB1_3_4/BUF_4  ( .I(\MC_ARK_ARC_1_2/buf_output[166] ), .Z(
        \SB1_3_4/i0_4 ) );
  CLKBUF_X4 \SB1_3_16/BUF_1  ( .I(\MC_ARK_ARC_1_2/buf_output[91] ), .Z(
        \SB1_3_16/i0[6] ) );
  CLKBUF_X4 U9013 ( .I(\MC_ARK_ARC_1_2/buf_output[152] ), .Z(\SB1_3_6/i0_0 )
         );
  CLKBUF_X4 \SB1_3_26/BUF_0  ( .I(\MC_ARK_ARC_1_2/buf_output[30] ), .Z(
        \SB1_3_26/i0[9] ) );
  NAND2_X2 \SB1_3_6/Component_Function_5/N1  ( .A1(\SB1_3_6/i0_0 ), .A2(
        \SB1_3_6/i3[0] ), .ZN(\SB1_3_6/Component_Function_5/NAND4_in[0] ) );
  CLKBUF_X4 U8866 ( .I(\MC_ARK_ARC_1_2/buf_output[159] ), .Z(\SB1_3_5/i0[10] )
         );
  CLKBUF_X4 U8562 ( .I(\MC_ARK_ARC_1_2/buf_output[29] ), .Z(\SB1_3_27/i0_3 )
         );
  CLKBUF_X4 U3637 ( .I(\MC_ARK_ARC_1_2/buf_output[169] ), .Z(\SB1_3_3/i0[6] )
         );
  CLKBUF_X4 U3646 ( .I(\MC_ARK_ARC_1_2/buf_output[168] ), .Z(\SB1_3_3/i0[9] )
         );
  CLKBUF_X4 U2908 ( .I(\MC_ARK_ARC_1_2/buf_output[189] ), .Z(\SB1_3_0/i0[10] )
         );
  CLKBUF_X4 U3252 ( .I(\MC_ARK_ARC_1_2/buf_output[174] ), .Z(\SB1_3_2/i0[9] )
         );
  CLKBUF_X4 U3247 ( .I(\MC_ARK_ARC_1_2/buf_output[164] ), .Z(\SB1_3_4/i0_0 )
         );
  CLKBUF_X4 \SB1_3_9/BUF_0  ( .I(\MC_ARK_ARC_1_2/buf_output[132] ), .Z(
        \SB1_3_9/i0[9] ) );
  NAND3_X2 \SB1_3_2/Component_Function_2/N4  ( .A1(\SB1_3_2/i1_5 ), .A2(
        \SB1_3_2/i0_0 ), .A3(\SB1_3_2/i0_4 ), .ZN(
        \SB1_3_2/Component_Function_2/NAND4_in[3] ) );
  BUF_X4 U4524 ( .I(\SB1_3_2/buf_output[3] ), .Z(\SB2_3_0/i0[10] ) );
  CLKBUF_X4 \SB2_3_16/BUF_2  ( .I(\SB1_3_19/buf_output[2] ), .Z(
        \SB2_3_16/i0_0 ) );
  CLKBUF_X4 U8487 ( .I(\SB1_3_3/buf_output[2] ), .Z(\SB2_3_0/i0_0 ) );
  CLKBUF_X4 \SB2_3_16/BUF_3  ( .I(\SB1_3_18/buf_output[3] ), .Z(
        \SB2_3_16/i0[10] ) );
  CLKBUF_X4 U1443 ( .I(\SB1_3_20/buf_output[2] ), .Z(\SB2_3_17/i0_0 ) );
  CLKBUF_X4 \SB2_3_29/BUF_1  ( .I(\SB1_3_1/buf_output[1] ), .Z(
        \SB2_3_29/i0[6] ) );
  CLKBUF_X2 U733 ( .I(\SB1_3_19/buf_output[0] ), .Z(\SB2_3_14/i0[9] ) );
  CLKBUF_X4 U732 ( .I(\SB1_3_12/buf_output[1] ), .Z(\SB2_3_8/i0[6] ) );
  CLKBUF_X4 U9024 ( .I(\SB1_3_8/buf_output[3] ), .Z(\SB2_3_6/i0[10] ) );
  CLKBUF_X4 \SB2_3_29/BUF_3  ( .I(\SB1_3_31/buf_output[3] ), .Z(
        \SB2_3_29/i0[10] ) );
  CLKBUF_X4 U4546 ( .I(\SB1_3_19/buf_output[3] ), .Z(\SB2_3_17/i0[10] ) );
  CLKBUF_X4 \SB2_3_13/BUF_1  ( .I(\SB1_3_17/buf_output[1] ), .Z(
        \SB2_3_13/i0[6] ) );
  CLKBUF_X4 U726 ( .I(\SB1_3_4/buf_output[1] ), .Z(\SB2_3_0/i0[6] ) );
  CLKBUF_X4 \SB2_3_22/BUF_1  ( .I(\SB1_3_26/buf_output[1] ), .Z(
        \SB2_3_22/i0[6] ) );
  CLKBUF_X4 U3237 ( .I(\SB1_3_29/buf_output[3] ), .Z(\SB2_3_27/i0[10] ) );
  CLKBUF_X4 \SB2_3_0/BUF_0  ( .I(\SB1_3_5/buf_output[0] ), .Z(\SB2_3_0/i0[9] )
         );
  CLKBUF_X4 \SB2_3_6/BUF_1  ( .I(\SB1_3_10/buf_output[1] ), .Z(\SB2_3_6/i0[6] ) );
  CLKBUF_X4 \SB2_3_28/BUF_1  ( .I(\SB1_3_0/buf_output[1] ), .Z(
        \SB2_3_28/i0[6] ) );
  CLKBUF_X4 \SB2_3_28/BUF_0  ( .I(\SB1_3_1/buf_output[0] ), .Z(
        \SB2_3_28/i0[9] ) );
  CLKBUF_X4 U4560 ( .I(\SB1_3_16/buf_output[2] ), .Z(\SB2_3_13/i0_0 ) );
  CLKBUF_X4 U2836 ( .I(\SB1_3_5/buf_output[4] ), .Z(\SB2_3_4/i0_4 ) );
  CLKBUF_X4 U8721 ( .I(\RI3[3][35] ), .Z(\SB2_3_26/i0_3 ) );
  CLKBUF_X4 \SB2_3_18/BUF_3  ( .I(\SB1_3_20/buf_output[3] ), .Z(
        \SB2_3_18/i0[10] ) );
  CLKBUF_X4 U2487 ( .I(\SB1_3_14/buf_output[5] ), .Z(\SB2_3_14/i0_3 ) );
  CLKBUF_X4 \SB2_3_10/BUF_1  ( .I(\SB1_3_14/buf_output[1] ), .Z(
        \SB2_3_10/i0[6] ) );
  CLKBUF_X4 U2033 ( .I(\SB1_3_26/buf_output[2] ), .Z(\SB2_3_23/i0_0 ) );
  CLKBUF_X4 \SB2_3_10/BUF_2  ( .I(\SB1_3_13/buf_output[2] ), .Z(
        \SB2_3_10/i0_0 ) );
  CLKBUF_X4 \SB2_3_23/BUF_1  ( .I(\SB1_3_27/buf_output[1] ), .Z(
        \SB2_3_23/i0[6] ) );
  CLKBUF_X4 \SB2_3_18/BUF_4  ( .I(\SB1_3_19/buf_output[4] ), .Z(
        \SB2_3_18/i0_4 ) );
  CLKBUF_X4 \SB2_3_25/BUF_5  ( .I(\SB1_3_25/buf_output[5] ), .Z(
        \SB2_3_25/i0_3 ) );
  CLKBUF_X4 U4602 ( .I(\SB1_3_7/buf_output[2] ), .Z(\SB2_3_4/i0_0 ) );
  CLKBUF_X4 U2446 ( .I(\SB1_3_19/buf_output[5] ), .Z(\SB2_3_19/i0_3 ) );
  CLKBUF_X4 U7958 ( .I(\SB1_3_0/buf_output[3] ), .Z(\SB2_3_30/i0[10] ) );
  CLKBUF_X4 \SB2_3_10/BUF_0  ( .I(\SB1_3_15/buf_output[0] ), .Z(
        \SB2_3_10/i0[9] ) );
  CLKBUF_X4 \SB2_3_18/BUF_1  ( .I(\SB1_3_22/buf_output[1] ), .Z(
        \SB2_3_18/i0[6] ) );
  CLKBUF_X4 U3699 ( .I(\SB1_3_23/buf_output[1] ), .Z(\SB2_3_19/i0[6] ) );
  CLKBUF_X4 \SB2_3_5/BUF_1  ( .I(\SB1_3_9/buf_output[1] ), .Z(\SB2_3_5/i0[6] )
         );
  CLKBUF_X4 U5202 ( .I(\SB1_3_14/buf_output[3] ), .Z(\SB2_3_12/i0[10] ) );
  CLKBUF_X4 U2296 ( .I(\SB1_3_8/buf_output[0] ), .Z(\SB2_3_3/i0[9] ) );
  CLKBUF_X4 U1831 ( .I(\SB1_3_4/buf_output[4] ), .Z(\SB2_3_3/i0_4 ) );
  CLKBUF_X4 \SB2_3_30/BUF_2  ( .I(\SB1_3_1/buf_output[2] ), .Z(\SB2_3_30/i0_0 ) );
  CLKBUF_X4 \SB2_3_5/BUF_0  ( .I(\SB1_3_10/buf_output[0] ), .Z(\SB2_3_5/i0[9] ) );
  CLKBUF_X4 \SB2_3_13/BUF_0  ( .I(\SB1_3_18/buf_output[0] ), .Z(
        \SB2_3_13/i0[9] ) );
  CLKBUF_X4 U4647 ( .I(\SB1_3_20/buf_output[5] ), .Z(\SB2_3_20/i0_3 ) );
  CLKBUF_X4 U759 ( .I(\SB1_3_13/buf_output[0] ), .Z(\SB2_3_8/i0[9] ) );
  CLKBUF_X4 \SB2_3_31/BUF_2  ( .I(\SB1_3_2/buf_output[2] ), .Z(\SB2_3_31/i0_0 ) );
  CLKBUF_X4 \SB2_3_2/BUF_2  ( .I(\SB1_3_5/buf_output[2] ), .Z(\SB2_3_2/i0_0 )
         );
  CLKBUF_X4 \SB2_3_11/BUF_1  ( .I(\SB1_3_15/buf_output[1] ), .Z(
        \SB2_3_11/i0[6] ) );
  CLKBUF_X4 U8667 ( .I(\SB1_3_0/buf_output[4] ), .Z(\SB2_3_31/i0_4 ) );
  NAND2_X1 U2692 ( .A1(\SB2_3_19/i0_0 ), .A2(\SB2_3_19/i3[0] ), .ZN(
        \SB2_3_19/Component_Function_5/NAND4_in[0] ) );
  CLKBUF_X4 U8846 ( .I(\SB2_3_4/buf_output[3] ), .Z(\RI5[3][177] ) );
  CLKBUF_X4 U4738 ( .I(\SB2_3_16/buf_output[3] ), .Z(\RI5[3][105] ) );
  CLKBUF_X4 U8838 ( .I(\SB2_3_19/buf_output[5] ), .Z(\RI5[3][77] ) );
  CLKBUF_X4 U4591 ( .I(\SB2_3_19/buf_output[3] ), .Z(\RI5[3][87] ) );
  BUF_X2 U3728 ( .I(\SB2_3_13/buf_output[3] ), .Z(n3658) );
  CLKBUF_X4 U3730 ( .I(\SB2_3_8/buf_output[5] ), .Z(\RI5[3][143] ) );
  CLKBUF_X4 U5728 ( .I(\SB2_3_20/buf_output[0] ), .Z(\RI5[3][96] ) );
  CLKBUF_X4 U1324 ( .I(\MC_ARK_ARC_1_3/buf_output[135] ), .Z(\SB3_9/i0[10] )
         );
  CLKBUF_X4 U1442 ( .I(\MC_ARK_ARC_1_3/buf_output[182] ), .Z(\SB3_1/i0_0 ) );
  CLKBUF_X4 U2552 ( .I(\MC_ARK_ARC_1_3/buf_output[158] ), .Z(\SB3_5/i0_0 ) );
  BUF_X2 U2148 ( .I(\MC_ARK_ARC_1_3/buf_output[133] ), .Z(\SB3_9/i0[6] ) );
  CLKBUF_X4 U1277 ( .I(\MC_ARK_ARC_1_3/buf_output[24] ), .Z(\SB3_27/i0[9] ) );
  CLKBUF_X4 U2190 ( .I(\MC_ARK_ARC_1_3/buf_output[58] ), .Z(\SB3_22/i0_4 ) );
  CLKBUF_X4 \SB3_31/BUF_1  ( .I(\MC_ARK_ARC_1_3/buf_output[1] ), .Z(
        \SB3_31/i0[6] ) );
  CLKBUF_X4 \SB3_15/BUF_2  ( .I(\MC_ARK_ARC_1_3/buf_output[98] ), .Z(
        \SB3_15/i0_0 ) );
  CLKBUF_X4 U657 ( .I(\MC_ARK_ARC_1_3/buf_output[40] ), .Z(\SB3_25/i0_4 ) );
  CLKBUF_X4 U2842 ( .I(\RI1[4][77] ), .Z(\SB3_19/i0_3 ) );
  CLKBUF_X4 U4669 ( .I(\MC_ARK_ARC_1_3/buf_output[15] ), .Z(\SB3_29/i0[10] )
         );
  CLKBUF_X4 \SB3_18/BUF_4  ( .I(\MC_ARK_ARC_1_3/buf_output[82] ), .Z(
        \SB3_18/i0_4 ) );
  CLKBUF_X4 U4545 ( .I(\MC_ARK_ARC_1_3/buf_output[60] ), .Z(\SB3_21/i0[9] ) );
  CLKBUF_X4 U2985 ( .I(\MC_ARK_ARC_1_3/buf_output[65] ), .Z(\RI1[4][65] ) );
  CLKBUF_X4 \SB3_2/BUF_4  ( .I(\MC_ARK_ARC_1_3/buf_output[178] ), .Z(
        \SB3_2/i0_4 ) );
  CLKBUF_X4 U1809 ( .I(n1401), .Z(\SB3_23/i0_0 ) );
  CLKBUF_X4 U1807 ( .I(\MC_ARK_ARC_1_3/buf_output[14] ), .Z(\SB3_29/i0_0 ) );
  CLKBUF_X4 \SB3_14/BUF_0  ( .I(\MC_ARK_ARC_1_3/buf_output[102] ), .Z(
        \SB3_14/i0[9] ) );
  CLKBUF_X4 U8809 ( .I(\SB3_31/buf_output[4] ), .Z(\SB4_30/i0_4 ) );
  CLKBUF_X4 U4537 ( .I(\SB3_28/buf_output[3] ), .Z(\SB4_26/i0[10] ) );
  CLKBUF_X4 U4920 ( .I(\SB3_25/buf_output[2] ), .Z(\SB4_22/i0_0 ) );
  BUF_X2 \SB4_23/BUF_0  ( .I(\SB3_28/buf_output[0] ), .Z(\SB4_23/i0[9] ) );
  CLKBUF_X4 U7385 ( .I(\SB3_19/buf_output[4] ), .Z(\SB4_18/i0_4 ) );
  CLKBUF_X4 U2158 ( .I(\SB3_8/buf_output[2] ), .Z(\SB4_5/i0_0 ) );
  CLKBUF_X4 U2417 ( .I(\SB3_22/buf_output[1] ), .Z(\SB4_18/i0[6] ) );
  CLKBUF_X4 U583 ( .I(\SB3_22/buf_output[0] ), .Z(\SB4_17/i0[9] ) );
  CLKBUF_X4 \SB4_4/BUF_0  ( .I(\SB3_9/buf_output[0] ), .Z(\SB4_4/i0[9] ) );
  CLKBUF_X4 U581 ( .I(\SB3_2/buf_output[4] ), .Z(\SB4_1/i0_4 ) );
  CLKBUF_X4 U1792 ( .I(\SB3_23/buf_output[5] ), .Z(\SB4_23/i0_3 ) );
  CLKBUF_X4 U4168 ( .I(\SB3_1/buf_output[1] ), .Z(\SB4_29/i0[6] ) );
  CLKBUF_X4 \SB4_24/BUF_0  ( .I(\SB3_29/buf_output[0] ), .Z(\SB4_24/i0[9] ) );
  BUF_X2 \SB4_15/BUF_3  ( .I(\SB3_17/buf_output[3] ), .Z(\SB4_15/i0[10] ) );
  CLKBUF_X4 U3189 ( .I(\SB3_6/buf_output[0] ), .Z(\SB4_1/i0[9] ) );
  BUF_X4 U1260 ( .I(\MC_ARK_ARC_1_3/buf_output[68] ), .Z(\SB3_20/i0_0 ) );
  BUF_X4 U8040 ( .I(\SB2_0_30/buf_output[4] ), .Z(\RI5[0][16] ) );
  NAND3_X2 \SB1_0_22/Component_Function_4/N2  ( .A1(\SB1_0_22/i3[0] ), .A2(
        \SB1_0_22/i0_0 ), .A3(\SB1_0_22/i1_7 ), .ZN(
        \SB1_0_22/Component_Function_4/NAND4_in[1] ) );
  AND2_X1 U1651 ( .A1(\MC_ARK_ARC_1_0/buf_output[51] ), .A2(
        \MC_ARK_ARC_1_0/buf_output[50] ), .Z(n2224) );
  NAND2_X2 U3610 ( .A1(\SB1_0_11/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_0_11/Component_Function_4/NAND4_in[0] ), .ZN(n1053) );
  BUF_X4 U4584 ( .I(\MC_ARK_ARC_1_1/buf_output[81] ), .Z(\SB1_2_18/i0[10] ) );
  INV_X2 U1261 ( .I(\MC_ARK_ARC_1_3/buf_output[68] ), .ZN(\SB3_20/i1[9] ) );
  NAND3_X2 \SB2_0_29/Component_Function_3/N2  ( .A1(\SB2_0_29/i0_0 ), .A2(
        \SB2_0_29/i0_3 ), .A3(\SB2_0_29/i0_4 ), .ZN(
        \SB2_0_29/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U8830 ( .A1(\SB2_3_22/i1_5 ), .A2(\SB2_3_22/i0[8] ), .A3(
        \SB2_3_22/i3[0] ), .ZN(\SB2_3_22/Component_Function_3/NAND4_in[3] ) );
  BUF_X2 \SB1_0_17/BUF_0  ( .I(n287), .Z(\SB1_0_17/i0[9] ) );
  BUF_X2 \SB1_0_10/BUF_4  ( .I(n384), .Z(\SB1_0_10/i0_4 ) );
  BUF_X2 \SB1_0_12/BUF_1  ( .I(n303), .Z(\SB1_0_12/i0[6] ) );
  INV_X1 \SB1_0_16/INV_4  ( .I(n4752), .ZN(\SB1_0_16/i0[7] ) );
  INV_X1 \SB1_0_10/INV_2  ( .I(n310), .ZN(\SB1_0_10/i1[9] ) );
  NAND3_X1 \SB1_0_3/Component_Function_4/N3  ( .A1(\SB1_0_3/i0[9] ), .A2(
        \SB1_0_3/i0[10] ), .A3(\SB1_0_3/i0_3 ), .ZN(
        \SB1_0_3/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U11038 ( .A1(\SB1_0_4/i1_5 ), .A2(\SB1_0_4/i3[0] ), .A3(
        \SB1_0_4/i0[8] ), .ZN(\SB1_0_4/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U10280 ( .A1(\SB1_0_27/i0[10] ), .A2(\SB1_0_27/i1[9] ), .A3(
        \SB1_0_27/i1_7 ), .ZN(n4244) );
  NAND3_X1 U1136 ( .A1(\SB1_0_4/i0_3 ), .A2(\SB1_0_4/i0[6] ), .A3(
        \SB1_0_4/i1[9] ), .ZN(n1667) );
  BUF_X2 \SB1_0_23/BUF_0  ( .I(n269), .Z(\SB1_0_23/i0[9] ) );
  CLKBUF_X2 \SB1_0_29/BUF_1  ( .I(n252), .Z(\SB1_0_29/i0[6] ) );
  BUF_X2 \SB1_0_21/BUF_4  ( .I(n362), .Z(\SB1_0_21/i0_4 ) );
  INV_X1 \SB1_0_8/INV_3  ( .I(n387), .ZN(\SB1_0_8/i0[8] ) );
  INV_X1 U1462 ( .I(n401), .ZN(\SB1_0_1/i0[8] ) );
  NAND3_X1 U4721 ( .A1(\SB1_0_7/i0_3 ), .A2(\SB1_0_7/i0[10] ), .A3(n390), .ZN(
        n1549) );
  NAND3_X1 U6962 ( .A1(\SB1_0_15/i0[10] ), .A2(\SB1_0_15/i1[9] ), .A3(
        \SB1_0_15/i1_7 ), .ZN(n2330) );
  NAND3_X1 \SB1_0_2/Component_Function_2/N3  ( .A1(\SB1_0_2/i0_3 ), .A2(
        \SB1_0_2/i0[8] ), .A3(\SB1_0_2/i0[9] ), .ZN(
        \SB1_0_2/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1944 ( .A1(\SB1_0_5/i0[10] ), .A2(\SB1_0_5/i0_3 ), .A3(
        \SB1_0_5/i0[9] ), .ZN(n2478) );
  NAND3_X1 U1698 ( .A1(\SB1_0_25/i0_3 ), .A2(\SB1_0_25/i0[10] ), .A3(
        \SB1_0_25/i0[9] ), .ZN(\SB1_0_25/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U9313 ( .A1(\SB1_0_1/i0_3 ), .A2(\SB1_0_1/i0[6] ), .A3(
        \SB1_0_1/i1[9] ), .ZN(\SB1_0_1/Component_Function_3/NAND4_in[0] ) );
  NAND2_X1 U5574 ( .A1(\SB1_0_17/Component_Function_4/NAND4_in[1] ), .A2(n2036), .ZN(n2035) );
  NAND2_X1 \SB1_0_29/Component_Function_5/N1  ( .A1(\SB1_0_29/i0_0 ), .A2(
        \SB1_0_29/i3[0] ), .ZN(\SB1_0_29/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U1126 ( .A1(\SB1_0_23/i0_3 ), .A2(\SB1_0_23/i0_4 ), .A3(
        \SB1_0_23/i1[9] ), .ZN(\SB1_0_23/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_3/Component_Function_1/N2  ( .A1(\SB1_0_3/i0_3 ), .A2(
        \SB1_0_3/i1_7 ), .A3(\SB1_0_3/i0[8] ), .ZN(
        \SB1_0_3/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U7708 ( .A1(\SB1_0_8/i0_0 ), .A2(\SB1_0_8/i1_5 ), .A3(
        \SB1_0_8/i0_4 ), .ZN(n2750) );
  NAND3_X1 \SB1_0_3/Component_Function_1/N4  ( .A1(\SB1_0_3/i1_7 ), .A2(
        \SB1_0_3/i0[8] ), .A3(\SB1_0_3/i0_4 ), .ZN(
        \SB1_0_3/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U3742 ( .A1(\SB1_0_14/i0_3 ), .A2(\SB1_0_14/i0[9] ), .A3(
        \SB1_0_14/i0[8] ), .ZN(n1105) );
  NAND3_X1 \SB1_0_1/Component_Function_3/N2  ( .A1(\SB1_0_1/i0_0 ), .A2(
        \SB1_0_1/i0_3 ), .A3(\SB1_0_1/i0_4 ), .ZN(
        \SB1_0_1/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U10279 ( .A1(\SB1_0_5/i0_0 ), .A2(\SB1_0_5/i0[9] ), .A3(
        \SB1_0_5/i0[8] ), .ZN(\SB1_0_5/Component_Function_4/NAND4_in[0] ) );
  NAND2_X1 \SB1_0_6/Component_Function_1/N1  ( .A1(\SB1_0_6/i0_3 ), .A2(
        \SB1_0_6/i1[9] ), .ZN(\SB1_0_6/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U1131 ( .A1(\SB1_0_25/i0_4 ), .A2(\SB1_0_25/i1[9] ), .A3(
        \SB1_0_25/i1_5 ), .ZN(n2554) );
  NAND2_X1 U3345 ( .A1(\SB1_0_28/i0_3 ), .A2(\SB1_0_28/i1[9] ), .ZN(
        \SB1_0_28/Component_Function_1/NAND4_in[0] ) );
  INV_X2 \SB1_0_1/INV_4  ( .I(\SB1_0_1/i0_4 ), .ZN(\SB1_0_1/i0[7] ) );
  NAND3_X1 \SB1_0_16/Component_Function_3/N1  ( .A1(\SB1_0_16/i1[9] ), .A2(
        \SB1_0_16/i0_3 ), .A3(\SB1_0_16/i0[6] ), .ZN(
        \SB1_0_16/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U9454 ( .A1(\SB1_0_16/i0_3 ), .A2(\SB1_0_16/i0_0 ), .A3(n4752), 
        .ZN(\SB1_0_16/Component_Function_3/NAND4_in[1] ) );
  INV_X1 \SB1_0_25/INV_4  ( .I(\SB1_0_25/i0_4 ), .ZN(\SB1_0_25/i0[7] ) );
  NAND3_X1 \SB1_0_8/Component_Function_2/N1  ( .A1(\SB1_0_8/i1_5 ), .A2(
        \SB1_0_8/i0[10] ), .A3(\SB1_0_8/i1[9] ), .ZN(
        \SB1_0_8/Component_Function_2/NAND4_in[0] ) );
  NAND2_X1 \SB1_0_9/Component_Function_5/N1  ( .A1(\SB1_0_9/i0_0 ), .A2(
        \SB1_0_9/i3[0] ), .ZN(\SB1_0_9/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB1_0_15/Component_Function_1/N1  ( .A1(\SB1_0_15/i0_3 ), .A2(
        \SB1_0_15/i1[9] ), .ZN(\SB1_0_15/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_25/Component_Function_3/N3  ( .A1(\SB1_0_25/i1[9] ), .A2(
        \SB1_0_25/i1_7 ), .A3(\SB1_0_25/i0[10] ), .ZN(
        \SB1_0_25/Component_Function_3/NAND4_in[2] ) );
  INV_X1 U1935 ( .I(\SB1_0_20/i0_4 ), .ZN(\SB1_0_20/i0[7] ) );
  NAND3_X1 \SB1_0_9/Component_Function_2/N3  ( .A1(\SB1_0_9/i0_3 ), .A2(
        \SB1_0_9/i0[8] ), .A3(\SB1_0_9/i0[9] ), .ZN(
        \SB1_0_9/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U4672 ( .A1(\SB1_0_19/i0_0 ), .A2(\SB1_0_19/i0[7] ), .A3(
        \SB1_0_19/i0_3 ), .ZN(n2201) );
  NAND3_X1 U10318 ( .A1(\SB1_0_13/i0_0 ), .A2(\SB1_0_13/i1_5 ), .A3(
        \SB1_0_13/i0_4 ), .ZN(n4260) );
  NAND2_X1 \SB1_0_26/Component_Function_5/N1  ( .A1(\SB1_0_26/i0_0 ), .A2(
        \SB1_0_26/i3[0] ), .ZN(\SB1_0_26/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U1642 ( .A1(\SB1_0_12/i0[10] ), .A2(\SB1_0_12/i0_3 ), .A3(
        \SB1_0_12/i0_4 ), .ZN(n3155) );
  NAND3_X1 U4661 ( .A1(\SB1_0_6/i0[10] ), .A2(\SB1_0_6/i0_4 ), .A3(
        \SB1_0_6/i0_3 ), .ZN(\SB1_0_6/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U1112 ( .A1(\SB1_0_15/i0[10] ), .A2(\SB1_0_15/i0_3 ), .A3(
        \SB1_0_15/i0[9] ), .ZN(n1121) );
  NAND3_X1 \SB1_0_21/Component_Function_2/N1  ( .A1(\SB1_0_21/i1_5 ), .A2(
        \SB1_0_21/i0[10] ), .A3(\SB1_0_21/i1[9] ), .ZN(
        \SB1_0_21/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_8/Component_Function_3/N3  ( .A1(\SB1_0_8/i1[9] ), .A2(
        \SB1_0_8/i1_7 ), .A3(\SB1_0_8/i0[10] ), .ZN(
        \SB1_0_8/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_7/Component_Function_1/N2  ( .A1(\SB1_0_7/i0_3 ), .A2(
        \SB1_0_7/i1_7 ), .A3(\SB1_0_7/i0[8] ), .ZN(
        \SB1_0_7/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_0_3/Component_Function_2/N3  ( .A1(\SB1_0_3/i0_3 ), .A2(
        \SB1_0_3/i0[8] ), .A3(\SB1_0_3/i0[9] ), .ZN(
        \SB1_0_3/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_7/Component_Function_2/N3  ( .A1(\SB1_0_7/i0_3 ), .A2(
        \SB1_0_7/i0[8] ), .A3(\SB1_0_7/i0[9] ), .ZN(
        \SB1_0_7/Component_Function_2/NAND4_in[2] ) );
  NAND2_X1 \SB1_0_10/Component_Function_5/N1  ( .A1(\SB1_0_10/i0_0 ), .A2(
        \SB1_0_10/i3[0] ), .ZN(\SB1_0_10/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_0_28/Component_Function_2/N3  ( .A1(\SB1_0_28/i0_3 ), .A2(
        \SB1_0_28/i0[8] ), .A3(\SB1_0_28/i0[9] ), .ZN(
        \SB1_0_28/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_0_1/Component_Function_5/N2  ( .A1(\SB1_0_1/i0_0 ), .A2(
        \SB1_0_1/i0[6] ), .A3(\SB1_0_1/i0[10] ), .ZN(
        \SB1_0_1/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1618 ( .A1(\SB1_0_1/i0[10] ), .A2(\SB1_0_1/i0_3 ), .A3(
        \SB1_0_1/i0[6] ), .ZN(\SB1_0_1/Component_Function_2/NAND4_in[1] ) );
  NAND2_X1 U11031 ( .A1(n1052), .A2(
        \SB1_0_11/Component_Function_4/NAND4_in[1] ), .ZN(n4675) );
  NAND3_X1 U5625 ( .A1(\SB1_0_25/i0_3 ), .A2(\SB1_0_25/i1[9] ), .A3(
        \SB1_0_25/i0_4 ), .ZN(\SB1_0_25/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1528 ( .A1(\SB1_0_3/i0_0 ), .A2(\SB1_0_3/i0[6] ), .A3(
        \SB1_0_3/i0[10] ), .ZN(\SB1_0_3/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U7405 ( .A1(\SB1_0_15/i0[10] ), .A2(\SB1_0_15/i1[9] ), .A3(
        \SB1_0_15/i1_5 ), .ZN(\SB1_0_15/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U4658 ( .A1(\SB1_0_6/i0_3 ), .A2(\SB1_0_6/i0[8] ), .A3(
        \SB1_0_6/i0[9] ), .ZN(\SB1_0_6/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1351 ( .A1(\SB1_0_6/i0_3 ), .A2(\SB1_0_6/i0_4 ), .A3(
        \SB1_0_6/i0_0 ), .ZN(n1917) );
  NAND3_X1 U9838 ( .A1(\SB1_0_9/i0_3 ), .A2(\SB1_0_9/i0[6] ), .A3(
        \SB1_0_9/i0[10] ), .ZN(n4028) );
  NAND3_X1 \SB1_0_6/Component_Function_2/N2  ( .A1(\SB1_0_6/i0_3 ), .A2(
        \SB1_0_6/i0[10] ), .A3(\SB1_0_6/i0[6] ), .ZN(
        \SB1_0_6/Component_Function_2/NAND4_in[1] ) );
  INV_X2 U5567 ( .I(n2682), .ZN(\SB2_0_16/i0_4 ) );
  BUF_X2 \SB2_0_23/BUF_0  ( .I(\RI3[0][48] ), .Z(\SB2_0_23/i0[9] ) );
  INV_X4 \SB2_0_2/INV_2  ( .I(\RI3[0][176] ), .ZN(\SB2_0_2/i1[9] ) );
  INV_X1 \SB2_0_27/INV_0  ( .I(n1091), .ZN(\SB2_0_27/i3[0] ) );
  CLKBUF_X2 \SB2_0_31/BUF_1  ( .I(\RI3[0][1] ), .Z(\SB2_0_31/i0[6] ) );
  INV_X2 U2688 ( .I(n2877), .ZN(\SB2_0_23/i0_4 ) );
  BUF_X2 \SB1_0_0/BUF_4_0  ( .I(\SB1_0_0/buf_output[4] ), .Z(\RI3[0][4] ) );
  BUF_X2 \SB2_0_2/BUF_1  ( .I(\RI3[0][175] ), .Z(\SB2_0_2/i0[6] ) );
  INV_X2 U3720 ( .I(n2237), .ZN(\SB2_0_27/i0_4 ) );
  NAND3_X1 U1611 ( .A1(\SB2_0_27/i0[10] ), .A2(\SB2_0_27/i0_0 ), .A3(
        \SB2_0_27/i0[6] ), .ZN(n2227) );
  NAND3_X1 U4312 ( .A1(\SB2_0_27/i0[6] ), .A2(\SB2_0_27/i0_4 ), .A3(n1091), 
        .ZN(n1895) );
  NAND3_X1 U6426 ( .A1(n3689), .A2(\SB2_0_5/i0_3 ), .A3(\RI3[0][160] ), .ZN(
        \SB2_0_5/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 U3413 ( .A1(\RI3[0][134] ), .A2(\SB2_0_9/i3[0] ), .ZN(
        \SB2_0_9/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_8/Component_Function_5/N1  ( .A1(\SB2_0_8/i0_0 ), .A2(
        \SB2_0_8/i3[0] ), .ZN(\SB2_0_8/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_0_17/Component_Function_5/N1  ( .A1(\SB2_0_17/i0_0 ), .A2(
        \SB2_0_17/i3[0] ), .ZN(\SB2_0_17/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U1526 ( .A1(\SB2_0_8/i0_3 ), .A2(\RI3[0][142] ), .A3(
        \SB2_0_8/i1[9] ), .ZN(\SB2_0_8/Component_Function_5/NAND4_in[2] ) );
  INV_X1 \SB2_0_3/INV_0  ( .I(\SB1_0_8/buf_output[0] ), .ZN(\SB2_0_3/i3[0] )
         );
  NAND3_X1 U9388 ( .A1(\SB2_0_16/i0[9] ), .A2(\SB2_0_16/i0_4 ), .A3(
        \SB2_0_16/i0[6] ), .ZN(n3819) );
  INV_X4 \SB2_0_2/INV_3  ( .I(\SB2_0_2/i0[10] ), .ZN(\SB2_0_2/i0[8] ) );
  BUF_X2 \SB2_0_15/BUF_0  ( .I(\RI3[0][96] ), .Z(\SB2_0_15/i0[9] ) );
  BUF_X2 \SB2_0_30/BUF_0  ( .I(\SB1_0_3/buf_output[0] ), .Z(\SB2_0_30/i0[9] )
         );
  BUF_X2 \SB2_0_0/BUF_0  ( .I(\SB1_0_5/buf_output[0] ), .Z(\SB2_0_0/i0[9] ) );
  BUF_X2 U3379 ( .I(\SB1_0_27/buf_output[4] ), .Z(\RI3[0][34] ) );
  CLKBUF_X2 \SB2_0_6/BUF_1  ( .I(\SB1_0_10/buf_output[1] ), .Z(\SB2_0_6/i0[6] ) );
  CLKBUF_X2 \SB2_0_4/BUF_0  ( .I(\RI3[0][162] ), .Z(\SB2_0_4/i0[9] ) );
  CLKBUF_X2 \SB2_0_12/BUF_1  ( .I(\SB1_0_16/buf_output[1] ), .Z(
        \SB2_0_12/i0[6] ) );
  BUF_X2 U1604 ( .I(\RI3[0][80] ), .Z(\SB2_0_18/i0_0 ) );
  CLKBUF_X2 \SB2_0_4/BUF_1  ( .I(\RI3[0][163] ), .Z(\SB2_0_4/i0[6] ) );
  BUF_X2 \SB2_0_0/BUF_1  ( .I(\SB1_0_4/buf_output[1] ), .Z(\SB2_0_0/i0[6] ) );
  BUF_X2 \SB2_0_20/BUF_2  ( .I(\RI3[0][68] ), .Z(\SB2_0_20/i0_0 ) );
  INV_X1 \SB2_0_4/INV_4  ( .I(\RI3[0][166] ), .ZN(\SB2_0_4/i0[7] ) );
  BUF_X2 \SB2_0_28/BUF_1  ( .I(\SB1_0_0/buf_output[1] ), .Z(\SB2_0_28/i0[6] )
         );
  INV_X2 U5705 ( .I(n2753), .ZN(\SB2_0_1/i0_4 ) );
  INV_X1 \SB2_0_18/INV_0  ( .I(\SB1_0_23/buf_output[0] ), .ZN(\SB2_0_18/i3[0] ) );
  INV_X1 U1530 ( .I(\RI3[0][180] ), .ZN(\SB2_0_1/i3[0] ) );
  INV_X1 U2514 ( .I(\RI3[0][61] ), .ZN(\SB2_0_21/i1_7 ) );
  INV_X1 \SB2_0_10/INV_1  ( .I(\RI3[0][127] ), .ZN(\SB2_0_10/i1_7 ) );
  INV_X1 \SB2_0_17/INV_1  ( .I(\SB1_0_21/buf_output[1] ), .ZN(\SB2_0_17/i1_7 )
         );
  INV_X1 U3012 ( .I(\SB1_0_11/buf_output[5] ), .ZN(\SB2_0_11/i1_5 ) );
  INV_X1 U1777 ( .I(\SB1_0_0/buf_output[5] ), .ZN(\SB2_0_0/i1_5 ) );
  INV_X1 \SB2_0_24/INV_5  ( .I(\SB1_0_24/buf_output[5] ), .ZN(\SB2_0_24/i1_5 )
         );
  INV_X1 U1959 ( .I(\RI3[0][142] ), .ZN(\SB2_0_8/i0[7] ) );
  NAND3_X1 \SB2_0_23/Component_Function_1/N2  ( .A1(\SB2_0_23/i0_3 ), .A2(
        \SB2_0_23/i1_7 ), .A3(\SB2_0_23/i0[8] ), .ZN(
        \SB2_0_23/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 U5089 ( .A1(\SB2_0_4/i0_3 ), .A2(\SB2_0_4/i1[9] ), .ZN(n1454) );
  NAND3_X1 \SB2_0_7/Component_Function_3/N3  ( .A1(\SB2_0_7/i1[9] ), .A2(
        \SB2_0_7/i1_7 ), .A3(\RI3[0][147] ), .ZN(
        \SB2_0_7/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_28/Component_Function_4/N2  ( .A1(\SB2_0_28/i3[0] ), .A2(
        \SB2_0_28/i0_0 ), .A3(\SB2_0_28/i1_7 ), .ZN(
        \SB2_0_28/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_16/Component_Function_2/N1  ( .A1(\SB2_0_16/i1_5 ), .A2(
        \SB2_0_16/i0[10] ), .A3(\SB2_0_16/i1[9] ), .ZN(
        \SB2_0_16/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U9534 ( .A1(\SB2_0_28/i0_3 ), .A2(\SB2_0_28/i0[10] ), .A3(
        \RI3[0][18] ), .ZN(\SB2_0_28/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_27/Component_Function_2/N1  ( .A1(\SB2_0_27/i1_5 ), .A2(
        \SB2_0_27/i0[10] ), .A3(\SB2_0_27/i1[9] ), .ZN(
        \SB2_0_27/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U9833 ( .A1(\SB2_0_9/i0_3 ), .A2(\RI3[0][134] ), .A3(\SB2_0_9/i0_4 ), .ZN(\SB2_0_9/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_1/Component_Function_4/N2  ( .A1(\SB2_0_1/i3[0] ), .A2(
        \SB2_0_1/i0_0 ), .A3(\SB2_0_1/i1_7 ), .ZN(
        \SB2_0_1/Component_Function_4/NAND4_in[1] ) );
  NAND2_X1 \SB2_0_24/Component_Function_1/N1  ( .A1(\SB2_0_24/i0_3 ), .A2(
        \SB2_0_24/i1[9] ), .ZN(\SB2_0_24/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_6/Component_Function_3/N4  ( .A1(\SB2_0_6/i1_5 ), .A2(
        \SB2_0_6/i0[8] ), .A3(\SB2_0_6/i3[0] ), .ZN(
        \SB2_0_6/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U9296 ( .A1(\SB2_0_26/i0[8] ), .A2(\SB2_0_26/i1_5 ), .A3(
        \SB2_0_26/i3[0] ), .ZN(\SB2_0_26/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_7/Component_Function_3/N4  ( .A1(\SB2_0_7/i1_5 ), .A2(
        \SB2_0_7/i0[8] ), .A3(\SB2_0_7/i3[0] ), .ZN(
        \SB2_0_7/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U4115 ( .A1(\SB2_0_15/i3[0] ), .A2(\SB2_0_15/i1_5 ), .A3(
        \SB2_0_15/i0[8] ), .ZN(\SB2_0_15/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U11185 ( .A1(\SB2_0_10/i0[10] ), .A2(\SB2_0_10/i1[9] ), .A3(
        \SB2_0_10/i1_7 ), .ZN(n4730) );
  NAND3_X1 \SB2_0_9/Component_Function_1/N4  ( .A1(\SB2_0_9/i1_7 ), .A2(
        \SB2_0_9/i0[8] ), .A3(\SB2_0_9/i0_4 ), .ZN(
        \SB2_0_9/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U1093 ( .A1(\SB2_0_23/i0_0 ), .A2(\SB2_0_23/i1_5 ), .A3(
        \SB2_0_23/i0_4 ), .ZN(\SB2_0_23/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U1982 ( .A1(\SB2_0_9/i1[9] ), .A2(n5518), .A3(\SB2_0_9/i0_4 ), .ZN(
        \SB2_0_9/Component_Function_4/NAND4_in[3] ) );
  NAND2_X1 \SB2_0_21/Component_Function_5/N1  ( .A1(\SB2_0_21/i0_0 ), .A2(
        \SB2_0_21/i3[0] ), .ZN(\SB2_0_21/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_10/Component_Function_0/N2  ( .A1(\SB2_0_10/i0[8] ), .A2(
        n2738), .A3(\SB2_0_10/i0[6] ), .ZN(
        \SB2_0_10/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_10/Component_Function_3/N2  ( .A1(\SB2_0_10/i0_0 ), .A2(
        \SB2_0_10/i0_3 ), .A3(\SB2_0_10/i0_4 ), .ZN(
        \SB2_0_10/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_26/Component_Function_2/N1  ( .A1(\SB2_0_26/i1_5 ), .A2(
        \SB2_0_26/i0[10] ), .A3(\SB2_0_26/i1[9] ), .ZN(
        \SB2_0_26/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U1090 ( .A1(\SB2_0_20/i0[9] ), .A2(\SB2_0_20/i0[6] ), .A3(
        \SB2_0_20/i1_5 ), .ZN(\SB2_0_20/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_8/Component_Function_1/N2  ( .A1(\SB2_0_8/i0_3 ), .A2(
        \SB2_0_8/i1_7 ), .A3(\SB2_0_8/i0[8] ), .ZN(
        \SB2_0_8/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U9964 ( .A1(\RI3[0][191] ), .A2(\SB2_0_0/i0[6] ), .A3(
        \SB2_0_0/i1[9] ), .ZN(n4078) );
  NAND3_X1 \SB2_0_25/Component_Function_3/N1  ( .A1(\SB2_0_25/i1[9] ), .A2(
        \SB2_0_25/i0_3 ), .A3(\RI3[0][37] ), .ZN(
        \SB2_0_25/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_20/Component_Function_1/N4  ( .A1(\SB2_0_20/i1_7 ), .A2(
        \SB2_0_20/i0[8] ), .A3(\SB2_0_20/i0_4 ), .ZN(
        \SB2_0_20/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U6240 ( .A1(\SB2_0_11/i0[8] ), .A2(\SB2_0_11/i0_3 ), .A3(n1911), 
        .ZN(\SB2_0_11/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_15/Component_Function_4/N4  ( .A1(\SB2_0_15/i1[9] ), .A2(
        \SB2_0_15/i1_5 ), .A3(\RI3[0][100] ), .ZN(
        \SB2_0_15/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U1144 ( .A1(\SB2_0_0/i0[9] ), .A2(\SB2_0_0/i0[6] ), .A3(
        \RI3[0][190] ), .ZN(\SB2_0_0/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_18/Component_Function_3/N4  ( .A1(\SB2_0_18/i1_5 ), .A2(
        \SB2_0_18/i0[8] ), .A3(\SB2_0_18/i3[0] ), .ZN(
        \SB2_0_18/Component_Function_3/NAND4_in[3] ) );
  INV_X2 \SB2_0_17/INV_4  ( .I(\RI3[0][88] ), .ZN(\SB2_0_17/i0[7] ) );
  NAND3_X1 U9295 ( .A1(\SB2_0_8/i0[6] ), .A2(\SB2_0_8/i1_5 ), .A3(
        \SB2_0_8/i0[9] ), .ZN(\SB2_0_8/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U3159 ( .A1(n2774), .A2(\SB2_0_19/i0[6] ), .A3(\SB2_0_19/i0_0 ), 
        .ZN(n885) );
  NAND3_X1 \SB2_0_19/Component_Function_5/N4  ( .A1(\SB2_0_19/i0[9] ), .A2(
        \SB2_0_19/i0[6] ), .A3(\RI3[0][76] ), .ZN(
        \SB2_0_19/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U3792 ( .A1(\SB2_0_21/i0[9] ), .A2(\SB2_0_21/i0_4 ), .A3(
        \SB2_0_21/i0[6] ), .ZN(n1125) );
  NAND3_X1 \SB2_0_17/Component_Function_1/N2  ( .A1(\SB2_0_17/i0_3 ), .A2(
        \SB2_0_17/i1_7 ), .A3(\SB2_0_17/i0[8] ), .ZN(
        \SB2_0_17/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_27/Component_Function_3/N2  ( .A1(\SB2_0_27/i0_0 ), .A2(
        \SB2_0_27/i0_3 ), .A3(\SB2_0_27/i0_4 ), .ZN(
        \SB2_0_27/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_28/Component_Function_1/N4  ( .A1(\SB2_0_28/i1_7 ), .A2(
        \SB2_0_28/i0[8] ), .A3(\RI3[0][22] ), .ZN(
        \SB2_0_28/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U1525 ( .A1(\SB2_0_8/i1_5 ), .A2(\SB2_0_8/i0[10] ), .A3(
        \SB2_0_8/i1[9] ), .ZN(\SB2_0_8/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_8/Component_Function_2/N4  ( .A1(\SB2_0_8/i1_5 ), .A2(
        \SB2_0_8/i0_0 ), .A3(\RI3[0][142] ), .ZN(
        \SB2_0_8/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_23/Component_Function_2/N1  ( .A1(\SB2_0_23/i1_5 ), .A2(
        \SB2_0_23/i0[10] ), .A3(\SB2_0_23/i1[9] ), .ZN(
        \SB2_0_23/Component_Function_2/NAND4_in[0] ) );
  INV_X1 \SB2_0_14/INV_1  ( .I(\RI3[0][103] ), .ZN(\SB2_0_14/i1_7 ) );
  NAND3_X1 \SB2_0_15/Component_Function_1/N2  ( .A1(\SB2_0_15/i0_3 ), .A2(
        \SB2_0_15/i1_7 ), .A3(\SB2_0_15/i0[8] ), .ZN(
        \SB2_0_15/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_23/Component_Function_1/N4  ( .A1(\SB2_0_23/i1_7 ), .A2(
        \SB2_0_23/i0[8] ), .A3(\SB2_0_23/i0_4 ), .ZN(
        \SB2_0_23/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_27/Component_Function_3/N3  ( .A1(\SB2_0_27/i1[9] ), .A2(
        \SB2_0_27/i1_7 ), .A3(\SB2_0_27/i0[10] ), .ZN(
        \SB2_0_27/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_28/Component_Function_1/N2  ( .A1(\SB2_0_28/i0_3 ), .A2(
        \SB2_0_28/i1_7 ), .A3(\SB2_0_28/i0[8] ), .ZN(
        \SB2_0_28/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U8627 ( .A1(\SB2_0_5/i0_3 ), .A2(\SB2_0_5/i0_0 ), .A3(\RI3[0][160] ), .ZN(\SB2_0_5/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3558 ( .A1(\SB2_0_24/i1_7 ), .A2(\SB2_0_24/i0_3 ), .A3(
        \SB2_0_24/i0[8] ), .ZN(n1688) );
  INV_X2 \SB2_0_15/INV_4  ( .I(\RI3[0][100] ), .ZN(\SB2_0_15/i0[7] ) );
  NAND3_X1 \SB2_0_24/Component_Function_0/N3  ( .A1(\SB2_0_24/i0[10] ), .A2(
        \RI3[0][46] ), .A3(\SB2_0_24/i0_3 ), .ZN(
        \SB2_0_24/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB2_0_9/Component_Function_1/N1  ( .A1(\SB2_0_9/i0_3 ), .A2(
        \SB2_0_9/i1[9] ), .ZN(\SB2_0_9/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_1/Component_Function_4/N1  ( .A1(\SB2_0_1/i0[9] ), .A2(
        \SB2_0_1/i0_0 ), .A3(\SB2_0_1/i0[8] ), .ZN(
        \SB2_0_1/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U10108 ( .A1(\SB2_0_15/i0_3 ), .A2(\SB2_0_15/i1[9] ), .A3(
        \SB2_0_15/i0[6] ), .ZN(\SB2_0_15/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U3268 ( .A1(\SB2_0_27/i0[10] ), .A2(\SB2_0_27/i0_3 ), .A3(n2679), 
        .ZN(n943) );
  NAND3_X1 U10856 ( .A1(\SB2_0_6/i0[9] ), .A2(\SB2_0_6/i1_5 ), .A3(
        \SB2_0_6/i0[6] ), .ZN(n4533) );
  NAND2_X1 \SB2_0_6/Component_Function_1/N1  ( .A1(\RI3[0][155] ), .A2(
        \SB2_0_6/i1[9] ), .ZN(\SB2_0_6/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U4227 ( .A1(\SB2_0_15/i0_3 ), .A2(\RI3[0][100] ), .A3(
        \SB2_0_15/i1[9] ), .ZN(n1306) );
  NAND3_X1 \SB2_0_10/Component_Function_1/N2  ( .A1(\SB2_0_10/i0_3 ), .A2(
        \SB2_0_10/i1_7 ), .A3(\SB2_0_10/i0[8] ), .ZN(
        \SB2_0_10/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_0_3/Component_Function_4/N4  ( .A1(\SB2_0_3/i1[9] ), .A2(
        \SB2_0_3/i1_5 ), .A3(\RI3[0][172] ), .ZN(
        \SB2_0_3/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U10700 ( .A1(\SB2_0_11/i0[7] ), .A2(\SB2_0_11/i0_0 ), .A3(
        \SB2_0_11/i0_3 ), .ZN(n4445) );
  NAND3_X1 U7348 ( .A1(\SB2_0_23/i3[0] ), .A2(\SB2_0_23/i1_5 ), .A3(
        \SB2_0_23/i0[8] ), .ZN(n2540) );
  NAND3_X1 \SB2_0_17/Component_Function_3/N2  ( .A1(\SB2_0_17/i0_0 ), .A2(
        \SB2_0_17/i0_3 ), .A3(\RI3[0][88] ), .ZN(
        \SB2_0_17/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U10147 ( .A1(\SB2_0_23/i0[10] ), .A2(\SB2_0_23/i1_7 ), .A3(
        \SB2_0_23/i1[9] ), .ZN(\SB2_0_23/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_0/Component_Function_1/N2  ( .A1(\RI3[0][191] ), .A2(
        \SB2_0_0/i1_7 ), .A3(\SB2_0_0/i0[8] ), .ZN(
        \SB2_0_0/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U1974 ( .A1(\SB2_0_20/i0[7] ), .A2(\SB2_0_20/i0[6] ), .A3(
        \SB2_0_20/i0[8] ), .ZN(n1270) );
  NAND3_X1 U9268 ( .A1(\SB2_0_14/i0[8] ), .A2(\SB2_0_14/i1_7 ), .A3(
        \RI3[0][106] ), .ZN(\SB2_0_14/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U1570 ( .A1(\SB2_0_18/i0[10] ), .A2(\SB2_0_18/i1_5 ), .A3(
        \SB2_0_18/i1[9] ), .ZN(\SB2_0_18/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_15/Component_Function_2/N1  ( .A1(\SB2_0_15/i1_5 ), .A2(
        \SB2_0_15/i0[10] ), .A3(\SB2_0_15/i1[9] ), .ZN(
        \SB2_0_15/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_30/Component_Function_4/N1  ( .A1(\SB2_0_30/i0[9] ), .A2(
        \SB2_0_30/i0_0 ), .A3(\SB2_0_30/i0[8] ), .ZN(
        \SB2_0_30/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U2969 ( .A1(\SB2_0_30/i3[0] ), .A2(\SB2_0_30/i1_5 ), .A3(
        \SB2_0_30/i0[8] ), .ZN(\SB2_0_30/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_0_22/Component_Function_1/N3  ( .A1(\SB2_0_22/i1_5 ), .A2(
        \SB2_0_22/i0[6] ), .A3(\RI3[0][54] ), .ZN(
        \SB2_0_22/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U2767 ( .A1(\SB2_0_1/i1_7 ), .A2(\SB2_0_1/i0[8] ), .A3(
        \SB2_0_1/i0_4 ), .ZN(\SB2_0_1/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U8408 ( .A1(\SB2_0_18/i0[9] ), .A2(\SB2_0_18/i0_3 ), .A3(
        \SB2_0_18/i0[8] ), .ZN(n3572) );
  NAND3_X1 U7510 ( .A1(\SB2_0_8/i0_3 ), .A2(\SB2_0_8/i0[9] ), .A3(
        \SB2_0_8/i0[10] ), .ZN(\SB2_0_8/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U8551 ( .A1(\SB2_0_23/i0_3 ), .A2(\SB2_0_23/i0_0 ), .A3(
        \SB2_0_23/i0_4 ), .ZN(n3618) );
  NAND3_X1 U6732 ( .A1(\SB2_0_2/i0[8] ), .A2(\RI3[0][176] ), .A3(
        \SB2_0_2/i0[9] ), .ZN(\SB2_0_2/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_28/Component_Function_3/N4  ( .A1(\SB2_0_28/i1_5 ), .A2(
        \SB2_0_28/i0[8] ), .A3(\SB2_0_28/i3[0] ), .ZN(
        \SB2_0_28/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U6508 ( .A1(\SB2_0_1/i0_3 ), .A2(\SB2_0_1/i0_0 ), .A3(n5054), .ZN(
        n3289) );
  NAND3_X1 U1524 ( .A1(\SB2_0_8/i1[9] ), .A2(\SB2_0_8/i1_7 ), .A3(
        \SB2_0_8/i0[10] ), .ZN(\SB2_0_8/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_31/Component_Function_4/N3  ( .A1(\SB2_0_31/i0[9] ), .A2(
        \SB2_0_31/i0[10] ), .A3(\SB2_0_31/i0_3 ), .ZN(
        \SB2_0_31/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U10312 ( .A1(\RI3[0][39] ), .A2(\SB2_0_25/i0[9] ), .A3(
        \SB2_0_25/i0_3 ), .ZN(\SB2_0_25/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_7/Component_Function_1/N4  ( .A1(\SB2_0_7/i1_7 ), .A2(
        \SB2_0_7/i0[8] ), .A3(\SB1_0_8/buf_output[4] ), .ZN(
        \SB2_0_7/Component_Function_1/NAND4_in[3] ) );
  NAND2_X1 \SB2_0_7/Component_Function_0/N1  ( .A1(\SB2_0_7/i0[10] ), .A2(
        \SB2_0_7/i0[9] ), .ZN(\SB2_0_7/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_0_2/Component_Function_0/N2  ( .A1(\SB2_0_2/i0[8] ), .A2(
        \SB2_0_2/i0[7] ), .A3(\SB2_0_2/i0[6] ), .ZN(
        \SB2_0_2/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U5214 ( .A1(\SB2_0_21/i0[6] ), .A2(\SB2_0_21/i1_5 ), .A3(
        \SB2_0_21/i0[9] ), .ZN(\SB2_0_21/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_0_28/Component_Function_3/N1  ( .A1(\SB2_0_28/i1[9] ), .A2(
        \SB2_0_28/i0_3 ), .A3(\SB2_0_28/i0[6] ), .ZN(
        \SB2_0_28/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U8601 ( .A1(\SB2_0_18/i0[9] ), .A2(\SB2_0_18/i0[6] ), .A3(
        \RI3[0][82] ), .ZN(n3633) );
  NAND3_X1 U3404 ( .A1(\SB2_0_15/i0[10] ), .A2(\RI3[0][100] ), .A3(
        \SB2_0_15/i0_3 ), .ZN(n904) );
  NAND3_X1 U6058 ( .A1(\SB2_0_1/i0[10] ), .A2(\SB2_0_1/i0[6] ), .A3(
        \SB2_0_1/i0_0 ), .ZN(\SB2_0_1/Component_Function_5/NAND4_in[1] ) );
  INV_X2 U6590 ( .I(\RI5[0][5] ), .ZN(n2673) );
  BUF_X2 U46 ( .I(Key[12]), .Z(n132) );
  NAND4_X1 U5723 ( .A1(\SB2_0_25/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_0_25/Component_Function_1/NAND4_in[0] ), .A3(n1804), .A4(
        \SB2_0_25/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_0_25/buf_output[1] ) );
  INV_X1 U6 ( .I(n25), .ZN(n548) );
  BUF_X2 \SB2_0_6/BUF_4_0  ( .I(\SB2_0_6/buf_output[4] ), .Z(\RI5[0][160] ) );
  INV_X1 \SB1_1_2/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[174] ), .ZN(
        \SB1_1_2/i3[0] ) );
  INV_X1 \SB1_1_23/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[48] ), .ZN(
        \SB1_1_23/i3[0] ) );
  INV_X1 \SB1_1_0/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[186] ), .ZN(
        \SB1_1_0/i3[0] ) );
  INV_X1 \SB1_1_8/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[138] ), .ZN(
        \SB1_1_8/i3[0] ) );
  INV_X1 \SB1_1_14/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[103] ), .ZN(
        \SB1_1_14/i1_7 ) );
  INV_X1 \SB1_1_11/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[121] ), .ZN(
        \SB1_1_11/i1_7 ) );
  NAND3_X1 \SB1_1_31/Component_Function_4/N2  ( .A1(\SB1_1_31/i3[0] ), .A2(
        \SB1_1_31/i0_0 ), .A3(\SB1_1_31/i1_7 ), .ZN(
        \SB1_1_31/Component_Function_4/NAND4_in[1] ) );
  INV_X1 \SB1_1_14/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[102] ), .ZN(
        \SB1_1_14/i3[0] ) );
  NAND3_X1 \SB1_1_31/Component_Function_4/N3  ( .A1(\SB1_1_31/i0[9] ), .A2(
        \SB1_1_31/i0[10] ), .A3(\SB1_1_31/i0_3 ), .ZN(
        \SB1_1_31/Component_Function_4/NAND4_in[2] ) );
  INV_X1 \SB1_1_12/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[114] ), .ZN(
        \SB1_1_12/i3[0] ) );
  INV_X1 \SB1_1_0/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[187] ), .ZN(
        \SB1_1_0/i1_7 ) );
  INV_X1 \SB1_1_2/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[179] ), .ZN(
        \SB1_1_2/i1_5 ) );
  BUF_X2 U9039 ( .I(\MC_ARK_ARC_1_0/buf_output[13] ), .Z(\SB1_1_29/i0[6] ) );
  INV_X1 \SB1_1_16/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[95] ), .ZN(
        \SB1_1_16/i1_5 ) );
  CLKBUF_X2 \SB1_1_15/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[97] ), .Z(
        \SB1_1_15/i0[6] ) );
  CLKBUF_X2 \SB1_1_25/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[40] ), .Z(
        \SB1_1_25/i0_4 ) );
  BUF_X2 \SB1_1_24/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[46] ), .Z(
        \SB1_1_24/i0_4 ) );
  BUF_X2 \SB1_1_14/BUF_4  ( .I(\MC_ARK_ARC_1_0/buf_output[106] ), .Z(
        \SB1_1_14/i0_4 ) );
  INV_X1 \SB1_1_29/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[12] ), .ZN(
        \SB1_1_29/i3[0] ) );
  INV_X1 U3150 ( .I(\MC_ARK_ARC_1_0/buf_output[45] ), .ZN(\SB1_1_24/i0[8] ) );
  INV_X1 \SB1_1_21/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[65] ), .ZN(
        \SB1_1_21/i1_5 ) );
  INV_X1 \SB1_1_3/INV_3  ( .I(\MC_ARK_ARC_1_0/buf_output[171] ), .ZN(
        \SB1_1_3/i0[8] ) );
  INV_X1 \SB1_1_6/INV_5  ( .I(\MC_ARK_ARC_1_0/buf_output[155] ), .ZN(
        \SB1_1_6/i1_5 ) );
  INV_X1 \SB1_1_16/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[91] ), .ZN(
        \SB1_1_16/i1_7 ) );
  NAND3_X1 U1061 ( .A1(\SB1_1_31/i0_0 ), .A2(\SB1_1_31/i0[9] ), .A3(
        \SB1_1_31/i0[8] ), .ZN(n2557) );
  NAND2_X1 \SB1_1_2/Component_Function_0/N1  ( .A1(\SB1_1_2/i0[10] ), .A2(
        \SB1_1_2/i0[9] ), .ZN(\SB1_1_2/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_14/Component_Function_1/N1  ( .A1(\SB1_1_14/i0_3 ), .A2(
        \SB1_1_14/i1[9] ), .ZN(\SB1_1_14/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_11/Component_Function_0/N3  ( .A1(\SB1_1_11/i0[10] ), .A2(
        \SB1_1_11/i0_4 ), .A3(\SB1_1_11/i0_3 ), .ZN(
        \SB1_1_11/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3464 ( .A1(\SB1_1_20/i1_5 ), .A2(\SB1_1_20/i0[8] ), .A3(
        \SB1_1_20/i3[0] ), .ZN(\SB1_1_20/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U1010 ( .A1(\SB1_1_0/i0[9] ), .A2(\SB1_1_0/i0[8] ), .A3(
        \SB1_1_0/i0_0 ), .ZN(n1358) );
  NAND3_X1 U6992 ( .A1(\SB1_1_9/i0[10] ), .A2(\SB1_1_9/i1[9] ), .A3(
        \SB1_1_9/i1_5 ), .ZN(n3369) );
  INV_X1 \SB1_1_15/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[97] ), .ZN(
        \SB1_1_15/i1_7 ) );
  NAND3_X1 U3662 ( .A1(\SB1_1_10/i1_5 ), .A2(\SB1_1_10/i0[6] ), .A3(
        \SB1_1_10/i0[9] ), .ZN(\SB1_1_10/Component_Function_1/NAND4_in[2] ) );
  INV_X1 \SB1_1_26/INV_0  ( .I(\MC_ARK_ARC_1_0/buf_output[30] ), .ZN(
        \SB1_1_26/i3[0] ) );
  INV_X1 U8878 ( .I(\MC_ARK_ARC_1_0/buf_output[84] ), .ZN(\SB1_1_17/i3[0] ) );
  INV_X1 \SB1_1_28/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[19] ), .ZN(
        \SB1_1_28/i1_7 ) );
  NAND2_X1 U10510 ( .A1(\SB1_1_12/i0_0 ), .A2(\SB1_1_12/i3[0] ), .ZN(n1668) );
  INV_X1 \SB1_1_23/INV_1  ( .I(\MC_ARK_ARC_1_0/buf_output[49] ), .ZN(
        \SB1_1_23/i1_7 ) );
  INV_X1 U1036 ( .I(\MC_ARK_ARC_1_0/buf_output[126] ), .ZN(\SB1_1_10/i3[0] )
         );
  NAND2_X1 \SB1_1_29/Component_Function_5/N1  ( .A1(\SB1_1_29/i0_0 ), .A2(
        \SB1_1_29/i3[0] ), .ZN(\SB1_1_29/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U1020 ( .A1(\SB1_1_14/i1_5 ), .A2(\SB1_1_14/i0[6] ), .A3(
        \SB1_1_14/i0[9] ), .ZN(\SB1_1_14/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U6693 ( .A1(\SB1_1_19/i0_0 ), .A2(\SB1_1_19/i0[8] ), .A3(
        \SB1_1_19/i0[9] ), .ZN(\SB1_1_19/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_9/Component_Function_2/N3  ( .A1(\SB1_1_9/i0_3 ), .A2(
        \SB1_1_9/i0[8] ), .A3(\SB1_1_9/i0[9] ), .ZN(
        \SB1_1_9/Component_Function_2/NAND4_in[2] ) );
  NAND2_X1 \SB1_1_27/Component_Function_1/N1  ( .A1(\SB1_1_27/i0_3 ), .A2(
        \SB1_1_27/i1[9] ), .ZN(\SB1_1_27/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_18/Component_Function_5/N2  ( .A1(\SB1_1_18/i0_0 ), .A2(
        \SB1_1_18/i0[6] ), .A3(\SB1_1_18/i0[10] ), .ZN(
        \SB1_1_18/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB1_1_23/Component_Function_0/N1  ( .A1(\SB1_1_23/i0[10] ), .A2(
        \SB1_1_23/i0[9] ), .ZN(\SB1_1_23/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_25/Component_Function_3/N2  ( .A1(\SB1_1_25/i0_0 ), .A2(
        \SB1_1_25/i0_3 ), .A3(\SB1_1_25/i0_4 ), .ZN(
        \SB1_1_25/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U4726 ( .A1(\SB1_1_7/i0[10] ), .A2(\SB1_1_7/i0[9] ), .A3(
        \SB1_1_7/i0_3 ), .ZN(n3035) );
  BUF_X2 \SB1_1_13/BUF_1  ( .I(\MC_ARK_ARC_1_0/buf_output[109] ), .Z(
        \SB1_1_13/i0[6] ) );
  NAND3_X1 U8141 ( .A1(\SB1_1_19/i0[9] ), .A2(\SB1_1_19/i0[10] ), .A3(
        \SB1_1_19/i0_3 ), .ZN(n1494) );
  NAND3_X1 U10825 ( .A1(\SB1_1_2/i0[10] ), .A2(\SB1_1_2/i0[6] ), .A3(
        \SB1_1_2/i0_3 ), .ZN(\SB1_1_2/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U8942 ( .A1(\SB1_1_11/i0[6] ), .A2(\SB1_1_11/i1[9] ), .A3(
        \SB1_1_11/i0_3 ), .ZN(n4667) );
  NAND3_X1 U10131 ( .A1(\SB1_1_15/i0[8] ), .A2(\SB1_1_15/i1_5 ), .A3(
        \SB1_1_15/i3[0] ), .ZN(n1203) );
  NAND3_X1 \SB1_1_23/Component_Function_3/N2  ( .A1(\SB1_1_23/i0_0 ), .A2(
        \SB1_1_23/i0_3 ), .A3(\SB1_1_23/i0_4 ), .ZN(
        \SB1_1_23/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1377 ( .A1(\SB1_1_5/i1_7 ), .A2(\SB1_1_5/i0[8] ), .A3(
        \SB1_1_5/i0_4 ), .ZN(\SB1_1_5/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U6084 ( .A1(\SB1_1_21/i3[0] ), .A2(\SB1_1_21/i0[8] ), .A3(
        \SB1_1_21/i1_5 ), .ZN(n3229) );
  NAND3_X1 U9959 ( .A1(\SB1_1_2/i0[9] ), .A2(\SB1_1_2/i0[8] ), .A3(
        \SB1_1_2/i0_3 ), .ZN(n4105) );
  NAND3_X1 \SB1_1_3/Component_Function_1/N3  ( .A1(\SB1_1_3/i1_5 ), .A2(
        \SB1_1_3/i0[6] ), .A3(\SB1_1_3/i0[9] ), .ZN(
        \SB1_1_3/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1435 ( .A1(\SB1_1_10/i0_3 ), .A2(\SB1_1_10/i0[9] ), .A3(
        \SB1_1_10/i0[10] ), .ZN(n4301) );
  NAND3_X1 \SB1_1_12/Component_Function_2/N1  ( .A1(\SB1_1_12/i1_5 ), .A2(
        \SB1_1_12/i0[10] ), .A3(\SB1_1_12/i1[9] ), .ZN(
        \SB1_1_12/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U9633 ( .A1(\SB1_1_22/i0[9] ), .A2(\SB1_1_22/i0[8] ), .A3(
        \SB1_1_22/i0_0 ), .ZN(n3940) );
  NAND3_X1 U1449 ( .A1(\SB1_1_27/i0[10] ), .A2(\SB1_1_27/i1[9] ), .A3(
        \SB1_1_27/i1_7 ), .ZN(\SB1_1_27/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U7372 ( .A1(\SB1_1_16/i0_3 ), .A2(\SB1_1_16/i0[8] ), .A3(
        \SB1_1_16/i0[9] ), .ZN(n3423) );
  NAND3_X1 \SB1_1_6/Component_Function_0/N4  ( .A1(\SB1_1_6/i0[7] ), .A2(
        \SB1_1_6/i0_3 ), .A3(\SB1_1_6/i0_0 ), .ZN(
        \SB1_1_6/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U6570 ( .A1(\SB1_1_22/i0[9] ), .A2(\RI1[1][59] ), .A3(
        \SB1_1_22/i0[10] ), .ZN(n4356) );
  NAND3_X1 \SB1_1_19/Component_Function_3/N4  ( .A1(\SB1_1_19/i1_5 ), .A2(
        \SB1_1_19/i0[8] ), .A3(\SB1_1_19/i3[0] ), .ZN(
        \SB1_1_19/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U7496 ( .A1(\SB1_1_7/i0[8] ), .A2(\SB1_1_7/i1_5 ), .A3(
        \SB1_1_7/i3[0] ), .ZN(n4718) );
  NAND3_X1 \SB1_1_9/Component_Function_1/N2  ( .A1(\SB1_1_9/i0_3 ), .A2(
        \SB1_1_9/i1_7 ), .A3(\SB1_1_9/i0[8] ), .ZN(
        \SB1_1_9/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U4075 ( .A1(\SB1_1_25/i0[8] ), .A2(\SB1_1_25/i0_3 ), .A3(
        \SB1_1_25/i1_7 ), .ZN(n3895) );
  NAND3_X1 \SB1_1_30/Component_Function_0/N2  ( .A1(\SB1_1_30/i0[8] ), .A2(
        \SB1_1_30/i0[7] ), .A3(\SB1_1_30/i0[6] ), .ZN(
        \SB1_1_30/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U4983 ( .A1(\SB1_1_26/i0[10] ), .A2(\SB1_1_26/i1[9] ), .A3(
        \SB1_1_26/i1_7 ), .ZN(n1407) );
  NAND3_X1 \SB1_1_21/Component_Function_1/N2  ( .A1(\SB1_1_21/i0_3 ), .A2(
        \SB1_1_21/i1_7 ), .A3(\SB1_1_21/i0[8] ), .ZN(
        \SB1_1_21/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U1023 ( .A1(\SB1_1_7/i0[10] ), .A2(\SB1_1_7/i1[9] ), .A3(
        \SB1_1_7/i1_7 ), .ZN(\SB1_1_7/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U10331 ( .A1(\SB1_1_20/i0[8] ), .A2(\SB1_1_20/i1_7 ), .A3(
        \RI1[1][71] ), .ZN(\SB1_1_20/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_8/Component_Function_1/N3  ( .A1(n3647), .A2(\SB1_1_8/i0[6] ), .A3(\SB1_1_8/i0[9] ), .ZN(\SB1_1_8/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_24/Component_Function_2/N4  ( .A1(\SB1_1_24/i1_5 ), .A2(
        \SB1_1_24/i0_0 ), .A3(\SB1_1_24/i0_4 ), .ZN(
        \SB1_1_24/Component_Function_2/NAND4_in[3] ) );
  NAND2_X1 \SB1_1_24/Component_Function_5/N1  ( .A1(\SB1_1_24/i0_0 ), .A2(
        \SB1_1_24/i3[0] ), .ZN(\SB1_1_24/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_17/Component_Function_5/N1  ( .A1(\SB1_1_17/i0_0 ), .A2(
        \SB1_1_17/i3[0] ), .ZN(\SB1_1_17/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 U4271 ( .A1(\SB1_1_25/i0_0 ), .A2(\SB1_1_25/i3[0] ), .ZN(n1324) );
  NAND2_X1 \SB1_1_19/Component_Function_5/N1  ( .A1(\SB1_1_19/i0_0 ), .A2(
        \SB1_1_19/i3[0] ), .ZN(\SB1_1_19/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 U1164 ( .A1(\SB1_1_31/i0_0 ), .A2(\SB1_1_31/i3[0] ), .ZN(
        \SB1_1_31/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U1668 ( .A1(\RI1[1][143] ), .A2(\SB1_1_8/i0[8] ), .A3(
        \SB1_1_8/i0[9] ), .ZN(\SB1_1_8/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2007 ( .A1(\SB1_1_20/i1_5 ), .A2(\SB1_1_20/i0_0 ), .A3(
        \SB1_1_20/i0_4 ), .ZN(\SB1_1_20/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U9490 ( .A1(\SB1_1_17/i0_3 ), .A2(\SB1_1_17/i0[8] ), .A3(
        \SB1_1_17/i1_7 ), .ZN(n3872) );
  NAND2_X1 U7062 ( .A1(\SB1_1_21/i0[10] ), .A2(\SB1_1_21/i0[9] ), .ZN(n3378)
         );
  NAND3_X1 U9600 ( .A1(\SB1_1_9/i0_0 ), .A2(\SB1_1_9/i0_3 ), .A3(
        \SB1_1_9/i0[7] ), .ZN(n3920) );
  NAND2_X1 \SB1_1_20/Component_Function_1/N1  ( .A1(\SB1_1_20/i0_3 ), .A2(
        \SB1_1_20/i1[9] ), .ZN(\SB1_1_20/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_17/Component_Function_1/N4  ( .A1(\SB1_1_17/i1_7 ), .A2(
        \SB1_1_17/i0[8] ), .A3(\SB1_1_17/i0_4 ), .ZN(
        \SB1_1_17/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U6299 ( .A1(\SB1_1_28/i0[10] ), .A2(\SB1_1_28/i1[9] ), .A3(
        \SB1_1_28/i1_5 ), .ZN(n3264) );
  NAND3_X1 U3447 ( .A1(\SB1_1_0/i0_3 ), .A2(\SB1_1_0/i0_4 ), .A3(
        \SB1_1_0/i1[9] ), .ZN(\SB1_1_0/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB1_1_17/Component_Function_5/N3  ( .A1(\SB1_1_17/i1[9] ), .A2(
        \SB1_1_17/i0_4 ), .A3(\SB1_1_17/i0_3 ), .ZN(
        \SB1_1_17/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U6929 ( .A1(\SB1_1_0/i0[9] ), .A2(\SB1_1_0/i0[6] ), .A3(
        \SB1_1_0/i0_4 ), .ZN(n2315) );
  NAND3_X1 U6579 ( .A1(\SB1_1_17/i0_4 ), .A2(\SB1_1_17/i0[6] ), .A3(
        \SB1_1_17/i0[9] ), .ZN(n3302) );
  NAND3_X1 U5157 ( .A1(\SB1_1_13/i0[6] ), .A2(\SB1_1_13/i0[9] ), .A3(
        \SB1_1_13/i0_4 ), .ZN(\SB1_1_13/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U6753 ( .A1(\SB1_1_7/i0[10] ), .A2(\SB1_1_7/i0_0 ), .A3(
        \SB1_1_7/i0[6] ), .ZN(\SB1_1_7/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1732 ( .A1(\SB1_1_7/i0[9] ), .A2(\SB1_1_7/i0[6] ), .A3(
        \SB1_1_7/i0_4 ), .ZN(\SB1_1_7/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_21/Component_Function_1/N4  ( .A1(\SB1_1_21/i1_7 ), .A2(
        \SB1_1_21/i0[8] ), .A3(\SB1_1_21/i0_4 ), .ZN(
        \SB1_1_21/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_3/Component_Function_3/N1  ( .A1(\SB1_1_3/i1[9] ), .A2(
        \SB1_1_3/i0_3 ), .A3(\SB1_1_3/i0[6] ), .ZN(
        \SB1_1_3/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U1498 ( .A1(\SB1_1_9/i1[9] ), .A2(\SB1_1_9/i0_3 ), .A3(
        \SB1_1_9/i0[6] ), .ZN(\SB1_1_9/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_29/Component_Function_4/N3  ( .A1(\SB1_1_29/i0[9] ), .A2(
        \SB1_1_29/i0[10] ), .A3(\SB1_1_29/i0_3 ), .ZN(
        \SB1_1_29/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U7583 ( .A1(\SB1_1_23/i0[10] ), .A2(\SB1_1_23/i0_3 ), .A3(
        \SB1_1_23/i0[6] ), .ZN(\SB1_1_23/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_31/Component_Function_2/N2  ( .A1(\SB1_1_31/i0_3 ), .A2(
        \SB1_1_31/i0[10] ), .A3(\SB1_1_31/i0[6] ), .ZN(
        \SB1_1_31/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_20/Component_Function_0/N2  ( .A1(\SB1_1_20/i0[8] ), .A2(
        \SB1_1_20/i0[7] ), .A3(\SB1_1_20/i0[6] ), .ZN(
        \SB1_1_20/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U6094 ( .A1(\SB1_1_5/i0[10] ), .A2(\SB1_1_5/i1_7 ), .A3(
        \SB1_1_5/i1[9] ), .ZN(\SB1_1_5/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U1422 ( .A1(\SB1_1_2/i0[8] ), .A2(\SB1_1_2/i1_5 ), .A3(
        \SB1_1_2/i3[0] ), .ZN(n4388) );
  NAND3_X1 \SB1_1_9/Component_Function_4/N4  ( .A1(\SB1_1_9/i1[9] ), .A2(
        \SB1_1_9/i1_5 ), .A3(\SB1_1_9/i0_4 ), .ZN(
        \SB1_1_9/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_17/Component_Function_3/N4  ( .A1(\SB1_1_17/i1_5 ), .A2(
        \SB1_1_17/i0[8] ), .A3(\SB1_1_17/i3[0] ), .ZN(
        \SB1_1_17/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_1_27/Component_Function_4/N2  ( .A1(\SB1_1_27/i3[0] ), .A2(
        \SB1_1_27/i0_0 ), .A3(\SB1_1_27/i1_7 ), .ZN(
        \SB1_1_27/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U1410 ( .A1(\SB1_1_24/i0_3 ), .A2(\SB1_1_24/i1[9] ), .A3(
        \SB1_1_24/i0[6] ), .ZN(\SB1_1_24/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U1737 ( .A1(\SB1_1_27/i1[9] ), .A2(\SB1_1_27/i1_5 ), .A3(
        \SB1_1_27/i0_4 ), .ZN(\SB1_1_27/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U9029 ( .A1(\SB1_1_17/i1_5 ), .A2(\SB1_1_17/i0[10] ), .A3(
        \SB1_1_17/i1[9] ), .ZN(\SB1_1_17/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U5620 ( .A1(\SB1_1_31/i0_4 ), .A2(\SB1_1_31/i1_7 ), .A3(
        \SB1_1_31/i0[8] ), .ZN(n1710) );
  NAND3_X1 U7434 ( .A1(\SB1_1_10/i3[0] ), .A2(\SB1_1_10/i1_5 ), .A3(
        \SB1_1_10/i0[8] ), .ZN(n3434) );
  NAND3_X1 U1403 ( .A1(\SB1_1_6/i0_0 ), .A2(\SB1_1_6/i0_4 ), .A3(
        \SB1_1_6/i1_5 ), .ZN(n3234) );
  NAND2_X1 \SB1_1_26/Component_Function_1/N1  ( .A1(\SB1_1_26/i0_3 ), .A2(
        \SB1_1_26/i1[9] ), .ZN(\SB1_1_26/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_10/Component_Function_3/N3  ( .A1(\SB1_1_10/i1[9] ), .A2(
        \SB1_1_10/i1_7 ), .A3(\SB1_1_10/i0[10] ), .ZN(
        \SB1_1_10/Component_Function_3/NAND4_in[2] ) );
  NAND2_X1 \SB1_1_3/Component_Function_5/N1  ( .A1(\SB1_1_3/i0_0 ), .A2(
        \SB1_1_3/i3[0] ), .ZN(\SB1_1_3/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 U1018 ( .A1(\SB1_1_22/i0_0 ), .A2(\SB1_1_22/i3[0] ), .ZN(n1044) );
  NAND2_X1 \SB1_1_15/Component_Function_5/N1  ( .A1(\SB1_1_15/i0_0 ), .A2(
        \SB1_1_15/i3[0] ), .ZN(\SB1_1_15/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_27/Component_Function_5/N1  ( .A1(\SB1_1_27/i0_0 ), .A2(
        \SB1_1_27/i3[0] ), .ZN(\SB1_1_27/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB1_1_30/Component_Function_1/N1  ( .A1(\SB1_1_30/i0_3 ), .A2(
        \SB1_1_30/i1[9] ), .ZN(\SB1_1_30/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_1_13/Component_Function_0/N4  ( .A1(\SB1_1_13/i0[7] ), .A2(
        \SB1_1_13/i0_3 ), .A3(\SB1_1_13/i0_0 ), .ZN(
        \SB1_1_13/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U1420 ( .A1(\SB1_1_30/i0[8] ), .A2(\SB1_1_30/i0_4 ), .A3(
        \SB1_1_30/i1_7 ), .ZN(n4218) );
  NAND3_X1 U7337 ( .A1(\SB1_1_7/i0[9] ), .A2(\SB1_1_7/i1_5 ), .A3(
        \SB1_1_7/i0[6] ), .ZN(n3415) );
  INV_X1 \SB2_1_2/INV_0  ( .I(\SB1_1_7/buf_output[0] ), .ZN(\SB2_1_2/i3[0] )
         );
  NAND3_X1 U2009 ( .A1(\SB1_1_5/i0[6] ), .A2(\SB1_1_5/i1[9] ), .A3(
        \SB1_1_5/i0_3 ), .ZN(n1164) );
  NAND3_X1 U1395 ( .A1(\SB1_1_23/i1_5 ), .A2(\SB1_1_23/i0_4 ), .A3(
        \SB1_1_23/i1[9] ), .ZN(n3532) );
  NAND3_X1 U10410 ( .A1(\SB1_1_10/i0_3 ), .A2(\SB1_1_10/i0_0 ), .A3(
        \SB1_1_10/i0_4 ), .ZN(\SB1_1_10/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_31/Component_Function_2/N4  ( .A1(\SB1_1_31/i1_5 ), .A2(
        \SB1_1_31/i0_0 ), .A3(\SB1_1_31/i0_4 ), .ZN(
        \SB1_1_31/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U7953 ( .A1(\SB1_1_19/i0[6] ), .A2(\SB1_1_19/i1_5 ), .A3(
        \SB1_1_19/i0[9] ), .ZN(n3508) );
  NAND3_X1 U4631 ( .A1(\SB1_1_3/i0_0 ), .A2(\SB1_1_3/i0[6] ), .A3(
        \SB1_1_3/i0[10] ), .ZN(\SB1_1_3/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_1_28/Component_Function_5/N2  ( .A1(\SB1_1_28/i0_0 ), .A2(
        \SB1_1_28/i0[6] ), .A3(\SB1_1_28/i0[10] ), .ZN(
        \SB1_1_28/Component_Function_5/NAND4_in[1] ) );
  BUF_X2 U1519 ( .I(\SB1_1_10/buf_output[1] ), .Z(\SB2_1_6/i0[6] ) );
  INV_X1 \SB2_1_12/INV_0  ( .I(\SB1_1_17/buf_output[0] ), .ZN(\SB2_1_12/i3[0] ) );
  INV_X1 U7978 ( .I(\SB1_1_2/buf_output[0] ), .ZN(\SB2_1_29/i3[0] ) );
  NAND3_X1 U1029 ( .A1(\SB1_1_23/i0[10] ), .A2(\SB1_1_23/i0[9] ), .A3(
        \SB1_1_23/i0_3 ), .ZN(\SB1_1_23/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U7924 ( .A1(\SB1_1_23/i0_0 ), .A2(\SB1_1_23/i1_5 ), .A3(
        \SB1_1_23/i0_4 ), .ZN(n2868) );
  NAND3_X1 U1999 ( .A1(\SB1_1_11/i0_0 ), .A2(\SB1_1_11/i0[6] ), .A3(
        \SB1_1_11/i0[10] ), .ZN(\SB1_1_11/Component_Function_5/NAND4_in[1] )
         );
  NAND3_X1 U1002 ( .A1(\SB1_1_29/i0_0 ), .A2(\SB1_1_29/i0_3 ), .A3(
        \SB1_1_29/i0_4 ), .ZN(\SB1_1_29/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1207 ( .A1(\SB1_1_20/i0_0 ), .A2(\SB1_1_20/i0[10] ), .A3(
        \SB1_1_20/i0[6] ), .ZN(\SB1_1_20/Component_Function_5/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_23/Component_Function_5/N1  ( .A1(\SB2_1_23/i0_0 ), .A2(
        \SB2_1_23/i3[0] ), .ZN(\SB2_1_23/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 U2259 ( .A1(\SB2_1_29/i0_0 ), .A2(\SB2_1_29/i3[0] ), .ZN(
        \SB2_1_29/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_2/Component_Function_5/N1  ( .A1(\SB2_1_2/i0_0 ), .A2(
        \SB2_1_2/i3[0] ), .ZN(\SB2_1_2/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_18/Component_Function_5/N1  ( .A1(\SB2_1_18/i0_0 ), .A2(
        \SB2_1_18/i3[0] ), .ZN(\SB2_1_18/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_1_6/Component_Function_5/N1  ( .A1(\SB2_1_6/i0_0 ), .A2(
        \SB2_1_6/i3[0] ), .ZN(\SB2_1_6/Component_Function_5/NAND4_in[0] ) );
  CLKBUF_X2 \SB2_1_4/BUF_0  ( .I(\SB1_1_9/buf_output[0] ), .Z(\SB2_1_4/i0[9] )
         );
  BUF_X2 \SB2_1_13/BUF_1  ( .I(\SB1_1_17/buf_output[1] ), .Z(\SB2_1_13/i0[6] )
         );
  CLKBUF_X2 \SB2_1_7/BUF_0  ( .I(\SB1_1_12/buf_output[0] ), .Z(\SB2_1_7/i0[9] ) );
  BUF_X2 \SB2_1_16/BUF_0  ( .I(\SB1_1_21/buf_output[0] ), .Z(\SB2_1_16/i0[9] )
         );
  CLKBUF_X2 \SB2_1_17/BUF_0  ( .I(\SB1_1_22/buf_output[0] ), .Z(
        \SB2_1_17/i0[9] ) );
  BUF_X2 \SB2_1_13/BUF_2  ( .I(\RI3[1][110] ), .Z(\SB2_1_13/i0_0 ) );
  INV_X2 U10090 ( .I(n4149), .ZN(n578) );
  NAND2_X1 \SB2_1_25/Component_Function_5/N1  ( .A1(\SB2_1_25/i0_0 ), .A2(
        \SB2_1_25/i3[0] ), .ZN(\SB2_1_25/Component_Function_5/NAND4_in[0] ) );
  INV_X1 \SB2_1_10/INV_1  ( .I(\SB1_1_14/buf_output[1] ), .ZN(\SB2_1_10/i1_7 )
         );
  NAND2_X1 \SB2_1_17/Component_Function_5/N1  ( .A1(\SB2_1_17/i0_0 ), .A2(
        \SB2_1_17/i3[0] ), .ZN(\SB2_1_17/Component_Function_5/NAND4_in[0] ) );
  BUF_X2 \SB2_1_23/BUF_0  ( .I(\SB1_1_28/buf_output[0] ), .Z(\SB2_1_23/i0[9] )
         );
  INV_X1 \SB2_1_13/INV_1  ( .I(\SB1_1_17/buf_output[1] ), .ZN(\SB2_1_13/i1_7 )
         );
  NAND3_X1 U971 ( .A1(\SB2_1_19/i0_3 ), .A2(n1396), .A3(n578), .ZN(
        \SB2_1_19/Component_Function_5/NAND4_in[2] ) );
  BUF_X2 \SB2_1_15/BUF_0  ( .I(\SB1_1_20/buf_output[0] ), .Z(\SB2_1_15/i0[9] )
         );
  BUF_X2 \SB2_1_29/BUF_0  ( .I(\SB1_1_2/buf_output[0] ), .Z(\SB2_1_29/i0[9] )
         );
  CLKBUF_X2 \SB2_1_15/BUF_2  ( .I(\SB1_1_18/buf_output[2] ), .Z(
        \SB2_1_15/i0_0 ) );
  INV_X2 U10555 ( .I(\SB2_1_11/i0[7] ), .ZN(\SB1_1_12/buf_output[4] ) );
  INV_X1 U3480 ( .I(\SB1_1_20/buf_output[0] ), .ZN(\SB2_1_15/i3[0] ) );
  INV_X1 U7618 ( .I(\SB1_1_23/buf_output[1] ), .ZN(\SB2_1_19/i1_7 ) );
  INV_X1 \SB2_1_26/INV_1  ( .I(\SB1_1_30/buf_output[1] ), .ZN(\SB2_1_26/i1_7 )
         );
  INV_X1 U2873 ( .I(\SB1_1_4/buf_output[5] ), .ZN(\SB2_1_4/i1_5 ) );
  INV_X1 U3974 ( .I(\SB1_1_11/buf_output[5] ), .ZN(\SB2_1_11/i1_5 ) );
  INV_X1 \SB2_1_21/INV_1  ( .I(\SB1_1_25/buf_output[1] ), .ZN(\SB2_1_21/i1_7 )
         );
  NAND2_X1 \SB2_1_28/Component_Function_1/N1  ( .A1(\SB2_1_28/i0_3 ), .A2(
        \SB2_1_28/i1[9] ), .ZN(\SB2_1_28/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_11/Component_Function_4/N2  ( .A1(\SB2_1_11/i3[0] ), .A2(
        \SB2_1_11/i0_0 ), .A3(\SB2_1_11/i1_7 ), .ZN(
        \SB2_1_11/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U2853 ( .A1(\SB2_1_23/i3[0] ), .A2(\SB2_1_23/i1_5 ), .A3(
        \SB2_1_23/i0[8] ), .ZN(\SB2_1_23/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_15/Component_Function_3/N2  ( .A1(\SB2_1_15/i0_0 ), .A2(
        \SB2_1_15/i0_3 ), .A3(\SB2_1_15/i0_4 ), .ZN(
        \SB2_1_15/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3003 ( .A1(\SB2_1_22/i0_3 ), .A2(\SB2_1_22/i1_7 ), .A3(
        \SB2_1_22/i0[8] ), .ZN(\SB2_1_22/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U1294 ( .A1(\SB2_1_16/i0_3 ), .A2(\SB2_1_16/i0[10] ), .A3(
        \SB2_1_16/i0[9] ), .ZN(\SB2_1_16/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1362 ( .A1(\SB2_1_18/i0_0 ), .A2(n1379), .A3(\SB2_1_18/i0_3 ), 
        .ZN(n3357) );
  NAND3_X1 \SB2_1_8/Component_Function_1/N2  ( .A1(\SB2_1_8/i0_3 ), .A2(
        \SB2_1_8/i1_7 ), .A3(\SB2_1_8/i0[8] ), .ZN(
        \SB2_1_8/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_15/Component_Function_3/N3  ( .A1(\SB2_1_15/i1[9] ), .A2(
        \SB2_1_15/i1_7 ), .A3(\SB2_1_15/i0[10] ), .ZN(
        \SB2_1_15/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U981 ( .A1(\SB2_1_7/i0[10] ), .A2(\SB2_1_7/i0_3 ), .A3(n5790), .ZN(
        \SB2_1_7/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U8036 ( .A1(\SB2_1_19/i0_3 ), .A2(\SB1_1_22/buf_output[2] ), .A3(
        n578), .ZN(\SB2_1_19/Component_Function_3/NAND4_in[1] ) );
  NAND2_X1 U1349 ( .A1(\SB2_1_26/i0_0 ), .A2(\SB2_1_26/i3[0] ), .ZN(n3392) );
  NAND3_X1 U6419 ( .A1(\SB2_1_9/i0[10] ), .A2(\SB2_1_9/i1[9] ), .A3(
        \SB2_1_9/i1_7 ), .ZN(\SB2_1_9/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_2/Component_Function_4/N2  ( .A1(\SB2_1_2/i3[0] ), .A2(
        \SB2_1_2/i0_0 ), .A3(\SB2_1_2/i1_7 ), .ZN(
        \SB2_1_2/Component_Function_4/NAND4_in[1] ) );
  NAND2_X1 \SB2_1_1/Component_Function_0/N1  ( .A1(\SB2_1_1/i0[10] ), .A2(
        \SB2_1_1/i0[9] ), .ZN(\SB2_1_1/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_21/Component_Function_0/N4  ( .A1(\SB2_1_21/i0[7] ), .A2(
        \SB2_1_21/i0_3 ), .A3(\SB2_1_21/i0_0 ), .ZN(
        \SB2_1_21/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_27/Component_Function_0/N4  ( .A1(\SB2_1_27/i0[7] ), .A2(
        \SB2_1_27/i0_3 ), .A3(\SB2_1_27/i0_0 ), .ZN(
        \SB2_1_27/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U6317 ( .A1(\SB2_1_13/i0[10] ), .A2(n1117), .A3(\SB2_1_13/i0_4 ), 
        .ZN(n2018) );
  NAND3_X1 \SB2_1_15/Component_Function_3/N4  ( .A1(\SB2_1_15/i1_5 ), .A2(
        \SB2_1_15/i0[8] ), .A3(\SB2_1_15/i3[0] ), .ZN(
        \SB2_1_15/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_7/Component_Function_3/N4  ( .A1(\SB2_1_7/i1_5 ), .A2(
        \SB2_1_7/i0[8] ), .A3(\SB2_1_7/i3[0] ), .ZN(
        \SB2_1_7/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_2/Component_Function_2/N3  ( .A1(\SB2_1_2/i0_3 ), .A2(
        \SB2_1_2/i0[8] ), .A3(\SB2_1_2/i0[9] ), .ZN(
        \SB2_1_2/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2988 ( .A1(\SB2_1_16/i1_5 ), .A2(\SB2_1_16/i0[8] ), .A3(
        \SB2_1_16/i3[0] ), .ZN(\SB2_1_16/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U1321 ( .A1(\SB2_1_18/i3[0] ), .A2(\SB2_1_18/i1_5 ), .A3(
        \SB2_1_18/i0[8] ), .ZN(n4349) );
  NAND3_X1 U1330 ( .A1(n2687), .A2(\SB2_1_0/i1_7 ), .A3(\SB2_1_0/i0[8] ), .ZN(
        n4387) );
  NAND3_X1 \SB2_1_12/Component_Function_2/N1  ( .A1(\SB2_1_12/i1_5 ), .A2(
        \SB2_1_12/i0[10] ), .A3(\SB2_1_12/i1[9] ), .ZN(
        \SB2_1_12/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U10513 ( .A1(\SB2_1_19/i0[8] ), .A2(\SB2_1_19/i1_5 ), .A3(
        \SB2_1_19/i3[0] ), .ZN(n4549) );
  NAND3_X1 \SB2_1_4/Component_Function_3/N3  ( .A1(n3660), .A2(\SB2_1_4/i1_7 ), 
        .A3(\SB2_1_4/i0[10] ), .ZN(\SB2_1_4/Component_Function_3/NAND4_in[2] )
         );
  NAND3_X1 U5920 ( .A1(\SB2_1_13/i0_3 ), .A2(\SB1_1_18/buf_output[0] ), .A3(
        \SB2_1_13/i0[8] ), .ZN(\SB2_1_13/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_11/Component_Function_2/N2  ( .A1(\SB2_1_11/i0_3 ), .A2(
        \SB2_1_11/i0[10] ), .A3(\SB2_1_11/i0[6] ), .ZN(
        \SB2_1_11/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U1636 ( .A1(\SB2_1_3/i1_7 ), .A2(\SB2_1_3/i0[8] ), .A3(n5208), .ZN(
        \SB2_1_3/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U3491 ( .A1(\SB2_1_20/i0_3 ), .A2(\SB2_1_20/i1_7 ), .A3(
        \SB2_1_20/i0[8] ), .ZN(\SB2_1_20/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_11/Component_Function_1/N2  ( .A1(\SB2_1_11/i0_3 ), .A2(
        \SB2_1_11/i1_7 ), .A3(\SB2_1_11/i0[8] ), .ZN(
        \SB2_1_11/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U1301 ( .A1(\SB2_1_2/i0_4 ), .A2(\SB2_1_2/i1[9] ), .A3(
        \SB2_1_2/i1_5 ), .ZN(n4323) );
  NAND3_X1 U8875 ( .A1(\SB2_1_5/i1_5 ), .A2(\SB2_1_5/i0[6] ), .A3(
        \SB2_1_5/i0[9] ), .ZN(\SB2_1_5/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_1_2/Component_Function_1/N3  ( .A1(\SB2_1_2/i1_5 ), .A2(
        \SB2_1_2/i0[6] ), .A3(\SB2_1_2/i0[9] ), .ZN(
        \SB2_1_2/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U6827 ( .A1(\SB2_1_1/i0[9] ), .A2(\SB2_1_1/i0[6] ), .A3(
        \SB2_1_1/i1_5 ), .ZN(\SB2_1_1/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1327 ( .A1(\SB2_1_25/i0[6] ), .A2(\SB2_1_25/i1_5 ), .A3(
        \SB2_1_25/i0[9] ), .ZN(n3002) );
  NAND3_X1 \SB2_1_10/Component_Function_1/N3  ( .A1(\SB2_1_10/i1_5 ), .A2(
        \SB2_1_10/i0[6] ), .A3(\SB2_1_10/i0[9] ), .ZN(
        \SB2_1_10/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U11181 ( .A1(\SB2_1_17/i0[10] ), .A2(\SB2_1_17/i1_5 ), .A3(
        \SB2_1_17/i1[9] ), .ZN(\SB2_1_17/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_31/Component_Function_0/N3  ( .A1(\SB2_1_31/i0[10] ), .A2(
        \SB2_1_31/i0_4 ), .A3(\SB2_1_31/i0_3 ), .ZN(
        \SB2_1_31/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB2_1_13/Component_Function_1/N1  ( .A1(\SB2_1_13/i0_3 ), .A2(
        \SB2_1_13/i1[9] ), .ZN(\SB2_1_13/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_18/Component_Function_4/N4  ( .A1(\SB2_1_18/i1[9] ), .A2(
        \SB2_1_18/i1_5 ), .A3(\SB2_1_18/i0_4 ), .ZN(
        \SB2_1_18/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_6/Component_Function_3/N4  ( .A1(\SB2_1_6/i1_5 ), .A2(
        \SB2_1_6/i0[8] ), .A3(\SB2_1_6/i3[0] ), .ZN(
        \SB2_1_6/Component_Function_3/NAND4_in[3] ) );
  NAND2_X1 \SB2_1_27/Component_Function_0/N1  ( .A1(\SB2_1_27/i0[10] ), .A2(
        \SB2_1_27/i0[9] ), .ZN(\SB2_1_27/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 U1319 ( .A1(n2745), .A2(\SB2_1_8/i0[10] ), .ZN(n4014) );
  NAND3_X1 \SB2_1_27/Component_Function_4/N4  ( .A1(\SB2_1_27/i1[9] ), .A2(
        \SB2_1_27/i1_5 ), .A3(\SB2_1_27/i0_4 ), .ZN(
        \SB2_1_27/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_3/Component_Function_2/N2  ( .A1(\SB2_1_3/i0_3 ), .A2(
        \SB2_1_3/i0[10] ), .A3(\SB2_1_3/i0[6] ), .ZN(
        \SB2_1_3/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_18/Component_Function_1/N3  ( .A1(\SB2_1_18/i1_5 ), .A2(
        \SB1_1_22/buf_output[1] ), .A3(\SB2_1_18/i0[9] ), .ZN(
        \SB2_1_18/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_1_4/Component_Function_1/N1  ( .A1(\SB2_1_4/i0_3 ), .A2(n3660), 
        .ZN(\SB2_1_4/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U10817 ( .A1(\SB2_1_25/i0[10] ), .A2(\SB2_1_25/i1_5 ), .A3(
        \SB2_1_25/i1[9] ), .ZN(n4517) );
  NAND3_X1 \SB2_1_12/Component_Function_4/N4  ( .A1(\SB2_1_12/i1[9] ), .A2(
        \SB2_1_12/i1_5 ), .A3(\SB2_1_12/i0_4 ), .ZN(
        \SB2_1_12/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U6586 ( .A1(n5790), .A2(\SB2_1_7/i1[9] ), .A3(\SB2_1_7/i1_5 ), .ZN(
        n2545) );
  NAND3_X1 U949 ( .A1(\SB2_1_6/i1[9] ), .A2(\SB2_1_6/i0_3 ), .A3(
        \SB2_1_6/i0[6] ), .ZN(\SB2_1_6/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_25/Component_Function_2/N2  ( .A1(\SB2_1_25/i0_3 ), .A2(
        \SB2_1_25/i0[10] ), .A3(\SB2_1_25/i0[6] ), .ZN(
        \SB2_1_25/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_1/Component_Function_4/N4  ( .A1(\SB2_1_1/i1[9] ), .A2(
        \SB2_1_1/i1_5 ), .A3(\SB2_1_1/i0_4 ), .ZN(
        \SB2_1_1/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U9752 ( .A1(\SB2_1_11/i0_0 ), .A2(\SB2_1_11/i0_3 ), .A3(n3885), 
        .ZN(n4506) );
  NAND3_X1 U3532 ( .A1(\SB2_1_19/i0_3 ), .A2(\SB2_1_19/i0[10] ), .A3(
        \SB2_1_19/i0[9] ), .ZN(n2472) );
  NAND3_X1 U1704 ( .A1(\SB2_1_20/i0[10] ), .A2(\SB2_1_20/i0_3 ), .A3(
        \SB2_1_20/i0_4 ), .ZN(n890) );
  NAND3_X1 U10849 ( .A1(\SB2_1_8/i0[10] ), .A2(\SB2_1_8/i0_3 ), .A3(
        \SB2_1_8/i0_4 ), .ZN(n4529) );
  NAND3_X1 \SB2_1_11/Component_Function_0/N2  ( .A1(\SB2_1_11/i0[8] ), .A2(
        n3885), .A3(\SB2_1_11/i0[6] ), .ZN(
        \SB2_1_11/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_21/Component_Function_1/N2  ( .A1(\SB2_1_21/i0_3 ), .A2(
        \SB2_1_21/i1_7 ), .A3(\SB2_1_21/i0[8] ), .ZN(
        \SB2_1_21/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U3524 ( .A1(\SB2_1_22/i1[9] ), .A2(\SB2_1_22/i1_5 ), .A3(
        \SB2_1_22/i0_4 ), .ZN(\SB2_1_22/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_19/Component_Function_3/N1  ( .A1(n1396), .A2(
        \SB2_1_19/i0_3 ), .A3(\SB2_1_19/i0[6] ), .ZN(
        \SB2_1_19/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U5582 ( .A1(\SB2_1_2/i0_0 ), .A2(\SB2_1_2/i1_5 ), .A3(
        \SB2_1_2/i0_4 ), .ZN(n1689) );
  NAND3_X1 U7537 ( .A1(\SB2_1_20/i0_0 ), .A2(\SB2_1_20/i1_5 ), .A3(
        \SB2_1_20/i0_4 ), .ZN(\SB2_1_20/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_1_4/Component_Function_2/N2  ( .A1(\SB2_1_4/i0_3 ), .A2(
        \SB2_1_4/i0[10] ), .A3(\SB2_1_4/i0[6] ), .ZN(
        \SB2_1_4/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U7159 ( .A1(n4149), .A2(\SB2_1_19/i0[6] ), .A3(\SB2_1_19/i0[8] ), 
        .ZN(\SB2_1_19/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 U5253 ( .A1(\SB2_1_9/i0[10] ), .A2(\SB2_1_9/i0[9] ), .ZN(n1528) );
  NAND3_X1 \SB2_1_3/Component_Function_3/N2  ( .A1(\SB2_1_3/i0_0 ), .A2(
        \SB2_1_3/i0_3 ), .A3(n5208), .ZN(
        \SB2_1_3/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_15/Component_Function_2/N1  ( .A1(\SB2_1_15/i1_5 ), .A2(
        \SB2_1_15/i0[10] ), .A3(\SB2_1_15/i1[9] ), .ZN(
        \SB2_1_15/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U2503 ( .A1(\SB2_1_19/i0_3 ), .A2(n578), .A3(\SB2_1_19/i0[10] ), 
        .ZN(\SB2_1_19/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB2_1_19/Component_Function_1/N1  ( .A1(\SB2_1_19/i0_3 ), .A2(
        n1396), .ZN(\SB2_1_19/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U1251 ( .A1(\SB2_1_25/i0_3 ), .A2(\SB2_1_25/i0[10] ), .A3(
        \SB2_1_25/i0[9] ), .ZN(\SB2_1_25/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U8618 ( .A1(\SB2_1_30/i1[9] ), .A2(n3690), .A3(\SB2_1_30/i1_5 ), 
        .ZN(\SB2_1_30/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_1_25/Component_Function_4/N2  ( .A1(\SB2_1_25/i3[0] ), .A2(
        \SB2_1_25/i0_0 ), .A3(\SB2_1_25/i1_7 ), .ZN(
        \SB2_1_25/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U4886 ( .A1(n3690), .A2(\SB2_1_30/i0_3 ), .A3(\SB2_1_30/i0[6] ), 
        .ZN(\SB2_1_30/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_1_28/Component_Function_4/N4  ( .A1(\SB2_1_28/i1[9] ), .A2(
        \SB2_1_28/i1_5 ), .A3(\SB2_1_28/i0_4 ), .ZN(
        \SB2_1_28/Component_Function_4/NAND4_in[3] ) );
  INV_X1 \SB1_2_16/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[90] ), .ZN(
        \SB1_2_16/i3[0] ) );
  INV_X1 \SB1_2_28/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[18] ), .ZN(
        \SB1_2_28/i3[0] ) );
  INV_X1 \SB1_2_5/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[156] ), .ZN(
        \SB1_2_5/i3[0] ) );
  INV_X1 U3550 ( .I(\MC_ARK_ARC_1_1/buf_output[162] ), .ZN(\SB1_2_4/i3[0] ) );
  CLKBUF_X2 \SB1_2_26/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[30] ), .Z(
        \SB1_2_26/i0[9] ) );
  INV_X1 \SB1_2_15/INV_5  ( .I(n5500), .ZN(\SB1_2_15/i1_5 ) );
  NAND3_X1 U6373 ( .A1(\SB1_2_15/i0_0 ), .A2(\SB1_2_15/i0[8] ), .A3(
        \SB1_2_15/i0[9] ), .ZN(n2047) );
  NOR2_X1 U5788 ( .A1(\SB1_2_26/i0[9] ), .A2(\RI1[2][35] ), .ZN(n3192) );
  INV_X1 \SB1_2_3/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[168] ), .ZN(
        \SB1_2_3/i3[0] ) );
  NAND3_X1 U9636 ( .A1(\SB1_2_5/i0_0 ), .A2(\SB1_2_5/i0[9] ), .A3(
        \SB1_2_5/i0[8] ), .ZN(\SB1_2_5/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U10787 ( .A1(\SB1_2_2/i0_0 ), .A2(\SB1_2_2/i0[8] ), .A3(
        \SB1_2_2/i0[9] ), .ZN(n4498) );
  NAND3_X1 \SB1_2_0/Component_Function_4/N2  ( .A1(\SB1_2_0/i3[0] ), .A2(
        \SB1_2_0/i0_0 ), .A3(\SB1_2_0/i1_7 ), .ZN(
        \SB1_2_0/Component_Function_4/NAND4_in[1] ) );
  INV_X1 \SB1_2_17/INV_5  ( .I(\MC_ARK_ARC_1_1/buf_output[89] ), .ZN(
        \SB1_2_17/i1_5 ) );
  BUF_X2 \SB1_2_23/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[48] ), .Z(
        \SB1_2_23/i0[9] ) );
  NAND3_X1 \SB1_2_5/Component_Function_4/N3  ( .A1(\SB1_2_5/i0[9] ), .A2(
        \SB1_2_5/i0[10] ), .A3(\SB1_2_5/i0_3 ), .ZN(
        \SB1_2_5/Component_Function_4/NAND4_in[2] ) );
  CLKBUF_X2 U2049 ( .I(\MC_ARK_ARC_1_1/buf_output[13] ), .Z(\SB1_2_29/i0[6] )
         );
  INV_X1 \SB1_2_8/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[138] ), .ZN(
        \SB1_2_8/i3[0] ) );
  INV_X1 \SB1_2_24/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[42] ), .ZN(
        \SB1_2_24/i3[0] ) );
  INV_X1 \SB1_2_25/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[36] ), .ZN(
        \SB1_2_25/i3[0] ) );
  INV_X1 U1162 ( .I(\MC_ARK_ARC_1_1/buf_output[61] ), .ZN(\SB1_2_21/i1_7 ) );
  INV_X1 U4717 ( .I(\MC_ARK_ARC_1_1/buf_output[37] ), .ZN(\SB1_2_25/i1_7 ) );
  INV_X1 \SB1_2_23/INV_1  ( .I(\MC_ARK_ARC_1_1/buf_output[49] ), .ZN(
        \SB1_2_23/i1_7 ) );
  BUF_X2 \SB1_2_20/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[67] ), .Z(
        \SB1_2_20/i0[6] ) );
  INV_X1 \SB1_2_12/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[114] ), .ZN(
        \SB1_2_12/i3[0] ) );
  INV_X1 \SB1_2_18/INV_0  ( .I(\MC_ARK_ARC_1_1/buf_output[78] ), .ZN(
        \SB1_2_18/i3[0] ) );
  BUF_X2 \SB1_2_6/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[151] ), .Z(
        \SB1_2_6/i0[6] ) );
  BUF_X2 \SB1_2_25/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[37] ), .Z(
        \SB1_2_25/i0[6] ) );
  NAND3_X1 U6171 ( .A1(\SB1_2_0/i0_4 ), .A2(\SB1_2_0/i1[9] ), .A3(
        \SB1_2_0/i1_5 ), .ZN(n1949) );
  BUF_X2 \SB1_2_2/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[175] ), .Z(
        \SB1_2_2/i0[6] ) );
  BUF_X2 U8860 ( .I(\MC_ARK_ARC_1_1/buf_output[72] ), .Z(\SB1_2_19/i0[9] ) );
  BUF_X2 \SB1_2_9/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[132] ), .Z(
        \SB1_2_9/i0[9] ) );
  BUF_X2 \SB1_2_5/BUF_1  ( .I(\MC_ARK_ARC_1_1/buf_output[157] ), .Z(
        \SB1_2_5/i0[6] ) );
  INV_X1 \SB1_2_1/INV_5  ( .I(\MC_ARK_ARC_1_1/buf_output[185] ), .ZN(
        \SB1_2_1/i1_5 ) );
  INV_X1 U3539 ( .I(\MC_ARK_ARC_1_1/buf_output[29] ), .ZN(\SB1_2_27/i1_5 ) );
  INV_X1 \SB1_2_22/INV_1  ( .I(\MC_ARK_ARC_1_1/buf_output[55] ), .ZN(
        \SB1_2_22/i1_7 ) );
  BUF_X2 \SB1_2_22/BUF_0  ( .I(\MC_ARK_ARC_1_1/buf_output[54] ), .Z(
        \SB1_2_22/i0[9] ) );
  NAND3_X1 U1221 ( .A1(\SB1_2_26/i0[8] ), .A2(\SB1_2_26/i0[9] ), .A3(
        \RI1[2][35] ), .ZN(\SB1_2_26/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_25/Component_Function_2/N3  ( .A1(\SB1_2_25/i0_3 ), .A2(
        \SB1_2_25/i0[8] ), .A3(\SB1_2_25/i0[9] ), .ZN(
        \SB1_2_25/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2065 ( .A1(\SB1_2_31/i0[9] ), .A2(\SB1_2_31/i0[10] ), .A3(
        \SB1_2_31/i0_3 ), .ZN(\SB1_2_31/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U4925 ( .A1(\SB1_2_3/i1[9] ), .A2(\SB1_2_3/i0_3 ), .A3(
        \SB1_2_3/i0[6] ), .ZN(\SB1_2_3/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U877 ( .A1(\SB1_2_11/i0_0 ), .A2(\SB1_2_11/i1_5 ), .A3(
        \SB1_2_11/i0_4 ), .ZN(n2843) );
  NAND3_X1 U1769 ( .A1(\SB1_2_31/i0[9] ), .A2(\SB1_2_31/i0_0 ), .A3(
        \SB1_2_31/i0[8] ), .ZN(n4474) );
  NAND3_X1 U924 ( .A1(\SB1_2_18/i0[10] ), .A2(\SB1_2_18/i1[9] ), .A3(
        \SB1_2_18/i1_7 ), .ZN(\SB1_2_18/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U1159 ( .A1(\RI1[2][47] ), .A2(\SB1_2_24/i1[9] ), .A3(
        \SB1_2_24/i0_4 ), .ZN(\SB1_2_24/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_8/Component_Function_2/N3  ( .A1(\SB1_2_8/i0_3 ), .A2(
        \SB1_2_8/i0[8] ), .A3(\SB1_2_8/i0[9] ), .ZN(
        \SB1_2_8/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U8822 ( .A1(\SB1_2_19/i0_3 ), .A2(\SB1_2_19/i0[8] ), .A3(
        \SB1_2_19/i1_7 ), .ZN(\SB1_2_19/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U8909 ( .A1(\SB1_2_6/i1[9] ), .A2(\SB1_2_6/i1_7 ), .A3(
        \SB1_2_6/i0[10] ), .ZN(\SB1_2_6/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U1211 ( .A1(\SB1_2_7/i0[10] ), .A2(\SB1_2_7/i0_3 ), .A3(
        \SB1_2_7/i0[9] ), .ZN(n3546) );
  NAND2_X1 \SB1_2_25/Component_Function_1/N1  ( .A1(\SB1_2_25/i0_3 ), .A2(
        \SB1_2_25/i1[9] ), .ZN(\SB1_2_25/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_27/Component_Function_3/N4  ( .A1(\SB1_2_27/i1_5 ), .A2(
        \SB1_2_27/i0[8] ), .A3(\SB1_2_27/i3[0] ), .ZN(
        \SB1_2_27/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_5/Component_Function_5/N2  ( .A1(\SB1_2_5/i0_0 ), .A2(
        \SB1_2_5/i0[6] ), .A3(\SB1_2_5/i0[10] ), .ZN(
        \SB1_2_5/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_23/Component_Function_2/N1  ( .A1(\SB1_2_23/i1_5 ), .A2(
        \SB1_2_23/i0[10] ), .A3(\SB1_2_23/i1[9] ), .ZN(
        \SB1_2_23/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_0/Component_Function_2/N1  ( .A1(\SB1_2_0/i1_5 ), .A2(
        \SB1_2_0/i0[10] ), .A3(\SB1_2_0/i1[9] ), .ZN(
        \SB1_2_0/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U898 ( .A1(\SB1_2_22/i1_5 ), .A2(\SB1_2_22/i0_4 ), .A3(
        \SB1_2_22/i1[9] ), .ZN(\SB1_2_22/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U903 ( .A1(\SB1_2_17/i0[10] ), .A2(\SB1_2_17/i0_3 ), .A3(
        \SB1_2_17/i0[6] ), .ZN(n1452) );
  NAND3_X1 \SB1_2_4/Component_Function_0/N2  ( .A1(\SB1_2_4/i0[8] ), .A2(
        \SB1_2_4/i0[7] ), .A3(\SB1_2_4/i0[6] ), .ZN(
        \SB1_2_4/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U1235 ( .A1(\SB1_2_6/i0[8] ), .A2(\SB1_2_6/i3[0] ), .A3(
        \SB1_2_6/i1_5 ), .ZN(n4559) );
  NAND3_X1 \SB1_2_0/Component_Function_0/N2  ( .A1(\SB1_2_0/i0[8] ), .A2(
        \SB1_2_0/i0[7] ), .A3(\SB1_2_0/i0[6] ), .ZN(
        \SB1_2_0/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_24/Component_Function_4/N2  ( .A1(\SB1_2_24/i3[0] ), .A2(
        \SB1_2_24/i0_0 ), .A3(\SB1_2_24/i1_7 ), .ZN(
        \SB1_2_24/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U7314 ( .A1(\SB1_2_2/i0_0 ), .A2(\SB1_2_2/i0_3 ), .A3(
        \SB1_2_2/i0[7] ), .ZN(n2647) );
  NAND3_X1 U7225 ( .A1(\SB1_2_1/i0[6] ), .A2(\SB1_2_1/i0[9] ), .A3(
        \SB1_2_1/i1_5 ), .ZN(n3404) );
  NAND3_X1 \SB1_2_1/Component_Function_0/N3  ( .A1(\SB1_2_1/i0[10] ), .A2(
        \SB1_2_1/i0_4 ), .A3(\SB1_2_1/i0_3 ), .ZN(
        \SB1_2_1/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U5716 ( .A1(\SB1_2_21/i0_0 ), .A2(\SB1_2_21/i1_7 ), .A3(
        \SB1_2_21/i3[0] ), .ZN(n1751) );
  NAND3_X1 U1165 ( .A1(\SB1_2_29/i0[8] ), .A2(\SB1_2_29/i1_7 ), .A3(
        \SB1_2_29/i0_4 ), .ZN(n4548) );
  NAND3_X1 U7050 ( .A1(\SB1_2_2/i0_0 ), .A2(\SB1_2_2/i1_5 ), .A3(
        \SB1_2_2/i0_4 ), .ZN(\SB1_2_2/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U1584 ( .A1(\SB1_2_5/i1[9] ), .A2(\SB1_2_5/i0_4 ), .A3(
        \SB1_2_5/i0_3 ), .ZN(\SB1_2_5/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_24/Component_Function_0/N2  ( .A1(\SB1_2_24/i0[8] ), .A2(
        \SB1_2_24/i0[7] ), .A3(\SB1_2_24/i0[6] ), .ZN(
        \SB1_2_24/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U1835 ( .A1(\SB1_2_12/i0[6] ), .A2(\SB1_2_12/i0[9] ), .A3(
        \SB1_2_12/i1_5 ), .ZN(n940) );
  NAND2_X1 U6893 ( .A1(\SB1_2_10/i0_0 ), .A2(\SB1_2_10/i3[0] ), .ZN(n3348) );
  NAND3_X1 \SB1_2_23/Component_Function_1/N3  ( .A1(\SB1_2_23/i1_5 ), .A2(
        \SB1_2_23/i0[6] ), .A3(\SB1_2_23/i0[9] ), .ZN(
        \SB1_2_23/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB1_2_2/Component_Function_5/N1  ( .A1(\SB1_2_2/i0_0 ), .A2(
        \SB1_2_2/i3[0] ), .ZN(\SB1_2_2/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB1_2_25/Component_Function_5/N1  ( .A1(\SB1_2_25/i0_0 ), .A2(
        \SB1_2_25/i3[0] ), .ZN(\SB1_2_25/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB1_2_14/Component_Function_5/N1  ( .A1(\SB1_2_14/i0_0 ), .A2(
        \SB1_2_14/i3[0] ), .ZN(\SB1_2_14/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_9/Component_Function_2/N3  ( .A1(\SB1_2_9/i0_3 ), .A2(
        \SB1_2_9/i0[8] ), .A3(\SB1_2_9/i0[9] ), .ZN(
        \SB1_2_9/Component_Function_2/NAND4_in[2] ) );
  NAND2_X1 \SB1_2_22/Component_Function_5/N1  ( .A1(\SB1_2_22/i0_0 ), .A2(
        \SB1_2_22/i3[0] ), .ZN(\SB1_2_22/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_21/Component_Function_1/N3  ( .A1(\SB1_2_21/i1_5 ), .A2(
        \SB1_2_21/i0[6] ), .A3(\SB1_2_21/i0[9] ), .ZN(
        \SB1_2_21/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB1_2_6/Component_Function_5/N1  ( .A1(\SB1_2_6/i0_0 ), .A2(
        \SB1_2_6/i3[0] ), .ZN(\SB1_2_6/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_10/Component_Function_5/N4  ( .A1(\SB1_2_10/i0[9] ), .A2(
        \SB1_2_10/i0[6] ), .A3(\SB1_2_10/i0_4 ), .ZN(
        \SB1_2_10/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 U5541 ( .A1(\SB1_2_26/i0_0 ), .A2(\SB1_2_26/i3[0] ), .ZN(
        \SB1_2_26/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U11077 ( .A1(\SB1_2_2/i0[8] ), .A2(\SB1_2_2/i0_3 ), .A3(
        \SB1_2_2/i0[9] ), .ZN(\SB1_2_2/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U7064 ( .A1(\SB1_2_3/i0_0 ), .A2(\SB1_2_3/i1_5 ), .A3(
        \SB1_2_3/i0_4 ), .ZN(\SB1_2_3/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U914 ( .A1(\SB1_2_15/i0_3 ), .A2(\SB1_2_15/i0[8] ), .A3(
        \SB1_2_15/i0[9] ), .ZN(\SB1_2_15/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U5032 ( .A1(\SB1_2_14/i0[6] ), .A2(\SB1_2_14/i0[9] ), .A3(
        \SB1_2_14/i0_4 ), .ZN(n1427) );
  NAND3_X1 U1409 ( .A1(\SB1_2_27/i0[9] ), .A2(\SB1_2_27/i0[10] ), .A3(
        \SB1_2_27/i0_3 ), .ZN(\SB1_2_27/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1183 ( .A1(\SB1_2_8/i0[10] ), .A2(\SB1_2_8/i1[9] ), .A3(
        \SB1_2_8/i1_7 ), .ZN(n2796) );
  NAND3_X1 U9727 ( .A1(\SB1_2_30/i0[9] ), .A2(\SB1_2_30/i0_4 ), .A3(
        \SB1_2_30/i0[6] ), .ZN(n3981) );
  NAND3_X1 U8586 ( .A1(\SB1_2_3/i1[9] ), .A2(\SB1_2_3/i1_5 ), .A3(
        \SB1_2_3/i0_4 ), .ZN(\SB1_2_3/Component_Function_4/NAND4_in[3] ) );
  NAND2_X1 \SB1_2_0/Component_Function_5/N1  ( .A1(\SB1_2_0/i0_0 ), .A2(
        \SB1_2_0/i3[0] ), .ZN(\SB1_2_0/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U3593 ( .A1(\SB1_2_26/i0[8] ), .A2(\SB1_2_26/i0_4 ), .A3(
        \SB1_2_26/i1_7 ), .ZN(n4531) );
  NAND3_X1 U11035 ( .A1(\SB1_2_3/i0[9] ), .A2(\SB1_2_3/i0[6] ), .A3(
        \SB1_2_3/i0_4 ), .ZN(n4644) );
  NAND3_X1 U5476 ( .A1(\SB1_2_30/i0_4 ), .A2(\SB1_2_30/i1[9] ), .A3(
        \SB1_2_30/i1_5 ), .ZN(n1639) );
  NAND3_X1 \SB1_2_21/Component_Function_4/N4  ( .A1(\SB1_2_21/i1[9] ), .A2(
        \SB1_2_21/i1_5 ), .A3(\SB1_2_21/i0_4 ), .ZN(
        \SB1_2_21/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_1/Component_Function_2/N4  ( .A1(\SB1_2_1/i1_5 ), .A2(
        \SB1_2_1/i0_0 ), .A3(\SB1_2_1/i0_4 ), .ZN(
        \SB1_2_1/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_18/Component_Function_1/N3  ( .A1(\SB1_2_18/i1_5 ), .A2(
        \SB1_2_18/i0[6] ), .A3(\SB1_2_18/i0[9] ), .ZN(
        \SB1_2_18/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_27/Component_Function_0/N3  ( .A1(\SB1_2_27/i0[10] ), .A2(
        \SB1_2_27/i0_4 ), .A3(\SB1_2_27/i0_3 ), .ZN(
        \SB1_2_27/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U7966 ( .A1(\SB1_2_13/i0_3 ), .A2(\SB1_2_13/i0[10] ), .A3(
        \SB1_2_13/i0[9] ), .ZN(n3510) );
  NAND3_X1 U10880 ( .A1(\SB1_2_6/i0[8] ), .A2(\SB1_2_6/i0_3 ), .A3(
        \SB1_2_6/i0[9] ), .ZN(n4552) );
  NAND2_X1 \SB1_2_2/Component_Function_0/N1  ( .A1(\SB1_2_2/i0[10] ), .A2(
        \SB1_2_2/i0[9] ), .ZN(\SB1_2_2/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 U2076 ( .A1(\SB1_2_13/i0[10] ), .A2(\SB1_2_13/i0[9] ), .ZN(
        \SB1_2_13/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 U6040 ( .A1(\SB1_2_2/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_2_2/Component_Function_4/NAND4_in[2] ), .ZN(n1894) );
  NAND3_X1 \SB1_2_13/Component_Function_4/N4  ( .A1(\SB1_2_13/i1[9] ), .A2(
        \SB1_2_13/i1_5 ), .A3(\SB1_2_13/i0_4 ), .ZN(
        \SB1_2_13/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_22/Component_Function_4/N3  ( .A1(\SB1_2_22/i0[9] ), .A2(
        \SB1_2_22/i0[10] ), .A3(\SB1_2_22/i0_3 ), .ZN(
        \SB1_2_22/Component_Function_4/NAND4_in[2] ) );
  NAND2_X1 U5607 ( .A1(\SB1_2_14/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_14/Component_Function_4/NAND4_in[2] ), .ZN(n1707) );
  NAND3_X1 U3569 ( .A1(\SB1_2_28/i1_7 ), .A2(\SB1_2_28/i0[8] ), .A3(
        \SB1_2_28/i0_4 ), .ZN(\SB1_2_28/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_25/Component_Function_0/N3  ( .A1(\SB1_2_25/i0[10] ), .A2(
        \SB1_2_25/i0_4 ), .A3(\SB1_2_25/i0_3 ), .ZN(
        \SB1_2_25/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_17/Component_Function_2/N3  ( .A1(\SB1_2_17/i0_3 ), .A2(
        \SB1_2_17/i0[8] ), .A3(\SB1_2_17/i0[9] ), .ZN(
        \SB1_2_17/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_23/Component_Function_5/N2  ( .A1(\SB1_2_23/i0_0 ), .A2(
        \SB1_2_23/i0[6] ), .A3(\SB1_2_23/i0[10] ), .ZN(
        \SB1_2_23/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U9724 ( .A1(\SB1_2_17/i0[8] ), .A2(\SB1_2_17/i0_4 ), .A3(
        \SB1_2_17/i1_7 ), .ZN(n3979) );
  NAND2_X1 U9795 ( .A1(\SB1_2_5/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_5/Component_Function_4/NAND4_in[2] ), .ZN(n4011) );
  NAND2_X1 U9796 ( .A1(\SB1_2_5/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_2_5/Component_Function_4/NAND4_in[1] ), .ZN(n4012) );
  NAND2_X1 U3270 ( .A1(\SB1_2_2/Component_Function_4/NAND4_in[1] ), .A2(n4498), 
        .ZN(n2168) );
  NAND3_X1 U7533 ( .A1(\SB1_2_0/i0_0 ), .A2(\SB1_2_0/i1_5 ), .A3(
        \SB1_2_0/i0_4 ), .ZN(n2644) );
  NAND3_X1 U7236 ( .A1(\SB1_2_1/i1[9] ), .A2(\SB1_2_1/i0_3 ), .A3(
        \SB1_2_1/i0[6] ), .ZN(\SB1_2_1/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U10243 ( .A1(\SB1_2_31/i0_0 ), .A2(\SB1_2_31/i0_4 ), .A3(
        \SB1_2_31/i1_5 ), .ZN(\SB1_2_31/Component_Function_2/NAND4_in[3] ) );
  NAND2_X1 U1879 ( .A1(\SB1_2_16/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_2_16/Component_Function_4/NAND4_in[2] ), .ZN(n1659) );
  NAND3_X1 U10567 ( .A1(\SB1_2_7/i0[10] ), .A2(\SB1_2_7/i0[6] ), .A3(
        \SB1_2_7/i0_3 ), .ZN(\SB1_2_7/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_1/Component_Function_3/N2  ( .A1(\SB1_2_1/i0_0 ), .A2(
        \SB1_2_1/i0_3 ), .A3(\SB1_2_1/i0_4 ), .ZN(
        \SB1_2_1/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_3/Component_Function_3/N2  ( .A1(\SB1_2_3/i0_0 ), .A2(
        \SB1_2_3/i0_3 ), .A3(\SB1_2_3/i0_4 ), .ZN(
        \SB1_2_3/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_1/Component_Function_5/N3  ( .A1(\SB1_2_1/i1[9] ), .A2(
        \SB1_2_1/i0_4 ), .A3(\SB1_2_1/i0_3 ), .ZN(
        \SB1_2_1/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U3591 ( .A1(\SB1_2_8/i0[10] ), .A2(\SB1_2_8/i0[9] ), .A3(
        \SB1_2_8/i0_3 ), .ZN(n2294) );
  NAND3_X1 U922 ( .A1(\SB1_2_31/i0[8] ), .A2(\SB1_2_31/i3[0] ), .A3(
        \SB1_2_31/i1_5 ), .ZN(n2689) );
  NAND3_X1 U8841 ( .A1(\RI1[2][47] ), .A2(\SB1_2_24/i0[8] ), .A3(
        \SB1_2_24/i0[9] ), .ZN(\SB1_2_24/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U11150 ( .A1(\SB1_2_23/i0[8] ), .A2(\SB1_2_23/i3[0] ), .A3(
        \SB1_2_23/i1_5 ), .ZN(n4712) );
  NAND2_X1 U858 ( .A1(\SB1_2_23/i0_3 ), .A2(\SB1_2_23/i1[9] ), .ZN(n1594) );
  NAND3_X1 \SB1_2_23/Component_Function_0/N3  ( .A1(\SB1_2_23/i0[10] ), .A2(
        \SB1_2_23/i0_4 ), .A3(\SB1_2_23/i0_3 ), .ZN(
        \SB1_2_23/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB1_2_11/Component_Function_5/N1  ( .A1(\SB1_2_11/i0_0 ), .A2(
        \SB1_2_11/i3[0] ), .ZN(\SB1_2_11/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U909 ( .A1(\SB1_2_10/i0_0 ), .A2(\SB1_2_10/i0[9] ), .A3(
        \SB1_2_10/i0[8] ), .ZN(n2457) );
  NAND3_X1 U10829 ( .A1(\SB1_2_30/i0_0 ), .A2(\SB1_2_30/i0_4 ), .A3(
        \SB1_2_30/i1_5 ), .ZN(n4521) );
  NAND3_X1 \SB1_2_21/Component_Function_4/N1  ( .A1(\SB1_2_21/i0[9] ), .A2(
        \SB1_2_21/i0_0 ), .A3(\SB1_2_21/i0[8] ), .ZN(
        \SB1_2_21/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_5/Component_Function_2/N3  ( .A1(\SB1_2_5/i0_3 ), .A2(
        \SB1_2_5/i0[8] ), .A3(\SB1_2_5/i0[9] ), .ZN(
        \SB1_2_5/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U9399 ( .A1(\SB1_2_18/i0[6] ), .A2(\SB1_2_18/i0_3 ), .A3(
        \SB1_2_18/i1[9] ), .ZN(n3828) );
  NAND3_X1 U5300 ( .A1(\SB1_2_30/i0[8] ), .A2(\SB1_2_30/i3[0] ), .A3(
        \SB1_2_30/i1_5 ), .ZN(n1547) );
  NAND3_X1 \SB1_2_24/Component_Function_1/N3  ( .A1(\SB1_2_24/i1_5 ), .A2(
        \SB1_2_24/i0[6] ), .A3(\SB1_2_24/i0[9] ), .ZN(
        \SB1_2_24/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U9334 ( .A1(\SB1_2_10/i0_0 ), .A2(\SB1_2_10/i1_7 ), .A3(
        \SB1_2_10/i3[0] ), .ZN(n4477) );
  NAND3_X1 U6773 ( .A1(\SB1_2_21/i0_0 ), .A2(\SB1_2_21/i1_5 ), .A3(
        \SB1_2_21/i0_4 ), .ZN(\SB1_2_21/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB1_2_28/Component_Function_2/N3  ( .A1(\SB1_2_28/i0_3 ), .A2(
        \SB1_2_28/i0[8] ), .A3(\SB1_2_28/i0[9] ), .ZN(
        \SB1_2_28/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1371 ( .A1(\SB1_2_28/i0[10] ), .A2(\SB1_2_28/i0_3 ), .A3(
        \SB1_2_28/i0[6] ), .ZN(\SB1_2_28/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_3/Component_Function_4/N3  ( .A1(\SB1_2_3/i0[9] ), .A2(
        \SB1_2_3/i0[10] ), .A3(\SB1_2_3/i0_3 ), .ZN(
        \SB1_2_3/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U7293 ( .A1(\SB1_2_1/i0_0 ), .A2(\SB1_2_1/i0[6] ), .A3(
        \SB1_2_1/i0[10] ), .ZN(\SB1_2_1/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 \SB1_2_23/Component_Function_3/N3  ( .A1(\SB1_2_23/i1[9] ), .A2(
        \SB1_2_23/i1_7 ), .A3(\SB1_2_23/i0[10] ), .ZN(
        \SB1_2_23/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U5301 ( .A1(\RI1[2][47] ), .A2(\SB1_2_24/i1[9] ), .A3(
        \SB1_2_24/i0[6] ), .ZN(\SB1_2_24/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U5838 ( .A1(\SB1_2_25/i0_0 ), .A2(\SB1_2_25/i0[8] ), .A3(
        \SB1_2_25/i0[9] ), .ZN(\SB1_2_25/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U8625 ( .A1(\RI1[2][47] ), .A2(\SB1_2_24/i0[9] ), .A3(
        \SB1_2_24/i0[10] ), .ZN(\SB1_2_24/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U2069 ( .A1(\RI1[2][47] ), .A2(\SB1_2_24/i0[7] ), .A3(
        \SB1_2_24/i0_0 ), .ZN(n2844) );
  NAND3_X1 U3931 ( .A1(\SB1_2_9/i0[8] ), .A2(\SB1_2_9/i3[0] ), .A3(
        \SB1_2_9/i1_5 ), .ZN(n2923) );
  NAND2_X1 \SB1_2_14/Component_Function_0/N1  ( .A1(\SB1_2_14/i0[10] ), .A2(
        \SB1_2_14/i0[9] ), .ZN(\SB1_2_14/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB1_2_13/Component_Function_1/N4  ( .A1(\SB1_2_13/i1_7 ), .A2(
        \SB1_2_13/i0[8] ), .A3(\SB1_2_13/i0_4 ), .ZN(
        \SB1_2_13/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U2066 ( .A1(\SB1_2_13/i1_5 ), .A2(\SB1_2_13/i0[6] ), .A3(
        \SB1_2_13/i0[9] ), .ZN(\SB1_2_13/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_2_9/Component_Function_3/N2  ( .A1(\SB1_2_9/i0_0 ), .A2(
        \SB1_2_9/i0_3 ), .A3(\SB1_2_9/i0_4 ), .ZN(
        \SB1_2_9/Component_Function_3/NAND4_in[1] ) );
  INV_X1 \SB2_2_13/INV_0  ( .I(\SB1_2_18/buf_output[0] ), .ZN(\SB2_2_13/i3[0] ) );
  INV_X1 U3024 ( .I(\SB1_2_13/buf_output[0] ), .ZN(\SB2_2_8/i3[0] ) );
  BUF_X2 \SB2_2_4/BUF_0  ( .I(\SB1_2_9/buf_output[0] ), .Z(\SB2_2_4/i0[9] ) );
  INV_X1 \SB2_2_27/INV_0  ( .I(\SB1_2_0/buf_output[0] ), .ZN(\SB2_2_27/i3[0] )
         );
  CLKBUF_X2 U1085 ( .I(\SB1_2_10/buf_output[1] ), .Z(\SB2_2_6/i0[6] ) );
  BUF_X2 \SB2_2_30/BUF_0  ( .I(\SB1_2_3/buf_output[0] ), .Z(\SB2_2_30/i0[9] )
         );
  BUF_X2 \SB2_2_12/BUF_0  ( .I(\SB1_2_17/buf_output[0] ), .Z(\SB2_2_12/i0[9] )
         );
  CLKBUF_X2 \SB2_2_0/BUF_0  ( .I(\SB1_2_5/buf_output[0] ), .Z(\SB2_2_0/i0[9] )
         );
  INV_X2 U5686 ( .I(n6073), .ZN(\SB1_2_28/buf_output[4] ) );
  INV_X1 U3314 ( .I(\SB1_2_8/buf_output[0] ), .ZN(\SB2_2_3/i3[0] ) );
  INV_X2 U6985 ( .I(n2342), .ZN(\SB1_2_4/buf_output[4] ) );
  INV_X2 U9384 ( .I(\SB2_2_13/i0[7] ), .ZN(n580) );
  INV_X1 \SB2_2_15/INV_1  ( .I(\SB1_2_19/buf_output[1] ), .ZN(\SB2_2_15/i1_7 )
         );
  INV_X1 U9017 ( .I(\SB1_2_26/buf_output[1] ), .ZN(\SB2_2_22/i1_7 ) );
  INV_X1 \SB2_2_21/INV_1  ( .I(\SB1_2_25/buf_output[1] ), .ZN(\SB2_2_21/i1_7 )
         );
  INV_X1 \SB2_2_5/INV_1  ( .I(\SB1_2_9/buf_output[1] ), .ZN(\SB2_2_5/i1_7 ) );
  NAND3_X1 U6326 ( .A1(\SB2_2_0/i0_3 ), .A2(\SB2_2_0/i0_0 ), .A3(
        \SB2_2_0/i0[7] ), .ZN(n3268) );
  NAND3_X1 \SB2_2_19/Component_Function_3/N4  ( .A1(\SB2_2_19/i1_5 ), .A2(
        \SB2_2_19/i0[8] ), .A3(\SB2_2_19/i3[0] ), .ZN(
        \SB2_2_19/Component_Function_3/NAND4_in[3] ) );
  NAND2_X1 \SB2_2_12/Component_Function_5/N1  ( .A1(\SB2_2_12/i0_0 ), .A2(
        \SB2_2_12/i3[0] ), .ZN(\SB2_2_12/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_31/Component_Function_1/N1  ( .A1(\SB2_2_31/i0_3 ), .A2(
        \SB2_2_31/i1[9] ), .ZN(\SB2_2_31/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_19/Component_Function_3/N2  ( .A1(\SB2_2_19/i0_0 ), .A2(
        \SB2_2_19/i0_3 ), .A3(\SB2_2_19/i0_4 ), .ZN(
        \SB2_2_19/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3874 ( .A1(\SB2_2_2/i0_3 ), .A2(\SB2_2_2/i0[10] ), .A3(
        \SB2_2_2/i0[9] ), .ZN(\SB2_2_2/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U6920 ( .A1(\SB2_2_21/i0_3 ), .A2(\SB2_2_21/i1[9] ), .A3(
        \SB2_2_21/i0_4 ), .ZN(\SB2_2_21/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 \SB2_2_6/Component_Function_5/N1  ( .A1(\SB2_2_6/i0_0 ), .A2(
        \SB2_2_6/i3[0] ), .ZN(\SB2_2_6/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_21/Component_Function_5/N1  ( .A1(\SB2_2_21/i0_0 ), .A2(
        \SB2_2_21/i3[0] ), .ZN(\SB2_2_21/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U828 ( .A1(\SB2_2_8/i0[10] ), .A2(\SB2_2_8/i1[9] ), .A3(
        \SB2_2_8/i1_7 ), .ZN(\SB2_2_8/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_18/Component_Function_4/N3  ( .A1(\SB2_2_18/i0[9] ), .A2(
        \SB2_2_18/i0[10] ), .A3(\SB2_2_18/i0_3 ), .ZN(
        \SB2_2_18/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_5/Component_Function_1/N3  ( .A1(\SB2_2_5/i1_5 ), .A2(
        \SB2_2_5/i0[6] ), .A3(\SB2_2_5/i0[9] ), .ZN(
        \SB2_2_5/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_2/Component_Function_4/N1  ( .A1(\SB2_2_2/i0[9] ), .A2(
        \SB2_2_2/i0_0 ), .A3(\SB2_2_2/i0[8] ), .ZN(
        \SB2_2_2/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_26/Component_Function_0/N2  ( .A1(\SB2_2_26/i0[8] ), .A2(
        \SB2_2_26/i0[7] ), .A3(\SB2_2_26/i0[6] ), .ZN(
        \SB2_2_26/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB2_2_31/Component_Function_1/N4  ( .A1(\SB2_2_31/i1_7 ), .A2(
        \SB2_2_31/i0[8] ), .A3(n569), .ZN(
        \SB2_2_31/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U4296 ( .A1(\SB2_2_24/i0_3 ), .A2(\SB2_2_24/i0[8] ), .A3(
        \SB2_2_24/i0[9] ), .ZN(\SB2_2_24/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U11189 ( .A1(\SB2_2_13/i0[10] ), .A2(\SB2_2_13/i0_3 ), .A3(
        \SB2_2_13/i0[9] ), .ZN(n4732) );
  NAND3_X1 U821 ( .A1(\SB2_2_17/i0_3 ), .A2(\SB2_2_17/i0_4 ), .A3(
        \SB2_2_17/i0[10] ), .ZN(n1199) );
  NAND2_X1 \SB2_2_22/Component_Function_0/N1  ( .A1(\SB2_2_22/i0[10] ), .A2(
        \SB2_2_22/i0[9] ), .ZN(\SB2_2_22/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_30/Component_Function_2/N4  ( .A1(\SB2_2_30/i1_5 ), .A2(
        \SB2_2_30/i0_0 ), .A3(n2343), .ZN(
        \SB2_2_30/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U5331 ( .A1(\SB2_2_26/i0[10] ), .A2(\SB2_2_26/i0_3 ), .A3(
        \SB2_2_26/i0_4 ), .ZN(\SB2_2_26/Component_Function_0/NAND4_in[2] ) );
  CLKBUF_X2 \SB2_2_3/BUF_0  ( .I(\SB1_2_8/buf_output[0] ), .Z(\SB2_2_3/i0[9] )
         );
  CLKBUF_X2 \SB2_2_29/BUF_0  ( .I(\SB1_2_2/buf_output[0] ), .Z(
        \SB2_2_29/i0[9] ) );
  INV_X2 U5224 ( .I(\SB2_2_7/i0[7] ), .ZN(\SB1_2_8/buf_output[4] ) );
  INV_X1 \SB2_2_26/INV_0  ( .I(\SB1_2_31/buf_output[0] ), .ZN(\SB2_2_26/i3[0] ) );
  INV_X1 U1630 ( .I(\SB1_2_30/buf_output[1] ), .ZN(\SB2_2_26/i1_7 ) );
  NAND3_X1 U7182 ( .A1(\SB2_2_13/i0_0 ), .A2(\SB2_2_13/i3[0] ), .A3(
        \SB2_2_13/i1_7 ), .ZN(\SB2_2_13/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U846 ( .A1(\SB2_2_23/i0_3 ), .A2(\SB2_2_23/i0[10] ), .A3(
        \SB2_2_23/i0_4 ), .ZN(n2524) );
  NAND3_X1 \SB2_2_7/Component_Function_4/N2  ( .A1(\SB2_2_7/i3[0] ), .A2(
        \SB2_2_7/i0_0 ), .A3(\SB2_2_7/i1_7 ), .ZN(
        \SB2_2_7/Component_Function_4/NAND4_in[1] ) );
  NAND2_X1 U987 ( .A1(\SB2_2_24/i0_0 ), .A2(\SB2_2_24/i3[0] ), .ZN(n3323) );
  NAND3_X1 \SB2_2_12/Component_Function_3/N4  ( .A1(\SB2_2_12/i1_5 ), .A2(
        \SB2_2_12/i0[8] ), .A3(\SB2_2_12/i3[0] ), .ZN(
        \SB2_2_12/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U855 ( .A1(\SB2_2_11/i0[8] ), .A2(\SB2_2_11/i3[0] ), .A3(
        \SB2_2_11/i1_5 ), .ZN(n2451) );
  NAND3_X1 \SB2_2_31/Component_Function_4/N2  ( .A1(\SB2_2_31/i3[0] ), .A2(
        \SB2_2_31/i0_0 ), .A3(\SB2_2_31/i1_7 ), .ZN(
        \SB2_2_31/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U6123 ( .A1(\SB2_2_18/i0_3 ), .A2(\SB2_2_18/i0[8] ), .A3(
        \SB2_2_18/i1_7 ), .ZN(\SB2_2_18/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 \SB2_2_29/Component_Function_5/N1  ( .A1(\SB2_2_29/i0_0 ), .A2(
        \SB2_2_29/i3[0] ), .ZN(\SB2_2_29/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_1/Component_Function_2/N1  ( .A1(\SB2_2_1/i1_5 ), .A2(
        \SB2_2_1/i0[10] ), .A3(\SB2_2_1/i1[9] ), .ZN(
        \SB2_2_1/Component_Function_2/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_30/Component_Function_5/N1  ( .A1(\SB2_2_30/i0_0 ), .A2(
        \SB2_2_30/i3[0] ), .ZN(\SB2_2_30/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U3584 ( .A1(\SB2_2_14/i0[8] ), .A2(n5932), .A3(\SB2_2_14/i1_7 ), 
        .ZN(\SB2_2_14/Component_Function_1/NAND4_in[3] ) );
  INV_X1 \SB2_2_1/INV_1  ( .I(\SB1_2_5/buf_output[1] ), .ZN(\SB2_2_1/i1_7 ) );
  NAND3_X1 \SB2_2_4/Component_Function_4/N4  ( .A1(\SB2_2_4/i1[9] ), .A2(
        \SB2_2_4/i1_5 ), .A3(\SB2_2_4/i0_4 ), .ZN(
        \SB2_2_4/Component_Function_4/NAND4_in[3] ) );
  NAND2_X1 U8633 ( .A1(\SB2_2_2/i0_0 ), .A2(\SB2_2_2/i3[0] ), .ZN(n1469) );
  NAND3_X1 \SB2_2_13/Component_Function_2/N3  ( .A1(\SB2_2_13/i0_3 ), .A2(
        \SB2_2_13/i0[8] ), .A3(\SB2_2_13/i0[9] ), .ZN(
        \SB2_2_13/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U6207 ( .A1(\SB2_2_14/i0[9] ), .A2(\SB2_2_14/i1_5 ), .A3(
        \SB2_2_14/i0[6] ), .ZN(n4452) );
  NAND3_X1 U2638 ( .A1(\SB2_2_29/i0_3 ), .A2(\SB2_2_29/i0[10] ), .A3(n1837), 
        .ZN(\SB2_2_29/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_31/Component_Function_4/N4  ( .A1(\SB2_2_31/i1[9] ), .A2(
        \SB2_2_31/i1_5 ), .A3(n569), .ZN(
        \SB2_2_31/Component_Function_4/NAND4_in[3] ) );
  INV_X1 U8254 ( .I(\SB1_2_10/buf_output[1] ), .ZN(\SB2_2_6/i1_7 ) );
  NAND2_X1 \SB2_2_3/Component_Function_5/N1  ( .A1(\SB2_2_3/i0_0 ), .A2(
        \SB2_2_3/i3[0] ), .ZN(\SB2_2_3/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_26/Component_Function_2/N3  ( .A1(\SB2_2_26/i0_3 ), .A2(
        \SB2_2_26/i0[8] ), .A3(\SB2_2_26/i0[9] ), .ZN(
        \SB2_2_26/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U7061 ( .A1(\SB2_2_0/i0[10] ), .A2(\SB2_2_0/i1_5 ), .A3(
        \SB2_2_0/i1[9] ), .ZN(\SB2_2_0/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_26/Component_Function_2/N1  ( .A1(\SB2_2_26/i1_5 ), .A2(
        \SB2_2_26/i0[10] ), .A3(\SB2_2_26/i1[9] ), .ZN(
        \SB2_2_26/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U8398 ( .A1(\SB2_2_0/i1_5 ), .A2(\SB2_2_0/i0_0 ), .A3(
        \SB2_2_0/i0_4 ), .ZN(\SB2_2_0/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U2088 ( .A1(n1394), .A2(\SB2_2_13/i0[6] ), .A3(\SB2_2_13/i0[9] ), 
        .ZN(\SB2_2_13/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U2755 ( .A1(\SB2_2_19/i1[9] ), .A2(\SB2_2_19/i1_5 ), .A3(
        \SB2_2_19/i0_4 ), .ZN(\SB2_2_19/Component_Function_4/NAND4_in[3] ) );
  INV_X1 \SB2_2_20/INV_1  ( .I(\SB1_2_24/buf_output[1] ), .ZN(\SB2_2_20/i1_7 )
         );
  NAND3_X1 \SB2_2_10/Component_Function_4/N1  ( .A1(\SB2_2_10/i0[9] ), .A2(
        \SB2_2_10/i0_0 ), .A3(\SB2_2_10/i0[8] ), .ZN(
        \SB2_2_10/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_13/Component_Function_0/N3  ( .A1(\SB2_2_13/i0[10] ), .A2(
        n580), .A3(\SB2_2_13/i0_3 ), .ZN(
        \SB2_2_13/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U2123 ( .A1(\SB2_2_6/i0[6] ), .A2(\SB2_2_6/i0_3 ), .A3(
        \SB2_2_6/i1[9] ), .ZN(\SB2_2_6/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2635 ( .A1(\SB2_2_29/i0_3 ), .A2(\SB2_2_29/i0[9] ), .A3(
        \SB2_2_29/i0[10] ), .ZN(\SB2_2_29/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U7789 ( .A1(\SB2_2_3/i1[9] ), .A2(\SB1_2_4/buf_output[4] ), .A3(
        \SB2_2_3/i1_5 ), .ZN(n2802) );
  NAND3_X1 U2095 ( .A1(\SB2_2_12/i1[9] ), .A2(\SB2_2_12/i1_5 ), .A3(
        \SB2_2_12/i0_4 ), .ZN(\SB2_2_12/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U1006 ( .A1(n5515), .A2(n4749), .A3(\SB2_2_11/i1_5 ), .ZN(n4626) );
  NAND3_X1 U7187 ( .A1(\SB2_2_17/i0_3 ), .A2(\SB2_2_17/i0[10] ), .A3(
        \SB2_2_17/i0[9] ), .ZN(n1278) );
  NAND3_X1 \SB2_2_2/Component_Function_0/N2  ( .A1(\SB2_2_2/i0[8] ), .A2(
        \SB2_2_2/i0[7] ), .A3(\SB2_2_2/i0[6] ), .ZN(
        \SB2_2_2/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U1810 ( .A1(\SB2_2_20/i0_3 ), .A2(\SB2_2_20/i0_4 ), .A3(
        \SB2_2_20/i1[9] ), .ZN(n1644) );
  NAND3_X1 U3774 ( .A1(\SB2_2_21/i0_3 ), .A2(\SB2_2_21/i0[6] ), .A3(
        \SB2_2_21/i1[9] ), .ZN(\SB2_2_21/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_1/Component_Function_3/N4  ( .A1(\SB2_2_1/i1_5 ), .A2(
        \SB2_2_1/i0[8] ), .A3(\SB2_2_1/i3[0] ), .ZN(
        \SB2_2_1/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_25/Component_Function_0/N2  ( .A1(\SB2_2_25/i0[8] ), .A2(
        \SB2_2_25/i0[7] ), .A3(\SB2_2_25/i0[6] ), .ZN(
        \SB2_2_25/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U5399 ( .A1(\SB2_2_20/i0_3 ), .A2(\SB2_2_20/i0[10] ), .A3(
        \SB2_2_20/i0[9] ), .ZN(n1598) );
  NAND3_X1 U4999 ( .A1(\SB2_2_1/i0[10] ), .A2(\SB2_2_1/i1_7 ), .A3(
        \SB2_2_1/i1[9] ), .ZN(\SB2_2_1/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U4133 ( .A1(\SB2_2_19/i1_7 ), .A2(\SB2_2_19/i0[8] ), .A3(
        \SB2_2_19/i0_4 ), .ZN(\SB2_2_19/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_1/Component_Function_1/N4  ( .A1(\SB2_2_1/i1_7 ), .A2(
        \SB2_2_1/i0[8] ), .A3(\SB2_2_1/i0_4 ), .ZN(
        \SB2_2_1/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_20/Component_Function_1/N4  ( .A1(\SB2_2_20/i1_7 ), .A2(
        \SB2_2_20/i0[8] ), .A3(\SB2_2_20/i0_4 ), .ZN(
        \SB2_2_20/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U7895 ( .A1(\SB2_2_10/i0_0 ), .A2(n581), .A3(\SB2_2_10/i1_5 ), .ZN(
        n3495) );
  NAND3_X1 U2405 ( .A1(\SB2_2_9/i0[9] ), .A2(\SB2_2_9/i0_3 ), .A3(
        \SB2_2_9/i0[10] ), .ZN(n639) );
  NAND3_X1 U5080 ( .A1(\SB2_2_27/i1[9] ), .A2(\SB2_2_27/i1_5 ), .A3(
        \SB1_2_28/buf_output[4] ), .ZN(
        \SB2_2_27/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U5926 ( .A1(\SB2_2_7/i3[0] ), .A2(\SB2_2_7/i0[8] ), .A3(
        \SB2_2_7/i1_5 ), .ZN(n3207) );
  NAND3_X1 U843 ( .A1(\SB2_2_29/i0[8] ), .A2(\SB2_2_29/i1_7 ), .A3(n1837), 
        .ZN(\SB2_2_29/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_4/Component_Function_1/N4  ( .A1(\SB2_2_4/i1_7 ), .A2(
        \SB2_2_4/i0[8] ), .A3(\SB2_2_4/i0_4 ), .ZN(
        \SB2_2_4/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_0/Component_Function_4/N4  ( .A1(\SB2_2_0/i1[9] ), .A2(
        \SB2_2_0/i1_5 ), .A3(\SB2_2_0/i0_4 ), .ZN(
        \SB2_2_0/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U6752 ( .A1(\SB2_2_1/i0_4 ), .A2(\SB2_2_1/i1[9] ), .A3(
        \SB2_2_1/i1_5 ), .ZN(n2236) );
  NAND3_X1 U2887 ( .A1(\SB2_2_21/i0[9] ), .A2(\SB2_2_21/i0[8] ), .A3(
        \SB2_2_21/i0_0 ), .ZN(n792) );
  NAND3_X1 U2085 ( .A1(\SB2_2_1/i0[9] ), .A2(\SB2_2_1/i0[6] ), .A3(
        \SB2_2_1/i1_5 ), .ZN(n1649) );
  NAND3_X1 U6086 ( .A1(\SB2_2_15/i0[6] ), .A2(\SB2_2_15/i1_5 ), .A3(
        \SB2_2_15/i0[9] ), .ZN(\SB2_2_15/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_2_27/Component_Function_1/N3  ( .A1(\SB2_2_27/i1_5 ), .A2(
        \SB2_2_27/i0[6] ), .A3(\SB2_2_27/i0[9] ), .ZN(
        \SB2_2_27/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_2_31/Component_Function_5/N1  ( .A1(\SB2_2_31/i0_0 ), .A2(
        \SB2_2_31/i3[0] ), .ZN(\SB2_2_31/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U977 ( .A1(\SB2_2_22/i0[10] ), .A2(\SB2_2_22/i0_0 ), .A3(
        \SB2_2_22/i0[6] ), .ZN(n3353) );
  NAND2_X1 \SB2_2_5/Component_Function_5/N1  ( .A1(\SB2_2_5/i0_0 ), .A2(
        \SB2_2_5/i3[0] ), .ZN(\SB2_2_5/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB2_2_9/Component_Function_1/N1  ( .A1(\SB2_2_9/i0_3 ), .A2(
        \SB2_2_9/i1[9] ), .ZN(\SB2_2_9/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 \SB2_2_11/Component_Function_1/N3  ( .A1(\SB2_2_11/i1_5 ), .A2(
        \SB2_2_11/i0[6] ), .A3(\SB2_2_11/i0[9] ), .ZN(
        \SB2_2_11/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U3128 ( .A1(\SB2_2_28/i0[10] ), .A2(\SB2_2_28/i1[9] ), .A3(
        \SB2_2_28/i1_7 ), .ZN(n874) );
  NAND3_X1 U3173 ( .A1(\SB2_2_20/i0[6] ), .A2(\SB2_2_20/i1_5 ), .A3(
        \SB2_2_20/i0[9] ), .ZN(\SB2_2_20/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U4695 ( .A1(\SB2_2_24/i0_3 ), .A2(\SB2_2_24/i0_0 ), .A3(
        \SB2_2_24/i0_4 ), .ZN(n3032) );
  NAND3_X1 \SB2_2_3/Component_Function_1/N4  ( .A1(\SB2_2_3/i1_7 ), .A2(
        \SB2_2_3/i0[8] ), .A3(\SB1_2_4/buf_output[4] ), .ZN(
        \SB2_2_3/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_2_20/Component_Function_4/N4  ( .A1(\SB2_2_20/i1[9] ), .A2(
        \SB2_2_20/i1_5 ), .A3(\SB2_2_20/i0_4 ), .ZN(
        \SB2_2_20/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U9129 ( .A1(\SB2_2_5/i0[6] ), .A2(\SB2_2_5/i0[10] ), .A3(
        \SB2_2_5/i0_0 ), .ZN(n3717) );
  NAND3_X1 \SB2_2_31/Component_Function_5/N2  ( .A1(\SB2_2_31/i0_0 ), .A2(
        \SB2_2_31/i0[6] ), .A3(\SB2_2_31/i0[10] ), .ZN(
        \SB2_2_31/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1034 ( .A1(\SB2_2_6/i0[10] ), .A2(\SB2_2_6/i0_3 ), .A3(
        \SB2_2_6/i0[9] ), .ZN(n4432) );
  NAND3_X1 U2636 ( .A1(\SB2_2_29/i0[10] ), .A2(\SB2_2_29/i0_3 ), .A3(
        \SB2_2_29/i0[6] ), .ZN(\SB2_2_29/Component_Function_2/NAND4_in[1] ) );
  BUF_X2 U8160 ( .I(\SB2_2_1/buf_output[4] ), .Z(\RI5[2][190] ) );
  BUF_X2 U3251 ( .I(\MC_ARK_ARC_1_2/buf_output[118] ), .Z(\SB1_3_12/i0_4 ) );
  BUF_X2 \SB1_3_26/BUF_1  ( .I(\MC_ARK_ARC_1_2/buf_output[31] ), .Z(
        \SB1_3_26/i0[6] ) );
  BUF_X2 \SB1_3_8/BUF_0  ( .I(\MC_ARK_ARC_1_2/buf_output[138] ), .Z(
        \SB1_3_8/i0[9] ) );
  INV_X1 U4789 ( .I(\MC_ARK_ARC_1_2/buf_output[139] ), .ZN(\SB1_3_8/i1_7 ) );
  NAND3_X1 U5603 ( .A1(\SB1_3_25/i3[0] ), .A2(\SB1_3_25/i0_0 ), .A3(
        \SB1_3_25/i1_7 ), .ZN(n1704) );
  INV_X1 \SB1_3_6/INV_1  ( .I(\MC_ARK_ARC_1_2/buf_output[151] ), .ZN(
        \SB1_3_6/i1_7 ) );
  INV_X1 \SB1_3_28/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[18] ), .ZN(
        \SB1_3_28/i3[0] ) );
  INV_X1 \SB1_3_24/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[42] ), .ZN(
        \SB1_3_24/i3[0] ) );
  INV_X1 U935 ( .I(\MC_ARK_ARC_1_2/buf_output[174] ), .ZN(\SB1_3_2/i3[0] ) );
  INV_X1 \SB1_3_3/INV_1  ( .I(\MC_ARK_ARC_1_2/buf_output[169] ), .ZN(
        \SB1_3_3/i1_7 ) );
  BUF_X2 U4808 ( .I(\MC_ARK_ARC_1_2/buf_output[145] ), .Z(\SB1_3_7/i0[6] ) );
  NAND3_X1 U4331 ( .A1(\SB1_3_11/i0_3 ), .A2(\SB1_3_11/i0[8] ), .A3(
        \SB1_3_11/i1_7 ), .ZN(\SB1_3_11/Component_Function_1/NAND4_in[1] ) );
  INV_X1 \SB1_3_7/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[144] ), .ZN(
        \SB1_3_7/i3[0] ) );
  INV_X1 \SB1_3_5/INV_0  ( .I(\MC_ARK_ARC_1_2/buf_output[156] ), .ZN(
        \SB1_3_5/i3[0] ) );
  NAND3_X1 U8645 ( .A1(\SB1_3_11/i0[9] ), .A2(\SB1_3_11/i0[6] ), .A3(n2908), 
        .ZN(\SB1_3_11/Component_Function_1/NAND4_in[2] ) );
  INV_X1 \SB1_3_2/INV_1  ( .I(\MC_ARK_ARC_1_2/buf_output[175] ), .ZN(
        \SB1_3_2/i1_7 ) );
  BUF_X2 \SB1_3_29/BUF_1  ( .I(\MC_ARK_ARC_1_2/buf_output[13] ), .Z(
        \SB1_3_29/i0[6] ) );
  NAND3_X1 U10928 ( .A1(\SB1_3_24/i0_4 ), .A2(\SB1_3_24/i1_5 ), .A3(
        \SB1_3_24/i0_0 ), .ZN(n4585) );
  NAND3_X1 U2457 ( .A1(\SB1_3_9/i1[9] ), .A2(\SB1_3_9/i0_3 ), .A3(
        \SB1_3_9/i0[6] ), .ZN(\SB1_3_9/Component_Function_3/NAND4_in[0] ) );
  BUF_X2 \SB1_3_20/BUF_0  ( .I(\MC_ARK_ARC_1_2/buf_output[66] ), .Z(
        \SB1_3_20/i0[9] ) );
  CLKBUF_X2 \SB1_3_19/BUF_0  ( .I(\MC_ARK_ARC_1_2/buf_output[72] ), .Z(
        \SB1_3_19/i0[9] ) );
  BUF_X2 U3249 ( .I(\MC_ARK_ARC_1_2/buf_output[73] ), .Z(\SB1_3_19/i0[6] ) );
  BUF_X2 U3248 ( .I(\MC_ARK_ARC_1_2/buf_output[171] ), .Z(\SB1_3_3/i0[10] ) );
  BUF_X2 U2105 ( .I(\MC_ARK_ARC_1_2/buf_output[157] ), .Z(\SB1_3_5/i0[6] ) );
  BUF_X2 U4788 ( .I(\MC_ARK_ARC_1_2/buf_output[139] ), .Z(\SB1_3_8/i0[6] ) );
  INV_X1 U2108 ( .I(\MC_ARK_ARC_1_2/buf_output[0] ), .ZN(\SB1_3_31/i3[0] ) );
  INV_X1 U1657 ( .I(\MC_ARK_ARC_1_2/buf_output[83] ), .ZN(\SB1_3_18/i1_5 ) );
  INV_X1 \SB1_3_2/INV_3  ( .I(n3673), .ZN(\SB1_3_2/i0[8] ) );
  INV_X1 \SB1_3_28/INV_5  ( .I(\MC_ARK_ARC_1_2/buf_output[23] ), .ZN(
        \SB1_3_28/i1_5 ) );
  INV_X1 \SB1_3_25/INV_4  ( .I(\SB1_3_25/i0_4 ), .ZN(\SB1_3_25/i0[7] ) );
  CLKBUF_X2 U810 ( .I(\MC_ARK_ARC_1_2/buf_output[126] ), .Z(\SB1_3_10/i0[9] )
         );
  NAND3_X1 U847 ( .A1(\SB1_3_7/i0_3 ), .A2(\SB1_3_7/i0_0 ), .A3(
        \SB1_3_7/i0[7] ), .ZN(n3805) );
  NAND3_X1 U3648 ( .A1(\SB1_3_1/i0_3 ), .A2(\SB1_3_1/i0_4 ), .A3(
        \SB1_3_1/i1[9] ), .ZN(n1106) );
  NAND3_X1 U2488 ( .A1(\SB1_3_18/i0_0 ), .A2(\SB1_3_18/i0_4 ), .A3(
        \SB1_3_18/i1_5 ), .ZN(n3752) );
  NAND2_X1 U9213 ( .A1(\SB1_3_6/i1[9] ), .A2(\SB1_3_6/i0_3 ), .ZN(n3753) );
  NAND3_X1 \SB1_3_13/Component_Function_1/N4  ( .A1(\SB1_3_13/i1_7 ), .A2(
        \SB1_3_13/i0[8] ), .A3(\SB1_3_13/i0_4 ), .ZN(
        \SB1_3_13/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U1434 ( .A1(\SB1_3_7/i0[9] ), .A2(\SB1_3_7/i0[10] ), .A3(
        \SB1_3_7/i0_3 ), .ZN(\SB1_3_7/Component_Function_4/NAND4_in[2] ) );
  NAND2_X1 \SB1_3_11/Component_Function_5/N1  ( .A1(\SB1_3_11/i0_0 ), .A2(
        \SB1_3_11/i3[0] ), .ZN(\SB1_3_11/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_2/Component_Function_0/N2  ( .A1(\SB1_3_2/i0[8] ), .A2(
        \SB1_3_2/i0[7] ), .A3(\SB1_3_2/i0[6] ), .ZN(
        \SB1_3_2/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_8/Component_Function_0/N3  ( .A1(\SB1_3_8/i0[10] ), .A2(
        \SB1_3_8/i0_4 ), .A3(\SB1_3_8/i0_3 ), .ZN(
        \SB1_3_8/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_30/Component_Function_0/N2  ( .A1(\SB1_3_30/i0[8] ), .A2(
        \SB1_3_30/i0[7] ), .A3(\SB1_3_30/i0[6] ), .ZN(
        \SB1_3_30/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_17/Component_Function_4/N2  ( .A1(\SB1_3_17/i3[0] ), .A2(
        \SB1_3_17/i0_0 ), .A3(\SB1_3_17/i1_7 ), .ZN(
        \SB1_3_17/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U778 ( .A1(\SB1_3_12/i0[8] ), .A2(\SB1_3_12/i1_5 ), .A3(
        \SB1_3_12/i3[0] ), .ZN(\SB1_3_12/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_9/Component_Function_0/N2  ( .A1(\SB1_3_9/i0[8] ), .A2(
        \SB1_3_9/i0[7] ), .A3(\SB1_3_9/i0[6] ), .ZN(
        \SB1_3_9/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U5651 ( .A1(\SB1_3_1/i0[8] ), .A2(\SB1_3_1/i3[0] ), .A3(
        \SB1_3_1/i1_5 ), .ZN(n1730) );
  NAND3_X1 U4421 ( .A1(\SB1_3_5/i1[9] ), .A2(\SB1_3_5/i1_5 ), .A3(
        \SB1_3_5/i0_4 ), .ZN(\SB1_3_5/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U4356 ( .A1(\SB1_3_21/i0[8] ), .A2(\SB1_3_21/i3[0] ), .A3(
        \SB1_3_21/i1_5 ), .ZN(n1350) );
  NAND3_X1 \SB1_3_3/Component_Function_0/N2  ( .A1(\SB1_3_3/i0[8] ), .A2(
        \SB1_3_3/i0[7] ), .A3(\SB1_3_3/i0[6] ), .ZN(
        \SB1_3_3/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U3110 ( .A1(\SB1_3_21/i0_0 ), .A2(\SB1_3_21/i3[0] ), .A3(
        \SB1_3_21/i1_7 ), .ZN(n2109) );
  NAND2_X1 \SB1_3_1/Component_Function_5/N1  ( .A1(\SB1_3_1/i0_0 ), .A2(
        \SB1_3_1/i3[0] ), .ZN(\SB1_3_1/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_30/Component_Function_1/N4  ( .A1(\SB1_3_30/i1_7 ), .A2(
        \SB1_3_30/i0[8] ), .A3(\SB1_3_30/i0_4 ), .ZN(
        \SB1_3_30/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U1673 ( .A1(\SB1_3_2/i0[9] ), .A2(\SB1_3_2/i0[10] ), .A3(
        \SB1_3_2/i0_3 ), .ZN(\SB1_3_2/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U895 ( .A1(\SB1_3_13/i0[6] ), .A2(\SB1_3_13/i1_5 ), .A3(
        \SB1_3_13/i0[9] ), .ZN(\SB1_3_13/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U5185 ( .A1(\SB1_3_24/i0_4 ), .A2(\SB1_3_24/i1_7 ), .A3(
        \SB1_3_24/i0[8] ), .ZN(n1498) );
  NAND3_X1 U1361 ( .A1(\SB1_3_15/i1_5 ), .A2(\SB1_3_15/i0[6] ), .A3(
        \SB1_3_15/i0[9] ), .ZN(\SB1_3_15/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U6932 ( .A1(\SB1_3_5/i0[8] ), .A2(\SB1_3_5/i1_5 ), .A3(
        \SB1_3_5/i3[0] ), .ZN(n2317) );
  NAND3_X1 U772 ( .A1(\SB1_3_10/i0_3 ), .A2(\SB1_3_10/i0[7] ), .A3(
        \SB1_3_10/i0_0 ), .ZN(\SB1_3_10/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2121 ( .A1(\SB1_3_22/i1_5 ), .A2(\SB1_3_22/i0[6] ), .A3(
        \SB1_3_22/i0[9] ), .ZN(\SB1_3_22/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB1_3_3/Component_Function_5/N1  ( .A1(\SB1_3_3/i0_0 ), .A2(
        \SB1_3_3/i3[0] ), .ZN(\SB1_3_3/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 U2485 ( .A1(\SB1_3_18/i0_0 ), .A2(\SB1_3_18/i3[0] ), .ZN(
        \SB1_3_18/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U1464 ( .A1(\SB1_3_27/i0_0 ), .A2(\SB1_3_27/i0[6] ), .A3(
        \SB1_3_27/i0[10] ), .ZN(\SB1_3_27/Component_Function_5/NAND4_in[1] )
         );
  NAND2_X1 \SB1_3_0/Component_Function_5/N1  ( .A1(\SB1_3_0/i0_0 ), .A2(
        \SB1_3_0/i3[0] ), .ZN(\SB1_3_0/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U3647 ( .A1(\SB1_3_5/i0[9] ), .A2(\SB1_3_5/i0[6] ), .A3(
        \SB1_3_5/i1_5 ), .ZN(n2185) );
  NAND3_X1 U11212 ( .A1(\SB1_3_5/i0[10] ), .A2(\SB1_3_5/i1[9] ), .A3(
        \SB1_3_5/i1_7 ), .ZN(\SB1_3_5/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_3/Component_Function_1/N3  ( .A1(\SB1_3_3/i1_5 ), .A2(
        \SB1_3_3/i0[6] ), .A3(\SB1_3_3/i0[9] ), .ZN(
        \SB1_3_3/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_8/Component_Function_1/N3  ( .A1(\SB1_3_8/i1_5 ), .A2(
        \SB1_3_8/i0[6] ), .A3(\SB1_3_8/i0[9] ), .ZN(
        \SB1_3_8/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U2133 ( .A1(\SB1_3_22/i0_0 ), .A2(\SB1_3_22/i1_5 ), .A3(
        \SB1_3_22/i0_4 ), .ZN(n1245) );
  NAND3_X1 U2867 ( .A1(\SB1_3_0/i0_4 ), .A2(\SB1_3_0/i1[9] ), .A3(
        \SB1_3_0/i0_3 ), .ZN(n806) );
  NAND3_X1 U9654 ( .A1(\SB1_3_0/i0[10] ), .A2(\SB1_3_0/i0[9] ), .A3(
        \SB1_3_0/i0_3 ), .ZN(n3945) );
  NAND3_X1 U7201 ( .A1(\SB1_3_2/i1_5 ), .A2(\SB1_3_2/i1[9] ), .A3(
        \SB1_3_2/i0_4 ), .ZN(\SB1_3_2/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_23/Component_Function_4/N4  ( .A1(\SB1_3_23/i1[9] ), .A2(
        \SB1_3_23/i1_5 ), .A3(\SB1_3_23/i0_4 ), .ZN(
        \SB1_3_23/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U8672 ( .A1(\SB1_3_31/i0[9] ), .A2(\SB1_3_31/i0_0 ), .A3(
        \SB1_3_31/i0[8] ), .ZN(\SB1_3_31/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_25/Component_Function_5/N2  ( .A1(\SB1_3_25/i0_0 ), .A2(
        \SB1_3_25/i0[6] ), .A3(\SB1_3_25/i0[10] ), .ZN(
        \SB1_3_25/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U2028 ( .A1(\SB1_3_9/i0[10] ), .A2(\SB1_3_9/i0_3 ), .A3(
        \SB1_3_9/i0[6] ), .ZN(\SB1_3_9/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_3/Component_Function_2/N4  ( .A1(\SB1_3_3/i1_5 ), .A2(
        \SB1_3_3/i0_0 ), .A3(\SB1_3_3/i0_4 ), .ZN(
        \SB1_3_3/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U814 ( .A1(\SB1_3_13/i0_3 ), .A2(\SB1_3_13/i0_0 ), .A3(
        \SB1_3_13/i0_4 ), .ZN(n841) );
  NAND2_X1 \SB1_3_9/Component_Function_0/N1  ( .A1(\SB1_3_9/i0[10] ), .A2(
        \SB1_3_9/i0[9] ), .ZN(\SB1_3_9/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U2118 ( .A1(\SB1_3_25/i0_0 ), .A2(\SB1_3_25/i0_4 ), .A3(
        \SB1_3_25/i1_5 ), .ZN(n1814) );
  NAND3_X1 \SB1_3_5/Component_Function_4/N3  ( .A1(\SB1_3_5/i0[9] ), .A2(
        \SB1_3_5/i0[10] ), .A3(\SB1_3_5/i0_3 ), .ZN(
        \SB1_3_5/Component_Function_4/NAND4_in[2] ) );
  NAND2_X1 U764 ( .A1(\SB1_3_4/i0_0 ), .A2(\SB1_3_4/i3[0] ), .ZN(n2054) );
  NAND3_X1 \SB1_3_9/Component_Function_1/N3  ( .A1(\SB1_3_9/i1_5 ), .A2(
        \SB1_3_9/i0[6] ), .A3(\SB1_3_9/i0[9] ), .ZN(
        \SB1_3_9/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 U3660 ( .A1(\SB1_3_0/i0_3 ), .A2(\SB1_3_0/i1[9] ), .ZN(
        \SB1_3_0/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U7810 ( .A1(\SB1_3_12/i0[6] ), .A2(\SB1_3_12/i0[9] ), .A3(
        \SB1_3_12/i1_5 ), .ZN(\SB1_3_12/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U5174 ( .A1(\SB1_3_24/i0_3 ), .A2(\SB1_3_24/i0[6] ), .A3(
        \SB1_3_24/i1[9] ), .ZN(\SB1_3_24/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2839 ( .A1(\SB1_3_4/i1_5 ), .A2(\SB1_3_4/i0[6] ), .A3(
        \SB1_3_4/i0[9] ), .ZN(\SB1_3_4/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U10375 ( .A1(\SB1_3_26/i0_3 ), .A2(\SB1_3_26/i0_4 ), .A3(
        \SB1_3_26/i1[9] ), .ZN(\SB1_3_26/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U751 ( .A1(\SB1_3_16/i0_4 ), .A2(\SB1_3_16/i0[9] ), .A3(
        \SB1_3_16/i0[6] ), .ZN(n2782) );
  NAND3_X1 U1156 ( .A1(\SB1_3_3/i0_0 ), .A2(\SB1_3_3/i0[6] ), .A3(
        \SB1_3_3/i0[10] ), .ZN(\SB1_3_3/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1219 ( .A1(\SB1_3_26/i0_0 ), .A2(\SB1_3_26/i0[6] ), .A3(
        \SB1_3_26/i0[10] ), .ZN(\SB1_3_26/Component_Function_5/NAND4_in[1] )
         );
  NAND3_X1 U781 ( .A1(\SB1_3_22/i0_0 ), .A2(\SB1_3_22/i0[6] ), .A3(
        \SB1_3_22/i0[10] ), .ZN(\SB1_3_22/Component_Function_5/NAND4_in[1] )
         );
  NAND3_X1 \SB1_3_1/Component_Function_0/N3  ( .A1(\SB1_3_1/i0[10] ), .A2(
        \SB1_3_1/i0_4 ), .A3(\SB1_3_1/i0_3 ), .ZN(
        \SB1_3_1/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 \SB1_3_6/Component_Function_0/N4  ( .A1(\SB1_3_6/i0[7] ), .A2(
        \SB1_3_6/i0_3 ), .A3(\SB1_3_6/i0_0 ), .ZN(
        \SB1_3_6/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 \SB1_3_7/Component_Function_4/N2  ( .A1(\SB1_3_7/i3[0] ), .A2(
        \SB1_3_7/i0_0 ), .A3(\SB1_3_7/i1_7 ), .ZN(
        \SB1_3_7/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 \SB1_3_2/Component_Function_3/N1  ( .A1(\SB1_3_2/i1[9] ), .A2(
        \SB1_3_2/i0_3 ), .A3(\SB1_3_2/i0[6] ), .ZN(
        \SB1_3_2/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U819 ( .A1(\SB1_3_7/i0[6] ), .A2(\SB1_3_7/i0[10] ), .A3(
        \SB1_3_7/i0_3 ), .ZN(\SB1_3_7/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U5342 ( .A1(\SB1_3_2/i0[10] ), .A2(\SB1_3_2/i0_0 ), .A3(
        \SB1_3_2/i0[6] ), .ZN(n1570) );
  NAND2_X1 \SB1_3_17/Component_Function_5/N1  ( .A1(\SB1_3_17/i0_0 ), .A2(
        \SB1_3_17/i3[0] ), .ZN(\SB1_3_17/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U908 ( .A1(\SB1_3_1/i0_0 ), .A2(\SB1_3_1/i0[7] ), .A3(
        \SB1_3_1/i0_3 ), .ZN(n4518) );
  NAND4_X1 U10894 ( .A1(\SB1_3_2/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_3_2/Component_Function_3/NAND4_in[0] ), .A3(n1658), .A4(n4563), 
        .ZN(\SB1_3_2/buf_output[3] ) );
  NAND2_X1 U774 ( .A1(n3949), .A2(\SB1_3_11/Component_Function_2/NAND4_in[0] ), 
        .ZN(n3119) );
  NAND3_X1 \SB1_3_26/Component_Function_3/N1  ( .A1(\SB1_3_26/i1[9] ), .A2(
        \SB1_3_26/i0_3 ), .A3(\SB1_3_26/i0[6] ), .ZN(
        \SB1_3_26/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB1_3_26/Component_Function_3/N2  ( .A1(\SB1_3_26/i0_0 ), .A2(
        \SB1_3_26/i0_3 ), .A3(\SB1_3_26/i0_4 ), .ZN(
        \SB1_3_26/Component_Function_3/NAND4_in[1] ) );
  INV_X1 \SB2_3_1/INV_1  ( .I(\SB1_3_5/buf_output[1] ), .ZN(\SB2_3_1/i1_7 ) );
  INV_X1 U9902 ( .I(\SB1_3_0/buf_output[1] ), .ZN(\SB2_3_28/i1_7 ) );
  CLKBUF_X2 \SB2_3_1/BUF_0  ( .I(\SB1_3_6/buf_output[0] ), .Z(\SB2_3_1/i0[9] )
         );
  CLKBUF_X2 \SB2_3_16/BUF_0  ( .I(\SB1_3_21/buf_output[0] ), .Z(
        \SB2_3_16/i0[9] ) );
  BUF_X2 \SB2_3_20/BUF_0  ( .I(\SB1_3_25/buf_output[0] ), .Z(\SB2_3_20/i0[9] )
         );
  BUF_X2 \SB2_3_24/BUF_1  ( .I(\SB1_3_28/buf_output[1] ), .Z(\SB2_3_24/i0[6] )
         );
  CLKBUF_X2 \SB2_3_22/BUF_0  ( .I(\SB1_3_27/buf_output[0] ), .Z(
        \SB2_3_22/i0[9] ) );
  CLKBUF_X2 \SB2_3_9/BUF_0  ( .I(\SB1_3_14/buf_output[0] ), .Z(\SB2_3_9/i0[9] ) );
  BUF_X2 \SB2_3_9/BUF_1  ( .I(\SB1_3_13/buf_output[1] ), .Z(\SB2_3_9/i0[6] )
         );
  CLKBUF_X2 \SB2_3_15/BUF_0  ( .I(\SB1_3_20/buf_output[0] ), .Z(
        \SB2_3_15/i0[9] ) );
  BUF_X2 \SB2_3_23/BUF_3  ( .I(\SB1_3_25/buf_output[3] ), .Z(\SB2_3_23/i0[10] ) );
  BUF_X2 \SB2_3_31/BUF_0  ( .I(\SB1_3_4/buf_output[0] ), .Z(\SB2_3_31/i0[9] )
         );
  INV_X2 U3710 ( .I(n2692), .ZN(\SB2_3_24/i0_4 ) );
  INV_X2 U736 ( .I(\SB2_3_13/i0[7] ), .ZN(\SB1_3_14/buf_output[4] ) );
  INV_X2 U9278 ( .I(n3678), .ZN(\SB2_3_7/i1[9] ) );
  INV_X1 U6336 ( .I(\SB1_3_6/buf_output[1] ), .ZN(\SB2_3_2/i1_7 ) );
  INV_X1 \SB2_3_16/INV_1  ( .I(\SB1_3_20/buf_output[1] ), .ZN(\SB2_3_16/i1_7 )
         );
  INV_X1 \SB2_3_25/INV_1  ( .I(\SB1_3_29/buf_output[1] ), .ZN(\SB2_3_25/i1_7 )
         );
  INV_X1 U8814 ( .I(\SB1_3_23/buf_output[3] ), .ZN(\SB2_3_21/i0[8] ) );
  INV_X1 U2569 ( .I(\SB1_3_12/buf_output[5] ), .ZN(\SB2_3_12/i1_5 ) );
  NAND3_X1 \SB2_3_21/Component_Function_5/N3  ( .A1(\SB2_3_21/i1[9] ), .A2(
        \SB1_3_22/buf_output[4] ), .A3(\SB2_3_21/i0_3 ), .ZN(
        \SB2_3_21/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_13/Component_Function_3/N4  ( .A1(\SB2_3_13/i1_5 ), .A2(
        \SB2_3_13/i0[8] ), .A3(\SB2_3_13/i3[0] ), .ZN(
        \SB2_3_13/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_3/Component_Function_4/N2  ( .A1(\SB2_3_3/i3[0] ), .A2(
        \SB2_3_3/i0_0 ), .A3(\SB2_3_3/i1_7 ), .ZN(
        \SB2_3_3/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U8457 ( .A1(\SB2_3_10/i0_3 ), .A2(\SB2_3_10/i0_0 ), .A3(
        \SB2_3_10/i0[7] ), .ZN(\SB2_3_10/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2970 ( .A1(\SB2_3_14/i0_3 ), .A2(\SB2_3_14/i0[9] ), .A3(
        \SB2_3_14/i0[8] ), .ZN(\SB2_3_14/Component_Function_2/NAND4_in[2] ) );
  NAND2_X1 \SB2_3_29/Component_Function_5/N1  ( .A1(\SB2_3_29/i0_0 ), .A2(
        \SB2_3_29/i3[0] ), .ZN(\SB2_3_29/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 U3666 ( .A1(\SB2_3_18/i0_0 ), .A2(\SB2_3_18/i3[0] ), .ZN(n1076) );
  NAND3_X1 \SB2_3_3/Component_Function_4/N3  ( .A1(\SB2_3_3/i0[9] ), .A2(
        \SB2_3_3/i0[10] ), .A3(\SB2_3_3/i0_3 ), .ZN(
        \SB2_3_3/Component_Function_4/NAND4_in[2] ) );
  NAND2_X1 \SB2_3_21/Component_Function_5/N1  ( .A1(\SB2_3_21/i0_0 ), .A2(
        \SB2_3_21/i3[0] ), .ZN(\SB2_3_21/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U3707 ( .A1(\SB2_3_16/i0[10] ), .A2(\SB2_3_16/i0_4 ), .A3(
        \SB2_3_16/i0_3 ), .ZN(\SB2_3_16/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 \SB2_3_9/Component_Function_5/N1  ( .A1(\SB2_3_9/i0_0 ), .A2(
        \SB2_3_9/i3[0] ), .ZN(\SB2_3_9/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_9/Component_Function_1/N4  ( .A1(\SB2_3_9/i1_7 ), .A2(
        \SB2_3_9/i0[8] ), .A3(\SB2_3_9/i0_4 ), .ZN(
        \SB2_3_9/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_17/Component_Function_2/N2  ( .A1(\SB2_3_17/i0_3 ), .A2(
        \SB2_3_17/i0[10] ), .A3(\SB2_3_17/i0[6] ), .ZN(
        \SB2_3_17/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U3744 ( .A1(\SB2_3_6/i0_0 ), .A2(\SB2_3_6/i0_3 ), .A3(
        \SB2_3_6/i0[7] ), .ZN(n2248) );
  NAND3_X1 U8955 ( .A1(\SB2_3_28/i0_3 ), .A2(n5490), .A3(n577), .ZN(
        \SB2_3_28/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_5/Component_Function_3/N1  ( .A1(n3671), .A2(\SB2_3_5/i0_3 ), 
        .A3(\SB2_3_5/i0[6] ), .ZN(\SB2_3_5/Component_Function_3/NAND4_in[0] )
         );
  NAND3_X1 U2497 ( .A1(n5491), .A2(\SB2_3_2/i3[0] ), .A3(\SB2_3_2/i1_5 ), .ZN(
        n3749) );
  NAND3_X1 U7088 ( .A1(\SB2_3_30/i0_4 ), .A2(\SB2_3_30/i1[9] ), .A3(
        \SB2_3_30/i1_5 ), .ZN(n2382) );
  NAND3_X1 \SB2_3_10/Component_Function_0/N2  ( .A1(\SB2_3_10/i0[8] ), .A2(
        \SB2_3_10/i0[7] ), .A3(\SB2_3_10/i0[6] ), .ZN(
        \SB2_3_10/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U2149 ( .A1(\SB2_3_16/i0_4 ), .A2(\SB2_3_16/i1_7 ), .A3(
        \SB2_3_16/i0[8] ), .ZN(n1828) );
  NAND3_X1 U3712 ( .A1(\SB2_3_31/i1_7 ), .A2(\SB2_3_31/i0[8] ), .A3(
        \SB2_3_31/i0_4 ), .ZN(\SB2_3_31/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U2164 ( .A1(\SB2_3_31/i0_3 ), .A2(\SB2_3_31/i1_7 ), .A3(
        \SB2_3_31/i0[8] ), .ZN(\SB2_3_31/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U8626 ( .A1(\SB2_3_23/i1_5 ), .A2(\SB2_3_23/i0[8] ), .A3(
        \SB2_3_23/i3[0] ), .ZN(\SB2_3_23/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U3039 ( .A1(\SB2_3_4/i0[10] ), .A2(\SB2_3_4/i0_3 ), .A3(
        \SB2_3_4/i0[9] ), .ZN(n3464) );
  NAND3_X1 U2559 ( .A1(\SB2_3_14/i0_0 ), .A2(\SB2_3_14/i0_4 ), .A3(
        \SB2_3_14/i1_5 ), .ZN(n4341) );
  NAND2_X1 U2145 ( .A1(\SB2_3_30/i0_0 ), .A2(\SB2_3_30/i3[0] ), .ZN(n1735) );
  NAND2_X1 \SB2_3_16/Component_Function_5/N1  ( .A1(\SB2_3_16/i0_0 ), .A2(
        \SB2_3_16/i3[0] ), .ZN(\SB2_3_16/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U3709 ( .A1(\SB2_3_7/i1[9] ), .A2(\SB2_3_7/i1_5 ), .A3(
        \SB1_3_8/buf_output[4] ), .ZN(
        \SB2_3_7/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U5204 ( .A1(\SB2_3_8/i0[10] ), .A2(\SB2_3_8/i1_7 ), .A3(n3669), 
        .ZN(n2408) );
  NAND3_X1 \SB2_3_6/Component_Function_5/N3  ( .A1(\SB2_3_6/i1[9] ), .A2(
        \SB2_3_6/i0_4 ), .A3(\SB2_3_6/i0_3 ), .ZN(
        \SB2_3_6/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1151 ( .A1(n2564), .A2(n5513), .A3(\SB2_3_0/i0[6] ), .ZN(n735) );
  NAND3_X1 U5616 ( .A1(\SB2_3_29/i0[6] ), .A2(\RI3[3][16] ), .A3(
        \SB2_3_29/i0[9] ), .ZN(n1734) );
  NAND3_X1 U673 ( .A1(\SB2_3_17/i0_3 ), .A2(\SB2_3_17/i0[8] ), .A3(
        \SB2_3_17/i0[9] ), .ZN(\SB2_3_17/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_7/Component_Function_1/N4  ( .A1(\SB2_3_7/i1_7 ), .A2(
        \SB2_3_7/i0[8] ), .A3(\SB1_3_8/buf_output[4] ), .ZN(
        \SB2_3_7/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U10296 ( .A1(\SB2_3_24/i0[9] ), .A2(\SB2_3_24/i0_4 ), .A3(
        \SB2_3_24/i0[6] ), .ZN(\SB2_3_24/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U8348 ( .A1(\SB2_3_1/i0_3 ), .A2(\SB2_3_1/i0_0 ), .A3(
        \SB2_3_1/i0_4 ), .ZN(\SB2_3_1/Component_Function_3/NAND4_in[1] ) );
  NAND2_X1 U3714 ( .A1(\SB2_3_15/i0[10] ), .A2(\SB2_3_15/i0[9] ), .ZN(
        \SB2_3_15/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U1780 ( .A1(\SB2_3_15/i0_3 ), .A2(\SB2_3_15/i0[10] ), .A3(
        \SB1_3_16/buf_output[4] ), .ZN(n3265) );
  NAND3_X1 U2998 ( .A1(n3670), .A2(\SB1_3_16/buf_output[4] ), .A3(
        \SB2_3_15/i1_7 ), .ZN(\SB2_3_15/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_14/Component_Function_2/N2  ( .A1(\SB2_3_14/i0_3 ), .A2(
        \SB2_3_14/i0[10] ), .A3(\SB2_3_14/i0[6] ), .ZN(
        \SB2_3_14/Component_Function_2/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_26/Component_Function_5/N1  ( .A1(\SB2_3_26/i0_0 ), .A2(
        \SB2_3_26/i3[0] ), .ZN(\SB2_3_26/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U676 ( .A1(\SB2_3_6/i0[10] ), .A2(\SB2_3_6/i0_3 ), .A3(
        \SB2_3_6/i0[6] ), .ZN(\SB2_3_6/Component_Function_2/NAND4_in[1] ) );
  NAND2_X1 \SB2_3_10/Component_Function_0/N1  ( .A1(\SB2_3_10/i0[10] ), .A2(
        \SB2_3_10/i0[9] ), .ZN(\SB2_3_10/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 \SB2_3_29/Component_Function_1/N1  ( .A1(\SB2_3_29/i0_3 ), .A2(
        \SB2_3_29/i1[9] ), .ZN(\SB2_3_29/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U1958 ( .A1(\SB2_3_4/i3[0] ), .A2(\SB2_3_4/i0[8] ), .A3(n5519), 
        .ZN(\SB2_3_4/Component_Function_3/NAND4_in[3] ) );
  NAND2_X1 U10517 ( .A1(\SB2_3_7/i0_0 ), .A2(n4354), .ZN(n4717) );
  NAND3_X1 U8675 ( .A1(\SB2_3_7/i0_3 ), .A2(n1670), .A3(\SB2_3_7/i1[9] ), .ZN(
        n4679) );
  NAND3_X1 \SB2_3_30/Component_Function_2/N1  ( .A1(\SB2_3_30/i1_5 ), .A2(
        \SB2_3_30/i0[10] ), .A3(\SB2_3_30/i1[9] ), .ZN(
        \SB2_3_30/Component_Function_2/NAND4_in[0] ) );
  NAND2_X1 U6406 ( .A1(\SB2_3_1/i0[10] ), .A2(\SB2_3_1/i0[6] ), .ZN(n3280) );
  INV_X1 U4782 ( .I(\SB1_3_4/buf_output[1] ), .ZN(\SB2_3_0/i1_7 ) );
  NAND3_X1 \SB2_3_13/Component_Function_3/N1  ( .A1(\SB2_3_13/i1[9] ), .A2(
        \SB2_3_13/i0_3 ), .A3(\SB2_3_13/i0[6] ), .ZN(
        \SB2_3_13/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 \SB2_3_15/Component_Function_1/N3  ( .A1(\SB2_3_15/i1_5 ), .A2(
        \SB2_3_15/i0[6] ), .A3(\SB2_3_15/i0[9] ), .ZN(
        \SB2_3_15/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U679 ( .A1(\SB2_3_29/i0[6] ), .A2(\SB2_3_29/i1_5 ), .A3(
        \SB2_3_29/i0[9] ), .ZN(n4334) );
  NAND3_X1 \SB2_3_5/Component_Function_2/N1  ( .A1(\SB2_3_5/i1_5 ), .A2(
        \SB2_3_5/i0[10] ), .A3(n3671), .ZN(
        \SB2_3_5/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U720 ( .A1(\SB2_3_21/i0[9] ), .A2(\SB1_3_22/buf_output[4] ), .A3(
        \SB2_3_21/i0[6] ), .ZN(\SB2_3_21/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U7139 ( .A1(\SB2_3_5/i0[9] ), .A2(\SB2_3_5/i1_5 ), .A3(
        \SB2_3_5/i0[6] ), .ZN(\SB2_3_5/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB2_3_2/Component_Function_4/N1  ( .A1(\SB2_3_2/i0[9] ), .A2(
        \SB2_3_2/i0_0 ), .A3(n5491), .ZN(
        \SB2_3_2/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U10102 ( .A1(\SB2_3_11/i0[6] ), .A2(n5240), .A3(n3645), .ZN(n4154)
         );
  NAND3_X1 U4710 ( .A1(\SB2_3_23/i0_3 ), .A2(\SB2_3_23/i1_7 ), .A3(
        \SB2_3_23/i0[8] ), .ZN(\SB2_3_23/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_16/Component_Function_2/N2  ( .A1(\SB2_3_16/i0_3 ), .A2(
        \SB2_3_16/i0[10] ), .A3(\SB2_3_16/i0[6] ), .ZN(
        \SB2_3_16/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 \SB2_3_29/Component_Function_4/N3  ( .A1(\SB2_3_29/i0[9] ), .A2(
        \SB2_3_29/i0[10] ), .A3(\SB2_3_29/i0_3 ), .ZN(
        \SB2_3_29/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U700 ( .A1(\SB2_3_19/i1_5 ), .A2(\SB2_3_19/i0[8] ), .A3(
        \SB2_3_19/i3[0] ), .ZN(\SB2_3_19/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2997 ( .A1(n3670), .A2(\SB2_3_15/i1_5 ), .A3(\SB2_3_15/i3[0] ), 
        .ZN(\SB2_3_15/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_20/Component_Function_3/N4  ( .A1(\SB2_3_20/i1_5 ), .A2(
        \SB2_3_20/i0[8] ), .A3(\SB2_3_20/i3[0] ), .ZN(
        \SB2_3_20/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U697 ( .A1(\SB2_3_0/i1_5 ), .A2(n5513), .A3(\SB2_3_0/i3[0] ), .ZN(
        \SB2_3_0/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U3702 ( .A1(\SB2_3_25/i3[0] ), .A2(\SB2_3_25/i0_0 ), .A3(
        \SB2_3_25/i1_7 ), .ZN(\SB2_3_25/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U10416 ( .A1(\SB2_3_22/i0[6] ), .A2(\SB2_3_22/i0[8] ), .A3(
        \SB2_3_22/i0[7] ), .ZN(\SB2_3_22/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U2475 ( .A1(\SB2_3_9/i0[10] ), .A2(\SB2_3_9/i1_7 ), .A3(
        \SB2_3_9/i1[9] ), .ZN(\SB2_3_9/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2910 ( .A1(\SB2_3_21/i0_3 ), .A2(\SB2_3_21/i0[9] ), .A3(
        \SB2_3_21/i0[8] ), .ZN(n3440) );
  NAND3_X1 \SB2_3_22/Component_Function_0/N4  ( .A1(\SB2_3_22/i0[7] ), .A2(
        \SB2_3_22/i0_3 ), .A3(\SB2_3_22/i0_0 ), .ZN(
        \SB2_3_22/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U5431 ( .A1(\SB2_3_27/i0_4 ), .A2(\SB2_3_27/i1_7 ), .A3(
        \SB2_3_27/i0[8] ), .ZN(n3140) );
  NAND3_X1 \SB2_3_30/Component_Function_3/N4  ( .A1(\SB2_3_30/i1_5 ), .A2(
        \SB2_3_30/i0[8] ), .A3(\SB2_3_30/i3[0] ), .ZN(
        \SB2_3_30/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U702 ( .A1(\SB2_3_26/i0_0 ), .A2(\SB2_3_26/i0_4 ), .A3(
        \SB2_3_26/i1_5 ), .ZN(n4628) );
  NAND3_X1 U5760 ( .A1(\SB2_3_21/i0_3 ), .A2(\SB2_3_21/i0[10] ), .A3(
        \SB2_3_21/i0[6] ), .ZN(n3185) );
  NAND3_X1 \SB2_3_17/Component_Function_1/N4  ( .A1(\SB2_3_17/i1_7 ), .A2(
        \SB2_3_17/i0[8] ), .A3(\SB2_3_17/i0_4 ), .ZN(
        \SB2_3_17/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_20/Component_Function_3/N1  ( .A1(\SB2_3_20/i1[9] ), .A2(
        \SB2_3_20/i0_3 ), .A3(\SB2_3_20/i0[6] ), .ZN(
        \SB2_3_20/Component_Function_3/NAND4_in[0] ) );
  NAND2_X1 U5108 ( .A1(\SB2_3_13/i0_0 ), .A2(\SB2_3_13/i3[0] ), .ZN(n1467) );
  NAND3_X1 U710 ( .A1(n2692), .A2(n2906), .A3(\SB2_3_24/i0[6] ), .ZN(n2312) );
  NAND3_X1 U9759 ( .A1(\SB2_3_11/i0[10] ), .A2(\SB2_3_11/i0_3 ), .A3(
        \SB2_3_11/i0[6] ), .ZN(\SB2_3_11/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U3726 ( .A1(\SB2_3_16/i1_5 ), .A2(\SB2_3_16/i0_0 ), .A3(
        \SB2_3_16/i0_4 ), .ZN(\SB2_3_16/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 \SB2_3_31/Component_Function_2/N1  ( .A1(\SB2_3_31/i1_5 ), .A2(
        \SB2_3_31/i0[10] ), .A3(\SB2_3_31/i1[9] ), .ZN(
        \SB2_3_31/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U8922 ( .A1(\SB2_3_2/i0[6] ), .A2(\SB2_3_2/i1_5 ), .A3(
        \SB2_3_2/i0[9] ), .ZN(\SB2_3_2/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 \SB2_3_4/Component_Function_0/N1  ( .A1(\SB2_3_4/i0[10] ), .A2(
        \SB2_3_4/i0[9] ), .ZN(\SB2_3_4/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U2292 ( .A1(\SB2_3_30/i0_0 ), .A2(\SB2_3_30/i0_3 ), .A3(
        \SB2_3_30/i0_4 ), .ZN(\SB2_3_30/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1644 ( .A1(\SB2_3_2/i1_5 ), .A2(\SB2_3_2/i0[10] ), .A3(
        \SB2_3_2/i1[9] ), .ZN(\SB2_3_2/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U690 ( .A1(\SB2_3_10/i0_0 ), .A2(\SB2_3_10/i0_4 ), .A3(
        \SB2_3_10/i1_5 ), .ZN(n2677) );
  NAND3_X1 U10217 ( .A1(\SB2_3_10/i0_3 ), .A2(\SB2_3_10/i1[9] ), .A3(
        \SB2_3_10/i0[6] ), .ZN(\SB2_3_10/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2159 ( .A1(\SB2_3_29/i0[10] ), .A2(\SB2_3_29/i0_3 ), .A3(
        \RI3[3][16] ), .ZN(n1402) );
  BUF_X2 U7907 ( .I(\SB2_3_26/buf_output[0] ), .Z(\RI5[3][60] ) );
  BUF_X2 U8900 ( .I(\SB2_3_14/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[132] ) );
  BUF_X2 \SB3_28/BUF_1  ( .I(\MC_ARK_ARC_1_3/buf_output[19] ), .Z(
        \SB3_28/i0[6] ) );
  BUF_X2 U1885 ( .I(\MC_ARK_ARC_1_3/buf_output[151] ), .Z(\SB3_6/i0[6] ) );
  BUF_X2 U4608 ( .I(\MC_ARK_ARC_1_3/buf_output[127] ), .Z(\SB3_10/i0[6] ) );
  BUF_X2 U4946 ( .I(\MC_ARK_ARC_1_3/buf_output[186] ), .Z(\SB3_0/i0[9] ) );
  NAND3_X1 U8768 ( .A1(\SB3_11/i0_3 ), .A2(\SB3_11/i0[8] ), .A3(\SB3_11/i0[9] ), .ZN(\SB3_11/Component_Function_2/NAND4_in[2] ) );
  BUF_X2 U8832 ( .I(\MC_ARK_ARC_1_3/buf_output[103] ), .Z(\SB3_14/i0[6] ) );
  INV_X1 \SB3_31/INV_0  ( .I(\MC_ARK_ARC_1_3/buf_output[0] ), .ZN(
        \SB3_31/i3[0] ) );
  BUF_X2 U1309 ( .I(\MC_ARK_ARC_1_3/buf_output[78] ), .Z(\SB3_18/i0[9] ) );
  BUF_X2 U4730 ( .I(\MC_ARK_ARC_1_3/buf_output[128] ), .Z(\SB3_10/i0_0 ) );
  CLKBUF_X2 U8902 ( .I(\MC_ARK_ARC_1_3/buf_output[75] ), .Z(\SB3_19/i0[10] )
         );
  BUF_X2 U3212 ( .I(\MC_ARK_ARC_1_3/buf_output[105] ), .Z(\SB3_14/i0[10] ) );
  BUF_X2 U4489 ( .I(\MC_ARK_ARC_1_3/buf_output[22] ), .Z(\SB3_28/i0_4 ) );
  CLKBUF_X2 U2172 ( .I(\MC_ARK_ARC_1_3/buf_output[16] ), .Z(\SB3_29/i0_4 ) );
  BUF_X2 \SB3_8/BUF_4  ( .I(\MC_ARK_ARC_1_3/buf_output[142] ), .Z(\SB3_8/i0_4 ) );
  BUF_X2 U663 ( .I(\MC_ARK_ARC_1_3/buf_output[13] ), .Z(\SB3_29/i0[6] ) );
  INV_X1 U8912 ( .I(\RI1[4][53] ), .ZN(\SB3_23/i1_5 ) );
  INV_X1 \SB3_10/INV_2  ( .I(\MC_ARK_ARC_1_3/buf_output[128] ), .ZN(
        \SB3_10/i1[9] ) );
  INV_X1 U4668 ( .I(\MC_ARK_ARC_1_3/buf_output[15] ), .ZN(\SB3_29/i0[8] ) );
  INV_X1 \SB3_13/INV_5  ( .I(\MC_ARK_ARC_1_3/buf_output[113] ), .ZN(
        \SB3_13/i1_5 ) );
  NAND3_X1 U8624 ( .A1(\SB3_13/i0_3 ), .A2(\SB3_13/i0[9] ), .A3(\SB3_13/i0[8] ), .ZN(n1079) );
  NAND3_X1 U637 ( .A1(\SB3_2/i0_0 ), .A2(\SB3_2/i0[7] ), .A3(\SB3_2/i0_3 ), 
        .ZN(n4431) );
  NAND3_X1 \SB3_31/Component_Function_2/N2  ( .A1(\SB3_31/i0_3 ), .A2(
        \SB3_31/i0[10] ), .A3(\SB3_31/i0[6] ), .ZN(
        \SB3_31/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U3751 ( .A1(\SB3_29/i1_5 ), .A2(\SB3_29/i0[10] ), .A3(
        \SB3_29/i1[9] ), .ZN(\SB3_29/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 \SB3_4/Component_Function_4/N4  ( .A1(\SB3_4/i1[9] ), .A2(n2910), 
        .A3(\SB3_4/i0_4 ), .ZN(\SB3_4/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 \SB3_27/Component_Function_1/N3  ( .A1(\SB3_27/i1_5 ), .A2(
        \SB3_27/i0[6] ), .A3(\SB3_27/i0[9] ), .ZN(
        \SB3_27/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 \SB3_18/Component_Function_1/N4  ( .A1(\SB3_18/i1_7 ), .A2(
        \SB3_18/i0[8] ), .A3(\SB3_18/i0_4 ), .ZN(
        \SB3_18/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_26/Component_Function_2/N1  ( .A1(\SB3_26/i1_5 ), .A2(
        \SB3_26/i0[10] ), .A3(\SB3_26/i1[9] ), .ZN(
        \SB3_26/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U2987 ( .A1(\SB3_23/i0_4 ), .A2(\SB3_23/i1[9] ), .A3(\SB3_23/i1_5 ), 
        .ZN(n823) );
  NAND3_X1 U1216 ( .A1(\SB3_18/i0_3 ), .A2(\SB3_18/i0[8] ), .A3(\SB3_18/i0[9] ), .ZN(\SB3_18/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1202 ( .A1(\SB3_6/i1_5 ), .A2(\SB3_6/i0[8] ), .A3(\SB3_6/i3[0] ), 
        .ZN(n774) );
  NAND2_X1 \SB3_17/Component_Function_5/N1  ( .A1(\SB3_17/i0_0 ), .A2(
        \SB3_17/i3[0] ), .ZN(\SB3_17/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 U4648 ( .A1(\SB3_8/i0_0 ), .A2(\SB3_8/i3[0] ), .ZN(
        \SB3_8/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB3_18/Component_Function_5/N1  ( .A1(\SB3_18/i0_0 ), .A2(
        \SB3_18/i3[0] ), .ZN(\SB3_18/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U8817 ( .A1(\SB3_9/i0_4 ), .A2(\SB3_9/i1[9] ), .A3(\SB3_9/i1_5 ), 
        .ZN(\SB3_9/Component_Function_4/NAND4_in[3] ) );
  NAND2_X1 \SB3_29/Component_Function_5/N1  ( .A1(\SB3_29/i0_0 ), .A2(
        \SB3_29/i3[0] ), .ZN(\SB3_29/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U10333 ( .A1(\SB3_17/i0[6] ), .A2(\SB3_17/i1_5 ), .A3(
        \SB3_17/i0[9] ), .ZN(\SB3_17/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U8963 ( .A1(\SB3_14/i0_3 ), .A2(\SB3_14/i0[8] ), .A3(\SB3_14/i0[9] ), .ZN(\SB3_14/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 \SB3_31/Component_Function_1/N3  ( .A1(\SB3_31/i1_5 ), .A2(
        \SB3_31/i0[6] ), .A3(\SB3_31/i0[9] ), .ZN(
        \SB3_31/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U2285 ( .A1(\SB3_10/i0[9] ), .A2(\SB3_10/i0[10] ), .A3(
        \SB3_10/i0_3 ), .ZN(\SB3_10/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2435 ( .A1(\SB3_17/i1_7 ), .A2(\SB3_17/i0[8] ), .A3(\SB3_17/i0_4 ), 
        .ZN(\SB3_17/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 \SB3_13/Component_Function_3/N1  ( .A1(\SB3_13/i1[9] ), .A2(
        \SB3_13/i0_3 ), .A3(\SB3_13/i0[6] ), .ZN(
        \SB3_13/Component_Function_3/NAND4_in[0] ) );
  NAND2_X1 \SB3_30/Component_Function_1/N1  ( .A1(\SB3_30/i0_3 ), .A2(
        \SB3_30/i1[9] ), .ZN(\SB3_30/Component_Function_1/NAND4_in[0] ) );
  NAND2_X1 \SB3_27/Component_Function_0/N1  ( .A1(\SB3_27/i0[10] ), .A2(
        \SB3_27/i0[9] ), .ZN(\SB3_27/Component_Function_0/NAND4_in[0] ) );
  NAND2_X1 U7706 ( .A1(\SB3_5/i0[9] ), .A2(\SB3_5/i0[10] ), .ZN(
        \SB3_5/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 \SB3_12/Component_Function_2/N1  ( .A1(\SB3_12/i1_5 ), .A2(
        \SB3_12/i0[10] ), .A3(\SB3_12/i1[9] ), .ZN(
        \SB3_12/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U598 ( .A1(\SB3_6/i1_5 ), .A2(\RI1[4][154] ), .A3(\SB3_6/i0_0 ), 
        .ZN(\SB3_6/Component_Function_2/NAND4_in[3] ) );
  NAND2_X1 U8781 ( .A1(\SB3_20/i3[0] ), .A2(\SB3_20/i0_0 ), .ZN(n3908) );
  NAND3_X1 U2609 ( .A1(\SB3_4/i0[6] ), .A2(\SB3_4/i0[9] ), .A3(\SB3_4/i0_4 ), 
        .ZN(n1863) );
  NAND3_X1 U6325 ( .A1(\SB3_29/i0[10] ), .A2(\SB3_29/i1[9] ), .A3(
        \SB3_29/i1_7 ), .ZN(n2023) );
  NAND3_X1 U1297 ( .A1(\SB3_12/i0_3 ), .A2(\SB3_12/i0[10] ), .A3(
        \SB3_12/i0[6] ), .ZN(\SB3_12/Component_Function_2/NAND4_in[1] ) );
  NAND2_X1 \SB3_1/Component_Function_0/N1  ( .A1(\SB3_1/i0[10] ), .A2(
        \SB3_1/i0[9] ), .ZN(\SB3_1/Component_Function_0/NAND4_in[0] ) );
  BUF_X2 U3765 ( .I(\SB3_13/buf_output[4] ), .Z(\SB4_12/i0_4 ) );
  CLKBUF_X2 \SB4_9/BUF_0  ( .I(\SB3_14/buf_output[0] ), .Z(\SB4_9/i0[9] ) );
  BUF_X2 U3187 ( .I(\SB3_13/buf_output[1] ), .Z(\SB4_9/i0[6] ) );
  CLKBUF_X2 U8707 ( .I(\SB3_18/buf_output[0] ), .Z(\SB4_13/i0[9] ) );
  BUF_X2 \SB4_7/BUF_1  ( .I(\SB3_11/buf_output[1] ), .Z(\SB4_7/i0[6] ) );
  BUF_X2 \SB4_29/BUF_0  ( .I(\SB3_2/buf_output[0] ), .Z(\SB4_29/i0[9] ) );
  CLKBUF_X2 U3090 ( .I(\SB3_30/buf_output[2] ), .Z(n2897) );
  BUF_X2 U4408 ( .I(\SB3_31/buf_output[1] ), .Z(\SB4_27/i0[6] ) );
  CLKBUF_X2 \SB4_8/BUF_0  ( .I(\SB3_13/buf_output[0] ), .Z(\SB4_8/i0[9] ) );
  CLKBUF_X2 \SB4_20/BUF_0  ( .I(\SB3_25/buf_output[0] ), .Z(\SB4_20/i0[9] ) );
  BUF_X2 \SB4_22/BUF_0  ( .I(\SB3_27/buf_output[0] ), .Z(\SB4_22/i0[9] ) );
  BUF_X2 U4576 ( .I(\SB3_16/buf_output[4] ), .Z(\SB4_15/i0_4 ) );
  BUF_X2 U580 ( .I(\SB3_5/buf_output[4] ), .Z(\SB4_4/i0_4 ) );
  INV_X1 \SB4_31/INV_0  ( .I(\SB3_4/buf_output[0] ), .ZN(\SB4_31/i3[0] ) );
  AND4_X1 U9025 ( .A1(n1490), .A2(\SB3_11/Component_Function_5/NAND4_in[2] ), 
        .A3(\SB3_11/Component_Function_5/NAND4_in[0] ), .A4(n3999), .Z(n3684)
         );
  NAND3_X1 U9415 ( .A1(\SB4_17/i1_7 ), .A2(\SB4_17/i0_4 ), .A3(n3661), .ZN(
        \SB4_17/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U8761 ( .A1(\SB4_22/i0_0 ), .A2(\SB4_22/i3[0] ), .A3(\SB4_22/i1_7 ), 
        .ZN(n4403) );
  NAND3_X1 \SB4_31/Component_Function_0/N2  ( .A1(n3652), .A2(\SB4_31/i0[7] ), 
        .A3(\SB4_31/i0[6] ), .ZN(\SB4_31/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U5862 ( .A1(\SB4_5/i0_4 ), .A2(\SB4_5/i1_7 ), .A3(\SB4_5/i0[8] ), 
        .ZN(n1816) );
  NAND3_X1 \SB4_2/Component_Function_3/N4  ( .A1(\SB4_2/i1_5 ), .A2(
        \SB4_2/i0[8] ), .A3(\SB4_2/i3[0] ), .ZN(
        \SB4_2/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U9443 ( .A1(\SB4_22/i0_3 ), .A2(\SB4_22/i0_0 ), .A3(\SB4_22/i0[7] ), 
        .ZN(\SB4_22/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 \SB4_22/Component_Function_5/N1  ( .A1(\SB4_22/i0_0 ), .A2(
        \SB4_22/i3[0] ), .ZN(\SB4_22/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 \SB4_2/Component_Function_0/N1  ( .A1(\SB4_2/i0[10] ), .A2(
        \SB4_2/i0[9] ), .ZN(\SB4_2/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U7252 ( .A1(\SB4_2/i0_3 ), .A2(\SB4_2/i0_4 ), .A3(\SB4_2/i1[9] ), 
        .ZN(\SB4_2/Component_Function_5/NAND4_in[2] ) );
  NAND4_X1 U12 ( .A1(n2607), .A2(\SB4_13/Component_Function_1/NAND4_in[2] ), 
        .A3(\SB4_13/Component_Function_1/NAND4_in[1] ), .A4(n3231), .ZN(n5028)
         );
  NAND3_X1 U26 ( .A1(\SB4_28/i0_0 ), .A2(\SB4_28/i0_3 ), .A3(\SB4_28/i0_4 ), 
        .ZN(n4646) );
  NAND3_X1 U65 ( .A1(\SB4_18/i0[6] ), .A2(\SB4_18/i0[9] ), .A3(\SB4_18/i0_4 ), 
        .ZN(n6082) );
  NAND3_X1 U66 ( .A1(\SB4_5/i0_4 ), .A2(\SB4_5/i0_3 ), .A3(\SB4_5/i1[9] ), 
        .ZN(\SB4_5/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U118 ( .A1(\SB4_22/i0_4 ), .A2(\SB4_22/i0_0 ), .A3(\SB4_22/i0_3 ), 
        .ZN(n5701) );
  NAND3_X1 U181 ( .A1(\SB4_31/i0_3 ), .A2(\SB4_31/i0[10] ), .A3(\SB4_31/i0[6] ), .ZN(n2529) );
  NAND3_X1 U182 ( .A1(\SB4_5/i0[10] ), .A2(\SB4_5/i0_3 ), .A3(\SB4_5/i0[9] ), 
        .ZN(\SB4_5/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U203 ( .A1(\SB4_31/i0_3 ), .A2(n3652), .A3(\SB4_31/i0[9] ), .ZN(
        \SB4_31/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U295 ( .A1(\SB4_22/i0_0 ), .A2(\SB4_22/i0[9] ), .A3(\SB4_22/i0[8] ), 
        .ZN(\SB4_22/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U314 ( .A1(\SB4_30/i0[6] ), .A2(\SB4_30/i0[8] ), .A3(\SB4_30/i0[7] ), .ZN(\SB4_30/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U323 ( .A1(\SB4_0/i0[10] ), .A2(\SB4_0/i0_3 ), .A3(\SB4_0/i0[6] ), 
        .ZN(n1031) );
  NAND3_X1 U573 ( .A1(\SB4_20/i0_4 ), .A2(\SB4_20/i0_0 ), .A3(\SB4_20/i0_3 ), 
        .ZN(n6217) );
  AND4_X1 U574 ( .A1(n2867), .A2(\SB3_30/Component_Function_5/NAND4_in[1] ), 
        .A3(\SB3_30/Component_Function_5/NAND4_in[0] ), .A4(n3110), .Z(n5525)
         );
  CLKBUF_X2 U582 ( .I(\SB3_10/buf_output[4] ), .Z(\SB4_9/i0_4 ) );
  CLKBUF_X2 U584 ( .I(\SB3_3/buf_output[0] ), .Z(\SB4_30/i0[9] ) );
  CLKBUF_X2 U585 ( .I(\SB3_8/buf_output[0] ), .Z(\SB4_3/i0[9] ) );
  CLKBUF_X2 U587 ( .I(\SB3_11/buf_output[0] ), .Z(\SB4_6/i0[9] ) );
  BUF_X2 U588 ( .I(\SB3_24/buf_output[1] ), .Z(\SB4_20/i0[6] ) );
  CLKBUF_X4 U589 ( .I(\SB3_30/buf_output[3] ), .Z(\SB4_28/i0[10] ) );
  NAND3_X1 U592 ( .A1(\SB3_2/i1[9] ), .A2(\SB3_2/i1_7 ), .A3(\SB3_2/i0[10] ), 
        .ZN(\SB3_2/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U593 ( .A1(\SB3_31/i0_3 ), .A2(\SB3_31/i0_0 ), .A3(\SB3_31/i0[7] ), 
        .ZN(n6537) );
  NAND3_X1 U595 ( .A1(\SB3_16/i0_0 ), .A2(\SB3_16/i0_3 ), .A3(\SB3_16/i0_4 ), 
        .ZN(\SB3_16/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U601 ( .A1(\SB3_20/i0[10] ), .A2(\SB3_20/i0_3 ), .A3(\SB3_20/i0[6] ), .ZN(n3106) );
  NAND3_X1 U602 ( .A1(\SB3_1/i0[10] ), .A2(\SB3_1/i1_5 ), .A3(n4765), .ZN(
        \SB3_1/Component_Function_2/NAND4_in[0] ) );
  NAND2_X1 U603 ( .A1(\SB3_11/i0_0 ), .A2(\SB3_11/i3[0] ), .ZN(
        \SB3_11/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U604 ( .A1(\SB3_30/i1[9] ), .A2(\SB3_30/i0[10] ), .A3(\SB3_30/i1_7 ), .ZN(n5798) );
  NAND3_X1 U606 ( .A1(\SB3_11/i0[6] ), .A2(n582), .A3(\SB3_11/i0[9] ), .ZN(
        \SB3_11/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 U611 ( .A1(\SB3_4/i0[9] ), .A2(\SB3_4/i0[10] ), .ZN(
        \SB3_4/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U612 ( .A1(\SB3_21/i0[9] ), .A2(\SB3_21/i0[8] ), .A3(\RI1[4][65] ), 
        .ZN(n5771) );
  NAND3_X1 U613 ( .A1(\SB3_0/i0_3 ), .A2(\SB3_0/i1[9] ), .A3(\SB3_0/i0[6] ), 
        .ZN(n6108) );
  NAND3_X1 U617 ( .A1(\SB3_31/i0[9] ), .A2(\SB3_31/i0_0 ), .A3(\SB3_31/i0[8] ), 
        .ZN(n4966) );
  NAND3_X1 U619 ( .A1(\SB3_2/i0[6] ), .A2(\SB3_2/i1_5 ), .A3(\SB3_2/i0[9] ), 
        .ZN(n5662) );
  NAND3_X1 U621 ( .A1(\SB3_16/i0_3 ), .A2(\SB3_16/i0[9] ), .A3(\SB3_16/i0[8] ), 
        .ZN(n5729) );
  NAND3_X1 U625 ( .A1(\SB3_12/i3[0] ), .A2(\SB3_12/i0_0 ), .A3(\SB3_12/i1_7 ), 
        .ZN(n6079) );
  NAND3_X1 U627 ( .A1(\SB3_12/i0[8] ), .A2(\SB3_12/i3[0] ), .A3(\SB3_12/i1_5 ), 
        .ZN(n3912) );
  NAND3_X1 U629 ( .A1(\SB3_1/i0[9] ), .A2(\SB3_1/i0[8] ), .A3(\SB3_1/i0_3 ), 
        .ZN(\SB3_1/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U630 ( .A1(\SB3_24/i0[8] ), .A2(\SB3_24/i1_5 ), .A3(\SB3_24/i3[0] ), 
        .ZN(n4530) );
  NAND3_X1 U632 ( .A1(\SB3_3/i0_4 ), .A2(\SB3_3/i0[8] ), .A3(\SB3_3/i1_7 ), 
        .ZN(\SB3_3/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U633 ( .A1(\SB3_0/i0[8] ), .A2(\SB3_0/i3[0] ), .A3(\SB3_0/i1_5 ), 
        .ZN(n5791) );
  NAND3_X1 U634 ( .A1(\SB3_25/i1[9] ), .A2(\SB3_25/i0[10] ), .A3(\SB3_25/i1_7 ), .ZN(n6001) );
  NAND3_X1 U636 ( .A1(\SB3_19/i0_3 ), .A2(\SB3_19/i1[9] ), .A3(\SB3_19/i0_4 ), 
        .ZN(\SB3_19/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U638 ( .A1(\SB3_14/i0[9] ), .A2(\SB3_14/i0[6] ), .A3(\SB3_14/i0_4 ), 
        .ZN(n5140) );
  NAND3_X1 U641 ( .A1(\SB3_2/i0[6] ), .A2(\SB3_2/i0_3 ), .A3(\SB3_2/i1[9] ), 
        .ZN(\SB3_2/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U642 ( .A1(\SB3_7/i0[10] ), .A2(\SB3_7/i0_3 ), .A3(\SB3_7/i0[9] ), 
        .ZN(n4870) );
  CLKBUF_X2 U644 ( .I(\MC_ARK_ARC_1_3/buf_output[99] ), .Z(\SB3_15/i0[10] ) );
  BUF_X2 U646 ( .I(\MC_ARK_ARC_1_3/buf_output[23] ), .Z(\SB3_28/i0_3 ) );
  BUF_X2 U648 ( .I(\MC_ARK_ARC_1_3/buf_output[118] ), .Z(\SB3_12/i0_4 ) );
  BUF_X2 U649 ( .I(\MC_ARK_ARC_1_3/buf_output[38] ), .Z(\SB3_25/i0_0 ) );
  INV_X1 U650 ( .I(\RI1[4][77] ), .ZN(\SB3_19/i1_5 ) );
  NAND3_X1 U653 ( .A1(\SB3_1/i3[0] ), .A2(\SB3_1/i0[8] ), .A3(\SB3_1/i1_5 ), 
        .ZN(n4668) );
  BUF_X2 U654 ( .I(\SB2_3_12/buf_output[5] ), .Z(n5503) );
  NAND3_X1 U655 ( .A1(\SB2_3_9/i0[9] ), .A2(\SB2_3_9/i0_0 ), .A3(
        \SB2_3_9/i0[8] ), .ZN(\SB2_3_9/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U658 ( .A1(\SB2_3_31/i0_4 ), .A2(\SB2_3_31/i0_0 ), .A3(
        \SB2_3_31/i1_5 ), .ZN(n5541) );
  NAND3_X1 U661 ( .A1(\SB2_3_22/i0_0 ), .A2(\SB2_3_22/i1_5 ), .A3(
        \SB2_3_22/i0_4 ), .ZN(n4671) );
  NAND3_X1 U665 ( .A1(\SB2_3_0/i0[6] ), .A2(\SB2_3_0/i0[9] ), .A3(
        \SB2_3_0/i1_5 ), .ZN(n4371) );
  NAND3_X1 U671 ( .A1(\SB2_3_4/i0_3 ), .A2(\SB2_3_4/i0_0 ), .A3(
        \SB2_3_4/i0[7] ), .ZN(n6057) );
  NAND3_X1 U675 ( .A1(\SB2_3_30/i0[10] ), .A2(\SB2_3_30/i1_7 ), .A3(
        \SB2_3_30/i1[9] ), .ZN(n918) );
  NAND3_X1 U677 ( .A1(\SB2_3_5/i0_3 ), .A2(\SB2_3_5/i0[10] ), .A3(
        \SB2_3_5/i0[9] ), .ZN(n1844) );
  NAND3_X1 U680 ( .A1(\SB2_3_9/i1_5 ), .A2(\SB2_3_9/i0[8] ), .A3(
        \SB2_3_9/i3[0] ), .ZN(\SB2_3_9/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U681 ( .A1(\SB2_3_10/i0_3 ), .A2(\SB2_3_10/i0_4 ), .A3(
        \SB2_3_10/i0_0 ), .ZN(n6431) );
  NAND3_X1 U682 ( .A1(\SB2_3_3/i0_0 ), .A2(\SB2_3_3/i0[7] ), .A3(
        \SB2_3_3/i0_3 ), .ZN(\SB2_3_3/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U693 ( .A1(\SB2_3_9/i0_3 ), .A2(\SB2_3_9/i0_0 ), .A3(
        \SB2_3_9/i0[7] ), .ZN(n6093) );
  NAND3_X1 U694 ( .A1(\RI3[3][16] ), .A2(\SB2_3_29/i0_0 ), .A3(\SB2_3_29/i1_5 ), .ZN(\SB2_3_29/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U698 ( .A1(\SB2_3_21/i0_0 ), .A2(\SB2_3_21/i0[10] ), .A3(
        \SB2_3_21/i0[6] ), .ZN(n5132) );
  NAND2_X1 U705 ( .A1(\SB2_3_3/i0_0 ), .A2(\SB2_3_3/i3[0] ), .ZN(n6020) );
  NAND3_X1 U706 ( .A1(\SB2_3_3/i0_0 ), .A2(\SB2_3_3/i0[6] ), .A3(
        \SB2_3_3/i0[10] ), .ZN(n6016) );
  NAND3_X1 U707 ( .A1(\SB2_3_5/i0_3 ), .A2(\SB2_3_5/i0_4 ), .A3(\SB2_3_5/i0_0 ), .ZN(\SB2_3_5/Component_Function_3/NAND4_in[1] ) );
  INV_X1 U708 ( .I(\SB2_3_20/i0_4 ), .ZN(\SB2_3_20/i0[7] ) );
  NAND3_X1 U709 ( .A1(\SB2_3_8/i0[7] ), .A2(\SB2_3_8/i0_0 ), .A3(
        \SB2_3_8/i0_3 ), .ZN(\SB2_3_8/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U711 ( .A1(\SB2_3_11/i0[9] ), .A2(\SB2_3_11/i0_3 ), .A3(
        \SB2_3_11/i0[10] ), .ZN(n5291) );
  NAND3_X1 U712 ( .A1(\SB2_3_3/i0_4 ), .A2(\SB2_3_3/i0[9] ), .A3(
        \SB2_3_3/i0[6] ), .ZN(n1477) );
  NAND3_X1 U713 ( .A1(\SB2_3_11/i0_3 ), .A2(\SB2_3_11/i0_0 ), .A3(n3645), .ZN(
        \SB2_3_11/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U717 ( .A1(\SB2_3_7/i0[9] ), .A2(\SB2_3_7/i1_5 ), .A3(n1670), .ZN(
        \SB2_3_7/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U718 ( .A1(\SB2_3_25/i0_0 ), .A2(\SB2_3_25/i1_5 ), .A3(
        \SB1_3_26/buf_output[4] ), .ZN(
        \SB2_3_25/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U719 ( .A1(\SB2_3_18/i0_3 ), .A2(\SB2_3_18/i0[8] ), .A3(
        \SB2_3_18/i1_7 ), .ZN(\SB2_3_18/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U721 ( .A1(\SB1_3_14/buf_output[4] ), .A2(\SB2_3_13/i0_0 ), .A3(
        \SB2_3_13/i1_5 ), .ZN(\SB2_3_13/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U725 ( .A1(\SB2_3_25/i0[9] ), .A2(\SB2_3_25/i0_3 ), .A3(
        \SB2_3_25/i0[8] ), .ZN(n4929) );
  NAND3_X1 U728 ( .A1(n5511), .A2(n2911), .A3(\SB2_3_28/i1_5 ), .ZN(n5637) );
  NAND3_X1 U729 ( .A1(\SB2_3_2/i0_3 ), .A2(\SB2_3_2/i0_4 ), .A3(
        \SB2_3_2/i0[10] ), .ZN(n5393) );
  NAND3_X1 U741 ( .A1(\SB2_3_11/i0_3 ), .A2(\SB2_3_11/i1[9] ), .A3(
        \SB2_3_11/i0[6] ), .ZN(\SB2_3_11/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U742 ( .A1(\SB2_3_8/i0_0 ), .A2(\SB2_3_8/i3[0] ), .A3(
        \SB2_3_8/i1_7 ), .ZN(n5468) );
  NAND3_X1 U743 ( .A1(\SB2_3_2/i0_0 ), .A2(\SB2_3_2/i3[0] ), .A3(
        \SB2_3_2/i1_7 ), .ZN(n5483) );
  NAND3_X1 U744 ( .A1(\SB2_3_0/i0_3 ), .A2(\SB2_3_0/i0[10] ), .A3(
        \SB1_3_1/buf_output[4] ), .ZN(
        \SB2_3_0/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U745 ( .A1(\SB2_3_13/i0[10] ), .A2(\SB2_3_13/i0_3 ), .A3(
        \SB2_3_13/i0[9] ), .ZN(\SB2_3_13/Component_Function_4/NAND4_in[2] ) );
  AND2_X1 U747 ( .A1(\SB1_3_8/buf_output[1] ), .A2(\SB1_3_6/buf_output[3] ), 
        .Z(n2261) );
  INV_X2 U749 ( .I(n5890), .ZN(\SB1_3_28/buf_output[3] ) );
  BUF_X2 U753 ( .I(\SB1_3_0/buf_output[0] ), .Z(\RI3[3][24] ) );
  INV_X1 U762 ( .I(\SB1_3_26/buf_output[1] ), .ZN(\SB2_3_22/i1_7 ) );
  NAND2_X1 U763 ( .A1(\SB1_3_4/Component_Function_3/NAND4_in[1] ), .A2(n5756), 
        .ZN(n4962) );
  NAND2_X1 U766 ( .A1(\SB1_3_18/i0_3 ), .A2(\SB1_3_18/i1[9] ), .ZN(n5342) );
  NAND2_X1 U767 ( .A1(\SB1_3_11/i0[6] ), .A2(n5539), .ZN(
        \SB1_3_11/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 U769 ( .A1(\SB1_3_24/i0[6] ), .A2(n5970), .ZN(n1341) );
  NAND2_X1 U779 ( .A1(\SB1_3_11/i0[9] ), .A2(\SB1_3_11/i0[10] ), .ZN(n4974) );
  NAND2_X1 U780 ( .A1(\SB1_3_4/i0_3 ), .A2(\SB1_3_4/i1[9] ), .ZN(n4394) );
  NAND3_X1 U782 ( .A1(\SB1_3_29/i0_3 ), .A2(\RI1[3][14] ), .A3(\SB1_3_29/i0_4 ), .ZN(\SB1_3_29/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U784 ( .A1(\SB1_3_4/i0[10] ), .A2(\SB1_3_4/i0_3 ), .A3(
        \SB1_3_4/i0[9] ), .ZN(n6279) );
  NAND3_X1 U795 ( .A1(\SB1_3_27/i0_4 ), .A2(\SB1_3_27/i1_7 ), .A3(
        \SB1_3_27/i0[8] ), .ZN(n1817) );
  NAND3_X1 U796 ( .A1(\SB1_3_18/i0[10] ), .A2(\SB1_3_18/i0[9] ), .A3(
        \SB1_3_18/i0_3 ), .ZN(\SB1_3_18/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U797 ( .A1(\SB1_3_26/i0_3 ), .A2(\SB1_3_26/i0[8] ), .A3(
        \SB1_3_26/i0[9] ), .ZN(n3931) );
  NAND3_X1 U799 ( .A1(\SB1_3_7/i0[9] ), .A2(\SB1_3_7/i0[6] ), .A3(
        \SB1_3_7/i0_4 ), .ZN(n6498) );
  NAND3_X1 U801 ( .A1(\SB1_3_2/i0[6] ), .A2(\SB1_3_2/i1_5 ), .A3(
        \SB1_3_2/i0[9] ), .ZN(\SB1_3_2/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U802 ( .A1(\SB1_3_14/i0_0 ), .A2(\SB1_3_14/i1_5 ), .A3(
        \SB1_3_14/i0_4 ), .ZN(n5355) );
  NAND2_X1 U803 ( .A1(\SB1_3_14/Component_Function_4/NAND4_in[2] ), .A2(n5992), 
        .ZN(n2602) );
  NAND2_X1 U804 ( .A1(\SB1_3_25/i0_0 ), .A2(\SB1_3_25/i3[0] ), .ZN(n5684) );
  NAND3_X1 U808 ( .A1(\SB1_3_19/i0_4 ), .A2(\SB1_3_19/i0[9] ), .A3(
        \SB1_3_19/i0[6] ), .ZN(n6252) );
  NAND2_X1 U809 ( .A1(\SB1_3_30/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_3_30/Component_Function_4/NAND4_in[2] ), .ZN(n5231) );
  NAND3_X1 U812 ( .A1(\SB1_3_6/i0[9] ), .A2(\SB1_3_6/i0[6] ), .A3(
        \SB1_3_6/i1_5 ), .ZN(n5720) );
  NAND3_X1 U815 ( .A1(\SB1_3_4/i0_3 ), .A2(\SB1_3_4/i1_7 ), .A3(
        \SB1_3_4/i0[8] ), .ZN(\SB1_3_4/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U816 ( .A1(\SB1_3_0/i0_0 ), .A2(\SB1_3_0/i0_3 ), .A3(
        \SB1_3_0/i0[7] ), .ZN(n5307) );
  NAND3_X1 U817 ( .A1(\SB1_3_21/i0_4 ), .A2(\SB1_3_21/i0[8] ), .A3(
        \SB1_3_21/i1_7 ), .ZN(n5708) );
  NAND3_X1 U818 ( .A1(\SB1_3_18/i0_3 ), .A2(\SB1_3_18/i0[8] ), .A3(
        \SB1_3_18/i1_7 ), .ZN(\SB1_3_18/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U820 ( .A1(\SB1_3_28/i0_0 ), .A2(\SB1_3_28/i0_4 ), .A3(
        \SB1_3_28/i1_5 ), .ZN(n5542) );
  NAND3_X1 U823 ( .A1(\SB1_3_27/i0[10] ), .A2(\SB1_3_27/i1[9] ), .A3(
        \SB1_3_27/i1_7 ), .ZN(n5379) );
  NAND3_X1 U825 ( .A1(\SB1_3_16/i1_7 ), .A2(\SB1_3_16/i0[10] ), .A3(
        \SB1_3_16/i1[9] ), .ZN(n6382) );
  NAND3_X1 U827 ( .A1(\SB1_3_3/i0[8] ), .A2(\SB1_3_3/i3[0] ), .A3(
        \SB1_3_3/i1_5 ), .ZN(n4782) );
  NAND3_X1 U829 ( .A1(\SB1_3_17/i0_4 ), .A2(\SB1_3_17/i1_7 ), .A3(
        \SB1_3_17/i0[8] ), .ZN(n6417) );
  NAND3_X1 U833 ( .A1(\SB1_3_14/i0[8] ), .A2(\SB1_3_14/i1_5 ), .A3(
        \SB1_3_14/i3[0] ), .ZN(n6036) );
  NAND3_X1 U836 ( .A1(\SB1_3_6/i0[8] ), .A2(\SB1_3_6/i3[0] ), .A3(
        \SB1_3_6/i1_5 ), .ZN(n5100) );
  NAND3_X1 U838 ( .A1(\SB1_3_20/i0_4 ), .A2(\SB1_3_20/i0[9] ), .A3(
        \SB1_3_20/i0[6] ), .ZN(n6406) );
  NAND3_X1 U839 ( .A1(\SB1_3_18/i0_3 ), .A2(\SB1_3_18/i1[9] ), .A3(
        \SB1_3_18/i0[6] ), .ZN(n5062) );
  NAND3_X1 U841 ( .A1(\SB1_3_29/i0[8] ), .A2(\SB1_3_29/i1_5 ), .A3(
        \SB1_3_29/i3[0] ), .ZN(\SB1_3_29/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U844 ( .A1(\SB1_3_3/i0[6] ), .A2(\SB1_3_3/i1[9] ), .A3(
        \SB1_3_3/i0_3 ), .ZN(n5154) );
  NAND3_X1 U845 ( .A1(\SB1_3_19/i0_3 ), .A2(\SB1_3_19/i1[9] ), .A3(
        \SB1_3_19/i0[6] ), .ZN(n5287) );
  NAND3_X1 U848 ( .A1(\SB1_3_14/i0[10] ), .A2(\SB1_3_14/i1[9] ), .A3(
        \SB1_3_14/i1_7 ), .ZN(n6216) );
  NAND3_X1 U860 ( .A1(\SB1_3_21/i0_3 ), .A2(\SB1_3_21/i0[10] ), .A3(
        \SB1_3_21/i0[9] ), .ZN(n1060) );
  NAND3_X1 U863 ( .A1(\SB1_3_16/i0_3 ), .A2(\SB1_3_16/i0[9] ), .A3(
        \SB1_3_16/i0[8] ), .ZN(n6037) );
  INV_X2 U864 ( .I(\RI1[3][131] ), .ZN(\SB1_3_10/i1_5 ) );
  INV_X1 U872 ( .I(n5550), .ZN(n2908) );
  BUF_X2 U878 ( .I(\RI1[3][41] ), .Z(\SB1_3_25/i0_3 ) );
  BUF_X2 U885 ( .I(\RI1[3][89] ), .Z(\SB1_3_17/i0_3 ) );
  NAND2_X1 U886 ( .A1(n6125), .A2(n4835), .ZN(n1508) );
  NAND3_X1 U889 ( .A1(\SB2_2_22/i0_0 ), .A2(\SB2_2_22/i0_3 ), .A3(
        \SB2_2_22/i0_4 ), .ZN(\SB2_2_22/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U890 ( .A1(\SB2_2_20/i0[6] ), .A2(\SB2_2_20/i0_3 ), .A3(
        \SB2_2_20/i1[9] ), .ZN(n6178) );
  NAND3_X1 U892 ( .A1(\SB2_2_20/i0[10] ), .A2(\SB2_2_20/i0_0 ), .A3(
        \SB2_2_20/i0[6] ), .ZN(\SB2_2_20/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U896 ( .A1(\SB2_2_29/i0_3 ), .A2(\SB2_2_29/i1_7 ), .A3(
        \SB2_2_29/i0[8] ), .ZN(\SB2_2_29/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U897 ( .A1(n2074), .A2(\SB2_2_6/i0_0 ), .A3(\SB2_2_6/i0_3 ), .ZN(
        \SB2_2_6/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U899 ( .A1(\SB2_2_22/i0_3 ), .A2(\SB2_2_22/i0[8] ), .A3(
        \SB2_2_22/i0[9] ), .ZN(\SB2_2_22/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U910 ( .A1(\SB2_2_3/i0_3 ), .A2(\SB2_2_3/i1_7 ), .A3(
        \SB2_2_3/i0[8] ), .ZN(n5256) );
  NAND3_X1 U911 ( .A1(\SB2_2_11/i0_3 ), .A2(\SB2_2_11/i0[9] ), .A3(
        \SB2_2_11/i0[8] ), .ZN(n5146) );
  NAND3_X1 U912 ( .A1(\SB2_2_28/i0[8] ), .A2(\SB2_2_28/i3[0] ), .A3(
        \SB2_2_28/i1_5 ), .ZN(n5863) );
  NAND3_X1 U916 ( .A1(\SB2_2_18/i0_4 ), .A2(\SB2_2_18/i0_3 ), .A3(
        \SB2_2_18/i0_0 ), .ZN(\SB2_2_18/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U918 ( .A1(\SB2_2_6/i0_0 ), .A2(\SB2_2_6/i0[9] ), .A3(
        \SB2_2_6/i0[8] ), .ZN(n5472) );
  NAND3_X1 U919 ( .A1(\SB2_2_4/i0[6] ), .A2(\SB2_2_4/i1_5 ), .A3(
        \SB2_2_4/i0[9] ), .ZN(n5762) );
  NAND3_X1 U923 ( .A1(\SB2_2_31/i0[10] ), .A2(\SB2_2_31/i1[9] ), .A3(
        \SB2_2_31/i1_7 ), .ZN(\SB2_2_31/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U928 ( .A1(\SB2_2_10/i0_0 ), .A2(\SB2_2_10/i0[7] ), .A3(
        \SB2_2_10/i0_3 ), .ZN(n4676) );
  NAND2_X1 U929 ( .A1(\SB2_2_11/i0_0 ), .A2(\SB2_2_11/i3[0] ), .ZN(n5987) );
  NAND3_X1 U930 ( .A1(\SB2_2_25/i1_5 ), .A2(\SB2_2_25/i0[10] ), .A3(
        \SB2_2_25/i1[9] ), .ZN(\SB2_2_25/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U934 ( .A1(\SB2_2_3/i0[9] ), .A2(\SB2_2_3/i1_5 ), .A3(
        \SB2_2_3/i0[6] ), .ZN(n5728) );
  NAND3_X1 U937 ( .A1(\SB2_2_25/i1_5 ), .A2(\SB2_2_25/i0[8] ), .A3(
        \SB2_2_25/i3[0] ), .ZN(\SB2_2_25/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U938 ( .A1(\SB2_2_17/i0_4 ), .A2(\SB2_2_17/i1_5 ), .A3(
        \SB2_2_17/i1[9] ), .ZN(n6467) );
  NAND3_X1 U939 ( .A1(\SB2_2_22/i0_3 ), .A2(\SB2_2_22/i0_4 ), .A3(
        \SB2_2_22/i1[9] ), .ZN(n1884) );
  NAND3_X1 U946 ( .A1(\SB2_2_8/i0_3 ), .A2(\SB2_2_8/i0[9] ), .A3(
        \SB2_2_8/i0[10] ), .ZN(\SB2_2_8/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U958 ( .A1(\SB2_2_26/i0_0 ), .A2(\SB2_2_26/i3[0] ), .A3(
        \SB2_2_26/i1_7 ), .ZN(\SB2_2_26/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U960 ( .A1(\SB2_2_26/i0[6] ), .A2(\SB2_2_26/i0_3 ), .A3(
        \SB2_2_26/i0[10] ), .ZN(\SB2_2_26/Component_Function_2/NAND4_in[1] )
         );
  AND2_X1 U963 ( .A1(n4749), .A2(\SB1_2_15/buf_output[1] ), .Z(n4754) );
  NAND3_X1 U967 ( .A1(\SB2_2_27/i0_3 ), .A2(\SB2_2_27/i0[9] ), .A3(
        \SB2_2_27/i0[8] ), .ZN(\SB2_2_27/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U968 ( .A1(\SB2_2_10/i0_0 ), .A2(\SB2_2_10/i3[0] ), .A3(
        \SB2_2_10/i1_7 ), .ZN(\SB2_2_10/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U969 ( .A1(\SB2_2_1/i0[6] ), .A2(\SB2_2_1/i0[9] ), .A3(
        \SB2_2_1/i0_4 ), .ZN(n5469) );
  NAND3_X1 U970 ( .A1(\SB2_2_3/i3[0] ), .A2(\SB2_2_3/i0[8] ), .A3(
        \SB2_2_3/i1_5 ), .ZN(\SB2_2_3/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U973 ( .A1(\SB2_2_23/i0[8] ), .A2(\SB2_2_23/i3[0] ), .A3(
        \SB2_2_23/i1_5 ), .ZN(\SB2_2_23/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U983 ( .A1(n5512), .A2(\SB2_2_28/i0[10] ), .A3(\SB2_2_28/i0[9] ), 
        .ZN(n5021) );
  NAND3_X1 U984 ( .A1(\SB2_2_24/i0_4 ), .A2(\SB2_2_24/i1_5 ), .A3(
        \SB2_2_24/i0_0 ), .ZN(n3201) );
  NAND3_X1 U985 ( .A1(\SB2_2_13/i0[9] ), .A2(\SB2_2_13/i0_0 ), .A3(
        \SB2_2_13/i0[8] ), .ZN(n5209) );
  NAND3_X1 U988 ( .A1(\SB2_2_29/i0[8] ), .A2(\SB2_2_29/i3[0] ), .A3(
        \SB2_2_29/i1_5 ), .ZN(n5438) );
  NAND3_X1 U989 ( .A1(\SB2_2_15/i0_0 ), .A2(\SB2_2_15/i0_3 ), .A3(
        \SB2_2_15/i0_4 ), .ZN(n4771) );
  NAND3_X1 U991 ( .A1(\SB2_2_22/i0[10] ), .A2(\SB2_2_22/i0[9] ), .A3(
        \SB2_2_22/i0_3 ), .ZN(n5182) );
  INV_X1 U998 ( .I(\SB2_2_28/i1_5 ), .ZN(n5512) );
  NOR2_X1 U1003 ( .A1(n5883), .A2(n5881), .ZN(n4015) );
  NAND3_X1 U1004 ( .A1(\SB1_2_9/i0[10] ), .A2(\SB1_2_9/i1[9] ), .A3(
        \SB1_2_9/i1_7 ), .ZN(n2922) );
  NAND3_X1 U1009 ( .A1(\SB1_2_14/i0_3 ), .A2(\SB1_2_14/i0_0 ), .A3(
        \SB1_2_14/i0[7] ), .ZN(n4578) );
  NAND3_X1 U1012 ( .A1(\SB1_2_22/i0[10] ), .A2(\SB1_2_22/i0_0 ), .A3(
        \SB1_2_22/i0[6] ), .ZN(\SB1_2_22/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1014 ( .A1(\SB1_2_22/i0[6] ), .A2(\SB1_2_22/i0[9] ), .A3(
        \SB1_2_22/i0_4 ), .ZN(n5982) );
  NAND3_X1 U1015 ( .A1(\SB1_2_28/i0_0 ), .A2(\SB1_2_28/i1_5 ), .A3(
        \SB1_2_28/i0_4 ), .ZN(n5419) );
  NAND3_X1 U1017 ( .A1(\SB1_2_1/i0[6] ), .A2(\SB1_2_1/i0_3 ), .A3(
        \SB1_2_1/i0[10] ), .ZN(n6461) );
  NAND3_X1 U1019 ( .A1(\SB1_2_17/i1[9] ), .A2(\SB1_2_17/i0_3 ), .A3(
        \SB1_2_17/i0[6] ), .ZN(\SB1_2_17/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U1021 ( .A1(\SB1_2_25/i0[10] ), .A2(\SB1_2_25/i1[9] ), .A3(
        \SB1_2_25/i1_5 ), .ZN(\SB1_2_25/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U1022 ( .A1(\SB1_2_25/i0[10] ), .A2(\SB1_2_25/i0_0 ), .A3(
        \SB1_2_25/i0[6] ), .ZN(\SB1_2_25/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1024 ( .A1(\SB1_2_17/i0_3 ), .A2(\SB1_2_17/i0[9] ), .A3(
        \SB1_2_17/i0[10] ), .ZN(n6308) );
  NAND2_X1 U1028 ( .A1(\SB1_2_29/Component_Function_4/NAND4_in[3] ), .A2(n6124), .ZN(n1071) );
  NAND3_X1 U1030 ( .A1(\SB1_2_13/i0_3 ), .A2(\SB1_2_13/i0[10] ), .A3(
        \SB1_2_13/i0[6] ), .ZN(\SB1_2_13/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U1031 ( .A1(\SB1_2_30/i0_4 ), .A2(\SB1_2_30/i0_3 ), .A3(
        \SB1_2_30/i1[9] ), .ZN(\SB1_2_30/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1033 ( .A1(\SB1_2_17/i1[9] ), .A2(\SB1_2_17/i1_7 ), .A3(
        \SB1_2_17/i0[10] ), .ZN(\SB1_2_17/Component_Function_3/NAND4_in[2] )
         );
  NAND3_X1 U1040 ( .A1(\SB1_2_9/i0[10] ), .A2(\SB1_2_9/i0[9] ), .A3(
        \SB1_2_9/i0_3 ), .ZN(n6458) );
  NAND3_X1 U1044 ( .A1(\SB1_2_8/i0_0 ), .A2(\SB1_2_8/i0[10] ), .A3(
        \SB1_2_8/i0[6] ), .ZN(\SB1_2_8/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1045 ( .A1(\SB1_2_18/i0_0 ), .A2(\SB1_2_18/i1_5 ), .A3(
        \SB1_2_18/i0_4 ), .ZN(\SB1_2_18/Component_Function_2/NAND4_in[3] ) );
  NAND2_X1 U1048 ( .A1(\SB1_2_16/i0[10] ), .A2(\SB1_2_16/i0[9] ), .ZN(
        \SB1_2_16/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U1053 ( .A1(\SB1_2_2/i0_0 ), .A2(\SB1_2_2/i0_3 ), .A3(
        \SB1_2_2/i0_4 ), .ZN(\SB1_2_2/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1054 ( .A1(\SB1_2_4/i0[6] ), .A2(\SB1_2_4/i0[9] ), .A3(
        \SB1_2_4/i1_5 ), .ZN(n5979) );
  NAND3_X1 U1057 ( .A1(\SB1_2_9/i0[6] ), .A2(\SB1_2_9/i0[9] ), .A3(
        \SB1_2_9/i1_5 ), .ZN(n6223) );
  NAND3_X1 U1059 ( .A1(\SB1_2_16/i0[10] ), .A2(\SB1_2_16/i0[6] ), .A3(
        \RI1[2][95] ), .ZN(\SB1_2_16/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U1065 ( .A1(\SB1_2_9/i1_7 ), .A2(\SB1_2_9/i0_3 ), .A3(
        \SB1_2_9/i0[8] ), .ZN(\SB1_2_9/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U1073 ( .A1(\SB1_2_21/i0[9] ), .A2(\SB1_2_21/i0[6] ), .A3(
        \SB1_2_21/i0_4 ), .ZN(n5000) );
  NAND2_X1 U1075 ( .A1(\SB1_2_16/i3[0] ), .A2(\SB1_2_16/i0_0 ), .ZN(
        \SB1_2_16/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U1076 ( .A1(\SB1_2_5/i0[6] ), .A2(\SB1_2_5/i0[9] ), .A3(
        \SB1_2_5/i1_5 ), .ZN(n5674) );
  NAND3_X1 U1081 ( .A1(\SB1_2_15/i0[10] ), .A2(\SB1_2_15/i1[9] ), .A3(
        \SB1_2_15/i1_7 ), .ZN(n5941) );
  NAND3_X1 U1086 ( .A1(\SB1_2_15/i0_4 ), .A2(\SB1_2_15/i0_0 ), .A3(
        \SB1_2_15/i1_5 ), .ZN(n5314) );
  NAND3_X1 U1088 ( .A1(\SB1_2_23/i0_4 ), .A2(\SB1_2_23/i0_3 ), .A3(
        \SB1_2_23/i0_0 ), .ZN(n6363) );
  NAND3_X1 U1092 ( .A1(\SB1_2_30/i0_3 ), .A2(\SB1_2_30/i0[8] ), .A3(
        \SB1_2_30/i1_7 ), .ZN(\SB1_2_30/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U1095 ( .A1(\SB1_2_14/i0[8] ), .A2(\SB1_2_14/i0_4 ), .A3(
        \SB1_2_14/i1_7 ), .ZN(n5984) );
  NAND3_X1 U1097 ( .A1(\SB1_2_13/i1_7 ), .A2(\SB1_2_13/i0_0 ), .A3(
        \SB1_2_13/i3[0] ), .ZN(\SB1_2_13/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U1101 ( .A1(\SB1_2_0/i0_4 ), .A2(\SB1_2_0/i0_0 ), .A3(
        \SB1_2_0/i0_3 ), .ZN(n6463) );
  NAND3_X1 U1106 ( .A1(\SB1_2_18/i0_0 ), .A2(\SB1_2_18/i3[0] ), .A3(
        \SB1_2_18/i1_7 ), .ZN(\SB1_2_18/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U1109 ( .A1(\SB1_2_3/i0_0 ), .A2(\SB1_2_3/i1_7 ), .A3(
        \SB1_2_3/i3[0] ), .ZN(n5263) );
  NAND3_X1 U1111 ( .A1(\SB1_2_5/i0[8] ), .A2(\SB1_2_5/i3[0] ), .A3(
        \SB1_2_5/i1_5 ), .ZN(n5452) );
  NAND3_X1 U1118 ( .A1(\SB1_2_12/i0_0 ), .A2(\SB1_2_12/i1_7 ), .A3(
        \SB1_2_12/i3[0] ), .ZN(n5709) );
  NAND3_X1 U1120 ( .A1(\SB1_2_28/i0_0 ), .A2(\SB1_2_28/i0_3 ), .A3(
        \SB1_2_28/i0_4 ), .ZN(\SB1_2_28/Component_Function_3/NAND4_in[1] ) );
  INV_X1 U1123 ( .I(\MC_ARK_ARC_1_1/buf_output[108] ), .ZN(\SB1_2_13/i3[0] )
         );
  BUF_X2 U1138 ( .I(\MC_ARK_ARC_1_1/buf_output[31] ), .Z(\SB1_2_26/i0[6] ) );
  NAND3_X1 U1142 ( .A1(\SB1_2_28/i0[10] ), .A2(\SB1_2_28/i0_0 ), .A3(
        \SB1_2_28/i0[6] ), .ZN(\SB1_2_28/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1143 ( .A1(\SB1_2_4/i1_5 ), .A2(\SB1_2_4/i0[8] ), .A3(
        \SB1_2_4/i3[0] ), .ZN(n5986) );
  NAND3_X1 U1145 ( .A1(\SB1_2_11/i0_4 ), .A2(\SB1_2_11/i1[9] ), .A3(
        \SB1_2_11/i1_5 ), .ZN(n1713) );
  INV_X1 U1146 ( .I(\MC_ARK_ARC_1_1/buf_output[174] ), .ZN(\SB1_2_2/i3[0] ) );
  NAND3_X1 U1147 ( .A1(\SB2_1_15/i0_3 ), .A2(\SB2_1_15/i0_4 ), .A3(
        \SB2_1_15/i1[9] ), .ZN(n5485) );
  NAND3_X1 U1158 ( .A1(\SB2_1_15/i0[9] ), .A2(\SB2_1_15/i0_3 ), .A3(
        \SB2_1_15/i0[8] ), .ZN(n5693) );
  NAND3_X1 U1163 ( .A1(\SB2_1_23/i0_3 ), .A2(\SB2_1_23/i1_7 ), .A3(
        \SB2_1_23/i0[8] ), .ZN(\SB2_1_23/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U1169 ( .A1(\SB2_1_15/i0[9] ), .A2(\SB2_1_15/i0_3 ), .A3(
        \SB2_1_15/i0[10] ), .ZN(\SB2_1_15/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U1171 ( .A1(\SB2_1_16/i0[10] ), .A2(\SB2_1_16/i0_4 ), .A3(
        \SB2_1_16/i0_3 ), .ZN(\SB2_1_16/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U1172 ( .A1(\SB2_1_5/i0_0 ), .A2(\SB2_1_5/i1_5 ), .A3(
        \SB1_1_6/buf_output[4] ), .ZN(n5364) );
  NAND3_X1 U1173 ( .A1(\SB2_1_8/i0_0 ), .A2(\SB2_1_8/i0[10] ), .A3(
        \SB2_1_8/i0[6] ), .ZN(n3723) );
  NAND3_X1 U1174 ( .A1(\SB2_1_29/i0[9] ), .A2(\SB2_1_29/i1_5 ), .A3(
        \SB2_1_29/i0[6] ), .ZN(n1632) );
  NAND3_X1 U1175 ( .A1(\SB2_1_23/i1[9] ), .A2(\SB2_1_23/i0_3 ), .A3(
        \SB2_1_23/i0[6] ), .ZN(\SB2_1_23/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U1176 ( .A1(\SB2_1_20/i0[9] ), .A2(\SB2_1_20/i0_4 ), .A3(
        \SB2_1_20/i0[6] ), .ZN(n5217) );
  NAND3_X1 U1184 ( .A1(\SB2_1_10/i0[6] ), .A2(\SB2_1_10/i0[7] ), .A3(
        \SB2_1_10/i0[8] ), .ZN(\SB2_1_10/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U1186 ( .A1(\SB2_1_16/i0[6] ), .A2(\SB2_1_16/i1_5 ), .A3(
        \SB2_1_16/i0[9] ), .ZN(\SB2_1_16/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1192 ( .A1(\SB2_1_6/i0[10] ), .A2(\SB2_1_6/i1[9] ), .A3(
        \SB2_1_6/i1_5 ), .ZN(\SB2_1_6/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U1194 ( .A1(\SB2_1_4/i0_3 ), .A2(\SB2_1_4/i0[9] ), .A3(
        \SB2_1_4/i0[8] ), .ZN(n6012) );
  NAND3_X1 U1197 ( .A1(\SB2_1_22/i0_4 ), .A2(\SB2_1_22/i1_7 ), .A3(
        \SB2_1_22/i0[8] ), .ZN(\SB2_1_22/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U1199 ( .A1(\SB2_1_28/i3[0] ), .A2(\SB2_1_28/i0[8] ), .A3(
        \SB2_1_28/i1_5 ), .ZN(n6440) );
  NAND3_X1 U1204 ( .A1(\SB2_1_19/i0[10] ), .A2(n1396), .A3(\SB2_1_19/i1_7 ), 
        .ZN(\SB2_1_19/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U1205 ( .A1(\SB2_1_9/i0_3 ), .A2(\SB2_1_9/i0[6] ), .A3(
        \SB2_1_9/i1[9] ), .ZN(n3982) );
  NAND3_X1 U1208 ( .A1(\SB2_1_3/i0_0 ), .A2(\SB2_1_3/i3[0] ), .A3(
        \SB2_1_3/i1_7 ), .ZN(\SB2_1_3/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U1212 ( .A1(\SB2_1_24/i0[10] ), .A2(\SB2_1_24/i0_3 ), .A3(
        \SB2_1_24/i0[9] ), .ZN(n4543) );
  NAND3_X1 U1213 ( .A1(\SB2_1_31/i0_0 ), .A2(\SB2_1_31/i0[8] ), .A3(
        \SB2_1_31/i0[9] ), .ZN(n5151) );
  NAND3_X1 U1214 ( .A1(\SB2_1_3/i1[9] ), .A2(n5208), .A3(\SB2_1_3/i1_5 ), .ZN(
        n5958) );
  NAND3_X1 U1215 ( .A1(\SB2_1_29/i0[10] ), .A2(\SB2_1_29/i0[9] ), .A3(
        \SB2_1_29/i0_3 ), .ZN(n5304) );
  INV_X1 U1220 ( .I(\SB1_1_6/buf_output[1] ), .ZN(\SB2_1_2/i1_7 ) );
  INV_X1 U1222 ( .I(\SB1_1_7/buf_output[1] ), .ZN(\SB2_1_3/i1_7 ) );
  INV_X1 U1229 ( .I(\SB2_1_3/i0_4 ), .ZN(\SB2_1_3/i0[7] ) );
  INV_X1 U1231 ( .I(\SB1_1_8/buf_output[1] ), .ZN(\SB2_1_4/i1_7 ) );
  NAND3_X1 U1232 ( .A1(\SB2_1_13/i0_3 ), .A2(\SB2_1_13/i0_4 ), .A3(
        \SB2_1_13/i1[9] ), .ZN(n990) );
  NAND2_X1 U1234 ( .A1(\SB2_1_5/i0_0 ), .A2(\SB2_1_5/i3[0] ), .ZN(n5938) );
  INV_X2 U1236 ( .I(\SB2_1_0/i0[7] ), .ZN(n2687) );
  NAND3_X1 U1238 ( .A1(\SB2_1_9/i3[0] ), .A2(\SB2_1_9/i0[8] ), .A3(
        \SB2_1_9/i1_5 ), .ZN(\SB2_1_9/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U1239 ( .A1(\SB2_1_18/i0_0 ), .A2(\SB2_1_18/i0[10] ), .A3(
        \SB1_1_22/buf_output[1] ), .ZN(n5230) );
  CLKBUF_X2 U1241 ( .I(\SB1_1_29/buf_output[0] ), .Z(\SB2_1_24/i0[9] ) );
  CLKBUF_X4 U1242 ( .I(\SB1_1_31/buf_output[5] ), .Z(\SB2_1_31/i0_3 ) );
  NAND3_X1 U1243 ( .A1(\SB1_1_20/i0_3 ), .A2(\SB1_1_20/i0_4 ), .A3(
        \SB1_1_20/i1[9] ), .ZN(n5299) );
  NAND3_X1 U1247 ( .A1(\SB1_1_3/i0[6] ), .A2(\SB1_1_3/i0_4 ), .A3(
        \SB1_1_3/i0[9] ), .ZN(n1524) );
  NAND3_X1 U1249 ( .A1(\SB1_1_8/i0[10] ), .A2(\SB1_1_8/i0[6] ), .A3(
        \SB1_1_8/i0_0 ), .ZN(\SB1_1_8/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1250 ( .A1(\SB1_1_30/i0_0 ), .A2(\SB1_1_30/i1_5 ), .A3(
        \SB1_1_30/i0_4 ), .ZN(n1414) );
  NAND3_X1 U1258 ( .A1(\SB1_1_30/i0[6] ), .A2(\SB1_1_30/i1_5 ), .A3(
        \SB1_1_30/i0[9] ), .ZN(\SB1_1_30/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1259 ( .A1(\SB1_1_14/i0[9] ), .A2(\SB1_1_14/i0[6] ), .A3(
        \SB1_1_14/i0_4 ), .ZN(n6349) );
  NAND3_X1 U1264 ( .A1(\SB1_1_14/i0[10] ), .A2(\SB1_1_14/i0[6] ), .A3(
        \SB1_1_14/i0_3 ), .ZN(n5201) );
  NAND2_X1 U1271 ( .A1(\SB1_1_1/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_1_1/Component_Function_4/NAND4_in[1] ), .ZN(n6524) );
  NAND3_X1 U1278 ( .A1(\SB1_1_9/i0_3 ), .A2(\SB1_1_9/i0[10] ), .A3(
        \SB1_1_9/i0[9] ), .ZN(\SB1_1_9/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1279 ( .A1(\SB1_1_28/i1[9] ), .A2(\SB1_1_28/i1_5 ), .A3(
        \SB1_1_28/i0_4 ), .ZN(\SB1_1_28/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U1283 ( .A1(\SB1_1_29/i0_0 ), .A2(\SB1_1_29/i0_4 ), .A3(
        \SB1_1_29/i1_5 ), .ZN(n5408) );
  NAND3_X1 U1286 ( .A1(\SB1_1_16/i0[8] ), .A2(\SB1_1_16/i0[7] ), .A3(
        \SB1_1_16/i0[6] ), .ZN(\SB1_1_16/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U1288 ( .A1(\SB1_1_2/i0[10] ), .A2(\SB1_1_2/i1[9] ), .A3(
        \SB1_1_2/i1_7 ), .ZN(\SB1_1_2/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U1289 ( .A1(\SB1_1_28/i0[10] ), .A2(\SB1_1_28/i1[9] ), .A3(
        \SB1_1_28/i1_7 ), .ZN(\SB1_1_28/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U1290 ( .A1(\SB1_1_22/i0[10] ), .A2(\SB1_1_22/i1[9] ), .A3(
        \SB1_1_22/i1_7 ), .ZN(n1514) );
  NAND3_X1 U1291 ( .A1(\SB1_1_24/i0[10] ), .A2(\SB1_1_24/i1[9] ), .A3(
        \SB1_1_24/i1_7 ), .ZN(n5955) );
  NAND2_X1 U1296 ( .A1(\SB1_1_20/i0[10] ), .A2(\SB1_1_20/i0[9] ), .ZN(n4001)
         );
  NAND3_X1 U1298 ( .A1(\SB1_1_11/i0_0 ), .A2(\SB1_1_11/i1_5 ), .A3(
        \SB1_1_11/i0_4 ), .ZN(n5788) );
  NAND3_X1 U1299 ( .A1(\SB1_1_11/i0[10] ), .A2(\SB1_1_11/i0[6] ), .A3(
        \SB1_1_11/i0_3 ), .ZN(n5785) );
  NAND3_X1 U1306 ( .A1(\SB1_1_23/i0_0 ), .A2(\SB1_1_23/i3[0] ), .A3(
        \SB1_1_23/i1_7 ), .ZN(\SB1_1_23/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U1316 ( .A1(\SB1_1_9/i0[6] ), .A2(\SB1_1_9/i0_4 ), .A3(
        \SB1_1_9/i0[9] ), .ZN(n2202) );
  NAND3_X1 U1317 ( .A1(\SB1_1_9/i0[6] ), .A2(\SB1_1_9/i0[8] ), .A3(
        \SB1_1_9/i0[7] ), .ZN(\SB1_1_9/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U1320 ( .A1(\SB1_1_9/i0[8] ), .A2(\SB1_1_9/i3[0] ), .A3(
        \SB1_1_9/i1_5 ), .ZN(n6107) );
  NAND2_X1 U1322 ( .A1(n1358), .A2(\SB1_1_0/Component_Function_4/NAND4_in[3] ), 
        .ZN(n5827) );
  NAND3_X1 U1325 ( .A1(\SB1_1_9/i0[6] ), .A2(\SB1_1_9/i1_5 ), .A3(
        \SB1_1_9/i0[9] ), .ZN(\SB1_1_9/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U1326 ( .A1(\SB1_1_4/i0_4 ), .A2(\SB1_1_4/i0[6] ), .A3(
        \SB1_1_4/i0[9] ), .ZN(n2993) );
  NAND3_X1 U1331 ( .A1(\SB1_1_23/i0[9] ), .A2(\SB1_1_23/i1_5 ), .A3(
        \SB1_1_23/i0[6] ), .ZN(\SB1_1_23/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 U1332 ( .A1(\SB1_1_7/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_1_7/Component_Function_2/NAND4_in[0] ), .ZN(n5447) );
  NAND3_X1 U1340 ( .A1(\SB1_1_29/i0[9] ), .A2(\SB1_1_29/i1_5 ), .A3(
        \SB1_1_29/i0[6] ), .ZN(n5969) );
  NAND3_X1 U1341 ( .A1(\SB1_1_23/i0[8] ), .A2(\SB1_1_23/i1_7 ), .A3(
        \SB1_1_23/i0_4 ), .ZN(n2582) );
  NAND3_X1 U1343 ( .A1(\SB1_1_30/i0_3 ), .A2(\SB1_1_30/i0_0 ), .A3(
        \SB1_1_30/i0[7] ), .ZN(n6251) );
  NAND3_X1 U1345 ( .A1(\SB1_1_12/i0[9] ), .A2(\SB1_1_12/i0_3 ), .A3(
        \SB1_1_12/i0[8] ), .ZN(n1627) );
  NAND3_X1 U1346 ( .A1(\SB1_1_20/i0[6] ), .A2(\SB1_1_20/i1_5 ), .A3(
        \SB1_1_20/i0[9] ), .ZN(n6233) );
  NAND3_X1 U1347 ( .A1(\SB1_1_15/i0_3 ), .A2(\SB1_1_15/i0_0 ), .A3(
        \MC_ARK_ARC_1_0/buf_output[100] ), .ZN(
        \SB1_1_15/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1356 ( .A1(\SB1_1_13/i0_0 ), .A2(\SB1_1_13/i1_5 ), .A3(
        \SB1_1_13/i0_4 ), .ZN(n6058) );
  NAND3_X1 U1357 ( .A1(\SB1_1_10/i1[9] ), .A2(\SB1_1_10/i0_4 ), .A3(
        \SB1_1_10/i1_5 ), .ZN(n5646) );
  NAND3_X1 U1369 ( .A1(\SB1_1_26/i0_0 ), .A2(\SB1_1_26/i1_5 ), .A3(
        \SB1_1_26/i0_4 ), .ZN(n5016) );
  NAND3_X1 U1376 ( .A1(\SB1_1_3/i0[10] ), .A2(\SB1_1_3/i0_3 ), .A3(
        \SB1_1_3/i0[9] ), .ZN(n5206) );
  NAND3_X1 U1378 ( .A1(\SB1_1_29/i0[9] ), .A2(\SB1_1_29/i0[6] ), .A3(
        \SB1_1_29/i0_4 ), .ZN(n5918) );
  NAND3_X1 U1380 ( .A1(\SB1_1_7/i0_0 ), .A2(\SB1_1_7/i0[9] ), .A3(
        \SB1_1_7/i0[8] ), .ZN(n5819) );
  NAND3_X1 U1381 ( .A1(\SB1_1_21/i0[8] ), .A2(\SB1_1_21/i0_3 ), .A3(
        \SB1_1_21/i0[9] ), .ZN(n2155) );
  NAND3_X1 U1386 ( .A1(\SB1_1_31/i0[8] ), .A2(\SB1_1_31/i3[0] ), .A3(
        \SB1_1_31/i1_5 ), .ZN(\SB1_1_31/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U1389 ( .A1(\SB1_1_6/i0_0 ), .A2(\SB1_1_6/i0[9] ), .A3(
        \SB1_1_6/i0[8] ), .ZN(n6104) );
  NAND3_X1 U1391 ( .A1(\SB1_1_30/i0_0 ), .A2(\SB1_1_30/i1_7 ), .A3(
        \SB1_1_30/i3[0] ), .ZN(n3366) );
  BUF_X2 U1392 ( .I(\MC_ARK_ARC_1_0/buf_output[94] ), .Z(\SB1_1_16/i0_4 ) );
  BUF_X2 U1393 ( .I(\MC_ARK_ARC_1_0/buf_output[24] ), .Z(\SB1_1_27/i0[9] ) );
  BUF_X2 U1394 ( .I(\SB2_0_30/buf_output[1] ), .Z(\RI5[0][31] ) );
  BUF_X2 U1396 ( .I(Key[97]), .Z(n187) );
  NAND3_X1 U1398 ( .A1(\SB2_0_1/i0[10] ), .A2(\SB2_0_1/i0_3 ), .A3(
        \SB2_0_1/i0_4 ), .ZN(\SB2_0_1/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U1401 ( .A1(\SB2_0_7/i0[10] ), .A2(\SB2_0_7/i0_3 ), .A3(
        \SB1_0_8/buf_output[4] ), .ZN(n6011) );
  NAND3_X1 U1405 ( .A1(\SB2_0_10/i0[10] ), .A2(\SB2_0_10/i0_3 ), .A3(n571), 
        .ZN(n6165) );
  NAND3_X1 U1406 ( .A1(n5054), .A2(\SB2_0_1/i0[8] ), .A3(\SB2_0_1/i0[6] ), 
        .ZN(n2536) );
  NAND3_X1 U1415 ( .A1(\RI3[0][155] ), .A2(n2765), .A3(\RI3[0][154] ), .ZN(
        \SB2_0_6/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U1416 ( .A1(\SB2_0_28/i0[10] ), .A2(\SB2_0_28/i1[9] ), .A3(
        \SB2_0_28/i1_7 ), .ZN(\SB2_0_28/Component_Function_3/NAND4_in[2] ) );
  NAND2_X1 U1417 ( .A1(\SB2_0_1/i0[9] ), .A2(\SB2_0_1/i0[10] ), .ZN(
        \SB2_0_1/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U1421 ( .A1(\SB2_0_11/i0_3 ), .A2(\SB2_0_11/i0[10] ), .A3(n1911), 
        .ZN(\SB2_0_11/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1424 ( .A1(\SB2_0_5/i0_3 ), .A2(\SB2_0_5/i0[10] ), .A3(
        \SB2_0_5/i0[6] ), .ZN(n3770) );
  NAND3_X1 U1425 ( .A1(\SB2_0_26/i0_0 ), .A2(\SB2_0_26/i0[10] ), .A3(
        \SB2_0_26/i0[6] ), .ZN(n5872) );
  NAND3_X1 U1431 ( .A1(\SB2_0_14/i0[6] ), .A2(\SB2_0_14/i0[9] ), .A3(
        \SB2_0_14/i1_5 ), .ZN(n5796) );
  NAND3_X1 U1433 ( .A1(\SB2_0_1/i0[9] ), .A2(\SB2_0_1/i1_5 ), .A3(
        \SB2_0_1/i0[6] ), .ZN(n5412) );
  NAND3_X1 U1439 ( .A1(\RI3[0][10] ), .A2(\SB2_0_30/i1_7 ), .A3(
        \SB2_0_30/i0[8] ), .ZN(n6356) );
  NAND3_X1 U1440 ( .A1(\SB2_0_15/i0_0 ), .A2(\RI3[0][100] ), .A3(
        \SB2_0_15/i1_5 ), .ZN(n5805) );
  NAND3_X1 U1441 ( .A1(\SB2_0_2/i0_3 ), .A2(\RI3[0][178] ), .A3(
        \SB2_0_2/i0[10] ), .ZN(n5297) );
  NAND3_X1 U1454 ( .A1(\SB2_0_12/i3[0] ), .A2(\SB2_0_12/i1_5 ), .A3(
        \SB2_0_12/i0[8] ), .ZN(n4910) );
  NAND3_X1 U1457 ( .A1(\SB2_0_20/i0_3 ), .A2(\SB2_0_20/i0_4 ), .A3(
        \SB2_0_20/i0[10] ), .ZN(\SB2_0_20/Component_Function_0/NAND4_in[2] )
         );
  NAND3_X1 U1460 ( .A1(\SB2_0_7/i0[10] ), .A2(\SB2_0_7/i0[9] ), .A3(
        \SB2_0_7/i0_3 ), .ZN(n6000) );
  NAND3_X1 U1468 ( .A1(\SB2_0_1/i0_3 ), .A2(\SB2_0_1/i0_0 ), .A3(
        \SB2_0_1/i0_4 ), .ZN(\SB2_0_1/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1482 ( .A1(\RI3[0][191] ), .A2(\SB2_0_0/i0_0 ), .A3(\RI3[0][190] ), 
        .ZN(n5854) );
  NAND3_X1 U1485 ( .A1(\SB2_0_28/i0[6] ), .A2(\SB2_0_28/i1_5 ), .A3(
        \RI3[0][18] ), .ZN(n5613) );
  NAND2_X1 U1487 ( .A1(\RI3[0][106] ), .A2(n4761), .ZN(n5754) );
  NAND3_X1 U1488 ( .A1(\SB2_0_2/i0[8] ), .A2(\SB2_0_2/i0_3 ), .A3(
        \SB2_0_2/i0[9] ), .ZN(n1958) );
  INV_X1 U1489 ( .I(\SB1_0_23/buf_output[1] ), .ZN(\SB2_0_19/i1_7 ) );
  NAND3_X1 U1493 ( .A1(\RI3[0][155] ), .A2(\RI3[0][154] ), .A3(\SB2_0_6/i0_0 ), 
        .ZN(\SB2_0_6/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1494 ( .A1(\SB2_0_5/i0[10] ), .A2(n3689), .A3(\SB2_0_5/i1_7 ), 
        .ZN(n6202) );
  NAND3_X1 U1500 ( .A1(\SB2_0_1/i0[9] ), .A2(\SB2_0_1/i0_3 ), .A3(
        \SB2_0_1/i0[10] ), .ZN(\SB2_0_1/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1505 ( .A1(\SB2_0_15/i0[9] ), .A2(\SB2_0_15/i0_3 ), .A3(
        \SB2_0_15/i0[10] ), .ZN(n3501) );
  NAND3_X1 U1507 ( .A1(\SB2_0_5/i0_3 ), .A2(n3689), .A3(\SB2_0_5/i0[6] ), .ZN(
        n5377) );
  INV_X1 U1520 ( .I(\RI3[0][91] ), .ZN(\SB2_0_16/i1_7 ) );
  INV_X2 U1523 ( .I(\SB2_0_6/i0[7] ), .ZN(\RI3[0][154] ) );
  INV_X2 U1527 ( .I(\SB2_0_19/i0[7] ), .ZN(\RI3[0][76] ) );
  NAND3_X1 U1529 ( .A1(\SB2_0_16/i0[10] ), .A2(\SB2_0_16/i0_0 ), .A3(
        \SB2_0_16/i0[6] ), .ZN(n5530) );
  NAND3_X1 U1534 ( .A1(\SB2_0_23/i0[10] ), .A2(\SB2_0_23/i0[6] ), .A3(
        \SB2_0_23/i0_0 ), .ZN(n5849) );
  INV_X2 U1535 ( .I(\SB2_0_5/i0[7] ), .ZN(\RI3[0][160] ) );
  NAND2_X1 U1541 ( .A1(\SB1_0_31/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_0_31/Component_Function_4/NAND4_in[0] ), .ZN(n6501) );
  NAND3_X1 U1542 ( .A1(\SB1_0_6/i0[10] ), .A2(\SB1_0_6/i1_5 ), .A3(
        \SB1_0_6/i1[9] ), .ZN(\SB1_0_6/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U1543 ( .A1(\SB1_0_29/i0_4 ), .A2(\SB1_0_29/i1_5 ), .A3(
        \SB1_0_29/i0_0 ), .ZN(n5871) );
  NAND3_X1 U1544 ( .A1(\SB1_0_20/i1_5 ), .A2(\SB1_0_20/i0[8] ), .A3(
        \SB1_0_20/i3[0] ), .ZN(n5207) );
  NAND2_X1 U1545 ( .A1(\SB1_0_4/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_0_4/Component_Function_3/NAND4_in[3] ), .ZN(n6436) );
  NAND2_X1 U1546 ( .A1(n1667), .A2(n6479), .ZN(n5657) );
  NAND2_X1 U1550 ( .A1(\SB1_0_10/Component_Function_4/NAND4_in[0] ), .A2(n5341), .ZN(n4641) );
  NAND3_X1 U1553 ( .A1(\SB1_0_9/i0_0 ), .A2(\SB1_0_9/i0[6] ), .A3(
        \SB1_0_9/i0[10] ), .ZN(\SB1_0_9/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1554 ( .A1(\SB1_0_23/i0_0 ), .A2(\SB1_0_23/i0[6] ), .A3(
        \SB1_0_23/i0[10] ), .ZN(\SB1_0_23/Component_Function_5/NAND4_in[1] )
         );
  NAND3_X1 U1557 ( .A1(\SB1_0_20/i0[8] ), .A2(\SB1_0_20/i0_4 ), .A3(
        \SB1_0_20/i1_7 ), .ZN(n6350) );
  NAND3_X1 U1560 ( .A1(\SB1_0_25/i0_0 ), .A2(\SB1_0_25/i1_5 ), .A3(
        \SB1_0_25/i0_4 ), .ZN(n2629) );
  NAND3_X1 U1561 ( .A1(\SB1_0_8/i0_3 ), .A2(\SB1_0_8/i0[10] ), .A3(
        \SB1_0_8/i0[6] ), .ZN(\SB1_0_8/Component_Function_2/NAND4_in[1] ) );
  BUF_X2 U1563 ( .I(n263), .Z(\SB1_0_25/i0[9] ) );
  NAND3_X1 U1564 ( .A1(\SB1_0_6/i0_3 ), .A2(\SB1_0_6/i0[10] ), .A3(
        \SB1_0_6/i0[9] ), .ZN(n6225) );
  NAND3_X1 U1567 ( .A1(\SB1_0_10/i0_0 ), .A2(\SB1_0_10/i1_7 ), .A3(
        \SB1_0_10/i3[0] ), .ZN(n5341) );
  BUF_X4 U1573 ( .I(\MC_ARK_ARC_1_1/buf_output[56] ), .Z(\SB1_2_22/i0_0 ) );
  NAND2_X2 U1574 ( .A1(\SB2_3_23/i0_0 ), .A2(\SB2_3_23/i3[0] ), .ZN(n4823) );
  NAND3_X2 U1575 ( .A1(\SB1_3_24/i0[10] ), .A2(\SB1_3_24/i1[9] ), .A3(
        \SB1_3_24/i1_5 ), .ZN(n4338) );
  NAND3_X2 U1576 ( .A1(\SB2_1_0/i0_3 ), .A2(\SB2_1_0/i0[8] ), .A3(
        \SB2_1_0/i0[9] ), .ZN(\SB2_1_0/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 U1577 ( .I(\SB1_1_28/buf_output[4] ), .Z(\SB2_1_27/i0_4 ) );
  BUF_X4 U1578 ( .I(\SB1_2_28/buf_output[5] ), .Z(\SB2_2_28/i0_3 ) );
  BUF_X2 U1579 ( .I(\MC_ARK_ARC_1_2/buf_output[115] ), .Z(\SB1_3_12/i0[6] ) );
  NAND3_X2 U1581 ( .A1(\SB1_1_7/i0_3 ), .A2(\SB1_1_7/i1_7 ), .A3(
        \SB1_1_7/i0[8] ), .ZN(\SB1_1_7/Component_Function_1/NAND4_in[1] ) );
  NAND3_X2 U1583 ( .A1(\SB1_0_29/i0[10] ), .A2(\SB1_0_29/i0_3 ), .A3(
        \SB1_0_29/i0[6] ), .ZN(n4228) );
  NAND3_X2 U1589 ( .A1(\SB1_0_25/i0_3 ), .A2(\SB1_0_25/i0_0 ), .A3(
        \SB1_0_25/i0_4 ), .ZN(\SB1_0_25/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U1590 ( .A1(\SB2_0_13/i0_4 ), .A2(\SB2_0_13/i0_3 ), .A3(
        \SB2_0_13/i1[9] ), .ZN(\SB2_0_13/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U1591 ( .A1(\SB1_0_26/i0_0 ), .A2(\SB1_0_26/i0_3 ), .A3(
        \SB1_0_26/i0_4 ), .ZN(\SB1_0_26/Component_Function_3/NAND4_in[1] ) );
  INV_X1 U1592 ( .I(\MC_ARK_ARC_1_3/buf_output[121] ), .ZN(\SB3_11/i1_7 ) );
  BUF_X2 U1593 ( .I(\MC_ARK_ARC_1_3/buf_output[121] ), .Z(\SB3_11/i0[6] ) );
  NAND3_X1 U1603 ( .A1(\SB3_10/i0[9] ), .A2(\SB3_10/i0[8] ), .A3(\SB3_10/i0_3 ), .ZN(n5733) );
  NAND3_X1 U1613 ( .A1(\SB3_6/i0[9] ), .A2(\SB3_6/i0[6] ), .A3(\RI1[4][154] ), 
        .ZN(\SB3_6/Component_Function_5/NAND4_in[3] ) );
  INV_X1 U1622 ( .I(\MC_ARK_ARC_1_2/buf_output[146] ), .ZN(\SB1_3_7/i1[9] ) );
  BUF_X2 U1637 ( .I(\MC_ARK_ARC_1_2/buf_output[146] ), .Z(\SB1_3_7/i0_0 ) );
  NAND3_X1 U1639 ( .A1(\SB3_28/i0_3 ), .A2(\SB3_28/i0_0 ), .A3(\SB3_28/i0_4 ), 
        .ZN(\SB3_28/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U1640 ( .A1(\SB3_28/i1[9] ), .A2(\SB3_28/i1_5 ), .A3(\SB3_28/i0_4 ), 
        .ZN(\SB3_28/Component_Function_4/NAND4_in[3] ) );
  CLKBUF_X4 U1643 ( .I(\SB1_3_12/buf_output[2] ), .Z(\SB2_3_9/i0_0 ) );
  CLKBUF_X4 U1655 ( .I(\SB3_8/buf_output[5] ), .Z(\SB4_8/i0_3 ) );
  NAND2_X1 U1659 ( .A1(\SB3_6/Component_Function_2/NAND4_in[3] ), .A2(
        \SB3_6/Component_Function_2/NAND4_in[2] ), .ZN(n5004) );
  NAND3_X1 U1671 ( .A1(\RI1[4][155] ), .A2(\SB3_6/i0[8] ), .A3(\SB3_6/i0[9] ), 
        .ZN(\SB3_6/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1672 ( .A1(\SB2_2_10/i0_3 ), .A2(\SB2_2_10/i0[8] ), .A3(
        \SB2_2_10/i0[9] ), .ZN(\SB2_2_10/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1680 ( .A1(\SB3_9/i1[9] ), .A2(\SB3_9/i0_3 ), .A3(\SB3_9/i0[6] ), 
        .ZN(\SB3_9/Component_Function_3/NAND4_in[0] ) );
  BUF_X2 U1684 ( .I(\MC_ARK_ARC_1_1/buf_output[117] ), .Z(\SB1_2_12/i0[10] )
         );
  INV_X1 U1686 ( .I(\MC_ARK_ARC_1_1/buf_output[117] ), .ZN(\SB1_2_12/i0[8] )
         );
  CLKBUF_X2 U1691 ( .I(\MC_ARK_ARC_1_3/buf_datainput[90] ), .Z(n2895) );
  CLKBUF_X4 U1694 ( .I(\SB1_2_24/buf_output[4] ), .Z(\SB2_2_23/i0_4 ) );
  NAND3_X1 U1710 ( .A1(\SB4_30/i0[6] ), .A2(\SB4_30/i0_4 ), .A3(\SB4_30/i0[9] ), .ZN(\SB4_30/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U1715 ( .A1(\SB4_3/i0_3 ), .A2(n5495), .A3(\SB4_3/i0[9] ), .ZN(
        \SB4_3/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1716 ( .A1(\SB3_3/i0[10] ), .A2(\SB3_3/i1_7 ), .A3(\SB3_3/i1[9] ), 
        .ZN(n5068) );
  NAND3_X1 U1718 ( .A1(\SB1_3_14/i0_3 ), .A2(\SB1_3_14/i1[9] ), .A3(
        \SB1_3_14/i0_4 ), .ZN(n941) );
  NAND3_X1 U1719 ( .A1(\SB1_3_14/i0_0 ), .A2(\SB1_3_14/i0_3 ), .A3(
        \SB1_3_14/i0[7] ), .ZN(n667) );
  NAND3_X1 U1720 ( .A1(\SB1_3_14/i0_3 ), .A2(\SB1_3_14/i0[8] ), .A3(
        \SB1_3_14/i0[9] ), .ZN(\SB1_3_14/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U1721 ( .A1(\SB1_3_14/i0[9] ), .A2(\SB1_3_14/i0[10] ), .A3(
        \SB1_3_14/i0_3 ), .ZN(\SB1_3_14/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U1722 ( .A1(\SB1_3_14/i1[9] ), .A2(\SB1_3_14/i0_3 ), .A3(
        \SB1_3_14/i0[6] ), .ZN(\SB1_3_14/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U1724 ( .A1(\SB3_26/i0_0 ), .A2(\SB3_26/i0_4 ), .A3(\SB3_26/i0_3 ), 
        .ZN(n4208) );
  NAND3_X1 U1726 ( .A1(\SB3_26/i0_4 ), .A2(\SB3_26/i1[9] ), .A3(\SB3_26/i0_3 ), 
        .ZN(n3585) );
  BUF_X2 U1727 ( .I(\MC_ARK_ARC_1_3/buf_output[34] ), .Z(\SB3_26/i0_4 ) );
  INV_X1 U1729 ( .I(\MC_ARK_ARC_1_3/buf_output[129] ), .ZN(\SB3_10/i0[8] ) );
  BUF_X2 U1731 ( .I(\MC_ARK_ARC_1_3/buf_output[129] ), .Z(\SB3_10/i0[10] ) );
  CLKBUF_X4 U1736 ( .I(\MC_ARK_ARC_1_0/buf_output[22] ), .Z(\SB1_1_28/i0_4 )
         );
  BUF_X2 U1738 ( .I(\MC_ARK_ARC_1_0/buf_output[44] ), .Z(\SB1_1_24/i0_0 ) );
  INV_X1 U1742 ( .I(\MC_ARK_ARC_1_0/buf_output[44] ), .ZN(\SB1_1_24/i1[9] ) );
  OR3_X1 U1743 ( .A1(n5501), .A2(\MC_ARK_ARC_1_2/buf_output[132] ), .A3(
        \MC_ARK_ARC_1_2/buf_output[137] ), .Z(n1926) );
  NAND3_X1 U1745 ( .A1(\SB4_30/i0[10] ), .A2(n4751), .A3(\SB4_30/i1_7 ), .ZN(
        \SB4_30/Component_Function_3/NAND4_in[2] ) );
  NAND2_X1 U1748 ( .A1(\SB3_6/i0_0 ), .A2(\SB3_6/i3[0] ), .ZN(
        \SB3_6/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U1749 ( .A1(\SB3_6/i0_0 ), .A2(\SB3_6/i0[10] ), .A3(\SB3_6/i0[6] ), 
        .ZN(\SB3_6/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U1750 ( .A1(\SB2_3_1/i3[0] ), .A2(\SB2_3_1/i1_5 ), .A3(
        \SB2_3_1/i0[8] ), .ZN(n4682) );
  NAND2_X1 U1754 ( .A1(\SB2_3_1/i0[9] ), .A2(\SB2_3_1/i0[8] ), .ZN(n3279) );
  NAND3_X1 U1760 ( .A1(\SB2_3_1/i0_3 ), .A2(\SB2_3_1/i1_7 ), .A3(
        \SB2_3_1/i0[8] ), .ZN(\SB2_3_1/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U1764 ( .A1(\SB2_3_1/i0_4 ), .A2(\SB2_3_1/i1_7 ), .A3(
        \SB2_3_1/i0[8] ), .ZN(n5349) );
  NAND3_X1 U1765 ( .A1(\SB4_30/i0_4 ), .A2(\SB4_30/i1_7 ), .A3(\SB4_30/i0[8] ), 
        .ZN(\SB4_30/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U1767 ( .A1(\SB4_10/i0[10] ), .A2(\SB4_10/i1_7 ), .A3(n3653), .ZN(
        \SB4_10/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U1768 ( .A1(\SB1_3_7/i1_5 ), .A2(\SB1_3_7/i0[6] ), .A3(
        \SB1_3_7/i0[9] ), .ZN(\SB1_3_7/Component_Function_1/NAND4_in[2] ) );
  CLKBUF_X4 U1770 ( .I(\MC_ARK_ARC_1_2/buf_output[121] ), .Z(\SB1_3_11/i0[6] )
         );
  CLKBUF_X4 U1772 ( .I(\SB1_3_6/buf_output[2] ), .Z(\SB2_3_3/i0_0 ) );
  CLKBUF_X4 U1774 ( .I(\SB1_1_23/buf_output[3] ), .Z(\SB2_1_21/i0[10] ) );
  NAND3_X1 U1775 ( .A1(\SB2_3_19/i0[10] ), .A2(\SB2_3_19/i1_7 ), .A3(n5494), 
        .ZN(\SB2_3_19/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U1779 ( .A1(\SB2_3_19/i0_3 ), .A2(n5494), .A3(\SB2_3_19/i0_4 ), 
        .ZN(n4968) );
  NAND3_X1 U1781 ( .A1(\SB2_3_19/i0[10] ), .A2(\SB2_3_19/i1_5 ), .A3(n5494), 
        .ZN(\SB2_3_19/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U1783 ( .A1(\SB4_23/i0[10] ), .A2(\SB4_23/i0_3 ), .A3(
        \SB4_23/i0[6] ), .ZN(n1578) );
  CLKBUF_X2 U1786 ( .I(\SB3_11/buf_output[2] ), .Z(\SB4_8/i0_0 ) );
  INV_X1 U1787 ( .I(\RI1[4][59] ), .ZN(\SB3_22/i1_5 ) );
  BUF_X2 U1789 ( .I(\RI1[4][59] ), .Z(\SB3_22/i0_3 ) );
  NAND2_X1 U1790 ( .A1(n1079), .A2(\SB3_13/Component_Function_2/NAND4_in[0] ), 
        .ZN(n6395) );
  NAND3_X1 U1791 ( .A1(\SB2_1_8/i1[9] ), .A2(\SB2_1_8/i0_4 ), .A3(
        \SB2_1_8/i0_3 ), .ZN(\SB2_1_8/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U1795 ( .A1(\SB2_1_8/i1_5 ), .A2(\SB2_1_8/i0[10] ), .A3(
        \SB2_1_8/i1[9] ), .ZN(\SB2_1_8/Component_Function_2/NAND4_in[0] ) );
  NAND2_X1 U1796 ( .A1(\SB2_1_8/i0_3 ), .A2(\SB2_1_8/i1[9] ), .ZN(
        \SB2_1_8/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U1797 ( .A1(\SB2_1_8/i0[6] ), .A2(\SB2_1_8/i1[9] ), .A3(
        \SB2_1_8/i0_3 ), .ZN(\SB2_1_8/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U1801 ( .A1(\SB2_1_8/i0[10] ), .A2(\SB2_1_8/i1_7 ), .A3(
        \SB2_1_8/i1[9] ), .ZN(n5864) );
  NAND3_X1 U1821 ( .A1(\SB3_22/i0_4 ), .A2(\SB3_22/i0[9] ), .A3(\SB3_22/i0[6] ), .ZN(n6047) );
  NAND3_X1 U1822 ( .A1(\SB3_22/i1_5 ), .A2(\SB3_22/i0[6] ), .A3(\SB3_22/i0[9] ), .ZN(\SB3_22/Component_Function_1/NAND4_in[2] ) );
  NAND4_X1 U1823 ( .A1(\SB4_30/Component_Function_1/NAND4_in[2] ), .A2(
        \SB4_30/Component_Function_1/NAND4_in[3] ), .A3(
        \SB4_30/Component_Function_1/NAND4_in[1] ), .A4(
        \SB4_30/Component_Function_1/NAND4_in[0] ), .ZN(n5561) );
  CLKBUF_X4 U1825 ( .I(\RI1[4][41] ), .Z(\SB3_25/i0_3 ) );
  NAND3_X1 U1829 ( .A1(\SB3_26/i0[9] ), .A2(\SB3_26/i1_5 ), .A3(\SB3_26/i0[6] ), .ZN(\SB3_26/Component_Function_1/NAND4_in[2] ) );
  INV_X1 U1830 ( .I(\SB3_18/buf_output[1] ), .ZN(\SB4_14/i1_7 ) );
  BUF_X2 U1833 ( .I(\SB3_18/buf_output[1] ), .Z(\SB4_14/i0[6] ) );
  NAND3_X1 U1836 ( .A1(\SB3_3/i0[10] ), .A2(\SB3_3/i0[6] ), .A3(\SB3_3/i0_3 ), 
        .ZN(n1687) );
  NAND3_X1 U1838 ( .A1(\SB3_3/i0_4 ), .A2(\SB3_3/i0_0 ), .A3(\SB3_3/i0_3 ), 
        .ZN(n4993) );
  INV_X1 U1839 ( .I(\MC_ARK_ARC_1_2/buf_output[191] ), .ZN(\SB1_3_0/i1_5 ) );
  NAND3_X1 U1840 ( .A1(\SB2_3_12/i0_4 ), .A2(\SB2_3_12/i0_3 ), .A3(
        \SB2_3_12/i0_0 ), .ZN(\SB2_3_12/Component_Function_3/NAND4_in[1] ) );
  NAND2_X1 U1843 ( .A1(\SB2_3_12/i3[0] ), .A2(\SB2_3_12/i0_0 ), .ZN(n3973) );
  NAND3_X1 U1844 ( .A1(\SB2_3_12/i0_4 ), .A2(\SB2_3_12/i0_0 ), .A3(
        \SB2_3_12/i1_5 ), .ZN(n6536) );
  BUF_X2 U1846 ( .I(\SB3_21/buf_output[0] ), .Z(\SB4_16/i0[9] ) );
  INV_X1 U1848 ( .I(\MC_ARK_ARC_1_3/buf_output[114] ), .ZN(\SB3_12/i3[0] ) );
  BUF_X2 U1850 ( .I(\MC_ARK_ARC_1_3/buf_output[114] ), .Z(\SB3_12/i0[9] ) );
  INV_X1 U1855 ( .I(\SB3_14/buf_output[5] ), .ZN(\SB4_14/i1_5 ) );
  BUF_X2 U1856 ( .I(\SB3_12/buf_output[1] ), .Z(\SB4_8/i0[6] ) );
  CLKBUF_X4 U1859 ( .I(\SB1_3_14/buf_output[2] ), .Z(\SB2_3_11/i0_0 ) );
  NAND3_X1 U1861 ( .A1(\SB3_22/i1_5 ), .A2(\SB3_22/i0[10] ), .A3(
        \SB3_22/i1[9] ), .ZN(\SB3_22/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U1864 ( .A1(\SB3_22/i0_4 ), .A2(\SB3_22/i0_3 ), .A3(\SB3_22/i1[9] ), 
        .ZN(\SB3_22/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 U1869 ( .A1(\SB3_22/i0_3 ), .A2(\SB3_22/i1[9] ), .ZN(
        \SB3_22/Component_Function_1/NAND4_in[0] ) );
  BUF_X2 U1873 ( .I(\MC_ARK_ARC_1_2/buf_output[69] ), .Z(\SB1_3_20/i0[10] ) );
  INV_X1 U1880 ( .I(\MC_ARK_ARC_1_2/buf_output[69] ), .ZN(\SB1_3_20/i0[8] ) );
  NAND3_X1 U1886 ( .A1(\SB2_2_11/i3[0] ), .A2(\SB2_2_11/i0_0 ), .A3(
        \SB2_2_11/i1_7 ), .ZN(\SB2_2_11/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U1887 ( .A1(\SB2_2_11/i0_4 ), .A2(\SB2_2_11/i1_7 ), .A3(
        \SB2_2_11/i0[8] ), .ZN(n1431) );
  NAND3_X1 U1890 ( .A1(n5515), .A2(\SB1_2_13/buf_output[3] ), .A3(
        \SB2_2_11/i1_7 ), .ZN(\SB2_2_11/Component_Function_3/NAND4_in[2] ) );
  CLKBUF_X4 U1897 ( .I(\SB3_3/buf_output[5] ), .Z(\SB4_3/i0_3 ) );
  NAND3_X1 U1900 ( .A1(\SB2_3_14/i1_5 ), .A2(\SB2_3_14/i0[10] ), .A3(
        \SB2_3_14/i1[9] ), .ZN(\SB2_3_14/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U1902 ( .A1(\SB1_3_20/i0_0 ), .A2(\SB1_3_20/i0_4 ), .A3(
        \SB1_3_20/i1_5 ), .ZN(\SB1_3_20/Component_Function_2/NAND4_in[3] ) );
  NAND2_X1 U1905 ( .A1(\SB1_3_20/i0_0 ), .A2(\SB1_3_20/i3[0] ), .ZN(
        \SB1_3_20/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U1906 ( .A1(\SB1_3_20/i0_0 ), .A2(\SB1_3_20/i0[6] ), .A3(
        \SB1_3_20/i0[10] ), .ZN(\SB1_3_20/Component_Function_5/NAND4_in[1] )
         );
  NAND3_X1 U1912 ( .A1(\SB4_30/i0[10] ), .A2(\SB4_30/i0[6] ), .A3(
        \SB4_30/i0_0 ), .ZN(n5172) );
  NAND3_X1 U1913 ( .A1(\SB4_30/i0_0 ), .A2(\SB4_30/i0_4 ), .A3(n5525), .ZN(
        n5424) );
  NAND3_X1 U1914 ( .A1(\SB4_30/i0_0 ), .A2(\SB4_30/i3[0] ), .A3(\SB4_30/i1_7 ), 
        .ZN(\SB4_30/Component_Function_4/NAND4_in[1] ) );
  BUF_X2 U1934 ( .I(\SB3_1/buf_output[2] ), .Z(\SB4_30/i0_0 ) );
  INV_X1 U1939 ( .I(\MC_ARK_ARC_1_3/buf_output[162] ), .ZN(\SB3_4/i3[0] ) );
  BUF_X2 U1941 ( .I(\MC_ARK_ARC_1_3/buf_output[162] ), .Z(\SB3_4/i0[9] ) );
  INV_X1 U1942 ( .I(\MC_ARK_ARC_1_3/buf_output[180] ), .ZN(\SB3_1/i3[0] ) );
  BUF_X2 U1947 ( .I(\MC_ARK_ARC_1_3/buf_output[180] ), .Z(\SB3_1/i0[9] ) );
  NAND3_X1 U1948 ( .A1(\SB4_22/i0_0 ), .A2(\SB4_22/i1_5 ), .A3(\SB4_22/i0_4 ), 
        .ZN(\SB4_22/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U1972 ( .A1(\SB3_14/i0_0 ), .A2(\SB3_14/i1_5 ), .A3(\SB3_14/i0_4 ), 
        .ZN(\SB3_14/Component_Function_2/NAND4_in[3] ) );
  BUF_X2 U1976 ( .I(\SB3_18/buf_output[4] ), .Z(\SB4_17/i0_4 ) );
  NAND3_X1 U1977 ( .A1(\SB3_23/i0_0 ), .A2(\SB3_23/i1_5 ), .A3(\SB3_23/i0_4 ), 
        .ZN(n4597) );
  NAND2_X1 U1985 ( .A1(\SB3_23/i0_0 ), .A2(\SB3_23/i3[0] ), .ZN(n5781) );
  NAND3_X1 U1986 ( .A1(\SB3_23/i3[0] ), .A2(\SB3_23/i0_0 ), .A3(\SB3_23/i1_7 ), 
        .ZN(\SB3_23/Component_Function_4/NAND4_in[1] ) );
  BUF_X2 U1987 ( .I(\SB3_13/buf_output[5] ), .Z(\SB4_13/i0_3 ) );
  INV_X1 U1989 ( .I(\SB3_13/buf_output[5] ), .ZN(\SB4_13/i1_5 ) );
  CLKBUF_X4 U1990 ( .I(\SB2_2_12/buf_output[2] ), .Z(\RI5[2][134] ) );
  CLKBUF_X4 U1996 ( .I(\SB3_4/buf_output[5] ), .Z(\SB4_4/i0_3 ) );
  NAND3_X1 U2002 ( .A1(\SB1_3_29/i0[10] ), .A2(\RI1[3][14] ), .A3(
        \SB1_3_29/i0[6] ), .ZN(\SB1_3_29/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U2004 ( .A1(\SB1_3_29/i0_3 ), .A2(\SB1_3_29/i0[10] ), .A3(
        \SB1_3_29/i0[9] ), .ZN(n2555) );
  NAND3_X1 U2005 ( .A1(\SB1_3_29/i0[10] ), .A2(\SB1_3_29/i0_3 ), .A3(
        \SB1_3_29/i0[6] ), .ZN(n5906) );
  INV_X1 U2008 ( .I(\MC_ARK_ARC_1_2/buf_output[15] ), .ZN(\SB1_3_29/i0[8] ) );
  BUF_X2 U2010 ( .I(\MC_ARK_ARC_1_2/buf_output[15] ), .Z(\SB1_3_29/i0[10] ) );
  BUF_X2 U2011 ( .I(\SB3_17/buf_output[0] ), .Z(\SB4_12/i0[9] ) );
  NAND2_X1 U2012 ( .A1(\SB1_2_20/i0_0 ), .A2(\SB1_2_20/i3[0] ), .ZN(
        \SB1_2_20/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U2018 ( .A1(\SB1_2_20/i0[7] ), .A2(\SB1_2_20/i0_3 ), .A3(
        \SB1_2_20/i0_0 ), .ZN(\SB1_2_20/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2020 ( .A1(\SB1_2_20/i0_0 ), .A2(\SB1_2_20/i0_4 ), .A3(n2909), 
        .ZN(n6465) );
  BUF_X2 U2024 ( .I(\MC_ARK_ARC_1_0/buf_output[81] ), .Z(\SB1_1_18/i0[10] ) );
  INV_X1 U2026 ( .I(\MC_ARK_ARC_1_0/buf_output[81] ), .ZN(\SB1_1_18/i0[8] ) );
  INV_X1 U2027 ( .I(\SB3_2/buf_output[1] ), .ZN(\SB4_30/i1_7 ) );
  BUF_X2 U2030 ( .I(\SB3_2/buf_output[1] ), .Z(\SB4_30/i0[6] ) );
  NAND3_X1 U2034 ( .A1(\SB4_13/i0_0 ), .A2(\SB4_13/i3[0] ), .A3(\SB4_13/i1_7 ), 
        .ZN(\SB4_13/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U2038 ( .A1(\SB3_20/i0_4 ), .A2(\SB3_20/i0_3 ), .A3(\SB3_20/i1[9] ), 
        .ZN(n4226) );
  NAND3_X1 U2045 ( .A1(\SB1_0_10/i0[10] ), .A2(\SB1_0_10/i0_3 ), .A3(
        \SB1_0_10/i0[6] ), .ZN(n2431) );
  NAND3_X1 U2046 ( .A1(\SB1_0_10/i0_0 ), .A2(\SB1_0_10/i0_3 ), .A3(
        \SB1_0_10/i0_4 ), .ZN(\SB1_0_10/Component_Function_3/NAND4_in[1] ) );
  CLKBUF_X4 U2048 ( .I(n426), .Z(\SB1_0_10/i0_3 ) );
  NAND3_X1 U2051 ( .A1(\SB4_14/i1[9] ), .A2(\SB4_14/i1_5 ), .A3(\SB4_14/i0_4 ), 
        .ZN(\SB4_14/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U2055 ( .A1(\SB4_14/i1_7 ), .A2(\SB4_14/i0[8] ), .A3(\SB4_14/i0_4 ), 
        .ZN(\SB4_14/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U2056 ( .A1(\SB4_14/i0_4 ), .A2(\SB4_14/i0_0 ), .A3(\SB4_14/i1_5 ), 
        .ZN(n6491) );
  NAND3_X1 U2062 ( .A1(\SB4_14/i0_0 ), .A2(\SB4_14/i0_3 ), .A3(\SB4_14/i0_4 ), 
        .ZN(n4053) );
  CLKBUF_X2 U2063 ( .I(\RI1[3][167] ), .Z(n5189) );
  INV_X1 U2068 ( .I(\MC_ARK_ARC_1_3/buf_output[86] ), .ZN(\SB3_17/i1[9] ) );
  BUF_X2 U2070 ( .I(\MC_ARK_ARC_1_3/buf_output[86] ), .Z(\SB3_17/i0_0 ) );
  CLKBUF_X4 U2072 ( .I(\SB3_0/buf_output[3] ), .Z(\SB4_30/i0[10] ) );
  NAND3_X1 U2075 ( .A1(\SB3_23/i0_3 ), .A2(\SB3_23/i1[9] ), .A3(\SB3_23/i0_4 ), 
        .ZN(\SB3_23/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2078 ( .A1(\SB3_23/i0_3 ), .A2(\SB3_23/i0[8] ), .A3(\SB3_23/i0[9] ), .ZN(n942) );
  NAND2_X1 U2079 ( .A1(\SB3_23/i0_3 ), .A2(\SB3_23/i1[9] ), .ZN(n6112) );
  NAND3_X1 U2081 ( .A1(\SB3_23/i0_0 ), .A2(\SB3_23/i0_3 ), .A3(\SB3_23/i0_4 ), 
        .ZN(\SB3_23/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2086 ( .A1(\SB3_23/i0_3 ), .A2(\SB3_23/i0_4 ), .A3(\SB3_23/i0[10] ), .ZN(\SB3_23/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U2089 ( .A1(\SB3_23/i0_3 ), .A2(\SB3_23/i1[9] ), .A3(\SB3_23/i0[6] ), .ZN(n5255) );
  CLKBUF_X4 U2094 ( .I(\SB2_2_9/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[162] ) );
  NAND3_X1 U2096 ( .A1(\SB3_24/i0_3 ), .A2(\SB3_24/i1[9] ), .A3(\SB3_24/i0[6] ), .ZN(n6529) );
  NAND3_X1 U2097 ( .A1(\SB3_24/i0_3 ), .A2(\SB3_24/i0[9] ), .A3(\SB3_24/i0[8] ), .ZN(n3888) );
  NAND3_X1 U2098 ( .A1(\SB2_1_5/i0_3 ), .A2(\SB1_1_6/buf_output[4] ), .A3(
        \SB2_1_5/i1[9] ), .ZN(\SB2_1_5/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2101 ( .A1(\SB2_1_5/i0_3 ), .A2(\SB2_1_5/i0[6] ), .A3(
        \SB2_1_5/i1[9] ), .ZN(n6301) );
  NAND3_X1 U2109 ( .A1(\SB2_1_5/i0[10] ), .A2(\SB2_1_5/i1_5 ), .A3(
        \SB2_1_5/i1[9] ), .ZN(\SB2_1_5/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U2116 ( .A1(\SB2_1_5/i0[10] ), .A2(\SB2_1_5/i1[9] ), .A3(
        \SB2_1_5/i1_7 ), .ZN(n1558) );
  NAND2_X1 U2117 ( .A1(\SB2_1_5/i0_3 ), .A2(\SB2_1_5/i1[9] ), .ZN(n3724) );
  NAND2_X1 U2119 ( .A1(\SB1_0_24/i0_0 ), .A2(\SB1_0_24/i3[0] ), .ZN(
        \SB1_0_24/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U2135 ( .A1(\SB1_0_24/i0_4 ), .A2(\SB1_0_24/i0_0 ), .A3(
        \SB1_0_24/i1_5 ), .ZN(n1167) );
  NAND3_X1 U2138 ( .A1(\SB1_0_24/i0_0 ), .A2(\SB1_0_24/i0[10] ), .A3(
        \SB1_0_24/i0[6] ), .ZN(\SB1_0_24/Component_Function_5/NAND4_in[1] ) );
  BUF_X2 U2143 ( .I(n374), .Z(\SB1_0_15/i0_4 ) );
  BUF_X4 U2150 ( .I(\MC_ARK_ARC_1_3/buf_output[119] ), .Z(\SB3_12/i0_3 ) );
  CLKBUF_X4 U2153 ( .I(\MC_ARK_ARC_1_3/buf_output[116] ), .Z(\SB3_12/i0_0 ) );
  CLKBUF_X4 U2154 ( .I(\MC_ARK_ARC_1_3/buf_output[63] ), .Z(\SB3_21/i0[10] )
         );
  NAND3_X1 U2157 ( .A1(\SB1_3_28/i0[9] ), .A2(\SB1_3_28/i0_3 ), .A3(
        \SB1_3_28/i0[8] ), .ZN(n5441) );
  NAND3_X1 U2160 ( .A1(\SB1_3_28/i1[9] ), .A2(\SB1_3_28/i0_3 ), .A3(
        \SB1_3_28/i0[6] ), .ZN(\SB1_3_28/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2163 ( .A1(\SB1_3_28/i0[10] ), .A2(\SB1_3_28/i0_3 ), .A3(
        \SB1_3_28/i0[6] ), .ZN(\SB1_3_28/Component_Function_2/NAND4_in[1] ) );
  INV_X1 U2167 ( .I(\MC_ARK_ARC_1_3/buf_output[150] ), .ZN(\SB3_6/i3[0] ) );
  BUF_X2 U2168 ( .I(\MC_ARK_ARC_1_3/buf_output[150] ), .Z(\SB3_6/i0[9] ) );
  CLKBUF_X4 U2170 ( .I(\SB3_10/buf_output[5] ), .Z(\SB4_10/i0_3 ) );
  NAND3_X1 U2173 ( .A1(\SB3_2/i0[9] ), .A2(\SB3_2/i0_3 ), .A3(\SB3_2/i0[8] ), 
        .ZN(n6215) );
  NAND3_X1 U2175 ( .A1(\SB3_2/i0_3 ), .A2(\SB3_2/i1_7 ), .A3(\SB3_2/i0[8] ), 
        .ZN(\SB3_2/Component_Function_1/NAND4_in[1] ) );
  CLKBUF_X4 U2176 ( .I(\SB2_1_10/buf_output[3] ), .Z(\RI5[1][141] ) );
  NAND3_X1 U2180 ( .A1(\SB1_3_12/i1[9] ), .A2(\SB1_3_12/i0_4 ), .A3(
        \SB1_3_12/i0_3 ), .ZN(\SB1_3_12/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2181 ( .A1(\SB1_3_12/i0_0 ), .A2(\SB1_3_12/i0_4 ), .A3(
        \SB1_3_12/i0_3 ), .ZN(n3360) );
  NAND3_X1 U2182 ( .A1(\SB1_3_12/i0_0 ), .A2(\SB1_3_12/i0_3 ), .A3(
        \SB1_3_12/i0[7] ), .ZN(\SB1_3_12/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2185 ( .A1(\SB1_3_12/i0_3 ), .A2(\SB1_3_12/i0[6] ), .A3(
        \SB1_3_12/i1[9] ), .ZN(n6462) );
  NAND3_X1 U2186 ( .A1(\SB1_3_12/i0_3 ), .A2(\SB1_3_12/i0[8] ), .A3(
        \SB1_3_12/i0[9] ), .ZN(\SB1_3_12/Component_Function_2/NAND4_in[2] ) );
  NAND2_X1 U2187 ( .A1(\SB1_3_12/i0_3 ), .A2(\SB1_3_12/i1[9] ), .ZN(n5942) );
  NAND3_X1 U2188 ( .A1(\SB1_3_12/i0[10] ), .A2(\SB1_3_12/i0_4 ), .A3(
        \SB1_3_12/i0_3 ), .ZN(\SB1_3_12/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U2191 ( .A1(\SB1_3_12/i0_3 ), .A2(\SB1_3_12/i0[9] ), .A3(
        \SB1_3_12/i0[10] ), .ZN(n6125) );
  CLKBUF_X4 U2192 ( .I(\SB2_1_22/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[74] ) );
  CLKBUF_X4 U2198 ( .I(\SB3_16/buf_output[2] ), .Z(\SB4_13/i0_0 ) );
  INV_X1 U2200 ( .I(\SB3_3/buf_output[1] ), .ZN(\SB4_31/i1_7 ) );
  BUF_X2 U2202 ( .I(\SB3_3/buf_output[1] ), .Z(\SB4_31/i0[6] ) );
  NAND3_X1 U2215 ( .A1(\SB3_24/i1_5 ), .A2(\SB3_24/i0_0 ), .A3(\SB3_24/i0_4 ), 
        .ZN(\SB3_24/Component_Function_2/NAND4_in[3] ) );
  NAND2_X1 U2217 ( .A1(\SB3_24/i0_0 ), .A2(\SB3_24/i3[0] ), .ZN(n1250) );
  NAND3_X1 U2222 ( .A1(\SB3_24/i0_0 ), .A2(\SB3_24/i0[8] ), .A3(\SB3_24/i0[9] ), .ZN(n5396) );
  NAND3_X1 U2223 ( .A1(\SB3_24/i0_0 ), .A2(\SB3_24/i0[10] ), .A3(
        \SB3_24/i0[6] ), .ZN(n4997) );
  INV_X1 U2224 ( .I(\SB3_26/buf_output[2] ), .ZN(\SB4_23/i1[9] ) );
  BUF_X2 U2225 ( .I(\SB3_26/buf_output[2] ), .Z(\SB4_23/i0_0 ) );
  BUF_X2 U2229 ( .I(\SB3_5/buf_output[1] ), .Z(\SB4_1/i0[6] ) );
  INV_X1 U2232 ( .I(\MC_ARK_ARC_1_3/buf_output[39] ), .ZN(\SB3_25/i0[8] ) );
  BUF_X2 U2234 ( .I(\MC_ARK_ARC_1_3/buf_output[39] ), .Z(\SB3_25/i0[10] ) );
  INV_X1 U2240 ( .I(\MC_ARK_ARC_1_3/buf_output[80] ), .ZN(\SB3_18/i1[9] ) );
  BUF_X2 U2246 ( .I(\MC_ARK_ARC_1_3/buf_output[80] ), .Z(\SB3_18/i0_0 ) );
  INV_X1 U2250 ( .I(\MC_ARK_ARC_1_3/buf_output[177] ), .ZN(\SB3_2/i0[8] ) );
  BUF_X2 U2256 ( .I(\MC_ARK_ARC_1_3/buf_output[177] ), .Z(\SB3_2/i0[10] ) );
  INV_X1 U2260 ( .I(\MC_ARK_ARC_1_3/buf_output[153] ), .ZN(\SB3_6/i0[8] ) );
  BUF_X2 U2261 ( .I(\MC_ARK_ARC_1_3/buf_output[153] ), .Z(\SB3_6/i0[10] ) );
  INV_X1 U2262 ( .I(\MC_ARK_ARC_1_2/buf_output[27] ), .ZN(\SB1_3_27/i0[8] ) );
  BUF_X2 U2263 ( .I(\MC_ARK_ARC_1_2/buf_output[27] ), .Z(\SB1_3_27/i0[10] ) );
  BUF_X2 U2264 ( .I(\SB3_17/buf_output[2] ), .Z(\SB4_14/i0_0 ) );
  INV_X1 U2265 ( .I(\SB3_17/buf_output[2] ), .ZN(\SB4_14/i1[9] ) );
  NAND2_X1 U2266 ( .A1(\SB4_30/i0_3 ), .A2(n4751), .ZN(
        \SB4_30/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U2268 ( .A1(\SB4_30/i0_3 ), .A2(\SB4_30/i0_0 ), .A3(\SB4_30/i0_4 ), 
        .ZN(n3935) );
  NAND3_X1 U2278 ( .A1(\SB4_30/i0_3 ), .A2(\SB4_30/i1_7 ), .A3(\SB4_30/i0[8] ), 
        .ZN(\SB4_30/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U2280 ( .A1(\SB4_30/i0_0 ), .A2(\SB4_30/i0[7] ), .A3(\SB4_30/i0_3 ), 
        .ZN(n5433) );
  NAND3_X1 U2281 ( .A1(\SB4_30/i0[10] ), .A2(\SB4_30/i0_4 ), .A3(\SB4_30/i0_3 ), .ZN(\SB4_30/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U2282 ( .A1(\SB4_30/i0[6] ), .A2(\SB4_30/i0_3 ), .A3(n4751), .ZN(
        n5339) );
  NAND3_X1 U2286 ( .A1(\SB4_30/i0[6] ), .A2(\SB4_30/i0[10] ), .A3(
        \SB4_30/i0_3 ), .ZN(n5312) );
  NAND3_X1 U2290 ( .A1(\SB4_30/i0[10] ), .A2(\SB4_30/i0[9] ), .A3(
        \SB4_30/i0_3 ), .ZN(n4851) );
  CLKBUF_X2 U2294 ( .I(\SB3_12/buf_output[3] ), .Z(\SB4_10/i0[10] ) );
  INV_X1 U2295 ( .I(\SB3_12/buf_output[3] ), .ZN(\SB4_10/i0[8] ) );
  NAND3_X1 U2298 ( .A1(\SB4_6/i0_0 ), .A2(\SB4_6/i0_3 ), .A3(\SB4_6/i0_4 ), 
        .ZN(\SB4_6/Component_Function_3/NAND4_in[1] ) );
  BUF_X2 U2299 ( .I(\MC_ARK_ARC_1_1/buf_output[146] ), .Z(\SB1_2_7/i0_0 ) );
  INV_X1 U2300 ( .I(\MC_ARK_ARC_1_1/buf_output[146] ), .ZN(\SB1_2_7/i1[9] ) );
  INV_X1 U2303 ( .I(\MC_ARK_ARC_1_0/buf_output[54] ), .ZN(\SB1_1_22/i3[0] ) );
  BUF_X2 U2304 ( .I(\MC_ARK_ARC_1_0/buf_output[54] ), .Z(\SB1_1_22/i0[9] ) );
  AND2_X1 U2305 ( .A1(\MC_ARK_ARC_1_0/buf_output[54] ), .A2(
        \MC_ARK_ARC_1_0/buf_output[55] ), .Z(n4522) );
  NAND3_X1 U2306 ( .A1(\SB2_3_18/i0_3 ), .A2(\SB2_3_18/i1[9] ), .A3(
        \SB2_3_18/i0_4 ), .ZN(n2576) );
  NAND3_X1 U2308 ( .A1(\SB2_3_18/i1[9] ), .A2(\SB2_3_18/i1_7 ), .A3(
        \SB2_3_18/i0[10] ), .ZN(\SB2_3_18/Component_Function_3/NAND4_in[2] )
         );
  NAND3_X1 U2309 ( .A1(\SB2_3_18/i0[10] ), .A2(\SB2_3_18/i1_5 ), .A3(
        \SB2_3_18/i1[9] ), .ZN(\SB2_3_18/Component_Function_2/NAND4_in[0] ) );
  CLKBUF_X4 U2310 ( .I(\SB3_7/buf_output[5] ), .Z(\SB4_7/i0_3 ) );
  NAND3_X1 U2311 ( .A1(\SB2_1_0/i0_3 ), .A2(\SB2_1_0/i0[10] ), .A3(n2687), 
        .ZN(n4535) );
  NAND3_X1 U2312 ( .A1(\SB2_1_0/i0[10] ), .A2(\SB2_1_0/i0_3 ), .A3(
        \SB2_1_0/i0[9] ), .ZN(n4422) );
  NAND3_X1 U2313 ( .A1(\SB2_1_0/i0[7] ), .A2(\SB2_1_0/i0_0 ), .A3(
        \SB2_1_0/i0_3 ), .ZN(n1708) );
  NAND3_X1 U2315 ( .A1(\SB2_1_0/i0_0 ), .A2(\SB2_1_0/i0_3 ), .A3(n2687), .ZN(
        \SB2_1_0/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2316 ( .A1(\SB2_1_0/i0[10] ), .A2(\SB2_1_0/i0_3 ), .A3(
        \SB2_1_0/i0[6] ), .ZN(n5108) );
  NAND3_X1 U2319 ( .A1(\SB4_18/i0_0 ), .A2(n3662), .A3(\SB4_18/i0[9] ), .ZN(
        n1220) );
  NAND3_X1 U2322 ( .A1(\SB2_3_12/i0_3 ), .A2(n1603), .A3(n3651), .ZN(
        \SB2_3_12/Component_Function_2/NAND4_in[2] ) );
  NAND2_X1 U2323 ( .A1(\SB2_0_13/i0_3 ), .A2(\SB2_0_13/i1[9] ), .ZN(
        \SB2_0_13/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U2324 ( .A1(\SB2_0_13/i1[9] ), .A2(\SB2_0_13/i0_3 ), .A3(
        \SB2_0_13/i0[6] ), .ZN(\SB2_0_13/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2326 ( .A1(\SB2_0_13/i1[9] ), .A2(n3663), .A3(\SB2_0_13/i0_4 ), 
        .ZN(\SB2_0_13/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U2329 ( .A1(\SB2_0_13/i0[10] ), .A2(n3663), .A3(\SB2_0_13/i1[9] ), 
        .ZN(\SB2_0_13/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U2330 ( .A1(\SB2_0_13/i1_7 ), .A2(\SB2_0_13/i0[10] ), .A3(
        \SB2_0_13/i1[9] ), .ZN(\SB2_0_13/Component_Function_3/NAND4_in[2] ) );
  INV_X1 U2333 ( .I(\MC_ARK_ARC_1_1/buf_output[144] ), .ZN(\SB1_2_7/i3[0] ) );
  BUF_X2 U2335 ( .I(\MC_ARK_ARC_1_1/buf_output[144] ), .Z(\SB1_2_7/i0[9] ) );
  INV_X1 U2337 ( .I(\MC_ARK_ARC_1_3/buf_output[93] ), .ZN(\SB3_16/i0[8] ) );
  BUF_X2 U2338 ( .I(\MC_ARK_ARC_1_3/buf_output[93] ), .Z(\SB3_16/i0[10] ) );
  CLKBUF_X4 U2339 ( .I(\SB2_3_28/buf_output[3] ), .Z(\RI5[3][33] ) );
  NAND3_X1 U2341 ( .A1(\SB1_2_1/i0[8] ), .A2(\SB1_2_1/i1_5 ), .A3(
        \SB1_2_1/i3[0] ), .ZN(\SB1_2_1/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2343 ( .A1(\SB1_2_1/i0[6] ), .A2(\SB1_2_1/i0[8] ), .A3(
        \SB1_2_1/i0[7] ), .ZN(\SB1_2_1/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U2345 ( .A1(\SB4_1/i0[6] ), .A2(\SB4_1/i0_0 ), .A3(\SB4_1/i0[10] ), 
        .ZN(n5196) );
  NAND3_X1 U2349 ( .A1(\SB4_1/i0_3 ), .A2(\SB4_1/i0[6] ), .A3(\SB4_1/i1[9] ), 
        .ZN(n2960) );
  BUF_X2 U2350 ( .I(\SB1_3_31/buf_output[0] ), .Z(\SB2_3_26/i0[9] ) );
  INV_X1 U2352 ( .I(\SB1_3_31/buf_output[0] ), .ZN(\SB2_3_26/i3[0] ) );
  INV_X1 U2357 ( .I(\MC_ARK_ARC_1_2/buf_output[43] ), .ZN(\SB1_3_24/i1_7 ) );
  BUF_X2 U2359 ( .I(\MC_ARK_ARC_1_2/buf_output[43] ), .Z(\SB1_3_24/i0[6] ) );
  BUF_X2 U2362 ( .I(\MC_ARK_ARC_1_0/buf_output[163] ), .Z(\SB1_1_4/i0[6] ) );
  INV_X1 U2364 ( .I(\MC_ARK_ARC_1_0/buf_output[163] ), .ZN(\SB1_1_4/i1_7 ) );
  NAND2_X1 U2366 ( .A1(\SB4_0/i0[10] ), .A2(\SB4_0/i0[9] ), .ZN(
        \SB4_0/Component_Function_0/NAND4_in[0] ) );
  BUF_X2 U2369 ( .I(\SB3_5/buf_output[0] ), .Z(\SB4_0/i0[9] ) );
  INV_X1 U2370 ( .I(\SB3_22/buf_output[3] ), .ZN(\SB4_20/i0[8] ) );
  BUF_X2 U2371 ( .I(\SB3_22/buf_output[3] ), .Z(\SB4_20/i0[10] ) );
  INV_X1 U2373 ( .I(\MC_ARK_ARC_1_3/buf_output[140] ), .ZN(\SB3_8/i1[9] ) );
  BUF_X2 U2379 ( .I(\MC_ARK_ARC_1_3/buf_output[140] ), .Z(\SB3_8/i0_0 ) );
  INV_X1 U2380 ( .I(\MC_ARK_ARC_1_3/buf_output[183] ), .ZN(\SB3_1/i0[8] ) );
  BUF_X2 U2381 ( .I(\MC_ARK_ARC_1_3/buf_output[183] ), .Z(\SB3_1/i0[10] ) );
  INV_X1 U2382 ( .I(\MC_ARK_ARC_1_0/buf_output[99] ), .ZN(\SB1_1_15/i0[8] ) );
  BUF_X2 U2383 ( .I(\MC_ARK_ARC_1_0/buf_output[99] ), .Z(\SB1_1_15/i0[10] ) );
  CLKBUF_X4 U2384 ( .I(\SB2_3_27/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[44] ) );
  NAND3_X1 U2389 ( .A1(\SB2_0_16/i0_3 ), .A2(\SB2_0_16/i0_0 ), .A3(
        \SB2_0_16/i0_4 ), .ZN(\SB2_0_16/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2393 ( .A1(\SB2_0_16/i0[9] ), .A2(\SB2_0_16/i0_3 ), .A3(
        \SB2_0_16/i0[10] ), .ZN(n4157) );
  NAND3_X1 U2400 ( .A1(\SB2_0_16/i1[9] ), .A2(\SB2_0_16/i0_3 ), .A3(
        \SB2_0_16/i0[6] ), .ZN(\SB2_0_16/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2401 ( .A1(\SB2_0_16/i0_3 ), .A2(\SB2_0_16/i0[9] ), .A3(
        \SB2_0_16/i0[8] ), .ZN(n4621) );
  NAND3_X1 U2403 ( .A1(\SB2_0_16/i0_3 ), .A2(\SB2_0_16/i0[10] ), .A3(
        \SB2_0_16/i0_4 ), .ZN(n4510) );
  NAND3_X1 U2406 ( .A1(\SB2_0_16/i0_3 ), .A2(\SB2_0_16/i0[10] ), .A3(
        \SB2_0_16/i0[6] ), .ZN(\SB2_0_16/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U2408 ( .A1(\SB3_21/i0[10] ), .A2(\SB3_21/i1[9] ), .A3(
        \SB3_21/i1_7 ), .ZN(n2005) );
  NAND3_X1 U2409 ( .A1(\SB3_21/i0_3 ), .A2(\SB3_21/i0[10] ), .A3(
        \SB3_21/i0[9] ), .ZN(n6459) );
  NAND3_X1 U2410 ( .A1(\SB3_21/i1_5 ), .A2(\SB3_21/i0[10] ), .A3(
        \SB3_21/i1[9] ), .ZN(\SB3_21/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U2411 ( .A1(\SB3_21/i0[10] ), .A2(\SB3_21/i0[6] ), .A3(\RI1[4][65] ), .ZN(n4002) );
  NAND3_X1 U2415 ( .A1(\SB1_2_29/i0[10] ), .A2(\RI1[2][17] ), .A3(
        \SB1_2_29/i0[9] ), .ZN(\SB1_2_29/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U2419 ( .A1(\SB1_2_29/i0[10] ), .A2(\RI1[2][17] ), .A3(
        \SB1_2_29/i0[6] ), .ZN(\SB1_2_29/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U2420 ( .A1(\SB1_2_29/i0[10] ), .A2(\SB1_2_29/i0_0 ), .A3(
        \SB1_2_29/i0[6] ), .ZN(\SB1_2_29/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U2421 ( .A1(\SB1_2_29/i1_5 ), .A2(\SB1_2_29/i0[10] ), .A3(
        \SB1_2_29/i1[9] ), .ZN(\SB1_2_29/Component_Function_2/NAND4_in[0] ) );
  INV_X1 U2422 ( .I(\MC_ARK_ARC_1_2/buf_output[19] ), .ZN(\SB1_3_28/i1_7 ) );
  BUF_X2 U2423 ( .I(\MC_ARK_ARC_1_2/buf_output[19] ), .Z(\SB1_3_28/i0[6] ) );
  BUF_X2 U2424 ( .I(\MC_ARK_ARC_1_3/buf_output[85] ), .Z(\SB3_17/i0[6] ) );
  INV_X1 U2425 ( .I(\MC_ARK_ARC_1_3/buf_output[85] ), .ZN(\SB3_17/i1_7 ) );
  INV_X1 U2426 ( .I(n307), .ZN(\SB1_0_11/i1[9] ) );
  BUF_X2 U2430 ( .I(n307), .Z(\SB1_0_11/i0_0 ) );
  NAND3_X1 U2431 ( .A1(\SB1_0_23/i1_5 ), .A2(\SB1_0_23/i0[8] ), .A3(
        \SB1_0_23/i3[0] ), .ZN(\SB1_0_23/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2436 ( .A1(\SB1_0_23/i1_5 ), .A2(\SB1_0_23/i0_0 ), .A3(
        \SB1_0_23/i0_4 ), .ZN(\SB1_0_23/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U2439 ( .A1(\SB1_0_23/i1[9] ), .A2(\SB1_0_23/i1_5 ), .A3(
        \SB1_0_23/i0_4 ), .ZN(\SB1_0_23/Component_Function_4/NAND4_in[3] ) );
  INV_X1 U2440 ( .I(\SB1_2_23/buf_output[1] ), .ZN(\SB2_2_19/i1_7 ) );
  BUF_X2 U2441 ( .I(\SB1_2_23/buf_output[1] ), .Z(\SB2_2_19/i0[6] ) );
  INV_X1 U2442 ( .I(\MC_ARK_ARC_1_2/buf_output[68] ), .ZN(\SB1_3_20/i1[9] ) );
  BUF_X2 U2444 ( .I(\MC_ARK_ARC_1_2/buf_output[68] ), .Z(\SB1_3_20/i0_0 ) );
  CLKBUF_X4 U2445 ( .I(\SB1_2_10/buf_output[5] ), .Z(\SB2_2_10/i0_3 ) );
  CLKBUF_X4 U2447 ( .I(\SB1_1_0/buf_output[5] ), .Z(\SB2_1_0/i0_3 ) );
  BUF_X2 U2449 ( .I(\MC_ARK_ARC_1_2/buf_output[55] ), .Z(\SB1_3_22/i0[6] ) );
  NAND2_X1 U2450 ( .A1(\SB1_0_18/i0_3 ), .A2(\SB1_0_18/i1[9] ), .ZN(n6499) );
  NAND3_X1 U2454 ( .A1(\SB1_0_18/i1[9] ), .A2(\SB1_0_18/i1_5 ), .A3(n4753), 
        .ZN(\SB1_0_18/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U2455 ( .A1(\SB1_0_18/i1[9] ), .A2(\SB1_0_18/i1_7 ), .A3(n1367), 
        .ZN(\SB1_0_18/Component_Function_3/NAND4_in[2] ) );
  INV_X1 U2456 ( .I(\MC_ARK_ARC_1_3/buf_output[189] ), .ZN(\SB3_0/i0[8] ) );
  BUF_X2 U2459 ( .I(\MC_ARK_ARC_1_3/buf_output[189] ), .Z(\SB3_0/i0[10] ) );
  INV_X1 U2460 ( .I(\MC_ARK_ARC_1_1/buf_output[133] ), .ZN(\SB1_2_9/i1_7 ) );
  BUF_X2 U2466 ( .I(\MC_ARK_ARC_1_1/buf_output[133] ), .Z(\SB1_2_9/i0[6] ) );
  INV_X1 U2474 ( .I(\MC_ARK_ARC_1_1/buf_output[97] ), .ZN(\SB1_2_15/i1_7 ) );
  BUF_X2 U2477 ( .I(\MC_ARK_ARC_1_1/buf_output[97] ), .Z(\SB1_2_15/i0[6] ) );
  INV_X1 U2479 ( .I(\MC_ARK_ARC_1_3/buf_output[165] ), .ZN(\SB3_4/i0[8] ) );
  BUF_X2 U2480 ( .I(\MC_ARK_ARC_1_3/buf_output[165] ), .Z(\SB3_4/i0[10] ) );
  INV_X2 U2482 ( .I(\SB2_1_15/i0_4 ), .ZN(n5493) );
  CLKBUF_X4 U2484 ( .I(n3686), .Z(\SB1_2_9/i0_0 ) );
  AND4_X2 U2494 ( .A1(\SB3_1/Component_Function_2/NAND4_in[1] ), .A2(
        \SB3_1/Component_Function_2/NAND4_in[2] ), .A3(
        \SB3_1/Component_Function_2/NAND4_in[0] ), .A4(n4092), .Z(n4751) );
  BUF_X4 U2495 ( .I(\SB1_3_3/buf_output[4] ), .Z(\SB2_3_2/i0_4 ) );
  BUF_X2 U2496 ( .I(\MC_ARK_ARC_1_3/buf_output[104] ), .Z(\SB3_14/i0_0 ) );
  INV_X1 U2504 ( .I(\MC_ARK_ARC_1_3/buf_output[104] ), .ZN(\SB3_14/i1[9] ) );
  INV_X1 U2512 ( .I(\RI1[3][41] ), .ZN(\SB1_3_25/i1_5 ) );
  NAND3_X1 U2513 ( .A1(\SB2_3_9/i0[9] ), .A2(\SB2_3_9/i0[10] ), .A3(
        \SB2_3_9/i0_3 ), .ZN(\SB2_3_9/Component_Function_4/NAND4_in[2] ) );
  BUF_X4 U2516 ( .I(\SB1_2_13/buf_output[2] ), .Z(\SB2_2_10/i0_0 ) );
  INV_X1 U2517 ( .I(\SB1_3_0/buf_output[0] ), .ZN(\SB2_3_27/i3[0] ) );
  AND2_X2 U2519 ( .A1(\SB1_3_0/buf_output[0] ), .A2(\SB1_3_28/buf_output[4] ), 
        .Z(n4272) );
  INV_X1 U2520 ( .I(\MC_ARK_ARC_1_2/buf_output[157] ), .ZN(\SB1_3_5/i1_7 ) );
  NAND3_X1 U2521 ( .A1(\SB2_2_11/i0_3 ), .A2(n5826), .A3(\SB2_2_11/i0_4 ), 
        .ZN(n3490) );
  NAND3_X1 U2522 ( .A1(n5826), .A2(\SB2_2_11/i0_3 ), .A3(\SB2_2_11/i0[9] ), 
        .ZN(n1561) );
  NAND3_X1 U2525 ( .A1(\SB2_2_25/i0_3 ), .A2(\SB2_2_25/i1_7 ), .A3(
        \SB2_2_25/i0[8] ), .ZN(\SB2_2_25/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U2529 ( .A1(\SB2_2_25/i0_3 ), .A2(\SB2_2_25/i0_0 ), .A3(
        \SB2_2_25/i0[7] ), .ZN(\SB2_2_25/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2531 ( .A1(\SB2_2_25/i1[9] ), .A2(\SB2_2_25/i0_3 ), .A3(
        \SB2_2_25/i0[6] ), .ZN(\SB2_2_25/Component_Function_3/NAND4_in[0] ) );
  NAND2_X1 U2533 ( .A1(\SB2_2_25/i0_3 ), .A2(\SB2_2_25/i1[9] ), .ZN(
        \SB2_2_25/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U2534 ( .A1(\SB2_2_25/i0_3 ), .A2(\SB2_2_25/i0[9] ), .A3(
        \SB2_2_25/i0[10] ), .ZN(\SB2_2_25/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U2536 ( .A1(\SB2_2_25/i0_3 ), .A2(\SB2_2_25/i0_4 ), .A3(
        \SB2_2_25/i0_0 ), .ZN(\SB2_2_25/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2538 ( .A1(\SB2_2_25/i0_3 ), .A2(\SB2_2_25/i0[8] ), .A3(
        \SB2_2_25/i0[9] ), .ZN(\SB2_2_25/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2539 ( .A1(\SB2_2_25/i0_3 ), .A2(\SB2_2_25/i0[10] ), .A3(
        \SB2_2_25/i0[6] ), .ZN(\SB2_2_25/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U2540 ( .A1(\SB2_2_25/i0_3 ), .A2(\SB2_2_25/i0_4 ), .A3(
        \SB2_2_25/i1[9] ), .ZN(\SB2_2_25/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2544 ( .A1(\SB2_2_25/i0[10] ), .A2(\SB2_2_25/i1[9] ), .A3(
        \SB2_2_25/i1_7 ), .ZN(\SB2_2_25/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2547 ( .A1(\SB1_2_8/i0[8] ), .A2(\SB1_2_8/i3[0] ), .A3(
        \SB1_2_8/i1_5 ), .ZN(\SB1_2_8/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U2554 ( .A1(\SB1_2_8/i0[9] ), .A2(\SB1_2_8/i0[6] ), .A3(
        \SB1_2_8/i1_5 ), .ZN(n4674) );
  NAND3_X1 U2557 ( .A1(\RI3[0][156] ), .A2(\SB2_0_5/i0[6] ), .A3(\RI3[0][160] ), .ZN(\SB2_0_5/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U2560 ( .A1(\SB2_0_5/i0_3 ), .A2(\SB2_0_5/i0[10] ), .A3(
        \RI3[0][156] ), .ZN(\SB2_0_5/Component_Function_4/NAND4_in[2] ) );
  INV_X1 U2561 ( .I(\MC_ARK_ARC_1_0/buf_output[7] ), .ZN(\SB1_1_30/i1_7 ) );
  BUF_X4 U2564 ( .I(\MC_ARK_ARC_1_0/buf_output[7] ), .Z(\SB1_1_30/i0[6] ) );
  OR3_X2 U2565 ( .A1(\SB1_2_7/buf_output[2] ), .A2(n5190), .A3(\SB2_2_4/i0[7] ), .Z(\SB2_2_4/Component_Function_5/NAND4_in[2] ) );
  INV_X1 U2570 ( .I(n337), .ZN(\SB1_0_1/i1[9] ) );
  BUF_X2 U2571 ( .I(n337), .Z(\SB1_0_1/i0_0 ) );
  BUF_X4 U2574 ( .I(\SB2_2_11/buf_output[2] ), .Z(\RI5[2][140] ) );
  CLKBUF_X4 U2575 ( .I(\SB1_1_11/buf_output[2] ), .Z(\SB2_1_8/i0_0 ) );
  NAND3_X1 U2582 ( .A1(n4765), .A2(\SB3_1/i0_3 ), .A3(\SB3_1/i0[6] ), .ZN(
        \SB3_1/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2585 ( .A1(\SB3_4/i1[9] ), .A2(\SB3_4/i0_3 ), .A3(\SB3_4/i0[6] ), 
        .ZN(\SB3_4/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2592 ( .A1(\SB3_4/i0_3 ), .A2(\SB3_4/i0[10] ), .A3(\SB3_4/i0[6] ), 
        .ZN(\SB3_4/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U2593 ( .A1(\SB3_4/i0_3 ), .A2(\SB3_4/i0_4 ), .A3(\SB3_4/i1[9] ), 
        .ZN(\SB3_4/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2595 ( .A1(\SB3_4/i0[9] ), .A2(\SB3_4/i0[10] ), .A3(\SB3_4/i0_3 ), 
        .ZN(\SB3_4/Component_Function_4/NAND4_in[2] ) );
  INV_X1 U2597 ( .I(n339), .ZN(\SB1_0_0/i1_7 ) );
  BUF_X1 U2598 ( .I(n339), .Z(n6028) );
  INV_X1 U2600 ( .I(\MC_ARK_ARC_1_1/buf_output[132] ), .ZN(\SB1_2_9/i3[0] ) );
  CLKBUF_X4 U2603 ( .I(\MC_ARK_ARC_1_1/buf_output[135] ), .Z(\SB1_2_9/i0[10] )
         );
  BUF_X4 U2604 ( .I(\MC_ARK_ARC_1_1/buf_output[136] ), .Z(\SB1_2_9/i0_4 ) );
  CLKBUF_X4 U2606 ( .I(\SB1_1_2/buf_output[3] ), .Z(\SB2_1_0/i0[10] ) );
  CLKBUF_X4 U2607 ( .I(\MC_ARK_ARC_1_0/buf_output[101] ), .Z(\SB1_1_15/i0_3 )
         );
  INV_X1 U2608 ( .I(\MC_ARK_ARC_1_1/buf_output[179] ), .ZN(\SB1_2_2/i1_5 ) );
  CLKBUF_X4 U2610 ( .I(\MC_ARK_ARC_1_2/buf_output[120] ), .Z(\SB1_3_11/i0[9] )
         );
  CLKBUF_X12 U2612 ( .I(Key[75]), .Z(n177) );
  CLKBUF_X4 U2615 ( .I(\SB2_0_16/buf_output[2] ), .Z(\RI5[0][110] ) );
  NAND3_X1 U2619 ( .A1(\SB1_1_16/i0[10] ), .A2(\SB1_1_16/i0_4 ), .A3(
        \SB1_1_16/i0_3 ), .ZN(\SB1_1_16/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U2620 ( .A1(\SB1_1_16/i0_4 ), .A2(\SB1_1_16/i1_7 ), .A3(
        \SB1_1_16/i0[8] ), .ZN(n2792) );
  NAND3_X1 U2624 ( .A1(\SB1_1_16/i0_4 ), .A2(\SB1_1_16/i1[9] ), .A3(
        \SB1_1_16/i0_3 ), .ZN(\SB1_1_16/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2625 ( .A1(\SB1_1_16/i0_0 ), .A2(\SB1_1_16/i0_3 ), .A3(
        \SB1_1_16/i0_4 ), .ZN(\SB1_1_16/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U2626 ( .A1(\SB1_1_16/i0_4 ), .A2(\SB1_1_16/i1[9] ), .A3(
        \SB1_1_16/i1_5 ), .ZN(\SB1_1_16/Component_Function_4/NAND4_in[3] ) );
  BUF_X4 U2630 ( .I(\SB1_3_28/buf_output[5] ), .Z(\SB2_3_28/i0_3 ) );
  CLKBUF_X4 U2634 ( .I(n419), .Z(\SB1_0_17/i0_3 ) );
  INV_X1 U2640 ( .I(\SB1_0_27/buf_output[5] ), .ZN(\SB2_0_27/i1_5 ) );
  CLKBUF_X4 U2643 ( .I(\SB1_0_27/buf_output[5] ), .Z(\SB2_0_27/i0_3 ) );
  INV_X1 U2651 ( .I(\MC_ARK_ARC_1_2/buf_output[39] ), .ZN(\SB1_3_25/i0[8] ) );
  BUF_X2 U2652 ( .I(\MC_ARK_ARC_1_2/buf_output[39] ), .Z(\SB1_3_25/i0[10] ) );
  INV_X1 U2656 ( .I(\SB1_3_21/buf_output[1] ), .ZN(\SB2_3_17/i1_7 ) );
  NAND3_X1 U2659 ( .A1(\SB1_3_7/i0_0 ), .A2(\SB1_3_7/i0[6] ), .A3(
        \SB1_3_7/i0[10] ), .ZN(\SB1_3_7/Component_Function_5/NAND4_in[1] ) );
  CLKBUF_X4 U2660 ( .I(\SB2_2_4/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[177] ) );
  NAND3_X1 U2661 ( .A1(\SB1_0_10/i0_3 ), .A2(\SB1_0_10/i0_0 ), .A3(
        \SB1_0_10/i0[7] ), .ZN(\SB1_0_10/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2662 ( .A1(\SB1_0_10/i1[9] ), .A2(\SB1_0_10/i0_4 ), .A3(
        \SB1_0_10/i0_3 ), .ZN(\SB1_0_10/Component_Function_5/NAND4_in[2] ) );
  INV_X1 U2664 ( .I(\MC_ARK_ARC_1_0/buf_output[13] ), .ZN(\SB1_1_29/i1_7 ) );
  BUF_X4 U2666 ( .I(\MC_ARK_ARC_1_0/buf_output[51] ), .Z(\SB1_1_23/i0[10] ) );
  INV_X1 U2671 ( .I(\SB2_2_8/i0_4 ), .ZN(\SB2_2_8/i0[7] ) );
  INV_X1 U2673 ( .I(\MC_ARK_ARC_1_1/buf_output[176] ), .ZN(\SB1_2_2/i1[9] ) );
  CLKBUF_X4 U2674 ( .I(\MC_ARK_ARC_1_1/buf_output[176] ), .Z(\SB1_2_2/i0_0 )
         );
  BUF_X4 U2675 ( .I(\SB1_1_13/buf_output[1] ), .Z(\SB2_1_9/i0[6] ) );
  INV_X1 U2676 ( .I(\SB1_3_24/buf_output[5] ), .ZN(\SB2_3_24/i1_5 ) );
  NAND3_X1 U2683 ( .A1(\SB1_2_12/i0[8] ), .A2(\SB1_2_12/i3[0] ), .A3(
        \SB1_2_12/i1_5 ), .ZN(n6091) );
  NAND3_X1 U2686 ( .A1(\SB1_2_12/i0_3 ), .A2(\SB1_2_12/i1_7 ), .A3(
        \SB1_2_12/i0[8] ), .ZN(\SB1_2_12/Component_Function_1/NAND4_in[1] ) );
  CLKBUF_X4 U2689 ( .I(n430), .Z(\SB1_0_6/i0_3 ) );
  INV_X1 U2691 ( .I(n430), .ZN(\SB1_0_6/i1_5 ) );
  NAND3_X1 U2693 ( .A1(\SB2_2_1/i0[10] ), .A2(\SB2_2_1/i0_3 ), .A3(
        \SB2_2_1/i0_4 ), .ZN(n6385) );
  NAND3_X1 U2695 ( .A1(\SB2_2_1/i0_3 ), .A2(\SB2_2_1/i1[9] ), .A3(
        \SB2_2_1/i0[6] ), .ZN(\SB2_2_1/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U2697 ( .A1(\SB2_2_1/i0_3 ), .A2(\SB2_2_1/i1_7 ), .A3(
        \SB2_2_1/i0[8] ), .ZN(\SB2_2_1/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 U2707 ( .A1(\SB2_2_1/i0_3 ), .A2(\SB2_2_1/i1[9] ), .ZN(
        \SB2_2_1/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U2708 ( .A1(\SB2_2_1/i0_3 ), .A2(\SB2_2_1/i0[8] ), .A3(
        \SB2_2_1/i0[9] ), .ZN(\SB2_2_1/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2710 ( .A1(\SB2_2_1/i0_3 ), .A2(\SB2_2_1/i0_0 ), .A3(
        \SB2_2_1/i0[7] ), .ZN(n5188) );
  NAND3_X1 U2711 ( .A1(\SB2_2_1/i0_3 ), .A2(\SB2_2_1/i0_4 ), .A3(
        \SB2_2_1/i0_0 ), .ZN(n3437) );
  NAND3_X1 U2716 ( .A1(\SB2_0_8/i0[9] ), .A2(\SB2_0_8/i0[6] ), .A3(
        \RI3[0][142] ), .ZN(\SB2_0_8/Component_Function_5/NAND4_in[3] ) );
  INV_X1 U2718 ( .I(\SB1_2_31/buf_output[1] ), .ZN(\SB2_2_27/i1_7 ) );
  BUF_X4 U2725 ( .I(\RI3[0][182] ), .Z(\SB2_0_1/i0_0 ) );
  INV_X1 U2726 ( .I(\RI1[3][89] ), .ZN(\SB1_3_17/i1_5 ) );
  NAND3_X1 U2727 ( .A1(\SB1_2_5/i3[0] ), .A2(\SB1_2_5/i0_0 ), .A3(
        \SB1_2_5/i1_7 ), .ZN(\SB1_2_5/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U2730 ( .A1(\SB1_2_5/i0_3 ), .A2(\SB1_2_5/i0[8] ), .A3(
        \SB1_2_5/i1_7 ), .ZN(\SB1_2_5/Component_Function_1/NAND4_in[1] ) );
  INV_X1 U2741 ( .I(\MC_ARK_ARC_1_1/buf_output[157] ), .ZN(\SB1_2_5/i1_7 ) );
  BUF_X2 U2743 ( .I(\MC_ARK_ARC_1_1/buf_output[140] ), .Z(\SB1_2_8/i0_0 ) );
  CLKBUF_X4 U2747 ( .I(\MC_ARK_ARC_1_1/buf_output[116] ), .Z(\SB1_2_12/i0_0 )
         );
  INV_X1 U2748 ( .I(n268), .ZN(\SB1_0_24/i1[9] ) );
  BUF_X2 U2749 ( .I(n268), .Z(\SB1_0_24/i0_0 ) );
  NAND3_X2 U2750 ( .A1(\SB2_0_29/i1_7 ), .A2(\SB2_0_29/i0[8] ), .A3(
        \SB2_0_29/i0_4 ), .ZN(\SB2_0_29/Component_Function_1/NAND4_in[3] ) );
  BUF_X2 U2751 ( .I(\MC_ARK_ARC_1_2/buf_output[96] ), .Z(\SB1_3_15/i0[9] ) );
  CLKBUF_X4 U2752 ( .I(\MC_ARK_ARC_1_1/buf_output[190] ), .Z(\SB1_2_0/i0_4 )
         );
  NAND3_X1 U2753 ( .A1(\SB2_2_16/i0_3 ), .A2(\SB2_2_16/i1_7 ), .A3(
        \SB2_2_16/i0[8] ), .ZN(\SB2_2_16/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 U2762 ( .A1(\SB2_2_16/i0_3 ), .A2(\SB2_2_16/i1[9] ), .ZN(
        \SB2_2_16/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U2765 ( .A1(\SB2_2_16/i0[9] ), .A2(\SB2_2_16/i0_3 ), .A3(
        \SB2_2_16/i0[10] ), .ZN(\SB2_2_16/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U2766 ( .A1(\SB2_2_16/i0_3 ), .A2(\SB2_2_16/i0_0 ), .A3(
        \SB2_2_16/i0_4 ), .ZN(n5638) );
  NAND3_X1 U2768 ( .A1(\SB2_2_16/i0_3 ), .A2(\SB2_2_16/i0_4 ), .A3(
        \SB2_2_16/i1[9] ), .ZN(\SB2_2_16/Component_Function_5/NAND4_in[2] ) );
  INV_X1 U2773 ( .I(\MC_ARK_ARC_1_0/buf_output[14] ), .ZN(\SB1_1_29/i1[9] ) );
  BUF_X4 U2777 ( .I(\MC_ARK_ARC_1_0/buf_output[14] ), .Z(\SB1_1_29/i0_0 ) );
  BUF_X2 U2778 ( .I(\MC_ARK_ARC_1_1/buf_output[60] ), .Z(\SB1_2_21/i0[9] ) );
  INV_X1 U2784 ( .I(\MC_ARK_ARC_1_1/buf_output[60] ), .ZN(\SB1_2_21/i3[0] ) );
  NAND3_X1 U2787 ( .A1(\SB1_3_11/i0_3 ), .A2(\SB1_3_11/i0[10] ), .A3(
        \SB1_3_11/i0[6] ), .ZN(\SB1_3_11/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U2788 ( .A1(\SB1_3_11/i0[9] ), .A2(\SB1_3_11/i0_3 ), .A3(
        \SB1_3_11/i0[10] ), .ZN(n5136) );
  NAND3_X1 U2789 ( .A1(\SB1_3_11/i0[9] ), .A2(\SB1_3_11/i0_3 ), .A3(
        \SB1_3_11/i0[8] ), .ZN(\SB1_3_11/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2792 ( .A1(\SB1_3_6/i1[9] ), .A2(\SB1_3_6/i0_3 ), .A3(
        \SB1_3_6/i0[6] ), .ZN(\SB1_3_6/Component_Function_3/NAND4_in[0] ) );
  CLKBUF_X4 U2800 ( .I(\MC_ARK_ARC_1_2/buf_output[134] ), .Z(\SB1_3_9/i0_0 )
         );
  BUF_X4 U2804 ( .I(\MC_ARK_ARC_1_2/buf_output[45] ), .Z(\SB1_3_24/i0[10] ) );
  BUF_X4 U2807 ( .I(n247), .Z(\SB1_0_31/i0_0 ) );
  INV_X1 U2808 ( .I(\MC_ARK_ARC_1_0/buf_output[55] ), .ZN(\SB1_1_22/i1_7 ) );
  BUF_X2 U2810 ( .I(\MC_ARK_ARC_1_0/buf_output[55] ), .Z(\SB1_1_22/i0[6] ) );
  INV_X1 U2811 ( .I(\MC_ARK_ARC_1_3/buf_output[175] ), .ZN(\SB3_2/i1_7 ) );
  BUF_X2 U2813 ( .I(\MC_ARK_ARC_1_3/buf_output[175] ), .Z(\SB3_2/i0[6] ) );
  BUF_X2 U2814 ( .I(\MC_ARK_ARC_1_2/buf_output[20] ), .Z(\SB1_3_28/i0_0 ) );
  INV_X1 U2815 ( .I(\MC_ARK_ARC_1_2/buf_output[20] ), .ZN(\SB1_3_28/i1[9] ) );
  NAND3_X1 U2816 ( .A1(\SB2_0_30/i0[7] ), .A2(\SB2_0_30/i0[6] ), .A3(
        \SB2_0_30/i0[8] ), .ZN(n4164) );
  NAND3_X1 U2820 ( .A1(\SB1_1_9/i0_3 ), .A2(\SB1_1_9/i0[10] ), .A3(
        \SB1_1_9/i0[6] ), .ZN(\SB1_1_9/Component_Function_2/NAND4_in[1] ) );
  INV_X1 U2823 ( .I(\MC_ARK_ARC_1_2/buf_output[118] ), .ZN(\SB1_3_12/i0[7] )
         );
  NAND3_X1 U2825 ( .A1(\SB1_0_0/i0[7] ), .A2(\SB1_0_0/i0_3 ), .A3(
        \SB1_0_0/i0_0 ), .ZN(\SB1_0_0/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U2830 ( .A1(\SB1_0_0/i0_3 ), .A2(\SB1_0_0/i0[10] ), .A3(n1376), 
        .ZN(\SB1_0_0/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U2832 ( .A1(\SB1_0_0/i0_3 ), .A2(\SB1_0_0/i0[8] ), .A3(
        \SB1_0_0/i1_7 ), .ZN(\SB1_0_0/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U2833 ( .A1(\SB1_0_0/i0_3 ), .A2(\SB1_0_0/i0[8] ), .A3(
        \SB1_0_0/i0[9] ), .ZN(\SB1_0_0/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U2843 ( .A1(\SB1_0_0/i0[10] ), .A2(\SB1_0_0/i0_3 ), .A3(
        \SB1_0_0/i0[9] ), .ZN(n1131) );
  NAND2_X1 U2844 ( .A1(\SB1_0_0/i0_3 ), .A2(\SB1_0_0/i1[9] ), .ZN(
        \SB1_0_0/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U2851 ( .A1(\SB1_0_0/i0_3 ), .A2(n1376), .A3(\SB1_0_0/i1[9] ), .ZN(
        n759) );
  NAND3_X1 U2852 ( .A1(\SB1_0_0/i0_4 ), .A2(\SB1_0_0/i0_3 ), .A3(
        \SB1_0_0/i1[9] ), .ZN(\SB1_0_0/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U2855 ( .A1(\SB1_0_18/i0[9] ), .A2(\SB1_0_18/i0_0 ), .A3(
        \SB1_0_18/i0[8] ), .ZN(\SB1_0_18/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U2856 ( .A1(\SB1_0_18/i0[8] ), .A2(\SB1_0_18/i0_3 ), .A3(
        \SB1_0_18/i1_7 ), .ZN(\SB1_0_18/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U2857 ( .A1(\SB1_3_25/i0_3 ), .A2(\SB1_3_25/i1[9] ), .A3(
        \SB1_3_25/i0_4 ), .ZN(n5683) );
  NAND3_X1 U2859 ( .A1(\SB1_3_25/i0[10] ), .A2(\SB1_3_25/i1[9] ), .A3(
        \SB1_3_25/i1_7 ), .ZN(\SB1_3_25/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U2860 ( .A1(\SB1_3_25/i0[10] ), .A2(\SB1_3_25/i1[9] ), .A3(
        \SB1_3_25/i1_5 ), .ZN(n5244) );
  NAND3_X1 U2861 ( .A1(\SB2_0_16/i0_3 ), .A2(\SB2_0_16/i0_4 ), .A3(
        \SB2_0_16/i1[9] ), .ZN(\SB2_0_16/Component_Function_5/NAND4_in[2] ) );
  INV_X1 U2868 ( .I(\RI3[0][161] ), .ZN(\SB2_0_5/i1_5 ) );
  BUF_X4 U2871 ( .I(n310), .Z(\SB1_0_10/i0_0 ) );
  INV_X1 U2877 ( .I(\MC_ARK_ARC_1_1/buf_output[143] ), .ZN(\SB1_2_8/i1_5 ) );
  CLKBUF_X4 U2879 ( .I(\MC_ARK_ARC_1_1/buf_output[143] ), .Z(\SB1_2_8/i0_3 )
         );
  NAND3_X1 U2881 ( .A1(\SB2_0_14/i0_3 ), .A2(\SB2_0_14/i0[9] ), .A3(
        \RI3[0][105] ), .ZN(n6473) );
  NAND3_X1 U2886 ( .A1(\SB2_0_14/i0[8] ), .A2(\SB2_0_14/i0_3 ), .A3(
        \SB2_0_14/i1_7 ), .ZN(\SB2_0_14/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U2891 ( .A1(\RI3[0][105] ), .A2(\RI3[0][106] ), .A3(\SB2_0_14/i0_3 ), .ZN(\SB2_0_14/Component_Function_0/NAND4_in[2] ) );
  BUF_X4 U2892 ( .I(\RI3[0][86] ), .Z(\SB2_0_17/i0_0 ) );
  INV_X1 U2896 ( .I(n395), .ZN(\SB1_0_4/i0[8] ) );
  BUF_X2 U2897 ( .I(n395), .Z(\SB1_0_4/i0[10] ) );
  INV_X1 U2898 ( .I(\SB3_25/buf_output[2] ), .ZN(\SB4_22/i1[9] ) );
  NAND3_X1 U2900 ( .A1(\SB1_1_6/i1[9] ), .A2(\SB1_1_6/i1_5 ), .A3(
        \SB1_1_6/i0_4 ), .ZN(\SB1_1_6/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U2902 ( .A1(\SB1_1_6/i0_3 ), .A2(\SB1_1_6/i0_4 ), .A3(
        \SB1_1_6/i1[9] ), .ZN(n5462) );
  NAND3_X1 U2903 ( .A1(\SB1_1_6/i0_3 ), .A2(\SB1_1_6/i1[9] ), .A3(
        \SB1_1_6/i0[6] ), .ZN(n5484) );
  NAND2_X1 U2904 ( .A1(\SB1_1_6/i0_3 ), .A2(\SB1_1_6/i1[9] ), .ZN(
        \SB1_1_6/Component_Function_1/NAND4_in[0] ) );
  AND2_X2 U2911 ( .A1(\MC_ARK_ARC_1_2/buf_output[166] ), .A2(
        \MC_ARK_ARC_1_2/buf_output[163] ), .Z(n3122) );
  INV_X1 U2913 ( .I(\MC_ARK_ARC_1_2/buf_output[163] ), .ZN(\SB1_3_4/i1_7 ) );
  BUF_X2 U2914 ( .I(\MC_ARK_ARC_1_2/buf_output[163] ), .Z(\SB1_3_4/i0[6] ) );
  CLKBUF_X4 U2923 ( .I(\MC_ARK_ARC_1_2/buf_output[53] ), .Z(\SB1_3_23/i0_3 )
         );
  CLKBUF_X4 U2924 ( .I(\MC_ARK_ARC_1_2/buf_output[119] ), .Z(\SB1_3_12/i0_3 )
         );
  AND2_X2 U2926 ( .A1(\MC_ARK_ARC_1_2/buf_output[120] ), .A2(
        \MC_ARK_ARC_1_2/buf_output[124] ), .Z(n5539) );
  INV_X1 U2939 ( .I(\MC_ARK_ARC_1_2/buf_output[120] ), .ZN(\SB1_3_11/i3[0] )
         );
  INV_X1 U2940 ( .I(n425), .ZN(\SB1_0_11/i1_5 ) );
  CLKBUF_X4 U2942 ( .I(\SB1_1_11/buf_output[3] ), .Z(\SB2_1_9/i0[10] ) );
  BUF_X2 U2943 ( .I(\MC_ARK_ARC_1_0/buf_output[104] ), .Z(\SB1_1_14/i0_0 ) );
  INV_X1 U2950 ( .I(\MC_ARK_ARC_1_1/buf_output[13] ), .ZN(\SB1_2_29/i1_7 ) );
  NAND2_X2 U2951 ( .A1(\SB1_3_12/i0[10] ), .A2(\SB1_3_12/i0[9] ), .ZN(
        \SB1_3_12/Component_Function_0/NAND4_in[0] ) );
  BUF_X2 U2953 ( .I(\MC_ARK_ARC_1_2/buf_output[114] ), .Z(\SB1_3_12/i0[9] ) );
  NAND2_X2 U2956 ( .A1(\SB3_1/i0_0 ), .A2(\SB3_1/i3[0] ), .ZN(
        \SB3_1/Component_Function_5/NAND4_in[0] ) );
  CLKBUF_X4 U2957 ( .I(\SB2_3_9/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[152] ) );
  INV_X1 U2961 ( .I(n298), .ZN(\SB1_0_14/i1[9] ) );
  BUF_X2 U2962 ( .I(n298), .Z(\SB1_0_14/i0_0 ) );
  CLKBUF_X4 U2964 ( .I(\SB3_5/buf_output[2] ), .Z(\SB4_2/i0_0 ) );
  CLKBUF_X4 U2966 ( .I(\SB3_23/buf_output[4] ), .Z(\SB4_22/i0_4 ) );
  BUF_X2 U2967 ( .I(\SB3_17/buf_output[1] ), .Z(\SB4_13/i0[6] ) );
  CLKBUF_X4 U2971 ( .I(\SB3_2/buf_output[2] ), .Z(\SB4_31/i0_0 ) );
  CLKBUF_X4 U2976 ( .I(\SB4_29/i0_4 ), .Z(n1793) );
  CLKBUF_X4 U2982 ( .I(\SB3_9/buf_output[5] ), .Z(\SB4_9/i0_3 ) );
  CLKBUF_X4 U2983 ( .I(\SB3_4/buf_output[3] ), .Z(\SB4_2/i0[10] ) );
  BUF_X2 U2989 ( .I(\SB3_10/buf_output[1] ), .Z(\SB4_6/i0[6] ) );
  CLKBUF_X4 U2994 ( .I(\SB3_0/buf_output[5] ), .Z(\SB4_0/i0_3 ) );
  BUF_X2 U3001 ( .I(\SB3_0/buf_output[1] ), .Z(\SB4_28/i0[6] ) );
  BUF_X2 U3002 ( .I(\SB3_28/buf_output[4] ), .Z(\SB4_27/i0_4 ) );
  INV_X4 U3005 ( .I(\RI1[4][155] ), .ZN(\SB3_6/i1_5 ) );
  CLKBUF_X8 U3010 ( .I(\RI1[4][65] ), .Z(\SB3_21/i0_3 ) );
  CLKBUF_X4 U3011 ( .I(\MC_ARK_ARC_1_3/buf_output[92] ), .Z(\SB3_16/i0_0 ) );
  CLKBUF_X4 U3013 ( .I(n5508), .Z(\SB3_30/i0_3 ) );
  CLKBUF_X4 U3022 ( .I(\SB2_3_13/buf_output[5] ), .Z(\RI5[3][113] ) );
  BUF_X4 U3023 ( .I(\SB2_3_11/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[135] ) );
  CLKBUF_X4 U3029 ( .I(\SB2_3_4/buf_output[0] ), .Z(\RI5[3][0] ) );
  NAND3_X2 U3032 ( .A1(\SB2_3_11/i0[6] ), .A2(n4768), .A3(n5240), .ZN(
        \SB2_3_11/Component_Function_1/NAND4_in[2] ) );
  CLKBUF_X2 U3033 ( .I(\SB1_3_16/buf_output[0] ), .Z(n5240) );
  CLKBUF_X4 U3035 ( .I(\SB1_3_7/buf_output[3] ), .Z(\SB2_3_5/i0[10] ) );
  BUF_X4 U3036 ( .I(\SB1_3_10/buf_output[2] ), .Z(\SB2_3_7/i0_0 ) );
  CLKBUF_X4 U3037 ( .I(\SB1_3_24/buf_output[5] ), .Z(\SB2_3_24/i0_3 ) );
  CLKBUF_X4 U3038 ( .I(\SB1_3_30/buf_output[2] ), .Z(\SB2_3_27/i0_0 ) );
  CLKBUF_X4 U3040 ( .I(\SB1_3_23/buf_output[3] ), .Z(\SB2_3_21/i0[10] ) );
  BUF_X2 U3041 ( .I(\SB1_3_3/buf_output[0] ), .Z(\SB2_3_30/i0[9] ) );
  BUF_X4 U3043 ( .I(\SB1_3_11/buf_output[5] ), .Z(\SB2_3_11/i0_3 ) );
  CLKBUF_X8 U3048 ( .I(\RI1[3][131] ), .Z(\SB1_3_10/i0_3 ) );
  BUF_X2 U3049 ( .I(\MC_ARK_ARC_1_2/buf_output[36] ), .Z(\SB1_3_25/i0[9] ) );
  CLKBUF_X4 U3054 ( .I(\MC_ARK_ARC_1_2/buf_output[26] ), .Z(\SB1_3_27/i0_0 )
         );
  CLKBUF_X4 U3059 ( .I(\MC_ARK_ARC_1_2/buf_output[98] ), .Z(\SB1_3_15/i0_0 )
         );
  CLKBUF_X4 U3060 ( .I(\MC_ARK_ARC_1_2/buf_output[57] ), .Z(\SB1_3_22/i0[10] )
         );
  CLKBUF_X4 U3067 ( .I(\MC_ARK_ARC_1_2/buf_output[0] ), .Z(\SB1_3_31/i0[9] )
         );
  BUF_X2 U3068 ( .I(\MC_ARK_ARC_1_2/buf_output[60] ), .Z(\SB1_3_21/i0[9] ) );
  CLKBUF_X4 U3070 ( .I(\MC_ARK_ARC_1_2/buf_output[21] ), .Z(\SB1_3_28/i0[10] )
         );
  CLKBUF_X4 U3075 ( .I(\MC_ARK_ARC_1_2/buf_output[142] ), .Z(\SB1_3_8/i0_4 )
         );
  CLKBUF_X4 U3077 ( .I(\SB2_2_3/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[183] ) );
  CLKBUF_X4 U3083 ( .I(\SB2_2_8/buf_output[5] ), .Z(\RI5[2][143] ) );
  BUF_X4 U3084 ( .I(\SB2_2_27/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[39] ) );
  CLKBUF_X4 U3086 ( .I(\SB2_2_25/buf_output[3] ), .Z(\RI5[2][51] ) );
  INV_X1 U3092 ( .I(n5057), .ZN(n2894) );
  BUF_X4 U3093 ( .I(\SB2_2_5/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[186] ) );
  CLKBUF_X4 U3094 ( .I(\SB2_2_31/buf_output[4] ), .Z(\RI5[2][10] ) );
  CLKBUF_X4 U3095 ( .I(\SB1_2_29/buf_output[1] ), .Z(\SB2_2_25/i0[6] ) );
  CLKBUF_X4 U3097 ( .I(\SB1_2_24/buf_output[1] ), .Z(\SB2_2_20/i0[6] ) );
  CLKBUF_X4 U3105 ( .I(\SB1_2_1/buf_output[1] ), .Z(\SB2_2_29/i0[6] ) );
  CLKBUF_X4 U3106 ( .I(\SB1_2_14/buf_output[3] ), .Z(\SB2_2_12/i0[10] ) );
  CLKBUF_X4 U3109 ( .I(\SB1_2_7/buf_output[1] ), .Z(\SB2_2_3/i0[6] ) );
  CLKBUF_X4 U3111 ( .I(\SB1_2_9/buf_output[2] ), .Z(\SB2_2_6/i0_0 ) );
  CLKBUF_X4 U3112 ( .I(\SB1_2_28/buf_output[2] ), .Z(\SB2_2_25/i0_0 ) );
  CLKBUF_X4 U3113 ( .I(\SB1_2_22/buf_output[3] ), .Z(\SB2_2_20/i0[10] ) );
  NAND2_X1 U3116 ( .A1(n1556), .A2(\SB1_2_4/Component_Function_4/NAND4_in[3] ), 
        .ZN(n1555) );
  CLKBUF_X4 U3118 ( .I(\SB1_2_10/buf_output[3] ), .Z(\SB2_2_8/i0[10] ) );
  NAND3_X2 U3119 ( .A1(\SB1_2_30/i0[9] ), .A2(\SB1_2_30/i0_0 ), .A3(
        \SB1_2_30/i0[8] ), .ZN(\SB1_2_30/Component_Function_4/NAND4_in[0] ) );
  CLKBUF_X4 U3121 ( .I(\MC_ARK_ARC_1_1/buf_output[183] ), .Z(\SB1_2_1/i0[10] )
         );
  CLKBUF_X4 U3124 ( .I(\MC_ARK_ARC_1_1/buf_output[9] ), .Z(\SB1_2_30/i0[10] )
         );
  CLKBUF_X4 U3133 ( .I(\MC_ARK_ARC_1_1/buf_output[122] ), .Z(\SB1_2_11/i0_0 )
         );
  CLKBUF_X4 U3141 ( .I(\MC_ARK_ARC_1_1/buf_output[87] ), .Z(\SB1_2_17/i0[10] )
         );
  CLKBUF_X4 U3143 ( .I(\MC_ARK_ARC_1_1/buf_output[162] ), .Z(\SB1_2_4/i0[9] )
         );
  CLKBUF_X4 U3144 ( .I(\SB2_1_10/buf_output[2] ), .Z(\RI5[1][146] ) );
  BUF_X4 U3145 ( .I(\SB2_1_25/buf_output[4] ), .Z(\RI5[1][46] ) );
  CLKBUF_X4 U3148 ( .I(\SB2_1_16/buf_output[1] ), .Z(\RI5[1][115] ) );
  CLKBUF_X4 U3153 ( .I(\SB1_1_30/buf_output[1] ), .Z(\SB2_1_26/i0[6] ) );
  BUF_X4 U3154 ( .I(\SB2_1_3/i0_4 ), .Z(n5208) );
  CLKBUF_X2 U3155 ( .I(\SB1_1_0/buf_output[5] ), .Z(n5042) );
  CLKBUF_X4 U3158 ( .I(\SB1_1_2/buf_output[4] ), .Z(\SB2_1_1/i0_4 ) );
  BUF_X4 U3162 ( .I(\SB1_1_26/buf_output[5] ), .Z(\SB2_1_26/i0_3 ) );
  NAND2_X1 U3163 ( .A1(\SB1_1_6/Component_Function_4/NAND4_in[2] ), .A2(n6104), 
        .ZN(n1190) );
  NAND3_X2 U3168 ( .A1(\SB1_1_30/i0_3 ), .A2(\SB1_1_30/i0[10] ), .A3(
        \SB1_1_30/i0[6] ), .ZN(\SB1_1_30/Component_Function_2/NAND4_in[1] ) );
  CLKBUF_X4 U3169 ( .I(\MC_ARK_ARC_1_0/buf_output[128] ), .Z(\SB1_1_10/i0_0 )
         );
  CLKBUF_X4 U3171 ( .I(\MC_ARK_ARC_1_0/buf_output[182] ), .Z(\SB1_1_1/i0_0 )
         );
  CLKBUF_X4 U3172 ( .I(\MC_ARK_ARC_1_0/buf_output[188] ), .Z(\SB1_1_0/i0_0 )
         );
  CLKBUF_X4 U3176 ( .I(\MC_ARK_ARC_1_0/buf_output[176] ), .Z(\SB1_1_2/i0_0 )
         );
  CLKBUF_X4 U3177 ( .I(\MC_ARK_ARC_1_0/buf_output[63] ), .Z(\SB1_1_21/i0[10] )
         );
  CLKBUF_X4 U3181 ( .I(\SB2_0_24/buf_output[3] ), .Z(\RI5[0][57] ) );
  CLKBUF_X4 U3182 ( .I(\SB2_0_14/buf_output[3] ), .Z(\RI5[0][117] ) );
  BUF_X4 U3188 ( .I(\SB2_0_26/buf_output[4] ), .Z(\RI5[0][40] ) );
  CLKBUF_X2 U3190 ( .I(n2753), .Z(n5054) );
  INV_X4 U3191 ( .I(n5644), .ZN(\SB2_0_2/i0[10] ) );
  CLKBUF_X4 U3194 ( .I(\SB1_0_12/buf_output[5] ), .Z(\SB2_0_12/i0_3 ) );
  NAND2_X1 U3196 ( .A1(\SB1_0_20/Component_Function_4/NAND4_in[2] ), .A2(n6347), .ZN(n6439) );
  NAND2_X1 U3197 ( .A1(\SB1_0_17/Component_Function_4/NAND4_in[3] ), .A2(n5673), .ZN(n2037) );
  CLKBUF_X4 U3201 ( .I(n365), .Z(\SB1_0_19/i0[10] ) );
  BUF_X2 U3202 ( .I(n320), .Z(\SB1_0_6/i0[9] ) );
  CLKBUF_X4 U3206 ( .I(n265), .Z(\SB1_0_25/i0_0 ) );
  BUF_X2 U3211 ( .I(n348), .Z(\SB1_0_28/i0_4 ) );
  CLKBUF_X4 U3219 ( .I(n388), .Z(\SB1_0_8/i0_4 ) );
  CLKBUF_X4 U3220 ( .I(n292), .Z(\SB1_0_16/i0_0 ) );
  BUF_X2 U3223 ( .I(n258), .Z(\SB1_0_27/i0[6] ) );
  BUF_X4 U3225 ( .I(n372), .Z(n4752) );
  CLKBUF_X4 U3226 ( .I(n368), .Z(n4753) );
  NAND3_X1 U3227 ( .A1(\SB1_0_3/i0[10] ), .A2(\SB1_0_3/i1_7 ), .A3(
        \SB1_0_3/i1[9] ), .ZN(n1646) );
  NAND3_X1 U3228 ( .A1(\SB1_0_8/i1[9] ), .A2(\SB1_0_8/i1_5 ), .A3(
        \SB1_0_8/i0_4 ), .ZN(\SB1_0_8/Component_Function_4/NAND4_in[3] ) );
  CLKBUF_X4 U3230 ( .I(n396), .Z(\SB1_0_4/i0_4 ) );
  CLKBUF_X4 U3246 ( .I(n328), .Z(\SB1_0_4/i0_0 ) );
  INV_X1 U3250 ( .I(n263), .ZN(\SB1_0_25/i3[0] ) );
  NAND3_X1 U3256 ( .A1(\SB1_0_11/i1[9] ), .A2(\SB1_0_11/i1_5 ), .A3(
        \SB1_0_11/i0_4 ), .ZN(\SB1_0_11/Component_Function_4/NAND4_in[3] ) );
  NAND2_X1 U3257 ( .A1(\SB1_0_11/i0_0 ), .A2(\SB1_0_11/i3[0] ), .ZN(
        \SB1_0_11/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 U3258 ( .A1(\SB1_0_12/i0_3 ), .A2(\SB1_0_12/i1[9] ), .ZN(n3733) );
  NAND3_X1 U3263 ( .A1(\SB1_0_4/i0[7] ), .A2(\SB1_0_4/i0_3 ), .A3(
        \SB1_0_4/i0_0 ), .ZN(\SB1_0_4/Component_Function_0/NAND4_in[3] ) );
  BUF_X2 U3271 ( .I(n338), .Z(\SB1_0_0/i0[9] ) );
  NAND2_X1 U3280 ( .A1(\SB1_0_8/i0_3 ), .A2(\SB1_0_8/i1[9] ), .ZN(
        \SB1_0_8/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U3281 ( .A1(\SB1_0_6/i0[6] ), .A2(\SB1_0_6/i1[9] ), .A3(
        \SB1_0_6/i0_3 ), .ZN(\SB1_0_6/Component_Function_3/NAND4_in[0] ) );
  NAND2_X1 U3288 ( .A1(\SB1_0_12/i0_0 ), .A2(\SB1_0_12/i3[0] ), .ZN(
        \SB1_0_12/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U3303 ( .A1(\SB1_0_8/i0_3 ), .A2(\SB1_0_8/i0_0 ), .A3(
        \SB1_0_8/i0_4 ), .ZN(n2534) );
  NAND3_X1 U3307 ( .A1(\SB1_0_28/i0_3 ), .A2(\SB1_0_28/i0_0 ), .A3(
        \SB1_0_28/i0_4 ), .ZN(\SB1_0_28/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3308 ( .A1(\SB1_0_18/i0_3 ), .A2(n1367), .A3(\SB1_0_18/i0[6] ), 
        .ZN(n1581) );
  NAND2_X1 U3321 ( .A1(\SB1_0_7/i0_3 ), .A2(\SB1_0_7/i1[9] ), .ZN(
        \SB1_0_7/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U3323 ( .A1(\SB1_0_25/i0[7] ), .A2(\SB1_0_25/i0_3 ), .A3(
        \SB1_0_25/i0_0 ), .ZN(\SB1_0_25/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 U3327 ( .A1(\SB1_0_25/i0_3 ), .A2(\SB1_0_25/i1[9] ), .ZN(
        \SB1_0_25/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U3330 ( .A1(\SB1_0_0/i0_0 ), .A2(\SB1_0_0/i0_4 ), .A3(
        \SB1_0_0/i1_5 ), .ZN(n6474) );
  NAND2_X1 U3340 ( .A1(\SB1_0_5/i0_3 ), .A2(\SB1_0_5/i1[9] ), .ZN(n6332) );
  CLKBUF_X4 U3342 ( .I(n386), .Z(\SB1_0_9/i0_4 ) );
  NAND3_X1 U3343 ( .A1(\SB1_0_3/i0[7] ), .A2(\SB1_0_3/i0_3 ), .A3(
        \SB1_0_3/i0_0 ), .ZN(\SB1_0_3/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U3359 ( .A1(\SB1_0_2/i0_4 ), .A2(\SB1_0_2/i0_0 ), .A3(
        \SB1_0_2/i0_3 ), .ZN(\SB1_0_2/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3362 ( .A1(\SB1_0_0/i0_4 ), .A2(\SB1_0_0/i0[9] ), .A3(n6028), .ZN(
        n6482) );
  NAND3_X1 U3369 ( .A1(\SB2_0_30/i0[9] ), .A2(\SB2_0_30/i0[6] ), .A3(
        \RI3[0][10] ), .ZN(n5279) );
  NAND3_X1 U3373 ( .A1(\SB2_0_15/i0_3 ), .A2(\SB2_0_15/i0_0 ), .A3(
        \RI3[0][100] ), .ZN(\SB2_0_15/Component_Function_3/NAND4_in[1] ) );
  NAND2_X1 U3374 ( .A1(\SB2_0_19/i0_0 ), .A2(\SB2_0_19/i3[0] ), .ZN(
        \SB2_0_19/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U3375 ( .A1(\SB2_0_30/i3[0] ), .A2(\SB2_0_30/i0_0 ), .A3(
        \SB2_0_30/i1_7 ), .ZN(\SB2_0_30/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U3376 ( .A1(\SB2_0_16/i1_7 ), .A2(\SB2_0_16/i0[8] ), .A3(
        \SB2_0_16/i0_4 ), .ZN(\SB2_0_16/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U3382 ( .A1(\SB2_0_9/i0_3 ), .A2(\SB2_0_9/i1_7 ), .A3(
        \SB2_0_9/i0[8] ), .ZN(\SB2_0_9/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U3383 ( .A1(n571), .A2(\SB2_0_10/i0_0 ), .A3(\SB2_0_10/i0[8] ), 
        .ZN(\SB2_0_10/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U3385 ( .A1(\SB2_0_31/i0[10] ), .A2(\SB2_0_31/i0_0 ), .A3(
        \SB2_0_31/i0[6] ), .ZN(\SB2_0_31/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U3386 ( .A1(\SB2_0_24/i0[10] ), .A2(\SB2_0_24/i0_3 ), .A3(
        \SB2_0_24/i0[9] ), .ZN(\SB2_0_24/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U3388 ( .A1(\SB2_0_11/i1_5 ), .A2(\SB2_0_11/i0[10] ), .A3(
        \SB2_0_11/i1[9] ), .ZN(\SB2_0_11/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U3389 ( .A1(\SB2_0_23/i0[10] ), .A2(\SB2_0_23/i0_3 ), .A3(
        \SB2_0_23/i0[9] ), .ZN(n3526) );
  NAND3_X1 U3390 ( .A1(\SB2_0_7/i0[9] ), .A2(\SB2_0_7/i0_0 ), .A3(
        \SB2_0_7/i0[8] ), .ZN(\SB2_0_7/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U3391 ( .A1(\SB2_0_8/i1[9] ), .A2(\SB2_0_8/i0_3 ), .A3(
        \SB2_0_8/i0[6] ), .ZN(\SB2_0_8/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U3395 ( .A1(\SB2_0_23/i0[8] ), .A2(n2877), .A3(\SB2_0_23/i0[6] ), 
        .ZN(\SB2_0_23/Component_Function_0/NAND4_in[1] ) );
  NAND2_X1 U3402 ( .A1(\SB2_0_27/i0[10] ), .A2(n2679), .ZN(
        \SB2_0_27/Component_Function_0/NAND4_in[0] ) );
  CLKBUF_X4 U3406 ( .I(\SB1_0_15/buf_output[4] ), .Z(\RI3[0][106] ) );
  NAND3_X1 U3408 ( .A1(\SB2_0_21/i0_3 ), .A2(\SB2_0_21/i0[10] ), .A3(
        \SB2_0_21/i0[6] ), .ZN(\SB2_0_21/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U3410 ( .A1(\RI3[0][160] ), .A2(n3689), .A3(\SB2_0_5/i1_5 ), .ZN(
        n6224) );
  NAND3_X1 U3416 ( .A1(\SB2_0_20/i0_3 ), .A2(\SB2_0_20/i1_7 ), .A3(
        \SB2_0_20/i0[8] ), .ZN(\SB2_0_20/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U3424 ( .A1(\SB2_0_9/i0[10] ), .A2(\SB2_0_9/i0_4 ), .A3(
        \SB2_0_9/i0_3 ), .ZN(\SB2_0_9/Component_Function_0/NAND4_in[2] ) );
  CLKBUF_X4 U3425 ( .I(\SB2_0_24/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[67] ) );
  CLKBUF_X4 U3430 ( .I(\SB2_0_17/buf_output[4] ), .Z(\RI5[0][94] ) );
  INV_X1 U3431 ( .I(\MC_ARK_ARC_1_0/buf_output[144] ), .ZN(\SB1_1_7/i3[0] ) );
  CLKBUF_X4 U3435 ( .I(\MC_ARK_ARC_1_0/buf_output[162] ), .Z(\SB1_1_4/i0[9] )
         );
  INV_X1 U3436 ( .I(\MC_ARK_ARC_1_0/buf_output[109] ), .ZN(\SB1_1_13/i1_7 ) );
  NAND3_X1 U3437 ( .A1(\SB1_1_31/i1[9] ), .A2(\SB1_1_31/i1_5 ), .A3(
        \SB1_1_31/i0_4 ), .ZN(\SB1_1_31/Component_Function_4/NAND4_in[3] ) );
  INV_X1 U3446 ( .I(\MC_ARK_ARC_1_0/buf_output[161] ), .ZN(\SB1_1_5/i1_5 ) );
  NAND3_X1 U3449 ( .A1(\SB1_1_25/i0[8] ), .A2(\SB1_1_25/i1_5 ), .A3(
        \SB1_1_25/i3[0] ), .ZN(n4691) );
  CLKBUF_X8 U3450 ( .I(\RI1[1][11] ), .Z(\SB1_1_30/i0_3 ) );
  NAND3_X1 U3452 ( .A1(\SB1_1_25/i0[8] ), .A2(\SB1_1_25/i0[9] ), .A3(
        \SB1_1_25/i0_3 ), .ZN(\SB1_1_25/Component_Function_2/NAND4_in[2] ) );
  CLKBUF_X4 U3454 ( .I(\MC_ARK_ARC_1_0/buf_output[180] ), .Z(\SB1_1_1/i0[9] )
         );
  NAND3_X1 U3458 ( .A1(\SB1_1_20/i0_3 ), .A2(\SB1_1_20/i0[8] ), .A3(
        \SB1_1_20/i0[9] ), .ZN(\SB1_1_20/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3459 ( .A1(\SB1_1_19/i0_0 ), .A2(\SB1_1_19/i0_3 ), .A3(
        \SB1_1_19/i0_4 ), .ZN(\SB1_1_19/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3461 ( .A1(\SB1_1_13/i0_0 ), .A2(\SB1_1_13/i1_7 ), .A3(
        \SB1_1_13/i3[0] ), .ZN(n1004) );
  NAND3_X1 U3462 ( .A1(\SB1_1_13/i0_3 ), .A2(\SB1_1_13/i0_4 ), .A3(
        \SB1_1_13/i1[9] ), .ZN(n5989) );
  NAND3_X1 U3466 ( .A1(\SB1_1_6/i0[10] ), .A2(\SB1_1_6/i0_4 ), .A3(
        \SB1_1_6/i0_3 ), .ZN(\SB1_1_6/Component_Function_0/NAND4_in[2] ) );
  CLKBUF_X4 U3476 ( .I(\MC_ARK_ARC_1_0/buf_output[186] ), .Z(\SB1_1_0/i0[9] )
         );
  NAND2_X1 U3478 ( .A1(\SB1_1_7/Component_Function_2/NAND4_in[3] ), .A2(
        \SB1_1_7/Component_Function_2/NAND4_in[1] ), .ZN(n5446) );
  NAND3_X1 U3481 ( .A1(\SB1_1_23/i0_3 ), .A2(\SB1_1_23/i1_7 ), .A3(
        \SB1_1_23/i0[8] ), .ZN(\SB1_1_23/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U3486 ( .A1(\SB1_1_16/i0[8] ), .A2(\SB1_1_16/i1_5 ), .A3(
        \SB1_1_16/i3[0] ), .ZN(n1342) );
  NAND3_X1 U3487 ( .A1(\SB1_1_27/i0[9] ), .A2(\SB1_1_27/i0[8] ), .A3(
        \SB1_1_27/i0_3 ), .ZN(n5867) );
  NAND3_X1 U3492 ( .A1(\SB1_1_3/i0[8] ), .A2(\SB1_1_3/i0[7] ), .A3(
        \SB1_1_3/i0[6] ), .ZN(\SB1_1_3/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U3493 ( .A1(\SB1_1_18/i0[10] ), .A2(\SB1_1_18/i1[9] ), .A3(
        \SB1_1_18/i1_7 ), .ZN(\SB1_1_18/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U3495 ( .A1(\SB1_1_28/i0[8] ), .A2(\SB1_1_28/i1_5 ), .A3(
        \SB1_1_28/i3[0] ), .ZN(n846) );
  NAND3_X1 U3499 ( .A1(\SB1_1_25/i0_4 ), .A2(\SB1_1_25/i0[8] ), .A3(
        \SB1_1_25/i1_7 ), .ZN(n1625) );
  NAND3_X1 U3500 ( .A1(\SB1_1_0/i0_0 ), .A2(\SB1_1_0/i0_3 ), .A3(
        \SB1_1_0/i0[7] ), .ZN(n1880) );
  CLKBUF_X4 U3502 ( .I(\SB1_1_8/buf_output[1] ), .Z(\SB2_1_4/i0[6] ) );
  CLKBUF_X4 U3506 ( .I(\SB1_1_30/buf_output[3] ), .Z(\SB2_1_28/i0[10] ) );
  NAND3_X1 U3509 ( .A1(\SB2_1_4/i0[9] ), .A2(\SB2_1_4/i0[6] ), .A3(
        \SB1_1_5/buf_output[4] ), .ZN(n3512) );
  CLKBUF_X4 U3510 ( .I(\SB1_1_26/buf_output[1] ), .Z(\SB2_1_22/i0[6] ) );
  CLKBUF_X4 U3511 ( .I(\SB1_1_17/buf_output[4] ), .Z(\SB2_1_16/i0_4 ) );
  CLKBUF_X4 U3517 ( .I(\SB1_1_20/buf_output[2] ), .Z(\SB2_1_17/i0_0 ) );
  CLKBUF_X4 U3522 ( .I(\SB1_1_12/buf_output[2] ), .Z(\SB2_1_9/i0_0 ) );
  NAND3_X1 U3528 ( .A1(\SB2_1_28/i0[8] ), .A2(\SB2_1_28/i0[7] ), .A3(
        \SB2_1_28/i0[6] ), .ZN(\SB2_1_28/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U3529 ( .A1(\SB2_1_23/i1_5 ), .A2(\SB2_1_23/i0[6] ), .A3(
        \SB2_1_23/i0[9] ), .ZN(\SB2_1_23/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U3531 ( .A1(\SB2_1_6/i1[9] ), .A2(\SB2_1_6/i1_5 ), .A3(
        \SB2_1_6/i0_4 ), .ZN(\SB2_1_6/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U3536 ( .A1(\SB2_1_21/i0[6] ), .A2(\RI3[1][60] ), .A3(
        \SB2_1_21/i1_5 ), .ZN(n4709) );
  NAND3_X1 U3538 ( .A1(\SB2_1_26/i0[8] ), .A2(\SB2_1_26/i0[7] ), .A3(
        \SB2_1_26/i0[6] ), .ZN(\SB2_1_26/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U3544 ( .A1(\SB2_1_30/i0_3 ), .A2(\SB2_1_30/i0[8] ), .A3(
        \SB2_1_30/i0[9] ), .ZN(\SB2_1_30/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3545 ( .A1(\SB2_1_30/i0_0 ), .A2(\SB2_1_30/i0_3 ), .A3(
        \SB2_1_30/i0_4 ), .ZN(\SB2_1_30/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3546 ( .A1(\SB2_1_11/i1_7 ), .A2(\SB2_1_11/i0[8] ), .A3(
        \SB1_1_12/buf_output[4] ), .ZN(
        \SB2_1_11/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U3552 ( .A1(\SB2_1_8/i0_4 ), .A2(\SB2_1_8/i1[9] ), .A3(
        \SB2_1_8/i1_5 ), .ZN(n6290) );
  NAND3_X1 U3556 ( .A1(\SB2_1_14/i1[9] ), .A2(\SB2_1_14/i1_5 ), .A3(
        \SB2_1_14/i0_4 ), .ZN(\SB2_1_14/Component_Function_4/NAND4_in[3] ) );
  NAND2_X1 U3562 ( .A1(\SB2_1_19/i0[10] ), .A2(\SB2_1_19/i0[9] ), .ZN(
        \SB2_1_19/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U3563 ( .A1(\SB2_1_3/i0[7] ), .A2(\SB2_1_3/i0_3 ), .A3(
        \SB2_1_3/i0_0 ), .ZN(\SB2_1_3/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U3564 ( .A1(\SB2_1_1/i0_3 ), .A2(\SB2_1_1/i0[9] ), .A3(
        \SB2_1_1/i0[8] ), .ZN(n1269) );
  NAND3_X1 U3565 ( .A1(n1579), .A2(\SB2_1_25/i1[9] ), .A3(\SB2_1_25/i1_5 ), 
        .ZN(n4382) );
  CLKBUF_X4 U3571 ( .I(\SB2_1_15/buf_output[1] ), .Z(\RI5[1][121] ) );
  NAND2_X1 U3572 ( .A1(\SB1_2_9/i3[0] ), .A2(\SB1_2_9/i1_7 ), .ZN(n5882) );
  INV_X1 U3579 ( .I(\MC_ARK_ARC_1_1/buf_output[163] ), .ZN(\SB1_2_4/i1_7 ) );
  CLKBUF_X4 U3581 ( .I(\MC_ARK_ARC_1_1/buf_output[70] ), .Z(\SB1_2_20/i0_4 )
         );
  NOR2_X1 U3583 ( .A1(\SB1_2_9/i1[9] ), .A2(n5882), .ZN(n5881) );
  NAND3_X1 U3587 ( .A1(\SB1_2_13/i0_0 ), .A2(\SB1_2_13/i0[7] ), .A3(
        \SB1_2_13/i0_3 ), .ZN(\SB1_2_13/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U3611 ( .A1(\SB1_2_16/i0[10] ), .A2(\SB1_2_16/i1[9] ), .A3(
        \SB1_2_16/i1_7 ), .ZN(n5622) );
  NAND3_X1 U3613 ( .A1(\SB1_2_2/i1_5 ), .A2(\SB1_2_2/i0[6] ), .A3(
        \SB1_2_2/i0[9] ), .ZN(\SB1_2_2/Component_Function_1/NAND4_in[2] ) );
  NAND2_X1 U3614 ( .A1(\SB1_2_13/i0_0 ), .A2(\SB1_2_13/i3[0] ), .ZN(
        \SB1_2_13/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U3620 ( .A1(\SB1_2_24/i1_5 ), .A2(\SB1_2_24/i1[9] ), .A3(
        \SB1_2_24/i0_4 ), .ZN(n1457) );
  NAND3_X1 U3621 ( .A1(\SB1_2_24/i0[8] ), .A2(\SB1_2_24/i3[0] ), .A3(n2913), 
        .ZN(n5957) );
  NAND3_X1 U3624 ( .A1(\SB1_2_29/i0[10] ), .A2(\SB1_2_29/i0_4 ), .A3(
        \RI1[2][17] ), .ZN(\SB1_2_29/Component_Function_0/NAND4_in[2] ) );
  NAND2_X1 U3625 ( .A1(\SB1_2_26/i0[8] ), .A2(n3192), .ZN(
        \SB1_2_26/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U3630 ( .A1(\SB1_2_27/i0_0 ), .A2(\SB1_2_27/i0_3 ), .A3(
        \SB1_2_27/i0_4 ), .ZN(\SB1_2_27/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3631 ( .A1(\SB1_2_22/i0[10] ), .A2(\SB1_2_22/i0_4 ), .A3(
        \SB1_2_22/i0_3 ), .ZN(\SB1_2_22/Component_Function_0/NAND4_in[2] ) );
  CLKBUF_X4 U3635 ( .I(\MC_ARK_ARC_1_1/buf_output[85] ), .Z(\SB1_2_17/i0[6] )
         );
  CLKBUF_X4 U3638 ( .I(\MC_ARK_ARC_1_1/buf_output[123] ), .Z(\SB1_2_11/i0[10] ) );
  NAND3_X1 U3639 ( .A1(\SB1_2_10/i0_0 ), .A2(\SB1_2_10/i0[7] ), .A3(
        \SB1_2_10/i0_3 ), .ZN(n2169) );
  NAND3_X1 U3643 ( .A1(\SB1_2_17/i0[8] ), .A2(\SB1_2_17/i1_5 ), .A3(
        \SB1_2_17/i3[0] ), .ZN(n1750) );
  NAND3_X1 U3650 ( .A1(\SB1_2_26/i0[8] ), .A2(\SB1_2_26/i0[7] ), .A3(
        \SB1_2_26/i0[6] ), .ZN(\SB1_2_26/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U3657 ( .A1(\SB1_2_3/i0[6] ), .A2(\SB1_2_3/i1_5 ), .A3(
        \SB1_2_3/i0[9] ), .ZN(n1465) );
  NAND3_X1 U3659 ( .A1(\SB1_2_27/i0_4 ), .A2(\SB1_2_27/i1[9] ), .A3(
        \SB1_2_27/i1_5 ), .ZN(n5413) );
  NAND3_X1 U3661 ( .A1(\SB1_2_15/i0[10] ), .A2(\SB1_2_15/i0_4 ), .A3(
        \SB1_2_15/i0_3 ), .ZN(\SB1_2_15/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3663 ( .A1(\SB1_2_29/i1[9] ), .A2(\RI1[2][17] ), .A3(
        \SB1_2_29/i0[6] ), .ZN(\SB1_2_29/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U3664 ( .A1(\SB1_2_12/i0[9] ), .A2(\SB1_2_12/i0_0 ), .A3(
        \SB1_2_12/i0[8] ), .ZN(\SB1_2_12/Component_Function_4/NAND4_in[0] ) );
  CLKBUF_X1 U3681 ( .I(\SB2_2_13/i0[7] ), .Z(n5779) );
  CLKBUF_X1 U3686 ( .I(\SB1_2_13/buf_output[0] ), .Z(n5880) );
  NAND3_X1 U3687 ( .A1(\SB2_2_6/i0[7] ), .A2(\SB2_2_6/i0_3 ), .A3(
        \SB2_2_6/i0_0 ), .ZN(\SB2_2_6/Component_Function_0/NAND4_in[3] ) );
  CLKBUF_X4 U3692 ( .I(\SB1_2_30/buf_output[0] ), .Z(\SB2_2_25/i0[9] ) );
  INV_X1 U3695 ( .I(\SB1_2_26/buf_output[0] ), .ZN(\SB2_2_21/i3[0] ) );
  NAND3_X1 U3697 ( .A1(n5779), .A2(\SB2_2_13/i0_3 ), .A3(\SB2_2_13/i0_0 ), 
        .ZN(\SB2_2_13/Component_Function_0/NAND4_in[3] ) );
  CLKBUF_X4 U3698 ( .I(\SB1_2_13/buf_output[4] ), .Z(\SB2_2_12/i0_4 ) );
  NAND3_X1 U3700 ( .A1(\SB2_2_6/i0[6] ), .A2(\SB2_2_6/i0_0 ), .A3(
        \SB2_2_6/i0[10] ), .ZN(n6427) );
  NAND3_X1 U3701 ( .A1(\SB2_2_31/i0[10] ), .A2(n569), .A3(\SB2_2_31/i0_3 ), 
        .ZN(\SB2_2_31/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3713 ( .A1(\SB2_2_22/i0[8] ), .A2(\SB2_2_22/i3[0] ), .A3(
        \SB2_2_22/i1_5 ), .ZN(n1820) );
  NAND3_X1 U3715 ( .A1(\SB2_2_19/i0[6] ), .A2(\SB2_2_19/i1_5 ), .A3(
        \SB2_2_19/i0[9] ), .ZN(n3701) );
  CLKBUF_X4 U3717 ( .I(\SB1_2_15/buf_output[2] ), .Z(\SB2_2_12/i0_0 ) );
  NAND3_X1 U3718 ( .A1(\SB2_2_18/i0[6] ), .A2(\SB2_2_18/i0_3 ), .A3(
        \SB2_2_18/i0[10] ), .ZN(n5010) );
  NAND3_X1 U3721 ( .A1(\SB2_2_21/i0_0 ), .A2(\SB2_2_21/i3[0] ), .A3(
        \SB2_2_21/i1_7 ), .ZN(n6444) );
  NAND3_X1 U3725 ( .A1(\SB2_2_3/i0_3 ), .A2(\SB2_2_3/i0_0 ), .A3(n5886), .ZN(
        n4494) );
  CLKBUF_X4 U3727 ( .I(\SB1_2_27/buf_output[4] ), .Z(\SB2_2_26/i0_4 ) );
  NAND3_X1 U3729 ( .A1(\SB2_2_12/i0[10] ), .A2(\SB2_2_12/i0_3 ), .A3(
        \SB2_2_12/i0[9] ), .ZN(n6517) );
  NAND2_X1 U3732 ( .A1(\SB2_2_10/i0_3 ), .A2(n5029), .ZN(n5985) );
  NAND3_X1 U3733 ( .A1(\SB2_2_10/i1_7 ), .A2(\SB2_2_10/i0[8] ), .A3(n581), 
        .ZN(n5245) );
  NAND3_X1 U3738 ( .A1(\SB2_2_15/i3[0] ), .A2(\SB2_2_15/i0[8] ), .A3(
        \SB2_2_15/i1_5 ), .ZN(n1748) );
  INV_X1 U3740 ( .I(n6), .ZN(n495) );
  NAND3_X1 U3743 ( .A1(\SB1_3_12/i0_4 ), .A2(\SB1_3_12/i1[9] ), .A3(
        \SB1_3_12/i1_5 ), .ZN(n6067) );
  INV_X1 U3746 ( .I(\MC_ARK_ARC_1_2/buf_output[55] ), .ZN(\SB1_3_22/i1_7 ) );
  INV_X1 U3749 ( .I(n6540), .ZN(\SB1_3_29/i1_5 ) );
  BUF_X2 U3750 ( .I(\MC_ARK_ARC_1_2/buf_output[187] ), .Z(\SB1_3_0/i0[6] ) );
  INV_X1 U3755 ( .I(\MC_ARK_ARC_1_2/buf_output[96] ), .ZN(\SB1_3_15/i3[0] ) );
  NAND3_X1 U3756 ( .A1(\SB1_3_1/i0[10] ), .A2(\SB1_3_1/i0_3 ), .A3(
        \SB1_3_1/i0[9] ), .ZN(n3984) );
  NAND2_X1 U3757 ( .A1(\SB1_3_10/i0_3 ), .A2(\SB1_3_10/i1[9] ), .ZN(
        \SB1_3_10/Component_Function_1/NAND4_in[0] ) );
  CLKBUF_X4 U3759 ( .I(n5501), .Z(\SB1_3_9/i0[10] ) );
  NAND2_X1 U3762 ( .A1(\SB1_3_26/i0_0 ), .A2(\SB1_3_26/i3[0] ), .ZN(
        \SB1_3_26/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U3766 ( .A1(\SB1_3_21/i0_0 ), .A2(\SB1_3_21/i0[8] ), .A3(
        \SB1_3_21/i0[9] ), .ZN(n1967) );
  CLKBUF_X4 U3769 ( .I(\MC_ARK_ARC_1_2/buf_output[49] ), .Z(\SB1_3_23/i0[6] )
         );
  NAND3_X1 U3772 ( .A1(\SB1_3_27/i0_0 ), .A2(\SB1_3_27/i0_3 ), .A3(
        \SB1_3_27/i0_4 ), .ZN(\SB1_3_27/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3773 ( .A1(\SB1_3_1/i1_7 ), .A2(\SB1_3_1/i0[8] ), .A3(
        \SB1_3_1/i0_4 ), .ZN(\SB1_3_1/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U3775 ( .A1(\SB1_3_0/i0_3 ), .A2(\SB1_3_0/i0[8] ), .A3(
        \SB1_3_0/i0[9] ), .ZN(\SB1_3_0/Component_Function_2/NAND4_in[2] ) );
  NAND2_X1 U3776 ( .A1(\SB1_3_23/i0_0 ), .A2(\SB1_3_23/i3[0] ), .ZN(
        \SB1_3_23/Component_Function_5/NAND4_in[0] ) );
  NAND2_X1 U3782 ( .A1(\SB1_3_21/i0_3 ), .A2(\SB1_3_21/i1[9] ), .ZN(
        \SB1_3_21/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U3785 ( .A1(\SB1_3_5/i1_7 ), .A2(\SB1_3_5/i0[8] ), .A3(
        \SB1_3_5/i0_4 ), .ZN(\SB1_3_5/Component_Function_1/NAND4_in[3] ) );
  CLKBUF_X4 U3787 ( .I(\MC_ARK_ARC_1_2/buf_output[117] ), .Z(\SB1_3_12/i0[10] ) );
  NAND3_X1 U3788 ( .A1(\SB1_3_19/i0_3 ), .A2(\SB1_3_19/i0[8] ), .A3(
        \SB1_3_19/i0[9] ), .ZN(\SB1_3_19/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U3793 ( .A1(\SB1_3_23/i0_0 ), .A2(\SB1_3_23/i3[0] ), .A3(
        \SB1_3_23/i1_7 ), .ZN(n3452) );
  NAND3_X1 U3804 ( .A1(\SB1_3_4/i0[9] ), .A2(\SB1_3_4/i0_0 ), .A3(
        \SB1_3_4/i0[8] ), .ZN(\SB1_3_4/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U3809 ( .A1(\SB1_3_4/i0[10] ), .A2(\SB1_3_4/i0_4 ), .A3(
        \SB1_3_4/i0_3 ), .ZN(\SB1_3_4/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3812 ( .A1(\SB1_3_30/i0_0 ), .A2(\SB1_3_30/i0[7] ), .A3(
        \SB1_3_30/i0_3 ), .ZN(\SB1_3_30/Component_Function_0/NAND4_in[3] ) );
  CLKBUF_X4 U3813 ( .I(\MC_ARK_ARC_1_2/buf_output[162] ), .Z(\SB1_3_4/i0[9] )
         );
  NAND3_X1 U3815 ( .A1(\SB1_3_6/i0[9] ), .A2(\SB1_3_6/i0[10] ), .A3(
        \SB1_3_6/i0_3 ), .ZN(\SB1_3_6/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U3816 ( .A1(\SB1_3_13/i0[10] ), .A2(\SB1_3_13/i0_3 ), .A3(
        \SB1_3_13/i0[9] ), .ZN(n4035) );
  NAND3_X1 U3818 ( .A1(\SB2_3_1/i1_5 ), .A2(\SB2_3_1/i0[10] ), .A3(
        \SB2_3_1/i1[9] ), .ZN(\SB2_3_1/Component_Function_2/NAND4_in[0] ) );
  CLKBUF_X4 U3820 ( .I(\SB1_3_7/buf_output[4] ), .Z(\SB2_3_6/i0_4 ) );
  CLKBUF_X4 U3821 ( .I(\SB1_3_3/buf_output[1] ), .Z(\SB2_3_31/i0[6] ) );
  CLKBUF_X4 U3822 ( .I(\SB1_3_15/buf_output[4] ), .Z(\SB2_3_14/i0_4 ) );
  CLKBUF_X4 U3824 ( .I(\SB1_3_6/buf_output[1] ), .Z(\SB2_3_2/i0[6] ) );
  BUF_X2 U3826 ( .I(\SB1_3_30/buf_output[1] ), .Z(\SB2_3_26/i0[6] ) );
  CLKBUF_X4 U3829 ( .I(\SB1_3_26/buf_output[0] ), .Z(\SB2_3_21/i0[9] ) );
  CLKBUF_X4 U3830 ( .I(\SB1_3_11/buf_output[3] ), .Z(\SB2_3_9/i0[10] ) );
  CLKBUF_X4 U3832 ( .I(\SB1_3_9/buf_output[0] ), .Z(\SB2_3_4/i0[9] ) );
  NAND3_X1 U3834 ( .A1(\SB2_3_26/i0[9] ), .A2(\SB2_3_26/i1_5 ), .A3(
        \SB2_3_26/i0[6] ), .ZN(\SB2_3_26/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U3836 ( .A1(\SB2_3_26/i0[9] ), .A2(\SB1_3_28/buf_output[3] ), .A3(
        \SB2_3_26/i0_3 ), .ZN(n6416) );
  NAND2_X1 U3837 ( .A1(\SB2_3_29/i0[10] ), .A2(\SB2_3_29/i0[9] ), .ZN(
        \SB2_3_29/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U3839 ( .A1(\SB2_3_14/i0[9] ), .A2(\SB2_3_14/i0[6] ), .A3(
        \SB2_3_14/i1_5 ), .ZN(\SB2_3_14/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U3854 ( .A1(\SB2_3_27/i0[10] ), .A2(\SB2_3_27/i0_3 ), .A3(
        \RI3[3][24] ), .ZN(n6526) );
  NAND3_X1 U3855 ( .A1(\SB2_3_19/i0_0 ), .A2(\SB2_3_19/i0_3 ), .A3(
        \SB2_3_19/i0[7] ), .ZN(n1271) );
  NAND3_X1 U3858 ( .A1(\SB2_3_12/i0[10] ), .A2(\SB2_3_12/i0_3 ), .A3(
        \SB2_3_12/i0_4 ), .ZN(\SB2_3_12/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U3860 ( .A1(\SB2_3_31/i0[9] ), .A2(\SB2_3_31/i1_5 ), .A3(
        \SB2_3_31/i0[6] ), .ZN(n5643) );
  NAND3_X1 U3861 ( .A1(\SB2_3_10/i0_3 ), .A2(\SB2_3_10/i1_7 ), .A3(
        \SB2_3_10/i0[8] ), .ZN(\SB2_3_10/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U3864 ( .A1(\SB2_3_17/i0_3 ), .A2(\SB2_3_17/i0_0 ), .A3(
        \SB2_3_17/i0_4 ), .ZN(\SB2_3_17/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U3865 ( .A1(\SB2_3_2/i0[10] ), .A2(\SB2_3_2/i1[9] ), .A3(
        \SB2_3_2/i1_7 ), .ZN(\SB2_3_2/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U3867 ( .A1(\SB2_3_1/i0_3 ), .A2(\SB2_3_1/i0[10] ), .A3(
        \SB2_3_1/i0[9] ), .ZN(\SB2_3_1/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U3873 ( .A1(\SB2_3_15/i0[10] ), .A2(\SB2_3_15/i1[9] ), .A3(
        \SB2_3_15/i1_7 ), .ZN(n1951) );
  NAND2_X1 U3875 ( .A1(\SB2_3_22/i0[10] ), .A2(\SB2_3_22/i0[9] ), .ZN(
        \SB2_3_22/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U3879 ( .A1(\SB2_3_10/i0_3 ), .A2(\SB2_3_10/i0[10] ), .A3(
        \SB2_3_10/i0[9] ), .ZN(n1872) );
  NAND2_X1 U3880 ( .A1(\SB2_3_17/i0_0 ), .A2(\SB2_3_17/i3[0] ), .ZN(
        \SB2_3_17/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U3884 ( .A1(\SB2_3_11/i0[9] ), .A2(\SB2_3_11/i0_3 ), .A3(
        \SB2_3_11/i0[8] ), .ZN(n5809) );
  NAND3_X1 U3885 ( .A1(\SB2_3_13/i1_7 ), .A2(\SB2_3_13/i0[8] ), .A3(
        \SB1_3_14/buf_output[4] ), .ZN(
        \SB2_3_13/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U3887 ( .A1(\SB2_3_17/i0_3 ), .A2(\SB2_3_17/i0[10] ), .A3(
        \SB2_3_17/i0[9] ), .ZN(n4021) );
  NAND3_X1 U3888 ( .A1(\SB2_3_27/i1_5 ), .A2(\SB2_3_27/i0[8] ), .A3(
        \SB2_3_27/i3[0] ), .ZN(\SB2_3_27/Component_Function_3/NAND4_in[3] ) );
  INV_X1 U3889 ( .I(n14), .ZN(n488) );
  NAND3_X1 U3890 ( .A1(\SB2_3_19/i0_0 ), .A2(\SB2_3_19/i1_5 ), .A3(
        \SB2_3_19/i0_4 ), .ZN(n6489) );
  CLKBUF_X4 U3891 ( .I(\SB2_3_19/buf_output[2] ), .Z(\RI5[3][92] ) );
  CLKBUF_X4 U3893 ( .I(\SB2_3_19/buf_output[1] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[97] ) );
  INV_X1 U3896 ( .I(n3), .ZN(n544) );
  INV_X1 U3897 ( .I(\RI1[4][179] ), .ZN(\SB3_2/i1_5 ) );
  BUF_X2 U3901 ( .I(\MC_ARK_ARC_1_3/buf_output[90] ), .Z(\SB3_16/i0[9] ) );
  CLKBUF_X2 U3904 ( .I(\MC_ARK_ARC_1_3/buf_output[132] ), .Z(\SB3_9/i0[9] ) );
  CLKBUF_X4 U3905 ( .I(\MC_ARK_ARC_1_3/buf_output[174] ), .Z(\SB3_2/i0[9] ) );
  CLKBUF_X4 U3907 ( .I(\MC_ARK_ARC_1_3/buf_output[84] ), .Z(\SB3_17/i0[9] ) );
  NAND3_X1 U3911 ( .A1(\SB3_6/i0[7] ), .A2(\SB3_6/i0_0 ), .A3(\RI1[4][155] ), 
        .ZN(n5618) );
  CLKBUF_X4 U3912 ( .I(\MC_ARK_ARC_1_3/buf_output[173] ), .Z(\SB3_3/i0_3 ) );
  NAND3_X1 U3916 ( .A1(\SB3_20/i1_7 ), .A2(\SB3_20/i0[8] ), .A3(\SB3_20/i0_4 ), 
        .ZN(\SB3_20/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U3918 ( .A1(\SB3_15/i0_0 ), .A2(\SB3_15/i1_5 ), .A3(\SB3_15/i0_4 ), 
        .ZN(\SB3_15/Component_Function_2/NAND4_in[3] ) );
  CLKBUF_X4 U3919 ( .I(\MC_ARK_ARC_1_3/buf_output[184] ), .Z(\SB3_1/i0_4 ) );
  NAND3_X1 U3925 ( .A1(\SB3_22/i1[9] ), .A2(\SB3_22/i1_7 ), .A3(
        \SB3_22/i0[10] ), .ZN(\SB3_22/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U3927 ( .A1(\SB3_17/i0_0 ), .A2(\SB3_17/i0_3 ), .A3(\SB3_17/i0_4 ), 
        .ZN(n3960) );
  NAND3_X1 U3929 ( .A1(\SB3_25/i0_3 ), .A2(\SB3_25/i1[9] ), .A3(\SB3_25/i0_4 ), 
        .ZN(n2850) );
  NAND3_X1 U3930 ( .A1(\SB3_1/i0_0 ), .A2(\SB3_1/i0_3 ), .A3(\SB3_1/i0[7] ), 
        .ZN(n3295) );
  NAND3_X1 U3941 ( .A1(\SB3_11/i0[10] ), .A2(\SB3_11/i1[9] ), .A3(
        \SB3_11/i1_7 ), .ZN(n6530) );
  NAND3_X1 U3942 ( .A1(\SB3_10/i0[8] ), .A2(\SB3_10/i3[0] ), .A3(\SB3_10/i1_5 ), .ZN(n2879) );
  NAND3_X1 U3944 ( .A1(\SB3_12/i1_7 ), .A2(\SB3_12/i0[8] ), .A3(\SB3_12/i0_4 ), 
        .ZN(\SB3_12/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U3945 ( .A1(\SB3_14/i0_3 ), .A2(\SB3_14/i1[9] ), .A3(\SB3_14/i0_4 ), 
        .ZN(n1875) );
  NAND3_X1 U3946 ( .A1(\SB3_17/i0[6] ), .A2(\SB3_17/i0[8] ), .A3(
        \SB3_17/i0[7] ), .ZN(\SB3_17/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U3947 ( .A1(\SB3_12/i0_4 ), .A2(\SB3_12/i1[9] ), .A3(\SB3_12/i1_5 ), 
        .ZN(n2720) );
  CLKBUF_X4 U3948 ( .I(\SB3_1/buf_output[5] ), .Z(\SB4_1/i0_3 ) );
  CLKBUF_X4 U3949 ( .I(\SB3_0/buf_output[4] ), .Z(\SB4_31/i0_4 ) );
  CLKBUF_X4 U3953 ( .I(\SB3_27/buf_output[1] ), .Z(\SB4_23/i0[6] ) );
  CLKBUF_X4 U3954 ( .I(\SB3_29/buf_output[4] ), .Z(\SB4_28/i0_4 ) );
  NAND3_X1 U3957 ( .A1(\SB4_26/i1_5 ), .A2(\SB4_26/i0_0 ), .A3(\SB4_26/i0_4 ), 
        .ZN(\SB4_26/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U3958 ( .A1(\SB4_1/i0_3 ), .A2(\SB4_1/i0[9] ), .A3(\SB4_1/i0[10] ), 
        .ZN(n6377) );
  NAND3_X1 U3959 ( .A1(\SB4_1/i0[9] ), .A2(\SB4_1/i0_3 ), .A3(\SB4_1/i0[8] ), 
        .ZN(n5160) );
  NAND3_X1 U3960 ( .A1(\SB4_16/i0[6] ), .A2(\SB4_16/i0[9] ), .A3(\SB4_16/i1_5 ), .ZN(\SB4_16/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U3962 ( .A1(\SB4_4/i0_4 ), .A2(\SB4_4/i0_3 ), .A3(
        \SB3_7/buf_output[2] ), .ZN(n5459) );
  NAND3_X1 U3964 ( .A1(\SB4_22/i0_3 ), .A2(\SB4_22/i0[9] ), .A3(\SB4_22/i0[8] ), .ZN(n6260) );
  NAND2_X1 U3965 ( .A1(\SB4_30/i0[10] ), .A2(\SB4_30/i0[9] ), .ZN(n4384) );
  NAND2_X1 U3972 ( .A1(\SB4_14/i0[9] ), .A2(\SB4_14/i0[10] ), .ZN(n784) );
  NAND3_X1 U3973 ( .A1(\SB4_13/i0_3 ), .A2(\SB4_13/i0_0 ), .A3(\SB4_13/i0_4 ), 
        .ZN(n6394) );
  NAND3_X1 U3978 ( .A1(\SB4_13/i0[9] ), .A2(\SB4_13/i0[6] ), .A3(\SB4_13/i0_4 ), .ZN(\SB4_13/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U3979 ( .A1(\SB4_16/i0[10] ), .A2(\SB4_16/i1[9] ), .A3(
        \SB4_16/i1_7 ), .ZN(\SB4_16/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U3980 ( .A1(\SB4_13/i0_0 ), .A2(\SB4_13/i0_4 ), .A3(\SB4_13/i1_5 ), 
        .ZN(n6365) );
  NAND3_X1 U3984 ( .A1(\SB4_26/i0_3 ), .A2(\SB4_26/i0[10] ), .A3(\SB4_26/i0_4 ), .ZN(n5357) );
  NAND3_X1 U3986 ( .A1(\SB4_28/i0_0 ), .A2(\SB4_28/i3[0] ), .A3(\SB4_28/i1_7 ), 
        .ZN(n6044) );
  NAND3_X1 U3989 ( .A1(\SB4_8/i0_3 ), .A2(\SB4_8/i0[10] ), .A3(\SB4_8/i0[9] ), 
        .ZN(n629) );
  NAND3_X1 U3992 ( .A1(\SB4_22/i0_4 ), .A2(\SB4_22/i0[9] ), .A3(\SB4_22/i0[6] ), .ZN(n5471) );
  NAND2_X1 U3993 ( .A1(\SB4_22/i0_3 ), .A2(\SB4_22/i1[9] ), .ZN(
        \SB4_22/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U3994 ( .A1(\SB4_9/i0_0 ), .A2(\SB4_9/i0_4 ), .A3(\SB4_9/i0_3 ), 
        .ZN(n6130) );
  AND2_X1 U3999 ( .A1(n6458), .A2(\SB1_2_9/Component_Function_4/NAND4_in[3] ), 
        .Z(n4755) );
  XNOR2_X1 U4005 ( .A1(\SB2_0_9/buf_output[5] ), .A2(n64), .ZN(n4756) );
  AND2_X1 U4007 ( .A1(n1956), .A2(\SB1_1_16/Component_Function_4/NAND4_in[3] ), 
        .Z(n4757) );
  AND2_X1 U4008 ( .A1(\SB1_1_16/i0[8] ), .A2(\SB1_1_16/i0[9] ), .Z(n4758) );
  AND2_X1 U4010 ( .A1(\SB2_1_9/i1_7 ), .A2(\SB2_1_9/i0[8] ), .Z(n4759) );
  AND2_X2 U4011 ( .A1(\SB2_1_9/Component_Function_3/NAND4_in[2] ), .A2(n3982), 
        .Z(n4760) );
  AND2_X2 U4013 ( .A1(\RI3[0][103] ), .A2(\SB1_0_19/buf_output[0] ), .Z(n4761)
         );
  XNOR2_X1 U4014 ( .A1(\MC_ARK_ARC_1_1/temp6[81] ), .A2(n4657), .ZN(n4762) );
  AND4_X2 U4018 ( .A1(\SB1_3_17/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_17/Component_Function_5/NAND4_in[3] ), .A3(n3976), .A4(
        \SB1_3_17/Component_Function_5/NAND4_in[0] ), .Z(n4763) );
  XNOR2_X1 U4019 ( .A1(n5811), .A2(n2461), .ZN(n4764) );
  XNOR2_X1 U4022 ( .A1(\MC_ARK_ARC_1_3/temp5[182] ), .A2(n2610), .ZN(n4765) );
  XNOR2_X1 U4023 ( .A1(\MC_ARK_ARC_1_3/temp5[149] ), .A2(
        \MC_ARK_ARC_1_3/temp6[149] ), .ZN(n4766) );
  XNOR2_X1 U4025 ( .A1(\SB2_3_13/buf_output[5] ), .A2(\SB2_3_14/buf_output[5] ), .ZN(n4767) );
  AND4_X2 U4026 ( .A1(n2598), .A2(\SB1_3_11/Component_Function_5/NAND4_in[3] ), 
        .A3(\SB1_3_11/Component_Function_5/NAND4_in[0] ), .A4(n6275), .Z(n4768) );
  AND4_X2 U4027 ( .A1(\SB1_2_18/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_18/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_2_18/Component_Function_5/NAND4_in[0] ), .A4(n2142), .Z(n4769) );
  NAND4_X2 U4028 ( .A1(\SB3_24/Component_Function_3/NAND4_in[1] ), .A2(n6529), 
        .A3(n4530), .A4(n4770), .ZN(\SB3_24/buf_output[3] ) );
  NAND3_X1 U4029 ( .A1(\SB3_24/i0[10] ), .A2(\SB3_24/i1_7 ), .A3(
        \SB3_24/i1[9] ), .ZN(n4770) );
  NAND4_X2 U4033 ( .A1(\SB2_2_12/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_12/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_2_12/Component_Function_3/NAND4_in[3] ), .A4(
        \SB2_2_12/Component_Function_3/NAND4_in[1] ), .ZN(
        \SB2_2_12/buf_output[3] ) );
  NAND4_X2 U4034 ( .A1(\SB2_2_15/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_15/Component_Function_3/NAND4_in[2] ), .A3(n1748), .A4(n4771), 
        .ZN(\SB2_2_15/buf_output[3] ) );
  XOR2_X1 U4035 ( .A1(n4772), .A2(n97), .Z(Ciphertext[189]) );
  NAND4_X2 U4036 ( .A1(\SB4_0/Component_Function_3/NAND4_in[3] ), .A2(n1322), 
        .A3(\SB4_0/Component_Function_3/NAND4_in[1] ), .A4(n5454), .ZN(n4772)
         );
  XOR2_X1 U4038 ( .A1(n4774), .A2(n4773), .Z(\MC_ARK_ARC_1_3/temp5[167] ) );
  XOR2_X1 U4040 ( .A1(\RI5[3][137] ), .A2(n1365), .Z(n4773) );
  XOR2_X1 U4047 ( .A1(\RI5[3][113] ), .A2(\RI5[3][161] ), .Z(n4774) );
  XOR2_X1 U4048 ( .A1(\MC_ARK_ARC_1_2/temp5[86] ), .A2(
        \MC_ARK_ARC_1_2/temp6[86] ), .Z(\MC_ARK_ARC_1_2/buf_output[86] ) );
  XOR2_X1 U4050 ( .A1(\MC_ARK_ARC_1_2/temp2[86] ), .A2(n5706), .Z(
        \MC_ARK_ARC_1_2/temp5[86] ) );
  INV_X2 U4052 ( .I(\SB1_2_17/buf_output[2] ), .ZN(\SB2_2_14/i1[9] ) );
  NAND4_X2 U4058 ( .A1(\SB1_2_17/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_17/Component_Function_2/NAND4_in[3] ), .A3(n1452), .A4(
        \SB1_2_17/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB1_2_17/buf_output[2] ) );
  NAND4_X2 U4059 ( .A1(n5010), .A2(\SB2_2_18/Component_Function_2/NAND4_in[0] ), .A3(\SB2_2_18/Component_Function_2/NAND4_in[2] ), .A4(n3616), .ZN(
        \SB2_2_18/buf_output[2] ) );
  XOR2_X1 U4060 ( .A1(n4775), .A2(n244), .Z(Ciphertext[118]) );
  NAND4_X2 U4061 ( .A1(n5535), .A2(\SB4_12/Component_Function_4/NAND4_in[0] ), 
        .A3(\SB4_12/Component_Function_4/NAND4_in[3] ), .A4(n4476), .ZN(n4775)
         );
  INV_X1 U4062 ( .I(\SB1_3_3/buf_output[1] ), .ZN(\SB2_3_31/i1_7 ) );
  NAND4_X2 U4063 ( .A1(\SB1_3_3/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_3_3/Component_Function_1/NAND4_in[2] ), .A3(n5075), .A4(n1684), 
        .ZN(\SB1_3_3/buf_output[1] ) );
  NAND3_X2 U4064 ( .A1(\SB1_3_8/i0_3 ), .A2(\SB1_3_8/i0[8] ), .A3(
        \SB1_3_8/i1_7 ), .ZN(\SB1_3_8/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 U4065 ( .A1(n2646), .A2(\SB1_3_26/Component_Function_4/NAND4_in[3] ), .ZN(n4862) );
  NAND4_X2 U4066 ( .A1(\SB1_3_7/Component_Function_5/NAND4_in[1] ), .A2(n6498), 
        .A3(\SB1_3_7/Component_Function_5/NAND4_in[0] ), .A4(n4776), .ZN(
        \SB1_3_7/buf_output[5] ) );
  NAND3_X2 U4068 ( .A1(\SB1_3_7/i1[9] ), .A2(\SB1_3_7/i0_4 ), .A3(
        \SB1_3_7/i0_3 ), .ZN(n4776) );
  NAND4_X2 U4069 ( .A1(\SB1_1_17/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_17/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_17/Component_Function_3/NAND4_in[3] ), .A4(
        \SB1_1_17/Component_Function_3/NAND4_in[2] ), .ZN(
        \SB1_1_17/buf_output[3] ) );
  XOR2_X1 U4070 ( .A1(n4778), .A2(n4777), .Z(\MC_ARK_ARC_1_1/temp6[29] ) );
  XOR2_X1 U4072 ( .A1(\RI5[1][131] ), .A2(n488), .Z(n4777) );
  XOR2_X1 U4073 ( .A1(\RI5[1][65] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[95] ), 
        .Z(n4778) );
  NAND4_X2 U4074 ( .A1(\SB1_3_21/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_3_21/Component_Function_2/NAND4_in[1] ), .A3(n5761), .A4(n4840), 
        .ZN(\SB1_3_21/buf_output[2] ) );
  NAND4_X2 U4077 ( .A1(\SB1_3_18/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_3_18/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_3_18/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_3_18/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB1_3_18/buf_output[4] ) );
  NAND4_X2 U4080 ( .A1(\SB1_0_12/Component_Function_2/NAND4_in[0] ), .A2(n1978), .A3(n5338), .A4(\SB1_0_12/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB1_0_12/buf_output[2] ) );
  XOR2_X1 U4085 ( .A1(n4779), .A2(n126), .Z(Ciphertext[55]) );
  NAND4_X2 U4086 ( .A1(n6261), .A2(\SB4_22/Component_Function_1/NAND4_in[3] ), 
        .A3(\SB4_22/Component_Function_1/NAND4_in[1] ), .A4(
        \SB4_22/Component_Function_1/NAND4_in[0] ), .ZN(n4779) );
  NAND4_X2 U4087 ( .A1(n5146), .A2(n5784), .A3(n5285), .A4(n4626), .ZN(
        \SB2_2_11/buf_output[2] ) );
  XOR2_X1 U4091 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[155] ), .A2(\RI5[3][131] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[185] ) );
  XOR2_X1 U4095 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[155] ), .A2(\RI5[3][161] ), 
        .Z(n2281) );
  NAND4_X2 U4096 ( .A1(\SB2_1_6/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_1_6/Component_Function_2/NAND4_in[0] ), .A3(n5476), .A4(n5803), 
        .ZN(\SB2_1_6/buf_output[2] ) );
  NAND4_X2 U4099 ( .A1(\SB1_1_17/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_1_17/Component_Function_4/NAND4_in[2] ), .A3(n5059), .A4(
        \SB1_1_17/Component_Function_4/NAND4_in[0] ), .ZN(
        \SB1_1_17/buf_output[4] ) );
  NAND3_X2 U4100 ( .A1(\SB1_3_15/i0_0 ), .A2(\SB1_3_15/i0[10] ), .A3(
        \SB1_3_15/i0[6] ), .ZN(\SB1_3_15/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U4101 ( .A1(\SB1_3_8/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_3_8/Component_Function_3/NAND4_in[0] ), .A3(n4296), .A4(
        \SB1_3_8/Component_Function_3/NAND4_in[2] ), .ZN(
        \SB1_3_8/buf_output[3] ) );
  NAND3_X2 U4106 ( .A1(\SB2_3_6/i0[10] ), .A2(\SB2_3_6/i0_0 ), .A3(
        \SB2_3_6/i0[6] ), .ZN(n5345) );
  NAND4_X2 U4107 ( .A1(\SB2_2_16/Component_Function_5/NAND4_in[2] ), .A2(n4022), .A3(n3041), .A4(n6488), .ZN(\SB2_2_16/buf_output[5] ) );
  NAND4_X2 U4108 ( .A1(\SB2_2_27/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_27/Component_Function_2/NAND4_in[2] ), .A3(n3198), .A4(n4455), 
        .ZN(\SB2_2_27/buf_output[2] ) );
  NAND4_X2 U4110 ( .A1(\SB2_0_23/Component_Function_5/NAND4_in[2] ), .A2(n950), 
        .A3(n5849), .A4(\SB2_0_23/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_0_23/buf_output[5] ) );
  NAND4_X2 U4113 ( .A1(\SB2_2_5/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_5/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_2_5/Component_Function_2/NAND4_in[1] ), .A4(n1881), .ZN(
        \SB2_2_5/buf_output[2] ) );
  NAND3_X2 U4114 ( .A1(\SB2_2_6/i0[10] ), .A2(\SB2_2_6/i1_7 ), .A3(
        \SB2_2_6/i1[9] ), .ZN(\SB2_2_6/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U4116 ( .A1(\SB1_2_27/i0_3 ), .A2(\SB1_2_27/i0_4 ), .A3(
        \SB1_2_27/i1[9] ), .ZN(n5110) );
  NAND4_X2 U4118 ( .A1(\SB1_3_21/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_3_21/Component_Function_1/NAND4_in[2] ), .A3(n5708), .A4(
        \SB1_3_21/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_3_21/buf_output[1] ) );
  XOR2_X1 U4119 ( .A1(\RI5[0][32] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[56] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[86] ) );
  NAND4_X2 U4123 ( .A1(\SB1_2_11/Component_Function_3/NAND4_in[2] ), .A2(
        \SB1_2_11/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_2_11/Component_Function_3/NAND4_in[1] ), .A4(
        \SB1_2_11/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_2_11/buf_output[3] ) );
  NAND3_X1 U4126 ( .A1(\SB3_5/i0_4 ), .A2(\SB3_5/i0_3 ), .A3(\SB3_5/i0[10] ), 
        .ZN(\SB3_5/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U4127 ( .A1(\SB1_3_12/i0_4 ), .A2(\SB1_3_12/i1_7 ), .A3(
        \SB1_3_12/i0[8] ), .ZN(\SB1_3_12/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U4131 ( .A1(\SB2_1_3/Component_Function_1/NAND4_in[1] ), .A2(n4802), 
        .A3(\SB2_1_3/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_1_3/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_1_3/buf_output[1] ) );
  NAND4_X2 U4134 ( .A1(\SB1_2_26/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_26/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_2_26/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_2_26/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_2_26/buf_output[0] ) );
  NAND4_X2 U4143 ( .A1(\SB1_2_16/Component_Function_5/NAND4_in[1] ), .A2(n715), 
        .A3(\SB1_2_16/Component_Function_5/NAND4_in[0] ), .A4(
        \SB1_2_16/Component_Function_5/NAND4_in[2] ), .ZN(
        \SB1_2_16/buf_output[5] ) );
  XOR2_X1 U4148 ( .A1(n4781), .A2(n4780), .Z(\MC_ARK_ARC_1_0/temp6[38] ) );
  XOR2_X1 U4149 ( .A1(\RI5[0][104] ), .A2(n89), .Z(n4780) );
  XOR2_X1 U4150 ( .A1(\RI5[0][140] ), .A2(\RI5[0][74] ), .Z(n4781) );
  NAND4_X2 U4152 ( .A1(\SB1_3_3/Component_Function_3/NAND4_in[1] ), .A2(n1546), 
        .A3(n5154), .A4(n4782), .ZN(\SB1_3_3/buf_output[3] ) );
  NAND4_X2 U4154 ( .A1(n1849), .A2(n3118), .A3(
        \SB1_2_15/Component_Function_5/NAND4_in[0] ), .A4(n4783), .ZN(
        \SB1_2_15/buf_output[5] ) );
  NAND3_X2 U4155 ( .A1(\SB1_2_15/i0[6] ), .A2(\SB1_2_15/i0_0 ), .A3(
        \SB1_2_15/i0[10] ), .ZN(n4783) );
  XOR2_X1 U4159 ( .A1(\MC_ARK_ARC_1_2/temp4[35] ), .A2(n4784), .Z(n5276) );
  XOR2_X1 U4160 ( .A1(\RI5[2][101] ), .A2(\RI5[2][137] ), .Z(n4784) );
  NAND4_X2 U4166 ( .A1(\SB4_29/Component_Function_4/NAND4_in[3] ), .A2(
        \SB4_29/Component_Function_4/NAND4_in[1] ), .A3(
        \SB4_29/Component_Function_4/NAND4_in[0] ), .A4(n4785), .ZN(n5615) );
  NAND3_X2 U4167 ( .A1(\SB4_29/i0[10] ), .A2(\SB4_29/i0_3 ), .A3(
        \SB4_29/i0[9] ), .ZN(n4785) );
  NAND4_X2 U4170 ( .A1(n2050), .A2(\SB2_3_26/Component_Function_5/NAND4_in[3] ), .A3(n4971), .A4(\SB2_3_26/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_3_26/buf_output[5] ) );
  XOR2_X1 U4171 ( .A1(\MC_ARK_ARC_1_1/temp2[97] ), .A2(n4786), .Z(
        \MC_ARK_ARC_1_1/temp5[97] ) );
  XOR2_X1 U4174 ( .A1(\RI5[1][97] ), .A2(\RI5[1][91] ), .Z(n4786) );
  XOR2_X1 U4175 ( .A1(n4788), .A2(n4787), .Z(\MC_ARK_ARC_1_2/temp5[125] ) );
  XOR2_X1 U4177 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[95] ), .A2(\RI5[2][119] ), 
        .Z(n4787) );
  XOR2_X1 U4181 ( .A1(\RI5[2][71] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[125] ), 
        .Z(n4788) );
  XOR2_X1 U4182 ( .A1(n4790), .A2(n4789), .Z(\MC_ARK_ARC_1_0/buf_output[20] )
         );
  XOR2_X1 U4189 ( .A1(\MC_ARK_ARC_1_0/temp4[20] ), .A2(
        \MC_ARK_ARC_1_0/temp2[20] ), .Z(n4789) );
  XOR2_X1 U4190 ( .A1(\MC_ARK_ARC_1_0/temp3[20] ), .A2(
        \MC_ARK_ARC_1_0/temp1[20] ), .Z(n4790) );
  XOR2_X1 U4191 ( .A1(n4791), .A2(n158), .Z(Ciphertext[33]) );
  NAND4_X2 U4193 ( .A1(n2419), .A2(\SB4_26/Component_Function_3/NAND4_in[3] ), 
        .A3(n2103), .A4(\SB4_26/Component_Function_3/NAND4_in[1] ), .ZN(n4791)
         );
  NAND4_X2 U4196 ( .A1(\SB1_2_29/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_2_29/Component_Function_2/NAND4_in[0] ), .A3(n3575), .A4(n5330), 
        .ZN(\SB1_2_29/buf_output[2] ) );
  BUF_X4 U4198 ( .I(\SB2_3_21/buf_output[2] ), .Z(\RI5[3][80] ) );
  NAND4_X2 U4199 ( .A1(\SB2_1_11/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_11/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_1_11/Component_Function_4/NAND4_in[1] ), .A4(n4792), .ZN(
        \SB2_1_11/buf_output[4] ) );
  NAND3_X2 U4201 ( .A1(\SB2_1_11/i0[9] ), .A2(\SB2_1_11/i0_3 ), .A3(
        \SB2_1_11/i0[10] ), .ZN(n4792) );
  BUF_X2 U4202 ( .I(\SB3_11/buf_output[3] ), .Z(\SB4_9/i0[10] ) );
  NAND4_X2 U4204 ( .A1(n2387), .A2(\SB2_3_30/Component_Function_5/NAND4_in[1] ), .A3(n4803), .A4(n1735), .ZN(\SB2_3_30/buf_output[5] ) );
  XOR2_X1 U4205 ( .A1(\MC_ARK_ARC_1_2/temp1[20] ), .A2(n4793), .Z(
        \MC_ARK_ARC_1_2/temp5[20] ) );
  XOR2_X1 U4208 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[158] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[182] ), .Z(n4793) );
  XOR2_X1 U4211 ( .A1(\MC_ARK_ARC_1_3/temp5[178] ), .A2(n4794), .Z(
        \MC_ARK_ARC_1_3/buf_output[178] ) );
  XOR2_X1 U4217 ( .A1(\MC_ARK_ARC_1_3/temp4[178] ), .A2(
        \MC_ARK_ARC_1_3/temp3[178] ), .Z(n4794) );
  XOR2_X1 U4218 ( .A1(n4795), .A2(n86), .Z(Ciphertext[32]) );
  NAND4_X2 U4219 ( .A1(\SB4_26/Component_Function_2/NAND4_in[1] ), .A2(
        \SB4_26/Component_Function_2/NAND4_in[0] ), .A3(
        \SB4_26/Component_Function_2/NAND4_in[3] ), .A4(n6421), .ZN(n4795) );
  NAND4_X2 U4223 ( .A1(\SB2_3_3/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_3_3/Component_Function_2/NAND4_in[3] ), .A3(n5634), .A4(
        \SB2_3_3/Component_Function_2/NAND4_in[1] ), .ZN(
        \SB2_3_3/buf_output[2] ) );
  NAND4_X2 U4224 ( .A1(\SB2_2_21/Component_Function_0/NAND4_in[1] ), .A2(n1086), .A3(\SB2_2_21/Component_Function_0/NAND4_in[2] ), .A4(n4796), .ZN(
        \SB2_2_21/buf_output[0] ) );
  NAND2_X1 U4225 ( .A1(\SB2_2_21/i0[10] ), .A2(\SB2_2_21/i0[9] ), .ZN(n4796)
         );
  NAND4_X2 U4226 ( .A1(\SB2_1_24/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_1_24/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_1_24/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_24/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_1_24/buf_output[1] ) );
  INV_X2 U4229 ( .I(\SB1_1_25/buf_output[2] ), .ZN(\SB2_1_22/i1[9] ) );
  NAND4_X2 U4230 ( .A1(n2865), .A2(\SB1_1_25/Component_Function_2/NAND4_in[1] ), .A3(\SB1_1_25/Component_Function_2/NAND4_in[0] ), .A4(
        \SB1_1_25/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB1_1_25/buf_output[2] ) );
  XOR2_X1 U4234 ( .A1(\MC_ARK_ARC_1_1/temp4[34] ), .A2(n4797), .Z(n4254) );
  XOR2_X1 U4235 ( .A1(\RI5[1][136] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[100] ), 
        .Z(n4797) );
  INV_X2 U4236 ( .I(n1603), .ZN(\SB2_3_12/i3[0] ) );
  NAND2_X2 U4237 ( .A1(n6185), .A2(n6513), .ZN(n1603) );
  XOR2_X1 U4241 ( .A1(\SB2_3_19/buf_output[5] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[41] ), .Z(n5094) );
  XOR2_X1 U4247 ( .A1(\MC_ARK_ARC_1_0/temp2[124] ), .A2(n4798), .Z(
        \MC_ARK_ARC_1_0/temp5[124] ) );
  XOR2_X1 U4250 ( .A1(\RI5[0][118] ), .A2(\RI5[0][124] ), .Z(n4798) );
  XOR2_X1 U4251 ( .A1(\MC_ARK_ARC_1_2/temp2[76] ), .A2(n4799), .Z(
        \MC_ARK_ARC_1_2/temp5[76] ) );
  XOR2_X1 U4253 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[70] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[76] ), .Z(n4799) );
  NAND3_X2 U4255 ( .A1(\SB1_1_0/i0[10] ), .A2(\SB1_1_0/i0_0 ), .A3(
        \SB1_1_0/i0[6] ), .ZN(n6299) );
  NAND3_X2 U4256 ( .A1(\SB1_3_12/i0[10] ), .A2(\SB1_3_12/i1[9] ), .A3(
        \SB1_3_12/i1_5 ), .ZN(\SB1_3_12/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U4258 ( .A1(\SB1_1_8/i0_4 ), .A2(\SB1_1_8/i1[9] ), .A3(
        \RI1[1][143] ), .ZN(\SB1_1_8/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U4260 ( .A1(\SB1_2_15/i0_4 ), .A2(\SB1_2_15/i0_0 ), .A3(
        \SB1_2_15/i0_3 ), .ZN(\SB1_2_15/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U4261 ( .A1(\SB1_3_9/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_9/Component_Function_3/NAND4_in[1] ), .A3(n4939), .A4(n1926), 
        .ZN(\SB1_3_9/buf_output[3] ) );
  NAND3_X2 U4263 ( .A1(\SB2_0_4/i0[10] ), .A2(\SB2_0_4/i0_3 ), .A3(
        \SB2_0_4/i0[6] ), .ZN(\SB2_0_4/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U4269 ( .A1(\SB2_1_0/i0[10] ), .A2(\SB2_1_0/i1_5 ), .A3(
        \SB2_1_0/i1[9] ), .ZN(\SB2_1_0/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U4273 ( .A1(\SB2_1_5/Component_Function_4/NAND4_in[3] ), .A2(n6285), 
        .A3(\SB2_1_5/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_1_5/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB2_1_5/buf_output[4] ) );
  XOR2_X1 U4274 ( .A1(n4801), .A2(n4800), .Z(n4066) );
  XOR2_X1 U4275 ( .A1(\RI5[1][45] ), .A2(n455), .Z(n4800) );
  XOR2_X1 U4276 ( .A1(\RI5[1][81] ), .A2(\RI5[1][15] ), .Z(n4801) );
  NAND3_X1 U4281 ( .A1(\SB2_1_3/i0[6] ), .A2(\SB2_1_3/i1_5 ), .A3(
        \SB2_1_3/i0[9] ), .ZN(n4802) );
  NAND2_X2 U4282 ( .A1(\SB2_2_22/i0_0 ), .A2(\SB2_2_22/i3[0] ), .ZN(n6433) );
  NAND3_X1 U4283 ( .A1(\SB2_3_30/i0[9] ), .A2(\SB2_3_30/i0[6] ), .A3(
        \SB1_3_31/buf_output[4] ), .ZN(n4803) );
  AND2_X1 U4285 ( .A1(n2047), .A2(n4804), .Z(n4036) );
  NAND3_X1 U4289 ( .A1(\SB1_2_15/i0_0 ), .A2(\SB1_2_15/i1_7 ), .A3(
        \SB1_2_15/i3[0] ), .ZN(n4804) );
  XOR2_X1 U4290 ( .A1(n5574), .A2(n4805), .Z(n2621) );
  XOR2_X1 U4291 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[129] ), .A2(
        \SB2_2_20/buf_output[3] ), .Z(n4805) );
  XOR2_X1 U4292 ( .A1(\SB2_0_14/buf_output[1] ), .A2(\RI5[0][103] ), .Z(
        \MC_ARK_ARC_1_0/temp2[157] ) );
  NAND3_X1 U4295 ( .A1(\RI3[0][82] ), .A2(\SB2_0_18/i0[8] ), .A3(
        \SB2_0_18/i1_7 ), .ZN(\SB2_0_18/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U4303 ( .A1(\SB2_2_28/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_2_28/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_2_28/Component_Function_1/NAND4_in[0] ), .A4(n4806), .ZN(
        \SB2_2_28/buf_output[1] ) );
  NAND3_X1 U4305 ( .A1(\SB2_2_28/i0[9] ), .A2(\SB2_2_28/i0[6] ), .A3(
        \SB2_2_28/i1_5 ), .ZN(n4806) );
  NAND2_X2 U4307 ( .A1(n4023), .A2(n4807), .ZN(n1158) );
  NAND3_X1 U4308 ( .A1(\SB1_1_5/i0_0 ), .A2(\SB1_1_5/i1_7 ), .A3(
        \SB1_1_5/i3[0] ), .ZN(n4807) );
  NAND3_X2 U4311 ( .A1(\SB1_1_25/i0[10] ), .A2(\SB1_1_25/i1[9] ), .A3(
        \SB1_1_25/i1_7 ), .ZN(n4873) );
  BUF_X4 U4316 ( .I(n429), .Z(\SB1_0_7/i0_3 ) );
  NAND3_X1 U4317 ( .A1(\SB2_1_10/i0[6] ), .A2(\SB2_1_10/i0_3 ), .A3(
        \SB2_1_10/i1[9] ), .ZN(\SB2_1_10/Component_Function_3/NAND4_in[0] ) );
  NAND4_X2 U4318 ( .A1(\SB1_1_2/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_2/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_1_2/Component_Function_2/NAND4_in[3] ), .A4(n4105), .ZN(
        \SB1_1_2/buf_output[2] ) );
  NAND3_X1 U4319 ( .A1(\SB2_2_15/i0_3 ), .A2(\SB2_2_15/i0[8] ), .A3(
        \SB2_2_15/i1_7 ), .ZN(\SB2_2_15/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U4321 ( .A1(\MC_ARK_ARC_1_1/temp4[97] ), .A2(n4808), .Z(n6392) );
  XOR2_X1 U4325 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[163] ), .A2(\RI5[1][7] ), 
        .Z(n4808) );
  XOR2_X1 U4332 ( .A1(\RI5[0][110] ), .A2(\RI5[0][104] ), .Z(
        \MC_ARK_ARC_1_0/temp1[110] ) );
  CLKBUF_X2 U4334 ( .I(Key[96]), .Z(n79) );
  NAND3_X1 U4336 ( .A1(\SB1_3_15/i0_3 ), .A2(\SB1_3_15/i0_4 ), .A3(
        \SB1_3_15/i1[9] ), .ZN(\SB1_3_15/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U4338 ( .A1(\SB2_3_7/i0[9] ), .A2(\SB2_3_7/i0[8] ), .A3(
        \SB2_3_7/i0_3 ), .ZN(n3882) );
  NAND4_X2 U4339 ( .A1(\SB2_2_10/Component_Function_3/NAND4_in[3] ), .A2(
        \SB2_2_10/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_2_10/Component_Function_3/NAND4_in[0] ), .A4(
        \SB2_2_10/Component_Function_3/NAND4_in[2] ), .ZN(
        \SB2_2_10/buf_output[3] ) );
  NAND4_X2 U4344 ( .A1(\SB1_2_5/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_5/Component_Function_3/NAND4_in[1] ), .A3(n5452), .A4(n6353), 
        .ZN(\SB1_2_5/buf_output[3] ) );
  NAND3_X2 U4346 ( .A1(\SB1_2_12/i0_3 ), .A2(\SB1_2_12/i0[10] ), .A3(
        \SB1_2_12/i0[6] ), .ZN(n4050) );
  NAND3_X1 U4350 ( .A1(\SB3_0/i0_3 ), .A2(\SB3_0/i0_0 ), .A3(\SB3_0/i0[7] ), 
        .ZN(\SB3_0/Component_Function_0/NAND4_in[3] ) );
  NAND4_X2 U4352 ( .A1(n806), .A2(\SB1_3_0/Component_Function_5/NAND4_in[3] ), 
        .A3(\SB1_3_0/Component_Function_5/NAND4_in[0] ), .A4(n6210), .ZN(
        \SB1_3_0/buf_output[5] ) );
  NAND3_X2 U4355 ( .A1(\SB2_1_6/i0_3 ), .A2(\SB2_1_6/i0_4 ), .A3(
        \SB2_1_6/i1[9] ), .ZN(n2392) );
  NAND3_X1 U4357 ( .A1(\SB4_2/i0_0 ), .A2(\SB4_2/i0_3 ), .A3(\SB4_2/i0_4 ), 
        .ZN(\SB4_2/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U4359 ( .A1(\SB2_2_27/i0_0 ), .A2(\SB2_2_27/i0[9] ), .A3(
        \SB2_2_27/i0[8] ), .ZN(n3775) );
  NAND4_X2 U4360 ( .A1(n5266), .A2(n3926), .A3(
        \SB4_3/Component_Function_4/NAND4_in[0] ), .A4(
        \SB4_3/Component_Function_4/NAND4_in[1] ), .ZN(n4843) );
  NAND4_X2 U4365 ( .A1(n2284), .A2(\SB1_3_4/Component_Function_5/NAND4_in[2] ), 
        .A3(\SB1_3_4/Component_Function_5/NAND4_in[3] ), .A4(n2054), .ZN(
        \SB1_3_4/buf_output[5] ) );
  INV_X1 U4366 ( .I(\SB3_7/buf_output[0] ), .ZN(\SB4_2/i3[0] ) );
  NAND4_X2 U4369 ( .A1(\SB3_7/Component_Function_0/NAND4_in[3] ), .A2(
        \SB3_7/Component_Function_0/NAND4_in[0] ), .A3(
        \SB3_7/Component_Function_0/NAND4_in[1] ), .A4(n4289), .ZN(
        \SB3_7/buf_output[0] ) );
  NAND3_X1 U4373 ( .A1(\SB3_12/i0_3 ), .A2(\SB3_12/i0[8] ), .A3(\SB3_12/i1_7 ), 
        .ZN(\SB3_12/Component_Function_1/NAND4_in[1] ) );
  NAND3_X2 U4374 ( .A1(\SB2_2_10/i0[6] ), .A2(\SB2_2_10/i0[10] ), .A3(
        \SB2_2_10/i0_0 ), .ZN(\SB2_2_10/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U4375 ( .A1(\SB1_3_21/Component_Function_3/NAND4_in[0] ), .A2(n1350), .A3(n4845), .A4(n1663), .ZN(\SB1_3_21/buf_output[3] ) );
  NAND4_X2 U4376 ( .A1(\SB1_3_3/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_3/Component_Function_2/NAND4_in[0] ), .A3(n4412), .A4(
        \SB1_3_3/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB1_3_3/buf_output[2] ) );
  XOR2_X1 U4377 ( .A1(n4810), .A2(n4809), .Z(\MC_ARK_ARC_1_1/temp5[185] ) );
  XOR2_X1 U4378 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[185] ), .A2(\RI5[1][131] ), 
        .Z(n4809) );
  XOR2_X1 U4383 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[179] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[155] ), .Z(n4810) );
  NAND4_X2 U4392 ( .A1(\SB1_1_3/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_3/Component_Function_4/NAND4_in[1] ), .A3(n5206), .A4(n1643), 
        .ZN(\SB1_1_3/buf_output[4] ) );
  NAND3_X1 U4393 ( .A1(\SB1_2_1/i0[10] ), .A2(\SB1_2_1/i0_3 ), .A3(
        \SB1_2_1/i0[9] ), .ZN(\SB1_2_1/Component_Function_4/NAND4_in[2] ) );
  XOR2_X1 U4394 ( .A1(n4811), .A2(n24), .Z(Ciphertext[138]) );
  NAND4_X2 U4400 ( .A1(\SB4_8/Component_Function_0/NAND4_in[3] ), .A2(
        \SB4_8/Component_Function_0/NAND4_in[2] ), .A3(
        \SB4_8/Component_Function_0/NAND4_in[1] ), .A4(
        \SB4_8/Component_Function_0/NAND4_in[0] ), .ZN(n4811) );
  NAND3_X1 U4406 ( .A1(\SB1_3_4/i1_7 ), .A2(\MC_ARK_ARC_1_2/buf_output[166] ), 
        .A3(\SB1_3_4/i0[8] ), .ZN(\SB1_3_4/Component_Function_1/NAND4_in[3] )
         );
  NAND4_X2 U4409 ( .A1(\SB4_8/Component_Function_5/NAND4_in[2] ), .A2(
        \SB4_8/Component_Function_5/NAND4_in[1] ), .A3(
        \SB4_8/Component_Function_5/NAND4_in[0] ), .A4(n4812), .ZN(n5698) );
  NAND3_X1 U4411 ( .A1(\SB4_8/i0[6] ), .A2(\SB4_8/i0_4 ), .A3(\SB4_8/i0[9] ), 
        .ZN(n4812) );
  NAND4_X2 U4414 ( .A1(n1156), .A2(\SB4_27/Component_Function_2/NAND4_in[1] ), 
        .A3(\SB4_27/Component_Function_2/NAND4_in[0] ), .A4(n4813), .ZN(n3249)
         );
  NAND3_X1 U4415 ( .A1(\SB4_27/i0[9] ), .A2(\SB4_27/i0_3 ), .A3(\SB4_27/i0[8] ), .ZN(n4813) );
  NAND3_X1 U4417 ( .A1(\SB1_2_1/i0_3 ), .A2(\SB1_2_1/i0[8] ), .A3(
        \SB1_2_1/i1_7 ), .ZN(\SB1_2_1/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U4420 ( .A1(\SB1_1_25/i0_0 ), .A2(\SB1_1_25/i0[7] ), .A3(
        \SB1_1_25/i0_3 ), .ZN(\SB1_1_25/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U4422 ( .A1(\SB2_2_29/i0[6] ), .A2(\SB1_2_2/buf_output[0] ), .A3(
        \SB2_2_29/i1_5 ), .ZN(\SB2_2_29/Component_Function_1/NAND4_in[2] ) );
  XOR2_X1 U4423 ( .A1(n4814), .A2(\MC_ARK_ARC_1_2/temp4[92] ), .Z(n3496) );
  XOR2_X1 U4428 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[158] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[2] ), .Z(n4814) );
  BUF_X2 U4429 ( .I(\SB3_27/buf_output[3] ), .Z(\SB4_25/i0[10] ) );
  BUF_X4 U4430 ( .I(\RI1[3][131] ), .Z(n1388) );
  XOR2_X1 U4436 ( .A1(n5585), .A2(n4815), .Z(n3042) );
  XOR2_X1 U4437 ( .A1(\RI5[0][183] ), .A2(\RI5[0][177] ), .Z(n4815) );
  NAND4_X2 U4440 ( .A1(\SB1_2_4/Component_Function_3/NAND4_in[0] ), .A2(n6126), 
        .A3(n5986), .A4(n4816), .ZN(\SB1_2_4/buf_output[3] ) );
  NAND3_X2 U4449 ( .A1(\SB1_2_4/i0_3 ), .A2(\SB1_2_4/i0_0 ), .A3(
        \SB1_2_4/i0_4 ), .ZN(n4816) );
  XOR2_X1 U4450 ( .A1(n4817), .A2(n46), .Z(Ciphertext[151]) );
  NAND4_X2 U4453 ( .A1(\SB4_6/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_6/Component_Function_1/NAND4_in[3] ), .A3(
        \SB4_6/Component_Function_1/NAND4_in[2] ), .A4(
        \SB4_6/Component_Function_1/NAND4_in[0] ), .ZN(n4817) );
  NOR2_X2 U4460 ( .A1(n1153), .A2(n4818), .ZN(\SB2_2_10/i0[7] ) );
  NAND2_X1 U4464 ( .A1(n1411), .A2(n1569), .ZN(n4818) );
  XOR2_X1 U4465 ( .A1(\SB2_3_8/buf_output[5] ), .A2(n1365), .Z(n2560) );
  NAND4_X2 U4472 ( .A1(\SB1_3_3/Component_Function_5/NAND4_in[1] ), .A2(n2258), 
        .A3(\SB1_3_3/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_3_3/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_3/buf_output[5] ) );
  XOR2_X1 U4474 ( .A1(n4819), .A2(n125), .Z(Ciphertext[25]) );
  NAND4_X2 U4476 ( .A1(\SB4_27/Component_Function_1/NAND4_in[2] ), .A2(
        \SB4_27/Component_Function_1/NAND4_in[1] ), .A3(
        \SB4_27/Component_Function_1/NAND4_in[3] ), .A4(n1921), .ZN(n4819) );
  NAND4_X2 U4477 ( .A1(\SB2_1_20/Component_Function_3/NAND4_in[0] ), .A2(n1236), .A3(\SB2_1_20/Component_Function_3/NAND4_in[3] ), .A4(n3079), .ZN(
        \SB2_1_20/buf_output[3] ) );
  INV_X1 U4479 ( .I(\SB3_5/buf_output[1] ), .ZN(\SB4_1/i1_7 ) );
  NAND4_X2 U4480 ( .A1(\SB3_5/Component_Function_1/NAND4_in[1] ), .A2(
        \SB3_5/Component_Function_1/NAND4_in[2] ), .A3(n2070), .A4(
        \SB3_5/Component_Function_1/NAND4_in[3] ), .ZN(\SB3_5/buf_output[1] )
         );
  XOR2_X1 U4481 ( .A1(n4820), .A2(n214), .Z(Ciphertext[181]) );
  NAND4_X2 U4482 ( .A1(\SB4_1/Component_Function_1/NAND4_in[1] ), .A2(n2153), 
        .A3(n4391), .A4(\SB4_1/Component_Function_1/NAND4_in[0] ), .ZN(n4820)
         );
  NAND4_X2 U4486 ( .A1(\SB4_28/Component_Function_2/NAND4_in[0] ), .A2(n2663), 
        .A3(\SB4_28/Component_Function_2/NAND4_in[2] ), .A4(n4821), .ZN(n5775)
         );
  NAND3_X1 U4490 ( .A1(\SB4_28/i0_3 ), .A2(\SB4_28/i0[6] ), .A3(
        \SB4_28/i0[10] ), .ZN(n4821) );
  XOR2_X1 U4491 ( .A1(\MC_ARK_ARC_1_2/temp1[160] ), .A2(n4822), .Z(
        \MC_ARK_ARC_1_2/temp5[160] ) );
  XOR2_X1 U4492 ( .A1(\RI5[2][130] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[106] ), 
        .Z(n4822) );
  INV_X2 U4493 ( .I(\SB1_2_8/buf_output[2] ), .ZN(\SB2_2_5/i1[9] ) );
  NAND4_X2 U4496 ( .A1(n5959), .A2(\SB1_2_8/Component_Function_2/NAND4_in[1] ), 
        .A3(\SB1_2_8/Component_Function_2/NAND4_in[2] ), .A4(n5281), .ZN(
        \SB1_2_8/buf_output[2] ) );
  NAND3_X1 U4497 ( .A1(\SB1_2_8/i0_3 ), .A2(\SB1_2_8/i0_0 ), .A3(
        \SB1_2_8/i0[7] ), .ZN(n1813) );
  INV_X2 U4498 ( .I(\SB1_2_1/buf_output[2] ), .ZN(\SB2_2_30/i1[9] ) );
  NAND4_X2 U4501 ( .A1(\SB1_2_1/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_2_1/Component_Function_2/NAND4_in[0] ), .A3(n6461), .A4(
        \SB1_2_1/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB1_2_1/buf_output[2] ) );
  AND2_X1 U4502 ( .A1(\SB2_3_6/i0[8] ), .A2(\SB1_3_11/buf_output[0] ), .Z(
        n3150) );
  NAND4_X2 U4504 ( .A1(\SB1_2_15/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_2_15/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_2_15/Component_Function_1/NAND4_in[3] ), .A4(
        \SB1_2_15/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_2_15/buf_output[1] ) );
  NAND3_X2 U4505 ( .A1(\SB2_2_16/i0_3 ), .A2(\SB2_2_16/i0[9] ), .A3(
        \SB2_2_16/i0[8] ), .ZN(\SB2_2_16/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U4508 ( .A1(\SB2_1_0/i1_5 ), .A2(\SB2_1_0/i0[8] ), .A3(
        \SB2_1_0/i3[0] ), .ZN(n2756) );
  NAND4_X2 U4511 ( .A1(n2615), .A2(n4725), .A3(n6258), .A4(n4823), .ZN(
        \SB2_3_23/buf_output[5] ) );
  XOR2_X1 U4513 ( .A1(\MC_ARK_ARC_1_1/temp2[56] ), .A2(n1132), .Z(n1885) );
  NAND4_X2 U4514 ( .A1(\SB1_3_26/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_3_26/Component_Function_5/NAND4_in[1] ), .A3(n1871), .A4(
        \SB1_3_26/Component_Function_5/NAND4_in[0] ), .ZN(\RI3[3][35] ) );
  NAND3_X1 U4515 ( .A1(\SB4_1/i0[6] ), .A2(\SB4_1/i0[9] ), .A3(\SB4_1/i1_5 ), 
        .ZN(n2153) );
  NAND4_X2 U4516 ( .A1(\SB2_1_30/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_30/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_1_30/Component_Function_2/NAND4_in[1] ), .A4(n4824), .ZN(
        \SB2_1_30/buf_output[2] ) );
  NAND3_X2 U4518 ( .A1(\SB2_1_30/i0_0 ), .A2(\SB2_1_30/i0_4 ), .A3(
        \SB2_1_30/i1_5 ), .ZN(n4824) );
  XOR2_X1 U4519 ( .A1(n3677), .A2(\RI5[2][32] ), .Z(\MC_ARK_ARC_1_2/temp1[32] ) );
  XOR2_X1 U4520 ( .A1(\MC_ARK_ARC_1_1/temp6[101] ), .A2(
        \MC_ARK_ARC_1_1/temp5[101] ), .Z(\MC_ARK_ARC_1_1/buf_output[101] ) );
  XOR2_X1 U4522 ( .A1(\MC_ARK_ARC_1_1/temp4[101] ), .A2(n5095), .Z(
        \MC_ARK_ARC_1_1/temp6[101] ) );
  XOR2_X1 U4523 ( .A1(\MC_ARK_ARC_1_2/temp5[45] ), .A2(
        \MC_ARK_ARC_1_2/temp6[45] ), .Z(\MC_ARK_ARC_1_2/buf_output[45] ) );
  XOR2_X1 U4530 ( .A1(\MC_ARK_ARC_1_2/temp2[45] ), .A2(n1500), .Z(
        \MC_ARK_ARC_1_2/temp5[45] ) );
  XOR2_X1 U4536 ( .A1(n2235), .A2(n4825), .Z(n6176) );
  XOR2_X1 U4538 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[149] ), .A2(\RI5[2][113] ), 
        .Z(n4825) );
  XOR2_X1 U4544 ( .A1(n4827), .A2(n4826), .Z(\MC_ARK_ARC_1_2/temp5[56] ) );
  XOR2_X1 U4550 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[2] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[56] ), .Z(n4826) );
  XOR2_X1 U4553 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[50] ), .A2(n3677), .Z(
        n4827) );
  XOR2_X1 U4559 ( .A1(n4828), .A2(n187), .Z(Ciphertext[180]) );
  NAND4_X2 U4561 ( .A1(\SB4_1/Component_Function_0/NAND4_in[3] ), .A2(
        \SB4_1/Component_Function_0/NAND4_in[2] ), .A3(n4853), .A4(n4954), 
        .ZN(n4828) );
  XOR2_X1 U4562 ( .A1(\MC_ARK_ARC_1_1/temp4[92] ), .A2(n4829), .Z(
        \MC_ARK_ARC_1_1/temp6[92] ) );
  XOR2_X1 U4563 ( .A1(\RI5[1][2] ), .A2(\RI5[1][158] ), .Z(n4829) );
  NAND4_X2 U4564 ( .A1(\SB2_2_0/Component_Function_5/NAND4_in[2] ), .A2(n1609), 
        .A3(n4987), .A4(n4121), .ZN(\SB2_2_0/buf_output[5] ) );
  NAND4_X2 U4565 ( .A1(\SB2_1_2/Component_Function_5/NAND4_in[2] ), .A2(n2583), 
        .A3(\SB2_1_2/Component_Function_5/NAND4_in[0] ), .A4(n4830), .ZN(
        \SB2_1_2/buf_output[5] ) );
  NAND3_X2 U4570 ( .A1(\SB2_1_2/i0[9] ), .A2(\SB2_1_2/i0[6] ), .A3(
        \SB2_1_2/i0_4 ), .ZN(n4830) );
  XOR2_X1 U4571 ( .A1(n4831), .A2(n230), .Z(Ciphertext[183]) );
  NAND4_X2 U4572 ( .A1(n6195), .A2(\SB4_1/Component_Function_3/NAND4_in[3] ), 
        .A3(n4891), .A4(n2960), .ZN(n4831) );
  XOR2_X1 U4574 ( .A1(n3718), .A2(\MC_ARK_ARC_1_2/temp5[125] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[125] ) );
  XOR2_X1 U4578 ( .A1(n4842), .A2(n4841), .Z(n3718) );
  XOR2_X1 U4579 ( .A1(n4832), .A2(n2530), .Z(n2610) );
  XOR2_X1 U4581 ( .A1(\RI5[3][26] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[56] ), 
        .Z(n4832) );
  XOR2_X1 U4583 ( .A1(\MC_ARK_ARC_1_2/temp4[63] ), .A2(n4833), .Z(n5056) );
  XOR2_X1 U4586 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[129] ), .A2(\RI5[2][165] ), 
        .Z(n4833) );
  NAND3_X2 U4587 ( .A1(\SB1_2_6/i0[10] ), .A2(\SB1_2_6/i1[9] ), .A3(
        \SB1_2_6/i1_5 ), .ZN(n5097) );
  NAND3_X2 U4588 ( .A1(\SB2_2_3/i0_0 ), .A2(\SB1_2_4/buf_output[4] ), .A3(
        \SB2_2_3/i1_5 ), .ZN(\SB2_2_3/Component_Function_2/NAND4_in[3] ) );
  NAND4_X2 U4589 ( .A1(n2429), .A2(\SB2_1_16/Component_Function_5/NAND4_in[1] ), .A3(n4846), .A4(\SB2_1_16/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_1_16/buf_output[5] ) );
  NAND3_X2 U4593 ( .A1(\SB1_3_31/i0_0 ), .A2(\SB1_3_31/i1_7 ), .A3(
        \SB1_3_31/i3[0] ), .ZN(\SB1_3_31/Component_Function_4/NAND4_in[1] ) );
  NAND3_X2 U4594 ( .A1(\RI3[0][15] ), .A2(\SB2_0_29/i1[9] ), .A3(
        \SB2_0_29/i1_5 ), .ZN(\SB2_0_29/Component_Function_2/NAND4_in[0] ) );
  INV_X2 U4598 ( .I(\SB1_1_13/buf_output[2] ), .ZN(\SB2_1_10/i1[9] ) );
  NAND4_X2 U4599 ( .A1(\SB1_1_13/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_13/Component_Function_2/NAND4_in[1] ), .A3(n6058), .A4(n4240), 
        .ZN(\SB1_1_13/buf_output[2] ) );
  NAND3_X2 U4603 ( .A1(\SB4_2/i0[10] ), .A2(\SB4_2/i1_5 ), .A3(\SB4_2/i1[9] ), 
        .ZN(n5272) );
  NAND3_X1 U4612 ( .A1(\SB2_3_7/i0_3 ), .A2(n3739), .A3(\SB2_3_7/i0_0 ), .ZN(
        \SB2_3_7/Component_Function_0/NAND4_in[3] ) );
  XOR2_X1 U4613 ( .A1(\MC_ARK_ARC_1_2/temp4[146] ), .A2(n4834), .Z(n5787) );
  XOR2_X1 U4614 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[116] ), .A2(
        \SB2_2_11/buf_output[2] ), .Z(n4834) );
  NAND3_X1 U4615 ( .A1(\SB1_3_12/i0[9] ), .A2(\SB1_3_12/i0_0 ), .A3(
        \SB1_3_12/i0[8] ), .ZN(n4835) );
  NAND4_X2 U4619 ( .A1(\SB2_2_3/Component_Function_2/NAND4_in[2] ), .A2(n3942), 
        .A3(n1149), .A4(\SB2_2_3/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_2_3/buf_output[2] ) );
  NAND4_X2 U4622 ( .A1(n3531), .A2(n4968), .A3(
        \SB2_3_19/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_3_19/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_3_19/buf_output[5] ) );
  NAND3_X2 U4629 ( .A1(\SB2_1_16/i0_0 ), .A2(\SB2_1_16/i0_3 ), .A3(
        \SB2_1_16/i0_4 ), .ZN(\SB2_1_16/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U4630 ( .A1(\SB1_3_19/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_19/Component_Function_5/NAND4_in[2] ), .A3(n6252), .A4(
        \SB1_3_19/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_19/buf_output[5] ) );
  NAND4_X2 U4633 ( .A1(\SB2_1_26/Component_Function_3/NAND4_in[3] ), .A2(
        \SB2_1_26/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_1_26/Component_Function_3/NAND4_in[0] ), .A4(
        \SB2_1_26/Component_Function_3/NAND4_in[1] ), .ZN(
        \SB2_1_26/buf_output[3] ) );
  XOR2_X1 U4637 ( .A1(\MC_ARK_ARC_1_3/temp1[143] ), .A2(n4836), .Z(
        \MC_ARK_ARC_1_3/temp5[143] ) );
  XOR2_X1 U4639 ( .A1(\RI5[3][113] ), .A2(\RI5[3][89] ), .Z(n4836) );
  XOR2_X1 U4640 ( .A1(\RI5[2][26] ), .A2(\SB2_2_24/buf_output[2] ), .Z(n6088)
         );
  NAND4_X2 U4656 ( .A1(\SB1_2_14/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_2_14/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_2_14/Component_Function_3/NAND4_in[3] ), .A4(n4837), .ZN(
        \SB1_2_14/buf_output[3] ) );
  NAND3_X2 U4659 ( .A1(\SB1_2_14/i0[10] ), .A2(\SB1_2_14/i1_7 ), .A3(
        \SB1_2_14/i1[9] ), .ZN(n4837) );
  XOR2_X1 U4664 ( .A1(n4839), .A2(n4838), .Z(n1655) );
  XOR2_X1 U4666 ( .A1(\RI5[0][15] ), .A2(n192), .Z(n4838) );
  XOR2_X1 U4667 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[105] ), .A2(\RI5[0][39] ), 
        .Z(n4839) );
  NAND3_X2 U4679 ( .A1(\SB1_3_21/i0_0 ), .A2(\SB1_3_21/i0_4 ), .A3(
        \SB1_3_21/i1_5 ), .ZN(n4840) );
  NAND3_X1 U4681 ( .A1(\SB3_28/i0[8] ), .A2(\SB3_28/i1_5 ), .A3(\SB3_28/i3[0] ), .ZN(n2319) );
  XOR2_X1 U4682 ( .A1(\MC_ARK_ARC_1_2/temp3[86] ), .A2(
        \MC_ARK_ARC_1_2/temp4[86] ), .Z(\MC_ARK_ARC_1_2/temp6[86] ) );
  XOR2_X1 U4683 ( .A1(\RI5[2][191] ), .A2(n463), .Z(n4841) );
  XOR2_X1 U4687 ( .A1(\RI5[2][35] ), .A2(\RI5[2][161] ), .Z(n4842) );
  XOR2_X1 U4689 ( .A1(n4843), .A2(n107), .Z(Ciphertext[172]) );
  NAND4_X2 U4692 ( .A1(n4681), .A2(\SB2_3_16/Component_Function_5/NAND4_in[0] ), .A3(\SB2_3_16/Component_Function_5/NAND4_in[2] ), .A4(n4844), .ZN(
        \SB2_3_16/buf_output[5] ) );
  NAND3_X2 U4701 ( .A1(\SB2_3_16/i0[10] ), .A2(\SB2_3_16/i0[6] ), .A3(
        \SB2_3_16/i0_0 ), .ZN(n4844) );
  NAND3_X2 U4702 ( .A1(\SB1_3_21/i0_0 ), .A2(\SB1_3_21/i0_3 ), .A3(
        \SB1_3_21/i0_4 ), .ZN(n4845) );
  NAND3_X2 U4707 ( .A1(\SB2_1_16/i0[6] ), .A2(\SB2_1_16/i0_4 ), .A3(
        \SB2_1_16/i0[9] ), .ZN(n4846) );
  NAND2_X2 U4708 ( .A1(n2891), .A2(n4847), .ZN(\SB2_1_7/i0_4 ) );
  AND2_X1 U4711 ( .A1(n4907), .A2(\SB1_1_8/Component_Function_4/NAND4_in[1] ), 
        .Z(n4847) );
  INV_X1 U4718 ( .I(\SB1_0_3/buf_output[0] ), .ZN(\SB2_0_30/i3[0] ) );
  NAND4_X2 U4719 ( .A1(\SB1_0_3/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_0_3/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_0_3/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_0_3/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_0_3/buf_output[0] ) );
  XOR2_X1 U4727 ( .A1(n3762), .A2(n4848), .Z(\MC_ARK_ARC_1_2/temp5[189] ) );
  XOR2_X1 U4732 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[183] ), .A2(n1390), .Z(
        n4848) );
  NAND3_X2 U4733 ( .A1(\SB2_1_22/i0_4 ), .A2(\SB2_1_22/i1_5 ), .A3(
        \SB2_1_22/i0_0 ), .ZN(n1798) );
  NAND3_X1 U4734 ( .A1(\SB2_3_25/i0[6] ), .A2(\SB1_3_30/buf_output[0] ), .A3(
        \SB1_3_26/buf_output[4] ), .ZN(
        \SB2_3_25/Component_Function_5/NAND4_in[3] ) );
  XOR2_X1 U4735 ( .A1(\MC_ARK_ARC_1_3/temp4[167] ), .A2(n5094), .Z(
        \MC_ARK_ARC_1_3/temp6[167] ) );
  NAND4_X2 U4736 ( .A1(\SB1_2_17/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_2_17/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_2_17/Component_Function_1/NAND4_in[0] ), .A4(n3979), .ZN(
        \SB1_2_17/buf_output[1] ) );
  NAND4_X2 U4737 ( .A1(n2217), .A2(\SB2_1_22/Component_Function_5/NAND4_in[3] ), .A3(\SB2_1_22/Component_Function_5/NAND4_in[0] ), .A4(n4849), .ZN(
        \SB2_1_22/buf_output[5] ) );
  NAND3_X2 U4740 ( .A1(\SB2_1_22/i0[6] ), .A2(\SB2_1_22/i0[10] ), .A3(
        \SB2_1_22/i0_0 ), .ZN(n4849) );
  XOR2_X1 U4742 ( .A1(\MC_ARK_ARC_1_1/temp3[89] ), .A2(n4850), .Z(n5081) );
  XOR2_X1 U4743 ( .A1(\RI5[1][59] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[35] ), 
        .Z(n4850) );
  NAND4_X2 U4744 ( .A1(n691), .A2(\SB4_30/Component_Function_4/NAND4_in[3] ), 
        .A3(\SB4_30/Component_Function_4/NAND4_in[1] ), .A4(n4851), .ZN(n5064)
         );
  NAND3_X2 U4745 ( .A1(\SB1_0_17/i0_3 ), .A2(n2899), .A3(\SB1_0_17/i1[9] ), 
        .ZN(\SB1_0_17/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U4750 ( .A1(n4852), .A2(n202), .Z(Ciphertext[171]) );
  NAND4_X2 U4751 ( .A1(n5133), .A2(\SB4_3/Component_Function_3/NAND4_in[3] ), 
        .A3(n2777), .A4(\SB4_3/Component_Function_3/NAND4_in[2] ), .ZN(n4852)
         );
  NAND3_X1 U4755 ( .A1(\SB4_1/i0[6] ), .A2(\SB4_1/i0[7] ), .A3(\SB4_1/i0[8] ), 
        .ZN(n4853) );
  NAND3_X1 U4756 ( .A1(n3662), .A2(\SB4_18/i1_5 ), .A3(\SB4_18/i3[0] ), .ZN(
        \SB4_18/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U4757 ( .A1(n1349), .A2(n4854), .Z(\MC_ARK_ARC_1_2/buf_output[19] )
         );
  XOR2_X1 U4762 ( .A1(\MC_ARK_ARC_1_2/temp4[19] ), .A2(n4470), .Z(n4854) );
  NAND4_X2 U4771 ( .A1(\SB2_2_1/Component_Function_5/NAND4_in[2] ), .A2(n5469), 
        .A3(\SB2_2_1/Component_Function_5/NAND4_in[0] ), .A4(n4855), .ZN(
        \SB2_2_1/buf_output[5] ) );
  NAND3_X2 U4772 ( .A1(\SB2_2_1/i0[6] ), .A2(\SB2_2_1/i0_0 ), .A3(
        \SB2_2_1/i0[10] ), .ZN(n4855) );
  XOR2_X1 U4774 ( .A1(n4857), .A2(n4856), .Z(\MC_ARK_ARC_1_2/buf_output[116] )
         );
  XOR2_X1 U4776 ( .A1(n6481), .A2(\MC_ARK_ARC_1_2/temp4[116] ), .Z(n4856) );
  XOR2_X1 U4777 ( .A1(n632), .A2(n4885), .Z(n4857) );
  INV_X2 U4779 ( .I(\SB1_2_11/buf_output[5] ), .ZN(\SB2_2_11/i1_5 ) );
  NAND4_X2 U4780 ( .A1(\SB1_2_11/Component_Function_5/NAND4_in[3] ), .A2(n5116), .A3(n3820), .A4(\SB1_2_11/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_2_11/buf_output[5] ) );
  BUF_X4 U4784 ( .I(\SB2_3_24/buf_output[1] ), .Z(\RI5[3][67] ) );
  NAND4_X2 U4785 ( .A1(n2880), .A2(\SB4_29/Component_Function_5/NAND4_in[2] ), 
        .A3(\SB4_29/Component_Function_5/NAND4_in[0] ), .A4(n4858), .ZN(n5431)
         );
  NAND3_X2 U4786 ( .A1(\SB4_29/i0[10] ), .A2(\SB4_29/i0[6] ), .A3(
        \SB4_29/i0_0 ), .ZN(n4858) );
  XOR2_X1 U4787 ( .A1(\MC_ARK_ARC_1_3/temp5[137] ), .A2(n4859), .Z(
        \MC_ARK_ARC_1_3/buf_output[137] ) );
  XOR2_X1 U4791 ( .A1(\MC_ARK_ARC_1_3/temp4[137] ), .A2(
        \MC_ARK_ARC_1_3/temp3[137] ), .Z(n4859) );
  NAND4_X2 U4793 ( .A1(\SB2_0_10/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_10/Component_Function_2/NAND4_in[3] ), .A3(n4861), .A4(n4860), 
        .ZN(\SB2_0_10/buf_output[2] ) );
  NAND3_X2 U4795 ( .A1(\SB2_0_10/i0[10] ), .A2(\SB2_0_10/i0[6] ), .A3(
        \SB2_0_10/i0_3 ), .ZN(n4860) );
  NAND3_X2 U4797 ( .A1(n571), .A2(\SB2_0_10/i0_3 ), .A3(\SB2_0_10/i0[8] ), 
        .ZN(n4861) );
  NAND3_X1 U4798 ( .A1(\SB2_2_15/i0_0 ), .A2(\SB2_2_15/i3[0] ), .A3(
        \SB2_2_15/i1_7 ), .ZN(\SB2_2_15/Component_Function_4/NAND4_in[1] ) );
  NOR2_X2 U4801 ( .A1(n4491), .A2(n4862), .ZN(\SB2_3_25/i0[7] ) );
  XOR2_X1 U4806 ( .A1(n4863), .A2(n40), .Z(Ciphertext[144]) );
  NAND4_X2 U4810 ( .A1(\SB4_7/Component_Function_0/NAND4_in[3] ), .A2(n3597), 
        .A3(\SB4_7/Component_Function_0/NAND4_in[1] ), .A4(
        \SB4_7/Component_Function_0/NAND4_in[0] ), .ZN(n4863) );
  XOR2_X1 U4811 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[9] ), .A2(
        \SB2_1_6/buf_output[3] ), .Z(n5777) );
  NAND3_X1 U4813 ( .A1(\SB4_14/i0_0 ), .A2(\SB4_14/i3[0] ), .A3(\SB4_14/i1_7 ), 
        .ZN(n1302) );
  NAND4_X2 U4814 ( .A1(n731), .A2(\SB2_0_23/Component_Function_2/NAND4_in[1] ), 
        .A3(\SB2_0_23/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_0_23/Component_Function_2/NAND4_in[0] ), .ZN(
        \SB2_0_23/buf_output[2] ) );
  NAND4_X2 U4816 ( .A1(\SB2_2_15/Component_Function_2/NAND4_in[3] ), .A2(n3615), .A3(\SB2_2_15/Component_Function_2/NAND4_in[0] ), .A4(n3152), .ZN(
        \SB2_2_15/buf_output[2] ) );
  NAND4_X2 U4821 ( .A1(\SB2_0_13/Component_Function_5/NAND4_in[2] ), .A2(n957), 
        .A3(\SB2_0_13/Component_Function_5/NAND4_in[0] ), .A4(n5668), .ZN(
        \SB2_0_13/buf_output[5] ) );
  XOR2_X1 U4823 ( .A1(n4865), .A2(n4864), .Z(\MC_ARK_ARC_1_1/temp5[164] ) );
  XOR2_X1 U4824 ( .A1(\RI5[1][134] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[110] ), 
        .Z(n4864) );
  XOR2_X1 U4826 ( .A1(\RI5[1][164] ), .A2(\RI5[1][158] ), .Z(n4865) );
  NAND3_X1 U4829 ( .A1(\SB2_3_15/i0_0 ), .A2(\SB1_3_16/buf_output[4] ), .A3(
        \SB2_3_15/i1_5 ), .ZN(\SB2_3_15/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 U4830 ( .A1(\SB1_3_2/i0[9] ), .A2(\SB1_3_2/i0[6] ), .A3(
        \SB1_3_2/i0_4 ), .ZN(n6345) );
  NAND3_X2 U4831 ( .A1(\SB2_0_11/i0_3 ), .A2(\SB2_0_11/i0[6] ), .A3(
        \SB2_0_11/i0[10] ), .ZN(\SB2_0_11/Component_Function_2/NAND4_in[1] )
         );
  NAND3_X1 U4833 ( .A1(\SB2_2_14/i0[7] ), .A2(\SB2_2_14/i0_0 ), .A3(
        \SB2_2_14/i0_3 ), .ZN(\SB2_2_14/Component_Function_0/NAND4_in[3] ) );
  XOR2_X1 U4837 ( .A1(\MC_ARK_ARC_1_1/temp6[57] ), .A2(
        \MC_ARK_ARC_1_1/temp5[57] ), .Z(\MC_ARK_ARC_1_1/buf_output[57] ) );
  NAND3_X1 U4839 ( .A1(\SB1_3_30/i0[10] ), .A2(\SB1_3_30/i0_3 ), .A3(
        \SB1_3_30/i0_4 ), .ZN(\SB1_3_30/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U4841 ( .A1(\SB4_23/i0_3 ), .A2(\SB4_23/i1[9] ), .A3(\SB4_23/i0[6] ), .ZN(\SB4_23/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U4847 ( .A1(\RI5[2][184] ), .A2(\RI5[2][28] ), .Z(n5067) );
  NAND3_X1 U4848 ( .A1(\SB1_2_16/i0[8] ), .A2(\RI1[2][95] ), .A3(
        \MC_ARK_ARC_1_1/buf_output[90] ), .ZN(
        \SB1_2_16/Component_Function_2/NAND4_in[2] ) );
  XOR2_X1 U4857 ( .A1(n4867), .A2(n4866), .Z(\MC_ARK_ARC_1_1/temp5[98] ) );
  XOR2_X1 U4859 ( .A1(\RI5[1][98] ), .A2(\RI5[1][68] ), .Z(n4866) );
  XOR2_X1 U4862 ( .A1(\RI5[1][44] ), .A2(\RI5[1][92] ), .Z(n4867) );
  NAND3_X1 U4863 ( .A1(\SB1_2_15/i0[10] ), .A2(\SB1_2_15/i1[9] ), .A3(
        \SB1_2_15/i1_5 ), .ZN(\SB1_2_15/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U4869 ( .A1(\SB2_0_15/i0[10] ), .A2(\SB2_0_15/i1_7 ), .A3(
        \SB2_0_15/i1[9] ), .ZN(n5679) );
  NAND4_X2 U4870 ( .A1(\SB2_1_25/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_25/Component_Function_3/NAND4_in[3] ), .A3(n4978), .A4(n2067), 
        .ZN(\SB2_1_25/buf_output[3] ) );
  NAND3_X2 U4875 ( .A1(\SB2_1_6/i0_3 ), .A2(\SB2_1_6/i0_0 ), .A3(
        \SB2_1_6/i0_4 ), .ZN(\SB2_1_6/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U4878 ( .A1(n3509), .A2(\SB2_3_9/Component_Function_5/NAND4_in[1] ), 
        .A3(\SB2_3_9/Component_Function_5/NAND4_in[0] ), .A4(n1403), .ZN(
        \SB2_3_9/buf_output[5] ) );
  XOR2_X1 U4880 ( .A1(n4869), .A2(n4868), .Z(\MC_ARK_ARC_1_3/buf_output[39] )
         );
  XOR2_X1 U4881 ( .A1(n5700), .A2(\MC_ARK_ARC_1_3/temp4[39] ), .Z(n4868) );
  XOR2_X1 U4887 ( .A1(\MC_ARK_ARC_1_3/temp2[39] ), .A2(
        \MC_ARK_ARC_1_3/temp3[39] ), .Z(n4869) );
  XOR2_X1 U4890 ( .A1(\MC_ARK_ARC_1_0/temp5[89] ), .A2(n4627), .Z(
        \MC_ARK_ARC_1_0/buf_output[89] ) );
  NAND4_X2 U4893 ( .A1(\SB3_7/Component_Function_4/NAND4_in[1] ), .A2(
        \SB3_7/Component_Function_4/NAND4_in[3] ), .A3(
        \SB3_7/Component_Function_4/NAND4_in[0] ), .A4(n4870), .ZN(
        \SB3_7/buf_output[4] ) );
  XOR2_X1 U4896 ( .A1(\MC_ARK_ARC_1_3/temp6[165] ), .A2(
        \MC_ARK_ARC_1_3/temp5[165] ), .Z(\MC_ARK_ARC_1_3/buf_output[165] ) );
  NAND4_X2 U4898 ( .A1(\SB2_1_18/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_1_18/Component_Function_2/NAND4_in[0] ), .A3(n4979), .A4(
        \SB2_1_18/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_1_18/buf_output[2] ) );
  NAND3_X1 U4900 ( .A1(\SB2_0_10/i0_0 ), .A2(\SB2_0_10/i0_4 ), .A3(
        \SB2_0_10/i1_5 ), .ZN(\SB2_0_10/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U4901 ( .A1(\SB1_2_7/i0[10] ), .A2(\SB1_2_7/i1_7 ), .A3(
        \SB1_2_7/i1[9] ), .ZN(n2856) );
  NAND4_X2 U4902 ( .A1(\SB2_3_2/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_3_2/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_2/Component_Function_2/NAND4_in[3] ), .A4(n5204), .ZN(
        \SB2_3_2/buf_output[2] ) );
  XOR2_X1 U4903 ( .A1(\RI5[1][55] ), .A2(\RI5[1][19] ), .Z(
        \MC_ARK_ARC_1_1/temp3[145] ) );
  NAND4_X2 U4905 ( .A1(\SB2_1_11/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_1_11/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_1_11/Component_Function_2/NAND4_in[3] ), .A4(n4871), .ZN(
        \SB2_1_11/buf_output[2] ) );
  NAND3_X2 U4906 ( .A1(\SB2_1_11/i0[10] ), .A2(\SB2_1_11/i1_5 ), .A3(
        \SB2_1_11/i1[9] ), .ZN(n4871) );
  NAND3_X1 U4907 ( .A1(\SB2_3_5/i0_4 ), .A2(\SB2_3_5/i1_7 ), .A3(
        \SB2_3_5/i0[8] ), .ZN(\SB2_3_5/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U4908 ( .A1(n2706), .A2(\SB1_1_19/Component_Function_5/NAND4_in[2] ), .A3(n5001), .A4(\SB1_1_19/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_19/buf_output[5] ) );
  XOR2_X1 U4909 ( .A1(\RI5[0][68] ), .A2(\RI5[0][62] ), .Z(n3247) );
  XOR2_X1 U4910 ( .A1(\RI5[3][55] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[49] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[55] ) );
  NAND3_X1 U4916 ( .A1(\SB4_23/i0_3 ), .A2(\SB4_23/i0[9] ), .A3(
        \SB4_23/i0[10] ), .ZN(\SB4_23/Component_Function_4/NAND4_in[2] ) );
  NAND4_X2 U4917 ( .A1(n2459), .A2(\SB2_3_6/Component_Function_3/NAND4_in[0] ), 
        .A3(\SB2_3_6/Component_Function_3/NAND4_in[3] ), .A4(n4872), .ZN(
        \SB2_3_6/buf_output[3] ) );
  NAND3_X2 U4918 ( .A1(\SB2_3_6/i0_4 ), .A2(\SB2_3_6/i0_0 ), .A3(
        \SB2_3_6/i0_3 ), .ZN(n4872) );
  INV_X1 U4919 ( .I(\SB3_17/buf_output[5] ), .ZN(\SB4_17/i1_5 ) );
  NAND4_X2 U4922 ( .A1(\SB3_17/Component_Function_5/NAND4_in[2] ), .A2(
        \SB3_17/Component_Function_5/NAND4_in[1] ), .A3(n5946), .A4(
        \SB3_17/Component_Function_5/NAND4_in[0] ), .ZN(\SB3_17/buf_output[5] ) );
  NAND4_X2 U4924 ( .A1(\SB1_1_25/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_1_25/Component_Function_3/NAND4_in[0] ), .A3(n4691), .A4(n4873), 
        .ZN(\SB1_1_25/buf_output[3] ) );
  XOR2_X1 U4930 ( .A1(\RI5[3][23] ), .A2(\RI5[3][47] ), .Z(n3422) );
  NAND4_X2 U4931 ( .A1(\SB1_2_13/Component_Function_3/NAND4_in[1] ), .A2(n2122), .A3(n2763), .A4(\SB1_2_13/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_2_13/buf_output[3] ) );
  NAND4_X2 U4933 ( .A1(\SB2_3_15/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_15/Component_Function_4/NAND4_in[3] ), .A3(n643), .A4(
        \SB2_3_15/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB2_3_15/buf_output[4] ) );
  NAND4_X2 U4941 ( .A1(\SB2_1_4/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_1_4/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_4/Component_Function_0/NAND4_in[0] ), .A4(n845), .ZN(
        \SB2_1_4/buf_output[0] ) );
  NAND3_X1 U4942 ( .A1(\SB2_2_11/i0_3 ), .A2(\SB2_2_11/i0[8] ), .A3(
        \SB2_2_11/i1_7 ), .ZN(\SB2_2_11/Component_Function_1/NAND4_in[1] ) );
  NAND4_X2 U4943 ( .A1(\SB2_0_14/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_0_14/Component_Function_1/NAND4_in[1] ), .A3(n5796), .A4(
        \SB2_0_14/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_0_14/buf_output[1] ) );
  NAND4_X2 U4955 ( .A1(\SB1_3_18/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_18/Component_Function_2/NAND4_in[2] ), .A3(
        \SB1_3_18/Component_Function_2/NAND4_in[0] ), .A4(n3752), .ZN(
        \SB1_3_18/buf_output[2] ) );
  XOR2_X1 U4956 ( .A1(\SB2_0_5/buf_output[3] ), .A2(\RI5[0][177] ), .Z(n5150)
         );
  NAND3_X2 U4958 ( .A1(\SB1_1_14/i0[10] ), .A2(\SB1_1_14/i1[9] ), .A3(
        \SB1_1_14/i1_5 ), .ZN(n5145) );
  NAND4_X2 U4962 ( .A1(\SB2_1_8/Component_Function_2/NAND4_in[0] ), .A2(n2379), 
        .A3(n3091), .A4(\SB2_1_8/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB2_1_8/buf_output[2] ) );
  NAND4_X2 U4965 ( .A1(\SB4_17/Component_Function_3/NAND4_in[3] ), .A2(
        \SB4_17/Component_Function_3/NAND4_in[2] ), .A3(n2098), .A4(n4874), 
        .ZN(n3172) );
  NAND3_X1 U4969 ( .A1(\SB4_17/i0[6] ), .A2(\SB4_17/i0_3 ), .A3(\SB4_17/i1[9] ), .ZN(n4874) );
  XOR2_X1 U4976 ( .A1(\MC_ARK_ARC_1_2/temp4[120] ), .A2(
        \MC_ARK_ARC_1_2/temp3[120] ), .Z(n2184) );
  NAND4_X2 U4977 ( .A1(\SB3_22/Component_Function_4/NAND4_in[1] ), .A2(
        \SB3_22/Component_Function_4/NAND4_in[0] ), .A3(
        \SB3_22/Component_Function_4/NAND4_in[3] ), .A4(
        \SB3_22/Component_Function_4/NAND4_in[2] ), .ZN(\SB3_22/buf_output[4] ) );
  NAND4_X2 U4982 ( .A1(\SB2_1_16/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_16/Component_Function_2/NAND4_in[1] ), .A3(n2998), .A4(n5461), 
        .ZN(\SB2_1_16/buf_output[2] ) );
  XOR2_X1 U4989 ( .A1(n1937), .A2(n4253), .Z(\MC_ARK_ARC_1_2/buf_output[183] )
         );
  NAND4_X2 U4991 ( .A1(\SB1_3_7/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_7/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_7/Component_Function_4/NAND4_in[3] ), .A4(
        \SB1_3_7/Component_Function_4/NAND4_in[2] ), .ZN(
        \SB1_3_7/buf_output[4] ) );
  NAND4_X2 U4993 ( .A1(\SB1_3_15/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_15/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_3_15/Component_Function_2/NAND4_in[3] ), .A4(n4906), .ZN(
        \SB1_3_15/buf_output[2] ) );
  NAND4_X2 U4997 ( .A1(\SB1_3_31/Component_Function_5/NAND4_in[2] ), .A2(n1251), .A3(\SB1_3_31/Component_Function_5/NAND4_in[1] ), .A4(
        \SB1_3_31/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_31/buf_output[5] ) );
  NAND2_X1 U4998 ( .A1(\SB1_3_26/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_26/Component_Function_4/NAND4_in[2] ), .ZN(n4491) );
  NAND4_X2 U5002 ( .A1(\SB1_3_11/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_11/Component_Function_4/NAND4_in[3] ), .A3(n5136), .A4(
        \SB1_3_11/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB1_3_11/buf_output[4] ) );
  NAND4_X2 U5003 ( .A1(n2351), .A2(\SB1_0_10/Component_Function_5/NAND4_in[2] ), .A3(\SB1_0_10/Component_Function_5/NAND4_in[0] ), .A4(
        \SB1_0_10/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[0][131] ) );
  XOR2_X1 U5006 ( .A1(\MC_ARK_ARC_1_0/temp6[61] ), .A2(
        \MC_ARK_ARC_1_0/temp5[61] ), .Z(\MC_ARK_ARC_1_0/buf_output[61] ) );
  NAND3_X1 U5012 ( .A1(\SB1_1_8/i0[9] ), .A2(\SB1_1_8/i0[8] ), .A3(
        \SB1_1_8/i0_0 ), .ZN(\SB1_1_8/Component_Function_4/NAND4_in[0] ) );
  NAND4_X1 U5013 ( .A1(\SB3_15/Component_Function_3/NAND4_in[1] ), .A2(
        \SB3_15/Component_Function_3/NAND4_in[0] ), .A3(n4423), .A4(n4137), 
        .ZN(\SB3_15/buf_output[3] ) );
  XOR2_X1 U5014 ( .A1(\RI5[0][101] ), .A2(\RI5[0][65] ), .Z(
        \MC_ARK_ARC_1_0/temp3[191] ) );
  NAND3_X1 U5020 ( .A1(\SB1_1_30/i0_3 ), .A2(\SB1_1_30/i0[8] ), .A3(
        \SB1_1_30/i1_7 ), .ZN(\SB1_1_30/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U5022 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[153] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[129] ), .Z(\MC_ARK_ARC_1_2/temp2[183] )
         );
  NAND4_X2 U5023 ( .A1(\SB4_27/Component_Function_5/NAND4_in[3] ), .A2(n2695), 
        .A3(\SB4_27/Component_Function_5/NAND4_in[1] ), .A4(
        \SB4_27/Component_Function_5/NAND4_in[0] ), .ZN(n6538) );
  XOR2_X1 U5025 ( .A1(\MC_ARK_ARC_1_1/temp2[95] ), .A2(n4875), .Z(n767) );
  XOR2_X1 U5036 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[89] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[95] ), .Z(n4875) );
  XOR2_X1 U5037 ( .A1(\RI5[1][128] ), .A2(\RI5[1][152] ), .Z(
        \MC_ARK_ARC_1_1/temp2[182] ) );
  XOR2_X1 U5040 ( .A1(n4336), .A2(\MC_ARK_ARC_1_3/temp6[71] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[71] ) );
  XOR2_X1 U5042 ( .A1(n4303), .A2(\MC_ARK_ARC_1_3/temp6[55] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[55] ) );
  XOR2_X1 U5046 ( .A1(n3877), .A2(n3876), .Z(n616) );
  NAND4_X2 U5048 ( .A1(\SB1_0_21/Component_Function_5/NAND4_in[2] ), .A2(n5672), .A3(\SB1_0_21/Component_Function_5/NAND4_in[3] ), .A4(
        \SB1_0_21/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_0_21/buf_output[5] ) );
  NAND4_X2 U5052 ( .A1(n3551), .A2(\SB1_1_27/Component_Function_1/NAND4_in[1] ), .A3(\SB1_1_27/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_1_27/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_1_27/buf_output[1] ) );
  NAND4_X2 U5053 ( .A1(n4188), .A2(n4156), .A3(
        \SB4_17/Component_Function_4/NAND4_in[0] ), .A4(n1679), .ZN(n6226) );
  XOR2_X1 U5054 ( .A1(n4876), .A2(n178), .Z(Ciphertext[70]) );
  NAND4_X2 U5055 ( .A1(\SB4_20/Component_Function_4/NAND4_in[3] ), .A2(
        \SB4_20/Component_Function_4/NAND4_in[1] ), .A3(
        \SB4_20/Component_Function_4/NAND4_in[0] ), .A4(n6269), .ZN(n4876) );
  NAND4_X2 U5063 ( .A1(\SB4_3/Component_Function_1/NAND4_in[2] ), .A2(
        \SB4_3/Component_Function_1/NAND4_in[3] ), .A3(
        \SB4_3/Component_Function_1/NAND4_in[1] ), .A4(
        \SB4_3/Component_Function_1/NAND4_in[0] ), .ZN(n4006) );
  NAND4_X2 U5067 ( .A1(\SB2_2_16/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_16/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_2_16/Component_Function_4/NAND4_in[1] ), .A4(
        \SB2_2_16/Component_Function_4/NAND4_in[2] ), .ZN(
        \SB2_2_16/buf_output[4] ) );
  NAND4_X2 U5075 ( .A1(n4983), .A2(\SB2_1_26/Component_Function_1/NAND4_in[3] ), .A3(\SB2_1_26/Component_Function_1/NAND4_in[1] ), .A4(
        \SB2_1_26/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_1_26/buf_output[1] ) );
  XOR2_X1 U5077 ( .A1(\MC_ARK_ARC_1_0/temp5[141] ), .A2(n6527), .Z(
        \MC_ARK_ARC_1_0/buf_output[141] ) );
  XOR2_X1 U5078 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[2] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[38] ), .Z(n4060) );
  NAND4_X2 U5079 ( .A1(\SB4_27/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_27/Component_Function_0/NAND4_in[1] ), .A3(n2071), .A4(n3271), 
        .ZN(n2010) );
  XOR2_X1 U5081 ( .A1(n4877), .A2(n147), .Z(Ciphertext[127]) );
  NAND4_X2 U5082 ( .A1(\SB4_10/Component_Function_1/NAND4_in[2] ), .A2(
        \SB4_10/Component_Function_1/NAND4_in[3] ), .A3(
        \SB4_10/Component_Function_1/NAND4_in[1] ), .A4(n2456), .ZN(n4877) );
  NAND4_X2 U5083 ( .A1(\SB2_2_9/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_9/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_2_9/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_2_9/Component_Function_2/NAND4_in[1] ), .ZN(
        \SB2_2_9/buf_output[2] ) );
  NAND4_X2 U5087 ( .A1(n3297), .A2(\SB1_3_30/Component_Function_2/NAND4_in[0] ), .A3(n5048), .A4(n6287), .ZN(\SB1_3_30/buf_output[2] ) );
  XOR2_X1 U5090 ( .A1(\MC_ARK_ARC_1_3/temp2[140] ), .A2(n4878), .Z(
        \MC_ARK_ARC_1_3/temp5[140] ) );
  XOR2_X1 U5091 ( .A1(\RI5[3][134] ), .A2(\RI5[3][140] ), .Z(n4878) );
  XOR2_X1 U5092 ( .A1(n4879), .A2(n191), .Z(Ciphertext[28]) );
  NAND4_X2 U5095 ( .A1(n3456), .A2(n4900), .A3(
        \SB4_27/Component_Function_4/NAND4_in[1] ), .A4(n2746), .ZN(n4879) );
  XOR2_X1 U5096 ( .A1(\MC_ARK_ARC_1_3/temp1[17] ), .A2(n4880), .Z(
        \MC_ARK_ARC_1_3/temp5[17] ) );
  XOR2_X1 U5097 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[155] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[179] ), .Z(n4880) );
  XOR2_X1 U5100 ( .A1(n4881), .A2(n159), .Z(Ciphertext[149]) );
  NAND4_X2 U5102 ( .A1(\SB4_7/Component_Function_5/NAND4_in[3] ), .A2(n6293), 
        .A3(\SB4_7/Component_Function_5/NAND4_in[1] ), .A4(
        \SB4_7/Component_Function_5/NAND4_in[0] ), .ZN(n4881) );
  XOR2_X1 U5103 ( .A1(n4883), .A2(n4882), .Z(\MC_ARK_ARC_1_3/temp5[182] ) );
  XOR2_X1 U5106 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[182] ), .A2(\RI5[3][128] ), 
        .Z(n4882) );
  XOR2_X1 U5109 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[152] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[176] ), .Z(n4883) );
  AND3_X1 U5110 ( .A1(\SB1_2_9/i0_0 ), .A2(\SB1_2_9/i0[9] ), .A3(
        \SB1_2_9/i0[8] ), .Z(n5883) );
  NAND2_X2 U5111 ( .A1(n6170), .A2(n4884), .ZN(\RI5[2][157] ) );
  AND2_X1 U5113 ( .A1(\SB2_2_9/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_9/Component_Function_1/NAND4_in[1] ), .Z(n4884) );
  XOR2_X1 U5115 ( .A1(\RI5[2][26] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[182] ), 
        .Z(n4885) );
  XOR2_X1 U5122 ( .A1(n4204), .A2(n4886), .Z(\MC_ARK_ARC_1_3/buf_output[93] )
         );
  XOR2_X1 U5124 ( .A1(\MC_ARK_ARC_1_3/temp4[93] ), .A2(n2547), .Z(n4886) );
  XOR2_X1 U5125 ( .A1(\MC_ARK_ARC_1_3/temp5[167] ), .A2(
        \MC_ARK_ARC_1_3/temp6[167] ), .Z(\MC_ARK_ARC_1_3/buf_output[167] ) );
  NAND4_X2 U5126 ( .A1(n826), .A2(\SB2_2_14/Component_Function_2/NAND4_in[0] ), 
        .A3(n3029), .A4(n4887), .ZN(\SB2_2_14/buf_output[2] ) );
  NAND3_X2 U5130 ( .A1(n5932), .A2(\SB2_2_14/i0_0 ), .A3(\SB2_2_14/i1_5 ), 
        .ZN(n4887) );
  XOR2_X1 U5131 ( .A1(n4888), .A2(\MC_ARK_ARC_1_2/temp6[46] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[46] ) );
  XOR2_X1 U5132 ( .A1(\MC_ARK_ARC_1_2/temp1[46] ), .A2(n4733), .Z(n4888) );
  XOR2_X1 U5133 ( .A1(n3874), .A2(n4889), .Z(n5619) );
  XOR2_X1 U5134 ( .A1(\RI5[2][11] ), .A2(\RI5[2][35] ), .Z(n4889) );
  XOR2_X1 U5135 ( .A1(\RI5[1][171] ), .A2(\RI5[1][165] ), .Z(
        \MC_ARK_ARC_1_1/temp1[171] ) );
  NAND4_X2 U5140 ( .A1(\SB1_2_3/Component_Function_5/NAND4_in[2] ), .A2(n4644), 
        .A3(n2933), .A4(n4890), .ZN(\SB1_2_3/buf_output[5] ) );
  NAND3_X2 U5142 ( .A1(\SB1_2_3/i0[6] ), .A2(\SB1_2_3/i0[10] ), .A3(
        \SB1_2_3/i0_0 ), .ZN(n4890) );
  NAND4_X2 U5144 ( .A1(\SB3_3/Component_Function_3/NAND4_in[0] ), .A2(n1799), 
        .A3(n4993), .A4(n5068), .ZN(\SB3_3/buf_output[3] ) );
  NAND3_X1 U5150 ( .A1(\SB4_1/i1_7 ), .A2(\SB4_1/i0[10] ), .A3(\SB4_1/i1[9] ), 
        .ZN(n4891) );
  NAND4_X2 U5151 ( .A1(\SB2_1_23/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_1_23/Component_Function_2/NAND4_in[2] ), .A3(n2223), .A4(n4892), 
        .ZN(\SB2_1_23/buf_output[2] ) );
  NAND3_X2 U5152 ( .A1(\SB2_1_23/i0[10] ), .A2(\SB2_1_23/i1_5 ), .A3(
        \SB2_1_23/i1[9] ), .ZN(n4892) );
  XOR2_X1 U5156 ( .A1(\MC_ARK_ARC_1_1/temp1[53] ), .A2(n4893), .Z(n1138) );
  XOR2_X1 U5158 ( .A1(\RI5[1][191] ), .A2(\RI5[1][23] ), .Z(n4893) );
  NAND4_X2 U5159 ( .A1(\SB2_2_23/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_23/Component_Function_3/NAND4_in[3] ), .A3(
        \SB2_2_23/Component_Function_3/NAND4_in[2] ), .A4(n5616), .ZN(
        \SB2_2_23/buf_output[3] ) );
  NAND4_X2 U5160 ( .A1(\SB1_3_29/Component_Function_1/NAND4_in[1] ), .A2(n1971), .A3(\SB1_3_29/Component_Function_1/NAND4_in[0] ), .A4(
        \SB1_3_29/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_3_29/buf_output[1] ) );
  XOR2_X1 U5161 ( .A1(\RI5[0][106] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[112] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[112] ) );
  NAND4_X2 U5162 ( .A1(\SB2_0_4/Component_Function_3/NAND4_in[3] ), .A2(
        \SB2_0_4/Component_Function_3/NAND4_in[2] ), .A3(n4970), .A4(n5141), 
        .ZN(\SB2_0_4/buf_output[3] ) );
  NAND3_X2 U5163 ( .A1(\SB2_2_21/i0[6] ), .A2(\SB2_2_21/i0[10] ), .A3(
        \SB2_2_21/i0_3 ), .ZN(\SB2_2_21/Component_Function_2/NAND4_in[1] ) );
  NAND4_X2 U5164 ( .A1(\SB1_0_18/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_0_18/Component_Function_2/NAND4_in[3] ), .A3(
        \SB1_0_18/Component_Function_2/NAND4_in[0] ), .A4(n1581), .ZN(
        \SB1_0_18/buf_output[2] ) );
  XOR2_X1 U5165 ( .A1(\RI5[2][63] ), .A2(\RI5[2][69] ), .Z(n2951) );
  NAND4_X2 U5167 ( .A1(\SB2_0_7/Component_Function_0/NAND4_in[1] ), .A2(n6011), 
        .A3(\SB2_0_7/Component_Function_0/NAND4_in[0] ), .A4(
        \SB2_0_7/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB2_0_7/buf_output[0] ) );
  NAND4_X2 U5168 ( .A1(\SB1_3_17/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_17/Component_Function_2/NAND4_in[2] ), .A3(n5144), .A4(n5937), 
        .ZN(\SB1_3_17/buf_output[2] ) );
  NAND4_X2 U5172 ( .A1(\SB2_1_12/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_12/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_12/Component_Function_1/NAND4_in[2] ), .A4(n4894), .ZN(
        \SB2_1_12/buf_output[1] ) );
  NAND3_X1 U5175 ( .A1(\SB2_1_12/i0_4 ), .A2(\SB2_1_12/i1_7 ), .A3(
        \SB2_1_12/i0[8] ), .ZN(n4894) );
  NAND3_X1 U5184 ( .A1(\SB1_3_20/i0[10] ), .A2(\SB1_3_20/i1[9] ), .A3(
        \SB1_3_20/i1_7 ), .ZN(\SB1_3_20/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U5186 ( .A1(\SB1_1_29/i0[10] ), .A2(\SB1_1_29/i0[6] ), .A3(
        \SB1_1_29/i0_0 ), .ZN(\SB1_1_29/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U5188 ( .A1(\MC_ARK_ARC_1_2/temp5[69] ), .A2(n5264), .Z(
        \MC_ARK_ARC_1_2/buf_output[69] ) );
  XOR2_X1 U5191 ( .A1(\RI5[0][137] ), .A2(\RI5[0][131] ), .Z(
        \MC_ARK_ARC_1_0/temp1[137] ) );
  XOR2_X1 U5192 ( .A1(\MC_ARK_ARC_1_2/temp6[191] ), .A2(n5543), .Z(
        \MC_ARK_ARC_1_2/buf_output[191] ) );
  NAND4_X2 U5193 ( .A1(n2540), .A2(\SB2_0_23/Component_Function_3/NAND4_in[0] ), .A3(n3618), .A4(\SB2_0_23/Component_Function_3/NAND4_in[2] ), .ZN(
        \SB2_0_23/buf_output[3] ) );
  NAND4_X2 U5194 ( .A1(\SB1_1_13/Component_Function_4/NAND4_in[0] ), .A2(n1328), .A3(n1004), .A4(n4895), .ZN(\SB1_1_13/buf_output[4] ) );
  NAND3_X1 U5195 ( .A1(\SB1_1_13/i0_4 ), .A2(\SB1_1_13/i1[9] ), .A3(
        \SB1_1_13/i1_5 ), .ZN(n4895) );
  XOR2_X1 U5197 ( .A1(n4896), .A2(n204), .Z(Ciphertext[182]) );
  NAND4_X2 U5198 ( .A1(n5193), .A2(n4350), .A3(n3809), .A4(n5160), .ZN(n4896)
         );
  CLKBUF_X4 U5205 ( .I(\SB2_0_0/buf_output[3] ), .Z(\RI5[0][9] ) );
  XOR2_X1 U5206 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[158] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[122] ), .Z(n5889) );
  NAND4_X2 U5207 ( .A1(\SB1_3_11/Component_Function_1/NAND4_in[2] ), .A2(n775), 
        .A3(n6368), .A4(\SB1_3_11/Component_Function_1/NAND4_in[1] ), .ZN(
        \SB1_3_11/buf_output[1] ) );
  NAND3_X1 U5208 ( .A1(\SB2_2_8/i0_3 ), .A2(\SB2_2_8/i0_4 ), .A3(
        \SB2_2_8/i0[10] ), .ZN(n1439) );
  XOR2_X1 U5209 ( .A1(\MC_ARK_ARC_1_3/temp5[152] ), .A2(n4897), .Z(
        \MC_ARK_ARC_1_3/buf_output[152] ) );
  XOR2_X1 U5211 ( .A1(\MC_ARK_ARC_1_3/temp4[152] ), .A2(
        \MC_ARK_ARC_1_3/temp3[152] ), .Z(n4897) );
  XOR2_X1 U5212 ( .A1(n4898), .A2(n117), .Z(Ciphertext[27]) );
  NAND4_X2 U5213 ( .A1(\SB4_27/Component_Function_3/NAND4_in[2] ), .A2(
        \SB4_27/Component_Function_3/NAND4_in[3] ), .A3(
        \SB4_27/Component_Function_3/NAND4_in[1] ), .A4(
        \SB4_27/Component_Function_3/NAND4_in[0] ), .ZN(n4898) );
  XOR2_X1 U5215 ( .A1(n4899), .A2(n199), .Z(Ciphertext[146]) );
  NAND4_X2 U5219 ( .A1(n1830), .A2(n5839), .A3(
        \SB4_7/Component_Function_2/NAND4_in[0] ), .A4(
        \SB4_7/Component_Function_2/NAND4_in[1] ), .ZN(n4899) );
  NAND3_X1 U5220 ( .A1(\SB4_27/i0_3 ), .A2(\SB4_27/i0[9] ), .A3(
        \SB4_27/i0[10] ), .ZN(n4900) );
  XOR2_X1 U5222 ( .A1(n4901), .A2(n236), .Z(Ciphertext[147]) );
  NAND4_X2 U5236 ( .A1(\SB4_7/Component_Function_3/NAND4_in[3] ), .A2(
        \SB4_7/Component_Function_3/NAND4_in[1] ), .A3(n3929), .A4(n3399), 
        .ZN(n4901) );
  NAND4_X2 U5237 ( .A1(n5353), .A2(\SB2_3_12/Component_Function_1/NAND4_in[1] ), .A3(\SB2_3_12/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_3_12/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_3_12/buf_output[1] ) );
  BUF_X4 U5239 ( .I(\SB2_1_30/buf_output[2] ), .Z(\RI5[1][26] ) );
  XOR2_X1 U5240 ( .A1(n5319), .A2(n4902), .Z(\MC_ARK_ARC_1_0/buf_output[138] )
         );
  XOR2_X1 U5241 ( .A1(n5239), .A2(\MC_ARK_ARC_1_0/temp4[138] ), .Z(n4902) );
  XOR2_X1 U5242 ( .A1(\MC_ARK_ARC_1_0/temp1[94] ), .A2(n4903), .Z(
        \MC_ARK_ARC_1_0/temp5[94] ) );
  XOR2_X1 U5244 ( .A1(\RI5[0][64] ), .A2(\RI5[0][40] ), .Z(n4903) );
  XOR2_X1 U5245 ( .A1(\MC_ARK_ARC_1_3/temp4[183] ), .A2(n4904), .Z(n6236) );
  XOR2_X1 U5246 ( .A1(\RI5[3][93] ), .A2(\SB2_3_24/buf_output[3] ), .Z(n4904)
         );
  XOR2_X1 U5247 ( .A1(\MC_ARK_ARC_1_3/temp5[95] ), .A2(n4905), .Z(
        \MC_ARK_ARC_1_3/buf_output[95] ) );
  XOR2_X1 U5248 ( .A1(\MC_ARK_ARC_1_3/temp4[95] ), .A2(
        \MC_ARK_ARC_1_3/temp3[95] ), .Z(n4905) );
  NAND3_X2 U5249 ( .A1(\SB1_3_15/i0[9] ), .A2(\SB1_3_15/i0_3 ), .A3(
        \SB1_3_15/i0[8] ), .ZN(n4906) );
  NAND3_X1 U5250 ( .A1(\SB2_2_5/i0[10] ), .A2(\SB2_2_5/i0_3 ), .A3(
        \SB2_2_5/i0_4 ), .ZN(\SB2_2_5/Component_Function_0/NAND4_in[2] ) );
  INV_X2 U5251 ( .I(\SB1_1_0/buf_output[2] ), .ZN(\SB2_1_29/i1[9] ) );
  NAND4_X2 U5257 ( .A1(n1318), .A2(\SB1_1_0/Component_Function_2/NAND4_in[3] ), 
        .A3(\SB1_1_0/Component_Function_2/NAND4_in[0] ), .A4(n1577), .ZN(
        \SB1_1_0/buf_output[2] ) );
  XOR2_X1 U5258 ( .A1(\SB2_1_1/buf_output[3] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[159] ), .Z(n1433) );
  INV_X1 U5259 ( .I(\SB3_13/buf_output[1] ), .ZN(\SB4_9/i1_7 ) );
  NAND4_X2 U5260 ( .A1(\SB3_13/Component_Function_1/NAND4_in[3] ), .A2(
        \SB3_13/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_13/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_13/Component_Function_1/NAND4_in[0] ), .ZN(\SB3_13/buf_output[1] ) );
  XOR2_X1 U5261 ( .A1(\RI5[2][110] ), .A2(\SB2_2_10/buf_output[2] ), .Z(n5076)
         );
  NAND3_X1 U5268 ( .A1(\SB1_1_8/i0_4 ), .A2(\SB1_1_8/i1[9] ), .A3(n3270), .ZN(
        n4907) );
  XOR2_X1 U5271 ( .A1(n4908), .A2(n83), .Z(Ciphertext[191]) );
  NAND4_X2 U5284 ( .A1(\SB4_0/Component_Function_5/NAND4_in[1] ), .A2(
        \SB4_0/Component_Function_5/NAND4_in[3] ), .A3(
        \SB4_0/Component_Function_5/NAND4_in[2] ), .A4(
        \SB4_0/Component_Function_5/NAND4_in[0] ), .ZN(n4908) );
  XOR2_X1 U5285 ( .A1(n2945), .A2(n4909), .Z(\MC_ARK_ARC_1_1/temp5[129] ) );
  XOR2_X1 U5287 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[123] ), .A2(
        \SB2_1_12/buf_output[3] ), .Z(n4909) );
  NAND4_X2 U5291 ( .A1(\SB2_0_12/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_12/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_0_12/Component_Function_3/NAND4_in[1] ), .A4(n4910), .ZN(
        \SB2_0_12/buf_output[3] ) );
  NAND3_X2 U5292 ( .A1(\SB2_2_7/i0_0 ), .A2(\SB2_2_7/i0[9] ), .A3(
        \SB2_2_7/i0[8] ), .ZN(\SB2_2_7/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U5295 ( .A1(\SB3_8/i0_0 ), .A2(\SB3_8/i0_3 ), .A3(\SB3_8/i0[7] ), 
        .ZN(n4052) );
  XOR2_X1 U5297 ( .A1(n4911), .A2(n53), .Z(Ciphertext[161]) );
  NAND4_X2 U5298 ( .A1(n2914), .A2(\SB4_5/Component_Function_5/NAND4_in[1] ), 
        .A3(\SB4_5/Component_Function_5/NAND4_in[0] ), .A4(
        \SB4_5/Component_Function_5/NAND4_in[2] ), .ZN(n4911) );
  XOR2_X1 U5299 ( .A1(n4912), .A2(n154), .Z(Ciphertext[139]) );
  NAND4_X2 U5302 ( .A1(\SB4_8/Component_Function_1/NAND4_in[3] ), .A2(
        \SB4_8/Component_Function_1/NAND4_in[2] ), .A3(
        \SB4_8/Component_Function_1/NAND4_in[1] ), .A4(n768), .ZN(n4912) );
  XOR2_X1 U5304 ( .A1(n4913), .A2(n196), .Z(Ciphertext[140]) );
  NAND4_X2 U5306 ( .A1(\SB4_8/Component_Function_2/NAND4_in[0] ), .A2(
        \SB4_8/Component_Function_2/NAND4_in[3] ), .A3(n6212), .A4(
        \SB4_8/Component_Function_2/NAND4_in[2] ), .ZN(n4913) );
  XOR2_X1 U5309 ( .A1(n4914), .A2(n239), .Z(Ciphertext[142]) );
  NAND4_X2 U5311 ( .A1(\SB4_8/Component_Function_4/NAND4_in[3] ), .A2(n3175), 
        .A3(n4018), .A4(n629), .ZN(n4914) );
  XOR2_X1 U5315 ( .A1(n4916), .A2(n4915), .Z(n5743) );
  XOR2_X1 U5316 ( .A1(\SB2_3_7/buf_output[2] ), .A2(n233), .Z(n4915) );
  XOR2_X1 U5322 ( .A1(\RI5[3][98] ), .A2(\RI5[3][128] ), .Z(n4916) );
  NAND4_X2 U5323 ( .A1(\SB3_6/Component_Function_4/NAND4_in[0] ), .A2(n2762), 
        .A3(n785), .A4(n4917), .ZN(\SB3_6/buf_output[4] ) );
  NAND3_X1 U5324 ( .A1(\SB3_6/i0_0 ), .A2(\SB3_6/i1_7 ), .A3(\SB3_6/i3[0] ), 
        .ZN(n4917) );
  NAND3_X2 U5326 ( .A1(\SB2_2_31/i0[10] ), .A2(\SB2_2_31/i1_5 ), .A3(
        \SB2_2_31/i1[9] ), .ZN(\SB2_2_31/Component_Function_2/NAND4_in[0] ) );
  INV_X2 U5333 ( .I(\SB1_3_29/buf_output[2] ), .ZN(\SB2_3_26/i1[9] ) );
  NAND4_X2 U5336 ( .A1(\SB1_3_29/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_29/Component_Function_2/NAND4_in[2] ), .A3(n5906), .A4(n2307), 
        .ZN(\SB1_3_29/buf_output[2] ) );
  NAND4_X2 U5337 ( .A1(\SB2_3_17/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_17/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_17/Component_Function_3/NAND4_in[3] ), .A4(n4918), .ZN(
        \SB2_3_17/buf_output[3] ) );
  NAND3_X2 U5338 ( .A1(\SB2_3_17/i0[10] ), .A2(\SB2_3_17/i1_7 ), .A3(
        \SB2_3_17/i1[9] ), .ZN(n4918) );
  NAND3_X1 U5339 ( .A1(\RI3[0][88] ), .A2(\SB2_0_17/i1[9] ), .A3(
        \SB2_0_17/i1_5 ), .ZN(\SB2_0_17/Component_Function_4/NAND4_in[3] ) );
  NAND2_X1 U5340 ( .A1(n1021), .A2(\SB3_1/Component_Function_3/NAND4_in[1] ), 
        .ZN(n5559) );
  XOR2_X1 U5341 ( .A1(\MC_ARK_ARC_1_3/temp2[159] ), .A2(n4125), .Z(
        \MC_ARK_ARC_1_3/temp5[159] ) );
  NAND4_X2 U5344 ( .A1(n1639), .A2(n2526), .A3(
        \SB1_2_30/Component_Function_4/NAND4_in[0] ), .A4(
        \SB1_2_30/Component_Function_4/NAND4_in[1] ), .ZN(\SB2_2_29/i0_4 ) );
  NAND4_X2 U5346 ( .A1(\SB2_0_0/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_0_0/Component_Function_0/NAND4_in[2] ), .A3(n760), .A4(
        \SB2_0_0/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_0_0/buf_output[0] ) );
  XOR2_X1 U5347 ( .A1(\RI5[0][24] ), .A2(\RI5[0][0] ), .Z(n1826) );
  XOR2_X1 U5348 ( .A1(\RI5[1][65] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[101] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[191] ) );
  NAND4_X2 U5356 ( .A1(\SB3_16/Component_Function_2/NAND4_in[1] ), .A2(n5729), 
        .A3(n6246), .A4(n6089), .ZN(\SB3_16/buf_output[2] ) );
  NAND4_X2 U5359 ( .A1(\SB1_3_8/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_3_8/Component_Function_5/NAND4_in[1] ), .A3(n6304), .A4(
        \SB1_3_8/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_8/buf_output[5] ) );
  XOR2_X1 U5362 ( .A1(\MC_ARK_ARC_1_3/temp5[162] ), .A2(n4919), .Z(
        \MC_ARK_ARC_1_3/buf_output[162] ) );
  XOR2_X1 U5364 ( .A1(\MC_ARK_ARC_1_3/temp4[162] ), .A2(n5156), .Z(n4919) );
  XOR2_X1 U5365 ( .A1(n4920), .A2(n241), .Z(Ciphertext[166]) );
  NAND4_X2 U5368 ( .A1(\SB4_4/Component_Function_4/NAND4_in[0] ), .A2(n3471), 
        .A3(n3180), .A4(\SB4_4/Component_Function_4/NAND4_in[1] ), .ZN(n4920)
         );
  XOR2_X1 U5369 ( .A1(\RI5[3][108] ), .A2(\RI5[3][102] ), .Z(
        \MC_ARK_ARC_1_3/temp1[108] ) );
  NAND2_X2 U5370 ( .A1(n2285), .A2(n5755), .ZN(\RI5[3][102] ) );
  NAND3_X1 U5371 ( .A1(\SB2_3_23/i0[9] ), .A2(\SB2_3_23/i0_3 ), .A3(
        \SB2_3_23/i0[10] ), .ZN(\SB2_3_23/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X2 U5372 ( .A1(\SB2_2_10/i0[10] ), .A2(\SB2_2_10/i0_3 ), .A3(
        \SB2_2_10/i0[9] ), .ZN(n6137) );
  NAND3_X2 U5374 ( .A1(\SB1_1_23/i0_3 ), .A2(\SB1_1_23/i0_4 ), .A3(
        \SB1_1_23/i1[9] ), .ZN(n1337) );
  NAND4_X2 U5378 ( .A1(\SB2_2_9/Component_Function_5/NAND4_in[2] ), .A2(n4935), 
        .A3(\SB2_2_9/Component_Function_5/NAND4_in[0] ), .A4(n4921), .ZN(
        \SB2_2_9/buf_output[5] ) );
  NAND3_X2 U5381 ( .A1(\SB2_2_9/i0[10] ), .A2(\SB2_2_9/i0_0 ), .A3(
        \SB2_2_9/i0[6] ), .ZN(n4921) );
  INV_X2 U5382 ( .I(\SB2_2_10/i0[7] ), .ZN(n581) );
  NAND3_X2 U5384 ( .A1(\SB1_2_15/i0_4 ), .A2(\SB1_2_15/i0[6] ), .A3(
        \SB1_2_15/i0[9] ), .ZN(n1849) );
  NAND4_X2 U5385 ( .A1(\SB4_4/Component_Function_2/NAND4_in[3] ), .A2(n6490), 
        .A3(n4931), .A4(n4922), .ZN(n5332) );
  NAND3_X1 U5386 ( .A1(\SB4_4/i0_3 ), .A2(\SB4_4/i0[9] ), .A3(\SB4_4/i0[8] ), 
        .ZN(n4922) );
  NAND3_X1 U5390 ( .A1(\SB2_0_0/i0[8] ), .A2(\SB2_0_0/i3[0] ), .A3(
        \SB2_0_0/i1_5 ), .ZN(\SB2_0_0/Component_Function_3/NAND4_in[3] ) );
  NAND4_X2 U5393 ( .A1(n3861), .A2(n2680), .A3(
        \SB4_16/Component_Function_4/NAND4_in[0] ), .A4(n4923), .ZN(n5533) );
  NAND3_X1 U5403 ( .A1(\SB4_16/i0[9] ), .A2(\SB4_16/i0[10] ), .A3(
        \SB4_16/i0_3 ), .ZN(n4923) );
  NAND3_X2 U5408 ( .A1(\SB4_2/i0[10] ), .A2(\SB4_2/i1_7 ), .A3(\SB4_2/i1[9] ), 
        .ZN(\SB4_2/Component_Function_3/NAND4_in[2] ) );
  XOR2_X1 U5409 ( .A1(\MC_ARK_ARC_1_1/temp1[38] ), .A2(n4924), .Z(
        \MC_ARK_ARC_1_1/temp5[38] ) );
  XOR2_X1 U5413 ( .A1(\RI5[1][8] ), .A2(\RI5[1][176] ), .Z(n4924) );
  XOR2_X1 U5414 ( .A1(n4925), .A2(n229), .Z(Ciphertext[100]) );
  NAND4_X2 U5415 ( .A1(n873), .A2(\SB4_15/Component_Function_4/NAND4_in[3] ), 
        .A3(n5443), .A4(n1235), .ZN(n4925) );
  NAND4_X2 U5416 ( .A1(\SB2_1_1/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_1_1/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_1/Component_Function_0/NAND4_in[0] ), .A4(n4926), .ZN(
        \SB2_1_1/buf_output[0] ) );
  NAND3_X2 U5420 ( .A1(\SB2_1_1/i0[10] ), .A2(\SB2_1_1/i0_4 ), .A3(
        \SB2_1_1/i0_3 ), .ZN(n4926) );
  NAND4_X2 U5421 ( .A1(\SB2_2_27/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_2_27/Component_Function_0/NAND4_in[0] ), .A3(
        \SB2_2_27/Component_Function_0/NAND4_in[2] ), .A4(n4927), .ZN(
        \SB2_2_27/buf_output[0] ) );
  NAND3_X1 U5423 ( .A1(\SB2_2_27/i0[6] ), .A2(\SB2_2_27/i0[8] ), .A3(n6073), 
        .ZN(n4927) );
  XOR2_X1 U5424 ( .A1(n4928), .A2(\MC_ARK_ARC_1_0/temp5[109] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[109] ) );
  XOR2_X1 U5428 ( .A1(\MC_ARK_ARC_1_0/temp3[109] ), .A2(
        \MC_ARK_ARC_1_0/temp4[109] ), .Z(n4928) );
  NAND4_X2 U5429 ( .A1(\SB2_3_25/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_3_25/Component_Function_2/NAND4_in[3] ), .A3(n4929), .A4(n4975), 
        .ZN(\SB2_3_25/buf_output[2] ) );
  XOR2_X1 U5435 ( .A1(\MC_ARK_ARC_1_1/temp1[174] ), .A2(n4930), .Z(
        \MC_ARK_ARC_1_1/temp5[174] ) );
  XOR2_X1 U5436 ( .A1(\RI5[1][120] ), .A2(\RI5[1][144] ), .Z(n4930) );
  NAND3_X1 U5439 ( .A1(\SB4_4/i0[10] ), .A2(n3655), .A3(\SB4_4/i1_5 ), .ZN(
        n4931) );
  BUF_X4 U5441 ( .I(n418), .Z(\SB1_0_18/i0_3 ) );
  XOR2_X1 U5442 ( .A1(n4932), .A2(n243), .Z(Ciphertext[34]) );
  NAND4_X2 U5443 ( .A1(n5609), .A2(n4742), .A3(
        \SB4_26/Component_Function_4/NAND4_in[1] ), .A4(n2372), .ZN(n4932) );
  NAND4_X2 U5447 ( .A1(\SB2_2_1/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_1/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_2_1/Component_Function_2/NAND4_in[1] ), .A4(n4933), .ZN(
        \SB2_2_1/buf_output[2] ) );
  NAND3_X2 U5448 ( .A1(\SB2_2_1/i0_4 ), .A2(\SB2_2_1/i0_0 ), .A3(
        \SB2_2_1/i1_5 ), .ZN(n4933) );
  NAND3_X2 U5449 ( .A1(\SB1_1_8/i0[9] ), .A2(\SB1_1_8/i0[6] ), .A3(
        \SB1_1_8/i0_4 ), .ZN(\SB1_1_8/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U5450 ( .A1(\SB2_2_4/i0_3 ), .A2(\SB2_2_4/i0_4 ), .A3(
        \SB2_2_4/i0[10] ), .ZN(\SB2_2_4/Component_Function_0/NAND4_in[2] ) );
  NAND4_X2 U5451 ( .A1(\SB2_3_9/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_3_9/Component_Function_2/NAND4_in[0] ), .A3(n5114), .A4(n5878), 
        .ZN(\SB2_3_9/buf_output[2] ) );
  NAND4_X2 U5455 ( .A1(\SB1_3_22/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_22/Component_Function_5/NAND4_in[3] ), .A3(n5033), .A4(
        \SB1_3_22/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_22/buf_output[5] ) );
  XOR2_X1 U5458 ( .A1(\MC_ARK_ARC_1_1/temp1[144] ), .A2(n6234), .Z(
        \MC_ARK_ARC_1_1/temp5[144] ) );
  XOR2_X1 U5459 ( .A1(\RI5[2][75] ), .A2(\RI5[2][111] ), .Z(n3068) );
  NAND3_X1 U5460 ( .A1(\SB2_0_10/i0[10] ), .A2(\SB2_0_10/i0[6] ), .A3(
        \SB2_0_10/i0_0 ), .ZN(\SB2_0_10/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U5470 ( .A1(\SB3_31/i0_0 ), .A2(\SB3_31/i3[0] ), .A3(\SB3_31/i1_7 ), 
        .ZN(\SB3_31/Component_Function_4/NAND4_in[1] ) );
  NAND3_X2 U5473 ( .A1(\SB2_2_19/i0_4 ), .A2(\SB2_2_19/i0_0 ), .A3(
        \SB2_2_19/i1_5 ), .ZN(n5910) );
  NAND3_X2 U5474 ( .A1(\SB1_2_7/i0[6] ), .A2(\SB1_2_7/i0[9] ), .A3(
        \SB1_2_7/i0_4 ), .ZN(n5180) );
  NAND4_X2 U5475 ( .A1(\SB2_1_27/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_1_27/Component_Function_4/NAND4_in[3] ), .A3(n5179), .A4(
        \SB2_1_27/Component_Function_4/NAND4_in[0] ), .ZN(
        \SB2_1_27/buf_output[4] ) );
  NAND4_X2 U5477 ( .A1(n2862), .A2(n5000), .A3(
        \SB1_2_21/Component_Function_5/NAND4_in[1] ), .A4(
        \SB1_2_21/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_2_21/buf_output[5] ) );
  NAND4_X2 U5478 ( .A1(n3954), .A2(n4715), .A3(n5577), .A4(n4560), .ZN(
        \SB2_3_22/buf_output[5] ) );
  NAND3_X1 U5480 ( .A1(\SB1_3_3/i0_3 ), .A2(\SB1_3_3/i0[10] ), .A3(
        \SB1_3_3/i0[9] ), .ZN(\SB1_3_3/Component_Function_4/NAND4_in[2] ) );
  NAND4_X2 U5481 ( .A1(n5485), .A2(\SB2_1_15/Component_Function_5/NAND4_in[1] ), .A3(\SB2_1_15/Component_Function_5/NAND4_in[0] ), .A4(n4934), .ZN(
        \SB2_1_15/buf_output[5] ) );
  NAND3_X2 U5482 ( .A1(\SB2_1_15/i0[9] ), .A2(\SB2_1_15/i0_4 ), .A3(
        \SB2_1_15/i0[6] ), .ZN(n4934) );
  NAND3_X2 U5483 ( .A1(\SB2_2_9/i0[9] ), .A2(\SB2_2_9/i0_4 ), .A3(
        \SB2_2_9/i0[6] ), .ZN(n4935) );
  XOR2_X1 U5484 ( .A1(\MC_ARK_ARC_1_1/temp4[161] ), .A2(n4936), .Z(n4960) );
  XOR2_X1 U5485 ( .A1(\RI5[1][71] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[35] ), 
        .Z(n4936) );
  XOR2_X1 U5486 ( .A1(n4938), .A2(n4937), .Z(\MC_ARK_ARC_1_1/temp6[75] ) );
  XOR2_X1 U5487 ( .A1(\RI5[1][177] ), .A2(n211), .Z(n4937) );
  XOR2_X1 U5491 ( .A1(\RI5[1][141] ), .A2(\RI5[1][111] ), .Z(n4938) );
  NAND3_X1 U5496 ( .A1(\SB4_30/i0[10] ), .A2(n4751), .A3(n5525), .ZN(
        \SB4_30/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U5503 ( .A1(\SB1_3_9/i1_7 ), .A2(\SB1_3_9/i1[9] ), .A3(n5502), .ZN(
        n4939) );
  NAND3_X1 U5505 ( .A1(\SB1_3_22/buf_output[4] ), .A2(\SB2_3_21/i0[8] ), .A3(
        \SB2_3_21/i1_7 ), .ZN(n3191) );
  NAND2_X2 U5507 ( .A1(n2718), .A2(n3329), .ZN(\SB1_3_22/buf_output[4] ) );
  NAND4_X2 U5508 ( .A1(\SB1_1_16/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_1_16/Component_Function_5/NAND4_in[1] ), .A3(n2713), .A4(
        \SB1_1_16/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_16/buf_output[5] ) );
  NAND4_X2 U5510 ( .A1(\SB3_23/Component_Function_1/NAND4_in[1] ), .A2(n3896), 
        .A3(n6112), .A4(n4940), .ZN(\SB3_23/buf_output[1] ) );
  NAND3_X1 U5511 ( .A1(\SB3_23/i0[9] ), .A2(\SB3_23/i0[6] ), .A3(\SB3_23/i1_5 ), .ZN(n4940) );
  XOR2_X1 U5513 ( .A1(\MC_ARK_ARC_1_0/temp2[81] ), .A2(n4941), .Z(n2170) );
  XOR2_X1 U5521 ( .A1(\RI5[0][75] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[81] ), 
        .Z(n4941) );
  XOR2_X1 U5524 ( .A1(n4942), .A2(n98), .Z(Ciphertext[77]) );
  NAND4_X2 U5526 ( .A1(\SB4_19/Component_Function_5/NAND4_in[1] ), .A2(
        \SB4_19/Component_Function_5/NAND4_in[3] ), .A3(
        \SB4_19/Component_Function_5/NAND4_in[2] ), .A4(
        \SB4_19/Component_Function_5/NAND4_in[0] ), .ZN(n4942) );
  XOR2_X1 U5527 ( .A1(\SB2_0_18/buf_output[3] ), .A2(\RI5[0][87] ), .Z(n5467)
         );
  XOR2_X1 U5529 ( .A1(n4943), .A2(\MC_ARK_ARC_1_1/temp2[161] ), .Z(n4959) );
  XOR2_X1 U5537 ( .A1(\RI5[1][161] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[155] ), 
        .Z(n4943) );
  NOR2_X2 U5538 ( .A1(n4945), .A2(n4944), .ZN(n5515) );
  NAND2_X1 U5539 ( .A1(\SB1_2_14/Component_Function_2/NAND4_in[2] ), .A2(n1225), .ZN(n4944) );
  NAND3_X2 U5540 ( .A1(\SB1_2_14/i0_0 ), .A2(\SB1_2_14/i0_4 ), .A3(
        \SB1_2_14/i1_5 ), .ZN(n1225) );
  NAND2_X1 U5543 ( .A1(\SB1_2_14/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_14/Component_Function_2/NAND4_in[1] ), .ZN(n4945) );
  XOR2_X1 U5545 ( .A1(n4947), .A2(n4946), .Z(\MC_ARK_ARC_1_1/temp5[124] ) );
  XOR2_X1 U5547 ( .A1(\RI5[1][124] ), .A2(\RI5[1][94] ), .Z(n4946) );
  XOR2_X1 U5548 ( .A1(\RI5[1][118] ), .A2(\RI5[1][70] ), .Z(n4947) );
  XOR2_X1 U5553 ( .A1(n4948), .A2(n210), .Z(Ciphertext[135]) );
  NAND4_X2 U5555 ( .A1(n4051), .A2(\SB4_9/Component_Function_3/NAND4_in[3] ), 
        .A3(n3922), .A4(n6130), .ZN(n4948) );
  XOR2_X1 U5556 ( .A1(\MC_ARK_ARC_1_2/temp4[45] ), .A2(n3880), .Z(
        \MC_ARK_ARC_1_2/temp6[45] ) );
  XOR2_X1 U5558 ( .A1(n4949), .A2(n220), .Z(Ciphertext[136]) );
  NAND4_X2 U5560 ( .A1(n3953), .A2(\SB4_9/Component_Function_4/NAND4_in[3] ), 
        .A3(n6381), .A4(n4558), .ZN(n4949) );
  INV_X1 U5562 ( .I(\SB3_11/buf_output[3] ), .ZN(\SB4_9/i0[8] ) );
  NAND4_X2 U5564 ( .A1(\SB3_11/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_11/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_11/Component_Function_3/NAND4_in[3] ), .A4(n6530), .ZN(
        \SB3_11/buf_output[3] ) );
  NAND3_X1 U5565 ( .A1(\SB4_1/i0_0 ), .A2(\SB4_1/i0_3 ), .A3(\SB4_1/i0[7] ), 
        .ZN(\SB4_1/Component_Function_0/NAND4_in[3] ) );
  NAND3_X2 U5570 ( .A1(\SB1_1_5/i0[6] ), .A2(\SB1_1_5/i0_3 ), .A3(
        \SB1_1_5/i0[10] ), .ZN(\SB1_1_5/Component_Function_2/NAND4_in[1] ) );
  XOR2_X1 U5571 ( .A1(n3577), .A2(n4743), .Z(\MC_ARK_ARC_1_2/buf_output[159] )
         );
  NAND4_X2 U5575 ( .A1(\SB2_0_22/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_22/Component_Function_2/NAND4_in[1] ), .A3(n5976), .A4(
        \SB2_0_22/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB2_0_22/buf_output[2] ) );
  XOR2_X1 U5576 ( .A1(\RI5[2][69] ), .A2(\RI5[2][33] ), .Z(
        \MC_ARK_ARC_1_2/temp3[159] ) );
  NAND3_X2 U5579 ( .A1(\SB1_1_9/i0[10] ), .A2(\SB1_1_9/i0[6] ), .A3(
        \SB1_1_9/i0_0 ), .ZN(\SB1_1_9/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U5580 ( .A1(\SB1_1_14/i0[10] ), .A2(\SB1_1_14/i1[9] ), .A3(
        \SB1_1_14/i1_7 ), .ZN(n3698) );
  NAND3_X2 U5581 ( .A1(\SB2_0_17/i0_3 ), .A2(\SB2_0_17/i0[9] ), .A3(
        \SB2_0_17/i0[8] ), .ZN(\SB2_0_17/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 U5583 ( .A1(\SB3_4/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_4/Component_Function_2/NAND4_in[1] ), .A3(n5098), .A4(
        \SB3_4/Component_Function_2/NAND4_in[3] ), .ZN(\SB3_4/buf_output[2] )
         );
  NAND4_X2 U5584 ( .A1(\SB1_2_31/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_2_31/Component_Function_2/NAND4_in[3] ), .A3(n5391), .A4(
        \SB1_2_31/Component_Function_2/NAND4_in[0] ), .ZN(
        \SB1_2_31/buf_output[2] ) );
  NAND3_X2 U5587 ( .A1(\SB1_3_18/i0_3 ), .A2(\SB1_3_18/i0_4 ), .A3(
        \SB1_3_18/i1[9] ), .ZN(n3754) );
  NAND4_X2 U5591 ( .A1(\SB1_0_23/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_0_23/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_23/Component_Function_0/NAND4_in[0] ), .A4(n4950), .ZN(
        \SB1_0_23/buf_output[0] ) );
  NAND3_X2 U5594 ( .A1(\SB1_0_23/i0[10] ), .A2(\SB1_0_23/i0_4 ), .A3(
        \SB1_0_23/i0_3 ), .ZN(n4950) );
  NAND2_X2 U5595 ( .A1(n2710), .A2(n6502), .ZN(\RI3[0][183] ) );
  NAND3_X1 U5598 ( .A1(\SB1_0_3/i0_0 ), .A2(\SB1_0_3/i0_4 ), .A3(
        \SB1_0_3/i0_3 ), .ZN(\SB1_0_3/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U5600 ( .A1(n4951), .A2(\MC_ARK_ARC_1_0/temp6[63] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[63] ) );
  XOR2_X1 U5602 ( .A1(n5399), .A2(\MC_ARK_ARC_1_0/temp1[63] ), .Z(n4951) );
  NAND3_X2 U5605 ( .A1(\SB3_4/i0[9] ), .A2(\SB3_4/i0_3 ), .A3(\SB3_4/i0[8] ), 
        .ZN(n5098) );
  NAND4_X2 U5608 ( .A1(\SB1_2_31/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_31/Component_Function_5/NAND4_in[2] ), .A3(n1444), .A4(n4271), 
        .ZN(\SB1_2_31/buf_output[5] ) );
  XOR2_X1 U5609 ( .A1(\MC_ARK_ARC_1_0/temp2[15] ), .A2(n4952), .Z(
        \MC_ARK_ARC_1_0/temp5[15] ) );
  XOR2_X1 U5611 ( .A1(\SB2_0_0/buf_output[3] ), .A2(\RI5[0][15] ), .Z(n4952)
         );
  NAND3_X1 U5613 ( .A1(\SB4_1/i0_0 ), .A2(\SB4_1/i0_4 ), .A3(\SB4_1/i1_5 ), 
        .ZN(n4350) );
  NAND4_X2 U5614 ( .A1(\SB2_3_24/Component_Function_0/NAND4_in[3] ), .A2(n2312), .A3(\SB2_3_24/Component_Function_0/NAND4_in[0] ), .A4(n4953), .ZN(
        \SB2_3_24/buf_output[0] ) );
  NAND3_X1 U5617 ( .A1(\SB2_3_24/i0_3 ), .A2(\SB2_3_24/i0_4 ), .A3(
        \SB1_3_26/buf_output[3] ), .ZN(n4953) );
  NAND2_X1 U5619 ( .A1(\SB4_1/i0[9] ), .A2(\SB4_1/i0[10] ), .ZN(n4954) );
  NOR2_X2 U5624 ( .A1(n4956), .A2(n4955), .ZN(n1389) );
  NAND2_X1 U5626 ( .A1(\SB3_30/Component_Function_2/NAND4_in[2] ), .A2(
        \SB3_30/Component_Function_2/NAND4_in[1] ), .ZN(n4955) );
  NAND2_X1 U5628 ( .A1(\SB3_30/Component_Function_2/NAND4_in[0] ), .A2(n1669), 
        .ZN(n4956) );
  NAND3_X2 U5629 ( .A1(\SB3_30/i0_4 ), .A2(\SB3_30/i0_0 ), .A3(\SB3_30/i1_5 ), 
        .ZN(n1669) );
  INV_X4 U5631 ( .I(\RI1[4][154] ), .ZN(\SB3_6/i0[7] ) );
  XOR2_X1 U5632 ( .A1(n4958), .A2(n4957), .Z(n1962) );
  XOR2_X1 U5633 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[110] ), .A2(n98), .Z(n4957) );
  XOR2_X1 U5635 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[74] ), .A2(\RI5[1][44] ), 
        .Z(n4958) );
  INV_X2 U5637 ( .I(\SB1_3_1/buf_output[2] ), .ZN(\SB2_3_30/i1[9] ) );
  NAND4_X2 U5638 ( .A1(\SB1_3_1/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_1/Component_Function_2/NAND4_in[2] ), .A3(
        \SB1_3_1/Component_Function_2/NAND4_in[1] ), .A4(n4286), .ZN(
        \SB1_3_1/buf_output[2] ) );
  XOR2_X1 U5643 ( .A1(n4960), .A2(n4959), .Z(\MC_ARK_ARC_1_1/buf_output[161] )
         );
  XOR2_X1 U5649 ( .A1(\MC_ARK_ARC_1_3/temp2[191] ), .A2(n4961), .Z(n6305) );
  XOR2_X1 U5650 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[191] ), .A2(\RI5[3][185] ), 
        .Z(n4961) );
  NAND3_X1 U5652 ( .A1(\SB2_3_2/i0_3 ), .A2(\SB2_3_2/i1_7 ), .A3(n5491), .ZN(
        \SB2_3_2/Component_Function_1/NAND4_in[1] ) );
  NOR2_X2 U5653 ( .A1(n4963), .A2(n4962), .ZN(n5491) );
  NAND2_X1 U5654 ( .A1(n5647), .A2(n1685), .ZN(n4963) );
  NAND3_X2 U5657 ( .A1(n4964), .A2(\SB2_1_9/Component_Function_1/NAND4_in[3] ), 
        .A3(\SB2_1_9/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_1_9/buf_output[1] ) );
  OAI21_X2 U5660 ( .A1(n4759), .A2(\SB2_1_9/i1[9] ), .B(\SB2_1_9/i0_3 ), .ZN(
        n4964) );
  INV_X1 U5661 ( .I(\SB1_0_29/buf_output[5] ), .ZN(\SB2_0_29/i1_5 ) );
  NAND4_X2 U5662 ( .A1(\SB1_0_29/Component_Function_5/NAND4_in[2] ), .A2(n1109), .A3(\SB1_0_29/Component_Function_5/NAND4_in[0] ), .A4(n5795), .ZN(
        \SB1_0_29/buf_output[5] ) );
  XOR2_X1 U5663 ( .A1(\RI5[0][188] ), .A2(\RI5[0][32] ), .Z(
        \MC_ARK_ARC_1_0/temp3[122] ) );
  NAND4_X2 U5664 ( .A1(\SB2_1_20/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_20/Component_Function_2/NAND4_in[3] ), .A3(
        \SB2_1_20/Component_Function_2/NAND4_in[2] ), .A4(n4965), .ZN(
        \SB2_1_20/buf_output[2] ) );
  NAND3_X2 U5665 ( .A1(\SB2_1_20/i0[10] ), .A2(\SB2_1_20/i0_3 ), .A3(
        \SB2_1_20/i0[6] ), .ZN(n4965) );
  NAND4_X2 U5669 ( .A1(\SB3_31/Component_Function_4/NAND4_in[2] ), .A2(
        \SB3_31/Component_Function_4/NAND4_in[1] ), .A3(
        \SB3_31/Component_Function_4/NAND4_in[3] ), .A4(n4966), .ZN(
        \SB3_31/buf_output[4] ) );
  XOR2_X1 U5671 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[74] ), .A2(
        \SB2_3_21/buf_output[2] ), .Z(n5776) );
  INV_X1 U5674 ( .I(\SB3_4/buf_output[5] ), .ZN(\SB4_4/i1_5 ) );
  NAND4_X2 U5676 ( .A1(\SB3_4/Component_Function_5/NAND4_in[1] ), .A2(
        \SB3_4/Component_Function_5/NAND4_in[2] ), .A3(n1863), .A4(n3475), 
        .ZN(\SB3_4/buf_output[5] ) );
  INV_X2 U5677 ( .I(\SB1_3_3/buf_output[3] ), .ZN(\SB2_3_1/i0[8] ) );
  XOR2_X1 U5678 ( .A1(\MC_ARK_ARC_1_3/temp1[157] ), .A2(n4967), .Z(
        \MC_ARK_ARC_1_3/temp5[157] ) );
  XOR2_X1 U5679 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[103] ), .A2(\RI5[3][127] ), 
        .Z(n4967) );
  NAND3_X2 U5690 ( .A1(\SB2_3_11/i0[10] ), .A2(\SB2_3_11/i1_7 ), .A3(
        \SB2_3_11/i1[9] ), .ZN(n6331) );
  XOR2_X1 U5693 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[163] ), .A2(\RI5[1][127] ), 
        .Z(\MC_ARK_ARC_1_1/temp3[61] ) );
  NAND2_X2 U5694 ( .A1(n3145), .A2(n5402), .ZN(
        \MC_ARK_ARC_1_1/buf_datainput[163] ) );
  INV_X2 U5696 ( .I(\SB1_0_25/buf_output[3] ), .ZN(\SB2_0_23/i0[8] ) );
  NAND4_X2 U5699 ( .A1(\SB1_0_25/Component_Function_3/NAND4_in[2] ), .A2(
        \SB1_0_25/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_0_25/Component_Function_3/NAND4_in[1] ), .A4(n3313), .ZN(
        \SB1_0_25/buf_output[3] ) );
  XOR2_X1 U5701 ( .A1(n5605), .A2(n4969), .Z(n5806) );
  XOR2_X1 U5710 ( .A1(\RI5[2][120] ), .A2(\RI5[2][114] ), .Z(n4969) );
  NAND3_X1 U5711 ( .A1(\SB2_1_15/i0[10] ), .A2(\SB2_1_15/i0_0 ), .A3(
        \SB1_1_19/buf_output[1] ), .ZN(
        \SB2_1_15/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U5714 ( .A1(\SB2_3_8/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_3_8/Component_Function_1/NAND4_in[3] ), .A3(n3059), .A4(
        \SB2_3_8/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_3_8/buf_output[1] ) );
  NAND3_X2 U5718 ( .A1(\SB2_0_4/i0_3 ), .A2(\SB2_0_4/i0[6] ), .A3(
        \SB2_0_4/i1[9] ), .ZN(n4970) );
  NAND3_X1 U5725 ( .A1(\SB1_2_18/i0_0 ), .A2(\SB1_2_18/i0[9] ), .A3(n4762), 
        .ZN(\SB1_2_18/Component_Function_4/NAND4_in[0] ) );
  NAND3_X2 U5727 ( .A1(\SB2_3_26/i0_0 ), .A2(\SB1_3_28/buf_output[3] ), .A3(
        \SB2_3_26/i0[6] ), .ZN(n4971) );
  NAND3_X1 U5730 ( .A1(\SB2_1_26/i0[6] ), .A2(\SB2_1_26/i0[9] ), .A3(
        \SB2_1_26/i1_5 ), .ZN(n4983) );
  NAND3_X1 U5731 ( .A1(\SB3_3/i0[6] ), .A2(\SB3_3/i0_3 ), .A3(\SB3_3/i1[9] ), 
        .ZN(\SB3_3/Component_Function_3/NAND4_in[0] ) );
  NAND4_X2 U5732 ( .A1(\SB2_3_18/Component_Function_3/NAND4_in[0] ), .A2(n2251), .A3(\SB2_3_18/Component_Function_3/NAND4_in[2] ), .A4(n4972), .ZN(
        \SB2_3_18/buf_output[3] ) );
  NAND3_X2 U5733 ( .A1(\SB2_3_18/i0_3 ), .A2(\SB2_3_18/i0_0 ), .A3(
        \SB2_3_18/i0_4 ), .ZN(n4972) );
  XOR2_X1 U5734 ( .A1(\RI5[3][69] ), .A2(\SB2_3_28/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_3/temp3[159] ) );
  NAND4_X2 U5735 ( .A1(\SB2_3_11/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_11/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_3_11/Component_Function_5/NAND4_in[0] ), .A4(n4154), .ZN(
        \SB2_3_11/buf_output[5] ) );
  NAND4_X2 U5736 ( .A1(\SB2_1_26/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_1_26/Component_Function_0/NAND4_in[1] ), .A3(n4075), .A4(n4973), 
        .ZN(\SB2_1_26/buf_output[0] ) );
  NAND3_X1 U5739 ( .A1(\SB2_1_26/i0_0 ), .A2(\SB2_1_26/i0_3 ), .A3(
        \SB2_1_26/i0[7] ), .ZN(n4973) );
  NAND4_X2 U5741 ( .A1(\SB1_3_11/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_3_11/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_3_11/Component_Function_0/NAND4_in[1] ), .A4(n4974), .ZN(
        \SB1_3_11/buf_output[0] ) );
  NAND3_X2 U5746 ( .A1(\SB2_2_25/i0_4 ), .A2(\SB2_2_25/i0_0 ), .A3(
        \SB2_2_25/i1_5 ), .ZN(\SB2_2_25/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U5755 ( .A1(\SB1_3_5/i0_3 ), .A2(\SB1_3_5/i0[8] ), .A3(
        \SB1_3_5/i1_7 ), .ZN(\SB1_3_5/Component_Function_1/NAND4_in[1] ) );
  NAND3_X2 U5761 ( .A1(\SB1_2_26/i1_5 ), .A2(\SB1_2_26/i1[9] ), .A3(
        \SB1_2_26/i0_4 ), .ZN(n4714) );
  NAND4_X2 U5762 ( .A1(\SB1_3_19/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_3_19/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_3_19/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_3_19/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_3_19/buf_output[0] ) );
  NAND4_X2 U5763 ( .A1(n657), .A2(n5031), .A3(n5637), .A4(n6509), .ZN(
        \SB2_3_28/buf_output[2] ) );
  NAND4_X2 U5764 ( .A1(\SB2_2_0/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_0/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_2_0/Component_Function_1/NAND4_in[1] ), .A4(
        \SB2_2_0/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB2_2_0/buf_output[1] ) );
  NAND2_X2 U5767 ( .A1(\SB1_3_29/i1[9] ), .A2(\SB1_3_29/i0_3 ), .ZN(
        \SB1_3_29/Component_Function_1/NAND4_in[0] ) );
  NAND4_X2 U5772 ( .A1(\SB4_21/Component_Function_1/NAND4_in[3] ), .A2(
        \SB4_21/Component_Function_1/NAND4_in[1] ), .A3(
        \SB4_21/Component_Function_1/NAND4_in[0] ), .A4(
        \SB4_21/Component_Function_1/NAND4_in[2] ), .ZN(n2775) );
  NAND4_X2 U5773 ( .A1(\SB2_0_15/Component_Function_5/NAND4_in[3] ), .A2(n1306), .A3(\SB2_0_15/Component_Function_5/NAND4_in[0] ), .A4(n5473), .ZN(
        \SB2_0_15/buf_output[5] ) );
  NAND3_X2 U5775 ( .A1(\SB1_0_15/i0[6] ), .A2(\SB1_0_15/i0[10] ), .A3(
        \SB1_0_15/i0_0 ), .ZN(\SB1_0_15/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U5776 ( .A1(\SB2_3_25/i0_3 ), .A2(\SB2_3_25/i0[6] ), .A3(
        \SB2_3_25/i0[10] ), .ZN(n4975) );
  NAND4_X2 U5777 ( .A1(\SB1_0_29/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_0_29/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_0_29/Component_Function_0/NAND4_in[0] ), .A4(n4976), .ZN(
        \SB1_0_29/buf_output[0] ) );
  NAND3_X1 U5779 ( .A1(\SB1_0_29/i0_4 ), .A2(\SB1_0_29/i0[10] ), .A3(
        \SB1_0_29/i0_3 ), .ZN(n4976) );
  XOR2_X1 U5780 ( .A1(n2371), .A2(n4977), .Z(\MC_ARK_ARC_1_2/buf_output[58] )
         );
  XOR2_X1 U5784 ( .A1(\MC_ARK_ARC_1_2/temp4[58] ), .A2(n3132), .Z(n4977) );
  NAND3_X1 U5785 ( .A1(\SB1_0_15/i0[6] ), .A2(\SB1_0_15/i0[8] ), .A3(
        \SB1_0_15/i0[7] ), .ZN(\SB1_0_15/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U5787 ( .A1(\SB2_3_19/i0_3 ), .A2(\SB2_3_19/i0[9] ), .A3(
        \SB2_3_19/i0[8] ), .ZN(\SB2_3_19/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U5789 ( .A1(\SB1_3_29/i1[9] ), .A2(\SB1_3_29/i0_3 ), .A3(
        \SB1_3_29/i0[6] ), .ZN(\SB1_3_29/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U5790 ( .A1(\SB2_1_25/i0[10] ), .A2(\SB2_1_25/i1_7 ), .A3(
        \SB2_1_25/i1[9] ), .ZN(n4978) );
  NAND3_X2 U5791 ( .A1(\SB2_1_18/i0_3 ), .A2(\SB2_1_18/i0[10] ), .A3(
        \SB1_1_22/buf_output[1] ), .ZN(n4979) );
  NAND4_X2 U5792 ( .A1(\SB2_0_24/Component_Function_3/NAND4_in[3] ), .A2(
        \SB2_0_24/Component_Function_3/NAND4_in[0] ), .A3(n800), .A4(n4980), 
        .ZN(\SB2_0_24/buf_output[3] ) );
  NAND3_X2 U5793 ( .A1(\SB2_0_24/i0_3 ), .A2(\SB2_0_24/i0_0 ), .A3(
        \RI3[0][46] ), .ZN(n4980) );
  NOR2_X2 U5796 ( .A1(n4981), .A2(n2334), .ZN(\SB2_3_28/i0[7] ) );
  NAND2_X1 U5797 ( .A1(n953), .A2(n2555), .ZN(n4981) );
  XOR2_X1 U5804 ( .A1(n4982), .A2(n198), .Z(Ciphertext[133]) );
  NAND4_X2 U5805 ( .A1(\SB4_9/Component_Function_1/NAND4_in[1] ), .A2(n3871), 
        .A3(n2693), .A4(\SB4_9/Component_Function_1/NAND4_in[0] ), .ZN(n4982)
         );
  INV_X2 U5808 ( .I(\SB1_2_29/buf_output[2] ), .ZN(\SB2_2_26/i1[9] ) );
  XOR2_X1 U5809 ( .A1(n4984), .A2(n215), .Z(Ciphertext[134]) );
  NAND4_X2 U5810 ( .A1(n6399), .A2(n927), .A3(n5006), .A4(n6379), .ZN(n4984)
         );
  XOR2_X1 U5811 ( .A1(\MC_ARK_ARC_1_2/temp5[115] ), .A2(n4985), .Z(
        \MC_ARK_ARC_1_2/buf_output[115] ) );
  XOR2_X1 U5812 ( .A1(\MC_ARK_ARC_1_2/temp4[115] ), .A2(
        \MC_ARK_ARC_1_2/temp3[115] ), .Z(n4985) );
  XOR2_X1 U5816 ( .A1(n6061), .A2(n4986), .Z(\MC_ARK_ARC_1_1/buf_output[181] )
         );
  XOR2_X1 U5817 ( .A1(n5629), .A2(n5630), .Z(n4986) );
  NAND3_X2 U5818 ( .A1(\SB2_2_0/i0_4 ), .A2(\SB2_2_0/i0[9] ), .A3(
        \SB2_2_0/i0[6] ), .ZN(n4987) );
  INV_X2 U5819 ( .I(\SB2_1_31/i0[7] ), .ZN(\SB2_1_31/i0_4 ) );
  NAND3_X1 U5820 ( .A1(\SB2_1_31/i0[6] ), .A2(\SB2_1_31/i0[7] ), .A3(
        \SB2_1_31/i0[8] ), .ZN(\SB2_1_31/Component_Function_0/NAND4_in[1] ) );
  NOR2_X2 U5823 ( .A1(n5999), .A2(n5827), .ZN(\SB2_1_31/i0[7] ) );
  XOR2_X1 U5824 ( .A1(n4988), .A2(n68), .Z(Ciphertext[187]) );
  NAND4_X2 U5825 ( .A1(\SB4_0/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_0/Component_Function_1/NAND4_in[2] ), .A3(
        \SB4_0/Component_Function_1/NAND4_in[3] ), .A4(n2038), .ZN(n4988) );
  INV_X1 U5826 ( .I(\SB3_31/buf_output[1] ), .ZN(\SB4_27/i1_7 ) );
  NAND4_X2 U5829 ( .A1(\SB3_31/Component_Function_1/NAND4_in[1] ), .A2(
        \SB3_31/Component_Function_1/NAND4_in[2] ), .A3(
        \SB3_31/Component_Function_1/NAND4_in[3] ), .A4(
        \SB3_31/Component_Function_1/NAND4_in[0] ), .ZN(\SB3_31/buf_output[1] ) );
  INV_X2 U5830 ( .I(\SB1_3_5/buf_output[2] ), .ZN(\SB2_3_2/i1[9] ) );
  NAND4_X2 U5831 ( .A1(\SB1_3_5/Component_Function_2/NAND4_in[0] ), .A2(n6228), 
        .A3(n5372), .A4(n2003), .ZN(\SB1_3_5/buf_output[2] ) );
  AND2_X1 U5832 ( .A1(n6270), .A2(n4989), .Z(n4305) );
  NAND3_X1 U5835 ( .A1(\SB2_3_3/i0[8] ), .A2(\SB2_3_3/i1_7 ), .A3(
        \SB1_3_4/buf_output[4] ), .ZN(n4989) );
  XOR2_X1 U5840 ( .A1(n4990), .A2(n135), .Z(Ciphertext[9]) );
  NAND4_X2 U5842 ( .A1(\SB4_30/Component_Function_3/NAND4_in[3] ), .A2(n3935), 
        .A3(n5339), .A4(\SB4_30/Component_Function_3/NAND4_in[2] ), .ZN(n4990)
         );
  XOR2_X1 U5843 ( .A1(n4992), .A2(n4991), .Z(\MC_ARK_ARC_1_2/buf_output[9] )
         );
  XOR2_X1 U5845 ( .A1(n5973), .A2(\MC_ARK_ARC_1_2/temp4[9] ), .Z(n4991) );
  XOR2_X1 U5848 ( .A1(n3068), .A2(n6068), .Z(n4992) );
  XOR2_X1 U5852 ( .A1(n4994), .A2(n216), .Z(Ciphertext[50]) );
  NAND4_X2 U5853 ( .A1(n2628), .A2(\SB4_23/Component_Function_2/NAND4_in[0] ), 
        .A3(\SB4_23/Component_Function_2/NAND4_in[2] ), .A4(n1578), .ZN(n4994)
         );
  XOR2_X1 U5854 ( .A1(n4995), .A2(n138), .Z(Ciphertext[44]) );
  NAND4_X2 U5856 ( .A1(\SB4_24/Component_Function_2/NAND4_in[0] ), .A2(
        \SB4_24/Component_Function_2/NAND4_in[3] ), .A3(
        \SB4_24/Component_Function_2/NAND4_in[2] ), .A4(
        \SB4_24/Component_Function_2/NAND4_in[1] ), .ZN(n4995) );
  NAND4_X2 U5857 ( .A1(\SB2_3_25/Component_Function_4/NAND4_in[0] ), .A2(n4492), .A3(\SB2_3_25/Component_Function_4/NAND4_in[1] ), .A4(n4996), .ZN(
        \SB2_3_25/buf_output[4] ) );
  NAND3_X1 U5859 ( .A1(\SB2_3_25/i0[9] ), .A2(\SB2_3_25/i0[10] ), .A3(
        \SB2_3_25/i0_3 ), .ZN(n4996) );
  NAND4_X2 U5860 ( .A1(\SB3_24/Component_Function_5/NAND4_in[3] ), .A2(n2578), 
        .A3(n1250), .A4(n4997), .ZN(\SB3_24/buf_output[5] ) );
  XOR2_X1 U5865 ( .A1(\MC_ARK_ARC_1_3/temp5[10] ), .A2(n4998), .Z(
        \MC_ARK_ARC_1_3/buf_output[10] ) );
  XOR2_X1 U5866 ( .A1(\MC_ARK_ARC_1_3/temp4[10] ), .A2(
        \MC_ARK_ARC_1_3/temp3[10] ), .Z(n4998) );
  XOR2_X1 U5876 ( .A1(n4999), .A2(\MC_ARK_ARC_1_1/temp4[163] ), .Z(n6424) );
  XOR2_X1 U5877 ( .A1(\RI5[1][73] ), .A2(\RI5[1][37] ), .Z(n4999) );
  NAND3_X1 U5879 ( .A1(\SB4_1/i0_4 ), .A2(\SB4_1/i0_3 ), .A3(\SB4_1/i0[10] ), 
        .ZN(\SB4_1/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U5880 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[67] ), .A2(\RI5[0][19] ), 
        .Z(n5385) );
  NAND4_X2 U5882 ( .A1(\SB2_2_10/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_10/Component_Function_2/NAND4_in[2] ), .A3(n3495), .A4(n5985), 
        .ZN(\SB2_2_10/buf_output[2] ) );
  NAND3_X2 U5886 ( .A1(\SB1_1_19/i0_0 ), .A2(\SB1_1_19/i0[6] ), .A3(
        \SB1_1_19/i0[10] ), .ZN(n5001) );
  NAND4_X2 U5888 ( .A1(n3725), .A2(\SB2_2_11/Component_Function_5/NAND4_in[2] ), .A3(n5987), .A4(n5002), .ZN(\SB2_2_11/buf_output[5] ) );
  NAND3_X2 U5889 ( .A1(\SB2_2_11/i0_4 ), .A2(\SB2_2_11/i0[6] ), .A3(
        \SB2_2_11/i0[9] ), .ZN(n5002) );
  XOR2_X1 U5890 ( .A1(n5003), .A2(n143), .Z(Ciphertext[11]) );
  NAND4_X2 U5894 ( .A1(\SB4_30/Component_Function_5/NAND4_in[2] ), .A2(
        \SB4_30/Component_Function_5/NAND4_in[0] ), .A3(n5172), .A4(
        \SB4_30/Component_Function_5/NAND4_in[3] ), .ZN(n5003) );
  INV_X2 U5895 ( .I(\SB1_3_18/buf_output[2] ), .ZN(\SB2_3_15/i1[9] ) );
  NAND3_X1 U5896 ( .A1(\SB4_3/i0_4 ), .A2(\SB4_3/i1_5 ), .A3(n1371), .ZN(n5266) );
  NOR2_X2 U5900 ( .A1(n5005), .A2(n5004), .ZN(n1371) );
  NAND2_X1 U5902 ( .A1(\SB3_6/Component_Function_2/NAND4_in[1] ), .A2(
        \SB3_6/Component_Function_2/NAND4_in[0] ), .ZN(n5005) );
  NAND4_X2 U5910 ( .A1(\SB2_2_25/Component_Function_5/NAND4_in[2] ), .A2(n2145), .A3(n5298), .A4(\SB2_2_25/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_2_25/buf_output[5] ) );
  INV_X2 U5912 ( .I(\SB1_2_15/buf_output[2] ), .ZN(\SB2_2_12/i1[9] ) );
  NAND4_X2 U5914 ( .A1(\SB1_2_15/Component_Function_2/NAND4_in[1] ), .A2(n5314), .A3(\SB1_2_15/Component_Function_2/NAND4_in[0] ), .A4(
        \SB1_2_15/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB1_2_15/buf_output[2] ) );
  NAND3_X2 U5917 ( .A1(\SB2_2_13/i0[6] ), .A2(\SB2_2_13/i0_3 ), .A3(
        \SB2_2_13/i1[9] ), .ZN(n5712) );
  XOR2_X1 U5921 ( .A1(\SB2_2_8/buf_output[5] ), .A2(\RI5[2][137] ), .Z(n5426)
         );
  NAND3_X1 U5928 ( .A1(\SB4_9/i0[9] ), .A2(\SB4_9/i0_3 ), .A3(\SB4_9/i0[8] ), 
        .ZN(n5006) );
  XOR2_X1 U5930 ( .A1(\MC_ARK_ARC_1_2/temp1[140] ), .A2(n5007), .Z(n1928) );
  XOR2_X1 U5931 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[86] ), .A2(\RI5[2][110] ), 
        .Z(n5007) );
  XOR2_X1 U5936 ( .A1(\MC_ARK_ARC_1_3/temp2[123] ), .A2(n5008), .Z(
        \MC_ARK_ARC_1_3/temp5[123] ) );
  XOR2_X1 U5938 ( .A1(\RI5[3][123] ), .A2(\RI5[3][117] ), .Z(n5008) );
  NAND3_X2 U5940 ( .A1(\SB1_2_13/i0[10] ), .A2(\SB1_2_13/i1_7 ), .A3(
        \SB1_2_13/i1[9] ), .ZN(n2763) );
  CLKBUF_X4 U5941 ( .I(\SB2_2_9/buf_output[2] ), .Z(\RI5[2][152] ) );
  NAND3_X1 U5942 ( .A1(\SB1_3_19/i0[10] ), .A2(\SB1_3_19/i0_3 ), .A3(
        \SB1_3_19/i0_4 ), .ZN(\SB1_3_19/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 U5943 ( .A1(\SB1_3_7/i0[9] ), .A2(\SB1_3_7/i0_3 ), .A3(
        \SB1_3_7/i0[8] ), .ZN(n5036) );
  NAND3_X1 U5946 ( .A1(\SB3_2/i0[10] ), .A2(\SB3_2/i1[9] ), .A3(\SB3_2/i1_5 ), 
        .ZN(n5669) );
  NAND3_X2 U5947 ( .A1(\SB1_2_9/i0[9] ), .A2(\SB1_2_9/i0[6] ), .A3(
        \SB1_2_9/i0_4 ), .ZN(n3886) );
  NAND4_X2 U5948 ( .A1(\SB2_1_5/Component_Function_5/NAND4_in[2] ), .A2(n5938), 
        .A3(n5326), .A4(\SB2_1_5/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB2_1_5/buf_output[5] ) );
  NAND3_X1 U5955 ( .A1(\SB2_3_6/i0[10] ), .A2(\SB2_3_6/i1[9] ), .A3(
        \SB2_3_6/i1_5 ), .ZN(\SB2_3_6/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U5958 ( .A1(\SB1_2_25/i0[10] ), .A2(\SB1_2_25/i1[9] ), .A3(
        \SB1_2_25/i1_7 ), .ZN(\SB1_2_25/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U5959 ( .A1(\SB4_19/i0[6] ), .A2(\SB3_21/buf_output[3] ), .A3(
        \SB4_19/i0_3 ), .ZN(\SB4_19/Component_Function_2/NAND4_in[1] ) );
  NAND4_X2 U5963 ( .A1(n1992), .A2(n5183), .A3(
        \SB2_1_23/Component_Function_5/NAND4_in[0] ), .A4(n5009), .ZN(
        \SB2_1_23/buf_output[5] ) );
  NAND3_X2 U5967 ( .A1(\SB2_1_23/i0[6] ), .A2(\SB2_1_23/i0[10] ), .A3(
        \SB2_1_23/i0_0 ), .ZN(n5009) );
  NAND3_X1 U5968 ( .A1(\SB3_27/i0[10] ), .A2(\SB3_27/i1_5 ), .A3(n4764), .ZN(
        \SB3_27/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U5969 ( .A1(\MC_ARK_ARC_1_0/temp2[29] ), .A2(n5011), .Z(
        \MC_ARK_ARC_1_0/temp5[29] ) );
  XOR2_X1 U5970 ( .A1(\RI5[0][29] ), .A2(\RI5[0][23] ), .Z(n5011) );
  NAND4_X2 U5971 ( .A1(\SB4_21/Component_Function_3/NAND4_in[3] ), .A2(n6455), 
        .A3(\SB4_21/Component_Function_3/NAND4_in[1] ), .A4(n5012), .ZN(n6183)
         );
  NAND3_X1 U5975 ( .A1(\SB4_21/i0[10] ), .A2(\SB4_21/i1_7 ), .A3(n3666), .ZN(
        n5012) );
  XOR2_X1 U5976 ( .A1(n5013), .A2(\MC_ARK_ARC_1_3/temp4[27] ), .Z(
        \MC_ARK_ARC_1_3/temp6[27] ) );
  XOR2_X1 U5980 ( .A1(\RI5[3][93] ), .A2(\RI5[3][129] ), .Z(n5013) );
  XOR2_X1 U5982 ( .A1(\SB2_0_25/buf_output[2] ), .A2(\RI5[0][50] ), .Z(n3126)
         );
  XOR2_X1 U5983 ( .A1(n5014), .A2(n152), .Z(Ciphertext[47]) );
  NAND4_X2 U5988 ( .A1(\SB4_24/Component_Function_5/NAND4_in[1] ), .A2(
        \SB4_24/Component_Function_5/NAND4_in[2] ), .A3(
        \SB4_24/Component_Function_5/NAND4_in[0] ), .A4(n3015), .ZN(n5014) );
  XOR2_X1 U5994 ( .A1(\MC_ARK_ARC_1_2/temp2[83] ), .A2(n5015), .Z(n817) );
  XOR2_X1 U5995 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[83] ), .A2(\RI5[2][77] ), 
        .Z(n5015) );
  NAND4_X2 U5996 ( .A1(n4284), .A2(\SB1_1_26/Component_Function_2/NAND4_in[2] ), .A3(n2405), .A4(n5016), .ZN(\SB1_1_26/buf_output[2] ) );
  XOR2_X1 U5997 ( .A1(n1198), .A2(\MC_ARK_ARC_1_0/temp6[75] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[75] ) );
  XOR2_X1 U6000 ( .A1(\MC_ARK_ARC_1_0/temp1[75] ), .A2(n1062), .Z(n1198) );
  XOR2_X1 U6002 ( .A1(n613), .A2(n5017), .Z(\MC_ARK_ARC_1_1/buf_output[114] )
         );
  XOR2_X1 U6003 ( .A1(\MC_ARK_ARC_1_1/temp4[114] ), .A2(
        \MC_ARK_ARC_1_1/temp3[114] ), .Z(n5017) );
  XOR2_X1 U6005 ( .A1(n1303), .A2(n5018), .Z(\MC_ARK_ARC_1_0/buf_output[189] )
         );
  XOR2_X1 U6007 ( .A1(\MC_ARK_ARC_1_0/temp4[189] ), .A2(n4337), .Z(n5018) );
  XOR2_X1 U6008 ( .A1(n5020), .A2(n5019), .Z(n6129) );
  XOR2_X1 U6009 ( .A1(\RI5[3][59] ), .A2(n130), .Z(n5019) );
  XOR2_X1 U6014 ( .A1(\RI5[3][29] ), .A2(\RI5[3][95] ), .Z(n5020) );
  NAND4_X2 U6020 ( .A1(\SB2_2_28/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_28/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_2_28/Component_Function_4/NAND4_in[1] ), .A4(n5021), .ZN(
        \SB2_2_28/buf_output[4] ) );
  XOR2_X1 U6022 ( .A1(n5023), .A2(n5022), .Z(\MC_ARK_ARC_1_0/temp5[8] ) );
  XOR2_X1 U6027 ( .A1(\RI5[0][170] ), .A2(\RI5[0][8] ), .Z(n5022) );
  XOR2_X1 U6031 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[2] ), .A2(\RI5[0][146] ), 
        .Z(n5023) );
  XOR2_X1 U6032 ( .A1(\MC_ARK_ARC_1_0/temp2[91] ), .A2(n5024), .Z(
        \MC_ARK_ARC_1_0/temp5[91] ) );
  XOR2_X1 U6034 ( .A1(\RI5[0][85] ), .A2(\RI5[0][91] ), .Z(n5024) );
  NAND3_X2 U6035 ( .A1(\SB2_3_28/i0[6] ), .A2(\SB2_3_28/i0[9] ), .A3(n577), 
        .ZN(n3430) );
  XOR2_X1 U6038 ( .A1(n5025), .A2(n137), .Z(Ciphertext[69]) );
  NAND4_X2 U6049 ( .A1(\SB4_20/Component_Function_3/NAND4_in[0] ), .A2(
        \SB4_20/Component_Function_3/NAND4_in[2] ), .A3(n6217), .A4(n1888), 
        .ZN(n5025) );
  NAND3_X2 U6050 ( .A1(\SB2_0_20/i0_3 ), .A2(\SB2_0_20/i0_0 ), .A3(
        \SB2_0_20/i0_4 ), .ZN(\SB2_0_20/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U6051 ( .A1(n5026), .A2(n170), .Z(Ciphertext[99]) );
  NAND4_X2 U6052 ( .A1(\SB4_15/Component_Function_3/NAND4_in[3] ), .A2(n3848), 
        .A3(n5088), .A4(n4605), .ZN(n5026) );
  XOR2_X1 U6055 ( .A1(\SB2_0_25/buf_output[3] ), .A2(\RI5[0][45] ), .Z(n3978)
         );
  XOR2_X1 U6056 ( .A1(\MC_ARK_ARC_1_0/temp4[137] ), .A2(n5027), .Z(n1877) );
  XOR2_X1 U6059 ( .A1(\RI5[0][11] ), .A2(\RI5[0][47] ), .Z(n5027) );
  XOR2_X1 U6061 ( .A1(\RI5[2][187] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[151] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[85] ) );
  NAND4_X2 U6063 ( .A1(n6355), .A2(\SB1_2_5/Component_Function_2/NAND4_in[2] ), 
        .A3(\SB1_2_5/Component_Function_2/NAND4_in[1] ), .A4(
        \SB1_2_5/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB1_2_5/buf_output[2] ) );
  XOR2_X1 U6065 ( .A1(n5028), .A2(n193), .Z(Ciphertext[109]) );
  NAND3_X1 U6066 ( .A1(\SB1_2_28/i0_4 ), .A2(\SB1_2_28/i1[9] ), .A3(
        \SB1_2_28/i1_5 ), .ZN(\SB1_2_28/Component_Function_4/NAND4_in[3] ) );
  BUF_X2 U6069 ( .I(\SB2_3_12/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[119] ) );
  INV_X1 U6073 ( .I(n5030), .ZN(n5029) );
  NAND2_X1 U6075 ( .A1(\SB1_2_14/buf_output[1] ), .A2(\SB1_2_12/buf_output[3] ), .ZN(n5030) );
  NAND3_X2 U6077 ( .A1(\SB2_3_28/i0[6] ), .A2(\SB2_3_28/i0_3 ), .A3(n5511), 
        .ZN(n5031) );
  XOR2_X1 U6082 ( .A1(\MC_ARK_ARC_1_2/temp5[20] ), .A2(n5032), .Z(
        \MC_ARK_ARC_1_2/buf_output[20] ) );
  XOR2_X1 U6085 ( .A1(\MC_ARK_ARC_1_2/temp4[20] ), .A2(n5578), .Z(n5032) );
  INV_X1 U6089 ( .I(\SB1_3_6/buf_output[5] ), .ZN(\SB2_3_6/i1_5 ) );
  NAND4_X2 U6090 ( .A1(\SB1_3_6/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_6/Component_Function_5/NAND4_in[3] ), .A3(n5222), .A4(
        \SB1_3_6/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_6/buf_output[5] ) );
  NAND3_X2 U6091 ( .A1(\SB1_3_22/i0_3 ), .A2(\SB1_3_22/i0_4 ), .A3(
        \SB1_3_22/i1[9] ), .ZN(n5033) );
  NAND4_X2 U6098 ( .A1(\SB3_0/Component_Function_1/NAND4_in[2] ), .A2(
        \SB3_0/Component_Function_1/NAND4_in[1] ), .A3(n962), .A4(n5034), .ZN(
        \SB3_0/buf_output[1] ) );
  NAND2_X1 U6100 ( .A1(\SB3_0/i0_3 ), .A2(\SB3_0/i1[9] ), .ZN(n5034) );
  NAND4_X2 U6101 ( .A1(\SB2_1_19/Component_Function_5/NAND4_in[1] ), .A2(
        \SB2_1_19/Component_Function_5/NAND4_in[2] ), .A3(n5035), .A4(
        \SB2_1_19/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_1_19/buf_output[5] ) );
  NAND3_X2 U6108 ( .A1(\SB2_1_19/i0[6] ), .A2(n578), .A3(\SB2_1_19/i0[9] ), 
        .ZN(n5035) );
  NAND4_X2 U6112 ( .A1(\SB1_3_7/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_7/Component_Function_2/NAND4_in[1] ), .A3(n6022), .A4(n5036), 
        .ZN(\SB1_3_7/buf_output[2] ) );
  NAND4_X2 U6114 ( .A1(\SB2_2_29/Component_Function_3/NAND4_in[1] ), .A2(n5438), .A3(\SB2_2_29/Component_Function_3/NAND4_in[0] ), .A4(n5037), .ZN(
        \SB2_2_29/buf_output[3] ) );
  NAND3_X1 U6119 ( .A1(\SB2_2_29/i0[10] ), .A2(\SB2_2_29/i1[9] ), .A3(
        \SB2_2_29/i1_7 ), .ZN(n5037) );
  XOR2_X1 U6120 ( .A1(n5039), .A2(n5038), .Z(n2803) );
  XOR2_X1 U6121 ( .A1(n6190), .A2(n575), .Z(n5038) );
  XOR2_X1 U6125 ( .A1(n2664), .A2(n3012), .Z(n5039) );
  XOR2_X1 U6126 ( .A1(\MC_ARK_ARC_1_3/temp2[185] ), .A2(n5040), .Z(
        \MC_ARK_ARC_1_3/temp5[185] ) );
  XOR2_X1 U6129 ( .A1(\RI5[3][185] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[179] ), 
        .Z(n5040) );
  NAND3_X1 U6130 ( .A1(\SB1_0_19/i0[10] ), .A2(\SB1_0_19/i0[9] ), .A3(
        \SB1_0_19/i0_3 ), .ZN(\SB1_0_19/Component_Function_4/NAND4_in[2] ) );
  NAND3_X2 U6131 ( .A1(\SB2_3_8/i0_3 ), .A2(\SB1_3_9/buf_output[4] ), .A3(
        \SB2_3_8/i0_0 ), .ZN(\SB2_3_8/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U6133 ( .A1(n2218), .A2(\SB2_0_22/Component_Function_5/NAND4_in[0] ), .A3(n5930), .A4(n3855), .ZN(\SB2_0_22/buf_output[5] ) );
  NAND4_X2 U6134 ( .A1(\SB1_2_18/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_2_18/Component_Function_0/NAND4_in[0] ), .A3(
        \SB1_2_18/Component_Function_0/NAND4_in[2] ), .A4(n5041), .ZN(
        \SB1_2_18/buf_output[0] ) );
  NAND3_X2 U6136 ( .A1(\SB1_2_18/i0_0 ), .A2(\SB1_2_18/i0[7] ), .A3(
        \SB1_2_18/i0_3 ), .ZN(n5041) );
  NAND3_X1 U6139 ( .A1(\SB2_0_17/i0_0 ), .A2(\SB2_0_17/i0[9] ), .A3(
        \SB2_0_17/i0[8] ), .ZN(\SB2_0_17/Component_Function_4/NAND4_in[0] ) );
  NAND3_X2 U6140 ( .A1(\SB2_2_5/i0[6] ), .A2(\SB2_2_5/i0_4 ), .A3(
        \SB2_2_5/i0[9] ), .ZN(\SB2_2_5/Component_Function_5/NAND4_in[3] ) );
  NAND3_X2 U6146 ( .A1(\SB1_1_21/i0[10] ), .A2(\SB1_1_21/i0[6] ), .A3(
        \SB1_1_21/i0_0 ), .ZN(\SB1_1_21/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U6148 ( .A1(n2408), .A2(\SB2_3_8/Component_Function_3/NAND4_in[0] ), 
        .A3(\SB2_3_8/Component_Function_3/NAND4_in[1] ), .A4(n4728), .ZN(
        \SB2_3_8/buf_output[3] ) );
  NAND3_X1 U6150 ( .A1(\SB2_0_25/i0_0 ), .A2(\SB2_0_25/i0[9] ), .A3(
        \SB2_0_25/i0[8] ), .ZN(\SB2_0_25/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U6152 ( .A1(\SB4_30/i0_4 ), .A2(n5525), .A3(n4751), .ZN(
        \SB4_30/Component_Function_4/NAND4_in[3] ) );
  NAND4_X2 U6153 ( .A1(\SB2_3_3/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_3/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_3_3/Component_Function_3/NAND4_in[3] ), .A4(
        \SB2_3_3/Component_Function_3/NAND4_in[1] ), .ZN(
        \SB2_3_3/buf_output[3] ) );
  NAND4_X2 U6156 ( .A1(\SB1_3_0/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_3_0/Component_Function_0/NAND4_in[1] ), .A3(n5307), .A4(
        \SB1_3_0/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_3_0/buf_output[0] ) );
  INV_X4 U6157 ( .I(n5042), .ZN(\SB2_1_0/i1_5 ) );
  XOR2_X1 U6165 ( .A1(\RI5[0][19] ), .A2(\RI5[0][13] ), .Z(n1307) );
  NAND4_X2 U6167 ( .A1(\SB2_2_28/Component_Function_5/NAND4_in[1] ), .A2(
        \SB2_2_28/Component_Function_5/NAND4_in[3] ), .A3(n1741), .A4(
        \SB2_2_28/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_2_28/buf_output[5] ) );
  NAND3_X2 U6168 ( .A1(\SB2_2_28/i0[10] ), .A2(\SB2_2_28/i0_0 ), .A3(
        \SB2_2_28/i0[6] ), .ZN(\SB2_2_28/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U6169 ( .A1(\SB3_1/Component_Function_1/NAND4_in[3] ), .A2(
        \SB3_1/Component_Function_1/NAND4_in[2] ), .A3(n5376), .A4(
        \SB3_1/Component_Function_1/NAND4_in[0] ), .ZN(\SB3_1/buf_output[1] )
         );
  XOR2_X1 U6170 ( .A1(n5043), .A2(n52), .Z(Ciphertext[13]) );
  NAND4_X2 U6173 ( .A1(\SB4_29/Component_Function_1/NAND4_in[1] ), .A2(n4096), 
        .A3(n5117), .A4(\SB4_29/Component_Function_1/NAND4_in[0] ), .ZN(n5043)
         );
  NAND3_X2 U6174 ( .A1(\SB2_1_16/i1[9] ), .A2(\SB2_1_16/i0_3 ), .A3(
        \SB2_1_16/i0[6] ), .ZN(\SB2_1_16/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U6175 ( .A1(\MC_ARK_ARC_1_2/temp2[44] ), .A2(n5044), .Z(
        \MC_ARK_ARC_1_2/temp5[44] ) );
  XOR2_X1 U6182 ( .A1(\RI5[2][44] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[38] ), 
        .Z(n5044) );
  XOR2_X1 U6184 ( .A1(n5045), .A2(n75), .Z(Ciphertext[160]) );
  NAND4_X2 U6185 ( .A1(n2766), .A2(\SB4_5/Component_Function_4/NAND4_in[0] ), 
        .A3(n5667), .A4(\SB4_5/Component_Function_4/NAND4_in[2] ), .ZN(n5045)
         );
  NAND4_X2 U6186 ( .A1(n5109), .A2(\SB2_2_27/Component_Function_5/NAND4_in[3] ), .A3(\SB2_2_27/Component_Function_5/NAND4_in[1] ), .A4(n5046), .ZN(
        \SB2_2_27/buf_output[5] ) );
  NAND2_X2 U6191 ( .A1(\SB2_2_27/i0_0 ), .A2(\SB2_2_27/i3[0] ), .ZN(n5046) );
  INV_X2 U6192 ( .I(n5047), .ZN(n5495) );
  NAND4_X2 U6193 ( .A1(\SB3_5/Component_Function_3/NAND4_in[3] ), .A2(
        \SB3_5/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_5/Component_Function_3/NAND4_in[2] ), .A4(n2249), .ZN(n5047) );
  NAND3_X2 U6194 ( .A1(\SB3_8/i0_0 ), .A2(\SB3_8/i1_5 ), .A3(\SB3_8/i0_4 ), 
        .ZN(\SB3_8/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U6196 ( .A1(\SB1_3_30/i0[10] ), .A2(\SB1_3_30/i0[6] ), .A3(
        \SB1_3_30/i0_3 ), .ZN(n5048) );
  XOR2_X1 U6197 ( .A1(\MC_ARK_ARC_1_0/temp2[191] ), .A2(n5049), .Z(n3821) );
  XOR2_X1 U6202 ( .A1(\RI5[0][185] ), .A2(\RI5[0][191] ), .Z(n5049) );
  AND2_X1 U6203 ( .A1(n1060), .A2(n5050), .Z(n1209) );
  NAND3_X1 U6204 ( .A1(\SB1_3_21/i1[9] ), .A2(\SB1_3_21/i1_5 ), .A3(
        \MC_ARK_ARC_1_2/buf_output[64] ), .ZN(n5050) );
  XOR2_X1 U6205 ( .A1(\RI5[3][4] ), .A2(\RI5[3][160] ), .Z(
        \MC_ARK_ARC_1_3/temp3[94] ) );
  NAND2_X2 U6206 ( .A1(n4017), .A2(n4016), .ZN(\RI5[3][160] ) );
  NAND4_X2 U6211 ( .A1(\SB3_16/Component_Function_5/NAND4_in[2] ), .A2(
        \SB3_16/Component_Function_5/NAND4_in[1] ), .A3(
        \SB3_16/Component_Function_5/NAND4_in[0] ), .A4(n5051), .ZN(
        \SB3_16/buf_output[5] ) );
  NAND3_X2 U6215 ( .A1(\SB3_16/i0[9] ), .A2(\SB3_16/i0_4 ), .A3(\SB3_16/i0[6] ), .ZN(n5051) );
  XOR2_X1 U6221 ( .A1(n2596), .A2(n5052), .Z(\MC_ARK_ARC_1_1/buf_output[63] )
         );
  XOR2_X1 U6222 ( .A1(\MC_ARK_ARC_1_1/temp2[63] ), .A2(
        \MC_ARK_ARC_1_1/temp1[63] ), .Z(n5052) );
  INV_X2 U6224 ( .I(\SB1_2_21/buf_output[2] ), .ZN(\SB2_2_18/i1[9] ) );
  NAND4_X2 U6230 ( .A1(\SB1_2_21/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_21/Component_Function_2/NAND4_in[2] ), .A3(n5416), .A4(
        \SB1_2_21/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB1_2_21/buf_output[2] ) );
  XOR2_X1 U6231 ( .A1(n5053), .A2(\MC_ARK_ARC_1_1/temp5[68] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[68] ) );
  XOR2_X1 U6232 ( .A1(\MC_ARK_ARC_1_1/temp3[68] ), .A2(
        \MC_ARK_ARC_1_1/temp4[68] ), .Z(n5053) );
  NAND4_X2 U6233 ( .A1(\SB2_2_21/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_2_21/Component_Function_3/NAND4_in[3] ), .A3(
        \SB2_2_21/Component_Function_3/NAND4_in[0] ), .A4(n5055), .ZN(
        \SB2_2_21/buf_output[3] ) );
  NAND3_X2 U6238 ( .A1(\SB2_2_21/i0_0 ), .A2(\SB2_2_21/i0_3 ), .A3(
        \SB2_2_21/i0_4 ), .ZN(n5055) );
  XOR2_X1 U6242 ( .A1(n2234), .A2(n5056), .Z(\MC_ARK_ARC_1_2/buf_output[63] )
         );
  NAND3_X2 U6246 ( .A1(\SB1_2_7/i0_0 ), .A2(\SB1_2_7/i1_5 ), .A3(
        \SB1_2_7/i0_4 ), .ZN(n6042) );
  NAND4_X2 U6252 ( .A1(\SB2_1_4/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_1_4/Component_Function_2/NAND4_in[0] ), .A3(n6012), .A4(
        \SB2_1_4/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_1_4/buf_output[2] ) );
  NAND4_X2 U6253 ( .A1(\SB2_3_21/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_3_21/Component_Function_1/NAND4_in[1] ), .A3(n3191), .A4(
        \SB2_3_21/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_3_21/buf_output[1] ) );
  NAND4_X2 U6254 ( .A1(\SB1_3_19/Component_Function_3/NAND4_in[1] ), .A2(n5287), .A3(n2373), .A4(n820), .ZN(\SB1_3_19/buf_output[3] ) );
  NAND3_X2 U6260 ( .A1(\SB1_2_8/i0_3 ), .A2(\SB1_2_8/i1_7 ), .A3(
        \SB1_2_8/i0[8] ), .ZN(n4589) );
  NAND4_X2 U6261 ( .A1(\SB2_2_28/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_2_28/Component_Function_2/NAND4_in[0] ), .A3(n5174), .A4(
        \SB2_2_28/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_2_28/buf_output[2] ) );
  XOR2_X1 U6262 ( .A1(\RI5[1][47] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[41] ), 
        .Z(n5389) );
  NAND4_X2 U6265 ( .A1(\SB2_3_21/Component_Function_5/NAND4_in[3] ), .A2(
        \SB2_3_21/Component_Function_5/NAND4_in[2] ), .A3(n5132), .A4(
        \SB2_3_21/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_3_21/buf_output[5] ) );
  NAND3_X1 U6268 ( .A1(\SB2_3_28/i0[6] ), .A2(\SB2_3_28/i0_3 ), .A3(n2911), 
        .ZN(\SB2_3_28/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U6272 ( .A1(\SB1_1_27/i0[10] ), .A2(\SB1_1_27/i1[9] ), .A3(
        \SB1_1_27/i1_5 ), .ZN(\SB1_1_27/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U6281 ( .A1(\MC_ARK_ARC_1_1/temp6[146] ), .A2(
        \MC_ARK_ARC_1_1/temp5[146] ), .Z(\MC_ARK_ARC_1_1/buf_output[146] ) );
  INV_X1 U6287 ( .I(\SB1_3_21/buf_output[5] ), .ZN(\SB2_3_21/i1_5 ) );
  NAND4_X2 U6288 ( .A1(n4072), .A2(n5252), .A3(
        \SB1_3_21/Component_Function_5/NAND4_in[1] ), .A4(
        \SB1_3_21/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_21/buf_output[5] ) );
  NAND4_X2 U6290 ( .A1(\SB1_2_24/Component_Function_5/NAND4_in[2] ), .A2(n887), 
        .A3(n5152), .A4(\SB1_2_24/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_2_24/buf_output[5] ) );
  NAND3_X2 U6298 ( .A1(\SB1_3_3/i0_3 ), .A2(\SB1_3_3/i1[9] ), .A3(
        \SB1_3_3/i0_4 ), .ZN(\SB1_3_3/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U6301 ( .A1(\SB1_3_7/i1_7 ), .A2(\SB1_3_7/i0_3 ), .A3(
        \SB1_3_7/i0[8] ), .ZN(n6271) );
  NAND2_X2 U6304 ( .A1(\SB2_2_12/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_2_12/Component_Function_1/NAND4_in[2] ), .ZN(n5057) );
  NAND4_X2 U6306 ( .A1(\SB2_2_23/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_23/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_23/Component_Function_5/NAND4_in[0] ), .A4(n5058), .ZN(
        \SB2_2_23/buf_output[5] ) );
  NAND3_X2 U6315 ( .A1(\SB2_2_23/i0[6] ), .A2(\SB2_2_23/i0_4 ), .A3(
        \SB2_2_23/i0[9] ), .ZN(n5058) );
  NAND3_X2 U6316 ( .A1(\SB1_1_17/i0_4 ), .A2(\SB1_1_17/i1[9] ), .A3(
        \SB1_1_17/i1_5 ), .ZN(n5059) );
  XOR2_X1 U6320 ( .A1(n3176), .A2(n4454), .Z(\MC_ARK_ARC_1_2/buf_output[110] )
         );
  XOR2_X1 U6321 ( .A1(n6408), .A2(n1050), .Z(n3176) );
  XOR2_X1 U6322 ( .A1(n3285), .A2(n5060), .Z(\MC_ARK_ARC_1_1/buf_output[115] )
         );
  XOR2_X1 U6323 ( .A1(n3000), .A2(n2999), .Z(n5060) );
  NAND3_X2 U6330 ( .A1(n1670), .A2(\SB1_3_12/buf_output[0] ), .A3(
        \SB1_3_8/buf_output[4] ), .ZN(
        \SB2_3_7/Component_Function_5/NAND4_in[3] ) );
  NAND4_X2 U6333 ( .A1(\SB2_3_24/Component_Function_1/NAND4_in[1] ), .A2(n1013), .A3(\SB2_3_24/Component_Function_1/NAND4_in[0] ), .A4(n5061), .ZN(
        \SB2_3_24/buf_output[1] ) );
  NAND3_X1 U6334 ( .A1(\SB2_3_24/i0_4 ), .A2(\SB2_3_24/i1_7 ), .A3(n2906), 
        .ZN(n5061) );
  NAND4_X2 U6335 ( .A1(\SB1_3_18/Component_Function_3/NAND4_in[1] ), .A2(n3077), .A3(\SB1_3_18/Component_Function_3/NAND4_in[2] ), .A4(n5062), .ZN(
        \SB1_3_18/buf_output[3] ) );
  XOR2_X1 U6344 ( .A1(n5063), .A2(n169), .Z(Ciphertext[21]) );
  NAND4_X2 U6345 ( .A1(n3266), .A2(\SB4_28/Component_Function_3/NAND4_in[3] ), 
        .A3(\SB4_28/Component_Function_3/NAND4_in[2] ), .A4(n4646), .ZN(n5063)
         );
  NAND4_X2 U6350 ( .A1(\SB2_3_10/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_3_10/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_3_10/Component_Function_0/NAND4_in[0] ), .A4(
        \SB2_3_10/Component_Function_0/NAND4_in[1] ), .ZN(
        \SB2_3_10/buf_output[0] ) );
  INV_X1 U6352 ( .I(\SB3_1/buf_output[5] ), .ZN(\SB4_1/i1_5 ) );
  NAND4_X2 U6355 ( .A1(n2958), .A2(\SB3_1/Component_Function_5/NAND4_in[1] ), 
        .A3(n6280), .A4(\SB3_1/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB3_1/buf_output[5] ) );
  XOR2_X1 U6357 ( .A1(n5064), .A2(n200), .Z(Ciphertext[10]) );
  NAND4_X2 U6358 ( .A1(\SB2_3_2/Component_Function_3/NAND4_in[0] ), .A2(n3749), 
        .A3(\SB2_3_2/Component_Function_3/NAND4_in[2] ), .A4(n5065), .ZN(
        \SB2_3_2/buf_output[3] ) );
  NAND3_X2 U6360 ( .A1(\SB2_3_2/i0_4 ), .A2(\SB2_3_2/i0_0 ), .A3(
        \SB2_3_2/i0_3 ), .ZN(n5065) );
  NAND3_X1 U6361 ( .A1(\SB2_2_16/i0_3 ), .A2(\SB2_2_16/i0[6] ), .A3(
        \SB2_2_16/i1[9] ), .ZN(\SB2_2_16/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U6362 ( .A1(\SB1_1_22/i0_0 ), .A2(\SB1_1_22/i0_4 ), .A3(
        \RI1[1][59] ), .ZN(\SB1_1_22/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U6363 ( .A1(\MC_ARK_ARC_1_3/temp2[74] ), .A2(n5066), .Z(
        \MC_ARK_ARC_1_3/temp5[74] ) );
  XOR2_X1 U6364 ( .A1(\RI5[3][68] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[74] ), 
        .Z(n5066) );
  XOR2_X1 U6370 ( .A1(n5067), .A2(\MC_ARK_ARC_1_2/temp4[118] ), .Z(
        \MC_ARK_ARC_1_2/temp6[118] ) );
  XOR2_X1 U6371 ( .A1(n5069), .A2(n115), .Z(Ciphertext[60]) );
  NAND4_X2 U6374 ( .A1(n6179), .A2(\SB4_21/Component_Function_0/NAND4_in[2] ), 
        .A3(n4402), .A4(\SB4_21/Component_Function_0/NAND4_in[3] ), .ZN(n5069)
         );
  XOR2_X1 U6375 ( .A1(n5070), .A2(n3), .Z(Ciphertext[185]) );
  NAND4_X2 U6376 ( .A1(\SB4_1/Component_Function_5/NAND4_in[3] ), .A2(
        \SB4_1/Component_Function_5/NAND4_in[2] ), .A3(
        \SB4_1/Component_Function_5/NAND4_in[0] ), .A4(n5196), .ZN(n5070) );
  XOR2_X1 U6377 ( .A1(n5072), .A2(n5071), .Z(n5650) );
  XOR2_X1 U6380 ( .A1(\RI5[3][89] ), .A2(\RI5[3][149] ), .Z(n5071) );
  XOR2_X1 U6390 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[53] ), .A2(\RI5[3][125] ), 
        .Z(n5072) );
  BUF_X4 U6392 ( .I(\SB2_3_31/buf_output[3] ), .Z(\RI5[3][15] ) );
  XOR2_X1 U6393 ( .A1(\MC_ARK_ARC_1_1/temp4[90] ), .A2(n5073), .Z(n727) );
  XOR2_X1 U6395 ( .A1(\RI5[1][156] ), .A2(\RI5[1][0] ), .Z(n5073) );
  NAND4_X2 U6398 ( .A1(\SB1_3_14/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_14/Component_Function_2/NAND4_in[2] ), .A3(n5355), .A4(n5074), 
        .ZN(\SB1_3_14/buf_output[2] ) );
  NAND3_X2 U6399 ( .A1(\SB1_3_14/i0[10] ), .A2(\SB1_3_14/i1[9] ), .A3(
        \SB1_3_14/i1_5 ), .ZN(n5074) );
  XOR2_X1 U6400 ( .A1(\RI5[0][182] ), .A2(\RI5[0][152] ), .Z(n6219) );
  NAND2_X1 U6403 ( .A1(\SB1_3_3/i0_3 ), .A2(\SB1_3_3/i1[9] ), .ZN(n5075) );
  XOR2_X1 U6407 ( .A1(\MC_ARK_ARC_1_2/temp4[44] ), .A2(n5076), .Z(n5398) );
  XOR2_X1 U6409 ( .A1(n5078), .A2(n5077), .Z(\MC_ARK_ARC_1_0/buf_output[100] )
         );
  XOR2_X1 U6410 ( .A1(n4466), .A2(\MC_ARK_ARC_1_0/temp4[100] ), .Z(n5077) );
  XOR2_X1 U6411 ( .A1(\MC_ARK_ARC_1_0/temp3[100] ), .A2(
        \MC_ARK_ARC_1_0/temp2[100] ), .Z(n5078) );
  NAND3_X1 U6413 ( .A1(\SB2_3_3/i0_3 ), .A2(\SB2_3_3/i0_4 ), .A3(
        \SB2_3_3/i0[10] ), .ZN(\SB2_3_3/Component_Function_0/NAND4_in[2] ) );
  NAND4_X2 U6416 ( .A1(\SB2_0_7/Component_Function_5/NAND4_in[1] ), .A2(n1440), 
        .A3(\SB2_0_7/Component_Function_5/NAND4_in[0] ), .A4(n5079), .ZN(
        \SB2_0_7/buf_output[5] ) );
  NAND3_X1 U6417 ( .A1(\SB2_0_7/i0[9] ), .A2(\SB1_0_8/buf_output[4] ), .A3(
        \SB2_0_7/i0[6] ), .ZN(n5079) );
  NAND3_X2 U6422 ( .A1(\SB2_3_2/i0_4 ), .A2(\SB2_3_2/i0[6] ), .A3(
        \SB2_3_2/i0[9] ), .ZN(n3783) );
  NAND3_X1 U6424 ( .A1(\SB1_2_7/i0[10] ), .A2(\SB1_2_7/i1[9] ), .A3(
        \SB1_2_7/i1_5 ), .ZN(\SB1_2_7/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U6427 ( .A1(\SB2_3_9/i0[10] ), .A2(\SB2_3_9/i1[9] ), .A3(
        \SB2_3_9/i1_5 ), .ZN(\SB2_3_9/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U6428 ( .A1(\SB3_5/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_5/Component_Function_4/NAND4_in[3] ), .A3(n5143), .A4(
        \SB3_5/Component_Function_4/NAND4_in[1] ), .ZN(\SB3_5/buf_output[4] )
         );
  NAND4_X2 U6430 ( .A1(\SB3_4/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_4/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_4/Component_Function_0/NAND4_in[0] ), .A4(n5080), .ZN(
        \SB3_4/buf_output[0] ) );
  NAND3_X2 U6435 ( .A1(\SB3_4/i0_0 ), .A2(\SB3_4/i0_3 ), .A3(\SB3_4/i0[7] ), 
        .ZN(n5080) );
  NAND3_X2 U6437 ( .A1(\SB1_3_18/i0[10] ), .A2(\SB1_3_18/i1_7 ), .A3(
        \SB1_3_18/i1[9] ), .ZN(\SB1_3_18/Component_Function_3/NAND4_in[2] ) );
  XOR2_X1 U6440 ( .A1(n5082), .A2(n5081), .Z(\MC_ARK_ARC_1_1/buf_output[89] )
         );
  XOR2_X1 U6454 ( .A1(\MC_ARK_ARC_1_1/temp1[89] ), .A2(
        \MC_ARK_ARC_1_1/temp4[89] ), .Z(n5082) );
  BUF_X2 U6455 ( .I(\RI3[0][121] ), .Z(\SB2_0_11/i0[6] ) );
  NAND3_X1 U6458 ( .A1(\SB4_30/i0_0 ), .A2(\SB4_30/i0[8] ), .A3(\SB4_30/i0[9] ), .ZN(n691) );
  XOR2_X1 U6473 ( .A1(\RI5[1][171] ), .A2(\RI5[1][147] ), .Z(
        \MC_ARK_ARC_1_1/temp2[9] ) );
  XOR2_X1 U6476 ( .A1(\RI5[0][128] ), .A2(\RI5[0][176] ), .Z(n1960) );
  NAND3_X1 U6481 ( .A1(\SB1_3_9/i0[8] ), .A2(\SB1_3_9/i1_7 ), .A3(
        \SB1_3_9/i0_3 ), .ZN(\SB1_3_9/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U6485 ( .A1(\SB1_2_4/i0[10] ), .A2(\SB1_2_4/i1_5 ), .A3(
        \SB1_2_4/i1[9] ), .ZN(\SB1_2_4/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U6488 ( .A1(\SB2_3_5/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_3_5/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_3_5/Component_Function_4/NAND4_in[3] ), .A4(n1844), .ZN(
        \SB2_3_5/buf_output[4] ) );
  XOR2_X1 U6490 ( .A1(\RI5[0][134] ), .A2(\RI5[0][158] ), .Z(n1762) );
  NAND4_X2 U6500 ( .A1(\SB1_1_20/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_20/Component_Function_3/NAND4_in[3] ), .A3(
        \SB1_1_20/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_1_20/Component_Function_3/NAND4_in[1] ), .ZN(
        \SB1_1_20/buf_output[3] ) );
  NAND3_X2 U6502 ( .A1(\SB2_2_4/i0[6] ), .A2(\SB2_2_4/i0_0 ), .A3(
        \SB2_2_4/i0[10] ), .ZN(\SB2_2_4/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U6509 ( .A1(\SB3_4/i0[10] ), .A2(\SB3_4/i1[9] ), .A3(\SB3_4/i1_7 ), 
        .ZN(n5978) );
  BUF_X4 U6512 ( .I(\MC_ARK_ARC_1_0/buf_output[2] ), .Z(\SB1_1_31/i0_0 ) );
  NAND2_X2 U6513 ( .A1(\SB2_2_30/i0_3 ), .A2(\SB2_2_30/i1[9] ), .ZN(
        \SB2_2_30/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 U6514 ( .A1(\SB1_2_11/i0[10] ), .A2(\SB1_2_11/i0_0 ), .A3(
        \SB1_2_11/i0[6] ), .ZN(n3820) );
  XOR2_X1 U6516 ( .A1(n1873), .A2(\MC_ARK_ARC_1_2/temp1[81] ), .Z(n5226) );
  BUF_X4 U6521 ( .I(\SB2_3_16/buf_output[5] ), .Z(\RI5[3][95] ) );
  NAND4_X2 U6523 ( .A1(\SB1_0_17/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_17/Component_Function_2/NAND4_in[2] ), .A3(n4193), .A4(
        \SB1_0_17/Component_Function_2/NAND4_in[1] ), .ZN(
        \SB1_0_17/buf_output[2] ) );
  NAND4_X2 U6531 ( .A1(\SB2_0_24/Component_Function_2/NAND4_in[2] ), .A2(n1790), .A3(n1789), .A4(\SB2_0_24/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_0_24/buf_output[2] ) );
  XOR2_X1 U6534 ( .A1(n5083), .A2(n225), .Z(Ciphertext[110]) );
  NAND4_X2 U6535 ( .A1(\SB4_13/Component_Function_2/NAND4_in[1] ), .A2(
        \SB4_13/Component_Function_2/NAND4_in[0] ), .A3(
        \SB4_13/Component_Function_2/NAND4_in[2] ), .A4(n6365), .ZN(n5083) );
  NAND4_X2 U6536 ( .A1(\SB1_1_2/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_1_2/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_1_2/Component_Function_4/NAND4_in[1] ), .A4(
        \SB1_1_2/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_1_2/buf_output[4] ) );
  NAND4_X2 U6541 ( .A1(n6486), .A2(n4129), .A3(n2367), .A4(n1765), .ZN(
        \SB3_10/buf_output[5] ) );
  NAND3_X2 U6542 ( .A1(\SB2_3_4/i0_0 ), .A2(\SB2_3_4/i0_4 ), .A3(
        \SB2_3_4/i0_3 ), .ZN(n2053) );
  NAND4_X2 U6544 ( .A1(\SB2_2_23/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_23/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_2_23/Component_Function_2/NAND4_in[1] ), .A4(n5084), .ZN(
        \SB2_2_23/buf_output[2] ) );
  NAND3_X2 U6549 ( .A1(\SB2_2_23/i0_0 ), .A2(\SB2_2_23/i0_4 ), .A3(
        \SB2_2_23/i1_5 ), .ZN(n5084) );
  BUF_X4 U6550 ( .I(\SB1_2_22/buf_output[5] ), .Z(\SB2_2_22/i0_3 ) );
  NAND4_X2 U6551 ( .A1(n2339), .A2(n6518), .A3(n5406), .A4(
        \SB2_3_31/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_3_31/buf_output[5] ) );
  XOR2_X1 U6553 ( .A1(n6309), .A2(n6310), .Z(\MC_ARK_ARC_1_0/buf_output[133] )
         );
  NAND4_X2 U6554 ( .A1(\SB1_2_18/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_18/Component_Function_2/NAND4_in[3] ), .A3(
        \SB1_2_18/Component_Function_2/NAND4_in[2] ), .A4(n5085), .ZN(
        \SB1_2_18/buf_output[2] ) );
  NAND3_X2 U6555 ( .A1(\SB1_2_18/i0[6] ), .A2(\SB1_2_18/i0_3 ), .A3(
        \SB1_2_18/i0[10] ), .ZN(n5085) );
  NAND4_X2 U6556 ( .A1(\SB1_1_9/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_9/Component_Function_3/NAND4_in[2] ), .A3(
        \SB1_1_9/Component_Function_3/NAND4_in[1] ), .A4(n6107), .ZN(
        \SB1_1_9/buf_output[3] ) );
  XOR2_X1 U6559 ( .A1(\RI5[2][80] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[74] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[80] ) );
  XOR2_X1 U6560 ( .A1(\MC_ARK_ARC_1_1/temp6[36] ), .A2(
        \MC_ARK_ARC_1_1/temp5[36] ), .Z(\MC_ARK_ARC_1_1/buf_output[36] ) );
  XOR2_X1 U6561 ( .A1(n761), .A2(n625), .Z(\MC_ARK_ARC_1_1/buf_output[79] ) );
  NAND4_X2 U6564 ( .A1(\SB2_1_11/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_11/Component_Function_5/NAND4_in[0] ), .A3(n5162), .A4(n3987), 
        .ZN(\SB2_1_11/buf_output[5] ) );
  NAND4_X2 U6567 ( .A1(\SB2_1_27/Component_Function_3/NAND4_in[0] ), .A2(n5280), .A3(\SB2_1_27/Component_Function_3/NAND4_in[1] ), .A4(
        \SB2_1_27/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_1_27/buf_output[3] ) );
  NAND4_X2 U6568 ( .A1(\SB2_0_13/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_13/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_0_13/Component_Function_2/NAND4_in[2] ), .A4(n4672), .ZN(
        \SB2_0_13/buf_output[2] ) );
  NAND4_X2 U6569 ( .A1(\SB2_3_1/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_3_1/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_3_1/Component_Function_4/NAND4_in[1] ), .A4(
        \SB2_3_1/Component_Function_4/NAND4_in[2] ), .ZN(
        \SB2_3_1/buf_output[4] ) );
  NAND4_X2 U6573 ( .A1(\SB4_10/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_10/Component_Function_0/NAND4_in[1] ), .A3(
        \SB4_10/Component_Function_0/NAND4_in[0] ), .A4(n5086), .ZN(n3008) );
  NAND3_X1 U6574 ( .A1(\SB4_10/i0_3 ), .A2(\SB3_13/buf_output[2] ), .A3(
        \SB4_10/i0[7] ), .ZN(n5086) );
  NAND4_X2 U6581 ( .A1(\SB2_2_13/Component_Function_2/NAND4_in[2] ), .A2(n1610), .A3(n4591), .A4(n5087), .ZN(\SB2_2_13/buf_output[2] ) );
  NAND3_X2 U6587 ( .A1(\SB2_2_13/i0[10] ), .A2(\SB2_2_13/i0[6] ), .A3(
        \SB2_2_13/i0_3 ), .ZN(n5087) );
  NAND3_X1 U6589 ( .A1(\SB4_15/i0[10] ), .A2(\SB4_15/i1[9] ), .A3(
        \SB4_15/i1_7 ), .ZN(n5088) );
  NAND3_X1 U6591 ( .A1(\SB2_3_22/i0[8] ), .A2(\SB2_3_22/i1_7 ), .A3(
        \SB1_3_23/buf_output[4] ), .ZN(
        \SB2_3_22/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 U6592 ( .A1(\SB2_1_0/i0_0 ), .A2(\SB2_1_0/i1_5 ), .A3(n2687), .ZN(
        \SB2_1_0/Component_Function_2/NAND4_in[3] ) );
  NAND4_X2 U6596 ( .A1(n4682), .A2(\SB2_3_1/Component_Function_3/NAND4_in[0] ), 
        .A3(\SB2_3_1/Component_Function_3/NAND4_in[1] ), .A4(n5089), .ZN(
        \SB2_3_1/buf_output[3] ) );
  NAND3_X2 U6597 ( .A1(\SB2_3_1/i0[10] ), .A2(\SB2_3_1/i1[9] ), .A3(
        \SB2_3_1/i1_7 ), .ZN(n5089) );
  NAND3_X1 U6600 ( .A1(\SB3_5/i0[6] ), .A2(\SB3_5/i0[10] ), .A3(
        \MC_ARK_ARC_1_3/buf_output[161] ), .ZN(n6361) );
  AND4_X2 U6601 ( .A1(\SB3_21/Component_Function_5/NAND4_in[1] ), .A2(
        \SB3_21/Component_Function_5/NAND4_in[0] ), .A3(n2606), .A4(
        \SB3_21/Component_Function_5/NAND4_in[3] ), .Z(\SB4_21/i1_5 ) );
  XOR2_X1 U6603 ( .A1(n5090), .A2(n206), .Z(Ciphertext[62]) );
  NAND4_X2 U6614 ( .A1(\SB4_21/Component_Function_2/NAND4_in[2] ), .A2(n1425), 
        .A3(n5170), .A4(n2279), .ZN(n5090) );
  NAND4_X2 U6622 ( .A1(n3791), .A2(\SB4_16/Component_Function_5/NAND4_in[1] ), 
        .A3(\SB4_16/Component_Function_5/NAND4_in[0] ), .A4(n5091), .ZN(n5131)
         );
  NAND3_X1 U6623 ( .A1(\SB4_16/i0[9] ), .A2(\SB4_16/i0_4 ), .A3(\SB4_16/i0[6] ), .ZN(n5091) );
  INV_X2 U6630 ( .I(\MC_ARK_ARC_1_2/buf_output[121] ), .ZN(\SB1_3_11/i1_7 ) );
  NAND3_X2 U6631 ( .A1(\RI1[2][95] ), .A2(\SB1_2_16/i1[9] ), .A3(
        \SB1_2_16/i0_4 ), .ZN(\SB1_2_16/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U6632 ( .A1(n2687), .A2(\SB2_1_0/i1[9] ), .A3(\SB2_1_0/i1_5 ), .ZN(
        \SB2_1_0/Component_Function_4/NAND4_in[3] ) );
  NAND3_X2 U6634 ( .A1(\SB2_3_7/i1_7 ), .A2(\SB2_3_7/i0_3 ), .A3(
        \SB2_3_7/i0[8] ), .ZN(n5565) );
  INV_X4 U6635 ( .I(\SB2_0_2/i0[7] ), .ZN(\RI3[0][178] ) );
  NAND2_X1 U6638 ( .A1(\SB1_0_3/Component_Function_4/NAND4_in[1] ), .A2(n5846), 
        .ZN(n6435) );
  INV_X1 U6641 ( .I(\SB3_23/buf_output[3] ), .ZN(\SB4_21/i0[8] ) );
  NAND4_X2 U6645 ( .A1(n2818), .A2(\SB3_23/Component_Function_3/NAND4_in[2] ), 
        .A3(\SB3_23/Component_Function_3/NAND4_in[1] ), .A4(n5255), .ZN(
        \SB3_23/buf_output[3] ) );
  XOR2_X1 U6649 ( .A1(n5092), .A2(\MC_ARK_ARC_1_2/temp6[17] ), .Z(n6540) );
  XOR2_X1 U6650 ( .A1(n5782), .A2(\MC_ARK_ARC_1_2/temp1[17] ), .Z(n5092) );
  XOR2_X1 U6652 ( .A1(n5093), .A2(\MC_ARK_ARC_1_3/temp5[41] ), .Z(\RI1[4][41] ) );
  XOR2_X1 U6653 ( .A1(\MC_ARK_ARC_1_3/temp3[41] ), .A2(
        \MC_ARK_ARC_1_3/temp4[41] ), .Z(n5093) );
  INV_X2 U6655 ( .I(\SB1_1_31/buf_output[2] ), .ZN(\SB2_1_28/i1[9] ) );
  NAND4_X2 U6657 ( .A1(\SB1_1_31/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_31/Component_Function_2/NAND4_in[3] ), .A3(
        \SB1_1_31/Component_Function_2/NAND4_in[1] ), .A4(n6205), .ZN(
        \SB1_1_31/buf_output[2] ) );
  NAND3_X2 U6666 ( .A1(\SB2_1_0/i0[9] ), .A2(\SB2_1_0/i1_5 ), .A3(
        \SB2_1_0/i0[6] ), .ZN(\SB2_1_0/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 U6667 ( .A1(\SB2_3_27/i0[10] ), .A2(n3680), .A3(\SB2_3_27/i0_0 ), 
        .ZN(\SB2_3_27/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U6668 ( .A1(\SB2_1_29/i0_3 ), .A2(\SB2_1_29/i0_4 ), .A3(
        \SB2_1_29/i1[9] ), .ZN(n5968) );
  XOR2_X1 U6669 ( .A1(\RI5[1][167] ), .A2(\RI5[1][11] ), .Z(n5095) );
  INV_X2 U6670 ( .I(\SB1_1_29/buf_output[5] ), .ZN(\SB2_1_29/i1_5 ) );
  NAND4_X2 U6672 ( .A1(\SB1_1_29/Component_Function_5/NAND4_in[2] ), .A2(n5918), .A3(\SB1_1_29/Component_Function_5/NAND4_in[1] ), .A4(
        \SB1_1_29/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_29/buf_output[5] ) );
  NAND3_X2 U6678 ( .A1(\SB2_2_22/i1[9] ), .A2(\SB2_2_22/i0_3 ), .A3(
        \SB2_2_22/i0[6] ), .ZN(\SB2_2_22/Component_Function_3/NAND4_in[0] ) );
  NAND4_X2 U6680 ( .A1(\SB1_1_6/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_6/Component_Function_2/NAND4_in[1] ), .A3(n3234), .A4(n5096), 
        .ZN(\SB1_1_6/buf_output[2] ) );
  NAND3_X2 U6681 ( .A1(\SB1_1_6/i0_3 ), .A2(\SB1_1_6/i0[8] ), .A3(
        \SB1_1_6/i0[9] ), .ZN(n5096) );
  NAND4_X2 U6683 ( .A1(\SB1_2_6/Component_Function_2/NAND4_in[3] ), .A2(n4552), 
        .A3(n4438), .A4(n5097), .ZN(\SB1_2_6/buf_output[2] ) );
  NAND3_X1 U6686 ( .A1(\SB1_2_31/i0[10] ), .A2(\SB1_2_31/i0_0 ), .A3(
        \MC_ARK_ARC_1_1/buf_output[1] ), .ZN(
        \SB1_2_31/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U6688 ( .A1(\SB1_2_7/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_2_7/Component_Function_2/NAND4_in[0] ), .A3(n6042), .A4(n5099), 
        .ZN(\SB1_2_7/buf_output[2] ) );
  NAND3_X2 U6689 ( .A1(\SB1_2_7/i0[9] ), .A2(\SB1_2_7/i0_3 ), .A3(
        \SB1_2_7/i0[8] ), .ZN(n5099) );
  NAND4_X2 U6691 ( .A1(\SB1_3_6/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_3_6/Component_Function_3/NAND4_in[1] ), .A3(n3262), .A4(n5100), 
        .ZN(\SB1_3_6/buf_output[3] ) );
  INV_X2 U6695 ( .I(\SB1_2_12/buf_output[3] ), .ZN(\SB2_2_10/i0[8] ) );
  NAND4_X2 U6700 ( .A1(\SB1_2_12/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_2_12/Component_Function_3/NAND4_in[2] ), .A3(n5185), .A4(n6091), 
        .ZN(\SB1_2_12/buf_output[3] ) );
  NAND2_X2 U6704 ( .A1(\SB2_0_2/i1[9] ), .A2(\SB2_0_2/i0_3 ), .ZN(
        \SB2_0_2/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 U6708 ( .A1(\SB2_3_15/i0_3 ), .A2(\SB1_3_16/buf_output[4] ), .A3(
        \SB2_3_15/i1[9] ), .ZN(\SB2_3_15/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U6710 ( .A1(\SB3_7/Component_Function_2/NAND4_in[1] ), .A2(
        \SB3_7/Component_Function_2/NAND4_in[3] ), .A3(n4727), .A4(
        \SB3_7/Component_Function_2/NAND4_in[0] ), .ZN(\SB3_7/buf_output[2] )
         );
  NAND3_X2 U6712 ( .A1(\SB3_7/i0[10] ), .A2(\SB3_7/i1[9] ), .A3(n4766), .ZN(
        \SB3_7/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U6714 ( .A1(n4489), .A2(n4225), .A3(n5778), .A4(n5101), .ZN(n5122)
         );
  NAND2_X2 U6716 ( .A1(\SB4_29/i0[10] ), .A2(\SB4_29/i0[9] ), .ZN(n5101) );
  NAND4_X2 U6718 ( .A1(\SB3_4/Component_Function_1/NAND4_in[1] ), .A2(
        \SB3_4/Component_Function_1/NAND4_in[3] ), .A3(
        \SB3_4/Component_Function_1/NAND4_in[0] ), .A4(n5102), .ZN(
        \SB3_4/buf_output[1] ) );
  NAND3_X1 U6720 ( .A1(\SB3_4/i0[6] ), .A2(\SB3_4/i0[9] ), .A3(n2910), .ZN(
        n5102) );
  XOR2_X1 U6724 ( .A1(\MC_ARK_ARC_1_3/temp1[162] ), .A2(n5103), .Z(
        \MC_ARK_ARC_1_3/temp5[162] ) );
  XOR2_X1 U6734 ( .A1(\RI5[3][108] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[132] ), 
        .Z(n5103) );
  NAND4_X2 U6737 ( .A1(\SB2_3_18/Component_Function_0/NAND4_in[1] ), .A2(n1082), .A3(\SB2_3_18/Component_Function_0/NAND4_in[0] ), .A4(n5104), .ZN(
        \SB2_3_18/buf_output[0] ) );
  NAND3_X1 U6747 ( .A1(\SB2_3_18/i0_3 ), .A2(\SB2_3_18/i0_0 ), .A3(
        \SB2_3_18/i0[7] ), .ZN(n5104) );
  XOR2_X1 U6748 ( .A1(n2727), .A2(n2726), .Z(\MC_ARK_ARC_1_3/buf_output[146] )
         );
  XOR2_X1 U6750 ( .A1(n2620), .A2(\MC_ARK_ARC_1_3/temp1[146] ), .Z(n2727) );
  NAND4_X2 U6751 ( .A1(\SB1_1_23/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_23/Component_Function_4/NAND4_in[2] ), .A3(
        \SB1_1_23/Component_Function_4/NAND4_in[1] ), .A4(n3532), .ZN(
        \SB1_1_23/buf_output[4] ) );
  NAND4_X2 U6754 ( .A1(\SB1_3_12/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_3_12/Component_Function_1/NAND4_in[1] ), .A3(n5942), .A4(
        \SB1_3_12/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB1_3_12/buf_output[1] ) );
  XOR2_X1 U6761 ( .A1(n3637), .A2(n3636), .Z(\MC_ARK_ARC_1_1/buf_output[170] )
         );
  XOR2_X1 U6762 ( .A1(n5895), .A2(\MC_ARK_ARC_1_1/temp4[170] ), .Z(n3637) );
  XOR2_X1 U6763 ( .A1(\RI5[0][125] ), .A2(\RI5[0][89] ), .Z(
        \MC_ARK_ARC_1_0/temp3[23] ) );
  NAND4_X2 U6764 ( .A1(n2756), .A2(\SB2_1_0/Component_Function_3/NAND4_in[2] ), 
        .A3(\SB2_1_0/Component_Function_3/NAND4_in[0] ), .A4(
        \SB2_1_0/Component_Function_3/NAND4_in[1] ), .ZN(
        \SB2_1_0/buf_output[3] ) );
  NAND4_X2 U6776 ( .A1(\SB2_0_5/Component_Function_3/NAND4_in[3] ), .A2(
        \SB2_0_5/Component_Function_3/NAND4_in[1] ), .A3(n5377), .A4(n6202), 
        .ZN(\SB2_0_5/buf_output[3] ) );
  NAND3_X1 U6777 ( .A1(\SB1_0_11/i0_3 ), .A2(n382), .A3(\SB1_0_11/i1[9] ), 
        .ZN(n1241) );
  XOR2_X1 U6779 ( .A1(\MC_ARK_ARC_1_0/temp6[177] ), .A2(
        \MC_ARK_ARC_1_0/temp5[177] ), .Z(\MC_ARK_ARC_1_0/buf_output[177] ) );
  NAND4_X2 U6780 ( .A1(\SB3_2/Component_Function_3/NAND4_in[1] ), .A2(n1777), 
        .A3(\SB3_2/Component_Function_3/NAND4_in[0] ), .A4(
        \SB3_2/Component_Function_3/NAND4_in[2] ), .ZN(\SB3_2/buf_output[3] )
         );
  BUF_X4 U6783 ( .I(\SB2_1_0/buf_output[5] ), .Z(\RI5[1][191] ) );
  NAND3_X2 U6784 ( .A1(\SB2_1_26/i0[6] ), .A2(\SB2_1_26/i0[10] ), .A3(
        \SB2_1_26/i0_3 ), .ZN(n6273) );
  XOR2_X1 U6788 ( .A1(n5105), .A2(n33), .Z(Ciphertext[188]) );
  NAND4_X2 U6790 ( .A1(n1174), .A2(n3173), .A3(n5301), .A4(n1031), .ZN(n5105)
         );
  NAND3_X2 U6792 ( .A1(\SB2_2_21/i0[6] ), .A2(\SB2_2_21/i0_4 ), .A3(
        \SB2_2_21/i0[9] ), .ZN(n1811) );
  BUF_X4 U6794 ( .I(\MC_ARK_ARC_1_3/buf_output[191] ), .Z(\SB3_0/i0_3 ) );
  XOR2_X1 U6798 ( .A1(n5607), .A2(n5608), .Z(\MC_ARK_ARC_1_3/buf_output[175] )
         );
  XOR2_X1 U6802 ( .A1(\MC_ARK_ARC_1_3/temp1[174] ), .A2(n5106), .Z(n3009) );
  XOR2_X1 U6803 ( .A1(\RI5[3][144] ), .A2(\RI5[3][120] ), .Z(n5106) );
  NAND4_X2 U6808 ( .A1(\SB1_0_16/Component_Function_2/NAND4_in[1] ), .A2(n4189), .A3(n673), .A4(\SB1_0_16/Component_Function_2/NAND4_in[0] ), .ZN(
        \SB1_0_16/buf_output[2] ) );
  XOR2_X1 U6813 ( .A1(n5107), .A2(\MC_ARK_ARC_1_3/temp2[163] ), .Z(
        \MC_ARK_ARC_1_3/temp5[163] ) );
  XOR2_X1 U6817 ( .A1(\RI5[3][163] ), .A2(\RI5[3][157] ), .Z(n5107) );
  XOR2_X1 U6818 ( .A1(\MC_ARK_ARC_1_1/temp6[105] ), .A2(
        \MC_ARK_ARC_1_1/temp5[105] ), .Z(\MC_ARK_ARC_1_1/buf_output[105] ) );
  XOR2_X1 U6820 ( .A1(\RI5[1][79] ), .A2(\RI5[1][103] ), .Z(
        \MC_ARK_ARC_1_1/temp2[133] ) );
  NAND4_X2 U6821 ( .A1(\SB2_1_0/Component_Function_2/NAND4_in[3] ), .A2(
        \SB2_1_0/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_1_0/Component_Function_2/NAND4_in[2] ), .A4(n5108), .ZN(
        \SB2_1_0/buf_output[2] ) );
  NAND4_X2 U6824 ( .A1(n4617), .A2(\SB3_0/Component_Function_5/NAND4_in[3] ), 
        .A3(n6510), .A4(\SB3_0/Component_Function_5/NAND4_in[1] ), .ZN(
        \SB3_0/buf_output[5] ) );
  NAND4_X2 U6825 ( .A1(\SB2_0_11/Component_Function_5/NAND4_in[0] ), .A2(n780), 
        .A3(\SB2_0_11/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_0_11/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB2_0_11/buf_output[5] ) );
  NAND4_X2 U6828 ( .A1(\SB1_0_11/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_0_11/Component_Function_3/NAND4_in[0] ), .A3(n6196), .A4(
        \SB1_0_11/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_0_11/buf_output[3] ) );
  XOR2_X1 U6839 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[65] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[29] ), .Z(\MC_ARK_ARC_1_2/temp3[155] )
         );
  NAND4_X2 U6840 ( .A1(\SB2_1_21/Component_Function_5/NAND4_in[2] ), .A2(n856), 
        .A3(n2439), .A4(\SB2_1_21/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_1_21/buf_output[5] ) );
  NAND4_X2 U6846 ( .A1(n933), .A2(n5110), .A3(n6045), .A4(
        \SB1_2_27/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_2_27/buf_output[5] ) );
  NAND3_X2 U6848 ( .A1(\SB2_2_27/i0_3 ), .A2(\SB2_2_27/i1[9] ), .A3(
        \SB1_2_28/buf_output[4] ), .ZN(n5109) );
  XOR2_X1 U6849 ( .A1(\RI5[3][143] ), .A2(n5503), .Z(
        \MC_ARK_ARC_1_3/temp2[173] ) );
  NAND3_X2 U6850 ( .A1(\SB1_3_11/i0_4 ), .A2(\SB1_3_11/i0_0 ), .A3(n2908), 
        .ZN(n3949) );
  XOR2_X1 U6862 ( .A1(\MC_ARK_ARC_1_3/temp5[172] ), .A2(n5111), .Z(
        \MC_ARK_ARC_1_3/buf_output[172] ) );
  XOR2_X1 U6871 ( .A1(\MC_ARK_ARC_1_3/temp3[172] ), .A2(
        \MC_ARK_ARC_1_3/temp4[172] ), .Z(n5111) );
  XOR2_X1 U6873 ( .A1(\MC_ARK_ARC_1_2/temp3[155] ), .A2(n5112), .Z(n6027) );
  XOR2_X1 U6874 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[125] ), .A2(\RI5[2][101] ), 
        .Z(n5112) );
  XOR2_X1 U6877 ( .A1(n3300), .A2(n5113), .Z(n4133) );
  XOR2_X1 U6878 ( .A1(\RI5[1][53] ), .A2(\RI5[1][59] ), .Z(n5113) );
  NAND3_X2 U6882 ( .A1(\SB2_3_9/i0_0 ), .A2(\SB2_3_9/i0_4 ), .A3(
        \SB2_3_9/i1_5 ), .ZN(n5114) );
  NAND3_X2 U6883 ( .A1(\SB2_1_14/i0_4 ), .A2(\SB2_1_14/i1_7 ), .A3(
        \SB2_1_14/i0[8] ), .ZN(\SB2_1_14/Component_Function_1/NAND4_in[3] ) );
  XOR2_X1 U6887 ( .A1(n4421), .A2(n5115), .Z(\MC_ARK_ARC_1_2/buf_output[111] )
         );
  XOR2_X1 U6888 ( .A1(\MC_ARK_ARC_1_2/temp1[111] ), .A2(
        \MC_ARK_ARC_1_2/temp4[111] ), .Z(n5115) );
  NAND3_X2 U6892 ( .A1(\SB1_2_11/i0_4 ), .A2(\SB1_2_11/i0_3 ), .A3(
        \SB1_2_11/i1[9] ), .ZN(n5116) );
  NAND3_X1 U6898 ( .A1(\SB4_29/i0[9] ), .A2(\SB4_29/i0[6] ), .A3(\SB4_29/i1_5 ), .ZN(n5117) );
  NAND4_X2 U6899 ( .A1(\SB2_3_7/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_7/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_3_7/Component_Function_4/NAND4_in[3] ), .A4(n5118), .ZN(
        \SB2_3_7/buf_output[4] ) );
  NAND3_X2 U6907 ( .A1(\SB2_3_7/i0[9] ), .A2(\SB2_3_7/i0[10] ), .A3(
        \SB2_3_7/i0_3 ), .ZN(n5118) );
  XOR2_X1 U6908 ( .A1(\MC_ARK_ARC_1_1/temp4[157] ), .A2(n5119), .Z(n1641) );
  XOR2_X1 U6911 ( .A1(\RI5[1][127] ), .A2(\RI5[1][103] ), .Z(n5119) );
  NAND3_X2 U6912 ( .A1(\SB1_1_15/i0_4 ), .A2(\SB1_1_15/i1[9] ), .A3(
        \SB1_1_15/i1_5 ), .ZN(\SB1_1_15/Component_Function_4/NAND4_in[3] ) );
  XOR2_X1 U6913 ( .A1(n5120), .A2(n217), .Z(Ciphertext[51]) );
  NAND4_X2 U6914 ( .A1(\SB4_23/Component_Function_3/NAND4_in[3] ), .A2(
        \SB4_23/Component_Function_3/NAND4_in[1] ), .A3(
        \SB4_23/Component_Function_3/NAND4_in[0] ), .A4(
        \SB4_23/Component_Function_3/NAND4_in[2] ), .ZN(n5120) );
  NAND3_X2 U6915 ( .A1(\SB2_3_28/i0[8] ), .A2(\SB2_3_28/i1_5 ), .A3(
        \SB2_3_28/i3[0] ), .ZN(\SB2_3_28/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 U6916 ( .A1(\SB2_0_22/i0_0 ), .A2(\SB2_0_22/i0_3 ), .A3(
        \SB2_0_22/i0[7] ), .ZN(n2366) );
  XOR2_X1 U6919 ( .A1(n5121), .A2(n237), .Z(Ciphertext[46]) );
  NAND4_X2 U6921 ( .A1(\SB4_24/Component_Function_4/NAND4_in[0] ), .A2(n6198), 
        .A3(\SB4_24/Component_Function_4/NAND4_in[3] ), .A4(n4545), .ZN(n5121)
         );
  NAND3_X2 U6925 ( .A1(\SB2_0_30/i0[10] ), .A2(\SB2_0_30/i1[9] ), .A3(
        \SB2_0_30/i1_7 ), .ZN(\SB2_0_30/Component_Function_3/NAND4_in[2] ) );
  XOR2_X1 U6927 ( .A1(\RI5[1][50] ), .A2(\RI5[1][44] ), .Z(
        \MC_ARK_ARC_1_1/temp1[50] ) );
  XOR2_X1 U6928 ( .A1(n5122), .A2(n48), .Z(Ciphertext[12]) );
  INV_X2 U6931 ( .I(\SB1_2_19/buf_output[2] ), .ZN(\SB2_2_16/i1[9] ) );
  NAND4_X2 U6935 ( .A1(\SB1_2_19/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_2_19/Component_Function_2/NAND4_in[3] ), .A3(n4499), .A4(
        \SB1_2_19/Component_Function_2/NAND4_in[1] ), .ZN(
        \SB1_2_19/buf_output[2] ) );
  NAND4_X2 U6936 ( .A1(\SB2_3_12/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_3_12/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_3_12/Component_Function_4/NAND4_in[0] ), .A4(n4000), .ZN(
        \SB2_3_12/buf_output[4] ) );
  XOR2_X1 U6939 ( .A1(n5123), .A2(n189), .Z(Ciphertext[57]) );
  NAND4_X2 U6940 ( .A1(n4579), .A2(\SB4_22/Component_Function_3/NAND4_in[0] ), 
        .A3(\SB4_22/Component_Function_3/NAND4_in[2] ), .A4(n5701), .ZN(n5123)
         );
  NAND4_X2 U6941 ( .A1(\SB2_1_5/Component_Function_2/NAND4_in[0] ), .A2(n5365), 
        .A3(n5364), .A4(\SB2_1_5/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB2_1_5/buf_output[2] ) );
  BUF_X4 U6944 ( .I(\RI3[0][131] ), .Z(\SB2_0_10/i0_3 ) );
  NAND3_X1 U6949 ( .A1(\SB2_3_10/i0_3 ), .A2(\SB2_3_10/i0[9] ), .A3(
        \SB2_3_10/i0[8] ), .ZN(\SB2_3_10/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U6950 ( .A1(\SB1_0_2/i0[10] ), .A2(\SB1_0_2/i0_0 ), .A3(
        \SB1_0_2/i0[6] ), .ZN(\SB1_0_2/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U6953 ( .A1(\SB1_2_25/Component_Function_2/NAND4_in[1] ), .A2(n4444), .A3(\SB1_2_25/Component_Function_2/NAND4_in[0] ), .A4(
        \SB1_2_25/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB1_2_25/buf_output[2] ) );
  XOR2_X1 U6959 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[183] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[27] ), .Z(\MC_ARK_ARC_1_2/temp3[117] )
         );
  NAND4_X2 U6960 ( .A1(\SB3_27/Component_Function_2/NAND4_in[0] ), .A2(n590), 
        .A3(n6404), .A4(n2976), .ZN(\SB3_27/buf_output[2] ) );
  XOR2_X1 U6961 ( .A1(n5124), .A2(n9), .Z(Ciphertext[54]) );
  NAND4_X2 U6963 ( .A1(\SB4_22/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_22/Component_Function_0/NAND4_in[1] ), .A3(
        \SB4_22/Component_Function_0/NAND4_in[3] ), .A4(
        \SB4_22/Component_Function_0/NAND4_in[0] ), .ZN(n5124) );
  XOR2_X1 U6964 ( .A1(n5611), .A2(n4726), .Z(\MC_ARK_ARC_1_2/buf_output[117] )
         );
  INV_X1 U6966 ( .I(\SB3_27/buf_output[5] ), .ZN(\SB4_27/i1_5 ) );
  NAND4_X2 U6968 ( .A1(n2723), .A2(\SB3_27/Component_Function_5/NAND4_in[3] ), 
        .A3(n6180), .A4(\SB3_27/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB3_27/buf_output[5] ) );
  NAND3_X2 U6973 ( .A1(\SB1_3_12/i0[10] ), .A2(\SB1_3_12/i0[6] ), .A3(
        \SB1_3_12/i0_0 ), .ZN(\SB1_3_12/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U6974 ( .A1(\SB3_11/i0_0 ), .A2(\SB3_11/i0_4 ), .A3(n582), .ZN(
        n3057) );
  XOR2_X1 U6975 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[179] ), .A2(\RI5[0][53] ), 
        .Z(n1184) );
  NAND4_X2 U6976 ( .A1(\SB2_3_10/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_3_10/Component_Function_3/NAND4_in[3] ), .A3(n6431), .A4(
        \SB2_3_10/Component_Function_3/NAND4_in[0] ), .ZN(
        \SB2_3_10/buf_output[3] ) );
  XOR2_X1 U6979 ( .A1(n1450), .A2(n2028), .Z(\MC_ARK_ARC_1_0/buf_output[126] )
         );
  NAND4_X2 U6983 ( .A1(\SB3_22/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_22/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_22/Component_Function_3/NAND4_in[2] ), .A4(n2215), .ZN(
        \SB3_22/buf_output[3] ) );
  NAND3_X1 U6986 ( .A1(n3653), .A2(\SB4_10/i0_3 ), .A3(\SB4_10/i0[6] ), .ZN(
        n4283) );
  XOR2_X1 U6990 ( .A1(n727), .A2(\MC_ARK_ARC_1_1/temp5[90] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[90] ) );
  XOR2_X1 U7000 ( .A1(\MC_ARK_ARC_1_3/temp1[124] ), .A2(
        \MC_ARK_ARC_1_3/temp2[124] ), .Z(\MC_ARK_ARC_1_3/temp5[124] ) );
  INV_X2 U7001 ( .I(n5125), .ZN(\MC_ARK_ARC_1_3/buf_output[110] ) );
  XNOR2_X1 U7003 ( .A1(n4740), .A2(n4739), .ZN(n5125) );
  NAND4_X2 U7008 ( .A1(\SB2_0_4/Component_Function_5/NAND4_in[2] ), .A2(n3004), 
        .A3(n1409), .A4(\SB2_0_4/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_0_4/buf_output[5] ) );
  XOR2_X1 U7014 ( .A1(n5126), .A2(n148), .Z(Ciphertext[141]) );
  NAND4_X2 U7016 ( .A1(\SB4_8/Component_Function_3/NAND4_in[2] ), .A2(n6369), 
        .A3(n6514), .A4(\SB4_8/Component_Function_3/NAND4_in[3] ), .ZN(n5126)
         );
  INV_X4 U7019 ( .I(\SB2_0_24/i0[7] ), .ZN(\RI3[0][46] ) );
  NAND3_X1 U7020 ( .A1(\RI3[0][43] ), .A2(\SB2_0_24/i0[7] ), .A3(
        \SB2_0_24/i0[8] ), .ZN(n5933) );
  NOR2_X2 U7021 ( .A1(n5128), .A2(n5127), .ZN(\SB2_0_24/i0[7] ) );
  NAND2_X2 U7022 ( .A1(\SB1_0_25/Component_Function_4/NAND4_in[2] ), .A2(n2554), .ZN(n5127) );
  NAND2_X1 U7025 ( .A1(\SB1_0_25/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_0_25/Component_Function_4/NAND4_in[1] ), .ZN(n5128) );
  XOR2_X1 U7029 ( .A1(\MC_ARK_ARC_1_3/temp5[82] ), .A2(n5129), .Z(
        \MC_ARK_ARC_1_3/buf_output[82] ) );
  XOR2_X1 U7032 ( .A1(\MC_ARK_ARC_1_3/temp3[82] ), .A2(
        \MC_ARK_ARC_1_3/temp4[82] ), .Z(n5129) );
  NAND4_X2 U7033 ( .A1(n4058), .A2(\SB3_18/Component_Function_2/NAND4_in[0] ), 
        .A3(\SB3_18/Component_Function_2/NAND4_in[2] ), .A4(n5130), .ZN(
        \SB3_18/buf_output[2] ) );
  NAND3_X1 U7042 ( .A1(\SB3_18/i0_0 ), .A2(\SB3_18/i0_4 ), .A3(\SB3_18/i1_5 ), 
        .ZN(n5130) );
  XOR2_X1 U7043 ( .A1(n5131), .A2(n47), .Z(Ciphertext[95]) );
  XOR2_X1 U7044 ( .A1(\MC_ARK_ARC_1_3/temp5[149] ), .A2(
        \MC_ARK_ARC_1_3/temp6[149] ), .Z(\MC_ARK_ARC_1_3/buf_output[149] ) );
  XOR2_X1 U7045 ( .A1(\MC_ARK_ARC_1_3/temp1[149] ), .A2(
        \MC_ARK_ARC_1_3/temp2[149] ), .Z(\MC_ARK_ARC_1_3/temp5[149] ) );
  BUF_X4 U7046 ( .I(\MC_ARK_ARC_1_3/buf_output[155] ), .Z(\RI1[4][155] ) );
  NAND3_X1 U7057 ( .A1(\SB4_3/i0_4 ), .A2(\SB3_6/buf_output[2] ), .A3(
        \SB4_3/i0_3 ), .ZN(n5133) );
  XOR2_X1 U7058 ( .A1(n5134), .A2(n180), .Z(Ciphertext[68]) );
  NAND4_X2 U7065 ( .A1(\SB4_20/Component_Function_2/NAND4_in[0] ), .A2(n6348), 
        .A3(\SB4_20/Component_Function_2/NAND4_in[2] ), .A4(
        \SB4_20/Component_Function_2/NAND4_in[1] ), .ZN(n5134) );
  NAND3_X1 U7066 ( .A1(\SB4_21/i0_4 ), .A2(\SB4_21/i0[9] ), .A3(\SB4_21/i0[6] ), .ZN(\SB4_21/Component_Function_5/NAND4_in[3] ) );
  NAND4_X2 U7067 ( .A1(\SB2_3_10/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_10/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_3_10/Component_Function_5/NAND4_in[0] ), .A4(n5135), .ZN(
        \SB2_3_10/buf_output[5] ) );
  NAND3_X2 U7068 ( .A1(\SB2_3_10/i0_4 ), .A2(\SB2_3_10/i0[6] ), .A3(
        \SB2_3_10/i0[9] ), .ZN(n5135) );
  NAND3_X2 U7069 ( .A1(\SB2_3_0/i0_3 ), .A2(n5513), .A3(\SB2_3_0/i1_7 ), .ZN(
        \SB2_3_0/Component_Function_1/NAND4_in[1] ) );
  NAND3_X2 U7072 ( .A1(\SB2_2_29/i0_3 ), .A2(\SB2_2_29/i0[8] ), .A3(
        \SB2_2_29/i0[9] ), .ZN(n6084) );
  XOR2_X1 U7073 ( .A1(\MC_ARK_ARC_1_1/temp6[4] ), .A2(n5137), .Z(
        \MC_ARK_ARC_1_1/buf_output[4] ) );
  XOR2_X1 U7074 ( .A1(\MC_ARK_ARC_1_1/temp2[4] ), .A2(
        \MC_ARK_ARC_1_1/temp1[4] ), .Z(n5137) );
  XOR2_X1 U7076 ( .A1(n5138), .A2(\MC_ARK_ARC_1_2/temp5[142] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[142] ) );
  XOR2_X1 U7077 ( .A1(\MC_ARK_ARC_1_2/temp4[142] ), .A2(
        \MC_ARK_ARC_1_2/temp3[142] ), .Z(n5138) );
  NAND4_X2 U7080 ( .A1(\SB1_2_30/Component_Function_5/NAND4_in[2] ), .A2(n3981), .A3(n2724), .A4(\SB1_2_30/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_2_30/buf_output[5] ) );
  NAND4_X2 U7081 ( .A1(n4195), .A2(\SB2_1_27/Component_Function_5/NAND4_in[0] ), .A3(\SB2_1_27/Component_Function_5/NAND4_in[3] ), .A4(n5139), .ZN(
        \SB2_1_27/buf_output[5] ) );
  NAND3_X2 U7082 ( .A1(\SB2_1_27/i0_0 ), .A2(\SB2_1_27/i0[10] ), .A3(
        \SB2_1_27/i0[6] ), .ZN(n5139) );
  NAND4_X2 U7084 ( .A1(\SB3_14/Component_Function_5/NAND4_in[1] ), .A2(n1875), 
        .A3(\SB3_14/Component_Function_5/NAND4_in[0] ), .A4(n5140), .ZN(
        \SB3_14/buf_output[5] ) );
  NAND3_X2 U7095 ( .A1(\SB2_0_4/i0_3 ), .A2(\SB2_0_4/i0_0 ), .A3(\RI3[0][166] ), .ZN(n5141) );
  NAND4_X2 U7096 ( .A1(\SB2_0_11/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_0_11/Component_Function_3/NAND4_in[0] ), .A3(n3693), .A4(n5142), 
        .ZN(\SB2_0_11/buf_output[3] ) );
  NAND3_X1 U7097 ( .A1(\SB2_0_11/i0_0 ), .A2(\SB2_0_11/i0_3 ), .A3(
        \SB2_0_11/i0_4 ), .ZN(n5142) );
  NAND3_X1 U7098 ( .A1(\SB2_3_24/i0[9] ), .A2(\SB2_3_24/i0_3 ), .A3(
        \SB1_3_26/buf_output[3] ), .ZN(n5654) );
  NAND3_X2 U7105 ( .A1(\SB3_5/i0[9] ), .A2(\SB3_5/i0_3 ), .A3(\SB3_5/i0[10] ), 
        .ZN(n5143) );
  NAND4_X2 U7108 ( .A1(\SB2_0_13/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_0_13/Component_Function_0/NAND4_in[1] ), .A3(n3171), .A4(
        \SB2_0_13/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_0_13/buf_output[0] ) );
  NAND3_X2 U7111 ( .A1(\SB1_3_17/i0_4 ), .A2(\SB1_3_17/i0_0 ), .A3(
        \SB1_3_17/i1_5 ), .ZN(n5144) );
  NAND4_X2 U7113 ( .A1(\SB1_1_14/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_1_14/Component_Function_2/NAND4_in[3] ), .A3(n5201), .A4(n5145), 
        .ZN(\SB1_1_14/buf_output[2] ) );
  NAND4_X2 U7114 ( .A1(\SB2_3_1/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_3_1/Component_Function_0/NAND4_in[0] ), .A3(
        \SB2_3_1/Component_Function_0/NAND4_in[2] ), .A4(n5147), .ZN(
        \SB2_3_1/buf_output[0] ) );
  NAND3_X1 U7118 ( .A1(\SB2_3_1/i0_3 ), .A2(\SB2_3_1/i0_0 ), .A3(
        \SB2_3_1/i0[7] ), .ZN(n5147) );
  INV_X2 U7119 ( .I(\SB1_1_20/buf_output[3] ), .ZN(\SB2_1_18/i0[8] ) );
  XOR2_X1 U7120 ( .A1(n5148), .A2(n1351), .Z(\MC_ARK_ARC_1_3/buf_output[48] )
         );
  XOR2_X1 U7121 ( .A1(\MC_ARK_ARC_1_3/temp2[48] ), .A2(
        \MC_ARK_ARC_1_3/temp4[48] ), .Z(n5148) );
  XOR2_X1 U7122 ( .A1(n2603), .A2(n5149), .Z(\MC_ARK_ARC_1_1/buf_output[130] )
         );
  XOR2_X1 U7129 ( .A1(n3543), .A2(\MC_ARK_ARC_1_1/temp2[130] ), .Z(n5149) );
  INV_X1 U7136 ( .I(\SB1_3_15/buf_output[3] ), .ZN(\SB2_3_13/i0[8] ) );
  NAND4_X2 U7137 ( .A1(\SB1_3_15/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_3_15/Component_Function_3/NAND4_in[0] ), .A3(n5920), .A4(n1037), 
        .ZN(\SB1_3_15/buf_output[3] ) );
  BUF_X4 U7141 ( .I(\MC_ARK_ARC_1_2/buf_output[62] ), .Z(\SB1_3_21/i0_0 ) );
  XOR2_X1 U7144 ( .A1(n5150), .A2(\MC_ARK_ARC_1_0/temp2[177] ), .Z(
        \MC_ARK_ARC_1_0/temp5[177] ) );
  NAND4_X2 U7150 ( .A1(\SB2_1_31/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_1_31/Component_Function_4/NAND4_in[2] ), .A3(n3792), .A4(n5151), 
        .ZN(\SB2_1_31/buf_output[4] ) );
  NAND3_X2 U7151 ( .A1(\SB1_2_24/i0[9] ), .A2(\SB1_2_24/i0[6] ), .A3(
        \SB1_2_24/i0_4 ), .ZN(n5152) );
  XOR2_X1 U7155 ( .A1(n5153), .A2(\MC_ARK_ARC_1_2/temp1[171] ), .Z(n2819) );
  XOR2_X1 U7157 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[117] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[141] ), .Z(n5153) );
  BUF_X4 U7160 ( .I(\SB2_2_22/buf_output[5] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[59] ) );
  XOR2_X1 U7161 ( .A1(n3454), .A2(\MC_ARK_ARC_1_0/temp5[68] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[68] ) );
  NAND3_X1 U7165 ( .A1(\SB4_2/i0_0 ), .A2(\SB4_2/i0[8] ), .A3(\SB4_2/i0[9] ), 
        .ZN(\SB4_2/Component_Function_4/NAND4_in[0] ) );
  BUF_X4 U7167 ( .I(\SB1_3_3/buf_output[3] ), .Z(\SB2_3_1/i0[10] ) );
  NAND4_X2 U7174 ( .A1(\SB1_1_20/Component_Function_5/NAND4_in[1] ), .A2(n5299), .A3(n1944), .A4(\SB1_1_20/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_20/buf_output[5] ) );
  NAND4_X2 U7183 ( .A1(\SB1_2_13/Component_Function_5/NAND4_in[2] ), .A2(n1523), .A3(\SB1_2_13/Component_Function_5/NAND4_in[0] ), .A4(
        \SB1_2_13/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB1_2_13/buf_output[5] ) );
  NAND3_X2 U7184 ( .A1(\SB1_2_13/i0_4 ), .A2(\SB1_2_13/i0[6] ), .A3(
        \SB1_2_13/i0[9] ), .ZN(\SB1_2_13/Component_Function_5/NAND4_in[3] ) );
  XOR2_X1 U7189 ( .A1(\SB2_1_16/buf_output[1] ), .A2(\RI5[1][91] ), .Z(
        \MC_ARK_ARC_1_1/temp2[145] ) );
  XOR2_X1 U7191 ( .A1(n5155), .A2(n122), .Z(Ciphertext[92]) );
  NAND4_X2 U7193 ( .A1(\SB4_16/Component_Function_2/NAND4_in[0] ), .A2(
        \SB4_16/Component_Function_2/NAND4_in[3] ), .A3(n4340), .A4(
        \SB4_16/Component_Function_2/NAND4_in[2] ), .ZN(n5155) );
  NAND4_X2 U7196 ( .A1(\SB1_2_7/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_2_7/Component_Function_5/NAND4_in[1] ), .A3(n5180), .A4(n5939), 
        .ZN(\SB1_2_7/buf_output[5] ) );
  XOR2_X1 U7197 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[36] ), .A2(\RI5[3][72] ), 
        .Z(n5156) );
  XOR2_X1 U7198 ( .A1(\MC_ARK_ARC_1_3/temp3[157] ), .A2(
        \MC_ARK_ARC_1_3/temp4[157] ), .Z(\MC_ARK_ARC_1_3/temp6[157] ) );
  XOR2_X1 U7205 ( .A1(\RI5[2][159] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[153] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[159] ) );
  NAND3_X1 U7206 ( .A1(\SB4_21/i0_4 ), .A2(\SB3_24/buf_output[2] ), .A3(
        \SB4_21/i0_3 ), .ZN(\SB4_21/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U7217 ( .A1(\MC_ARK_ARC_1_1/temp5[28] ), .A2(
        \MC_ARK_ARC_1_1/temp6[28] ), .Z(\MC_ARK_ARC_1_1/buf_output[28] ) );
  NAND4_X2 U7222 ( .A1(\SB1_3_31/Component_Function_4/NAND4_in[0] ), .A2(n6466), .A3(\SB1_3_31/Component_Function_4/NAND4_in[1] ), .A4(
        \SB1_3_31/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB1_3_31/buf_output[4] ) );
  NAND4_X2 U7223 ( .A1(n1099), .A2(n3409), .A3(
        \SB2_2_22/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_2_22/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_2_22/buf_output[1] ) );
  NAND4_X2 U7224 ( .A1(\SB2_1_29/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_1_29/Component_Function_4/NAND4_in[0] ), .A3(n5304), .A4(
        \SB2_1_29/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_1_29/buf_output[4] ) );
  XOR2_X1 U7231 ( .A1(\MC_ARK_ARC_1_1/temp3[112] ), .A2(
        \MC_ARK_ARC_1_1/temp4[112] ), .Z(n2798) );
  XOR2_X1 U7232 ( .A1(n5158), .A2(n5157), .Z(n5168) );
  XOR2_X1 U7233 ( .A1(\RI5[3][32] ), .A2(\RI5[3][158] ), .Z(n5157) );
  XOR2_X1 U7234 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[152] ), .A2(\RI5[3][68] ), 
        .Z(n5158) );
  NAND4_X2 U7235 ( .A1(n1445), .A2(\SB1_1_15/Component_Function_1/NAND4_in[1] ), .A3(\SB1_1_15/Component_Function_1/NAND4_in[0] ), .A4(n5159), .ZN(
        \SB1_1_15/buf_output[1] ) );
  NAND3_X2 U7237 ( .A1(\SB1_1_15/i0_4 ), .A2(\SB1_1_15/i0[8] ), .A3(
        \SB1_1_15/i1_7 ), .ZN(n5159) );
  XOR2_X1 U7244 ( .A1(\MC_ARK_ARC_1_3/temp4[102] ), .A2(n5161), .Z(
        \MC_ARK_ARC_1_3/temp6[102] ) );
  XOR2_X1 U7245 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[168] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[12] ), .Z(n5161) );
  NAND3_X2 U7247 ( .A1(\SB2_1_11/i0[6] ), .A2(\SB2_1_11/i0_0 ), .A3(
        \SB2_1_11/i0[10] ), .ZN(n5162) );
  NAND4_X2 U7254 ( .A1(n1766), .A2(\SB1_1_23/Component_Function_2/NAND4_in[1] ), .A3(n2868), .A4(n5163), .ZN(\SB1_1_23/buf_output[2] ) );
  NAND3_X2 U7257 ( .A1(\SB1_1_23/i0[10] ), .A2(\SB1_1_23/i1[9] ), .A3(
        \SB1_1_23/i1_5 ), .ZN(n5163) );
  NAND3_X2 U7259 ( .A1(\SB2_1_20/i0_4 ), .A2(\SB2_1_20/i0_3 ), .A3(
        \SB2_1_20/i1[9] ), .ZN(n2890) );
  XOR2_X1 U7260 ( .A1(n6105), .A2(n5164), .Z(\MC_ARK_ARC_1_3/temp5[50] ) );
  XOR2_X1 U7261 ( .A1(\RI5[3][188] ), .A2(\RI5[3][50] ), .Z(n5164) );
  XOR2_X1 U7262 ( .A1(n5165), .A2(n2467), .Z(n1568) );
  XOR2_X1 U7263 ( .A1(\RI5[1][81] ), .A2(\RI5[1][57] ), .Z(n5165) );
  NAND3_X2 U7266 ( .A1(\SB1_2_14/i1_5 ), .A2(\SB1_2_14/i0[8] ), .A3(
        \SB1_2_14/i3[0] ), .ZN(\SB1_2_14/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U7273 ( .A1(n5340), .A2(n5166), .Z(\MC_ARK_ARC_1_1/buf_output[131] )
         );
  XOR2_X1 U7277 ( .A1(\MC_ARK_ARC_1_1/temp3[131] ), .A2(n3443), .Z(n5166) );
  XOR2_X1 U7278 ( .A1(n6505), .A2(n6303), .Z(\MC_ARK_ARC_1_1/temp5[101] ) );
  XOR2_X1 U7281 ( .A1(n5168), .A2(n5167), .Z(\MC_ARK_ARC_1_3/buf_output[158] )
         );
  XOR2_X1 U7284 ( .A1(n1933), .A2(\MC_ARK_ARC_1_3/temp4[158] ), .Z(n5167) );
  XOR2_X1 U7285 ( .A1(\MC_ARK_ARC_1_2/temp1[42] ), .A2(n5169), .Z(n4306) );
  XOR2_X1 U7287 ( .A1(\RI5[2][12] ), .A2(\RI5[2][180] ), .Z(n5169) );
  NAND3_X1 U7298 ( .A1(\SB4_21/i0_4 ), .A2(\SB3_24/buf_output[2] ), .A3(
        \SB4_21/i1_5 ), .ZN(n5170) );
  XOR2_X1 U7299 ( .A1(\RI5[2][51] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[45] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[51] ) );
  XOR2_X1 U7300 ( .A1(n5171), .A2(n15), .Z(Ciphertext[179]) );
  NAND4_X2 U7301 ( .A1(\SB4_2/Component_Function_5/NAND4_in[2] ), .A2(
        \SB4_2/Component_Function_5/NAND4_in[3] ), .A3(n5194), .A4(
        \SB4_2/Component_Function_5/NAND4_in[0] ), .ZN(n5171) );
  XOR2_X1 U7302 ( .A1(n3806), .A2(\MC_ARK_ARC_1_3/temp6[177] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[177] ) );
  NAND4_X2 U7305 ( .A1(\SB2_3_26/Component_Function_2/NAND4_in[0] ), .A2(n5996), .A3(\SB2_3_26/Component_Function_2/NAND4_in[1] ), .A4(n4628), .ZN(
        \SB2_3_26/buf_output[2] ) );
  NAND3_X2 U7306 ( .A1(\SB1_3_31/i0[7] ), .A2(\SB1_3_31/i0_3 ), .A3(
        \SB1_3_31/i0_0 ), .ZN(n3555) );
  NAND4_X2 U7312 ( .A1(\SB2_0_8/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_8/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_0_8/Component_Function_5/NAND4_in[0] ), .A4(n5173), .ZN(
        \SB2_0_8/buf_output[5] ) );
  NAND3_X2 U7315 ( .A1(\SB2_0_8/i0[6] ), .A2(\SB2_0_8/i0_0 ), .A3(
        \SB2_0_8/i0[10] ), .ZN(n5173) );
  NAND3_X2 U7319 ( .A1(\SB2_2_28/i0[10] ), .A2(\SB2_2_28/i0_3 ), .A3(
        \SB2_2_28/i0[6] ), .ZN(n5174) );
  NAND4_X2 U7320 ( .A1(\SB2_1_29/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_1_29/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_1_29/Component_Function_2/NAND4_in[1] ), .A4(n5175), .ZN(
        \SB2_1_29/buf_output[2] ) );
  NAND3_X1 U7321 ( .A1(\SB2_1_29/i0_0 ), .A2(\SB2_1_29/i0_4 ), .A3(
        \SB2_1_29/i1_5 ), .ZN(n5175) );
  XOR2_X1 U7324 ( .A1(n1419), .A2(n5176), .Z(n2939) );
  XOR2_X1 U7330 ( .A1(\RI5[1][5] ), .A2(n3650), .Z(n5176) );
  XOR2_X1 U7332 ( .A1(n5177), .A2(\MC_ARK_ARC_1_1/temp4[14] ), .Z(
        \MC_ARK_ARC_1_1/temp6[14] ) );
  XOR2_X1 U7333 ( .A1(\RI5[1][116] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[80] ), 
        .Z(n5177) );
  XOR2_X1 U7334 ( .A1(\RI5[1][128] ), .A2(\RI5[1][134] ), .Z(
        \MC_ARK_ARC_1_1/temp1[134] ) );
  XOR2_X1 U7336 ( .A1(\MC_ARK_ARC_1_2/temp5[164] ), .A2(n5178), .Z(
        \MC_ARK_ARC_1_2/buf_output[164] ) );
  XOR2_X1 U7339 ( .A1(n3382), .A2(n3381), .Z(n5178) );
  NAND3_X2 U7340 ( .A1(\SB2_1_27/i0[9] ), .A2(\SB2_1_27/i0_3 ), .A3(
        \SB2_1_27/i0[10] ), .ZN(n5179) );
  BUF_X4 U7342 ( .I(\SB2_2_3/buf_output[2] ), .Z(\RI5[2][188] ) );
  XOR2_X1 U7343 ( .A1(\MC_ARK_ARC_1_1/temp6[134] ), .A2(n4708), .Z(n3686) );
  XOR2_X1 U7344 ( .A1(\MC_ARK_ARC_1_1/temp4[134] ), .A2(
        \MC_ARK_ARC_1_1/temp3[134] ), .Z(\MC_ARK_ARC_1_1/temp6[134] ) );
  XOR2_X1 U7346 ( .A1(\MC_ARK_ARC_1_0/temp6[125] ), .A2(n5181), .Z(
        \MC_ARK_ARC_1_0/buf_output[125] ) );
  XOR2_X1 U7351 ( .A1(\MC_ARK_ARC_1_0/temp1[125] ), .A2(n2278), .Z(n5181) );
  NAND3_X2 U7354 ( .A1(\SB1_2_22/i0_3 ), .A2(\SB1_2_22/i1[9] ), .A3(
        \SB1_2_22/i0[6] ), .ZN(\SB1_2_22/Component_Function_3/NAND4_in[0] ) );
  NAND4_X2 U7358 ( .A1(\SB2_2_22/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_2_22/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_2_22/Component_Function_4/NAND4_in[1] ), .A4(n5182), .ZN(
        \SB2_2_22/buf_output[4] ) );
  NAND3_X1 U7359 ( .A1(\SB1_1_27/buf_output[1] ), .A2(\SB1_1_24/buf_output[4] ), .A3(\SB1_1_28/buf_output[0] ), .ZN(n5183) );
  NAND3_X1 U7361 ( .A1(\SB1_1_27/i0_3 ), .A2(\SB1_1_27/i0[8] ), .A3(
        \SB1_1_27/i1_7 ), .ZN(\SB1_1_27/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U7363 ( .A1(n4287), .A2(n5184), .Z(\MC_ARK_ARC_1_1/buf_output[7] )
         );
  XOR2_X1 U7364 ( .A1(\MC_ARK_ARC_1_1/temp4[7] ), .A2(
        \MC_ARK_ARC_1_1/temp3[7] ), .Z(n5184) );
  INV_X2 U7366 ( .I(\SB1_1_27/buf_output[1] ), .ZN(\SB2_1_23/i1_7 ) );
  NAND3_X2 U7368 ( .A1(\SB1_2_12/i0_3 ), .A2(\SB1_2_12/i1[9] ), .A3(
        \SB1_2_12/i0[6] ), .ZN(n5185) );
  NAND4_X2 U7373 ( .A1(n2353), .A2(n1125), .A3(n5186), .A4(
        \SB2_0_21/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_0_21/buf_output[5] ) );
  NAND3_X2 U7374 ( .A1(\SB2_0_21/i0[6] ), .A2(\SB2_0_21/i0[10] ), .A3(
        \SB2_0_21/i0_0 ), .ZN(n5186) );
  XOR2_X1 U7375 ( .A1(n570), .A2(\RI5[2][20] ), .Z(\MC_ARK_ARC_1_2/temp1[20] )
         );
  XOR2_X1 U7383 ( .A1(\MC_ARK_ARC_1_1/temp4[188] ), .A2(n5187), .Z(n5579) );
  XOR2_X1 U7390 ( .A1(\RI5[1][62] ), .A2(\RI5[1][98] ), .Z(n5187) );
  NAND4_X2 U7398 ( .A1(n6385), .A2(\SB2_2_1/Component_Function_0/NAND4_in[1] ), 
        .A3(\SB2_2_1/Component_Function_0/NAND4_in[0] ), .A4(n5188), .ZN(
        \SB2_2_1/buf_output[0] ) );
  NAND3_X2 U7399 ( .A1(\SB1_0_25/i0[10] ), .A2(\SB1_0_25/i0_0 ), .A3(
        \SB1_0_25/i0[6] ), .ZN(\SB1_0_25/Component_Function_5/NAND4_in[1] ) );
  INV_X2 U7414 ( .I(\MC_ARK_ARC_1_1/buf_output[149] ), .ZN(\SB1_2_7/i1_5 ) );
  INV_X4 U7415 ( .I(n5189), .ZN(\SB1_3_4/i1_5 ) );
  INV_X1 U7416 ( .I(\SB1_2_4/buf_output[5] ), .ZN(n5190) );
  NAND4_X2 U7419 ( .A1(\SB1_1_24/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_1_24/Component_Function_5/NAND4_in[0] ), .A3(
        \SB1_1_24/Component_Function_5/NAND4_in[3] ), .A4(n5191), .ZN(
        \SB1_1_24/buf_output[5] ) );
  NAND3_X2 U7427 ( .A1(\SB1_1_24/i0[10] ), .A2(\SB1_1_24/i0_0 ), .A3(
        \SB1_1_24/i0[6] ), .ZN(n5191) );
  NAND4_X2 U7429 ( .A1(\SB2_0_9/Component_Function_2/NAND4_in[0] ), .A2(n4373), 
        .A3(\SB2_0_9/Component_Function_2/NAND4_in[3] ), .A4(n5192), .ZN(
        \SB2_0_9/buf_output[2] ) );
  NAND3_X2 U7432 ( .A1(\SB2_0_9/i0[9] ), .A2(\SB2_0_9/i0_3 ), .A3(
        \SB2_0_9/i0[8] ), .ZN(n5192) );
  XOR2_X1 U7433 ( .A1(\RI5[0][70] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[46] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[100] ) );
  NAND3_X2 U7435 ( .A1(\SB1_1_15/i0_4 ), .A2(\SB1_1_15/i0[9] ), .A3(
        \SB1_1_15/i0[6] ), .ZN(n6070) );
  XOR2_X1 U7438 ( .A1(n5912), .A2(n5911), .Z(n3636) );
  INV_X2 U7439 ( .I(\SB1_2_7/buf_output[1] ), .ZN(\SB2_2_3/i1_7 ) );
  NAND4_X2 U7440 ( .A1(n2202), .A2(\SB1_1_9/Component_Function_5/NAND4_in[1] ), 
        .A3(n3936), .A4(\SB1_1_9/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_9/buf_output[5] ) );
  INV_X2 U7441 ( .I(\SB1_2_6/buf_output[2] ), .ZN(\SB2_2_3/i1[9] ) );
  NAND3_X2 U7443 ( .A1(\SB2_1_9/i0_3 ), .A2(\SB2_1_9/i0_4 ), .A3(
        \SB2_1_9/i0[10] ), .ZN(\SB2_1_9/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U7446 ( .A1(\SB4_1/i0[6] ), .A2(\SB4_1/i0[10] ), .A3(\SB4_1/i0_3 ), 
        .ZN(n5193) );
  NAND3_X2 U7449 ( .A1(\SB4_2/i0[10] ), .A2(\SB4_2/i0_0 ), .A3(\SB4_2/i0[6] ), 
        .ZN(n5194) );
  XOR2_X1 U7450 ( .A1(\SB2_0_24/buf_output[3] ), .A2(\SB2_0_28/buf_output[3] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[87] ) );
  NAND4_X2 U7451 ( .A1(n652), .A2(\SB1_0_11/Component_Function_2/NAND4_in[1] ), 
        .A3(\SB1_0_11/Component_Function_2/NAND4_in[2] ), .A4(n5195), .ZN(
        \SB1_0_11/buf_output[2] ) );
  NAND3_X2 U7454 ( .A1(\SB1_0_11/i0_4 ), .A2(\SB1_0_11/i0_0 ), .A3(
        \SB1_0_11/i1_5 ), .ZN(n5195) );
  XOR2_X1 U7455 ( .A1(\MC_ARK_ARC_1_1/temp4[146] ), .A2(n5197), .Z(
        \MC_ARK_ARC_1_1/temp6[146] ) );
  XOR2_X1 U7456 ( .A1(\RI5[1][20] ), .A2(\RI5[1][56] ), .Z(n5197) );
  NAND3_X2 U7460 ( .A1(\SB2_1_31/i0[10] ), .A2(\SB2_1_31/i0_3 ), .A3(
        \SB2_1_31/i0[6] ), .ZN(\SB2_1_31/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U7462 ( .A1(\SB3_5/i0[8] ), .A2(\SB3_5/i0[9] ), .A3(\SB3_5/i0_0 ), 
        .ZN(\SB3_5/Component_Function_4/NAND4_in[0] ) );
  INV_X2 U7464 ( .I(\MC_ARK_ARC_1_0/buf_output[182] ), .ZN(\SB1_1_1/i1[9] ) );
  NAND3_X2 U7467 ( .A1(\RI1[2][47] ), .A2(\SB1_2_24/i0[8] ), .A3(
        \SB1_2_24/i1_7 ), .ZN(\SB1_2_24/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U7469 ( .A1(n5199), .A2(n5198), .Z(\MC_ARK_ARC_1_2/buf_output[75] )
         );
  XOR2_X1 U7472 ( .A1(\MC_ARK_ARC_1_2/temp2[75] ), .A2(
        \MC_ARK_ARC_1_2/temp4[75] ), .Z(n5198) );
  XOR2_X1 U7479 ( .A1(\MC_ARK_ARC_1_2/temp3[75] ), .A2(n1532), .Z(n5199) );
  XOR2_X1 U7488 ( .A1(n5200), .A2(\MC_ARK_ARC_1_3/temp6[166] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[166] ) );
  XOR2_X1 U7492 ( .A1(n6288), .A2(\MC_ARK_ARC_1_3/temp2[166] ), .Z(n5200) );
  NAND3_X2 U7493 ( .A1(\SB2_2_4/i0[6] ), .A2(\SB2_2_4/i0_3 ), .A3(
        \SB2_2_4/i1[9] ), .ZN(\SB2_2_4/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U7497 ( .A1(\SB4_3/i0_4 ), .A2(\SB4_3/i1_7 ), .A3(n5495), .ZN(
        \SB4_3/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U7499 ( .A1(\SB4_3/Component_Function_0/NAND4_in[1] ), .A2(
        \SB4_3/Component_Function_0/NAND4_in[2] ), .A3(
        \SB4_3/Component_Function_0/NAND4_in[3] ), .A4(n6274), .ZN(n3692) );
  NAND3_X2 U7500 ( .A1(\SB2_0_23/i0[10] ), .A2(\SB2_0_23/i0_3 ), .A3(
        \SB2_0_23/i0[6] ), .ZN(\SB2_0_23/Component_Function_2/NAND4_in[1] ) );
  INV_X2 U7507 ( .I(\SB1_1_11/buf_output[3] ), .ZN(\SB2_1_9/i0[8] ) );
  NAND4_X2 U7508 ( .A1(\SB1_1_11/Component_Function_3/NAND4_in[1] ), .A2(n4667), .A3(n2200), .A4(n3704), .ZN(\SB1_1_11/buf_output[3] ) );
  XOR2_X1 U7509 ( .A1(n5202), .A2(n182), .Z(Ciphertext[58]) );
  NAND4_X2 U7512 ( .A1(\SB4_22/Component_Function_4/NAND4_in[3] ), .A2(n2808), 
        .A3(n4403), .A4(\SB4_22/Component_Function_4/NAND4_in[0] ), .ZN(n5202)
         );
  NAND4_X2 U7514 ( .A1(\SB1_3_15/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_15/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_15/Component_Function_4/NAND4_in[3] ), .A4(n5203), .ZN(
        \SB1_3_15/buf_output[4] ) );
  NAND3_X2 U7522 ( .A1(\SB1_3_15/i0[9] ), .A2(\SB1_3_15/i0[10] ), .A3(
        \SB1_3_15/i0_3 ), .ZN(n5203) );
  NAND3_X2 U7525 ( .A1(\SB2_1_11/i0_3 ), .A2(\SB2_1_11/i1[9] ), .A3(
        \SB2_1_11/i0[6] ), .ZN(\SB2_1_11/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U7526 ( .A1(\SB1_3_4/i0[10] ), .A2(\SB1_3_4/i1_7 ), .A3(
        \SB1_3_4/i1[9] ), .ZN(n1685) );
  NAND3_X2 U7529 ( .A1(\SB2_3_2/i0_3 ), .A2(\SB2_3_2/i0[9] ), .A3(n5491), .ZN(
        n5204) );
  NAND3_X1 U7530 ( .A1(\SB1_3_9/i1_5 ), .A2(\SB1_3_9/i1[9] ), .A3(n5501), .ZN(
        n5346) );
  NAND4_X2 U7531 ( .A1(\SB1_0_2/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_0_2/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_2/Component_Function_1/NAND4_in[3] ), .A4(n5205), .ZN(
        \RI3[0][7] ) );
  NAND2_X1 U7532 ( .A1(\SB1_0_2/i0_3 ), .A2(\SB1_0_2/i1[9] ), .ZN(n5205) );
  INV_X2 U7534 ( .I(\SB1_3_4/buf_output[2] ), .ZN(\SB2_3_1/i1[9] ) );
  NAND4_X2 U7539 ( .A1(n6432), .A2(\SB1_3_4/Component_Function_2/NAND4_in[1] ), 
        .A3(\SB1_3_4/Component_Function_2/NAND4_in[2] ), .A4(n2670), .ZN(
        \SB1_3_4/buf_output[2] ) );
  NAND4_X2 U7541 ( .A1(\SB1_0_20/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_0_20/Component_Function_3/NAND4_in[2] ), .A3(
        \SB1_0_20/Component_Function_3/NAND4_in[0] ), .A4(n5207), .ZN(
        \RI3[0][81] ) );
  NAND3_X1 U7547 ( .A1(\SB2_0_30/i0[6] ), .A2(\SB2_0_30/i1_5 ), .A3(
        \SB1_0_3/buf_output[0] ), .ZN(
        \SB2_0_30/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 U7552 ( .A1(\SB3_5/i1[9] ), .A2(\SB3_5/i1_5 ), .A3(\SB3_5/i0[10] ), 
        .ZN(n5745) );
  NAND4_X2 U7553 ( .A1(\SB2_2_13/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_2_13/Component_Function_4/NAND4_in[1] ), .A3(n4732), .A4(n5209), 
        .ZN(\SB2_2_13/buf_output[4] ) );
  XOR2_X1 U7554 ( .A1(\RI5[2][159] ), .A2(\RI5[2][123] ), .Z(
        \MC_ARK_ARC_1_2/temp3[57] ) );
  NAND4_X2 U7558 ( .A1(\SB2_3_21/Component_Function_3/NAND4_in[3] ), .A2(n4089), .A3(\SB2_3_21/Component_Function_3/NAND4_in[0] ), .A4(n5210), .ZN(
        \SB2_3_21/buf_output[3] ) );
  NAND3_X1 U7564 ( .A1(\SB2_3_21/i0_0 ), .A2(\SB1_3_22/buf_output[4] ), .A3(
        \SB2_3_21/i0_3 ), .ZN(n5210) );
  XOR2_X1 U7565 ( .A1(n5211), .A2(n34), .Z(Ciphertext[156]) );
  NAND4_X2 U7566 ( .A1(\SB4_5/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_5/Component_Function_0/NAND4_in[1] ), .A3(
        \SB4_5/Component_Function_0/NAND4_in[0] ), .A4(n2030), .ZN(n5211) );
  NAND2_X2 U7570 ( .A1(\SB1_3_15/i3[0] ), .A2(\SB1_3_15/i0_0 ), .ZN(n5213) );
  NAND3_X2 U7572 ( .A1(\SB3_5/i1_7 ), .A2(\SB3_5/i1[9] ), .A3(\SB3_5/i0[10] ), 
        .ZN(\SB3_5/Component_Function_3/NAND4_in[2] ) );
  BUF_X4 U7577 ( .I(n428), .Z(\SB1_0_8/i0_3 ) );
  XOR2_X1 U7578 ( .A1(\MC_ARK_ARC_1_2/temp4[15] ), .A2(n5212), .Z(n2831) );
  XOR2_X1 U7586 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[81] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[117] ), .Z(n5212) );
  NAND3_X2 U7587 ( .A1(\SB1_1_2/i0_0 ), .A2(\SB1_1_2/i1_7 ), .A3(
        \SB1_1_2/i3[0] ), .ZN(\SB1_1_2/Component_Function_4/NAND4_in[1] ) );
  NAND4_X2 U7588 ( .A1(\SB1_3_15/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_3_15/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_3_15/Component_Function_5/NAND4_in[1] ), .A4(n5213), .ZN(
        \SB1_3_15/buf_output[5] ) );
  AND2_X1 U7591 ( .A1(\SB1_1_8/Component_Function_4/NAND4_in[0] ), .A2(n5214), 
        .Z(n2891) );
  NAND3_X2 U7592 ( .A1(\SB1_1_8/i0[10] ), .A2(\SB1_1_8/i0[9] ), .A3(
        \RI1[1][143] ), .ZN(n5214) );
  NAND4_X2 U7593 ( .A1(\SB1_1_21/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_1_21/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_1_21/Component_Function_4/NAND4_in[1] ), .A4(n5215), .ZN(
        \SB1_1_21/buf_output[4] ) );
  NAND3_X1 U7595 ( .A1(\SB1_1_21/i0[10] ), .A2(\SB1_1_21/i0_3 ), .A3(n3131), 
        .ZN(n5215) );
  XOR2_X1 U7597 ( .A1(n5216), .A2(n227), .Z(Ciphertext[157]) );
  NAND4_X2 U7599 ( .A1(\SB4_5/Component_Function_1/NAND4_in[2] ), .A2(
        \SB4_5/Component_Function_1/NAND4_in[1] ), .A3(
        \SB4_5/Component_Function_1/NAND4_in[0] ), .A4(n1816), .ZN(n5216) );
  NAND3_X1 U7602 ( .A1(\SB2_1_21/i0_4 ), .A2(\SB2_1_21/i1_7 ), .A3(
        \SB2_1_21/i0[8] ), .ZN(\SB2_1_21/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U7607 ( .A1(n2890), .A2(\SB2_1_20/Component_Function_5/NAND4_in[1] ), .A3(\SB2_1_20/Component_Function_5/NAND4_in[0] ), .A4(n5217), .ZN(
        \SB2_1_20/buf_output[5] ) );
  XOR2_X1 U7608 ( .A1(\MC_ARK_ARC_1_1/temp2[85] ), .A2(n5218), .Z(n6480) );
  XOR2_X1 U7609 ( .A1(\RI5[1][85] ), .A2(\RI5[1][79] ), .Z(n5218) );
  XOR2_X1 U7610 ( .A1(n5219), .A2(n6320), .Z(n706) );
  XOR2_X1 U7611 ( .A1(\RI5[0][134] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[86] ), 
        .Z(n5219) );
  NAND3_X2 U7612 ( .A1(\SB2_1_7/i0[7] ), .A2(\SB2_1_7/i0_0 ), .A3(
        \SB2_1_7/i0_3 ), .ZN(\SB2_1_7/Component_Function_0/NAND4_in[3] ) );
  NAND3_X2 U7615 ( .A1(\SB1_0_17/i0_3 ), .A2(\SB1_0_17/i1_7 ), .A3(
        \SB1_0_17/i0[8] ), .ZN(\SB1_0_17/Component_Function_1/NAND4_in[1] ) );
  NAND3_X2 U7616 ( .A1(\SB2_2_15/i1_5 ), .A2(\SB2_2_15/i0[10] ), .A3(
        \SB2_2_15/i1[9] ), .ZN(\SB2_2_15/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U7619 ( .A1(\SB3_4/i0_0 ), .A2(n2910), .A3(\SB3_4/i0_4 ), .ZN(
        \SB3_4/Component_Function_2/NAND4_in[3] ) );
  NAND4_X2 U7620 ( .A1(\SB2_1_16/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_16/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_16/Component_Function_3/NAND4_in[3] ), .A4(n6403), .ZN(
        \SB2_1_16/buf_output[3] ) );
  XOR2_X1 U7621 ( .A1(n6211), .A2(n5220), .Z(n5366) );
  XOR2_X1 U7623 ( .A1(\RI5[2][188] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[182] ), 
        .Z(n5220) );
  XOR2_X1 U7628 ( .A1(n5221), .A2(\MC_ARK_ARC_1_2/temp4[155] ), .Z(n5460) );
  XOR2_X1 U7633 ( .A1(\RI5[2][155] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[149] ), 
        .Z(n5221) );
  NAND3_X2 U7635 ( .A1(\SB1_3_6/i0_3 ), .A2(\SB1_3_6/i0_4 ), .A3(
        \SB1_3_6/i1[9] ), .ZN(n5222) );
  XOR2_X1 U7638 ( .A1(\MC_ARK_ARC_1_1/temp6[75] ), .A2(n5223), .Z(
        \MC_ARK_ARC_1_1/buf_output[75] ) );
  XOR2_X1 U7645 ( .A1(\MC_ARK_ARC_1_1/temp2[75] ), .A2(
        \MC_ARK_ARC_1_1/temp1[75] ), .Z(n5223) );
  BUF_X4 U7646 ( .I(\SB1_3_9/buf_output[5] ), .Z(\SB2_3_9/i0_3 ) );
  NAND4_X2 U7647 ( .A1(\SB2_2_12/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_2_12/Component_Function_2/NAND4_in[0] ), .A3(n3892), .A4(n5224), 
        .ZN(\SB2_2_12/buf_output[2] ) );
  NAND3_X1 U7649 ( .A1(\SB2_2_12/i0_0 ), .A2(\SB1_2_13/buf_output[4] ), .A3(
        \SB2_2_12/i1_5 ), .ZN(n5224) );
  INV_X8 U7651 ( .I(n2913), .ZN(\RI1[2][47] ) );
  XOR2_X1 U7656 ( .A1(n4314), .A2(n3921), .Z(\MC_ARK_ARC_1_0/buf_output[164] )
         );
  NAND4_X2 U7661 ( .A1(\SB1_3_31/Component_Function_3/NAND4_in[0] ), .A2(n3420), .A3(n6456), .A4(n5225), .ZN(\SB1_3_31/buf_output[3] ) );
  NAND3_X2 U7662 ( .A1(\SB1_3_31/i0[8] ), .A2(\SB1_3_31/i3[0] ), .A3(
        \SB1_3_31/i1_5 ), .ZN(n5225) );
  XOR2_X1 U7663 ( .A1(n5226), .A2(\MC_ARK_ARC_1_2/temp6[81] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[81] ) );
  NAND3_X1 U7666 ( .A1(\SB1_2_25/i0[8] ), .A2(\MC_ARK_ARC_1_1/buf_output[40] ), 
        .A3(\SB1_2_25/i1_7 ), .ZN(n5926) );
  BUF_X4 U7670 ( .I(\SB2_0_24/buf_output[2] ), .Z(\RI5[0][62] ) );
  NAND2_X2 U7671 ( .A1(\SB1_3_9/i3[0] ), .A2(\SB1_3_9/i0_0 ), .ZN(
        \SB1_3_9/Component_Function_5/NAND4_in[0] ) );
  XOR2_X1 U7672 ( .A1(n5227), .A2(n234), .Z(Ciphertext[159]) );
  NAND4_X2 U7674 ( .A1(\SB4_5/Component_Function_3/NAND4_in[3] ), .A2(n3424), 
        .A3(n5260), .A4(n5581), .ZN(n5227) );
  NAND4_X2 U7677 ( .A1(\SB1_1_21/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_1_21/Component_Function_2/NAND4_in[3] ), .A3(n2155), .A4(n5228), 
        .ZN(\SB1_1_21/buf_output[2] ) );
  NAND3_X2 U7679 ( .A1(\SB1_1_21/i0[10] ), .A2(\SB1_1_21/i1[9] ), .A3(
        \SB1_1_21/i1_5 ), .ZN(n5228) );
  NAND3_X2 U7683 ( .A1(\SB2_2_12/i0_4 ), .A2(\SB2_2_12/i0_3 ), .A3(
        \SB2_2_12/i0_0 ), .ZN(\SB2_2_12/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U7686 ( .A1(\RI5[0][10] ), .A2(\RI5[0][16] ), .Z(
        \MC_ARK_ARC_1_0/temp1[16] ) );
  NAND3_X2 U7688 ( .A1(\SB3_5/i0_0 ), .A2(\SB3_5/i0_3 ), .A3(\SB3_5/i0[7] ), 
        .ZN(n5794) );
  XOR2_X1 U7689 ( .A1(\MC_ARK_ARC_1_3/temp4[168] ), .A2(n5229), .Z(
        \MC_ARK_ARC_1_3/temp6[168] ) );
  XOR2_X1 U7691 ( .A1(\RI5[3][42] ), .A2(\RI5[3][78] ), .Z(n5229) );
  NAND2_X2 U7694 ( .A1(n4015), .A2(n4755), .ZN(\SB2_2_8/i0_4 ) );
  NAND4_X2 U7695 ( .A1(\SB2_1_18/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_18/Component_Function_5/NAND4_in[0] ), .A3(n5845), .A4(n5230), 
        .ZN(\SB2_1_18/buf_output[5] ) );
  INV_X4 U7698 ( .I(\SB2_3_29/i0[7] ), .ZN(\RI3[3][16] ) );
  NAND3_X1 U7702 ( .A1(\SB2_3_29/i0[6] ), .A2(\SB2_3_29/i0[8] ), .A3(
        \SB2_3_29/i0[7] ), .ZN(\SB2_3_29/Component_Function_0/NAND4_in[1] ) );
  NOR2_X2 U7703 ( .A1(n5232), .A2(n5231), .ZN(\SB2_3_29/i0[7] ) );
  NAND2_X1 U7704 ( .A1(\SB1_3_30/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_30/Component_Function_4/NAND4_in[1] ), .ZN(n5232) );
  BUF_X4 U7705 ( .I(n3664), .Z(\SB1_3_14/i0_3 ) );
  NAND3_X1 U7711 ( .A1(\SB4_3/i0_3 ), .A2(\SB4_3/i0[7] ), .A3(
        \SB3_6/buf_output[2] ), .ZN(\SB4_3/Component_Function_0/NAND4_in[3] )
         );
  NOR2_X2 U7712 ( .A1(n5789), .A2(n599), .ZN(n3689) );
  NAND3_X2 U7716 ( .A1(\SB2_1_3/i0[7] ), .A2(\SB2_1_3/i0[6] ), .A3(
        \SB2_1_3/i0[8] ), .ZN(n5584) );
  NAND2_X2 U7719 ( .A1(n5234), .A2(n5233), .ZN(
        \SB3_5/Component_Function_3/NAND4_in[3] ) );
  NOR2_X1 U7720 ( .A1(\SB3_5/i0[10] ), .A2(\MC_ARK_ARC_1_3/buf_output[156] ), 
        .ZN(n5233) );
  INV_X2 U7721 ( .I(\SB3_5/i0_3 ), .ZN(n5234) );
  XOR2_X1 U7723 ( .A1(n4160), .A2(\MC_ARK_ARC_1_1/temp2[6] ), .Z(
        \MC_ARK_ARC_1_1/temp5[6] ) );
  INV_X2 U7724 ( .I(\SB1_3_2/buf_output[2] ), .ZN(\SB2_3_31/i1[9] ) );
  NAND4_X2 U7726 ( .A1(\SB1_3_2/Component_Function_2/NAND4_in[2] ), .A2(n5694), 
        .A3(\SB1_3_2/Component_Function_2/NAND4_in[0] ), .A4(
        \SB1_3_2/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB1_3_2/buf_output[2] ) );
  NAND3_X1 U7727 ( .A1(\SB1_3_5/i0_3 ), .A2(\SB1_3_5/i1[9] ), .A3(
        \MC_ARK_ARC_1_2/buf_output[160] ), .ZN(
        \SB1_3_5/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U7733 ( .A1(\SB3_23/Component_Function_0/NAND4_in[3] ), .A2(n946), 
        .A3(\SB3_23/Component_Function_0/NAND4_in[2] ), .A4(n5235), .ZN(
        \SB3_23/buf_output[0] ) );
  NAND2_X1 U7734 ( .A1(\SB3_23/i0[9] ), .A2(\SB3_23/i0[10] ), .ZN(n5235) );
  XOR2_X1 U7736 ( .A1(\SB2_3_4/buf_output[0] ), .A2(\RI5[3][186] ), .Z(
        \MC_ARK_ARC_1_3/temp1[0] ) );
  XOR2_X1 U7737 ( .A1(\RI5[1][3] ), .A2(\RI5[1][39] ), .Z(
        \MC_ARK_ARC_1_1/temp3[129] ) );
  BUF_X4 U7738 ( .I(\MC_ARK_ARC_1_0/buf_output[8] ), .Z(\SB1_1_30/i0_0 ) );
  XOR2_X1 U7745 ( .A1(n5236), .A2(n188), .Z(Ciphertext[3]) );
  NAND4_X2 U7747 ( .A1(n1472), .A2(\SB4_31/Component_Function_3/NAND4_in[3] ), 
        .A3(\SB4_31/Component_Function_3/NAND4_in[2] ), .A4(
        \SB4_31/Component_Function_3/NAND4_in[1] ), .ZN(n5236) );
  XOR2_X1 U7754 ( .A1(n5237), .A2(n2560), .Z(n1601) );
  XOR2_X1 U7755 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[191] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[5] ), .Z(n5237) );
  XOR2_X1 U7756 ( .A1(\MC_ARK_ARC_1_2/temp2[29] ), .A2(n5238), .Z(
        \MC_ARK_ARC_1_2/temp5[29] ) );
  XOR2_X1 U7757 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[29] ), .A2(\RI5[2][23] ), 
        .Z(n5238) );
  XOR2_X1 U7766 ( .A1(\RI5[0][108] ), .A2(\SB2_0_2/buf_output[0] ), .Z(n5239)
         );
  NAND4_X2 U7768 ( .A1(\SB1_1_6/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_1_6/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_1_6/Component_Function_0/NAND4_in[3] ), .A4(
        \SB1_1_6/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_1_6/buf_output[0] ) );
  NAND3_X2 U7770 ( .A1(\SB2_3_21/i0_0 ), .A2(\SB1_3_22/buf_output[4] ), .A3(
        \SB2_3_21/i1_5 ), .ZN(n5552) );
  NAND3_X2 U7772 ( .A1(\SB1_2_17/i0[6] ), .A2(\SB1_2_17/i0[9] ), .A3(
        \SB1_2_17/i0_4 ), .ZN(n4316) );
  XOR2_X1 U7780 ( .A1(\RI5[1][116] ), .A2(\RI5[1][152] ), .Z(n5465) );
  NAND3_X2 U7781 ( .A1(\SB1_0_2/i0_4 ), .A2(\SB1_0_2/i1[9] ), .A3(
        \SB1_0_2/i0_3 ), .ZN(\SB1_0_2/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U7783 ( .A1(n5248), .A2(\SB2_2_21/Component_Function_5/NAND4_in[2] ), .A3(n1811), .A4(\SB2_2_21/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_2_21/buf_output[5] ) );
  XOR2_X1 U7792 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[166] ), .A2(\RI5[0][190] ), 
        .Z(n2073) );
  NAND3_X2 U7797 ( .A1(\SB1_1_29/i0[9] ), .A2(\SB1_1_29/i0_3 ), .A3(
        \SB1_1_29/i0[8] ), .ZN(n1567) );
  CLKBUF_X4 U7799 ( .I(\SB1_3_12/buf_output[0] ), .Z(\SB2_3_7/i0[9] ) );
  NAND2_X2 U7800 ( .A1(\SB1_1_30/i0_0 ), .A2(\SB1_1_30/i3[0] ), .ZN(
        \SB1_1_30/Component_Function_5/NAND4_in[0] ) );
  XOR2_X1 U7805 ( .A1(\MC_ARK_ARC_1_2/temp6[114] ), .A2(
        \MC_ARK_ARC_1_2/temp5[114] ), .Z(\MC_ARK_ARC_1_2/buf_output[114] ) );
  NAND4_X2 U7816 ( .A1(\SB1_2_23/Component_Function_3/NAND4_in[0] ), .A2(n6363), .A3(\SB1_2_23/Component_Function_3/NAND4_in[2] ), .A4(n4712), .ZN(
        \SB1_2_23/buf_output[3] ) );
  XOR2_X1 U7821 ( .A1(\RI5[2][114] ), .A2(\RI5[2][108] ), .Z(
        \MC_ARK_ARC_1_2/temp1[114] ) );
  XOR2_X1 U7825 ( .A1(\RI5[1][151] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[187] ), 
        .Z(n5842) );
  XOR2_X1 U7827 ( .A1(n5313), .A2(n650), .Z(\MC_ARK_ARC_1_3/temp5[160] ) );
  NAND4_X2 U7828 ( .A1(n1538), .A2(n1451), .A3(
        \SB2_1_9/Component_Function_2/NAND4_in[2] ), .A4(n3514), .ZN(
        \SB2_1_9/buf_output[2] ) );
  NAND3_X2 U7835 ( .A1(\SB2_3_23/i0_3 ), .A2(\SB2_3_23/i0[10] ), .A3(
        \SB2_3_23/i0[6] ), .ZN(n6268) );
  BUF_X4 U7836 ( .I(\SB2_3_15/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[116] ) );
  NAND4_X2 U7841 ( .A1(\SB2_3_13/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_3_13/Component_Function_0/NAND4_in[0] ), .A3(
        \SB2_3_13/Component_Function_0/NAND4_in[3] ), .A4(n3162), .ZN(
        \SB2_3_13/buf_output[0] ) );
  NAND2_X1 U7842 ( .A1(n1311), .A2(\SB1_3_16/Component_Function_4/NAND4_in[3] ), .ZN(n6418) );
  XOR2_X1 U7844 ( .A1(n6030), .A2(n5241), .Z(n6003) );
  XOR2_X1 U7845 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[36] ), .A2(\RI5[2][60] ), 
        .Z(n5241) );
  XOR2_X1 U7846 ( .A1(\RI5[0][176] ), .A2(\RI5[0][152] ), .Z(
        \MC_ARK_ARC_1_0/temp2[14] ) );
  XOR2_X1 U7847 ( .A1(n5242), .A2(\MC_ARK_ARC_1_3/temp4[80] ), .Z(n3052) );
  XOR2_X1 U7849 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[182] ), .A2(\RI5[3][146] ), 
        .Z(n5242) );
  NAND3_X2 U7853 ( .A1(\SB1_3_4/i0[8] ), .A2(\SB1_3_4/i3[0] ), .A3(
        \SB1_3_4/i1_5 ), .ZN(n5756) );
  NAND4_X2 U7855 ( .A1(\SB2_2_21/Component_Function_4/NAND4_in[3] ), .A2(n2473), .A3(n792), .A4(n6444), .ZN(\SB2_2_21/buf_output[4] ) );
  NAND4_X2 U7856 ( .A1(n1326), .A2(\SB1_0_2/Component_Function_2/NAND4_in[0] ), 
        .A3(\SB1_0_2/Component_Function_2/NAND4_in[2] ), .A4(n5243), .ZN(
        \RI3[0][2] ) );
  NAND3_X2 U7862 ( .A1(\SB1_0_2/i0[10] ), .A2(\SB1_0_2/i0_3 ), .A3(
        \SB1_0_2/i0[6] ), .ZN(n5243) );
  XOR2_X1 U7863 ( .A1(\SB2_3_13/buf_output[1] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[109] ), .Z(\MC_ARK_ARC_1_3/temp2[163] )
         );
  NAND3_X1 U7866 ( .A1(\SB1_1_26/i0_0 ), .A2(\SB1_1_26/i3[0] ), .A3(
        \SB1_1_26/i1_7 ), .ZN(\SB1_1_26/Component_Function_4/NAND4_in[1] ) );
  NAND3_X2 U7867 ( .A1(\SB2_3_11/i0[10] ), .A2(n4768), .A3(\SB2_3_11/i1[9] ), 
        .ZN(\SB2_3_11/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U7868 ( .A1(\SB3_23/i0_3 ), .A2(\SB3_23/i0[6] ), .A3(
        \SB3_23/i0[10] ), .ZN(\SB3_23/Component_Function_2/NAND4_in[1] ) );
  NAND4_X2 U7869 ( .A1(\SB1_3_25/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_25/Component_Function_2/NAND4_in[2] ), .A3(n1814), .A4(n5244), 
        .ZN(\SB1_3_25/buf_output[2] ) );
  BUF_X4 U7873 ( .I(\SB2_3_22/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[74] ) );
  NAND4_X2 U7875 ( .A1(\SB2_2_10/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_2_10/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_10/Component_Function_1/NAND4_in[0] ), .A4(n5245), .ZN(
        \SB2_2_10/buf_output[1] ) );
  XOR2_X1 U7878 ( .A1(\RI5[2][10] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[34] ), 
        .Z(n5591) );
  XOR2_X1 U7879 ( .A1(n5246), .A2(\MC_ARK_ARC_1_0/temp4[26] ), .Z(
        \MC_ARK_ARC_1_0/temp6[26] ) );
  XOR2_X1 U7881 ( .A1(\SB2_0_13/buf_output[2] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[92] ), .Z(n5246) );
  XOR2_X1 U7885 ( .A1(n626), .A2(n5247), .Z(\RI1[4][89] ) );
  XOR2_X1 U7886 ( .A1(n5905), .A2(\MC_ARK_ARC_1_3/temp1[89] ), .Z(n5247) );
  NAND3_X2 U7889 ( .A1(\SB2_2_21/i0_0 ), .A2(\SB2_2_21/i0[6] ), .A3(
        \SB2_2_21/i0[10] ), .ZN(n5248) );
  XOR2_X1 U7890 ( .A1(n5249), .A2(n242), .Z(Ciphertext[76]) );
  NAND4_X2 U7891 ( .A1(\SB4_19/Component_Function_4/NAND4_in[0] ), .A2(
        \SB4_19/Component_Function_4/NAND4_in[2] ), .A3(
        \SB4_19/Component_Function_4/NAND4_in[3] ), .A4(
        \SB4_19/Component_Function_4/NAND4_in[1] ), .ZN(n5249) );
  XOR2_X1 U7893 ( .A1(n5250), .A2(n213), .Z(Ciphertext[74]) );
  NAND4_X2 U7894 ( .A1(\SB4_19/Component_Function_2/NAND4_in[2] ), .A2(
        \SB4_19/Component_Function_2/NAND4_in[1] ), .A3(n2049), .A4(
        \SB4_19/Component_Function_2/NAND4_in[0] ), .ZN(n5250) );
  XOR2_X1 U7897 ( .A1(\MC_ARK_ARC_1_0/temp1[110] ), .A2(n5251), .Z(n1654) );
  XOR2_X1 U7898 ( .A1(\RI5[0][176] ), .A2(\RI5[0][20] ), .Z(n5251) );
  XOR2_X1 U7902 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[2] ), .A2(\RI5[0][188] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[2] ) );
  NAND3_X2 U7910 ( .A1(\SB1_3_21/i0_4 ), .A2(\SB1_3_21/i0_3 ), .A3(
        \SB1_3_21/i1[9] ), .ZN(n5252) );
  XOR2_X1 U7911 ( .A1(n5253), .A2(\MC_ARK_ARC_1_1/temp6[162] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[162] ) );
  XOR2_X1 U7912 ( .A1(n5635), .A2(n6423), .Z(n5253) );
  NAND4_X2 U7921 ( .A1(\SB2_1_0/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_1_0/Component_Function_1/NAND4_in[1] ), .A3(n4387), .A4(
        \SB2_1_0/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_1_0/buf_output[1] ) );
  NAND4_X2 U7923 ( .A1(\SB3_17/Component_Function_2/NAND4_in[3] ), .A2(
        \SB3_17/Component_Function_2/NAND4_in[0] ), .A3(n5599), .A4(
        \SB3_17/Component_Function_2/NAND4_in[2] ), .ZN(\SB3_17/buf_output[2] ) );
  NAND4_X2 U7929 ( .A1(\SB1_1_31/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_1_31/Component_Function_0/NAND4_in[0] ), .A3(
        \SB1_1_31/Component_Function_0/NAND4_in[2] ), .A4(n5254), .ZN(
        \SB1_1_31/buf_output[0] ) );
  NAND3_X2 U7931 ( .A1(\SB1_1_31/i0_0 ), .A2(\SB1_1_31/i0[7] ), .A3(
        \SB1_1_31/i0_3 ), .ZN(n5254) );
  NAND3_X2 U7934 ( .A1(\SB2_2_5/i0[10] ), .A2(\SB2_2_5/i1_5 ), .A3(
        \SB2_2_5/i1[9] ), .ZN(\SB2_2_5/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U7935 ( .A1(\SB2_2_3/Component_Function_1/NAND4_in[0] ), .A2(n5728), 
        .A3(\SB2_2_3/Component_Function_1/NAND4_in[3] ), .A4(n5256), .ZN(
        \SB2_2_3/buf_output[1] ) );
  XOR2_X1 U7937 ( .A1(\MC_ARK_ARC_1_2/temp6[101] ), .A2(n5257), .Z(
        \MC_ARK_ARC_1_2/buf_output[101] ) );
  XOR2_X1 U7939 ( .A1(n5726), .A2(\MC_ARK_ARC_1_2/temp1[101] ), .Z(n5257) );
  XOR2_X1 U7940 ( .A1(n5259), .A2(n5258), .Z(n1478) );
  XOR2_X1 U7941 ( .A1(\RI5[3][37] ), .A2(n216), .Z(n5258) );
  XOR2_X1 U7967 ( .A1(\RI5[3][7] ), .A2(\RI5[3][73] ), .Z(n5259) );
  NAND3_X1 U7969 ( .A1(\SB4_5/i0_3 ), .A2(\SB4_5/i0[6] ), .A3(\SB4_5/i1[9] ), 
        .ZN(n5260) );
  BUF_X4 U7970 ( .I(\SB2_3_18/buf_output[3] ), .Z(\RI5[3][93] ) );
  NAND3_X2 U7972 ( .A1(\SB2_2_8/i0_3 ), .A2(\SB2_2_8/i0[6] ), .A3(
        \SB2_2_8/i0[10] ), .ZN(n1249) );
  NAND4_X2 U7973 ( .A1(\SB1_2_22/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_2_22/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_2_22/Component_Function_2/NAND4_in[2] ), .A4(n5261), .ZN(
        \SB1_2_22/buf_output[2] ) );
  NAND3_X1 U7974 ( .A1(\SB1_2_22/i0_0 ), .A2(\SB1_2_22/i1_5 ), .A3(
        \SB1_2_22/i0_4 ), .ZN(n5261) );
  NAND4_X2 U7975 ( .A1(\SB2_3_23/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_3_23/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_3_23/Component_Function_1/NAND4_in[0] ), .A4(n5262), .ZN(
        \SB2_3_23/buf_output[1] ) );
  NAND3_X1 U7979 ( .A1(\SB2_3_23/i0[9] ), .A2(\SB2_3_23/i0[6] ), .A3(
        \SB2_3_23/i1_5 ), .ZN(n5262) );
  NAND4_X2 U7984 ( .A1(\SB1_2_3/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_3/Component_Function_4/NAND4_in[3] ), .A3(
        \SB1_2_3/Component_Function_4/NAND4_in[2] ), .A4(n5263), .ZN(
        \SB1_2_3/buf_output[4] ) );
  NAND3_X2 U7994 ( .A1(\SB2_3_29/i0[10] ), .A2(\SB2_3_29/i1_5 ), .A3(
        \SB2_3_29/i1[9] ), .ZN(\SB2_3_29/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U8003 ( .A1(\MC_ARK_ARC_1_2/temp4[69] ), .A2(
        \MC_ARK_ARC_1_2/temp3[69] ), .Z(n5264) );
  XOR2_X1 U8007 ( .A1(n5265), .A2(n134), .Z(Ciphertext[96]) );
  NAND4_X2 U8012 ( .A1(\SB4_15/Component_Function_0/NAND4_in[3] ), .A2(
        \SB4_15/Component_Function_0/NAND4_in[1] ), .A3(
        \SB4_15/Component_Function_0/NAND4_in[2] ), .A4(n3854), .ZN(n5265) );
  NAND3_X1 U8013 ( .A1(\SB3_2/i0[6] ), .A2(\SB3_2/i0[8] ), .A3(\SB3_2/i0[7] ), 
        .ZN(\SB3_2/Component_Function_0/NAND4_in[1] ) );
  NAND4_X2 U8014 ( .A1(\SB2_0_0/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_0/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_0_0/Component_Function_5/NAND4_in[0] ), .A4(n5267), .ZN(
        \SB2_0_0/buf_output[5] ) );
  NAND3_X2 U8018 ( .A1(\SB2_0_0/i0[10] ), .A2(\SB2_0_0/i0_0 ), .A3(
        \SB2_0_0/i0[6] ), .ZN(n5267) );
  NAND4_X2 U8019 ( .A1(\SB2_2_2/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_2_2/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_2_2/Component_Function_4/NAND4_in[2] ), .A4(n5268), .ZN(
        \SB2_2_2/buf_output[4] ) );
  NAND3_X2 U8020 ( .A1(\SB2_2_2/i0_4 ), .A2(\SB2_2_2/i1[9] ), .A3(
        \SB2_2_2/i1_5 ), .ZN(n5268) );
  XOR2_X1 U8022 ( .A1(n5269), .A2(n205), .Z(Ciphertext[31]) );
  NAND4_X2 U8024 ( .A1(\SB4_26/Component_Function_1/NAND4_in[2] ), .A2(
        \SB4_26/Component_Function_1/NAND4_in[3] ), .A3(
        \SB4_26/Component_Function_1/NAND4_in[0] ), .A4(
        \SB4_26/Component_Function_1/NAND4_in[1] ), .ZN(n5269) );
  NAND3_X1 U8026 ( .A1(\SB1_3_4/i0[6] ), .A2(\SB1_3_4/i0[8] ), .A3(
        \SB1_3_4/i0[7] ), .ZN(\SB1_3_4/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U8029 ( .A1(n5270), .A2(n59), .Z(Ciphertext[184]) );
  NAND4_X2 U8031 ( .A1(\SB4_1/Component_Function_4/NAND4_in[3] ), .A2(n5640), 
        .A3(n3469), .A4(n6377), .ZN(n5270) );
  XOR2_X1 U8039 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[74] ), .A2(\RI5[1][50] ), 
        .Z(n3102) );
  INV_X2 U8045 ( .I(\SB1_2_23/buf_output[3] ), .ZN(\SB2_2_21/i0[8] ) );
  XOR2_X1 U8046 ( .A1(n1665), .A2(n5271), .Z(\MC_ARK_ARC_1_2/buf_output[23] )
         );
  XOR2_X1 U8048 ( .A1(n3961), .A2(n882), .Z(n5271) );
  NAND4_X2 U8049 ( .A1(n2469), .A2(\SB4_2/Component_Function_2/NAND4_in[2] ), 
        .A3(\SB4_2/Component_Function_2/NAND4_in[3] ), .A4(n5272), .ZN(n6471)
         );
  XOR2_X1 U8051 ( .A1(n5273), .A2(\MC_ARK_ARC_1_2/temp4[131] ), .Z(
        \MC_ARK_ARC_1_2/temp6[131] ) );
  XOR2_X1 U8052 ( .A1(\RI5[2][5] ), .A2(\RI5[2][41] ), .Z(n5273) );
  NAND4_X2 U8054 ( .A1(\SB2_2_31/Component_Function_5/NAND4_in[1] ), .A2(
        \SB2_2_31/Component_Function_5/NAND4_in[3] ), .A3(
        \SB2_2_31/Component_Function_5/NAND4_in[0] ), .A4(n5274), .ZN(
        \SB2_2_31/buf_output[5] ) );
  NAND3_X2 U8055 ( .A1(\SB2_2_31/i0_3 ), .A2(n569), .A3(\SB2_2_31/i1[9] ), 
        .ZN(n5274) );
  NAND3_X1 U8056 ( .A1(\SB4_31/i0[9] ), .A2(\SB4_31/i0_4 ), .A3(\SB4_31/i0[6] ), .ZN(n1238) );
  NAND3_X2 U8063 ( .A1(\SB1_0_20/i0_3 ), .A2(\SB1_0_20/i0_4 ), .A3(
        \SB1_0_20/i1[9] ), .ZN(n804) );
  NAND4_X2 U8064 ( .A1(\SB2_2_20/Component_Function_5/NAND4_in[1] ), .A2(n1644), .A3(n669), .A4(\SB2_2_20/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_2_20/buf_output[5] ) );
  NAND3_X2 U8066 ( .A1(\SB1_1_30/i0_3 ), .A2(\SB1_1_30/i1[9] ), .A3(
        \SB1_1_30/i0[6] ), .ZN(\SB1_1_30/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U8069 ( .A1(\SB1_2_8/i0[10] ), .A2(\SB1_2_8/i1[9] ), .A3(
        \SB1_2_8/i1_5 ), .ZN(n5281) );
  NAND3_X2 U8070 ( .A1(\SB1_1_12/i0_4 ), .A2(\SB1_1_12/i0_3 ), .A3(
        \SB1_1_12/i1[9] ), .ZN(n6328) );
  BUF_X4 U8083 ( .I(\MC_ARK_ARC_1_3/buf_output[160] ), .Z(\SB3_5/i0_4 ) );
  XOR2_X1 U8088 ( .A1(\RI5[2][171] ), .A2(\SB2_2_9/buf_output[3] ), .Z(n5973)
         );
  NAND4_X2 U8089 ( .A1(n1620), .A2(\SB2_2_9/Component_Function_0/NAND4_in[2] ), 
        .A3(\SB2_2_9/Component_Function_0/NAND4_in[3] ), .A4(
        \SB2_2_9/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_2_9/buf_output[0] ) );
  NAND3_X1 U8090 ( .A1(\SB2_3_15/i0_3 ), .A2(\SB2_3_15/i0[9] ), .A3(
        \SB1_3_17/buf_output[3] ), .ZN(n643) );
  NAND3_X2 U8111 ( .A1(\SB2_2_5/i0[10] ), .A2(\SB2_2_5/i1_7 ), .A3(
        \SB2_2_5/i1[9] ), .ZN(\SB2_2_5/Component_Function_3/NAND4_in[2] ) );
  INV_X2 U8116 ( .I(\MC_ARK_ARC_1_1/buf_output[122] ), .ZN(\SB1_2_11/i1[9] )
         );
  NAND4_X2 U8118 ( .A1(\SB1_3_27/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_3_27/Component_Function_5/NAND4_in[1] ), .A3(n4459), .A4(n5275), 
        .ZN(\SB1_3_27/buf_output[5] ) );
  NAND3_X2 U8123 ( .A1(\SB1_3_27/i0[9] ), .A2(\SB1_3_27/i0[6] ), .A3(
        \SB1_3_27/i0_4 ), .ZN(n5275) );
  NAND3_X1 U8127 ( .A1(\SB1_2_15/i0_3 ), .A2(\SB1_2_15/i0[8] ), .A3(
        \SB1_2_15/i1_7 ), .ZN(\SB1_2_15/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U8128 ( .A1(n4298), .A2(n5276), .Z(\MC_ARK_ARC_1_2/buf_output[35] )
         );
  XOR2_X1 U8129 ( .A1(\RI5[3][39] ), .A2(\RI5[3][75] ), .Z(
        \MC_ARK_ARC_1_3/temp3[165] ) );
  XOR2_X1 U8131 ( .A1(\MC_ARK_ARC_1_3/temp4[22] ), .A2(
        \MC_ARK_ARC_1_3/temp3[22] ), .Z(\MC_ARK_ARC_1_3/temp6[22] ) );
  XOR2_X1 U8133 ( .A1(\MC_ARK_ARC_1_2/temp4[96] ), .A2(
        \MC_ARK_ARC_1_2/temp3[96] ), .Z(\MC_ARK_ARC_1_2/temp6[96] ) );
  NAND4_X2 U8138 ( .A1(\SB1_3_12/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_12/Component_Function_2/NAND4_in[2] ), .A3(
        \SB1_3_12/Component_Function_2/NAND4_in[0] ), .A4(n5277), .ZN(
        \SB1_3_12/buf_output[2] ) );
  NAND3_X2 U8140 ( .A1(\SB1_3_12/i0_4 ), .A2(\SB1_3_12/i1_5 ), .A3(
        \SB1_3_12/i0_0 ), .ZN(n5277) );
  XOR2_X1 U8144 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[67] ), .A2(\RI5[0][31] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[157] ) );
  BUF_X4 U8149 ( .I(\SB1_1_5/buf_output[1] ), .Z(\SB2_1_1/i0[6] ) );
  NAND4_X2 U8151 ( .A1(\SB2_0_30/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_30/Component_Function_5/NAND4_in[0] ), .A3(n5279), .A4(n5278), 
        .ZN(\SB2_0_30/buf_output[5] ) );
  NAND3_X2 U8152 ( .A1(\SB2_0_30/i0[10] ), .A2(\SB2_0_30/i0_0 ), .A3(
        \SB2_0_30/i0[6] ), .ZN(n5278) );
  NAND3_X2 U8153 ( .A1(\SB2_1_27/i0[10] ), .A2(\SB2_1_27/i1_7 ), .A3(
        \SB2_1_27/i1[9] ), .ZN(n5280) );
  NAND4_X2 U8156 ( .A1(\SB2_0_19/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_19/Component_Function_3/NAND4_in[2] ), .A3(n1239), .A4(n5282), 
        .ZN(\SB2_0_19/buf_output[3] ) );
  NAND3_X2 U8166 ( .A1(\SB2_0_19/i0_3 ), .A2(\SB2_0_19/i0_0 ), .A3(
        \RI3[0][76] ), .ZN(n5282) );
  XOR2_X1 U8169 ( .A1(n926), .A2(n5283), .Z(\MC_ARK_ARC_1_1/temp5[143] ) );
  XOR2_X1 U8175 ( .A1(\RI5[1][137] ), .A2(\RI5[1][143] ), .Z(n5283) );
  NAND3_X2 U8177 ( .A1(\SB2_2_5/i0_3 ), .A2(\SB2_2_5/i0_4 ), .A3(
        \SB2_2_5/i1[9] ), .ZN(n4003) );
  XOR2_X1 U8178 ( .A1(\MC_ARK_ARC_1_1/temp3[157] ), .A2(n5284), .Z(n1642) );
  XOR2_X1 U8179 ( .A1(\RI5[1][157] ), .A2(\RI5[1][151] ), .Z(n5284) );
  NAND3_X2 U8181 ( .A1(\SB1_1_30/i0_0 ), .A2(\SB1_1_30/i0[8] ), .A3(
        \SB1_1_30/i0[9] ), .ZN(n2725) );
  NAND2_X2 U8182 ( .A1(\SB2_2_11/i0_3 ), .A2(n4754), .ZN(n5285) );
  XOR2_X1 U8183 ( .A1(\MC_ARK_ARC_1_0/temp4[111] ), .A2(n5286), .Z(n1964) );
  XOR2_X1 U8184 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[21] ), .A2(\RI5[0][177] ), 
        .Z(n5286) );
  XOR2_X1 U8190 ( .A1(n5289), .A2(n5288), .Z(\MC_ARK_ARC_1_1/buf_output[122] )
         );
  XOR2_X1 U8193 ( .A1(n3149), .A2(n4345), .Z(n5288) );
  XOR2_X1 U8195 ( .A1(n2502), .A2(n4111), .Z(n5289) );
  XOR2_X1 U8197 ( .A1(\MC_ARK_ARC_1_0/temp4[163] ), .A2(n5290), .Z(
        \MC_ARK_ARC_1_0/temp6[163] ) );
  XOR2_X1 U8201 ( .A1(\RI5[0][37] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[73] ), 
        .Z(n5290) );
  NAND3_X2 U8202 ( .A1(\SB3_31/i1_5 ), .A2(\SB3_31/i0[8] ), .A3(\SB3_31/i3[0] ), .ZN(\SB3_31/Component_Function_3/NAND4_in[3] ) );
  NAND4_X2 U8203 ( .A1(\SB2_3_11/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_11/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_3_11/Component_Function_4/NAND4_in[1] ), .A4(n5291), .ZN(
        \SB2_3_11/buf_output[4] ) );
  NAND3_X2 U8205 ( .A1(\SB2_1_23/i0_3 ), .A2(\SB2_1_23/i0[9] ), .A3(
        \SB2_1_23/i0[8] ), .ZN(\SB2_1_23/Component_Function_2/NAND4_in[2] ) );
  XOR2_X1 U8207 ( .A1(n5292), .A2(n90), .Z(Ciphertext[120]) );
  NAND4_X2 U8208 ( .A1(\SB4_11/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_11/Component_Function_0/NAND4_in[3] ), .A3(
        \SB4_11/Component_Function_0/NAND4_in[1] ), .A4(n4216), .ZN(n5292) );
  NAND4_X2 U8214 ( .A1(n3957), .A2(\SB1_3_8/Component_Function_1/NAND4_in[1] ), 
        .A3(\SB1_3_8/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_3_8/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_3_8/buf_output[1] ) );
  BUF_X4 U8215 ( .I(\SB1_3_4/buf_output[3] ), .Z(\SB2_3_2/i0[10] ) );
  NAND3_X2 U8218 ( .A1(\SB3_2/i0_3 ), .A2(\SB3_2/i0_4 ), .A3(\SB3_2/i1[9] ), 
        .ZN(n5572) );
  XOR2_X1 U8219 ( .A1(\MC_ARK_ARC_1_1/temp1[114] ), .A2(
        \MC_ARK_ARC_1_1/temp2[114] ), .Z(n613) );
  NAND3_X1 U8220 ( .A1(\SB2_3_4/i0[6] ), .A2(\SB2_3_4/i0[8] ), .A3(
        \SB2_3_4/i0[7] ), .ZN(\SB2_3_4/Component_Function_0/NAND4_in[1] ) );
  NAND3_X2 U8224 ( .A1(\SB2_3_7/i0_3 ), .A2(\SB1_3_8/buf_output[4] ), .A3(
        \SB2_3_7/i0_0 ), .ZN(n6106) );
  NAND4_X2 U8225 ( .A1(\SB1_1_18/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_18/Component_Function_2/NAND4_in[2] ), .A3(
        \SB1_1_18/Component_Function_2/NAND4_in[1] ), .A4(n5293), .ZN(
        \SB1_1_18/buf_output[2] ) );
  NAND3_X2 U8227 ( .A1(\SB1_1_18/i0_4 ), .A2(\SB1_1_18/i0_0 ), .A3(
        \SB1_1_18/i1_5 ), .ZN(n5293) );
  XOR2_X1 U8228 ( .A1(n4357), .A2(n5294), .Z(\MC_ARK_ARC_1_1/buf_output[117] )
         );
  XOR2_X1 U8230 ( .A1(n1560), .A2(\MC_ARK_ARC_1_1/temp2[117] ), .Z(n5294) );
  XOR2_X1 U8231 ( .A1(n3694), .A2(\MC_ARK_ARC_1_3/temp4[187] ), .Z(
        \MC_ARK_ARC_1_3/temp6[187] ) );
  NAND3_X2 U8232 ( .A1(\SB2_3_25/i0[9] ), .A2(\SB2_3_25/i1_5 ), .A3(
        \SB2_3_25/i0[6] ), .ZN(\SB2_3_25/Component_Function_1/NAND4_in[2] ) );
  BUF_X4 U8238 ( .I(n422), .Z(\SB1_0_14/i0_3 ) );
  XOR2_X1 U8244 ( .A1(n5296), .A2(n5295), .Z(\MC_ARK_ARC_1_1/temp5[2] ) );
  XOR2_X1 U8248 ( .A1(\RI5[1][2] ), .A2(\RI5[1][140] ), .Z(n5295) );
  XOR2_X1 U8252 ( .A1(\RI5[1][188] ), .A2(\RI5[1][164] ), .Z(n5296) );
  NAND4_X2 U8255 ( .A1(\SB2_0_2/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_0_2/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_0_2/Component_Function_0/NAND4_in[0] ), .A4(n5297), .ZN(
        \SB2_0_2/buf_output[0] ) );
  NAND3_X2 U8256 ( .A1(\SB2_2_25/i0[10] ), .A2(\SB2_2_25/i0[6] ), .A3(
        \SB2_2_25/i0_0 ), .ZN(n5298) );
  NAND4_X2 U8271 ( .A1(\SB2_2_10/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_10/Component_Function_5/NAND4_in[1] ), .A3(n5300), .A4(
        \SB2_2_10/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_2_10/buf_output[5] ) );
  NAND3_X2 U8276 ( .A1(\SB2_2_10/i0[6] ), .A2(n581), .A3(\SB2_2_10/i0[9] ), 
        .ZN(n5300) );
  NAND3_X1 U8280 ( .A1(\SB4_0/i0[9] ), .A2(\SB4_0/i0_3 ), .A3(\SB4_0/i0[8] ), 
        .ZN(n5301) );
  NAND3_X2 U8293 ( .A1(\SB1_3_17/i0[10] ), .A2(\SB1_3_17/i0_3 ), .A3(
        \SB1_3_17/i0[6] ), .ZN(n5937) );
  XOR2_X1 U8294 ( .A1(\MC_ARK_ARC_1_3/temp5[164] ), .A2(n5302), .Z(
        \MC_ARK_ARC_1_3/buf_output[164] ) );
  XOR2_X1 U8295 ( .A1(\MC_ARK_ARC_1_3/temp4[164] ), .A2(n3037), .Z(n5302) );
  NAND3_X2 U8296 ( .A1(\SB2_1_25/i3[0] ), .A2(\SB2_1_25/i0[8] ), .A3(
        \SB2_1_25/i1_5 ), .ZN(\SB2_1_25/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U8298 ( .A1(n5303), .A2(n45), .Z(Ciphertext[59]) );
  NAND4_X2 U8300 ( .A1(\SB4_22/Component_Function_5/NAND4_in[1] ), .A2(
        \SB4_22/Component_Function_5/NAND4_in[2] ), .A3(
        \SB4_22/Component_Function_5/NAND4_in[0] ), .A4(n5471), .ZN(n5303) );
  INV_X2 U8304 ( .I(\MC_ARK_ARC_1_3/buf_output[38] ), .ZN(\SB3_25/i1[9] ) );
  NAND3_X1 U8307 ( .A1(\SB1_1_30/i0_3 ), .A2(\SB1_1_30/i0[10] ), .A3(
        \SB1_1_30/i0_4 ), .ZN(\SB1_1_30/Component_Function_0/NAND4_in[2] ) );
  BUF_X4 U8308 ( .I(\SB2_2_10/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[141] ) );
  INV_X1 U8309 ( .I(\SB3_24/buf_output[1] ), .ZN(\SB4_20/i1_7 ) );
  NAND4_X2 U8312 ( .A1(n4173), .A2(\SB3_24/Component_Function_1/NAND4_in[1] ), 
        .A3(\SB3_24/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_24/Component_Function_1/NAND4_in[0] ), .ZN(\SB3_24/buf_output[1] ) );
  XOR2_X1 U8313 ( .A1(n5305), .A2(n160), .Z(Ciphertext[22]) );
  NAND4_X2 U8315 ( .A1(n2671), .A2(n4482), .A3(n5589), .A4(n6044), .ZN(n5305)
         );
  NAND3_X2 U8316 ( .A1(n2605), .A2(\SB2_0_29/i0_4 ), .A3(\SB2_0_29/i0[6] ), 
        .ZN(n3439) );
  NAND3_X2 U8319 ( .A1(\SB1_3_26/i0_3 ), .A2(\SB1_3_26/i1_7 ), .A3(
        \SB1_3_26/i0[8] ), .ZN(\SB1_3_26/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U8323 ( .A1(n5306), .A2(n3009), .Z(\MC_ARK_ARC_1_3/buf_output[174] )
         );
  XOR2_X1 U8326 ( .A1(\MC_ARK_ARC_1_3/temp3[174] ), .A2(
        \MC_ARK_ARC_1_3/temp4[174] ), .Z(n5306) );
  BUF_X4 U8329 ( .I(\MC_ARK_ARC_1_2/buf_output[129] ), .Z(\SB1_3_10/i0[10] )
         );
  NAND4_X2 U8333 ( .A1(\SB1_0_17/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_0_17/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_17/Component_Function_1/NAND4_in[3] ), .A4(n5904), .ZN(
        \SB1_0_17/buf_output[1] ) );
  NAND3_X2 U8334 ( .A1(\SB1_2_20/i0[10] ), .A2(\SB1_2_20/i1[9] ), .A3(n2909), 
        .ZN(n5699) );
  NAND3_X2 U8337 ( .A1(\SB2_3_4/i0[6] ), .A2(\SB2_3_4/i0_3 ), .A3(
        \SB2_3_4/i1[9] ), .ZN(n2128) );
  XOR2_X1 U8341 ( .A1(\RI5[0][143] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[179] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[77] ) );
  XOR2_X1 U8342 ( .A1(n5308), .A2(n153), .Z(Ciphertext[8]) );
  NAND4_X2 U8344 ( .A1(\SB4_30/Component_Function_2/NAND4_in[2] ), .A2(
        \SB4_30/Component_Function_2/NAND4_in[0] ), .A3(n5312), .A4(n5424), 
        .ZN(n5308) );
  XOR2_X1 U8345 ( .A1(n5309), .A2(n51), .Z(Ciphertext[56]) );
  NAND4_X2 U8346 ( .A1(n4242), .A2(\SB4_22/Component_Function_2/NAND4_in[1] ), 
        .A3(\SB4_22/Component_Function_2/NAND4_in[3] ), .A4(n6260), .ZN(n5309)
         );
  XOR2_X1 U8347 ( .A1(n5310), .A2(n17), .Z(Ciphertext[6]) );
  NAND4_X2 U8349 ( .A1(n5433), .A2(\SB4_30/Component_Function_0/NAND4_in[2] ), 
        .A3(n4384), .A4(\SB4_30/Component_Function_0/NAND4_in[1] ), .ZN(n5310)
         );
  NAND3_X2 U8350 ( .A1(\SB2_2_1/i0_3 ), .A2(\SB2_2_1/i0_4 ), .A3(
        \SB2_2_1/i1[9] ), .ZN(\SB2_2_1/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U8352 ( .A1(\SB2_3_9/i0_4 ), .A2(\SB2_3_9/i0[6] ), .A3(
        \SB2_3_9/i0[9] ), .ZN(n1403) );
  NAND3_X1 U8353 ( .A1(\SB4_31/i0_0 ), .A2(\SB4_31/i0[7] ), .A3(\SB4_31/i0_3 ), 
        .ZN(\SB4_31/Component_Function_0/NAND4_in[3] ) );
  NAND4_X2 U8354 ( .A1(\SB1_0_22/Component_Function_5/NAND4_in[2] ), .A2(n5415), .A3(\SB1_0_22/Component_Function_5/NAND4_in[0] ), .A4(n2773), .ZN(
        \SB1_0_22/buf_output[5] ) );
  NAND3_X1 U8355 ( .A1(\SB2_3_19/i0[6] ), .A2(\SB2_3_19/i0_3 ), .A3(n5494), 
        .ZN(\SB2_3_19/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U8356 ( .A1(\SB4_1/i1[9] ), .A2(\SB4_1/i0[10] ), .A3(\SB4_1/i1_5 ), 
        .ZN(n3809) );
  NAND4_X2 U8359 ( .A1(\SB1_1_19/Component_Function_2/NAND4_in[3] ), .A2(
        \SB1_1_19/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_1_19/Component_Function_2/NAND4_in[0] ), .A4(n4101), .ZN(
        \SB1_1_19/buf_output[2] ) );
  BUF_X4 U8361 ( .I(\SB2_3_7/buf_output[3] ), .Z(\RI5[3][159] ) );
  XOR2_X1 U8362 ( .A1(n5311), .A2(n4416), .Z(\MC_ARK_ARC_1_2/temp5[131] ) );
  XOR2_X1 U8363 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[125] ), .A2(\RI5[2][101] ), 
        .Z(n5311) );
  XOR2_X1 U8364 ( .A1(\MC_ARK_ARC_1_1/temp5[159] ), .A2(n6470), .Z(
        \MC_ARK_ARC_1_1/buf_output[159] ) );
  NAND4_X2 U8366 ( .A1(\SB2_0_31/Component_Function_5/NAND4_in[1] ), .A2(n5386), .A3(n2920), .A4(\SB2_0_31/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_0_31/buf_output[5] ) );
  NAND4_X2 U8367 ( .A1(\SB2_3_22/Component_Function_2/NAND4_in[0] ), .A2(n4671), .A3(n5423), .A4(\SB2_3_22/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB2_3_22/buf_output[2] ) );
  NAND4_X2 U8369 ( .A1(\SB1_3_25/Component_Function_5/NAND4_in[1] ), .A2(n1761), .A3(n5683), .A4(n5684), .ZN(\SB1_3_25/buf_output[5] ) );
  NAND3_X2 U8370 ( .A1(\SB1_0_17/i0_0 ), .A2(n2899), .A3(\SB1_0_17/i1_5 ), 
        .ZN(n4193) );
  NAND3_X2 U8373 ( .A1(\SB2_2_31/i0_0 ), .A2(\SB2_2_31/i0_3 ), .A3(n569), .ZN(
        \SB2_2_31/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U8374 ( .A1(\SB1_3_28/i0_3 ), .A2(\SB1_3_28/i0_4 ), .A3(
        \SB1_3_28/i1[9] ), .ZN(n4308) );
  NAND3_X2 U8376 ( .A1(\SB1_3_10/i0_3 ), .A2(\SB1_3_10/i0[10] ), .A3(
        \SB1_3_10/i0[9] ), .ZN(\SB1_3_10/Component_Function_4/NAND4_in[2] ) );
  XOR2_X1 U8377 ( .A1(\MC_ARK_ARC_1_1/temp6[78] ), .A2(
        \MC_ARK_ARC_1_1/temp5[78] ), .Z(\MC_ARK_ARC_1_1/buf_output[78] ) );
  NAND4_X2 U8378 ( .A1(n5401), .A2(\SB1_2_3/Component_Function_1/NAND4_in[1] ), 
        .A3(n1465), .A4(\SB1_2_3/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_2_3/buf_output[1] ) );
  NAND4_X2 U8383 ( .A1(\SB1_2_30/Component_Function_3/NAND4_in[1] ), .A2(n5343), .A3(\SB1_2_30/Component_Function_3/NAND4_in[0] ), .A4(n1547), .ZN(
        \SB1_2_30/buf_output[3] ) );
  XOR2_X1 U8384 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[154] ), .A2(\RI5[3][160] ), 
        .Z(n5313) );
  BUF_X4 U8385 ( .I(\SB2_2_31/buf_output[3] ), .Z(\RI5[2][15] ) );
  NAND4_X2 U8387 ( .A1(\SB2_1_17/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_1_17/Component_Function_4/NAND4_in[0] ), .A3(n3334), .A4(n5315), 
        .ZN(\SB2_1_17/buf_output[4] ) );
  NAND3_X1 U8388 ( .A1(\SB2_1_17/i0_0 ), .A2(\SB2_1_17/i3[0] ), .A3(
        \SB2_1_17/i1_7 ), .ZN(n5315) );
  NAND3_X2 U8389 ( .A1(\SB1_2_9/i0_3 ), .A2(\SB1_2_9/i0_4 ), .A3(
        \SB1_2_9/i1[9] ), .ZN(\SB1_2_9/Component_Function_5/NAND4_in[2] ) );
  INV_X2 U8390 ( .I(\RI3[0][93] ), .ZN(\SB2_0_16/i0[8] ) );
  NAND4_X2 U8391 ( .A1(\SB1_0_18/Component_Function_3/NAND4_in[3] ), .A2(
        \SB1_0_18/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_0_18/Component_Function_3/NAND4_in[1] ), .A4(
        \SB1_0_18/Component_Function_3/NAND4_in[2] ), .ZN(\RI3[0][93] ) );
  XOR2_X1 U8394 ( .A1(n5317), .A2(n5316), .Z(n5319) );
  XOR2_X1 U8396 ( .A1(\RI5[0][84] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[48] ), 
        .Z(n5316) );
  XOR2_X1 U8397 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[132] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[138] ), .Z(n5317) );
  NAND4_X2 U8402 ( .A1(n1331), .A2(\SB1_3_10/Component_Function_5/NAND4_in[2] ), .A3(n1329), .A4(n5318), .ZN(\SB1_3_10/buf_output[5] ) );
  NAND3_X2 U8403 ( .A1(\SB1_3_10/i0[10] ), .A2(\SB1_3_10/i0_0 ), .A3(
        \SB1_3_10/i0[6] ), .ZN(n5318) );
  NAND3_X1 U8404 ( .A1(\SB2_1_12/i0_3 ), .A2(\SB2_1_12/i1_7 ), .A3(
        \SB2_1_12/i0[8] ), .ZN(\SB2_1_12/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U8405 ( .A1(n5320), .A2(n63), .Z(Ciphertext[1]) );
  NAND4_X2 U8406 ( .A1(\SB4_31/Component_Function_1/NAND4_in[2] ), .A2(
        \SB4_31/Component_Function_1/NAND4_in[3] ), .A3(
        \SB4_31/Component_Function_1/NAND4_in[1] ), .A4(
        \SB4_31/Component_Function_1/NAND4_in[0] ), .ZN(n5320) );
  NAND4_X2 U8407 ( .A1(\SB2_0_4/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_4/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_4/Component_Function_4/NAND4_in[3] ), .A4(n5321), .ZN(
        \SB2_0_4/buf_output[4] ) );
  NAND3_X2 U8412 ( .A1(\SB2_0_4/i0[10] ), .A2(\SB2_0_4/i0[9] ), .A3(
        \SB2_0_4/i0_3 ), .ZN(n5321) );
  XOR2_X1 U8415 ( .A1(n2798), .A2(n5322), .Z(\MC_ARK_ARC_1_1/buf_output[112] )
         );
  XOR2_X1 U8416 ( .A1(\MC_ARK_ARC_1_1/temp2[112] ), .A2(
        \MC_ARK_ARC_1_1/temp1[112] ), .Z(n5322) );
  XOR2_X1 U8418 ( .A1(n5323), .A2(n38), .Z(Ciphertext[5]) );
  NAND4_X2 U8419 ( .A1(\SB4_31/Component_Function_5/NAND4_in[2] ), .A2(n1238), 
        .A3(n6051), .A4(n2179), .ZN(n5323) );
  XOR2_X1 U8423 ( .A1(\MC_ARK_ARC_1_2/temp1[32] ), .A2(n5324), .Z(n3787) );
  XOR2_X1 U8428 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[68] ), .A2(\RI5[2][98] ), 
        .Z(n5324) );
  XOR2_X1 U8429 ( .A1(n6097), .A2(n5325), .Z(\MC_ARK_ARC_1_1/buf_output[50] )
         );
  XOR2_X1 U8430 ( .A1(\MC_ARK_ARC_1_1/temp4[50] ), .A2(n5465), .Z(n5325) );
  NAND2_X2 U8431 ( .A1(\SB1_3_26/i0_3 ), .A2(\SB1_3_26/i1[9] ), .ZN(
        \SB1_3_26/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 U8432 ( .A1(\SB2_1_5/i0_0 ), .A2(\SB2_1_5/i0[10] ), .A3(
        \SB2_1_5/i0[6] ), .ZN(n5326) );
  XOR2_X1 U8434 ( .A1(\RI5[1][40] ), .A2(\RI5[1][4] ), .Z(
        \MC_ARK_ARC_1_1/temp3[130] ) );
  XOR2_X1 U8435 ( .A1(n5327), .A2(n113), .Z(Ciphertext[23]) );
  NAND4_X2 U8437 ( .A1(\SB4_28/Component_Function_5/NAND4_in[2] ), .A2(n2394), 
        .A3(\SB4_28/Component_Function_5/NAND4_in[1] ), .A4(
        \SB4_28/Component_Function_5/NAND4_in[0] ), .ZN(n5327) );
  XOR2_X1 U8438 ( .A1(\MC_ARK_ARC_1_0/temp5[23] ), .A2(n5328), .Z(
        \MC_ARK_ARC_1_0/buf_output[23] ) );
  XOR2_X1 U8439 ( .A1(\MC_ARK_ARC_1_0/temp4[23] ), .A2(
        \MC_ARK_ARC_1_0/temp3[23] ), .Z(n5328) );
  XOR2_X1 U8441 ( .A1(n5329), .A2(n106), .Z(Ciphertext[115]) );
  NAND4_X2 U8442 ( .A1(\SB4_12/Component_Function_1/NAND4_in[2] ), .A2(
        \SB4_12/Component_Function_1/NAND4_in[1] ), .A3(n2032), .A4(
        \SB4_12/Component_Function_1/NAND4_in[0] ), .ZN(n5329) );
  NAND3_X2 U8445 ( .A1(\SB1_2_29/i1_5 ), .A2(\SB1_2_29/i0_4 ), .A3(
        \SB1_2_29/i0_0 ), .ZN(n5330) );
  XOR2_X1 U8446 ( .A1(\MC_ARK_ARC_1_3/temp4[173] ), .A2(n5331), .Z(n1892) );
  XOR2_X1 U8447 ( .A1(\RI5[3][83] ), .A2(\RI5[3][47] ), .Z(n5331) );
  NAND3_X1 U8448 ( .A1(\SB4_3/i0_3 ), .A2(n5495), .A3(\SB4_3/i1_7 ), .ZN(
        \SB4_3/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U8453 ( .A1(n5332), .A2(n108), .Z(Ciphertext[164]) );
  XOR2_X1 U8454 ( .A1(\MC_ARK_ARC_1_1/temp2[32] ), .A2(n5333), .Z(
        \MC_ARK_ARC_1_1/temp5[32] ) );
  XOR2_X1 U8456 ( .A1(\RI5[1][26] ), .A2(\RI5[1][32] ), .Z(n5333) );
  BUF_X4 U8459 ( .I(\RI1[3][167] ), .Z(\SB1_3_4/i0_3 ) );
  XOR2_X1 U8463 ( .A1(n1568), .A2(n5334), .Z(\MC_ARK_ARC_1_1/buf_output[111] )
         );
  XOR2_X1 U8464 ( .A1(\MC_ARK_ARC_1_1/temp3[111] ), .A2(
        \MC_ARK_ARC_1_1/temp4[111] ), .Z(n5334) );
  NAND4_X2 U8465 ( .A1(\SB3_3/Component_Function_1/NAND4_in[1] ), .A2(
        \SB3_3/Component_Function_1/NAND4_in[0] ), .A3(
        \SB3_3/Component_Function_1/NAND4_in[3] ), .A4(n5335), .ZN(
        \SB3_3/buf_output[1] ) );
  NAND3_X2 U8466 ( .A1(\SB3_3/i0[9] ), .A2(\SB3_3/i1_5 ), .A3(\SB3_3/i0[6] ), 
        .ZN(n5335) );
  NAND2_X2 U8470 ( .A1(\SB1_0_17/i0_3 ), .A2(\SB1_0_17/i1[9] ), .ZN(n5904) );
  NAND4_X2 U8475 ( .A1(\SB1_3_31/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_31/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_3_31/Component_Function_2/NAND4_in[2] ), .A4(n4662), .ZN(n6330)
         );
  NAND3_X2 U8478 ( .A1(\SB1_3_31/i0_4 ), .A2(\SB1_3_31/i0_0 ), .A3(
        \SB1_3_31/i1_5 ), .ZN(n4662) );
  XOR2_X1 U8479 ( .A1(n5337), .A2(n5336), .Z(\MC_ARK_ARC_1_0/temp5[152] ) );
  XOR2_X1 U8481 ( .A1(\RI5[0][98] ), .A2(\RI5[0][152] ), .Z(n5336) );
  XOR2_X1 U8482 ( .A1(\RI5[0][122] ), .A2(\RI5[0][146] ), .Z(n5337) );
  NAND3_X1 U8483 ( .A1(n5495), .A2(\SB4_3/i0[9] ), .A3(\SB3_6/buf_output[2] ), 
        .ZN(\SB4_3/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U8485 ( .A1(n5495), .A2(\SB4_3/i1_5 ), .A3(\SB4_3/i3[0] ), .ZN(
        \SB4_3/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 U8488 ( .A1(\SB2_2_7/i1[9] ), .A2(\SB1_2_8/buf_output[4] ), .A3(
        \SB2_2_7/i0_3 ), .ZN(\SB2_2_7/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U8489 ( .A1(\SB1_0_12/i0[10] ), .A2(\SB1_0_12/i0_3 ), .A3(
        \SB1_0_12/i0[6] ), .ZN(n5338) );
  NAND3_X2 U8490 ( .A1(\SB1_1_12/i0[10] ), .A2(\SB1_1_12/i1_7 ), .A3(
        \SB1_1_12/i1[9] ), .ZN(\SB1_1_12/Component_Function_3/NAND4_in[2] ) );
  NAND4_X2 U8491 ( .A1(\SB1_0_16/Component_Function_5/NAND4_in[2] ), .A2(n3505), .A3(n4315), .A4(\SB1_0_16/Component_Function_5/NAND4_in[0] ), .ZN(
        \RI3[0][95] ) );
  BUF_X4 U8492 ( .I(\SB3_5/buf_output[5] ), .Z(\SB4_5/i0_3 ) );
  NAND4_X2 U8493 ( .A1(\SB1_3_5/Component_Function_5/NAND4_in[2] ), .A2(n5566), 
        .A3(n5481), .A4(\SB1_3_5/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_5/buf_output[5] ) );
  NAND3_X2 U8495 ( .A1(\SB1_1_30/i0_3 ), .A2(\SB1_1_30/i0_0 ), .A3(
        \SB1_1_30/i0_4 ), .ZN(\SB1_1_30/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U8496 ( .A1(n2207), .A2(\MC_ARK_ARC_1_1/temp4[131] ), .Z(n5340) );
  NAND3_X2 U8497 ( .A1(\SB2_2_6/i0[10] ), .A2(n2074), .A3(\SB2_2_6/i0_3 ), 
        .ZN(n3292) );
  NAND4_X2 U8498 ( .A1(\SB1_3_18/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_3_18/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_3_18/Component_Function_1/NAND4_in[3] ), .A4(n5342), .ZN(
        \SB1_3_18/buf_output[1] ) );
  INV_X2 U8499 ( .I(\SB1_2_28/buf_output[3] ), .ZN(\SB2_2_26/i0[8] ) );
  NAND4_X2 U8502 ( .A1(\SB1_2_28/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_28/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_28/Component_Function_3/NAND4_in[3] ), .A4(n3899), .ZN(
        \SB1_2_28/buf_output[3] ) );
  NAND3_X1 U8504 ( .A1(\SB2_2_28/i0_3 ), .A2(\SB2_2_28/i0[8] ), .A3(
        \SB1_2_1/buf_output[0] ), .ZN(
        \SB2_2_28/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U8505 ( .A1(\SB1_2_14/i0_3 ), .A2(\SB1_2_14/i1_7 ), .A3(
        \SB1_2_14/i0[8] ), .ZN(\SB1_2_14/Component_Function_1/NAND4_in[1] ) );
  NAND3_X2 U8506 ( .A1(\SB1_2_30/i0[10] ), .A2(\SB1_2_30/i1[9] ), .A3(
        \SB1_2_30/i1_7 ), .ZN(n5343) );
  NAND4_X2 U8507 ( .A1(\SB4_31/Component_Function_0/NAND4_in[3] ), .A2(
        \SB4_31/Component_Function_0/NAND4_in[2] ), .A3(
        \SB4_31/Component_Function_0/NAND4_in[0] ), .A4(
        \SB4_31/Component_Function_0/NAND4_in[1] ), .ZN(n5354) );
  XOR2_X1 U8508 ( .A1(\MC_ARK_ARC_1_3/temp1[175] ), .A2(n5344), .Z(n5607) );
  XOR2_X1 U8509 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[49] ), .A2(\RI5[3][85] ), 
        .Z(n5344) );
  NAND4_X2 U8510 ( .A1(\SB2_3_6/Component_Function_5/NAND4_in[0] ), .A2(
        \SB2_3_6/Component_Function_5/NAND4_in[2] ), .A3(n5855), .A4(n5345), 
        .ZN(\SB2_3_6/buf_output[5] ) );
  NAND4_X2 U8511 ( .A1(\SB1_3_9/Component_Function_2/NAND4_in[3] ), .A2(n4106), 
        .A3(\SB1_3_9/Component_Function_2/NAND4_in[1] ), .A4(n5346), .ZN(
        \SB1_3_9/buf_output[2] ) );
  NAND4_X2 U8514 ( .A1(\SB2_3_1/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_1/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_3_1/Component_Function_5/NAND4_in[0] ), .A4(n5347), .ZN(
        \SB2_3_1/buf_output[5] ) );
  NAND3_X2 U8516 ( .A1(\SB2_3_1/i0[6] ), .A2(\SB2_3_1/i0_4 ), .A3(
        \SB2_3_1/i0[9] ), .ZN(n5347) );
  NAND3_X2 U8517 ( .A1(\SB1_1_5/i0[6] ), .A2(\SB1_1_5/i1_5 ), .A3(
        \SB1_1_5/i0[9] ), .ZN(\SB1_1_5/Component_Function_1/NAND4_in[2] ) );
  NAND4_X2 U8518 ( .A1(\SB2_3_2/Component_Function_5/NAND4_in[2] ), .A2(n3783), 
        .A3(\SB2_3_2/Component_Function_5/NAND4_in[0] ), .A4(n5348), .ZN(
        \SB2_3_2/buf_output[5] ) );
  NAND3_X2 U8519 ( .A1(\SB2_3_2/i0_0 ), .A2(\SB2_3_2/i0[6] ), .A3(
        \SB2_3_2/i0[10] ), .ZN(n5348) );
  NAND4_X2 U8520 ( .A1(\SB2_3_1/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_3_1/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_3_1/Component_Function_1/NAND4_in[1] ), .A4(n5349), .ZN(
        \SB2_3_1/buf_output[1] ) );
  INV_X1 U8525 ( .I(\SB3_14/buf_output[3] ), .ZN(\SB4_12/i0[8] ) );
  NAND4_X2 U8526 ( .A1(\SB3_14/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_14/Component_Function_3/NAND4_in[1] ), .A3(n5537), .A4(n1979), 
        .ZN(\SB3_14/buf_output[3] ) );
  NAND3_X2 U8532 ( .A1(\SB3_1/i0_0 ), .A2(\SB3_1/i0_4 ), .A3(\SB3_1/i0_3 ), 
        .ZN(\SB3_1/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U8533 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[154] ), .A2(\RI5[3][130] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[184] ) );
  XOR2_X1 U8534 ( .A1(n5350), .A2(n197), .Z(Ciphertext[158]) );
  NAND4_X2 U8536 ( .A1(\SB4_5/Component_Function_2/NAND4_in[0] ), .A2(n2522), 
        .A3(n6114), .A4(n5663), .ZN(n5350) );
  NAND3_X2 U8539 ( .A1(\SB1_2_30/i1[9] ), .A2(\SB1_2_30/i0_3 ), .A3(
        \SB1_2_30/i0[6] ), .ZN(\SB1_2_30/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U8544 ( .A1(\SB2_0_5/i0_3 ), .A2(\SB2_0_5/i0[8] ), .A3(
        \RI3[0][156] ), .ZN(\SB2_0_5/Component_Function_2/NAND4_in[2] ) );
  BUF_X4 U8545 ( .I(\SB3_7/buf_output[0] ), .Z(\SB4_2/i0[9] ) );
  NAND3_X1 U8547 ( .A1(\SB2_0_27/i0[10] ), .A2(\SB2_0_27/i0_3 ), .A3(
        \SB2_0_27/i0_4 ), .ZN(n2189) );
  XOR2_X1 U8548 ( .A1(\RI5[1][175] ), .A2(\RI5[1][55] ), .Z(n5629) );
  NAND4_X2 U8550 ( .A1(\SB1_2_4/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_2_4/Component_Function_2/NAND4_in[0] ), .A3(n5375), .A4(n4326), 
        .ZN(\SB1_2_4/buf_output[2] ) );
  NAND3_X2 U8553 ( .A1(\SB2_3_17/i0[6] ), .A2(\SB2_3_17/i0_4 ), .A3(
        \SB2_3_17/i0[9] ), .ZN(\SB2_3_17/Component_Function_5/NAND4_in[3] ) );
  XOR2_X1 U8555 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[185] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[149] ), .Z(n3129) );
  NAND4_X2 U8560 ( .A1(\SB3_2/Component_Function_5/NAND4_in[1] ), .A2(n5572), 
        .A3(n4136), .A4(\SB3_2/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB3_2/buf_output[5] ) );
  NAND3_X1 U8563 ( .A1(\SB2_0_27/i0_3 ), .A2(\SB2_0_27/i1[9] ), .A3(
        \SB2_0_27/i0[6] ), .ZN(\SB2_0_27/Component_Function_3/NAND4_in[0] ) );
  NAND4_X2 U8565 ( .A1(\SB1_2_25/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_2_25/Component_Function_5/NAND4_in[0] ), .A3(
        \SB1_2_25/Component_Function_5/NAND4_in[1] ), .A4(n5351), .ZN(
        \SB1_2_25/buf_output[5] ) );
  NAND3_X2 U8566 ( .A1(\SB1_2_25/i0_4 ), .A2(\SB1_2_25/i0[9] ), .A3(
        \SB1_2_25/i0[6] ), .ZN(n5351) );
  NAND3_X2 U8567 ( .A1(\SB2_3_7/i0_3 ), .A2(\SB1_3_8/buf_output[4] ), .A3(
        \SB2_3_7/i1[9] ), .ZN(\SB2_3_7/Component_Function_5/NAND4_in[2] ) );
  INV_X2 U8568 ( .I(\SB1_2_25/buf_output[5] ), .ZN(\SB2_2_25/i1_5 ) );
  NAND3_X2 U8572 ( .A1(\SB1_2_27/i0[10] ), .A2(\SB1_2_27/i1[9] ), .A3(
        \SB1_2_27/i1_7 ), .ZN(n3522) );
  NAND4_X2 U8573 ( .A1(\SB2_1_29/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_1_29/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_1_29/Component_Function_3/NAND4_in[3] ), .A4(n5352), .ZN(
        \SB2_1_29/buf_output[3] ) );
  NAND3_X2 U8574 ( .A1(\SB2_1_29/i0[10] ), .A2(\SB2_1_29/i1[9] ), .A3(
        \SB2_1_29/i1_7 ), .ZN(n5352) );
  NAND3_X1 U8575 ( .A1(\SB2_3_12/i0_4 ), .A2(\SB2_3_12/i1_7 ), .A3(n3651), 
        .ZN(n5353) );
  NAND3_X2 U8576 ( .A1(\SB4_5/i0_0 ), .A2(\SB4_5/i0_3 ), .A3(\SB4_5/i0[7] ), 
        .ZN(n2030) );
  XOR2_X1 U8577 ( .A1(n5354), .A2(n60), .Z(Ciphertext[0]) );
  NAND4_X2 U8578 ( .A1(n3224), .A2(\SB4_23/Component_Function_4/NAND4_in[2] ), 
        .A3(n2705), .A4(n5356), .ZN(n5604) );
  NAND3_X1 U8579 ( .A1(\SB4_23/i0_0 ), .A2(\SB4_23/i0[9] ), .A3(\SB4_23/i0[8] ), .ZN(n5356) );
  BUF_X4 U8581 ( .I(\MC_ARK_ARC_1_1/buf_output[179] ), .Z(\SB1_2_2/i0_3 ) );
  NAND4_X2 U8583 ( .A1(\SB4_26/Component_Function_0/NAND4_in[1] ), .A2(
        \SB4_26/Component_Function_0/NAND4_in[3] ), .A3(n1709), .A4(n5357), 
        .ZN(n3112) );
  XOR2_X1 U8587 ( .A1(n5358), .A2(n67), .Z(Ciphertext[41]) );
  NAND4_X2 U8588 ( .A1(\SB4_25/Component_Function_5/NAND4_in[3] ), .A2(
        \SB4_25/Component_Function_5/NAND4_in[2] ), .A3(
        \SB4_25/Component_Function_5/NAND4_in[1] ), .A4(
        \SB4_25/Component_Function_5/NAND4_in[0] ), .ZN(n5358) );
  XOR2_X1 U8590 ( .A1(\MC_ARK_ARC_1_3/temp6[32] ), .A2(
        \MC_ARK_ARC_1_3/temp5[32] ), .Z(n1384) );
  XOR2_X1 U8591 ( .A1(\MC_ARK_ARC_1_3/temp4[32] ), .A2(
        \MC_ARK_ARC_1_3/temp3[32] ), .Z(\MC_ARK_ARC_1_3/temp6[32] ) );
  XOR2_X1 U8593 ( .A1(n5359), .A2(n109), .Z(Ciphertext[40]) );
  NAND4_X2 U8594 ( .A1(\SB4_25/Component_Function_4/NAND4_in[3] ), .A2(n2839), 
        .A3(\SB4_25/Component_Function_4/NAND4_in[1] ), .A4(
        \SB4_25/Component_Function_4/NAND4_in[0] ), .ZN(n5359) );
  NAND3_X1 U8596 ( .A1(\SB2_3_20/i0[7] ), .A2(\SB2_3_20/i0[6] ), .A3(
        \SB2_3_20/i0[8] ), .ZN(\SB2_3_20/Component_Function_0/NAND4_in[1] ) );
  BUF_X4 U8597 ( .I(\MC_ARK_ARC_1_1/buf_output[111] ), .Z(\SB1_2_13/i0[10] )
         );
  XOR2_X1 U8599 ( .A1(\MC_ARK_ARC_1_1/temp2[100] ), .A2(n5360), .Z(n3486) );
  XOR2_X1 U8600 ( .A1(\RI5[1][94] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[100] ), 
        .Z(n5360) );
  NAND2_X1 U8604 ( .A1(\SB3_10/i3[0] ), .A2(\SB3_10/i0_0 ), .ZN(n1765) );
  XOR2_X1 U8607 ( .A1(n5361), .A2(n235), .Z(Ciphertext[129]) );
  NAND4_X2 U8608 ( .A1(n6428), .A2(\SB4_10/Component_Function_3/NAND4_in[3] ), 
        .A3(n4283), .A4(\SB4_10/Component_Function_3/NAND4_in[2] ), .ZN(n5361)
         );
  NAND3_X2 U8609 ( .A1(\SB2_3_20/i1[9] ), .A2(\SB2_3_20/i0_4 ), .A3(
        \SB2_3_20/i0_3 ), .ZN(\SB2_3_20/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U8629 ( .A1(n5362), .A2(n6457), .Z(\MC_ARK_ARC_1_2/temp5[161] ) );
  XOR2_X1 U8638 ( .A1(\RI5[2][161] ), .A2(\RI5[2][155] ), .Z(n5362) );
  XOR2_X1 U8639 ( .A1(n5363), .A2(n136), .Z(Ciphertext[73]) );
  NAND4_X2 U8640 ( .A1(\SB4_19/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_19/Component_Function_1/NAND4_in[3] ), .A3(
        \SB4_19/Component_Function_1/NAND4_in[2] ), .A4(
        \SB4_19/Component_Function_1/NAND4_in[0] ), .ZN(n5363) );
  NAND3_X2 U8648 ( .A1(\SB1_3_29/i1_7 ), .A2(\SB1_3_29/i0[8] ), .A3(
        \SB1_3_29/i0_4 ), .ZN(\SB1_3_29/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 U8651 ( .A1(\SB2_1_5/i0[10] ), .A2(\SB2_1_5/i0_3 ), .A3(
        \SB2_1_5/i0[6] ), .ZN(n5365) );
  XOR2_X1 U8652 ( .A1(n5366), .A2(n2470), .Z(\MC_ARK_ARC_1_2/buf_output[188] )
         );
  XOR2_X1 U8657 ( .A1(\MC_ARK_ARC_1_1/temp3[9] ), .A2(
        \MC_ARK_ARC_1_1/temp4[9] ), .Z(n6076) );
  NAND3_X2 U8659 ( .A1(\SB2_3_22/i0_3 ), .A2(\SB2_3_22/i0[6] ), .A3(
        \SB2_3_22/i1[9] ), .ZN(\SB2_3_22/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U8660 ( .A1(n6520), .A2(\MC_ARK_ARC_1_1/temp6[176] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[176] ) );
  NAND3_X1 U8662 ( .A1(\SB1_2_25/i0_3 ), .A2(\SB1_2_25/i0[8] ), .A3(
        \SB1_2_25/i1_7 ), .ZN(\SB1_2_25/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U8670 ( .A1(n5751), .A2(n5367), .Z(n5453) );
  XOR2_X1 U8671 ( .A1(\RI5[1][39] ), .A2(\RI5[1][45] ), .Z(n5367) );
  XOR2_X1 U8674 ( .A1(\MC_ARK_ARC_1_1/temp4[22] ), .A2(n5368), .Z(
        \MC_ARK_ARC_1_1/temp6[22] ) );
  XOR2_X1 U8676 ( .A1(\RI5[1][124] ), .A2(\RI5[1][88] ), .Z(n5368) );
  NAND3_X2 U8678 ( .A1(\SB2_2_22/i0[10] ), .A2(\SB2_2_22/i0_3 ), .A3(
        \SB2_2_22/i0_4 ), .ZN(n5556) );
  NAND3_X2 U8683 ( .A1(\SB2_0_12/i0_3 ), .A2(\SB2_0_12/i0_4 ), .A3(
        \SB2_0_12/i1[9] ), .ZN(n3089) );
  NAND4_X2 U8688 ( .A1(\SB1_1_4/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_1_4/Component_Function_1/NAND4_in[0] ), .A3(
        \SB1_1_4/Component_Function_1/NAND4_in[3] ), .A4(n5369), .ZN(
        \SB1_1_4/buf_output[1] ) );
  NAND3_X1 U8690 ( .A1(\SB1_1_4/i0[6] ), .A2(\SB1_1_4/i1_5 ), .A3(
        \SB1_1_4/i0[9] ), .ZN(n5369) );
  NAND3_X1 U8691 ( .A1(\SB2_0_5/i0_3 ), .A2(\SB2_0_5/i0[10] ), .A3(
        \RI3[0][160] ), .ZN(\SB2_0_5/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U8692 ( .A1(\MC_ARK_ARC_1_2/temp1[152] ), .A2(n5370), .Z(n4145) );
  XOR2_X1 U8696 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[122] ), .A2(\RI5[2][98] ), 
        .Z(n5370) );
  NAND4_X2 U8698 ( .A1(\SB1_1_21/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_1_21/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_1_21/Component_Function_5/NAND4_in[0] ), .A4(n5371), .ZN(
        \SB1_1_21/buf_output[5] ) );
  NAND3_X2 U8699 ( .A1(\SB1_1_21/i0_4 ), .A2(\SB1_1_21/i0[6] ), .A3(
        \SB1_1_21/i0[9] ), .ZN(n5371) );
  NAND3_X2 U8703 ( .A1(\SB1_3_5/i0[9] ), .A2(\SB1_3_5/i0[8] ), .A3(
        \SB1_3_5/i0_3 ), .ZN(n5372) );
  XOR2_X1 U8704 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[166] ), .A2(\RI5[0][130] ), 
        .Z(n6267) );
  XOR2_X1 U8710 ( .A1(n5374), .A2(n5373), .Z(n2509) );
  XOR2_X1 U8718 ( .A1(\RI5[0][75] ), .A2(n214), .Z(n5373) );
  XOR2_X1 U8723 ( .A1(\RI5[0][9] ), .A2(\RI5[0][39] ), .Z(n5374) );
  NAND3_X2 U8724 ( .A1(\SB1_2_4/i0_3 ), .A2(\SB1_2_4/i0[6] ), .A3(
        \SB1_2_4/i0[10] ), .ZN(n5375) );
  NAND3_X1 U8725 ( .A1(\SB3_1/i0_3 ), .A2(\SB3_1/i0[8] ), .A3(\SB3_1/i1_7 ), 
        .ZN(n5376) );
  NAND3_X1 U8733 ( .A1(\SB1_1_3/i0[8] ), .A2(\SB1_1_3/i3[0] ), .A3(
        \SB1_1_3/i1_5 ), .ZN(\SB1_1_3/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U8736 ( .A1(n3052), .A2(n5378), .Z(\MC_ARK_ARC_1_3/buf_output[80] )
         );
  XOR2_X1 U8742 ( .A1(n5873), .A2(n5776), .Z(n5378) );
  NAND3_X1 U8744 ( .A1(\SB1_3_0/i0_4 ), .A2(\SB1_3_0/i1_7 ), .A3(
        \SB1_3_0/i0[8] ), .ZN(\SB1_3_0/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U8747 ( .A1(n4471), .A2(\SB1_3_27/Component_Function_3/NAND4_in[1] ), .A3(n4383), .A4(n5379), .ZN(\SB1_3_27/buf_output[3] ) );
  NAND3_X2 U8748 ( .A1(\SB4_2/i0_3 ), .A2(\SB4_2/i0_0 ), .A3(\SB4_2/i0[7] ), 
        .ZN(n6075) );
  XOR2_X1 U8751 ( .A1(\MC_ARK_ARC_1_2/temp1[58] ), .A2(n5380), .Z(n2371) );
  XOR2_X1 U8752 ( .A1(\RI5[2][28] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[4] ), 
        .Z(n5380) );
  XOR2_X1 U8753 ( .A1(n5381), .A2(n129), .Z(Ciphertext[67]) );
  NAND4_X2 U8754 ( .A1(\SB4_20/Component_Function_1/NAND4_in[3] ), .A2(
        \SB4_20/Component_Function_1/NAND4_in[1] ), .A3(
        \SB4_20/Component_Function_1/NAND4_in[0] ), .A4(
        \SB4_20/Component_Function_1/NAND4_in[2] ), .ZN(n5381) );
  NAND3_X2 U8757 ( .A1(\SB1_2_20/i0[10] ), .A2(\SB1_2_20/i1[9] ), .A3(
        \SB1_2_20/i1_7 ), .ZN(n5482) );
  NAND4_X2 U8762 ( .A1(n1211), .A2(n3631), .A3(
        \SB2_1_17/Component_Function_5/NAND4_in[0] ), .A4(n5382), .ZN(
        \SB2_1_17/buf_output[5] ) );
  NAND3_X2 U8765 ( .A1(\SB2_1_17/i0_0 ), .A2(\SB2_1_17/i0[10] ), .A3(
        \SB2_1_17/i0[6] ), .ZN(n5382) );
  NAND4_X2 U8766 ( .A1(\SB2_1_1/Component_Function_2/NAND4_in[0] ), .A2(n1269), 
        .A3(n3244), .A4(n5383), .ZN(\SB2_1_1/buf_output[2] ) );
  NAND3_X2 U8770 ( .A1(\SB2_1_1/i0[10] ), .A2(\SB2_1_1/i0_3 ), .A3(
        \SB2_1_1/i0[6] ), .ZN(n5383) );
  INV_X2 U8771 ( .I(\SB1_3_1/buf_output[3] ), .ZN(\SB2_3_31/i0[8] ) );
  NAND4_X2 U8776 ( .A1(\SB1_3_1/Component_Function_3/NAND4_in[0] ), .A2(n3934), 
        .A3(\SB1_3_1/Component_Function_3/NAND4_in[1] ), .A4(n1730), .ZN(
        \SB1_3_1/buf_output[3] ) );
  XOR2_X1 U8777 ( .A1(n5385), .A2(n5384), .Z(n2435) );
  XOR2_X1 U8779 ( .A1(\RI5[0][43] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[73] ), 
        .Z(n5384) );
  NAND3_X1 U8785 ( .A1(\SB1_1_25/i0[10] ), .A2(\SB1_1_25/i0_3 ), .A3(
        \SB1_1_25/i0[6] ), .ZN(\SB1_1_25/Component_Function_2/NAND4_in[1] ) );
  BUF_X4 U8786 ( .I(\SB1_2_30/buf_output[5] ), .Z(\SB2_2_30/i0_3 ) );
  NAND3_X2 U8787 ( .A1(\SB2_0_22/i0_3 ), .A2(\SB2_0_22/i0[8] ), .A3(
        \RI3[0][54] ), .ZN(\SB2_0_22/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U8788 ( .A1(\SB2_3_4/i0[10] ), .A2(\SB2_3_4/i0_3 ), .A3(
        \SB2_3_4/i0_4 ), .ZN(\SB2_3_4/Component_Function_0/NAND4_in[2] ) );
  NAND3_X2 U8792 ( .A1(\RI3[0][4] ), .A2(\SB2_0_31/i0[6] ), .A3(
        \SB2_0_31/i0[9] ), .ZN(n5386) );
  NAND4_X2 U8795 ( .A1(\SB1_3_24/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_3_24/Component_Function_1/NAND4_in[1] ), .A3(n1498), .A4(n5387), 
        .ZN(\SB1_3_24/buf_output[1] ) );
  NAND2_X1 U8796 ( .A1(\SB1_3_24/i0_3 ), .A2(\SB1_3_24/i1[9] ), .ZN(n5387) );
  NAND4_X2 U8797 ( .A1(\SB2_0_31/Component_Function_3/NAND4_in[3] ), .A2(
        \SB2_0_31/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_0_31/Component_Function_3/NAND4_in[0] ), .A4(n5388), .ZN(
        \SB2_0_31/buf_output[3] ) );
  NAND3_X1 U8798 ( .A1(\RI3[0][4] ), .A2(\SB2_0_31/i0_0 ), .A3(\SB2_0_31/i0_3 ), .ZN(n5388) );
  XOR2_X1 U8799 ( .A1(n6442), .A2(n5389), .Z(n1354) );
  XOR2_X1 U8803 ( .A1(n5390), .A2(n31), .Z(Ciphertext[137]) );
  NAND4_X2 U8805 ( .A1(\SB4_9/Component_Function_5/NAND4_in[1] ), .A2(
        \SB4_9/Component_Function_5/NAND4_in[2] ), .A3(
        \SB4_9/Component_Function_5/NAND4_in[0] ), .A4(
        \SB4_9/Component_Function_5/NAND4_in[3] ), .ZN(n5390) );
  XOR2_X1 U8806 ( .A1(\RI5[2][15] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[183] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[45] ) );
  NAND3_X2 U8807 ( .A1(\SB1_2_31/i0_3 ), .A2(\SB1_2_31/i0[8] ), .A3(
        \SB1_2_31/i0[9] ), .ZN(n5391) );
  NAND3_X2 U8808 ( .A1(\SB4_2/i1_5 ), .A2(\SB4_2/i0_0 ), .A3(\SB4_2/i0_4 ), 
        .ZN(\SB4_2/Component_Function_2/NAND4_in[3] ) );
  XOR2_X1 U8810 ( .A1(\RI5[0][26] ), .A2(\RI5[0][62] ), .Z(
        \MC_ARK_ARC_1_0/temp3[152] ) );
  NAND3_X2 U8815 ( .A1(\SB1_2_30/i0_0 ), .A2(\SB1_2_30/i0[10] ), .A3(
        \SB1_2_30/i0[6] ), .ZN(n2724) );
  XOR2_X1 U8816 ( .A1(n2355), .A2(n6244), .Z(\MC_ARK_ARC_1_3/buf_output[188] )
         );
  BUF_X4 U8824 ( .I(\SB1_1_8/buf_output[2] ), .Z(\SB2_1_5/i0_0 ) );
  NAND3_X1 U8829 ( .A1(\SB1_2_26/i0_0 ), .A2(\MC_ARK_ARC_1_1/buf_output[34] ), 
        .A3(\RI1[2][35] ), .ZN(n4488) );
  NAND4_X2 U8831 ( .A1(n2095), .A2(n699), .A3(n5462), .A4(
        \SB1_1_6/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_6/buf_output[5] ) );
  NAND4_X2 U8835 ( .A1(\SB3_5/Component_Function_2/NAND4_in[2] ), .A2(
        \SB3_5/Component_Function_2/NAND4_in[3] ), .A3(n5745), .A4(n6361), 
        .ZN(\SB3_5/buf_output[2] ) );
  NAND4_X2 U8836 ( .A1(n2519), .A2(n2529), .A3(
        \SB4_31/Component_Function_2/NAND4_in[2] ), .A4(n5392), .ZN(n5685) );
  NAND3_X1 U8840 ( .A1(\SB4_31/i0[10] ), .A2(\SB4_31/i1[9] ), .A3(
        \SB4_31/i1_5 ), .ZN(n5392) );
  NAND4_X2 U8849 ( .A1(n2239), .A2(n2189), .A3(
        \SB2_0_27/Component_Function_0/NAND4_in[3] ), .A4(
        \SB2_0_27/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_0_27/buf_output[0] ) );
  XOR2_X1 U8851 ( .A1(n3635), .A2(n3634), .Z(\MC_ARK_ARC_1_2/buf_output[26] )
         );
  NAND3_X2 U8853 ( .A1(\SB2_3_30/i0_3 ), .A2(\SB2_3_30/i0[8] ), .A3(
        \SB2_3_30/i0[9] ), .ZN(\SB2_3_30/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 U8854 ( .A1(\SB2_3_2/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_3_2/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_3_2/Component_Function_0/NAND4_in[0] ), .A4(n5393), .ZN(
        \SB2_3_2/buf_output[0] ) );
  NAND4_X2 U8857 ( .A1(n1951), .A2(\SB2_3_15/Component_Function_3/NAND4_in[3] ), .A3(\SB2_3_15/Component_Function_3/NAND4_in[1] ), .A4(
        \SB2_3_15/Component_Function_3/NAND4_in[0] ), .ZN(
        \SB2_3_15/buf_output[3] ) );
  NAND4_X2 U8864 ( .A1(\SB1_2_25/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_25/Component_Function_3/NAND4_in[1] ), .A3(n6062), .A4(
        \SB1_2_25/Component_Function_3/NAND4_in[2] ), .ZN(
        \SB1_2_25/buf_output[3] ) );
  XOR2_X1 U8865 ( .A1(n6041), .A2(\MC_ARK_ARC_1_3/temp4[161] ), .Z(n1729) );
  NAND3_X2 U8869 ( .A1(\SB2_3_4/i0[6] ), .A2(n5519), .A3(\SB2_3_4/i0[9] ), 
        .ZN(n4139) );
  NAND4_X2 U8870 ( .A1(\SB3_3/Component_Function_5/NAND4_in[1] ), .A2(n2191), 
        .A3(\SB3_3/Component_Function_5/NAND4_in[2] ), .A4(
        \SB3_3/Component_Function_5/NAND4_in[0] ), .ZN(\SB3_3/buf_output[5] )
         );
  XOR2_X1 U8876 ( .A1(\RI5[1][166] ), .A2(\RI5[1][10] ), .Z(
        \MC_ARK_ARC_1_1/temp3[100] ) );
  NAND3_X1 U8880 ( .A1(\SB3_24/i0_4 ), .A2(\SB3_24/i1_7 ), .A3(\SB3_24/i0[8] ), 
        .ZN(n4173) );
  NAND3_X2 U8887 ( .A1(\SB2_2_30/i0_3 ), .A2(\SB2_2_30/i0_0 ), .A3(n2343), 
        .ZN(\SB2_2_30/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U8890 ( .A1(\SB2_3_23/i0_3 ), .A2(\SB2_3_23/i1[9] ), .A3(
        \SB2_3_23/i0[6] ), .ZN(\SB2_3_23/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U8891 ( .A1(\SB2_2_23/i0[10] ), .A2(\SB2_2_23/i0[6] ), .A3(
        \SB2_2_23/i0_0 ), .ZN(\SB2_2_23/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U8893 ( .A1(n5395), .A2(n5394), .Z(n4309) );
  XOR2_X1 U8897 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[110] ), .A2(n31), .Z(n5394) );
  XOR2_X1 U8898 ( .A1(\RI5[1][146] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[80] ), 
        .Z(n5395) );
  XOR2_X1 U8904 ( .A1(n1531), .A2(\MC_ARK_ARC_1_3/temp5[44] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[44] ) );
  XOR2_X1 U8907 ( .A1(\MC_ARK_ARC_1_3/temp4[44] ), .A2(n4211), .Z(n1531) );
  NAND4_X2 U8911 ( .A1(\SB3_24/Component_Function_4/NAND4_in[2] ), .A2(
        \SB3_24/Component_Function_4/NAND4_in[1] ), .A3(n2633), .A4(n5396), 
        .ZN(\SB3_24/buf_output[4] ) );
  NAND3_X2 U8914 ( .A1(\SB1_1_12/i0_3 ), .A2(\SB1_1_12/i1[9] ), .A3(
        \SB1_1_12/i0[6] ), .ZN(n6157) );
  XOR2_X1 U8915 ( .A1(n5397), .A2(n186), .Z(Ciphertext[14]) );
  NAND4_X2 U8917 ( .A1(\SB4_29/Component_Function_2/NAND4_in[0] ), .A2(
        \SB4_29/Component_Function_2/NAND4_in[3] ), .A3(
        \SB4_29/Component_Function_2/NAND4_in[2] ), .A4(n6140), .ZN(n5397) );
  XOR2_X1 U8918 ( .A1(\MC_ARK_ARC_1_2/temp5[44] ), .A2(n5398), .Z(
        \MC_ARK_ARC_1_2/buf_output[44] ) );
  XOR2_X1 U8932 ( .A1(\MC_ARK_ARC_1_2/temp4[42] ), .A2(
        \MC_ARK_ARC_1_2/temp3[42] ), .Z(\MC_ARK_ARC_1_2/temp6[42] ) );
  XOR2_X1 U8933 ( .A1(\RI5[0][9] ), .A2(\RI5[0][33] ), .Z(n5399) );
  XOR2_X1 U8936 ( .A1(n4041), .A2(n5400), .Z(\MC_ARK_ARC_1_3/buf_output[85] )
         );
  XOR2_X1 U8941 ( .A1(\MC_ARK_ARC_1_3/temp2[85] ), .A2(
        \MC_ARK_ARC_1_3/temp1[85] ), .Z(n5400) );
  NAND3_X1 U8946 ( .A1(\SB1_2_3/i0_4 ), .A2(\SB1_2_3/i1_7 ), .A3(
        \SB1_2_3/i0[8] ), .ZN(n5401) );
  NAND3_X2 U8947 ( .A1(\SB2_3_22/i0[10] ), .A2(\SB2_3_22/i1[9] ), .A3(
        \SB2_3_22/i1_7 ), .ZN(\SB2_3_22/Component_Function_3/NAND4_in[2] ) );
  AND2_X1 U8948 ( .A1(\SB2_1_8/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_8/Component_Function_1/NAND4_in[2] ), .Z(n5402) );
  XOR2_X1 U8952 ( .A1(\MC_ARK_ARC_1_1/temp4[177] ), .A2(n5403), .Z(n2854) );
  XOR2_X1 U8954 ( .A1(\RI5[1][87] ), .A2(\RI5[1][51] ), .Z(n5403) );
  NAND2_X2 U8957 ( .A1(\SB2_2_14/i0_3 ), .A2(\SB2_2_14/i1[9] ), .ZN(
        \SB2_2_14/Component_Function_1/NAND4_in[0] ) );
  NAND3_X2 U8958 ( .A1(\SB1_2_2/i0_0 ), .A2(\SB1_2_2/i0[6] ), .A3(
        \SB1_2_2/i0[10] ), .ZN(\SB1_2_2/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U8960 ( .A1(\MC_ARK_ARC_1_1/temp5[175] ), .A2(n5404), .Z(
        \MC_ARK_ARC_1_1/buf_output[175] ) );
  XOR2_X1 U8971 ( .A1(\MC_ARK_ARC_1_1/temp3[175] ), .A2(
        \MC_ARK_ARC_1_1/temp4[175] ), .Z(n5404) );
  BUF_X4 U8974 ( .I(\MC_ARK_ARC_1_3/buf_output[161] ), .Z(\SB3_5/i0_3 ) );
  NAND3_X2 U8977 ( .A1(\SB1_3_15/i0[9] ), .A2(\SB1_3_15/i0[6] ), .A3(
        \SB1_3_15/i0_4 ), .ZN(\SB1_3_15/Component_Function_5/NAND4_in[3] ) );
  XOR2_X1 U8978 ( .A1(\RI5[1][157] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[163] ), 
        .Z(n3039) );
  NAND2_X2 U8991 ( .A1(\SB4_18/i0_3 ), .A2(\SB4_18/i1[9] ), .ZN(
        \SB4_18/Component_Function_1/NAND4_in[0] ) );
  XOR2_X1 U8999 ( .A1(\MC_ARK_ARC_1_2/temp6[96] ), .A2(n5405), .Z(
        \MC_ARK_ARC_1_2/buf_output[96] ) );
  XOR2_X1 U9000 ( .A1(\MC_ARK_ARC_1_2/temp1[96] ), .A2(
        \MC_ARK_ARC_1_2/temp2[96] ), .Z(n5405) );
  NAND3_X1 U9003 ( .A1(\SB2_3_31/i0[6] ), .A2(\SB1_3_4/buf_output[0] ), .A3(
        \SB1_3_0/buf_output[4] ), .ZN(n5406) );
  NAND3_X2 U9006 ( .A1(\SB3_0/i0_3 ), .A2(\SB3_0/i0[8] ), .A3(\SB3_0/i0[9] ), 
        .ZN(n675) );
  XOR2_X1 U9007 ( .A1(\MC_ARK_ARC_1_2/temp5[172] ), .A2(
        \MC_ARK_ARC_1_2/temp6[172] ), .Z(\MC_ARK_ARC_1_2/buf_output[172] ) );
  NAND3_X2 U9010 ( .A1(\SB2_2_30/i0_3 ), .A2(\SB2_2_30/i0[10] ), .A3(n2343), 
        .ZN(n6478) );
  XOR2_X1 U9014 ( .A1(n3344), .A2(n5407), .Z(\MC_ARK_ARC_1_1/buf_output[191] )
         );
  XOR2_X1 U9019 ( .A1(n5451), .A2(n5760), .Z(n5407) );
  INV_X2 U9022 ( .I(\SB1_2_12/buf_output[2] ), .ZN(\SB2_2_9/i1[9] ) );
  NAND4_X2 U9023 ( .A1(n2260), .A2(n4050), .A3(
        \SB1_2_12/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_2_12/Component_Function_2/NAND4_in[0] ), .ZN(
        \SB1_2_12/buf_output[2] ) );
  NAND4_X2 U9038 ( .A1(\SB1_1_29/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_1_29/Component_Function_2/NAND4_in[0] ), .A3(n1567), .A4(n5408), 
        .ZN(\SB1_1_29/buf_output[2] ) );
  INV_X2 U9042 ( .I(\SB1_3_16/buf_output[3] ), .ZN(\SB2_3_14/i0[8] ) );
  NAND4_X2 U9043 ( .A1(\SB1_3_16/Component_Function_3/NAND4_in[1] ), .A2(n6382), .A3(n4616), .A4(\SB1_3_16/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_3_16/buf_output[3] ) );
  NAND4_X2 U9044 ( .A1(\SB2_0_18/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_0_18/Component_Function_0/NAND4_in[2] ), .A3(n836), .A4(n5409), 
        .ZN(\SB2_0_18/buf_output[0] ) );
  NAND2_X2 U9045 ( .A1(\SB2_0_18/i0[9] ), .A2(\SB2_0_18/i0[10] ), .ZN(n5409)
         );
  NAND4_X2 U9047 ( .A1(\SB3_2/Component_Function_2/NAND4_in[1] ), .A2(n5669), 
        .A3(n2313), .A4(n6215), .ZN(\SB3_2/buf_output[2] ) );
  NAND3_X2 U9048 ( .A1(\SB2_2_14/i0_3 ), .A2(\SB2_2_14/i0[10] ), .A3(
        \SB2_2_14/i0[6] ), .ZN(n3029) );
  XOR2_X1 U9053 ( .A1(\MC_ARK_ARC_1_3/temp1[35] ), .A2(n5410), .Z(
        \MC_ARK_ARC_1_3/temp5[35] ) );
  XOR2_X1 U9055 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[5] ), .A2(\RI5[3][173] ), 
        .Z(n5410) );
  NAND4_X2 U9059 ( .A1(\SB4_23/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_23/Component_Function_0/NAND4_in[3] ), .A3(
        \SB4_23/Component_Function_0/NAND4_in[0] ), .A4(
        \SB4_23/Component_Function_0/NAND4_in[1] ), .ZN(n5916) );
  XOR2_X1 U9061 ( .A1(n5411), .A2(n176), .Z(Ciphertext[64]) );
  NAND4_X2 U9064 ( .A1(n4643), .A2(\SB4_21/Component_Function_4/NAND4_in[3] ), 
        .A3(\SB4_21/Component_Function_4/NAND4_in[1] ), .A4(n1517), .ZN(n5411)
         );
  INV_X1 U9067 ( .I(\SB1_1_22/buf_output[0] ), .ZN(\SB2_1_17/i3[0] ) );
  NAND4_X2 U9071 ( .A1(\SB1_1_22/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_1_22/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_1_22/Component_Function_0/NAND4_in[0] ), .A4(
        \SB1_1_22/Component_Function_0/NAND4_in[3] ), .ZN(
        \SB1_1_22/buf_output[0] ) );
  NAND4_X2 U9072 ( .A1(\SB2_0_1/Component_Function_1/NAND4_in[1] ), .A2(n5412), 
        .A3(\SB2_0_1/Component_Function_1/NAND4_in[3] ), .A4(
        \SB2_0_1/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_0_1/buf_output[1] ) );
  INV_X2 U9073 ( .I(\SB1_1_8/buf_output[5] ), .ZN(\SB2_1_8/i1_5 ) );
  NAND4_X2 U9074 ( .A1(\SB1_2_27/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_2_27/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_2_27/Component_Function_4/NAND4_in[2] ), .A4(n5413), .ZN(
        \SB1_2_27/buf_output[4] ) );
  XOR2_X1 U9076 ( .A1(n5414), .A2(n208), .Z(Ciphertext[86]) );
  NAND4_X2 U9079 ( .A1(\SB4_17/Component_Function_2/NAND4_in[1] ), .A2(n4352), 
        .A3(n3564), .A4(\SB4_17/Component_Function_2/NAND4_in[2] ), .ZN(n5414)
         );
  NAND3_X2 U9080 ( .A1(\SB1_0_22/i0_0 ), .A2(\SB1_0_22/i0[10] ), .A3(
        \SB1_0_22/i0[6] ), .ZN(n5415) );
  NAND3_X2 U9081 ( .A1(\SB1_2_21/i0[6] ), .A2(\SB1_2_21/i0_3 ), .A3(
        \SB1_2_21/i0[10] ), .ZN(n5416) );
  NAND3_X2 U9082 ( .A1(\SB2_1_8/i3[0] ), .A2(\SB2_1_8/i0[8] ), .A3(
        \SB2_1_8/i1_5 ), .ZN(\SB2_1_8/Component_Function_3/NAND4_in[3] ) );
  INV_X1 U9083 ( .I(\SB3_6/buf_output[3] ), .ZN(\SB4_4/i0[8] ) );
  NAND4_X2 U9084 ( .A1(\SB3_6/Component_Function_3/NAND4_in[1] ), .A2(n774), 
        .A3(\SB3_6/Component_Function_3/NAND4_in[0] ), .A4(
        \SB3_6/Component_Function_3/NAND4_in[2] ), .ZN(\SB3_6/buf_output[3] )
         );
  NAND3_X1 U9085 ( .A1(\SB4_1/i0_0 ), .A2(\SB4_1/i1_7 ), .A3(\SB4_1/i3[0] ), 
        .ZN(n3469) );
  NAND4_X2 U9086 ( .A1(n2449), .A2(\SB2_1_1/Component_Function_5/NAND4_in[1] ), 
        .A3(\SB2_1_1/Component_Function_5/NAND4_in[0] ), .A4(n5417), .ZN(
        \SB2_1_1/buf_output[5] ) );
  NAND3_X2 U9087 ( .A1(\SB2_1_1/i0_4 ), .A2(\SB2_1_1/i0[6] ), .A3(
        \SB2_1_1/i0[9] ), .ZN(n5417) );
  INV_X2 U9090 ( .I(\SB1_2_18/buf_output[3] ), .ZN(\SB2_2_16/i0[8] ) );
  NAND4_X2 U9091 ( .A1(\SB1_2_18/Component_Function_3/NAND4_in[1] ), .A2(n3828), .A3(\SB1_2_18/Component_Function_3/NAND4_in[2] ), .A4(n2318), .ZN(
        \SB1_2_18/buf_output[3] ) );
  BUF_X4 U9096 ( .I(\SB3_29/buf_output[5] ), .Z(\SB4_29/i0_3 ) );
  INV_X1 U9097 ( .I(\SB1_3_21/buf_output[0] ), .ZN(\SB2_3_16/i3[0] ) );
  NAND4_X2 U9098 ( .A1(\SB1_3_21/Component_Function_0/NAND4_in[3] ), .A2(
        \SB1_3_21/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_3_21/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_3_21/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_3_21/buf_output[0] ) );
  XOR2_X1 U9100 ( .A1(n5418), .A2(n80), .Z(Ciphertext[15]) );
  NAND4_X2 U9101 ( .A1(n3161), .A2(n6372), .A3(
        \SB4_29/Component_Function_3/NAND4_in[3] ), .A4(n3504), .ZN(n5418) );
  NAND4_X2 U9102 ( .A1(\SB1_2_28/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_2_28/Component_Function_2/NAND4_in[2] ), .A3(
        \SB1_2_28/Component_Function_2/NAND4_in[0] ), .A4(n5419), .ZN(
        \SB1_2_28/buf_output[2] ) );
  XOR2_X1 U9104 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[133] ), .A2(\RI5[2][109] ), 
        .Z(n838) );
  XOR2_X1 U9105 ( .A1(n5420), .A2(\MC_ARK_ARC_1_3/temp6[148] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[148] ) );
  XOR2_X1 U9106 ( .A1(\MC_ARK_ARC_1_3/temp1[148] ), .A2(
        \MC_ARK_ARC_1_3/temp2[148] ), .Z(n5420) );
  INV_X2 U9107 ( .I(\SB1_2_7/buf_output[2] ), .ZN(\SB2_2_4/i1[9] ) );
  XOR2_X1 U9110 ( .A1(\MC_ARK_ARC_1_2/temp2[74] ), .A2(n5421), .Z(
        \MC_ARK_ARC_1_2/temp5[74] ) );
  XOR2_X1 U9112 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[68] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[74] ), .Z(n5421) );
  INV_X2 U9113 ( .I(\SB1_3_0/buf_output[3] ), .ZN(\SB2_3_30/i0[8] ) );
  NAND4_X2 U9115 ( .A1(\SB1_3_0/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_3_0/Component_Function_3/NAND4_in[0] ), .A3(n5742), .A4(
        \SB1_3_0/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_3_0/buf_output[3] ) );
  NAND4_X2 U9127 ( .A1(\SB4_16/Component_Function_0/NAND4_in[1] ), .A2(
        \SB4_16/Component_Function_0/NAND4_in[2] ), .A3(n3838), .A4(n5422), 
        .ZN(n3779) );
  NAND2_X1 U9128 ( .A1(\SB4_16/i0[10] ), .A2(\SB4_16/i0[9] ), .ZN(n5422) );
  NAND3_X2 U9130 ( .A1(\SB2_3_22/i0[10] ), .A2(\SB2_3_22/i0_3 ), .A3(
        \SB2_3_22/i0[6] ), .ZN(n5423) );
  NAND3_X2 U9131 ( .A1(\SB2_2_7/i0_3 ), .A2(\SB2_2_7/i0[10] ), .A3(
        \SB2_2_7/i0[9] ), .ZN(n5551) );
  INV_X2 U9132 ( .I(\SB1_2_3/buf_output[3] ), .ZN(\SB2_2_1/i0[8] ) );
  NAND4_X2 U9133 ( .A1(n880), .A2(\SB1_2_3/Component_Function_3/NAND4_in[0] ), 
        .A3(\SB1_2_3/Component_Function_3/NAND4_in[1] ), .A4(
        \SB1_2_3/Component_Function_3/NAND4_in[2] ), .ZN(
        \SB1_2_3/buf_output[3] ) );
  XOR2_X1 U9135 ( .A1(n5425), .A2(n156), .Z(Ciphertext[148]) );
  NAND4_X2 U9136 ( .A1(\SB4_7/Component_Function_4/NAND4_in[2] ), .A2(n6333), 
        .A3(n4329), .A4(n4567), .ZN(n5425) );
  NAND3_X2 U9137 ( .A1(\SB1_3_4/i0[6] ), .A2(\SB1_3_4/i1[9] ), .A3(
        \SB1_3_4/i0_3 ), .ZN(n5647) );
  NAND3_X2 U9138 ( .A1(\SB1_3_8/i0[6] ), .A2(\SB1_3_8/i0[7] ), .A3(
        \SB1_3_8/i0[8] ), .ZN(\SB1_3_8/Component_Function_0/NAND4_in[1] ) );
  NAND4_X2 U9140 ( .A1(n2287), .A2(n4318), .A3(n1097), .A4(
        \SB2_0_9/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_0_9/buf_output[5] ) );
  NAND3_X1 U9141 ( .A1(n5880), .A2(\SB2_2_8/i0[6] ), .A3(\SB2_2_8/i1_5 ), .ZN(
        \SB2_2_8/Component_Function_1/NAND4_in[2] ) );
  XOR2_X1 U9148 ( .A1(n5427), .A2(n5426), .Z(\MC_ARK_ARC_1_2/temp5[143] ) );
  XOR2_X1 U9149 ( .A1(\RI5[2][89] ), .A2(\RI5[2][113] ), .Z(n5427) );
  NAND4_X2 U9151 ( .A1(\SB2_0_17/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_17/Component_Function_5/NAND4_in[0] ), .A3(n2618), .A4(n5428), 
        .ZN(\SB2_0_17/buf_output[5] ) );
  NAND3_X2 U9153 ( .A1(\SB2_0_17/i0[10] ), .A2(\SB2_0_17/i0_0 ), .A3(
        \SB2_0_17/i0[6] ), .ZN(n5428) );
  XOR2_X1 U9154 ( .A1(n5430), .A2(n5429), .Z(\MC_ARK_ARC_1_1/temp6[107] ) );
  XOR2_X1 U9155 ( .A1(\RI5[1][17] ), .A2(n42), .Z(n5429) );
  XOR2_X1 U9159 ( .A1(\RI5[1][173] ), .A2(\RI5[1][143] ), .Z(n5430) );
  XOR2_X1 U9162 ( .A1(n5431), .A2(n132), .Z(Ciphertext[17]) );
  NAND3_X2 U9164 ( .A1(\SB2_1_16/i0_4 ), .A2(\SB2_1_16/i0_3 ), .A3(
        \SB2_1_16/i1[9] ), .ZN(n2429) );
  NAND3_X2 U9165 ( .A1(\SB2_2_14/i3[0] ), .A2(\SB2_2_14/i1_5 ), .A3(
        \SB2_2_14/i0[8] ), .ZN(\SB2_2_14/Component_Function_3/NAND4_in[3] ) );
  OAI21_X2 U9167 ( .A1(n2904), .A2(\SB2_3_3/i1[9] ), .B(\SB2_3_3/i0_3 ), .ZN(
        n4304) );
  NAND3_X2 U9170 ( .A1(\SB3_30/i0[10] ), .A2(\SB3_30/i0_0 ), .A3(
        \SB3_30/i0[6] ), .ZN(\SB3_30/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U9173 ( .A1(\MC_ARK_ARC_1_2/temp5[144] ), .A2(n5432), .Z(
        \MC_ARK_ARC_1_2/buf_output[144] ) );
  XOR2_X1 U9177 ( .A1(n4063), .A2(\MC_ARK_ARC_1_2/temp4[144] ), .Z(n5432) );
  NOR2_X2 U9178 ( .A1(n2027), .A2(n2025), .ZN(n6073) );
  NAND4_X2 U9181 ( .A1(n4497), .A2(\SB2_2_26/Component_Function_3/NAND4_in[1] ), .A3(\SB2_2_26/Component_Function_3/NAND4_in[3] ), .A4(n5434), .ZN(
        \SB2_2_26/buf_output[3] ) );
  NAND3_X2 U9190 ( .A1(\SB2_2_26/i0[6] ), .A2(\SB2_2_26/i0_3 ), .A3(
        \SB2_2_26/i1[9] ), .ZN(n5434) );
  BUF_X4 U9193 ( .I(\MC_ARK_ARC_1_1/buf_output[5] ), .Z(\SB1_2_31/i0_3 ) );
  NAND3_X2 U9194 ( .A1(\SB4_29/i0[10] ), .A2(\SB4_29/i0[6] ), .A3(
        \SB4_29/i0_3 ), .ZN(n6140) );
  NAND3_X2 U9198 ( .A1(\SB3_12/i0_3 ), .A2(\SB3_12/i0_0 ), .A3(\SB3_12/i0_4 ), 
        .ZN(n6512) );
  NAND4_X2 U9200 ( .A1(\SB3_5/Component_Function_5/NAND4_in[3] ), .A2(n2158), 
        .A3(n2135), .A4(n5435), .ZN(\SB3_5/buf_output[5] ) );
  NAND3_X2 U9201 ( .A1(\SB3_5/i0[6] ), .A2(\SB3_5/i0_0 ), .A3(\SB3_5/i0[10] ), 
        .ZN(n5435) );
  NAND4_X2 U9210 ( .A1(\SB1_2_9/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_2_9/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_2_9/Component_Function_5/NAND4_in[0] ), .A4(n3886), .ZN(
        \SB1_2_9/buf_output[5] ) );
  BUF_X2 U9211 ( .I(\SB3_10/buf_output[2] ), .Z(\SB4_7/i0_0 ) );
  XOR2_X1 U9212 ( .A1(\MC_ARK_ARC_1_2/temp1[57] ), .A2(n5436), .Z(
        \MC_ARK_ARC_1_2/temp5[57] ) );
  XOR2_X1 U9215 ( .A1(\RI5[2][3] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[27] ), 
        .Z(n5436) );
  NAND3_X2 U9216 ( .A1(\SB3_0/i0[10] ), .A2(\SB3_0/i0_0 ), .A3(\SB3_0/i0[6] ), 
        .ZN(\SB3_0/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U9217 ( .A1(\MC_ARK_ARC_1_2/temp1[187] ), .A2(n5437), .Z(
        \MC_ARK_ARC_1_2/temp5[187] ) );
  XOR2_X1 U9218 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[133] ), .A2(\RI5[2][157] ), 
        .Z(n5437) );
  INV_X2 U9222 ( .I(\MC_ARK_ARC_1_1/buf_output[5] ), .ZN(\SB1_2_31/i1_5 ) );
  NAND3_X2 U9226 ( .A1(\SB2_3_0/i0_3 ), .A2(\SB2_3_0/i0[9] ), .A3(
        \SB2_3_0/i0[10] ), .ZN(n6053) );
  NAND3_X2 U9233 ( .A1(\SB2_3_12/i3[0] ), .A2(n3651), .A3(\SB2_3_12/i1_5 ), 
        .ZN(\SB2_3_12/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U9234 ( .A1(\RI5[3][57] ), .A2(\RI5[3][21] ), .Z(
        \MC_ARK_ARC_1_3/temp3[147] ) );
  XOR2_X1 U9238 ( .A1(\MC_ARK_ARC_1_2/temp1[27] ), .A2(
        \MC_ARK_ARC_1_2/temp2[27] ), .Z(\MC_ARK_ARC_1_2/temp5[27] ) );
  NAND4_X2 U9239 ( .A1(n4155), .A2(\SB2_1_1/Component_Function_3/NAND4_in[3] ), 
        .A3(\SB2_1_1/Component_Function_3/NAND4_in[1] ), .A4(n5439), .ZN(
        \SB2_1_1/buf_output[3] ) );
  NAND3_X2 U9246 ( .A1(\SB2_1_1/i0_3 ), .A2(\SB2_1_1/i0[6] ), .A3(
        \SB2_1_1/i1[9] ), .ZN(n5439) );
  NAND4_X2 U9248 ( .A1(\SB1_2_25/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_25/Component_Function_0/NAND4_in[0] ), .A3(
        \SB1_2_25/Component_Function_0/NAND4_in[1] ), .A4(n5440), .ZN(
        \SB1_2_25/buf_output[0] ) );
  NAND3_X1 U9249 ( .A1(\SB1_2_25/i0[7] ), .A2(\SB1_2_25/i0_0 ), .A3(
        \SB1_2_25/i0_3 ), .ZN(n5440) );
  NAND4_X2 U9254 ( .A1(\SB1_3_28/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_28/Component_Function_2/NAND4_in[1] ), .A3(n5542), .A4(n5441), 
        .ZN(\SB1_3_28/buf_output[2] ) );
  NAND3_X2 U9256 ( .A1(\SB2_1_30/i0_3 ), .A2(\SB2_1_30/i0_4 ), .A3(
        \SB2_1_30/i1[9] ), .ZN(\SB2_1_30/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U9258 ( .A1(\SB2_3_5/Component_Function_5/NAND4_in[1] ), .A2(n4372), 
        .A3(\SB2_3_5/Component_Function_5/NAND4_in[0] ), .A4(n5442), .ZN(
        \SB2_3_5/buf_output[5] ) );
  NAND3_X2 U9265 ( .A1(\SB2_3_5/i0[6] ), .A2(\SB2_3_5/i0_4 ), .A3(
        \SB2_3_5/i0[9] ), .ZN(n5442) );
  NAND3_X1 U9266 ( .A1(\SB2_2_9/i1_7 ), .A2(\SB1_2_9/buf_output[5] ), .A3(
        \SB2_2_9/i0[8] ), .ZN(\SB2_2_9/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U9269 ( .A1(\SB4_15/i0[10] ), .A2(\SB4_15/i0_3 ), .A3(
        \SB4_15/i0[9] ), .ZN(n5443) );
  NAND3_X2 U9273 ( .A1(\SB3_12/i0_3 ), .A2(\SB3_12/i0[8] ), .A3(\SB3_12/i0[9] ), .ZN(\SB3_12/Component_Function_2/NAND4_in[2] ) );
  BUF_X2 U9276 ( .I(\SB3_15/buf_output[0] ), .Z(\SB4_10/i0[9] ) );
  NAND3_X2 U9279 ( .A1(\SB1_3_8/i0_3 ), .A2(\SB1_3_8/i1[9] ), .A3(
        \SB1_3_8/i0[6] ), .ZN(\SB1_3_8/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U9281 ( .A1(\MC_ARK_ARC_1_3/temp5[114] ), .A2(n5444), .Z(
        \MC_ARK_ARC_1_3/buf_output[114] ) );
  XOR2_X1 U9283 ( .A1(\MC_ARK_ARC_1_3/temp3[114] ), .A2(
        \MC_ARK_ARC_1_3/temp4[114] ), .Z(n5444) );
  NAND3_X1 U9285 ( .A1(\SB3_1/i0[9] ), .A2(\SB3_1/i1_5 ), .A3(\SB3_1/i0[6] ), 
        .ZN(\SB3_1/Component_Function_1/NAND4_in[2] ) );
  XOR2_X1 U9286 ( .A1(n1232), .A2(n5445), .Z(n5645) );
  XOR2_X1 U9287 ( .A1(\RI5[2][101] ), .A2(\RI5[2][107] ), .Z(n5445) );
  NOR2_X2 U9290 ( .A1(n5447), .A2(n5446), .ZN(n6194) );
  NAND3_X2 U9291 ( .A1(\SB1_1_7/i0[10] ), .A2(\SB1_1_7/i0_3 ), .A3(
        \SB1_1_7/i0[6] ), .ZN(\SB1_1_7/Component_Function_2/NAND4_in[1] ) );
  XOR2_X1 U9299 ( .A1(n817), .A2(n5448), .Z(\MC_ARK_ARC_1_2/buf_output[83] )
         );
  XOR2_X1 U9301 ( .A1(n3129), .A2(\MC_ARK_ARC_1_2/temp4[83] ), .Z(n5448) );
  XOR2_X1 U9303 ( .A1(n5449), .A2(n74), .Z(Ciphertext[111]) );
  NAND4_X2 U9304 ( .A1(n2228), .A2(\SB4_13/Component_Function_3/NAND4_in[3] ), 
        .A3(\SB4_13/Component_Function_3/NAND4_in[0] ), .A4(n6394), .ZN(n5449)
         );
  XOR2_X1 U9306 ( .A1(n5450), .A2(\MC_ARK_ARC_1_0/temp4[170] ), .Z(
        \MC_ARK_ARC_1_0/temp6[170] ) );
  XOR2_X1 U9309 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[44] ), .A2(\RI5[0][80] ), 
        .Z(n5450) );
  XOR2_X1 U9310 ( .A1(\RI5[1][137] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[35] ), 
        .Z(n5451) );
  NAND3_X1 U9312 ( .A1(\SB1_1_22/i1[9] ), .A2(\SB1_1_22/i0_4 ), .A3(
        \RI1[1][59] ), .ZN(n5554) );
  XOR2_X1 U9315 ( .A1(\MC_ARK_ARC_1_1/temp6[45] ), .A2(n5453), .Z(
        \MC_ARK_ARC_1_1/buf_output[45] ) );
  NAND3_X1 U9316 ( .A1(\SB4_0/i0[6] ), .A2(\SB4_0/i0_3 ), .A3(n1386), .ZN(
        n5454) );
  NAND3_X1 U9320 ( .A1(\SB1_1_1/i0_3 ), .A2(\SB1_1_1/i0_0 ), .A3(
        \SB1_1_1/i0[7] ), .ZN(n2100) );
  NAND4_X2 U9321 ( .A1(\SB1_2_1/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_2_1/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_2_1/Component_Function_4/NAND4_in[2] ), .A4(n5455), .ZN(
        \SB1_2_1/buf_output[4] ) );
  NAND3_X1 U9324 ( .A1(\SB1_2_1/i0_4 ), .A2(\SB1_2_1/i1[9] ), .A3(
        \SB1_2_1/i1_5 ), .ZN(n5455) );
  NAND4_X2 U9327 ( .A1(\SB1_1_4/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_4/Component_Function_5/NAND4_in[2] ), .A3(n2993), .A4(
        \SB1_1_4/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_4/buf_output[5] ) );
  INV_X2 U9329 ( .I(\SB1_1_23/buf_output[2] ), .ZN(\SB2_1_20/i1[9] ) );
  XOR2_X1 U9330 ( .A1(n5829), .A2(n5456), .Z(n5875) );
  XOR2_X1 U9332 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[86] ), .A2(\RI5[0][152] ), 
        .Z(n5456) );
  NAND2_X1 U9333 ( .A1(\SB4_31/i0[9] ), .A2(\SB4_31/i0[10] ), .ZN(
        \SB4_31/Component_Function_0/NAND4_in[0] ) );
  XOR2_X1 U9341 ( .A1(\MC_ARK_ARC_1_1/temp1[39] ), .A2(n5457), .Z(n864) );
  XOR2_X1 U9342 ( .A1(\RI5[1][177] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[9] ), 
        .Z(n5457) );
  BUF_X4 U9344 ( .I(\SB2_0_14/buf_output[2] ), .Z(\RI5[0][122] ) );
  NAND3_X2 U9346 ( .A1(\SB1_2_4/i0[6] ), .A2(\SB1_2_4/i0_0 ), .A3(
        \SB1_2_4/i0[10] ), .ZN(\SB1_2_4/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U9347 ( .A1(\SB4_31/i0_4 ), .A2(\SB4_31/i0_3 ), .A3(\SB4_31/i0[10] ), .ZN(\SB4_31/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U9349 ( .A1(\SB1_3_9/i0_3 ), .A2(\SB1_3_9/i1[9] ), .A3(
        \MC_ARK_ARC_1_2/buf_output[136] ), .ZN(
        \SB1_3_9/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U9351 ( .A1(\SB2_1_28/Component_Function_2/NAND4_in[0] ), .A2(n6429), .A3(\SB2_1_28/Component_Function_2/NAND4_in[1] ), .A4(n5458), .ZN(
        \SB2_1_28/buf_output[2] ) );
  NAND3_X2 U9352 ( .A1(\SB2_1_28/i0_4 ), .A2(\SB2_1_28/i0_0 ), .A3(
        \SB2_1_28/i1_5 ), .ZN(n5458) );
  NAND3_X1 U9355 ( .A1(\SB4_31/i0_3 ), .A2(\SB4_31/i0[6] ), .A3(\SB4_31/i1[9] ), .ZN(n1472) );
  NAND4_X2 U9356 ( .A1(\SB4_4/Component_Function_3/NAND4_in[3] ), .A2(n5570), 
        .A3(\SB4_4/Component_Function_3/NAND4_in[2] ), .A4(n5459), .ZN(n6243)
         );
  NAND3_X2 U9357 ( .A1(\SB2_0_24/i0_3 ), .A2(\SB2_0_24/i0[10] ), .A3(
        \RI3[0][43] ), .ZN(n1789) );
  XOR2_X1 U9358 ( .A1(n6027), .A2(n5460), .Z(\MC_ARK_ARC_1_2/buf_output[155] )
         );
  NAND3_X2 U9359 ( .A1(\SB2_1_16/i0_0 ), .A2(\SB2_1_16/i0_4 ), .A3(
        \SB2_1_16/i1_5 ), .ZN(n5461) );
  NAND3_X2 U9360 ( .A1(\SB2_1_11/i0_3 ), .A2(\SB2_1_11/i0_0 ), .A3(
        \SB1_1_12/buf_output[4] ), .ZN(
        \SB2_1_11/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U9361 ( .A1(\RI5[2][62] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[86] ), 
        .Z(n632) );
  XOR2_X1 U9362 ( .A1(\MC_ARK_ARC_1_0/temp5[155] ), .A2(
        \MC_ARK_ARC_1_0/temp6[155] ), .Z(\MC_ARK_ARC_1_0/buf_output[155] ) );
  XOR2_X1 U9364 ( .A1(n2069), .A2(\MC_ARK_ARC_1_3/temp6[2] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[2] ) );
  XOR2_X1 U9370 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[170] ), .A2(\RI5[1][146] ), 
        .Z(n2739) );
  NAND3_X2 U9373 ( .A1(\SB4_31/i0[10] ), .A2(\SB4_31/i0[9] ), .A3(
        \SB4_31/i0_3 ), .ZN(n2531) );
  XOR2_X1 U9374 ( .A1(\RI5[3][113] ), .A2(\RI5[3][77] ), .Z(
        \MC_ARK_ARC_1_3/temp3[11] ) );
  NAND3_X2 U9375 ( .A1(\SB4_29/i0_0 ), .A2(n1793), .A3(\SB4_29/i0_3 ), .ZN(
        n3504) );
  BUF_X4 U9376 ( .I(\MC_ARK_ARC_1_0/buf_output[134] ), .Z(\SB1_1_9/i0_0 ) );
  XOR2_X1 U9386 ( .A1(\MC_ARK_ARC_1_0/temp6[99] ), .A2(n5463), .Z(
        \MC_ARK_ARC_1_0/buf_output[99] ) );
  XOR2_X1 U9387 ( .A1(\MC_ARK_ARC_1_0/temp1[99] ), .A2(n2022), .Z(n5463) );
  BUF_X4 U9389 ( .I(\MC_ARK_ARC_1_1/buf_output[112] ), .Z(\SB1_2_13/i0_4 ) );
  XOR2_X1 U9391 ( .A1(n5627), .A2(n5464), .Z(n5583) );
  XOR2_X1 U9392 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[92] ), .A2(\RI5[2][98] ), 
        .Z(n5464) );
  BUF_X4 U9394 ( .I(\SB2_2_15/buf_output[2] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[116] ) );
  XOR2_X1 U9396 ( .A1(n2309), .A2(n5466), .Z(\MC_ARK_ARC_1_2/buf_output[95] )
         );
  XOR2_X1 U9397 ( .A1(n6038), .A2(\MC_ARK_ARC_1_2/temp4[95] ), .Z(n5466) );
  XOR2_X1 U9398 ( .A1(n3905), .A2(n5467), .Z(n5479) );
  XOR2_X1 U9408 ( .A1(\RI5[1][50] ), .A2(\RI5[1][14] ), .Z(
        \MC_ARK_ARC_1_1/temp3[140] ) );
  NAND4_X2 U9409 ( .A1(\SB2_3_8/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_8/Component_Function_4/NAND4_in[3] ), .A3(n4282), .A4(n5468), 
        .ZN(\SB2_3_8/buf_output[4] ) );
  XOR2_X1 U9412 ( .A1(\MC_ARK_ARC_1_1/temp2[116] ), .A2(n5470), .Z(n5843) );
  XOR2_X1 U9414 ( .A1(\RI5[1][116] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[110] ), 
        .Z(n5470) );
  NAND4_X2 U9420 ( .A1(\SB2_2_6/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_2_6/Component_Function_4/NAND4_in[3] ), .A3(n4432), .A4(n5472), 
        .ZN(\SB2_2_6/buf_output[4] ) );
  NAND3_X2 U9421 ( .A1(\SB2_0_15/i0[10] ), .A2(\SB2_0_15/i0_0 ), .A3(
        \SB2_0_15/i0[6] ), .ZN(n5473) );
  NAND4_X2 U9422 ( .A1(\SB1_2_19/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_2_19/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_19/Component_Function_1/NAND4_in[0] ), .A4(n5474), .ZN(
        \SB1_2_19/buf_output[1] ) );
  NAND3_X2 U9425 ( .A1(\SB1_2_19/i0_4 ), .A2(\SB1_2_19/i0[8] ), .A3(
        \SB1_2_19/i1_7 ), .ZN(n5474) );
  XOR2_X1 U9426 ( .A1(n5475), .A2(\MC_ARK_ARC_1_2/temp6[118] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[118] ) );
  XOR2_X1 U9429 ( .A1(\MC_ARK_ARC_1_2/temp2[118] ), .A2(
        \MC_ARK_ARC_1_2/temp1[118] ), .Z(n5475) );
  NAND3_X1 U9432 ( .A1(\SB2_0_27/i0_3 ), .A2(n2237), .A3(\SB2_0_27/i0_0 ), 
        .ZN(\SB2_0_27/Component_Function_0/NAND4_in[3] ) );
  NAND3_X2 U9433 ( .A1(\SB1_0_17/i0_3 ), .A2(\SB1_0_17/i0_0 ), .A3(n2899), 
        .ZN(n4685) );
  NAND3_X1 U9436 ( .A1(\SB3_23/i0_3 ), .A2(\SB3_23/i0[9] ), .A3(
        \SB3_23/i0[10] ), .ZN(\SB3_23/Component_Function_4/NAND4_in[2] ) );
  INV_X1 U9438 ( .I(\SB1_1_26/buf_output[5] ), .ZN(\SB2_1_26/i1_5 ) );
  NAND4_X2 U9442 ( .A1(\SB1_1_26/Component_Function_5/NAND4_in[1] ), .A2(n1940), .A3(\SB1_1_26/Component_Function_5/NAND4_in[3] ), .A4(
        \SB1_1_26/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_26/buf_output[5] ) );
  BUF_X4 U9444 ( .I(\MC_ARK_ARC_1_0/buf_output[144] ), .Z(\SB1_1_7/i0[9] ) );
  NAND3_X2 U9445 ( .A1(\SB2_1_6/i0_3 ), .A2(\SB2_1_6/i0[8] ), .A3(
        \SB2_1_6/i0[9] ), .ZN(n5476) );
  XOR2_X1 U9446 ( .A1(n5477), .A2(n5478), .Z(\MC_ARK_ARC_1_2/temp5[158] ) );
  XOR2_X1 U9447 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[158] ), .A2(\RI5[2][104] ), 
        .Z(n5477) );
  XOR2_X1 U9448 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[128] ), .A2(\RI5[2][152] ), 
        .Z(n5478) );
  NAND3_X2 U9449 ( .A1(\SB1_1_1/i0_3 ), .A2(\SB1_1_1/i1[9] ), .A3(
        \SB1_1_1/i0_4 ), .ZN(n6232) );
  XOR2_X1 U9452 ( .A1(n3559), .A2(n5479), .Z(\MC_ARK_ARC_1_0/buf_output[93] )
         );
  BUF_X4 U9453 ( .I(\RI1[4][179] ), .Z(\SB3_2/i0_3 ) );
  XOR2_X1 U9456 ( .A1(n5480), .A2(n92), .Z(Ciphertext[178]) );
  NAND4_X2 U9460 ( .A1(\SB4_2/Component_Function_4/NAND4_in[1] ), .A2(
        \SB4_2/Component_Function_4/NAND4_in[0] ), .A3(n4592), .A4(n5593), 
        .ZN(n5480) );
  NAND3_X2 U9461 ( .A1(\SB1_3_5/i0[6] ), .A2(\SB1_3_5/i0_0 ), .A3(
        \SB1_3_5/i0[10] ), .ZN(n5481) );
  NAND4_X2 U9462 ( .A1(\SB1_2_20/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_2_20/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_2_20/Component_Function_3/NAND4_in[3] ), .A4(n5482), .ZN(
        \SB1_2_20/buf_output[3] ) );
  NAND3_X2 U9466 ( .A1(\SB1_2_18/i0_0 ), .A2(\SB1_2_18/i0[6] ), .A3(
        \SB1_2_18/i0[10] ), .ZN(\SB1_2_18/Component_Function_5/NAND4_in[1] )
         );
  NAND4_X2 U9467 ( .A1(\SB2_3_2/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_3_2/Component_Function_4/NAND4_in[0] ), .A3(n679), .A4(n5483), 
        .ZN(\SB2_3_2/buf_output[4] ) );
  NAND4_X2 U9468 ( .A1(\SB1_1_6/Component_Function_3/NAND4_in[1] ), .A2(n4293), 
        .A3(n2700), .A4(n5484), .ZN(\SB1_1_6/buf_output[3] ) );
  NAND3_X1 U9469 ( .A1(\SB1_1_1/i0_3 ), .A2(\SB1_1_1/i0[6] ), .A3(
        \SB1_1_1/i1[9] ), .ZN(\SB1_1_1/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U9473 ( .A1(\SB2_1_31/i0[10] ), .A2(\SB2_1_31/i0_0 ), .A3(
        \SB2_1_31/i0[6] ), .ZN(\SB2_1_31/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U9474 ( .A1(\SB1_3_16/i0_0 ), .A2(\SB1_3_16/i0_4 ), .A3(
        \SB1_3_16/i1_5 ), .ZN(n5770) );
  NAND3_X2 U9475 ( .A1(\SB2_2_4/i0_3 ), .A2(\SB2_2_4/i0_0 ), .A3(
        \SB2_2_4/i0_4 ), .ZN(\SB2_2_4/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U9476 ( .A1(\SB1_0_8/i0_3 ), .A2(\SB1_0_8/i0_4 ), .A3(
        \SB1_0_8/i1[9] ), .ZN(n2539) );
  BUF_X4 U9477 ( .I(\SB1_2_25/buf_output[2] ), .Z(\SB2_2_22/i0_0 ) );
  BUF_X4 U9479 ( .I(\SB3_22/buf_output[5] ), .Z(\SB4_22/i0_3 ) );
  NAND3_X2 U9480 ( .A1(\SB1_3_8/i0_3 ), .A2(\SB1_3_8/i0[9] ), .A3(
        \SB1_3_8/i0[8] ), .ZN(\SB1_3_8/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U9482 ( .A1(\SB4_16/i0[10] ), .A2(\SB4_16/i0_3 ), .A3(
        \SB4_16/i0[6] ), .ZN(n4340) );
  CLKBUF_X4 U9483 ( .I(\SB3_14/buf_output[5] ), .Z(\SB4_14/i0_3 ) );
  CLKBUF_X4 U9485 ( .I(\SB3_6/buf_output[5] ), .Z(\SB4_6/i0_3 ) );
  NAND3_X1 U9488 ( .A1(\SB2_3_30/i1_5 ), .A2(\SB2_3_30/i0[6] ), .A3(
        \SB2_3_30/i0[9] ), .ZN(\SB2_3_30/Component_Function_1/NAND4_in[2] ) );
  CLKBUF_X4 U9491 ( .I(\SB3_24/buf_output[5] ), .Z(\SB4_24/i0_3 ) );
  NAND3_X1 U9492 ( .A1(\SB2_3_1/i0_0 ), .A2(\SB2_3_1/i1_5 ), .A3(
        \SB2_3_1/i0_4 ), .ZN(\SB2_3_1/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U9494 ( .A1(\SB4_8/i0[6] ), .A2(\SB4_8/i0_3 ), .A3(\SB4_8/i0[10] ), 
        .ZN(n6212) );
  CLKBUF_X4 U9497 ( .I(\SB3_26/buf_output[4] ), .Z(\SB4_25/i0_4 ) );
  CLKBUF_X4 U9498 ( .I(\RI3[4][23] ), .Z(\SB4_28/i0_3 ) );
  CLKBUF_X4 U9499 ( .I(\SB2_2_7/buf_output[3] ), .Z(\RI5[2][159] ) );
  NAND3_X1 U9500 ( .A1(\SB2_3_18/i0_4 ), .A2(\SB2_3_18/i1[9] ), .A3(
        \SB2_3_18/i1_5 ), .ZN(n4694) );
  NAND3_X1 U9501 ( .A1(\SB2_3_18/i1[9] ), .A2(\SB2_3_18/i0_3 ), .A3(
        \SB2_3_18/i0[6] ), .ZN(\SB2_3_18/Component_Function_3/NAND4_in[0] ) );
  CLKBUF_X4 U9502 ( .I(\SB1_3_21/buf_output[5] ), .Z(\SB2_3_21/i0_3 ) );
  CLKBUF_X4 U9504 ( .I(\SB3_7/buf_output[4] ), .Z(\SB4_6/i0_4 ) );
  CLKBUF_X4 U9505 ( .I(\SB2_3_13/buf_output[1] ), .Z(\RI5[3][133] ) );
  NAND3_X1 U9508 ( .A1(\SB4_6/i0_3 ), .A2(\SB4_6/i0[9] ), .A3(n579), .ZN(n5724) );
  NAND3_X1 U9512 ( .A1(\SB4_6/i0_3 ), .A2(\SB4_6/i0[10] ), .A3(\SB4_6/i0[9] ), 
        .ZN(\SB4_6/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U9513 ( .A1(\SB3_3/i0[7] ), .A2(\SB3_3/i0_3 ), .A3(\SB3_3/i0_0 ), 
        .ZN(\SB3_3/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 U9514 ( .A1(\SB3_3/i0_0 ), .A2(\SB3_3/i3[0] ), .ZN(
        \SB3_3/Component_Function_5/NAND4_in[0] ) );
  CLKBUF_X4 U9515 ( .I(\SB3_26/buf_output[5] ), .Z(\SB4_26/i0_3 ) );
  NAND2_X1 U9516 ( .A1(\SB4_13/i0_3 ), .A2(\SB4_13/i1[9] ), .ZN(n3231) );
  INV_X1 U9517 ( .I(n5505), .ZN(\SB4_15/i0[8] ) );
  BUF_X4 U9518 ( .I(\SB2_3_6/buf_output[0] ), .Z(\RI5[3][180] ) );
  CLKBUF_X4 U9519 ( .I(\SB3_25/buf_output[4] ), .Z(\SB4_24/i0_4 ) );
  CLKBUF_X4 U9520 ( .I(\SB2_2_9/buf_output[3] ), .Z(\RI5[2][147] ) );
  BUF_X2 U9525 ( .I(\SB3_24/buf_output[4] ), .Z(\SB4_23/i0_4 ) );
  NAND3_X1 U9526 ( .A1(\SB4_6/i0_4 ), .A2(\SB4_6/i0[10] ), .A3(\SB4_6/i0_3 ), 
        .ZN(n3461) );
  NAND2_X1 U9527 ( .A1(\SB1_3_17/i0_3 ), .A2(\SB1_3_17/i1[9] ), .ZN(n6135) );
  NAND3_X1 U9528 ( .A1(\SB1_3_17/i0_0 ), .A2(\SB1_3_17/i0_3 ), .A3(
        \SB1_3_17/i0[7] ), .ZN(n2520) );
  CLKBUF_X4 U9529 ( .I(\SB3_16/buf_output[0] ), .Z(\SB4_11/i0[9] ) );
  NAND2_X1 U9536 ( .A1(\SB4_6/i0[10] ), .A2(\SB4_6/i0[9] ), .ZN(
        \SB4_6/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U9538 ( .A1(\SB3_30/i0_3 ), .A2(\SB3_30/i0[10] ), .A3(
        \SB3_30/i0[6] ), .ZN(\SB3_30/Component_Function_2/NAND4_in[1] ) );
  CLKBUF_X4 U9539 ( .I(\RI1[4][89] ), .Z(\SB3_17/i0_3 ) );
  INV_X1 U9542 ( .I(\RI1[4][89] ), .ZN(\SB3_17/i1_5 ) );
  INV_X1 U9545 ( .I(\SB3_17/buf_output[1] ), .ZN(\SB4_13/i1_7 ) );
  NAND3_X1 U9548 ( .A1(\SB1_3_26/i0_0 ), .A2(\SB1_3_26/i0_3 ), .A3(
        \SB1_3_26/i0[7] ), .ZN(n2769) );
  NAND3_X1 U9549 ( .A1(\SB1_3_26/i0_4 ), .A2(\SB1_3_26/i0_3 ), .A3(
        \SB1_3_26/i0[10] ), .ZN(n6163) );
  NAND3_X1 U9551 ( .A1(\SB4_6/i0_3 ), .A2(\SB4_6/i0[10] ), .A3(\SB4_6/i0[6] ), 
        .ZN(n5844) );
  CLKBUF_X4 U9554 ( .I(\SB1_2_16/buf_output[0] ), .Z(\SB2_2_11/i0[9] ) );
  NAND3_X1 U9555 ( .A1(\SB3_11/i0[7] ), .A2(\SB3_11/i0_3 ), .A3(\SB3_11/i0_0 ), 
        .ZN(\SB3_11/Component_Function_0/NAND4_in[3] ) );
  CLKBUF_X4 U9556 ( .I(\MC_ARK_ARC_1_3/buf_output[122] ), .Z(\SB3_11/i0_0 ) );
  NAND3_X1 U9557 ( .A1(\SB4_16/i0_0 ), .A2(\SB4_16/i0[9] ), .A3(\SB4_16/i0[8] ), .ZN(\SB4_16/Component_Function_4/NAND4_in[0] ) );
  BUF_X2 U9559 ( .I(\SB1_3_8/buf_output[1] ), .Z(\SB2_3_4/i0[6] ) );
  INV_X1 U9560 ( .I(\SB1_3_8/buf_output[1] ), .ZN(\SB2_3_4/i1_7 ) );
  CLKBUF_X4 U9565 ( .I(\SB2_3_25/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[51] ) );
  CLKBUF_X4 U9567 ( .I(\SB3_12/buf_output[4] ), .Z(\SB4_11/i0_4 ) );
  NAND3_X1 U9574 ( .A1(\SB2_3_21/i0[10] ), .A2(\SB2_3_21/i0_3 ), .A3(
        \SB1_3_22/buf_output[4] ), .ZN(
        \SB2_3_21/Component_Function_0/NAND4_in[2] ) );
  NOR2_X1 U9577 ( .A1(\SB2_3_21/i0[10] ), .A2(\SB2_3_21/i1_7 ), .ZN(n971) );
  CLKBUF_X4 U9582 ( .I(\MC_ARK_ARC_1_2/buf_output[122] ), .Z(\SB1_3_11/i0_0 )
         );
  INV_X1 U9583 ( .I(\SB4_19/i0[7] ), .ZN(n5486) );
  CLKBUF_X12 U9584 ( .I(\SB3_20/buf_output[4] ), .Z(\SB4_19/i0_4 ) );
  NAND3_X1 U9585 ( .A1(\SB1_3_29/i1_5 ), .A2(\SB1_3_29/i0_4 ), .A3(
        \RI1[3][14] ), .ZN(n2307) );
  NAND3_X1 U9586 ( .A1(\SB1_3_28/i3[0] ), .A2(\SB1_3_28/i0[8] ), .A3(
        \SB1_3_28/i1_5 ), .ZN(\SB1_3_28/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U9587 ( .A1(\SB1_3_28/i0_4 ), .A2(\SB1_3_28/i1_7 ), .A3(
        \SB1_3_28/i0[8] ), .ZN(n1295) );
  CLKBUF_X4 U9590 ( .I(\MC_ARK_ARC_1_2/buf_output[18] ), .Z(\SB1_3_28/i0[9] )
         );
  NAND3_X1 U9591 ( .A1(\SB4_11/i0[10] ), .A2(\SB4_11/i0_4 ), .A3(\SB4_11/i0_3 ), .ZN(\SB4_11/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U9593 ( .A1(\SB4_11/i0_0 ), .A2(\SB4_11/i0_3 ), .A3(\SB4_11/i0[7] ), 
        .ZN(\SB4_11/Component_Function_0/NAND4_in[3] ) );
  CLKBUF_X4 U9594 ( .I(\SB3_11/buf_output[5] ), .Z(\SB4_11/i0_3 ) );
  BUF_X2 U9596 ( .I(\SB3_20/buf_output[2] ), .Z(\SB4_17/i0_0 ) );
  NAND3_X1 U9597 ( .A1(\SB4_17/i0_0 ), .A2(\SB4_17/i1_7 ), .A3(\SB4_17/i3[0] ), 
        .ZN(n1679) );
  NAND3_X1 U9598 ( .A1(\SB4_17/i0_4 ), .A2(\SB4_17/i0_0 ), .A3(\SB4_17/i0_3 ), 
        .ZN(n2098) );
  XOR2_X1 U9601 ( .A1(n3636), .A2(n3637), .Z(n5487) );
  NAND3_X1 U9605 ( .A1(\SB2_2_15/i0_4 ), .A2(\SB2_2_15/i1_7 ), .A3(
        \SB2_2_15/i0[8] ), .ZN(\SB2_2_15/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U9612 ( .A1(\SB2_2_15/i0_3 ), .A2(\SB2_2_15/i0[9] ), .A3(
        \SB2_2_15/i0[8] ), .ZN(n3615) );
  CLKBUF_X4 U9613 ( .I(\SB1_3_6/buf_output[4] ), .Z(\SB2_3_5/i0_4 ) );
  INV_X1 U9617 ( .I(\SB1_1_5/buf_output[1] ), .ZN(\SB2_1_1/i1_7 ) );
  BUF_X2 U9621 ( .I(\MC_ARK_ARC_1_1/buf_output[84] ), .Z(\SB1_2_17/i0[9] ) );
  INV_X1 U9622 ( .I(\MC_ARK_ARC_1_1/buf_output[84] ), .ZN(\SB1_2_17/i3[0] ) );
  NAND3_X1 U9624 ( .A1(\SB1_0_29/i0[6] ), .A2(\SB1_0_29/i0_3 ), .A3(
        \SB1_0_29/i1[9] ), .ZN(n4631) );
  NAND3_X1 U9626 ( .A1(\SB1_0_29/i0_4 ), .A2(\SB1_0_29/i0_3 ), .A3(
        \SB1_0_29/i1[9] ), .ZN(\SB1_0_29/Component_Function_5/NAND4_in[2] ) );
  BUF_X2 U9627 ( .I(n346), .Z(\SB1_0_29/i0_4 ) );
  NAND3_X1 U9629 ( .A1(\SB1_0_29/i0_4 ), .A2(\SB1_0_29/i0[9] ), .A3(
        \SB1_0_29/i0[6] ), .ZN(n1109) );
  NAND3_X1 U9630 ( .A1(\SB4_28/i0[9] ), .A2(\SB4_28/i0[10] ), .A3(
        \SB4_28/i0_3 ), .ZN(n5589) );
  NAND3_X1 U9634 ( .A1(\SB1_2_7/i0_3 ), .A2(\SB1_2_7/i0_4 ), .A3(
        \SB1_2_7/i1[9] ), .ZN(\SB1_2_7/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 U9638 ( .A1(\SB1_2_7/i0_3 ), .A2(\SB1_2_7/i1[9] ), .ZN(
        \SB1_2_7/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U9639 ( .A1(\SB1_2_7/i1[9] ), .A2(\SB1_2_7/i0_3 ), .A3(
        \MC_ARK_ARC_1_1/buf_output[145] ), .ZN(
        \SB1_2_7/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U9640 ( .A1(n1501), .A2(\MC_ARK_ARC_1_3/temp6[8] ), .Z(n5488) );
  CLKBUF_X4 U9641 ( .I(\MC_ARK_ARC_1_3/buf_output[7] ), .Z(\SB3_30/i0[6] ) );
  NAND3_X1 U9642 ( .A1(\SB4_12/i0_0 ), .A2(\SB4_12/i0_4 ), .A3(\SB4_12/i1_5 ), 
        .ZN(n4562) );
  BUF_X2 U9644 ( .I(\MC_ARK_ARC_1_3/buf_output[138] ), .Z(\SB3_8/i0[9] ) );
  NAND3_X1 U9645 ( .A1(\SB3_8/i0[9] ), .A2(\SB3_8/i0[6] ), .A3(\SB3_8/i0_4 ), 
        .ZN(\SB3_8/Component_Function_5/NAND4_in[3] ) );
  NAND3_X1 U9647 ( .A1(\SB3_8/i0_3 ), .A2(\SB3_8/i0[8] ), .A3(\SB3_8/i0[9] ), 
        .ZN(\SB3_8/Component_Function_2/NAND4_in[2] ) );
  CLKBUF_X4 U9649 ( .I(\SB1_2_5/buf_output[3] ), .Z(\SB2_2_3/i0[10] ) );
  NAND3_X1 U9661 ( .A1(\SB3_11/i0_3 ), .A2(\SB3_11/i0[6] ), .A3(\SB3_11/i1[9] ), .ZN(\SB3_11/Component_Function_3/NAND4_in[0] ) );
  CLKBUF_X4 U9662 ( .I(\MC_ARK_ARC_1_3/buf_output[120] ), .Z(\SB3_11/i0[9] )
         );
  CLKBUF_X4 U9663 ( .I(\MC_ARK_ARC_1_3/buf_output[25] ), .Z(\SB3_27/i0[6] ) );
  INV_X1 U9664 ( .I(\MC_ARK_ARC_1_3/buf_output[43] ), .ZN(\SB3_24/i1_7 ) );
  BUF_X2 U9666 ( .I(\MC_ARK_ARC_1_3/buf_output[43] ), .Z(\SB3_24/i0[6] ) );
  NAND4_X1 U9673 ( .A1(\SB1_3_31/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_31/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_3_31/Component_Function_2/NAND4_in[2] ), .A4(n4662), .ZN(n5489)
         );
  NAND4_X1 U9674 ( .A1(\SB1_3_31/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_31/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_3_31/Component_Function_2/NAND4_in[2] ), .A4(n4662), .ZN(n5490)
         );
  NAND4_X1 U9676 ( .A1(\SB1_3_31/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_31/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_3_31/Component_Function_2/NAND4_in[2] ), .A4(n4662), .ZN(
        \SB2_3_28/i0_0 ) );
  NAND3_X2 U9678 ( .A1(\SB1_3_31/i1_5 ), .A2(\SB1_3_31/i0[10] ), .A3(
        \SB1_3_31/i1[9] ), .ZN(\SB1_3_31/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U9685 ( .A1(\SB2_3_19/i0[10] ), .A2(\SB2_3_19/i0_3 ), .A3(
        \SB2_3_19/i0[9] ), .ZN(n3291) );
  NAND3_X2 U9688 ( .A1(\SB3_11/i0[9] ), .A2(\SB3_11/i0_3 ), .A3(
        \SB3_11/i0[10] ), .ZN(n3556) );
  BUF_X2 U9689 ( .I(\SB3_11/buf_output[4] ), .Z(\SB4_10/i0_4 ) );
  BUF_X4 U9690 ( .I(\SB2_3_6/buf_output[2] ), .Z(\RI5[3][170] ) );
  NAND3_X1 U9695 ( .A1(\SB1_2_12/i0_0 ), .A2(\SB1_2_12/i0_3 ), .A3(
        \SB1_2_12/i0_4 ), .ZN(\SB1_2_12/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U9696 ( .A1(\SB2_2_10/i0[10] ), .A2(n581), .A3(\SB2_2_10/i0_3 ), 
        .ZN(\SB2_2_10/Component_Function_0/NAND4_in[2] ) );
  CLKBUF_X4 U9697 ( .I(\MC_ARK_ARC_1_3/buf_output[137] ), .Z(\SB3_9/i0_3 ) );
  NAND3_X1 U9698 ( .A1(\SB3_9/i1[9] ), .A2(\SB3_9/i0_4 ), .A3(\SB3_9/i0_3 ), 
        .ZN(\SB3_9/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U9699 ( .A1(\RI1[3][143] ), .A2(\SB1_3_8/i0_0 ), .A3(
        \SB1_3_8/i0[7] ), .ZN(\SB1_3_8/Component_Function_0/NAND4_in[3] ) );
  CLKBUF_X4 U9705 ( .I(\MC_ARK_ARC_1_3/buf_output[108] ), .Z(\SB3_13/i0[9] )
         );
  NAND3_X1 U9710 ( .A1(\SB1_2_20/i0[9] ), .A2(\SB1_2_20/i0[10] ), .A3(
        \SB1_2_20/i0_3 ), .ZN(\SB1_2_20/Component_Function_4/NAND4_in[2] ) );
  NAND4_X1 U9712 ( .A1(\SB4_19/Component_Function_3/NAND4_in[1] ), .A2(
        \SB4_19/Component_Function_3/NAND4_in[3] ), .A3(n870), .A4(n1228), 
        .ZN(n729) );
  NAND3_X1 U9714 ( .A1(\SB3_27/i0[9] ), .A2(\SB3_27/i0_3 ), .A3(\SB3_27/i0[8] ), .ZN(n2976) );
  NAND3_X1 U9717 ( .A1(\SB3_27/i0_3 ), .A2(\SB3_27/i0_0 ), .A3(\SB3_27/i0[7] ), 
        .ZN(n6264) );
  BUF_X2 U9720 ( .I(\MC_ARK_ARC_1_1/buf_output[180] ), .Z(\SB1_2_1/i0[9] ) );
  INV_X1 U9723 ( .I(\MC_ARK_ARC_1_1/buf_output[180] ), .ZN(\SB1_2_1/i3[0] ) );
  INV_X1 U9728 ( .I(\SB4_8/i1[9] ), .ZN(n5492) );
  NAND3_X1 U9735 ( .A1(\SB3_19/i0_3 ), .A2(\SB3_19/i0[8] ), .A3(\SB3_19/i0[9] ), .ZN(\SB3_19/Component_Function_2/NAND4_in[2] ) );
  CLKBUF_X4 U9736 ( .I(\MC_ARK_ARC_1_0/buf_output[119] ), .Z(\SB1_1_12/i0_3 )
         );
  NAND3_X1 U9737 ( .A1(\SB4_23/i0_0 ), .A2(\SB4_23/i0_3 ), .A3(\SB4_23/i0_4 ), 
        .ZN(\SB4_23/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U9738 ( .A1(\SB1_2_4/i0_0 ), .A2(\SB1_2_4/i0[9] ), .A3(
        \SB1_2_4/i0[8] ), .ZN(n1556) );
  NAND3_X1 U9739 ( .A1(\SB1_2_4/i0_3 ), .A2(\SB1_2_4/i0[8] ), .A3(
        \SB1_2_4/i0[9] ), .ZN(\SB1_2_4/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U9740 ( .A1(\SB2_3_20/i0_3 ), .A2(\SB2_3_20/i0[10] ), .A3(
        \SB2_3_20/i0[9] ), .ZN(n3708) );
  INV_X1 U9742 ( .I(\MC_ARK_ARC_1_1/buf_output[171] ), .ZN(\SB1_2_3/i0[8] ) );
  NAND3_X1 U9743 ( .A1(\SB1_2_3/i0[9] ), .A2(\SB1_2_3/i0_3 ), .A3(
        \SB1_2_3/i0[8] ), .ZN(n4252) );
  NAND3_X1 U9744 ( .A1(\SB1_2_3/i0[8] ), .A2(\SB1_2_3/i3[0] ), .A3(
        \SB1_2_3/i1_5 ), .ZN(n880) );
  INV_X1 U9746 ( .I(n355), .ZN(\SB1_0_24/i0[8] ) );
  BUF_X2 U9748 ( .I(n355), .Z(\SB1_0_24/i0[10] ) );
  NAND3_X1 U9749 ( .A1(\SB4_13/i0_3 ), .A2(n3683), .A3(\SB4_13/i0[9] ), .ZN(
        \SB4_13/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U9750 ( .A1(\SB3_15/i1[9] ), .A2(\SB3_15/i1_5 ), .A3(
        \SB3_15/i0[10] ), .ZN(\SB3_15/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U9751 ( .A1(\SB3_15/i0_3 ), .A2(\SB3_15/i1[9] ), .A3(\SB3_15/i0[6] ), .ZN(\SB3_15/Component_Function_3/NAND4_in[0] ) );
  NAND2_X1 U9755 ( .A1(\SB3_1/Component_Function_3/NAND4_in[0] ), .A2(n4668), 
        .ZN(n5558) );
  BUF_X2 U9757 ( .I(\SB3_26/buf_output[0] ), .Z(\SB4_21/i0[9] ) );
  NAND2_X1 U9758 ( .A1(\SB2_3_24/i0_3 ), .A2(\SB2_3_24/i1[9] ), .ZN(
        \SB2_3_24/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U9761 ( .A1(\SB2_3_24/i0_3 ), .A2(\SB2_3_24/i1[9] ), .A3(
        \SB2_3_24/i0_4 ), .ZN(\SB2_3_24/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U9769 ( .A1(\SB2_3_24/i0_3 ), .A2(\SB2_3_24/i1[9] ), .A3(
        \SB2_3_24/i0[6] ), .ZN(\SB2_3_24/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U9771 ( .A1(\SB1_3_26/buf_output[3] ), .A2(\SB2_3_24/i1[9] ), .A3(
        \SB2_3_24/i1_7 ), .ZN(n3435) );
  NAND3_X1 U9774 ( .A1(\SB2_3_24/i1_5 ), .A2(\SB1_3_26/buf_output[3] ), .A3(
        \SB2_3_24/i1[9] ), .ZN(\SB2_3_24/Component_Function_2/NAND4_in[0] ) );
  CLKBUF_X4 U9776 ( .I(\MC_ARK_ARC_1_3/buf_output[74] ), .Z(\SB3_19/i0_0 ) );
  NAND3_X1 U9777 ( .A1(\SB4_4/i1_5 ), .A2(\SB3_7/buf_output[2] ), .A3(
        \SB4_4/i0_4 ), .ZN(\SB4_4/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U9781 ( .A1(\SB3_16/i0[8] ), .A2(\SB3_16/i3[0] ), .A3(\SB3_16/i1_5 ), .ZN(n2131) );
  CLKBUF_X4 U9782 ( .I(\MC_ARK_ARC_1_3/buf_output[95] ), .Z(\SB3_16/i0_3 ) );
  BUF_X2 U9783 ( .I(\SB3_23/buf_output[2] ), .Z(\SB4_20/i0_0 ) );
  NAND3_X1 U9784 ( .A1(\SB4_8/i0_0 ), .A2(\SB4_8/i0_4 ), .A3(\SB4_8/i0_3 ), 
        .ZN(n6369) );
  CLKBUF_X4 U9789 ( .I(\MC_ARK_ARC_1_1/buf_output[80] ), .Z(\SB1_2_18/i0_0 )
         );
  NAND3_X1 U9793 ( .A1(\SB3_24/i0_4 ), .A2(\SB3_24/i0_3 ), .A3(\SB3_24/i1[9] ), 
        .ZN(n2578) );
  NAND3_X1 U9798 ( .A1(\SB4_8/i0[6] ), .A2(\SB4_8/i0_3 ), .A3(\SB4_8/i1[9] ), 
        .ZN(n6514) );
  NAND3_X1 U9801 ( .A1(\SB3_14/i0[10] ), .A2(\SB3_14/i1[9] ), .A3(
        \SB3_14/i1_7 ), .ZN(n5537) );
  NAND3_X1 U9802 ( .A1(\SB3_14/i0[10] ), .A2(\SB3_14/i0_3 ), .A3(
        \SB3_14/i0[6] ), .ZN(n6174) );
  NAND3_X1 U9806 ( .A1(\SB3_14/i0_3 ), .A2(\SB3_14/i0[10] ), .A3(
        \SB3_14/i0[9] ), .ZN(n6134) );
  NAND3_X1 U9807 ( .A1(\SB4_27/i0_3 ), .A2(\SB4_27/i0[10] ), .A3(
        \SB4_27/i0[6] ), .ZN(\SB4_27/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U9809 ( .A1(\SB3_18/i0[7] ), .A2(\SB3_18/i0_3 ), .A3(\SB3_18/i0_0 ), 
        .ZN(\SB3_18/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U9813 ( .A1(\SB4_21/i0[6] ), .A2(n3666), .A3(\SB4_21/i0_3 ), .ZN(
        n6455) );
  CLKBUF_X4 U9815 ( .I(\SB1_1_30/buf_output[5] ), .Z(\SB2_1_30/i0_3 ) );
  NAND3_X1 U9816 ( .A1(\SB1_2_17/i1_5 ), .A2(\SB1_2_17/i0[10] ), .A3(
        \SB1_2_17/i1[9] ), .ZN(\SB1_2_17/Component_Function_2/NAND4_in[0] ) );
  CLKBUF_X4 U9817 ( .I(\MC_ARK_ARC_1_3/buf_output[152] ), .Z(\SB3_6/i0_0 ) );
  INV_X1 U9818 ( .I(\MC_ARK_ARC_1_3/buf_output[57] ), .ZN(\SB3_22/i0[8] ) );
  BUF_X2 U9819 ( .I(\MC_ARK_ARC_1_3/buf_output[57] ), .Z(\SB3_22/i0[10] ) );
  CLKBUF_X4 U9821 ( .I(\SB3_22/buf_output[4] ), .Z(\SB4_21/i0_4 ) );
  NAND2_X1 U9824 ( .A1(\SB1_3_28/i0_3 ), .A2(\SB1_3_28/i1[9] ), .ZN(
        \SB1_3_28/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U9825 ( .A1(\SB1_3_28/i0[10] ), .A2(\SB1_3_28/i1[9] ), .A3(
        \SB1_3_28/i1_7 ), .ZN(n2316) );
  CLKBUF_X4 U9826 ( .I(\MC_ARK_ARC_1_2/buf_output[22] ), .Z(\SB1_3_28/i0_4 )
         );
  NAND3_X1 U9831 ( .A1(\SB1_1_12/i0_3 ), .A2(\SB1_1_12/i0[8] ), .A3(
        \SB1_1_12/i1_7 ), .ZN(\SB1_1_12/Component_Function_1/NAND4_in[1] ) );
  CLKBUF_X8 U9832 ( .I(\SB1_0_16/buf_output[3] ), .Z(\RI3[0][105] ) );
  CLKBUF_X4 U9836 ( .I(\SB1_2_20/buf_output[3] ), .Z(\SB2_2_18/i0[10] ) );
  CLKBUF_X4 U9842 ( .I(\SB3_4/buf_output[2] ), .Z(\SB4_1/i0_0 ) );
  BUF_X2 U9843 ( .I(n363), .Z(\SB1_0_20/i0[10] ) );
  INV_X1 U9844 ( .I(n363), .ZN(\SB1_0_20/i0[8] ) );
  INV_X1 U9845 ( .I(\SB3_20/buf_output[2] ), .ZN(\SB4_17/i1[9] ) );
  BUF_X4 U9846 ( .I(\SB2_2_6/buf_output[3] ), .Z(\RI5[2][165] ) );
  AND4_X2 U9851 ( .A1(\SB1_3_22/Component_Function_2/NAND4_in[0] ), .A2(n1245), 
        .A3(\SB1_3_22/Component_Function_2/NAND4_in[2] ), .A4(n5902), .Z(n5494) );
  NAND3_X1 U9853 ( .A1(\SB1_3_18/i0[10] ), .A2(\SB1_3_18/i0_4 ), .A3(
        \SB1_3_18/i0_3 ), .ZN(\SB1_3_18/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U9854 ( .A1(\SB2_0_26/i3[0] ), .A2(\SB2_0_26/i0_0 ), .A3(
        \SB2_0_26/i1_7 ), .ZN(\SB2_0_26/Component_Function_4/NAND4_in[1] ) );
  NAND2_X1 U9855 ( .A1(\SB2_0_26/i0_0 ), .A2(\SB2_0_26/i3[0] ), .ZN(n1795) );
  NAND3_X1 U9859 ( .A1(\SB2_0_26/i0_0 ), .A2(\SB2_0_26/i1_5 ), .A3(
        \RI3[0][34] ), .ZN(\SB2_0_26/Component_Function_2/NAND4_in[3] ) );
  NAND3_X1 U9861 ( .A1(\SB2_0_26/i0_3 ), .A2(\SB2_0_26/i0_0 ), .A3(
        \RI3[0][34] ), .ZN(\SB2_0_26/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U9862 ( .A1(\SB3_8/i0_3 ), .A2(\SB3_8/i0[9] ), .A3(\SB3_8/i0[10] ), 
        .ZN(n5838) );
  NAND3_X1 U9866 ( .A1(\SB3_8/i0_3 ), .A2(\SB3_8/i0[10] ), .A3(\SB3_8/i0[6] ), 
        .ZN(\SB3_8/Component_Function_2/NAND4_in[1] ) );
  CLKBUF_X4 U9867 ( .I(\MC_ARK_ARC_1_1/buf_output[174] ), .Z(\SB1_2_2/i0[9] )
         );
  BUF_X2 U9869 ( .I(\MC_ARK_ARC_1_3/buf_output[190] ), .Z(\SB3_0/i0_4 ) );
  INV_X1 U9870 ( .I(\MC_ARK_ARC_1_3/buf_output[190] ), .ZN(\SB3_0/i0[7] ) );
  CLKBUF_X4 U9876 ( .I(\MC_ARK_ARC_1_3/buf_output[26] ), .Z(\SB3_27/i0_0 ) );
  CLKBUF_X12 U9877 ( .I(Key[191]), .Z(n241) );
  BUF_X2 U9879 ( .I(\MC_ARK_ARC_1_1/buf_output[115] ), .Z(\SB1_2_12/i0[6] ) );
  BUF_X2 U9881 ( .I(\SB1_2_12/buf_output[1] ), .Z(\SB2_2_8/i0[6] ) );
  NAND3_X1 U9886 ( .A1(n3651), .A2(\SB2_3_12/i0[7] ), .A3(\SB2_3_12/i0[6] ), 
        .ZN(\SB2_3_12/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U9889 ( .A1(\SB2_2_31/i1_5 ), .A2(\SB2_2_31/i0[8] ), .A3(
        \SB2_2_31/i3[0] ), .ZN(\SB2_2_31/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U9890 ( .A1(\SB3_16/i0[7] ), .A2(\SB3_16/i0_3 ), .A3(\SB3_16/i0_0 ), 
        .ZN(\SB3_16/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U9891 ( .A1(\SB3_16/i1[9] ), .A2(\SB3_16/i0_4 ), .A3(\SB3_16/i0_3 ), 
        .ZN(\SB3_16/Component_Function_5/NAND4_in[2] ) );
  BUF_X2 U9892 ( .I(\SB3_24/buf_output[3] ), .Z(\SB4_22/i0[10] ) );
  CLKBUF_X4 U9893 ( .I(\SB3_12/buf_output[5] ), .Z(\SB4_12/i0_3 ) );
  XOR2_X1 U9896 ( .A1(Key[148]), .A2(Plaintext[148]), .Z(n5496) );
  CLKBUF_X4 U9905 ( .I(\SB3_6/buf_output[4] ), .Z(\SB4_5/i0_4 ) );
  CLKBUF_X4 U9906 ( .I(\SB1_3_2/buf_output[1] ), .Z(\SB2_3_30/i0[6] ) );
  INV_X1 U9907 ( .I(\SB3_10/buf_output[2] ), .ZN(\SB4_7/i1[9] ) );
  NAND3_X1 U9912 ( .A1(\SB2_3_14/i1[9] ), .A2(\SB2_3_14/i0_3 ), .A3(
        \SB2_3_14/i0[6] ), .ZN(\SB2_3_14/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U9914 ( .A1(\SB2_3_14/i0[10] ), .A2(\SB2_3_14/i1_7 ), .A3(
        \SB2_3_14/i1[9] ), .ZN(n2657) );
  NAND3_X1 U9918 ( .A1(\SB1_3_17/i0[10] ), .A2(\SB1_3_17/i0_3 ), .A3(
        \SB1_3_17/i0[9] ), .ZN(n6397) );
  NAND3_X1 U9922 ( .A1(\SB1_3_17/i0_4 ), .A2(\SB1_3_17/i0[10] ), .A3(
        \SB1_3_17/i0_3 ), .ZN(n4098) );
  NAND3_X1 U9925 ( .A1(\SB1_3_17/i0[10] ), .A2(\SB1_3_17/i1[9] ), .A3(
        \SB1_3_17/i1_7 ), .ZN(n2226) );
  CLKBUF_X4 U9930 ( .I(\MC_ARK_ARC_1_2/buf_output[87] ), .Z(\SB1_3_17/i0[10] )
         );
  CLKBUF_X12 U9934 ( .I(\SB2_0_0/buf_output[2] ), .Z(n5497) );
  CLKBUF_X12 U9936 ( .I(\SB2_0_0/buf_output[2] ), .Z(\RI5[0][14] ) );
  CLKBUF_X4 U9938 ( .I(\SB2_2_4/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_2/buf_datainput[0] ) );
  NAND3_X1 U9940 ( .A1(\SB4_8/i1_7 ), .A2(\SB4_8/i0[8] ), .A3(\SB4_8/i0_4 ), 
        .ZN(\SB4_8/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U9945 ( .A1(\SB4_8/i0[10] ), .A2(\SB4_8/i0_3 ), .A3(\SB4_8/i0_4 ), 
        .ZN(\SB4_8/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U9946 ( .A1(Key[41]), .A2(Plaintext[41]), .Z(n5498) );
  BUF_X4 U9947 ( .I(\MC_ARK_ARC_1_0/buf_output[88] ), .Z(\SB1_1_17/i0_4 ) );
  XOR2_X1 U9948 ( .A1(\MC_ARK_ARC_1_3/temp6[134] ), .A2(
        \MC_ARK_ARC_1_3/temp5[134] ), .Z(n5499) );
  NAND3_X1 U9952 ( .A1(\SB3_9/i0[9] ), .A2(\SB3_9/i0[10] ), .A3(\SB3_9/i0_3 ), 
        .ZN(\SB3_9/Component_Function_4/NAND4_in[2] ) );
  CLKBUF_X4 U9953 ( .I(\RI3[0][57] ), .Z(\SB2_0_22/i0[10] ) );
  NAND3_X1 U9954 ( .A1(\SB4_22/i0[10] ), .A2(\SB4_22/i1_5 ), .A3(
        \SB4_22/i1[9] ), .ZN(n4242) );
  NAND3_X1 U9957 ( .A1(\SB1_3_31/i0[10] ), .A2(\SB1_3_31/i1[9] ), .A3(
        \SB1_3_31/i1_7 ), .ZN(n3420) );
  NAND3_X1 U9958 ( .A1(\SB1_3_31/i1[9] ), .A2(\SB1_3_31/i1_5 ), .A3(
        \MC_ARK_ARC_1_2/buf_output[4] ), .ZN(
        \SB1_3_31/Component_Function_4/NAND4_in[3] ) );
  INV_X1 U9960 ( .I(\SB3_22/buf_output[2] ), .ZN(\SB4_19/i1[9] ) );
  CLKBUF_X2 U9962 ( .I(\SB3_22/buf_output[2] ), .Z(\SB4_19/i0_0 ) );
  NAND3_X1 U9963 ( .A1(\SB2_3_14/i0_3 ), .A2(\SB1_3_19/buf_output[0] ), .A3(
        \SB2_3_14/i0[10] ), .ZN(\SB2_3_14/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U9966 ( .A1(\SB3_23/i0[9] ), .A2(\SB3_23/i0[6] ), .A3(\SB3_23/i0_4 ), .ZN(n954) );
  NAND3_X1 U9967 ( .A1(\SB1_2_8/i0_0 ), .A2(\SB1_2_8/i0_4 ), .A3(
        \SB1_2_8/i1_5 ), .ZN(n5959) );
  CLKBUF_X4 U9970 ( .I(\MC_ARK_ARC_1_2/buf_output[176] ), .Z(\SB1_3_2/i0_0 )
         );
  CLKBUF_X4 U9971 ( .I(\SB1_2_31/buf_output[2] ), .Z(\SB2_2_28/i0_0 ) );
  CLKBUF_X4 U9980 ( .I(\MC_ARK_ARC_1_1/buf_output[154] ), .Z(\SB1_2_6/i0_4 )
         );
  NAND3_X1 U9981 ( .A1(\SB4_22/i1_7 ), .A2(\SB4_22/i0[8] ), .A3(\SB4_22/i0_4 ), 
        .ZN(\SB4_22/Component_Function_1/NAND4_in[3] ) );
  INV_X1 U9987 ( .I(\SB1_0_30/i0_4 ), .ZN(\SB1_0_30/i0[7] ) );
  NAND3_X1 U9988 ( .A1(\SB1_3_23/i0_0 ), .A2(\SB1_3_23/i0_3 ), .A3(
        \SB1_3_23/i0_4 ), .ZN(\SB1_3_23/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U9994 ( .A1(\SB2_2_24/i0[10] ), .A2(\SB2_2_24/i0[9] ), .A3(
        \SB2_2_24/i0_3 ), .ZN(n2665) );
  CLKBUF_X4 U9996 ( .I(\SB1_2_26/buf_output[3] ), .Z(\SB2_2_24/i0[10] ) );
  NAND3_X1 U9997 ( .A1(\SB1_2_24/i0[10] ), .A2(\SB1_2_24/i1[9] ), .A3(n2913), 
        .ZN(\SB1_2_24/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U9998 ( .A1(\MC_ARK_ARC_1_1/temp5[101] ), .A2(
        \MC_ARK_ARC_1_1/temp6[101] ), .Z(n5500) );
  CLKBUF_X4 U10001 ( .I(\MC_ARK_ARC_1_2/buf_output[58] ), .Z(\SB1_3_22/i0_4 )
         );
  NAND3_X1 U10003 ( .A1(\SB3_19/i0_0 ), .A2(\SB3_19/i1_5 ), .A3(\SB3_19/i0_4 ), 
        .ZN(n3863) );
  NAND2_X1 U10004 ( .A1(\SB2_2_22/i0_3 ), .A2(\SB2_2_22/i1[9] ), .ZN(
        \SB2_2_22/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U10005 ( .A1(\SB1_0_17/i0_3 ), .A2(\SB1_0_17/i0[8] ), .A3(
        \SB1_0_17/i0[9] ), .ZN(\SB1_0_17/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U10006 ( .A1(\SB1_0_17/i0[10] ), .A2(n2899), .A3(\SB1_0_17/i0_3 ), 
        .ZN(\SB1_0_17/Component_Function_0/NAND4_in[2] ) );
  CLKBUF_X4 U10007 ( .I(\SB1_0_16/buf_output[2] ), .Z(\SB2_0_13/i0_0 ) );
  CLKBUF_X4 U10008 ( .I(\SB1_0_30/buf_output[5] ), .Z(\SB2_0_30/i0_3 ) );
  INV_X1 U10010 ( .I(\SB1_0_30/buf_output[5] ), .ZN(\SB2_0_30/i1_5 ) );
  INV_X1 U10011 ( .I(n388), .ZN(\SB1_0_8/i0[7] ) );
  NAND3_X1 U10013 ( .A1(\SB2_3_9/i0_3 ), .A2(\SB2_3_9/i1_7 ), .A3(
        \SB2_3_9/i0[8] ), .ZN(\SB2_3_9/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U10016 ( .A1(\SB2_3_11/i0[8] ), .A2(\SB2_3_11/i1_7 ), .A3(n3645), 
        .ZN(\SB2_3_11/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U10017 ( .A1(\SB2_3_11/i0_3 ), .A2(\SB2_3_11/i1_7 ), .A3(
        \SB2_3_11/i0[8] ), .ZN(\SB2_3_11/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U10022 ( .A1(\SB2_1_0/i0_3 ), .A2(\SB2_1_0/i1[9] ), .A3(n2687), 
        .ZN(\SB2_1_0/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 U10024 ( .A1(\SB2_1_0/i0_3 ), .A2(\SB2_1_0/i1[9] ), .ZN(
        \SB2_1_0/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U10025 ( .A1(\SB2_1_0/i1[9] ), .A2(\SB2_1_0/i0_3 ), .A3(
        \SB2_1_0/i0[6] ), .ZN(\SB2_1_0/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U10026 ( .A1(\SB2_1_0/i0[10] ), .A2(\SB2_1_0/i1[9] ), .A3(
        \SB2_1_0/i1_7 ), .ZN(\SB2_1_0/Component_Function_3/NAND4_in[2] ) );
  BUF_X4 U10027 ( .I(\MC_ARK_ARC_1_1/buf_output[137] ), .Z(\SB1_2_9/i0_3 ) );
  CLKBUF_X4 U10031 ( .I(\SB2_1_1/buf_output[3] ), .Z(\RI5[1][3] ) );
  CLKBUF_X4 U10032 ( .I(\SB2_0_29/buf_output[1] ), .Z(\RI5[0][37] ) );
  NAND3_X1 U10033 ( .A1(\SB2_0_13/i3[0] ), .A2(\SB2_0_13/i0_0 ), .A3(
        \SB2_0_13/i1_7 ), .ZN(\SB2_0_13/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U10038 ( .A1(n2621), .A2(\MC_ARK_ARC_1_2/temp6[135] ), .Z(n5501) );
  XOR2_X1 U10039 ( .A1(\MC_ARK_ARC_1_2/temp6[135] ), .A2(n2621), .Z(n5502) );
  NAND3_X1 U10040 ( .A1(\SB1_0_25/i0_0 ), .A2(\SB1_0_25/i0[9] ), .A3(
        \SB1_0_25/i0[8] ), .ZN(\SB1_0_25/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U10041 ( .A1(\SB2_0_1/i0_3 ), .A2(\SB2_0_1/i1_7 ), .A3(
        \SB2_0_1/i0[8] ), .ZN(\SB2_0_1/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U10048 ( .A1(\SB2_0_1/i0_3 ), .A2(\SB2_0_1/i1[9] ), .A3(
        \SB2_0_1/i0_4 ), .ZN(\SB2_0_1/Component_Function_5/NAND4_in[2] ) );
  CLKBUF_X4 U10053 ( .I(\SB1_2_18/buf_output[4] ), .Z(\SB2_2_17/i0_4 ) );
  CLKBUF_X4 U10058 ( .I(\RI1[4][143] ), .Z(\SB3_8/i0_3 ) );
  INV_X1 U10060 ( .I(\RI1[4][143] ), .ZN(\SB3_8/i1_5 ) );
  NAND3_X1 U10061 ( .A1(\SB3_8/i1[9] ), .A2(\SB3_8/i0_3 ), .A3(\SB3_8/i0[6] ), 
        .ZN(\SB3_8/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U10062 ( .A1(\SB3_8/i0_3 ), .A2(\SB3_8/i1[9] ), .A3(\SB3_8/i0_4 ), 
        .ZN(n2889) );
  NAND3_X1 U10065 ( .A1(\SB3_8/i0_3 ), .A2(\SB3_8/i0_4 ), .A3(\SB3_8/i0_0 ), 
        .ZN(\SB3_8/Component_Function_3/NAND4_in[1] ) );
  CLKBUF_X4 U10068 ( .I(\SB3_9/buf_output[4] ), .Z(\SB4_8/i0_4 ) );
  NAND3_X1 U10076 ( .A1(\SB2_0_11/i0[8] ), .A2(\SB2_0_11/i0[7] ), .A3(
        \SB2_0_11/i0[6] ), .ZN(\SB2_0_11/Component_Function_0/NAND4_in[1] ) );
  CLKBUF_X4 U10077 ( .I(n5488), .Z(\SB3_30/i0_0 ) );
  NAND2_X1 U10082 ( .A1(\SB1_3_10/i0[10] ), .A2(\SB1_3_10/i0[9] ), .ZN(
        \SB1_3_10/Component_Function_0/NAND4_in[0] ) );
  NAND3_X1 U10083 ( .A1(n1388), .A2(\SB1_3_10/i0[10] ), .A3(\SB1_3_10/i0_4 ), 
        .ZN(\SB1_3_10/Component_Function_0/NAND4_in[2] ) );
  INV_X1 U10084 ( .I(\SB1_3_24/buf_output[1] ), .ZN(\SB2_3_20/i1_7 ) );
  NAND3_X1 U10085 ( .A1(\SB2_2_27/i0_3 ), .A2(\SB2_2_27/i1_7 ), .A3(
        \SB2_2_27/i0[8] ), .ZN(\SB2_2_27/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U10086 ( .A1(\SB1_2_28/buf_output[4] ), .A2(\SB2_2_27/i1_7 ), .A3(
        \SB2_2_27/i0[8] ), .ZN(n3917) );
  NAND3_X1 U10092 ( .A1(\SB2_2_27/i0[8] ), .A2(\SB2_2_27/i3[0] ), .A3(
        \SB2_2_27/i1_5 ), .ZN(\SB2_2_27/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U10095 ( .A1(\SB2_0_3/i1_5 ), .A2(\SB2_0_3/i0[8] ), .A3(
        \SB2_0_3/i3[0] ), .ZN(\SB2_0_3/Component_Function_3/NAND4_in[3] ) );
  CLKBUF_X8 U10096 ( .I(\SB2_2_14/i0_4 ), .Z(n5932) );
  CLKBUF_X4 U10098 ( .I(\SB1_3_24/buf_output[3] ), .Z(\SB2_3_22/i0[10] ) );
  BUF_X2 U10099 ( .I(\MC_ARK_ARC_1_3/buf_output[79] ), .Z(\SB3_18/i0[6] ) );
  NAND3_X1 U10101 ( .A1(\SB3_11/i0_3 ), .A2(\SB3_11/i0[10] ), .A3(
        \SB3_11/i0[6] ), .ZN(\SB3_11/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U10103 ( .A1(\SB3_11/i0[10] ), .A2(\SB3_11/i0_4 ), .A3(
        \SB3_11/i0_3 ), .ZN(\SB3_11/Component_Function_0/NAND4_in[2] ) );
  CLKBUF_X4 U10107 ( .I(\MC_ARK_ARC_1_3/buf_output[123] ), .Z(\SB3_11/i0[10] )
         );
  NAND3_X1 U10109 ( .A1(\SB1_1_19/i0_3 ), .A2(\SB1_1_19/i0[10] ), .A3(
        \SB1_1_19/i0[6] ), .ZN(\SB1_1_19/Component_Function_2/NAND4_in[1] ) );
  CLKBUF_X4 U10110 ( .I(\MC_ARK_ARC_1_3/buf_output[69] ), .Z(\SB3_20/i0[10] )
         );
  BUF_X2 U10111 ( .I(\SB3_20/buf_output[1] ), .Z(\SB4_16/i0[6] ) );
  INV_X1 U10114 ( .I(\SB3_20/buf_output[1] ), .ZN(\SB4_16/i1_7 ) );
  NAND3_X1 U10121 ( .A1(\SB4_8/i1[9] ), .A2(\SB4_8/i1_5 ), .A3(\SB4_8/i0_4 ), 
        .ZN(\SB4_8/Component_Function_4/NAND4_in[3] ) );
  BUF_X2 U10123 ( .I(\MC_ARK_ARC_1_1/buf_output[91] ), .Z(\SB1_2_16/i0[6] ) );
  INV_X1 U10126 ( .I(\MC_ARK_ARC_1_1/buf_output[91] ), .ZN(\SB1_2_16/i1_7 ) );
  BUF_X2 U10129 ( .I(\SB3_1/buf_output[0] ), .Z(\SB4_28/i0[9] ) );
  INV_X1 U10133 ( .I(\SB3_1/buf_output[0] ), .ZN(\SB4_28/i3[0] ) );
  NAND3_X1 U10136 ( .A1(\SB3_24/i0_4 ), .A2(\SB3_24/i0_3 ), .A3(
        \SB3_24/i0[10] ), .ZN(n4331) );
  NAND3_X1 U10137 ( .A1(\SB3_24/i0[10] ), .A2(\SB3_24/i1[9] ), .A3(
        \SB3_24/i1_5 ), .ZN(n3759) );
  NAND3_X1 U10139 ( .A1(\SB2_2_25/i0_4 ), .A2(\SB2_2_25/i1_5 ), .A3(
        \SB2_2_25/i1[9] ), .ZN(n796) );
  NAND3_X1 U10140 ( .A1(\SB1_1_8/i0_0 ), .A2(\RI1[1][143] ), .A3(
        \SB1_1_8/i0_4 ), .ZN(\SB1_1_8/Component_Function_3/NAND4_in[1] ) );
  NAND2_X1 U10143 ( .A1(\SB1_1_8/i0_0 ), .A2(\SB1_1_8/i3[0] ), .ZN(
        \SB1_1_8/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U10144 ( .A1(\SB1_1_8/i3[0] ), .A2(\SB1_1_8/i0_0 ), .A3(
        \SB1_1_8/i1_7 ), .ZN(\SB1_1_8/Component_Function_4/NAND4_in[1] ) );
  INV_X4 U10145 ( .I(n2738), .ZN(\SB2_0_10/i0_4 ) );
  NAND2_X1 U10146 ( .A1(n1687), .A2(\SB3_3/Component_Function_2/NAND4_in[2] ), 
        .ZN(n5563) );
  NAND3_X1 U10152 ( .A1(\SB1_1_18/i0_4 ), .A2(\SB1_1_18/i1[9] ), .A3(
        \SB1_1_18/i1_5 ), .ZN(n2637) );
  CLKBUF_X4 U10153 ( .I(\SB2_2_24/buf_output[3] ), .Z(\RI5[2][57] ) );
  NAND3_X1 U10154 ( .A1(\SB3_3/i0[9] ), .A2(\SB3_3/i0_3 ), .A3(\SB3_3/i0[8] ), 
        .ZN(\SB3_3/Component_Function_2/NAND4_in[2] ) );
  CLKBUF_X4 U10159 ( .I(\MC_ARK_ARC_1_3/buf_output[172] ), .Z(\SB3_3/i0_4 ) );
  NAND3_X1 U10160 ( .A1(\SB2_3_19/i0[10] ), .A2(\SB2_3_19/i0_3 ), .A3(
        \SB2_3_19/i0_4 ), .ZN(n2112) );
  NAND3_X1 U10161 ( .A1(\SB2_3_19/i0_3 ), .A2(\SB2_3_19/i0_0 ), .A3(
        \SB2_3_19/i0_4 ), .ZN(\SB2_3_19/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U10162 ( .A1(\SB2_3_19/i0[6] ), .A2(\SB2_3_19/i0[9] ), .A3(
        \SB2_3_19/i0_4 ), .ZN(n3531) );
  NAND3_X1 U10163 ( .A1(\SB1_2_26/i0[10] ), .A2(\SB1_2_26/i0_4 ), .A3(
        \RI1[2][35] ), .ZN(\SB1_2_26/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U10167 ( .A1(n3569), .A2(n3568), .Z(n5504) );
  NAND4_X1 U10170 ( .A1(\SB3_17/Component_Function_3/NAND4_in[0] ), .A2(n4551), 
        .A3(n3963), .A4(n3960), .ZN(n5505) );
  NAND4_X1 U10171 ( .A1(\SB3_17/Component_Function_3/NAND4_in[0] ), .A2(n4551), 
        .A3(n3963), .A4(n3960), .ZN(\SB3_17/buf_output[3] ) );
  CLKBUF_X4 U10172 ( .I(\MC_ARK_ARC_1_3/buf_output[188] ), .Z(\SB3_0/i0_0 ) );
  XOR2_X1 U10173 ( .A1(n4115), .A2(n4114), .Z(n5506) );
  CLKBUF_X4 U10174 ( .I(\MC_ARK_ARC_1_3/buf_output[94] ), .Z(\SB3_16/i0_4 ) );
  NAND3_X1 U10178 ( .A1(\SB4_16/i0_3 ), .A2(\SB4_16/i0_4 ), .A3(\SB4_16/i1[9] ), .ZN(n3791) );
  NAND3_X1 U10179 ( .A1(\SB4_16/i0[9] ), .A2(\SB4_16/i0_3 ), .A3(
        \SB4_16/i0[8] ), .ZN(\SB4_16/Component_Function_2/NAND4_in[2] ) );
  CLKBUF_X4 U10180 ( .I(\SB2_0_30/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[21] ) );
  CLKBUF_X4 U10181 ( .I(\SB3_16/buf_output[5] ), .Z(\SB4_16/i0_3 ) );
  NAND3_X1 U10182 ( .A1(\SB1_2_16/i1_5 ), .A2(\SB1_2_16/i1[9] ), .A3(
        \SB1_2_16/i0[10] ), .ZN(\SB1_2_16/Component_Function_2/NAND4_in[0] )
         );
  NAND3_X1 U10183 ( .A1(\SB1_2_16/i0[10] ), .A2(\RI1[2][95] ), .A3(
        \SB1_2_16/i0_4 ), .ZN(\SB1_2_16/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U10184 ( .A1(\SB1_2_16/i0_0 ), .A2(\SB1_2_16/i0[6] ), .A3(
        \SB1_2_16/i0[10] ), .ZN(\SB1_2_16/Component_Function_5/NAND4_in[1] )
         );
  CLKBUF_X4 U10185 ( .I(\MC_ARK_ARC_1_1/buf_output[93] ), .Z(\SB1_2_16/i0[10] ) );
  XOR2_X1 U10186 ( .A1(\MC_ARK_ARC_1_2/temp5[51] ), .A2(n6013), .Z(n5507) );
  INV_X1 U10187 ( .I(\MC_ARK_ARC_1_2/buf_output[6] ), .ZN(\SB1_3_30/i3[0] ) );
  NAND3_X1 U10188 ( .A1(\SB1_2_30/i0[10] ), .A2(\SB1_2_30/i0_4 ), .A3(
        \SB1_2_30/i0_3 ), .ZN(\SB1_2_30/Component_Function_0/NAND4_in[2] ) );
  CLKBUF_X4 U10189 ( .I(\MC_ARK_ARC_1_2/buf_output[92] ), .Z(\SB1_3_16/i0_0 )
         );
  INV_X1 U10191 ( .I(\MC_ARK_ARC_1_3/buf_output[107] ), .ZN(\SB3_14/i1_5 ) );
  CLKBUF_X4 U10192 ( .I(\MC_ARK_ARC_1_3/buf_output[107] ), .Z(\SB3_14/i0_3 )
         );
  XOR2_X1 U10195 ( .A1(\MC_ARK_ARC_1_3/temp6[11] ), .A2(
        \MC_ARK_ARC_1_3/temp5[11] ), .Z(n5508) );
  XOR2_X1 U10198 ( .A1(\MC_ARK_ARC_1_3/temp5[11] ), .A2(
        \MC_ARK_ARC_1_3/temp6[11] ), .Z(n5509) );
  NAND3_X1 U10200 ( .A1(\SB1_3_29/i0_3 ), .A2(\SB1_3_29/i0[8] ), .A3(
        \SB1_3_29/i0[9] ), .ZN(\SB1_3_29/Component_Function_2/NAND4_in[2] ) );
  BUF_X2 U10207 ( .I(\SB1_3_15/buf_output[3] ), .Z(\SB2_3_13/i0[10] ) );
  NAND3_X1 U10211 ( .A1(\SB2_3_24/i1_5 ), .A2(\SB2_3_24/i0_0 ), .A3(
        \SB2_3_24/i0_4 ), .ZN(\SB2_3_24/Component_Function_2/NAND4_in[3] ) );
  CLKBUF_X4 U10216 ( .I(\SB2_3_17/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_3/buf_datainput[114] ) );
  CLKBUF_X4 U10218 ( .I(\MC_ARK_ARC_1_2/buf_output[32] ), .Z(\SB1_3_26/i0_0 )
         );
  NAND3_X1 U10221 ( .A1(\SB1_3_16/i0[9] ), .A2(\SB1_3_16/i1_5 ), .A3(
        \SB1_3_16/i0[6] ), .ZN(n6358) );
  CLKBUF_X4 U10222 ( .I(\MC_ARK_ARC_1_2/buf_output[10] ), .Z(\SB1_3_30/i0_4 )
         );
  AND4_X2 U10223 ( .A1(\SB1_1_31/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_31/Component_Function_5/NAND4_in[3] ), .A3(n6024), .A4(
        \SB1_1_31/Component_Function_5/NAND4_in[0] ), .Z(n5510) );
  NAND4_X2 U10228 ( .A1(\SB1_3_30/Component_Function_3/NAND4_in[1] ), .A2(
        n4664), .A3(n6257), .A4(n6146), .ZN(n5511) );
  CLKBUF_X4 U10229 ( .I(\MC_ARK_ARC_1_1/buf_output[77] ), .Z(\SB1_2_19/i0_3 )
         );
  INV_X1 U10233 ( .I(\MC_ARK_ARC_1_1/buf_output[77] ), .ZN(\SB1_2_19/i1_5 ) );
  CLKBUF_X4 U10236 ( .I(\SB1_2_19/buf_output[3] ), .Z(\SB2_2_17/i0[10] ) );
  CLKBUF_X4 U10237 ( .I(\SB1_3_28/buf_output[4] ), .Z(\SB2_3_27/i0_4 ) );
  BUF_X4 U10240 ( .I(\MC_ARK_ARC_1_2/buf_output[95] ), .Z(\SB1_3_16/i0_3 ) );
  INV_X1 U10241 ( .I(\MC_ARK_ARC_1_2/buf_output[90] ), .ZN(\SB1_3_16/i3[0] )
         );
  BUF_X2 U10249 ( .I(\MC_ARK_ARC_1_2/buf_output[90] ), .Z(\SB1_3_16/i0[9] ) );
  INV_X1 U10250 ( .I(\MC_ARK_ARC_1_2/buf_output[109] ), .ZN(\SB1_3_13/i1_7 )
         );
  BUF_X2 U10255 ( .I(\MC_ARK_ARC_1_2/buf_output[109] ), .Z(\SB1_3_13/i0[6] )
         );
  NAND3_X1 U10258 ( .A1(\SB4_5/i0[10] ), .A2(\SB4_5/i0_4 ), .A3(\SB4_5/i0_3 ), 
        .ZN(\SB4_5/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U10259 ( .A1(\SB2_1_23/i0_3 ), .A2(\SB2_1_23/i0[10] ), .A3(
        \SB2_1_23/i0[9] ), .ZN(\SB2_1_23/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U10262 ( .A1(\SB2_1_23/i0_3 ), .A2(\SB2_1_23/i0_0 ), .A3(
        \SB2_1_23/i0_4 ), .ZN(\SB2_1_23/Component_Function_3/NAND4_in[1] ) );
  BUF_X2 U10264 ( .I(\MC_ARK_ARC_1_3/buf_output[170] ), .Z(\SB3_3/i0_0 ) );
  INV_X1 U10265 ( .I(\MC_ARK_ARC_1_3/buf_output[170] ), .ZN(\SB3_3/i1[9] ) );
  NAND3_X1 U10266 ( .A1(\SB4_1/i0_0 ), .A2(\SB4_1/i0[8] ), .A3(\SB4_1/i0[9] ), 
        .ZN(n5640) );
  NAND3_X1 U10267 ( .A1(\SB3_6/i1_5 ), .A2(\SB3_6/i0[6] ), .A3(\SB3_6/i0[9] ), 
        .ZN(\SB3_6/Component_Function_1/NAND4_in[2] ) );
  CLKBUF_X4 U10269 ( .I(\MC_ARK_ARC_1_3/buf_output[17] ), .Z(\SB3_29/i0_3 ) );
  NAND3_X1 U10271 ( .A1(\SB1_0_16/i0[9] ), .A2(\SB1_0_16/i0_3 ), .A3(
        \SB1_0_16/i0[10] ), .ZN(\SB1_0_16/Component_Function_4/NAND4_in[2] )
         );
  NAND3_X1 U10282 ( .A1(\SB1_0_16/i0[7] ), .A2(\SB1_0_16/i0_3 ), .A3(
        \SB1_0_16/i0_0 ), .ZN(\SB1_0_16/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U10286 ( .A1(\SB1_0_16/i0_3 ), .A2(\SB1_0_16/i1_7 ), .A3(
        \SB1_0_16/i0[8] ), .ZN(\SB1_0_16/Component_Function_1/NAND4_in[1] ) );
  NAND2_X1 U10289 ( .A1(\SB1_0_16/i0_3 ), .A2(\SB1_0_16/i1[9] ), .ZN(
        \SB1_0_16/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U10290 ( .A1(\SB1_0_16/i0_3 ), .A2(\SB1_0_16/i0[9] ), .A3(
        \SB1_0_16/i0[8] ), .ZN(n4189) );
  NAND3_X1 U10292 ( .A1(\SB1_0_16/i0_3 ), .A2(\SB1_0_16/i1[9] ), .A3(n4752), 
        .ZN(\SB1_0_16/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U10298 ( .A1(\SB2_0_22/i0_3 ), .A2(\SB2_0_22/i0[10] ), .A3(
        \SB2_0_22/i0[6] ), .ZN(\SB2_0_22/Component_Function_2/NAND4_in[1] ) );
  NAND3_X1 U10300 ( .A1(\SB4_2/i0_0 ), .A2(\SB4_2/i3[0] ), .A3(\SB4_2/i1_7 ), 
        .ZN(\SB4_2/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U10303 ( .A1(\SB1_2_16/i0[6] ), .A2(\SB1_2_16/i1[9] ), .A3(
        \RI1[2][95] ), .ZN(n6511) );
  NAND3_X1 U10307 ( .A1(\SB2_0_23/i0[10] ), .A2(\SB2_0_23/i0_3 ), .A3(
        \SB2_0_23/i0_4 ), .ZN(n3034) );
  NAND3_X1 U10308 ( .A1(\SB2_0_23/i0_3 ), .A2(\SB2_0_23/i0_4 ), .A3(
        \SB2_0_23/i1[9] ), .ZN(\SB2_0_23/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U10309 ( .A1(\SB2_0_23/i1[9] ), .A2(\SB2_0_23/i0_3 ), .A3(
        \SB2_0_23/i0[6] ), .ZN(\SB2_0_23/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U10311 ( .A1(\SB2_0_12/i1[9] ), .A2(\SB2_0_12/i0_3 ), .A3(
        \SB2_0_12/i0[6] ), .ZN(\SB2_0_12/Component_Function_3/NAND4_in[0] ) );
  BUF_X2 U10317 ( .I(\MC_ARK_ARC_1_2/buf_output[7] ), .Z(\SB1_3_30/i0[6] ) );
  INV_X1 U10319 ( .I(\MC_ARK_ARC_1_2/buf_output[7] ), .ZN(\SB1_3_30/i1_7 ) );
  INV_X1 U10320 ( .I(\MC_ARK_ARC_1_0/buf_output[24] ), .ZN(\SB1_1_27/i3[0] )
         );
  CLKBUF_X4 U10321 ( .I(\SB2_0_0/buf_output[1] ), .Z(\RI5[0][19] ) );
  NAND3_X1 U10328 ( .A1(\SB2_3_3/i0[10] ), .A2(\SB2_3_3/i1_5 ), .A3(
        \SB2_3_3/i1[9] ), .ZN(\SB2_3_3/Component_Function_2/NAND4_in[0] ) );
  NAND3_X1 U10329 ( .A1(\SB2_3_3/i0_4 ), .A2(\SB2_3_3/i1[9] ), .A3(
        \SB2_3_3/i1_5 ), .ZN(n6282) );
  NAND3_X1 U10335 ( .A1(\SB2_3_3/i1[9] ), .A2(\SB2_3_3/i0_3 ), .A3(
        \SB2_3_3/i0[6] ), .ZN(\SB2_3_3/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U10336 ( .A1(\SB2_3_3/i1[9] ), .A2(\SB2_3_3/i1_7 ), .A3(
        \SB2_3_3/i0[10] ), .ZN(\SB2_3_3/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U10338 ( .A1(\SB2_3_3/i0_4 ), .A2(\SB2_3_3/i0_3 ), .A3(
        \SB2_3_3/i1[9] ), .ZN(\SB2_3_3/Component_Function_5/NAND4_in[2] ) );
  CLKBUF_X4 U10339 ( .I(\SB3_0/buf_output[2] ), .Z(\SB4_29/i0_0 ) );
  NAND3_X1 U10340 ( .A1(\SB4_1/i0_0 ), .A2(\SB4_1/i0_3 ), .A3(\SB4_1/i0_4 ), 
        .ZN(n6195) );
  NAND3_X1 U10343 ( .A1(\SB3_12/i1[9] ), .A2(\SB3_12/i0_4 ), .A3(\SB3_12/i0_3 ), .ZN(\SB3_12/Component_Function_5/NAND4_in[2] ) );
  NAND2_X1 U10344 ( .A1(\SB3_12/i0_3 ), .A2(\SB3_12/i1[9] ), .ZN(
        \SB3_12/Component_Function_1/NAND4_in[0] ) );
  NAND3_X1 U10345 ( .A1(\SB3_12/i0[10] ), .A2(\SB3_12/i0_3 ), .A3(
        \SB3_12/i0[9] ), .ZN(\SB3_12/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U10347 ( .A1(\SB4_20/i1[9] ), .A2(n3674), .A3(\SB4_20/i0_4 ), .ZN(
        \SB4_20/Component_Function_4/NAND4_in[3] ) );
  CLKBUF_X4 U10349 ( .I(\SB2_0_16/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_0/buf_datainput[105] ) );
  INV_X1 U10351 ( .I(\MC_ARK_ARC_1_3/buf_output[91] ), .ZN(\SB3_16/i1_7 ) );
  BUF_X2 U10353 ( .I(\MC_ARK_ARC_1_3/buf_output[91] ), .Z(\SB3_16/i0[6] ) );
  INV_X1 U10355 ( .I(n418), .ZN(\SB1_0_18/i1_5 ) );
  NAND3_X1 U10361 ( .A1(\SB2_2_19/i0[9] ), .A2(\SB1_2_23/buf_output[1] ), .A3(
        \SB1_2_20/buf_output[4] ), .ZN(
        \SB2_2_19/Component_Function_5/NAND4_in[3] ) );
  CLKBUF_X4 U10362 ( .I(\SB3_7/buf_output[3] ), .Z(\SB4_5/i0[10] ) );
  AND4_X2 U10366 ( .A1(\SB1_3_2/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_3_2/Component_Function_3/NAND4_in[0] ), .A3(n1658), .A4(n4563), 
        .Z(n5513) );
  AND4_X2 U10367 ( .A1(\SB3_31/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_31/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_31/Component_Function_2/NAND4_in[2] ), .A4(
        \SB3_31/Component_Function_2/NAND4_in[3] ), .Z(n5514) );
  NAND3_X1 U10369 ( .A1(\SB2_3_27/i0[7] ), .A2(\SB2_3_27/i0_3 ), .A3(
        \SB2_3_27/i0_0 ), .ZN(\SB2_3_27/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 U10372 ( .A1(\SB2_3_27/i0_0 ), .A2(\SB2_3_27/i3[0] ), .ZN(
        \SB2_3_27/Component_Function_5/NAND4_in[0] ) );
  BUF_X2 U10376 ( .I(\MC_ARK_ARC_1_2/buf_output[6] ), .Z(\SB1_3_30/i0[9] ) );
  XOR2_X1 U10377 ( .A1(n4454), .A2(n3176), .Z(n5516) );
  CLKBUF_X4 U10378 ( .I(\MC_ARK_ARC_1_2/buf_output[112] ), .Z(\SB1_3_13/i0_4 )
         );
  NAND3_X1 U10379 ( .A1(\SB1_1_31/i0_0 ), .A2(\SB1_1_31/i0[6] ), .A3(
        \SB1_1_31/i0[10] ), .ZN(\SB1_1_31/Component_Function_5/NAND4_in[1] )
         );
  XOR2_X1 U10381 ( .A1(Key[134]), .A2(Plaintext[134]), .Z(n5517) );
  AND4_X2 U10390 ( .A1(\SB1_0_9/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_9/Component_Function_5/NAND4_in[3] ), .A3(n1812), .A4(
        \SB1_0_9/Component_Function_5/NAND4_in[0] ), .Z(n5518) );
  NAND3_X1 U10391 ( .A1(\SB2_2_22/i0_0 ), .A2(\SB2_2_22/i1_5 ), .A3(
        \SB2_2_22/i0_4 ), .ZN(n4568) );
  NAND3_X1 U10392 ( .A1(\SB2_2_22/i3[0] ), .A2(\SB2_2_22/i0_0 ), .A3(
        \SB2_2_22/i1_7 ), .ZN(\SB2_2_22/Component_Function_4/NAND4_in[1] ) );
  NAND3_X1 U10394 ( .A1(\SB2_2_22/i0[7] ), .A2(\SB2_2_22/i0_3 ), .A3(
        \SB2_2_22/i0_0 ), .ZN(\SB2_2_22/Component_Function_0/NAND4_in[3] ) );
  INV_X1 U10397 ( .I(n429), .ZN(\SB1_0_7/i1_5 ) );
  NAND3_X1 U10398 ( .A1(\SB3_30/i1[9] ), .A2(\SB3_30/i0[6] ), .A3(n5509), .ZN(
        n3451) );
  INV_X1 U10399 ( .I(\RI3[0][131] ), .ZN(\SB2_0_10/i1_5 ) );
  INV_X1 U10400 ( .I(\SB3_22/buf_output[5] ), .ZN(\SB4_22/i1_5 ) );
  BUF_X2 U10401 ( .I(\MC_ARK_ARC_1_1/buf_output[150] ), .Z(\SB1_2_6/i0[9] ) );
  INV_X1 U10402 ( .I(\MC_ARK_ARC_1_1/buf_output[150] ), .ZN(\SB1_2_6/i3[0] )
         );
  CLKBUF_X4 U10403 ( .I(\SB3_30/buf_output[0] ), .Z(\SB4_25/i0[9] ) );
  NAND3_X1 U10406 ( .A1(\SB2_2_20/i0[7] ), .A2(\SB2_2_20/i0_3 ), .A3(
        \SB2_2_20/i0_0 ), .ZN(\SB2_2_20/Component_Function_0/NAND4_in[3] ) );
  NAND2_X1 U10412 ( .A1(\SB2_2_20/i0_0 ), .A2(\SB2_2_20/i3[0] ), .ZN(
        \SB2_2_20/Component_Function_5/NAND4_in[0] ) );
  CLKBUF_X4 U10417 ( .I(\SB1_2_23/buf_output[2] ), .Z(\SB2_2_20/i0_0 ) );
  BUF_X4 U10422 ( .I(\SB2_1_23/buf_output[3] ), .Z(
        \MC_ARK_ARC_1_1/buf_datainput[63] ) );
  NAND3_X1 U10424 ( .A1(\SB1_2_20/i0_4 ), .A2(n2909), .A3(\SB1_2_20/i1[9] ), 
        .ZN(\SB1_2_20/Component_Function_4/NAND4_in[3] ) );
  AND4_X2 U10428 ( .A1(\SB1_3_4/Component_Function_5/NAND4_in[2] ), .A2(n2284), 
        .A3(\SB1_3_4/Component_Function_5/NAND4_in[3] ), .A4(n2054), .Z(n5519)
         );
  NAND4_X1 U10430 ( .A1(\SB3_1/Component_Function_2/NAND4_in[1] ), .A2(
        \SB3_1/Component_Function_2/NAND4_in[2] ), .A3(
        \SB3_1/Component_Function_2/NAND4_in[0] ), .A4(n4092), .ZN(
        \SB3_1/buf_output[2] ) );
  INV_X1 U10432 ( .I(\SB1_2_29/buf_output[1] ), .ZN(\SB2_2_25/i1_7 ) );
  CLKBUF_X4 U10438 ( .I(\MC_ARK_ARC_1_1/buf_output[12] ), .Z(\SB1_2_29/i0[9] )
         );
  CLKBUF_X4 U10439 ( .I(\MC_ARK_ARC_1_0/buf_output[113] ), .Z(\SB1_1_13/i0_3 )
         );
  INV_X1 U10441 ( .I(\MC_ARK_ARC_1_0/buf_output[113] ), .ZN(\SB1_1_13/i1_5 )
         );
  CLKBUF_X4 U10444 ( .I(\SB1_1_13/buf_output[3] ), .Z(\SB2_1_11/i0[10] ) );
  CLKBUF_X4 U10446 ( .I(\MC_ARK_ARC_1_2/buf_output[44] ), .Z(\SB1_3_24/i0_0 )
         );
  CLKBUF_X4 U10447 ( .I(\RI1[4][87] ), .Z(\SB3_17/i0[10] ) );
  CLKBUF_X4 U10448 ( .I(\MC_ARK_ARC_1_1/buf_output[51] ), .Z(\SB1_2_23/i0[10] ) );
  XOR2_X1 U10450 ( .A1(n2820), .A2(\MC_ARK_ARC_1_3/temp6[63] ), .Z(n5520) );
  BUF_X2 U10451 ( .I(\SB3_30/buf_output[1] ), .Z(\SB4_26/i0[6] ) );
  CLKBUF_X4 U10453 ( .I(\RI3[0][32] ), .Z(\SB2_0_26/i0_0 ) );
  NAND3_X1 U10455 ( .A1(\SB3_0/i0_0 ), .A2(\SB3_0/i0_3 ), .A3(\SB3_0/i0_4 ), 
        .ZN(\SB3_0/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U10456 ( .A1(\SB3_0/i0[9] ), .A2(\SB3_0/i0[10] ), .A3(\SB3_0/i0_3 ), 
        .ZN(\SB3_0/Component_Function_4/NAND4_in[2] ) );
  NAND3_X1 U10457 ( .A1(\SB3_0/i0_4 ), .A2(\SB3_0/i0_3 ), .A3(\SB3_0/i1[9] ), 
        .ZN(n4617) );
  CLKBUF_X4 U10461 ( .I(\MC_ARK_ARC_1_2/buf_output[50] ), .Z(\SB1_3_23/i0_0 )
         );
  CLKBUF_X4 U10463 ( .I(\MC_ARK_ARC_1_3/buf_output[134] ), .Z(\SB3_9/i0_0 ) );
  CLKBUF_X4 U10472 ( .I(\MC_ARK_ARC_1_0/buf_output[56] ), .Z(\SB1_1_22/i0_0 )
         );
  NAND3_X1 U10473 ( .A1(\RI1[1][59] ), .A2(\SB1_1_22/i1[9] ), .A3(
        \SB1_1_22/i0[6] ), .ZN(\SB1_1_22/Component_Function_3/NAND4_in[0] ) );
  NAND2_X2 U10479 ( .A1(n3913), .A2(n4760), .ZN(n5521) );
  XOR2_X1 U10480 ( .A1(n4553), .A2(\MC_ARK_ARC_1_1/temp5[153] ), .Z(n5522) );
  NAND3_X1 U10482 ( .A1(\SB1_0_8/i0_3 ), .A2(\SB1_0_8/i0_0 ), .A3(
        \SB1_0_8/i0[7] ), .ZN(\SB1_0_8/Component_Function_0/NAND4_in[3] ) );
  NAND3_X1 U10484 ( .A1(\SB1_0_8/i0[10] ), .A2(\SB1_0_8/i0_4 ), .A3(
        \SB1_0_8/i0_3 ), .ZN(\SB1_0_8/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U10485 ( .A1(\SB1_0_8/i0_3 ), .A2(\SB1_0_8/i0[6] ), .A3(
        \SB1_0_8/i1[9] ), .ZN(\SB1_0_8/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U10486 ( .A1(\SB1_0_8/i0_3 ), .A2(\SB1_0_8/i0[8] ), .A3(
        \SB1_0_8/i0[9] ), .ZN(\SB1_0_8/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U10492 ( .A1(\SB1_0_8/i0_3 ), .A2(\SB1_0_8/i0[10] ), .A3(
        \SB1_0_8/i0[9] ), .ZN(\SB1_0_8/Component_Function_4/NAND4_in[2] ) );
  NAND3_X2 U10493 ( .A1(\SB1_3_1/i0_3 ), .A2(\SB1_3_1/i0[10] ), .A3(
        \SB1_3_1/i0[6] ), .ZN(\SB1_3_1/Component_Function_2/NAND4_in[1] ) );
  XOR2_X1 U10494 ( .A1(n1146), .A2(\MC_ARK_ARC_1_1/temp5[86] ), .Z(n5523) );
  NAND3_X1 U10496 ( .A1(\SB3_31/i0_4 ), .A2(\SB3_31/i0[8] ), .A3(\SB3_31/i1_7 ), .ZN(\SB3_31/Component_Function_1/NAND4_in[3] ) );
  NAND3_X1 U10502 ( .A1(\SB3_31/i0_3 ), .A2(\SB3_31/i1_7 ), .A3(\SB3_31/i0[8] ), .ZN(\SB3_31/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U10504 ( .A1(\MC_ARK_ARC_1_2/temp6[86] ), .A2(
        \MC_ARK_ARC_1_2/temp5[86] ), .Z(n5524) );
  CLKBUF_X4 U10507 ( .I(\SB3_21/buf_output[2] ), .Z(\SB4_18/i0_0 ) );
  CLKBUF_X4 U10512 ( .I(\SB1_3_27/buf_output[2] ), .Z(\SB2_3_24/i0_0 ) );
  XOR2_X1 U10514 ( .A1(n6327), .A2(n5917), .Z(n5526) );
  XOR2_X1 U10515 ( .A1(\MC_ARK_ARC_1_2/temp6[80] ), .A2(
        \MC_ARK_ARC_1_2/temp5[80] ), .Z(n5527) );
  INV_X1 U10516 ( .I(\MC_ARK_ARC_1_1/buf_output[19] ), .ZN(\SB1_2_28/i1_7 ) );
  BUF_X2 U10524 ( .I(\MC_ARK_ARC_1_1/buf_output[19] ), .Z(\SB1_2_28/i0[6] ) );
  BUF_X2 U10525 ( .I(\MC_ARK_ARC_1_0/buf_output[50] ), .Z(\SB1_1_23/i0_0 ) );
  BUF_X2 U10529 ( .I(\MC_ARK_ARC_1_2/buf_output[25] ), .Z(\SB1_3_27/i0[6] ) );
  INV_X1 U10535 ( .I(\MC_ARK_ARC_1_2/buf_output[25] ), .ZN(\SB1_3_27/i1_7 ) );
  CLKBUF_X4 U10536 ( .I(\MC_ARK_ARC_1_0/buf_output[116] ), .Z(\SB1_1_12/i0_0 )
         );
  NAND4_X2 U10542 ( .A1(n4202), .A2(
        \SB2_2_20/Component_Function_2/NAND4_in[0] ), .A3(n5736), .A4(
        \SB2_2_20/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB2_2_20/buf_output[2] ) );
  XOR2_X1 U10545 ( .A1(\RI5[1][76] ), .A2(\RI5[1][70] ), .Z(
        \MC_ARK_ARC_1_1/temp1[76] ) );
  NAND4_X2 U10546 ( .A1(n4528), .A2(
        \SB2_1_10/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_1_10/Component_Function_0/NAND4_in[3] ), .A4(n5528), .ZN(
        \SB2_1_10/buf_output[0] ) );
  NAND2_X1 U10548 ( .A1(\SB2_1_10/i0[10] ), .A2(\SB2_1_10/i0[9] ), .ZN(n5528)
         );
  NAND3_X1 U10549 ( .A1(\SB3_4/i0[10] ), .A2(\SB3_4/i0_3 ), .A3(\SB3_4/i0_4 ), 
        .ZN(\SB3_4/Component_Function_0/NAND4_in[2] ) );
  NAND4_X2 U10553 ( .A1(\SB4_15/Component_Function_2/NAND4_in[0] ), .A2(n1867), 
        .A3(\SB4_15/Component_Function_2/NAND4_in[1] ), .A4(n3248), .ZN(n6344)
         );
  NAND4_X2 U10557 ( .A1(n3968), .A2(\SB3_0/Component_Function_2/NAND4_in[3] ), 
        .A3(n675), .A4(n6378), .ZN(\SB3_0/buf_output[2] ) );
  NAND4_X2 U10563 ( .A1(\SB3_4/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_4/Component_Function_3/NAND4_in[1] ), .A3(n5978), .A4(n6278), 
        .ZN(\SB3_4/buf_output[3] ) );
  XOR2_X1 U10565 ( .A1(\RI5[1][156] ), .A2(\RI5[1][108] ), .Z(n6423) );
  NAND3_X1 U10566 ( .A1(\SB4_16/i0_0 ), .A2(\SB4_16/i0_4 ), .A3(\SB4_16/i1_5 ), 
        .ZN(\SB4_16/Component_Function_2/NAND4_in[3] ) );
  NAND4_X2 U10568 ( .A1(\SB4_14/Component_Function_5/NAND4_in[2] ), .A2(n2572), 
        .A3(\SB4_14/Component_Function_5/NAND4_in[0] ), .A4(
        \SB4_14/Component_Function_5/NAND4_in[1] ), .ZN(n3988) );
  XOR2_X1 U10569 ( .A1(\RI5[3][83] ), .A2(\RI5[3][89] ), .Z(
        \MC_ARK_ARC_1_3/temp1[89] ) );
  XOR2_X1 U10570 ( .A1(\RI5[3][85] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[91] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[91] ) );
  XOR2_X1 U10572 ( .A1(\SB2_1_22/buf_output[2] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[38] ), .Z(\MC_ARK_ARC_1_1/temp3[164] )
         );
  NAND3_X2 U10575 ( .A1(\SB2_3_18/i0[6] ), .A2(\SB2_3_18/i0[9] ), .A3(
        \SB2_3_18/i0_4 ), .ZN(n4692) );
  XOR2_X1 U10578 ( .A1(n5529), .A2(n231), .Z(Ciphertext[190]) );
  NAND4_X2 U10580 ( .A1(n5767), .A2(\SB4_0/Component_Function_4/NAND4_in[2] ), 
        .A3(n2658), .A4(\SB4_0/Component_Function_4/NAND4_in[0] ), .ZN(n5529)
         );
  NAND4_X2 U10581 ( .A1(\SB1_3_22/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_3_22/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_3_22/Component_Function_1/NAND4_in[0] ), .A4(
        \SB1_3_22/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_3_22/buf_output[1] ) );
  NAND4_X2 U10582 ( .A1(\SB1_1_12/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_12/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_1_12/Component_Function_1/NAND4_in[3] ), .A4(
        \SB1_1_12/Component_Function_1/NAND4_in[1] ), .ZN(
        \SB1_1_12/buf_output[1] ) );
  NAND4_X2 U10583 ( .A1(\SB2_0_16/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_0_16/Component_Function_5/NAND4_in[0] ), .A3(n3819), .A4(n5530), 
        .ZN(\SB2_0_16/buf_output[5] ) );
  INV_X2 U10584 ( .I(\SB3_16/buf_output[2] ), .ZN(\SB4_13/i1[9] ) );
  NAND4_X2 U10585 ( .A1(n6397), .A2(
        \SB1_3_17/Component_Function_4/NAND4_in[1] ), .A3(n6306), .A4(n5531), 
        .ZN(\SB1_3_17/buf_output[4] ) );
  NAND3_X2 U10586 ( .A1(\SB1_3_17/i0_0 ), .A2(\SB1_3_17/i0[9] ), .A3(
        \SB1_3_17/i0[8] ), .ZN(n5531) );
  NAND4_X2 U10588 ( .A1(\SB2_3_21/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_3_21/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_3_21/Component_Function_4/NAND4_in[1] ), .A4(n5532), .ZN(
        \SB2_3_21/buf_output[4] ) );
  NAND3_X1 U10589 ( .A1(\SB2_3_21/i1[9] ), .A2(\SB2_3_21/i1_5 ), .A3(
        \SB1_3_22/buf_output[4] ), .ZN(n5532) );
  NAND3_X1 U10597 ( .A1(\SB3_14/i0[10] ), .A2(\SB3_14/i1_5 ), .A3(
        \SB3_14/i1[9] ), .ZN(\SB3_14/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U10599 ( .A1(n5533), .A2(n240), .Z(Ciphertext[94]) );
  XOR2_X1 U10603 ( .A1(n5534), .A2(n177), .Z(Ciphertext[122]) );
  NAND4_X2 U10604 ( .A1(n2686), .A2(n2635), .A3(
        \SB4_11/Component_Function_2/NAND4_in[3] ), .A4(
        \SB4_11/Component_Function_2/NAND4_in[2] ), .ZN(n5534) );
  NAND3_X1 U10607 ( .A1(\SB4_12/i0[10] ), .A2(\SB4_12/i0_3 ), .A3(
        \SB3_17/buf_output[0] ), .ZN(n5535) );
  XOR2_X1 U10608 ( .A1(n4214), .A2(n5536), .Z(\MC_ARK_ARC_1_3/buf_output[105] ) );
  XOR2_X1 U10612 ( .A1(n4392), .A2(n6307), .Z(n5536) );
  XOR2_X1 U10616 ( .A1(n5538), .A2(n131), .Z(Ciphertext[119]) );
  NAND4_X2 U10617 ( .A1(\SB4_12/Component_Function_5/NAND4_in[3] ), .A2(
        \SB4_12/Component_Function_5/NAND4_in[1] ), .A3(n2518), .A4(n3203), 
        .ZN(n5538) );
  NAND4_X2 U10618 ( .A1(\SB2_3_0/Component_Function_2/NAND4_in[2] ), .A2(n2300), .A3(n6214), .A4(n5540), .ZN(\SB2_3_0/buf_output[2] ) );
  NAND3_X2 U10631 ( .A1(\SB2_3_0/i0_3 ), .A2(\SB2_3_0/i0[6] ), .A3(
        \SB2_3_0/i0[10] ), .ZN(n5540) );
  NAND4_X2 U10632 ( .A1(\SB2_3_31/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_3_31/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_3_31/Component_Function_2/NAND4_in[1] ), .A4(n5541), .ZN(
        \SB2_3_31/buf_output[2] ) );
  XOR2_X1 U10633 ( .A1(\MC_ARK_ARC_1_2/temp2[191] ), .A2(n2967), .Z(n5543) );
  NOR2_X2 U10641 ( .A1(n1048), .A2(n5544), .ZN(\SB2_0_28/i0[7] ) );
  NAND2_X2 U10642 ( .A1(n3092), .A2(
        \SB1_0_29/Component_Function_4/NAND4_in[1] ), .ZN(n5544) );
  XOR2_X1 U10643 ( .A1(n5545), .A2(n66), .Z(Ciphertext[117]) );
  NAND4_X2 U10644 ( .A1(\SB4_12/Component_Function_3/NAND4_in[3] ), .A2(n2465), 
        .A3(n965), .A4(n6515), .ZN(n5545) );
  XOR2_X1 U10649 ( .A1(n5546), .A2(\MC_ARK_ARC_1_3/temp6[57] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[57] ) );
  XOR2_X1 U10650 ( .A1(\MC_ARK_ARC_1_3/temp1[57] ), .A2(
        \MC_ARK_ARC_1_3/temp2[57] ), .Z(n5546) );
  NAND4_X2 U10656 ( .A1(\SB3_13/Component_Function_4/NAND4_in[1] ), .A2(
        \SB3_13/Component_Function_4/NAND4_in[2] ), .A3(n2600), .A4(n5547), 
        .ZN(\SB3_13/buf_output[4] ) );
  NAND3_X1 U10658 ( .A1(\SB3_13/i0[9] ), .A2(\SB3_13/i0[8] ), .A3(
        \MC_ARK_ARC_1_3/buf_output[110] ), .ZN(n5547) );
  XOR2_X1 U10659 ( .A1(n5808), .A2(n5548), .Z(\MC_ARK_ARC_1_1/temp5[140] ) );
  XOR2_X1 U10661 ( .A1(\RI5[1][134] ), .A2(\RI5[1][140] ), .Z(n5548) );
  INV_X2 U10663 ( .I(n5549), .ZN(n3913) );
  NAND2_X2 U10667 ( .A1(\SB2_1_9/Component_Function_3/NAND4_in[3] ), .A2(n5710), .ZN(n5549) );
  NAND4_X2 U10669 ( .A1(\SB2_2_27/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_2_27/Component_Function_4/NAND4_in[3] ), .A3(n3775), .A4(n6121), 
        .ZN(\SB2_2_27/buf_output[4] ) );
  XOR2_X1 U10676 ( .A1(n701), .A2(n700), .Z(\RI1[3][167] ) );
  NAND4_X2 U10677 ( .A1(\SB2_3_27/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_3_27/Component_Function_2/NAND4_in[0] ), .A3(n5703), .A4(n4598), 
        .ZN(\SB2_3_27/buf_output[2] ) );
  INV_X2 U10687 ( .I(\SB1_3_11/buf_output[3] ), .ZN(\SB2_3_9/i0[8] ) );
  NAND4_X2 U10690 ( .A1(n4377), .A2(
        \SB1_3_11/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_3_11/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_3_11/Component_Function_3/NAND4_in[0] ), .ZN(
        \SB1_3_11/buf_output[3] ) );
  NAND4_X2 U10691 ( .A1(\SB3_30/Component_Function_1/NAND4_in[1] ), .A2(
        \SB3_30/Component_Function_1/NAND4_in[2] ), .A3(n2101), .A4(
        \SB3_30/Component_Function_1/NAND4_in[0] ), .ZN(\SB3_30/buf_output[1] ) );
  NAND4_X2 U10693 ( .A1(n3283), .A2(
        \SB2_2_12/Component_Function_5/NAND4_in[1] ), .A3(n5802), .A4(
        \SB2_2_12/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_2_12/buf_output[5] ) );
  XOR2_X1 U10697 ( .A1(\MC_ARK_ARC_1_2/temp5[125] ), .A2(n3718), .Z(n5550) );
  XOR2_X1 U10701 ( .A1(\RI5[2][11] ), .A2(\RI5[2][17] ), .Z(
        \MC_ARK_ARC_1_2/temp1[17] ) );
  XOR2_X1 U10705 ( .A1(\MC_ARK_ARC_1_1/temp5[44] ), .A2(n4309), .Z(
        \MC_ARK_ARC_1_1/buf_output[44] ) );
  XOR2_X1 U10706 ( .A1(n1718), .A2(n5602), .Z(n2562) );
  NAND4_X2 U10707 ( .A1(\SB2_2_7/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_2_7/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_2_7/Component_Function_4/NAND4_in[0] ), .A4(n5551), .ZN(
        \SB2_2_7/buf_output[4] ) );
  NAND4_X2 U10708 ( .A1(\SB2_3_21/Component_Function_2/NAND4_in[0] ), .A2(
        n3440), .A3(n3185), .A4(n5552), .ZN(\SB2_3_21/buf_output[2] ) );
  NAND4_X2 U10709 ( .A1(\SB1_2_28/Component_Function_5/NAND4_in[1] ), .A2(
        n4652), .A3(\SB1_2_28/Component_Function_5/NAND4_in[0] ), .A4(n5553), 
        .ZN(\SB1_2_28/buf_output[5] ) );
  NAND3_X2 U10714 ( .A1(\SB1_2_28/i0[6] ), .A2(\SB1_2_28/i0[9] ), .A3(
        \SB1_2_28/i0_4 ), .ZN(n5553) );
  NAND3_X1 U10717 ( .A1(\SB4_6/i0[10] ), .A2(\SB4_6/i1_5 ), .A3(\SB4_6/i1[9] ), 
        .ZN(\SB4_6/Component_Function_2/NAND4_in[0] ) );
  NAND2_X2 U10719 ( .A1(n5840), .A2(n5841), .ZN(\SB4_6/i0[10] ) );
  XOR2_X1 U10723 ( .A1(\RI5[2][121] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[115] ), .Z(\MC_ARK_ARC_1_2/temp1[121] ) );
  INV_X2 U10726 ( .I(\RI3[0][32] ), .ZN(\SB2_0_26/i1[9] ) );
  NAND4_X2 U10729 ( .A1(n4095), .A2(n834), .A3(n5871), .A4(n4228), .ZN(
        \RI3[0][32] ) );
  NAND4_X2 U10733 ( .A1(n6528), .A2(
        \SB1_1_22/Component_Function_5/NAND4_in[3] ), .A3(n1044), .A4(n5554), 
        .ZN(\SB1_1_22/buf_output[5] ) );
  XOR2_X1 U10735 ( .A1(\MC_ARK_ARC_1_3/temp1[91] ), .A2(n5555), .Z(
        \MC_ARK_ARC_1_3/temp5[91] ) );
  XOR2_X1 U10741 ( .A1(\SB2_3_25/buf_output[1] ), .A2(\RI5[3][37] ), .Z(n5555)
         );
  NAND4_X2 U10744 ( .A1(\SB2_2_22/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_2_22/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_2_22/Component_Function_0/NAND4_in[0] ), .A4(n5556), .ZN(
        \SB2_2_22/buf_output[0] ) );
  NAND4_X2 U10745 ( .A1(\SB2_1_21/Component_Function_0/NAND4_in[1] ), .A2(
        n4697), .A3(\SB2_1_21/Component_Function_0/NAND4_in[3] ), .A4(n5557), 
        .ZN(\SB2_1_21/buf_output[0] ) );
  NAND2_X2 U10746 ( .A1(\SB2_1_21/i0[10] ), .A2(\RI3[1][60] ), .ZN(n5557) );
  NAND3_X1 U10749 ( .A1(\SB3_25/i0[10] ), .A2(\SB3_25/i0_0 ), .A3(
        \SB3_25/i0[6] ), .ZN(\SB3_25/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U10751 ( .A1(\SB3_2/i0[6] ), .A2(\SB3_2/i0[10] ), .A3(\SB3_2/i0_0 ), 
        .ZN(\SB3_2/Component_Function_5/NAND4_in[1] ) );
  NOR2_X2 U10752 ( .A1(n5559), .A2(n5558), .ZN(n6025) );
  NAND4_X2 U10753 ( .A1(n6009), .A2(
        \SB2_2_22/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_2_22/Component_Function_3/NAND4_in[1] ), .A4(n1820), .ZN(
        \SB2_2_22/buf_output[3] ) );
  NAND4_X2 U10758 ( .A1(\SB2_1_7/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_7/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_1_7/Component_Function_3/NAND4_in[3] ), .A4(n5560), .ZN(
        \SB2_1_7/buf_output[3] ) );
  NAND3_X2 U10759 ( .A1(\SB2_1_7/i0_3 ), .A2(\SB2_1_7/i0_0 ), .A3(n5790), .ZN(
        n5560) );
  XOR2_X1 U10764 ( .A1(n5561), .A2(n114), .Z(Ciphertext[7]) );
  NAND4_X2 U10766 ( .A1(\SB2_1_10/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_1_10/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_1_10/Component_Function_2/NAND4_in[0] ), .A4(n5562), .ZN(
        \SB2_1_10/buf_output[2] ) );
  NAND3_X2 U10775 ( .A1(\SB1_1_11/buf_output[4] ), .A2(\SB2_1_10/i0_0 ), .A3(
        \SB2_1_10/i1_5 ), .ZN(n5562) );
  NOR2_X2 U10776 ( .A1(n5564), .A2(n5563), .ZN(n1386) );
  NAND2_X1 U10777 ( .A1(n2108), .A2(\SB3_3/Component_Function_2/NAND4_in[0] ), 
        .ZN(n5564) );
  NAND4_X2 U10780 ( .A1(\SB2_3_7/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_3_7/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_3_7/Component_Function_1/NAND4_in[2] ), .A4(n5565), .ZN(
        \SB2_3_7/buf_output[1] ) );
  NAND3_X2 U10782 ( .A1(\SB1_3_5/i0[9] ), .A2(\SB1_3_5/i0[6] ), .A3(
        \SB1_3_5/i0_4 ), .ZN(n5566) );
  NAND4_X2 U10784 ( .A1(n959), .A2(n2171), .A3(
        \SB3_16/Component_Function_1/NAND4_in[0] ), .A4(n5567), .ZN(
        \SB3_16/buf_output[1] ) );
  NAND3_X1 U10788 ( .A1(\SB3_16/i0[6] ), .A2(\SB3_16/i0[9] ), .A3(
        \SB3_16/i1_5 ), .ZN(n5567) );
  NAND3_X1 U10789 ( .A1(\SB3_8/i0_0 ), .A2(\SB3_8/i3[0] ), .A3(\SB3_8/i1_7 ), 
        .ZN(\SB3_8/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U10790 ( .A1(n5568), .A2(n84), .Z(Ciphertext[114]) );
  NAND4_X2 U10791 ( .A1(\SB4_12/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_12/Component_Function_0/NAND4_in[1] ), .A3(n3388), .A4(n4515), 
        .ZN(n5568) );
  NAND4_X2 U10792 ( .A1(\SB3_8/Component_Function_1/NAND4_in[1] ), .A2(
        \SB3_8/Component_Function_1/NAND4_in[3] ), .A3(
        \SB3_8/Component_Function_1/NAND4_in[2] ), .A4(n5569), .ZN(
        \SB3_8/buf_output[1] ) );
  NAND2_X1 U10793 ( .A1(\SB3_8/i0_3 ), .A2(\SB3_8/i1[9] ), .ZN(n5569) );
  NAND3_X2 U10796 ( .A1(\SB2_3_4/i0[10] ), .A2(\SB2_3_4/i1[9] ), .A3(n5519), 
        .ZN(n6362) );
  NAND3_X1 U10803 ( .A1(\SB4_4/i0[6] ), .A2(\SB4_4/i0_3 ), .A3(n3655), .ZN(
        n5570) );
  XOR2_X1 U10804 ( .A1(\MC_ARK_ARC_1_2/temp1[156] ), .A2(n5571), .Z(n2186) );
  XOR2_X1 U10806 ( .A1(\RI5[2][126] ), .A2(\RI5[2][102] ), .Z(n5571) );
  NAND4_X2 U10809 ( .A1(n3450), .A2(n3058), .A3(n6279), .A4(
        \SB1_3_4/Component_Function_4/NAND4_in[0] ), .ZN(
        \SB1_3_4/buf_output[4] ) );
  NAND4_X2 U10810 ( .A1(\SB1_2_23/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_2_23/Component_Function_1/NAND4_in[2] ), .A3(n1594), .A4(
        \SB1_2_23/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_2_23/buf_output[1] ) );
  NAND4_X2 U10815 ( .A1(\SB2_0_14/Component_Function_0/NAND4_in[0] ), .A2(
        \SB2_0_14/Component_Function_0/NAND4_in[3] ), .A3(n5573), .A4(
        \SB2_0_14/Component_Function_0/NAND4_in[2] ), .ZN(
        \SB2_0_14/buf_output[0] ) );
  NAND3_X2 U10816 ( .A1(\SB2_0_14/i0[8] ), .A2(\SB2_0_14/i0[7] ), .A3(
        \SB2_0_14/i0[6] ), .ZN(n5573) );
  NAND3_X2 U10821 ( .A1(\SB2_2_21/i0[6] ), .A2(\SB2_2_21/i0[9] ), .A3(
        \SB2_2_21/i1_5 ), .ZN(\SB2_2_21/Component_Function_1/NAND4_in[2] ) );
  NAND3_X1 U10823 ( .A1(\SB4_16/i0_4 ), .A2(\SB4_16/i1[9] ), .A3(\SB4_16/i1_5 ), .ZN(n3861) );
  NAND3_X1 U10830 ( .A1(\SB2_2_11/i0[6] ), .A2(\SB2_2_11/i0_3 ), .A3(n5515), 
        .ZN(\SB2_2_11/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U10831 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[105] ), .A2(\RI5[2][135] ), .Z(n5574) );
  NAND4_X2 U10833 ( .A1(\SB2_1_10/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_1_10/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_1_10/Component_Function_1/NAND4_in[2] ), .A4(
        \SB2_1_10/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB2_1_10/buf_output[1] ) );
  NAND4_X2 U10835 ( .A1(\SB1_2_31/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_31/Component_Function_3/NAND4_in[2] ), .A3(n2689), .A4(n5575), 
        .ZN(\SB1_2_31/buf_output[3] ) );
  NAND3_X2 U10836 ( .A1(\SB1_2_31/i0_0 ), .A2(\SB1_2_31/i0_3 ), .A3(
        \SB1_2_31/i0_4 ), .ZN(n5575) );
  XOR2_X1 U10846 ( .A1(n4629), .A2(n5576), .Z(n2385) );
  XOR2_X1 U10847 ( .A1(\SB2_3_21/buf_output[5] ), .A2(\RI5[3][59] ), .Z(n5576)
         );
  NAND3_X2 U10850 ( .A1(\SB2_3_22/i0[6] ), .A2(\SB2_3_22/i0_4 ), .A3(
        \SB2_3_22/i0[9] ), .ZN(n5577) );
  NAND2_X1 U10853 ( .A1(\SB1_3_8/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_8/Component_Function_2/NAND4_in[1] ), .ZN(n3413) );
  AND2_X1 U10857 ( .A1(n3075), .A2(n1861), .Z(n2718) );
  XOR2_X1 U10859 ( .A1(\MC_ARK_ARC_1_2/temp6[140] ), .A2(n1928), .Z(
        \MC_ARK_ARC_1_2/buf_output[140] ) );
  NAND3_X2 U10860 ( .A1(\SB1_1_4/i0[10] ), .A2(\SB1_1_4/i0_3 ), .A3(
        \SB1_1_4/i0[9] ), .ZN(\SB1_1_4/Component_Function_4/NAND4_in[2] ) );
  XOR2_X1 U10861 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[122] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[86] ), .Z(n5578) );
  NAND3_X1 U10863 ( .A1(\SB2_2_6/i0_3 ), .A2(\SB2_2_6/i0[8] ), .A3(
        \SB2_2_6/i1_7 ), .ZN(\SB2_2_6/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U10868 ( .A1(\RI5[1][86] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[110] ), 
        .Z(n5808) );
  NAND4_X2 U10874 ( .A1(\SB1_1_2/Component_Function_3/NAND4_in[2] ), .A2(
        \SB1_1_2/Component_Function_3/NAND4_in[1] ), .A3(n6010), .A4(n4388), 
        .ZN(\SB1_1_2/buf_output[3] ) );
  XOR2_X1 U10882 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[175] ), .A2(\RI5[2][169] ), .Z(\MC_ARK_ARC_1_2/temp1[175] ) );
  OR2_X2 U10885 ( .A1(n5789), .A2(n599), .Z(\SB2_0_5/i0_0 ) );
  XOR2_X1 U10891 ( .A1(n3540), .A2(n5579), .Z(\MC_ARK_ARC_1_1/buf_output[188] ) );
  XOR2_X1 U10895 ( .A1(n5580), .A2(n58), .Z(Ciphertext[154]) );
  NAND4_X2 U10897 ( .A1(\SB4_6/Component_Function_4/NAND4_in[0] ), .A2(
        \SB4_6/Component_Function_4/NAND4_in[3] ), .A3(n5817), .A4(
        \SB4_6/Component_Function_4/NAND4_in[2] ), .ZN(n5580) );
  NAND3_X2 U10898 ( .A1(\SB4_5/i0_0 ), .A2(\SB4_5/i0_4 ), .A3(\SB4_5/i0_3 ), 
        .ZN(n5581) );
  XOR2_X1 U10901 ( .A1(n5583), .A2(n5582), .Z(\MC_ARK_ARC_1_2/buf_output[98] )
         );
  XOR2_X1 U10911 ( .A1(n3166), .A2(n5626), .Z(n5582) );
  NAND4_X2 U10915 ( .A1(\SB2_1_3/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_1_3/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_1_3/Component_Function_0/NAND4_in[0] ), .A4(n5584), .ZN(
        \SB2_1_3/buf_output[0] ) );
  XOR2_X1 U10916 ( .A1(\RI5[0][153] ), .A2(\RI5[0][129] ), .Z(n5585) );
  NAND4_X2 U10920 ( .A1(\SB2_1_19/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_1_19/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_1_19/Component_Function_1/NAND4_in[0] ), .A4(n5586), .ZN(
        \SB2_1_19/buf_output[1] ) );
  NAND3_X2 U10924 ( .A1(\SB2_1_19/i0[6] ), .A2(\SB2_1_19/i0[9] ), .A3(
        \SB2_1_19/i1_5 ), .ZN(n5586) );
  AND2_X1 U10925 ( .A1(\SB1_1_4/Component_Function_4/NAND4_in[2] ), .A2(n2584), 
        .Z(n6539) );
  NAND4_X2 U10926 ( .A1(\SB2_2_31/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_31/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_2_31/Component_Function_4/NAND4_in[3] ), .A4(n5587), .ZN(
        \SB2_2_31/buf_output[4] ) );
  NAND3_X2 U10931 ( .A1(\SB2_2_31/i0[9] ), .A2(\SB2_2_31/i0_3 ), .A3(
        \SB2_2_31/i0[10] ), .ZN(n5587) );
  NAND3_X1 U10933 ( .A1(\SB3_31/i0[9] ), .A2(\SB3_31/i0_3 ), .A3(
        \SB3_31/i0[10] ), .ZN(\SB3_31/Component_Function_4/NAND4_in[2] ) );
  XOR2_X1 U10938 ( .A1(n5588), .A2(n5737), .Z(n5874) );
  XOR2_X1 U10939 ( .A1(\RI5[0][188] ), .A2(\RI5[0][116] ), .Z(n5588) );
  XOR2_X1 U10940 ( .A1(\MC_ARK_ARC_1_1/temp4[4] ), .A2(n5590), .Z(
        \MC_ARK_ARC_1_1/temp6[4] ) );
  XOR2_X1 U10943 ( .A1(\RI5[1][70] ), .A2(\RI5[1][106] ), .Z(n5590) );
  XOR2_X1 U10944 ( .A1(n5591), .A2(n3799), .Z(n4073) );
  NAND4_X2 U10945 ( .A1(\SB3_8/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_8/Component_Function_2/NAND4_in[2] ), .A3(
        \SB3_8/Component_Function_2/NAND4_in[1] ), .A4(
        \SB3_8/Component_Function_2/NAND4_in[3] ), .ZN(\SB3_8/buf_output[2] )
         );
  NAND4_X2 U10946 ( .A1(\SB1_1_17/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_1_17/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_1_17/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_1_17/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_1_17/buf_output[0] ) );
  NAND4_X2 U10947 ( .A1(n2015), .A2(
        \SB2_0_26/Component_Function_5/NAND4_in[3] ), .A3(n5872), .A4(n1795), 
        .ZN(\SB2_0_26/buf_output[5] ) );
  INV_X8 U10948 ( .I(n5592), .ZN(\RI1[2][17] ) );
  INV_X2 U10949 ( .I(\MC_ARK_ARC_1_1/buf_output[17] ), .ZN(n5592) );
  NAND4_X2 U10952 ( .A1(\SB3_25/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_25/Component_Function_2/NAND4_in[2] ), .A3(n5596), .A4(n5642), 
        .ZN(\SB3_25/buf_output[2] ) );
  NAND4_X2 U10953 ( .A1(\SB2_2_16/Component_Function_0/NAND4_in[1] ), .A2(
        n5719), .A3(n2650), .A4(\SB2_2_16/Component_Function_0/NAND4_in[0] ), 
        .ZN(\SB2_2_16/buf_output[0] ) );
  NAND3_X1 U10954 ( .A1(\SB1_3_7/i0_0 ), .A2(\SB1_3_7/i0_4 ), .A3(
        \SB1_3_7/i0_3 ), .ZN(\SB1_3_7/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U10955 ( .A1(\SB4_2/i0[10] ), .A2(\SB4_2/i0_3 ), .A3(\SB4_2/i0[9] ), 
        .ZN(n5593) );
  NAND4_X1 U10956 ( .A1(\SB2_0_25/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_0_25/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_0_25/Component_Function_4/NAND4_in[2] ), .A4(n5594), .ZN(
        \SB2_0_25/buf_output[4] ) );
  NAND3_X2 U10957 ( .A1(\SB2_0_25/i0_0 ), .A2(\SB2_0_25/i3[0] ), .A3(
        \SB2_0_25/i1_7 ), .ZN(n5594) );
  XOR2_X1 U10962 ( .A1(\MC_ARK_ARC_1_3/temp2[165] ), .A2(n5595), .Z(
        \MC_ARK_ARC_1_3/temp5[165] ) );
  XOR2_X1 U10963 ( .A1(\RI5[3][159] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[165] ), .Z(n5595) );
  INV_X2 U10966 ( .I(\SB1_3_19/buf_output[2] ), .ZN(\SB2_3_16/i1[9] ) );
  NAND4_X2 U10968 ( .A1(\SB1_3_19/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_19/Component_Function_2/NAND4_in[2] ), .A3(
        \SB1_3_19/Component_Function_2/NAND4_in[0] ), .A4(n2301), .ZN(
        \SB1_3_19/buf_output[2] ) );
  NAND3_X2 U10969 ( .A1(\SB2_1_21/i0[10] ), .A2(\SB2_1_21/i0_3 ), .A3(
        \SB2_1_21/i0[6] ), .ZN(n6283) );
  NAND3_X2 U10974 ( .A1(\SB2_3_30/i0_4 ), .A2(\SB2_3_30/i1[9] ), .A3(
        \SB2_3_30/i0_3 ), .ZN(n2387) );
  XOR2_X1 U10975 ( .A1(n6410), .A2(\MC_ARK_ARC_1_0/temp4[74] ), .Z(
        \MC_ARK_ARC_1_0/temp6[74] ) );
  NAND4_X2 U10977 ( .A1(n1436), .A2(n5692), .A3(
        \SB2_1_9/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_1_9/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_1_9/buf_output[5] ) );
  NAND3_X2 U10979 ( .A1(\SB3_25/i0[10] ), .A2(\SB3_25/i0_3 ), .A3(
        \SB3_25/i0[6] ), .ZN(n5596) );
  XOR2_X1 U10980 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[80] ), .A2(\RI5[1][44] ), 
        .Z(n5895) );
  XOR2_X1 U10984 ( .A1(\RI5[0][158] ), .A2(\RI5[0][182] ), .Z(
        \MC_ARK_ARC_1_0/temp2[20] ) );
  XOR2_X1 U10986 ( .A1(n3737), .A2(\MC_ARK_ARC_1_2/temp5[121] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[121] ) );
  XOR2_X1 U10988 ( .A1(\MC_ARK_ARC_1_1/temp2[107] ), .A2(n3903), .Z(
        \MC_ARK_ARC_1_1/temp5[107] ) );
  XOR2_X1 U10991 ( .A1(\RI5[3][184] ), .A2(\RI5[3][148] ), .Z(
        \MC_ARK_ARC_1_3/temp3[82] ) );
  XOR2_X1 U10993 ( .A1(\RI5[2][87] ), .A2(\RI5[2][93] ), .Z(n3105) );
  NAND3_X2 U11000 ( .A1(\SB2_2_19/i0[6] ), .A2(\SB2_2_19/i1[9] ), .A3(
        \SB2_2_19/i0_3 ), .ZN(\SB2_2_19/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U11001 ( .A1(\RI5[2][173] ), .A2(\RI5[2][179] ), .Z(
        \MC_ARK_ARC_1_2/temp1[179] ) );
  NAND4_X2 U11002 ( .A1(\SB2_2_3/Component_Function_5/NAND4_in[2] ), .A2(n2757), .A3(\SB2_2_3/Component_Function_5/NAND4_in[1] ), .A4(
        \SB2_2_3/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_2_3/buf_output[5] ) );
  XOR2_X1 U11004 ( .A1(n5598), .A2(n5597), .Z(n700) );
  XOR2_X1 U11007 ( .A1(\RI5[2][41] ), .A2(n459), .Z(n5597) );
  XOR2_X1 U11008 ( .A1(\RI5[2][77] ), .A2(\RI5[2][11] ), .Z(n5598) );
  NAND3_X2 U11009 ( .A1(\SB3_17/i0[6] ), .A2(\SB3_17/i0[10] ), .A3(
        \SB3_17/i0_3 ), .ZN(n5599) );
  AND2_X1 U11011 ( .A1(\SB2_3_19/Component_Function_0/NAND4_in[0] ), .A2(n1271), .Z(n5755) );
  NAND4_X2 U11012 ( .A1(\SB3_13/Component_Function_5/NAND4_in[1] ), .A2(n6254), 
        .A3(\SB3_13/Component_Function_5/NAND4_in[2] ), .A4(n5600), .ZN(
        \SB3_13/buf_output[5] ) );
  NAND3_X2 U11016 ( .A1(\SB3_13/i0[9] ), .A2(\SB3_13/i0[6] ), .A3(
        \SB3_13/i0_4 ), .ZN(n5600) );
  XOR2_X1 U11019 ( .A1(n5601), .A2(n104), .Z(Ciphertext[106]) );
  NAND4_X2 U11021 ( .A1(\SB4_14/Component_Function_4/NAND4_in[2] ), .A2(
        \SB4_14/Component_Function_4/NAND4_in[0] ), .A3(n1302), .A4(
        \SB4_14/Component_Function_4/NAND4_in[3] ), .ZN(n5601) );
  XOR2_X1 U11027 ( .A1(\RI5[3][164] ), .A2(\RI5[3][170] ), .Z(n5602) );
  NAND4_X2 U11044 ( .A1(\SB1_3_31/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_3_31/Component_Function_0/NAND4_in[1] ), .A3(n3555), .A4(n5603), 
        .ZN(\SB1_3_31/buf_output[0] ) );
  NAND2_X1 U11051 ( .A1(\SB1_3_31/i0[9] ), .A2(\SB1_3_31/i0[10] ), .ZN(n5603)
         );
  NAND3_X1 U11052 ( .A1(\RI3[0][155] ), .A2(\SB2_0_6/i0[7] ), .A3(
        \SB2_0_6/i0_0 ), .ZN(\SB2_0_6/Component_Function_0/NAND4_in[3] ) );
  XOR2_X1 U11054 ( .A1(n5604), .A2(n118), .Z(Ciphertext[52]) );
  XOR2_X1 U11055 ( .A1(\RI5[2][66] ), .A2(\RI5[2][90] ), .Z(n5605) );
  XOR2_X1 U11057 ( .A1(\RI5[1][26] ), .A2(\RI5[1][2] ), .Z(
        \MC_ARK_ARC_1_1/temp2[56] ) );
  NAND3_X1 U11058 ( .A1(\SB3_11/i0[6] ), .A2(\SB3_11/i0[8] ), .A3(
        \SB3_11/i0[7] ), .ZN(\SB3_11/Component_Function_0/NAND4_in[1] ) );
  NAND4_X2 U11060 ( .A1(\SB2_0_20/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_20/Component_Function_4/NAND4_in[1] ), .A3(n6166), .A4(n5606), 
        .ZN(\SB2_0_20/buf_output[4] ) );
  NAND3_X1 U11061 ( .A1(\SB2_0_20/i1[9] ), .A2(\SB2_0_20/i0_4 ), .A3(
        \SB2_0_20/i1_5 ), .ZN(n5606) );
  XOR2_X1 U11062 ( .A1(\MC_ARK_ARC_1_3/temp2[175] ), .A2(
        \MC_ARK_ARC_1_3/temp4[175] ), .Z(n5608) );
  NAND3_X1 U11063 ( .A1(\SB3_31/i0_3 ), .A2(\SB3_31/i0[10] ), .A3(
        \SB3_31/i0_4 ), .ZN(\SB3_31/Component_Function_0/NAND4_in[2] ) );
  NAND3_X1 U11066 ( .A1(\SB4_26/i0[9] ), .A2(\SB4_26/i0_0 ), .A3(
        \SB4_26/i0[8] ), .ZN(n5609) );
  NAND4_X2 U11069 ( .A1(\SB2_0_20/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_20/Component_Function_3/NAND4_in[3] ), .A3(
        \SB2_0_20/Component_Function_3/NAND4_in[1] ), .A4(n5610), .ZN(
        \SB2_0_20/buf_output[3] ) );
  NAND3_X1 U11072 ( .A1(\SB2_0_20/i0[10] ), .A2(\SB2_0_20/i1[9] ), .A3(
        \SB2_0_20/i1_7 ), .ZN(n5610) );
  XOR2_X1 U11073 ( .A1(n1230), .A2(\MC_ARK_ARC_1_2/temp2[117] ), .Z(n5611) );
  XOR2_X1 U11075 ( .A1(n5612), .A2(\MC_ARK_ARC_1_0/temp2[87] ), .Z(
        \MC_ARK_ARC_1_0/temp5[87] ) );
  XOR2_X1 U11076 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[81] ), .A2(\RI5[0][87] ), 
        .Z(n5612) );
  NAND4_X2 U11081 ( .A1(\SB2_0_28/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_0_28/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_0_28/Component_Function_1/NAND4_in[0] ), .A4(n5613), .ZN(
        \SB2_0_28/buf_output[1] ) );
  NAND4_X2 U11082 ( .A1(\SB1_2_31/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_31/Component_Function_0/NAND4_in[1] ), .A3(
        \SB1_2_31/Component_Function_0/NAND4_in[0] ), .A4(n5614), .ZN(
        \SB1_2_31/buf_output[0] ) );
  NAND3_X1 U11084 ( .A1(\SB1_2_31/i0_0 ), .A2(\SB1_2_31/i0_3 ), .A3(
        \SB1_2_31/i0[7] ), .ZN(n5614) );
  NAND3_X1 U11086 ( .A1(\SB3_0/i0_4 ), .A2(\SB3_0/i1_5 ), .A3(\SB3_0/i0_0 ), 
        .ZN(\SB3_0/Component_Function_2/NAND4_in[3] ) );
  XOR2_X1 U11087 ( .A1(n5615), .A2(n190), .Z(Ciphertext[16]) );
  NAND3_X2 U11092 ( .A1(\SB2_2_23/i0_3 ), .A2(\SB2_2_23/i0_0 ), .A3(
        \SB2_2_23/i0_4 ), .ZN(n5616) );
  XOR2_X1 U11093 ( .A1(n1762), .A2(n5617), .Z(n3276) );
  XOR2_X1 U11094 ( .A1(\RI5[0][62] ), .A2(\RI5[0][98] ), .Z(n5617) );
  NAND4_X2 U11098 ( .A1(\SB3_6/Component_Function_0/NAND4_in[1] ), .A2(n2527), 
        .A3(\SB3_6/Component_Function_0/NAND4_in[0] ), .A4(n5618), .ZN(
        \SB3_6/buf_output[0] ) );
  INV_X2 U11099 ( .I(\SB1_2_5/buf_output[3] ), .ZN(\SB2_2_3/i0[8] ) );
  XOR2_X1 U11102 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[90] ), .A2(n1375), .Z(
        \MC_ARK_ARC_1_0/temp2[144] ) );
  XOR2_X1 U11104 ( .A1(\MC_ARK_ARC_1_2/temp6[65] ), .A2(n5619), .Z(
        \MC_ARK_ARC_1_2/buf_output[65] ) );
  XOR2_X1 U11107 ( .A1(n5620), .A2(n2611), .Z(n3837) );
  XOR2_X1 U11108 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[50] ), .A2(\RI5[2][44] ), 
        .Z(n5620) );
  XOR2_X1 U11110 ( .A1(\MC_ARK_ARC_1_0/temp1[176] ), .A2(n5621), .Z(n6493) );
  XOR2_X1 U11111 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[86] ), .A2(\RI5[0][50] ), 
        .Z(n5621) );
  NAND4_X2 U11112 ( .A1(\SB1_2_16/Component_Function_3/NAND4_in[3] ), .A2(
        \SB1_2_16/Component_Function_3/NAND4_in[1] ), .A3(n6511), .A4(n5622), 
        .ZN(\SB1_2_16/buf_output[3] ) );
  NAND3_X1 U11113 ( .A1(\SB3_29/i0[10] ), .A2(\SB3_29/i0_3 ), .A3(
        \SB3_29/i0[9] ), .ZN(\SB3_29/Component_Function_4/NAND4_in[2] ) );
  XOR2_X1 U11114 ( .A1(\MC_ARK_ARC_1_0/temp5[147] ), .A2(
        \MC_ARK_ARC_1_0/temp6[147] ), .Z(n3659) );
  XOR2_X1 U11115 ( .A1(n6259), .A2(n2612), .Z(\MC_ARK_ARC_1_0/temp5[147] ) );
  XOR2_X1 U11121 ( .A1(n4624), .A2(n5623), .Z(n6340) );
  XOR2_X1 U11126 ( .A1(\RI5[0][35] ), .A2(\RI5[0][29] ), .Z(n5623) );
  XOR2_X1 U11127 ( .A1(n5624), .A2(n162), .Z(Ciphertext[19]) );
  NAND4_X2 U11129 ( .A1(\SB4_28/Component_Function_1/NAND4_in[2] ), .A2(
        \SB4_28/Component_Function_1/NAND4_in[3] ), .A3(
        \SB4_28/Component_Function_1/NAND4_in[1] ), .A4(n4291), .ZN(n5624) );
  XOR2_X1 U11130 ( .A1(\MC_ARK_ARC_1_3/temp5[154] ), .A2(n5625), .Z(
        \MC_ARK_ARC_1_3/buf_output[154] ) );
  XOR2_X1 U11132 ( .A1(\MC_ARK_ARC_1_3/temp4[154] ), .A2(
        \MC_ARK_ARC_1_3/temp3[154] ), .Z(n5625) );
  XOR2_X1 U11133 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[68] ), .A2(n496), .Z(
        n5626) );
  XOR2_X1 U11135 ( .A1(\RI5[2][134] ), .A2(\RI5[2][44] ), .Z(n5627) );
  NAND4_X2 U11136 ( .A1(n4426), .A2(n3406), .A3(n6173), .A4(
        \SB3_29/Component_Function_5/NAND4_in[0] ), .ZN(\SB3_29/buf_output[5] ) );
  NAND3_X2 U11146 ( .A1(\SB1_3_2/i0[10] ), .A2(\SB1_3_2/i0[6] ), .A3(
        \SB1_3_2/i0_3 ), .ZN(n5694) );
  NAND4_X2 U11148 ( .A1(n5876), .A2(n4655), .A3(n5631), .A4(
        \SB2_0_2/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_0_2/buf_output[3] ) );
  NAND4_X2 U11149 ( .A1(\SB2_1_10/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_10/Component_Function_3/NAND4_in[3] ), .A3(n6015), .A4(
        \SB2_1_10/Component_Function_3/NAND4_in[2] ), .ZN(
        \SB2_1_10/buf_output[3] ) );
  NAND3_X1 U11151 ( .A1(\SB2_0_2/i0_3 ), .A2(\RI3[0][175] ), .A3(
        \SB2_0_2/i0[10] ), .ZN(\SB2_0_2/Component_Function_2/NAND4_in[1] ) );
  NAND4_X2 U11153 ( .A1(\SB2_1_31/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_1_31/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_1_31/Component_Function_3/NAND4_in[1] ), .A4(
        \SB2_1_31/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_1_31/buf_output[3] ) );
  NAND4_X2 U11155 ( .A1(\SB2_2_7/Component_Function_2/NAND4_in[3] ), .A2(
        \SB2_2_7/Component_Function_2/NAND4_in[2] ), .A3(n2970), .A4(n5628), 
        .ZN(\SB2_2_7/buf_output[2] ) );
  NAND3_X2 U11158 ( .A1(\SB2_2_7/i0_3 ), .A2(\SB2_2_7/i0[10] ), .A3(
        \SB2_2_7/i0[6] ), .ZN(n5628) );
  XOR2_X1 U11164 ( .A1(\RI5[1][91] ), .A2(\RI5[1][181] ), .Z(n5630) );
  NAND3_X2 U11165 ( .A1(\SB2_0_2/i0[6] ), .A2(\SB2_0_2/i1[9] ), .A3(
        \SB2_0_2/i0_3 ), .ZN(n5631) );
  XOR2_X1 U11167 ( .A1(\RI5[0][91] ), .A2(\RI5[0][97] ), .Z(
        \MC_ARK_ARC_1_0/temp1[97] ) );
  XOR2_X1 U11172 ( .A1(\MC_ARK_ARC_1_1/temp2[142] ), .A2(n5632), .Z(
        \MC_ARK_ARC_1_1/temp5[142] ) );
  XOR2_X1 U11173 ( .A1(\RI5[1][136] ), .A2(\RI5[1][142] ), .Z(n5632) );
  NAND4_X2 U11176 ( .A1(\SB3_6/Component_Function_2/NAND4_in[3] ), .A2(
        \SB3_6/Component_Function_2/NAND4_in[0] ), .A3(
        \SB3_6/Component_Function_2/NAND4_in[1] ), .A4(
        \SB3_6/Component_Function_2/NAND4_in[2] ), .ZN(\SB3_6/buf_output[2] )
         );
  XOR2_X1 U11178 ( .A1(\MC_ARK_ARC_1_1/temp1[146] ), .A2(n5633), .Z(
        \MC_ARK_ARC_1_1/temp5[146] ) );
  XOR2_X1 U11179 ( .A1(\RI5[1][116] ), .A2(\RI5[1][92] ), .Z(n5633) );
  NAND3_X2 U11180 ( .A1(\SB2_3_3/i0[9] ), .A2(\SB2_3_3/i0_3 ), .A3(
        \SB2_3_3/i0[8] ), .ZN(n5634) );
  INV_X2 U11182 ( .I(\SB1_1_15/buf_output[2] ), .ZN(\SB2_1_12/i1[9] ) );
  NAND4_X2 U11183 ( .A1(\SB1_1_15/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_1_15/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_1_15/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_1_15/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB1_1_15/buf_output[2] ) );
  NAND3_X2 U11186 ( .A1(n5790), .A2(n2852), .A3(\SB2_1_7/i0[9] ), .ZN(n3308)
         );
  XOR2_X1 U11187 ( .A1(\RI5[1][132] ), .A2(\RI5[1][162] ), .Z(n5635) );
  XOR2_X1 U11188 ( .A1(n5836), .A2(n5636), .Z(\MC_ARK_ARC_1_2/buf_output[175] ) );
  XOR2_X1 U11190 ( .A1(\MC_ARK_ARC_1_2/temp4[175] ), .A2(
        \MC_ARK_ARC_1_2/temp3[175] ), .Z(n5636) );
  NAND3_X2 U11193 ( .A1(\SB2_2_19/i0[6] ), .A2(\SB2_2_19/i0_3 ), .A3(
        \SB2_2_19/i0[10] ), .ZN(\SB2_2_19/Component_Function_2/NAND4_in[1] )
         );
  NAND3_X2 U11194 ( .A1(\SB2_3_0/i0[6] ), .A2(\SB2_3_0/i0[10] ), .A3(
        \SB2_3_0/i0_0 ), .ZN(\SB2_3_0/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U11197 ( .A1(\SB1_0_4/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_4/Component_Function_2/NAND4_in[3] ), .A3(
        \SB1_0_4/Component_Function_2/NAND4_in[1] ), .A4(
        \SB1_0_4/Component_Function_2/NAND4_in[2] ), .ZN(\RI3[0][182] ) );
  NAND4_X2 U11198 ( .A1(\SB2_2_16/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_2_16/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_2_16/Component_Function_3/NAND4_in[3] ), .A4(n5638), .ZN(
        \SB2_2_16/buf_output[3] ) );
  XOR2_X1 U11199 ( .A1(\MC_ARK_ARC_1_0/temp1[2] ), .A2(n5639), .Z(
        \MC_ARK_ARC_1_0/temp5[2] ) );
  XOR2_X1 U11200 ( .A1(\RI5[0][140] ), .A2(\RI5[0][164] ), .Z(n5639) );
  INV_X2 U11203 ( .I(\SB1_2_29/buf_output[3] ), .ZN(\SB2_2_27/i0[8] ) );
  NAND4_X2 U11204 ( .A1(\SB1_2_29/Component_Function_3/NAND4_in[2] ), .A2(
        n4071), .A3(\SB1_2_29/Component_Function_3/NAND4_in[0] ), .A4(n6255), 
        .ZN(\SB1_2_29/buf_output[3] ) );
  XOR2_X1 U11207 ( .A1(n5641), .A2(\MC_ARK_ARC_1_1/temp5[49] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[49] ) );
  XOR2_X1 U11211 ( .A1(\MC_ARK_ARC_1_1/temp3[49] ), .A2(
        \MC_ARK_ARC_1_1/temp4[49] ), .Z(n5641) );
  NAND3_X2 U11214 ( .A1(\SB3_25/i0_0 ), .A2(\SB3_25/i0_4 ), .A3(\SB3_25/i1_5 ), 
        .ZN(n5642) );
  NAND4_X2 U11216 ( .A1(\SB2_3_31/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_3_31/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_3_31/Component_Function_1/NAND4_in[3] ), .A4(n5643), .ZN(
        \SB2_3_31/buf_output[1] ) );
  NOR2_X2 U11217 ( .A1(n5657), .A2(n6436), .ZN(n5644) );
  XOR2_X1 U11218 ( .A1(n2609), .A2(n5645), .Z(n3664) );
  NAND4_X2 U11219 ( .A1(\SB1_1_10/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_1_10/Component_Function_4/NAND4_in[1] ), .A3(n4301), .A4(n5646), 
        .ZN(\SB1_1_10/buf_output[4] ) );
  NAND4_X2 U11220 ( .A1(\SB1_3_4/Component_Function_3/NAND4_in[1] ), .A2(n1685), .A3(n5756), .A4(n5647), .ZN(\SB1_3_4/buf_output[3] ) );
  NAND4_X2 U11221 ( .A1(\SB1_1_29/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_1_29/Component_Function_1/NAND4_in[3] ), .A3(n5969), .A4(n5648), 
        .ZN(\SB1_1_29/buf_output[1] ) );
  NAND3_X2 U11222 ( .A1(\SB1_1_29/i0_3 ), .A2(\SB1_1_29/i0[8] ), .A3(
        \SB1_1_29/i1_7 ), .ZN(n5648) );
  NAND4_X2 U11223 ( .A1(n2498), .A2(\SB3_18/Component_Function_3/NAND4_in[1] ), 
        .A3(\SB3_18/Component_Function_3/NAND4_in[0] ), .A4(n5649), .ZN(
        \SB3_18/buf_output[3] ) );
  NAND3_X1 U11224 ( .A1(\SB3_18/i1_7 ), .A2(\SB3_18/i1[9] ), .A3(
        \SB3_18/i0[10] ), .ZN(n5649) );
  XOR2_X1 U11225 ( .A1(\RI5[3][39] ), .A2(\RI5[3][45] ), .Z(
        \MC_ARK_ARC_1_3/temp1[45] ) );
  NAND3_X1 U11226 ( .A1(\SB2_1_10/i0_3 ), .A2(\SB2_1_10/i0_0 ), .A3(
        \SB2_1_10/i0[7] ), .ZN(\SB2_1_10/Component_Function_0/NAND4_in[3] ) );
  XOR2_X1 U11227 ( .A1(n5651), .A2(n5650), .Z(\RI1[4][179] ) );
  XOR2_X1 U11228 ( .A1(n1217), .A2(\MC_ARK_ARC_1_3/temp4[179] ), .Z(n5651) );
  NAND4_X2 U11229 ( .A1(\SB4_18/Component_Function_4/NAND4_in[3] ), .A2(n1220), 
        .A3(n2627), .A4(n5652), .ZN(n3747) );
  NAND3_X2 U11230 ( .A1(\SB4_18/i0[10] ), .A2(\SB4_18/i0_3 ), .A3(
        \SB4_18/i0[9] ), .ZN(n5652) );
  XOR2_X1 U11231 ( .A1(n5653), .A2(n101), .Z(Ciphertext[174]) );
  NAND4_X2 U11232 ( .A1(\SB4_2/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_2/Component_Function_0/NAND4_in[1] ), .A3(n6075), .A4(
        \SB4_2/Component_Function_0/NAND4_in[0] ), .ZN(n5653) );
  NAND4_X2 U11233 ( .A1(\SB2_3_24/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_3_24/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_3_24/Component_Function_4/NAND4_in[0] ), .A4(n5654), .ZN(
        \SB2_3_24/buf_output[4] ) );
  NAND4_X2 U11234 ( .A1(\SB1_2_24/Component_Function_2/NAND4_in[3] ), .A2(
        \SB1_2_24/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_2_24/Component_Function_2/NAND4_in[2] ), .A4(n5655), .ZN(
        \SB1_2_24/buf_output[2] ) );
  NAND3_X2 U11235 ( .A1(\RI1[2][47] ), .A2(\SB1_2_24/i0[10] ), .A3(
        \SB1_2_24/i0[6] ), .ZN(n5655) );
  XOR2_X1 U11236 ( .A1(n5656), .A2(\MC_ARK_ARC_1_3/temp6[52] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[52] ) );
  XOR2_X1 U11237 ( .A1(\MC_ARK_ARC_1_3/temp2[52] ), .A2(
        \MC_ARK_ARC_1_3/temp1[52] ), .Z(n5656) );
  NAND4_X2 U11238 ( .A1(n2137), .A2(
        \SB1_3_10/Component_Function_3/NAND4_in[0] ), .A3(n4264), .A4(
        \SB1_3_10/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_3_10/buf_output[3] ) );
  NAND3_X2 U11239 ( .A1(\SB1_3_24/i0_4 ), .A2(\SB1_3_24/i0_3 ), .A3(
        \SB1_3_24/i1[9] ), .ZN(\SB1_3_24/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U11240 ( .A1(\RI5[2][32] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[56] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[86] ) );
  XOR2_X1 U11241 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[56] ), .A2(\RI5[2][8] ), 
        .Z(n2930) );
  XOR2_X1 U11242 ( .A1(\MC_ARK_ARC_1_3/temp6[121] ), .A2(n2987), .Z(
        \MC_ARK_ARC_1_3/buf_output[121] ) );
  XOR2_X1 U11243 ( .A1(\MC_ARK_ARC_1_2/temp4[47] ), .A2(n4375), .Z(n6175) );
  NAND4_X2 U11244 ( .A1(\SB2_2_21/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_2_21/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_2_21/Component_Function_2/NAND4_in[1] ), .A4(n5705), .ZN(
        \SB2_2_21/buf_output[2] ) );
  XOR2_X1 U11245 ( .A1(n5658), .A2(n218), .Z(Ciphertext[105]) );
  NAND4_X2 U11246 ( .A1(n2267), .A2(n2363), .A3(n4053), .A4(
        \SB4_14/Component_Function_3/NAND4_in[3] ), .ZN(n5658) );
  XOR2_X1 U11247 ( .A1(n5659), .A2(n226), .Z(Ciphertext[104]) );
  NAND4_X2 U11248 ( .A1(n3190), .A2(\SB4_14/Component_Function_2/NAND4_in[1] ), 
        .A3(\SB4_14/Component_Function_2/NAND4_in[2] ), .A4(n6491), .ZN(n5659)
         );
  XOR2_X1 U11249 ( .A1(n5660), .A2(\MC_ARK_ARC_1_0/temp4[98] ), .Z(n2460) );
  XOR2_X1 U11250 ( .A1(\RI5[0][8] ), .A2(\RI5[0][164] ), .Z(n5660) );
  XOR2_X1 U11251 ( .A1(n5661), .A2(\MC_ARK_ARC_1_0/temp4[149] ), .Z(n5964) );
  XOR2_X1 U11252 ( .A1(\RI5[0][143] ), .A2(\RI5[0][149] ), .Z(n5661) );
  NAND3_X2 U11253 ( .A1(\SB2_2_28/i0_3 ), .A2(\SB2_2_28/i0_4 ), .A3(
        \SB2_2_28/i0_0 ), .ZN(\SB2_2_28/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U11254 ( .A1(n3462), .A2(\SB3_2/Component_Function_1/NAND4_in[0] ), 
        .A3(\SB3_2/Component_Function_1/NAND4_in[1] ), .A4(n5662), .ZN(
        \SB3_2/buf_output[1] ) );
  NAND3_X2 U11255 ( .A1(\SB4_5/i0_0 ), .A2(\SB4_5/i0_4 ), .A3(\SB4_5/i1_5 ), 
        .ZN(n5663) );
  XOR2_X1 U11256 ( .A1(n5664), .A2(\MC_ARK_ARC_1_2/temp4[123] ), .Z(
        \MC_ARK_ARC_1_2/temp6[123] ) );
  XOR2_X1 U11257 ( .A1(\SB2_2_28/buf_output[3] ), .A2(\RI5[2][189] ), .Z(n5664) );
  NAND4_X2 U11258 ( .A1(\SB1_0_18/Component_Function_4/NAND4_in[1] ), .A2(
        \SB1_0_18/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_0_18/Component_Function_4/NAND4_in[3] ), .A4(n5665), .ZN(
        \SB1_0_18/buf_output[4] ) );
  NAND3_X1 U11259 ( .A1(\SB1_0_18/i0_3 ), .A2(\SB1_0_18/i0[9] ), .A3(n1367), 
        .ZN(n5665) );
  XOR2_X1 U11260 ( .A1(n5891), .A2(n5666), .Z(n5807) );
  XOR2_X1 U11261 ( .A1(\RI5[1][76] ), .A2(\RI5[1][178] ), .Z(n5666) );
  NAND3_X2 U11262 ( .A1(\SB4_5/i0_0 ), .A2(\SB4_5/i3[0] ), .A3(\SB4_5/i1_7 ), 
        .ZN(n5667) );
  INV_X2 U11263 ( .I(\SB1_1_11/buf_output[2] ), .ZN(\SB2_1_8/i1[9] ) );
  NAND4_X2 U11264 ( .A1(\SB1_1_11/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_11/Component_Function_2/NAND4_in[2] ), .A3(n5785), .A4(n5788), 
        .ZN(\SB1_1_11/buf_output[2] ) );
  NAND3_X2 U11265 ( .A1(\SB1_3_4/i0_4 ), .A2(\SB1_3_4/i0_0 ), .A3(
        \SB1_3_4/i0_3 ), .ZN(\SB1_3_4/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U11266 ( .A1(\SB1_1_4/i0_0 ), .A2(\SB1_1_4/i3[0] ), .A3(
        \SB1_1_4/i1_7 ), .ZN(n4719) );
  NAND4_X2 U11267 ( .A1(\SB2_0_29/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_0_29/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_0_29/Component_Function_3/NAND4_in[1] ), .A4(n2093), .ZN(
        \SB2_0_29/buf_output[3] ) );
  NAND4_X2 U11268 ( .A1(n3374), .A2(\SB2_3_0/Component_Function_5/NAND4_in[1] ), .A3(n5676), .A4(\SB2_3_0/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_3_0/buf_output[5] ) );
  NAND3_X1 U11269 ( .A1(\SB4_8/i0[10] ), .A2(\SB4_8/i1[9] ), .A3(\SB4_8/i1_5 ), 
        .ZN(\SB4_8/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U11270 ( .A1(\SB2_0_13/i0[6] ), .A2(\SB2_0_13/i0[9] ), .A3(
        \SB2_0_13/i0_4 ), .ZN(n5668) );
  NAND3_X1 U11271 ( .A1(\SB1_0_18/i0_3 ), .A2(\SB1_0_18/i1[9] ), .A3(
        \SB1_0_18/i0[6] ), .ZN(\SB1_0_18/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U11272 ( .A1(n6158), .A2(n833), .Z(\MC_ARK_ARC_1_0/buf_output[119] )
         );
  INV_X2 U11273 ( .I(\SB1_0_0/buf_output[2] ), .ZN(\SB2_0_29/i1[9] ) );
  NAND4_X2 U11274 ( .A1(\SB1_0_0/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_0/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_0/Component_Function_2/NAND4_in[2] ), .A4(n6474), .ZN(
        \SB1_0_0/buf_output[2] ) );
  NAND3_X1 U11275 ( .A1(\SB1_0_18/i0_3 ), .A2(n4753), .A3(n1367), .ZN(
        \SB1_0_18/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U11276 ( .A1(\MC_ARK_ARC_1_1/temp1[12] ), .A2(
        \MC_ARK_ARC_1_1/temp2[12] ), .Z(\MC_ARK_ARC_1_1/temp5[12] ) );
  NAND4_X2 U11277 ( .A1(\SB2_2_8/Component_Function_2/NAND4_in[2] ), .A2(n1249), .A3(\SB2_2_8/Component_Function_2/NAND4_in[0] ), .A4(
        \SB2_2_8/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_2_8/buf_output[2] ) );
  NAND4_X2 U11278 ( .A1(\SB1_0_18/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_0_18/Component_Function_5/NAND4_in[1] ), .A3(n1939), .A4(
        \SB1_0_18/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_0_18/buf_output[5] ) );
  NAND3_X2 U11279 ( .A1(\SB2_0_18/i0_3 ), .A2(\SB2_0_18/i1[9] ), .A3(
        \SB2_0_18/i0[6] ), .ZN(n4663) );
  XOR2_X1 U11280 ( .A1(\MC_ARK_ARC_1_3/temp6[125] ), .A2(
        \MC_ARK_ARC_1_3/temp5[125] ), .Z(n1381) );
  XOR2_X1 U11281 ( .A1(\MC_ARK_ARC_1_3/temp4[125] ), .A2(
        \MC_ARK_ARC_1_3/temp3[125] ), .Z(\MC_ARK_ARC_1_3/temp6[125] ) );
  XOR2_X1 U11282 ( .A1(\RI5[3][86] ), .A2(\RI5[3][92] ), .Z(
        \MC_ARK_ARC_1_3/temp1[92] ) );
  NAND3_X2 U11283 ( .A1(\SB1_3_4/i0[6] ), .A2(\SB1_3_4/i0_3 ), .A3(
        \SB1_3_4/i0[10] ), .ZN(\SB1_3_4/Component_Function_2/NAND4_in[1] ) );
  INV_X2 U11284 ( .I(\SB1_0_18/buf_output[2] ), .ZN(\SB2_0_15/i1[9] ) );
  NAND3_X2 U11285 ( .A1(\SB2_2_20/i0[10] ), .A2(\SB2_2_20/i1[9] ), .A3(
        \SB2_2_20/i1_7 ), .ZN(n1907) );
  INV_X2 U11286 ( .I(\SB3_24/buf_output[3] ), .ZN(\SB4_22/i0[8] ) );
  XOR2_X1 U11287 ( .A1(n4127), .A2(n5670), .Z(\MC_ARK_ARC_1_3/buf_output[155] ) );
  XOR2_X1 U11288 ( .A1(\MC_ARK_ARC_1_3/temp2[155] ), .A2(n1192), .Z(n5670) );
  XOR2_X1 U11289 ( .A1(n4236), .A2(n5671), .Z(n2195) );
  XOR2_X1 U11290 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[153] ), .A2(\RI5[2][189] ), .Z(n5671) );
  NAND3_X2 U11291 ( .A1(\SB1_0_21/i0[10] ), .A2(\SB1_0_21/i0_0 ), .A3(
        \SB1_0_21/i0[6] ), .ZN(n5672) );
  NAND3_X1 U11292 ( .A1(\SB1_0_17/i0[10] ), .A2(\SB1_0_17/i0_3 ), .A3(
        \SB1_0_17/i0[9] ), .ZN(n5673) );
  NAND4_X2 U11293 ( .A1(\SB1_2_5/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_2_5/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_5/Component_Function_1/NAND4_in[0] ), .A4(n5674), .ZN(
        \SB1_2_5/buf_output[1] ) );
  INV_X1 U11294 ( .I(\SB3_12/buf_output[1] ), .ZN(\SB4_8/i1_7 ) );
  NAND4_X2 U11295 ( .A1(n6213), .A2(\SB3_12/Component_Function_1/NAND4_in[1] ), 
        .A3(\SB3_12/Component_Function_1/NAND4_in[3] ), .A4(
        \SB3_12/Component_Function_1/NAND4_in[0] ), .ZN(\SB3_12/buf_output[1] ) );
  XOR2_X1 U11296 ( .A1(n5675), .A2(n593), .Z(\MC_ARK_ARC_1_2/buf_output[43] )
         );
  XOR2_X1 U11297 ( .A1(\MC_ARK_ARC_1_2/temp2[43] ), .A2(n584), .Z(n5675) );
  NAND4_X2 U11298 ( .A1(\SB1_1_10/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_1_10/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_1_10/Component_Function_3/NAND4_in[2] ), .A4(n3434), .ZN(
        \SB1_1_10/buf_output[3] ) );
  NAND3_X2 U11299 ( .A1(\SB2_3_0/i0[6] ), .A2(\SB1_3_1/buf_output[4] ), .A3(
        \SB2_3_0/i0[9] ), .ZN(n5676) );
  XOR2_X1 U11300 ( .A1(n5677), .A2(\MC_ARK_ARC_1_0/temp5[132] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[132] ) );
  XOR2_X1 U11301 ( .A1(\MC_ARK_ARC_1_0/temp4[132] ), .A2(
        \MC_ARK_ARC_1_0/temp3[132] ), .Z(n5677) );
  XOR2_X1 U11302 ( .A1(\MC_ARK_ARC_1_1/temp2[9] ), .A2(n5678), .Z(
        \MC_ARK_ARC_1_1/temp5[9] ) );
  XOR2_X1 U11303 ( .A1(\RI5[1][3] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[9] ), 
        .Z(n5678) );
  NAND3_X2 U11304 ( .A1(\SB2_0_14/i1[9] ), .A2(\RI3[0][106] ), .A3(
        \SB2_0_14/i0_3 ), .ZN(n1092) );
  XOR2_X1 U11305 ( .A1(\MC_ARK_ARC_1_0/temp3[75] ), .A2(
        \MC_ARK_ARC_1_0/temp4[75] ), .Z(\MC_ARK_ARC_1_0/temp6[75] ) );
  NAND4_X2 U11306 ( .A1(\SB2_0_15/Component_Function_3/NAND4_in[3] ), .A2(
        \SB2_0_15/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_0_15/Component_Function_3/NAND4_in[1] ), .A4(n5679), .ZN(
        \SB2_0_15/buf_output[3] ) );
  NAND3_X1 U11307 ( .A1(\SB2_2_17/i0[8] ), .A2(\SB2_2_17/i1_7 ), .A3(
        \SB1_2_18/buf_output[4] ), .ZN(
        \SB2_2_17/Component_Function_1/NAND4_in[3] ) );
  XOR2_X1 U11308 ( .A1(n5680), .A2(n10), .Z(Ciphertext[175]) );
  NAND4_X2 U11309 ( .A1(\SB4_2/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_2/Component_Function_1/NAND4_in[0] ), .A3(n2569), .A4(
        \SB4_2/Component_Function_1/NAND4_in[2] ), .ZN(n5680) );
  NAND3_X2 U11310 ( .A1(\SB1_1_0/i0[10] ), .A2(\SB1_1_0/i1[9] ), .A3(
        \SB1_1_0/i1_5 ), .ZN(\SB1_1_0/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U11311 ( .A1(n1457), .A2(
        \SB1_2_24/Component_Function_4/NAND4_in[0] ), .A3(
        \SB1_2_24/Component_Function_4/NAND4_in[2] ), .A4(
        \SB1_2_24/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB1_2_24/buf_output[4] ) );
  XOR2_X1 U11312 ( .A1(n4134), .A2(n5681), .Z(\MC_ARK_ARC_1_3/buf_output[156] ) );
  XOR2_X1 U11313 ( .A1(\MC_ARK_ARC_1_3/temp4[156] ), .A2(n805), .Z(n5681) );
  NAND4_X2 U11314 ( .A1(\SB2_0_22/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_0_22/Component_Function_3/NAND4_in[0] ), .A3(n2274), .A4(n5682), 
        .ZN(\SB2_0_22/buf_output[3] ) );
  NAND3_X2 U11315 ( .A1(\SB2_0_22/i0_4 ), .A2(\SB2_0_22/i0_0 ), .A3(
        \SB2_0_22/i0_3 ), .ZN(n5682) );
  NAND3_X2 U11316 ( .A1(\SB2_1_28/i0_4 ), .A2(\SB2_1_28/i0_3 ), .A3(
        \SB2_1_28/i1[9] ), .ZN(\SB2_1_28/Component_Function_5/NAND4_in[2] ) );
  INV_X1 U11317 ( .I(\SB1_3_4/buf_output[0] ), .ZN(\SB2_3_31/i3[0] ) );
  NAND4_X2 U11318 ( .A1(\SB1_3_4/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_3_4/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_3_4/Component_Function_0/NAND4_in[2] ), .A4(
        \SB1_3_4/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_3_4/buf_output[0] ) );
  XOR2_X1 U11319 ( .A1(n5685), .A2(n219), .Z(Ciphertext[2]) );
  NAND4_X2 U11320 ( .A1(\SB2_2_22/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_22/Component_Function_2/NAND4_in[2] ), .A3(n4568), .A4(n5686), 
        .ZN(\SB2_2_22/buf_output[2] ) );
  NAND3_X2 U11321 ( .A1(\SB2_2_22/i0[10] ), .A2(\SB2_2_22/i0_3 ), .A3(
        \SB2_2_22/i0[6] ), .ZN(n5686) );
  INV_X1 U11322 ( .I(\SB1_2_24/buf_output[5] ), .ZN(\SB2_2_24/i1_5 ) );
  XOR2_X1 U11323 ( .A1(n5687), .A2(\MC_ARK_ARC_1_3/temp4[35] ), .Z(n3728) );
  XOR2_X1 U11324 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[101] ), .A2(\RI5[3][137] ), .Z(n5687) );
  NAND3_X2 U11325 ( .A1(\SB2_3_15/i0[6] ), .A2(\SB2_3_15/i0[9] ), .A3(
        \SB1_3_16/buf_output[4] ), .ZN(n4485) );
  XOR2_X1 U11326 ( .A1(n877), .A2(n5688), .Z(\MC_ARK_ARC_1_2/temp5[123] ) );
  XOR2_X1 U11327 ( .A1(\RI5[2][69] ), .A2(\RI5[2][93] ), .Z(n5688) );
  XOR2_X1 U11328 ( .A1(\MC_ARK_ARC_1_2/temp5[165] ), .A2(n5689), .Z(
        \MC_ARK_ARC_1_2/buf_output[165] ) );
  XOR2_X1 U11329 ( .A1(n6004), .A2(\MC_ARK_ARC_1_2/temp4[165] ), .Z(n5689) );
  INV_X2 U11330 ( .I(n5690), .ZN(n3660) );
  NAND4_X2 U11331 ( .A1(\SB1_1_7/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_7/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_1_7/Component_Function_2/NAND4_in[2] ), .A4(
        \SB1_1_7/Component_Function_2/NAND4_in[3] ), .ZN(n5690) );
  NAND3_X2 U11332 ( .A1(\SB2_1_26/i0_3 ), .A2(\SB2_1_26/i0[9] ), .A3(
        \SB2_1_26/i0[8] ), .ZN(\SB2_1_26/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 U11333 ( .A1(\SB1_1_3/Component_Function_2/NAND4_in[0] ), .A2(n741), 
        .A3(\SB1_1_3/Component_Function_2/NAND4_in[2] ), .A4(n5691), .ZN(
        \SB1_1_3/buf_output[2] ) );
  NAND3_X2 U11334 ( .A1(\SB1_1_3/i0[10] ), .A2(\SB1_1_3/i0[6] ), .A3(
        \SB1_1_3/i0_3 ), .ZN(n5691) );
  NAND3_X2 U11335 ( .A1(\SB2_1_9/i0[6] ), .A2(\SB2_1_9/i0_4 ), .A3(
        \SB2_1_9/i0[9] ), .ZN(n5692) );
  NAND4_X2 U11336 ( .A1(n2842), .A2(
        \SB2_1_15/Component_Function_2/NAND4_in[0] ), .A3(n5848), .A4(n5693), 
        .ZN(\SB2_1_15/buf_output[2] ) );
  NAND4_X2 U11337 ( .A1(\SB4_18/Component_Function_2/NAND4_in[2] ), .A2(n3468), 
        .A3(n3948), .A4(n5695), .ZN(n5707) );
  NAND3_X2 U11338 ( .A1(\SB4_18/i0_0 ), .A2(\SB4_18/i0_4 ), .A3(\SB4_18/i1_5 ), 
        .ZN(n5695) );
  XOR2_X1 U11339 ( .A1(n5696), .A2(n212), .Z(Ciphertext[38]) );
  NAND4_X2 U11340 ( .A1(\SB4_25/Component_Function_2/NAND4_in[1] ), .A2(
        \SB4_25/Component_Function_2/NAND4_in[3] ), .A3(n3137), .A4(
        \SB4_25/Component_Function_2/NAND4_in[2] ), .ZN(n5696) );
  NAND3_X1 U11341 ( .A1(\SB3_26/i0_4 ), .A2(\SB3_26/i0_0 ), .A3(\SB3_26/i1_5 ), 
        .ZN(n4566) );
  NAND3_X1 U11342 ( .A1(\SB3_26/i0_4 ), .A2(\SB3_26/i1_7 ), .A3(\SB3_26/i0[8] ), .ZN(\SB3_26/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U11343 ( .A1(\SB3_26/Component_Function_4/NAND4_in[1] ), .A2(
        \SB3_26/Component_Function_4/NAND4_in[0] ), .A3(
        \SB3_26/Component_Function_4/NAND4_in[2] ), .A4(n5697), .ZN(
        \SB3_26/buf_output[4] ) );
  NAND3_X1 U11344 ( .A1(\SB3_26/i0_4 ), .A2(\SB3_26/i1[9] ), .A3(\SB3_26/i1_5 ), .ZN(n5697) );
  INV_X2 U11345 ( .I(\SB1_2_16/buf_output[3] ), .ZN(\SB2_2_14/i0[8] ) );
  NAND4_X2 U11346 ( .A1(\SB2_2_14/Component_Function_3/NAND4_in[3] ), .A2(
        \SB2_2_14/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_2_14/Component_Function_3/NAND4_in[2] ), .A4(n1597), .ZN(
        \SB2_2_14/buf_output[3] ) );
  NAND3_X1 U11347 ( .A1(\SB3_12/i0_3 ), .A2(\SB3_12/i1[9] ), .A3(
        \SB3_12/i0[6] ), .ZN(\SB3_12/Component_Function_3/NAND4_in[0] ) );
  NAND4_X2 U11348 ( .A1(\SB2_2_20/Component_Function_3/NAND4_in[3] ), .A2(
        n6178), .A3(n1907), .A4(n6475), .ZN(\SB2_2_20/buf_output[3] ) );
  NAND4_X2 U11349 ( .A1(n3973), .A2(
        \SB2_3_12/Component_Function_5/NAND4_in[2] ), .A3(n6391), .A4(n2099), 
        .ZN(\SB2_3_12/buf_output[5] ) );
  NAND4_X2 U11350 ( .A1(\SB2_3_29/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_3_29/Component_Function_2/NAND4_in[3] ), .A3(n6063), .A4(
        \SB2_3_29/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB2_3_29/buf_output[2] ) );
  XOR2_X1 U11351 ( .A1(n5698), .A2(n222), .Z(Ciphertext[143]) );
  NAND4_X2 U11352 ( .A1(\SB3_14/Component_Function_2/NAND4_in[0] ), .A2(n6174), 
        .A3(\SB3_14/Component_Function_2/NAND4_in[2] ), .A4(
        \SB3_14/Component_Function_2/NAND4_in[3] ), .ZN(\SB3_14/buf_output[2] ) );
  NAND3_X2 U11353 ( .A1(\SB1_3_18/i0[8] ), .A2(\SB1_3_18/i0_4 ), .A3(
        \SB1_3_18/i1_7 ), .ZN(\SB1_3_18/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U11354 ( .A1(\SB2_3_22/Component_Function_3/NAND4_in[3] ), .A2(
        \SB2_3_22/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_3_22/Component_Function_3/NAND4_in[1] ), .A4(
        \SB2_3_22/Component_Function_3/NAND4_in[2] ), .ZN(
        \SB2_3_22/buf_output[3] ) );
  NAND4_X2 U11355 ( .A1(\SB2_3_17/Component_Function_5/NAND4_in[2] ), .A2(
        n3584), .A3(\SB2_3_17/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_3_17/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_3_17/buf_output[5] ) );
  NAND4_X2 U11356 ( .A1(\SB1_2_20/Component_Function_2/NAND4_in[1] ), .A2(
        n4152), .A3(n6465), .A4(n5699), .ZN(\SB1_2_20/buf_output[2] ) );
  XOR2_X1 U11357 ( .A1(\RI5[3][39] ), .A2(\RI5[3][33] ), .Z(n5700) );
  NAND3_X2 U11358 ( .A1(\SB2_3_22/i0_3 ), .A2(\SB2_3_22/i0[9] ), .A3(
        \SB2_3_22/i0[8] ), .ZN(\SB2_3_22/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U11359 ( .A1(\SB1_3_27/i0[6] ), .A2(\SB1_3_27/i0[8] ), .A3(
        \SB1_3_27/i0[7] ), .ZN(\SB1_3_27/Component_Function_0/NAND4_in[1] ) );
  XOR2_X1 U11360 ( .A1(\MC_ARK_ARC_1_1/temp4[69] ), .A2(n5702), .Z(
        \MC_ARK_ARC_1_1/temp6[69] ) );
  XOR2_X1 U11361 ( .A1(\RI5[1][171] ), .A2(\RI5[1][135] ), .Z(n5702) );
  NAND3_X2 U11362 ( .A1(\SB2_3_27/i0_3 ), .A2(\SB2_3_27/i0[10] ), .A3(n3680), 
        .ZN(n5703) );
  NAND4_X2 U11363 ( .A1(\SB2_1_5/Component_Function_0/NAND4_in[3] ), .A2(n2078), .A3(\SB2_1_5/Component_Function_0/NAND4_in[0] ), .A4(n5704), .ZN(
        \SB2_1_5/buf_output[0] ) );
  NAND3_X1 U11364 ( .A1(\SB2_1_5/i0[10] ), .A2(\SB2_1_5/i0_3 ), .A3(
        \SB1_1_6/buf_output[4] ), .ZN(n5704) );
  NAND3_X2 U11365 ( .A1(\SB2_2_21/i0_0 ), .A2(\SB2_2_21/i1_5 ), .A3(
        \SB2_2_21/i0_4 ), .ZN(n5705) );
  NAND3_X1 U11366 ( .A1(\SB1_0_16/i0_0 ), .A2(\SB1_0_16/i1_7 ), .A3(
        \SB1_0_16/i3[0] ), .ZN(\SB1_0_16/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U11367 ( .A1(\RI5[2][80] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[86] ), 
        .Z(n5706) );
  XOR2_X1 U11368 ( .A1(n5707), .A2(n203), .Z(Ciphertext[80]) );
  XOR2_X1 U11369 ( .A1(\RI5[2][121] ), .A2(\RI5[2][157] ), .Z(n3130) );
  NAND4_X2 U11370 ( .A1(\SB1_2_12/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_2_12/Component_Function_4/NAND4_in[3] ), .A3(
        \SB1_2_12/Component_Function_4/NAND4_in[0] ), .A4(n5709), .ZN(
        \SB1_2_12/buf_output[4] ) );
  NAND3_X2 U11371 ( .A1(\SB2_3_27/i0_3 ), .A2(\SB1_3_31/buf_output[1] ), .A3(
        \SB2_3_27/i1[9] ), .ZN(\SB2_3_27/Component_Function_3/NAND4_in[0] ) );
  NAND3_X2 U11372 ( .A1(\SB1_3_11/i0[6] ), .A2(\SB1_3_11/i0[10] ), .A3(
        \SB1_3_11/i0_0 ), .ZN(n6275) );
  XOR2_X1 U11373 ( .A1(\RI5[3][11] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[5] ), 
        .Z(n3156) );
  NAND3_X1 U11374 ( .A1(\SB2_2_9/i0[6] ), .A2(\SB1_2_14/buf_output[0] ), .A3(
        n3687), .ZN(\SB2_2_9/Component_Function_1/NAND4_in[2] ) );
  NAND3_X2 U11375 ( .A1(\SB2_3_8/i0[6] ), .A2(\SB2_3_8/i0[10] ), .A3(
        \SB2_3_8/i0_0 ), .ZN(n3544) );
  NAND4_X2 U11376 ( .A1(\SB3_23/Component_Function_2/NAND4_in[1] ), .A2(
        \SB3_23/Component_Function_2/NAND4_in[0] ), .A3(n942), .A4(n4597), 
        .ZN(\SB3_23/buf_output[2] ) );
  NAND4_X2 U11377 ( .A1(n4003), .A2(n3717), .A3(
        \SB2_2_5/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_2_5/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_2_5/buf_output[5] ) );
  INV_X1 U11378 ( .I(\SB3_23/buf_output[2] ), .ZN(\SB4_20/i1[9] ) );
  NAND3_X2 U11379 ( .A1(\SB2_1_9/i0_4 ), .A2(\SB2_1_9/i0_0 ), .A3(
        \SB2_1_9/i0_3 ), .ZN(n5710) );
  XOR2_X1 U11380 ( .A1(\MC_ARK_ARC_1_1/temp2[70] ), .A2(n5711), .Z(n4524) );
  XOR2_X1 U11381 ( .A1(\RI5[1][70] ), .A2(\RI5[1][64] ), .Z(n5711) );
  NAND4_X2 U11382 ( .A1(n2152), .A2(
        \SB2_2_13/Component_Function_3/NAND4_in[2] ), .A3(n5983), .A4(n5712), 
        .ZN(\SB2_2_13/buf_output[3] ) );
  XOR2_X1 U11383 ( .A1(\RI5[2][165] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[141] ), .Z(n4469) );
  XOR2_X1 U11384 ( .A1(n5713), .A2(n2927), .Z(\MC_ARK_ARC_1_1/temp5[135] ) );
  XOR2_X1 U11385 ( .A1(\RI5[1][81] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[105] ), 
        .Z(n5713) );
  XOR2_X1 U11386 ( .A1(n5714), .A2(n130), .Z(Ciphertext[108]) );
  NAND4_X2 U11387 ( .A1(n4746), .A2(\SB4_13/Component_Function_0/NAND4_in[2] ), 
        .A3(\SB4_13/Component_Function_0/NAND4_in[1] ), .A4(
        \SB4_13/Component_Function_0/NAND4_in[0] ), .ZN(n5714) );
  XOR2_X1 U11388 ( .A1(n5715), .A2(n232), .Z(Ciphertext[4]) );
  NAND4_X2 U11389 ( .A1(n4565), .A2(\SB4_31/Component_Function_4/NAND4_in[3] ), 
        .A3(n2428), .A4(n2531), .ZN(n5715) );
  XOR2_X1 U11390 ( .A1(n5716), .A2(n1518), .Z(\RI1[4][53] ) );
  XOR2_X1 U11391 ( .A1(n914), .A2(\MC_ARK_ARC_1_3/temp2[53] ), .Z(n5716) );
  NAND4_X2 U11392 ( .A1(\SB1_2_16/Component_Function_1/NAND4_in[2] ), .A2(
        n4024), .A3(\SB1_2_16/Component_Function_1/NAND4_in[1] ), .A4(n5717), 
        .ZN(\SB1_2_16/buf_output[1] ) );
  NAND2_X1 U11393 ( .A1(\SB1_2_16/i1[9] ), .A2(\RI1[2][95] ), .ZN(n5717) );
  XOR2_X1 U11394 ( .A1(n5718), .A2(n2937), .Z(\MC_ARK_ARC_1_3/temp6[176] ) );
  XOR2_X1 U11395 ( .A1(\RI5[3][20] ), .A2(\RI5[3][50] ), .Z(n5718) );
  XOR2_X1 U11396 ( .A1(n3730), .A2(\MC_ARK_ARC_1_2/temp6[177] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[177] ) );
  XOR2_X1 U11397 ( .A1(\MC_ARK_ARC_1_2/temp2[177] ), .A2(
        \MC_ARK_ARC_1_2/temp1[177] ), .Z(n3730) );
  NAND3_X1 U11398 ( .A1(\SB2_2_16/i0_3 ), .A2(\SB1_2_17/buf_output[4] ), .A3(
        \SB2_2_16/i0[10] ), .ZN(n5719) );
  NAND3_X2 U11399 ( .A1(\SB1_2_16/i0[9] ), .A2(\SB1_2_16/i0[6] ), .A3(
        \SB1_2_16/i0_4 ), .ZN(n715) );
  NAND4_X2 U11400 ( .A1(\SB1_3_6/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_3_6/Component_Function_1/NAND4_in[3] ), .A3(n3753), .A4(n5720), 
        .ZN(\SB1_3_6/buf_output[1] ) );
  NAND4_X2 U11401 ( .A1(n5809), .A2(
        \SB2_3_11/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_11/Component_Function_2/NAND4_in[0] ), .A4(
        \SB2_3_11/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_3_11/buf_output[2] ) );
  XOR2_X1 U11402 ( .A1(n5875), .A2(n5874), .Z(\MC_ARK_ARC_1_0/buf_output[50] )
         );
  XOR2_X1 U11403 ( .A1(n5722), .A2(n5721), .Z(\MC_ARK_ARC_1_0/buf_output[144] ) );
  XOR2_X1 U11404 ( .A1(\MC_ARK_ARC_1_0/temp4[144] ), .A2(
        \MC_ARK_ARC_1_0/temp2[144] ), .Z(n5721) );
  XOR2_X1 U11405 ( .A1(n6080), .A2(\MC_ARK_ARC_1_0/temp1[144] ), .Z(n5722) );
  XOR2_X1 U11406 ( .A1(n1054), .A2(n5723), .Z(\MC_ARK_ARC_1_1/temp5[169] ) );
  XOR2_X1 U11407 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[163] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[169] ), .Z(n5723) );
  NAND3_X2 U11408 ( .A1(\SB1_2_16/i0[10] ), .A2(\SB1_2_16/i0[9] ), .A3(
        \RI1[2][95] ), .ZN(\SB1_2_16/Component_Function_4/NAND4_in[2] ) );
  NAND4_X2 U11409 ( .A1(\SB1_0_8/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_0_8/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_0_8/Component_Function_0/NAND4_in[0] ), .A4(
        \SB1_0_8/Component_Function_0/NAND4_in[1] ), .ZN(
        \SB1_0_8/buf_output[0] ) );
  NAND3_X1 U11410 ( .A1(\SB2_1_23/i0_3 ), .A2(\SB2_1_23/i0[6] ), .A3(
        \SB2_1_23/i0[10] ), .ZN(\SB2_1_23/Component_Function_2/NAND4_in[1] )
         );
  NAND4_X2 U11411 ( .A1(\SB4_6/Component_Function_2/NAND4_in[3] ), .A2(
        \SB4_6/Component_Function_2/NAND4_in[0] ), .A3(n5844), .A4(n5724), 
        .ZN(n5850) );
  XOR2_X1 U11412 ( .A1(\RI5[3][2] ), .A2(\RI5[3][158] ), .Z(
        \MC_ARK_ARC_1_3/temp3[92] ) );
  XOR2_X1 U11413 ( .A1(\MC_ARK_ARC_1_1/temp5[135] ), .A2(n2117), .Z(
        \MC_ARK_ARC_1_1/buf_output[135] ) );
  NAND3_X2 U11414 ( .A1(\SB2_2_7/i0_3 ), .A2(\SB2_2_7/i0[9] ), .A3(
        \SB2_2_7/i0[8] ), .ZN(\SB2_2_7/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 U11415 ( .A1(n2575), .A2(n4311), .A3(
        \SB1_2_26/Component_Function_5/NAND4_in[1] ), .A4(
        \SB1_2_26/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_2_26/buf_output[5] ) );
  NAND2_X2 U11416 ( .A1(n3913), .A2(n4760), .ZN(\RI5[1][147] ) );
  NAND3_X2 U11417 ( .A1(\SB2_3_12/i0_3 ), .A2(\SB2_3_12/i0_4 ), .A3(
        \SB2_3_12/i1[9] ), .ZN(\SB2_3_12/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U11418 ( .A1(\MC_ARK_ARC_1_2/temp5[10] ), .A2(n5725), .Z(
        \MC_ARK_ARC_1_2/buf_output[10] ) );
  XOR2_X1 U11419 ( .A1(\MC_ARK_ARC_1_2/temp4[10] ), .A2(
        \MC_ARK_ARC_1_2/temp3[10] ), .Z(n5725) );
  XOR2_X1 U11420 ( .A1(\RI5[2][71] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[47] ), 
        .Z(n5726) );
  XOR2_X1 U11421 ( .A1(n5727), .A2(n13), .Z(Ciphertext[131]) );
  NAND4_X2 U11422 ( .A1(\SB4_10/Component_Function_5/NAND4_in[1] ), .A2(n4604), 
        .A3(\SB4_10/Component_Function_5/NAND4_in[2] ), .A4(
        \SB4_10/Component_Function_5/NAND4_in[0] ), .ZN(n5727) );
  XOR2_X1 U11423 ( .A1(n5730), .A2(n16), .Z(Ciphertext[155]) );
  NAND4_X2 U11424 ( .A1(\SB4_6/Component_Function_5/NAND4_in[1] ), .A2(
        \SB4_6/Component_Function_5/NAND4_in[2] ), .A3(
        \SB4_6/Component_Function_5/NAND4_in[3] ), .A4(
        \SB4_6/Component_Function_5/NAND4_in[0] ), .ZN(n5730) );
  XOR2_X1 U11425 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[44] ), .A2(\RI5[0][128] ), 
        .Z(n1416) );
  NAND4_X2 U11426 ( .A1(\SB2_2_29/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_29/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_29/Component_Function_5/NAND4_in[0] ), .A4(n5731), .ZN(
        \SB2_2_29/buf_output[5] ) );
  NAND3_X2 U11427 ( .A1(n1837), .A2(\SB2_2_29/i0[9] ), .A3(\SB2_2_29/i0[6] ), 
        .ZN(n5731) );
  XOR2_X1 U11428 ( .A1(n6071), .A2(n5732), .Z(\MC_ARK_ARC_1_1/buf_output[179] ) );
  XOR2_X1 U11429 ( .A1(\MC_ARK_ARC_1_1/temp3[179] ), .A2(
        \MC_ARK_ARC_1_1/temp4[179] ), .Z(n5732) );
  NAND4_X2 U11430 ( .A1(\SB3_10/Component_Function_2/NAND4_in[1] ), .A2(
        \SB3_10/Component_Function_2/NAND4_in[0] ), .A3(
        \SB3_10/Component_Function_2/NAND4_in[3] ), .A4(n5733), .ZN(
        \SB3_10/buf_output[2] ) );
  NAND3_X2 U11431 ( .A1(\SB2_1_21/i0[10] ), .A2(\SB2_1_21/i0[6] ), .A3(
        \SB2_1_21/i0_0 ), .ZN(n856) );
  XOR2_X1 U11432 ( .A1(n2344), .A2(n5734), .Z(n3513) );
  XOR2_X1 U11433 ( .A1(\RI5[0][20] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[44] ), 
        .Z(n5734) );
  NAND3_X1 U11434 ( .A1(\SB3_10/i0[8] ), .A2(\SB3_10/i1_7 ), .A3(\SB3_10/i0_3 ), .ZN(n1575) );
  NAND4_X2 U11435 ( .A1(\SB2_2_24/Component_Function_2/NAND4_in[0] ), .A2(
        n3201), .A3(\SB2_2_24/Component_Function_2/NAND4_in[2] ), .A4(n5735), 
        .ZN(\SB2_2_24/buf_output[2] ) );
  NAND3_X2 U11436 ( .A1(\SB2_2_24/i0[10] ), .A2(\SB2_2_24/i0_3 ), .A3(
        \SB2_2_24/i0[6] ), .ZN(n5735) );
  XOR2_X1 U11437 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[38] ), .A2(\RI5[1][44] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[44] ) );
  NAND3_X2 U11438 ( .A1(\SB2_2_20/i0[6] ), .A2(\SB2_2_20/i0[10] ), .A3(
        \SB2_2_20/i0_3 ), .ZN(n5736) );
  NAND3_X1 U11439 ( .A1(\SB4_31/i0_0 ), .A2(n3652), .A3(\SB4_31/i0[9] ), .ZN(
        n4565) );
  NAND3_X2 U11440 ( .A1(\SB2_1_20/i0[10] ), .A2(\SB2_1_20/i1_5 ), .A3(
        \SB2_1_20/i1[9] ), .ZN(\SB2_1_20/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U11441 ( .A1(\SB2_0_8/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_8/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_0_8/Component_Function_2/NAND4_in[1] ), .A4(
        \SB2_0_8/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_0_8/buf_output[2] ) );
  XOR2_X1 U11442 ( .A1(\RI5[1][86] ), .A2(\RI5[1][92] ), .Z(n5772) );
  XOR2_X1 U11443 ( .A1(\RI5[0][158] ), .A2(\RI5[0][152] ), .Z(
        \MC_ARK_ARC_1_0/temp1[158] ) );
  XOR2_X1 U11444 ( .A1(\MC_ARK_ARC_1_1/temp6[116] ), .A2(n5843), .Z(
        \MC_ARK_ARC_1_1/buf_output[116] ) );
  XOR2_X1 U11445 ( .A1(\SB2_0_31/buf_output[2] ), .A2(n141), .Z(n5737) );
  XOR2_X1 U11446 ( .A1(\RI5[1][142] ), .A2(n193), .Z(n6231) );
  NAND2_X2 U11447 ( .A1(n6301), .A2(n5738), .ZN(n6300) );
  NAND3_X2 U11448 ( .A1(\SB2_1_5/i0_0 ), .A2(\SB2_1_5/i0_3 ), .A3(
        \SB1_1_6/buf_output[4] ), .ZN(n5738) );
  NAND4_X2 U11449 ( .A1(\SB2_3_14/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_3_14/Component_Function_4/NAND4_in[0] ), .A3(n5739), .A4(
        \SB2_3_14/Component_Function_4/NAND4_in[2] ), .ZN(
        \SB2_3_14/buf_output[4] ) );
  NAND3_X1 U11450 ( .A1(\SB2_3_14/i0_4 ), .A2(\SB2_3_14/i1_5 ), .A3(
        \SB2_3_14/i1[9] ), .ZN(n5739) );
  NAND3_X1 U11451 ( .A1(\SB1_3_17/i0_0 ), .A2(\MC_ARK_ARC_1_2/buf_output[88] ), 
        .A3(\SB1_3_17/i0_3 ), .ZN(\SB1_3_17/Component_Function_3/NAND4_in[1] )
         );
  NAND4_X2 U11452 ( .A1(\SB2_1_12/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_12/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_1_12/Component_Function_5/NAND4_in[0] ), .A4(n5740), .ZN(
        \SB2_1_12/buf_output[5] ) );
  NAND3_X2 U11453 ( .A1(\SB2_1_12/i0[9] ), .A2(\SB2_1_12/i0_4 ), .A3(
        \SB2_1_12/i0[6] ), .ZN(n5740) );
  NAND2_X2 U11454 ( .A1(n5764), .A2(n567), .ZN(\RI5[1][171] ) );
  NAND4_X2 U11455 ( .A1(\SB2_0_26/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_26/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_0_26/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_0_26/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB2_0_26/buf_output[2] ) );
  NAND4_X2 U11456 ( .A1(\SB2_3_15/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_3_15/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_15/Component_Function_2/NAND4_in[3] ), .A4(n5741), .ZN(
        \SB2_3_15/buf_output[2] ) );
  NAND3_X2 U11457 ( .A1(\SB2_3_15/i0_3 ), .A2(\SB2_3_15/i0[9] ), .A3(n3670), 
        .ZN(n5741) );
  NAND3_X2 U11458 ( .A1(\SB1_3_0/i1[9] ), .A2(\SB1_3_0/i0[10] ), .A3(
        \SB1_3_0/i1_7 ), .ZN(n5742) );
  XOR2_X1 U11459 ( .A1(\MC_ARK_ARC_1_0/temp6[139] ), .A2(n1424), .Z(
        \MC_ARK_ARC_1_0/buf_output[139] ) );
  BUF_X4 U11460 ( .I(\SB2_1_7/i0_4 ), .Z(n5790) );
  NAND4_X1 U11461 ( .A1(\SB2_0_30/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_0_30/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_0_30/Component_Function_1/NAND4_in[2] ), .A4(n6356), .ZN(
        \SB2_0_30/buf_output[1] ) );
  XOR2_X1 U11462 ( .A1(\MC_ARK_ARC_1_3/temp5[62] ), .A2(n5743), .Z(
        \MC_ARK_ARC_1_3/buf_output[62] ) );
  INV_X2 U11463 ( .I(\SB1_3_21/buf_output[2] ), .ZN(\SB2_3_18/i1[9] ) );
  NAND4_X2 U11464 ( .A1(\SB2_1_9/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_1_9/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_1_9/Component_Function_4/NAND4_in[1] ), .A4(n5744), .ZN(
        \SB2_1_9/buf_output[4] ) );
  NAND3_X1 U11465 ( .A1(\SB2_1_9/i0_0 ), .A2(\SB2_1_9/i0[9] ), .A3(
        \SB2_1_9/i0[8] ), .ZN(n5744) );
  NAND3_X2 U11466 ( .A1(\SB1_1_27/i0[9] ), .A2(\SB1_1_27/i0[6] ), .A3(
        \SB1_1_27/i0_4 ), .ZN(n1745) );
  NAND4_X2 U11467 ( .A1(\SB1_1_5/Component_Function_3/NAND4_in[1] ), .A2(n1164), .A3(\SB1_1_5/Component_Function_3/NAND4_in[2] ), .A4(n5746), .ZN(
        \SB1_1_5/buf_output[3] ) );
  NAND3_X2 U11468 ( .A1(\SB1_1_5/i0[8] ), .A2(\SB1_1_5/i3[0] ), .A3(
        \SB1_1_5/i1_5 ), .ZN(n5746) );
  XOR2_X1 U11469 ( .A1(n5747), .A2(n5748), .Z(\MC_ARK_ARC_1_0/buf_output[57] )
         );
  XOR2_X1 U11470 ( .A1(n4619), .A2(\MC_ARK_ARC_1_0/temp4[57] ), .Z(n5747) );
  XOR2_X1 U11471 ( .A1(\MC_ARK_ARC_1_0/temp1[57] ), .A2(
        \MC_ARK_ARC_1_0/temp3[57] ), .Z(n5748) );
  NAND4_X2 U11472 ( .A1(\SB2_3_4/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_3_4/Component_Function_0/NAND4_in[2] ), .A3(n6057), .A4(
        \SB2_3_4/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_3_4/buf_output[0] ) );
  XOR2_X1 U11473 ( .A1(\MC_ARK_ARC_1_1/temp5[174] ), .A2(n5749), .Z(
        \MC_ARK_ARC_1_1/buf_output[174] ) );
  XOR2_X1 U11474 ( .A1(\MC_ARK_ARC_1_1/temp3[174] ), .A2(
        \MC_ARK_ARC_1_1/temp4[174] ), .Z(n5749) );
  XOR2_X1 U11475 ( .A1(n5750), .A2(n105), .Z(Ciphertext[89]) );
  NAND4_X2 U11476 ( .A1(n1695), .A2(\SB4_17/Component_Function_5/NAND4_in[1] ), 
        .A3(n4344), .A4(\SB4_17/Component_Function_5/NAND4_in[0] ), .ZN(n5750)
         );
  NAND3_X1 U11477 ( .A1(\SB3_21/i0_4 ), .A2(\SB3_21/i1_7 ), .A3(\SB3_21/i0[8] ), .ZN(\SB3_21/Component_Function_1/NAND4_in[3] ) );
  XOR2_X1 U11478 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[50] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[74] ), .Z(\MC_ARK_ARC_1_2/temp2[104] )
         );
  XOR2_X1 U11479 ( .A1(\RI5[1][183] ), .A2(\RI5[1][15] ), .Z(n5751) );
  NAND4_X2 U11480 ( .A1(\SB1_2_2/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_2/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_2_2/Component_Function_5/NAND4_in[0] ), .A4(n5752), .ZN(
        \SB1_2_2/buf_output[5] ) );
  NAND3_X2 U11481 ( .A1(\SB1_2_2/i0[9] ), .A2(\SB1_2_2/i0_4 ), .A3(
        \SB1_2_2/i0[6] ), .ZN(n5752) );
  NAND4_X2 U11482 ( .A1(\SB1_1_12/Component_Function_5/NAND4_in[3] ), .A2(
        n6328), .A3(n1668), .A4(\SB1_1_12/Component_Function_5/NAND4_in[1] ), 
        .ZN(\SB1_1_12/buf_output[5] ) );
  XOR2_X1 U11483 ( .A1(\RI5[1][83] ), .A2(\RI5[1][137] ), .Z(n5847) );
  NAND3_X1 U11484 ( .A1(\SB1_1_4/i0[10] ), .A2(\SB1_1_4/i0[6] ), .A3(
        \SB1_1_4/i0_0 ), .ZN(\SB1_1_4/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U11485 ( .A1(\SB1_1_8/Component_Function_3/NAND4_in[2] ), .A2(
        \SB1_1_8/Component_Function_3/NAND4_in[3] ), .A3(
        \SB1_1_8/Component_Function_3/NAND4_in[1] ), .A4(
        \SB1_1_8/Component_Function_3/NAND4_in[0] ), .ZN(
        \SB1_1_8/buf_output[3] ) );
  NAND3_X2 U11486 ( .A1(\SB1_2_14/i0_3 ), .A2(\SB1_2_14/i1[9] ), .A3(
        \SB1_2_14/i0_4 ), .ZN(n1847) );
  NAND3_X1 U11487 ( .A1(\SB1_3_31/i0[6] ), .A2(\SB1_3_31/i0_3 ), .A3(
        \SB1_3_31/i1[9] ), .ZN(\SB1_3_31/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U11488 ( .A1(\MC_ARK_ARC_1_1/temp6[41] ), .A2(
        \MC_ARK_ARC_1_1/temp5[41] ), .Z(\MC_ARK_ARC_1_1/buf_output[41] ) );
  NAND3_X1 U11489 ( .A1(\SB4_16/i0_3 ), .A2(\SB4_16/i1_7 ), .A3(\SB4_16/i0[8] ), .ZN(\SB4_16/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U11490 ( .A1(\RI5[1][143] ), .A2(\RI5[1][107] ), .Z(n4495) );
  XOR2_X1 U11491 ( .A1(\MC_ARK_ARC_1_0/temp5[2] ), .A2(n5753), .Z(
        \MC_ARK_ARC_1_0/buf_output[2] ) );
  XOR2_X1 U11492 ( .A1(\MC_ARK_ARC_1_0/temp4[2] ), .A2(
        \MC_ARK_ARC_1_0/temp3[2] ), .Z(n5753) );
  NAND4_X2 U11493 ( .A1(\SB2_1_8/Component_Function_5/NAND4_in[2] ), .A2(n3723), .A3(n1853), .A4(\SB2_1_8/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_1_8/buf_output[5] ) );
  NAND3_X1 U11494 ( .A1(\SB2_1_6/i0[10] ), .A2(\SB2_1_6/i0[6] ), .A3(
        \SB2_1_6/i0_3 ), .ZN(\SB2_1_6/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U11495 ( .A1(\SB2_2_20/i0[6] ), .A2(\SB2_2_20/i0[9] ), .A3(
        \SB2_2_20/i0_4 ), .ZN(n669) );
  NAND4_X2 U11496 ( .A1(n1092), .A2(
        \SB2_0_14/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_0_14/Component_Function_5/NAND4_in[0] ), .A4(n5754), .ZN(
        \SB2_0_14/buf_output[5] ) );
  NAND4_X2 U11497 ( .A1(\SB1_0_29/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_0_29/Component_Function_3/NAND4_in[3] ), .A3(n4631), .A4(n1277), 
        .ZN(\RI3[0][27] ) );
  XOR2_X1 U11498 ( .A1(\RI5[0][107] ), .A2(\RI5[0][173] ), .Z(n6443) );
  NAND3_X2 U11499 ( .A1(\SB2_1_31/i0_0 ), .A2(\SB2_1_31/i0_3 ), .A3(
        \SB2_1_31/i0_4 ), .ZN(\SB2_1_31/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U11500 ( .A1(\SB2_3_2/i0_3 ), .A2(\SB2_3_2/i0_4 ), .A3(
        \SB2_3_2/i1[9] ), .ZN(\SB2_3_2/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U11501 ( .A1(\SB2_0_17/Component_Function_3/NAND4_in[3] ), .A2(
        \SB2_0_17/Component_Function_3/NAND4_in[1] ), .A3(n705), .A4(
        \SB2_0_17/Component_Function_3/NAND4_in[2] ), .ZN(
        \SB2_0_17/buf_output[3] ) );
  XOR2_X1 U11502 ( .A1(n5758), .A2(n5757), .Z(\MC_ARK_ARC_1_0/buf_output[122] ) );
  XOR2_X1 U11503 ( .A1(\MC_ARK_ARC_1_0/temp3[122] ), .A2(n4665), .Z(n5757) );
  XOR2_X1 U11504 ( .A1(\MC_ARK_ARC_1_0/temp1[122] ), .A2(
        \MC_ARK_ARC_1_0/temp4[122] ), .Z(n5758) );
  XOR2_X1 U11505 ( .A1(\MC_ARK_ARC_1_2/temp4[121] ), .A2(n5759), .Z(n3737) );
  XOR2_X1 U11506 ( .A1(\RI5[2][187] ), .A2(\RI5[2][31] ), .Z(n5759) );
  XOR2_X1 U11507 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[185] ), .A2(
        \MC_ARK_ARC_1_2/buf_keyinput[54] ), .Z(n5760) );
  NAND3_X1 U11508 ( .A1(\SB1_3_21/i0[10] ), .A2(\SB1_3_21/i1[9] ), .A3(
        \SB1_3_21/i1_5 ), .ZN(n5761) );
  NAND4_X2 U11509 ( .A1(\SB2_2_4/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_2_4/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_2_4/Component_Function_1/NAND4_in[0] ), .A4(n5762), .ZN(
        \SB2_2_4/buf_output[1] ) );
  NAND4_X2 U11510 ( .A1(\SB1_2_14/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_14/Component_Function_0/NAND4_in[1] ), .A3(n4578), .A4(
        \SB1_2_14/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_2_14/buf_output[0] ) );
  XOR2_X1 U11511 ( .A1(\MC_ARK_ARC_1_1/temp4[113] ), .A2(n5763), .Z(n5917) );
  XOR2_X1 U11512 ( .A1(\RI5[1][107] ), .A2(\RI5[1][59] ), .Z(n5763) );
  AND2_X1 U11513 ( .A1(\SB2_1_5/Component_Function_3/NAND4_in[3] ), .A2(n1558), 
        .Z(n5764) );
  XOR2_X1 U11514 ( .A1(\RI5[3][87] ), .A2(n1392), .Z(n4313) );
  XOR2_X1 U11515 ( .A1(\MC_ARK_ARC_1_3/temp1[151] ), .A2(n5765), .Z(
        \MC_ARK_ARC_1_3/temp5[151] ) );
  XOR2_X1 U11516 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[97] ), .A2(\RI5[3][121] ), 
        .Z(n5765) );
  NAND4_X2 U11517 ( .A1(\SB2_1_27/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_1_27/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_1_27/Component_Function_1/NAND4_in[0] ), .A4(n5766), .ZN(
        \SB2_1_27/buf_output[1] ) );
  NAND3_X1 U11518 ( .A1(\SB1_1_28/buf_output[4] ), .A2(\SB2_1_27/i1_7 ), .A3(
        \SB2_1_27/i0[8] ), .ZN(n5766) );
  NAND3_X1 U11519 ( .A1(\SB4_0/i0_4 ), .A2(n1386), .A3(\SB4_0/i1_5 ), .ZN(
        n5767) );
  XOR2_X1 U11520 ( .A1(\MC_ARK_ARC_1_0/temp2[67] ), .A2(n5768), .Z(
        \MC_ARK_ARC_1_0/temp5[67] ) );
  XOR2_X1 U11521 ( .A1(\SB2_0_24/buf_output[1] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[61] ), .Z(n5768) );
  XOR2_X1 U11522 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[61] ), .A2(\RI5[0][97] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[187] ) );
  NAND4_X2 U11523 ( .A1(\SB1_1_10/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_10/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_1_10/Component_Function_2/NAND4_in[3] ), .A4(n6018), .ZN(
        \SB1_1_10/buf_output[2] ) );
  XOR2_X1 U11524 ( .A1(\RI5[0][128] ), .A2(\RI5[0][98] ), .Z(n4081) );
  NAND3_X1 U11525 ( .A1(\SB1_1_28/i0_0 ), .A2(\SB1_1_28/i3[0] ), .A3(
        \SB1_1_28/i1_7 ), .ZN(\SB1_1_28/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U11526 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[136] ), .A2(\RI5[2][172] ), .Z(\MC_ARK_ARC_1_2/temp3[70] ) );
  XOR2_X1 U11527 ( .A1(\RI5[2][134] ), .A2(\RI5[2][140] ), .Z(
        \MC_ARK_ARC_1_2/temp1[140] ) );
  NAND3_X1 U11528 ( .A1(\SB3_1/i0_4 ), .A2(n4765), .A3(\SB3_1/i1_5 ), .ZN(
        \SB3_1/Component_Function_4/NAND4_in[3] ) );
  XOR2_X1 U11529 ( .A1(n5769), .A2(n89), .Z(Ciphertext[150]) );
  NAND4_X2 U11530 ( .A1(\SB4_6/Component_Function_0/NAND4_in[3] ), .A2(
        \SB4_6/Component_Function_0/NAND4_in[1] ), .A3(
        \SB4_6/Component_Function_0/NAND4_in[0] ), .A4(n3461), .ZN(n5769) );
  XOR2_X1 U11531 ( .A1(n3777), .A2(\MC_ARK_ARC_1_1/temp4[52] ), .Z(n2812) );
  NAND4_X2 U11532 ( .A1(\SB1_3_16/Component_Function_2/NAND4_in[1] ), .A2(
        n6037), .A3(\SB1_3_16/Component_Function_2/NAND4_in[0] ), .A4(n5770), 
        .ZN(\SB1_3_16/buf_output[2] ) );
  INV_X2 U11533 ( .I(\SB1_3_9/buf_output[2] ), .ZN(\SB2_3_6/i1[9] ) );
  NAND4_X2 U11534 ( .A1(n878), .A2(\SB3_21/Component_Function_2/NAND4_in[0] ), 
        .A3(n4002), .A4(n5771), .ZN(\SB3_21/buf_output[2] ) );
  XOR2_X1 U11535 ( .A1(n3010), .A2(n5772), .Z(n3018) );
  NAND4_X2 U11536 ( .A1(n2097), .A2(\SB1_2_8/Component_Function_5/NAND4_in[1] ), .A3(n976), .A4(\SB1_2_8/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_2_8/buf_output[5] ) );
  NAND4_X2 U11537 ( .A1(n4688), .A2(
        \SB2_3_14/Component_Function_5/NAND4_in[0] ), .A3(n6043), .A4(
        \SB2_3_14/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB2_3_14/buf_output[5] ) );
  CLKBUF_X12 U11538 ( .I(\SB1_2_4/buf_output[3] ), .Z(n5818) );
  XOR2_X1 U11539 ( .A1(\MC_ARK_ARC_1_2/temp6[82] ), .A2(n5773), .Z(
        \MC_ARK_ARC_1_2/buf_output[82] ) );
  XOR2_X1 U11540 ( .A1(\MC_ARK_ARC_1_2/temp2[82] ), .A2(
        \MC_ARK_ARC_1_2/temp1[82] ), .Z(n5773) );
  NAND3_X2 U11541 ( .A1(\SB1_3_9/i0[10] ), .A2(\SB1_3_9/i0[6] ), .A3(
        \SB1_3_9/i0_0 ), .ZN(\SB1_3_9/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U11542 ( .A1(\SB2_2_11/Component_Function_3/NAND4_in[0] ), .A2(
        n2451), .A3(\SB2_2_11/Component_Function_3/NAND4_in[2] ), .A4(n5774), 
        .ZN(\SB2_2_11/buf_output[3] ) );
  NAND3_X2 U11543 ( .A1(\SB2_2_11/i0_4 ), .A2(\SB2_2_11/i0_0 ), .A3(
        \SB2_2_11/i0_3 ), .ZN(n5774) );
  XOR2_X1 U11544 ( .A1(n5775), .A2(n76), .Z(Ciphertext[20]) );
  INV_X2 U11545 ( .I(\SB1_1_9/buf_output[2] ), .ZN(\SB2_1_6/i1[9] ) );
  NAND4_X2 U11546 ( .A1(\SB1_1_9/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_1_9/Component_Function_2/NAND4_in[1] ), .A3(n3369), .A4(n1221), 
        .ZN(\SB1_1_9/buf_output[2] ) );
  XOR2_X1 U11547 ( .A1(n5777), .A2(\MC_ARK_ARC_1_1/temp4[99] ), .Z(n2250) );
  NAND3_X2 U11548 ( .A1(\SB2_0_18/i0[10] ), .A2(\SB2_0_18/i1[9] ), .A3(
        \SB2_0_18/i1_7 ), .ZN(\SB2_0_18/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U11549 ( .A1(\SB4_29/i0[6] ), .A2(\SB4_29/i0[7] ), .A3(
        \SB4_29/i0[8] ), .ZN(n5778) );
  NAND4_X2 U11550 ( .A1(\SB2_0_21/Component_Function_2/NAND4_in[1] ), .A2(
        n1674), .A3(\SB2_0_21/Component_Function_2/NAND4_in[0] ), .A4(
        \SB2_0_21/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_0_21/buf_output[2] ) );
  XOR2_X1 U11551 ( .A1(\MC_ARK_ARC_1_1/temp6[39] ), .A2(n864), .Z(
        \MC_ARK_ARC_1_1/buf_output[39] ) );
  NAND4_X2 U11552 ( .A1(\SB1_2_25/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_2_25/Component_Function_1/NAND4_in[1] ), .A3(n5926), .A4(
        \SB1_2_25/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_2_25/buf_output[1] ) );
  NAND4_X2 U11553 ( .A1(n3614), .A2(\SB1_2_6/Component_Function_5/NAND4_in[1] ), .A3(\SB1_2_6/Component_Function_5/NAND4_in[0] ), .A4(n5780), .ZN(
        \SB1_2_6/buf_output[5] ) );
  NAND3_X2 U11554 ( .A1(\SB1_2_6/i0[9] ), .A2(\SB1_2_6/i0[6] ), .A3(
        \SB1_2_6/i0_4 ), .ZN(n5780) );
  XOR2_X1 U11555 ( .A1(\RI5[0][80] ), .A2(\RI5[0][104] ), .Z(
        \MC_ARK_ARC_1_0/temp2[134] ) );
  XOR2_X1 U11556 ( .A1(n740), .A2(\MC_ARK_ARC_1_3/temp6[180] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[180] ) );
  XOR2_X1 U11557 ( .A1(\RI5[2][41] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[65] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[95] ) );
  NAND4_X2 U11558 ( .A1(\SB3_23/Component_Function_5/NAND4_in[1] ), .A2(n954), 
        .A3(\SB3_23/Component_Function_5/NAND4_in[2] ), .A4(n5781), .ZN(
        \SB3_23/buf_output[5] ) );
  XOR2_X1 U11559 ( .A1(\MC_ARK_ARC_1_1/temp5[17] ), .A2(n2391), .Z(
        \MC_ARK_ARC_1_1/buf_output[17] ) );
  NAND4_X2 U11560 ( .A1(\SB2_2_2/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_2/Component_Function_5/NAND4_in[1] ), .A3(n5813), .A4(n1469), 
        .ZN(\SB2_2_2/buf_output[5] ) );
  XOR2_X1 U11561 ( .A1(\RI5[2][179] ), .A2(\RI5[2][155] ), .Z(n5782) );
  NAND4_X2 U11562 ( .A1(\SB2_1_6/Component_Function_5/NAND4_in[1] ), .A2(n2392), .A3(\SB2_1_6/Component_Function_5/NAND4_in[0] ), .A4(n6298), .ZN(
        \SB2_1_6/buf_output[5] ) );
  NAND4_X2 U11563 ( .A1(\SB4_0/Component_Function_0/NAND4_in[2] ), .A2(
        \SB4_0/Component_Function_0/NAND4_in[1] ), .A3(n3868), .A4(
        \SB4_0/Component_Function_0/NAND4_in[0] ), .ZN(n6272) );
  NAND3_X2 U11564 ( .A1(\SB3_1/i0[9] ), .A2(\SB3_1/i0_4 ), .A3(\SB3_1/i0[6] ), 
        .ZN(n6280) );
  XOR2_X1 U11565 ( .A1(\MC_ARK_ARC_1_2/temp6[185] ), .A2(n5783), .Z(
        \MC_ARK_ARC_1_2/buf_output[185] ) );
  XOR2_X1 U11566 ( .A1(n6508), .A2(n2574), .Z(n5783) );
  NAND3_X2 U11567 ( .A1(\SB2_2_11/i0_4 ), .A2(\SB2_2_11/i0_0 ), .A3(
        \SB2_2_11/i1_5 ), .ZN(n5784) );
  NOR2_X2 U11568 ( .A1(n1707), .A2(n5786), .ZN(\SB2_2_13/i0[7] ) );
  NAND2_X2 U11569 ( .A1(n5921), .A2(n1706), .ZN(n5786) );
  XOR2_X1 U11570 ( .A1(n6326), .A2(n5787), .Z(\MC_ARK_ARC_1_2/buf_output[146] ) );
  NAND2_X2 U11571 ( .A1(\SB1_0_8/Component_Function_2/NAND4_in[2] ), .A2(n2750), .ZN(n5789) );
  NAND3_X1 U11572 ( .A1(\SB4_30/i0_3 ), .A2(\SB4_30/i0[9] ), .A3(
        \SB4_30/i0[8] ), .ZN(\SB4_30/Component_Function_2/NAND4_in[2] ) );
  NAND4_X2 U11573 ( .A1(\SB3_0/Component_Function_3/NAND4_in[1] ), .A2(n6108), 
        .A3(n3282), .A4(n5791), .ZN(\SB3_0/buf_output[3] ) );
  NAND4_X2 U11574 ( .A1(\SB1_2_2/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_2/Component_Function_3/NAND4_in[2] ), .A3(
        \SB1_2_2/Component_Function_3/NAND4_in[1] ), .A4(n5792), .ZN(
        \SB1_2_2/buf_output[3] ) );
  NAND3_X2 U11575 ( .A1(\SB1_2_2/i3[0] ), .A2(\SB1_2_2/i0[8] ), .A3(
        \SB1_2_2/i1_5 ), .ZN(n5792) );
  NAND3_X2 U11576 ( .A1(\SB2_2_0/i0[10] ), .A2(\SB2_2_0/i0_0 ), .A3(
        \SB2_2_0/i0[6] ), .ZN(n1609) );
  XOR2_X1 U11577 ( .A1(\MC_ARK_ARC_1_0/temp6[142] ), .A2(n5793), .Z(
        \MC_ARK_ARC_1_0/buf_output[142] ) );
  XOR2_X1 U11578 ( .A1(\MC_ARK_ARC_1_0/temp1[142] ), .A2(
        \MC_ARK_ARC_1_0/temp2[142] ), .Z(n5793) );
  NAND4_X2 U11579 ( .A1(\SB3_5/Component_Function_0/NAND4_in[1] ), .A2(
        \SB3_5/Component_Function_0/NAND4_in[2] ), .A3(
        \SB3_5/Component_Function_0/NAND4_in[0] ), .A4(n5794), .ZN(
        \SB3_5/buf_output[0] ) );
  NAND3_X2 U11580 ( .A1(\SB1_0_29/i0_0 ), .A2(\SB1_0_29/i0[10] ), .A3(
        \SB1_0_29/i0[6] ), .ZN(n5795) );
  NAND3_X1 U11581 ( .A1(\SB2_2_8/i0_4 ), .A2(\SB2_2_8/i1[9] ), .A3(
        \SB1_2_8/buf_output[5] ), .ZN(
        \SB2_2_8/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U11582 ( .A1(\SB2_2_10/i0_0 ), .A2(\SB2_2_10/i0_3 ), .A3(n581), 
        .ZN(\SB2_2_10/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U11583 ( .A1(\MC_ARK_ARC_1_1/temp1[14] ), .A2(n5797), .Z(
        \MC_ARK_ARC_1_1/temp5[14] ) );
  XOR2_X1 U11584 ( .A1(\RI5[1][152] ), .A2(\RI5[1][176] ), .Z(n5797) );
  NAND4_X2 U11585 ( .A1(\SB3_30/Component_Function_3/NAND4_in[1] ), .A2(n807), 
        .A3(n3451), .A4(n5798), .ZN(\SB3_30/buf_output[3] ) );
  XOR2_X1 U11586 ( .A1(\MC_ARK_ARC_1_0/temp2[154] ), .A2(n5799), .Z(
        \MC_ARK_ARC_1_0/temp5[154] ) );
  XOR2_X1 U11587 ( .A1(\RI5[0][148] ), .A2(\RI5[0][154] ), .Z(n5799) );
  XOR2_X1 U11588 ( .A1(n5847), .A2(n5800), .Z(\MC_ARK_ARC_1_1/temp5[137] ) );
  XOR2_X1 U11589 ( .A1(\RI5[1][107] ), .A2(\RI5[1][131] ), .Z(n5800) );
  NAND3_X1 U11590 ( .A1(\SB2_3_0/i0_3 ), .A2(\SB2_3_0/i0_0 ), .A3(
        \SB1_3_1/buf_output[4] ), .ZN(
        \SB2_3_0/Component_Function_3/NAND4_in[1] ) );
  INV_X2 U11591 ( .I(\SB1_2_30/buf_output[3] ), .ZN(\SB2_2_28/i0[8] ) );
  XOR2_X1 U11592 ( .A1(n5801), .A2(n6090), .Z(n6110) );
  XOR2_X1 U11593 ( .A1(\SB2_0_7/buf_output[3] ), .A2(\RI5[0][153] ), .Z(n5801)
         );
  XOR2_X1 U11594 ( .A1(n6060), .A2(n3547), .Z(n2028) );
  NAND3_X2 U11595 ( .A1(\SB2_2_12/i0_4 ), .A2(\SB2_2_12/i0[6] ), .A3(
        \SB2_2_12/i0[9] ), .ZN(n5802) );
  NAND3_X2 U11596 ( .A1(\SB2_0_14/i0[8] ), .A2(\SB2_0_14/i0[9] ), .A3(
        \SB2_0_14/i0_3 ), .ZN(\SB2_0_14/Component_Function_2/NAND4_in[2] ) );
  NAND3_X2 U11597 ( .A1(\SB2_1_6/i0_0 ), .A2(\SB2_1_6/i0_4 ), .A3(
        \SB2_1_6/i1_5 ), .ZN(n5803) );
  AND2_X1 U11598 ( .A1(n2520), .A2(n5804), .Z(n6185) );
  NAND3_X1 U11599 ( .A1(\SB1_3_17/i0[7] ), .A2(\SB1_3_17/i0[8] ), .A3(
        \SB1_3_17/i0[6] ), .ZN(n5804) );
  XOR2_X1 U11600 ( .A1(\MC_ARK_ARC_1_3/temp1[154] ), .A2(
        \MC_ARK_ARC_1_3/temp2[154] ), .Z(\MC_ARK_ARC_1_3/temp5[154] ) );
  XOR2_X1 U11601 ( .A1(\RI5[1][164] ), .A2(\RI5[1][140] ), .Z(n5911) );
  XOR2_X1 U11602 ( .A1(\RI5[2][1] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[7] ), 
        .Z(\MC_ARK_ARC_1_2/temp1[7] ) );
  NAND3_X1 U11603 ( .A1(\SB1_0_18/i1[9] ), .A2(\SB1_0_18/i1_5 ), .A3(n1367), 
        .ZN(\SB1_0_18/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U11604 ( .A1(\SB1_3_30/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_30/Component_Function_5/NAND4_in[2] ), .A3(n5824), .A4(
        \SB1_3_30/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_30/buf_output[5] ) );
  NAND4_X2 U11605 ( .A1(\SB2_0_15/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_15/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_0_15/Component_Function_2/NAND4_in[1] ), .A4(n5805), .ZN(
        \SB2_0_15/buf_output[2] ) );
  XOR2_X1 U11606 ( .A1(n2184), .A2(n5806), .Z(\MC_ARK_ARC_1_2/buf_output[120] ) );
  XOR2_X1 U11607 ( .A1(n5807), .A2(n6102), .Z(\MC_ARK_ARC_1_1/buf_output[40] )
         );
  NAND3_X1 U11608 ( .A1(\SB2_0_27/i0_4 ), .A2(\SB2_0_27/i1[9] ), .A3(
        \SB2_0_27/i1_5 ), .ZN(\SB2_0_27/Component_Function_4/NAND4_in[3] ) );
  NAND4_X2 U11609 ( .A1(\SB2_3_23/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_3_23/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_3_23/Component_Function_0/NAND4_in[0] ), .A4(n5810), .ZN(
        \SB2_3_23/buf_output[0] ) );
  NAND3_X2 U11610 ( .A1(\SB2_3_23/i0_3 ), .A2(\SB2_3_23/i0_0 ), .A3(
        \SB2_3_23/i0[7] ), .ZN(n5810) );
  XOR2_X1 U11611 ( .A1(n2461), .A2(n5811), .Z(\MC_ARK_ARC_1_3/buf_output[26] )
         );
  XOR2_X1 U11612 ( .A1(n1925), .A2(n3051), .Z(n5811) );
  XOR2_X1 U11613 ( .A1(n5812), .A2(\MC_ARK_ARC_1_1/temp6[76] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[76] ) );
  XOR2_X1 U11614 ( .A1(\MC_ARK_ARC_1_1/temp1[76] ), .A2(
        \MC_ARK_ARC_1_1/temp2[76] ), .Z(n5812) );
  NAND3_X2 U11615 ( .A1(\SB1_2_3/buf_output[4] ), .A2(\SB2_2_2/i0[6] ), .A3(
        \SB2_2_2/i0[9] ), .ZN(n5813) );
  NAND4_X2 U11616 ( .A1(\SB1_2_6/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_2_6/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_6/Component_Function_1/NAND4_in[0] ), .A4(n5814), .ZN(
        \SB1_2_6/buf_output[1] ) );
  NAND3_X1 U11617 ( .A1(\SB1_2_6/i0[8] ), .A2(\SB1_2_6/i0_4 ), .A3(
        \SB1_2_6/i1_7 ), .ZN(n5814) );
  XOR2_X1 U11618 ( .A1(\MC_ARK_ARC_1_1/temp2[68] ), .A2(n5815), .Z(
        \MC_ARK_ARC_1_1/temp5[68] ) );
  XOR2_X1 U11619 ( .A1(\RI5[1][68] ), .A2(\RI5[1][62] ), .Z(n5815) );
  INV_X2 U11620 ( .I(\RI3[0][92] ), .ZN(\SB2_0_16/i1[9] ) );
  NAND4_X2 U11621 ( .A1(\SB1_0_19/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_19/Component_Function_2/NAND4_in[3] ), .A3(n1287), .A4(
        \SB1_0_19/Component_Function_2/NAND4_in[2] ), .ZN(\RI3[0][92] ) );
  XOR2_X1 U11622 ( .A1(\MC_ARK_ARC_1_3/temp2[1] ), .A2(n5816), .Z(n6453) );
  XOR2_X1 U11623 ( .A1(\RI5[3][187] ), .A2(\RI5[3][1] ), .Z(n5816) );
  NAND2_X2 U11624 ( .A1(\SB1_2_7/i0_0 ), .A2(\SB1_2_7/i3[0] ), .ZN(n5939) );
  NAND2_X1 U11625 ( .A1(\SB1_0_6/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_0_6/Component_Function_4/NAND4_in[0] ), .ZN(n5857) );
  NAND3_X1 U11626 ( .A1(\SB4_6/i0_0 ), .A2(\SB4_6/i1_7 ), .A3(\SB4_6/i3[0] ), 
        .ZN(n5817) );
  INV_X4 U11627 ( .I(n5818), .ZN(\SB2_2_2/i0[8] ) );
  NAND3_X2 U11628 ( .A1(\SB1_2_4/i0[6] ), .A2(\SB1_2_4/i0_3 ), .A3(
        \SB1_2_4/i1[9] ), .ZN(\SB1_2_4/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U11629 ( .A1(\SB2_1_8/i0[6] ), .A2(\SB1_1_13/buf_output[0] ), .A3(
        \SB2_1_8/i1_5 ), .ZN(\SB2_1_8/Component_Function_1/NAND4_in[2] ) );
  NAND4_X2 U11630 ( .A1(\SB2_1_26/Component_Function_2/NAND4_in[0] ), .A2(
        n6273), .A3(n3778), .A4(\SB2_1_26/Component_Function_2/NAND4_in[2] ), 
        .ZN(\SB2_1_26/buf_output[2] ) );
  NAND4_X2 U11631 ( .A1(\SB2_2_2/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_2_2/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_2/Component_Function_1/NAND4_in[0] ), .A4(
        \SB2_2_2/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_2_2/buf_output[1] ) );
  XOR2_X1 U11632 ( .A1(n4614), .A2(n6424), .Z(\MC_ARK_ARC_1_1/buf_output[163] ) );
  NAND4_X2 U11633 ( .A1(n3035), .A2(\SB1_1_7/Component_Function_4/NAND4_in[1] ), .A3(\SB1_1_7/Component_Function_4/NAND4_in[3] ), .A4(n5819), .ZN(
        \SB1_1_7/buf_output[4] ) );
  XOR2_X1 U11634 ( .A1(\MC_ARK_ARC_1_0/temp5[146] ), .A2(n5820), .Z(
        \MC_ARK_ARC_1_0/buf_output[146] ) );
  XOR2_X1 U11635 ( .A1(n3293), .A2(n3294), .Z(n5820) );
  NAND4_X2 U11636 ( .A1(\SB2_0_19/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_19/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_0_19/Component_Function_2/NAND4_in[3] ), .A4(n5821), .ZN(
        \SB2_0_19/buf_output[2] ) );
  NAND3_X2 U11637 ( .A1(\SB2_0_19/i0_3 ), .A2(\SB2_0_19/i0[9] ), .A3(
        \SB2_0_19/i0[8] ), .ZN(n5821) );
  XOR2_X1 U11638 ( .A1(n5823), .A2(n5822), .Z(\MC_ARK_ARC_1_2/temp5[6] ) );
  XOR2_X1 U11639 ( .A1(\RI5[2][144] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[6] ), 
        .Z(n5822) );
  XOR2_X1 U11640 ( .A1(\RI5[2][168] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[0] ), 
        .Z(n5823) );
  NAND3_X2 U11641 ( .A1(\SB1_3_30/i0[9] ), .A2(\SB1_3_30/i0[6] ), .A3(
        \SB1_3_30/i0_4 ), .ZN(n5824) );
  INV_X2 U11642 ( .I(\SB3_11/buf_output[2] ), .ZN(\SB4_8/i1[9] ) );
  XOR2_X1 U11643 ( .A1(n6029), .A2(n5825), .Z(\MC_ARK_ARC_1_0/buf_output[53] )
         );
  XOR2_X1 U11644 ( .A1(n6265), .A2(\MC_ARK_ARC_1_0/temp4[53] ), .Z(n5825) );
  BUF_X2 U11645 ( .I(n4749), .Z(n5826) );
  NAND4_X2 U11646 ( .A1(\SB1_0_21/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_0_21/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_21/Component_Function_1/NAND4_in[3] ), .A4(
        \SB1_0_21/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_0_21/buf_output[1] ) );
  NAND3_X1 U11647 ( .A1(\SB1_2_12/i0_3 ), .A2(\SB1_2_12/i0_0 ), .A3(
        \SB1_2_12/i0[7] ), .ZN(\SB1_2_12/Component_Function_0/NAND4_in[3] ) );
  NAND3_X2 U11648 ( .A1(\SB2_1_14/i0_3 ), .A2(\SB2_1_14/i0_4 ), .A3(
        \SB2_1_14/i1[9] ), .ZN(\SB2_1_14/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U11649 ( .A1(\SB3_9/Component_Function_1/NAND4_in[3] ), .A2(
        \SB3_9/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_9/Component_Function_1/NAND4_in[0] ), .A4(n5828), .ZN(
        \SB3_9/buf_output[1] ) );
  NAND3_X1 U11650 ( .A1(\SB3_9/i0[9] ), .A2(\SB3_9/i0[6] ), .A3(\SB3_9/i1_5 ), 
        .ZN(n5828) );
  NAND4_X2 U11651 ( .A1(n3695), .A2(
        \SB2_1_31/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_1_31/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_1_31/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_1_31/buf_output[5] ) );
  XOR2_X1 U11652 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[44] ), .A2(\RI5[0][50] ), 
        .Z(n5829) );
  NAND3_X2 U11653 ( .A1(\SB1_1_17/i0[10] ), .A2(\SB1_1_17/i0_3 ), .A3(
        \SB1_1_17/i0[6] ), .ZN(n1984) );
  NAND3_X2 U11654 ( .A1(\SB1_2_13/i1_5 ), .A2(\SB1_2_13/i0[8] ), .A3(
        \SB1_2_13/i3[0] ), .ZN(\SB1_2_13/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U11655 ( .A1(\RI5[1][30] ), .A2(\RI5[1][36] ), .Z(
        \MC_ARK_ARC_1_1/temp1[36] ) );
  NAND4_X2 U11656 ( .A1(\SB2_3_20/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_3_20/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_20/Component_Function_3/NAND4_in[3] ), .A4(n5830), .ZN(
        \SB2_3_20/buf_output[3] ) );
  NAND3_X2 U11657 ( .A1(\SB2_3_20/i0[10] ), .A2(\SB2_3_20/i1[9] ), .A3(
        \SB2_3_20/i1_7 ), .ZN(n5830) );
  NAND3_X2 U11658 ( .A1(\SB2_1_1/i0_4 ), .A2(\SB2_1_1/i0_0 ), .A3(
        \SB2_1_1/i1_5 ), .ZN(n3244) );
  NAND3_X2 U11659 ( .A1(\SB2_2_2/i0_3 ), .A2(\SB2_2_2/i0[9] ), .A3(
        \SB2_2_2/i0[8] ), .ZN(\SB2_2_2/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U11660 ( .A1(\SB4_6/i0_3 ), .A2(\SB4_6/i0[6] ), .A3(\SB4_6/i1[9] ), 
        .ZN(n821) );
  NAND4_X2 U11661 ( .A1(\SB3_31/Component_Function_3/NAND4_in[1] ), .A2(
        \SB3_31/Component_Function_3/NAND4_in[0] ), .A3(n2072), .A4(
        \SB3_31/Component_Function_3/NAND4_in[3] ), .ZN(\SB3_31/buf_output[3] ) );
  NAND2_X1 U11662 ( .A1(\SB1_3_7/i1[9] ), .A2(\SB1_3_7/i0_3 ), .ZN(
        \SB1_3_7/Component_Function_1/NAND4_in[0] ) );
  XOR2_X1 U11663 ( .A1(\RI5[2][64] ), .A2(\RI5[2][88] ), .Z(
        \MC_ARK_ARC_1_2/temp2[118] ) );
  NAND4_X2 U11664 ( .A1(\SB1_1_31/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_31/Component_Function_5/NAND4_in[3] ), .A3(n6024), .A4(
        \SB1_1_31/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_31/buf_output[5] ) );
  XOR2_X1 U11665 ( .A1(\MC_ARK_ARC_1_0/temp2[4] ), .A2(n5831), .Z(
        \MC_ARK_ARC_1_0/temp5[4] ) );
  XOR2_X1 U11666 ( .A1(\RI5[0][190] ), .A2(\RI5[0][4] ), .Z(n5831) );
  XOR2_X1 U11667 ( .A1(\RI5[2][9] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[45] ), 
        .Z(\MC_ARK_ARC_1_2/temp3[135] ) );
  XOR2_X1 U11668 ( .A1(\RI5[1][165] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[159] ), .Z(\MC_ARK_ARC_1_1/temp1[165] ) );
  XOR2_X1 U11669 ( .A1(n3784), .A2(n6493), .Z(\MC_ARK_ARC_1_0/buf_output[176] ) );
  NAND2_X1 U11670 ( .A1(n2444), .A2(n1201), .ZN(n1014) );
  NAND4_X2 U11671 ( .A1(\SB1_3_12/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_3_12/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_3_12/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_3_12/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_3_12/buf_output[0] ) );
  NAND4_X2 U11672 ( .A1(\SB1_0_28/Component_Function_5/NAND4_in[1] ), .A2(
        n6249), .A3(\SB1_0_28/Component_Function_5/NAND4_in[0] ), .A4(
        \SB1_0_28/Component_Function_5/NAND4_in[3] ), .ZN(\RI3[0][23] ) );
  NAND3_X1 U11673 ( .A1(\SB2_2_9/i0_3 ), .A2(\SB2_2_9/i0[10] ), .A3(
        \SB2_2_9/i0_4 ), .ZN(\SB2_2_9/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U11674 ( .A1(n2886), .A2(\MC_ARK_ARC_1_3/temp5[129] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[129] ) );
  NAND3_X1 U11675 ( .A1(\SB1_3_7/i0_0 ), .A2(\SB1_3_7/i0[9] ), .A3(
        \SB1_3_7/i0[8] ), .ZN(\SB1_3_7/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U11676 ( .A1(\SB4_5/i0[6] ), .A2(\SB4_5/i0[8] ), .A3(\SB4_5/i0[7] ), 
        .ZN(\SB4_5/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U11677 ( .A1(\SB1_0_20/i0_0 ), .A2(\SB1_0_20/i0_4 ), .A3(
        \SB1_0_20/i0_3 ), .ZN(\SB1_0_20/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U11678 ( .A1(\SB2_0_7/Component_Function_2/NAND4_in[1] ), .A2(n6484), .A3(\SB2_0_7/Component_Function_2/NAND4_in[0] ), .A4(n4292), .ZN(
        \SB2_0_7/buf_output[2] ) );
  INV_X4 U11679 ( .I(n5832), .ZN(\RI3[0][147] ) );
  NOR2_X2 U11680 ( .A1(n5931), .A2(n5833), .ZN(n5832) );
  NAND2_X2 U11681 ( .A1(n3897), .A2(\SB1_0_9/Component_Function_3/NAND4_in[3] ), .ZN(n5833) );
  XOR2_X1 U11682 ( .A1(n5834), .A2(n4465), .Z(n2233) );
  XOR2_X1 U11683 ( .A1(\RI5[0][68] ), .A2(\RI5[0][98] ), .Z(n5834) );
  XOR2_X1 U11684 ( .A1(n5835), .A2(n172), .Z(Ciphertext[81]) );
  NAND4_X2 U11685 ( .A1(\SB4_18/Component_Function_3/NAND4_in[1] ), .A2(
        \SB4_18/Component_Function_3/NAND4_in[3] ), .A3(n3480), .A4(
        \SB4_18/Component_Function_3/NAND4_in[2] ), .ZN(n5835) );
  XOR2_X1 U11686 ( .A1(n1797), .A2(\MC_ARK_ARC_1_2/temp1[175] ), .Z(n5836) );
  XOR2_X1 U11687 ( .A1(\MC_ARK_ARC_1_1/temp2[126] ), .A2(n5837), .Z(n2161) );
  XOR2_X1 U11688 ( .A1(\RI5[1][0] ), .A2(\RI5[1][36] ), .Z(n5837) );
  NAND4_X2 U11689 ( .A1(\SB3_8/Component_Function_4/NAND4_in[3] ), .A2(
        \SB3_8/Component_Function_4/NAND4_in[0] ), .A3(
        \SB3_8/Component_Function_4/NAND4_in[1] ), .A4(n5838), .ZN(
        \SB3_8/buf_output[4] ) );
  NAND3_X1 U11690 ( .A1(\SB4_7/i0_4 ), .A2(\SB4_7/i0_0 ), .A3(\SB4_7/i1_5 ), 
        .ZN(n5839) );
  AND2_X1 U11691 ( .A1(\SB3_8/Component_Function_3/NAND4_in[2] ), .A2(n2113), 
        .Z(n5840) );
  AND2_X1 U11692 ( .A1(\SB3_8/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_8/Component_Function_3/NAND4_in[1] ), .Z(n5841) );
  INV_X1 U11693 ( .I(\SB3_9/buf_output[2] ), .ZN(\SB4_6/i1[9] ) );
  NAND4_X2 U11694 ( .A1(\SB3_9/Component_Function_2/NAND4_in[2] ), .A2(n5851), 
        .A3(\SB3_9/Component_Function_2/NAND4_in[1] ), .A4(
        \SB3_9/Component_Function_2/NAND4_in[0] ), .ZN(\SB3_9/buf_output[2] )
         );
  XOR2_X1 U11695 ( .A1(n5842), .A2(\MC_ARK_ARC_1_1/temp4[85] ), .Z(
        \MC_ARK_ARC_1_1/temp6[85] ) );
  NAND3_X2 U11696 ( .A1(\SB2_0_22/i0_3 ), .A2(\SB2_0_22/i0[6] ), .A3(
        \SB2_0_22/i1[9] ), .ZN(\SB2_0_22/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U11697 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[31] ), .A2(\RI5[1][55] ), 
        .Z(\MC_ARK_ARC_1_1/temp2[85] ) );
  NAND4_X2 U11698 ( .A1(\SB1_0_16/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_0_16/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_0_16/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_0_16/Component_Function_0/NAND4_in[0] ), .ZN(\SB2_0_11/i0[9] ) );
  NAND3_X1 U11699 ( .A1(\SB2_1_14/i0_0 ), .A2(\SB2_1_14/i0[9] ), .A3(
        \SB2_1_14/i0[8] ), .ZN(\SB2_1_14/Component_Function_4/NAND4_in[0] ) );
  NAND3_X1 U11700 ( .A1(\SB3_10/i0_4 ), .A2(\SB3_10/i1[9] ), .A3(\SB3_10/i1_5 ), .ZN(\SB3_10/Component_Function_4/NAND4_in[3] ) );
  NAND3_X1 U11701 ( .A1(\SB1_2_4/i0[10] ), .A2(\SB1_2_4/i1[9] ), .A3(
        \SB1_2_4/i1_7 ), .ZN(n6126) );
  NAND3_X2 U11702 ( .A1(\SB2_2_9/i0[9] ), .A2(\SB2_2_9/i0_3 ), .A3(
        \SB2_2_9/i0[8] ), .ZN(\SB2_2_9/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U11703 ( .A1(\SB2_2_3/i0_3 ), .A2(\SB1_2_8/buf_output[0] ), .A3(
        \SB2_2_3/i0[8] ), .ZN(\SB2_2_3/Component_Function_2/NAND4_in[2] ) );
  XOR2_X1 U11704 ( .A1(\RI5[0][189] ), .A2(\RI5[0][33] ), .Z(
        \MC_ARK_ARC_1_0/temp3[123] ) );
  NAND4_X2 U11705 ( .A1(n1742), .A2(n2079), .A3(
        \SB1_1_2/Component_Function_5/NAND4_in[3] ), .A4(
        \SB1_1_2/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_2/buf_output[5] ) );
  NAND3_X1 U11706 ( .A1(\SB1_0_18/i0_3 ), .A2(\SB1_0_18/i1[9] ), .A3(n4753), 
        .ZN(\SB1_0_18/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U11707 ( .A1(\SB2_2_8/i0_4 ), .A2(\SB2_2_8/i0[8] ), .A3(
        \SB2_2_8/i1_7 ), .ZN(\SB2_2_8/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 U11708 ( .A1(\SB2_1_18/i0[9] ), .A2(\SB1_1_22/buf_output[1] ), .A3(
        \SB2_1_18/i0_4 ), .ZN(n5845) );
  NAND3_X1 U11709 ( .A1(\SB1_0_3/i0_0 ), .A2(\SB1_0_3/i0[9] ), .A3(
        \SB1_0_3/i0[8] ), .ZN(n5846) );
  NAND3_X2 U11710 ( .A1(\SB2_1_15/i0[10] ), .A2(\SB2_1_15/i0_3 ), .A3(
        \SB2_1_15/i0[6] ), .ZN(n5848) );
  XOR2_X1 U11711 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[105] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[81] ), .Z(\MC_ARK_ARC_1_0/temp2[135] )
         );
  XOR2_X1 U11712 ( .A1(n5850), .A2(n56), .Z(Ciphertext[152]) );
  XOR2_X1 U11713 ( .A1(\RI5[1][43] ), .A2(\RI5[1][79] ), .Z(
        \MC_ARK_ARC_1_1/temp3[169] ) );
  NAND3_X1 U11714 ( .A1(\SB3_9/i0_0 ), .A2(\SB3_9/i0_4 ), .A3(\SB3_9/i1_5 ), 
        .ZN(n5851) );
  NAND4_X2 U11715 ( .A1(n5864), .A2(\SB2_1_8/Component_Function_3/NAND4_in[0] ), .A3(\SB2_1_8/Component_Function_3/NAND4_in[3] ), .A4(n5852), .ZN(
        \SB2_1_8/buf_output[3] ) );
  NAND3_X2 U11716 ( .A1(\SB2_1_8/i0_4 ), .A2(\SB2_1_8/i0_0 ), .A3(
        \SB2_1_8/i0_3 ), .ZN(n5852) );
  XOR2_X1 U11717 ( .A1(\MC_ARK_ARC_1_0/temp2[185] ), .A2(n5853), .Z(n1345) );
  XOR2_X1 U11718 ( .A1(\RI5[0][185] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[179] ), .Z(n5853) );
  NAND4_X2 U11719 ( .A1(n4130), .A2(\SB2_0_0/Component_Function_3/NAND4_in[3] ), .A3(n4078), .A4(n5854), .ZN(\SB2_0_0/buf_output[3] ) );
  XOR2_X1 U11720 ( .A1(\RI5[1][121] ), .A2(\RI5[1][85] ), .Z(
        \MC_ARK_ARC_1_1/temp3[19] ) );
  NAND3_X2 U11721 ( .A1(\SB2_3_6/i0[9] ), .A2(\SB2_3_6/i0_4 ), .A3(
        \SB2_3_6/i0[6] ), .ZN(n5855) );
  INV_X1 U11722 ( .I(\SB3_9/buf_output[5] ), .ZN(\SB4_9/i1_5 ) );
  NAND4_X2 U11723 ( .A1(n4366), .A2(\SB3_9/Component_Function_5/NAND4_in[2] ), 
        .A3(n6149), .A4(\SB3_9/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB3_9/buf_output[5] ) );
  NAND4_X2 U11724 ( .A1(\SB3_11/Component_Function_2/NAND4_in[1] ), .A2(
        \SB3_11/Component_Function_2/NAND4_in[2] ), .A3(n3057), .A4(n6111), 
        .ZN(\SB3_11/buf_output[2] ) );
  XOR2_X1 U11725 ( .A1(\MC_ARK_ARC_1_1/temp5[18] ), .A2(n5856), .Z(
        \MC_ARK_ARC_1_1/buf_output[18] ) );
  XOR2_X1 U11726 ( .A1(\MC_ARK_ARC_1_1/temp3[18] ), .A2(
        \MC_ARK_ARC_1_1/temp4[18] ), .Z(n5856) );
  NAND3_X1 U11727 ( .A1(\SB2_0_5/i0_3 ), .A2(\SB2_0_5/i0[7] ), .A3(
        \SB2_0_5/i0_0 ), .ZN(\SB2_0_5/Component_Function_0/NAND4_in[3] ) );
  NOR2_X2 U11728 ( .A1(n5858), .A2(n5857), .ZN(\SB2_0_5/i0[7] ) );
  NAND2_X2 U11729 ( .A1(n6225), .A2(n1310), .ZN(n5858) );
  XOR2_X1 U11730 ( .A1(n5859), .A2(\MC_ARK_ARC_1_3/temp5[124] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[124] ) );
  XOR2_X1 U11731 ( .A1(\MC_ARK_ARC_1_3/temp4[124] ), .A2(
        \MC_ARK_ARC_1_3/temp3[124] ), .Z(n5859) );
  XOR2_X1 U11732 ( .A1(n5860), .A2(n65), .Z(Ciphertext[153]) );
  NAND4_X2 U11733 ( .A1(\SB4_6/Component_Function_3/NAND4_in[2] ), .A2(n821), 
        .A3(\SB4_6/Component_Function_3/NAND4_in[3] ), .A4(
        \SB4_6/Component_Function_3/NAND4_in[1] ), .ZN(n5860) );
  XOR2_X1 U11734 ( .A1(n5861), .A2(\MC_ARK_ARC_1_3/temp6[135] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[135] ) );
  XOR2_X1 U11735 ( .A1(\MC_ARK_ARC_1_3/temp1[135] ), .A2(
        \MC_ARK_ARC_1_3/temp2[135] ), .Z(n5861) );
  NAND4_X2 U11736 ( .A1(\SB2_1_27/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_1_27/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_1_27/Component_Function_0/NAND4_in[1] ), .A4(
        \SB2_1_27/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_1_27/buf_output[0] ) );
  NAND4_X2 U11737 ( .A1(n5989), .A2(
        \SB1_1_13/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_1_13/Component_Function_5/NAND4_in[3] ), .A4(n5862), .ZN(
        \SB1_1_13/buf_output[5] ) );
  NAND2_X2 U11738 ( .A1(\SB1_1_13/i0_0 ), .A2(\SB1_1_13/i3[0] ), .ZN(n5862) );
  XOR2_X1 U11739 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[159] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[153] ), .Z(\MC_ARK_ARC_1_1/temp1[159] )
         );
  NAND4_X2 U11740 ( .A1(n874), .A2(\SB2_2_28/Component_Function_3/NAND4_in[0] ), .A3(\SB2_2_28/Component_Function_3/NAND4_in[1] ), .A4(n5863), .ZN(
        \SB2_2_28/buf_output[3] ) );
  NAND3_X2 U11741 ( .A1(\SB2_0_29/i0_4 ), .A2(\SB2_0_29/i0_3 ), .A3(
        \SB2_0_29/i1[9] ), .ZN(n4610) );
  NAND3_X1 U11742 ( .A1(\SB2_1_30/i0[8] ), .A2(\SB2_1_30/i3[0] ), .A3(
        \SB2_1_30/i1_5 ), .ZN(\SB2_1_30/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U11743 ( .A1(\RI5[1][128] ), .A2(\RI5[1][92] ), .Z(n1686) );
  NAND2_X1 U11744 ( .A1(\SB3_7/i0_0 ), .A2(\SB3_7/i3[0] ), .ZN(n1680) );
  XOR2_X1 U11745 ( .A1(\RI5[2][188] ), .A2(\RI5[2][164] ), .Z(
        \MC_ARK_ARC_1_2/temp2[26] ) );
  XOR2_X1 U11746 ( .A1(n2752), .A2(\MC_ARK_ARC_1_0/temp5[135] ), .Z(n1377) );
  XOR2_X1 U11747 ( .A1(\MC_ARK_ARC_1_0/temp1[135] ), .A2(
        \MC_ARK_ARC_1_0/temp2[135] ), .Z(\MC_ARK_ARC_1_0/temp5[135] ) );
  NAND3_X2 U11748 ( .A1(\SB4_18/i0[6] ), .A2(\SB4_18/i1[9] ), .A3(
        \SB4_18/i0_3 ), .ZN(n3480) );
  NAND4_X2 U11749 ( .A1(n5945), .A2(\SB2_0_1/Component_Function_2/NAND4_in[0] ), .A3(n6338), .A4(n5865), .ZN(\SB2_0_1/buf_output[2] ) );
  NAND3_X2 U11750 ( .A1(\SB2_0_1/i0_0 ), .A2(\SB2_0_1/i1_5 ), .A3(
        \SB2_0_1/i0_4 ), .ZN(n5865) );
  XOR2_X1 U11751 ( .A1(\MC_ARK_ARC_1_2/temp5[39] ), .A2(n5866), .Z(
        \MC_ARK_ARC_1_2/buf_output[39] ) );
  XOR2_X1 U11752 ( .A1(\MC_ARK_ARC_1_2/temp4[39] ), .A2(
        \MC_ARK_ARC_1_2/temp3[39] ), .Z(n5866) );
  NAND4_X2 U11753 ( .A1(\SB1_1_27/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_1_27/Component_Function_2/NAND4_in[0] ), .A3(n3128), .A4(n5867), 
        .ZN(\SB1_1_27/buf_output[2] ) );
  XOR2_X1 U11754 ( .A1(\MC_ARK_ARC_1_0/temp4[125] ), .A2(n5868), .Z(
        \MC_ARK_ARC_1_0/temp6[125] ) );
  XOR2_X1 U11755 ( .A1(\RI5[0][35] ), .A2(\RI5[0][191] ), .Z(n5868) );
  XOR2_X1 U11756 ( .A1(n5870), .A2(n5869), .Z(\MC_ARK_ARC_1_0/buf_output[92] )
         );
  XOR2_X1 U11757 ( .A1(\MC_ARK_ARC_1_0/temp2[92] ), .A2(n2266), .Z(n5869) );
  XOR2_X1 U11758 ( .A1(n3925), .A2(n3924), .Z(n5870) );
  XOR2_X1 U11759 ( .A1(\MC_ARK_ARC_1_1/temp6[69] ), .A2(
        \MC_ARK_ARC_1_1/temp5[69] ), .Z(\MC_ARK_ARC_1_1/buf_output[69] ) );
  XOR2_X1 U11760 ( .A1(\RI5[1][40] ), .A2(\RI5[1][16] ), .Z(
        \MC_ARK_ARC_1_1/temp2[70] ) );
  XOR2_X1 U11761 ( .A1(\MC_ARK_ARC_1_2/temp3[59] ), .A2(
        \MC_ARK_ARC_1_2/temp4[59] ), .Z(n6008) );
  NAND3_X1 U11762 ( .A1(\SB3_20/i0[10] ), .A2(\SB3_20/i1_7 ), .A3(
        \SB3_20/i1[9] ), .ZN(n2577) );
  NAND4_X2 U11763 ( .A1(\SB2_3_30/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_3_30/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_3_30/Component_Function_2/NAND4_in[3] ), .A4(
        \SB2_3_30/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB2_3_30/buf_output[2] ) );
  XOR2_X1 U11764 ( .A1(\RI5[1][167] ), .A2(\RI5[1][143] ), .Z(
        \MC_ARK_ARC_1_1/temp2[5] ) );
  XOR2_X1 U11765 ( .A1(\RI5[3][50] ), .A2(\RI5[3][26] ), .Z(n5873) );
  NAND4_X2 U11766 ( .A1(\SB2_0_3/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_0_3/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_0_3/Component_Function_3/NAND4_in[3] ), .A4(
        \SB2_0_3/Component_Function_3/NAND4_in[1] ), .ZN(
        \SB2_0_3/buf_output[3] ) );
  NAND3_X1 U11767 ( .A1(\SB3_17/i0_3 ), .A2(\SB3_17/i0[8] ), .A3(\SB3_17/i1_7 ), .ZN(\SB3_17/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U11768 ( .A1(\SB2_0_2/i0_3 ), .A2(\RI3[0][176] ), .A3(\RI3[0][178] ), .ZN(n5876) );
  NAND4_X2 U11769 ( .A1(\SB3_16/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_16/Component_Function_3/NAND4_in[1] ), .A3(n2131), .A4(n5877), 
        .ZN(\RI3[4][105] ) );
  NAND3_X2 U11770 ( .A1(\SB3_16/i0[10] ), .A2(\SB3_16/i1[9] ), .A3(
        \SB3_16/i1_7 ), .ZN(n5877) );
  NAND3_X2 U11771 ( .A1(\SB2_3_9/i0_3 ), .A2(\SB2_3_9/i0[10] ), .A3(
        \SB2_3_9/i0[6] ), .ZN(n5878) );
  XOR2_X1 U11772 ( .A1(n5879), .A2(\MC_ARK_ARC_1_2/temp5[132] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[132] ) );
  XOR2_X1 U11773 ( .A1(\MC_ARK_ARC_1_2/temp4[132] ), .A2(
        \MC_ARK_ARC_1_2/temp3[132] ), .Z(n5879) );
  NAND3_X1 U11774 ( .A1(\SB1_3_18/i0_4 ), .A2(\SB1_3_18/i1[9] ), .A3(
        \SB1_3_18/i1_5 ), .ZN(\SB1_3_18/Component_Function_4/NAND4_in[3] ) );
  NAND3_X2 U11775 ( .A1(\SB2_2_8/i0[6] ), .A2(\SB2_2_8/i0_4 ), .A3(n5880), 
        .ZN(\SB2_2_8/Component_Function_5/NAND4_in[3] ) );
  NAND4_X2 U11776 ( .A1(n1958), .A2(\SB2_0_2/Component_Function_2/NAND4_in[0] ), .A3(\SB2_0_2/Component_Function_2/NAND4_in[1] ), .A4(
        \SB2_0_2/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_0_2/buf_output[2] ) );
  NAND3_X2 U11777 ( .A1(\SB2_0_2/i0[6] ), .A2(\SB2_0_2/i0[9] ), .A3(
        \SB2_0_2/i1_5 ), .ZN(\SB2_0_2/Component_Function_1/NAND4_in[2] ) );
  XOR2_X1 U11778 ( .A1(n5885), .A2(n5884), .Z(n4298) );
  XOR2_X1 U11779 ( .A1(\RI5[2][173] ), .A2(\RI5[2][5] ), .Z(n5884) );
  XOR2_X1 U11780 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[29] ), .A2(\RI5[2][35] ), 
        .Z(n5885) );
  BUF_X2 U11781 ( .I(n2342), .Z(n5886) );
  INV_X2 U11782 ( .I(\SB1_2_20/buf_output[3] ), .ZN(\SB2_2_18/i0[8] ) );
  NAND4_X2 U11783 ( .A1(\SB2_1_15/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_1_15/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_15/Component_Function_3/NAND4_in[3] ), .A4(n5887), .ZN(
        \SB2_1_15/buf_output[3] ) );
  NAND3_X2 U11784 ( .A1(\SB2_1_15/i0_3 ), .A2(\SB2_1_15/i0[6] ), .A3(
        \SB2_1_15/i1[9] ), .ZN(n5887) );
  XOR2_X1 U11785 ( .A1(\RI5[0][148] ), .A2(\RI5[0][184] ), .Z(
        \MC_ARK_ARC_1_0/temp3[82] ) );
  XOR2_X1 U11786 ( .A1(n5889), .A2(n5888), .Z(n3069) );
  XOR2_X1 U11787 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[116] ), .A2(n511), .Z(
        n5888) );
  NAND3_X2 U11788 ( .A1(\SB2_1_28/i1_7 ), .A2(\SB2_1_28/i0[10] ), .A3(
        \SB2_1_28/i1[9] ), .ZN(\SB2_1_28/Component_Function_3/NAND4_in[2] ) );
  AND4_X2 U11789 ( .A1(\SB1_3_28/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_3_28/Component_Function_3/NAND4_in[0] ), .A3(
        \SB1_3_28/Component_Function_3/NAND4_in[3] ), .A4(n2316), .Z(n5890) );
  XOR2_X1 U11790 ( .A1(\RI5[1][10] ), .A2(\RI5[1][106] ), .Z(n5891) );
  XOR2_X1 U11791 ( .A1(n2433), .A2(n5892), .Z(\MC_ARK_ARC_1_1/buf_output[35] )
         );
  XOR2_X1 U11792 ( .A1(n624), .A2(\MC_ARK_ARC_1_1/temp1[35] ), .Z(n5892) );
  XOR2_X1 U11793 ( .A1(n5894), .A2(n5893), .Z(n2476) );
  XOR2_X1 U11794 ( .A1(\RI5[1][158] ), .A2(\RI5[1][20] ), .Z(n5893) );
  XOR2_X1 U11795 ( .A1(\RI5[1][182] ), .A2(\RI5[1][14] ), .Z(n5894) );
  XOR2_X1 U11796 ( .A1(\RI5[1][182] ), .A2(\RI5[1][146] ), .Z(
        \MC_ARK_ARC_1_1/temp3[80] ) );
  NAND4_X2 U11797 ( .A1(n1265), .A2(\SB1_0_0/Component_Function_5/NAND4_in[2] ), .A3(\SB1_0_0/Component_Function_5/NAND4_in[0] ), .A4(n6482), .ZN(
        \SB1_0_0/buf_output[5] ) );
  INV_X2 U11798 ( .I(\SB1_1_28/buf_output[2] ), .ZN(\SB2_1_25/i1[9] ) );
  NAND4_X2 U11799 ( .A1(n3264), .A2(
        \SB1_1_28/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_1_28/Component_Function_2/NAND4_in[2] ), .A4(n1130), .ZN(
        \SB1_1_28/buf_output[2] ) );
  INV_X1 U11800 ( .I(\SB3_9/buf_output[3] ), .ZN(\SB4_7/i0[8] ) );
  NAND4_X2 U11801 ( .A1(\SB3_9/Component_Function_3/NAND4_in[2] ), .A2(
        \SB3_9/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_9/Component_Function_3/NAND4_in[0] ), .A4(n2480), .ZN(
        \SB3_9/buf_output[3] ) );
  XOR2_X1 U11802 ( .A1(\MC_ARK_ARC_1_1/temp3[15] ), .A2(n1645), .Z(n1839) );
  XOR2_X1 U11803 ( .A1(\MC_ARK_ARC_1_0/temp2[104] ), .A2(n5896), .Z(n949) );
  XOR2_X1 U11804 ( .A1(\RI5[0][104] ), .A2(\RI5[0][98] ), .Z(n5896) );
  NAND4_X2 U11805 ( .A1(n1661), .A2(\SB2_2_5/Component_Function_3/NAND4_in[3] ), .A3(\SB2_2_5/Component_Function_3/NAND4_in[2] ), .A4(n3793), .ZN(
        \SB2_2_5/buf_output[3] ) );
  XOR2_X1 U11806 ( .A1(n5898), .A2(n5897), .Z(\MC_ARK_ARC_1_3/temp6[166] ) );
  XOR2_X1 U11807 ( .A1(\RI5[3][76] ), .A2(n113), .Z(n5897) );
  XOR2_X1 U11808 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[40] ), .A2(\RI5[3][10] ), 
        .Z(n5898) );
  XOR2_X1 U11809 ( .A1(n5899), .A2(\MC_ARK_ARC_1_0/temp4[113] ), .Z(n6240) );
  XOR2_X1 U11810 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[179] ), .A2(\RI5[0][23] ), 
        .Z(n5899) );
  XOR2_X1 U11811 ( .A1(n5901), .A2(n5900), .Z(n6244) );
  XOR2_X1 U11812 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[182] ), .A2(n110), .Z(
        n5900) );
  XOR2_X1 U11813 ( .A1(\RI5[3][32] ), .A2(\RI5[3][188] ), .Z(n5901) );
  NAND4_X2 U11814 ( .A1(\SB1_3_22/Component_Function_2/NAND4_in[0] ), .A2(
        n1245), .A3(\SB1_3_22/Component_Function_2/NAND4_in[2] ), .A4(n5902), 
        .ZN(\SB1_3_22/buf_output[2] ) );
  NAND3_X2 U11815 ( .A1(\SB1_3_22/i0[10] ), .A2(\SB1_3_22/i0[6] ), .A3(
        \SB1_3_22/i0_3 ), .ZN(n5902) );
  NAND4_X2 U11816 ( .A1(\SB2_2_17/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_17/Component_Function_3/NAND4_in[3] ), .A3(
        \SB2_2_17/Component_Function_3/NAND4_in[1] ), .A4(n5903), .ZN(
        \SB2_2_17/buf_output[3] ) );
  NAND3_X2 U11817 ( .A1(\SB2_2_17/i0[10] ), .A2(\SB2_2_17/i1_7 ), .A3(
        \SB2_2_17/i1[9] ), .ZN(n5903) );
  XOR2_X1 U11818 ( .A1(\RI5[3][59] ), .A2(\RI5[3][35] ), .Z(n5905) );
  NAND4_X2 U11819 ( .A1(\SB3_14/Component_Function_1/NAND4_in[2] ), .A2(
        \SB3_14/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_14/Component_Function_1/NAND4_in[0] ), .A4(n5907), .ZN(
        \SB3_14/buf_output[1] ) );
  NAND3_X1 U11820 ( .A1(\SB3_14/i1_7 ), .A2(\SB3_14/i0_4 ), .A3(\SB3_14/i0[8] ), .ZN(n5907) );
  XOR2_X1 U11821 ( .A1(n5909), .A2(n5908), .Z(\MC_ARK_ARC_1_2/temp5[2] ) );
  XOR2_X1 U11822 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[2] ), .A2(\RI5[2][164] ), 
        .Z(n5908) );
  XOR2_X1 U11823 ( .A1(\RI5[2][188] ), .A2(\RI5[2][140] ), .Z(n5909) );
  NAND4_X2 U11824 ( .A1(\SB2_2_19/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_19/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_2_19/Component_Function_2/NAND4_in[2] ), .A4(n5910), .ZN(
        \SB2_2_19/buf_output[2] ) );
  XOR2_X1 U11825 ( .A1(\SB2_1_6/buf_output[2] ), .A2(\RI5[1][116] ), .Z(n5912)
         );
  XOR2_X1 U11826 ( .A1(n5913), .A2(n4256), .Z(n3786) );
  XOR2_X1 U11827 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[2] ), .A2(\RI5[2][170] ), 
        .Z(n5913) );
  XOR2_X1 U11828 ( .A1(\MC_ARK_ARC_1_0/temp5[179] ), .A2(n5914), .Z(
        \MC_ARK_ARC_1_0/buf_output[179] ) );
  XOR2_X1 U11829 ( .A1(\MC_ARK_ARC_1_0/temp3[179] ), .A2(
        \MC_ARK_ARC_1_0/temp4[179] ), .Z(n5914) );
  XOR2_X1 U11830 ( .A1(\MC_ARK_ARC_1_3/temp2[56] ), .A2(n5915), .Z(
        \MC_ARK_ARC_1_3/temp5[56] ) );
  XOR2_X1 U11831 ( .A1(\RI5[3][50] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[56] ), 
        .Z(n5915) );
  XOR2_X1 U11832 ( .A1(n5916), .A2(n2), .Z(Ciphertext[48]) );
  NAND4_X2 U11833 ( .A1(n4690), .A2(
        \SB2_1_22/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_1_22/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_1_22/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB2_1_22/buf_output[4] ) );
  XOR2_X1 U11834 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[153] ), .A2(n5521), .Z(
        \MC_ARK_ARC_1_1/temp1[153] ) );
  INV_X2 U11835 ( .I(\SB1_0_0/buf_output[1] ), .ZN(\SB2_0_28/i1_7 ) );
  NAND4_X2 U11836 ( .A1(\SB1_1_1/Component_Function_5/NAND4_in[1] ), .A2(n6232), .A3(n4744), .A4(\SB1_1_1/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_1/buf_output[5] ) );
  NAND3_X1 U11837 ( .A1(\SB3_17/i0[10] ), .A2(\SB3_17/i1[9] ), .A3(
        \SB3_17/i1_7 ), .ZN(n3963) );
  NAND3_X2 U11838 ( .A1(\SB2_0_7/i0_3 ), .A2(\SB2_0_7/i1_7 ), .A3(
        \SB2_0_7/i0[8] ), .ZN(\SB2_0_7/Component_Function_1/NAND4_in[1] ) );
  NAND3_X2 U11839 ( .A1(\SB1_3_13/i0[6] ), .A2(\SB1_3_13/i0[10] ), .A3(
        \SB1_3_13/i0_0 ), .ZN(n6494) );
  NAND4_X2 U11840 ( .A1(\SB2_3_3/Component_Function_5/NAND4_in[2] ), .A2(n1477), .A3(n6016), .A4(n6020), .ZN(\SB2_3_3/buf_output[5] ) );
  XOR2_X1 U11841 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[191] ), .A2(\RI5[3][23] ), 
        .Z(\MC_ARK_ARC_1_3/temp2[53] ) );
  NAND3_X2 U11842 ( .A1(\SB2_3_7/i0[10] ), .A2(\SB2_3_7/i1_5 ), .A3(
        \SB2_3_7/i1[9] ), .ZN(\SB2_3_7/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U11843 ( .A1(n5917), .A2(n6327), .Z(\MC_ARK_ARC_1_1/buf_output[113] ) );
  XOR2_X1 U11844 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[95] ), .A2(\RI5[1][161] ), 
        .Z(n3956) );
  XOR2_X1 U11845 ( .A1(\MC_ARK_ARC_1_2/temp4[43] ), .A2(
        \MC_ARK_ARC_1_2/temp3[43] ), .Z(n593) );
  NAND4_X2 U11846 ( .A1(\SB1_1_20/Component_Function_1/NAND4_in[3] ), .A2(
        n6233), .A3(\SB1_1_20/Component_Function_1/NAND4_in[1] ), .A4(
        \SB1_1_20/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_1_20/buf_output[1] ) );
  XOR2_X1 U11847 ( .A1(\MC_ARK_ARC_1_2/temp2[133] ), .A2(
        \MC_ARK_ARC_1_2/temp1[133] ), .Z(n6128) );
  NAND4_X2 U11848 ( .A1(\SB2_3_14/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_3_14/Component_Function_2/NAND4_in[2] ), .A3(n4341), .A4(
        \SB2_3_14/Component_Function_2/NAND4_in[1] ), .ZN(
        \SB2_3_14/buf_output[2] ) );
  NAND4_X2 U11849 ( .A1(\SB1_2_22/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_2_22/Component_Function_5/NAND4_in[1] ), .A3(n5982), .A4(
        \SB1_2_22/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_2_22/buf_output[5] ) );
  NAND4_X2 U11850 ( .A1(\SB1_0_2/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_0_2/Component_Function_5/NAND4_in[1] ), .A3(n1715), .A4(n5919), 
        .ZN(\RI3[0][179] ) );
  NAND3_X1 U11851 ( .A1(\SB1_0_2/i0[6] ), .A2(\SB1_0_2/i0[9] ), .A3(n400), 
        .ZN(n5919) );
  NAND3_X2 U11852 ( .A1(\SB1_3_15/i0[10] ), .A2(\SB1_3_15/i1[9] ), .A3(
        \SB1_3_15/i1_7 ), .ZN(n5920) );
  NAND3_X1 U11853 ( .A1(\SB1_2_14/i1_5 ), .A2(\SB1_2_14/i1[9] ), .A3(
        \SB1_2_14/i0_4 ), .ZN(n5921) );
  NAND4_X2 U11854 ( .A1(\SB2_2_13/Component_Function_1/NAND4_in[2] ), .A2(
        \SB2_2_13/Component_Function_1/NAND4_in[1] ), .A3(
        \SB2_2_13/Component_Function_1/NAND4_in[0] ), .A4(n5922), .ZN(
        \SB2_2_13/buf_output[1] ) );
  NAND3_X2 U11855 ( .A1(n580), .A2(\SB2_2_13/i0[8] ), .A3(\SB2_2_13/i1_7 ), 
        .ZN(n5922) );
  XOR2_X1 U11856 ( .A1(\MC_ARK_ARC_1_1/temp4[135] ), .A2(n5923), .Z(n2117) );
  XOR2_X1 U11857 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[9] ), .A2(\RI5[1][45] ), 
        .Z(n5923) );
  XOR2_X1 U11858 ( .A1(n5924), .A2(n3834), .Z(\MC_ARK_ARC_1_0/buf_output[59] )
         );
  XOR2_X1 U11859 ( .A1(\MC_ARK_ARC_1_0/temp3[59] ), .A2(n1869), .Z(n5924) );
  XOR2_X1 U11860 ( .A1(\MC_ARK_ARC_1_1/temp2[136] ), .A2(
        \MC_ARK_ARC_1_1/temp4[136] ), .Z(n1347) );
  NAND3_X1 U11861 ( .A1(\SB2_3_20/i0[10] ), .A2(\SB2_3_20/i0_3 ), .A3(
        \SB2_3_20/i0_4 ), .ZN(\SB2_3_20/Component_Function_0/NAND4_in[2] ) );
  NAND2_X2 U11862 ( .A1(n2634), .A2(n1209), .ZN(\SB2_3_20/i0_4 ) );
  NAND4_X2 U11863 ( .A1(\SB2_1_19/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_19/Component_Function_4/NAND4_in[1] ), .A3(n2472), .A4(n5925), 
        .ZN(\SB2_1_19/buf_output[4] ) );
  NAND3_X1 U11864 ( .A1(n578), .A2(n1396), .A3(\SB2_1_19/i1_5 ), .ZN(n5925) );
  NAND3_X1 U11865 ( .A1(\SB2_1_30/i0[6] ), .A2(\SB2_1_30/i0[9] ), .A3(
        \SB2_1_30/i1_5 ), .ZN(\SB2_1_30/Component_Function_1/NAND4_in[2] ) );
  XOR2_X1 U11866 ( .A1(\MC_ARK_ARC_1_1/temp5[37] ), .A2(
        \MC_ARK_ARC_1_1/temp6[37] ), .Z(\MC_ARK_ARC_1_1/buf_output[37] ) );
  XOR2_X1 U11867 ( .A1(\RI5[3][159] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[135] ), .Z(n2780) );
  XOR2_X1 U11868 ( .A1(n5928), .A2(n5927), .Z(n6029) );
  XOR2_X1 U11869 ( .A1(\RI5[0][47] ), .A2(\RI5[0][119] ), .Z(n5927) );
  XOR2_X1 U11870 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[155] ), .A2(\RI5[0][53] ), 
        .Z(n5928) );
  XOR2_X1 U11871 ( .A1(n6477), .A2(n5929), .Z(\MC_ARK_ARC_1_1/temp6[116] ) );
  XOR2_X1 U11872 ( .A1(\RI5[1][26] ), .A2(\RI5[1][152] ), .Z(n5929) );
  INV_X2 U11873 ( .I(\SB1_3_6/buf_output[2] ), .ZN(\SB2_3_3/i1[9] ) );
  NAND4_X2 U11874 ( .A1(\SB1_3_6/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_6/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_3_6/Component_Function_2/NAND4_in[2] ), .A4(n1210), .ZN(
        \SB1_3_6/buf_output[2] ) );
  NAND3_X2 U11875 ( .A1(\SB2_0_22/i0_0 ), .A2(\SB2_0_22/i0[6] ), .A3(
        \SB2_0_22/i0[10] ), .ZN(n5930) );
  NAND2_X2 U11876 ( .A1(\SB1_0_9/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_9/Component_Function_3/NAND4_in[1] ), .ZN(n5931) );
  XOR2_X1 U11877 ( .A1(n1392), .A2(\RI5[3][147] ), .Z(
        \MC_ARK_ARC_1_3/temp3[45] ) );
  NAND3_X1 U11878 ( .A1(\SB2_2_15/i0_4 ), .A2(\SB2_2_15/i0[9] ), .A3(
        \SB1_2_19/buf_output[1] ), .ZN(
        \SB2_2_15/Component_Function_5/NAND4_in[3] ) );
  NAND4_X2 U11879 ( .A1(\SB2_0_24/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_0_24/Component_Function_0/NAND4_in[0] ), .A3(
        \SB2_0_24/Component_Function_0/NAND4_in[2] ), .A4(n5933), .ZN(
        \SB2_0_24/buf_output[0] ) );
  NAND3_X2 U11880 ( .A1(\SB1_1_20/i0[6] ), .A2(\SB1_1_20/i0[9] ), .A3(
        \SB1_1_20/i0_4 ), .ZN(n1944) );
  NAND4_X2 U11881 ( .A1(\SB2_1_2/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_2/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_1_2/Component_Function_2/NAND4_in[1] ), .A4(n1689), .ZN(
        \SB2_1_2/buf_output[2] ) );
  NAND4_X2 U11882 ( .A1(\SB2_2_15/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_2_15/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_2_15/Component_Function_0/NAND4_in[0] ), .A4(n5934), .ZN(
        \SB2_2_15/buf_output[0] ) );
  NAND3_X2 U11883 ( .A1(\SB2_2_15/i0_3 ), .A2(\SB2_2_15/i0_0 ), .A3(n722), 
        .ZN(n5934) );
  XOR2_X1 U11884 ( .A1(\MC_ARK_ARC_1_1/temp1[83] ), .A2(n5935), .Z(
        \MC_ARK_ARC_1_1/temp5[83] ) );
  XOR2_X1 U11885 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[29] ), .A2(\RI5[1][53] ), 
        .Z(n5935) );
  XOR2_X1 U11886 ( .A1(n5936), .A2(n100), .Z(Ciphertext[91]) );
  NAND4_X2 U11887 ( .A1(\SB4_16/Component_Function_1/NAND4_in[3] ), .A2(
        \SB4_16/Component_Function_1/NAND4_in[1] ), .A3(
        \SB4_16/Component_Function_1/NAND4_in[2] ), .A4(
        \SB4_16/Component_Function_1/NAND4_in[0] ), .ZN(n5936) );
  INV_X2 U11888 ( .I(\SB3_18/buf_output[3] ), .ZN(\SB4_16/i0[8] ) );
  XOR2_X1 U11889 ( .A1(\RI5[3][73] ), .A2(\RI5[3][79] ), .Z(
        \MC_ARK_ARC_1_3/temp1[79] ) );
  XOR2_X1 U11890 ( .A1(\RI5[0][53] ), .A2(\RI5[0][89] ), .Z(
        \MC_ARK_ARC_1_0/temp3[179] ) );
  XOR2_X1 U11891 ( .A1(n5940), .A2(\MC_ARK_ARC_1_3/temp4[83] ), .Z(n757) );
  XOR2_X1 U11892 ( .A1(\RI5[3][185] ), .A2(\RI5[3][149] ), .Z(n5940) );
  NAND3_X2 U11893 ( .A1(\SB2_3_27/i0[10] ), .A2(\SB2_3_27/i1_7 ), .A3(
        \SB2_3_27/i1[9] ), .ZN(\SB2_3_27/Component_Function_3/NAND4_in[2] ) );
  NAND4_X2 U11894 ( .A1(\SB1_2_15/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_15/Component_Function_3/NAND4_in[1] ), .A3(n4085), .A4(n5941), 
        .ZN(\SB1_2_15/buf_output[3] ) );
  NAND3_X2 U11895 ( .A1(\SB1_1_2/i0_3 ), .A2(\SB1_1_2/i0[6] ), .A3(
        \SB1_1_2/i1[9] ), .ZN(n6010) );
  XOR2_X1 U11896 ( .A1(\RI5[0][13] ), .A2(\RI5[0][169] ), .Z(
        \MC_ARK_ARC_1_0/temp3[103] ) );
  NAND4_X2 U11897 ( .A1(n4544), .A2(n6494), .A3(
        \SB1_3_13/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_3_13/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_13/buf_output[5] ) );
  XOR2_X1 U11898 ( .A1(n5944), .A2(n5943), .Z(\MC_ARK_ARC_1_2/temp5[109] ) );
  XOR2_X1 U11899 ( .A1(\RI5[2][109] ), .A2(\RI5[2][55] ), .Z(n5943) );
  XOR2_X1 U11900 ( .A1(\RI5[2][103] ), .A2(\RI5[2][79] ), .Z(n5944) );
  NAND3_X2 U11901 ( .A1(\SB2_0_1/i0[9] ), .A2(\SB2_0_1/i0[8] ), .A3(
        \SB2_0_1/i0_3 ), .ZN(n5945) );
  NAND3_X2 U11902 ( .A1(\SB3_17/i0[6] ), .A2(\SB3_17/i0_4 ), .A3(
        \SB3_17/i0[9] ), .ZN(n5946) );
  NAND4_X2 U11903 ( .A1(\SB4_18/Component_Function_0/NAND4_in[1] ), .A2(
        \SB4_18/Component_Function_0/NAND4_in[3] ), .A3(
        \SB4_18/Component_Function_0/NAND4_in[0] ), .A4(n5947), .ZN(n6171) );
  NAND3_X2 U11904 ( .A1(\SB4_18/i0_4 ), .A2(\SB4_18/i0_3 ), .A3(
        \SB4_18/i0[10] ), .ZN(n5947) );
  NAND2_X2 U11905 ( .A1(\SB1_1_0/Component_Function_4/NAND4_in[1] ), .A2(n5948), .ZN(n5999) );
  NAND3_X2 U11906 ( .A1(\SB1_1_0/i0[10] ), .A2(\SB1_1_0/i0[9] ), .A3(
        \SB1_1_0/i0_3 ), .ZN(n5948) );
  NAND3_X1 U11907 ( .A1(\SB3_23/i1[9] ), .A2(\SB3_23/i0[10] ), .A3(
        \SB3_23/i1_5 ), .ZN(\SB3_23/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U11908 ( .A1(n5950), .A2(n5949), .Z(\MC_ARK_ARC_1_2/temp6[14] ) );
  XOR2_X1 U11909 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[116] ), .A2(n502), .Z(
        n5949) );
  XOR2_X1 U11910 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[50] ), .A2(\RI5[2][80] ), 
        .Z(n5950) );
  NAND3_X2 U11911 ( .A1(\SB1_3_17/i0_4 ), .A2(\SB1_3_17/i0[6] ), .A3(
        \SB1_3_17/i0[9] ), .ZN(\SB1_3_17/Component_Function_5/NAND4_in[3] ) );
  NAND2_X1 U11912 ( .A1(\RI1[3][14] ), .A2(\SB1_3_29/i3[0] ), .ZN(
        \SB1_3_29/Component_Function_5/NAND4_in[0] ) );
  NAND3_X1 U11913 ( .A1(\SB1_2_14/i0_3 ), .A2(\SB1_2_14/i0_0 ), .A3(
        \SB1_2_14/i0_4 ), .ZN(\SB1_2_14/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U11914 ( .A1(\SB2_3_15/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_3_15/Component_Function_1/NAND4_in[0] ), .A3(
        \SB2_3_15/Component_Function_1/NAND4_in[2] ), .A4(n5951), .ZN(
        \SB2_3_15/buf_output[1] ) );
  NAND3_X2 U11915 ( .A1(\SB2_3_15/i0_3 ), .A2(\SB2_3_15/i1_7 ), .A3(n3670), 
        .ZN(n5951) );
  XOR2_X1 U11916 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[99] ), .A2(\RI5[1][75] ), 
        .Z(n2945) );
  NAND3_X2 U11917 ( .A1(\SB1_2_15/i0_4 ), .A2(\SB1_2_15/i1_7 ), .A3(
        \SB1_2_15/i0[8] ), .ZN(\SB1_2_15/Component_Function_1/NAND4_in[3] ) );
  XOR2_X1 U11918 ( .A1(n3486), .A2(n5952), .Z(\MC_ARK_ARC_1_1/buf_output[100] ) );
  XOR2_X1 U11919 ( .A1(\MC_ARK_ARC_1_1/temp3[100] ), .A2(
        \MC_ARK_ARC_1_1/temp4[100] ), .Z(n5952) );
  NAND4_X2 U11920 ( .A1(\SB2_1_21/Component_Function_3/NAND4_in[2] ), .A2(
        n1208), .A3(n3227), .A4(n4748), .ZN(\SB2_1_21/buf_output[3] ) );
  NAND3_X1 U11921 ( .A1(\SB2_3_23/i0_4 ), .A2(\SB2_3_23/i0_3 ), .A3(
        \SB2_3_23/i0[10] ), .ZN(\SB2_3_23/Component_Function_0/NAND4_in[2] )
         );
  NAND3_X2 U11922 ( .A1(\SB2_1_31/i0_3 ), .A2(\SB2_1_31/i0[6] ), .A3(
        \SB2_1_31/i1[9] ), .ZN(\SB2_1_31/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U11923 ( .A1(n5953), .A2(n5954), .Z(\MC_ARK_ARC_1_3/temp5[78] ) );
  XOR2_X1 U11924 ( .A1(\RI5[3][24] ), .A2(\RI5[3][72] ), .Z(n5953) );
  XOR2_X1 U11925 ( .A1(\RI5[3][78] ), .A2(\RI5[3][48] ), .Z(n5954) );
  XOR2_X1 U11926 ( .A1(\RI5[0][117] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[141] ), .Z(\MC_ARK_ARC_1_0/temp2[171] ) );
  NAND3_X2 U11927 ( .A1(\SB2_2_19/i0[10] ), .A2(\SB2_2_19/i1_7 ), .A3(
        \SB2_2_19/i1[9] ), .ZN(n6383) );
  INV_X2 U11928 ( .I(\SB1_1_24/buf_output[2] ), .ZN(\SB2_1_21/i1[9] ) );
  NAND4_X2 U11929 ( .A1(\SB1_1_24/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_1_24/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_1_24/Component_Function_2/NAND4_in[0] ), .A4(
        \SB1_1_24/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB1_1_24/buf_output[2] ) );
  NAND4_X2 U11930 ( .A1(\SB1_2_6/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_6/Component_Function_3/NAND4_in[2] ), .A3(
        \SB1_2_6/Component_Function_3/NAND4_in[1] ), .A4(n4559), .ZN(
        \SB1_2_6/buf_output[3] ) );
  NAND4_X2 U11931 ( .A1(\SB1_1_24/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_1_24/Component_Function_3/NAND4_in[0] ), .A3(n2876), .A4(n5955), 
        .ZN(\SB1_1_24/buf_output[3] ) );
  NAND3_X1 U11932 ( .A1(\SB4_8/i1_7 ), .A2(\SB4_8/i0_3 ), .A3(\SB4_8/i0[8] ), 
        .ZN(\SB4_8/Component_Function_1/NAND4_in[1] ) );
  NAND3_X2 U11933 ( .A1(\SB1_1_10/i0[9] ), .A2(\SB1_1_10/i0_3 ), .A3(
        \SB1_1_10/i0[8] ), .ZN(n6018) );
  XOR2_X1 U11934 ( .A1(n3808), .A2(\MC_ARK_ARC_1_1/temp6[155] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[155] ) );
  XOR2_X1 U11935 ( .A1(\RI5[0][77] ), .A2(\RI5[0][101] ), .Z(
        \MC_ARK_ARC_1_0/temp2[131] ) );
  INV_X4 U11936 ( .I(n5956), .ZN(n3645) );
  NOR2_X2 U11937 ( .A1(n1508), .A2(n1370), .ZN(n5956) );
  XOR2_X1 U11938 ( .A1(\RI5[0][163] ), .A2(\RI5[0][187] ), .Z(
        \MC_ARK_ARC_1_0/temp2[25] ) );
  XOR2_X1 U11939 ( .A1(n4299), .A2(n4300), .Z(\MC_ARK_ARC_1_0/buf_output[131] ) );
  NAND4_X2 U11940 ( .A1(\SB1_2_24/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_2_24/Component_Function_3/NAND4_in[0] ), .A3(n4413), .A4(n5957), 
        .ZN(\SB1_2_24/buf_output[3] ) );
  XOR2_X1 U11941 ( .A1(n4435), .A2(\MC_ARK_ARC_1_2/temp5[4] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[4] ) );
  NAND4_X2 U11942 ( .A1(n885), .A2(n6343), .A3(
        \SB2_0_19/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_0_19/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_0_19/buf_output[5] ) );
  NAND4_X2 U11943 ( .A1(\SB2_1_3/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_3/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_1_3/Component_Function_4/NAND4_in[1] ), .A4(n5958), .ZN(
        \SB2_1_3/buf_output[4] ) );
  NAND4_X2 U11944 ( .A1(\SB2_1_0/Component_Function_5/NAND4_in[2] ), .A2(n968), 
        .A3(n3756), .A4(\SB2_1_0/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_1_0/buf_output[5] ) );
  XOR2_X1 U11945 ( .A1(n5961), .A2(n5960), .Z(\MC_ARK_ARC_1_2/buf_output[8] )
         );
  XOR2_X1 U11946 ( .A1(\MC_ARK_ARC_1_2/temp1[8] ), .A2(
        \MC_ARK_ARC_1_2/temp3[8] ), .Z(n5960) );
  XOR2_X1 U11947 ( .A1(\MC_ARK_ARC_1_2/temp2[8] ), .A2(
        \MC_ARK_ARC_1_2/temp4[8] ), .Z(n5961) );
  XOR2_X1 U11948 ( .A1(n5962), .A2(\MC_ARK_ARC_1_0/temp2[153] ), .Z(
        \MC_ARK_ARC_1_0/temp5[153] ) );
  XOR2_X1 U11949 ( .A1(\RI5[0][147] ), .A2(\RI5[0][153] ), .Z(n5962) );
  INV_X2 U11950 ( .I(\SB1_2_8/i0[7] ), .ZN(\SB1_2_8/i0_4 ) );
  XNOR2_X1 U11951 ( .A1(\MC_ARK_ARC_1_1/temp5[142] ), .A2(
        \MC_ARK_ARC_1_1/temp6[142] ), .ZN(\SB1_2_8/i0[7] ) );
  INV_X2 U11952 ( .I(\SB3_18/buf_output[5] ), .ZN(\SB4_18/i1_5 ) );
  NAND3_X2 U11953 ( .A1(\SB2_0_7/i0[10] ), .A2(n2593), .A3(\SB2_0_7/i0_0 ), 
        .ZN(\SB2_0_7/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U11954 ( .A1(n5964), .A2(n5963), .Z(\MC_ARK_ARC_1_0/buf_output[149] ) );
  XOR2_X1 U11955 ( .A1(\MC_ARK_ARC_1_0/temp3[149] ), .A2(n6354), .Z(n5963) );
  XOR2_X1 U11956 ( .A1(\MC_ARK_ARC_1_0/temp2[170] ), .A2(n5965), .Z(n744) );
  XOR2_X1 U11957 ( .A1(\RI5[0][170] ), .A2(\RI5[0][164] ), .Z(n5965) );
  NAND3_X2 U11958 ( .A1(\SB1_1_3/i0_4 ), .A2(\SB1_1_3/i1[9] ), .A3(
        \SB1_1_3/i1_5 ), .ZN(n1643) );
  XOR2_X1 U11959 ( .A1(n5967), .A2(n5966), .Z(\MC_ARK_ARC_1_2/temp6[50] ) );
  XOR2_X1 U11960 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[116] ), .A2(n461), .Z(
        n5966) );
  XOR2_X1 U11961 ( .A1(\RI5[2][152] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[86] ), 
        .Z(n5967) );
  NAND4_X2 U11962 ( .A1(\SB2_1_29/Component_Function_5/NAND4_in[3] ), .A2(
        \SB2_1_29/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_1_29/Component_Function_5/NAND4_in[0] ), .A4(n5968), .ZN(
        \SB2_1_29/buf_output[5] ) );
  XOR2_X1 U11963 ( .A1(\MC_ARK_ARC_1_1/temp5[71] ), .A2(n4150), .Z(
        \MC_ARK_ARC_1_1/buf_output[71] ) );
  XOR2_X1 U11964 ( .A1(\MC_ARK_ARC_1_1/temp1[71] ), .A2(
        \MC_ARK_ARC_1_1/temp2[71] ), .Z(\MC_ARK_ARC_1_1/temp5[71] ) );
  AND2_X1 U11965 ( .A1(\MC_ARK_ARC_1_2/buf_output[46] ), .A2(
        \MC_ARK_ARC_1_2/buf_output[42] ), .Z(n5970) );
  XOR2_X1 U11966 ( .A1(n5972), .A2(n5971), .Z(\MC_ARK_ARC_1_1/buf_output[88] )
         );
  XOR2_X1 U11967 ( .A1(\MC_ARK_ARC_1_1/temp3[88] ), .A2(
        \MC_ARK_ARC_1_1/temp4[88] ), .Z(n5971) );
  XOR2_X1 U11968 ( .A1(\MC_ARK_ARC_1_1/temp2[88] ), .A2(
        \MC_ARK_ARC_1_1/temp1[88] ), .Z(n5972) );
  XOR2_X1 U11969 ( .A1(n5975), .A2(n5974), .Z(\MC_ARK_ARC_1_2/temp6[38] ) );
  XOR2_X1 U11970 ( .A1(\RI5[2][140] ), .A2(n519), .Z(n5974) );
  XOR2_X1 U11971 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[74] ), .A2(\RI5[2][104] ), 
        .Z(n5975) );
  NAND3_X2 U11972 ( .A1(\SB2_0_22/i0_4 ), .A2(\SB2_0_22/i0_0 ), .A3(
        \SB2_0_22/i1_5 ), .ZN(n5976) );
  XOR2_X1 U11973 ( .A1(n3416), .A2(n5977), .Z(\MC_ARK_ARC_1_0/buf_output[80] )
         );
  XOR2_X1 U11974 ( .A1(n1429), .A2(\MC_ARK_ARC_1_0/temp2[80] ), .Z(n5977) );
  INV_X1 U11975 ( .I(\SB3_12/buf_output[5] ), .ZN(\SB4_12/i1_5 ) );
  NAND4_X2 U11976 ( .A1(\SB3_12/Component_Function_5/NAND4_in[2] ), .A2(n913), 
        .A3(\SB3_12/Component_Function_5/NAND4_in[1] ), .A4(n1613), .ZN(
        \SB3_12/buf_output[5] ) );
  NAND4_X2 U11977 ( .A1(\SB2_1_3/Component_Function_5/NAND4_in[2] ), .A2(n5994), .A3(n1421), .A4(n6085), .ZN(\SB2_1_3/buf_output[5] ) );
  NAND3_X1 U11978 ( .A1(\SB1_1_2/i0[10] ), .A2(\SB1_1_2/i1[9] ), .A3(
        \SB1_1_2/i1_5 ), .ZN(\SB1_1_2/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U11979 ( .A1(n5503), .A2(\RI5[3][65] ), .Z(n6132) );
  XOR2_X1 U11980 ( .A1(\RI5[3][26] ), .A2(\RI5[3][2] ), .Z(
        \MC_ARK_ARC_1_3/temp2[56] ) );
  NAND4_X2 U11981 ( .A1(n1570), .A2(n6345), .A3(
        \SB1_3_2/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_3_2/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_2/buf_output[5] ) );
  NAND4_X2 U11982 ( .A1(n6358), .A2(
        \SB1_3_16/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_3_16/Component_Function_1/NAND4_in[1] ), .A4(
        \SB1_3_16/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_3_16/buf_output[1] ) );
  INV_X2 U11983 ( .I(\SB1_3_14/buf_output[5] ), .ZN(\SB2_3_14/i1_5 ) );
  NAND4_X2 U11984 ( .A1(n3746), .A2(n6023), .A3(n941), .A4(
        \SB1_3_14/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_14/buf_output[5] ) );
  NAND3_X2 U11985 ( .A1(\SB1_2_14/i0_3 ), .A2(\SB1_2_14/i1[9] ), .A3(
        \SB1_2_14/i0[6] ), .ZN(\SB1_2_14/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U11986 ( .A1(\SB3_22/i3[0] ), .A2(\SB3_22/i1_5 ), .A3(
        \SB3_22/i0[8] ), .ZN(n2215) );
  NAND3_X2 U11987 ( .A1(\SB2_2_27/i0[10] ), .A2(\SB2_2_27/i1_5 ), .A3(
        \SB2_2_27/i1[9] ), .ZN(\SB2_2_27/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U11988 ( .A1(\SB1_2_4/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_2_4/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_4/Component_Function_1/NAND4_in[0] ), .A4(n5979), .ZN(
        \SB1_2_4/buf_output[1] ) );
  XOR2_X1 U11989 ( .A1(n5981), .A2(n5980), .Z(n2568) );
  XOR2_X1 U11990 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[83] ), .A2(\RI5[2][89] ), 
        .Z(n5980) );
  XOR2_X1 U11991 ( .A1(\RI5[2][35] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[59] ), 
        .Z(n5981) );
  NAND3_X2 U11992 ( .A1(\SB2_2_13/i0_0 ), .A2(n580), .A3(\SB2_2_13/i0_3 ), 
        .ZN(n5983) );
  NAND4_X2 U11993 ( .A1(\SB1_2_14/Component_Function_1/NAND4_in[0] ), .A2(
        \SB1_2_14/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_2_14/Component_Function_1/NAND4_in[2] ), .A4(n5984), .ZN(
        \SB1_2_14/buf_output[1] ) );
  XOR2_X1 U11994 ( .A1(\RI5[1][172] ), .A2(\RI5[1][16] ), .Z(
        \MC_ARK_ARC_1_1/temp3[106] ) );
  XOR2_X1 U11995 ( .A1(n3826), .A2(n5988), .Z(\MC_ARK_ARC_1_3/temp5[10] ) );
  XOR2_X1 U11996 ( .A1(\RI5[3][4] ), .A2(\RI5[3][172] ), .Z(n5988) );
  NAND3_X1 U11997 ( .A1(\SB1_3_22/i0[6] ), .A2(\SB1_3_22/i0[8] ), .A3(
        \SB1_3_22/i0[7] ), .ZN(\SB1_3_22/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U11998 ( .A1(\RI3[0][178] ), .A2(\RI3[0][176] ), .A3(\SB2_0_2/i1_5 ), .ZN(\SB2_0_2/Component_Function_2/NAND4_in[3] ) );
  XOR2_X1 U11999 ( .A1(\MC_ARK_ARC_1_2/temp3[177] ), .A2(
        \MC_ARK_ARC_1_2/temp4[177] ), .Z(\MC_ARK_ARC_1_2/temp6[177] ) );
  NAND4_X2 U12000 ( .A1(\SB2_3_31/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_3_31/Component_Function_4/NAND4_in[3] ), .A3(n6049), .A4(n5990), 
        .ZN(\SB2_3_31/buf_output[4] ) );
  NAND3_X1 U12001 ( .A1(\SB2_3_31/i0_0 ), .A2(\SB2_3_31/i3[0] ), .A3(
        \SB2_3_31/i1_7 ), .ZN(n5990) );
  XOR2_X1 U12002 ( .A1(n3039), .A2(\MC_ARK_ARC_1_1/temp2[163] ), .Z(n4614) );
  NAND4_X2 U12003 ( .A1(\SB3_6/Component_Function_1/NAND4_in[2] ), .A2(
        \SB3_6/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_6/Component_Function_1/NAND4_in[3] ), .A4(n5991), .ZN(
        \SB3_6/buf_output[1] ) );
  NAND2_X1 U12004 ( .A1(\RI1[4][155] ), .A2(\SB3_6/i1[9] ), .ZN(n5991) );
  NAND4_X2 U12005 ( .A1(\SB1_2_4/Component_Function_0/NAND4_in[2] ), .A2(
        \SB1_2_4/Component_Function_0/NAND4_in[3] ), .A3(
        \SB1_2_4/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_2_4/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_2_4/buf_output[0] ) );
  NAND4_X2 U12006 ( .A1(\SB1_3_24/Component_Function_5/NAND4_in[0] ), .A2(
        \SB1_3_24/Component_Function_5/NAND4_in[2] ), .A3(n6074), .A4(n1341), 
        .ZN(\SB1_3_24/buf_output[5] ) );
  NAND4_X2 U12007 ( .A1(\SB1_1_8/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_8/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_1_8/Component_Function_5/NAND4_in[3] ), .A4(
        \SB1_1_8/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_8/buf_output[5] ) );
  NAND3_X1 U12008 ( .A1(\SB1_3_14/i0_0 ), .A2(\SB1_3_14/i0[8] ), .A3(
        \SB1_3_14/i0[9] ), .ZN(n5992) );
  XOR2_X1 U12009 ( .A1(n5993), .A2(n5), .Z(Ciphertext[72]) );
  NAND4_X2 U12010 ( .A1(\SB4_19/Component_Function_0/NAND4_in[1] ), .A2(
        \SB4_19/Component_Function_0/NAND4_in[2] ), .A3(n6098), .A4(
        \SB4_19/Component_Function_0/NAND4_in[0] ), .ZN(n5993) );
  NAND3_X1 U12011 ( .A1(\SB3_13/i0_4 ), .A2(\SB3_13/i1_5 ), .A3(
        \MC_ARK_ARC_1_3/buf_output[110] ), .ZN(
        \SB3_13/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 U12012 ( .A1(\SB2_1_3/i0[6] ), .A2(\SB2_1_3/i0_0 ), .A3(
        \SB2_1_3/i0[10] ), .ZN(n5994) );
  NAND4_X2 U12013 ( .A1(\SB2_3_29/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_3_29/Component_Function_1/NAND4_in[0] ), .A3(n4334), .A4(n5995), 
        .ZN(\SB2_3_29/buf_output[1] ) );
  NAND3_X2 U12014 ( .A1(\SB2_3_29/i0_3 ), .A2(\SB2_3_29/i0[8] ), .A3(
        \SB2_3_29/i1_7 ), .ZN(n5995) );
  INV_X2 U12015 ( .I(\SB1_2_17/buf_output[3] ), .ZN(\SB2_2_15/i0[8] ) );
  NAND4_X2 U12016 ( .A1(\SB1_2_17/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_17/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_2_17/Component_Function_3/NAND4_in[2] ), .A4(n1750), .ZN(
        \SB1_2_17/buf_output[3] ) );
  NAND3_X2 U12017 ( .A1(\SB2_3_26/i0[9] ), .A2(n4750), .A3(\SB2_3_26/i0_3 ), 
        .ZN(n5996) );
  XOR2_X1 U12018 ( .A1(n5998), .A2(n5997), .Z(n6238) );
  XOR2_X1 U12019 ( .A1(\RI5[1][17] ), .A2(\RI5[1][59] ), .Z(n5997) );
  XOR2_X1 U12020 ( .A1(\RI5[1][23] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[89] ), 
        .Z(n5998) );
  NAND3_X2 U12021 ( .A1(\SB2_1_3/i0[6] ), .A2(\SB2_1_3/i0_3 ), .A3(
        \SB2_1_3/i1[9] ), .ZN(\SB2_1_3/Component_Function_3/NAND4_in[0] ) );
  INV_X2 U12022 ( .I(\SB1_3_7/buf_output[3] ), .ZN(\SB2_3_5/i0[8] ) );
  NAND4_X2 U12023 ( .A1(\SB1_3_7/Component_Function_3/NAND4_in[1] ), .A2(n3972), .A3(n6297), .A4(\SB1_3_7/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_3_7/buf_output[3] ) );
  NAND4_X2 U12024 ( .A1(\SB1_0_23/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_0_23/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_0_23/Component_Function_1/NAND4_in[1] ), .A4(
        \SB1_0_23/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_0_23/buf_output[1] ) );
  NAND4_X2 U12025 ( .A1(\SB2_0_7/Component_Function_4/NAND4_in[0] ), .A2(n6000), .A3(\SB2_0_7/Component_Function_4/NAND4_in[3] ), .A4(
        \SB2_0_7/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB2_0_7/buf_output[4] ) );
  NAND4_X2 U12026 ( .A1(\SB3_25/Component_Function_3/NAND4_in[1] ), .A2(n6160), 
        .A3(n6446), .A4(n6001), .ZN(\SB3_25/buf_output[3] ) );
  NAND4_X2 U12027 ( .A1(\SB2_1_7/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_7/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_1_7/Component_Function_2/NAND4_in[1] ), .A4(n6002), .ZN(
        \SB2_1_7/buf_output[2] ) );
  NAND3_X2 U12028 ( .A1(\SB2_1_7/i0_0 ), .A2(n5790), .A3(\SB2_1_7/i1_5 ), .ZN(
        n6002) );
  XOR2_X1 U12029 ( .A1(n2751), .A2(n6003), .Z(\MC_ARK_ARC_1_2/buf_output[90] )
         );
  NAND2_X1 U12030 ( .A1(n2221), .A2(
        \SB1_3_27/Component_Function_4/NAND4_in[1] ), .ZN(n2244) );
  NAND3_X1 U12031 ( .A1(\SB3_2/i0[6] ), .A2(\SB3_2/i0[10] ), .A3(\SB3_2/i0_3 ), 
        .ZN(\SB3_2/Component_Function_2/NAND4_in[1] ) );
  XOR2_X1 U12032 ( .A1(\MC_ARK_ARC_1_3/temp3[89] ), .A2(
        \MC_ARK_ARC_1_3/temp4[89] ), .Z(n626) );
  XOR2_X1 U12033 ( .A1(n2895), .A2(\SB2_3_22/buf_output[0] ), .Z(
        \MC_ARK_ARC_1_3/temp1[90] ) );
  XOR2_X1 U12034 ( .A1(\MC_ARK_ARC_1_2/temp4[110] ), .A2(
        \MC_ARK_ARC_1_2/temp3[110] ), .Z(n4454) );
  NAND4_X2 U12035 ( .A1(\SB1_1_6/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_1_6/Component_Function_1/NAND4_in[2] ), .A3(
        \SB1_1_6/Component_Function_1/NAND4_in[3] ), .A4(
        \SB1_1_6/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_1_6/buf_output[1] ) );
  XOR2_X1 U12036 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[39] ), .A2(\RI5[2][75] ), 
        .Z(n6004) );
  NAND4_X2 U12037 ( .A1(\SB1_3_30/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_3_30/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_3_30/Component_Function_1/NAND4_in[0] ), .A4(n6005), .ZN(
        \SB1_3_30/buf_output[1] ) );
  NAND3_X1 U12038 ( .A1(\SB1_3_30/i0[6] ), .A2(\SB1_3_30/i0[9] ), .A3(
        \SB1_3_30/i1_5 ), .ZN(n6005) );
  XOR2_X1 U12039 ( .A1(\RI5[2][63] ), .A2(\RI5[2][87] ), .Z(
        \MC_ARK_ARC_1_2/temp2[117] ) );
  NAND4_X2 U12040 ( .A1(\SB1_1_8/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_1_8/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_1_8/Component_Function_1/NAND4_in[3] ), .A4(
        \SB1_1_8/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_1_8/buf_output[1] ) );
  NAND3_X1 U12041 ( .A1(\SB2_1_18/i0_3 ), .A2(\SB1_1_22/buf_output[1] ), .A3(
        \SB2_1_18/i1[9] ), .ZN(\SB2_1_18/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U12042 ( .A1(\SB3_13/i0[6] ), .A2(\SB3_13/i0[10] ), .A3(
        \MC_ARK_ARC_1_3/buf_output[110] ), .ZN(
        \SB3_13/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U12043 ( .A1(n3782), .A2(n6006), .Z(\MC_ARK_ARC_1_2/buf_output[33] )
         );
  XOR2_X1 U12044 ( .A1(\MC_ARK_ARC_1_2/temp4[33] ), .A2(
        \MC_ARK_ARC_1_2/temp3[33] ), .Z(n6006) );
  INV_X2 U12045 ( .I(\SB1_3_12/buf_output[3] ), .ZN(\SB2_3_10/i0[8] ) );
  NAND4_X2 U12046 ( .A1(\SB1_3_12/Component_Function_3/NAND4_in[2] ), .A2(
        n3360), .A3(n6462), .A4(\SB1_3_12/Component_Function_3/NAND4_in[3] ), 
        .ZN(\SB1_3_12/buf_output[3] ) );
  NAND3_X2 U12047 ( .A1(\SB2_2_28/i0_3 ), .A2(\SB2_2_28/i1[9] ), .A3(
        \SB2_2_28/i0_4 ), .ZN(n1741) );
  NAND4_X2 U12048 ( .A1(\SB2_2_16/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_16/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_2_16/Component_Function_2/NAND4_in[1] ), .A4(n6007), .ZN(
        \SB2_2_16/buf_output[2] ) );
  NAND3_X2 U12049 ( .A1(\SB2_2_16/i0_0 ), .A2(\SB2_2_16/i1_5 ), .A3(
        \SB2_2_16/i0_4 ), .ZN(n6007) );
  XOR2_X1 U12050 ( .A1(\MC_ARK_ARC_1_2/temp5[59] ), .A2(n6008), .Z(
        \RI1[3][59] ) );
  NAND4_X2 U12051 ( .A1(\SB1_2_24/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_2_24/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_2_24/Component_Function_1/NAND4_in[0] ), .A4(
        \SB1_2_24/Component_Function_1/NAND4_in[1] ), .ZN(
        \SB1_2_24/buf_output[1] ) );
  NAND3_X2 U12052 ( .A1(\SB2_2_22/i0[10] ), .A2(\SB2_2_22/i1[9] ), .A3(
        \SB2_2_22/i1_7 ), .ZN(n6009) );
  XOR2_X1 U12053 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[45] ), .A2(\RI5[2][69] ), 
        .Z(n4067) );
  NAND4_X2 U12054 ( .A1(\SB2_1_2/Component_Function_1/NAND4_in[3] ), .A2(n1851), .A3(n3710), .A4(\SB2_1_2/Component_Function_1/NAND4_in[2] ), .ZN(
        \SB2_1_2/buf_output[1] ) );
  XOR2_X1 U12055 ( .A1(\RI5[0][174] ), .A2(\RI5[0][168] ), .Z(
        \MC_ARK_ARC_1_0/temp1[174] ) );
  XOR2_X1 U12056 ( .A1(\MC_ARK_ARC_1_1/temp6[47] ), .A2(n1354), .Z(
        \MC_ARK_ARC_1_1/buf_output[47] ) );
  XOR2_X1 U12057 ( .A1(n6389), .A2(n3213), .Z(\MC_ARK_ARC_1_0/buf_output[174] ) );
  NAND3_X2 U12058 ( .A1(\SB2_1_25/i0_3 ), .A2(\SB2_1_25/i0[9] ), .A3(
        \SB2_1_25/i0[8] ), .ZN(n3612) );
  XOR2_X1 U12059 ( .A1(\MC_ARK_ARC_1_0/temp2[36] ), .A2(
        \MC_ARK_ARC_1_0/temp1[36] ), .Z(\MC_ARK_ARC_1_0/temp5[36] ) );
  NAND3_X2 U12060 ( .A1(\SB2_1_15/i1_5 ), .A2(\SB2_1_15/i1[9] ), .A3(
        \SB2_1_15/i0_4 ), .ZN(n6081) );
  XOR2_X1 U12061 ( .A1(\MC_ARK_ARC_1_2/temp5[51] ), .A2(n6013), .Z(
        \MC_ARK_ARC_1_2/buf_output[51] ) );
  XOR2_X1 U12062 ( .A1(\MC_ARK_ARC_1_2/temp3[51] ), .A2(
        \MC_ARK_ARC_1_2/temp4[51] ), .Z(n6013) );
  NAND3_X2 U12063 ( .A1(\SB2_2_8/i0_3 ), .A2(\SB2_2_8/i0_4 ), .A3(
        \SB2_2_8/i0_0 ), .ZN(\SB2_2_8/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U12064 ( .A1(\SB2_0_29/buf_output[3] ), .A2(\RI5[0][183] ), .Z(
        \MC_ARK_ARC_1_0/temp3[117] ) );
  XOR2_X1 U12065 ( .A1(n2587), .A2(n6014), .Z(\MC_ARK_ARC_1_1/buf_output[60] )
         );
  XOR2_X1 U12066 ( .A1(\MC_ARK_ARC_1_1/temp3[60] ), .A2(
        \MC_ARK_ARC_1_1/temp4[60] ), .Z(n6014) );
  XOR2_X1 U12067 ( .A1(\RI5[2][155] ), .A2(\RI5[2][119] ), .Z(
        \MC_ARK_ARC_1_2/temp3[53] ) );
  NAND3_X2 U12068 ( .A1(\SB2_1_10/i0_3 ), .A2(\SB2_1_10/i0_0 ), .A3(
        \SB1_1_11/buf_output[4] ), .ZN(n6015) );
  NAND4_X2 U12069 ( .A1(\SB2_1_7/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_7/Component_Function_5/NAND4_in[0] ), .A3(n3308), .A4(n6017), 
        .ZN(\SB2_1_7/buf_output[5] ) );
  NAND3_X2 U12070 ( .A1(\SB2_1_7/i0[10] ), .A2(\SB2_1_7/i0_0 ), .A3(n2852), 
        .ZN(n6017) );
  NAND4_X2 U12071 ( .A1(\SB2_3_7/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_3_7/Component_Function_0/NAND4_in[0] ), .A3(
        \SB2_3_7/Component_Function_0/NAND4_in[3] ), .A4(n6019), .ZN(
        \SB2_3_7/buf_output[0] ) );
  NAND3_X1 U12072 ( .A1(\SB2_3_7/i0_3 ), .A2(\SB2_3_7/i0[10] ), .A3(
        \SB1_3_8/buf_output[4] ), .ZN(n6019) );
  NAND3_X2 U12073 ( .A1(\SB2_0_22/i0[10] ), .A2(\SB2_0_22/i1_5 ), .A3(
        \SB2_0_22/i1[9] ), .ZN(\SB2_0_22/Component_Function_2/NAND4_in[0] ) );
  INV_X2 U12074 ( .I(\SB1_1_19/buf_output[2] ), .ZN(\SB2_1_16/i1[9] ) );
  XOR2_X1 U12075 ( .A1(n2062), .A2(n6021), .Z(\MC_ARK_ARC_1_1/buf_output[74] )
         );
  XOR2_X1 U12076 ( .A1(\MC_ARK_ARC_1_1/temp4[74] ), .A2(n6069), .Z(n6021) );
  NAND3_X1 U12077 ( .A1(\SB1_3_7/i0_4 ), .A2(\SB1_3_7/i1_5 ), .A3(
        \MC_ARK_ARC_1_2/buf_output[146] ), .ZN(n6022) );
  NAND3_X2 U12078 ( .A1(\SB1_3_14/i0[10] ), .A2(\SB1_3_14/i0[6] ), .A3(
        \SB1_3_14/i0_0 ), .ZN(n6023) );
  XOR2_X1 U12079 ( .A1(\RI5[0][19] ), .A2(\RI5[0][55] ), .Z(
        \MC_ARK_ARC_1_0/temp3[145] ) );
  BUF_X4 U12080 ( .I(\SB2_1_19/buf_output[2] ), .Z(\RI5[1][92] ) );
  NAND3_X2 U12081 ( .A1(\SB1_2_2/i0_3 ), .A2(\SB1_2_2/i0_4 ), .A3(
        \SB1_2_2/i1[9] ), .ZN(\SB1_2_2/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U12082 ( .A1(\SB2_2_25/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_2_25/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_2_25/Component_Function_2/NAND4_in[1] ), .A4(
        \SB2_2_25/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_2_25/buf_output[2] ) );
  XOR2_X1 U12083 ( .A1(\RI5[1][5] ), .A2(\RI5[1][161] ), .Z(
        \MC_ARK_ARC_1_1/temp3[95] ) );
  NAND3_X2 U12084 ( .A1(\SB1_1_31/i1[9] ), .A2(\SB1_1_31/i0_4 ), .A3(
        \SB1_1_31/i0_3 ), .ZN(n6024) );
  INV_X4 U12085 ( .I(n6025), .ZN(\SB4_31/i0[10] ) );
  XOR2_X1 U12086 ( .A1(\MC_ARK_ARC_1_3/temp2[82] ), .A2(n6026), .Z(
        \MC_ARK_ARC_1_3/temp5[82] ) );
  XOR2_X1 U12087 ( .A1(\RI5[3][76] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[82] ), 
        .Z(n6026) );
  NAND4_X2 U12088 ( .A1(n4200), .A2(\SB3_18/Component_Function_5/NAND4_in[2] ), 
        .A3(n6426), .A4(\SB3_18/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB3_18/buf_output[5] ) );
  NAND3_X1 U12089 ( .A1(\SB1_2_20/i0_4 ), .A2(\SB1_2_20/i0_0 ), .A3(
        \SB1_2_20/i0_3 ), .ZN(\SB1_2_20/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U12090 ( .A1(\SB2_3_29/i0[10] ), .A2(\SB2_3_29/i1[9] ), .A3(
        \SB2_3_29/i1_7 ), .ZN(\SB2_3_29/Component_Function_3/NAND4_in[2] ) );
  NAND3_X1 U12091 ( .A1(\SB1_2_2/i0_3 ), .A2(\SB1_2_2/i0[6] ), .A3(
        \SB1_2_2/i1[9] ), .ZN(\SB1_2_2/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U12092 ( .A1(\SB3_1/i1_5 ), .A2(\MC_ARK_ARC_1_3/buf_output[182] ), 
        .A3(\MC_ARK_ARC_1_3/buf_output[184] ), .ZN(n4092) );
  XOR2_X1 U12093 ( .A1(\RI5[2][84] ), .A2(\RI5[2][90] ), .Z(n6030) );
  XOR2_X1 U12094 ( .A1(n6031), .A2(n133), .Z(Ciphertext[65]) );
  NAND4_X2 U12095 ( .A1(\SB4_21/Component_Function_5/NAND4_in[1] ), .A2(
        \SB4_21/Component_Function_5/NAND4_in[2] ), .A3(
        \SB4_21/Component_Function_5/NAND4_in[3] ), .A4(
        \SB4_21/Component_Function_5/NAND4_in[0] ), .ZN(n6031) );
  NAND4_X2 U12096 ( .A1(\SB1_0_30/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_30/Component_Function_3/NAND4_in[1] ), .A3(
        \SB1_0_30/Component_Function_3/NAND4_in[3] ), .A4(n6032), .ZN(
        \SB1_0_30/buf_output[3] ) );
  NAND3_X1 U12097 ( .A1(\SB1_0_30/i0[10] ), .A2(\SB1_0_30/i1[9] ), .A3(
        \SB1_0_30/i1_7 ), .ZN(n6032) );
  XOR2_X1 U12098 ( .A1(\RI5[1][141] ), .A2(\RI5[1][117] ), .Z(
        \MC_ARK_ARC_1_1/temp2[171] ) );
  NAND3_X2 U12099 ( .A1(\SB2_1_14/i0_3 ), .A2(\SB2_1_14/i1[9] ), .A3(
        \SB2_1_14/i0[6] ), .ZN(\SB2_1_14/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U12100 ( .A1(\MC_ARK_ARC_1_3/temp1[152] ), .A2(
        \MC_ARK_ARC_1_3/temp2[152] ), .Z(\MC_ARK_ARC_1_3/temp5[152] ) );
  XOR2_X1 U12101 ( .A1(n6033), .A2(n949), .Z(\MC_ARK_ARC_1_0/buf_output[104] )
         );
  XOR2_X1 U12102 ( .A1(\MC_ARK_ARC_1_0/temp4[104] ), .A2(n3309), .Z(n6033) );
  XOR2_X1 U12103 ( .A1(\MC_ARK_ARC_1_3/temp1[79] ), .A2(n6034), .Z(
        \MC_ARK_ARC_1_3/temp5[79] ) );
  XOR2_X1 U12104 ( .A1(\RI5[3][25] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[49] ), 
        .Z(n6034) );
  XOR2_X1 U12105 ( .A1(n6035), .A2(n61), .Z(Ciphertext[93]) );
  NAND4_X2 U12106 ( .A1(\SB4_16/Component_Function_3/NAND4_in[3] ), .A2(n2411), 
        .A3(n3622), .A4(\SB4_16/Component_Function_3/NAND4_in[2] ), .ZN(n6035)
         );
  NAND3_X1 U12107 ( .A1(\SB3_21/i0_3 ), .A2(\SB3_21/i0[10] ), .A3(
        \SB3_21/i0_4 ), .ZN(\SB3_21/Component_Function_0/NAND4_in[2] ) );
  NAND4_X2 U12108 ( .A1(\SB1_3_14/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_3_14/Component_Function_3/NAND4_in[0] ), .A3(n6216), .A4(n6036), 
        .ZN(\SB1_3_14/buf_output[3] ) );
  NAND3_X1 U12109 ( .A1(\SB1_2_20/i0[10] ), .A2(\SB1_2_20/i0_0 ), .A3(
        \SB1_2_20/i0[6] ), .ZN(\SB1_2_20/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U12110 ( .A1(\SB2_3_20/i1_7 ), .A2(\SB2_3_20/i0[8] ), .A3(
        \SB2_3_20/i0_4 ), .ZN(n3054) );
  XOR2_X1 U12111 ( .A1(\MC_ARK_ARC_1_0/temp1[175] ), .A2(
        \MC_ARK_ARC_1_0/temp2[175] ), .Z(\MC_ARK_ARC_1_0/temp5[175] ) );
  XOR2_X1 U12112 ( .A1(\RI5[2][5] ), .A2(\RI5[2][161] ), .Z(n6038) );
  XOR2_X1 U12113 ( .A1(n6039), .A2(\MC_ARK_ARC_1_3/temp3[188] ), .Z(n2355) );
  XOR2_X1 U12114 ( .A1(\RI5[3][158] ), .A2(\RI5[3][134] ), .Z(n6039) );
  XOR2_X1 U12115 ( .A1(n6040), .A2(\MC_ARK_ARC_1_3/temp4[25] ), .Z(n1998) );
  XOR2_X1 U12116 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[91] ), .A2(\RI5[3][127] ), 
        .Z(n6040) );
  XOR2_X1 U12117 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[71] ), .A2(\RI5[3][35] ), 
        .Z(n6041) );
  XOR2_X1 U12118 ( .A1(n6095), .A2(\MC_ARK_ARC_1_0/temp4[105] ), .Z(
        \MC_ARK_ARC_1_0/temp6[105] ) );
  XOR2_X1 U12119 ( .A1(n2752), .A2(\MC_ARK_ARC_1_0/temp5[135] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[135] ) );
  XOR2_X1 U12120 ( .A1(\MC_ARK_ARC_1_0/temp4[135] ), .A2(
        \MC_ARK_ARC_1_0/temp3[135] ), .Z(n2752) );
  NAND3_X1 U12121 ( .A1(\SB2_2_10/i0_3 ), .A2(n581), .A3(\SB2_2_10/i1[9] ), 
        .ZN(\SB2_2_10/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U12122 ( .A1(\SB2_1_2/i0_4 ), .A2(\SB2_1_2/i0_0 ), .A3(
        \SB2_1_2/i0_3 ), .ZN(\SB2_1_2/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U12123 ( .A1(\SB1_3_15/i0_0 ), .A2(\SB1_3_15/i0_4 ), .A3(
        \SB1_3_15/i0_3 ), .ZN(\SB1_3_15/Component_Function_3/NAND4_in[1] ) );
  NAND4_X2 U12124 ( .A1(\SB1_0_11/Component_Function_5/NAND4_in[1] ), .A2(
        n1241), .A3(\SB1_0_11/Component_Function_5/NAND4_in[0] ), .A4(
        \SB1_0_11/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB1_0_11/buf_output[5] ) );
  NAND4_X2 U12125 ( .A1(\SB4_12/Component_Function_2/NAND4_in[0] ), .A2(
        \SB4_12/Component_Function_2/NAND4_in[2] ), .A3(n2406), .A4(n4562), 
        .ZN(n6144) );
  XOR2_X1 U12126 ( .A1(\RI5[1][126] ), .A2(\RI5[1][132] ), .Z(
        \MC_ARK_ARC_1_1/temp1[132] ) );
  NAND4_X2 U12127 ( .A1(n1696), .A2(n6070), .A3(
        \SB1_1_15/Component_Function_5/NAND4_in[1] ), .A4(
        \SB1_1_15/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_15/buf_output[5] ) );
  NAND3_X1 U12128 ( .A1(\SB4_18/i0_0 ), .A2(\SB4_18/i0_3 ), .A3(\SB4_18/i0[7] ), .ZN(\SB4_18/Component_Function_0/NAND4_in[3] ) );
  NAND4_X2 U12129 ( .A1(\SB3_31/Component_Function_5/NAND4_in[3] ), .A2(
        \SB3_31/Component_Function_5/NAND4_in[1] ), .A3(
        \SB3_31/Component_Function_5/NAND4_in[2] ), .A4(
        \SB3_31/Component_Function_5/NAND4_in[0] ), .ZN(\SB3_31/buf_output[5] ) );
  NAND3_X2 U12130 ( .A1(\SB3_31/i0_3 ), .A2(\SB3_31/i1[9] ), .A3(
        \SB3_31/i0[6] ), .ZN(\SB3_31/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U12131 ( .A1(\SB4_12/i0_4 ), .A2(\SB4_12/i1[9] ), .A3(\SB4_12/i1_5 ), .ZN(\SB4_12/Component_Function_4/NAND4_in[3] ) );
  NAND3_X2 U12132 ( .A1(\SB2_3_14/i0[10] ), .A2(\SB2_3_14/i0_0 ), .A3(
        \SB2_3_14/i0[6] ), .ZN(n6043) );
  NAND4_X2 U12133 ( .A1(\SB2_3_13/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_3_13/Component_Function_2/NAND4_in[0] ), .A3(
        \SB2_3_13/Component_Function_2/NAND4_in[3] ), .A4(n3236), .ZN(
        \SB2_3_13/buf_output[2] ) );
  NAND4_X2 U12134 ( .A1(\SB1_3_9/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_3_9/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_3_9/Component_Function_5/NAND4_in[3] ), .A4(
        \SB1_3_9/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_9/buf_output[5] ) );
  XOR2_X1 U12135 ( .A1(n1257), .A2(\MC_ARK_ARC_1_3/temp5[115] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[115] ) );
  NAND4_X2 U12136 ( .A1(\SB1_1_12/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_1_12/Component_Function_3/NAND4_in[2] ), .A3(n6157), .A4(n1120), 
        .ZN(\SB1_1_12/buf_output[3] ) );
  NAND4_X2 U12137 ( .A1(n4582), .A2(\SB2_2_2/Component_Function_2/NAND4_in[2] ), .A3(n6150), .A4(n3771), .ZN(\SB2_2_2/buf_output[2] ) );
  NAND3_X2 U12138 ( .A1(\SB3_12/i0[9] ), .A2(\SB3_12/i0[6] ), .A3(
        \SB3_12/i0_4 ), .ZN(n913) );
  NAND3_X2 U12139 ( .A1(\SB1_2_27/i0_4 ), .A2(\SB1_2_27/i0[6] ), .A3(
        \SB1_2_27/i0[9] ), .ZN(n6045) );
  XOR2_X1 U12140 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[59] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[53] ), .Z(\MC_ARK_ARC_1_2/temp1[59] ) );
  XOR2_X1 U12141 ( .A1(\RI5[1][40] ), .A2(\RI5[1][64] ), .Z(
        \MC_ARK_ARC_1_1/temp2[94] ) );
  XOR2_X1 U12142 ( .A1(\RI5[2][10] ), .A2(\RI5[2][46] ), .Z(
        \MC_ARK_ARC_1_2/temp3[136] ) );
  NAND3_X1 U12143 ( .A1(\SB3_14/i0_3 ), .A2(\SB3_14/i0_0 ), .A3(\SB3_14/i0_4 ), 
        .ZN(\SB3_14/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U12144 ( .A1(\MC_ARK_ARC_1_3/temp1[176] ), .A2(
        \MC_ARK_ARC_1_3/temp2[176] ), .Z(\MC_ARK_ARC_1_3/temp5[176] ) );
  XOR2_X1 U12145 ( .A1(n1299), .A2(\MC_ARK_ARC_1_1/temp6[25] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[25] ) );
  XOR2_X1 U12146 ( .A1(\MC_ARK_ARC_1_3/temp5[116] ), .A2(
        \MC_ARK_ARC_1_3/temp6[116] ), .Z(\MC_ARK_ARC_1_3/buf_output[116] ) );
  XOR2_X1 U12147 ( .A1(\MC_ARK_ARC_1_2/temp6[124] ), .A2(
        \MC_ARK_ARC_1_2/temp5[124] ), .Z(\MC_ARK_ARC_1_2/buf_output[124] ) );
  NAND3_X2 U12148 ( .A1(\SB2_1_11/i0[10] ), .A2(\SB2_1_11/i1[9] ), .A3(
        \SB2_1_11/i1_7 ), .ZN(\SB2_1_11/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U12149 ( .A1(\SB2_2_17/i3[0] ), .A2(\SB2_2_17/i0[8] ), .A3(
        \SB2_2_17/i1_5 ), .ZN(\SB2_2_17/Component_Function_3/NAND4_in[3] ) );
  NAND3_X1 U12150 ( .A1(\SB1_2_7/i0_3 ), .A2(\SB1_2_7/i0[8] ), .A3(
        \SB1_2_7/i1_7 ), .ZN(\SB1_2_7/Component_Function_1/NAND4_in[1] ) );
  NAND3_X2 U12151 ( .A1(\SB3_2/i0[6] ), .A2(\SB3_2/i0[9] ), .A3(\SB3_2/i0_4 ), 
        .ZN(n4136) );
  NAND4_X2 U12152 ( .A1(\SB2_1_23/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_1_23/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_1_23/Component_Function_0/NAND4_in[1] ), .A4(
        \SB2_1_23/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_1_23/buf_output[0] ) );
  NAND2_X1 U12153 ( .A1(\SB4_7/i0[9] ), .A2(\SB4_7/i0[10] ), .ZN(
        \SB4_7/Component_Function_0/NAND4_in[0] ) );
  NAND4_X2 U12154 ( .A1(\SB3_12/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_12/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_12/Component_Function_0/NAND4_in[0] ), .A4(n6046), .ZN(
        \SB3_12/buf_output[0] ) );
  NAND3_X1 U12155 ( .A1(\SB3_12/i0_3 ), .A2(\SB3_12/i0_0 ), .A3(\SB3_12/i0[7] ), .ZN(n6046) );
  NAND3_X2 U12156 ( .A1(\SB2_1_6/i0[10] ), .A2(\SB2_1_6/i1_7 ), .A3(
        \SB2_1_6/i1[9] ), .ZN(\SB2_1_6/Component_Function_3/NAND4_in[2] ) );
  NAND4_X2 U12157 ( .A1(\SB3_22/Component_Function_5/NAND4_in[1] ), .A2(
        \SB3_22/Component_Function_5/NAND4_in[2] ), .A3(
        \SB3_22/Component_Function_5/NAND4_in[0] ), .A4(n6047), .ZN(
        \SB3_22/buf_output[5] ) );
  XOR2_X1 U12158 ( .A1(\MC_ARK_ARC_1_3/temp6[58] ), .A2(n6048), .Z(
        \MC_ARK_ARC_1_3/buf_output[58] ) );
  XOR2_X1 U12159 ( .A1(\MC_ARK_ARC_1_3/temp1[58] ), .A2(
        \MC_ARK_ARC_1_3/temp2[58] ), .Z(n6048) );
  NAND3_X1 U12160 ( .A1(\SB2_3_31/i0_0 ), .A2(\SB2_3_31/i0[9] ), .A3(
        \SB2_3_31/i0[8] ), .ZN(n6049) );
  XOR2_X1 U12161 ( .A1(\MC_ARK_ARC_1_1/temp2[84] ), .A2(n6050), .Z(n799) );
  XOR2_X1 U12162 ( .A1(\RI5[1][78] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[84] ), 
        .Z(n6050) );
  NAND3_X2 U12163 ( .A1(\SB4_31/i0_0 ), .A2(\SB4_31/i0[10] ), .A3(
        \SB4_31/i0[6] ), .ZN(n6051) );
  XOR2_X1 U12164 ( .A1(\MC_ARK_ARC_1_1/temp1[134] ), .A2(n1292), .Z(n4708) );
  NAND3_X2 U12165 ( .A1(\SB1_0_13/i0_0 ), .A2(\SB1_0_13/i0_3 ), .A3(
        \SB1_0_13/i0_4 ), .ZN(n6405) );
  NAND4_X2 U12166 ( .A1(\SB3_16/Component_Function_4/NAND4_in[1] ), .A2(
        \SB3_16/Component_Function_4/NAND4_in[0] ), .A3(
        \SB3_16/Component_Function_4/NAND4_in[2] ), .A4(n6052), .ZN(
        \SB3_16/buf_output[4] ) );
  NAND3_X1 U12167 ( .A1(\SB3_16/i0_4 ), .A2(\SB3_16/i1[9] ), .A3(\SB3_16/i1_5 ), .ZN(n6052) );
  NAND4_X2 U12168 ( .A1(\SB2_3_0/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_3_0/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_3_0/Component_Function_4/NAND4_in[1] ), .A4(n6053), .ZN(
        \SB2_3_0/buf_output[4] ) );
  NAND4_X2 U12169 ( .A1(\SB4_15/Component_Function_1/NAND4_in[2] ), .A2(
        \SB4_15/Component_Function_1/NAND4_in[1] ), .A3(
        \SB4_15/Component_Function_1/NAND4_in[0] ), .A4(n6054), .ZN(n4620) );
  NAND3_X1 U12170 ( .A1(\SB4_15/i0_4 ), .A2(\SB4_15/i1_7 ), .A3(\SB4_15/i0[8] ), .ZN(n6054) );
  XOR2_X1 U12171 ( .A1(n6055), .A2(\MC_ARK_ARC_1_3/temp4[116] ), .Z(
        \MC_ARK_ARC_1_3/temp6[116] ) );
  XOR2_X1 U12172 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[182] ), .A2(\RI5[3][26] ), 
        .Z(n6055) );
  XOR2_X1 U12173 ( .A1(n6056), .A2(n30), .Z(Ciphertext[83]) );
  NAND4_X2 U12174 ( .A1(\SB4_18/Component_Function_5/NAND4_in[2] ), .A2(n4251), 
        .A3(n6082), .A4(n876), .ZN(n6056) );
  XOR2_X1 U12175 ( .A1(\MC_ARK_ARC_1_3/temp3[90] ), .A2(
        \MC_ARK_ARC_1_3/temp4[90] ), .Z(n4146) );
  NAND3_X2 U12176 ( .A1(\SB2_1_13/i0[10] ), .A2(\SB2_1_13/i0_0 ), .A3(
        \SB2_1_13/i0[6] ), .ZN(\SB2_1_13/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U12177 ( .A1(\SB3_13/i0_3 ), .A2(\SB3_13/i0_4 ), .A3(
        \MC_ARK_ARC_1_3/buf_output[110] ), .ZN(n1420) );
  XOR2_X1 U12178 ( .A1(\MC_ARK_ARC_1_1/temp1[46] ), .A2(n6059), .Z(n3158) );
  XOR2_X1 U12179 ( .A1(\RI5[1][184] ), .A2(\RI5[1][16] ), .Z(n6059) );
  XOR2_X1 U12180 ( .A1(\RI5[0][0] ), .A2(\RI5[0][162] ), .Z(n6060) );
  NAND4_X2 U12181 ( .A1(\SB1_2_1/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_2_1/Component_Function_5/NAND4_in[1] ), .A3(n2972), .A4(
        \SB1_2_1/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_2_1/buf_output[5] ) );
  XOR2_X1 U12182 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[82] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[106] ), .Z(\MC_ARK_ARC_1_2/temp2[136] )
         );
  XOR2_X1 U12183 ( .A1(\RI5[3][67] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[103] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[1] ) );
  XOR2_X1 U12184 ( .A1(\MC_ARK_ARC_1_1/temp4[181] ), .A2(n4342), .Z(n6061) );
  NAND3_X2 U12185 ( .A1(\SB1_2_25/i3[0] ), .A2(\SB1_2_25/i1_5 ), .A3(
        \SB1_2_25/i0[8] ), .ZN(n6062) );
  NAND3_X1 U12186 ( .A1(\SB1_1_6/i0[8] ), .A2(\SB1_1_6/i0_3 ), .A3(
        \SB1_1_6/i1_7 ), .ZN(\SB1_1_6/Component_Function_1/NAND4_in[1] ) );
  NAND4_X2 U12187 ( .A1(n6315), .A2(n2236), .A3(
        \SB2_2_1/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_2_1/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB2_2_1/buf_output[4] ) );
  NAND3_X2 U12188 ( .A1(\SB1_1_14/i0[6] ), .A2(\SB1_1_14/i0_0 ), .A3(
        \SB1_1_14/i0[10] ), .ZN(\SB1_1_14/Component_Function_5/NAND4_in[1] )
         );
  NAND3_X2 U12189 ( .A1(\SB2_3_29/i0[10] ), .A2(\SB2_3_29/i0_3 ), .A3(
        \SB2_3_29/i0[6] ), .ZN(n6063) );
  INV_X2 U12190 ( .I(\SB3_0/buf_output[3] ), .ZN(\SB4_30/i0[8] ) );
  XOR2_X1 U12191 ( .A1(n6064), .A2(\MC_ARK_ARC_1_3/temp2[114] ), .Z(
        \MC_ARK_ARC_1_3/temp5[114] ) );
  XOR2_X1 U12192 ( .A1(\RI5[3][108] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[114] ), .Z(n6064) );
  NAND4_X2 U12193 ( .A1(n4056), .A2(\SB2_0_3/Component_Function_5/NAND4_in[1] ), .A3(\SB2_0_3/Component_Function_5/NAND4_in[0] ), .A4(n6065), .ZN(
        \SB2_0_3/buf_output[5] ) );
  NAND3_X2 U12194 ( .A1(\SB2_0_3/i0[9] ), .A2(\RI3[0][172] ), .A3(
        \SB2_0_3/i0[6] ), .ZN(n6065) );
  XOR2_X1 U12195 ( .A1(n6066), .A2(\MC_ARK_ARC_1_2/temp5[55] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[55] ) );
  XOR2_X1 U12196 ( .A1(\MC_ARK_ARC_1_2/temp4[55] ), .A2(n3130), .Z(n6066) );
  XOR2_X1 U12197 ( .A1(\RI5[1][121] ), .A2(\RI5[1][157] ), .Z(
        \MC_ARK_ARC_1_1/temp3[55] ) );
  NAND2_X1 U12198 ( .A1(\SB1_3_12/Component_Function_4/NAND4_in[1] ), .A2(
        n6067), .ZN(n1370) );
  XOR2_X1 U12199 ( .A1(\RI5[2][9] ), .A2(\RI5[2][3] ), .Z(n6068) );
  XOR2_X1 U12200 ( .A1(\RI5[1][140] ), .A2(\RI5[1][176] ), .Z(n6069) );
  NAND3_X2 U12201 ( .A1(\SB2_3_20/i0[10] ), .A2(\SB2_3_20/i1[9] ), .A3(
        \SB2_3_20/i1_5 ), .ZN(\SB2_3_20/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U12202 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[74] ), .A2(\RI5[1][68] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[74] ) );
  XOR2_X1 U12203 ( .A1(\MC_ARK_ARC_1_1/temp1[179] ), .A2(
        \MC_ARK_ARC_1_1/temp2[179] ), .Z(n6071) );
  XOR2_X1 U12204 ( .A1(n6072), .A2(n207), .Z(Ciphertext[79]) );
  NAND4_X2 U12205 ( .A1(\SB4_18/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_18/Component_Function_1/NAND4_in[3] ), .A3(n6096), .A4(
        \SB4_18/Component_Function_1/NAND4_in[0] ), .ZN(n6072) );
  XOR2_X1 U12206 ( .A1(\RI5[3][67] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[91] ), 
        .Z(n1796) );
  INV_X2 U12207 ( .I(\SB1_3_24/buf_output[3] ), .ZN(\SB2_3_22/i0[8] ) );
  NAND4_X2 U12208 ( .A1(\SB1_3_24/Component_Function_3/NAND4_in[0] ), .A2(
        n6375), .A3(\SB1_3_24/Component_Function_3/NAND4_in[2] ), .A4(
        \SB1_3_24/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_3_24/buf_output[3] ) );
  NAND3_X2 U12209 ( .A1(\SB1_3_24/i0_0 ), .A2(\SB1_3_24/i0[10] ), .A3(
        \SB1_3_24/i0[6] ), .ZN(n6074) );
  NAND3_X1 U12210 ( .A1(\SB2_2_30/i0_3 ), .A2(\SB2_2_30/i0_0 ), .A3(
        \SB2_2_30/i0[7] ), .ZN(\SB2_2_30/Component_Function_0/NAND4_in[3] ) );
  NAND3_X2 U12211 ( .A1(\SB1_1_15/i0_4 ), .A2(\SB1_1_15/i0_0 ), .A3(
        \SB1_1_15/i1_5 ), .ZN(\SB1_1_15/Component_Function_2/NAND4_in[3] ) );
  NAND4_X2 U12212 ( .A1(\SB3_12/Component_Function_3/NAND4_in[0] ), .A2(
        \SB3_12/Component_Function_3/NAND4_in[2] ), .A3(n6512), .A4(n3912), 
        .ZN(\SB3_12/buf_output[3] ) );
  XOR2_X1 U12213 ( .A1(\MC_ARK_ARC_1_1/temp5[9] ), .A2(n6076), .Z(
        \MC_ARK_ARC_1_1/buf_output[9] ) );
  XOR2_X1 U12214 ( .A1(n6077), .A2(n94), .Z(Ciphertext[130]) );
  NAND4_X2 U12215 ( .A1(\SB4_10/Component_Function_4/NAND4_in[0] ), .A2(
        \SB4_10/Component_Function_4/NAND4_in[2] ), .A3(
        \SB4_10/Component_Function_4/NAND4_in[3] ), .A4(
        \SB4_10/Component_Function_4/NAND4_in[1] ), .ZN(n6077) );
  INV_X2 U12216 ( .I(\SB1_0_13/buf_output[2] ), .ZN(\SB2_0_10/i1[9] ) );
  NAND4_X2 U12217 ( .A1(\SB1_0_13/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_13/Component_Function_2/NAND4_in[1] ), .A3(n4260), .A4(
        \SB1_0_13/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB1_0_13/buf_output[2] ) );
  XOR2_X1 U12218 ( .A1(n6078), .A2(n3097), .Z(\MC_ARK_ARC_1_2/buf_output[163] ) );
  XOR2_X1 U12219 ( .A1(\MC_ARK_ARC_1_2/temp1[163] ), .A2(
        \MC_ARK_ARC_1_2/temp4[163] ), .Z(n6078) );
  NAND4_X2 U12220 ( .A1(\SB3_12/Component_Function_4/NAND4_in[0] ), .A2(
        \SB3_12/Component_Function_4/NAND4_in[2] ), .A3(n2720), .A4(n6079), 
        .ZN(\SB3_12/buf_output[4] ) );
  NAND3_X1 U12221 ( .A1(\SB1_2_11/i0[8] ), .A2(\SB1_2_11/i1_5 ), .A3(
        \SB1_2_11/i3[0] ), .ZN(\SB1_2_11/Component_Function_3/NAND4_in[3] ) );
  NAND3_X2 U12222 ( .A1(\RI3[0][155] ), .A2(n2765), .A3(\SB2_0_6/i0[9] ), .ZN(
        n3729) );
  XOR2_X1 U12223 ( .A1(\RI5[0][54] ), .A2(\RI5[0][18] ), .Z(n6080) );
  XOR2_X1 U12224 ( .A1(\RI5[0][134] ), .A2(\RI5[0][170] ), .Z(
        \MC_ARK_ARC_1_0/temp3[68] ) );
  XOR2_X1 U12225 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[128] ), .A2(\RI5[2][164] ), .Z(\MC_ARK_ARC_1_2/temp3[62] ) );
  XOR2_X1 U12226 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[128] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[92] ), .Z(n1584) );
  XOR2_X1 U12227 ( .A1(\SB2_3_25/buf_output[3] ), .A2(\RI5[3][87] ), .Z(
        \MC_ARK_ARC_1_3/temp3[177] ) );
  NAND4_X2 U12228 ( .A1(\SB1_0_6/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_0_6/Component_Function_2/NAND4_in[2] ), .A3(n1279), .A4(
        \SB1_0_6/Component_Function_2/NAND4_in[0] ), .ZN(
        \SB1_0_6/buf_output[2] ) );
  XOR2_X1 U12229 ( .A1(n3023), .A2(\MC_ARK_ARC_1_2/temp6[93] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[93] ) );
  NAND4_X2 U12230 ( .A1(\SB2_1_15/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_1_15/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_15/Component_Function_4/NAND4_in[2] ), .A4(n6081), .ZN(
        \SB2_1_15/buf_output[4] ) );
  NAND3_X1 U12231 ( .A1(\SB2_2_8/i0[9] ), .A2(\SB2_2_8/i0[8] ), .A3(
        \SB2_2_8/i0_0 ), .ZN(\SB2_2_8/Component_Function_4/NAND4_in[0] ) );
  XOR2_X1 U12232 ( .A1(n6083), .A2(\MC_ARK_ARC_1_0/temp2[167] ), .Z(
        \MC_ARK_ARC_1_0/temp5[167] ) );
  XOR2_X1 U12233 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[167] ), .A2(\RI5[0][161] ), .Z(n6083) );
  NAND3_X1 U12234 ( .A1(\SB2_3_26/i1_7 ), .A2(\SB2_3_26/i1[9] ), .A3(
        \SB1_3_28/buf_output[3] ), .ZN(
        \SB2_3_26/Component_Function_3/NAND4_in[2] ) );
  NAND4_X2 U12235 ( .A1(\SB2_2_29/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_2_29/Component_Function_2/NAND4_in[0] ), .A3(n4501), .A4(n6084), 
        .ZN(\SB2_2_29/buf_output[2] ) );
  NAND2_X2 U12236 ( .A1(\SB2_1_3/i0_0 ), .A2(\SB2_1_3/i3[0] ), .ZN(n6085) );
  XOR2_X1 U12237 ( .A1(n6087), .A2(n6086), .Z(\MC_ARK_ARC_1_0/buf_output[117] ) );
  XOR2_X1 U12238 ( .A1(\MC_ARK_ARC_1_0/temp3[117] ), .A2(
        \MC_ARK_ARC_1_0/temp2[117] ), .Z(n6086) );
  XOR2_X1 U12239 ( .A1(n3944), .A2(\MC_ARK_ARC_1_0/temp4[117] ), .Z(n6087) );
  XOR2_X1 U12240 ( .A1(n6088), .A2(\MC_ARK_ARC_1_2/temp4[152] ), .Z(
        \MC_ARK_ARC_1_2/temp6[152] ) );
  NAND2_X2 U12241 ( .A1(\SB1_1_31/Component_Function_4/NAND4_in[2] ), .A2(
        \SB1_1_31/Component_Function_4/NAND4_in[3] ), .ZN(n6203) );
  NAND3_X1 U12242 ( .A1(\SB3_2/i0[8] ), .A2(\SB3_2/i1_5 ), .A3(\SB3_2/i3[0] ), 
        .ZN(n1777) );
  NAND3_X2 U12243 ( .A1(\SB3_16/i0[10] ), .A2(\SB3_16/i1[9] ), .A3(
        \SB3_16/i1_5 ), .ZN(n6089) );
  XOR2_X1 U12244 ( .A1(\SB2_0_12/buf_output[3] ), .A2(\SB2_0_16/buf_output[3] ), .Z(n6090) );
  XOR2_X1 U12245 ( .A1(n6092), .A2(\MC_ARK_ARC_1_3/temp4[118] ), .Z(
        \MC_ARK_ARC_1_3/temp6[118] ) );
  XOR2_X1 U12246 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[28] ), .A2(\RI5[3][184] ), 
        .Z(n6092) );
  NAND4_X2 U12247 ( .A1(n3184), .A2(\SB2_3_9/Component_Function_0/NAND4_in[1] ), .A3(\SB2_3_9/Component_Function_0/NAND4_in[0] ), .A4(n6093), .ZN(
        \SB2_3_9/buf_output[0] ) );
  NAND3_X2 U12248 ( .A1(\SB1_2_14/i0[10] ), .A2(\SB1_2_14/i0_3 ), .A3(
        \SB1_2_14/i0[9] ), .ZN(\SB1_2_14/Component_Function_4/NAND4_in[2] ) );
  XOR2_X1 U12249 ( .A1(n6094), .A2(n1334), .Z(\MC_ARK_ARC_1_2/temp6[21] ) );
  XOR2_X1 U12250 ( .A1(\RI5[2][123] ), .A2(\RI5[2][87] ), .Z(n6094) );
  XOR2_X1 U12251 ( .A1(\RI5[0][171] ), .A2(\RI5[0][15] ), .Z(n6095) );
  NAND3_X2 U12252 ( .A1(\SB4_18/i0[6] ), .A2(\SB4_18/i1_5 ), .A3(
        \SB4_18/i0[9] ), .ZN(n6096) );
  NAND4_X2 U12253 ( .A1(n6155), .A2(n947), .A3(
        \SB3_22/Component_Function_1/NAND4_in[2] ), .A4(
        \SB3_22/Component_Function_1/NAND4_in[0] ), .ZN(\SB3_22/buf_output[1] ) );
  XOR2_X1 U12254 ( .A1(\RI5[3][161] ), .A2(\RI5[3][125] ), .Z(n3331) );
  XOR2_X1 U12255 ( .A1(n3956), .A2(n3955), .Z(\MC_ARK_ARC_1_1/temp6[59] ) );
  XOR2_X1 U12256 ( .A1(\MC_ARK_ARC_1_3/temp5[59] ), .A2(
        \MC_ARK_ARC_1_3/temp6[59] ), .Z(\RI1[4][59] ) );
  XOR2_X1 U12257 ( .A1(n6241), .A2(n6240), .Z(\MC_ARK_ARC_1_0/buf_output[113] ) );
  XOR2_X1 U12258 ( .A1(\MC_ARK_ARC_1_1/temp1[50] ), .A2(n1551), .Z(n6097) );
  NAND3_X1 U12259 ( .A1(\SB4_19/i0_0 ), .A2(\SB4_19/i0[7] ), .A3(\SB4_19/i0_3 ), .ZN(n6098) );
  NAND3_X1 U12260 ( .A1(\SB2_0_7/i0_3 ), .A2(\SB2_0_7/i1[9] ), .A3(n2593), 
        .ZN(\SB2_0_7/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U12261 ( .A1(\MC_ARK_ARC_1_1/temp5[141] ), .A2(n6099), .Z(
        \MC_ARK_ARC_1_1/buf_output[141] ) );
  XOR2_X1 U12262 ( .A1(\MC_ARK_ARC_1_1/temp3[141] ), .A2(
        \MC_ARK_ARC_1_1/temp4[141] ), .Z(n6099) );
  NAND3_X2 U12263 ( .A1(\SB2_0_13/i0[10] ), .A2(\SB2_0_13/i0_3 ), .A3(
        \SB2_0_13/i0[6] ), .ZN(\SB2_0_13/Component_Function_2/NAND4_in[1] ) );
  XOR2_X1 U12264 ( .A1(n6101), .A2(n6100), .Z(\MC_ARK_ARC_1_2/buf_output[62] )
         );
  XOR2_X1 U12265 ( .A1(n2930), .A2(\MC_ARK_ARC_1_2/temp4[62] ), .Z(n6100) );
  XOR2_X1 U12266 ( .A1(n2931), .A2(\MC_ARK_ARC_1_2/temp3[62] ), .Z(n6101) );
  XOR2_X1 U12267 ( .A1(n6231), .A2(\MC_ARK_ARC_1_1/temp1[40] ), .Z(n6102) );
  XOR2_X1 U12268 ( .A1(n6103), .A2(n195), .Z(Ciphertext[121]) );
  NAND4_X2 U12269 ( .A1(\SB4_11/Component_Function_1/NAND4_in[3] ), .A2(n6118), 
        .A3(\SB4_11/Component_Function_1/NAND4_in[1] ), .A4(n3796), .ZN(n6103)
         );
  INV_X2 U12270 ( .I(\SB1_3_30/buf_output[2] ), .ZN(\SB2_3_27/i1[9] ) );
  NAND3_X2 U12271 ( .A1(\SB1_1_11/i0_0 ), .A2(\SB1_1_11/i0[7] ), .A3(
        \SB1_1_11/i0_3 ), .ZN(\SB1_1_11/Component_Function_0/NAND4_in[3] ) );
  XOR2_X1 U12272 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[44] ), .A2(\RI5[3][20] ), 
        .Z(n6105) );
  NAND4_X2 U12273 ( .A1(\SB2_3_7/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_3_7/Component_Function_3/NAND4_in[3] ), .A3(n4679), .A4(n6106), 
        .ZN(\SB2_3_7/buf_output[3] ) );
  INV_X2 U12274 ( .I(\SB1_1_5/buf_output[2] ), .ZN(\SB2_1_2/i1[9] ) );
  NAND4_X2 U12275 ( .A1(\SB1_1_5/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_1_5/Component_Function_2/NAND4_in[3] ), .A3(
        \SB1_1_5/Component_Function_2/NAND4_in[1] ), .A4(
        \SB1_1_5/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB1_1_5/buf_output[2] ) );
  XOR2_X1 U12276 ( .A1(\MC_ARK_ARC_1_3/temp2[116] ), .A2(n6109), .Z(
        \MC_ARK_ARC_1_3/temp5[116] ) );
  XOR2_X1 U12277 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[116] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[110] ), .Z(n6109) );
  NAND3_X2 U12278 ( .A1(\SB2_2_27/i0_3 ), .A2(\SB2_2_27/i0[6] ), .A3(
        \SB2_2_27/i1[9] ), .ZN(\SB2_2_27/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U12279 ( .A1(n2512), .A2(n6110), .Z(\MC_ARK_ARC_1_0/buf_output[159] ) );
  NAND3_X2 U12280 ( .A1(\SB3_11/i0[10] ), .A2(\SB3_11/i1[9] ), .A3(n582), .ZN(
        n6111) );
  NAND3_X1 U12281 ( .A1(\MC_ARK_ARC_1_2/buf_output[114] ), .A2(
        \MC_ARK_ARC_1_2/buf_output[115] ), .A3(
        \MC_ARK_ARC_1_2/buf_output[118] ), .ZN(n6533) );
  BUF_X2 U12282 ( .I(\SB2_0_7/i0[7] ), .Z(n6113) );
  NAND3_X1 U12283 ( .A1(\SB4_5/i0_3 ), .A2(\SB4_5/i0[9] ), .A3(\SB4_5/i0[8] ), 
        .ZN(n6114) );
  NAND4_X2 U12284 ( .A1(\SB1_0_28/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_28/Component_Function_2/NAND4_in[1] ), .A3(
        \SB1_0_28/Component_Function_2/NAND4_in[2] ), .A4(n6115), .ZN(
        \SB1_0_28/buf_output[2] ) );
  NAND3_X2 U12285 ( .A1(\SB1_0_28/i0_0 ), .A2(\SB1_0_28/i0_4 ), .A3(
        \SB1_0_28/i1_5 ), .ZN(n6115) );
  NAND3_X2 U12286 ( .A1(\SB2_3_17/i0[6] ), .A2(\SB2_3_17/i0_3 ), .A3(
        \SB2_3_17/i1[9] ), .ZN(\SB2_3_17/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U12287 ( .A1(n6117), .A2(n6116), .Z(n6327) );
  XOR2_X1 U12288 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[179] ), .A2(\RI5[1][83] ), 
        .Z(n6116) );
  XOR2_X1 U12289 ( .A1(\RI5[1][113] ), .A2(\RI5[1][23] ), .Z(n6117) );
  NAND4_X2 U12290 ( .A1(\SB1_0_12/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_0_12/Component_Function_5/NAND4_in[2] ), .A3(n2286), .A4(
        \SB1_0_12/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_0_12/buf_output[5] ) );
  NAND4_X2 U12291 ( .A1(\SB1_2_12/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_2_12/Component_Function_5/NAND4_in[2] ), .A3(n6371), .A4(
        \SB1_2_12/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_2_12/buf_output[5] ) );
  NAND3_X1 U12292 ( .A1(\SB4_11/i0[9] ), .A2(\SB4_11/i0[6] ), .A3(n3684), .ZN(
        n6118) );
  NAND3_X2 U12293 ( .A1(\SB3_0/i0[10] ), .A2(\SB3_0/i1[9] ), .A3(\SB3_0/i1_7 ), 
        .ZN(n3282) );
  XOR2_X1 U12294 ( .A1(n2435), .A2(n6119), .Z(\MC_ARK_ARC_1_0/buf_output[73] )
         );
  XOR2_X1 U12295 ( .A1(\MC_ARK_ARC_1_0/temp3[73] ), .A2(
        \MC_ARK_ARC_1_0/temp4[73] ), .Z(n6119) );
  NAND3_X2 U12296 ( .A1(\SB2_1_28/i0[6] ), .A2(\SB2_1_28/i0_3 ), .A3(
        \SB2_1_28/i1[9] ), .ZN(\SB2_1_28/Component_Function_3/NAND4_in[0] ) );
  NAND4_X2 U12297 ( .A1(\SB2_0_0/Component_Function_2/NAND4_in[1] ), .A2(
        \SB2_0_0/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_0_0/Component_Function_2/NAND4_in[0] ), .A4(
        \SB2_0_0/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB2_0_0/buf_output[2] ) );
  XOR2_X1 U12298 ( .A1(n3189), .A2(n6120), .Z(\MC_ARK_ARC_1_1/buf_output[77] )
         );
  XOR2_X1 U12299 ( .A1(\MC_ARK_ARC_1_1/temp3[77] ), .A2(n4118), .Z(n6120) );
  NAND3_X2 U12300 ( .A1(\SB2_2_27/i0[10] ), .A2(\SB2_2_27/i0_3 ), .A3(
        \SB2_2_27/i0[9] ), .ZN(n6121) );
  NAND3_X2 U12301 ( .A1(\SB1_1_28/i1[9] ), .A2(\SB1_1_28/i0_3 ), .A3(
        \SB1_1_28/i0_4 ), .ZN(\SB1_1_28/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U12302 ( .A1(\MC_ARK_ARC_1_2/temp3[160] ), .A2(
        \MC_ARK_ARC_1_2/temp4[160] ), .Z(\MC_ARK_ARC_1_2/temp6[160] ) );
  XOR2_X1 U12303 ( .A1(n6122), .A2(\MC_ARK_ARC_1_1/temp6[58] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[58] ) );
  XOR2_X1 U12304 ( .A1(\MC_ARK_ARC_1_1/temp2[58] ), .A2(
        \MC_ARK_ARC_1_1/temp1[58] ), .Z(n6122) );
  NAND3_X1 U12305 ( .A1(n3993), .A2(\SB2_3_11/i0_0 ), .A3(\SB2_3_11/i0_3 ), 
        .ZN(\SB2_3_11/Component_Function_0/NAND4_in[3] ) );
  XOR2_X1 U12306 ( .A1(n6123), .A2(n3939), .Z(\MC_ARK_ARC_1_2/buf_output[119] ) );
  XOR2_X1 U12307 ( .A1(n6206), .A2(\MC_ARK_ARC_1_2/temp1[119] ), .Z(n6123) );
  NAND3_X2 U12308 ( .A1(\SB1_2_29/i0[9] ), .A2(\SB1_2_29/i0[8] ), .A3(
        \SB1_2_29/i0_0 ), .ZN(n6124) );
  XOR2_X1 U12309 ( .A1(n6128), .A2(n6127), .Z(\MC_ARK_ARC_1_2/buf_output[133] ) );
  XOR2_X1 U12310 ( .A1(n6409), .A2(\MC_ARK_ARC_1_2/temp4[133] ), .Z(n6127) );
  XOR2_X1 U12311 ( .A1(\MC_ARK_ARC_1_3/temp5[185] ), .A2(n6129), .Z(
        \MC_ARK_ARC_1_3/buf_output[185] ) );
  XOR2_X1 U12312 ( .A1(n6132), .A2(n6131), .Z(\MC_ARK_ARC_1_3/temp5[119] ) );
  XOR2_X1 U12313 ( .A1(\RI5[3][113] ), .A2(\RI5[3][89] ), .Z(n6131) );
  NAND3_X1 U12314 ( .A1(\SB4_11/i0_0 ), .A2(\SB4_11/i1_7 ), .A3(\SB4_11/i3[0] ), .ZN(n4547) );
  XOR2_X1 U12315 ( .A1(n6133), .A2(n55), .Z(Ciphertext[125]) );
  NAND4_X2 U12316 ( .A1(n3127), .A2(\SB4_11/Component_Function_5/NAND4_in[1] ), 
        .A3(\SB4_11/Component_Function_5/NAND4_in[2] ), .A4(
        \SB4_11/Component_Function_5/NAND4_in[0] ), .ZN(n6133) );
  NAND4_X2 U12317 ( .A1(\SB3_14/Component_Function_4/NAND4_in[1] ), .A2(
        \SB3_14/Component_Function_4/NAND4_in[3] ), .A3(n4212), .A4(n6134), 
        .ZN(\SB3_14/buf_output[4] ) );
  NAND4_X2 U12318 ( .A1(\SB1_3_17/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_3_17/Component_Function_1/NAND4_in[2] ), .A3(n6417), .A4(n6135), 
        .ZN(\SB1_3_17/buf_output[1] ) );
  NAND4_X2 U12319 ( .A1(\SB1_0_8/Component_Function_3/NAND4_in[0] ), .A2(n2534), .A3(\SB1_0_8/Component_Function_3/NAND4_in[2] ), .A4(n1142), .ZN(
        \SB2_0_6/i0[10] ) );
  NAND4_X2 U12320 ( .A1(n3736), .A2(\SB2_0_0/Component_Function_4/NAND4_in[3] ), .A3(\SB2_0_0/Component_Function_4/NAND4_in[0] ), .A4(n6136), .ZN(
        \SB2_0_0/buf_output[4] ) );
  NAND3_X1 U12321 ( .A1(\SB2_0_0/i0_0 ), .A2(\SB2_0_0/i3[0] ), .A3(
        \SB2_0_0/i1_7 ), .ZN(n6136) );
  NAND4_X2 U12322 ( .A1(\SB2_2_10/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_2_10/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_2_10/Component_Function_4/NAND4_in[1] ), .A4(n6137), .ZN(
        \SB2_2_10/buf_output[4] ) );
  XOR2_X1 U12323 ( .A1(n6139), .A2(n6138), .Z(\MC_ARK_ARC_1_0/buf_output[127] ) );
  XOR2_X1 U12324 ( .A1(\MC_ARK_ARC_1_0/temp3[127] ), .A2(
        \MC_ARK_ARC_1_0/temp2[127] ), .Z(n6138) );
  XOR2_X1 U12325 ( .A1(\MC_ARK_ARC_1_0/temp1[127] ), .A2(
        \MC_ARK_ARC_1_0/temp4[127] ), .Z(n6139) );
  NAND3_X2 U12326 ( .A1(\SB2_2_2/i0_3 ), .A2(\SB2_2_2/i0[6] ), .A3(
        \SB2_2_2/i0[10] ), .ZN(n6150) );
  XOR2_X1 U12327 ( .A1(n6142), .A2(n6141), .Z(n6158) );
  XOR2_X1 U12328 ( .A1(\RI5[0][29] ), .A2(n210), .Z(n6141) );
  XOR2_X1 U12329 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[155] ), .A2(\RI5[0][185] ), .Z(n6142) );
  XOR2_X1 U12330 ( .A1(n6143), .A2(\MC_ARK_ARC_1_0/temp4[130] ), .Z(
        \MC_ARK_ARC_1_0/temp6[130] ) );
  XOR2_X1 U12331 ( .A1(\RI5[0][4] ), .A2(\RI5[0][40] ), .Z(n6143) );
  XOR2_X1 U12332 ( .A1(n6144), .A2(n194), .Z(Ciphertext[116]) );
  XOR2_X1 U12333 ( .A1(n6145), .A2(\MC_ARK_ARC_1_2/temp1[63] ), .Z(n2234) );
  XOR2_X1 U12334 ( .A1(\RI5[2][9] ), .A2(\RI5[2][33] ), .Z(n6145) );
  NAND4_X2 U12335 ( .A1(\SB1_3_30/Component_Function_3/NAND4_in[1] ), .A2(
        n4664), .A3(n6257), .A4(n6146), .ZN(\SB1_3_30/buf_output[3] ) );
  NAND3_X2 U12336 ( .A1(\SB1_3_30/i0[6] ), .A2(\SB1_3_30/i1[9] ), .A3(
        \SB1_3_30/i0_3 ), .ZN(n6146) );
  NAND4_X2 U12337 ( .A1(\SB2_0_2/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_0_2/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_0_2/Component_Function_4/NAND4_in[3] ), .A4(n6147), .ZN(
        \SB2_0_2/buf_output[4] ) );
  NAND3_X1 U12338 ( .A1(\SB2_0_2/i0[9] ), .A2(\SB2_0_2/i0_3 ), .A3(
        \SB2_0_2/i0[10] ), .ZN(n6147) );
  XOR2_X1 U12339 ( .A1(\RI5[0][184] ), .A2(\RI5[0][16] ), .Z(
        \MC_ARK_ARC_1_0/temp2[46] ) );
  NAND4_X2 U12340 ( .A1(\SB1_0_3/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_3/Component_Function_2/NAND4_in[3] ), .A3(
        \SB1_0_3/Component_Function_2/NAND4_in[2] ), .A4(n6148), .ZN(
        \RI3[0][188] ) );
  NAND3_X2 U12341 ( .A1(\SB1_0_3/i0[10] ), .A2(\SB1_0_3/i0_3 ), .A3(
        \SB1_0_3/i0[6] ), .ZN(n6148) );
  INV_X2 U12342 ( .I(\SB2_0_19/i0[10] ), .ZN(\SB2_0_19/i0[8] ) );
  NAND4_X2 U12343 ( .A1(n869), .A2(n719), .A3(
        \SB1_0_21/Component_Function_3/NAND4_in[3] ), .A4(n832), .ZN(
        \SB2_0_19/i0[10] ) );
  NAND3_X2 U12344 ( .A1(\SB3_9/i0[10] ), .A2(\SB3_9/i0[6] ), .A3(\SB3_9/i0_0 ), 
        .ZN(n6149) );
  NAND3_X1 U12345 ( .A1(\SB2_0_2/i0[6] ), .A2(\RI3[0][176] ), .A3(
        \SB2_0_2/i0[10] ), .ZN(\SB2_0_2/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U12346 ( .A1(\RI5[1][141] ), .A2(\RI5[1][135] ), .Z(
        \MC_ARK_ARC_1_1/temp1[141] ) );
  XOR2_X1 U12347 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[135] ), .A2(\RI5[3][99] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[33] ) );
  XOR2_X1 U12348 ( .A1(n2033), .A2(n3943), .Z(\MC_ARK_ARC_1_3/buf_output[43] )
         );
  XOR2_X1 U12349 ( .A1(\MC_ARK_ARC_1_1/temp2[149] ), .A2(n6151), .Z(n6162) );
  XOR2_X1 U12350 ( .A1(\RI5[1][23] ), .A2(\RI5[1][59] ), .Z(n6151) );
  NAND4_X2 U12351 ( .A1(\SB2_1_31/Component_Function_2/NAND4_in[0] ), .A2(n597), .A3(\SB2_1_31/Component_Function_2/NAND4_in[1] ), .A4(n6152), .ZN(
        \SB2_1_31/buf_output[2] ) );
  NAND3_X2 U12352 ( .A1(\SB2_1_31/i0_0 ), .A2(\SB2_1_31/i0_4 ), .A3(n5510), 
        .ZN(n6152) );
  NAND3_X1 U12353 ( .A1(\SB4_29/i0[10] ), .A2(\SB4_29/i1_7 ), .A3(
        \SB4_29/i1[9] ), .ZN(n3161) );
  XOR2_X1 U12354 ( .A1(n6154), .A2(n6153), .Z(\MC_ARK_ARC_1_3/buf_output[189] ) );
  XOR2_X1 U12355 ( .A1(n693), .A2(\MC_ARK_ARC_1_3/temp4[189] ), .Z(n6153) );
  XOR2_X1 U12356 ( .A1(n2780), .A2(n6197), .Z(n6154) );
  NAND3_X1 U12357 ( .A1(\SB3_22/i0_3 ), .A2(\SB3_22/i0[8] ), .A3(\SB3_22/i1_7 ), .ZN(n6155) );
  XOR2_X1 U12358 ( .A1(n6156), .A2(n221), .Z(Ciphertext[112]) );
  NAND4_X2 U12359 ( .A1(n2759), .A2(\SB4_13/Component_Function_4/NAND4_in[0] ), 
        .A3(n901), .A4(\SB4_13/Component_Function_4/NAND4_in[1] ), .ZN(n6156)
         );
  NAND4_X2 U12360 ( .A1(\SB1_3_23/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_3_23/Component_Function_2/NAND4_in[1] ), .A3(n2778), .A4(n2493), 
        .ZN(\SB2_3_20/i0_0 ) );
  NAND3_X2 U12361 ( .A1(\SB1_3_23/i0_3 ), .A2(\SB1_3_23/i0[9] ), .A3(
        \SB1_3_23/i0[8] ), .ZN(n2493) );
  NAND3_X2 U12362 ( .A1(\SB2_3_27/i0_4 ), .A2(\SB2_3_27/i0_0 ), .A3(
        \SB2_3_27/i1_5 ), .ZN(n4598) );
  NAND3_X1 U12363 ( .A1(\RI3[0][155] ), .A2(\SB2_0_6/i1[9] ), .A3(
        \SB2_0_6/i0[6] ), .ZN(\SB2_0_6/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U12364 ( .A1(\MC_ARK_ARC_1_0/temp3[157] ), .A2(n6159), .Z(n2499) );
  XOR2_X1 U12365 ( .A1(\SB2_0_10/buf_output[1] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[157] ), .Z(n6159) );
  NAND3_X2 U12366 ( .A1(\SB1_1_28/i0[6] ), .A2(\SB1_1_28/i0_4 ), .A3(
        \SB1_1_28/i0[9] ), .ZN(n3405) );
  XOR2_X1 U12367 ( .A1(n1392), .A2(\MC_ARK_ARC_1_3/buf_datainput[135] ), .Z(
        \MC_ARK_ARC_1_3/temp2[165] ) );
  NAND3_X1 U12368 ( .A1(\SB3_25/i1[9] ), .A2(\SB3_25/i0_3 ), .A3(
        \SB3_25/i0[6] ), .ZN(n6160) );
  NAND3_X2 U12369 ( .A1(\SB1_1_5/i0[6] ), .A2(\SB1_1_5/i0[10] ), .A3(
        \SB1_1_5/i0_0 ), .ZN(\SB1_1_5/Component_Function_5/NAND4_in[1] ) );
  XOR2_X1 U12370 ( .A1(n6162), .A2(n6161), .Z(\MC_ARK_ARC_1_1/buf_output[149] ) );
  XOR2_X1 U12371 ( .A1(\MC_ARK_ARC_1_1/temp1[149] ), .A2(
        \MC_ARK_ARC_1_1/temp4[149] ), .Z(n6161) );
  NAND4_X2 U12372 ( .A1(\SB1_3_26/Component_Function_0/NAND4_in[1] ), .A2(
        n2769), .A3(\SB1_3_26/Component_Function_0/NAND4_in[0] ), .A4(n6163), 
        .ZN(\SB1_3_26/buf_output[0] ) );
  XOR2_X1 U12373 ( .A1(\SB2_2_17/buf_output[1] ), .A2(\RI5[2][73] ), .Z(
        \MC_ARK_ARC_1_2/temp3[7] ) );
  NAND3_X1 U12374 ( .A1(n5511), .A2(\SB2_3_28/i0_3 ), .A3(n577), .ZN(
        \SB2_3_28/Component_Function_0/NAND4_in[2] ) );
  NAND4_X2 U12375 ( .A1(\SB1_2_7/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_2_7/Component_Function_1/NAND4_in[1] ), .A3(n1733), .A4(
        \SB1_2_7/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_2_7/buf_output[1] ) );
  XOR2_X1 U12376 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[76] ), .A2(\RI5[0][100] ), 
        .Z(\MC_ARK_ARC_1_0/temp2[130] ) );
  XOR2_X1 U12377 ( .A1(n3345), .A2(n6164), .Z(n894) );
  XOR2_X1 U12378 ( .A1(\SB2_2_10/buf_output[4] ), .A2(\RI5[2][112] ), .Z(n6164) );
  XOR2_X1 U12379 ( .A1(\MC_ARK_ARC_1_2/temp6[113] ), .A2(n3991), .Z(
        \MC_ARK_ARC_1_2/buf_output[113] ) );
  NAND3_X1 U12380 ( .A1(\SB1_1_23/i0_3 ), .A2(\SB1_1_23/i0_0 ), .A3(
        \SB1_1_23/i0[7] ), .ZN(n3124) );
  XOR2_X1 U12381 ( .A1(\MC_ARK_ARC_1_2/temp1[7] ), .A2(
        \MC_ARK_ARC_1_2/temp2[7] ), .Z(n1987) );
  NAND3_X1 U12382 ( .A1(\SB2_1_7/i0_4 ), .A2(\SB2_1_7/i1_7 ), .A3(
        \SB2_1_7/i0[8] ), .ZN(n1650) );
  INV_X2 U12383 ( .I(\SB1_3_20/buf_output[2] ), .ZN(\SB2_3_17/i1[9] ) );
  NAND4_X2 U12384 ( .A1(\SB1_3_20/Component_Function_2/NAND4_in[1] ), .A2(
        \SB1_3_20/Component_Function_2/NAND4_in[0] ), .A3(
        \SB1_3_20/Component_Function_2/NAND4_in[3] ), .A4(
        \SB1_3_20/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB1_3_20/buf_output[2] ) );
  NAND4_X2 U12385 ( .A1(\SB2_0_10/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_10/Component_Function_4/NAND4_in[3] ), .A3(
        \SB2_0_10/Component_Function_4/NAND4_in[1] ), .A4(n6165), .ZN(
        \SB2_0_10/buf_output[4] ) );
  INV_X2 U12386 ( .I(\SB1_3_14/buf_output[3] ), .ZN(n3651) );
  INV_X1 U12387 ( .I(\SB1_1_31/buf_output[1] ), .ZN(\SB2_1_27/i1_7 ) );
  NAND4_X2 U12388 ( .A1(\SB1_1_31/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_1_31/Component_Function_1/NAND4_in[2] ), .A3(n1710), .A4(
        \SB1_1_31/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_1_31/buf_output[1] ) );
  NAND3_X2 U12389 ( .A1(\SB3_29/i0[10] ), .A2(\SB3_29/i0_3 ), .A3(
        \SB3_29/i0[6] ), .ZN(n6172) );
  XOR2_X1 U12390 ( .A1(\MC_ARK_ARC_1_3/temp6[37] ), .A2(
        \MC_ARK_ARC_1_3/temp5[37] ), .Z(\MC_ARK_ARC_1_3/buf_output[37] ) );
  XOR2_X1 U12391 ( .A1(\MC_ARK_ARC_1_3/temp5[44] ), .A2(n1531), .Z(n3657) );
  NAND3_X2 U12392 ( .A1(\SB2_0_20/i0[9] ), .A2(\SB2_0_20/i0_3 ), .A3(
        \SB2_0_20/i0[10] ), .ZN(n6166) );
  XOR2_X1 U12393 ( .A1(\SB2_2_15/buf_output[0] ), .A2(\RI5[2][102] ), .Z(n3483) );
  NAND4_X2 U12394 ( .A1(\SB2_1_16/Component_Function_1/NAND4_in[0] ), .A2(
        \SB2_1_16/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_1_16/Component_Function_1/NAND4_in[1] ), .A4(n6167), .ZN(
        \SB2_1_16/buf_output[1] ) );
  NAND3_X1 U12395 ( .A1(\SB2_1_16/i0[8] ), .A2(\SB2_1_16/i1_7 ), .A3(
        \SB1_1_17/buf_output[4] ), .ZN(n6167) );
  NAND4_X2 U12396 ( .A1(n4561), .A2(n6168), .A3(n4250), .A4(
        \SB2_2_19/Component_Function_5/NAND4_in[3] ), .ZN(
        \SB2_2_19/buf_output[5] ) );
  NAND3_X2 U12397 ( .A1(\SB2_2_19/i0[6] ), .A2(\SB2_2_19/i0[10] ), .A3(
        \SB2_2_19/i0_0 ), .ZN(n6168) );
  XOR2_X1 U12398 ( .A1(\MC_ARK_ARC_1_2/temp2[92] ), .A2(n6169), .Z(
        \MC_ARK_ARC_1_2/temp5[92] ) );
  XOR2_X1 U12399 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[92] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[86] ), .Z(n6169) );
  NAND3_X2 U12400 ( .A1(\SB3_29/i0[10] ), .A2(\SB3_29/i0_0 ), .A3(
        \SB3_29/i0[6] ), .ZN(n6173) );
  AND2_X1 U12401 ( .A1(\SB2_2_9/Component_Function_1/NAND4_in[3] ), .A2(
        \SB2_2_9/Component_Function_1/NAND4_in[2] ), .Z(n6170) );
  NAND3_X2 U12402 ( .A1(n1388), .A2(\SB1_3_10/i0_0 ), .A3(\SB1_3_10/i0_4 ), 
        .ZN(n4264) );
  XOR2_X1 U12403 ( .A1(n6171), .A2(n93), .Z(Ciphertext[78]) );
  XOR2_X1 U12404 ( .A1(\MC_ARK_ARC_1_1/temp6[109] ), .A2(n6334), .Z(
        \MC_ARK_ARC_1_1/buf_output[109] ) );
  NAND4_X2 U12405 ( .A1(\SB3_29/Component_Function_2/NAND4_in[2] ), .A2(
        \SB3_29/Component_Function_2/NAND4_in[0] ), .A3(
        \SB3_29/Component_Function_2/NAND4_in[3] ), .A4(n6172), .ZN(
        \SB3_29/buf_output[2] ) );
  NAND4_X2 U12406 ( .A1(n6427), .A2(n4429), .A3(
        \SB2_2_6/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_2_6/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_2_6/buf_output[5] ) );
  XOR2_X1 U12407 ( .A1(n6175), .A2(n6176), .Z(\MC_ARK_ARC_1_2/buf_output[47] )
         );
  XOR2_X1 U12408 ( .A1(\MC_ARK_ARC_1_3/temp1[84] ), .A2(n6177), .Z(
        \MC_ARK_ARC_1_3/temp5[84] ) );
  XOR2_X1 U12409 ( .A1(\RI5[3][54] ), .A2(\RI5[3][30] ), .Z(n6177) );
  XOR2_X1 U12410 ( .A1(\RI5[0][182] ), .A2(\RI5[0][146] ), .Z(
        \MC_ARK_ARC_1_0/temp3[80] ) );
  XOR2_X1 U12411 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[128] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[122] ), .Z(\MC_ARK_ARC_1_2/temp1[128] )
         );
  NAND3_X1 U12412 ( .A1(\SB4_21/i0[6] ), .A2(\SB4_21/i0[7] ), .A3(
        \SB4_21/i0[8] ), .ZN(n6179) );
  XOR2_X1 U12413 ( .A1(\MC_ARK_ARC_1_3/temp3[36] ), .A2(
        \MC_ARK_ARC_1_3/temp4[36] ), .Z(\MC_ARK_ARC_1_3/temp6[36] ) );
  NAND3_X2 U12414 ( .A1(\SB3_27/i0_0 ), .A2(\SB3_27/i0[10] ), .A3(
        \SB3_27/i0[6] ), .ZN(n6180) );
  NAND3_X2 U12415 ( .A1(\SB2_3_31/i0_0 ), .A2(\SB2_3_31/i0[10] ), .A3(
        \SB2_3_31/i0[6] ), .ZN(n6518) );
  NAND4_X2 U12416 ( .A1(n3882), .A2(n1059), .A3(n3765), .A4(
        \SB2_3_7/Component_Function_2/NAND4_in[0] ), .ZN(
        \SB2_3_7/buf_output[2] ) );
  NAND3_X2 U12417 ( .A1(\SB2_3_7/i0_3 ), .A2(\SB2_3_7/i0[10] ), .A3(n1670), 
        .ZN(n1059) );
  XOR2_X1 U12418 ( .A1(\RI5[3][164] ), .A2(\RI5[3][158] ), .Z(
        \MC_ARK_ARC_1_3/temp1[164] ) );
  XOR2_X1 U12419 ( .A1(n6181), .A2(\MC_ARK_ARC_1_3/temp5[84] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[84] ) );
  XOR2_X1 U12420 ( .A1(\MC_ARK_ARC_1_3/temp3[84] ), .A2(
        \MC_ARK_ARC_1_3/temp4[84] ), .Z(n6181) );
  XOR2_X1 U12421 ( .A1(n6182), .A2(n146), .Z(Ciphertext[163]) );
  NAND4_X2 U12422 ( .A1(\SB4_4/Component_Function_1/NAND4_in[2] ), .A2(n1506), 
        .A3(\SB4_4/Component_Function_1/NAND4_in[1] ), .A4(
        \SB4_4/Component_Function_1/NAND4_in[0] ), .ZN(n6182) );
  XOR2_X1 U12423 ( .A1(n6183), .A2(n233), .Z(Ciphertext[63]) );
  XOR2_X1 U12424 ( .A1(\MC_ARK_ARC_1_3/temp1[101] ), .A2(n6184), .Z(
        \MC_ARK_ARC_1_3/temp5[101] ) );
  XOR2_X1 U12425 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[71] ), .A2(\RI5[3][47] ), 
        .Z(n6184) );
  NAND3_X1 U12426 ( .A1(\SB3_22/i0[9] ), .A2(\SB3_22/i0_3 ), .A3(
        \SB3_22/i0[10] ), .ZN(\SB3_22/Component_Function_4/NAND4_in[2] ) );
  XOR2_X1 U12427 ( .A1(n960), .A2(n6186), .Z(n4336) );
  XOR2_X1 U12428 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[41] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[17] ), .Z(n6186) );
  XOR2_X1 U12429 ( .A1(\MC_ARK_ARC_1_1/temp2[155] ), .A2(n6187), .Z(n3808) );
  XOR2_X1 U12430 ( .A1(\RI5[1][149] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[155] ), .Z(n6187) );
  NAND4_X2 U12431 ( .A1(\SB1_3_20/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_3_20/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_3_20/Component_Function_4/NAND4_in[3] ), .A4(n6188), .ZN(
        \SB1_3_20/buf_output[4] ) );
  NAND3_X1 U12432 ( .A1(\SB1_3_20/i0[9] ), .A2(\SB1_3_20/i0[10] ), .A3(
        \SB1_3_20/i0_3 ), .ZN(n6188) );
  XOR2_X1 U12433 ( .A1(\MC_ARK_ARC_1_0/temp2[43] ), .A2(n6189), .Z(n6193) );
  XOR2_X1 U12434 ( .A1(\RI5[0][37] ), .A2(\RI5[0][43] ), .Z(n6189) );
  XOR2_X1 U12435 ( .A1(\RI5[1][161] ), .A2(\RI5[1][167] ), .Z(n6190) );
  INV_X2 U12436 ( .I(\SB1_1_24/buf_output[3] ), .ZN(\SB2_1_22/i0[8] ) );
  NAND4_X2 U12437 ( .A1(n828), .A2(\SB1_3_20/Component_Function_1/NAND4_in[1] ), .A3(\SB1_3_20/Component_Function_1/NAND4_in[0] ), .A4(n6191), .ZN(
        \SB1_3_20/buf_output[1] ) );
  NAND3_X1 U12438 ( .A1(\SB1_3_20/i0[9] ), .A2(\SB1_3_20/i0[6] ), .A3(
        \SB1_3_20/i1_5 ), .ZN(n6191) );
  INV_X2 U12439 ( .I(\SB1_2_5/buf_output[2] ), .ZN(\SB2_2_2/i1[9] ) );
  NAND4_X2 U12440 ( .A1(\SB3_20/Component_Function_1/NAND4_in[2] ), .A2(
        \SB3_20/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_20/Component_Function_1/NAND4_in[3] ), .A4(
        \SB3_20/Component_Function_1/NAND4_in[0] ), .ZN(\SB3_20/buf_output[1] ) );
  XOR2_X1 U12441 ( .A1(\MC_ARK_ARC_1_1/temp3[132] ), .A2(n6192), .Z(n3764) );
  XOR2_X1 U12442 ( .A1(\RI5[1][78] ), .A2(\RI5[1][102] ), .Z(n6192) );
  XOR2_X1 U12443 ( .A1(n3177), .A2(\MC_ARK_ARC_1_3/temp2[63] ), .Z(n2820) );
  NAND3_X1 U12444 ( .A1(\SB1_1_21/i0_3 ), .A2(\SB1_1_21/i1[9] ), .A3(
        \MC_ARK_ARC_1_0/buf_output[64] ), .ZN(
        \SB1_1_21/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U12445 ( .A1(n2046), .A2(\MC_ARK_ARC_1_2/temp4[64] ), .Z(n3974) );
  NAND4_X2 U12446 ( .A1(\SB2_3_26/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_3_26/Component_Function_4/NAND4_in[0] ), .A3(n6416), .A4(
        \SB2_3_26/Component_Function_4/NAND4_in[3] ), .ZN(
        \SB2_3_26/buf_output[4] ) );
  NAND3_X2 U12447 ( .A1(\SB3_18/i0[9] ), .A2(\SB3_18/i0[6] ), .A3(
        \SB3_18/i0_4 ), .ZN(n6426) );
  XOR2_X1 U12448 ( .A1(\RI5[1][86] ), .A2(\RI5[1][122] ), .Z(
        \MC_ARK_ARC_1_1/temp3[20] ) );
  XOR2_X1 U12449 ( .A1(n6193), .A2(\MC_ARK_ARC_1_0/temp6[43] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[43] ) );
  NAND4_X2 U12450 ( .A1(\SB2_3_24/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_3_24/Component_Function_5/NAND4_in[3] ), .A3(n6218), .A4(
        \SB2_3_24/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_3_24/buf_output[5] ) );
  NAND4_X2 U12451 ( .A1(n6349), .A2(
        \SB1_1_14/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_1_14/Component_Function_5/NAND4_in[2] ), .A4(
        \SB1_1_14/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_1_14/buf_output[5] ) );
  INV_X4 U12452 ( .I(n6194), .ZN(\SB1_1_7/buf_output[2] ) );
  XOR2_X1 U12453 ( .A1(\MC_ARK_ARC_1_3/temp1[94] ), .A2(n4059), .Z(n4184) );
  XOR2_X1 U12454 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[9] ), .A2(\RI5[1][15] ), 
        .Z(n4177) );
  NAND4_X2 U12455 ( .A1(\SB1_0_6/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_0_6/Component_Function_3/NAND4_in[2] ), .A3(n1917), .A4(n1916), 
        .ZN(\RI3[0][165] ) );
  XOR2_X1 U12456 ( .A1(\MC_ARK_ARC_1_1/temp1[78] ), .A2(
        \MC_ARK_ARC_1_1/temp2[78] ), .Z(\MC_ARK_ARC_1_1/temp5[78] ) );
  XOR2_X1 U12457 ( .A1(\RI5[3][83] ), .A2(\RI5[3][59] ), .Z(
        \MC_ARK_ARC_1_3/temp2[113] ) );
  XOR2_X1 U12458 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[167] ), .A2(\RI5[0][101] ), .Z(n2989) );
  NAND4_X2 U12459 ( .A1(\SB3_20/Component_Function_4/NAND4_in[1] ), .A2(
        \SB3_20/Component_Function_4/NAND4_in[2] ), .A3(n3748), .A4(
        \SB3_20/Component_Function_4/NAND4_in[0] ), .ZN(\SB3_20/buf_output[4] ) );
  XOR2_X1 U12460 ( .A1(\MC_ARK_ARC_1_3/temp6[113] ), .A2(n1699), .Z(n2291) );
  NAND3_X2 U12461 ( .A1(\SB1_3_2/i0[10] ), .A2(\SB1_3_2/i1[9] ), .A3(
        \SB1_3_2/i1_7 ), .ZN(n4563) );
  NAND4_X2 U12462 ( .A1(\SB2_3_23/Component_Function_3/NAND4_in[1] ), .A2(
        \SB2_3_23/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_3_23/Component_Function_3/NAND4_in[2] ), .A4(
        \SB2_3_23/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB2_3_23/buf_output[3] ) );
  XOR2_X1 U12463 ( .A1(\MC_ARK_ARC_1_0/temp6[65] ), .A2(n3727), .Z(
        \MC_ARK_ARC_1_0/buf_output[65] ) );
  NAND4_X2 U12464 ( .A1(\SB3_20/Component_Function_2/NAND4_in[3] ), .A2(
        \SB3_20/Component_Function_2/NAND4_in[0] ), .A3(n3106), .A4(n3830), 
        .ZN(\SB3_20/buf_output[2] ) );
  NAND4_X2 U12465 ( .A1(\SB2_1_21/Component_Function_2/NAND4_in[0] ), .A2(
        n6283), .A3(\SB2_1_21/Component_Function_2/NAND4_in[2] ), .A4(n711), 
        .ZN(\SB2_1_21/buf_output[2] ) );
  NAND3_X1 U12466 ( .A1(\SB1_0_11/i0[10] ), .A2(\SB1_0_11/i1_7 ), .A3(
        \SB1_0_11/i1[9] ), .ZN(n6196) );
  XOR2_X1 U12467 ( .A1(\RI5[3][63] ), .A2(\RI5[3][99] ), .Z(n6197) );
  NAND3_X1 U12468 ( .A1(\SB4_24/i0_0 ), .A2(\SB4_24/i3[0] ), .A3(\SB4_24/i1_7 ), .ZN(n6198) );
  NAND4_X2 U12469 ( .A1(n4720), .A2(
        \SB2_1_10/Component_Function_5/NAND4_in[3] ), .A3(n977), .A4(n6199), 
        .ZN(\SB2_1_10/buf_output[5] ) );
  NAND2_X1 U12470 ( .A1(\SB2_1_10/i0_0 ), .A2(n6200), .ZN(n6199) );
  INV_X1 U12471 ( .I(n6201), .ZN(n6200) );
  NAND2_X1 U12472 ( .A1(\SB1_1_12/buf_output[3] ), .A2(
        \SB1_1_14/buf_output[1] ), .ZN(n6201) );
  XOR2_X1 U12473 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[165] ), .A2(\RI5[0][171] ), .Z(n6364) );
  NOR2_X2 U12474 ( .A1(n2556), .A2(n6203), .ZN(n2828) );
  XOR2_X1 U12475 ( .A1(n6204), .A2(\MC_ARK_ARC_1_2/temp6[28] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[28] ) );
  XOR2_X1 U12476 ( .A1(\MC_ARK_ARC_1_2/temp2[28] ), .A2(
        \MC_ARK_ARC_1_2/temp1[28] ), .Z(n6204) );
  NAND3_X2 U12477 ( .A1(\SB1_1_31/i0[8] ), .A2(\SB1_1_31/i0[9] ), .A3(
        \SB1_1_31/i0_3 ), .ZN(n6205) );
  XOR2_X1 U12478 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[65] ), .A2(\RI5[2][89] ), 
        .Z(n6206) );
  NAND3_X1 U12479 ( .A1(\SB3_15/i0[6] ), .A2(\SB3_15/i0[9] ), .A3(
        \SB3_15/i1_5 ), .ZN(\SB3_15/Component_Function_1/NAND4_in[2] ) );
  XOR2_X1 U12480 ( .A1(\MC_ARK_ARC_1_1/temp6[65] ), .A2(n2807), .Z(n3681) );
  XOR2_X1 U12481 ( .A1(\MC_ARK_ARC_1_1/temp3[65] ), .A2(
        \MC_ARK_ARC_1_1/temp4[65] ), .Z(\MC_ARK_ARC_1_1/temp6[65] ) );
  INV_X2 U12482 ( .I(\SB1_3_9/buf_output[3] ), .ZN(\SB2_3_7/i0[8] ) );
  XOR2_X1 U12483 ( .A1(n4463), .A2(n6207), .Z(n3049) );
  XOR2_X1 U12484 ( .A1(\RI5[0][101] ), .A2(\RI5[0][95] ), .Z(n6207) );
  XOR2_X1 U12485 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[174] ), .A2(\RI5[3][18] ), 
        .Z(\MC_ARK_ARC_1_3/temp3[108] ) );
  XOR2_X1 U12486 ( .A1(n6208), .A2(\MC_ARK_ARC_1_0/temp1[189] ), .Z(n1303) );
  XOR2_X1 U12487 ( .A1(\RI5[0][159] ), .A2(\RI5[0][135] ), .Z(n6208) );
  XOR2_X1 U12488 ( .A1(n6209), .A2(n81), .Z(Ciphertext[18]) );
  NAND4_X2 U12489 ( .A1(n1918), .A2(n6485), .A3(n1703), .A4(
        \SB4_28/Component_Function_0/NAND4_in[0] ), .ZN(n6209) );
  XOR2_X1 U12490 ( .A1(\RI5[3][63] ), .A2(\RI5[3][93] ), .Z(n4054) );
  XOR2_X1 U12491 ( .A1(\MC_ARK_ARC_1_0/temp5[147] ), .A2(
        \MC_ARK_ARC_1_0/temp6[147] ), .Z(\MC_ARK_ARC_1_0/buf_output[147] ) );
  NAND3_X2 U12492 ( .A1(\SB1_3_0/i0_0 ), .A2(\SB1_3_0/i0[10] ), .A3(
        \SB1_3_0/i0[6] ), .ZN(n6210) );
  XOR2_X1 U12493 ( .A1(\RI5[2][134] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[158] ), .Z(n6211) );
  NAND3_X1 U12494 ( .A1(\SB3_12/i0[9] ), .A2(\SB3_12/i0[6] ), .A3(
        \SB3_12/i1_5 ), .ZN(n6213) );
  NAND4_X2 U12495 ( .A1(n3011), .A2(n2749), .A3(
        \SB1_3_26/Component_Function_1/NAND4_in[1] ), .A4(
        \SB1_3_26/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_3_26/buf_output[1] ) );
  NAND3_X2 U12496 ( .A1(\SB2_3_0/i0[10] ), .A2(\SB2_3_0/i1[9] ), .A3(
        \SB2_3_0/i1_5 ), .ZN(n6214) );
  NAND3_X2 U12497 ( .A1(\SB2_3_24/i0_0 ), .A2(\SB1_3_26/buf_output[3] ), .A3(
        \SB2_3_24/i0[6] ), .ZN(n6218) );
  NAND3_X2 U12498 ( .A1(\SB2_1_19/i0[10] ), .A2(n1396), .A3(\SB2_1_19/i1_5 ), 
        .ZN(n4381) );
  XOR2_X1 U12499 ( .A1(n1960), .A2(n6219), .Z(n1909) );
  INV_X1 U12500 ( .I(\SB1_2_10/buf_output[5] ), .ZN(\SB2_2_10/i1_5 ) );
  NAND4_X2 U12501 ( .A1(n3591), .A2(
        \SB1_2_10/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_2_10/Component_Function_5/NAND4_in[1] ), .A4(n3348), .ZN(
        \SB1_2_10/buf_output[5] ) );
  XOR2_X1 U12502 ( .A1(n6221), .A2(n6220), .Z(\MC_ARK_ARC_1_1/temp6[152] ) );
  XOR2_X1 U12503 ( .A1(\RI5[1][62] ), .A2(n55), .Z(n6220) );
  XOR2_X1 U12504 ( .A1(\RI5[1][188] ), .A2(\RI5[1][26] ), .Z(n6221) );
  XOR2_X1 U12505 ( .A1(\RI5[2][16] ), .A2(\RI5[2][52] ), .Z(
        \MC_ARK_ARC_1_2/temp3[142] ) );
  NAND4_X2 U12506 ( .A1(n611), .A2(\SB1_2_10/Component_Function_2/NAND4_in[1] ), .A3(\SB1_2_10/Component_Function_2/NAND4_in[2] ), .A4(n6222), .ZN(
        \SB1_2_10/buf_output[2] ) );
  NAND3_X2 U12507 ( .A1(\SB1_2_10/i0[10] ), .A2(\SB1_2_10/i1_5 ), .A3(
        \SB1_2_10/i1[9] ), .ZN(n6222) );
  NAND4_X2 U12508 ( .A1(n4710), .A2(\SB1_2_9/Component_Function_1/NAND4_in[1] ), .A3(\SB1_2_9/Component_Function_1/NAND4_in[0] ), .A4(n6223), .ZN(
        \SB1_2_9/buf_output[1] ) );
  NAND3_X1 U12509 ( .A1(\SB2_2_30/i0_3 ), .A2(\SB2_2_30/i0[10] ), .A3(
        \SB2_2_30/i0[9] ), .ZN(n1694) );
  NAND4_X2 U12510 ( .A1(\SB2_0_5/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_5/Component_Function_4/NAND4_in[2] ), .A3(
        \SB2_0_5/Component_Function_4/NAND4_in[1] ), .A4(n6224), .ZN(
        \SB2_0_5/buf_output[4] ) );
  XOR2_X1 U12511 ( .A1(n6226), .A2(n184), .Z(Ciphertext[88]) );
  NAND4_X2 U12512 ( .A1(\SB2_0_3/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_3/Component_Function_2/NAND4_in[1] ), .A3(
        \SB2_0_3/Component_Function_2/NAND4_in[2] ), .A4(n3016), .ZN(
        \SB2_0_3/buf_output[2] ) );
  NAND4_X2 U12513 ( .A1(\SB2_3_12/Component_Function_2/NAND4_in[2] ), .A2(
        \SB2_3_12/Component_Function_2/NAND4_in[0] ), .A3(n6536), .A4(n4113), 
        .ZN(\SB2_3_12/buf_output[2] ) );
  NAND3_X1 U12514 ( .A1(\SB3_14/i0[10] ), .A2(\SB3_14/i0_0 ), .A3(
        \SB3_14/i0[6] ), .ZN(\SB3_14/Component_Function_5/NAND4_in[1] ) );
  NAND3_X1 U12515 ( .A1(\SB2_2_10/i0_3 ), .A2(\SB2_2_10/i0[6] ), .A3(
        \SB2_2_10/i1[9] ), .ZN(\SB2_2_10/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U12516 ( .A1(\SB2_1_20/i0_0 ), .A2(\SB2_1_20/i0[9] ), .A3(
        \SB2_1_20/i0[8] ), .ZN(\SB2_1_20/Component_Function_4/NAND4_in[0] ) );
  NAND4_X2 U12517 ( .A1(\SB4_14/Component_Function_1/NAND4_in[1] ), .A2(
        \SB4_14/Component_Function_1/NAND4_in[2] ), .A3(
        \SB4_14/Component_Function_1/NAND4_in[0] ), .A4(
        \SB4_14/Component_Function_1/NAND4_in[3] ), .ZN(n6388) );
  XOR2_X1 U12518 ( .A1(n6266), .A2(\MC_ARK_ARC_1_0/temp1[52] ), .Z(n3215) );
  NAND3_X1 U12519 ( .A1(\SB2_0_3/i0_0 ), .A2(\SB2_0_3/i3[0] ), .A3(
        \SB2_0_3/i1_7 ), .ZN(\SB2_0_3/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U12520 ( .A1(n3356), .A2(n6534), .Z(n4461) );
  XOR2_X1 U12521 ( .A1(\MC_ARK_ARC_1_1/temp5[86] ), .A2(n1146), .Z(
        \MC_ARK_ARC_1_1/buf_output[86] ) );
  XOR2_X1 U12522 ( .A1(\MC_ARK_ARC_1_0/temp3[152] ), .A2(
        \MC_ARK_ARC_1_0/temp4[152] ), .Z(\MC_ARK_ARC_1_0/temp6[152] ) );
  NAND3_X2 U12523 ( .A1(\SB2_2_30/i0_3 ), .A2(\SB2_2_30/i0[10] ), .A3(
        \SB2_2_30/i0[6] ), .ZN(n4556) );
  XOR2_X1 U12524 ( .A1(\SB2_2_26/buf_output[2] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[86] ), .Z(\MC_ARK_ARC_1_2/temp3[176] )
         );
  NAND3_X1 U12525 ( .A1(\SB3_8/i0[10] ), .A2(\SB3_8/i1[9] ), .A3(\SB3_8/i1_7 ), 
        .ZN(\SB3_8/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U12526 ( .A1(\SB2_1_14/i0_3 ), .A2(\SB2_1_14/i0[10] ), .A3(
        \SB2_1_14/i0[6] ), .ZN(n4201) );
  NAND4_X2 U12527 ( .A1(\SB1_2_3/Component_Function_2/NAND4_in[1] ), .A2(n4252), .A3(\SB1_2_3/Component_Function_2/NAND4_in[3] ), .A4(n6227), .ZN(
        \SB1_2_3/buf_output[2] ) );
  NAND3_X2 U12528 ( .A1(\SB1_2_3/i0[10] ), .A2(\SB1_2_3/i1[9] ), .A3(
        \SB1_2_3/i1_5 ), .ZN(n6227) );
  NAND3_X1 U12529 ( .A1(\SB1_3_5/i0[6] ), .A2(\SB1_3_5/i0[10] ), .A3(
        \SB1_3_5/i0_3 ), .ZN(n6228) );
  XOR2_X1 U12530 ( .A1(n6229), .A2(\MC_ARK_ARC_1_3/temp1[41] ), .Z(
        \MC_ARK_ARC_1_3/temp5[41] ) );
  XOR2_X1 U12531 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[179] ), .A2(\RI5[3][11] ), 
        .Z(n6229) );
  XOR2_X1 U12532 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[135] ), .A2(\RI5[3][171] ), .Z(\MC_ARK_ARC_1_3/temp3[69] ) );
  BUF_X2 U12533 ( .I(\SB2_2_4/i0[7] ), .Z(n6230) );
  INV_X1 U12534 ( .I(\SB1_3_17/buf_output[1] ), .ZN(\SB2_3_13/i1_7 ) );
  XOR2_X1 U12535 ( .A1(\RI5[1][114] ), .A2(\RI5[1][90] ), .Z(n6234) );
  XOR2_X1 U12536 ( .A1(\MC_ARK_ARC_1_2/temp5[5] ), .A2(n6235), .Z(\RI1[3][5] )
         );
  XOR2_X1 U12537 ( .A1(\MC_ARK_ARC_1_2/temp3[5] ), .A2(
        \MC_ARK_ARC_1_2/temp4[5] ), .Z(n6235) );
  XOR2_X1 U12538 ( .A1(\MC_ARK_ARC_1_3/temp5[183] ), .A2(n6236), .Z(
        \MC_ARK_ARC_1_3/buf_output[183] ) );
  XOR2_X1 U12539 ( .A1(n6237), .A2(n6238), .Z(\MC_ARK_ARC_1_1/buf_output[23] )
         );
  XOR2_X1 U12540 ( .A1(n1063), .A2(n4268), .Z(n6237) );
  NAND4_X2 U12541 ( .A1(\SB2_1_14/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_1_14/Component_Function_5/NAND4_in[1] ), .A3(n2834), .A4(
        \SB2_1_14/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_1_14/buf_output[5] ) );
  NAND3_X2 U12542 ( .A1(\SB2_0_22/i0_3 ), .A2(\SB2_0_22/i0_4 ), .A3(
        \SB2_0_22/i1[9] ), .ZN(n2218) );
  XOR2_X1 U12543 ( .A1(\MC_ARK_ARC_1_0/temp1[83] ), .A2(n6239), .Z(
        \MC_ARK_ARC_1_0/temp5[83] ) );
  XOR2_X1 U12544 ( .A1(\RI5[0][53] ), .A2(\RI5[0][29] ), .Z(n6239) );
  NAND3_X1 U12545 ( .A1(\SB1_1_17/i0_3 ), .A2(\SB1_1_17/i0_0 ), .A3(
        \SB1_1_17/i0_4 ), .ZN(\SB1_1_17/Component_Function_3/NAND4_in[1] ) );
  XOR2_X1 U12546 ( .A1(n1095), .A2(\MC_ARK_ARC_1_0/temp2[113] ), .Z(n6241) );
  XOR2_X1 U12547 ( .A1(n6242), .A2(\MC_ARK_ARC_1_2/temp4[73] ), .Z(n3865) );
  XOR2_X1 U12548 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[175] ), .A2(\RI5[2][139] ), .Z(n6242) );
  XOR2_X1 U12549 ( .A1(n6243), .A2(n163), .Z(Ciphertext[165]) );
  XOR2_X1 U12550 ( .A1(\RI5[3][141] ), .A2(\RI5[3][147] ), .Z(n2240) );
  NAND4_X2 U12551 ( .A1(\SB2_1_3/Component_Function_2/NAND4_in[0] ), .A2(n1852), .A3(\SB2_1_3/Component_Function_2/NAND4_in[2] ), .A4(
        \SB2_1_3/Component_Function_2/NAND4_in[1] ), .ZN(
        \SB2_1_3/buf_output[2] ) );
  XOR2_X1 U12552 ( .A1(n2094), .A2(n6245), .Z(\MC_ARK_ARC_1_0/buf_output[86] )
         );
  XOR2_X1 U12553 ( .A1(n4523), .A2(\MC_ARK_ARC_1_0/temp4[86] ), .Z(n6245) );
  NAND3_X2 U12554 ( .A1(\SB3_16/i0_0 ), .A2(\SB3_16/i1_5 ), .A3(\SB3_16/i0_4 ), 
        .ZN(n6246) );
  INV_X1 U12555 ( .I(\SB1_2_13/buf_output[1] ), .ZN(\SB2_2_9/i1_7 ) );
  NAND4_X2 U12556 ( .A1(\SB1_2_13/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_2_13/Component_Function_1/NAND4_in[0] ), .A3(
        \SB1_2_13/Component_Function_1/NAND4_in[2] ), .A4(
        \SB1_2_13/Component_Function_1/NAND4_in[3] ), .ZN(
        \SB1_2_13/buf_output[1] ) );
  NAND3_X2 U12557 ( .A1(\SB2_0_12/i0[10] ), .A2(\SB2_0_12/i0[6] ), .A3(
        \SB2_0_12/i0_3 ), .ZN(\SB2_0_12/Component_Function_2/NAND4_in[1] ) );
  XOR2_X1 U12558 ( .A1(\RI5[3][39] ), .A2(\RI5[3][63] ), .Z(n3780) );
  NAND4_X2 U12559 ( .A1(\SB3_27/Component_Function_3/NAND4_in[2] ), .A2(n6412), 
        .A3(n1640), .A4(\SB3_27/Component_Function_3/NAND4_in[1] ), .ZN(
        \SB3_27/buf_output[3] ) );
  NAND4_X2 U12560 ( .A1(\SB2_2_30/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_2_30/Component_Function_1/NAND4_in[2] ), .A3(
        \SB2_2_30/Component_Function_1/NAND4_in[0] ), .A4(n6247), .ZN(
        \SB2_2_30/buf_output[1] ) );
  NAND3_X1 U12561 ( .A1(n2343), .A2(\SB2_2_30/i1_7 ), .A3(\SB2_2_30/i0[8] ), 
        .ZN(n6247) );
  NAND3_X2 U12562 ( .A1(\SB2_1_17/i0_3 ), .A2(\SB2_1_17/i0[6] ), .A3(
        \SB2_1_17/i1[9] ), .ZN(\SB2_1_17/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U12563 ( .A1(\MC_ARK_ARC_1_2/temp4[157] ), .A2(n6248), .Z(n683) );
  XOR2_X1 U12564 ( .A1(\RI5[2][31] ), .A2(\RI5[2][67] ), .Z(n6248) );
  NAND3_X2 U12565 ( .A1(\SB1_0_28/i0_3 ), .A2(\SB1_0_28/i0_4 ), .A3(
        \SB1_0_28/i1[9] ), .ZN(n6249) );
  NAND3_X2 U12566 ( .A1(\SB2_1_3/i0_3 ), .A2(\SB2_1_3/i1[9] ), .A3(n5208), 
        .ZN(\SB2_1_3/Component_Function_5/NAND4_in[2] ) );
  NAND4_X2 U12567 ( .A1(n1866), .A2(
        \SB2_2_15/Component_Function_5/NAND4_in[3] ), .A3(n6250), .A4(
        \SB2_2_15/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_2_15/buf_output[5] ) );
  NAND3_X2 U12568 ( .A1(\SB2_2_15/i0[6] ), .A2(\SB2_2_15/i0_0 ), .A3(
        \SB2_2_15/i0[10] ), .ZN(n6250) );
  NAND4_X2 U12569 ( .A1(\SB1_1_30/Component_Function_0/NAND4_in[1] ), .A2(
        \SB1_1_30/Component_Function_0/NAND4_in[2] ), .A3(
        \SB1_1_30/Component_Function_0/NAND4_in[0] ), .A4(n6251), .ZN(
        \SB1_1_30/buf_output[0] ) );
  XOR2_X1 U12570 ( .A1(n6253), .A2(n3126), .Z(\MC_ARK_ARC_1_0/temp5[56] ) );
  XOR2_X1 U12571 ( .A1(\SB2_0_2/buf_output[2] ), .A2(\RI5[0][26] ), .Z(n6253)
         );
  NAND2_X1 U12572 ( .A1(\SB3_13/i3[0] ), .A2(\MC_ARK_ARC_1_3/buf_output[110] ), 
        .ZN(n6254) );
  NAND3_X1 U12573 ( .A1(\SB2_2_18/i0_3 ), .A2(\SB2_2_18/i0_0 ), .A3(
        \SB2_2_18/i0[7] ), .ZN(\SB2_2_18/Component_Function_0/NAND4_in[3] ) );
  NAND2_X2 U12574 ( .A1(\SB1_2_29/i1_5 ), .A2(n1721), .ZN(n6255) );
  NAND3_X1 U12575 ( .A1(\SB1_3_6/i0_3 ), .A2(\MC_ARK_ARC_1_2/buf_output[150] ), 
        .A3(\SB1_3_6/i0[8] ), .ZN(\SB1_3_6/Component_Function_2/NAND4_in[2] )
         );
  NAND4_X2 U12576 ( .A1(\SB2_2_26/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_26/Component_Function_5/NAND4_in[1] ), .A3(n6448), .A4(
        \SB2_2_26/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_2_26/buf_output[5] ) );
  XOR2_X1 U12577 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[39] ), .A2(\RI5[2][63] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[93] ) );
  NAND3_X2 U12578 ( .A1(\SB2_2_5/i3[0] ), .A2(\SB2_2_5/i1_5 ), .A3(
        \SB2_2_5/i0[8] ), .ZN(\SB2_2_5/Component_Function_3/NAND4_in[3] ) );
  NAND4_X2 U12579 ( .A1(\SB2_0_29/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_29/Component_Function_2/NAND4_in[3] ), .A3(n3141), .A4(n1903), 
        .ZN(\SB2_0_29/buf_output[2] ) );
  XOR2_X1 U12580 ( .A1(\RI5[2][57] ), .A2(\RI5[2][93] ), .Z(
        \MC_ARK_ARC_1_2/temp3[183] ) );
  NAND3_X2 U12581 ( .A1(\SB2_1_12/i0_3 ), .A2(\SB2_1_12/i0_4 ), .A3(
        \SB2_1_12/i1[9] ), .ZN(\SB2_1_12/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U12582 ( .A1(\MC_ARK_ARC_1_2/temp4[23] ), .A2(
        \MC_ARK_ARC_1_2/temp3[23] ), .Z(n1665) );
  NAND4_X2 U12583 ( .A1(n2985), .A2(
        \SB2_2_27/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_2_27/Component_Function_3/NAND4_in[3] ), .A4(n3947), .ZN(
        \SB2_2_27/buf_output[3] ) );
  NAND3_X2 U12584 ( .A1(\SB2_3_28/i0[9] ), .A2(\SB2_3_28/i0_3 ), .A3(
        \SB2_3_28/i0[8] ), .ZN(n6509) );
  NAND4_X2 U12585 ( .A1(\SB2_2_24/Component_Function_3/NAND4_in[3] ), .A2(
        \SB2_2_24/Component_Function_3/NAND4_in[0] ), .A3(n3032), .A4(n4408), 
        .ZN(\SB2_2_24/buf_output[3] ) );
  XOR2_X1 U12586 ( .A1(\MC_ARK_ARC_1_1/temp2[165] ), .A2(
        \MC_ARK_ARC_1_1/temp1[165] ), .Z(n6496) );
  NAND3_X1 U12587 ( .A1(\SB3_6/i0[9] ), .A2(\RI1[4][155] ), .A3(\SB3_6/i0[10] ), .ZN(n2762) );
  NAND4_X2 U12588 ( .A1(\SB2_2_0/Component_Function_3/NAND4_in[3] ), .A2(n1773), .A3(\SB2_2_0/Component_Function_3/NAND4_in[1] ), .A4(n2553), .ZN(
        \SB2_2_0/buf_output[3] ) );
  NAND4_X2 U12589 ( .A1(\SB1_1_11/Component_Function_5/NAND4_in[1] ), .A2(
        \SB1_1_11/Component_Function_5/NAND4_in[2] ), .A3(
        \SB1_1_11/Component_Function_5/NAND4_in[0] ), .A4(n2624), .ZN(
        \SB1_1_11/buf_output[5] ) );
  XOR2_X1 U12590 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[38] ), .A2(\RI5[1][32] ), 
        .Z(\MC_ARK_ARC_1_1/temp1[38] ) );
  NAND3_X2 U12591 ( .A1(\SB2_1_16/i0_4 ), .A2(\SB2_1_16/i1[9] ), .A3(
        \SB2_1_16/i1_5 ), .ZN(\SB2_1_16/Component_Function_4/NAND4_in[3] ) );
  NAND4_X2 U12592 ( .A1(\SB2_2_4/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_2_4/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_2_4/Component_Function_0/NAND4_in[0] ), .A4(n6256), .ZN(
        \SB2_2_4/buf_output[0] ) );
  NAND3_X2 U12593 ( .A1(\SB2_2_4/i0_3 ), .A2(\SB2_2_4/i0_0 ), .A3(n6230), .ZN(
        n6256) );
  XOR2_X1 U12594 ( .A1(\RI5[2][35] ), .A2(\RI5[2][71] ), .Z(
        \MC_ARK_ARC_1_2/temp3[161] ) );
  NAND4_X2 U12595 ( .A1(\SB2_3_28/Component_Function_4/NAND4_in[2] ), .A2(
        \SB2_3_28/Component_Function_4/NAND4_in[0] ), .A3(n1320), .A4(
        \SB2_3_28/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB2_3_28/buf_output[4] ) );
  NAND3_X2 U12596 ( .A1(\SB2_1_12/i0_0 ), .A2(\SB2_1_12/i0_4 ), .A3(
        \SB2_1_12/i1_5 ), .ZN(n1009) );
  NAND3_X1 U12597 ( .A1(\SB2_3_5/i0_3 ), .A2(\SB2_3_5/i0[10] ), .A3(
        \SB2_3_5/i0_4 ), .ZN(\SB2_3_5/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U12598 ( .A1(n1571), .A2(\MC_ARK_ARC_1_2/temp1[39] ), .Z(
        \MC_ARK_ARC_1_2/temp5[39] ) );
  NAND3_X2 U12599 ( .A1(\SB1_3_30/i0[8] ), .A2(\SB1_3_30/i3[0] ), .A3(
        \SB1_3_30/i1_5 ), .ZN(n6257) );
  NAND3_X2 U12600 ( .A1(\SB2_3_23/i0[10] ), .A2(\SB2_3_23/i0_0 ), .A3(
        \SB2_3_23/i0[6] ), .ZN(n6258) );
  NAND4_X2 U12601 ( .A1(\SB3_5/Component_Function_3/NAND4_in[3] ), .A2(
        \SB3_5/Component_Function_3/NAND4_in[1] ), .A3(
        \SB3_5/Component_Function_3/NAND4_in[2] ), .A4(n2249), .ZN(
        \SB3_5/buf_output[3] ) );
  NAND3_X2 U12602 ( .A1(\SB1_3_30/i0[9] ), .A2(\SB1_3_30/i0[8] ), .A3(
        \SB1_3_30/i0_3 ), .ZN(n6287) );
  XOR2_X1 U12603 ( .A1(\RI5[0][117] ), .A2(\RI5[0][93] ), .Z(n6259) );
  NAND3_X1 U12604 ( .A1(\SB4_22/i0[9] ), .A2(\SB4_22/i1_5 ), .A3(
        \SB4_22/i0[6] ), .ZN(n6261) );
  XOR2_X1 U12605 ( .A1(\MC_ARK_ARC_1_3/temp6[29] ), .A2(n6262), .Z(
        \RI1[4][29] ) );
  XOR2_X1 U12606 ( .A1(\MC_ARK_ARC_1_3/temp1[29] ), .A2(n3230), .Z(n6262) );
  XOR2_X1 U12607 ( .A1(\MC_ARK_ARC_1_2/temp5[6] ), .A2(n6263), .Z(
        \MC_ARK_ARC_1_2/buf_output[6] ) );
  XOR2_X1 U12608 ( .A1(\MC_ARK_ARC_1_2/temp3[6] ), .A2(
        \MC_ARK_ARC_1_2/temp4[6] ), .Z(n6263) );
  NAND4_X2 U12609 ( .A1(\SB3_27/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_27/Component_Function_0/NAND4_in[1] ), .A3(
        \SB3_27/Component_Function_0/NAND4_in[0] ), .A4(n6264), .ZN(
        \SB3_27/buf_output[0] ) );
  XOR2_X1 U12610 ( .A1(\RI5[0][23] ), .A2(\RI5[0][191] ), .Z(n6265) );
  XOR2_X1 U12611 ( .A1(\RI5[0][190] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[22] ), 
        .Z(n6266) );
  NAND2_X1 U12612 ( .A1(\SB1_1_1/Component_Function_4/NAND4_in[3] ), .A2(n6276), .ZN(n6525) );
  XOR2_X1 U12613 ( .A1(n6267), .A2(\MC_ARK_ARC_1_0/temp4[64] ), .Z(
        \MC_ARK_ARC_1_0/temp6[64] ) );
  NAND4_X2 U12614 ( .A1(\SB2_3_23/Component_Function_2/NAND4_in[0] ), .A2(
        n3900), .A3(n4576), .A4(n6268), .ZN(\SB2_3_23/buf_output[2] ) );
  NAND3_X1 U12615 ( .A1(\SB4_20/i0[10] ), .A2(\SB4_20/i0_3 ), .A3(
        \SB4_20/i0[9] ), .ZN(n6269) );
  NAND3_X1 U12616 ( .A1(\SB1_3_7/buf_output[1] ), .A2(\SB1_3_8/buf_output[0] ), 
        .A3(\SB2_3_3/i1_5 ), .ZN(n6270) );
  NAND4_X2 U12617 ( .A1(\SB1_3_7/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_3_7/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_3_7/Component_Function_1/NAND4_in[0] ), .A4(n6271), .ZN(
        \SB1_3_7/buf_output[1] ) );
  NAND3_X1 U12618 ( .A1(\SB3_22/i0[6] ), .A2(\SB3_22/i1[9] ), .A3(
        \SB3_22/i0_3 ), .ZN(\SB3_22/Component_Function_3/NAND4_in[0] ) );
  XOR2_X1 U12619 ( .A1(\MC_ARK_ARC_1_2/temp5[145] ), .A2(
        \MC_ARK_ARC_1_2/temp6[145] ), .Z(\MC_ARK_ARC_1_2/buf_output[145] ) );
  XOR2_X1 U12620 ( .A1(n6272), .A2(n26), .Z(Ciphertext[186]) );
  NAND3_X2 U12621 ( .A1(\SB1_2_12/i0[10] ), .A2(\SB1_2_12/i1[9] ), .A3(
        \SB1_2_12/i1_5 ), .ZN(\SB1_2_12/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U12622 ( .A1(\RI5[2][147] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[141] ), .Z(\MC_ARK_ARC_1_2/temp1[147] ) );
  INV_X1 U12623 ( .I(\SB3_25/buf_output[3] ), .ZN(\SB4_23/i0[8] ) );
  XOR2_X1 U12624 ( .A1(n4145), .A2(\MC_ARK_ARC_1_2/temp6[152] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[152] ) );
  NAND4_X2 U12625 ( .A1(\SB2_2_8/Component_Function_5/NAND4_in[2] ), .A2(
        \SB2_2_8/Component_Function_5/NAND4_in[1] ), .A3(
        \SB2_2_8/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_2_8/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_2_8/buf_output[5] ) );
  XOR2_X1 U12626 ( .A1(\MC_ARK_ARC_1_3/temp5[75] ), .A2(
        \MC_ARK_ARC_1_3/temp6[75] ), .Z(\MC_ARK_ARC_1_3/buf_output[75] ) );
  NAND3_X2 U12627 ( .A1(\SB2_1_10/i0[10] ), .A2(\SB2_1_10/i1[9] ), .A3(
        \SB2_1_10/i1_7 ), .ZN(\SB2_1_10/Component_Function_3/NAND4_in[2] ) );
  NAND2_X1 U12628 ( .A1(\SB3_5/buf_output[3] ), .A2(\SB4_3/i0[9] ), .ZN(n6274)
         );
  NAND4_X2 U12629 ( .A1(n2598), .A2(
        \SB1_3_11/Component_Function_5/NAND4_in[3] ), .A3(
        \SB1_3_11/Component_Function_5/NAND4_in[0] ), .A4(n6275), .ZN(
        \SB1_3_11/buf_output[5] ) );
  NAND3_X1 U12630 ( .A1(\SB1_1_1/i0_0 ), .A2(\SB1_1_1/i0[9] ), .A3(
        \SB1_1_1/i0[8] ), .ZN(n6276) );
  NAND3_X2 U12631 ( .A1(\RI3[0][39] ), .A2(\SB2_0_25/i1[9] ), .A3(
        \SB2_0_25/i1_5 ), .ZN(\SB2_0_25/Component_Function_2/NAND4_in[0] ) );
  NAND4_X2 U12632 ( .A1(\SB2_1_18/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_1_18/Component_Function_3/NAND4_in[1] ), .A3(n4349), .A4(n6277), 
        .ZN(\SB2_1_18/buf_output[3] ) );
  NAND3_X2 U12633 ( .A1(\SB2_1_18/i1_7 ), .A2(\SB2_1_18/i0[10] ), .A3(
        \SB2_1_18/i1[9] ), .ZN(n6277) );
  NAND3_X2 U12634 ( .A1(\SB3_4/i0[8] ), .A2(n2910), .A3(\SB3_4/i3[0] ), .ZN(
        n6278) );
  INV_X2 U12635 ( .I(\RI3[0][86] ), .ZN(\SB2_0_17/i1[9] ) );
  NAND4_X2 U12636 ( .A1(\SB1_0_20/Component_Function_2/NAND4_in[3] ), .A2(
        \SB1_0_20/Component_Function_2/NAND4_in[2] ), .A3(
        \SB1_0_20/Component_Function_2/NAND4_in[0] ), .A4(n3442), .ZN(
        \RI3[0][86] ) );
  NAND3_X2 U12637 ( .A1(\SB2_3_11/i0_3 ), .A2(n3645), .A3(\SB2_3_11/i1[9] ), 
        .ZN(\SB2_3_11/Component_Function_5/NAND4_in[2] ) );
  NAND3_X1 U12638 ( .A1(\SB2_3_24/i0[6] ), .A2(\SB1_3_29/buf_output[0] ), .A3(
        \SB2_3_24/i1_5 ), .ZN(n1013) );
  XOR2_X1 U12639 ( .A1(\RI5[3][145] ), .A2(\RI5[3][181] ), .Z(
        \MC_ARK_ARC_1_3/temp3[79] ) );
  XOR2_X1 U12640 ( .A1(n6281), .A2(\MC_ARK_ARC_1_1/temp5[98] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[98] ) );
  XOR2_X1 U12641 ( .A1(\MC_ARK_ARC_1_1/temp3[98] ), .A2(
        \MC_ARK_ARC_1_1/temp4[98] ), .Z(n6281) );
  NAND4_X2 U12642 ( .A1(\SB2_3_3/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_3/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_3_3/Component_Function_4/NAND4_in[2] ), .A4(n6282), .ZN(
        \SB2_3_3/buf_output[4] ) );
  NAND3_X1 U12643 ( .A1(\SB4_15/i0[10] ), .A2(\SB4_15/i1[9] ), .A3(
        \SB4_15/i1_5 ), .ZN(\SB4_15/Component_Function_2/NAND4_in[0] ) );
  NAND2_X2 U12644 ( .A1(n4036), .A2(n6284), .ZN(\SB2_2_14/i0_4 ) );
  AND2_X1 U12645 ( .A1(n6302), .A2(\SB1_2_15/Component_Function_4/NAND4_in[3] ), .Z(n6284) );
  NAND3_X1 U12646 ( .A1(\SB3_18/i0[6] ), .A2(\SB3_18/i1_5 ), .A3(
        \SB3_18/i0[9] ), .ZN(n4057) );
  NAND3_X1 U12647 ( .A1(\SB1_1_23/i0_3 ), .A2(\SB1_1_23/i0[9] ), .A3(
        \SB1_1_23/i0[8] ), .ZN(n1766) );
  NAND3_X1 U12648 ( .A1(\SB2_1_5/i0[10] ), .A2(\SB2_1_5/i0_3 ), .A3(
        \SB2_1_5/i0[9] ), .ZN(n6285) );
  XOR2_X1 U12649 ( .A1(n6286), .A2(\MC_ARK_ARC_1_0/temp4[188] ), .Z(n3964) );
  XOR2_X1 U12650 ( .A1(\RI5[0][188] ), .A2(\RI5[0][182] ), .Z(n6286) );
  INV_X2 U12651 ( .I(\SB1_1_0/buf_output[3] ), .ZN(\SB2_1_30/i0[8] ) );
  NAND4_X2 U12652 ( .A1(\SB1_1_0/Component_Function_3/NAND4_in[0] ), .A2(n2599), .A3(n2211), .A4(\SB1_1_0/Component_Function_3/NAND4_in[1] ), .ZN(
        \SB1_1_0/buf_output[3] ) );
  NAND3_X1 U12653 ( .A1(\SB1_0_20/i0[8] ), .A2(\SB1_0_20/i0_3 ), .A3(
        \SB1_0_20/i1_7 ), .ZN(\SB1_0_20/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U12654 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[166] ), .A2(\RI5[3][160] ), .Z(n6288) );
  NAND4_X2 U12655 ( .A1(\SB2_2_4/Component_Function_2/NAND4_in[3] ), .A2(n6376), .A3(\SB2_2_4/Component_Function_2/NAND4_in[0] ), .A4(n6289), .ZN(
        \SB2_2_4/buf_output[2] ) );
  NAND3_X2 U12656 ( .A1(\SB2_2_4/i0_3 ), .A2(\SB2_2_4/i0[8] ), .A3(
        \SB2_2_4/i0[9] ), .ZN(n6289) );
  NAND4_X2 U12657 ( .A1(\SB2_3_15/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_3_15/Component_Function_0/NAND4_in[3] ), .A3(n3265), .A4(
        \SB2_3_15/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_3_15/buf_output[0] ) );
  NAND3_X1 U12658 ( .A1(\SB3_0/i0_3 ), .A2(\SB3_0/i0[8] ), .A3(\SB3_0/i1_7 ), 
        .ZN(\SB3_0/Component_Function_1/NAND4_in[1] ) );
  NAND3_X1 U12659 ( .A1(\SB4_5/i0_0 ), .A2(\SB4_5/i0[9] ), .A3(\SB4_5/i0[8] ), 
        .ZN(\SB4_5/Component_Function_4/NAND4_in[0] ) );
  XOR2_X1 U12660 ( .A1(\RI5[3][126] ), .A2(\RI5[3][102] ), .Z(
        \MC_ARK_ARC_1_3/temp2[156] ) );
  XOR2_X1 U12661 ( .A1(\RI5[1][77] ), .A2(\RI5[1][53] ), .Z(
        \MC_ARK_ARC_1_1/temp2[107] ) );
  NAND3_X1 U12662 ( .A1(\SB1_1_21/i0[6] ), .A2(\SB1_1_21/i0_3 ), .A3(
        \SB1_1_21/i1[9] ), .ZN(\SB1_1_21/Component_Function_3/NAND4_in[0] ) );
  NAND4_X2 U12663 ( .A1(\SB1_3_17/Component_Function_5/NAND4_in[3] ), .A2(
        n3976), .A3(\SB1_3_17/Component_Function_5/NAND4_in[1] ), .A4(
        \SB1_3_17/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_3_17/buf_output[5] ) );
  NAND4_X2 U12664 ( .A1(\SB2_2_30/Component_Function_5/NAND4_in[1] ), .A2(
        n3485), .A3(\SB2_2_30/Component_Function_5/NAND4_in[3] ), .A4(
        \SB2_2_30/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB2_2_30/buf_output[5] ) );
  NAND4_X2 U12665 ( .A1(\SB1_2_19/Component_Function_5/NAND4_in[3] ), .A2(
        n3277), .A3(\SB1_2_19/Component_Function_5/NAND4_in[0] ), .A4(
        \SB1_2_19/Component_Function_5/NAND4_in[1] ), .ZN(
        \SB1_2_19/buf_output[5] ) );
  NAND4_X2 U12666 ( .A1(\SB3_31/Component_Function_2/NAND4_in[0] ), .A2(
        \SB3_31/Component_Function_2/NAND4_in[1] ), .A3(
        \SB3_31/Component_Function_2/NAND4_in[2] ), .A4(
        \SB3_31/Component_Function_2/NAND4_in[3] ), .ZN(\SB3_31/buf_output[2] ) );
  XOR2_X1 U12667 ( .A1(\MC_ARK_ARC_1_2/temp3[82] ), .A2(
        \MC_ARK_ARC_1_2/temp4[82] ), .Z(\MC_ARK_ARC_1_2/temp6[82] ) );
  XOR2_X1 U12668 ( .A1(\RI5[2][51] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[27] ), 
        .Z(n1873) );
  NAND4_X2 U12669 ( .A1(\SB2_1_8/Component_Function_4/NAND4_in[1] ), .A2(
        \SB2_1_8/Component_Function_4/NAND4_in[0] ), .A3(
        \SB2_1_8/Component_Function_4/NAND4_in[2] ), .A4(n6290), .ZN(
        \SB2_1_8/buf_output[4] ) );
  XOR2_X1 U12670 ( .A1(\MC_ARK_ARC_1_1/temp5[2] ), .A2(n6291), .Z(
        \MC_ARK_ARC_1_1/buf_output[2] ) );
  XOR2_X1 U12671 ( .A1(\MC_ARK_ARC_1_1/temp3[2] ), .A2(
        \MC_ARK_ARC_1_1/temp4[2] ), .Z(n6291) );
  NAND3_X2 U12672 ( .A1(\SB1_3_15/i0_0 ), .A2(\SB1_3_15/i0_4 ), .A3(
        \SB1_3_15/i1_5 ), .ZN(\SB1_3_15/Component_Function_2/NAND4_in[3] ) );
  XOR2_X1 U12673 ( .A1(n2110), .A2(n6292), .Z(n4658) );
  XOR2_X1 U12674 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[132] ), .A2(\RI5[3][138] ), .Z(n6292) );
  NAND3_X1 U12675 ( .A1(\SB4_7/i0_4 ), .A2(\SB4_7/i0_3 ), .A3(\SB4_7/i1[9] ), 
        .ZN(n6293) );
  NAND4_X2 U12676 ( .A1(\SB2_3_14/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_3_14/Component_Function_0/NAND4_in[3] ), .A3(
        \SB2_3_14/Component_Function_0/NAND4_in[0] ), .A4(n6294), .ZN(
        \SB2_3_14/buf_output[0] ) );
  NAND3_X1 U12677 ( .A1(\SB2_3_14/i0_3 ), .A2(\SB2_3_14/i0[10] ), .A3(
        \SB2_3_14/i0_4 ), .ZN(n6294) );
  XOR2_X1 U12678 ( .A1(\RI5[1][143] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[179] ), .Z(\MC_ARK_ARC_1_1/temp3[77] ) );
  XOR2_X1 U12679 ( .A1(n6295), .A2(\MC_ARK_ARC_1_2/temp4[179] ), .Z(
        \MC_ARK_ARC_1_2/temp6[179] ) );
  XOR2_X1 U12680 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[53] ), .A2(\RI5[2][89] ), 
        .Z(n6295) );
  NAND3_X2 U12681 ( .A1(\SB2_1_8/i0_4 ), .A2(n2745), .A3(\SB2_1_8/i0[6] ), 
        .ZN(n1853) );
  NAND3_X2 U12682 ( .A1(\SB2_3_27/i0_4 ), .A2(\SB2_3_27/i0_3 ), .A3(
        \SB2_3_27/i0_0 ), .ZN(\SB2_3_27/Component_Function_3/NAND4_in[1] ) );
  NAND3_X2 U12683 ( .A1(\SB2_3_5/i0_3 ), .A2(n3671), .A3(\SB2_3_5/i0_4 ), .ZN(
        n4372) );
  NAND3_X1 U12684 ( .A1(\SB4_13/i0_0 ), .A2(\SB4_13/i0[9] ), .A3(n3683), .ZN(
        \SB4_13/Component_Function_4/NAND4_in[0] ) );
  NAND4_X2 U12685 ( .A1(\SB2_0_1/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_0_1/Component_Function_3/NAND4_in[0] ), .A3(
        \SB2_0_1/Component_Function_3/NAND4_in[1] ), .A4(n6296), .ZN(
        \SB2_0_1/buf_output[3] ) );
  NAND3_X2 U12686 ( .A1(\SB2_0_1/i3[0] ), .A2(\SB2_0_1/i1_5 ), .A3(
        \SB2_0_1/i0[8] ), .ZN(n6296) );
  XOR2_X1 U12687 ( .A1(\RI5[1][37] ), .A2(\RI5[1][61] ), .Z(n1628) );
  NAND3_X1 U12688 ( .A1(\SB1_3_28/i0_0 ), .A2(\SB1_3_28/i1_7 ), .A3(
        \SB1_3_28/i3[0] ), .ZN(\SB1_3_28/Component_Function_4/NAND4_in[1] ) );
  XOR2_X1 U12689 ( .A1(\MC_ARK_ARC_1_1/temp2[21] ), .A2(
        \MC_ARK_ARC_1_1/temp1[21] ), .Z(\MC_ARK_ARC_1_1/temp5[21] ) );
  XOR2_X1 U12690 ( .A1(\MC_ARK_ARC_1_0/temp6[169] ), .A2(
        \MC_ARK_ARC_1_0/temp5[169] ), .Z(\MC_ARK_ARC_1_0/buf_output[169] ) );
  NAND3_X1 U12691 ( .A1(\SB1_3_7/i0[6] ), .A2(\SB1_3_7/i1[9] ), .A3(
        \SB1_3_7/i0_3 ), .ZN(n6297) );
  NAND3_X2 U12692 ( .A1(\SB2_1_6/i0_4 ), .A2(\SB2_1_6/i0[6] ), .A3(
        \SB2_1_6/i0[9] ), .ZN(n6298) );
  INV_X1 U12693 ( .I(\SB3_0/buf_output[5] ), .ZN(\SB4_0/i1_5 ) );
  NAND3_X2 U12694 ( .A1(\SB1_3_13/i0[8] ), .A2(\SB1_3_13/i1_5 ), .A3(
        \SB1_3_13/i3[0] ), .ZN(n1426) );
  NAND4_X2 U12695 ( .A1(\SB1_1_0/Component_Function_5/NAND4_in[2] ), .A2(n2315), .A3(\SB1_1_0/Component_Function_5/NAND4_in[0] ), .A4(n6299), .ZN(
        \SB1_1_0/buf_output[5] ) );
  NAND4_X2 U12696 ( .A1(\SB3_22/Component_Function_2/NAND4_in[1] ), .A2(
        \SB3_22/Component_Function_2/NAND4_in[2] ), .A3(
        \SB3_22/Component_Function_2/NAND4_in[0] ), .A4(n3494), .ZN(
        \SB3_22/buf_output[2] ) );
  INV_X2 U12697 ( .I(n6300), .ZN(n567) );
  NAND3_X2 U12698 ( .A1(\SB1_2_15/i0[10] ), .A2(\SB1_2_15/i0_3 ), .A3(
        \SB1_2_15/i0[9] ), .ZN(n6302) );
  XOR2_X1 U12699 ( .A1(\RI5[1][71] ), .A2(\RI5[1][47] ), .Z(n6303) );
  NAND3_X1 U12700 ( .A1(n2074), .A2(\SB2_2_6/i1_7 ), .A3(\SB2_2_6/i0[8] ), 
        .ZN(\SB2_2_6/Component_Function_1/NAND4_in[3] ) );
  NAND3_X2 U12701 ( .A1(\SB1_3_8/i0[6] ), .A2(\SB1_3_8/i0_4 ), .A3(
        \SB1_3_8/i0[9] ), .ZN(n6304) );
  XOR2_X1 U12702 ( .A1(\MC_ARK_ARC_1_3/temp6[191] ), .A2(n6305), .Z(
        \MC_ARK_ARC_1_3/buf_output[191] ) );
  NAND3_X2 U12703 ( .A1(\SB1_3_17/i0_4 ), .A2(\SB1_3_17/i1[9] ), .A3(
        \SB1_3_17/i1_5 ), .ZN(n6306) );
  XOR2_X1 U12704 ( .A1(\RI5[3][105] ), .A2(\RI5[3][99] ), .Z(n6307) );
  NAND3_X2 U12705 ( .A1(\SB2_3_31/i0_3 ), .A2(\SB2_3_31/i1[9] ), .A3(
        \SB2_3_31/i0_4 ), .ZN(n2339) );
  NAND4_X2 U12706 ( .A1(\SB1_2_17/Component_Function_4/NAND4_in[0] ), .A2(
        \SB1_2_17/Component_Function_4/NAND4_in[1] ), .A3(
        \SB1_2_17/Component_Function_4/NAND4_in[3] ), .A4(n6308), .ZN(
        \SB1_2_17/buf_output[4] ) );
  NAND2_X1 U12707 ( .A1(\SB1_0_7/Component_Function_4/NAND4_in[1] ), .A2(n1671), .ZN(n6360) );
  XOR2_X1 U12708 ( .A1(n2199), .A2(\MC_ARK_ARC_1_0/temp4[133] ), .Z(n6309) );
  XOR2_X1 U12709 ( .A1(\MC_ARK_ARC_1_0/temp3[133] ), .A2(n2198), .Z(n6310) );
  NAND3_X1 U12710 ( .A1(\SB2_1_9/i0_4 ), .A2(\SB2_1_9/i1[9] ), .A3(
        \SB2_1_9/i1_5 ), .ZN(\SB2_1_9/Component_Function_4/NAND4_in[3] ) );
  XOR2_X1 U12711 ( .A1(n6311), .A2(\MC_ARK_ARC_1_2/temp6[179] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[179] ) );
  XOR2_X1 U12712 ( .A1(\MC_ARK_ARC_1_2/temp1[179] ), .A2(
        \MC_ARK_ARC_1_2/temp2[179] ), .Z(n6311) );
  NAND4_X2 U12713 ( .A1(n4716), .A2(\SB1_0_5/Component_Function_2/NAND4_in[0] ), .A3(n4241), .A4(\SB1_0_5/Component_Function_2/NAND4_in[2] ), .ZN(
        \SB1_0_5/buf_output[2] ) );
  NAND3_X1 U12714 ( .A1(n5492), .A2(\SB4_8/i1_7 ), .A3(\SB4_8/i3[0] ), .ZN(
        n3175) );
  XOR2_X1 U12715 ( .A1(n3156), .A2(n3901), .Z(\MC_ARK_ARC_1_3/temp5[11] ) );
  NAND3_X1 U12716 ( .A1(\SB1_0_0/i1_7 ), .A2(\SB1_0_0/i0[10] ), .A3(
        \SB1_0_0/i1[9] ), .ZN(\SB1_0_0/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U12717 ( .A1(\SB1_1_5/i0[6] ), .A2(\SB1_1_5/i0[8] ), .A3(
        \SB1_1_5/i0[7] ), .ZN(\SB1_1_5/Component_Function_0/NAND4_in[1] ) );
  NAND3_X2 U12718 ( .A1(\SB2_1_16/i0_3 ), .A2(\SB2_1_16/i0[8] ), .A3(
        \SB2_1_16/i1_7 ), .ZN(\SB2_1_16/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U12719 ( .A1(n6313), .A2(n6312), .Z(n6520) );
  XOR2_X1 U12720 ( .A1(\RI5[1][122] ), .A2(\RI5[1][176] ), .Z(n6312) );
  XOR2_X1 U12721 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[170] ), .A2(\RI5[1][146] ), .Z(n6313) );
  INV_X2 U12722 ( .I(\SB3_0/buf_output[2] ), .ZN(\SB4_29/i1[9] ) );
  BUF_X2 U12723 ( .I(n348), .Z(n6314) );
  NAND3_X1 U12724 ( .A1(\SB2_2_1/i0[10] ), .A2(\SB2_2_1/i0_3 ), .A3(
        \SB2_2_1/i0[9] ), .ZN(n6315) );
  NAND4_X2 U12725 ( .A1(\SB1_0_20/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_0_20/Component_Function_1/NAND4_in[1] ), .A3(n6350), .A4(
        \SB1_0_20/Component_Function_1/NAND4_in[0] ), .ZN(\RI3[0][91] ) );
  XOR2_X1 U12726 ( .A1(n6317), .A2(n6316), .Z(n1527) );
  XOR2_X1 U12727 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[185] ), .A2(n177), .Z(
        n6316) );
  XOR2_X1 U12728 ( .A1(\RI5[1][149] ), .A2(\RI5[1][119] ), .Z(n6317) );
  NOR2_X2 U12729 ( .A1(n3993), .A2(n4768), .ZN(n3992) );
  NAND3_X1 U12730 ( .A1(\SB1_1_15/i0_4 ), .A2(\SB1_1_15/i0[10] ), .A3(
        \SB1_1_15/i0_3 ), .ZN(\SB1_1_15/Component_Function_0/NAND4_in[2] ) );
  XOR2_X1 U12731 ( .A1(n4657), .A2(\MC_ARK_ARC_1_1/temp6[81] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[81] ) );
  XOR2_X1 U12732 ( .A1(\MC_ARK_ARC_1_1/temp1[81] ), .A2(
        \MC_ARK_ARC_1_1/temp2[81] ), .Z(n4657) );
  NAND4_X2 U12733 ( .A1(\SB2_0_30/Component_Function_2/NAND4_in[3] ), .A2(
        \SB2_0_30/Component_Function_2/NAND4_in[1] ), .A3(n3098), .A4(n6318), 
        .ZN(\SB2_0_30/buf_output[2] ) );
  NAND3_X2 U12734 ( .A1(\SB2_0_30/i0[9] ), .A2(\SB2_0_30/i0_3 ), .A3(
        \SB2_0_30/i0[8] ), .ZN(n6318) );
  XOR2_X1 U12735 ( .A1(n6319), .A2(\MC_ARK_ARC_1_0/temp5[116] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[116] ) );
  XOR2_X1 U12736 ( .A1(n6516), .A2(\MC_ARK_ARC_1_0/temp4[116] ), .Z(n6319) );
  INV_X1 U12737 ( .I(\SB3_6/buf_output[5] ), .ZN(\SB4_6/i1_5 ) );
  NAND4_X2 U12738 ( .A1(\SB3_6/Component_Function_5/NAND4_in[2] ), .A2(
        \SB3_6/Component_Function_5/NAND4_in[3] ), .A3(
        \SB3_6/Component_Function_5/NAND4_in[1] ), .A4(
        \SB3_6/Component_Function_5/NAND4_in[0] ), .ZN(\SB3_6/buf_output[5] )
         );
  XOR2_X1 U12739 ( .A1(\SB2_0_16/buf_output[2] ), .A2(\SB2_0_11/buf_output[2] ), .Z(n6320) );
  XOR2_X1 U12740 ( .A1(n6322), .A2(n6321), .Z(\MC_ARK_ARC_1_0/buf_output[158] ) );
  XOR2_X1 U12741 ( .A1(n2846), .A2(n4197), .Z(n6321) );
  XOR2_X1 U12742 ( .A1(n4198), .A2(\MC_ARK_ARC_1_0/temp1[158] ), .Z(n6322) );
  XOR2_X1 U12743 ( .A1(n6324), .A2(n6323), .Z(n6326) );
  XOR2_X1 U12744 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[56] ), .A2(\RI5[2][20] ), 
        .Z(n6323) );
  XOR2_X1 U12745 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[146] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[92] ), .Z(n6324) );
  NAND4_X2 U12746 ( .A1(\SB2_1_14/Component_Function_0/NAND4_in[1] ), .A2(
        \SB2_1_14/Component_Function_0/NAND4_in[2] ), .A3(
        \SB2_1_14/Component_Function_0/NAND4_in[0] ), .A4(n6325), .ZN(
        \SB2_1_14/buf_output[0] ) );
  NAND3_X2 U12747 ( .A1(\SB2_1_14/i0_3 ), .A2(\SB2_1_14/i0_0 ), .A3(
        \SB2_1_14/i0[7] ), .ZN(n6325) );
  NAND3_X2 U12748 ( .A1(\SB1_2_5/i0[10] ), .A2(\SB1_2_5/i1[9] ), .A3(
        \SB1_2_5/i1_7 ), .ZN(n6353) );
  XOR2_X1 U12749 ( .A1(\RI5[3][10] ), .A2(\RI5[3][148] ), .Z(n3826) );
  XOR2_X1 U12750 ( .A1(\RI5[0][6] ), .A2(\RI5[0][30] ), .Z(
        \MC_ARK_ARC_1_0/temp2[60] ) );
  NAND3_X2 U12751 ( .A1(\SB1_2_13/i0[6] ), .A2(\SB1_2_13/i0_3 ), .A3(
        \SB1_2_13/i1[9] ), .ZN(n2122) );
  NAND4_X2 U12752 ( .A1(\SB1_1_14/Component_Function_3/NAND4_in[1] ), .A2(
        n3698), .A3(\SB1_1_14/Component_Function_3/NAND4_in[3] ), .A4(n6329), 
        .ZN(\SB1_1_14/buf_output[3] ) );
  NAND3_X2 U12753 ( .A1(\SB1_1_14/i0[6] ), .A2(\SB1_1_14/i1[9] ), .A3(
        \SB1_1_14/i0_3 ), .ZN(n6329) );
  INV_X2 U12754 ( .I(n6330), .ZN(n2911) );
  NAND4_X2 U12755 ( .A1(\SB2_3_11/Component_Function_3/NAND4_in[3] ), .A2(
        \SB2_3_11/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_3_11/Component_Function_3/NAND4_in[0] ), .A4(n6331), .ZN(
        \SB2_3_11/buf_output[3] ) );
  NAND4_X2 U12756 ( .A1(\SB1_0_5/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_0_5/Component_Function_1/NAND4_in[2] ), .A3(n6337), .A4(n6332), 
        .ZN(\SB1_0_5/buf_output[1] ) );
  XOR2_X1 U12757 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[136] ), .A2(\RI5[2][142] ), .Z(\MC_ARK_ARC_1_2/temp1[142] ) );
  NAND3_X1 U12758 ( .A1(\SB4_7/i0_4 ), .A2(\SB4_7/i1[9] ), .A3(\SB4_7/i1_5 ), 
        .ZN(n6333) );
  XOR2_X1 U12759 ( .A1(\MC_ARK_ARC_1_1/temp2[109] ), .A2(
        \MC_ARK_ARC_1_1/temp1[109] ), .Z(n6334) );
  XOR2_X1 U12760 ( .A1(\MC_ARK_ARC_1_1/temp5[32] ), .A2(n6335), .Z(
        \MC_ARK_ARC_1_1/buf_output[32] ) );
  XOR2_X1 U12761 ( .A1(\MC_ARK_ARC_1_1/temp4[32] ), .A2(
        \MC_ARK_ARC_1_1/temp3[32] ), .Z(n6335) );
  XOR2_X1 U12762 ( .A1(n6336), .A2(n3919), .Z(\MC_ARK_ARC_1_0/buf_output[88] )
         );
  XOR2_X1 U12763 ( .A1(\MC_ARK_ARC_1_0/temp3[88] ), .A2(
        \MC_ARK_ARC_1_0/temp4[88] ), .Z(n6336) );
  NAND3_X1 U12764 ( .A1(\SB1_0_5/i0[8] ), .A2(\SB1_0_5/i1_7 ), .A3(
        \SB1_0_5/i0_4 ), .ZN(n6337) );
  NAND3_X2 U12765 ( .A1(\SB2_0_1/i0[10] ), .A2(\SB2_0_1/i0[6] ), .A3(
        \SB2_0_1/i0_3 ), .ZN(n6338) );
  XOR2_X1 U12766 ( .A1(n1416), .A2(n6339), .Z(n1634) );
  XOR2_X1 U12767 ( .A1(\RI5[0][134] ), .A2(\RI5[0][8] ), .Z(n6339) );
  NAND3_X1 U12768 ( .A1(\SB2_1_9/i0[9] ), .A2(\SB2_1_9/i0[6] ), .A3(
        \SB2_1_9/i1_5 ), .ZN(\SB2_1_9/Component_Function_1/NAND4_in[2] ) );
  XOR2_X1 U12769 ( .A1(n1682), .A2(n6340), .Z(\MC_ARK_ARC_1_0/buf_output[35] )
         );
  NAND4_X2 U12770 ( .A1(\SB2_1_14/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_1_14/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_1_14/Component_Function_4/NAND4_in[0] ), .A4(n6341), .ZN(
        \SB2_1_14/buf_output[4] ) );
  NAND3_X2 U12771 ( .A1(\SB2_1_14/i0_3 ), .A2(\SB2_1_14/i0[10] ), .A3(
        \SB2_1_14/i0[9] ), .ZN(n6341) );
  XOR2_X1 U12772 ( .A1(n3996), .A2(\MC_ARK_ARC_1_0/temp1[72] ), .Z(
        \MC_ARK_ARC_1_0/temp5[72] ) );
  NAND4_X2 U12773 ( .A1(\SB3_0/Component_Function_4/NAND4_in[3] ), .A2(
        \SB3_0/Component_Function_4/NAND4_in[0] ), .A3(
        \SB3_0/Component_Function_4/NAND4_in[2] ), .A4(
        \SB3_0/Component_Function_4/NAND4_in[1] ), .ZN(\SB3_0/buf_output[4] )
         );
  XOR2_X1 U12774 ( .A1(\MC_ARK_ARC_1_2/temp5[18] ), .A2(n6342), .Z(
        \MC_ARK_ARC_1_2/buf_output[18] ) );
  XOR2_X1 U12775 ( .A1(\MC_ARK_ARC_1_2/temp3[18] ), .A2(
        \MC_ARK_ARC_1_2/temp4[18] ), .Z(n6342) );
  NAND3_X2 U12776 ( .A1(\SB2_1_10/i0[10] ), .A2(\SB2_1_10/i1[9] ), .A3(
        \SB2_1_10/i1_5 ), .ZN(\SB2_1_10/Component_Function_2/NAND4_in[0] ) );
  NAND3_X2 U12777 ( .A1(\RI3[0][76] ), .A2(\SB2_0_19/i0_3 ), .A3(
        \SB2_0_19/i1[9] ), .ZN(n6343) );
  XOR2_X1 U12778 ( .A1(n6344), .A2(n42), .Z(Ciphertext[98]) );
  XOR2_X1 U12779 ( .A1(\MC_ARK_ARC_1_3/temp4[123] ), .A2(n6346), .Z(
        \MC_ARK_ARC_1_3/temp6[123] ) );
  XOR2_X1 U12780 ( .A1(\RI5[3][33] ), .A2(\RI5[3][189] ), .Z(n6346) );
  NAND3_X1 U12781 ( .A1(\SB1_0_20/i0_0 ), .A2(\SB1_0_20/i0[8] ), .A3(
        \SB1_0_20/i0[9] ), .ZN(n6347) );
  NAND3_X1 U12782 ( .A1(\SB4_20/i0_4 ), .A2(n3674), .A3(\SB4_20/i0_0 ), .ZN(
        n6348) );
  XOR2_X1 U12783 ( .A1(n6351), .A2(n36), .Z(Ciphertext[124]) );
  NAND4_X2 U12784 ( .A1(\SB4_11/Component_Function_4/NAND4_in[3] ), .A2(n2636), 
        .A3(n3626), .A4(n4547), .ZN(n6351) );
  XOR2_X1 U12785 ( .A1(\MC_ARK_ARC_1_0/temp5[107] ), .A2(n6352), .Z(
        \MC_ARK_ARC_1_0/buf_output[107] ) );
  XOR2_X1 U12786 ( .A1(\MC_ARK_ARC_1_0/temp4[107] ), .A2(
        \MC_ARK_ARC_1_0/temp3[107] ), .Z(n6352) );
  NAND3_X2 U12787 ( .A1(\SB2_1_2/i0[10] ), .A2(\SB2_1_2/i1_5 ), .A3(
        \SB2_1_2/i1[9] ), .ZN(\SB2_1_2/Component_Function_2/NAND4_in[0] ) );
  XOR2_X1 U12788 ( .A1(\RI5[0][95] ), .A2(\RI5[0][119] ), .Z(n6354) );
  NAND3_X2 U12789 ( .A1(\SB2_2_2/i1[9] ), .A2(\SB2_2_2/i0[10] ), .A3(
        \SB2_2_2/i1_5 ), .ZN(n4582) );
  NAND3_X1 U12790 ( .A1(\SB1_2_5/i0[10] ), .A2(\SB1_2_5/i1[9] ), .A3(
        \SB1_2_5/i1_5 ), .ZN(n6355) );
  NAND3_X1 U12791 ( .A1(\SB2_1_5/i0[8] ), .A2(\SB2_1_5/i3[0] ), .A3(
        \SB2_1_5/i1_5 ), .ZN(\SB2_1_5/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U12792 ( .A1(\RI5[3][107] ), .A2(\RI5[3][131] ), .Z(
        \MC_ARK_ARC_1_3/temp2[161] ) );
  NAND4_X2 U12793 ( .A1(\SB2_3_31/Component_Function_0/NAND4_in[2] ), .A2(
        \SB2_3_31/Component_Function_0/NAND4_in[1] ), .A3(n924), .A4(
        \SB2_3_31/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_3_31/buf_output[0] ) );
  NAND3_X1 U12794 ( .A1(\SB4_8/i0_0 ), .A2(\SB4_8/i0[6] ), .A3(\SB4_8/i0[10] ), 
        .ZN(\SB4_8/Component_Function_5/NAND4_in[1] ) );
  NAND4_X2 U12795 ( .A1(n6463), .A2(\SB1_2_0/Component_Function_3/NAND4_in[0] ), .A3(\SB1_2_0/Component_Function_3/NAND4_in[2] ), .A4(n6357), .ZN(
        \SB1_2_0/buf_output[3] ) );
  NAND3_X2 U12796 ( .A1(\SB1_2_0/i1_5 ), .A2(\SB1_2_0/i3[0] ), .A3(
        \SB1_2_0/i0[8] ), .ZN(n6357) );
  NOR2_X2 U12797 ( .A1(n6360), .A2(n6359), .ZN(\SB2_0_6/i0[7] ) );
  NAND2_X1 U12798 ( .A1(n3621), .A2(\SB1_0_7/Component_Function_4/NAND4_in[0] ), .ZN(n6359) );
  NAND4_X2 U12799 ( .A1(\SB2_3_4/Component_Function_2/NAND4_in[1] ), .A2(n3465), .A3(n1896), .A4(n6362), .ZN(\SB2_3_4/buf_output[2] ) );
  XOR2_X1 U12800 ( .A1(n6364), .A2(\MC_ARK_ARC_1_0/temp2[171] ), .Z(
        \MC_ARK_ARC_1_0/temp5[171] ) );
  NAND4_X2 U12801 ( .A1(\SB2_2_0/Component_Function_0/NAND4_in[1] ), .A2(n3268), .A3(n3269), .A4(\SB2_2_0/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB2_2_0/buf_output[0] ) );
  NAND3_X1 U12802 ( .A1(\SB1_0_20/i0[8] ), .A2(\SB1_0_20/i0_3 ), .A3(
        \SB1_0_20/i0[9] ), .ZN(\SB1_0_20/Component_Function_2/NAND4_in[2] ) );
  INV_X2 U12803 ( .I(\SB1_3_31/buf_output[1] ), .ZN(\SB2_3_27/i1_7 ) );
  NAND4_X2 U12804 ( .A1(\SB1_3_31/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_3_31/Component_Function_1/NAND4_in[1] ), .A3(n3731), .A4(
        \SB1_3_31/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_3_31/buf_output[1] ) );
  XOR2_X1 U12805 ( .A1(n4146), .A2(n6366), .Z(\MC_ARK_ARC_1_3/buf_output[90] )
         );
  XOR2_X1 U12806 ( .A1(\MC_ARK_ARC_1_3/temp1[90] ), .A2(n4457), .Z(n6366) );
  XOR2_X1 U12807 ( .A1(n6367), .A2(n1325), .Z(\MC_ARK_ARC_1_1/buf_output[186] ) );
  XOR2_X1 U12808 ( .A1(\MC_ARK_ARC_1_1/temp2[186] ), .A2(
        \MC_ARK_ARC_1_1/temp1[186] ), .Z(n6367) );
  NAND2_X1 U12809 ( .A1(\SB1_0_20/Component_Function_4/NAND4_in[1] ), .A2(
        n2613), .ZN(n6438) );
  NAND2_X2 U12810 ( .A1(\SB1_3_11/i0_3 ), .A2(\SB1_3_11/i1[9] ), .ZN(n6368) );
  XOR2_X1 U12811 ( .A1(n6370), .A2(\MC_ARK_ARC_1_2/temp5[103] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[103] ) );
  XOR2_X1 U12812 ( .A1(\MC_ARK_ARC_1_2/temp4[103] ), .A2(
        \MC_ARK_ARC_1_2/temp3[103] ), .Z(n6370) );
  NAND3_X2 U12813 ( .A1(\SB1_2_12/i0[9] ), .A2(\SB1_2_12/i0[6] ), .A3(
        \SB1_2_12/i0_4 ), .ZN(n6371) );
  NAND3_X2 U12814 ( .A1(\SB2_1_22/i0_4 ), .A2(\SB2_1_22/i0_3 ), .A3(
        \SB2_1_22/i0_0 ), .ZN(\SB2_1_22/Component_Function_3/NAND4_in[1] ) );
  NAND3_X1 U12815 ( .A1(\SB4_29/i0_3 ), .A2(\SB4_29/i1[9] ), .A3(
        \SB4_29/i0[6] ), .ZN(n6372) );
  NAND4_X2 U12816 ( .A1(\SB2_1_26/Component_Function_5/NAND4_in[3] ), .A2(
        \SB2_1_26/Component_Function_5/NAND4_in[1] ), .A3(n3392), .A4(n6373), 
        .ZN(\SB2_1_26/buf_output[5] ) );
  NAND3_X2 U12817 ( .A1(\SB2_1_26/i0_4 ), .A2(\SB2_1_26/i0_3 ), .A3(
        \SB2_1_26/i1[9] ), .ZN(n6373) );
  NAND4_X2 U12818 ( .A1(n1831), .A2(\SB2_2_8/Component_Function_4/NAND4_in[2] ), .A3(\SB2_2_8/Component_Function_4/NAND4_in[0] ), .A4(
        \SB2_2_8/Component_Function_4/NAND4_in[1] ), .ZN(
        \SB2_2_8/buf_output[4] ) );
  NAND3_X2 U12819 ( .A1(\SB2_2_16/i0_4 ), .A2(\SB2_2_16/i0[9] ), .A3(
        \SB2_2_16/i0[6] ), .ZN(n4022) );
  NAND3_X2 U12820 ( .A1(\SB2_0_18/i0[10] ), .A2(\SB2_0_18/i0_3 ), .A3(
        \SB2_0_18/i0[6] ), .ZN(n6411) );
  XOR2_X1 U12821 ( .A1(\MC_ARK_ARC_1_3/temp2[15] ), .A2(
        \MC_ARK_ARC_1_3/temp1[15] ), .Z(\MC_ARK_ARC_1_3/temp5[15] ) );
  XOR2_X1 U12822 ( .A1(n6374), .A2(n165), .Z(Ciphertext[177]) );
  NAND4_X2 U12823 ( .A1(\SB4_2/Component_Function_3/NAND4_in[1] ), .A2(
        \SB4_2/Component_Function_3/NAND4_in[0] ), .A3(
        \SB4_2/Component_Function_3/NAND4_in[2] ), .A4(
        \SB4_2/Component_Function_3/NAND4_in[3] ), .ZN(n6374) );
  XOR2_X1 U12824 ( .A1(\RI5[3][69] ), .A2(\RI5[3][93] ), .Z(
        \MC_ARK_ARC_1_3/temp2[123] ) );
  NAND3_X2 U12825 ( .A1(\SB1_3_24/i0_4 ), .A2(\SB1_3_24/i0_3 ), .A3(
        \SB1_3_24/i0_0 ), .ZN(n6375) );
  NAND3_X2 U12826 ( .A1(\SB2_2_4/i0[6] ), .A2(\SB2_2_4/i0_3 ), .A3(
        \SB2_2_4/i0[10] ), .ZN(n6376) );
  NAND3_X2 U12827 ( .A1(\SB3_0/i0[10] ), .A2(\SB3_0/i1[9] ), .A3(\SB3_0/i1_5 ), 
        .ZN(n6378) );
  NAND3_X1 U12828 ( .A1(\SB4_9/i0[10] ), .A2(\SB4_9/i0_3 ), .A3(\SB4_9/i0[6] ), 
        .ZN(n6379) );
  NAND4_X2 U12829 ( .A1(n2440), .A2(\SB1_1_0/Component_Function_1/NAND4_in[3] ), .A3(n1980), .A4(n6380), .ZN(\SB1_1_0/buf_output[1] ) );
  NAND3_X1 U12830 ( .A1(\SB1_1_0/i0_3 ), .A2(\SB1_1_0/i0[8] ), .A3(
        \SB1_1_0/i1_7 ), .ZN(n6380) );
  NAND3_X1 U12831 ( .A1(\SB4_9/i0[10] ), .A2(\SB4_9/i0_3 ), .A3(\SB4_9/i0[9] ), 
        .ZN(n6381) );
  XOR2_X1 U12832 ( .A1(\MC_ARK_ARC_1_2/temp1[103] ), .A2(
        \MC_ARK_ARC_1_2/temp2[103] ), .Z(\MC_ARK_ARC_1_2/temp5[103] ) );
  XOR2_X1 U12833 ( .A1(\SB2_2_10/buf_output[0] ), .A2(\RI5[2][180] ), .Z(
        \MC_ARK_ARC_1_2/temp2[18] ) );
  XOR2_X1 U12834 ( .A1(\RI5[2][51] ), .A2(\RI5[2][75] ), .Z(
        \MC_ARK_ARC_1_2/temp2[105] ) );
  NAND3_X1 U12835 ( .A1(\SB1_3_13/i0_3 ), .A2(\SB1_3_13/i0_0 ), .A3(
        \SB1_3_13/i0[7] ), .ZN(n2492) );
  NAND4_X2 U12836 ( .A1(\SB2_2_19/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_19/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_2_19/Component_Function_3/NAND4_in[3] ), .A4(n6383), .ZN(
        \SB2_2_19/buf_output[3] ) );
  XOR2_X1 U12837 ( .A1(\MC_ARK_ARC_1_1/temp2[172] ), .A2(n6384), .Z(
        \MC_ARK_ARC_1_1/temp5[172] ) );
  XOR2_X1 U12838 ( .A1(\RI5[1][172] ), .A2(\RI5[1][166] ), .Z(n6384) );
  NAND4_X2 U12839 ( .A1(\SB2_2_25/Component_Function_1/NAND4_in[1] ), .A2(
        \SB2_2_25/Component_Function_1/NAND4_in[3] ), .A3(
        \SB2_2_25/Component_Function_1/NAND4_in[0] ), .A4(n6386), .ZN(
        \SB2_2_25/buf_output[1] ) );
  NAND3_X1 U12840 ( .A1(\SB2_2_25/i0[6] ), .A2(\SB2_2_25/i0[9] ), .A3(
        \SB2_2_25/i1_5 ), .ZN(n6386) );
  XOR2_X1 U12841 ( .A1(\MC_ARK_ARC_1_2/temp5[76] ), .A2(n6387), .Z(
        \MC_ARK_ARC_1_2/buf_output[76] ) );
  XOR2_X1 U12842 ( .A1(\MC_ARK_ARC_1_2/temp3[76] ), .A2(
        \MC_ARK_ARC_1_2/temp4[76] ), .Z(n6387) );
  XOR2_X1 U12843 ( .A1(n6388), .A2(n166), .Z(Ciphertext[103]) );
  XOR2_X1 U12844 ( .A1(\MC_ARK_ARC_1_0/temp1[174] ), .A2(
        \MC_ARK_ARC_1_0/temp2[174] ), .Z(n6389) );
  NAND4_X2 U12845 ( .A1(\SB2_1_14/Component_Function_2/NAND4_in[2] ), .A2(
        n4201), .A3(n1151), .A4(n6390), .ZN(\SB2_1_14/buf_output[2] ) );
  NAND3_X2 U12846 ( .A1(\SB2_1_14/i0[10] ), .A2(\SB2_1_14/i1_5 ), .A3(
        \SB2_1_14/i1[9] ), .ZN(n6390) );
  NAND3_X1 U12847 ( .A1(\SB2_3_12/i0_0 ), .A2(\SB2_3_12/i0[6] ), .A3(
        \SB1_3_14/buf_output[3] ), .ZN(n6391) );
  XOR2_X1 U12848 ( .A1(n6392), .A2(\MC_ARK_ARC_1_1/temp5[97] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[97] ) );
  XOR2_X1 U12849 ( .A1(n6393), .A2(n14), .Z(Ciphertext[128]) );
  NAND4_X2 U12850 ( .A1(n2730), .A2(\SB4_10/Component_Function_2/NAND4_in[0] ), 
        .A3(n1511), .A4(n4554), .ZN(n6393) );
  XOR2_X1 U12851 ( .A1(\RI5[0][187] ), .A2(\RI5[0][181] ), .Z(
        \MC_ARK_ARC_1_0/temp1[187] ) );
  XOR2_X1 U12852 ( .A1(n4374), .A2(n2019), .Z(\MC_ARK_ARC_1_2/buf_output[105] ) );
  NAND3_X1 U12853 ( .A1(\SB4_13/i0_3 ), .A2(\SB4_13/i0[10] ), .A3(
        \SB4_13/i0_4 ), .ZN(\SB4_13/Component_Function_0/NAND4_in[2] ) );
  NOR2_X2 U12854 ( .A1(n6396), .A2(n6395), .ZN(n3653) );
  NAND2_X1 U12855 ( .A1(\SB3_13/Component_Function_2/NAND4_in[3] ), .A2(
        \SB3_13/Component_Function_2/NAND4_in[1] ), .ZN(n6396) );
  NAND3_X2 U12856 ( .A1(\SB2_0_14/i0[8] ), .A2(\SB2_0_14/i0[9] ), .A3(
        \RI3[0][104] ), .ZN(\SB2_0_14/Component_Function_4/NAND4_in[0] ) );
  NAND4_X2 U12857 ( .A1(\SB2_1_20/Component_Function_0/NAND4_in[3] ), .A2(n890), .A3(\SB2_1_20/Component_Function_0/NAND4_in[0] ), .A4(
        \SB2_1_20/Component_Function_0/NAND4_in[1] ), .ZN(
        \SB2_1_20/buf_output[0] ) );
  XOR2_X1 U12858 ( .A1(\MC_ARK_ARC_1_1/temp5[30] ), .A2(n6398), .Z(
        \MC_ARK_ARC_1_1/buf_output[30] ) );
  XOR2_X1 U12859 ( .A1(n2691), .A2(\MC_ARK_ARC_1_1/temp4[30] ), .Z(n6398) );
  NAND3_X1 U12860 ( .A1(\SB1_0_24/i0_3 ), .A2(n266), .A3(\SB1_0_24/i0[8] ), 
        .ZN(\SB1_0_24/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U12861 ( .A1(\SB1_3_17/i0_3 ), .A2(\SB1_3_17/i0[6] ), .A3(
        \SB1_3_17/i1[9] ), .ZN(\SB1_3_17/Component_Function_3/NAND4_in[0] ) );
  NAND3_X1 U12862 ( .A1(\SB4_9/i0[10] ), .A2(\SB4_9/i1_5 ), .A3(\SB4_9/i1[9] ), 
        .ZN(n6399) );
  XOR2_X1 U12863 ( .A1(\MC_ARK_ARC_1_1/temp2[123] ), .A2(
        \MC_ARK_ARC_1_1/temp1[123] ), .Z(\MC_ARK_ARC_1_1/temp5[123] ) );
  XOR2_X1 U12864 ( .A1(n6401), .A2(n6400), .Z(n1977) );
  XOR2_X1 U12865 ( .A1(\MC_ARK_ARC_1_0/temp2[71] ), .A2(n4756), .Z(n6400) );
  XOR2_X1 U12866 ( .A1(n6443), .A2(n2415), .Z(n6401) );
  XOR2_X1 U12867 ( .A1(\MC_ARK_ARC_1_0/temp1[141] ), .A2(n6402), .Z(
        \MC_ARK_ARC_1_0/temp5[141] ) );
  XOR2_X1 U12868 ( .A1(\RI5[0][111] ), .A2(\RI5[0][87] ), .Z(n6402) );
  NAND3_X2 U12869 ( .A1(\SB2_1_16/i0[10] ), .A2(\SB2_1_16/i1[9] ), .A3(
        \SB2_1_16/i1_7 ), .ZN(n6403) );
  NAND3_X2 U12870 ( .A1(\SB3_27/i0[10] ), .A2(\SB3_27/i0[6] ), .A3(
        \SB3_27/i0_3 ), .ZN(n6404) );
  NAND4_X2 U12871 ( .A1(\SB1_0_13/Component_Function_3/NAND4_in[2] ), .A2(
        \SB1_0_13/Component_Function_3/NAND4_in[3] ), .A3(
        \SB1_0_13/Component_Function_3/NAND4_in[0] ), .A4(n6405), .ZN(
        \RI3[0][123] ) );
  NAND4_X2 U12872 ( .A1(n4328), .A2(
        \SB1_3_20/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_3_20/Component_Function_5/NAND4_in[0] ), .A4(n6406), .ZN(
        \SB1_3_20/buf_output[5] ) );
  XOR2_X1 U12873 ( .A1(\MC_ARK_ARC_1_0/temp4[171] ), .A2(n6407), .Z(
        \MC_ARK_ARC_1_0/temp6[171] ) );
  XOR2_X1 U12874 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[81] ), .A2(\RI5[0][45] ), 
        .Z(n6407) );
  NAND3_X1 U12875 ( .A1(\SB1_0_20/i0[10] ), .A2(\SB1_0_20/i1[9] ), .A3(
        \SB1_0_20/i1_7 ), .ZN(\SB1_0_20/Component_Function_3/NAND4_in[2] ) );
  XOR2_X1 U12876 ( .A1(\RI5[2][80] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[56] ), 
        .Z(n6408) );
  XOR2_X1 U12877 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[7] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[43] ), .Z(n6409) );
  XOR2_X1 U12878 ( .A1(\RI5[0][140] ), .A2(\RI5[0][176] ), .Z(n6410) );
  NAND4_X2 U12879 ( .A1(\SB2_0_18/Component_Function_2/NAND4_in[0] ), .A2(
        n3572), .A3(n1638), .A4(n6411), .ZN(\SB2_0_18/buf_output[2] ) );
  NAND3_X1 U12880 ( .A1(\SB3_27/i0[6] ), .A2(\SB3_27/i0_3 ), .A3(n4764), .ZN(
        n6412) );
  NAND4_X2 U12881 ( .A1(n1438), .A2(\SB2_2_8/Component_Function_0/NAND4_in[1] ), .A3(n1439), .A4(n6413), .ZN(\SB2_2_8/buf_output[0] ) );
  NAND2_X1 U12882 ( .A1(\SB2_2_8/i0[9] ), .A2(\SB2_2_8/i0[10] ), .ZN(n6413) );
  NAND4_X2 U12883 ( .A1(\SB2_2_5/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_2_5/Component_Function_0/NAND4_in[0] ), .A3(
        \SB2_2_5/Component_Function_0/NAND4_in[2] ), .A4(n6414), .ZN(
        \SB2_2_5/buf_output[0] ) );
  NAND3_X2 U12884 ( .A1(\SB2_2_5/i0[7] ), .A2(\SB2_2_5/i0[8] ), .A3(
        \SB2_2_5/i0[6] ), .ZN(n6414) );
  XOR2_X1 U12885 ( .A1(n6415), .A2(\MC_ARK_ARC_1_3/temp5[97] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[97] ) );
  XOR2_X1 U12886 ( .A1(\MC_ARK_ARC_1_3/temp3[97] ), .A2(
        \MC_ARK_ARC_1_3/temp4[97] ), .Z(n6415) );
  XOR2_X1 U12887 ( .A1(\MC_ARK_ARC_1_2/temp1[0] ), .A2(
        \MC_ARK_ARC_1_2/temp2[0] ), .Z(\MC_ARK_ARC_1_2/temp5[0] ) );
  XOR2_X1 U12888 ( .A1(\RI5[1][171] ), .A2(n480), .Z(
        \MC_ARK_ARC_1_1/temp4[135] ) );
  NAND4_X2 U12889 ( .A1(\SB1_2_9/Component_Function_3/NAND4_in[0] ), .A2(
        \SB1_2_9/Component_Function_3/NAND4_in[1] ), .A3(n2922), .A4(n2923), 
        .ZN(\SB1_2_9/buf_output[3] ) );
  XOR2_X1 U12890 ( .A1(\RI5[2][143] ), .A2(\RI5[2][119] ), .Z(
        \MC_ARK_ARC_1_2/temp2[173] ) );
  NOR2_X2 U12891 ( .A1(n2241), .A2(n6418), .ZN(\SB2_3_15/i0[7] ) );
  NAND4_X2 U12892 ( .A1(\SB2_0_25/Component_Function_5/NAND4_in[3] ), .A2(
        \SB2_0_25/Component_Function_5/NAND4_in[0] ), .A3(
        \SB2_0_25/Component_Function_5/NAND4_in[1] ), .A4(n6419), .ZN(
        \SB2_0_25/buf_output[5] ) );
  NAND3_X2 U12893 ( .A1(\RI3[0][40] ), .A2(\SB2_0_25/i0_3 ), .A3(
        \SB2_0_25/i1[9] ), .ZN(n6419) );
  XOR2_X1 U12894 ( .A1(n6420), .A2(\MC_ARK_ARC_1_0/temp6[26] ), .Z(
        \MC_ARK_ARC_1_0/buf_output[26] ) );
  XOR2_X1 U12895 ( .A1(\MC_ARK_ARC_1_0/temp1[26] ), .A2(n3168), .Z(n6420) );
  INV_X2 U12896 ( .I(\SB1_2_28/buf_output[2] ), .ZN(\SB2_2_25/i1[9] ) );
  XOR2_X1 U12897 ( .A1(\RI5[1][34] ), .A2(\RI5[1][58] ), .Z(
        \MC_ARK_ARC_1_1/temp2[88] ) );
  NAND3_X1 U12898 ( .A1(\SB3_31/i0[6] ), .A2(\SB3_31/i0[8] ), .A3(
        \SB3_31/i0[7] ), .ZN(\SB3_31/Component_Function_0/NAND4_in[1] ) );
  NAND3_X1 U12899 ( .A1(\SB4_26/i0[9] ), .A2(\SB4_26/i0_3 ), .A3(
        \SB4_26/i0[8] ), .ZN(n6421) );
  XOR2_X1 U12900 ( .A1(\MC_ARK_ARC_1_0/temp5[18] ), .A2(
        \MC_ARK_ARC_1_0/temp6[18] ), .Z(\MC_ARK_ARC_1_0/buf_output[18] ) );
  NAND3_X2 U12901 ( .A1(\SB1_2_25/i0_4 ), .A2(\SB1_2_25/i0_3 ), .A3(
        \SB1_2_25/i1[9] ), .ZN(\SB1_2_25/Component_Function_5/NAND4_in[2] ) );
  NAND3_X2 U12902 ( .A1(\SB1_2_23/i0_4 ), .A2(\SB1_2_23/i1_5 ), .A3(
        \SB1_2_23/i0_0 ), .ZN(\SB1_2_23/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 U12903 ( .A1(\SB2_0_17/i0_0 ), .A2(\SB2_0_17/i1_5 ), .A3(
        \RI3[0][88] ), .ZN(n6504) );
  XOR2_X1 U12904 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[78] ), .A2(\RI5[0][114] ), 
        .Z(\MC_ARK_ARC_1_0/temp3[12] ) );
  XOR2_X1 U12905 ( .A1(\MC_ARK_ARC_1_1/temp2[27] ), .A2(n6422), .Z(
        \MC_ARK_ARC_1_1/temp5[27] ) );
  XOR2_X1 U12906 ( .A1(\RI5[1][21] ), .A2(\RI5[1][27] ), .Z(n6422) );
  XOR2_X1 U12907 ( .A1(\MC_ARK_ARC_1_0/temp5[128] ), .A2(
        \MC_ARK_ARC_1_0/temp6[128] ), .Z(\MC_ARK_ARC_1_0/buf_output[128] ) );
  XOR2_X1 U12908 ( .A1(n2385), .A2(\MC_ARK_ARC_1_3/temp6[65] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[65] ) );
  NAND4_X2 U12909 ( .A1(\SB1_0_12/Component_Function_3/NAND4_in[3] ), .A2(
        \SB1_0_12/Component_Function_3/NAND4_in[1] ), .A3(n3790), .A4(n2655), 
        .ZN(\RI3[0][129] ) );
  NAND4_X2 U12910 ( .A1(\SB1_2_4/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_2_4/Component_Function_5/NAND4_in[1] ), .A3(n6492), .A4(
        \SB1_2_4/Component_Function_5/NAND4_in[0] ), .ZN(
        \SB1_2_4/buf_output[5] ) );
  NAND4_X2 U12911 ( .A1(\SB1_0_0/Component_Function_1/NAND4_in[2] ), .A2(
        \SB1_0_0/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_0/Component_Function_1/NAND4_in[3] ), .A4(
        \SB1_0_0/Component_Function_1/NAND4_in[0] ), .ZN(
        \SB1_0_0/buf_output[1] ) );
  NAND4_X2 U12912 ( .A1(\SB3_21/Component_Function_4/NAND4_in[3] ), .A2(
        \SB3_21/Component_Function_4/NAND4_in[0] ), .A3(n6459), .A4(
        \SB3_21/Component_Function_4/NAND4_in[1] ), .ZN(\SB3_21/buf_output[4] ) );
  XOR2_X1 U12913 ( .A1(\RI5[0][122] ), .A2(\RI5[0][128] ), .Z(
        \MC_ARK_ARC_1_0/temp1[128] ) );
  NAND3_X1 U12914 ( .A1(\SB1_3_17/i0[8] ), .A2(\SB1_3_17/i0_3 ), .A3(
        \SB1_3_17/i1_7 ), .ZN(\SB1_3_17/Component_Function_1/NAND4_in[1] ) );
  XOR2_X1 U12915 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[0] ), .A2(
        \MC_ARK_ARC_1_2/buf_datainput[156] ), .Z(\MC_ARK_ARC_1_2/temp3[90] )
         );
  NAND3_X1 U12916 ( .A1(\SB4_20/i0_4 ), .A2(\SB4_20/i1_7 ), .A3(\SB4_20/i0[8] ), .ZN(\SB4_20/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U12917 ( .A1(\SB1_2_10/Component_Function_1/NAND4_in[1] ), .A2(
        \SB1_2_10/Component_Function_1/NAND4_in[3] ), .A3(
        \SB1_2_10/Component_Function_1/NAND4_in[0] ), .A4(n6425), .ZN(
        \SB1_2_10/buf_output[1] ) );
  NAND3_X2 U12918 ( .A1(\SB1_2_10/i0[9] ), .A2(\SB1_2_10/i0[6] ), .A3(
        \SB1_2_10/i1_5 ), .ZN(n6425) );
  INV_X2 U12919 ( .I(\SB1_0_14/buf_output[2] ), .ZN(\SB2_0_11/i1[9] ) );
  NAND4_X2 U12920 ( .A1(\SB1_0_14/Component_Function_2/NAND4_in[0] ), .A2(
        \SB1_0_14/Component_Function_2/NAND4_in[1] ), .A3(n1105), .A4(
        \SB1_0_14/Component_Function_2/NAND4_in[3] ), .ZN(
        \SB1_0_14/buf_output[2] ) );
  NAND3_X1 U12921 ( .A1(\SB4_10/i0_4 ), .A2(\SB3_13/buf_output[2] ), .A3(
        \SB4_10/i0_3 ), .ZN(n6428) );
  NAND3_X1 U12922 ( .A1(\SB4_11/i0_0 ), .A2(\SB3_12/buf_output[4] ), .A3(n3684), .ZN(\SB4_11/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 U12923 ( .A1(\SB2_1_28/i0_3 ), .A2(\SB2_1_28/i0[9] ), .A3(
        \SB2_1_28/i0[8] ), .ZN(n6429) );
  XOR2_X1 U12924 ( .A1(\MC_ARK_ARC_1_3/temp4[70] ), .A2(n6430), .Z(
        \MC_ARK_ARC_1_3/temp6[70] ) );
  XOR2_X1 U12925 ( .A1(\RI5[3][136] ), .A2(\RI5[3][172] ), .Z(n6430) );
  NAND3_X1 U12926 ( .A1(\SB1_3_4/i0[10] ), .A2(\SB1_3_4/i1_5 ), .A3(
        \SB1_3_4/i1[9] ), .ZN(n6432) );
  NAND3_X1 U12927 ( .A1(\SB3_11/i0_0 ), .A2(\SB3_11/i3[0] ), .A3(\SB3_11/i1_7 ), .ZN(\SB3_11/Component_Function_4/NAND4_in[1] ) );
  NAND4_X2 U12928 ( .A1(n1884), .A2(n3353), .A3(
        \SB2_2_22/Component_Function_5/NAND4_in[3] ), .A4(n6433), .ZN(
        \SB2_2_22/buf_output[5] ) );
  XOR2_X1 U12929 ( .A1(\RI5[1][115] ), .A2(\RI5[1][109] ), .Z(n3744) );
  XOR2_X1 U12930 ( .A1(\RI5[3][0] ), .A2(\RI5[3][24] ), .Z(
        \MC_ARK_ARC_1_3/temp2[54] ) );
  NAND3_X1 U12931 ( .A1(\SB2_0_2/i0_3 ), .A2(\RI3[0][176] ), .A3(
        \SB2_0_2/i0[7] ), .ZN(\SB2_0_2/Component_Function_0/NAND4_in[3] ) );
  NOR2_X2 U12932 ( .A1(n6435), .A2(n6434), .ZN(\SB2_0_2/i0[7] ) );
  NAND2_X2 U12933 ( .A1(\SB1_0_3/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_0_3/Component_Function_4/NAND4_in[2] ), .ZN(n6434) );
  XOR2_X1 U12934 ( .A1(n6437), .A2(\MC_ARK_ARC_1_1/temp5[43] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[43] ) );
  XOR2_X1 U12935 ( .A1(\MC_ARK_ARC_1_1/temp3[43] ), .A2(
        \MC_ARK_ARC_1_1/temp4[43] ), .Z(n6437) );
  NAND3_X1 U12936 ( .A1(\SB3_2/i0_4 ), .A2(\SB3_2/i1_7 ), .A3(\SB3_2/i0[8] ), 
        .ZN(n3462) );
  NAND3_X1 U12937 ( .A1(\SB2_0_19/i0[6] ), .A2(\SB2_0_19/i0[8] ), .A3(
        \SB2_0_19/i0[7] ), .ZN(\SB2_0_19/Component_Function_0/NAND4_in[1] ) );
  NOR2_X2 U12938 ( .A1(n6439), .A2(n6438), .ZN(\SB2_0_19/i0[7] ) );
  XOR2_X1 U12939 ( .A1(\SB2_1_27/buf_output[4] ), .A2(\SB2_1_26/buf_output[4] ), .Z(\MC_ARK_ARC_1_1/temp1[40] ) );
  NAND4_X2 U12940 ( .A1(\SB2_1_28/Component_Function_3/NAND4_in[2] ), .A2(
        \SB2_1_28/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_1_28/Component_Function_3/NAND4_in[0] ), .A4(n6440), .ZN(
        \SB2_1_28/buf_output[3] ) );
  XOR2_X1 U12941 ( .A1(\MC_ARK_ARC_1_0/temp2[86] ), .A2(n6441), .Z(n2094) );
  XOR2_X1 U12942 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[86] ), .A2(\RI5[0][80] ), 
        .Z(n6441) );
  XOR2_X1 U12943 ( .A1(\RI5[1][17] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[185] ), 
        .Z(n6442) );
  INV_X2 U12944 ( .I(\RI3[0][183] ), .ZN(\SB2_0_1/i0[8] ) );
  XOR2_X1 U12945 ( .A1(\RI5[2][147] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[153] ), .Z(\MC_ARK_ARC_1_2/temp1[153] ) );
  NAND4_X2 U12946 ( .A1(\SB2_1_17/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_1_17/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_1_17/Component_Function_2/NAND4_in[3] ), .A4(n6445), .ZN(
        \SB2_1_17/buf_output[2] ) );
  NAND3_X2 U12947 ( .A1(\SB2_1_17/i0_3 ), .A2(\SB2_1_17/i0[10] ), .A3(
        \SB2_1_17/i0[6] ), .ZN(n6445) );
  NAND4_X2 U12948 ( .A1(\SB1_2_22/Component_Function_3/NAND4_in[1] ), .A2(
        \SB1_2_22/Component_Function_3/NAND4_in[0] ), .A3(n1496), .A4(
        \SB1_2_22/Component_Function_3/NAND4_in[3] ), .ZN(
        \SB1_2_22/buf_output[3] ) );
  XOR2_X1 U12949 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[81] ), .A2(\RI5[2][57] ), 
        .Z(n4190) );
  NAND3_X1 U12950 ( .A1(\SB3_25/i1_5 ), .A2(\SB3_25/i3[0] ), .A3(
        \SB3_25/i0[8] ), .ZN(n6446) );
  XOR2_X1 U12951 ( .A1(\MC_ARK_ARC_1_1/temp2[33] ), .A2(
        \MC_ARK_ARC_1_1/temp3[33] ), .Z(n3870) );
  INV_X2 U12952 ( .I(\SB1_1_2/buf_output[2] ), .ZN(\SB2_1_31/i1[9] ) );
  XOR2_X1 U12953 ( .A1(n6447), .A2(n2669), .Z(\MC_ARK_ARC_1_0/buf_output[34] )
         );
  XOR2_X1 U12954 ( .A1(\MC_ARK_ARC_1_0/temp2[34] ), .A2(
        \MC_ARK_ARC_1_0/temp1[34] ), .Z(n6447) );
  XOR2_X1 U12955 ( .A1(\RI5[2][168] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[162] ), .Z(\MC_ARK_ARC_1_2/temp1[168] ) );
  INV_X1 U12956 ( .I(\SB3_25/buf_output[5] ), .ZN(\SB4_25/i1_5 ) );
  NAND4_X2 U12957 ( .A1(\SB3_25/Component_Function_5/NAND4_in[1] ), .A2(
        \SB3_25/Component_Function_5/NAND4_in[3] ), .A3(n2850), .A4(
        \SB3_25/Component_Function_5/NAND4_in[0] ), .ZN(\SB3_25/buf_output[5] ) );
  XOR2_X1 U12958 ( .A1(n4532), .A2(\MC_ARK_ARC_1_3/temp4[113] ), .Z(
        \MC_ARK_ARC_1_3/temp6[113] ) );
  NAND3_X1 U12959 ( .A1(n5511), .A2(n5489), .A3(\SB2_3_28/i0[6] ), .ZN(
        \SB2_3_28/Component_Function_5/NAND4_in[1] ) );
  NAND3_X2 U12960 ( .A1(\SB2_2_26/i0[6] ), .A2(\SB2_2_26/i0_4 ), .A3(
        \SB2_2_26/i0[9] ), .ZN(n6448) );
  NAND3_X1 U12961 ( .A1(\SB4_28/i0_0 ), .A2(\SB4_28/i0_3 ), .A3(\SB4_28/i0[7] ), .ZN(n1703) );
  NAND4_X2 U12962 ( .A1(\SB1_1_7/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_1_7/Component_Function_1/NAND4_in[0] ), .A3(n3415), .A4(
        \SB1_1_7/Component_Function_1/NAND4_in[1] ), .ZN(
        \SB1_1_7/buf_output[1] ) );
  XOR2_X1 U12963 ( .A1(n6450), .A2(n6449), .Z(\MC_ARK_ARC_1_2/temp6[72] ) );
  XOR2_X1 U12964 ( .A1(\RI5[2][174] ), .A2(n553), .Z(n6449) );
  XOR2_X1 U12965 ( .A1(\RI5[2][138] ), .A2(\RI5[2][108] ), .Z(n6450) );
  XOR2_X1 U12966 ( .A1(\MC_ARK_ARC_1_2/temp2[144] ), .A2(n6451), .Z(
        \MC_ARK_ARC_1_2/temp5[144] ) );
  XOR2_X1 U12967 ( .A1(\RI5[2][138] ), .A2(\RI5[2][144] ), .Z(n6451) );
  XOR2_X1 U12968 ( .A1(\MC_ARK_ARC_1_3/temp2[3] ), .A2(n6452), .Z(
        \MC_ARK_ARC_1_3/temp5[3] ) );
  XOR2_X1 U12969 ( .A1(\RI5[3][189] ), .A2(\RI5[3][3] ), .Z(n6452) );
  XOR2_X1 U12970 ( .A1(n6453), .A2(\MC_ARK_ARC_1_3/temp6[1] ), .Z(
        \MC_ARK_ARC_1_3/buf_output[1] ) );
  INV_X1 U12971 ( .I(\SB1_3_7/buf_output[1] ), .ZN(\SB2_3_3/i1_7 ) );
  XOR2_X1 U12972 ( .A1(\MC_ARK_ARC_1_0/temp3[147] ), .A2(
        \MC_ARK_ARC_1_0/temp4[147] ), .Z(\MC_ARK_ARC_1_0/temp6[147] ) );
  XOR2_X1 U12973 ( .A1(\MC_ARK_ARC_1_0/buf_datainput[138] ), .A2(
        \MC_ARK_ARC_1_0/buf_datainput[144] ), .Z(\MC_ARK_ARC_1_0/temp1[144] )
         );
  NAND4_X2 U12974 ( .A1(\SB3_25/Component_Function_1/NAND4_in[2] ), .A2(
        \SB3_25/Component_Function_1/NAND4_in[1] ), .A3(
        \SB3_25/Component_Function_1/NAND4_in[0] ), .A4(n6454), .ZN(
        \SB3_25/buf_output[1] ) );
  NAND3_X1 U12975 ( .A1(\SB3_25/i0_4 ), .A2(\SB3_25/i1_7 ), .A3(\SB3_25/i0[8] ), .ZN(n6454) );
  NAND3_X2 U12976 ( .A1(\SB1_3_31/i0_3 ), .A2(\SB1_3_31/i0_0 ), .A3(
        \SB1_3_31/i0_4 ), .ZN(n6456) );
  XOR2_X1 U12977 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[131] ), .A2(\RI5[2][107] ), .Z(n6457) );
  NAND3_X2 U12978 ( .A1(\SB1_3_13/i0_3 ), .A2(\SB1_3_13/i0_4 ), .A3(
        \SB1_3_13/i1[9] ), .ZN(\SB1_3_13/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U12979 ( .A1(\MC_ARK_ARC_1_3/temp5[112] ), .A2(n6460), .Z(
        \MC_ARK_ARC_1_3/buf_output[112] ) );
  XOR2_X1 U12980 ( .A1(\MC_ARK_ARC_1_3/temp3[112] ), .A2(
        \MC_ARK_ARC_1_3/temp4[112] ), .Z(n6460) );
  XOR2_X1 U12981 ( .A1(\RI5[0][65] ), .A2(\RI5[0][71] ), .Z(n2415) );
  INV_X1 U12982 ( .I(n413), .ZN(\SB1_0_23/i1_5 ) );
  XOR2_X1 U12983 ( .A1(n3541), .A2(n6464), .Z(\MC_ARK_ARC_1_1/buf_output[190] ) );
  XOR2_X1 U12984 ( .A1(\MC_ARK_ARC_1_1/temp1[190] ), .A2(
        \MC_ARK_ARC_1_1/temp2[190] ), .Z(n6464) );
  NAND3_X2 U12985 ( .A1(\SB3_11/i0_0 ), .A2(\SB3_11/i0[6] ), .A3(
        \SB3_11/i0[10] ), .ZN(n3999) );
  XOR2_X1 U12986 ( .A1(\RI5[0][15] ), .A2(\RI5[0][183] ), .Z(
        \MC_ARK_ARC_1_0/temp2[45] ) );
  NAND3_X2 U12987 ( .A1(\SB1_3_31/i0_3 ), .A2(\SB1_3_31/i0[10] ), .A3(
        \SB1_3_31/i0[9] ), .ZN(n6466) );
  NAND4_X2 U12988 ( .A1(\SB2_2_17/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_2_17/Component_Function_4/NAND4_in[1] ), .A3(n1278), .A4(n6467), 
        .ZN(\SB2_2_17/buf_output[4] ) );
  XOR2_X1 U12989 ( .A1(n6468), .A2(\MC_ARK_ARC_1_2/temp1[91] ), .Z(
        \MC_ARK_ARC_1_2/temp5[91] ) );
  XOR2_X1 U12990 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[61] ), .A2(\RI5[2][37] ), 
        .Z(n6468) );
  XOR2_X1 U12991 ( .A1(n4524), .A2(n6469), .Z(\MC_ARK_ARC_1_1/buf_output[70] )
         );
  XOR2_X1 U12992 ( .A1(\MC_ARK_ARC_1_1/temp4[70] ), .A2(
        \MC_ARK_ARC_1_1/temp3[70] ), .Z(n6469) );
  NAND3_X1 U12993 ( .A1(n5511), .A2(\SB2_3_28/i0_3 ), .A3(\SB2_3_28/i0[9] ), 
        .ZN(\SB2_3_28/Component_Function_4/NAND4_in[2] ) );
  NAND4_X2 U12994 ( .A1(\SB2_0_13/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_0_13/Component_Function_3/NAND4_in[2] ), .A3(
        \SB2_0_13/Component_Function_3/NAND4_in[3] ), .A4(
        \SB2_0_13/Component_Function_3/NAND4_in[1] ), .ZN(
        \SB2_0_13/buf_output[3] ) );
  XOR2_X1 U12995 ( .A1(\MC_ARK_ARC_1_1/temp4[159] ), .A2(n3050), .Z(n6470) );
  NAND3_X1 U12996 ( .A1(\SB1_3_26/i0[6] ), .A2(\SB1_3_26/i0_3 ), .A3(
        \SB1_3_26/i0[10] ), .ZN(\SB1_3_26/Component_Function_2/NAND4_in[1] )
         );
  XOR2_X1 U12997 ( .A1(n1023), .A2(n2389), .Z(\MC_ARK_ARC_1_2/buf_output[31] )
         );
  NOR2_X2 U12998 ( .A1(n1659), .A2(n1660), .ZN(n722) );
  XOR2_X1 U12999 ( .A1(n6471), .A2(n183), .Z(Ciphertext[176]) );
  XOR2_X1 U13000 ( .A1(\MC_ARK_ARC_1_2/temp6[41] ), .A2(n6472), .Z(
        \RI1[3][41] ) );
  XOR2_X1 U13001 ( .A1(\MC_ARK_ARC_1_2/temp2[41] ), .A2(
        \MC_ARK_ARC_1_2/temp1[41] ), .Z(n6472) );
  NAND3_X1 U13002 ( .A1(\SB2_2_26/i0[6] ), .A2(\SB2_2_26/i1_5 ), .A3(
        \SB2_2_26/i0[9] ), .ZN(\SB2_2_26/Component_Function_1/NAND4_in[2] ) );
  XOR2_X1 U13003 ( .A1(\MC_ARK_ARC_1_0/temp1[166] ), .A2(
        \MC_ARK_ARC_1_0/temp2[166] ), .Z(\MC_ARK_ARC_1_0/temp5[166] ) );
  NAND4_X2 U13004 ( .A1(\SB2_0_14/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_0_14/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_0_14/Component_Function_4/NAND4_in[3] ), .A4(n6473), .ZN(
        \SB2_0_14/buf_output[4] ) );
  NAND3_X2 U13005 ( .A1(\SB2_2_20/i0_3 ), .A2(\SB2_2_20/i0_0 ), .A3(
        \SB2_2_20/i0_4 ), .ZN(n6475) );
  XOR2_X1 U13006 ( .A1(n6476), .A2(\MC_ARK_ARC_1_1/temp4[138] ), .Z(
        \MC_ARK_ARC_1_1/temp6[138] ) );
  XOR2_X1 U13007 ( .A1(\RI5[1][12] ), .A2(\RI5[1][48] ), .Z(n6476) );
  XOR2_X1 U13008 ( .A1(\RI5[1][182] ), .A2(n133), .Z(n6477) );
  NAND4_X2 U13009 ( .A1(\SB2_2_30/Component_Function_0/NAND4_in[3] ), .A2(
        \SB2_2_30/Component_Function_0/NAND4_in[1] ), .A3(
        \SB2_2_30/Component_Function_0/NAND4_in[0] ), .A4(n6478), .ZN(
        \SB2_2_30/buf_output[0] ) );
  INV_X2 U13010 ( .I(\SB1_1_1/buf_output[2] ), .ZN(\SB2_1_30/i1[9] ) );
  NAND4_X2 U13011 ( .A1(\SB1_1_1/Component_Function_2/NAND4_in[0] ), .A2(n3386), .A3(\SB1_1_1/Component_Function_2/NAND4_in[2] ), .A4(n1906), .ZN(
        \SB1_1_1/buf_output[2] ) );
  NAND3_X2 U13012 ( .A1(\SB2_1_13/i0[10] ), .A2(\SB2_1_13/i0_3 ), .A3(
        \SB2_1_13/i0[6] ), .ZN(\SB2_1_13/Component_Function_2/NAND4_in[1] ) );
  NAND3_X2 U13013 ( .A1(\SB1_0_4/i0[10] ), .A2(\SB1_0_4/i1[9] ), .A3(
        \SB1_0_4/i1_7 ), .ZN(n6479) );
  XOR2_X1 U13014 ( .A1(n6480), .A2(\MC_ARK_ARC_1_1/temp6[85] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[85] ) );
  XOR2_X1 U13015 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[116] ), .A2(\RI5[2][110] ), .Z(n6481) );
  XOR2_X1 U13016 ( .A1(\RI5[2][62] ), .A2(\MC_ARK_ARC_1_2/buf_datainput[38] ), 
        .Z(\MC_ARK_ARC_1_2/temp2[92] ) );
  XOR2_X1 U13017 ( .A1(\RI5[2][167] ), .A2(\RI5[2][143] ), .Z(n3196) );
  XOR2_X1 U13018 ( .A1(n6483), .A2(\MC_ARK_ARC_1_1/temp5[133] ), .Z(
        \MC_ARK_ARC_1_1/buf_output[133] ) );
  XOR2_X1 U13019 ( .A1(\MC_ARK_ARC_1_1/temp3[133] ), .A2(
        \MC_ARK_ARC_1_1/temp4[133] ), .Z(n6483) );
  NAND3_X2 U13020 ( .A1(n390), .A2(\SB1_0_7/i0_0 ), .A3(\SB1_0_7/i1_5 ), .ZN(
        \SB1_0_7/Component_Function_2/NAND4_in[3] ) );
  NAND3_X2 U13021 ( .A1(\SB2_0_7/i0_3 ), .A2(\SB2_0_7/i0[9] ), .A3(
        \SB2_0_7/i0[8] ), .ZN(n6484) );
  NAND3_X1 U13022 ( .A1(\SB4_28/i0[6] ), .A2(\SB4_28/i0[8] ), .A3(
        \SB4_28/i0[7] ), .ZN(n6485) );
  NAND3_X2 U13023 ( .A1(\SB2_3_31/i0_3 ), .A2(\SB2_3_31/i0[8] ), .A3(
        \SB2_3_31/i0[9] ), .ZN(\SB2_3_31/Component_Function_2/NAND4_in[2] ) );
  NAND3_X1 U13024 ( .A1(\SB3_10/i0[9] ), .A2(\SB3_10/i0_4 ), .A3(
        \SB3_10/i0[6] ), .ZN(n6486) );
  XOR2_X1 U13025 ( .A1(n4067), .A2(n6487), .Z(n4183) );
  XOR2_X1 U13026 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[99] ), .A2(\RI5[2][93] ), 
        .Z(n6487) );
  NAND2_X2 U13027 ( .A1(\SB2_2_16/i0_0 ), .A2(\SB2_2_16/i3[0] ), .ZN(n6488) );
  NAND4_X2 U13028 ( .A1(n1683), .A2(
        \SB2_3_19/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_3_19/Component_Function_2/NAND4_in[0] ), .A4(n6489), .ZN(
        \SB2_3_19/buf_output[2] ) );
  NAND3_X1 U13029 ( .A1(\SB4_4/i0[10] ), .A2(\SB4_4/i0_3 ), .A3(\SB4_4/i0[6] ), 
        .ZN(n6490) );
  NAND3_X2 U13030 ( .A1(\SB1_1_13/i0[10] ), .A2(\SB1_1_13/i1[9] ), .A3(
        \SB1_1_13/i1_7 ), .ZN(\SB1_1_13/Component_Function_3/NAND4_in[2] ) );
  NAND3_X2 U13031 ( .A1(\SB1_2_4/i0[6] ), .A2(\SB1_2_4/i0_4 ), .A3(
        \SB1_2_4/i0[9] ), .ZN(n6492) );
  XOR2_X1 U13032 ( .A1(n6496), .A2(n6495), .Z(\MC_ARK_ARC_1_1/buf_output[165] ) );
  XOR2_X1 U13033 ( .A1(\MC_ARK_ARC_1_1/temp3[165] ), .A2(
        \MC_ARK_ARC_1_1/temp4[165] ), .Z(n6495) );
  NAND4_X2 U13034 ( .A1(\SB2_2_18/Component_Function_5/NAND4_in[2] ), .A2(
        n4039), .A3(\SB2_2_18/Component_Function_5/NAND4_in[0] ), .A4(n6497), 
        .ZN(\SB2_2_18/buf_output[5] ) );
  NAND3_X2 U13035 ( .A1(\SB2_2_18/i0[6] ), .A2(\SB2_2_18/i0[10] ), .A3(
        \SB2_2_18/i0_0 ), .ZN(n6497) );
  NAND4_X2 U13036 ( .A1(\SB1_0_18/Component_Function_1/NAND4_in[3] ), .A2(
        \SB1_0_18/Component_Function_1/NAND4_in[1] ), .A3(
        \SB1_0_18/Component_Function_1/NAND4_in[2] ), .A4(n6499), .ZN(
        \RI3[0][103] ) );
  NAND3_X1 U13037 ( .A1(\SB2_1_1/i1_7 ), .A2(\SB2_1_1/i0[8] ), .A3(
        \SB1_1_2/buf_output[4] ), .ZN(n4322) );
  INV_X4 U13038 ( .I(\SB2_0_30/i0[7] ), .ZN(\RI3[0][10] ) );
  NAND3_X1 U13039 ( .A1(\SB2_0_30/i0_0 ), .A2(\SB2_0_30/i0_3 ), .A3(
        \SB2_0_30/i0[7] ), .ZN(\SB2_0_30/Component_Function_0/NAND4_in[3] ) );
  NOR2_X2 U13040 ( .A1(n6501), .A2(n6500), .ZN(\SB2_0_30/i0[7] ) );
  NAND2_X2 U13041 ( .A1(\SB1_0_31/Component_Function_4/NAND4_in[3] ), .A2(
        \SB1_0_31/Component_Function_4/NAND4_in[2] ), .ZN(n6500) );
  AND2_X1 U13042 ( .A1(\SB1_0_3/Component_Function_3/NAND4_in[3] ), .A2(n1646), 
        .Z(n6502) );
  XOR2_X1 U13043 ( .A1(\MC_ARK_ARC_1_1/temp6[178] ), .A2(n6503), .Z(
        \MC_ARK_ARC_1_1/buf_output[178] ) );
  XOR2_X1 U13044 ( .A1(\MC_ARK_ARC_1_1/temp2[178] ), .A2(
        \MC_ARK_ARC_1_1/temp1[178] ), .Z(n6503) );
  INV_X2 U13045 ( .I(\SB1_1_17/buf_output[2] ), .ZN(\SB2_1_14/i1[9] ) );
  NAND4_X2 U13046 ( .A1(\SB1_1_17/Component_Function_2/NAND4_in[2] ), .A2(
        \SB1_1_17/Component_Function_2/NAND4_in[0] ), .A3(n1984), .A4(n2013), 
        .ZN(\SB1_1_17/buf_output[2] ) );
  NAND4_X2 U13047 ( .A1(\SB2_0_17/Component_Function_2/NAND4_in[0] ), .A2(
        \SB2_0_17/Component_Function_2/NAND4_in[2] ), .A3(
        \SB2_0_17/Component_Function_2/NAND4_in[1] ), .A4(n6504), .ZN(
        \SB2_0_17/buf_output[2] ) );
  XOR2_X1 U13048 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[101] ), .A2(
        \MC_ARK_ARC_1_1/buf_datainput[95] ), .Z(n6505) );
  NAND3_X1 U13049 ( .A1(\SB1_0_20/i0[10] ), .A2(\SB1_0_20/i0[9] ), .A3(
        \SB1_0_20/i0_3 ), .ZN(\SB1_0_20/Component_Function_4/NAND4_in[2] ) );
  XOR2_X1 U13050 ( .A1(\MC_ARK_ARC_1_0/temp5[130] ), .A2(
        \MC_ARK_ARC_1_0/temp6[130] ), .Z(\MC_ARK_ARC_1_0/buf_output[130] ) );
  NAND3_X2 U13051 ( .A1(\SB3_31/i0_3 ), .A2(\SB3_31/i1[9] ), .A3(\SB3_31/i0_4 ), .ZN(\SB3_31/Component_Function_5/NAND4_in[2] ) );
  XOR2_X1 U13052 ( .A1(\RI5[3][11] ), .A2(\MC_ARK_ARC_1_3/buf_datainput[17] ), 
        .Z(\MC_ARK_ARC_1_3/temp1[17] ) );
  XOR2_X1 U13053 ( .A1(\MC_ARK_ARC_1_3/temp5[122] ), .A2(n6506), .Z(
        \MC_ARK_ARC_1_3/buf_output[122] ) );
  XOR2_X1 U13054 ( .A1(\MC_ARK_ARC_1_3/temp3[122] ), .A2(
        \MC_ARK_ARC_1_3/temp4[122] ), .Z(n6506) );
  NAND3_X1 U13055 ( .A1(\SB3_29/i0_3 ), .A2(\SB3_29/i0_4 ), .A3(\SB3_29/i1[9] ), .ZN(n4426) );
  XOR2_X1 U13056 ( .A1(\MC_ARK_ARC_1_1/temp1[52] ), .A2(n6507), .Z(
        \MC_ARK_ARC_1_1/temp5[52] ) );
  XOR2_X1 U13057 ( .A1(\RI5[1][190] ), .A2(\MC_ARK_ARC_1_1/buf_datainput[22] ), 
        .Z(n6507) );
  NAND3_X2 U13058 ( .A1(\SB2_2_21/i0[8] ), .A2(\SB2_2_21/i1_5 ), .A3(
        \SB2_2_21/i3[0] ), .ZN(\SB2_2_21/Component_Function_3/NAND4_in[3] ) );
  XOR2_X1 U13059 ( .A1(\MC_ARK_ARC_1_2/buf_datainput[185] ), .A2(\RI5[2][179] ), .Z(n6508) );
  NAND3_X1 U13060 ( .A1(\SB2_0_29/i0_4 ), .A2(\SB2_0_29/i1[9] ), .A3(
        \SB2_0_29/i1_5 ), .ZN(\SB2_0_29/Component_Function_4/NAND4_in[3] ) );
  XOR2_X1 U13061 ( .A1(\MC_ARK_ARC_1_0/temp5[28] ), .A2(n1746), .Z(
        \MC_ARK_ARC_1_0/buf_output[28] ) );
  NAND2_X1 U13062 ( .A1(\SB3_0/i3[0] ), .A2(\SB3_0/i0_0 ), .ZN(n6510) );
  AND2_X1 U13063 ( .A1(n4098), .A2(\SB1_3_17/Component_Function_0/NAND4_in[0] ), .Z(n6513) );
  XOR2_X1 U13064 ( .A1(n2726), .A2(n2727), .Z(n3654) );
  XOR2_X1 U13065 ( .A1(\MC_ARK_ARC_1_3/temp2[146] ), .A2(
        \MC_ARK_ARC_1_3/temp4[146] ), .Z(n2726) );
  INV_X2 U13066 ( .I(\SB1_1_6/buf_output[2] ), .ZN(\SB2_1_3/i1[9] ) );
  NAND3_X1 U13067 ( .A1(\SB4_12/i0[10] ), .A2(\SB4_12/i1_7 ), .A3(
        \SB4_12/i1[9] ), .ZN(n6515) );
  XOR2_X1 U13068 ( .A1(\RI5[0][182] ), .A2(\RI5[0][26] ), .Z(n6516) );
  NAND4_X2 U13069 ( .A1(\SB2_2_12/Component_Function_4/NAND4_in[3] ), .A2(
        \SB2_2_12/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_2_12/Component_Function_4/NAND4_in[0] ), .A4(n6517), .ZN(
        \SB2_2_12/buf_output[4] ) );
  NAND3_X1 U13070 ( .A1(\RI3[0][40] ), .A2(\SB2_0_25/i1[9] ), .A3(
        \SB2_0_25/i1_5 ), .ZN(\SB2_0_25/Component_Function_4/NAND4_in[3] ) );
  NAND4_X2 U13071 ( .A1(\SB3_25/Component_Function_4/NAND4_in[2] ), .A2(
        \SB3_25/Component_Function_4/NAND4_in[0] ), .A3(
        \SB3_25/Component_Function_4/NAND4_in[1] ), .A4(n6519), .ZN(
        \SB3_25/buf_output[4] ) );
  NAND3_X1 U13072 ( .A1(\SB3_25/i0_4 ), .A2(\SB3_25/i1[9] ), .A3(\SB3_25/i1_5 ), .ZN(n6519) );
  XOR2_X1 U13073 ( .A1(\MC_ARK_ARC_1_2/temp5[56] ), .A2(n6521), .Z(
        \MC_ARK_ARC_1_2/buf_output[56] ) );
  XOR2_X1 U13074 ( .A1(n2983), .A2(\MC_ARK_ARC_1_2/temp4[56] ), .Z(n6521) );
  NAND4_X2 U13075 ( .A1(n1548), .A2(n1549), .A3(
        \SB1_0_7/Component_Function_0/NAND4_in[1] ), .A4(
        \SB1_0_7/Component_Function_0/NAND4_in[0] ), .ZN(
        \SB1_0_7/buf_output[0] ) );
  XOR2_X1 U13076 ( .A1(n2388), .A2(n6522), .Z(\MC_ARK_ARC_1_1/buf_output[91] )
         );
  XOR2_X1 U13077 ( .A1(\MC_ARK_ARC_1_1/temp1[91] ), .A2(n1628), .Z(n6522) );
  XOR2_X1 U13078 ( .A1(n6523), .A2(n228), .Z(Ciphertext[45]) );
  NAND4_X2 U13079 ( .A1(\SB4_24/Component_Function_3/NAND4_in[1] ), .A2(
        \SB4_24/Component_Function_3/NAND4_in[3] ), .A3(
        \SB4_24/Component_Function_3/NAND4_in[2] ), .A4(
        \SB4_24/Component_Function_3/NAND4_in[0] ), .ZN(n6523) );
  NAND3_X1 U13080 ( .A1(\SB2_1_0/i0[6] ), .A2(\SB2_1_0/i0[7] ), .A3(
        \SB2_1_0/i0[8] ), .ZN(\SB2_1_0/Component_Function_0/NAND4_in[1] ) );
  NOR2_X2 U13081 ( .A1(n6525), .A2(n6524), .ZN(\SB2_1_0/i0[7] ) );
  NAND2_X2 U13082 ( .A1(n4757), .A2(n2256), .ZN(\SB2_1_15/i0_4 ) );
  NAND4_X2 U13083 ( .A1(\SB2_3_27/Component_Function_4/NAND4_in[0] ), .A2(
        \SB2_3_27/Component_Function_4/NAND4_in[1] ), .A3(
        \SB2_3_27/Component_Function_4/NAND4_in[3] ), .A4(n6526), .ZN(
        \SB2_3_27/buf_output[4] ) );
  XOR2_X1 U13084 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[53] ), .A2(\RI5[3][59] ), 
        .Z(n1522) );
  XOR2_X1 U13085 ( .A1(\MC_ARK_ARC_1_1/buf_datainput[163] ), .A2(n237), .Z(
        \MC_ARK_ARC_1_1/temp4[127] ) );
  XOR2_X1 U13086 ( .A1(n618), .A2(\MC_ARK_ARC_1_0/temp4[141] ), .Z(n6527) );
  NAND2_X2 U13087 ( .A1(n6539), .A2(n2282), .ZN(\SB2_1_3/i0_4 ) );
  NAND3_X2 U13088 ( .A1(\SB1_1_22/i0[6] ), .A2(\SB1_1_22/i0[10] ), .A3(
        \SB1_1_22/i0_0 ), .ZN(n6528) );
  INV_X2 U13089 ( .I(\SB1_3_30/buf_output[5] ), .ZN(\SB2_3_30/i1_5 ) );
  XOR2_X1 U13090 ( .A1(\RI5[0][57] ), .A2(\MC_ARK_ARC_1_0/buf_datainput[51] ), 
        .Z(\MC_ARK_ARC_1_0/temp1[57] ) );
  XOR2_X1 U13091 ( .A1(n6531), .A2(\MC_ARK_ARC_1_2/temp6[148] ), .Z(
        \MC_ARK_ARC_1_2/buf_output[148] ) );
  XOR2_X1 U13092 ( .A1(\MC_ARK_ARC_1_2/temp1[148] ), .A2(
        \MC_ARK_ARC_1_2/temp2[148] ), .Z(n6531) );
  INV_X2 U13093 ( .I(\SB1_2_25/buf_output[2] ), .ZN(\SB2_2_22/i1[9] ) );
  NAND4_X2 U13094 ( .A1(\SB2_2_3/Component_Function_3/NAND4_in[0] ), .A2(
        \SB2_2_3/Component_Function_3/NAND4_in[1] ), .A3(
        \SB2_2_3/Component_Function_3/NAND4_in[3] ), .A4(n6532), .ZN(
        \SB2_2_3/buf_output[3] ) );
  NAND3_X2 U13095 ( .A1(\SB2_2_3/i0[10] ), .A2(\SB2_2_3/i1[9] ), .A3(
        \SB2_2_3/i1_7 ), .ZN(n6532) );
  NAND4_X2 U13096 ( .A1(\SB1_3_12/Component_Function_5/NAND4_in[2] ), .A2(
        \SB1_3_12/Component_Function_5/NAND4_in[1] ), .A3(
        \SB1_3_12/Component_Function_5/NAND4_in[0] ), .A4(n6533), .ZN(
        \SB1_3_12/buf_output[5] ) );
  XOR2_X1 U13097 ( .A1(\MC_ARK_ARC_1_3/buf_datainput[14] ), .A2(
        \MC_ARK_ARC_1_3/buf_datainput[38] ), .Z(n6534) );
  XOR2_X1 U13098 ( .A1(n3049), .A2(n6535), .Z(\MC_ARK_ARC_1_0/buf_output[101] ) );
  XOR2_X1 U13099 ( .A1(n4462), .A2(\MC_ARK_ARC_1_0/temp2[101] ), .Z(n6535) );
  NAND3_X2 U13100 ( .A1(\SB2_0_4/i0[10] ), .A2(\SB2_0_4/i0_0 ), .A3(
        \SB2_0_4/i0[6] ), .ZN(n3004) );
  NAND3_X1 U13101 ( .A1(n3668), .A2(\SB4_19/i1_7 ), .A3(\SB4_19/i0_4 ), .ZN(
        \SB4_19/Component_Function_1/NAND4_in[3] ) );
  NAND4_X2 U13102 ( .A1(\SB3_31/Component_Function_0/NAND4_in[2] ), .A2(
        \SB3_31/Component_Function_0/NAND4_in[0] ), .A3(
        \SB3_31/Component_Function_0/NAND4_in[1] ), .A4(n6537), .ZN(
        \SB3_31/buf_output[0] ) );
  XOR2_X1 U13103 ( .A1(n6538), .A2(n79), .Z(Ciphertext[29]) );
  INV_X1 U13104 ( .I(\MC_ARK_ARC_1_0/buf_output[18] ), .ZN(\SB1_1_28/i3[0] )
         );
  CLKBUF_X4 U13105 ( .I(\MC_ARK_ARC_1_0/buf_output[18] ), .Z(\SB1_1_28/i0[9] )
         );
  CLKBUF_X4 U13106 ( .I(\SB2_2_29/i0_4 ), .Z(n1837) );
endmodule


module SPEEDY_Top ( clk, Plaintext, Key, Ciphertext );
  input [191:0] Plaintext;
  input [191:0] Key;
  output [191:0] Ciphertext;
  input clk;

  wire   [191:0] reg_in;
  wire   [191:0] reg_key;
  wire   [191:0] reg_out;

  DFFSNQ_X1 \reg_in_reg[191]  ( .D(Plaintext[191]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[191]) );
  DFFSNQ_X1 \reg_in_reg[190]  ( .D(Plaintext[190]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[190]) );
  DFFSNQ_X1 \reg_in_reg[189]  ( .D(Plaintext[189]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[189]) );
  DFFSNQ_X1 \reg_in_reg[188]  ( .D(Plaintext[188]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[188]) );
  DFFSNQ_X1 \reg_in_reg[187]  ( .D(Plaintext[187]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[187]) );
  DFFSNQ_X1 \reg_in_reg[186]  ( .D(Plaintext[186]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[186]) );
  DFFSNQ_X1 \reg_in_reg[185]  ( .D(Plaintext[185]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[185]) );
  DFFSNQ_X1 \reg_in_reg[184]  ( .D(Plaintext[184]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[184]) );
  DFFSNQ_X1 \reg_in_reg[183]  ( .D(Plaintext[183]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[183]) );
  DFFSNQ_X1 \reg_in_reg[182]  ( .D(Plaintext[182]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[182]) );
  DFFSNQ_X1 \reg_in_reg[181]  ( .D(Plaintext[181]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[181]) );
  DFFSNQ_X1 \reg_in_reg[180]  ( .D(Plaintext[180]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[180]) );
  DFFSNQ_X1 \reg_in_reg[179]  ( .D(Plaintext[179]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[179]) );
  DFFSNQ_X1 \reg_in_reg[178]  ( .D(Plaintext[178]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[178]) );
  DFFSNQ_X1 \reg_in_reg[177]  ( .D(Plaintext[177]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[177]) );
  DFFSNQ_X1 \reg_in_reg[176]  ( .D(Plaintext[176]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[176]) );
  DFFSNQ_X1 \reg_in_reg[175]  ( .D(Plaintext[175]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[175]) );
  DFFSNQ_X1 \reg_in_reg[174]  ( .D(Plaintext[174]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[174]) );
  DFFSNQ_X1 \reg_in_reg[173]  ( .D(Plaintext[173]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[173]) );
  DFFSNQ_X1 \reg_in_reg[172]  ( .D(Plaintext[172]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[172]) );
  DFFSNQ_X1 \reg_in_reg[171]  ( .D(Plaintext[171]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[171]) );
  DFFSNQ_X1 \reg_in_reg[170]  ( .D(Plaintext[170]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[170]) );
  DFFSNQ_X1 \reg_in_reg[169]  ( .D(Plaintext[169]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[169]) );
  DFFSNQ_X1 \reg_in_reg[168]  ( .D(Plaintext[168]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[168]) );
  DFFSNQ_X1 \reg_in_reg[167]  ( .D(Plaintext[167]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[167]) );
  DFFSNQ_X1 \reg_in_reg[166]  ( .D(Plaintext[166]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[166]) );
  DFFSNQ_X1 \reg_in_reg[165]  ( .D(Plaintext[165]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[165]) );
  DFFSNQ_X1 \reg_in_reg[164]  ( .D(Plaintext[164]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[164]) );
  DFFSNQ_X1 \reg_in_reg[163]  ( .D(Plaintext[163]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[163]) );
  DFFSNQ_X1 \reg_in_reg[162]  ( .D(Plaintext[162]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[162]) );
  DFFSNQ_X1 \reg_in_reg[161]  ( .D(Plaintext[161]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[161]) );
  DFFSNQ_X1 \reg_in_reg[160]  ( .D(Plaintext[160]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[160]) );
  DFFSNQ_X1 \reg_in_reg[159]  ( .D(Plaintext[159]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[159]) );
  DFFSNQ_X1 \reg_in_reg[158]  ( .D(Plaintext[158]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[158]) );
  DFFSNQ_X1 \reg_in_reg[157]  ( .D(Plaintext[157]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[157]) );
  DFFSNQ_X1 \reg_in_reg[156]  ( .D(Plaintext[156]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[156]) );
  DFFSNQ_X1 \reg_in_reg[155]  ( .D(Plaintext[155]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[155]) );
  DFFSNQ_X1 \reg_in_reg[154]  ( .D(Plaintext[154]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[154]) );
  DFFSNQ_X1 \reg_in_reg[153]  ( .D(Plaintext[153]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[153]) );
  DFFSNQ_X1 \reg_in_reg[152]  ( .D(Plaintext[152]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[152]) );
  DFFSNQ_X1 \reg_in_reg[151]  ( .D(Plaintext[151]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[151]) );
  DFFSNQ_X1 \reg_in_reg[150]  ( .D(Plaintext[150]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[150]) );
  DFFSNQ_X1 \reg_in_reg[149]  ( .D(Plaintext[149]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[149]) );
  DFFSNQ_X1 \reg_in_reg[148]  ( .D(Plaintext[148]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[148]) );
  DFFSNQ_X1 \reg_in_reg[147]  ( .D(Plaintext[147]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[147]) );
  DFFSNQ_X1 \reg_in_reg[146]  ( .D(Plaintext[146]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[146]) );
  DFFSNQ_X1 \reg_in_reg[145]  ( .D(Plaintext[145]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[145]) );
  DFFSNQ_X1 \reg_in_reg[144]  ( .D(Plaintext[144]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[144]) );
  DFFSNQ_X1 \reg_in_reg[143]  ( .D(Plaintext[143]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[143]) );
  DFFSNQ_X1 \reg_in_reg[142]  ( .D(Plaintext[142]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[142]) );
  DFFSNQ_X1 \reg_in_reg[141]  ( .D(Plaintext[141]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[141]) );
  DFFSNQ_X1 \reg_in_reg[140]  ( .D(Plaintext[140]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[140]) );
  DFFSNQ_X1 \reg_in_reg[139]  ( .D(Plaintext[139]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[139]) );
  DFFSNQ_X1 \reg_in_reg[138]  ( .D(Plaintext[138]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[138]) );
  DFFSNQ_X1 \reg_in_reg[137]  ( .D(Plaintext[137]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[137]) );
  DFFSNQ_X1 \reg_in_reg[136]  ( .D(Plaintext[136]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[136]) );
  DFFSNQ_X1 \reg_in_reg[135]  ( .D(Plaintext[135]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[135]) );
  DFFSNQ_X1 \reg_in_reg[134]  ( .D(Plaintext[134]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[134]) );
  DFFSNQ_X1 \reg_in_reg[133]  ( .D(Plaintext[133]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[133]) );
  DFFSNQ_X1 \reg_in_reg[132]  ( .D(Plaintext[132]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[132]) );
  DFFSNQ_X1 \reg_in_reg[131]  ( .D(Plaintext[131]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[131]) );
  DFFSNQ_X1 \reg_in_reg[130]  ( .D(Plaintext[130]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[130]) );
  DFFSNQ_X1 \reg_in_reg[129]  ( .D(Plaintext[129]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[129]) );
  DFFSNQ_X1 \reg_in_reg[128]  ( .D(Plaintext[128]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[128]) );
  DFFSNQ_X1 \reg_in_reg[127]  ( .D(Plaintext[127]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[127]) );
  DFFSNQ_X1 \reg_in_reg[126]  ( .D(Plaintext[126]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[126]) );
  DFFSNQ_X1 \reg_in_reg[125]  ( .D(Plaintext[125]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[125]) );
  DFFSNQ_X1 \reg_in_reg[124]  ( .D(Plaintext[124]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[124]) );
  DFFSNQ_X1 \reg_in_reg[123]  ( .D(Plaintext[123]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[123]) );
  DFFSNQ_X1 \reg_in_reg[122]  ( .D(Plaintext[122]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[122]) );
  DFFSNQ_X1 \reg_in_reg[121]  ( .D(Plaintext[121]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[121]) );
  DFFSNQ_X1 \reg_in_reg[120]  ( .D(Plaintext[120]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[120]) );
  DFFSNQ_X1 \reg_in_reg[119]  ( .D(Plaintext[119]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[119]) );
  DFFSNQ_X1 \reg_in_reg[118]  ( .D(Plaintext[118]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[118]) );
  DFFSNQ_X1 \reg_in_reg[117]  ( .D(Plaintext[117]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[117]) );
  DFFSNQ_X1 \reg_in_reg[116]  ( .D(Plaintext[116]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[116]) );
  DFFSNQ_X1 \reg_in_reg[115]  ( .D(Plaintext[115]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[115]) );
  DFFSNQ_X1 \reg_in_reg[114]  ( .D(Plaintext[114]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[114]) );
  DFFSNQ_X1 \reg_in_reg[113]  ( .D(Plaintext[113]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[113]) );
  DFFSNQ_X1 \reg_in_reg[112]  ( .D(Plaintext[112]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[112]) );
  DFFSNQ_X1 \reg_in_reg[111]  ( .D(Plaintext[111]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[111]) );
  DFFSNQ_X1 \reg_in_reg[110]  ( .D(Plaintext[110]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[110]) );
  DFFSNQ_X1 \reg_in_reg[109]  ( .D(Plaintext[109]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[109]) );
  DFFSNQ_X1 \reg_in_reg[108]  ( .D(Plaintext[108]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[108]) );
  DFFSNQ_X1 \reg_in_reg[107]  ( .D(Plaintext[107]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[107]) );
  DFFSNQ_X1 \reg_in_reg[106]  ( .D(Plaintext[106]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[106]) );
  DFFSNQ_X1 \reg_in_reg[105]  ( .D(Plaintext[105]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[105]) );
  DFFSNQ_X1 \reg_in_reg[104]  ( .D(Plaintext[104]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[104]) );
  DFFSNQ_X1 \reg_in_reg[103]  ( .D(Plaintext[103]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[103]) );
  DFFSNQ_X1 \reg_in_reg[102]  ( .D(Plaintext[102]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[102]) );
  DFFSNQ_X1 \reg_in_reg[101]  ( .D(Plaintext[101]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[101]) );
  DFFSNQ_X1 \reg_in_reg[100]  ( .D(Plaintext[100]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[100]) );
  DFFSNQ_X1 \reg_in_reg[99]  ( .D(Plaintext[99]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[99]) );
  DFFSNQ_X1 \reg_in_reg[98]  ( .D(Plaintext[98]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[98]) );
  DFFSNQ_X1 \reg_in_reg[97]  ( .D(Plaintext[97]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[97]) );
  DFFSNQ_X1 \reg_in_reg[96]  ( .D(Plaintext[96]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[96]) );
  DFFSNQ_X1 \reg_in_reg[95]  ( .D(Plaintext[95]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[95]) );
  DFFSNQ_X1 \reg_in_reg[94]  ( .D(Plaintext[94]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[94]) );
  DFFSNQ_X1 \reg_in_reg[93]  ( .D(Plaintext[93]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[93]) );
  DFFSNQ_X1 \reg_in_reg[92]  ( .D(Plaintext[92]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[92]) );
  DFFSNQ_X1 \reg_in_reg[91]  ( .D(Plaintext[91]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[91]) );
  DFFSNQ_X1 \reg_in_reg[90]  ( .D(Plaintext[90]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[90]) );
  DFFSNQ_X1 \reg_in_reg[89]  ( .D(Plaintext[89]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[89]) );
  DFFSNQ_X1 \reg_in_reg[88]  ( .D(Plaintext[88]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[88]) );
  DFFSNQ_X1 \reg_in_reg[87]  ( .D(Plaintext[87]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[87]) );
  DFFSNQ_X1 \reg_in_reg[86]  ( .D(Plaintext[86]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[86]) );
  DFFSNQ_X1 \reg_in_reg[85]  ( .D(Plaintext[85]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[85]) );
  DFFSNQ_X1 \reg_in_reg[84]  ( .D(Plaintext[84]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[84]) );
  DFFSNQ_X1 \reg_in_reg[83]  ( .D(Plaintext[83]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[83]) );
  DFFSNQ_X1 \reg_in_reg[82]  ( .D(Plaintext[82]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[82]) );
  DFFSNQ_X1 \reg_in_reg[81]  ( .D(Plaintext[81]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[81]) );
  DFFSNQ_X1 \reg_in_reg[80]  ( .D(Plaintext[80]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[80]) );
  DFFSNQ_X1 \reg_in_reg[79]  ( .D(Plaintext[79]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[79]) );
  DFFSNQ_X1 \reg_in_reg[78]  ( .D(Plaintext[78]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[78]) );
  DFFSNQ_X1 \reg_in_reg[77]  ( .D(Plaintext[77]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[77]) );
  DFFSNQ_X1 \reg_in_reg[76]  ( .D(Plaintext[76]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[76]) );
  DFFSNQ_X1 \reg_in_reg[75]  ( .D(Plaintext[75]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[75]) );
  DFFSNQ_X1 \reg_in_reg[74]  ( .D(Plaintext[74]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[74]) );
  DFFSNQ_X1 \reg_in_reg[73]  ( .D(Plaintext[73]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[73]) );
  DFFSNQ_X1 \reg_in_reg[72]  ( .D(Plaintext[72]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[72]) );
  DFFSNQ_X1 \reg_in_reg[71]  ( .D(Plaintext[71]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[71]) );
  DFFSNQ_X1 \reg_in_reg[70]  ( .D(Plaintext[70]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[70]) );
  DFFSNQ_X1 \reg_in_reg[69]  ( .D(Plaintext[69]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[69]) );
  DFFSNQ_X1 \reg_in_reg[68]  ( .D(Plaintext[68]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[68]) );
  DFFSNQ_X1 \reg_in_reg[67]  ( .D(Plaintext[67]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[67]) );
  DFFSNQ_X1 \reg_in_reg[66]  ( .D(Plaintext[66]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[66]) );
  DFFSNQ_X1 \reg_in_reg[65]  ( .D(Plaintext[65]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[65]) );
  DFFSNQ_X1 \reg_in_reg[64]  ( .D(Plaintext[64]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[64]) );
  DFFSNQ_X1 \reg_in_reg[63]  ( .D(Plaintext[63]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[63]) );
  DFFSNQ_X1 \reg_in_reg[62]  ( .D(Plaintext[62]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[62]) );
  DFFSNQ_X1 \reg_in_reg[61]  ( .D(Plaintext[61]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[61]) );
  DFFSNQ_X1 \reg_in_reg[60]  ( .D(Plaintext[60]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[60]) );
  DFFSNQ_X1 \reg_in_reg[59]  ( .D(Plaintext[59]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[59]) );
  DFFSNQ_X1 \reg_in_reg[58]  ( .D(Plaintext[58]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[58]) );
  DFFSNQ_X1 \reg_in_reg[57]  ( .D(Plaintext[57]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[57]) );
  DFFSNQ_X1 \reg_in_reg[56]  ( .D(Plaintext[56]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[56]) );
  DFFSNQ_X1 \reg_in_reg[55]  ( .D(Plaintext[55]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[55]) );
  DFFSNQ_X1 \reg_in_reg[54]  ( .D(Plaintext[54]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[54]) );
  DFFSNQ_X1 \reg_in_reg[53]  ( .D(Plaintext[53]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[53]) );
  DFFSNQ_X1 \reg_in_reg[52]  ( .D(Plaintext[52]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[52]) );
  DFFSNQ_X1 \reg_in_reg[51]  ( .D(Plaintext[51]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[51]) );
  DFFSNQ_X1 \reg_in_reg[50]  ( .D(Plaintext[50]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[50]) );
  DFFSNQ_X1 \reg_in_reg[49]  ( .D(Plaintext[49]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[49]) );
  DFFSNQ_X1 \reg_in_reg[48]  ( .D(Plaintext[48]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[48]) );
  DFFSNQ_X1 \reg_in_reg[47]  ( .D(Plaintext[47]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[47]) );
  DFFSNQ_X1 \reg_in_reg[46]  ( .D(Plaintext[46]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[46]) );
  DFFSNQ_X1 \reg_in_reg[45]  ( .D(Plaintext[45]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[45]) );
  DFFSNQ_X1 \reg_in_reg[44]  ( .D(Plaintext[44]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[44]) );
  DFFSNQ_X1 \reg_in_reg[43]  ( .D(Plaintext[43]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[43]) );
  DFFSNQ_X1 \reg_in_reg[42]  ( .D(Plaintext[42]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[42]) );
  DFFSNQ_X1 \reg_in_reg[41]  ( .D(Plaintext[41]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[41]) );
  DFFSNQ_X1 \reg_in_reg[40]  ( .D(Plaintext[40]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[40]) );
  DFFSNQ_X1 \reg_in_reg[39]  ( .D(Plaintext[39]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[39]) );
  DFFSNQ_X1 \reg_in_reg[38]  ( .D(Plaintext[38]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[38]) );
  DFFSNQ_X1 \reg_in_reg[37]  ( .D(Plaintext[37]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[37]) );
  DFFSNQ_X1 \reg_in_reg[36]  ( .D(Plaintext[36]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[36]) );
  DFFSNQ_X1 \reg_in_reg[35]  ( .D(Plaintext[35]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[35]) );
  DFFSNQ_X1 \reg_in_reg[34]  ( .D(Plaintext[34]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[34]) );
  DFFSNQ_X1 \reg_in_reg[33]  ( .D(Plaintext[33]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[33]) );
  DFFSNQ_X1 \reg_in_reg[32]  ( .D(Plaintext[32]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[32]) );
  DFFSNQ_X1 \reg_in_reg[31]  ( .D(Plaintext[31]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[31]) );
  DFFSNQ_X1 \reg_in_reg[30]  ( .D(Plaintext[30]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[30]) );
  DFFSNQ_X1 \reg_in_reg[29]  ( .D(Plaintext[29]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[29]) );
  DFFSNQ_X1 \reg_in_reg[28]  ( .D(Plaintext[28]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[28]) );
  DFFSNQ_X1 \reg_in_reg[27]  ( .D(Plaintext[27]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[27]) );
  DFFSNQ_X1 \reg_in_reg[26]  ( .D(Plaintext[26]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[26]) );
  DFFSNQ_X1 \reg_in_reg[25]  ( .D(Plaintext[25]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[25]) );
  DFFSNQ_X1 \reg_in_reg[24]  ( .D(Plaintext[24]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[24]) );
  DFFSNQ_X1 \reg_in_reg[23]  ( .D(Plaintext[23]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[23]) );
  DFFSNQ_X1 \reg_in_reg[22]  ( .D(Plaintext[22]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[22]) );
  DFFSNQ_X1 \reg_in_reg[21]  ( .D(Plaintext[21]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[21]) );
  DFFSNQ_X1 \reg_in_reg[20]  ( .D(Plaintext[20]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[20]) );
  DFFSNQ_X1 \reg_in_reg[19]  ( .D(Plaintext[19]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[19]) );
  DFFSNQ_X1 \reg_in_reg[18]  ( .D(Plaintext[18]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[18]) );
  DFFSNQ_X1 \reg_in_reg[17]  ( .D(Plaintext[17]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[17]) );
  DFFSNQ_X1 \reg_in_reg[16]  ( .D(Plaintext[16]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[16]) );
  DFFSNQ_X1 \reg_in_reg[15]  ( .D(Plaintext[15]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[15]) );
  DFFSNQ_X1 \reg_in_reg[14]  ( .D(Plaintext[14]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[14]) );
  DFFSNQ_X1 \reg_in_reg[13]  ( .D(Plaintext[13]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[13]) );
  DFFSNQ_X1 \reg_in_reg[12]  ( .D(Plaintext[12]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[12]) );
  DFFSNQ_X1 \reg_in_reg[11]  ( .D(Plaintext[11]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[11]) );
  DFFSNQ_X1 \reg_in_reg[10]  ( .D(Plaintext[10]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[10]) );
  DFFSNQ_X1 \reg_in_reg[9]  ( .D(Plaintext[9]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[9]) );
  DFFSNQ_X1 \reg_in_reg[8]  ( .D(Plaintext[8]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[8]) );
  DFFSNQ_X1 \reg_in_reg[7]  ( .D(Plaintext[7]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[7]) );
  DFFSNQ_X1 \reg_in_reg[6]  ( .D(Plaintext[6]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[6]) );
  DFFSNQ_X1 \reg_in_reg[5]  ( .D(Plaintext[5]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[5]) );
  DFFSNQ_X1 \reg_in_reg[4]  ( .D(Plaintext[4]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[4]) );
  DFFSNQ_X1 \reg_in_reg[3]  ( .D(Plaintext[3]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[3]) );
  DFFSNQ_X1 \reg_in_reg[2]  ( .D(Plaintext[2]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[2]) );
  DFFSNQ_X1 \reg_in_reg[1]  ( .D(Plaintext[1]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[1]) );
  DFFSNQ_X1 \reg_in_reg[0]  ( .D(Plaintext[0]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[0]) );
  DFFSNQ_X1 \reg_key_reg[191]  ( .D(Key[191]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[191]) );
  DFFSNQ_X1 \reg_key_reg[190]  ( .D(Key[190]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[190]) );
  DFFSNQ_X1 \reg_key_reg[189]  ( .D(Key[189]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[189]) );
  DFFSNQ_X1 \reg_key_reg[188]  ( .D(Key[188]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[188]) );
  DFFSNQ_X1 \reg_key_reg[187]  ( .D(Key[187]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[187]) );
  DFFSNQ_X1 \reg_key_reg[186]  ( .D(Key[186]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[186]) );
  DFFSNQ_X1 \reg_key_reg[185]  ( .D(Key[185]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[185]) );
  DFFSNQ_X1 \reg_key_reg[184]  ( .D(Key[184]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[184]) );
  DFFSNQ_X1 \reg_key_reg[183]  ( .D(Key[183]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[183]) );
  DFFSNQ_X1 \reg_key_reg[182]  ( .D(Key[182]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[182]) );
  DFFSNQ_X1 \reg_key_reg[181]  ( .D(Key[181]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[181]) );
  DFFSNQ_X1 \reg_key_reg[180]  ( .D(Key[180]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[180]) );
  DFFSNQ_X1 \reg_key_reg[179]  ( .D(Key[179]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[179]) );
  DFFSNQ_X1 \reg_key_reg[178]  ( .D(Key[178]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[178]) );
  DFFSNQ_X1 \reg_key_reg[177]  ( .D(Key[177]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[177]) );
  DFFSNQ_X1 \reg_key_reg[176]  ( .D(Key[176]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[176]) );
  DFFSNQ_X1 \reg_key_reg[175]  ( .D(Key[175]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[175]) );
  DFFSNQ_X1 \reg_key_reg[174]  ( .D(Key[174]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[174]) );
  DFFSNQ_X1 \reg_key_reg[173]  ( .D(Key[173]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[173]) );
  DFFSNQ_X1 \reg_key_reg[172]  ( .D(Key[172]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[172]) );
  DFFSNQ_X1 \reg_key_reg[171]  ( .D(Key[171]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[171]) );
  DFFSNQ_X1 \reg_key_reg[170]  ( .D(Key[170]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[170]) );
  DFFSNQ_X1 \reg_key_reg[169]  ( .D(Key[169]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[169]) );
  DFFSNQ_X1 \reg_key_reg[168]  ( .D(Key[168]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[168]) );
  DFFSNQ_X1 \reg_key_reg[167]  ( .D(Key[167]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[167]) );
  DFFSNQ_X1 \reg_key_reg[166]  ( .D(Key[166]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[166]) );
  DFFSNQ_X1 \reg_key_reg[165]  ( .D(Key[165]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[165]) );
  DFFSNQ_X1 \reg_key_reg[164]  ( .D(Key[164]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[164]) );
  DFFSNQ_X1 \reg_key_reg[163]  ( .D(Key[163]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[163]) );
  DFFSNQ_X1 \reg_key_reg[162]  ( .D(Key[162]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[162]) );
  DFFSNQ_X1 \reg_key_reg[161]  ( .D(Key[161]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[161]) );
  DFFSNQ_X1 \reg_key_reg[160]  ( .D(Key[160]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[160]) );
  DFFSNQ_X1 \reg_key_reg[159]  ( .D(Key[159]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[159]) );
  DFFSNQ_X1 \reg_key_reg[158]  ( .D(Key[158]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[158]) );
  DFFSNQ_X1 \reg_key_reg[157]  ( .D(Key[157]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[157]) );
  DFFSNQ_X1 \reg_key_reg[156]  ( .D(Key[156]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[156]) );
  DFFSNQ_X1 \reg_key_reg[155]  ( .D(Key[155]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[155]) );
  DFFSNQ_X1 \reg_key_reg[154]  ( .D(Key[154]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[154]) );
  DFFSNQ_X1 \reg_key_reg[153]  ( .D(Key[153]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[153]) );
  DFFSNQ_X1 \reg_key_reg[152]  ( .D(Key[152]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[152]) );
  DFFSNQ_X1 \reg_key_reg[151]  ( .D(Key[151]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[151]) );
  DFFSNQ_X1 \reg_key_reg[150]  ( .D(Key[150]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[150]) );
  DFFSNQ_X1 \reg_key_reg[149]  ( .D(Key[149]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[149]) );
  DFFSNQ_X1 \reg_key_reg[148]  ( .D(Key[148]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[148]) );
  DFFSNQ_X1 \reg_key_reg[147]  ( .D(Key[147]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[147]) );
  DFFSNQ_X1 \reg_key_reg[146]  ( .D(Key[146]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[146]) );
  DFFSNQ_X1 \reg_key_reg[145]  ( .D(Key[145]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[145]) );
  DFFSNQ_X1 \reg_key_reg[144]  ( .D(Key[144]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[144]) );
  DFFSNQ_X1 \reg_key_reg[143]  ( .D(Key[143]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[143]) );
  DFFSNQ_X1 \reg_key_reg[142]  ( .D(Key[142]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[142]) );
  DFFSNQ_X1 \reg_key_reg[141]  ( .D(Key[141]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[141]) );
  DFFSNQ_X1 \reg_key_reg[140]  ( .D(Key[140]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[140]) );
  DFFSNQ_X1 \reg_key_reg[139]  ( .D(Key[139]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[139]) );
  DFFSNQ_X1 \reg_key_reg[138]  ( .D(Key[138]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[138]) );
  DFFSNQ_X1 \reg_key_reg[137]  ( .D(Key[137]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[137]) );
  DFFSNQ_X1 \reg_key_reg[136]  ( .D(Key[136]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[136]) );
  DFFSNQ_X1 \reg_key_reg[135]  ( .D(Key[135]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[135]) );
  DFFSNQ_X1 \reg_key_reg[134]  ( .D(Key[134]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[134]) );
  DFFSNQ_X1 \reg_key_reg[133]  ( .D(Key[133]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[133]) );
  DFFSNQ_X1 \reg_key_reg[132]  ( .D(Key[132]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[132]) );
  DFFSNQ_X1 \reg_key_reg[131]  ( .D(Key[131]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[131]) );
  DFFSNQ_X1 \reg_key_reg[130]  ( .D(Key[130]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[130]) );
  DFFSNQ_X1 \reg_key_reg[129]  ( .D(Key[129]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[129]) );
  DFFSNQ_X1 \reg_key_reg[128]  ( .D(Key[128]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[128]) );
  DFFSNQ_X1 \reg_key_reg[127]  ( .D(Key[127]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[127]) );
  DFFSNQ_X1 \reg_key_reg[126]  ( .D(Key[126]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[126]) );
  DFFSNQ_X1 \reg_key_reg[125]  ( .D(Key[125]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[125]) );
  DFFSNQ_X1 \reg_key_reg[124]  ( .D(Key[124]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[124]) );
  DFFSNQ_X1 \reg_key_reg[123]  ( .D(Key[123]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[123]) );
  DFFSNQ_X1 \reg_key_reg[122]  ( .D(Key[122]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[122]) );
  DFFSNQ_X1 \reg_key_reg[121]  ( .D(Key[121]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[121]) );
  DFFSNQ_X1 \reg_key_reg[120]  ( .D(Key[120]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[120]) );
  DFFSNQ_X1 \reg_key_reg[119]  ( .D(Key[119]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[119]) );
  DFFSNQ_X1 \reg_key_reg[118]  ( .D(Key[118]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[118]) );
  DFFSNQ_X1 \reg_key_reg[117]  ( .D(Key[117]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[117]) );
  DFFSNQ_X1 \reg_key_reg[116]  ( .D(Key[116]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[116]) );
  DFFSNQ_X1 \reg_key_reg[115]  ( .D(Key[115]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[115]) );
  DFFSNQ_X1 \reg_key_reg[114]  ( .D(Key[114]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[114]) );
  DFFSNQ_X1 \reg_key_reg[113]  ( .D(Key[113]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[113]) );
  DFFSNQ_X1 \reg_key_reg[112]  ( .D(Key[112]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[112]) );
  DFFSNQ_X1 \reg_key_reg[111]  ( .D(Key[111]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[111]) );
  DFFSNQ_X1 \reg_key_reg[110]  ( .D(Key[110]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[110]) );
  DFFSNQ_X1 \reg_key_reg[109]  ( .D(Key[109]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[109]) );
  DFFSNQ_X1 \reg_key_reg[108]  ( .D(Key[108]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[108]) );
  DFFSNQ_X1 \reg_key_reg[107]  ( .D(Key[107]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[107]) );
  DFFSNQ_X1 \reg_key_reg[106]  ( .D(Key[106]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[106]) );
  DFFSNQ_X1 \reg_key_reg[105]  ( .D(Key[105]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[105]) );
  DFFSNQ_X1 \reg_key_reg[104]  ( .D(Key[104]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[104]) );
  DFFSNQ_X1 \reg_key_reg[103]  ( .D(Key[103]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[103]) );
  DFFSNQ_X1 \reg_key_reg[102]  ( .D(Key[102]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[102]) );
  DFFSNQ_X1 \reg_key_reg[101]  ( .D(Key[101]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[101]) );
  DFFSNQ_X1 \reg_key_reg[100]  ( .D(Key[100]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[100]) );
  DFFSNQ_X1 \reg_key_reg[99]  ( .D(Key[99]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[99]) );
  DFFSNQ_X1 \reg_key_reg[98]  ( .D(Key[98]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[98]) );
  DFFSNQ_X1 \reg_key_reg[97]  ( .D(Key[97]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[97]) );
  DFFSNQ_X1 \reg_key_reg[96]  ( .D(Key[96]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[96]) );
  DFFSNQ_X1 \reg_key_reg[95]  ( .D(Key[95]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[95]) );
  DFFSNQ_X1 \reg_key_reg[94]  ( .D(Key[94]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[94]) );
  DFFSNQ_X1 \reg_key_reg[93]  ( .D(Key[93]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[93]) );
  DFFSNQ_X1 \reg_key_reg[92]  ( .D(Key[92]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[92]) );
  DFFSNQ_X1 \reg_key_reg[91]  ( .D(Key[91]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[91]) );
  DFFSNQ_X1 \reg_key_reg[90]  ( .D(Key[90]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[90]) );
  DFFSNQ_X1 \reg_key_reg[89]  ( .D(Key[89]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[89]) );
  DFFSNQ_X1 \reg_key_reg[88]  ( .D(Key[88]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[88]) );
  DFFSNQ_X1 \reg_key_reg[87]  ( .D(Key[87]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[87]) );
  DFFSNQ_X1 \reg_key_reg[86]  ( .D(Key[86]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[86]) );
  DFFSNQ_X1 \reg_key_reg[85]  ( .D(Key[85]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[85]) );
  DFFSNQ_X1 \reg_key_reg[84]  ( .D(Key[84]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[84]) );
  DFFSNQ_X1 \reg_key_reg[83]  ( .D(Key[83]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[83]) );
  DFFSNQ_X1 \reg_key_reg[82]  ( .D(Key[82]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[82]) );
  DFFSNQ_X1 \reg_key_reg[81]  ( .D(Key[81]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[81]) );
  DFFSNQ_X1 \reg_key_reg[80]  ( .D(Key[80]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[80]) );
  DFFSNQ_X1 \reg_key_reg[79]  ( .D(Key[79]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[79]) );
  DFFSNQ_X1 \reg_key_reg[78]  ( .D(Key[78]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[78]) );
  DFFSNQ_X1 \reg_key_reg[77]  ( .D(Key[77]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[77]) );
  DFFSNQ_X1 \reg_key_reg[76]  ( .D(Key[76]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[76]) );
  DFFSNQ_X1 \reg_key_reg[75]  ( .D(Key[75]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[75]) );
  DFFSNQ_X1 \reg_key_reg[74]  ( .D(Key[74]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[74]) );
  DFFSNQ_X1 \reg_key_reg[73]  ( .D(Key[73]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[73]) );
  DFFSNQ_X1 \reg_key_reg[72]  ( .D(Key[72]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[72]) );
  DFFSNQ_X1 \reg_key_reg[71]  ( .D(Key[71]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[71]) );
  DFFSNQ_X1 \reg_key_reg[70]  ( .D(Key[70]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[70]) );
  DFFSNQ_X1 \reg_key_reg[69]  ( .D(Key[69]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[69]) );
  DFFSNQ_X1 \reg_key_reg[68]  ( .D(Key[68]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[68]) );
  DFFSNQ_X1 \reg_key_reg[67]  ( .D(Key[67]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[67]) );
  DFFSNQ_X1 \reg_key_reg[66]  ( .D(Key[66]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[66]) );
  DFFSNQ_X1 \reg_key_reg[65]  ( .D(Key[65]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[65]) );
  DFFSNQ_X1 \reg_key_reg[64]  ( .D(Key[64]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[64]) );
  DFFSNQ_X1 \reg_key_reg[63]  ( .D(Key[63]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[63]) );
  DFFSNQ_X1 \reg_key_reg[62]  ( .D(Key[62]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[62]) );
  DFFSNQ_X1 \reg_key_reg[61]  ( .D(Key[61]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[61]) );
  DFFSNQ_X1 \reg_key_reg[60]  ( .D(Key[60]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[60]) );
  DFFSNQ_X1 \reg_key_reg[59]  ( .D(Key[59]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[59]) );
  DFFSNQ_X1 \reg_key_reg[58]  ( .D(Key[58]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[58]) );
  DFFSNQ_X1 \reg_key_reg[57]  ( .D(Key[57]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[57]) );
  DFFSNQ_X1 \reg_key_reg[56]  ( .D(Key[56]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[56]) );
  DFFSNQ_X1 \reg_key_reg[55]  ( .D(Key[55]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[55]) );
  DFFSNQ_X1 \reg_key_reg[54]  ( .D(Key[54]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[54]) );
  DFFSNQ_X1 \reg_key_reg[53]  ( .D(Key[53]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[53]) );
  DFFSNQ_X1 \reg_key_reg[52]  ( .D(Key[52]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[52]) );
  DFFSNQ_X1 \reg_key_reg[51]  ( .D(Key[51]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[51]) );
  DFFSNQ_X1 \reg_key_reg[50]  ( .D(Key[50]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[50]) );
  DFFSNQ_X1 \reg_key_reg[49]  ( .D(Key[49]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[49]) );
  DFFSNQ_X1 \reg_key_reg[48]  ( .D(Key[48]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[48]) );
  DFFSNQ_X1 \reg_key_reg[47]  ( .D(Key[47]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[47]) );
  DFFSNQ_X1 \reg_key_reg[46]  ( .D(Key[46]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[46]) );
  DFFSNQ_X1 \reg_key_reg[45]  ( .D(Key[45]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[45]) );
  DFFSNQ_X1 \reg_key_reg[44]  ( .D(Key[44]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[44]) );
  DFFSNQ_X1 \reg_key_reg[43]  ( .D(Key[43]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[43]) );
  DFFSNQ_X1 \reg_key_reg[42]  ( .D(Key[42]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[42]) );
  DFFSNQ_X1 \reg_key_reg[41]  ( .D(Key[41]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[41]) );
  DFFSNQ_X1 \reg_key_reg[40]  ( .D(Key[40]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[40]) );
  DFFSNQ_X1 \reg_key_reg[39]  ( .D(Key[39]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[39]) );
  DFFSNQ_X1 \reg_key_reg[38]  ( .D(Key[38]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[38]) );
  DFFSNQ_X1 \reg_key_reg[37]  ( .D(Key[37]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[37]) );
  DFFSNQ_X1 \reg_key_reg[36]  ( .D(Key[36]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[36]) );
  DFFSNQ_X1 \reg_key_reg[35]  ( .D(Key[35]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[35]) );
  DFFSNQ_X1 \reg_key_reg[34]  ( .D(Key[34]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[34]) );
  DFFSNQ_X1 \reg_key_reg[33]  ( .D(Key[33]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[33]) );
  DFFSNQ_X1 \reg_key_reg[32]  ( .D(Key[32]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[32]) );
  DFFSNQ_X1 \reg_key_reg[31]  ( .D(Key[31]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[31]) );
  DFFSNQ_X1 \reg_key_reg[30]  ( .D(Key[30]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[30]) );
  DFFSNQ_X1 \reg_key_reg[29]  ( .D(Key[29]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[29]) );
  DFFSNQ_X1 \reg_key_reg[28]  ( .D(Key[28]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[28]) );
  DFFSNQ_X1 \reg_key_reg[27]  ( .D(Key[27]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[27]) );
  DFFSNQ_X1 \reg_key_reg[26]  ( .D(Key[26]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[26]) );
  DFFSNQ_X1 \reg_key_reg[25]  ( .D(Key[25]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[25]) );
  DFFSNQ_X1 \reg_key_reg[24]  ( .D(Key[24]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[24]) );
  DFFSNQ_X1 \reg_key_reg[23]  ( .D(Key[23]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[23]) );
  DFFSNQ_X1 \reg_key_reg[22]  ( .D(Key[22]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[22]) );
  DFFSNQ_X1 \reg_key_reg[21]  ( .D(Key[21]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[21]) );
  DFFSNQ_X1 \reg_key_reg[20]  ( .D(Key[20]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[20]) );
  DFFSNQ_X1 \reg_key_reg[19]  ( .D(Key[19]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[19]) );
  DFFSNQ_X1 \reg_key_reg[18]  ( .D(Key[18]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[18]) );
  DFFSNQ_X1 \reg_key_reg[17]  ( .D(Key[17]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[17]) );
  DFFSNQ_X1 \reg_key_reg[16]  ( .D(Key[16]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[16]) );
  DFFSNQ_X1 \reg_key_reg[15]  ( .D(Key[15]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[15]) );
  DFFSNQ_X1 \reg_key_reg[14]  ( .D(Key[14]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[14]) );
  DFFSNQ_X1 \reg_key_reg[13]  ( .D(Key[13]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[13]) );
  DFFSNQ_X1 \reg_key_reg[12]  ( .D(Key[12]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[12]) );
  DFFSNQ_X1 \reg_key_reg[11]  ( .D(Key[11]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[11]) );
  DFFSNQ_X1 \reg_key_reg[10]  ( .D(Key[10]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[10]) );
  DFFSNQ_X1 \reg_key_reg[9]  ( .D(Key[9]), .CLK(clk), .SN(1'b1), .Q(reg_key[9]) );
  DFFSNQ_X1 \reg_key_reg[8]  ( .D(Key[8]), .CLK(clk), .SN(1'b1), .Q(reg_key[8]) );
  DFFSNQ_X1 \reg_key_reg[7]  ( .D(Key[7]), .CLK(clk), .SN(1'b1), .Q(reg_key[7]) );
  DFFSNQ_X1 \reg_key_reg[6]  ( .D(Key[6]), .CLK(clk), .SN(1'b1), .Q(reg_key[6]) );
  DFFSNQ_X1 \reg_key_reg[5]  ( .D(Key[5]), .CLK(clk), .SN(1'b1), .Q(reg_key[5]) );
  DFFSNQ_X1 \reg_key_reg[4]  ( .D(Key[4]), .CLK(clk), .SN(1'b1), .Q(reg_key[4]) );
  DFFSNQ_X1 \reg_key_reg[3]  ( .D(Key[3]), .CLK(clk), .SN(1'b1), .Q(reg_key[3]) );
  DFFSNQ_X1 \reg_key_reg[2]  ( .D(Key[2]), .CLK(clk), .SN(1'b1), .Q(reg_key[2]) );
  DFFSNQ_X1 \reg_key_reg[1]  ( .D(Key[1]), .CLK(clk), .SN(1'b1), .Q(reg_key[1]) );
  DFFSNQ_X1 \reg_key_reg[0]  ( .D(Key[0]), .CLK(clk), .SN(1'b1), .Q(reg_key[0]) );
  DFFRNQ_X1 \Ciphertext_reg[127]  ( .D(reg_out[127]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[127]) );
  DFFRNQ_X1 \Ciphertext_reg[145]  ( .D(reg_out[145]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[145]) );
  DFFRNQ_X1 \Ciphertext_reg[171]  ( .D(reg_out[171]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[171]) );
  DFFRNQ_X1 \Ciphertext_reg[60]  ( .D(reg_out[60]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[60]) );
  DFFRNQ_X1 \Ciphertext_reg[63]  ( .D(reg_out[63]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[63]) );
  DFFRNQ_X1 \Ciphertext_reg[147]  ( .D(reg_out[147]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[147]) );
  DFFRNQ_X1 \Ciphertext_reg[103]  ( .D(reg_out[103]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[103]) );
  DFFRNQ_X1 \Ciphertext_reg[13]  ( .D(reg_out[13]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[13]) );
  DFFRNQ_X1 \Ciphertext_reg[172]  ( .D(reg_out[172]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[172]) );
  DFFRNQ_X1 \Ciphertext_reg[143]  ( .D(reg_out[143]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[143]) );
  DFFRNQ_X1 \Ciphertext_reg[135]  ( .D(reg_out[135]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[135]) );
  DFFRNQ_X1 \Ciphertext_reg[174]  ( .D(reg_out[174]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[174]) );
  DFFRNQ_X1 \Ciphertext_reg[138]  ( .D(reg_out[138]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[138]) );
  DFFRNQ_X1 \Ciphertext_reg[141]  ( .D(reg_out[141]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[141]) );
  DFFRNQ_X1 \Ciphertext_reg[146]  ( .D(reg_out[146]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[146]) );
  DFFRNQ_X1 \Ciphertext_reg[58]  ( .D(reg_out[58]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[58]) );
  DFFRNQ_X1 \Ciphertext_reg[169]  ( .D(reg_out[169]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[169]) );
  DFFRNQ_X1 \Ciphertext_reg[173]  ( .D(reg_out[173]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[173]) );
  DFFRNQ_X1 \Ciphertext_reg[87]  ( .D(reg_out[87]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[87]) );
  DFFRNQ_X1 \Ciphertext_reg[149]  ( .D(reg_out[149]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[149]) );
  DFFRNQ_X1 \Ciphertext_reg[55]  ( .D(reg_out[55]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[55]) );
  DFFRNQ_X1 \Ciphertext_reg[144]  ( .D(reg_out[144]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[144]) );
  DFFRNQ_X1 \Ciphertext_reg[45]  ( .D(reg_out[45]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[45]) );
  DFFRNQ_X1 \Ciphertext_reg[86]  ( .D(reg_out[86]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[86]) );
  DFFRNQ_X1 \Ciphertext_reg[126]  ( .D(reg_out[126]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[126]) );
  DFFRNQ_X1 \Ciphertext_reg[21]  ( .D(reg_out[21]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[21]) );
  DFFRNQ_X1 \Ciphertext_reg[37]  ( .D(reg_out[37]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[37]) );
  DFFRNQ_X1 \Ciphertext_reg[133]  ( .D(reg_out[133]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[133]) );
  DFFRNQ_X1 \Ciphertext_reg[108]  ( .D(reg_out[108]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[108]) );
  DFFRNQ_X1 \Ciphertext_reg[54]  ( .D(reg_out[54]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[54]) );
  DFFRNQ_X1 \Ciphertext_reg[79]  ( .D(reg_out[79]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[79]) );
  DFFRNQ_X1 \Ciphertext_reg[20]  ( .D(reg_out[20]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[20]) );
  DFFRNQ_X1 \Ciphertext_reg[128]  ( .D(reg_out[128]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[128]) );
  DFFRNQ_X1 \Ciphertext_reg[11]  ( .D(reg_out[11]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[11]) );
  DFFRNQ_X1 \Ciphertext_reg[148]  ( .D(reg_out[148]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[148]) );
  DFFRNQ_X1 \Ciphertext_reg[59]  ( .D(reg_out[59]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[59]) );
  DFFRNQ_X1 \Ciphertext_reg[19]  ( .D(reg_out[19]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[19]) );
  DFFRNQ_X1 \Ciphertext_reg[84]  ( .D(reg_out[84]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[84]) );
  DFFRNQ_X1 \Ciphertext_reg[51]  ( .D(reg_out[51]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[51]) );
  DFFRNQ_X1 \Ciphertext_reg[77]  ( .D(reg_out[77]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[77]) );
  DFFRNQ_X1 \Ciphertext_reg[97]  ( .D(reg_out[97]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[97]) );
  DFFRNQ_X1 \Ciphertext_reg[164]  ( .D(reg_out[164]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[164]) );
  DFFRNQ_X1 \Ciphertext_reg[150]  ( .D(reg_out[150]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[150]) );
  DFFRNQ_X1 \Ciphertext_reg[100]  ( .D(reg_out[100]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[100]) );
  DFFRNQ_X1 \Ciphertext_reg[175]  ( .D(reg_out[175]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[175]) );
  DFFRNQ_X1 \Ciphertext_reg[96]  ( .D(reg_out[96]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[96]) );
  DFFRNQ_X1 \Ciphertext_reg[107]  ( .D(reg_out[107]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[107]) );
  DFFRNQ_X1 \Ciphertext_reg[142]  ( .D(reg_out[142]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[142]) );
  DFFRNQ_X1 \Ciphertext_reg[22]  ( .D(reg_out[22]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[22]) );
  DFFRNQ_X1 \Ciphertext_reg[23]  ( .D(reg_out[23]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[23]) );
  DFFRNQ_X1 \Ciphertext_reg[66]  ( .D(reg_out[66]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[66]) );
  DFFRNQ_X1 \Ciphertext_reg[163]  ( .D(reg_out[163]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[163]) );
  DFFRNQ_X1 \Ciphertext_reg[1]  ( .D(reg_out[1]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[1]) );
  DFFRNQ_X1 \Ciphertext_reg[7]  ( .D(reg_out[7]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[7]) );
  DFFRNQ_X1 \Ciphertext_reg[80]  ( .D(reg_out[80]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[80]) );
  DFFRNQ_X1 \Ciphertext_reg[18]  ( .D(reg_out[18]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[18]) );
  DFFRNQ_X1 \Ciphertext_reg[85]  ( .D(reg_out[85]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[85]) );
  DFFRNQ_X1 \Ciphertext_reg[69]  ( .D(reg_out[69]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[69]) );
  DFFRNQ_X1 \Ciphertext_reg[9]  ( .D(reg_out[9]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[9]) );
  DFFRNQ_X1 \Ciphertext_reg[10]  ( .D(reg_out[10]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[10]) );
  DFFRNQ_X1 \Ciphertext_reg[65]  ( .D(reg_out[65]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[65]) );
  DFFRNQ_X1 \Ciphertext_reg[179]  ( .D(reg_out[179]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[179]) );
  DFFRNQ_X1 \Ciphertext_reg[167]  ( .D(reg_out[167]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[167]) );
  DFFRNQ_X1 \Ciphertext_reg[88]  ( .D(reg_out[88]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[88]) );
  DFFRNQ_X1 \Ciphertext_reg[153]  ( .D(reg_out[153]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[153]) );
  DFFRNQ_X1 \Ciphertext_reg[140]  ( .D(reg_out[140]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[140]) );
  DFFRNQ_X1 \Ciphertext_reg[81]  ( .D(reg_out[81]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[81]) );
  DFFRNQ_X1 \Ciphertext_reg[130]  ( .D(reg_out[130]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[130]) );
  DFFRNQ_X1 \Ciphertext_reg[177]  ( .D(reg_out[177]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[177]) );
  DFFRNQ_X1 \Ciphertext_reg[104]  ( .D(reg_out[104]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[104]) );
  DFFRNQ_X1 \Ciphertext_reg[62]  ( .D(reg_out[62]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[62]) );
  DFFRNQ_X1 \Ciphertext_reg[42]  ( .D(reg_out[42]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[42]) );
  DFFRNQ_X1 \Ciphertext_reg[170]  ( .D(reg_out[170]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[170]) );
  DFFRNQ_X1 \Ciphertext_reg[129]  ( .D(reg_out[129]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[129]) );
  DFFRNQ_X1 \Ciphertext_reg[16]  ( .D(reg_out[16]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[16]) );
  DFFRNQ_X1 \Ciphertext_reg[41]  ( .D(reg_out[41]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[41]) );
  DFFRNQ_X1 \Ciphertext_reg[155]  ( .D(reg_out[155]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[155]) );
  DFFRNQ_X1 \Ciphertext_reg[57]  ( .D(reg_out[57]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[57]) );
  DFFRNQ_X1 \Ciphertext_reg[134]  ( .D(reg_out[134]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[134]) );
  DFFRNQ_X1 \Ciphertext_reg[30]  ( .D(reg_out[30]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[30]) );
  DFFRNQ_X1 \Ciphertext_reg[68]  ( .D(reg_out[68]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[68]) );
  DFFRNQ_X1 \Ciphertext_reg[98]  ( .D(reg_out[98]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[98]) );
  DFFRNQ_X1 \Ciphertext_reg[110]  ( .D(reg_out[110]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[110]) );
  DFFRNQ_X1 \Ciphertext_reg[132]  ( .D(reg_out[132]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[132]) );
  DFFRNQ_X1 \Ciphertext_reg[139]  ( .D(reg_out[139]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[139]) );
  DFFRNQ_X1 \Ciphertext_reg[64]  ( .D(reg_out[64]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[64]) );
  DFFRNQ_X1 \Ciphertext_reg[123]  ( .D(reg_out[123]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[123]) );
  DFFRNQ_X1 \Ciphertext_reg[71]  ( .D(reg_out[71]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[71]) );
  DFFRNQ_X1 \Ciphertext_reg[48]  ( .D(reg_out[48]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[48]) );
  DFFRNQ_X1 \Ciphertext_reg[116]  ( .D(reg_out[116]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[116]) );
  DFFRNQ_X1 \Ciphertext_reg[136]  ( .D(reg_out[136]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[136]) );
  DFFRNQ_X1 \Ciphertext_reg[61]  ( .D(reg_out[61]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[61]) );
  DFFRNQ_X1 \Ciphertext_reg[93]  ( .D(reg_out[93]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[93]) );
  DFFRNQ_X1 \Ciphertext_reg[186]  ( .D(reg_out[186]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[186]) );
  DFFRNQ_X1 \Ciphertext_reg[109]  ( .D(reg_out[109]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[109]) );
  DFFRNQ_X1 \Ciphertext_reg[113]  ( .D(reg_out[113]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[113]) );
  DFFRNQ_X1 \Ciphertext_reg[166]  ( .D(reg_out[166]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[166]) );
  DFFRNQ_X1 \Ciphertext_reg[74]  ( .D(reg_out[74]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[74]) );
  DFFRNQ_X1 \Ciphertext_reg[190]  ( .D(reg_out[190]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[190]) );
  DFFRNQ_X1 \Ciphertext_reg[101]  ( .D(reg_out[101]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[101]) );
  DFFRNQ_X1 \Ciphertext_reg[161]  ( .D(reg_out[161]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[161]) );
  DFFRNQ_X1 \Ciphertext_reg[90]  ( .D(reg_out[90]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[90]) );
  DFFRNQ_X1 \Ciphertext_reg[14]  ( .D(reg_out[14]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[14]) );
  DFFRNQ_X1 \Ciphertext_reg[157]  ( .D(reg_out[157]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[157]) );
  DFFRNQ_X1 \Ciphertext_reg[67]  ( .D(reg_out[67]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[67]) );
  DFFRNQ_X1 \Ciphertext_reg[112]  ( .D(reg_out[112]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[112]) );
  DFFRNQ_X1 \Ciphertext_reg[158]  ( .D(reg_out[158]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[158]) );
  DFFRNQ_X1 \Ciphertext_reg[188]  ( .D(reg_out[188]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[188]) );
  DFFRNQ_X1 \Ciphertext_reg[106]  ( .D(reg_out[106]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[106]) );
  DFFRNQ_X1 \Ciphertext_reg[99]  ( .D(reg_out[99]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[99]) );
  DFFRNQ_X1 \Ciphertext_reg[17]  ( .D(reg_out[17]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[17]) );
  DFFRNQ_X1 \Ciphertext_reg[12]  ( .D(reg_out[12]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[12]) );
  DFFRNQ_X1 \Ciphertext_reg[151]  ( .D(reg_out[151]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[151]) );
  DFFRNQ_X1 \Ciphertext_reg[152]  ( .D(reg_out[152]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[152]) );
  DFFRNQ_X1 \Ciphertext_reg[111]  ( .D(reg_out[111]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[111]) );
  DFFRNQ_X1 \Ciphertext_reg[76]  ( .D(reg_out[76]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[76]) );
  DFFRNQ_X1 \Ciphertext_reg[154]  ( .D(reg_out[154]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[154]) );
  DFFRNQ_X1 \Ciphertext_reg[102]  ( .D(reg_out[102]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[102]) );
  DFFRNQ_X1 \Ciphertext_reg[137]  ( .D(reg_out[137]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[137]) );
  DFFRNQ_X1 \Ciphertext_reg[189]  ( .D(reg_out[189]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[189]) );
  DFFRNQ_X1 \Ciphertext_reg[72]  ( .D(reg_out[72]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[72]) );
  DFFRNQ_X1 \Ciphertext_reg[44]  ( .D(reg_out[44]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[44]) );
  DFFRNQ_X1 \Ciphertext_reg[105]  ( .D(reg_out[105]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[105]) );
  DFFRNQ_X1 \Ciphertext_reg[6]  ( .D(reg_out[6]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[6]) );
  DFFRNQ_X1 \Ciphertext_reg[0]  ( .D(reg_out[0]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[0]) );
  DFFRNQ_X1 \Ciphertext_reg[78]  ( .D(reg_out[78]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[78]) );
  DFFRNQ_X1 \Ciphertext_reg[82]  ( .D(reg_out[82]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[82]) );
  DFFRNQ_X1 \Ciphertext_reg[83]  ( .D(reg_out[83]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[83]) );
  DFFRNQ_X1 \Ciphertext_reg[52]  ( .D(reg_out[52]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[52]) );
  DFFRNQ_X1 \Ciphertext_reg[162]  ( .D(reg_out[162]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[162]) );
  DFFRNQ_X1 \Ciphertext_reg[31]  ( .D(reg_out[31]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[31]) );
  DFFRNQ_X1 \Ciphertext_reg[15]  ( .D(reg_out[15]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[15]) );
  DFFRNQ_X1 \Ciphertext_reg[56]  ( .D(reg_out[56]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[56]) );
  DFFRNQ_X1 \Ciphertext_reg[120]  ( .D(reg_out[120]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[120]) );
  DFFRNQ_X1 \Ciphertext_reg[121]  ( .D(reg_out[121]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[121]) );
  DFFRNQ_X1 \Ciphertext_reg[75]  ( .D(reg_out[75]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[75]) );
  DFFRNQ_X1 \Ciphertext_reg[178]  ( .D(reg_out[178]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[178]) );
  DFFRNQ_X1 \Ciphertext_reg[73]  ( .D(reg_out[73]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[73]) );
  DFFRNQ_X1 \Ciphertext_reg[181]  ( .D(reg_out[181]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[181]) );
  DFFRNQ_X1 \Ciphertext_reg[187]  ( .D(reg_out[187]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[187]) );
  DFFRNQ_X1 \Ciphertext_reg[5]  ( .D(reg_out[5]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[5]) );
  DFFRNQ_X1 \Ciphertext_reg[165]  ( .D(reg_out[165]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[165]) );
  DFFRNQ_X1 \Ciphertext_reg[89]  ( .D(reg_out[89]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[89]) );
  DFFRNQ_X1 \Ciphertext_reg[124]  ( .D(reg_out[124]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[124]) );
  DFFRNQ_X1 \Ciphertext_reg[50]  ( .D(reg_out[50]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[50]) );
  DFFRNQ_X1 \Ciphertext_reg[191]  ( .D(reg_out[191]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[191]) );
  DFFRNQ_X1 \Ciphertext_reg[125]  ( .D(reg_out[125]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[125]) );
  DFFRNQ_X1 \Ciphertext_reg[160]  ( .D(reg_out[160]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[160]) );
  DFFRNQ_X1 \Ciphertext_reg[131]  ( .D(reg_out[131]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[131]) );
  DFFRNQ_X1 \Ciphertext_reg[91]  ( .D(reg_out[91]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[91]) );
  DFFRNQ_X1 \Ciphertext_reg[122]  ( .D(reg_out[122]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[122]) );
  DFFRNQ_X1 \Ciphertext_reg[27]  ( .D(reg_out[27]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[27]) );
  DFFRNQ_X1 \Ciphertext_reg[43]  ( .D(reg_out[43]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[43]) );
  DFFRNQ_X1 \Ciphertext_reg[35]  ( .D(reg_out[35]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[35]) );
  DFFRNQ_X1 \Ciphertext_reg[94]  ( .D(reg_out[94]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[94]) );
  DFFRNQ_X1 \Ciphertext_reg[53]  ( .D(reg_out[53]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[53]) );
  DFFRNQ_X1 \Ciphertext_reg[159]  ( .D(reg_out[159]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[159]) );
  DFFRNQ_X1 \Ciphertext_reg[117]  ( .D(reg_out[117]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[117]) );
  DFFRNQ_X1 \Ciphertext_reg[4]  ( .D(reg_out[4]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[4]) );
  DFFRNQ_X1 \Ciphertext_reg[3]  ( .D(reg_out[3]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[3]) );
  DFFRNQ_X1 \Ciphertext_reg[70]  ( .D(reg_out[70]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[70]) );
  DFFRNQ_X1 \Ciphertext_reg[47]  ( .D(reg_out[47]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[47]) );
  DFFRNQ_X1 \Ciphertext_reg[183]  ( .D(reg_out[183]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[183]) );
  DFFRNQ_X1 \Ciphertext_reg[92]  ( .D(reg_out[92]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[92]) );
  DFFRNQ_X1 \Ciphertext_reg[95]  ( .D(reg_out[95]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[95]) );
  DFFRNQ_X1 \Ciphertext_reg[8]  ( .D(reg_out[8]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[8]) );
  DFFRNQ_X1 \Ciphertext_reg[182]  ( .D(reg_out[182]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[182]) );
  DFFRNQ_X1 \Ciphertext_reg[115]  ( .D(reg_out[115]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[115]) );
  DFFRNQ_X1 \Ciphertext_reg[26]  ( .D(reg_out[26]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[26]) );
  DFFRNQ_X1 \Ciphertext_reg[114]  ( .D(reg_out[114]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[114]) );
  DFFRNQ_X1 \Ciphertext_reg[119]  ( .D(reg_out[119]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[119]) );
  DFFRNQ_X1 \Ciphertext_reg[29]  ( .D(reg_out[29]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[29]) );
  DFFRNQ_X1 \Ciphertext_reg[156]  ( .D(reg_out[156]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[156]) );
  DFFRNQ_X1 \Ciphertext_reg[38]  ( .D(reg_out[38]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[38]) );
  DFFRNQ_X1 \Ciphertext_reg[184]  ( .D(reg_out[184]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[184]) );
  DFFRNQ_X1 \Ciphertext_reg[180]  ( .D(reg_out[180]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[180]) );
  DFFRNQ_X1 \Ciphertext_reg[40]  ( .D(reg_out[40]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[40]) );
  DFFRNQ_X1 \Ciphertext_reg[36]  ( .D(reg_out[36]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[36]) );
  DFFRNQ_X1 \Ciphertext_reg[118]  ( .D(reg_out[118]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[118]) );
  DFFRNQ_X1 \Ciphertext_reg[49]  ( .D(reg_out[49]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[49]) );
  DFFRNQ_X1 \Ciphertext_reg[2]  ( .D(reg_out[2]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[2]) );
  DFFRNQ_X1 \Ciphertext_reg[24]  ( .D(reg_out[24]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[24]) );
  DFFRNQ_X1 \Ciphertext_reg[34]  ( .D(reg_out[34]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[34]) );
  DFFRNQ_X1 \Ciphertext_reg[168]  ( .D(reg_out[168]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[168]) );
  DFFRNQ_X1 \Ciphertext_reg[46]  ( .D(reg_out[46]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[46]) );
  DFFRNQ_X1 \Ciphertext_reg[33]  ( .D(reg_out[33]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[33]) );
  DFFRNQ_X1 \Ciphertext_reg[176]  ( .D(reg_out[176]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[176]) );
  DFFRNQ_X1 \Ciphertext_reg[185]  ( .D(reg_out[185]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[185]) );
  DFFRNQ_X1 \Ciphertext_reg[32]  ( .D(reg_out[32]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[32]) );
  DFFRNQ_X1 \Ciphertext_reg[39]  ( .D(reg_out[39]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[39]) );
  DFFRNQ_X1 \Ciphertext_reg[28]  ( .D(reg_out[28]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[28]) );
  DFFRNQ_X1 \Ciphertext_reg[25]  ( .D(reg_out[25]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[25]) );
  SPEEDY_Rounds5_0 SPEEDY_instance ( .Plaintext(reg_in), .Key(reg_key), 
        .Ciphertext(reg_out) );
endmodule

