module SPEEDY_Rounds6_0 ( Plaintext, Key, Ciphertext );
  input [191:0] Plaintext;
  input [191:0] Key;
  output [191:0] Ciphertext;
  wire   n1, n4, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n21, n22, n24,
         n25, n27, n28, n29, n31, n32, n34, n36, n37, n38, n39, n42, n44, n46,
         n47, n50, n51, n52, n53, n54, n57, n60, n61, n62, n66, n67, n71, n72,
         n73, n75, n78, n79, n81, n84, n85, n86, n87, n91, n92, n94, n97, n98,
         n100, n101, n102, n107, n110, n111, n112, n115, n118, n119, n120,
         n123, n124, n125, n128, n135, n136, n137, n138, n139, n144, n146,
         n149, n151, n152, n153, n154, n155, n156, n161, n162, n164, n168,
         n169, n170, n171, n175, n179, n180, n183, n184, n185, n187, n188,
         n193, n196, n204, n205, n206, n207, n210, n214, n215, n219, n221,
         n224, n225, n227, n229, n230, n231, n233, n236, n239, n242, n245,
         n250, n252, n253, n254, n258, n259, n261, n262, n263, n265, n266,
         n268, n270, n273, n274, n275, n276, n277, n279, n281, n283, n284,
         n285, n287, n292, n293, n294, n295, n297, n298, n299, n300, n304,
         n305, n308, n313, n314, n315, n317, n319, n320, n321, n322, n327,
         n328, n329, n330, n335, n337, n338, n339, n342, n343, n347, n348,
         n349, n354, n355, n356, n358, n363, n365, n367, n371, n375, n376,
         n379, n380, n384, n385, n386, n387, n388, n391, n392, n393, n396,
         n397, n398, n400, n401, n402, n405, n406, n408, n410, n412, n413,
         n414, n415, n416, n417, n419, n420, n421, n423, n424, n425, n431,
         n432, n433, n434, n436, n437, n438, n439, n440, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n452, n453, n454, n456, n457,
         n458, n460, n461, n462, n463, n465, n467, n468, n469, n470, n471,
         n474, n475, n476, n477, n478, n479, n480, n481, n485, n487, n488,
         n489, n490, n493, n494, n495, n496, n497, n498, n499, n500, n502,
         n503, n505, n506, n507, n508, n509, n510, n511, n513, n514, n515,
         n516, n517, n518, n519, n521, n522, n524, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n553,
         n554, n556, n560, n561, n562, n563, n564, n565, n567, n568, n570,
         n571, n572, n575, n576, n577, n578, n579, n580, n582, n583, n584,
         n586, n587, n589, n590, n591, n595, n596, n598, n599, n600, n601,
         n602, n603, n606, n607, n609, n610, n612, n613, n615, n616, n618,
         n620, n621, n622, n623, n624, n625, n627, n628, n629, n630, n632,
         n634, n635, n636, n637, n639, n641, n642, n643, n645, n646, n647,
         n651, n652, n654, n655, n657, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n671, n673, n675, n676, n678, n679, n680, n681,
         n686, n689, n690, n691, n692, n693, n694, n695, n696, n698, n699,
         n700, n701, n702, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n721, n722, n723, n724,
         n725, n727, n728, n729, n730, n732, n733, n734, n736, n737, n738,
         n739, n741, n742, n743, n744, n745, n746, n747, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n760, n761, n763, n764,
         n765, n767, n769, n770, n772, n773, n776, n777, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n801, n802, n803, n805, n806,
         n808, n809, n810, n812, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n836, n837, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n855, n856, n857, n858,
         n859, n861, n862, n864, n865, n867, n868, n870, n871, n873, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n893, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n924, n925, n926, n927, n929, n930, n931, n932, n933, n935,
         n936, n937, n938, n939, n940, n941, n942, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n972, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n985, n986, n987, n989, n990, n992, n994, n995, n996, n998,
         n1000, n1001, n1003, n1004, n1007, n1008, n1009, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1022, n1023, n1024, n1026,
         n1028, n1030, n1032, n1034, n1035, n1036, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1059, n1060, n1063, n1064, n1065,
         n1067, n1069, n1070, n1071, n1074, n1075, n1076, n1077, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1092, n1093, n1094, n1096, n1098, n1099, n1100, n1101, n1102, n1104,
         n1106, n1107, n1108, n1109, n1112, n1113, n1116, n1117, n1119, n1120,
         n1122, n1124, n1125, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1145, n1146, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1172, n1173, n1175, n1177, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1196, n1197, n1198, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1211, n1212, n1213, n1214,
         n1215, n1216, n1218, n1219, n1221, n1223, n1224, n1225, n1226, n1227,
         n1228, n1230, n1231, n1232, n1233, n1235, n1237, n1238, n1239, n1240,
         n1241, n1243, n1244, n1245, n1246, n1247, n1249, n1250, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1269, n1271, n1274, n1275, n1277, n1278,
         n1279, n1280, n1281, n1282, n1284, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1294, n1296, n1297, n1298, n1299, n1300, n1302, n1303,
         n1305, n1306, n1307, n1308, n1309, n1310, n1312, n1313, n1315, n1316,
         n1317, n1318, n1319, n1321, n1322, n1323, n1325, n1326, n1327, n1328,
         n1329, n1331, n1332, n1333, n1334, n1335, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1372, n1373, n1374, n1376, n1377, n1378, n1379, n1380, n1382, n1384,
         n1385, n1386, n1387, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1402, n1403, n1404, n1405, n1406, n1407, n1409,
         n1410, n1411, n1413, n1414, n1415, n1416, n1417, n1419, n1420, n1421,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1436, n1438, n1439, n1441, n1445, n1446, n1449, n1450,
         n1451, n1452, n1453, n1454, n1456, n1457, n1458, n1462, n1463, n1464,
         n1465, n1466, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1489, n1490,
         n1491, n1492, n1494, n1496, n1497, n1499, n1500, n1504, n1506, n1507,
         n1508, n1511, n1513, n1516, n1519, n1521, n1522, n1523, n1524, n1525,
         n1528, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1540,
         n1541, n1543, n1544, n1545, n1546, n1547, n1549, n1550, n1553, n1555,
         n1557, n1559, n1560, n1561, n1563, n1564, n1565, n1567, n1571, n1572,
         n1573, n1577, n1579, n1580, n1581, n1587, n1588, n1589, n1590, n1592,
         n1594, n1595, n1596, n1597, n1600, n1601, n1602, n1603, n1604, n1607,
         n1609, n1610, n1612, n1613, n1615, n1616, n1617, n1619, n1620, n1621,
         n1622, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1640, n1641, n1642, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1658, n1659, n1661, n1663,
         n1664, n1668, n1669, n1671, n1672, n1673, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1690,
         n1694, n1695, n1696, n1698, n1699, n1700, n1702, n1703, n1704, n1707,
         n1708, n1709, n1710, n1712, n1713, n1714, n1716, n1718, n1719, n1720,
         n1726, n1727, n1728, n1730, n1731, n1732, n1733, n1734, n1736, n1741,
         n1742, n1745, n1746, n1749, n1751, n1756, n1757, n1758, n1760, n1761,
         n1762, n1763, n1764, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1778, n1779, n1780, n1781, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1791, n1792, n1793, n1794, n1795,
         n1796, n1799, n1800, n1801, n1803, n1805, n1807, n1808, n1811, n1812,
         n1813, n1814, n1815, n1816, n1818, n1819, n1820, n1825, n1826, n1828,
         n1830, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1842, n1844,
         n1845, n1848, n1850, n1851, n1853, n1857, n1858, n1859, n1861, n1862,
         n1863, n1864, n1865, n1867, n1868, n1869, n1870, n1871, n1873, n1874,
         n1875, n1876, n1877, n1878, n1881, n1882, n1883, n1884, n1886, n1887,
         n1889, n1890, n1892, n1896, n1897, n1898, n1900, n1902, n1903, n1905,
         n1908, n1909, n1910, n1911, n1913, n1914, n1915, n1916, n1917, n1920,
         n1923, n1926, n1927, n1928, n1929, n1930, n1931, n1933, n1934, n1935,
         n1936, n1937, n1938, n1940, n1941, n1942, n1944, n1945, n1946, n1948,
         n1949, n1950, n1951, n1954, n1955, n1956, n1957, n1960, n1961, n1962,
         n1963, n1964, n1965, n1967, n1968, n1970, n1971, n1973, n1974, n1976,
         n1978, n1979, n1980, n1982, n1983, n1984, n1986, n1988, n1990, n1991,
         n1992, n1993, n1994, n1995, n1997, n1998, n2000, n2001, n2002, n2003,
         n2004, n2005, n2009, n2012, n2013, n2015, n2016, n2017, n2018, n2019,
         n2021, n2022, n2023, n2024, n2028, n2029, n2031, n2032, n2036, n2037,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2048, n2049, n2052,
         n2053, n2054, n2055, n2060, n2061, n2064, n2066, n2069, n2070, n2072,
         n2073, n2074, n2075, n2076, n2078, n2080, n2081, n2082, n2084, n2085,
         n2086, n2088, n2089, n2092, n2095, n2097, n2098, n2099, n2100, n2101,
         n2103, n2104, n2105, n2107, n2108, n2111, n2112, n2113, n2114, n2117,
         n2118, n2122, n2123, n2124, n2125, n2126, n2128, n2129, n2130, n2132,
         n2134, n2135, n2137, n2138, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2152, n2153, n2154, n2155, n2156, n2158,
         n2161, n2162, n2163, n2164, n2166, n2167, n2169, n2172, n2173, n2174,
         n2176, n2177, n2178, n2180, n2182, n2186, n2190, n2191, n2192, n2197,
         n2198, n2200, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2214, n2215, n2217, n2219, n2221, n2222, n2225,
         n2226, n2229, n2230, n2233, n2234, n2236, n2237, n2239, n2241, n2242,
         n2245, n2247, n2250, n2251, n2252, n2253, n2256, n2257, n2258, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2270, n2271, n2272,
         n2275, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2285, n2288,
         n2289, n2290, n2291, n2292, n2293, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2304, n2305, n2306, n2308, n2309, n2311, n2312, n2315,
         n2316, n2317, n2318, n2319, n2320, n2324, n2325, n2330, n2331, n2333,
         n2334, n2335, n2337, n2338, n2339, n2342, n2345, n2347, n2348, n2349,
         n2351, n2352, n2353, n2355, n2356, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2375, n2378, n2380,
         n2381, n2383, n2384, n2386, n2387, n2388, n2389, n2390, n2391, n2393,
         n2394, n2395, n2396, n2398, n2400, n2401, n2404, n2405, n2407, n2408,
         n2409, n2410, n2411, n2412, n2414, n2415, n2417, n2418, n2420, n2421,
         n2423, n2424, n2427, n2430, n2432, n2435, n2436, n2440, n2441, n2442,
         n2443, n2444, n2447, n2448, n2449, n2450, n2452, n2455, n2456, n2458,
         n2460, n2463, n2464, n2466, n2468, n2469, n2470, n2471, n2472, n2473,
         n2476, n2477, n2479, n2480, n2483, n2484, n2486, n2489, n2490, n2491,
         n2492, n2495, n2497, n2498, n2499, n2500, n2501, n2502, n2507, n2508,
         n2509, n2512, n2513, n2514, n2517, n2518, n2519, n2520, n2522, n2523,
         n2524, n2525, n2526, n2529, n2534, n2535, n2536, n2537, n2538, n2539,
         n2547, n2548, n2549, n2550, n2551, n2554, n2556, n2557, n2558, n2560,
         n2561, n2563, n2564, n2565, n2566, n2568, n2569, n2570, n2574, n2575,
         n2576, n2577, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2587,
         n2589, n2590, n2591, n2592, n2593, n2595, n2596, n2598, n2599, n2600,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2616, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2628, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2642, n2643, n2646, n2647, n2648, n2649,
         n2650, n2651, n2653, n2654, n2655, n2656, n2657, n2661, n2664, n2665,
         n2666, n2667, n2668, n2671, n2672, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2682, n2683, n2684, n2686, n2687, n2689, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2712, n2713, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2724, n2725, n2726, n2727, n2728,
         n2729, n2731, n2732, n2733, n2734, n2738, n2739, n2741, n2743, n2744,
         n2745, n2746, n2747, n2750, n2752, n2753, n2754, n2756, n2757, n2758,
         n2759, n2761, n2763, n2764, n2766, n2767, n2770, n2771, n2773, n2775,
         n2777, n2778, n2780, n2784, n2785, n2786, n2788, n2789, n2790, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2801, n2802, n2803, n2808,
         n2809, n2812, n2813, n2818, n2819, n2820, n2821, n2822, n2824, n2825,
         n2826, n2831, n2833, n2834, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2847, n2848, n2849, n2851, n2852, n2853, n2854, n2855,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2883, n2886, n2888, n2889, n2890, n2891, n2894,
         n2896, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2908, n2909, n2911, n2912, n2913, n2915, n2917, n2918, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2933,
         n2934, n2935, n2936, n2937, n2939, n2940, n2941, n2943, n2944, n2945,
         n2946, n2948, n2949, n2951, n2952, n2953, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2964, n2965, n2967, n2968, n2969, n2970, n2971,
         n2972, n2974, n2975, n2976, n2978, n2980, n2981, n2982, n2983, n2986,
         n2987, n2989, n2990, n2992, n2993, n2996, n2997, n2998, n2999, n3001,
         n3003, n3004, n3005, n3006, n3007, n3009, n3010, n3012, n3013, n3014,
         n3016, n3018, n3019, n3021, n3022, n3023, n3024, n3026, n3027, n3028,
         n3030, n3032, n3033, n3035, n3036, n3038, n3039, n3041, n3042, n3043,
         n3045, n3047, n3048, n3049, n3050, n3051, n3052, n3055, n3056, n3057,
         n3059, n3060, n3061, n3063, n3065, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3076, n3077, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3090, n3091, n3092, n3093, n3094, n3096, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3109, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3122, n3123,
         n3124, n3126, n3128, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3140, n3142, n3143, n3144, n3146, n3147, n3148, n3149, n3152, n3155,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3168, n3169, n3170, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3183, n3184, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3211, n3212,
         n3213, n3214, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3247, n3248, n3250, n3251, n3253, n3255, n3256, n3257, n3258, n3259,
         n3260, n3266, n3267, n3269, n3270, n3271, n3272, n3275, n3280, n3281,
         n3282, n3283, n3285, n3286, n3288, n3289, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3300, n3303, n3304, n3305, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3322, n3324, n3325, n3327, n3328, n3329, n3332, n3334, n3336, n3339,
         n3340, n3341, n3343, n3344, n3345, n3348, n3350, n3351, n3352, n3353,
         n3354, n3355, n3357, n3358, n3360, n3361, n3364, n3365, n3366, n3368,
         n3369, n3371, n3375, n3376, n3378, n3379, n3380, n3382, n3384, n3385,
         n3388, n3389, n3390, n3391, n3392, n3393, n3395, n3396, n3399, n3401,
         n3402, n3403, n3405, n3407, n3408, n3410, n3411, n3412, n3415, n3416,
         n3417, n3418, n3420, n3421, n3424, n3425, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3439, n3440, n3441, n3442,
         n3443, n3445, n3446, n3447, n3448, n3449, n3451, n3454, n3455, n3461,
         n3462, n3463, n3465, n3467, n3468, n3469, n3472, n3475, n3476, n3477,
         n3480, n3481, n3482, n3483, n3484, n3486, n3487, n3489, n3491, n3493,
         n3494, n3495, n3497, n3499, n3501, n3502, n3503, n3504, n3506, n3508,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3525, n3526, n3527, n3529, n3530, n3535, n3536, n3539,
         n3540, n3541, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3552,
         n3553, n3554, n3556, n3558, n3559, n3562, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3574, n3575, n3576, n3578, n3579, n3580, n3581,
         n3583, n3584, n3586, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3596, n3597, n3598, n3599, n3600, n3601, n3603, n3604, n3605, n3606,
         n3614, n3617, n3618, n3619, n3620, n3621, n3622, n3624, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3638, n3639,
         n3643, n3644, n3646, n3648, n3650, n3651, n3652, n3653, n3654, n3656,
         n3657, n3658, n3659, n3663, n3665, n3667, n3668, n3669, n3670, n3672,
         n3673, n3677, n3678, n3680, n3682, n3683, n3685, n3686, n3687, n3689,
         n3692, n3694, n3695, n3696, n3698, n3702, n3703, n3704, n3705, n3706,
         n3708, n3711, n3717, n3718, n3722, n3723, n3724, n3725, n3727, n3728,
         n3729, n3730, n3731, n3732, n3735, n3736, n3737, n3739, n3742, n3744,
         n3746, n3748, n3750, n3751, n3755, n3756, n3757, n3759, n3760, n3767,
         n3769, n3770, n3771, n3772, n3773, n3774, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3786, n3787, n3788, n3790, n3791, n3792,
         n3793, n3794, n3796, n3797, n3798, n3799, n3800, n3801, n3807, n3809,
         n3810, n3812, n3815, n3816, n3819, n3820, n3821, n3822, n3824, n3825,
         n3826, n3827, n3828, n3830, n3835, n3836, n3840, n3842, n3843, n3844,
         n3845, n3846, n3847, n3851, n3852, n3854, n3856, n3860, n3861, n3862,
         n3866, n3867, n3868, n3870, n3873, n3874, n3879, n3880, n3883, n3884,
         n3885, n3888, n3889, n3891, n3893, n3894, n3896, n3898, n3900, n3901,
         n3902, n3903, n3904, n3905, n3908, n3909, n3911, n3915, n3916, n3918,
         n3919, n3920, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3940, n3941,
         n3944, n3945, n3946, n3947, n3950, n3951, n3954, n3955, n3957, n3958,
         n3962, n3963, n3964, n3967, n3970, n3972, n3973, n3977, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4003, n4004, n4006,
         n4008, n4013, n4014, n4015, n4016, n4017, n4019, n4020, n4021, n4024,
         n4025, n4026, n4028, n4029, n4034, n4035, n4036, n4040, n4041, n4042,
         n4043, n4045, n4047, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4059, n4060, n4061, n4062, n4063, n4065, n4066, n4067,
         n4069, n4070, n4071, n4075, n4076, n4077, n4079, n4082, n4084, n4086,
         n4087, n4088, n4089, n4091, n4095, n4097, n4098, n4099, n4100, n4101,
         n4102, n4106, n4107, n4110, n4111, n4112, n4113, n4114, n4117, n4118,
         n4119, n4123, n4124, n4130, n4131, n4133, n4134, n4135, n4136, n4140,
         n4142, n4143, n4145, n4146, n4150, n4151, n4154, n4155, n4156, n4157,
         n4158, n4161, n4162, n4163, n4164, n4167, n4168, n4169, n4173, n4174,
         n4176, n4177, n4178, n4179, n4180, n4182, n4183, n4184, n4186, n4187,
         n4188, n4191, n4192, n4193, n4194, n4196, n4197, n4200, n4201, n4202,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4224, n4225, n4226,
         n4228, n4230, n4231, n4232, n4233, n4234, n4236, n4240, n4241, n4243,
         n4244, n4245, n4246, n4248, n4251, n4253, n4254, n4255, n4259, n4260,
         n4261, n4262, n4263, n4266, n4267, n4268, n4269, n4273, n4274, n4279,
         n4280, n4281, n4283, n4284, n4285, n4286, n4287, n4289, n4290, n4291,
         n4293, n4295, n4299, n4300, n4301, n4302, n4305, n4306, n4308, n4310,
         n4311, n4312, n4314, n4315, n4318, n4319, n4321, n4324, n4325, n4327,
         n4329, n4330, n4331, n4332, n4335, n4337, n4338, n4339, n4340, n4341,
         n4342, n4349, n4350, n4352, n4353, n4354, n4355, n4356, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4370,
         n4371, n4373, n4374, n4375, n4378, n4379, n4380, n4381, n4382, n4384,
         n4385, n4386, n4387, n4390, n4391, n4392, n4393, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4403, n4405, n4407, n4408, n4409, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4422,
         n4423, n4425, n4427, n4432, n4433, n4434, n4435, n4436, n4437, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4456, n4458, n4459, n4460, n4464, n4465, n4466, n4467,
         n4468, n4469, n4471, n4472, n4474, n4476, n4477, n4481, n4483, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4494, n4496, n4497, n4498,
         n4500, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4510, n4511,
         n4514, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4524, n4525,
         n4529, n4530, n4531, n4533, n4534, n4535, n4536, n4538, n4539, n4542,
         n4543, n4547, n4550, n4551, n4552, n4554, n4555, n4556, n4557, n4559,
         n4560, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4571,
         n4572, n4574, n4577, n4578, n4579, n4580, n4581, n4583, n4585, n4586,
         n4587, n4589, n4590, n4591, n4592, n4594, n4595, n4596, n4599, n4601,
         n4602, n4604, n4607, n4609, n4610, n4611, n4613, n4614, n4616, n4617,
         n4618, n4619, n4622, n4624, n4626, n4627, n4628, n4629, n4631, n4632,
         n4633, n4635, n4636, n4637, n4638, n4639, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4655, n4656, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4668, n4669, n4671,
         n4672, n4674, n4675, n4677, n4678, n4680, n4681, n4682, n4683, n4685,
         n4686, n4687, n4688, n4689, n4693, n4699, n4700, n4701, n4704, n4706,
         n4708, n4709, n4710, n4711, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4739, n4740, n4741, n4743, n4744,
         n4746, n4747, n4749, n4750, n4755, n4756, n4758, n4759, n4760, n4761,
         n4762, n4763, n4765, n4767, n4768, n4769, n4770, n4771, n4772, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4788, n4789, n4790, n4791, n4792, n4794, n4797, n4798,
         n4800, n4801, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4814, n4816, n4820, n4821, n4822, n4823, n4824, n4831,
         n4833, n4834, n4835, n4840, n4841, n4842, n4843, n4845, n4846, n4847,
         n4849, n4850, n4854, n4855, n4856, n4857, n4858, n4859, n4861, n4862,
         n4863, n4865, n4867, n4868, n4869, n4871, n4872, n4873, n4878, n4879,
         n4880, n4881, n4883, n4884, n4885, n4886, n4891, n4892, n4893, n4894,
         n4895, n4897, n4898, n4899, n4900, n4903, n4906, n4908, n4909, n4913,
         n4914, n4915, n4916, n4918, n4919, n4920, n4922, n4925, n4926, n4927,
         n4928, n4930, n4931, n4932, n4935, n4936, n4937, n4938, n4942, n4944,
         n4949, n4951, n4952, n4953, n4955, n4956, n4959, n4960, n4961, n4964,
         n4965, n4967, n4968, n4971, n4972, n4975, n4976, n4980, n4982, n4983,
         n4984, n4985, n4986, n4988, n4989, n4991, n4992, n4993, n4994, n4996,
         n4997, n4999, n5000, n5002, n5003, n5004, n5009, n5011, n5012, n5013,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5038,
         n5039, n5040, n5041, n5043, n5045, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5058, n5059, n5061, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5086, n5089, n5090, n5091, n5092,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5103, n5104, n5105,
         n5106, n5107, n5109, n5111, n5112, n5113, n5115, n5116, n5118, n5119,
         n5121, n5122, n5124, n5126, n5127, n5128, n5129, n5130, n5132, n5133,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5154, n5155, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5166, n5169, n5170, n5172, n5173, n5174,
         n5177, n5178, n5182, n5184, n5185, n5186, n5187, n5188, n5190, n5191,
         n5194, n5196, n5197, n5199, n5202, n5203, n5205, n5206, n5207, n5209,
         n5210, n5211, n5212, n5215, n5216, n5217, n5218, n5219, n5221, n5222,
         n5223, n5225, n5226, n5227, n5228, n5229, n5231, n5233, n5236, n5237,
         n5238, n5239, n5240, n5241, n5243, n5244, n5248, n5250, n5252, n5253,
         n5254, n5255, n5256, n5258, n5259, n5260, n5261, n5263, n5264, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5277,
         n5278, n5279, n5280, n5282, n5284, n5286, n5287, n5288, n5289, n5292,
         n5296, n5297, n5300, n5301, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5311, n5314, n5315, n5316, n5317, n5318, n5321, n5322, n5324,
         n5327, n5328, n5329, n5332, n5333, n5335, n5336, n5337, n5338, n5339,
         n5340, n5342, n5343, n5345, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5356, n5357, n5358, n5361, n5366, n5367, n5371, n5372, n5373,
         n5374, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5387, n5389, n5392, n5394, n5395, n5396, n5399, n5400, n5401,
         n5402, n5405, n5407, n5408, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5421, n5422, n5424, n5425, n5428, n5429, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5440, n5441, n5445,
         n5448, n5449, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5462, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5476, n5477, n5478, n5480, n5481, n5482, n5483, n5484,
         n5485, n5487, n5488, n5490, n5491, n5492, n5494, n5495, n5496, n5497,
         n5498, n5500, n5501, n5503, n5504, n5505, n5508, n5509, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5520, n5522, n5523, n5525,
         n5526, n5527, n5529, n5530, n5532, n5533, n5534, n5535, n5539, n5543,
         n5544, n5545, n5546, n5548, n5549, n5550, n5553, n5555, n5556, n5558,
         n5560, n5561, n5562, n5563, n5568, n5570, n5571, n5572, n5573, n5575,
         n5577, n5578, n5581, n5582, n5583, n5586, n5587, n5588, n5589, n5590,
         n5592, n5593, n5594, n5595, n5597, n5598, n5600, n5601, n5602, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5615, n5616,
         n5618, n5619, n5620, n5621, n5622, n5624, n5625, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5640,
         n5641, n5642, n5644, n5645, n5646, n5647, n5648, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5662, n5663, n5666, n5668, n5669, n5670,
         n5671, n5672, n5673, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5687, n5689, n5690, n5691, n5692, n5693,
         n5694, n5696, n5697, n5698, n5699, n5700, n5702, n5703, n5704, n5707,
         n5708, n5709, n5710, n5712, n5713, n5714, n5717, n5718, n5722, n5724,
         n5725, n5726, n5730, n5732, n5733, n5734, n5735, n5736, n5737, n5741,
         n5742, n5743, n5744, n5745, n5748, n5751, n5752, n5753, n5754, n5755,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5779, n5781, n5782, n5784, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5795, n5796, n5801, n5804, n5805, n5810, n5812, n5813,
         n5814, n5817, n5820, n5821, n5822, n5825, n5826, n5827, n5828, n5830,
         n5832, n5834, n5835, n5836, n5837, n5838, n5839, n5842, n5843, n5844,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5869,
         n5870, n5871, n5872, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5888, n5889, n5890, n5891,
         n5892, n5893, n5895, n5896, n5897, n5900, n5901, n5903, n5904, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5925, n5926, n5929, n5930, n5931,
         n5932, n5933, n5935, n5936, n5937, n5939, n5940, n5941, n5942, n5944,
         n5945, n5946, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5958,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5968, n5969, n5970,
         n5971, n5972, n5973, n5975, n5976, n5978, n5979, n5980, n5981, n5982,
         n5983, n5988, n5989, n5990, n5991, n5993, n5994, n5995, n5996, n5997,
         n5999, n6001, n6003, n6005, n6006, n6007, n6008, n6009, n6010, n6012,
         n6013, n6014, n6016, n6018, n6020, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6037,
         n6039, n6041, n6042, n6043, n6047, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6058, n6059, n6061, n6062, n6063, n6064, n6067, n6068,
         n6069, n6071, n6072, n6073, n6074, n6075, n6076, n6078, n6079, n6081,
         n6082, n6083, n6086, n6087, n6088, n6090, n6091, n6092, n6093, n6094,
         n6095, n6097, n6098, n6099, n6101, n6102, n6103, n6104, n6105, n6106,
         n6108, n6109, n6110, n6111, n6114, n6115, n6116, n6117, n6118, n6119,
         n6121, n6123, n6127, n6129, n6131, n6132, n6133, n6134, n6138, n6142,
         n6143, n6144, n6145, n6146, n6148, n6149, n6150, n6151, n6152, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6165, n6166,
         n6167, n6168, n6169, n6170, n6172, n6173, n6175, n6176, n6177, n6178,
         n6179, n6181, n6182, n6183, n6185, n6186, n6187, n6188, n6189, n6190,
         n6192, n6193, n6198, n6199, n6200, n6203, n6204, n6205, n6206, n6207,
         n6209, n6211, n6212, n6213, n6215, n6216, n6218, n6219, n6221, n6223,
         n6225, n6227, n6228, n6229, n6230, n6231, n6232, n6234, n6235, n6236,
         n6237, n6238, n6242, n6244, n6245, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6259, n6262, n6263, n6265,
         n6266, n6267, n6268, n6272, n6273, n6275, n6277, n6280, n6281, n6282,
         n6283, n6285, n6286, n6287, n6288, n6290, n6293, n6294, n6295, n6297,
         n6298, n6299, n6300, n6303, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6316, n6318, n6319, n6320, n6321, n6322, n6324, n6325, n6326,
         n6327, n6328, n6329, n6332, n6334, n6336, n6337, n6338, n6341, n6342,
         n6343, n6344, n6345, n6346, n6348, n6350, n6351, n6354, n6357, n6359,
         n6360, n6362, n6363, n6364, n6365, n6366, n6369, n6370, n6371, n6373,
         n6376, n6377, n6380, n6382, n6384, n6386, n6387, n6388, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6405, n6407, n6408, n6409, n6411, n6414, n6416, n6417, n6420, n6421,
         n6424, n6425, n6426, n6427, n6428, n6429, n6431, n6432, n6433, n6434,
         n6435, n6440, n6442, n6444, n6445, n6446, n6447, n6451, n6452, n6453,
         n6454, n6455, n6457, n6458, n6461, n6462, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6482, n6483, n6484, n6485, n6488, n6489, n6490, n6491, n6493,
         n6494, n6497, n6500, n6501, n6502, n6503, n6504, n6505, n6507, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6519, n6520, n6524, n6526,
         n6530, n6531, n6532, n6533, n6536, n6539, n6540, n6543, n6544, n6545,
         n6547, n6548, n6549, n6551, n6552, n6553, n6555, n6556, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6584, n6587, n6590, n6591, n6592, n6593, n6595, n6597, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6607, n6608, n6609, n6610, n6611,
         n6612, n6614, n6615, n6616, n6618, n6619, n6620, n6621, n6624, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6637, n6638,
         n6639, n6640, n6641, n6643, n6644, n6645, n6646, n6647, n6649, n6650,
         n6651, n6654, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6666, n6667, n6668, n6669, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6691, n6693, n6694, n6696, n6698, n6699, n6700,
         n6701, n6702, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6716, n6718, n6719, n6720, n6721, n6722, n6723, n6725,
         n6726, n6728, n6730, n6731, n6733, n6735, n6737, n6739, n6741, n6743,
         n6745, n6746, n6748, n6749, n6750, n6751, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6775, n6776, n6777,
         n6778, n6779, n6780, n6782, n6783, n6784, n6786, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6797, n6798, n6799, n6800, n6801, n6802,
         n6807, n6808, n6809, n6810, n6811, n6812, n6814, n6816, n6817, n6818,
         n6819, n6820, n6822, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6833, n6835, n6836, n6837, n6840, n6841, n6842, n6843, n6846,
         n6848, n6849, n6850, n6851, n6852, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6862, n6863, n6864, n6865, n6866, n6867, n6869, n6872,
         n6873, n6874, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6893, n6894, n6895, n6897,
         n6898, n6899, n6901, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6913, n6914, n6915, n6918, n6919, n6920, n6921, n6923,
         n6924, n6925, n6926, n6929, n6930, n6931, n6932, n6935, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6945, n6948, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6973, n6974, n6975,
         n6976, n6978, n6980, n6981, n6982, n6985, n6990, n6992, n6994, n6995,
         n6996, n6997, n6999, n7001, n7003, n7004, n7005, n7007, n7008, n7011,
         n7012, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7022, n7023,
         n7024, n7025, n7027, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7059, n7060, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7080, n7081,
         n7083, n7084, n7085, n7086, n7087, n7088, n7090, n7091, n7093, n7094,
         n7095, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7105, n7107,
         n7108, n7109, n7110, n7113, n7114, n7115, n7116, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7129, n7131, n7132, n7133,
         n7134, n7135, n7137, n7138, n7139, n7140, n7141, n7143, n7144, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7157, n7160,
         n7161, n7162, n7163, n7164, n7167, n7169, n7170, n7171, n7173, n7176,
         n7178, n7179, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7190, n7191, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7203, n7204, n7205, n7206, n7207, n7211, n7212, n7213, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7224, n7225, n7226, n7228,
         n7229, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7244, n7245, n7246, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7261, n7262, n7263, n7265, n7266,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7307, n7308, n7309,
         n7310, n7312, n7316, n7317, n7318, n7319, n7320, n7323, n7324, n7325,
         n7326, n7327, n7328, n7330, n7331, n7332, n7334, n7335, n7336, n7339,
         n7341, n7343, n7344, n7345, n7348, n7349, n7350, n7352, n7356, n7357,
         n7358, n7360, n7361, n7363, n7365, n7366, n7368, n7369, n7370, n7371,
         n7373, n7374, n7375, n7376, n7377, n7378, n7380, n7381, n7382, n7383,
         n7384, n7386, n7387, n7388, n7392, n7394, n7395, n7396, n7397, n7398,
         n7400, n7402, n7403, n7406, n7407, n7411, n7412, n7413, n7415, n7417,
         n7418, n7419, n7420, n7425, n7426, n7427, n7429, n7430, n7431, n7432,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7444, n7446, n7447,
         n7450, n7452, n7453, n7454, n7457, n7458, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7483, n7485, n7486, n7488,
         n7490, n7492, n7493, n7495, n7496, n7497, n7501, n7502, n7503, n7504,
         n7505, n7511, n7512, n7513, n7515, n7516, n7517, n7518, n7520, n7524,
         n7525, n7526, n7528, n7529, n7530, n7532, n7535, n7537, n7538, n7541,
         n7543, n7544, n7545, n7546, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7557, n7559, n7560, n7561, n7562, n7565, n7566, n7568, n7569,
         n7570, n7572, n7573, n7574, n7575, n7576, n7577, n7579, n7580, n7581,
         n7582, n7584, n7586, n7589, n7590, n7591, n7592, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7602, n7603, n7604, n7605, n7606, n7607,
         n7609, n7610, n7611, n7613, n7614, n7615, n7616, n7619, n7620, n7622,
         n7623, n7624, n7625, n7626, n7628, n7630, n7631, n7633, n7634, n7635,
         n7636, n7638, n7639, n7640, n7641, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7651, n7652, n7653, n7655, n7656, n7657, n7658, n7659,
         n7660, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7693, n7694, n7695,
         n7698, n7699, n7700, n7701, n7702, n7703, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7716, n7717, n7719, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7729, n7730, n7731, n7732,
         n7733, n7736, n7737, n7738, n7741, n7744, n7745, n7746, n7747, n7748,
         n7749, n7751, n7753, n7754, n7756, n7757, n7759, n7761, n7762, n7765,
         n7767, n7768, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7785, n7786, n7787, n7789, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7802, n7803, n7804,
         n7806, n7808, n7809, n7810, n7811, n7813, n7815, n7817, n7819, n7820,
         n7822, n7823, n7825, n7826, n7828, n7829, n7830, n7831, n7832, n7834,
         n7836, n7837, n7838, n7839, n7842, n7843, n7845, n7848, n7850, n7851,
         n7852, n7853, n7854, n7855, n7857, n7859, n7860, n7861, n7862, n7865,
         n7866, n7867, n7868, n7870, n7871, n7872, n7873, n7874, n7875, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7904, n7905, n7908, n7909, n7910, n7911, n7912, n7913, n7915, n7916,
         n7917, n7918, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7928,
         n7929, n7931, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7945, n7946, n7947, n7949, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7971, n7973, n7974, n7977, n7978, n7984,
         n7986, n7987, n7988, n7989, n7990, n7991, n7993, n7994, n7995, n7997,
         n7998, n7999, n8000, n8001, n8003, n8004, n8005, n8006, n8007, n8010,
         n8011, n8012, n8013, n8015, n8016, n8018, n8020, n8021, n8022, n8024,
         n8026, n8028, n8029, n8030, n8031, n8033, n8035, n8036, n8037, n8038,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8049, n8050, n8051,
         n8053, n8054, n8055, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8073, n8074,
         n8076, n8077, n8078, n8079, n8081, n8082, n8083, n8084, n8086, n8087,
         n8088, n8089, n8091, n8092, n8093, n8094, n8095, n8098, n8099, n8100,
         n8105, n8106, n8107, n8108, n8109, n8110, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8125, n8126, n8127,
         n8129, n8130, n8131, n8132, n8133, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8152, n8154, n8156, n8160, n8164, n8165, n8166, n8167, n8168, n8170,
         n8171, n8174, n8175, n8176, n8178, n8181, n8182, n8183, n8184, n8186,
         n8189, n8190, n8192, n8193, n8194, n8195, n8196, n8197, n8199, n8200,
         n8201, n8202, n8203, n8204, n8206, n8207, n8208, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8219, n8222, n8226, n8227, n8228,
         n8230, n8232, n8233, n8235, n8236, n8237, n8238, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8251, n8252, n8253, n8256,
         n8257, n8258, n8259, n8260, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8282, n8283, n8284, n8285, n8286, n8287, n8290, n8291, n8292, n8293,
         n8294, n8295, n8298, n8299, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8312, n8313, n8314, n8315, n8317, n8318, n8320,
         n8323, n8324, n8325, n8327, n8328, n8330, n8331, n8332, n8334, n8335,
         n8336, n8337, n8339, n8340, n8341, n8343, n8344, n8345, n8347, n8348,
         n8349, n8352, n8353, n8354, n8356, n8358, n8359, n8360, n8361, n8364,
         n8365, n8366, n8370, n8371, n8372, n8373, n8374, n8376, n8378, n8379,
         n8380, n8381, n8382, n8383, n8386, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8405, n8406,
         n8408, n8409, n8411, n8412, n8413, n8415, n8416, n8418, n8420, n8421,
         n8422, n8424, n8425, n8427, n8431, n8432, n8433, n8434, n8435, n8437,
         n8438, n8440, n8442, n8443, n8444, n8450, n8452, n8453, n8454, n8455,
         n8456, n8457, n8459, n8461, n8463, n8464, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8475, n8478, n8479, n8480, n8481, n8482,
         n8485, n8487, n8488, n8489, n8490, n8491, n8492, n8494, n8496, n8497,
         n8499, n8500, n8502, n8504, n8505, n8506, n8507, n8515, n8519, n8522,
         n8523, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8535, n8536, n8537, n8539, n8541, n8542, n8543, n8544, n8545, n8547,
         n8548, n8549, n8550, n8551, n8553, n8554, n8555, n8556, n8557, n8558,
         n8560, n8561, n8562, n8567, n8568, n8569, n8570, n8571, n8573, n8575,
         n8576, n8577, n8578, n8579, n8581, n8582, n8583, n8584, n8587, n8589,
         n8591, n8592, n8593, n8594, n8595, n8596, n8601, n8602, n8603, n8604,
         n8605, n8606, n8608, n8609, n8611, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8622, n8625, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8639, n8645, n8648, n8650, n8651,
         n8653, n8654, n8655, n8656, n8657, n8659, n8662, n8663, n8664, n8665,
         n8666, n8667, n8671, n8672, n8674, n8675, n8676, n8678, n8680, n8681,
         n8682, n8683, n8684, n8685, n8687, n8689, n8691, n8692, n8694, n8695,
         n8700, n8701, n8702, n8703, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8726, n8727, n8728, n8731, n8733, n8734, n8735,
         n8736, n8737, n8739, n8740, n8741, n8742, n8743, n8745, n8746, n8747,
         n8750, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8780, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8790, n8791, n8792, n8794, n8795, n8797, n8799,
         n8800, n8801, n8802, n8804, n8805, n8806, n8808, n8809, n8810, n8811,
         n8812, n8813, n8816, n8817, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8831, n8832, n8834, n8835, n8836,
         n8838, n8840, n8841, n8843, n8844, n8845, n8846, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8875, n8876,
         n8882, n8883, n8885, n8886, n8892, n8893, n8894, n8895, n8896, n8897,
         n8899, n8901, n8902, n8903, n8905, n8906, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8937, n8939, n8940, n8941, n8942, n8943, n8944,
         n8946, n8948, n8949, n8950, n8951, n8953, n8954, n8955, n8957, n8958,
         n8959, n8960, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8970,
         n8972, n8973, n8974, n8975, n8976, n8979, n8980, n8983, n8984, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n9000, n9002, n9003, n9004, n9005, n9006, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9020, n9021, n9022, n9025,
         n9026, n9027, n9028, n9030, n9031, n9032, n9033, n9037, n9038, n9040,
         n9041, n9042, n9044, n9045, n9046, n9050, n9052, n9055, n9057, n9058,
         n9059, n9062, n9064, n9065, n9066, n9068, n9071, n9073, n9075, n9076,
         n9078, n9080, n9083, n9085, n9087, n9088, n9090, n9092, n9093, n9095,
         n9097, n9098, n9099, n9101, n9102, n9103, n9105, n9106, n9107, n9108,
         n9110, n9111, n9113, n9114, n9115, n9116, n9118, n9119, n9120, n9121,
         n9123, n9125, n9126, n9127, n9129, n9131, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9141, n9145, n9146, n9147, n9148, n9149, n9151,
         n9152, n9153, n9154, n9155, n9156, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9166, n9167, n9168, n9170, n9171, n9172, n9173, n9174,
         n9176, n9177, n9178, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9189, n9191, n9192, n9193, n9195, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9211, n9212,
         n9213, n9214, n9215, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9227, n9228, n9230, n9231, n9232, n9233, n9234, n9235,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9247, n9248,
         n9249, n9251, n9252, n9255, n9256, n9257, n9258, n9259, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9277, n9278, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9292, n9293, n9294, n9296, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9334,
         n9335, n9338, n9339, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9349, n9350, n9351, n9352, n9353, n9356, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9373, n9374, n9375, n9377,
         n9378, n9379, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9390, n9391, n9392, n9393, n9395, n9396, n9397, n9398, n9399, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9411, n9412, n9413,
         n9414, n9418, n9419, n9420, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9430, n9432, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9456, n9459, n9460, n9462, n9464, n9467, n9468,
         n9469, n9472, n9473, n9474, n9475, n9476, n9478, n9479, n9480, n9481,
         n9483, n9484, n9485, n9486, n9487, n9488, n9490, n9493, n9495, n9496,
         n9500, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9521, n9522,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9535, n9536,
         n9538, n9539, n9540, n9542, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9555, n9558, n9560, n9561, n9563, n9564,
         n9567, n9568, n9569, n9571, n9573, n9574, n9575, n9577, n9578, n9579,
         n9580, n9581, n9582, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9597, n9599, n9601, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9615, n9616, n9617, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9629, n9630,
         n9631, n9634, n9635, n9636, n9637, n9640, n9641, n9644, n9645, n9646,
         n9647, n9648, n9650, n9651, n9652, n9653, n9654, n9655, n9658, n9659,
         n9660, n9661, n9663, n9664, n9665, n9666, n9667, n9668, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9681, n9683,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9701, n9703, n9704, n9705, n9706, n9708,
         n9709, n9710, n9711, n9714, n9717, n9718, n9719, n9721, n9724, n9725,
         n9728, n9729, n9731, n9732, n9733, n9734, n9736, n9737, n9738, n9739,
         n9740, n9741, n9744, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9757, n9758, n9759, n9760, n9761, n9762, n9764, n9766, n9768,
         n9769, n9770, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9780,
         n9781, n9782, n9783, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9796, n9797, n9798, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9828, n9831, n9832, n9833, n9835, n9836, n9837, n9838,
         n9839, n9840, n9842, n9843, n9844, n9846, n9847, n9848, n9852, n9854,
         n9855, n9856, n9857, n9858, n9859, n9861, n9862, n9863, n9865, n9866,
         n9867, n9868, n9870, n9871, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9884, n9885, n9886, n9887, n9889, n9890, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9936, n9937, n9939, n9941, n9943, n9945, n9946, n9949,
         n9950, n9951, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9973,
         n9975, n9976, n9977, n9978, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9988, n9990, n9991, n9992, n9993, n9994, n9995, n9998, n9999,
         n10000, n10001, n10003, n10004, n10005, n10006, n10007, n10009,
         n10010, n10011, n10012, n10013, n10015, n10017, n10018, n10019,
         n10020, n10024, n10026, n10028, n10030, n10031, n10033, n10035,
         n10038, n10039, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10051, n10052, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10062, n10063, n10064, n10066, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10079, n10080, n10081, n10082, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10092, n10093, n10095, n10096, n10097,
         n10098, n10099, n10100, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10116,
         n10117, n10118, n10119, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10140, n10142, n10143, n10145,
         n10146, n10148, n10149, n10150, n10152, n10154, n10155, n10157,
         n10159, n10160, n10163, n10164, n10165, n10166, n10167, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10186,
         n10187, n10188, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10205, n10206,
         n10207, n10208, n10209, n10210, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10224, n10226, n10227,
         n10228, n10229, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10241, n10243, n10244, n10247, n10248, n10249, n10251,
         n10252, n10254, n10255, n10257, n10258, n10259, n10260, n10261,
         n10262, n10264, n10265, n10266, n10268, n10270, n10271, n10272,
         n10273, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10310,
         n10312, n10313, n10314, n10315, n10316, n10317, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10335, n10337, n10339, n10340, n10342,
         n10343, n10344, n10345, n10346, n10347, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10357, n10358, n10359, n10360,
         n10361, n10364, n10365, n10366, n10367, n10369, n10370, n10371,
         n10372, n10373, n10374, n10376, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10401, n10402, n10404, n10405, n10409, n10410, n10411,
         n10412, n10413, n10414, n10416, n10419, n10420, n10421, n10422,
         n10423, n10424, n10426, n10427, n10428, n10429, n10430, n10431,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10446, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10456, n10459, n10460, n10461,
         n10462, n10463, n10465, n10466, n10467, n10468, n10469, n10470,
         n10472, n10473, n10474, n10475, n10478, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10488, n10489, n10490, n10491,
         n10492, n10493, n10495, n10496, n10497, n10498, n10500, n10501,
         n10504, n10505, n10507, n10508, n10510, n10511, n10513, n10514,
         n10515, n10516, n10519, n10522, n10523, n10524, n10525, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10535, n10536,
         n10537, n10539, n10542, n10546, n10547, n10548, n10549, n10550,
         n10552, n10553, n10555, n10556, n10557, n10558, n10560, n10561,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10576, n10578, n10579, n10581, n10582,
         n10583, n10584, n10585, n10587, n10588, n10589, n10598, n10599,
         n10600, n10603, n10604, n10605, n10606, n10608, n10609, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10619, n10620,
         n10621, n10622, n10623, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10637, n10638, n10639, n10640, n10641,
         n10643, n10644, n10645, n10646, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10669, n10670,
         n10671, n10673, n10674, n10675, n10679, n10680, n10681, n10683,
         n10685, n10686, n10687, n10689, n10693, n10694, n10695, n10696,
         n10697, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10707, n10708, n10710, n10713, n10714, n10715, n10716, n10717,
         n10718, n10720, n10721, n10722, n10723, n10724, n10725, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10735, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10747, n10748, n10749, n10750, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10762, n10763, n10764,
         n10765, n10766, n10768, n10769, n10770, n10772, n10773, n10775,
         n10776, n10777, n10778, n10780, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10796,
         n10797, n10798, n10799, n10800, n10804, n10805, n10806, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10821, n10822, n10823, n10824, n10825, n10827, n10828, n10829,
         n10831, n10832, n10833, n10834, n10835, n10837, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10877, n10878,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10895, n10896, n10897, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10907, n10908, n10909, n10910, n10914,
         n10915, n10916, n10917, n10921, n10922, n10923, n10924, n10925,
         n10926, n10928, n10931, n10932, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10951, n10953, n10954, n10955,
         n10959, n10960, n10961, n10963, n10964, n10965, n10966, n10967,
         n10968, n10970, n10971, n10972, n10973, n10974, n10975, n10977,
         n10978, n10979, n10980, n10985, n10986, n10987, n10989, n10990,
         n10991, n10992, n10993, n10999, n11000, n11003, n11004, n11005,
         n11006, n11008, n11010, n11011, n11012, n11013, n11017, n11018,
         n11019, n11020, n11022, n11023, n11027, n11028, n11031, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11041, n11042,
         n11045, n11046, n11048, n11049, n11050, n11051, n11052, n11053,
         n11055, n11057, n11058, n11059, n11061, n11062, n11063, n11064,
         n11066, n11067, n11068, n11069, n11070, n11072, n11074, n11075,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11089, n11090, n11091, n11092, n11093, n11095,
         n11096, n11097, n11098, n11100, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11126,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11155, n11156, n11157, n11158, n11159, n11161, n11162, n11164,
         n11166, n11167, n11169, n11170, n11171, n11172, n11173, n11175,
         n11177, n11178, n11179, n11180, n11181, n11182, n11185, n11186,
         n11187, n11192, n11193, n11194, n11195, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11208, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11225, n11227, n11228,
         n11229, n11231, n11232, n11235, n11236, n11238, n11240, n11241,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11253, n11254, n11255, n11257, n11258, n11259, n11261,
         n11262, n11263, n11264, n11265, n11266, n11268, n11269, n11270,
         n11271, n11272, n11276, n11278, n11280, n11281, n11282, n11285,
         n11287, n11289, n11290, n11291, n11292, n11294, n11295, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11306,
         n11308, n11309, n11310, n11311, n11312, n11315, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11330, n11331, n11332, n11333, n11334, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11346, n11347, n11348,
         n11349, n11350, n11351, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11364, n11365, n11366,
         n11368, n11370, n11372, n11374, n11376, n11378, n11379, n11380,
         n11381, n11382, n11383, n11385, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11396, n11397, n11398, n11399,
         n11401, n11402, n11405, n11406, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11416, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11426, n11427, n11428, n11429, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11450, n11451, n11452, n11453, n11454, n11456, n11457, n11458,
         n11459, n11460, n11461, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11474, n11475, n11476, n11477, n11480,
         n11481, n11483, n11484, n11485, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11497, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11507, n11508, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11542, n11543, n11544, n11545,
         n11548, n11551, n11552, n11555, n11556, n11557, n11558, n11559,
         n11560, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11574, n11575, n11576, n11577, n11578,
         n11580, n11581, n11582, n11584, n11585, n11586, n11587, n11589,
         n11590, n11591, n11593, n11595, n11596, n11597, n11599, n11600,
         n11601, n11603, n11604, n11605, n11608, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11626, n11627, n11628, n11629,
         n11630, n11631, n11633, n11634, n11635, n11636, n11637, n11640,
         n11641, n11643, n11644, n11645, n11646, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11663, n11665, n11666, n11667, n11668, n11669, n11670, n11673,
         n11675, n11676, n11677, n11678, n11680, n11681, n11682, n11683,
         n11684, n11686, n11687, n11688, n11689, n11690, n11691, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11732, n11733, n11734, n11735, n11736, n11737,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11748,
         n11749, n11750, n11751, n11752, n11754, n11755, n11756, n11757,
         n11759, n11760, n11761, n11762, n11765, n11766, n11767, n11768,
         n11769, n11770, n11773, n11774, n11775, n11776, n11777, n11778,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11788,
         n11789, n11792, n11795, n11796, n11797, n11798, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11812, n11814, n11815, n11816, n11817, n11819, n11820, n11821,
         n11822, n11823, n11824, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11847,
         n11848, n11850, n11852, n11853, n11854, n11855, n11856, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11880, n11883, n11884, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11895, n11897, n11898, n11899, n11900,
         n11902, n11903, n11904, n11905, n11907, n11909, n11910, n11911,
         n11912, n11913, n11915, n11916, n11917, n11918, n11919, n11920,
         n11922, n11923, n11924, n11925, n11926, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11966,
         n11967, n11968, n11969, n11970, n11971, n11973, n11974, n11975,
         n11976, n11977, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11990, n11991, n11992, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12002, n12004,
         n12005, n12006, n12008, n12010, n12011, n12013, n12014, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12048, n12049, n12051, n12052, n12053,
         n12054, n12055, n12057, n12058, n12059, n12060, n12061, n12062,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12074, n12075, n12076, n12077, n12078, n12080, n12082, n12083,
         n12084, n12085, n12086, n12088, n12089, n12090, n12091, n12093,
         n12094, n12095, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12107, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12127, n12128, n12130, n12131, n12132, n12133,
         n12135, n12136, n12137, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12147, n12148, n12149, n12150, n12151, n12153,
         n12154, n12156, n12157, n12159, n12160, n12161, n12163, n12164,
         n12165, n12166, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12208, n12209, n12211, n12212,
         n12213, n12214, n12215, n12217, n12218, n12220, n12221, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12243, n12244, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12256, n12257, n12258, n12259, n12260, n12262,
         n12263, n12264, n12265, n12266, n12268, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12290, n12291, n12293, n12295, n12296, n12297, n12300, n12302,
         n12304, n12308, n12309, n12310, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12340, n12341,
         n12342, n12343, n12344, n12345, n12347, n12348, n12351, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12379, n12380, n12381,
         n12382, n12383, n12384, n12386, n12387, n12390, n12391, n12392,
         n12394, n12395, n12396, n12397, n12398, n12399, n12402, n12403,
         n12407, n12408, n12409, n12410, n12411, n12413, n12414, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12429, n12430, n12431, n12432, n12433, n12434, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12448, n12449,
         n12450, n12452, n12453, n12454, n12456, n12457, n12458, n12459,
         n12461, n12462, n12465, n12467, n12468, n12469, n12471, n12472,
         n12473, n12474, n12475, n12476, n12478, n12479, n12482, n12485,
         n12486, n12487, n12488, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12500, n12502, n12504, n12505,
         n12506, n12507, n12508, n12509, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12519, n12520, n12521, n12522, n12525,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12538, n12539, n12540, n12541, n12542, n12545,
         n12546, n12547, n12548, n12549, n12551, n12552, n12553, n12556,
         n12557, n12559, n12561, n12562, n12563, n12564, n12565, n12567,
         n12568, n12570, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12582, n12583, n12584, n12585, n12586,
         n12587, n12590, n12592, n12593, n12594, n12595, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12609, n12610, n12611, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12624, n12625, n12626,
         n12627, n12628, n12629, n12632, n12634, n12636, n12637, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12657, n12658, n12659,
         n12662, n12663, n12665, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12704, n12705, n12707, n12708, n12711, n12712,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12724, n12725, n12726, n12727, n12728, n12729, n12731,
         n12732, n12733, n12735, n12736, n12738, n12742, n12743, n12744,
         n12746, n12747, n12748, n12749, n12750, n12751, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12762, n12763,
         n12764, n12765, n12768, n12770, n12771, n12774, n12775, n12777,
         n12779, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12803, n12804, n12805,
         n12807, n12808, n12809, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12821, n12823, n12824, n12826, n12827, n12828,
         n12830, n12831, n12832, n12836, n12837, n12840, n12841, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12855, n12856, n12858, n12861, n12862, n12863,
         n12864, n12865, n12866, n12868, n12869, n12871, n12872, n12873,
         n12875, n12876, n12877, n12878, n12879, n12880, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12891, n12892, n12894,
         n12895, n12896, n12898, n12899, n12900, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12915, n12916, n12917, n12918, n12919, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12939,
         n12942, n12943, n12944, n12945, n12947, n12948, n12950, n12951,
         n12952, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12962, n12966, n12968, n12969, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12980, n12981, n12982, n12983, n12985,
         n12986, n12987, n12989, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13006, n13008, n13009, n13011, n13012, n13013, n13014,
         n13015, n13016, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13040, n13041, n13042, n13043, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13055, n13056, n13058, n13059, n13060, n13061, n13063, n13065,
         n13066, n13067, n13068, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13082, n13083,
         n13084, n13085, n13086, n13087, n13089, n13090, n13091, n13092,
         n13093, n13095, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13120, n13121, n13122, n13123, n13124,
         n13125, n13127, n13129, n13130, n13131, n13132, n13133, n13136,
         n13137, n13138, n13139, n13140, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13154,
         n13157, n13159, n13160, n13161, n13162, n13163, n13167, n13168,
         n13169, n13170, n13172, n13173, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13204, n13205, n13208, n13209,
         n13210, n13212, n13213, n13214, n13216, n13217, n13219, n13222,
         n13223, n13224, n13226, n13227, n13230, n13231, n13232, n13234,
         n13235, n13236, n13237, n13238, n13239, n13242, n13243, n13245,
         n13246, n13247, n13248, n13249, n13251, n13252, n13253, n13254,
         n13255, n13258, n13260, n13261, n13262, n13263, n13265, n13266,
         n13267, n13268, n13272, n13273, n13274, n13275, n13276, n13279,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13308, n13309, n13310, n13312, n13313, n13314, n13315,
         n13316, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13334, n13336, n13338, n13339, n13340, n13341, n13342, n13343,
         n13345, n13346, n13347, n13348, n13349, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13363, n13364,
         n13365, n13366, n13367, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13377, n13378, n13379, n13380, n13381, n13382,
         n13384, n13386, n13388, n13389, n13390, n13391, n13393, n13394,
         n13395, n13396, n13397, n13401, n13402, n13403, n13404, n13405,
         n13407, n13408, n13409, n13411, n13412, n13413, n13414, n13415,
         n13417, n13419, n13421, n13422, n13423, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13444, n13445,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13464,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13485, n13488, n13489, n13490, n13491, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13506, n13507, n13508, n13509, n13510, n13511, n13513,
         n13514, n13517, n13519, n13520, n13521, n13524, n13525, n13526,
         n13527, n13528, n13529, n13530, n13531, n13532, n13534, n13535,
         n13537, n13538, n13539, n13540, n13541, n13544, n13545, n13546,
         n13547, n13548, n13549, n13551, n13552, n13553, n13554, n13555,
         n13556, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13578, n13579, n13580, n13581,
         n13582, n13583, n13585, n13586, n13587, n13589, n13590, n13591,
         n13592, n13593, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13605, n13606, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13621, n13622, n13623, n13624, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13635, n13636, n13637, n13638,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13673,
         n13677, n13678, n13679, n13680, n13681, n13682, n13684, n13685,
         n13686, n13689, n13690, n13692, n13693, n13694, n13695, n13696,
         n13698, n13700, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13712, n13716, n13719, n13720, n13721,
         n13723, n13724, n13725, n13727, n13730, n13732, n13733, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13745, n13746, n13747, n13748, n13751, n13752, n13759, n13760,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13770,
         n13771, n13772, n13773, n13774, n13777, n13778, n13780, n13782,
         n13783, n13784, n13785, n13786, n13787, n13788, n13791, n13792,
         n13793, n13794, n13796, n13800, n13802, n13803, n13804, n13806,
         n13807, n13809, n13810, n13811, n13812, n13814, n13815, n13816,
         n13817, n13819, n13822, n13824, n13825, n13826, n13828, n13829,
         n13830, n13831, n13833, n13834, n13835, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13867, n13869, n13872, n13873, n13874, n13876, n13877, n13878,
         n13879, n13880, n13881, n13883, n13884, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13898, n13899, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13920, n13921, n13922, n13924, n13925,
         n13927, n13928, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13943, n13944,
         n13945, n13946, n13947, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13960, n13962, n13963, n13965,
         n13966, n13968, n13969, n13970, n13971, n13972, n13973, n13974,
         n13975, n13977, n13978, n13979, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13989, n13993, n13994, n13995, n13996,
         n13998, n14000, n14001, n14002, n14004, n14005, n14008, n14009,
         n14010, n14011, n14012, n14014, n14016, n14017, n14019, n14020,
         n14021, n14022, n14023, n14024, n14027, n14029, n14030, n14031,
         n14032, n14033, n14034, n14036, n14037, n14038, n14039, n14041,
         n14042, n14043, n14044, n14045, n14047, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14058, n14060, n14062,
         n14065, n14066, n14067, n14069, n14070, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14086, n14087, n14088, n14091, n14092, n14093, n14094, n14095,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14106,
         n14107, n14108, n14110, n14111, n14112, n14113, n14114, n14117,
         n14118, n14119, n14120, n14122, n14123, n14124, n14125, n14126,
         n14129, n14130, n14131, n14132, n14133, n14134, n14136, n14137,
         n14138, n14139, n14142, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14153, n14154, n14155, n14156, n14157, n14159,
         n14160, n14161, n14162, n14163, n14164, n14166, n14168, n14170,
         n14171, n14172, n14173, n14174, n14176, n14177, n14178, n14179,
         n14181, n14183, n14184, n14187, n14188, n14189, n14190, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14201,
         n14202, n14203, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14219, n14220,
         n14221, n14222, n14223, n14227, n14228, n14230, n14231, n14232,
         n14233, n14234, n14236, n14237, n14238, n14239, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14255, n14257, n14258, n14259, n14261, n14262,
         n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
         n14271, n14272, n14273, n14274, n14276, n14277, n14279, n14280,
         n14281, n14282, n14283, n14284, n14288, n14289, n14290, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14305, n14306, n14307, n14308, n14309, n14311, n14312,
         n14314, n14315, n14316, n14318, n14320, n14321, n14322, n14325,
         n14326, n14327, n14328, n14329, n14331, n14332, n14334, n14335,
         n14336, n14337, n14339, n14340, n14342, n14344, n14346, n14348,
         n14349, n14350, n14352, n14354, n14355, n14359, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14373, n14375, n14376, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14391, n14392, n14393, n14394,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14404,
         n14407, n14409, n14410, n14411, n14412, n14415, n14416, n14417,
         n14418, n14419, n14420, n14422, n14423, n14424, n14425, n14426,
         n14428, n14429, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14442, n14443, n14444, n14445, n14447,
         n14449, n14450, n14451, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14463, n14464, n14465, n14466,
         n14470, n14471, n14472, n14473, n14478, n14479, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14509, n14510, n14511, n14513, n14514, n14516, n14517,
         n14518, n14519, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14529, n14530, n14531, n14532, n14533, n14534, n14536,
         n14537, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14550, n14551, n14552, n14555, n14556,
         n14557, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14597, n14598, n14600, n14601,
         n14602, n14603, n14605, n14606, n14607, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14671, n14673, n14674,
         n14676, n14677, n14678, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14701, n14702, n14703,
         n14704, n14705, n14706, n14708, n14709, n14710, n14711, n14712,
         n14713, n14716, n14717, n14719, n14720, n14721, n14722, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14772, n14773, n14774, n14775, n14776,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14791, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14801, n14802, n14803, n14805,
         n14806, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14817, n14818, n14819, n14820, n14821, n14822, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14851, n14853, n14854, n14855,
         n14856, n14858, n14859, n14860, n14861, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14878, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14895, n14896, n14897, n14898, n14899, n14901, n14902,
         n14903, n14905, n14906, n14907, n14908, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14920, n14922, n14924,
         n14925, n14926, n14927, n14930, n14931, n14932, n14933, n14934,
         n14935, n14937, n14938, n14939, n14940, n14942, n14943, n14944,
         n14945, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14957, n14959, n14960, n14964, n14965, n14966, n14967,
         n14968, n14969, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14983, n14985, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15002, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15031, n15032, n15033,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15077, n15078, n15079,
         n15083, n15084, n15085, n15086, n15089, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15101, n15103,
         n15106, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15119, n15120, n15121, n15123, n15124,
         n15126, n15127, n15129, n15130, n15132, n15133, n15134, n15135,
         n15136, n15137, n15139, n15140, n15141, n15142, n15143, n15144,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15160, n15161, n15162,
         n15165, n15166, n15167, n15168, n15169, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15179, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15198, n15204, n15205, n15206, n15207,
         n15208, n15211, n15212, n15213, n15215, n15216, n15217, n15219,
         n15220, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15234, n15235, n15236, n15237, n15238,
         n15239, n15240, n15241, n15242, n15243, n15245, n15246, n15247,
         n15249, n15250, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15264, n15265, n15266, n15267, n15268,
         n15270, n15271, n15272, n15274, n15275, n15276, n15277, n15278,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15321, n15322, n15323, n15324,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15334,
         n15335, n15337, n15338, n15339, n15340, n15341, n15343, n15344,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15362,
         n15364, n15365, n15366, n15367, n15368, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15381,
         n15382, n15383, n15384, n15385, n15386, n15389, n15390, n15391,
         n15393, n15394, n15395, n15396, n15397, n15399, n15400, n15401,
         n15402, n15404, n15405, n15406, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15441, n15442, n15443, n15444, n15446, n15448,
         n15449, n15450, n15451, n15452, n15455, n15456, n15457, n15458,
         n15459, n15460, n15462, n15464, n15465, n15466, n15467, n15468,
         n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
         n15478, n15479, n15480, n15481, n15483, n15484, n15485, n15486,
         n15487, n15489, n15490, n15494, n15495, n15496, n15497, n15498,
         n15500, n15501, n15502, n15505, n15506, n15507, n15508, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15534, n15536, n15537, n15538, n15539, n15540, n15543,
         n15544, n15546, n15548, n15550, n15551, n15553, n15555, n15556,
         n15557, n15559, n15560, n15561, n15562, n15564, n15565, n15566,
         n15569, n15570, n15571, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15583, n15584, n15585, n15588,
         n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15597,
         n15598, n15599, n15600, n15601, n15602, n15606, n15607, n15608,
         n15609, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15621, n15622, n15623, n15624, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15635, n15636, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15646, n15650, n15652,
         n15653, n15655, n15658, n15659, n15660, n15661, n15662, n15663,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15679, n15680, n15681,
         n15682, n15683, n15685, n15686, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15701, n15702,
         n15704, n15705, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15740, n15742, n15743, n15744, n15745, n15746, n15747, n15748,
         n15749, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
         n15759, n15761, n15763, n15765, n15768, n15769, n15770, n15771,
         n15772, n15774, n15775, n15776, n15777, n15778, n15779, n15780,
         n15781, n15783, n15785, n15786, n15787, n15788, n15789, n15790,
         n15791, n15792, n15793, n15795, n15796, n15797, n15798, n15799,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15827,
         n15828, n15829, n15830, n15831, n15832, n15833, n15835, n15836,
         n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844,
         n15845, n15846, n15847, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15857, n15858, n15859, n15860, n15861, n15862,
         n15863, n15864, n15865, n15867, n15869, n15870, n15872, n15873,
         n15874, n15875, n15876, n15877, n15880, n15882, n15883, n15885,
         n15886, n15887, n15888, n15889, n15890, n15891, n15893, n15894,
         n15896, n15897, n15898, n15899, n15900, n15902, n15904, n15905,
         n15906, n15907, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15917, n15919, n15920, n15923, n15925, n15927, n15928,
         n15929, n15930, n15931, n15932, n15934, n15935, n15936, n15939,
         n15941, n15942, n15943, n15944, n15946, n15947, n15948, n15949,
         n15950, n15951, n15953, n15954, n15955, n15956, n15957, n15959,
         n15960, n15961, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15971, n15973, n15974, n15976, n15977, n15978, n15979,
         n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15990,
         n15991, n15992, n15993, n15994, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16004, n16005, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16016, n16017, n16018,
         n16021, n16022, n16023, n16024, n16025, n16027, n16028, n16029,
         n16030, n16033, n16034, n16035, n16036, n16038, n16039, n16041,
         n16042, n16045, n16046, n16047, n16048, n16050, n16051, n16052,
         n16053, n16054, n16058, n16059, n16060, n16062, n16065, n16066,
         n16068, n16070, n16072, n16073, n16076, n16077, n16078, n16080,
         n16081, n16083, n16084, n16085, n16086, n16088, n16090, n16091,
         n16092, n16093, n16094, n16096, n16097, n16098, n16099, n16100,
         n16104, n16105, n16106, n16108, n16109, n16110, n16111, n16112,
         n16113, n16115, n16117, n16118, n16120, n16121, n16122, n16123,
         n16124, n16125, n16127, n16128, n16129, n16132, n16133, n16134,
         n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16144,
         n16146, n16147, n16148, n16149, n16150, n16152, n16154, n16155,
         n16156, n16157, n16158, n16159, n16160, n16162, n16163, n16164,
         n16165, n16166, n16167, n16169, n16170, n16173, n16174, n16175,
         n16176, n16178, n16180, n16181, n16182, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16200, n16202, n16203, n16204,
         n16205, n16207, n16209, n16210, n16211, n16212, n16215, n16216,
         n16217, n16218, n16220, n16221, n16222, n16224, n16225, n16226,
         n16228, n16229, n16231, n16232, n16235, n16236, n16237, n16238,
         n16239, n16240, n16241, n16242, n16243, n16246, n16247, n16248,
         n16249, n16251, n16253, n16254, n16257, n16258, n16259, n16260,
         n16261, n16262, n16263, n16265, n16266, n16267, n16269, n16271,
         n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279,
         n16280, n16281, n16282, n16283, n16284, n16286, n16287, n16288,
         n16290, n16291, n16292, n16293, n16295, n16297, n16298, n16300,
         n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308,
         n16309, n16310, n16311, n16313, n16315, n16317, n16318, n16319,
         n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
         n16328, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16343, n16344, n16345, n16346, n16347, n16348,
         n16349, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
         n16358, n16359, n16361, n16363, n16364, n16366, n16367, n16370,
         n16371, n16372, n16373, n16374, n16375, n16377, n16378, n16380,
         n16381, n16382, n16383, n16384, n16386, n16387, n16388, n16389,
         n16390, n16392, n16393, n16394, n16395, n16397, n16398, n16400,
         n16401, n16402, n16403, n16406, n16408, n16409, n16410, n16411,
         n16412, n16413, n16414, n16416, n16417, n16418, n16420, n16421,
         n16422, n16423, n16424, n16425, n16426, n16429, n16430, n16431,
         n16432, n16434, n16435, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16447, n16448, n16450, n16451,
         n16452, n16453, n16454, n16457, n16458, n16459, n16461, n16462,
         n16463, n16464, n16466, n16467, n16468, n16469, n16472, n16473,
         n16474, n16477, n16479, n16481, n16482, n16483, n16484, n16485,
         n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493,
         n16494, n16496, n16497, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16509, n16510, n16512, n16513, n16514, n16515,
         n16516, n16518, n16519, n16520, n16522, n16523, n16525, n16526,
         n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534,
         n16535, n16536, n16538, n16539, n16540, n16541, n16543, n16544,
         n16545, n16546, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16566, n16567, n16568, n16569, n16570, n16572,
         n16573, n16574, n16575, n16577, n16578, n16579, n16581, n16582,
         n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590,
         n16591, n16592, n16595, n16596, n16597, n16598, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16611, n16612, n16613, n16614, n16615, n16617, n16618, n16619,
         n16620, n16621, n16622, n16623, n16624, n16625, n16627, n16628,
         n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636,
         n16637, n16639, n16640, n16641, n16642, n16643, n16646, n16647,
         n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655,
         n16657, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16668, n16669, n16670, n16671, n16672, n16673, n16674,
         n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,
         n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690,
         n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698,
         n16699, n16700, n16701, n16703, n16704, n16705, n16708, n16710,
         n16711, n16712, n16713, n16716, n16717, n16718, n16719, n16722,
         n16723, n16724, n16725, n16727, n16728, n16729, n16730, n16732,
         n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740,
         n16741, n16743, n16745, n16747, n16748, n16749, n16750, n16751,
         n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759,
         n16762, n16763, n16766, n16767, n16768, n16769, n16770, n16773,
         n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781,
         n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789,
         n16790, n16792, n16793, n16795, n16796, n16797, n16798, n16799,
         n16800, n16801, n16803, n16804, n16805, n16806, n16807, n16809,
         n16810, n16811, n16812, n16815, n16816, n16817, n16818, n16819,
         n16820, n16823, n16824, n16826, n16827, n16828, n16829, n16831,
         n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16841,
         n16842, n16844, n16845, n16847, n16848, n16849, n16850, n16851,
         n16852, n16853, n16854, n16855, n16857, n16858, n16859, n16861,
         n16862, n16863, n16864, n16866, n16867, n16868, n16869, n16870,
         n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16879,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16891, n16893, n16896, n16897, n16898, n16899, n16901,
         n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911,
         n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919,
         n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927,
         n16928, n16930, n16933, n16934, n16937, n16938, n16939, n16940,
         n16943, n16945, n16946, n16947, n16948, n16949, n16950, n16951,
         n16952, n16953, n16954, n16955, n16957, n16958, n16959, n16960,
         n16961, n16962, n16963, n16964, n16966, n16969, n16971, n16972,
         n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980,
         n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16989,
         n16992, n16993, n16995, n16996, n16997, n16998, n17001, n17002,
         n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010,
         n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018,
         n17019, n17021, n17022, n17023, n17026, n17028, n17029, n17030,
         n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042,
         n17043, n17044, n17046, n17047, n17048, n17049, n17050, n17051,
         n17052, n17053, n17054, n17055, n17056, n17058, n17060, n17061,
         n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069,
         n17072, n17073, n17074, n17076, n17077, n17078, n17079, n17083,
         n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091,
         n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
         n17100, n17101, n17102, n17104, n17105, n17106, n17108, n17109,
         n17110, n17112, n17113, n17114, n17115, n17117, n17118, n17119,
         n17120, n17122, n17123, n17124, n17125, n17126, n17127, n17128,
         n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136,
         n17139, n17140, n17141, n17143, n17144, n17145, n17146, n17147,
         n17148, n17149, n17150, n17151, n17153, n17155, n17156, n17157,
         n17159, n17161, n17162, n17163, n17164, n17165, n17166, n17167,
         n17168, n17169, n17171, n17172, n17174, n17175, n17177, n17178,
         n17180, n17181, n17183, n17184, n17185, n17186, n17187, n17188,
         n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196,
         n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206,
         n17207, n17211, n17212, n17213, n17214, n17215, n17217, n17218,
         n17219, n17220, n17222, n17223, n17224, n17225, n17226, n17227,
         n17228, n17231, n17232, n17233, n17234, n17235, n17236, n17237,
         n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245,
         n17247, n17248, n17249, n17251, n17253, n17254, n17255, n17257,
         n17258, n17259, n17260, n17261, n17263, n17266, n17268, n17269,
         n17270, n17271, n17272, n17273, n17274, n17277, n17278, n17280,
         n17281, n17282, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17293, n17295, n17296, n17297, n17298, n17299,
         n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
         n17308, n17309, n17310, n17311, n17313, n17316, n17317, n17318,
         n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17327,
         n17328, n17329, n17330, n17331, n17333, n17334, n17335, n17336,
         n17338, n17339, n17341, n17342, n17346, n17347, n17348, n17350,
         n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17359,
         n17360, n17361, n17362, n17363, n17364, n17365, n17367, n17368,
         n17369, n17370, n17371, n17373, n17374, n17375, n17377, n17378,
         n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386,
         n17387, n17389, n17392, n17393, n17394, n17395, n17396, n17398,
         n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406,
         n17407, n17408, n17409, n17411, n17414, n17415, n17416, n17418,
         n17419, n17420, n17422, n17423, n17424, n17425, n17426, n17428,
         n17429, n17430, n17431, n17432, n17434, n17435, n17436, n17437,
         n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445,
         n17446, n17448, n17450, n17452, n17453, n17455, n17456, n17457,
         n17458, n17460, n17462, n17463, n17464, n17465, n17466, n17467,
         n17472, n17473, n17475, n17476, n17477, n17478, n17479, n17480,
         n17481, n17482, n17483, n17485, n17486, n17487, n17488, n17489,
         n17490, n17492, n17493, n17494, n17495, n17496, n17497, n17498,
         n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
         n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
         n17515, n17516, n17517, n17518, n17519, n17520, n17522, n17523,
         n17524, n17525, n17526, n17527, n17528, n17529, n17531, n17532,
         n17535, n17537, n17538, n17540, n17541, n17542, n17543, n17544,
         n17546, n17547, n17548, n17549, n17551, n17552, n17553, n17554,
         n17555, n17556, n17557, n17558, n17559, n17561, n17562, n17563,
         n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571,
         n17572, n17573, n17574, n17575, n17576, n17578, n17579, n17580,
         n17581, n17582, n17584, n17585, n17586, n17587, n17588, n17589,
         n17590, n17591, n17592, n17593, n17594, n17595, n17597, n17598,
         n17599, n17600, n17601, n17602, n17604, n17605, n17606, n17608,
         n17609, n17612, n17613, n17616, n17617, n17618, n17621, n17622,
         n17623, n17624, n17625, n17626, n17627, n17628, n17630, n17631,
         n17633, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17647, n17649, n17650, n17651, n17652,
         n17653, n17655, n17658, n17659, n17661, n17662, n17663, n17664,
         n17665, n17666, n17668, n17669, n17670, n17672, n17673, n17675,
         n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683,
         n17684, n17685, n17687, n17688, n17689, n17691, n17692, n17693,
         n17694, n17696, n17697, n17698, n17699, n17701, n17703, n17704,
         n17705, n17707, n17708, n17709, n17711, n17712, n17713, n17714,
         n17715, n17716, n17717, n17718, n17720, n17721, n17722, n17723,
         n17725, n17726, n17728, n17729, n17730, n17731, n17732, n17734,
         n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742,
         n17743, n17744, n17745, n17746, n17747, n17748, n17750, n17752,
         n17753, n17754, n17755, n17756, n17758, n17759, n17760, n17762,
         n17764, n17765, n17766, n17767, n17768, n17770, n17771, n17773,
         n17774, n17775, n17777, n17778, n17779, n17781, n17782, n17784,
         n17785, n17786, n17787, n17790, n17791, n17792, n17793, n17797,
         n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805,
         n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813,
         n17814, n17815, n17816, n17817, n17819, n17820, n17821, n17822,
         n17824, n17826, n17828, n17829, n17830, n17832, n17833, n17834,
         n17835, n17837, n17838, n17839, n17840, n17841, n17843, n17844,
         n17845, n17849, n17850, n17853, n17855, n17857, n17858, n17859,
         n17860, n17861, n17863, n17865, n17866, n17867, n17869, n17871,
         n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879,
         n17880, n17881, n17882, n17883, n17884, n17886, n17887, n17888,
         n17889, n17890, n17891, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17903, n17904, n17905, n17906, n17907,
         n17910, n17912, n17913, n17914, n17915, n17916, n17917, n17918,
         n17919, n17922, n17923, n17924, n17925, n17926, n17927, n17928,
         n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,
         n17937, n17938, n17939, n17940, n17941, n17943, n17944, n17945,
         n17947, n17948, n17949, n17950, n17953, n17954, n17955, n17956,
         n17957, n17958, n17959, n17960, n17963, n17964, n17967, n17968,
         n17970, n17971, n17973, n17974, n17975, n17977, n17978, n17980,
         n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17991,
         n17992, n17993, n17995, n17996, n17997, n17998, n17999, n18001,
         n18002, n18003, n18005, n18006, n18007, n18010, n18011, n18012,
         n18013, n18015, n18017, n18018, n18019, n18020, n18021, n18022,
         n18024, n18025, n18026, n18028, n18029, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18041, n18042,
         n18043, n18044, n18047, n18048, n18049, n18050, n18051, n18054,
         n18055, n18056, n18058, n18059, n18062, n18064, n18065, n18068,
         n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078,
         n18079, n18080, n18082, n18083, n18084, n18085, n18088, n18089,
         n18090, n18091, n18094, n18095, n18096, n18098, n18099, n18100,
         n18101, n18102, n18103, n18105, n18106, n18107, n18108, n18109,
         n18110, n18112, n18113, n18114, n18117, n18118, n18119, n18120,
         n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,
         n18129, n18130, n18131, n18132, n18133, n18135, n18136, n18137,
         n18138, n18139, n18141, n18142, n18143, n18144, n18145, n18146,
         n18147, n18148, n18149, n18150, n18151, n18152, n18154, n18155,
         n18156, n18159, n18160, n18161, n18162, n18163, n18165, n18166,
         n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174,
         n18175, n18177, n18179, n18180, n18181, n18182, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18192, n18194, n18195,
         n18196, n18197, n18198, n18199, n18200, n18204, n18205, n18206,
         n18207, n18208, n18209, n18210, n18213, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18224, n18225, n18226, n18227,
         n18228, n18230, n18231, n18235, n18236, n18237, n18238, n18239,
         n18240, n18241, n18242, n18246, n18251, n18254, n18256, n18257,
         n18259, n18260, n18261, n18264, n18265, n18266, n18267, n18268,
         n18269, n18270, n18274, n18275, n18276, n18277, n18278, n18279,
         n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287,
         n18288, n18289, n18290, n18292, n18293, n18294, n18295, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18307,
         n18308, n18309, n18310, n18311, n18313, n18314, n18315, n18316,
         n18317, n18318, n18320, n18321, n18322, n18323, n18324, n18326,
         n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334,
         n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18344,
         n18345, n18346, n18347, n18348, n18349, n18350, n18352, n18354,
         n18356, n18357, n18359, n18360, n18361, n18362, n18363, n18364,
         n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372,
         n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18381,
         n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389,
         n18390, n18391, n18392, n18393, n18395, n18396, n18397, n18398,
         n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406,
         n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18415,
         n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423,
         n18424, n18425, n18426, n18427, n18428, n18429, n18431, n18432,
         n18433, n18434, n18435, n18437, n18438, n18439, n18440, n18441,
         n18443, n18444, n18445, n18446, n18447, n18449, n18450, n18452,
         n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460,
         n18462, n18463, n18464, n18467, n18468, n18469, n18470, n18471,
         n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479,
         n18480, n18481, n18482, n18483, n18485, n18486, n18487, n18488,
         n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496,
         n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504,
         n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512,
         n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520,
         n18521, n18522, n18524, n18525, n18526, n18527, n18528, n18530,
         n18531, n18532, n18534, n18535, n18536, n18537, n18538, n18539,
         n18540, n18541, n18543, n18546, n18548, n18549, n18550, n18551,
         n18553, n18554, n18555, n18556, n18557, n18559, n18560, n18561,
         n18563, n18565, n18566, n18567, n18569, n18571, n18572, n18573,
         n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581,
         n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18590,
         n18591, n18593, n18594, n18595, n18596, n18598, n18599, n18600,
         n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608,
         n18609, n18613, n18615, n18616, n18617, n18618, n18619, n18621,
         n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629,
         n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638,
         n18639, n18640, n18641, n18642, n18643, n18647, n18648, n18649,
         n18650, n18651, n18653, n18654, n18655, n18656, n18657, n18658,
         n18659, n18660, n18662, n18663, n18664, n18665, n18666, n18667,
         n18668, n18669, n18671, n18672, n18674, n18676, n18677, n18678,
         n18679, n18680, n18681, n18682, n18683, n18686, n18687, n18688,
         n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698,
         n18699, n18700, n18701, n18702, n18704, n18705, n18706, n18707,
         n18708, n18709, n18710, n18711, n18714, n18715, n18716, n18717,
         n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18726,
         n18727, n18729, n18730, n18731, n18732, n18733, n18734, n18735,
         n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743,
         n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751,
         n18752, n18753, n18754, n18755, n18756, n18757, n18759, n18760,
         n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768,
         n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776,
         n18777, n18778, n18779, n18780, n18781, n18782, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18835,
         n18836, n18838, n18839, n18840, n18841, n18842, n18843, n18844,
         n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18853,
         n18854, n18855, n18856, n18858, n18859, n18860, n18861, n18862,
         n18863, n18864, n18865, n18866, n18867, n18869, n18870, n18871,
         n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880,
         n18881, n18882, n18884, n18885, n18886, n18887, n18888, n18889,
         n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898,
         n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18907,
         n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
         n18916, n18917, n18919, n18920, n18921, n18922, n18923, n18924,
         n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932,
         n18935, n18937, n18938, n18939, n18940, n18941, n18942, n18943,
         n18944, n18945, n18946, n18947, n18948, n18949, n18952, n18953,
         n18955, n18956, n18957, n18958, n18959, n18960, n18962, n18963,
         n18964, n18965, n18966, n18967, n18969, n18970, n18971, n18973,
         n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18982,
         n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990,
         n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18999,
         n19000, n19002, n19003, n19004, n19006, n19007, n19008, n19009,
         n19010, n19011, n19013, n19014, n19016, n19017, n19020, n19021,
         n19022, n19023, n19024, n19026, n19027, n19028, n19029, n19030,
         n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038,
         n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046,
         n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19056,
         n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064,
         n19065, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19084,
         n19085, n19087, n19088, n19089, n19090, n19091, n19092, n19093,
         n19094, n19095, n19096, n19097, n19098, n19100, n19101, n19102,
         n19103, n19104, n19105, n19107, n19108, n19109, n19110, n19111,
         n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119,
         n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19128,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19139, n19140, n19141, n19142, n19143, n19144, n19146, n19147,
         n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155,
         n19156, n19158, n19160, n19161, n19162, n19163, n19164, n19165,
         n19167, n19168, n19170, n19171, n19172, n19173, n19174, n19175,
         n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183,
         n19185, n19186, n19188, n19189, n19190, n19193, n19195, n19196,
         n19197, n19198, n19199, n19200, n19202, n19203, n19204, n19205,
         n19206, n19209, n19210, n19211, n19212, n19214, n19215, n19216,
         n19217, n19218, n19219, n19220, n19222, n19224, n19225, n19226,
         n19227, n19228, n19229, n19230, n19232, n19233, n19234, n19235,
         n19236, n19238, n19239, n19240, n19241, n19242, n19243, n19244,
         n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252,
         n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260,
         n19261, n19262, n19263, n19265, n19267, n19268, n19269, n19270,
         n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278,
         n19280, n19281, n19282, n19283, n19284, n19285, n19287, n19288,
         n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296,
         n19297, n19298, n19300, n19301, n19302, n19303, n19305, n19307,
         n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
         n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323,
         n19324, n19325, n19326, n19328, n19329, n19330, n19331, n19332,
         n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340,
         n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348,
         n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356,
         n19357, n19359, n19360, n19361, n19362, n19363, n19364, n19365,
         n19366, n19367, n19368, n19370, n19371, n19372, n19373, n19374,
         n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382,
         n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391,
         n19394, n19395, n19397, n19398, n19399, n19400, n19401, n19402,
         n19403, n19405, n19406, n19407, n19408, n19409, n19411, n19412,
         n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420,
         n19421, n19422, n19423, n19424, n19426, n19427, n19428, n19429,
         n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19438,
         n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446,
         n19447, n19448, n19449, n19450, n19451, n19453, n19454, n19455,
         n19456, n19457, n19459, n19460, n19461, n19462, n19463, n19464,
         n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19473,
         n19474, n19475, n19476, n19479, n19480, n19481, n19482, n19483,
         n19484, n19485, n19486, n19487, n19490, n19491, n19492, n19493,
         n19494, n19495, n19496, n19497, n19498, n19500, n19501, n19502,
         n19503, n19504, n19505, n19507, n19508, n19509, n19510, n19511,
         n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519,
         n19520, n19522, n19523, n19524, n19525, n19526, n19527, n19528,
         n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536,
         n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544,
         n19545, n19546, n19547, n19549, n19550, n19551, n19552, n19554,
         n19555, n19556, n19557, n19558, n19559, n19561, n19562, n19564,
         n19565, n19566, n19567, n19568, n19570, n19571, n19573, n19574,
         n19575, n19577, n19578, n19579, n19580, n19582, n19583, n19584,
         n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592,
         n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19609, n19610,
         n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618,
         n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626,
         n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634,
         n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642,
         n19644, n19647, n19648, n19649, n19651, n19653, n19654, n19655,
         n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664,
         n19666, n19667, n19668, n19669, n19671, n19672, n19673, n19675,
         n19676, n19677, n19679, n19680, n19681, n19682, n19683, n19684,
         n19685, n19686, n19687, n19689, n19690, n19691, n19693, n19694,
         n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702,
         n19703, n19705, n19706, n19707, n19708, n19709, n19710, n19711,
         n19712, n19713, n19716, n19717, n19718, n19719, n19721, n19722,
         n19723, n19724, n19726, n19727, n19728, n19729, n19730, n19731,
         n19732, n19733, n19734, n19735, n19736, n19737, n19739, n19740,
         n19741, n19742, n19743, n19744, n19746, n19748, n19749, n19750,
         n19751, n19752, n19754, n19755, n19757, n19759, n19761, n19763,
         n19764, n19766, n19767, n19768, n19769, n19770, n19771, n19772,
         n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780,
         n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789,
         n19790, n19791, n19792, n19794, n19796, n19798, n19799, n19800,
         n19801, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19814, n19816, n19817, n19818, n19819,
         n19820, n19822, n19823, n19824, n19825, n19826, n19827, n19828,
         n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19837,
         n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845,
         n19846, n19847, n19849, n19850, n19851, n19853, n19854, n19855,
         n19856, n19857, n19861, n19862, n19863, n19864, n19865, n19866,
         n19867, n19868, n19869, n19871, n19872, n19874, n19875, n19876,
         n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885,
         n19886, n19888, n19889, n19891, n19892, n19893, n19894, n19896,
         n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904,
         n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912,
         n19913, n19914, n19915, n19916, n19917, n19918, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19938,
         n19939, n19940, n19941, n19942, n19943, n19944, n19947, n19948,
         n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956,
         n19957, n19958, n19959, n19960, n19961, n19962, n19964, n19965,
         n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19974,
         n19975, n19976, n19977, n19979, n19984, n19986, n19987, n19990,
         n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998,
         n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007,
         n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015,
         n20017, n20018, n20019, n20020, n20021, n20022, n20024, n20025,
         n20026, n20028, n20029, n20032, n20033, n20034, n20035, n20036,
         n20037, n20038, n20039, n20040, n20042, n20043, n20044, n20045,
         n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054,
         n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062,
         n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070,
         n20071, n20072, n20073, n20075, n20076, n20077, n20078, n20079,
         n20080, n20081, n20083, n20084, n20085, n20086, n20087, n20088,
         n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096,
         n20097, n20098, n20099, n20100, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123,
         n20124, n20125, n20126, n20127, n20128, n20130, n20132, n20133,
         n20134, n20135, n20136, n20137, n20138, n20139, n20141, n20142,
         n20143, n20144, n20147, n20148, n20149, n20150, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20186, n20187,
         n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20196,
         n20197, n20199, n20200, n20201, n20202, n20203, n20204, n20205,
         n20206, n20207, n20208, n20209, n20210, n20213, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20233, n20234,
         n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242,
         n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20251,
         n20252, n20254, n20255, n20256, n20257, n20258, n20259, n20261,
         n20263, n20266, n20267, n20268, n20269, n20270, n20271, n20272,
         n20273, n20274, n20275, n20276, n20277, n20278, n20280, n20281,
         n20282, n20283, n20284, n20285, n20287, n20288, n20289, n20290,
         n20291, n20292, n20293, n20294, n20296, n20297, n20298, n20299,
         n20300, n20301, n20302, n20304, n20305, n20306, n20308, n20309,
         n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317,
         n20318, n20319, n20321, n20322, n20323, n20324, n20325, n20327,
         n20328, n20329, n20330, n20332, n20333, n20334, n20335, n20336,
         n20337, n20338, n20339, n20340, n20341, n20342, n20344, n20345,
         n20347, n20349, n20350, n20351, n20352, n20353, n20354, n20356,
         n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364,
         n20366, n20367, n20368, n20371, n20373, n20374, n20375, n20376,
         n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384,
         n20385, n20386, n20387, n20389, n20390, n20392, n20393, n20395,
         n20396, n20397, n20399, n20400, n20401, n20403, n20404, n20405,
         n20406, n20407, n20408, n20410, n20411, n20412, n20413, n20414,
         n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422,
         n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430,
         n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438,
         n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446,
         n20447, n20449, n20450, n20451, n20452, n20453, n20454, n20455,
         n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463,
         n20464, n20466, n20467, n20468, n20471, n20472, n20475, n20476,
         n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486,
         n20487, n20489, n20490, n20492, n20493, n20494, n20495, n20496,
         n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504,
         n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512,
         n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520,
         n20521, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20531, n20533, n20534, n20535, n20536, n20537, n20538, n20540,
         n20541, n20542, n20545, n20546, n20547, n20548, n20549, n20550,
         n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558,
         n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20568,
         n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576,
         n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584,
         n20585, n20586, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20598, n20599, n20600, n20601, n20602, n20603,
         n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20612,
         n20613, n20614, n20615, n20616, n20617, n20619, n20620, n20621,
         n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629,
         n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20639,
         n20640, n20641, n20642, n20644, n20645, n20647, n20648, n20649,
         n20650, n20651, n20652, n20654, n20657, n20658, n20659, n20660,
         n20661, n20662, n20663, n20664, n20667, n20668, n20669, n20670,
         n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678,
         n20679, n20680, n20682, n20684, n20686, n20687, n20688, n20690,
         n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698,
         n20699, n20700, n20702, n20703, n20704, n20705, n20706, n20707,
         n20708, n20709, n20710, n20711, n20712, n20713, n20715, n20716,
         n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724,
         n20726, n20727, n20729, n20730, n20731, n20732, n20733, n20736,
         n20737, n20738, n20739, n20740, n20742, n20743, n20744, n20746,
         n20747, n20748, n20749, n20751, n20752, n20753, n20754, n20755,
         n20756, n20757, n20758, n20759, n20762, n20764, n20765, n20766,
         n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774,
         n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782,
         n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790,
         n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798,
         n20799, n20801, n20802, n20803, n20804, n20806, n20807, n20808,
         n20809, n20810, n20813, n20815, n20816, n20818, n20819, n20820,
         n20821, n20822, n20823, n20824, n20825, n20827, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20848, n20849, n20850,
         n20851, n20852, n20853, n20855, n20856, n20857, n20858, n20859,
         n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867,
         n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875,
         n20877, n20879, n20880, n20881, n20882, n20883, n20884, n20885,
         n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893,
         n20894, n20895, n20896, n20897, n20899, n20900, n20902, n20904,
         n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912,
         n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920,
         n20921, n20922, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20938,
         n20939, n20940, n20941, n20944, n20945, n20946, n20947, n20949,
         n20950, n20951, n20953, n20954, n20955, n20956, n20957, n20958,
         n20959, n20960, n20961, n20962, n20963, n20964, n20966, n20967,
         n20968, n20970, n20971, n20972, n20974, n20975, n20976, n20977,
         n20978, n20979, n20982, n20983, n20984, n20985, n20986, n20987,
         n20988, n20989, n20990, n20992, n20993, n20994, n20995, n20996,
         n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004,
         n21005, n21006, n21007, n21009, n21010, n21011, n21012, n21014,
         n21015, n21016, n21017, n21018, n21019, n21020, n21022, n21023,
         n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031,
         n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039,
         n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047,
         n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055,
         n21056, n21057, n21058, n21059, n21060, n21061, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21093, n21095, n21096, n21097, n21098, n21099,
         n21100, n21101, n21104, n21107, n21109, n21110, n21112, n21113,
         n21114, n21115, n21117, n21118, n21119, n21120, n21121, n21122,
         n21123, n21125, n21126, n21127, n21129, n21131, n21132, n21134,
         n21136, n21137, n21138, n21139, n21140, n21141, n21143, n21145,
         n21146, n21147, n21148, n21149, n21151, n21152, n21153, n21154,
         n21155, n21156, n21158, n21159, n21160, n21161, n21162, n21163,
         n21164, n21165, n21167, n21168, n21169, n21170, n21171, n21172,
         n21173, n21175, n21176, n21178, n21179, n21180, n21181, n21182,
         n21183, n21184, n21187, n21188, n21189, n21190, n21191, n21192,
         n21193, n21195, n21196, n21198, n21199, n21200, n21202, n21203,
         n21204, n21206, n21207, n21209, n21210, n21211, n21212, n21213,
         n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221,
         n21222, n21223, n21224, n21225, n21226, n21228, n21230, n21232,
         n21233, n21234, n21235, n21237, n21239, n21240, n21241, n21243,
         n21244, n21247, n21248, n21249, n21251, n21252, n21253, n21254,
         n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21263,
         n21264, n21265, n21266, n21267, n21269, n21270, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21289, n21291, n21292,
         n21295, n21297, n21298, n21299, n21300, n21302, n21303, n21304,
         n21305, n21306, n21307, n21308, n21309, n21310, n21311, n21312,
         n21313, n21314, n21315, n21316, n21317, n21320, n21321, n21322,
         n21323, n21324, n21325, n21326, n21328, n21330, n21331, n21332,
         n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341,
         n21343, n21345, n21346, n21347, n21348, n21349, n21350, n21351,
         n21353, n21354, n21356, n21357, n21358, n21359, n21361, n21362,
         n21363, n21365, n21366, n21367, n21368, n21369, n21370, n21372,
         n21373, n21374, n21375, n21377, n21378, n21379, n21381, n21382,
         n21383, n21385, n21386, n21387, n21389, n21390, n21391, n21392,
         n21393, n21394, n21395, n21396, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21410,
         n21411, n21412, n21413, n21414, n21415, n21416, n21418, n21419,
         n21420, n21421, n21423, n21424, n21426, n21427, n21428, n21429,
         n21430, n21431, n21432, n21433, n21434, n21437, n21438, n21439,
         n21440, n21441, n21442, n21443, n21445, n21447, n21448, n21449,
         n21451, n21452, n21453, n21454, n21455, n21457, n21458, n21459,
         n21460, n21461, n21462, n21463, n21465, n21466, n21467, n21468,
         n21469, n21470, n21471, n21472, n21473, n21475, n21477, n21478,
         n21479, n21480, n21481, n21482, n21483, n21484, n21485, n21487,
         n21488, n21489, n21490, n21491, n21492, n21494, n21495, n21496,
         n21497, n21498, n21499, n21500, n21501, n21502, n21503, n21504,
         n21505, n21506, n21509, n21510, n21512, n21514, n21517, n21518,
         n21519, n21520, n21521, n21522, n21523, n21524, n21525, n21527,
         n21529, n21530, n21531, n21532, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21542, n21544, n21545, n21546, n21548,
         n21549, n21550, n21551, n21553, n21554, n21555, n21556, n21558,
         n21559, n21560, n21561, n21562, n21564, n21566, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21576, n21577, n21579,
         n21580, n21581, n21582, n21583, n21585, n21586, n21587, n21588,
         n21589, n21590, n21591, n21592, n21594, n21595, n21596, n21597,
         n21599, n21600, n21601, n21602, n21603, n21604, n21606, n21607,
         n21608, n21609, n21610, n21612, n21613, n21614, n21615, n21616,
         n21617, n21618, n21619, n21620, n21621, n21622, n21623, n21624,
         n21625, n21626, n21627, n21628, n21629, n21630, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21655, n21656, n21657, n21658,
         n21659, n21660, n21661, n21662, n21663, n21664, n21665, n21666,
         n21667, n21668, n21669, n21671, n21672, n21673, n21674, n21676,
         n21678, n21680, n21681, n21682, n21683, n21684, n21685, n21686,
         n21687, n21688, n21690, n21691, n21692, n21693, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21704, n21705, n21706,
         n21707, n21708, n21709, n21710, n21711, n21712, n21713, n21715,
         n21716, n21717, n21719, n21720, n21721, n21722, n21723, n21724,
         n21725, n21726, n21727, n21728, n21730, n21731, n21732, n21733,
         n21736, n21737, n21738, n21739, n21740, n21741, n21742, n21743,
         n21744, n21746, n21747, n21748, n21749, n21750, n21752, n21753,
         n21754, n21755, n21756, n21757, n21759, n21760, n21761, n21762,
         n21763, n21764, n21765, n21766, n21767, n21768, n21769, n21771,
         n21772, n21775, n21776, n21777, n21778, n21779, n21780, n21781,
         n21785, n21786, n21789, n21790, n21791, n21792, n21793, n21794,
         n21795, n21796, n21797, n21799, n21800, n21801, n21804, n21805,
         n21806, n21808, n21809, n21811, n21812, n21813, n21814, n21815,
         n21816, n21817, n21818, n21819, n21820, n21821, n21823, n21824,
         n21825, n21826, n21827, n21828, n21829, n21830, n21831, n21832,
         n21833, n21834, n21835, n21836, n21837, n21838, n21839, n21840,
         n21841, n21842, n21843, n21844, n21846, n21847, n21848, n21849,
         n21850, n21852, n21853, n21854, n21855, n21856, n21857, n21858,
         n21859, n21860, n21861, n21862, n21863, n21864, n21865, n21866,
         n21867, n21869, n21870, n21871, n21872, n21873, n21874, n21875,
         n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883,
         n21884, n21885, n21886, n21887, n21888, n21889, n21891, n21892,
         n21893, n21894, n21896, n21898, n21899, n21900, n21901, n21902,
         n21903, n21905, n21906, n21907, n21909, n21910, n21911, n21912,
         n21913, n21915, n21916, n21918, n21919, n21920, n21921, n21923,
         n21924, n21925, n21926, n21927, n21929, n21930, n21931, n21932,
         n21933, n21934, n21935, n21936, n21937, n21938, n21939, n21940,
         n21941, n21944, n21945, n21946, n21947, n21948, n21949, n21950,
         n21951, n21952, n21953, n21956, n21957, n21958, n21959, n21960,
         n21961, n21962, n21963, n21964, n21965, n21967, n21968, n21970,
         n21971, n21972, n21974, n21975, n21979, n21980, n21981, n21983,
         n21984, n21985, n21986, n21988, n21990, n21992, n21993, n21994,
         n21995, n21996, n21997, n21998, n21999, n22000, n22002, n22003,
         n22004, n22005, n22006, n22008, n22011, n22012, n22013, n22014,
         n22015, n22016, n22017, n22018, n22019, n22020, n22021, n22022,
         n22023, n22024, n22025, n22026, n22027, n22028, n22029, n22030,
         n22031, n22032, n22033, n22034, n22035, n22036, n22037, n22038,
         n22039, n22040, n22041, n22042, n22043, n22044, n22045, n22046,
         n22047, n22048, n22049, n22051, n22053, n22054, n22055, n22056,
         n22057, n22058, n22059, n22060, n22061, n22062, n22063, n22064,
         n22066, n22067, n22070, n22071, n22072, n22075, n22076, n22078,
         n22079, n22080, n22081, n22082, n22083, n22084, n22085, n22086,
         n22087, n22088, n22089, n22090, n22091, n22092, n22093, n22094,
         n22096, n22098, n22099, n22100, n22102, n22103, n22104, n22105,
         n22107, n22108, n22109, n22110, n22111, n22112, n22113, n22114,
         n22115, n22118, n22119, n22120, n22121, n22123, n22125, n22126,
         n22127, n22128, n22130, n22131, n22132, n22133, n22134, n22136,
         n22137, n22138, n22139, n22140, n22141, n22142, n22143, n22144,
         n22145, n22146, n22147, n22148, n22149, n22150, n22151, n22152,
         n22153, n22154, n22155, n22156, n22157, n22158, n22160, n22161,
         n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169,
         n22171, n22172, n22173, n22174, n22175, n22176, n22177, n22178,
         n22179, n22180, n22181, n22182, n22183, n22185, n22186, n22187,
         n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195,
         n22196, n22197, n22198, n22199, n22200, n22201, n22202, n22203,
         n22205, n22206, n22208, n22210, n22211, n22213, n22214, n22216,
         n22217, n22218, n22220, n22221, n22222, n22223, n22224, n22225,
         n22226, n22227, n22229, n22230, n22231, n22232, n22233, n22235,
         n22237, n22238, n22239, n22240, n22241, n22242, n22243, n22244,
         n22246, n22247, n22248, n22249, n22250, n22251, n22252, n22253,
         n22254, n22255, n22256, n22258, n22259, n22260, n22261, n22264,
         n22265, n22266, n22267, n22268, n22269, n22271, n22273, n22274,
         n22275, n22276, n22277, n22280, n22282, n22283, n22284, n22285,
         n22286, n22287, n22288, n22289, n22291, n22292, n22293, n22294,
         n22295, n22296, n22297, n22299, n22300, n22301, n22302, n22303,
         n22305, n22306, n22307, n22308, n22309, n22310, n22311, n22312,
         n22313, n22314, n22315, n22317, n22318, n22319, n22320, n22322,
         n22324, n22325, n22326, n22327, n22328, n22329, n22330, n22332,
         n22333, n22335, n22336, n22337, n22338, n22339, n22340, n22342,
         n22343, n22344, n22348, n22350, n22351, n22353, n22356, n22357,
         n22358, n22359, n22360, n22361, n22362, n22363, n22364, n22366,
         n22367, n22368, n22369, n22372, n22375, n22377, n22379, n22380,
         n22382, n22383, n22384, n22385, n22386, n22387, n22388, n22389,
         n22390, n22391, n22392, n22393, n22394, n22396, n22397, n22398,
         n22399, n22400, n22401, n22402, n22403, n22404, n22406, n22407,
         n22408, n22409, n22410, n22411, n22412, n22413, n22414, n22415,
         n22416, n22418, n22420, n22421, n22422, n22424, n22425, n22426,
         n22427, n22428, n22429, n22430, n22431, n22433, n22434, n22435,
         n22436, n22437, n22438, n22439, n22441, n22442, n22443, n22444,
         n22446, n22448, n22449, n22450, n22452, n22454, n22455, n22457,
         n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22466,
         n22467, n22468, n22470, n22471, n22472, n22473, n22474, n22475,
         n22476, n22477, n22478, n22479, n22480, n22482, n22483, n22484,
         n22486, n22487, n22488, n22489, n22490, n22491, n22495, n22496,
         n22497, n22498, n22499, n22500, n22502, n22503, n22504, n22505,
         n22508, n22509, n22510, n22511, n22512, n22513, n22515, n22516,
         n22517, n22518, n22521, n22522, n22523, n22524, n22526, n22527,
         n22529, n22530, n22531, n22534, n22535, n22536, n22537, n22539,
         n22540, n22542, n22543, n22544, n22546, n22547, n22549, n22550,
         n22551, n22552, n22553, n22555, n22556, n22557, n22558, n22560,
         n22561, n22562, n22563, n22564, n22565, n22566, n22567, n22568,
         n22569, n22570, n22571, n22572, n22573, n22574, n22575, n22576,
         n22577, n22578, n22579, n22580, n22581, n22582, n22583, n22584,
         n22585, n22586, n22587, n22588, n22589, n22590, n22591, n22592,
         n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22602,
         n22603, n22604, n22605, n22606, n22607, n22608, n22610, n22612,
         n22613, n22614, n22615, n22616, n22617, n22618, n22619, n22620,
         n22621, n22622, n22623, n22624, n22625, n22626, n22627, n22628,
         n22629, n22631, n22633, n22634, n22635, n22636, n22637, n22638,
         n22639, n22640, n22641, n22642, n22643, n22644, n22645, n22646,
         n22647, n22648, n22650, n22651, n22652, n22653, n22654, n22655,
         n22656, n22657, n22658, n22659, n22660, n22662, n22663, n22664,
         n22665, n22666, n22667, n22669, n22670, n22671, n22672, n22673,
         n22674, n22677, n22678, n22679, n22680, n22681, n22682, n22683,
         n22685, n22686, n22688, n22689, n22690, n22691, n22692, n22693,
         n22694, n22697, n22698, n22699, n22701, n22704, n22705, n22706,
         n22707, n22709, n22710, n22711, n22712, n22714, n22715, n22716,
         n22717, n22719, n22720, n22721, n22722, n22723, n22724, n22725,
         n22726, n22728, n22729, n22730, n22731, n22732, n22737, n22738,
         n22739, n22740, n22741, n22743, n22744, n22745, n22747, n22748,
         n22749, n22750, n22751, n22752, n22753, n22754, n22755, n22756,
         n22757, n22758, n22759, n22760, n22761, n22762, n22765, n22766,
         n22767, n22768, n22769, n22770, n22772, n22773, n22774, n22775,
         n22776, n22777, n22778, n22779, n22780, n22781, n22783, n22784,
         n22785, n22786, n22789, n22790, n22791, n22792, n22795, n22798,
         n22799, n22800, n22801, n22803, n22804, n22805, n22806, n22807,
         n22808, n22809, n22810, n22811, n22813, n22814, n22815, n22816,
         n22817, n22818, n22819, n22820, n22822, n22823, n22824, n22825,
         n22826, n22827, n22828, n22830, n22831, n22832, n22833, n22834,
         n22835, n22836, n22837, n22838, n22839, n22840, n22841, n22842,
         n22843, n22845, n22848, n22849, n22851, n22852, n22853, n22855,
         n22856, n22857, n22859, n22860, n22861, n22862, n22863, n22864,
         n22865, n22866, n22867, n22868, n22869, n22870, n22871, n22872,
         n22873, n22874, n22875, n22876, n22877, n22878, n22879, n22880,
         n22881, n22882, n22883, n22884, n22885, n22886, n22888, n22889,
         n22890, n22892, n22893, n22894, n22895, n22896, n22897, n22899,
         n22900, n22901, n22904, n22905, n22906, n22907, n22908, n22909,
         n22910, n22913, n22914, n22915, n22916, n22919, n22920, n22921,
         n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929,
         n22931, n22932, n22933, n22934, n22935, n22936, n22937, n22938,
         n22940, n22942, n22943, n22944, n22945, n22946, n22948, n22949,
         n22950, n22951, n22952, n22953, n22954, n22955, n22956, n22957,
         n22959, n22960, n22961, n22962, n22963, n22964, n22965, n22966,
         n22967, n22968, n22969, n22970, n22971, n22972, n22973, n22974,
         n22977, n22978, n22979, n22981, n22982, n22983, n22984, n22985,
         n22986, n22988, n22990, n22992, n22993, n22996, n22997, n22999,
         n23000, n23002, n23003, n23004, n23005, n23006, n23007, n23008,
         n23009, n23010, n23011, n23012, n23013, n23014, n23015, n23016,
         n23017, n23018, n23021, n23022, n23023, n23024, n23025, n23026,
         n23027, n23028, n23029, n23030, n23031, n23032, n23033, n23034,
         n23035, n23037, n23038, n23039, n23040, n23041, n23042, n23043,
         n23045, n23046, n23047, n23048, n23049, n23050, n23051, n23052,
         n23053, n23054, n23055, n23056, n23057, n23058, n23060, n23062,
         n23064, n23065, n23066, n23067, n23068, n23069, n23070, n23071,
         n23072, n23073, n23074, n23075, n23076, n23077, n23079, n23080,
         n23081, n23082, n23083, n23084, n23085, n23086, n23087, n23088,
         n23089, n23090, n23092, n23093, n23094, n23096, n23100, n23101,
         n23103, n23104, n23105, n23106, n23107, n23108, n23109, n23110,
         n23111, n23112, n23113, n23115, n23116, n23117, n23118, n23119,
         n23120, n23121, n23122, n23123, n23124, n23125, n23126, n23127,
         n23128, n23130, n23131, n23132, n23136, n23137, n23138, n23139,
         n23140, n23143, n23144, n23145, n23146, n23150, n23151, n23152,
         n23153, n23154, n23155, n23156, n23157, n23158, n23162, n23163,
         n23164, n23165, n23166, n23167, n23168, n23169, n23170, n23171,
         n23173, n23174, n23176, n23177, n23178, n23179, n23180, n23181,
         n23182, n23183, n23184, n23185, n23186, n23188, n23189, n23190,
         n23191, n23192, n23194, n23196, n23197, n23198, n23199, n23200,
         n23201, n23202, n23203, n23205, n23206, n23207, n23209, n23210,
         n23211, n23212, n23213, n23216, n23217, n23218, n23219, n23220,
         n23221, n23222, n23223, n23224, n23226, n23227, n23228, n23229,
         n23230, n23231, n23232, n23233, n23234, n23236, n23237, n23238,
         n23239, n23240, n23241, n23242, n23243, n23244, n23245, n23246,
         n23247, n23248, n23249, n23250, n23251, n23253, n23254, n23255,
         n23256, n23257, n23258, n23259, n23260, n23261, n23262, n23263,
         n23264, n23265, n23266, n23267, n23268, n23269, n23270, n23271,
         n23272, n23273, n23274, n23275, n23276, n23277, n23278, n23279,
         n23280, n23282, n23283, n23284, n23285, n23286, n23287, n23288,
         n23289, n23290, n23291, n23292, n23293, n23294, n23295, n23296,
         n23297, n23298, n23299, n23300, n23301, n23302, n23303, n23304,
         n23306, n23307, n23308, n23310, n23311, n23312, n23313, n23314,
         n23315, n23316, n23318, n23319, n23320, n23321, n23322, n23324,
         n23326, n23328, n23329, n23330, n23331, n23332, n23333, n23334,
         n23335, n23336, n23337, n23338, n23340, n23341, n23342, n23343,
         n23344, n23346, n23347, n23348, n23349, n23350, n23351, n23352,
         n23353, n23354, n23355, n23356, n23358, n23359, n23361, n23362,
         n23363, n23364, n23366, n23367, n23368, n23369, n23370, n23371,
         n23372, n23373, n23374, n23375, n23376, n23377, n23382, n23383,
         n23384, n23385, n23386, n23387, n23388, n23389, n23390, n23391,
         n23393, n23395, n23396, n23397, n23398, n23399, n23400, n23402,
         n23403, n23404, n23405, n23406, n23407, n23408, n23411, n23412,
         n23413, n23414, n23415, n23417, n23419, n23420, n23421, n23422,
         n23424, n23425, n23426, n23427, n23429, n23430, n23431, n23432,
         n23433, n23435, n23436, n23437, n23438, n23439, n23440, n23441,
         n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449,
         n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457,
         n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465,
         n23467, n23468, n23469, n23470, n23471, n23472, n23473, n23474,
         n23475, n23476, n23478, n23479, n23480, n23481, n23482, n23483,
         n23484, n23485, n23486, n23487, n23488, n23489, n23490, n23491,
         n23493, n23494, n23495, n23496, n23497, n23498, n23499, n23501,
         n23502, n23503, n23504, n23505, n23506, n23507, n23508, n23509,
         n23510, n23511, n23512, n23513, n23514, n23516, n23517, n23518,
         n23519, n23520, n23521, n23522, n23523, n23524, n23525, n23526,
         n23527, n23528, n23529, n23530, n23532, n23533, n23534, n23535,
         n23536, n23537, n23538, n23539, n23540, n23542, n23543, n23544,
         n23547, n23548, n23549, n23550, n23551, n23552, n23553, n23554,
         n23555, n23556, n23558, n23559, n23560, n23561, n23562, n23564,
         n23565, n23566, n23567, n23569, n23570, n23571, n23572, n23573,
         n23574, n23575, n23576, n23577, n23578, n23579, n23581, n23582,
         n23583, n23584, n23586, n23587, n23588, n23590, n23593, n23594,
         n23595, n23597, n23598, n23600, n23601, n23602, n23603, n23604,
         n23605, n23606, n23608, n23609, n23610, n23611, n23612, n23613,
         n23616, n23618, n23620, n23621, n23622, n23623, n23624, n23625,
         n23626, n23627, n23628, n23629, n23631, n23632, n23633, n23634,
         n23635, n23636, n23637, n23638, n23639, n23640, n23642, n23643,
         n23644, n23646, n23647, n23649, n23650, n23651, n23653, n23654,
         n23655, n23656, n23657, n23658, n23659, n23660, n23663, n23664,
         n23665, n23666, n23668, n23669, n23670, n23671, n23672, n23675,
         n23676, n23677, n23679, n23680, n23681, n23682, n23683, n23684,
         n23685, n23688, n23689, n23690, n23691, n23692, n23694, n23695,
         n23696, n23697, n23698, n23699, n23701, n23702, n23703, n23704,
         n23705, n23706, n23707, n23708, n23709, n23710, n23711, n23712,
         n23713, n23714, n23715, n23717, n23718, n23719, n23720, n23721,
         n23722, n23723, n23724, n23726, n23727, n23728, n23729, n23730,
         n23731, n23735, n23736, n23737, n23738, n23739, n23740, n23741,
         n23742, n23745, n23746, n23747, n23748, n23749, n23750, n23752,
         n23753, n23754, n23755, n23756, n23757, n23758, n23759, n23760,
         n23763, n23764, n23765, n23766, n23767, n23768, n23769, n23770,
         n23771, n23772, n23773, n23775, n23776, n23777, n23778, n23780,
         n23781, n23782, n23784, n23785, n23786, n23787, n23788, n23790,
         n23791, n23792, n23793, n23794, n23795, n23796, n23797, n23798,
         n23799, n23800, n23801, n23802, n23803, n23804, n23805, n23806,
         n23807, n23808, n23809, n23811, n23812, n23813, n23815, n23816,
         n23817, n23818, n23819, n23821, n23822, n23823, n23824, n23825,
         n23826, n23827, n23828, n23832, n23833, n23834, n23835, n23840,
         n23841, n23842, n23843, n23847, n23848, n23849, n23850, n23851,
         n23852, n23853, n23855, n23856, n23857, n23858, n23859, n23860,
         n23862, n23864, n23866, n23867, n23868, n23869, n23870, n23871,
         n23872, n23873, n23874, n23875, n23876, n23877, n23878, n23880,
         n23881, n23882, n23884, n23885, n23886, n23887, n23888, n23889,
         n23891, n23892, n23894, n23895, n23896, n23897, n23899, n23901,
         n23902, n23903, n23904, n23905, n23906, n23910, n23912, n23914,
         n23915, n23916, n23917, n23918, n23919, n23920, n23921, n23922,
         n23923, n23924, n23925, n23927, n23928, n23929, n23930, n23931,
         n23932, n23933, n23934, n23935, n23936, n23938, n23939, n23940,
         n23942, n23943, n23944, n23945, n23946, n23947, n23949, n23950,
         n23951, n23952, n23953, n23954, n23955, n23956, n23957, n23958,
         n23959, n23960, n23961, n23962, n23964, n23965, n23966, n23967,
         n23968, n23969, n23970, n23971, n23972, n23973, n23974, n23975,
         n23976, n23978, n23981, n23982, n23984, n23987, n23988, n23989,
         n23990, n23991, n23992, n23994, n23995, n23996, n23997, n23998,
         n23999, n24000, n24001, n24002, n24004, n24005, n24007, n24008,
         n24009, n24010, n24011, n24012, n24013, n24014, n24015, n24016,
         n24017, n24018, n24020, n24021, n24024, n24025, n24027, n24029,
         n24030, n24031, n24032, n24033, n24034, n24035, n24036, n24038,
         n24039, n24040, n24041, n24042, n24043, n24044, n24046, n24047,
         n24048, n24049, n24050, n24051, n24052, n24053, n24056, n24057,
         n24059, n24060, n24061, n24062, n24063, n24064, n24065, n24066,
         n24067, n24069, n24071, n24072, n24073, n24074, n24075, n24076,
         n24077, n24078, n24079, n24080, n24081, n24082, n24083, n24084,
         n24085, n24086, n24087, n24089, n24090, n24091, n24092, n24093,
         n24094, n24095, n24096, n24097, n24098, n24099, n24101, n24102,
         n24103, n24104, n24106, n24107, n24108, n24109, n24110, n24111,
         n24112, n24114, n24115, n24116, n24117, n24118, n24119, n24120,
         n24121, n24123, n24124, n24125, n24126, n24127, n24128, n24129,
         n24130, n24131, n24132, n24133, n24134, n24135, n24137, n24138,
         n24139, n24140, n24141, n24142, n24143, n24144, n24147, n24148,
         n24149, n24150, n24152, n24153, n24154, n24156, n24157, n24158,
         n24159, n24161, n24162, n24163, n24164, n24165, n24166, n24167,
         n24168, n24169, n24171, n24172, n24173, n24174, n24176, n24177,
         n24178, n24179, n24180, n24181, n24182, n24183, n24185, n24186,
         n24187, n24188, n24189, n24190, n24191, n24193, n24194, n24195,
         n24196, n24197, n24198, n24199, n24200, n24201, n24202, n24204,
         n24205, n24206, n24207, n24208, n24209, n24210, n24211, n24212,
         n24213, n24214, n24215, n24216, n24217, n24218, n24219, n24220,
         n24221, n24222, n24223, n24224, n24225, n24226, n24227, n24228,
         n24229, n24230, n24231, n24232, n24233, n24234, n24235, n24236,
         n24237, n24238, n24239, n24240, n24241, n24242, n24243, n24244,
         n24245, n24246, n24248, n24249, n24250, n24251, n24253, n24254,
         n24255, n24256, n24257, n24259, n24260, n24262, n24263, n24265,
         n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273,
         n24275, n24276, n24277, n24278, n24279, n24280, n24281, n24283,
         n24284, n24285, n24286, n24288, n24289, n24290, n24292, n24293,
         n24294, n24295, n24296, n24297, n24299, n24300, n24301, n24302,
         n24304, n24305, n24306, n24308, n24309, n24310, n24311, n24312,
         n24313, n24314, n24315, n24316, n24317, n24318, n24319, n24321,
         n24322, n24324, n24325, n24326, n24327, n24328, n24329, n24330,
         n24331, n24332, n24333, n24334, n24335, n24336, n24337, n24338,
         n24339, n24340, n24341, n24342, n24343, n24344, n24346, n24347,
         n24348, n24349, n24350, n24351, n24353, n24354, n24355, n24356,
         n24357, n24358, n24359, n24360, n24361, n24362, n24364, n24365,
         n24368, n24369, n24370, n24371, n24372, n24373, n24374, n24375,
         n24376, n24377, n24378, n24379, n24382, n24383, n24384, n24385,
         n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393,
         n24394, n24395, n24398, n24399, n24401, n24402, n24403, n24404,
         n24405, n24407, n24408, n24409, n24410, n24411, n24412, n24413,
         n24415, n24416, n24417, n24418, n24419, n24421, n24422, n24423,
         n24424, n24425, n24426, n24427, n24428, n24429, n24430, n24431,
         n24432, n24433, n24434, n24435, n24436, n24437, n24438, n24439,
         n24440, n24441, n24442, n24443, n24444, n24445, n24446, n24447,
         n24448, n24449, n24450, n24451, n24452, n24453, n24454, n24455,
         n24456, n24457, n24459, n24460, n24461, n24462, n24463, n24466,
         n24467, n24469, n24470, n24471, n24472, n24473, n24474, n24475,
         n24476, n24477, n24478, n24479, n24481, n24482, n24484, n24485,
         n24486, n24487, n24488, n24489, n24491, n24492, n24493, n24494,
         n24495, n24496, n24497, n24498, n24499, n24500, n24501, n24502,
         n24503, n24504, n24505, n24506, n24507, n24508, n24511, n24512,
         n24513, n24514, n24515, n24516, n24517, n24518, n24519, n24520,
         n24521, n24522, n24523, n24524, n24525, n24526, n24527, n24528,
         n24529, n24531, n24532, n24533, n24536, n24537, n24538, n24539,
         n24540, n24541, n24542, n24543, n24544, n24545, n24546, n24547,
         n24548, n24549, n24551, n24552, n24553, n24554, n24556, n24557,
         n24559, n24560, n24561, n24562, n24563, n24564, n24565, n24567,
         n24568, n24569, n24570, n24572, n24573, n24574, n24575, n24576,
         n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585,
         n24587, n24588, n24590, n24591, n24592, n24593, n24595, n24596,
         n24597, n24598, n24600, n24602, n24603, n24604, n24605, n24606,
         n24607, n24609, n24610, n24611, n24613, n24615, n24616, n24617,
         n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625,
         n24626, n24628, n24629, n24631, n24632, n24633, n24634, n24635,
         n24636, n24637, n24638, n24639, n24642, n24643, n24644, n24645,
         n24646, n24647, n24648, n24649, n24650, n24651, n24652, n24653,
         n24654, n24655, n24656, n24657, n24658, n24659, n24660, n24662,
         n24664, n24665, n24666, n24667, n24668, n24671, n24672, n24673,
         n24674, n24675, n24676, n24678, n24679, n24680, n24681, n24682,
         n24683, n24684, n24685, n24686, n24687, n24688, n24689, n24691,
         n24692, n24693, n24695, n24696, n24697, n24698, n24699, n24701,
         n24702, n24703, n24704, n24705, n24707, n24708, n24709, n24710,
         n24711, n24712, n24713, n24714, n24715, n24716, n24717, n24718,
         n24719, n24720, n24721, n24723, n24724, n24725, n24726, n24728,
         n24729, n24730, n24732, n24733, n24734, n24735, n24737, n24738,
         n24740, n24741, n24742, n24743, n24744, n24745, n24746, n24747,
         n24748, n24749, n24750, n24751, n24752, n24753, n24754, n24755,
         n24756, n24757, n24758, n24759, n24760, n24761, n24762, n24763,
         n24764, n24766, n24768, n24769, n24770, n24771, n24773, n24774,
         n24776, n24777, n24778, n24779, n24780, n24781, n24782, n24783,
         n24785, n24786, n24787, n24788, n24789, n24790, n24792, n24793,
         n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801,
         n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809,
         n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817,
         n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825,
         n24826, n24828, n24829, n24830, n24831, n24832, n24833, n24834,
         n24835, n24836, n24837, n24838, n24839, n24840, n24841, n24842,
         n24843, n24845, n24846, n24847, n24848, n24849, n24852, n24853,
         n24854, n24855, n24856, n24857, n24860, n24861, n24862, n24863,
         n24864, n24865, n24866, n24867, n24869, n24870, n24873, n24874,
         n24875, n24876, n24877, n24878, n24879, n24880, n24881, n24882,
         n24883, n24884, n24885, n24886, n24888, n24889, n24892, n24893,
         n24894, n24895, n24896, n24897, n24899, n24901, n24902, n24903,
         n24904, n24905, n24906, n24907, n24908, n24909, n24910, n24911,
         n24912, n24913, n24914, n24915, n24916, n24917, n24918, n24919,
         n24920, n24921, n24922, n24923, n24924, n24925, n24926, n24927,
         n24928, n24929, n24930, n24931, n24932, n24933, n24934, n24936,
         n24937, n24938, n24939, n24940, n24941, n24942, n24943, n24944,
         n24945, n24946, n24947, n24948, n24949, n24950, n24953, n24954,
         n24955, n24956, n24957, n24958, n24959, n24960, n24961, n24962,
         n24964, n24965, n24966, n24967, n24968, n24969, n24970, n24972,
         n24973, n24974, n24975, n24976, n24977, n24981, n24983, n24984,
         n24985, n24988, n24989, n24991, n24992, n24993, n24994, n24995,
         n24996, n24997, n24998, n24999, n25000, n25001, n25002, n25003,
         n25004, n25005, n25006, n25007, n25008, n25009, n25010, n25012,
         n25013, n25014, n25015, n25017, n25019, n25020, n25021, n25022,
         n25023, n25024, n25025, n25026, n25027, n25028, n25029, n25031,
         n25033, n25034, n25035, n25036, n25037, n25038, n25040, n25041,
         n25042, n25043, n25044, n25045, n25046, n25048, n25049, n25050,
         n25051, n25052, n25053, n25054, n25055, n25057, n25058, n25059,
         n25060, n25062, n25063, n25064, n25065, n25066, n25067, n25068,
         n25069, n25070, n25071, n25072, n25074, n25076, n25078, n25079,
         n25081, n25082, n25083, n25084, n25086, n25087, n25088, n25089,
         n25090, n25091, n25093, n25094, n25095, n25097, n25098, n25100,
         n25102, n25104, n25105, n25106, n25107, n25108, n25109, n25110,
         n25111, n25112, n25113, n25114, n25115, n25116, n25117, n25118,
         n25119, n25120, n25121, n25123, n25124, n25125, n25126, n25127,
         n25128, n25129, n25130, n25131, n25132, n25133, n25134, n25135,
         n25136, n25138, n25140, n25141, n25142, n25143, n25144, n25145,
         n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153,
         n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161,
         n25162, n25163, n25165, n25166, n25167, n25168, n25169, n25170,
         n25171, n25172, n25173, n25174, n25175, n25176, n25177, n25179,
         n25180, n25181, n25182, n25183, n25184, n25185, n25186, n25187,
         n25188, n25189, n25190, n25191, n25192, n25193, n25194, n25195,
         n25196, n25197, n25198, n25199, n25200, n25201, n25202, n25203,
         n25204, n25205, n25206, n25207, n25208, n25210, n25211, n25213,
         n25214, n25215, n25216, n25217, n25218, n25219, n25220, n25221,
         n25222, n25223, n25224, n25225, n25227, n25228, n25229, n25231,
         n25232, n25233, n25234, n25235, n25236, n25237, n25238, n25239,
         n25242, n25243, n25245, n25246, n25247, n25248, n25249, n25250,
         n25251, n25252, n25253, n25254, n25255, n25256, n25257, n25258,
         n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266,
         n25267, n25268, n25271, n25272, n25273, n25274, n25276, n25277,
         n25278, n25279, n25280, n25281, n25282, n25284, n25285, n25286,
         n25288, n25289, n25290, n25291, n25292, n25293, n25294, n25295,
         n25296, n25297, n25299, n25302, n25303, n25306, n25308, n25309,
         n25311, n25312, n25313, n25314, n25315, n25316, n25317, n25318,
         n25319, n25320, n25322, n25323, n25324, n25325, n25326, n25328,
         n25329, n25330, n25331, n25332, n25334, n25336, n25337, n25338,
         n25339, n25340, n25341, n25342, n25343, n25344, n25345, n25346,
         n25347, n25348, n25349, n25350, n25352, n25353, n25354, n25355,
         n25356, n25357, n25358, n25360, n25361, n25362, n25364, n25365,
         n25366, n25367, n25368, n25369, n25370, n25371, n25372, n25373,
         n25375, n25376, n25377, n25378, n25379, n25380, n25382, n25383,
         n25385, n25387, n25388, n25390, n25391, n25392, n25394, n25396,
         n25397, n25398, n25399, n25400, n25401, n25402, n25403, n25404,
         n25405, n25406, n25409, n25410, n25411, n25412, n25415, n25416,
         n25417, n25418, n25419, n25420, n25424, n25425, n25427, n25428,
         n25429, n25430, n25432, n25433, n25434, n25436, n25437, n25439,
         n25440, n25441, n25442, n25443, n25444, n25445, n25446, n25447,
         n25449, n25450, n25452, n25453, n25454, n25455, n25456, n25457,
         n25458, n25459, n25460, n25462, n25463, n25464, n25465, n25466,
         n25467, n25468, n25470, n25471, n25472, n25473, n25474, n25475,
         n25476, n25477, n25478, n25479, n25480, n25481, n25482, n25485,
         n25486, n25487, n25488, n25490, n25492, n25493, n25494, n25495,
         n25496, n25497, n25498, n25499, n25500, n25501, n25504, n25506,
         n25507, n25509, n25510, n25511, n25513, n25514, n25515, n25516,
         n25517, n25518, n25519, n25520, n25521, n25522, n25523, n25526,
         n25527, n25529, n25530, n25531, n25534, n25535, n25536, n25537,
         n25539, n25541, n25542, n25543, n25544, n25545, n25546, n25547,
         n25548, n25549, n25550, n25552, n25554, n25555, n25556, n25557,
         n25559, n25560, n25561, n25562, n25563, n25564, n25565, n25566,
         n25567, n25568, n25569, n25570, n25571, n25572, n25573, n25575,
         n25577, n25578, n25579, n25580, n25581, n25582, n25583, n25584,
         n25585, n25586, n25587, n25588, n25589, n25590, n25591, n25592,
         n25593, n25594, n25598, n25600, n25602, n25604, n25605, n25606,
         n25607, n25608, n25609, n25610, n25611, n25612, n25613, n25615,
         n25617, n25618, n25619, n25620, n25621, n25624, n25627, n25628,
         n25630, n25632, n25633, n25634, n25636, n25637, n25638, n25639,
         n25640, n25641, n25642, n25643, n25644, n25645, n25646, n25648,
         n25650, n25651, n25653, n25654, n25657, n25658, n25659, n25660,
         n25664, n25665, n25666, n25667, n25668, n25669, n25670, n25671,
         n25672, n25673, n25675, n25676, n25677, n25678, n25679, n25680,
         n25681, n25682, n25683, n25684, n25685, n25686, n25687, n25689,
         n25691, n25692, n25693, n25694, n25695, n25696, n25697, n25699,
         n25700, n25701, n25702, n25703, n25704, n25705, n25706, n25707,
         n25708, n25709, n25710, n25711, n25712, n25713, n25714, n25715,
         n25716, n25717, n25718, n25719, n25720, n25721, n25722, n25723,
         n25724, n25725, n25726, n25727, n25728, n25729, n25730, n25731,
         n25732, n25733, n25734, n25735, n25736, n25737, n25738, n25739,
         n25740, n25741, n25742, n25743, n25744, n25745, n25746, n25747,
         n25748, n25749, n25750, n25751, n25752, n25753, n25755, n25756,
         n25757, n25760, n25761, n25762, n25763, n25764, n25765, n25766,
         n25767, n25768, n25769, n25770, n25772, n25773, n25774, n25775,
         n25776, n25777, n25778, n25779, n25780, n25781, n25782, n25783,
         n25784, n25785, n25786, n25787, n25788, n25789, n25790, n25791,
         n25792, n25793, n25795, n25796, n25797, n25798, n25799, n25800,
         n25801, n25802, n25803, n25804, n25805, n25806, n25807, n25808,
         n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817,
         n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825,
         n25826, n25827, n25828, n25829, n25830, n25832, n25833, n25834,
         n25835, n25836, n25837, n25838, n25839, n25840, n25841, n25843,
         n25844, n25845, n25846, n25847, n25848, n25849, n25851, n25852,
         n25853, n25854, n25855, n25856, n25857, n25858, n25859, n25860,
         n25861, n25863, n25864, n25865, n25866, n25867, n25868, n25870,
         n25871, n25872, n25874, n25875, n25876, n25877, n25878, n25879,
         n25880, n25881, n25882, n25883, n25884, n25885, n25886, n25887,
         n25889, n25890, n25891, n25892, n25893, n25894, n25896, n25897,
         n25899, n25900, n25901, n25902, n25903, n25904, n25905, n25906,
         n25907, n25908, n25909, n25910, n25911, n25912, n25913, n25914,
         n25915, n25916, n25917, n25918, n25919, n25920, n25922, n25923,
         n25924, n25925, n25926, n25927, n25929, n25941, n25942, n25943,
         n25944, n25945, n25947, n25951, n25954, n25959, n25960, n25961,
         n25962, n25963, n25966, n25967, n25968, n25969, n25971, n25973,
         n25974, n25975, n25977, n25979, n25980, n25981, n25985, n25987,
         n25988, n25990, n25991, n25993, n25994, n25995, n25996, n25997,
         n25998, n25999, n26000, n26001, n26002, n26003, n26004, n26005,
         n26006, n26007, n26008, n26012, n26013, n26014, n26015, n26016,
         n26018, n26020, n26021, n26022, n26023, n26025, n26026, n26027,
         n26028, n26029, n26030, n26031, n26032, n26033, n26035, n26036,
         n26037, n26038, n26040, n26041, n26043, n26045, n26046, n26047,
         n26049, n26051, n26053, n26054, n26055, n26056, n26057, n26058,
         n26059, n26060, n26061, n26065, n26067, n26068, n26069, n26070,
         n26072, n26073, n26074, n26075, n26076, n26078, n26079, n26081,
         n26082, n26083, n26084, n26085, n26087, n26088, n26089, n26093,
         n26094, n26096, n26097, n26098, n26100, n26101, n26102, n26103,
         n26104, n26106, n26108, n26109, n26111, n26113, n26114, n26115,
         n26116, n26118, n26120, n26121, n26123, n26124, n26125, n26126,
         n26127, n26130, n26133, n26140, n26142, n26144, n26145, n26150,
         n26152, n26153, n26154, n26155, n26156, n26157, n26158, n26160,
         n26161, n26162, n26163, n26164, n26165, n26166, n26167, n26168,
         n26169, n26170, n26172, n26173, n26175, n26176, n26178, n26181,
         n26182, n26185, n26193, n26194, n26195, n26197, n26198, n26199,
         n26202, n26203, n26204, n26206, n26207, n26208, n26211, n26212,
         n26214, n26215, n26216, n26217, n26220, n26221, n26222, n26224,
         n26228, n26230, n26231, n26232, n26233, n26236, n26237, n26238,
         n26239, n26241, n26242, n26243, n26244, n26247, n26249, n26250,
         n26251, n26253, n26255, n26256, n26257, n26261, n26262, n26265,
         n26268, n26270, n26272, n26274, n26275, n26276, n26277, n26278,
         n26279, n26281, n26282, n26283, n26284, n26288, n26289, n26290,
         n26291, n26292, n26293, n26294, n26295, n26296, n26298, n26300,
         n26301, n26302, n26304, n26305, n26307, n26311, n26312, n26314,
         n26317, n26318, n26320, n26322, n26324, n26325, n26326, n26328,
         n26330, n26333, n26334, n26336, n26337, n26338, n26340, n26341,
         n26343, n26345, n26347, n26350, n26351, n26355, n26357, n26358,
         n26362, n26363, n26365, n26367, n26368, n26369, n26370, n26371,
         n26373, n26374, n26375, n26376, n26378, n26380, n26383, n26384,
         n26385, n26386, n26387, n26388, n26389, n26390, n26391, n26392,
         n26393, n26394, n26397, n26398, n26399, n26400, n26401, n26404,
         n26406, n26407, n26408, n26409, n26410, n26411, n26412, n26413,
         n26415, n26416, n26417, n26418, n26422, n26423, n26424, n26426,
         n26429, n26431, n26432, n26433, n26435, n26436, n26438, n26439,
         n26440, n26442, n26443, n26444, n26445, n26447, n26448, n26451,
         n26452, n26453, n26455, n26456, n26458, n26459, n26462, n26464,
         n26465, n26466, n26468, n26469, n26471, n26472, n26474, n26478,
         n26479, n26484, n26485, n26487, n26488, n26490, n26492, n26493,
         n26494, n26497, n26499, n26501, n26502, n26503, n26504, n26505,
         n26506, n26507, n26511, n26513, n26515, n26516, n26518, n26520,
         n26521, n26522, n26524, n26525, n26526, n26527, n26528, n26529,
         n26530, n26533, n26534, n26537, n26540, n26542, n26543, n26544,
         n26545, n26547, n26550, n26551, n26552, n26553, n26554, n26555,
         n26556, n26557, n26562, n26563, n26566, n26567, n26568, n26569,
         n26570, n26571, n26572, n26573, n26575, n26576, n26579, n26580,
         n26581, n26582, n26583, n26585, n26587, n26588, n26589, n26590,
         n26591, n26593, n26594, n26595, n26597, n26600, n26603, n26606,
         n26607, n26608, n26609, n26611, n26612, n26614, n26615, n26617,
         n26622, n26623, n26625, n26627, n26628, n26630, n26631, n26632,
         n26633, n26635, n26637, n26640, n26641, n26642, n26643, n26644,
         n26646, n26647, n26648, n26655, n26656, n26660, n26663, n26665,
         n26666, n26667, n26671, n26674, n26677, n26679, n26680, n26682,
         n26683, n26688, n26690, n26691, n26692, n26693, n26696, n26699,
         n26701, n26702, n26705, n26708, n26709, n26710, n26711, n26712,
         n26713, n26715, n26716, n26717, n26720, n26722, n26724, n26725,
         n26726, n26727, n26728, n26730, n26731, n26732, n26733, n26735,
         n26736, n26738, n26739, n26740, n26741, n26742, n26744, n26745,
         n26747, n26750, n26751, n26753, n26754, n26755, n26756, n26758,
         n26761, n26762, n26765, n26766, n26767, n26768, n26769, n26772,
         n26774, n26775, n26777, n26778, n26780, n26782, n26784, n26785,
         n26787, n26790, n26791, n26793, n26794, n26795, n26796, n26798,
         n26799, n26800, n26801, n26803, n26806, n26807, n26808, n26810,
         n26812, n26813, n26814, n26815, n26817, n26818, n26821, n26822,
         n26823, n26825, n26827, n26829, n26830, n26834, n26835, n26836,
         n26837, n26842, n26844, n26845, n26846, n26848, n26851, n26854,
         n26855, n26856, n26858, n26861, n26862, n26863, n26865, n26867,
         n26868, n26869, n26872, n26873, n26874, n26875, n26877, n26878,
         n26881, n26882, n26883, n26884, n26885, n26886, n26887, n26888,
         n26889, n26890, n26891, n26892, n26896, n26897, n26898, n26899,
         n26900, n26903, n26904, n26907, n26909, n26912, n26913, n26914,
         n26915, n26916, n26917, n26918, n26920, n26921, n26922, n26923,
         n26924, n26925, n26927, n26929, n26930, n26931, n26933, n26934,
         n26936, n26937, n26938, n26941, n26942, n26945, n26947, n26948,
         n26949, n26950, n26953, n26954, n26955, n26956, n26957, n26958,
         n26960, n26961, n26962, n26965, n26966, n26967, n26969, n26971,
         n26974, n26976, n26977, n26978, n26979, n26980, n26983, n26986,
         n26987, n26988, n26990, n26991, n26992, n26993, n26994, n26995,
         n26996, n26997, n26998, n27000, n27004, n27005, n27007, n27008,
         n27010, n27011, n27012, n27014, n27015, n27016, n27018, n27019,
         n27020, n27021, n27023, n27024, n27026, n27028, n27033, n27034,
         n27038, n27041, n27042, n27044, n27046, n27047, n27049, n27050,
         n27052, n27053, n27054, n27055, n27057, n27058, n27060, n27062,
         n27063, n27064, n27065, n27066, n27067, n27070, n27072, n27073,
         n27075, n27076, n27077, n27078, n27079, n27080, n27081, n27082,
         n27088, n27090, n27091, n27092, n27094, n27097, n27098, n27099,
         n27100, n27101, n27103, n27104, n27105, n27106, n27110, n27111,
         n27113, n27114, n27115, n27117, n27118, n27119, n27120, n27121,
         n27122, n27123, n27125, n27126, n27127, n27128, n27129, n27130,
         n27131, n27132, n27134, n27135, n27136, n27137, n27138, n27139,
         n27142, n27143, n27144, n27145, n27146, n27147, n27148, n27149,
         n27150, n27151, n27152, n27153, n27154, n27155, n27156, n27157,
         n27159, n27160, n27162, n27163, n27164, n27165, n27166, n27167,
         n27168, n27169, n27170, n27171, n27173, n27174, n27175, n27176,
         n27177, n27178, n27179, n27180, n27181, n27182, n27183, n27184,
         n27185, n27186, n27188, n27189, n27190, n27191, n27192, n27193,
         n27196, n27198, n27200, n27201, n27202, n27203, n27207, n27208,
         n27211, n27212, n27214, n27215, n27217, n27218, n27219, n27220,
         n27225, n27226, n27227, n27228, n27230, n27232, n27233, n27234,
         n27236, n27237, n27238, n27240, n27242, n27243, n27244, n27245,
         n27246, n27248, n27249, n27252, n27253, n27257, n27259, n27261,
         n27262, n27263, n27265, n27266, n27267, n27268, n27269, n27270,
         n27271, n27272, n27273, n27274, n27275, n27276, n27277, n27279,
         n27281, n27282, n27283, n27284, n27285, n27289, n27290, n27294,
         n27296, n27297, n27298, n27299, n27300, n27301, n27302, n27303,
         n27305, n27307, n27308, n27309, n27311, n27312, n27314, n27315,
         n27316, n27317, n27318, n27320, n27321, n27324, n27326, n27329,
         n27330, n27332, n27334, n27336, n27337, n27338, n27340, n27341,
         n27342, n27343, n27344, n27345, n27349, n27352, n27353, n27354,
         n27357, n27358, n27359, n27360, n27361, n27362, n27363, n27365,
         n27367, n27368, n27369, n27372, n27373, n27374, n27375, n27376,
         n27377, n27378, n27379, n27381, n27382, n27383, n27384, n27385,
         n27386, n27387, n27388, n27389, n27390, n27391, n27392, n27395,
         n27396, n27397, n27398, n27401, n27402, n27403, n27406, n27408,
         n27409, n27410, n27411, n27412, n27413, n27415, n27416, n27419,
         n27420, n27423, n27424, n27426, n27428, n27429, n27430, n27431,
         n27432, n27435, n27436, n27437, n27439, n27440, n27441, n27442,
         n27443, n27444, n27445, n27446, n27450, n27451, n27453, n27454,
         n27455, n27456, n27457, n27458, n27459, n27460, n27461, n27462,
         n27466, n27471, n27472, n27474, n27475, n27478, n27479, n27480,
         n27481, n27482, n27485, n27486, n27487, n27490, n27491, n27495,
         n27500, n27501, n27503, n27504, n27505, n27506, n27509, n27514,
         n27515, n27516, n27517, n27518, n27520, n27523, n27525, n27526,
         n27528, n27529, n27531, n27532, n27534, n27535, n27537, n27538,
         n27539, n27541, n27542, n27543, n27544, n27545, n27548, n27550,
         n27551, n27552, n27553, n27555, n27556, n27560, n27561, n27563,
         n27565, n27566, n27567, n27569, n27570, n27571, n27573, n27574,
         n27575, n27577, n27580, n27582, n27583, n27585, n27586, n27587,
         n27588, n27589, n27590, n27591, n27592, n27593, n27594, n27595,
         n27596, n27597, n27599, n27600, n27601, n27604, n27605, n27607,
         n27608, n27609, n27610, n27611, n27612, n27613, n27615, n27616,
         n27617, n27618, n27619, n27620, n27621, n27622, n27624, n27625,
         n27627, n27628, n27629, n27630, n27631, n27633, n27635, n27637,
         n27638, n27639, n27641, n27642, n27643, n27645, n27646, n27648,
         n27649, n27650, n27651, n27652, n27654, n27655, n27658, n27659,
         n27660, n27661, n27662, n27664, n27667, n27668, n27669, n27670,
         n27672, n27673, n27676, n27678, n27679, n27680, n27683, n27684,
         n27685, n27686, n27687, n27688, n27689, n27690, n27691, n27693,
         n27694, n27695, n27696, n27697, n27698, n27699, n27701, n27703,
         n27704, n27706, n27707, n27708, n27709, n27711, n27714, n27715,
         n27716, n27717, n27718, n27719, n27720, n27721, n27724, n27726,
         n27728, n27729, n27731, n27732, n27733, n27734, n27735, n27736,
         n27737, n27738, n27739, n27741, n27743, n27745, n27747, n27748,
         n27750, n27752, n27753, n27754, n27755, n27756, n27757, n27758,
         n27759, n27760, n27761, n27762, n27763, n27764, n27765, n27766,
         n27767, n27768, n27769, n27771, n27773, n27775, n27776, n27778,
         n27779, n27781, n27785, n27786, n27787, n27788, n27790, n27791,
         n27792, n27793, n27797, n27798, n27799, n27801, n27802, n27804,
         n27805, n27806, n27807, n27808, n27811, n27812, n27814, n27816,
         n27818, n27819, n27823, n27824, n27825, n27826, n27828, n27829,
         n27830, n27831, n27832, n27833, n27834, n27835, n27836, n27837,
         n27838, n27840, n27841, n27842, n27845, n27846, n27850, n27851,
         n27852, n27854, n27856, n27857, n27860, n27861, n27862, n27863,
         n27864, n27865, n27866, n27867, n27868, n27872, n27873, n27875,
         n27876, n27877, n27878, n27879, n27880, n27881, n27882, n27883,
         n27884, n27886, n27887, n27889, n27893, n27894, n27895, n27896,
         n27897, n27899, n27900, n27901, n27902, n27904, n27907, n27908,
         n27909, n27910, n27911, n27912, n27914, n27916, n27919, n27920,
         n27921, n27922, n27923, n27925, n27926, n27929, n27930, n27931,
         n27933, n27934, n27936, n27937, n27938, n27939, n27940, n27941,
         n27942, n27943, n27946, n27947, n27950, n27951, n27952, n27953,
         n27954, n27955, n27957, n27958, n27959, n27960, n27961, n27962,
         n27963, n27965, n27968, n27969, n27970, n27971, n27972, n27973,
         n27975, n27976, n27977, n27980, n27981, n27982, n27984, n27987,
         n27988, n27990, n27991, n27992, n27993, n27994, n27995, n27996,
         n27998, n28000, n28001, n28002, n28003, n28004, n28005, n28009,
         n28010, n28011, n28012, n28014, n28016, n28017, n28018, n28019,
         n28020, n28021, n28022, n28025, n28027, n28028, n28029, n28030,
         n28031, n28034, n28035, n28037, n28038, n28039, n28040, n28043,
         n28052, n28056, n28057, n28058, n28059, n28061, n28062, n28064,
         n28067, n28068, n28069, n28070, n28071, n28072, n28073, n28074,
         n28077, n28078, n28081, n28082, n28083, n28084, n28085, n28086,
         n28087, n28091, n28093, n28096, n28097, n28098, n28099, n28100,
         n28101, n28102, n28104, n28105, n28107, n28108, n28109, n28110,
         n28111, n28113, n28114, n28116, n28117, n28118, n28119, n28120,
         n28121, n28123, n28124, n28126, n28128, n28130, n28131, n28132,
         n28133, n28134, n28135, n28136, n28137, n28138, n28139, n28141,
         n28142, n28144, n28147, n28150, n28151, n28152, n28153, n28154,
         n28155, n28156, n28157, n28158, n28159, n28160, n28162, n28163,
         n28166, n28167, n28170, n28171, n28172, n28174, n28175, n28177,
         n28178, n28179, n28181, n28183, n28186, n28188, n28190, n28194,
         n28196, n28197, n28199, n28200, n28202, n28203, n28205, n28206,
         n28208, n28209, n28210, n28211, n28214, n28216, n28217, n28218,
         n28219, n28220, n28222, n28223, n28225, n28226, n28227, n28228,
         n28231, n28232, n28234, n28235, n28236, n28237, n28238, n28239,
         n28240, n28242, n28243, n28244, n28245, n28246, n28251, n28252,
         n28253, n28254, n28255, n28256, n28257, n28258, n28260, n28261,
         n28262, n28263, n28265, n28266, n28268, n28269, n28270, n28273,
         n28275, n28276, n28277, n28278, n28279, n28281, n28283, n28285,
         n28286, n28287, n28288, n28289, n28293, n28295, n28296, n28297,
         n28298, n28299, n28300, n28302, n28303, n28304, n28306, n28307,
         n28308, n28309, n28311, n28312, n28313, n28314, n28315, n28316,
         n28318, n28320, n28321, n28323, n28324, n28327, n28328, n28329,
         n28330, n28331, n28332, n28338, n28340, n28342, n28343, n28344,
         n28345, n28347, n28348, n28349, n28350, n28351, n28353, n28354,
         n28355, n28356, n28357, n28358, n28361, n28364, n28365, n28366,
         n28367, n28371, n28372, n28373, n28374, n28375, n28376, n28378,
         n28379, n28380, n28381, n28382, n28383, n28385, n28386, n28387,
         n28388, n28390, n28391, n28393, n28395, n28396, n28397, n28399,
         n28400, n28401, n28402, n28403, n28404, n28405, n28406, n28407,
         n28408, n28409, n28410, n28411, n28413, n28414, n28415, n28416,
         n28418, n28419, n28420, n28421, n28422, n28423, n28424, n28425,
         n28426, n28427, n28428, n28429, n28430, n28431, n28432, n28435,
         n28436, n28437, n28438, n28439, n28441, n28442, n28443, n28444,
         n28446, n28447, n28448, n28449, n28450, n28451, n28452, n28453,
         n28454, n28455, n28456, n28457, n28458, n28459, n28460, n28461,
         n28462, n28463, n28465, n28466, n28467, n28469, n28470, n28471,
         n28472, n28473, n28474, n28475, n28478, n28479, n28480, n28482,
         n28483, n28484, n28485, n28486, n28487, n28488, n28489, n28490,
         n28491, n28492, n28493, n28494, n28495, n28496, n28497, n28498,
         n28501, n28502, n28503, n28504, n28505, n28506, n28507, n28509,
         n28510, n28513, n28514, n28516, n28517, n28519, n28520, n28522,
         n28523, n28524, n28525, n28526, n28527, n28528, n28530, n28531,
         n28532, n28534, n28536, n28538, n28539, n28540, n28541, n28542,
         n28543, n28544, n28545, n28548, n28549, n28552, n28553, n28554,
         n28555, n28557, n28560, n28562, n28564, n28565, n28566, n28567,
         n28568, n28571, n28573, n28574, n28575, n28578, n28579, n28580,
         n28581, n28584, n28585, n28586, n28587, n28589, n28590, n28591,
         n28592, n28593, n28594, n28595, n28600, n28601, n28602, n28603,
         n28605, n28606, n28607, n28608, n28611, n28612, n28613, n28614,
         n28615, n28616, n28617, n28618, n28621, n28622, n28623, n28624,
         n28625, n28626, n28627, n28631, n28632, n28633, n28634, n28635,
         n28636, n28637, n28638, n28639, n28640, n28641, n28642, n28644,
         n28645, n28647, n28648, n28649, n28651, n28652, n28654, n28655,
         n28657, n28658, n28659, n28660, n28661, n28662, n28663, n28664,
         n28665, n28668, n28669, n28670, n28671, n28672, n28673, n28674,
         n28675, n28676, n28680, n28681, n28683, n28684, n28685, n28686,
         n28687, n28688, n28689, n28691, n28692, n28694, n28696, n28697,
         n28698, n28699, n28700, n28701, n28702, n28703, n28704, n28705,
         n28706, n28707, n28708, n28709, n28710, n28711, n28712, n28714,
         n28715, n28721, n28722, n28723, n28724, n28725, n28726, n28728,
         n28729, n28730, n28731, n28733, n28734, n28735, n28736, n28737,
         n28738, n28740, n28743, n28744, n28745, n28746, n28747, n28748,
         n28750, n28751, n28752, n28753, n28754, n28755, n28757, n28758,
         n28759, n28760, n28761, n28762, n28763, n28765, n28767, n28769,
         n28770, n28771, n28773, n28775, n28776, n28777, n28778, n28779,
         n28781, n28782, n28783, n28784, n28786, n28788, n28789, n28791,
         n28796, n28797, n28799, n28800, n28801, n28802, n28803, n28806,
         n28807, n28811, n28812, n28813, n28814, n28815, n28816, n28817,
         n28818, n28819, n28821, n28822, n28823, n28824, n28825, n28826,
         n28827, n28829, n28830, n28831, n28833, n28835, n28836, n28837,
         n28838, n28839, n28840, n28844, n28846, n28847, n28848, n28849,
         n28850, n28852, n28853, n28854, n28855, n28856, n28857, n28859,
         n28860, n28861, n28862, n28863, n28864, n28865, n28866, n28867,
         n28868, n28869, n28870, n28872, n28873, n28875, n28876, n28877,
         n28878, n28880, n28882, n28883, n28885, n28886, n28887, n28888,
         n28889, n28891, n28893, n28894, n28895, n28896, n28897, n28898,
         n28899, n28900, n28902, n28903, n28904, n28908, n28909, n28910,
         n28911, n28912, n28913, n28914, n28915, n28916, n28917, n28918,
         n28921, n28922, n28923, n28924, n28926, n28927, n28929, n28931,
         n28932, n28933, n28934, n28935, n28937, n28938, n28939, n28940,
         n28941, n28942, n28943, n28944, n28945, n28946, n28947, n28948,
         n28949, n28950, n28951, n28952, n28953, n28954, n28956, n28957,
         n28958, n28964, n28967, n28968, n28970, n28972, n28973, n28974,
         n28975, n28977, n28978, n28979, n28981, n28982, n28983, n28987,
         n28989, n28990, n28992, n28993, n28995, n28996, n28998, n28999,
         n29000, n29001, n29002, n29003, n29004, n29007, n29008, n29009,
         n29010, n29011, n29012, n29013, n29018, n29020, n29021, n29022,
         n29026, n29027, n29028, n29029, n29030, n29032, n29033, n29034,
         n29035, n29037, n29039, n29040, n29042, n29043, n29044, n29046,
         n29047, n29048, n29049, n29050, n29051, n29052, n29054, n29056,
         n29057, n29060, n29061, n29062, n29063, n29064, n29068, n29069,
         n29070, n29071, n29072, n29073, n29074, n29075, n29076, n29077,
         n29078, n29079, n29080, n29081, n29082, n29084, n29085, n29087,
         n29088, n29089, n29090, n29093, n29094, n29095, n29098, n29099,
         n29101, n29102, n29106, n29107, n29108, n29110, n29111, n29114,
         n29115, n29116, n29118, n29119, n29120, n29121, n29122, n29123,
         n29124, n29127, n29130, n29131, n29133, n29134, n29135, n29137,
         n29138, n29139, n29140, n29141, n29142, n29143, n29146, n29147,
         n29148, n29149, n29152, n29153, n29155, n29156, n29157, n29158,
         n29159, n29160, n29162, n29167, n29168, n29169, n29170, n29172,
         n29173, n29174, n29175, n29176, n29178, n29180, n29182, n29184,
         n29185, n29187, n29189, n29190, n29194, n29196, n29198, n29200,
         n29201, n29202, n29203, n29205, n29206, n29207, n29208, n29209,
         n29211, n29212, n29213, n29214, n29215, n29216, n29217, n29218,
         n29220, n29221, n29222, n29223, n29224, n29225, n29227, n29228,
         n29230, n29231, n29232, n29233, n29234, n29235, n29236, n29239,
         n29240, n29241, n29242, n29243, n29244, n29245, n29246, n29250,
         n29252, n29253, n29254, n29255, n29256, n29258, n29259, n29260,
         n29261, n29262, n29263, n29266, n29268, n29269, n29270, n29271,
         n29272, n29273, n29274, n29275, n29277, n29278, n29279, n29280,
         n29281, n29282, n29283, n29284, n29285, n29286, n29287, n29288,
         n29291, n29292, n29293, n29294, n29296, n29299, n29302, n29303,
         n29304, n29305, n29306, n29307, n29308, n29309, n29312, n29313,
         n29314, n29315, n29317, n29318, n29320, n29321, n29322, n29323,
         n29325, n29328, n29329, n29330, n29331, n29334, n29335, n29336,
         n29337, n29338, n29339, n29341, n29342, n29343, n29344, n29345,
         n29346, n29347, n29348, n29349, n29350, n29351, n29352, n29353,
         n29354, n29355, n29356, n29357, n29358, n29359, n29360, n29361,
         n29362, n29363, n29364, n29365, n29366, n29367, n29368, n29369,
         n29370, n29371, n29372, n29373, n29375, n29376, n29378, n29379,
         n29380, n29382, n29383, n29384, n29385, n29386, n29387, n29388,
         n29389, n29390, n29391, n29392, n29393, n29394, n29395, n29396,
         n29397, n29398, n29400, n29401, n29402, n29404, n29405, n29406,
         n29407, n29408, n29409, n29412, n29413, n29415, n29416, n29417,
         n29418, n29420, n29421, n29422, n29423, n29424, n29426, n29427,
         n29428, n29430, n29431, n29432, n29433, n29434, n29435, n29437,
         n29438, n29440, n29441, n29442, n29443, n29444, n29445, n29446,
         n29447, n29448, n29450, n29451, n29453, n29454, n29455, n29457,
         n29458, n29460, n29461, n29462, n29463, n29464, n29467, n29469,
         n29470, n29471, n29472, n29473, n29474, n29475, n29476, n29477,
         n29480, n29481, n29482, n29483, n29485, n29486, n29487, n29488,
         n29489, n29492, n29494, n29495, n29497, n29498, n29499, n29501,
         n29502, n29503, n29507, n29508, n29509, n29510, n29512, n29514,
         n29515, n29517, n29518, n29520, n29521, n29522, n29523, n29525,
         n29526, n29527, n29528, n29531, n29532, n29534, n29536, n29537,
         n29538, n29539, n29540, n29541, n29543, n29545, n29547, n29548,
         n29550, n29551, n29552, n29553, n29554, n29555, n29557, n29559,
         n29560, n29561, n29562, n29563, n29566, n29567, n29568, n29570,
         n29572, n29573, n29574, n29575, n29576, n29577, n29578, n29580,
         n29581, n29582, n29583, n29584, n29586, n29588, n29589, n29590,
         n29593, n29594, n29595, n29597, n29598, n29600, n29602, n29603,
         n29605, n29606, n29607, n29608, n29609, n29610, n29614, n29615,
         n29618, n29620, n29621, n29623, n29624, n29626, n29628, n29629,
         n29630, n29631, n29632, n29633, n29634, n29635, n29636, n29638,
         n29639, n29642, n29643, n29644, n29645, n29646, n29648, n29650,
         n29651, n29652, n29653, n29654, n29655, n29656, n29657, n29658,
         n29659, n29660, n29661, n29662, n29663, n29664, n29666, n29667,
         n29668, n29670, n29671, n29672, n29673, n29674, n29675, n29676,
         n29678, n29679, n29680, n29681, n29682, n29683, n29684, n29687,
         n29688, n29689, n29690, n29692, n29693, n29695, n29696, n29699,
         n29702, n29704, n29705, n29706, n29707, n29708, n29709, n29711,
         n29712, n29714, n29715, n29717, n29718, n29719, n29720, n29721,
         n29722, n29723, n29724, n29725, n29726, n29727, n29728, n29729,
         n29730, n29731, n29732, n29733, n29734, n29736, n29737, n29738,
         n29739, n29740, n29741, n29742, n29743, n29748, n29750, n29751,
         n29753, n29754, n29755, n29757, n29758, n29759, n29761, n29762,
         n29763, n29765, n29767, n29768, n29769, n29771, n29772, n29773,
         n29774, n29776, n29777, n29778, n29780, n29781, n29784, n29785,
         n29787, n29788, n29789, n29790, n29791, n29792, n29795, n29796,
         n29799, n29800, n29801, n29802, n29803, n29804, n29806, n29807,
         n29808, n29809, n29810, n29811, n29812, n29813, n29814, n29815,
         n29817, n29818, n29819, n29820, n29821, n29823, n29825, n29827,
         n29828, n29829, n29830, n29832, n29833, n29834, n29835, n29836,
         n29837, n29838, n29839, n29840, n29841, n29843, n29844, n29845,
         n29846, n29847, n29848, n29849, n29850, n29851, n29853, n29854,
         n29855, n29856, n29858, n29863, n29864, n29865, n29866, n29867,
         n29868, n29870, n29872, n29873, n29875, n29876, n29877, n29878,
         n29879, n29880, n29882, n29883, n29885, n29888, n29890, n29895,
         n29896, n29898, n29899, n29900, n29901, n29903, n29904, n29905,
         n29906, n29907, n29908, n29909, n29911, n29912, n29913, n29914,
         n29915, n29916, n29918, n29919, n29920, n29921, n29922, n29924,
         n29927, n29928, n29930, n29931, n29932, n29933, n29934, n29936,
         n29937, n29938, n29943, n29944, n29946, n29947, n29949, n29951,
         n29952, n29953, n29954, n29955, n29957, n29958, n29960, n29962,
         n29963, n29964, n29965, n29967, n29969, n29970, n29972, n29973,
         n29975, n29976, n29977, n29978, n29980, n29981, n29982, n29983,
         n29985, n29986, n29987, n29988, n29989, n29993, n29994, n29995,
         n29997, n30000, n30001, n30003, n30004, n30005, n30006, n30007,
         n30008, n30010, n30011, n30012, n30013, n30014, n30015, n30016,
         n30017, n30018, n30019, n30020, n30021, n30022, n30025, n30028,
         n30029, n30031, n30032, n30033, n30036, n30038, n30039, n30041,
         n30042, n30044, n30045, n30047, n30048, n30049, n30050, n30054,
         n30057, n30058, n30059, n30060, n30061, n30062, n30063, n30064,
         n30065, n30066, n30067, n30069, n30070, n30071, n30072, n30074,
         n30075, n30076, n30078, n30079, n30080, n30081, n30082, n30083,
         n30084, n30085, n30086, n30087, n30088, n30089, n30090, n30091,
         n30093, n30094, n30096, n30097, n30098, n30099, n30102, n30104,
         n30105, n30106, n30107, n30109, n30110, n30111, n30112, n30114,
         n30115, n30116, n30117, n30118, n30119, n30121, n30122, n30123,
         n30124, n30125, n30126, n30127, n30129, n30130, n30131, n30134,
         n30135, n30136, n30137, n30138, n30139, n30140, n30142, n30143,
         n30144, n30145, n30146, n30148, n30149, n30151, n30152, n30154,
         n30155, n30156, n30157, n30159, n30163, n30165, n30167, n30168,
         n30169, n30171, n30172, n30173, n30174, n30175, n30176, n30177,
         n30180, n30181, n30182, n30183, n30185, n30186, n30187, n30188,
         n30189, n30190, n30191, n30192, n30193, n30195, n30197, n30198,
         n30199, n30200, n30202, n30203, n30204, n30205, n30207, n30209,
         n30212, n30214, n30215, n30216, n30218, n30219, n30220, n30221,
         n30222, n30223, n30224, n30225, n30226, n30227, n30229, n30230,
         n30231, n30232, n30233, n30234, n30235, n30236, n30237, n30240,
         n30241, n30243, n30246, n30247, n30248, n30250, n30251, n30252,
         n30255, n30257, n30258, n30259, n30262, n30265, n30267, n30269,
         n30270, n30271, n30272, n30273, n30274, n30275, n30276, n30277,
         n30278, n30279, n30280, n30281, n30282, n30283, n30284, n30285,
         n30288, n30289, n30290, n30291, n30293, n30294, n30295, n30296,
         n30297, n30301, n30302, n30303, n30304, n30305, n30306, n30307,
         n30308, n30309, n30311, n30313, n30314, n30315, n30316, n30317,
         n30318, n30319, n30320, n30321, n30322, n30323, n30326, n30327,
         n30328, n30329, n30330, n30331, n30332, n30333, n30334, n30336,
         n30338, n30339, n30340, n30341, n30342, n30344, n30345, n30346,
         n30348, n30349, n30353, n30354, n30355, n30356, n30357, n30358,
         n30359, n30360, n30362, n30364, n30365, n30366, n30367, n30368,
         n30369, n30370, n30371, n30372, n30374, n30375, n30379, n30380,
         n30381, n30382, n30383, n30384, n30385, n30386, n30387, n30388,
         n30389, n30390, n30391, n30393, n30394, n30396, n30398, n30400,
         n30401, n30402, n30403, n30404, n30405, n30407, n30408, n30409,
         n30410, n30411, n30412, n30413, n30414, n30417, n30418, n30420,
         n30421, n30423, n30425, n30426, n30427, n30428, n30429, n30430,
         n30433, n30435, n30436, n30437, n30439, n30440, n30441, n30442,
         n30443, n30444, n30445, n30446, n30447, n30448, n30449, n30450,
         n30453, n30454, n30455, n30458, n30459, n30461, n30462, n30463,
         n30464, n30465, n30466, n30467, n30469, n30470, n30471, n30472,
         n30473, n30474, n30475, n30476, n30477, n30479, n30480, n30482,
         n30483, n30486, n30487, n30488, n30489, n30492, n30493, n30494,
         n30495, n30496, n30497, n30498, n30501, n30502, n30503, n30504,
         n30505, n30506, n30507, n30508, n30509, n30510, n30511, n30512,
         n30513, n30514, n30515, n30517, n30521, n30522, n30523, n30524,
         n30526, n30527, n30528, n30529, n30530, n30532, n30535, n30536,
         n30537, n30538, n30539, n30540, n30541, n30542, n30543, n30544,
         n30545, n30546, n30547, n30548, n30549, n30550, n30551, n30552,
         n30553, n30554, n30555, n30556, n30557, n30558, n30559, n30560,
         n30561, n30562, n30563, n30564, n30565, n30568, n30569, n30570,
         n30571, n30572, n30573, n30574, n30575, n30578, n30579, n30583,
         n30584, n30586, n30587, n30592, n30593, n30594, n30595, n30596,
         n30597, n30598, n30600, n30601, n30602, n30603, n30607, n30608,
         n30610, n30612, n30614, n30615, n30616, n30617, n30618, n30619,
         n30620, n30621, n30622, n30623, n30624, n30625, n30626, n30627,
         n30628, n30631, n30632, n30633, n30634, n30635, n30636, n30637,
         n30638, n30639, n30640, n30641, n30643, n30644, n30645, n30646,
         n30648, n30649, n30651, n30652, n30653, n30654, n30656, n30658,
         n30660, n30661, n30663, n30664, n30666, n30668, n30669, n30670,
         n30671, n30673, n30676, n30677, n30678, n30679, n30681, n30682,
         n30685, n30686, n30687, n30688, n30690, n30691, n30692, n30693,
         n30694, n30695, n30696, n30697, n30698, n30699, n30700, n30702,
         n30703, n30705, n30706, n30707, n30708, n30710, n30711, n30712,
         n30713, n30714, n30715, n30716, n30717, n30718, n30720, n30721,
         n30722, n30723, n30724, n30725, n30726, n30727, n30728, n30729,
         n30730, n30731, n30732, n30733, n30734, n30736, n30737, n30740,
         n30741, n30742, n30743, n30744, n30745, n30746, n30747, n30748,
         n30749, n30753, n30754, n30755, n30757, n30758, n30760, n30762,
         n30763, n30765, n30766, n30767, n30768, n30769, n30770, n30771,
         n30774, n30776, n30777, n30778, n30779, n30780, n30781, n30783,
         n30784, n30789, n30790, n30792, n30793, n30794, n30795, n30798,
         n30800, n30802, n30803, n30805, n30806, n30807, n30808, n30810,
         n30811, n30813, n30815, n30816, n30817, n30818, n30819, n30820,
         n30822, n30824, n30825, n30826, n30828, n30830, n30831, n30832,
         n30833, n30837, n30838, n30840, n30843, n30844, n30845, n30846,
         n30849, n30850, n30852, n30853, n30854, n30855, n30856, n30857,
         n30858, n30861, n30862, n30863, n30865, n30866, n30867, n30868,
         n30869, n30870, n30871, n30872, n30873, n30875, n30876, n30877,
         n30878, n30879, n30880, n30881, n30882, n30883, n30885, n30886,
         n30887, n30888, n30889, n30892, n30894, n30895, n30898, n30899,
         n30900, n30901, n30902, n30904, n30905, n30906, n30907, n30908,
         n30909, n30912, n30913, n30914, n30915, n30917, n30919, n30922,
         n30923, n30924, n30925, n30926, n30928, n30929, n30930, n30931,
         n30932, n30933, n30934, n30935, n30936, n30937, n30938, n30940,
         n30942, n30943, n30945, n30946, n30948, n30949, n30951, n30952,
         n30953, n30954, n30955, n30957, n30958, n30959, n30960, n30961,
         n30962, n30963, n30964, n30965, n30966, n30967, n30968, n30969,
         n30970, n30971, n30972, n30973, n30976, n30978, n30979, n30980,
         n30981, n30982, n30983, n30984, n30985, n30986, n30987, n30988,
         n30989, n30990, n30991, n30992, n30993, n30994, n30995, n30996,
         n30997, n30998, n30999, n31001, n31002, n31003, n31004, n31005,
         n31006, n31007, n31009, n31012, n31015, n31016, n31017, n31019,
         n31021, n31022, n31025, n31026, n31028, n31029, n31030, n31032,
         n31033, n31034, n31036, n31037, n31039, n31040, n31041, n31042,
         n31043, n31044, n31046, n31047, n31048, n31051, n31052, n31054,
         n31055, n31056, n31057, n31058, n31059, n31060, n31062, n31063,
         n31065, n31066, n31070, n31071, n31072, n31073, n31074, n31075,
         n31077, n31078, n31079, n31080, n31081, n31082, n31083, n31084,
         n31085, n31086, n31087, n31088, n31089, n31090, n31091, n31092,
         n31093, n31094, n31095, n31096, n31097, n31098, n31099, n31100,
         n31101, n31102, n31103, n31104, n31105, n31106, n31108, n31109,
         n31110, n31111, n31112, n31113, n31114, n31115, n31116, n31117,
         n31118, n31120, n31121, n31122, n31123, n31124, n31126, n31127,
         n31128, n31129, n31132, n31133, n31135, n31136, n31137, n31138,
         n31139, n31140, n31141, n31142, n31143, n31144, n31145, n31146,
         n31147, n31148, n31149, n31150, n31151, n31152, n31155, n31156,
         n31157, n31158, n31159, n31160, n31161, n31162, n31163, n31164,
         n31165, n31167, n31168, n31169, n31170, n31171, n31173, n31174,
         n31175, n31177, n31178, n31179, n31180, n31181, n31182, n31184,
         n31185, n31186, n31188, n31189, n31190, n31191, n31194, n31195,
         n31197, n31200, n31201, n31202, n31203, n31205, n31206, n31207,
         n31208, n31209, n31210, n31211, n31213, n31214, n31215, n31216,
         n31217, n31218, n31220, n31221, n31223, n31225, n31226, n31228,
         n31229, n31231, n31232, n31233, n31234, n31235, n31236, n31237,
         n31238, n31239, n31241, n31242, n31243, n31244, n31245, n31246,
         n31247, n31248, n31250, n31251, n31252, n31253, n31254, n31258,
         n31259, n31260, n31262, n31263, n31264, n31265, n31266, n31267,
         n31268, n31269, n31271, n31272, n31273, n31274, n31275, n31277,
         n31279, n31280, n31281, n31282, n31284, n31285, n31286, n31287,
         n31288, n31290, n31291, n31292, n31293, n31294, n31295, n31296,
         n31297, n31301, n31303, n31306, n31308, n31309, n31311, n31312,
         n31314, n31315, n31316, n31317, n31318, n31319, n31320, n31321,
         n31323, n31324, n31325, n31327, n31329, n31330, n31331, n31333,
         n31334, n31335, n31336, n31338, n31339, n31340, n31341, n31342,
         n31344, n31345, n31346, n31348, n31349, n31350, n31351, n31352,
         n31354, n31355, n31356, n31357, n31358, n31359, n31360, n31361,
         n31363, n31365, n31366, n31367, n31368, n31369, n31370, n31371,
         n31372, n31373, n31374, n31377, n31378, n31379, n31380, n31381,
         n31385, n31387, n31389, n31390, n31393, n31394, n31395, n31396,
         n31397, n31398, n31399, n31400, n31401, n31402, n31403, n31404,
         n31405, n31406, n31407, n31408, n31409, n31410, n31411, n31414,
         n31415, n31416, n31417, n31418, n31419, n31421, n31422, n31423,
         n31424, n31426, n31427, n31428, n31429, n31432, n31434, n31435,
         n31437, n31438, n31440, n31442, n31443, n31444, n31445, n31448,
         n31450, n31451, n31453, n31454, n31455, n31456, n31457, n31458,
         n31459, n31461, n31463, n31464, n31467, n31468, n31469, n31470,
         n31471, n31473, n31474, n31475, n31476, n31477, n31478, n31479,
         n31483, n31484, n31485, n31486, n31487, n31488, n31489, n31490,
         n31491, n31492, n31493, n31495, n31496, n31497, n31498, n31499,
         n31500, n31503, n31504, n31505, n31506, n31507, n31508, n31509,
         n31510, n31511, n31512, n31513, n31514, n31516, n31519, n31521,
         n31522, n31523, n31524, n31525, n31526, n31527, n31528, n31529,
         n31531, n31532, n31533, n31534, n31538, n31539, n31542, n31543,
         n31544, n31545, n31547, n31548, n31549, n31551, n31552, n31553,
         n31554, n31557, n31559, n31560, n31561, n31562, n31563, n31564,
         n31566, n31567, n31568, n31569, n31570, n31571, n31572, n31573,
         n31574, n31575, n31576, n31579, n31583, n31584, n31585, n31588,
         n31590, n31591, n31593, n31594, n31596, n31597, n31598, n31599,
         n31601, n31602, n31603, n31604, n31606, n31607, n31608, n31611,
         n31612, n31613, n31614, n31615, n31616, n31617, n31618, n31619,
         n31622, n31623, n31626, n31627, n31629, n31630, n31634, n31635,
         n31636, n31637, n31638, n31639, n31640, n31642, n31643, n31644,
         n31645, n31646, n31647, n31649, n31650, n31653, n31654, n31655,
         n31656, n31657, n31658, n31660, n31661, n31662, n31663, n31664,
         n31666, n31667, n31668, n31669, n31670, n31671, n31673, n31674,
         n31675, n31676, n31677, n31678, n31679, n31682, n31683, n31684,
         n31686, n31687, n31689, n31690, n31691, n31692, n31693, n31694,
         n31695, n31696, n31697, n31698, n31699, n31701, n31702, n31703,
         n31704, n31706, n31707, n31709, n31710, n31711, n31712, n31713,
         n31714, n31715, n31716, n31718, n31719, n31720, n31721, n31722,
         n31724, n31725, n31726, n31727, n31728, n31729, n31730, n31731,
         n31732, n31734, n31736, n31737, n31738, n31739, n31742, n31745,
         n31746, n31747, n31748, n31749, n31750, n31751, n31753, n31754,
         n31755, n31756, n31757, n31758, n31759, n31760, n31761, n31762,
         n31763, n31765, n31766, n31767, n31768, n31769, n31770, n31771,
         n31772, n31773, n31776, n31777, n31778, n31779, n31780, n31781,
         n31783, n31784, n31785, n31786, n31787, n31788, n31790, n31793,
         n31795, n31796, n31797, n31798, n31799, n31800, n31801, n31803,
         n31804, n31805, n31807, n31810, n31811, n31813, n31814, n31815,
         n31819, n31820, n31821, n31822, n31823, n31824, n31825, n31826,
         n31827, n31828, n31830, n31833, n31834, n31835, n31836, n31837,
         n31838, n31839, n31841, n31843, n31844, n31848, n31849, n31850,
         n31852, n31853, n31854, n31856, n31857, n31859, n31860, n31861,
         n31862, n31863, n31866, n31867, n31868, n31869, n31871, n31872,
         n31873, n31874, n31875, n31876, n31878, n31880, n31882, n31883,
         n31884, n31885, n31886, n31887, n31888, n31889, n31890, n31891,
         n31892, n31893, n31894, n31895, n31898, n31899, n31900, n31901,
         n31902, n31903, n31904, n31906, n31907, n31908, n31909, n31910,
         n31911, n31912, n31913, n31914, n31915, n31916, n31918, n31919,
         n31920, n31921, n31922, n31923, n31924, n31925, n31926, n31927,
         n31928, n31929, n31930, n31931, n31932, n31933, n31934, n31935,
         n31936, n31937, n31938, n31939, n31940, n31941, n31942, n31943,
         n31945, n31946, n31947, n31948, n31949, n31950, n31951, n31953,
         n31954, n31956, n31957, n31958, n31959, n31960, n31961, n31962,
         n31963, n31964, n31965, n31966, n31967, n31968, n31969, n31970,
         n31971, n31972, n31973, n31974, n31975, n31976, n31977, n31978,
         n31979, n31980, n31981, n31982, n31983, n31984, n31985, n31986,
         n31987, n31988, n31989, n31990, n31991, n31992, n31993, n31994,
         n31995, n31996, n31997, n31998, n31999, n32000, n32001, n32002,
         n32003, n32004, n32005, n32006, n32007, n32008, n32009, n32010,
         n32011, n32012, n32013, n32014, n32015, n32016, n32017, n32018,
         n32019, n32020, n32021, n32022, n32023, n32024, n32025, n32026,
         n32027, n32028, n32029, n32030, n32031, n32032, n32033, n32034,
         n32035, n32036, n32037, n32038, n32039, n32040, n32041, n32042,
         n32043, n32044, n32045, n32046, n32047, n32048, n32049, n32050,
         n32051, n32052, n32053, n32054, n32055, n32056, n32057, n32058,
         n32059, n32060, n32061, n32062, n32063, n32064, n32065, n32066,
         n32067, n32068, n32069, n32070, n32071, n32072, n32073, n32074,
         n32075, n32076, n32077, n32078, n32079, n32080, n32081, n32082,
         n32083, n32084, n32085, n32086, n32087, n32088, n32089, n32090,
         n32091, n32092, n32093, n32094, n32095, n32096, n32097, n32098,
         n32099, n32100, n32101, n32102, n32103, n32104, n32105, n32106,
         n32107, n32108, n32109, n32110, n32111, n32112, n32113, n32114,
         n32115, n32116, n32117, n32118, n32119, n32120, n32121, n32122,
         n32123, n32124, n32125, n32126, n32127, n32128, n32129, n32130,
         n32131, n32132, n32133, n32134, n32135, n32136, n32137, n32138,
         n32139, n32140, n32141, n32142, n32143, n32144, n32145, n32146,
         n32147, n32148, n32149, n32150, n32151, n32152, n32153, n32154,
         n32155, n32156, n32157, n32158, n32159, n32160, n32161, n32162,
         n32163, n32164, n32165, n32166, n32167, n32168, n32169, n32170,
         n32171, n32172, n32173, n32174, n32175, n32176, n32177, n32178,
         n32179, n32180, n32181, n32182, n32183, n32184, n32185, n32186,
         n32187, n32188, n32189, n32190, n32191, n32192, n32193, n32194,
         n32195, n32196, n32197, n32198, n32199, n32200, n32201, n32202,
         n32203, n32204, n32205, n32206, n32207, n32208, n32209, n32210,
         n32211, n32212, n32213, n32214, n32215, n32216, n32217, n32218,
         n32219, n32220, n32221, n32222, n32223, n32224, n32225, n32226,
         n32227, n32228, n32229, n32230, n32231, n32232, n32233, n32234,
         n32235, n32236, n32237, n32238, n32239, n32240, n32241, n32242,
         n32243, n32244, n32245, n32246, n32247, n32248, n32249, n32250,
         n32251, n32252, n32253, n32254, n32255, n32256, n32257, n32258,
         n32259, n32260, n32261, n32262, n32263, n32264, n32265, n32266,
         n32267, n32268, n32269, n32270, n32271, n32272, n32273, n32274,
         n32275, n32276, n32277, n32278, n32279, n32280, n32281, n32282,
         n32283, n32284, n32285, n32286, n32287, n32288, n32289, n32290,
         n32291, n32292, n32293, n32294, n32295, n32296, n32297, n32298,
         n32299, n32300, n32301, n32302, n32303, n32304, n32305, n32306,
         n32307, n32308, n32309, n32310, n32311, n32312, n32313, n32314,
         n32315, n32316, n32317, n32318, n32319, n32320, n32321, n32322,
         n32323, n32324, n32325, n32326, n32327, n32328, n32329, n32330,
         n32331, n32332, n32333, n32334, n32335, n32336, n32337, n32338,
         n32339, n32340, n32341, n32342, n32343, n32344, n32345, n32346,
         n32347, n32348, n32349, n32350, n32351, n32352, n32353, n32354,
         n32355, n32356, n32357, n32358, n32359, n32360, n32361, n32362,
         n32363, n32364, n32365, n32366, n32367, n32368, n32369, n32370,
         n32371, n32372, n32373, n32374, n32375, n32376, n32377, n32378,
         n32379, n32380, n32381, n32382, n32383, n32384, n32385, n32386,
         n32387, n32388, n32389, n32390, n32391, n32392, n32393, n32394,
         n32395, n32396, n32397, n32398, n32399, n32400, n32401, n32402,
         n32403, n32404, n32405, n32406, n32407, n32408, n32409, n32410,
         n32411, n32412, n32413, n32414, n32415, n32416, n32417, n32418,
         n32419, n32420, n32421, n32422, n32423, n32424, n32425, n32426,
         n32427, n32428, n32429, n32430, n32431, n32432, n32433, n32434,
         n32435, n32436, n32437, n32438, n32439, n32440, n32441, n32442,
         n32443, n32444, n32445, n32446, n32447, n32448, n32449, n32450,
         n32451, n32452, n32453, n32454, n32455, n32456, n32457, n32458,
         n32459, n32460, n32461, n32462, n32463, n32464, n32465, n32466,
         n32467, n32468, n32469, n32470, n32471, n32472, n32473, n32474,
         n32475, n32476, n32477, n32478, n32479, n32480, n32481, n32482,
         n32483, n32484, n32485, n32486, n32487, n32488, n32489, n32490,
         n32491, n32492, n32493, n32494, n32495, n32496, n32497, n32498,
         n32499, n32500, n32501, n32502, n32503, n32504, n32505, n32506,
         n32507, n32508, n32509, n32510, n32511, n32512, n32513, n32514,
         n32515, n32516, n32517, n32518, n32519, n32520, n32521, n32522,
         n32523, n32524, n32525, n32526, n32527, n32528, n32529, n32530,
         n32531, n32532, n32533, n32534, n32535, n32536, n32537, n32538,
         n32539, n32540, n32541, n32542, n32543, n32544, n32545, n32546,
         n32547, n32548, n32549, n32550, n32551, n32552, n32553, n32554,
         n32555, n32556, n32557, n32558, n32559, n32560, n32561, n32562,
         n32563, n32564, n32565, n32566, n32567, n32568, n32569, n32570,
         n32571, n32572, n32573, n32574, n32575, n32576, n32577, n32578,
         n32579, n32580, n32581, n32582, n32583, n32584, n32585, n32586,
         n32587, n32588, n32589, n32590, n32591, n32592, n32593, n32594,
         n32595, n32596, n32597, n32598, n32599, n32600, n32601, n32602,
         n32603, n32604, n32605, n32606, n32607, n32608, n32609, n32610,
         n32611, n32612, n32613, n32614, n32615, n32616, n32617, n32618,
         n32619, n32620, n32621, n32622, n32623, n32624, n32625, n32626,
         n32627, n32628, n32629, n32630, n32631, n32632, n32633, n32634,
         n32635, n32636, n32637, n32638, n32639, n32640, n32641, n32642,
         n32643, n32644, n32645, n32646, n32647, n32648, n32649, n32650,
         n32651, n32652, n32653, n32654, n32655, n32656, n32657, n32658,
         n32659, n32660, n32661, n32662, n32663, n32664, n32665, n32666,
         n32667, n32668, n32669, n32670, n32671, n32672, n32673, n32674,
         n32675, n32676, n32677, n32678, n32679, n32680, n32681, n32682,
         n32683, n32684, n32685, n32686, n32687, n32688, n32689, n32690,
         n32691, n32692, n32693, n32694, n32695, n32696, n32697, n32698,
         n32699, n32700, n32701, n32702, n32703, n32704, n32705, n32706,
         n32707, n32708, n32709, n32710, n32711, n32712, n32713, n32714,
         n32715, n32716, n32717, n32718, n32719, n32720, n32721, n32722,
         n32723, n32724, n32725, n32726, n32727, n32728, n32729, n32730,
         n32731, n32732, n32733, n32734, n32735, n32736, n32737, n32738,
         n32739, n32740, n32741, n32742, n32743, n32744, n32745, n32746,
         n32747, n32748, n32749, n32750, n32751, n32752, n32753, n32754,
         n32755, n32756, n32757, n32758, n32759, n32760, n32761, n32762,
         n32763, n32764, n32765, n32766, n32767, n32768, n32769, n32770,
         n32771, n32772, n32773, n32774, n32775, n32776, n32777, n32778,
         n32779, n32780, n32781, n32782, n32783, n32784, n32785, n32786,
         n32787, n32788, n32789, n32790, n32791, n32792, n32793, n32794,
         n32795, n32796, n32797, n32798, n32799, n32800, n32801, n32802,
         n32803, n32804, n32805, n32806, n32807, n32808, n32809, n32810,
         n32811, n32812, n32813, n32814, n32815, n32816, n32817, n32818,
         n32819, n32820, n32821, n32822, n32823, n32824, n32825, n32826,
         n32827, n32828, n32829, n32830, n32831, n32832, n32833, n32834,
         n32835, n32836, n32837, n32838, n32839, n32840, n32841, n32842,
         n32843, n32844, n32845, n32846, n32847, n32848, n32849, n32850,
         n32851, n32852, n32853, n32854, n32855, n32856, n32857, n32858,
         n32859, n32860, n32861, n32862, n32863, n32864, n32865, n32866,
         n32867, n32868, n32869, n32870, n32871, n32872, n32873, n32874,
         n32875, n32876, n32877, n32878, n32879, n32880, n32881, n32882,
         n32883, n32884, n32885, n32886, n32887, n32888, n32889, n32890,
         n32891, n32892, n32893, n32894, n32895, n32896, n32897, n32898,
         n32899, n32900, n32901, n32902, n32903, n32904, n32905, n32906,
         n32907, n32908, n32909, n32910, n32911, n32912, n32913, n32914,
         n32915, n32916, n32917, n32918, n32919, n32920, n32921, n32922,
         n32923, n32924, n32925, n32926, n32927, n32928, n32929, n32930,
         n32931, n32932, n32933, n32934, n32935, n32936, n32937, n32938,
         n32939, n32940, n32941, n32942, n32943, n32945, n32946, n32947,
         n32948, n32949, n32950, n32951, n32952, n32953, n32954, n32955,
         n32956, n32957, n32958, n32959, n32960, n32961, n32962, n32963,
         n32964, n32965, n32966, n32967, n32968, n32969, n32970, n32971,
         n32972, n32973, n32974, n32975, n32976, n32977, n32978, n32979,
         n32980, n32981, n32983, n32984, n32985, n32986, n32987, n32988,
         n32989, n32990, n32991, n32992, n32993, n32994, n32995, n32996,
         n32997, n32998, n32999, n33001, n33002, n33003, n33004, n33005,
         n33006, n33007, n33008, n33009, n33010, n33011, n33012, n33013,
         n33014, n33015, n33016, n33017, n33018, n33019, n33020, n33021,
         n33022, n33023, n33024, n33025, n33026, n33027, n33028, n33029,
         n33030, n33031, n33032, n33033, n33034, n33035, n33036, n33037,
         n33038, n33039, n33040, n33041, n33042, n33043, n33044, n33045,
         n33046, n33047, n33048, n33049, n33050, n33051, n33052, n33053,
         n33054, n33055, n33056, n33057, n33058, n33059, n33060, n33061,
         n33062, n33063, n33064, n33065, n33066, n33067, n33068, n33069,
         n33070, n33071, n33072, n33073, n33074, n33075, n33076, n33077,
         n33078, n33079, n33080, n33081, n33082, n33083, n33084, n33085,
         n33086, n33087, n33088, n33089, n33090, n33091, n33092, n33093,
         n33094, n33095, n33096, n33097, n33098, n33099, n33100, n33101,
         n33102, n33103, n33104, n33105, n33106, n33107, n33108, n33109,
         n33110, n33111, n33112, n33113, n33114, n33115, n33116, n33117,
         n33118, n33119, n33120, n33121, n33122, n33123, n33124, n33125,
         n33126, n33127, n33128, n33129, n33130, n33131, n33132, n33133,
         n33134, n33135, n33136, n33137, n33138, n33139, n33140, n33141,
         n33142, n33143, n33144, n33145, n33146, n33147, n33148, n33149,
         n33150, n33151, n33152, n33153, n33154, n33155, n33156, n33157,
         n33158, n33159, n33160, n33161, n33162, n33163, n33164, n33165,
         n33166, n33167, n33168, n33169, n33170, n33171, n33172, n33173,
         n33174, n33175, n33176, n33177, n33178, n33179, n33180, n33181,
         n33182, n33183, n33184, n33185, n33186, n33187, n33188, n33189,
         n33190, n33191, n33192, n33193, n33194, n33195, n33196, n33197,
         n33198, n33199, n33200, n33201, n33202, n33203, n33204, n33205,
         n33206, n33207, n33208, n33209, n33210, n33211, n33212, n33213,
         n33214, n33215, n33216, n33217, n33218, n33219, n33220, n33221,
         n33222, n33223, n33224, n33225, n33226, n33227, n33228, n33229,
         n33230, n33231, n33232, n33233, n33234, n33235, n33236, n33237,
         n33238, n33239, n33240, n33241, n33242, n33243, n33244, n33245,
         n33246, n33247, n33248, n33249, n33250, n33251, n33252, n33253,
         n33254, n33255, n33256, n33257, n33258, n33259, n33260, n33261,
         n33262, n33263, n33264, n33265, n33266, n33267, n33268, n33269,
         n33270, n33271, n33272, n33273, n33274, n33275, n33276, n33277,
         n33278, n33279, n33280, n33281, n33282, n33283, n33284, n33285,
         n33286, n33287, n33288, n33289, n33290, n33291, n33292, n33293,
         n33294, n33295, n33296, n33297, n33298, n33299, n33300, n33301,
         n33302, n33303, n33304, n33305, n33306, n33307, n33308, n33309,
         n33310, n33311, n33312, n33313, n33314, n33315, n33316, n33317,
         n33318, n33319, n33320, n33321, n33322, n33323, n33324, n33325,
         n33326, n33327, n33328, n33329, n33330, n33331, n33332, n33333,
         n33334, n33335, n33336, n33337, n33338, n33339, n33340, n33341,
         n33342, n33343, n33344, n33345, n33346, n33347, n33348, n33349,
         n33350, n33351, n33352, n33353, n33354, n33355, n33356, n33357,
         n33358, n33359, n33360, n33361, n33362, n33363, n33364, n33365,
         n33366, n33367, n33368, n33369, n33370, n33371, n33372, n33373,
         n33374, n33375, n33376, n33377, n33378, n33379, n33380, n33381,
         n33382, n33383, n33384, n33385, n33386, n33387, n33388, n33389,
         n33390, n33391, n33392, n33393, n33394, n33395, n33396, n33397,
         n33398, n33399, n33400, n33401, n33402, n33403, n33404, n33405,
         n33406, n33407, n33408, n33409, n33410, n33411, n33412, n33413,
         n33414, n33415, n33416, n33417, n33418, n33419, n33420, n33421,
         n33422, n33423, n33424, n33425, n33426, n33427, n33428, n33429,
         n33430, n33431, n33432, n33433, n33434, n33435, n33436, n33437,
         n33438, n33439, n33440, n33441, n33442, n33443, n33444, n33445,
         n33446, n33447, n33448, n33449, n33450, n33451, n33452, n33453,
         n33454, n33455, n33456, n33457, n33458, n33459, n33460, n33461,
         n33462, n33463, n33464, n33465, n33466, n33467, n33468, n33469,
         n33470, n33471, n33472, n33473, n33474, n33475, n33476, n33477,
         n33478, n33479, n33480, n33481, n33482, n33483, n33484, n33485,
         n33486, n33487, n33488, n33489, n33490, n33491, n33492, n33493,
         n33494, n33495, n33496, n33497, n33498, n33499, n33500, n33501,
         n33502, n33503, n33504, n33505, n33506, n33507, n33508, n33509,
         n33510, n33511, n33512, n33513, n33514, n33515, n33516, n33517,
         n33518, n33519, n33520, n33521, n33522, n33523, n33524, n33525,
         n33526, n33527, n33528, n33529, n33530, n33531, n33532, n33533,
         n33534, n33535, n33536, n33537, n33538, n33539, n33540, n33541,
         n33542, n33543, n33544, n33545, n33546, n33547, n33548, n33549,
         n33550, n33551, n33552, n33553, n33554, n33555, n33556, n33557,
         n33558, n33559, n33560, n33561, n33562, n33563, n33564, n33565,
         n33566, n33567, n33568, n33569, n33570, n33571, n33572, n33573,
         n33574, n33575, n33576, n33577, n33578, n33579, n33580, n33581,
         n33582, n33583, n33584, n33585, n33586, n33587, n33588, n33589,
         n33590, n33591, n33593, n33594, n33595, n33596, n33597, n33598,
         n33599, n33600, n33601, n33602, n33603, n33604, n33605, n33606,
         n33607, n33608, n33609, n33610, n33611, n33612, n33613, n33614,
         n33615, n33616, n33617, n33618, n33619, n33620, n33621, n33622,
         n33623, n33624, n33625, n33626, n33627, n33628, n33629, n33630,
         n33631, n33632, n33633, n33634, n33635, n33636, n33637, n33638,
         n33639, n33640, n33641, n33642, n33643, n33644, n33645, n33646,
         n33647, n33648, n33649, n33650, n33651, n33652, n33653, n33654,
         n33655, n33656, n33657, n33658, n33659, n33660, n33661, n33662,
         n33663, n33664, n33665, n33666, n33667, n33668, n33669, n33670,
         n33671, n33672, n33673, n33674, n33675, n33676, n33677, n33678,
         n33679, n33680, n33681, n33682, n33683, n33684, n33685, n33686,
         n33687, n33688, n33689, n33690, n33691, n33692, n33693, n33694,
         n33695, n33696, n33697, n33698, n33699, n33700, n33701, n33702,
         n33703, n33704, n33705, n33706, n33707, n33708, n33709, n33710,
         n33711, n33712, n33713, n33714, n33715, n33716, n33717, n33718,
         n33719, n33720, n33721, n33722, n33723, n33724, n33725, n33726,
         n33727, n33728, n33729, n33730, n33731, n33732, n33733, n33734,
         n33735, n33736, n33737, n33738, n33739, n33740, n33741, n33742,
         n33743, n33744, n33745, n33746, n33747, n33748, n33749, n33750,
         n33751, n33752, n33753, n33754, n33755, n33756, n33757, n33758,
         n33759, n33760, n33761, n33762, n33763, n33764, n33765, n33766,
         n33767, n33768, n33769, n33770, n33771, n33772, n33773, n33774,
         n33775, n33776, n33777, n33778, n33779, n33780, n33781, n33782,
         n33783, n33784, n33785, n33786, n33787, n33788, n33789, n33790,
         n33791, n33792, n33793, n33794, n33795, n33796, n33797, n33798,
         n33799, n33800, n33801, n33802, n33803, n33804, n33805, n33806,
         n33807, n33808, n33809, n33810, n33811, n33812, n33813, n33814,
         n33815, n33816, n33817, n33818, n33819, n33820, n33821, n33822,
         n33823, n33824, n33825, n33826, n33827, n33828, n33829, n33830,
         n33831, n33832, n33833, n33834, n33835, n33836, n33837, n33838,
         n33839, n33840, n33841, n33842, n33843, n33844, n33845, n33846,
         n33847, n33848, n33849, n33850, n33851, n33852, n33853, n33854,
         n33855, n33856, n33857, n33858, n33859, n33860, n33861, n33862,
         n33863, n33864, n33865, n33866, n33867, n33868, n33869, n33870,
         n33871, n33872, n33873, n33874, n33875, n33876, n33877, n33878,
         n33879, n33880, n33881, n33882, n33883, n33884, n33885, n33886,
         n33887, n33888, n33889, n33890, n33891, n33892, n33893, n33894,
         n33895, n33896, n33897, n33898, n33899, n33900, n33901, n33902,
         n33903, n33904, n33905, n33906, n33907, n33908, n33909, n33910,
         n33911, n33912, n33913, n33914, n33915, n33916, n33917, n33918,
         n33919, n33920, n33921, n33922, n33923, n33924, n33925, n33926,
         n33927, n33928, n33929, n33930, n33931, n33932, n33933, n33934,
         n33935, n33936, n33937, n33938, n33939, n33940, n33941, n33942,
         n33943, n33944, n33945, n33946, n33947, n33948, n33949, n33950,
         n33951, n33952, n33953, n33954, n33955, n33956, n33957, n33958,
         n33959, n33960, n33961, n33962, n33963, n33964, n33965, n33966,
         n33967, n33968, n33969, n33970, n33971, n33972, n33973, n33974,
         n33975, n33976, n33977, n33978, n33979, n33980, n33981, n33982,
         n33983, n33984, n33985, n33986, n33987, n33988, n33989, n33990,
         n33991, n33992, n33993, n33994, n33995, n33996, n33997, n33998,
         n33999, n34000, n34001, n34002, n34003, n34004, n34005, n34006,
         n34007, n34008, n34009, n34010, n34011, n34012, n34013, n34014,
         n34015, n34016, n34017, n34018, n34019, n34020, n34021, n34022,
         n34023, n34024, n34025, n34026, n34027, n34028, n34029, n34030,
         n34031, n34032, n34033, n34034, n34035, n34036, n34037, n34038,
         n34039, n34040, n34041, n34042, n34043, n34044, n34045, n34046,
         n34047, n34048, n34049, n34050, n34051, n34052, n34053, n34054,
         n34055, n34056, n34057, n34058, n34059, n34060, n34061, n34062,
         n34063, n34064, n34065, n34066, n34067, n34068, n34069, n34070,
         n34071, n34072, n34073, n34074, n34075, n34076, n34077, n34078,
         n34079, n34080, n34081, n34082, n34083, n34084, n34085, n34086,
         n34087, n34088, n34089, n34090, n34091, n34092, n34093, n34094,
         n34095, n34096, n34097, n34098, n34099, n34100, n34101, n34102,
         n34103, n34104, n34105, n34106, n34107, n34108, n34109, n34110,
         n34111, n34112, n34113, n34114, n34115, n34116, n34117, n34118,
         n34119, n34120, n34121, n34122, n34123, n34124, n34125, n34126,
         n34127, n34128, n34129, n34130, n34131, n34132, n34133, n34134,
         n34135, n34136, n34137, n34138, n34139, n34140, n34141, n34142,
         n34143, n34144, n34145, n34146, n34147, n34148, n34149, n34150,
         n34151, n34152, n34153, n34154, n34155, n34156, n34157, n34158,
         n34159, n34160, n34161, n34162, n34163, n34164, n34165, n34166,
         n34167, n34168, n34169, n34170;

  NAND2_X1 U2 ( .A1(n5901), .A2(n964), .ZN(n433) );
  NOR2_X1 U10 ( .A1(n17637), .A2(n25517), .ZN(n25509) );
  NAND3_X1 U35 ( .A1(n24584), .A2(n24583), .A3(n24582), .ZN(n10608) );
  NAND2_X1 U39 ( .A1(n10174), .A2(n32856), .ZN(n10173) );
  INV_X1 U130 ( .I(n13236), .ZN(n24592) );
  INV_X1 U138 ( .I(n5284), .ZN(n24782) );
  NAND2_X1 U145 ( .A1(n2444), .A2(n23618), .ZN(n214) );
  NOR2_X1 U192 ( .A1(n24271), .A2(n29307), .ZN(n2923) );
  NAND2_X1 U251 ( .A1(n16676), .A2(n13549), .ZN(n7504) );
  INV_X2 U278 ( .I(n33722), .ZN(n16786) );
  INV_X1 U313 ( .I(n23450), .ZN(n169) );
  INV_X1 U317 ( .I(n24386), .ZN(n12797) );
  INV_X1 U320 ( .I(n23534), .ZN(n23227) );
  INV_X1 U325 ( .I(n16703), .ZN(n18122) );
  INV_X1 U330 ( .I(n29885), .ZN(n8883) );
  INV_X1 U371 ( .I(n13679), .ZN(n13751) );
  INV_X1 U390 ( .I(n12729), .ZN(n11308) );
  INV_X2 U429 ( .I(n2860), .ZN(n1106) );
  NAND2_X1 U438 ( .A1(n11250), .A2(n29287), .ZN(n22685) );
  AOI21_X1 U442 ( .A1(n22672), .A2(n29304), .B(n9753), .ZN(n22673) );
  INV_X1 U447 ( .I(n17151), .ZN(n22577) );
  OR2_X1 U452 ( .A1(n639), .A2(n9953), .Z(n22682) );
  NAND2_X1 U487 ( .A1(n22562), .A2(n22403), .ZN(n6384) );
  INV_X1 U489 ( .I(n22679), .ZN(n22562) );
  INV_X1 U512 ( .I(n21958), .ZN(n1306) );
  OR2_X1 U554 ( .A1(n31511), .A2(n21651), .Z(n21641) );
  INV_X1 U577 ( .I(n21708), .ZN(n9119) );
  NAND2_X1 U586 ( .A1(n21491), .A2(n21568), .ZN(n21492) );
  NOR2_X1 U680 ( .A1(n21374), .A2(n4145), .ZN(n15814) );
  INV_X2 U695 ( .I(n21203), .ZN(n21400) );
  OAI21_X1 U738 ( .A1(n27177), .A2(n1034), .B(n3787), .ZN(n3558) );
  NAND3_X1 U752 ( .A1(n20591), .A2(n20589), .A3(n384), .ZN(n20173) );
  CLKBUF_X2 U760 ( .I(n15230), .Z(n8353) );
  INV_X2 U780 ( .I(n17544), .ZN(n20486) );
  OAI21_X1 U802 ( .A1(n11909), .A2(n16065), .B(n6644), .ZN(n10056) );
  NAND2_X1 U804 ( .A1(n1826), .A2(n402), .ZN(n9015) );
  NOR2_X1 U815 ( .A1(n10086), .A2(n6200), .ZN(n402) );
  NAND3_X1 U818 ( .A1(n25997), .A2(n16), .A3(n13747), .ZN(n15435) );
  INV_X2 U876 ( .I(n28951), .ZN(n1044) );
  INV_X1 U882 ( .I(n25208), .ZN(n293) );
  INV_X1 U884 ( .I(n15960), .ZN(n876) );
  INV_X1 U891 ( .I(n2581), .ZN(n18840) );
  INV_X2 U954 ( .I(n9319), .ZN(n7687) );
  INV_X1 U958 ( .I(n6846), .ZN(n18913) );
  NAND2_X1 U963 ( .A1(n7900), .A2(n30744), .ZN(n436) );
  INV_X1 U970 ( .I(n31971), .ZN(n952) );
  NAND2_X1 U994 ( .A1(n18515), .A2(n13663), .ZN(n16086) );
  INV_X1 U1011 ( .I(n18700), .ZN(n18007) );
  INV_X2 U1014 ( .I(n494), .ZN(n1188) );
  NAND2_X2 U1027 ( .A1(n34037), .A2(n1333), .ZN(n1915) );
  NOR2_X2 U1061 ( .A1(n21715), .A2(n21601), .ZN(n21710) );
  NAND2_X2 U1070 ( .A1(n29185), .A2(n23721), .ZN(n13342) );
  INV_X2 U1088 ( .I(n18018), .ZN(n18616) );
  NAND2_X2 U1102 ( .A1(n14246), .A2(n27182), .ZN(n25404) );
  INV_X2 U1162 ( .I(n13442), .ZN(n13816) );
  NOR2_X2 U1167 ( .A1(n20361), .A2(n27887), .ZN(n20451) );
  NOR2_X2 U1178 ( .A1(n25891), .A2(n25890), .ZN(n9941) );
  INV_X2 U1299 ( .I(n10335), .ZN(n17456) );
  NOR2_X2 U1317 ( .A1(n3455), .A2(n9800), .ZN(n3124) );
  OAI22_X2 U1353 ( .A1(n1143), .A2(n21237), .B1(n424), .B2(n780), .ZN(n12836)
         );
  INV_X2 U1384 ( .I(n16748), .ZN(n14198) );
  INV_X4 U1415 ( .I(n4656), .ZN(n19301) );
  AOI22_X2 U1424 ( .A1(n3189), .A2(n1720), .B1(n3188), .B2(n1120), .ZN(n3187)
         );
  NAND2_X2 U1440 ( .A1(n1384), .A2(n18990), .ZN(n19091) );
  NAND2_X2 U1452 ( .A1(n7600), .A2(n19255), .ZN(n2177) );
  INV_X2 U1465 ( .I(n17352), .ZN(n23904) );
  INV_X2 U1470 ( .I(n18674), .ZN(n18881) );
  BUF_X2 U1482 ( .I(n22535), .Z(n16434) );
  INV_X2 U1517 ( .I(n18990), .ZN(n878) );
  BUF_X4 U1528 ( .I(n16801), .Z(n10828) );
  NAND2_X2 U1536 ( .A1(n8787), .A2(n19115), .ZN(n19186) );
  BUF_X2 U1543 ( .I(n29781), .Z(n2582) );
  AOI21_X2 U1548 ( .A1(n18347), .A2(n18346), .B(n18345), .ZN(n2331) );
  NOR2_X1 U1557 ( .A1(n25971), .A2(n16740), .ZN(n16876) );
  NAND3_X1 U1559 ( .A1(n1358), .A2(n13327), .A3(n19949), .ZN(n20191) );
  OAI21_X1 U1569 ( .A1(n31407), .A2(n1074), .B(n694), .ZN(n66) );
  NAND2_X1 U1571 ( .A1(n14764), .A2(n712), .ZN(n14763) );
  INV_X1 U1616 ( .I(n5492), .ZN(n5113) );
  NOR2_X1 U1624 ( .A1(n33563), .A2(n268), .ZN(n17336) );
  INV_X2 U1625 ( .I(n11984), .ZN(n13499) );
  NAND2_X2 U1630 ( .A1(n14311), .A2(n11831), .ZN(n24548) );
  NAND2_X1 U1648 ( .A1(n16800), .A2(n29866), .ZN(n363) );
  NAND3_X1 U1651 ( .A1(n4770), .A2(n786), .A3(n4782), .ZN(n3433) );
  AOI21_X1 U1678 ( .A1(n21669), .A2(n21672), .B(n16345), .ZN(n21278) );
  NAND2_X1 U1685 ( .A1(n22919), .A2(n8365), .ZN(n268) );
  INV_X2 U1727 ( .I(n19641), .ZN(n1045) );
  NAND2_X1 U1736 ( .A1(n3722), .A2(n3723), .ZN(n15796) );
  OR2_X2 U1749 ( .A1(n5392), .A2(n11847), .Z(n21202) );
  INV_X1 U1766 ( .I(n18310), .ZN(n1184) );
  NAND2_X2 U1771 ( .A1(n17334), .A2(n17335), .ZN(n23346) );
  OAI21_X2 U1779 ( .A1(n827), .A2(n29), .B(n19050), .ZN(n13448) );
  XOR2_X1 U1788 ( .A1(n2278), .A2(n31259), .Z(n12011) );
  NOR2_X2 U1806 ( .A1(n12074), .A2(n16766), .ZN(n14284) );
  NAND2_X1 U1807 ( .A1(n24138), .A2(n16286), .ZN(n6980) );
  INV_X2 U1810 ( .I(n9436), .ZN(n11372) );
  NAND2_X1 U1820 ( .A1(n9695), .A2(n9697), .ZN(n13065) );
  NOR2_X1 U1821 ( .A1(n27123), .A2(n10858), .ZN(n9696) );
  INV_X2 U1830 ( .I(n12241), .ZN(n13852) );
  NAND2_X2 U1836 ( .A1(n11), .A2(n4209), .ZN(n20468) );
  BUF_X2 U1844 ( .I(n24117), .Z(n13) );
  INV_X2 U1849 ( .I(n5837), .ZN(n17495) );
  AOI21_X2 U1876 ( .A1(n17371), .A2(n28219), .B(n15366), .ZN(n9099) );
  INV_X1 U1877 ( .I(n25985), .ZN(n8450) );
  XOR2_X1 U1890 ( .A1(n18948), .A2(n17613), .Z(n367) );
  BUF_X2 U1898 ( .I(n18700), .Z(n22) );
  XOR2_X1 U1901 ( .A1(n24837), .A2(n16504), .Z(n13849) );
  AOI21_X2 U1908 ( .A1(n15585), .A2(n17234), .B(n14778), .ZN(n15584) );
  AOI21_X2 U1913 ( .A1(n6069), .A2(n761), .B(n4162), .ZN(n6068) );
  NAND2_X2 U1920 ( .A1(n6074), .A2(n21581), .ZN(n21666) );
  XOR2_X1 U1923 ( .A1(n8861), .A2(n10328), .Z(n3304) );
  AOI21_X2 U1936 ( .A1(n22607), .A2(n9155), .B(n5958), .ZN(n23110) );
  AND2_X1 U1943 ( .A1(n28338), .A2(n29279), .Z(n696) );
  XOR2_X1 U1954 ( .A1(n29277), .A2(n31), .Z(n4951) );
  XOR2_X1 U1955 ( .A1(n24538), .A2(n14079), .Z(n31) );
  XOR2_X1 U1957 ( .A1(n23473), .A2(n11667), .Z(n4661) );
  XOR2_X1 U1960 ( .A1(n7566), .A2(n34), .Z(n606) );
  XOR2_X1 U1961 ( .A1(n7565), .A2(n29413), .Z(n34) );
  BUF_X2 U1982 ( .I(Key[54]), .Z(n16690) );
  INV_X4 U1987 ( .I(n18683), .ZN(n1659) );
  XOR2_X1 U1996 ( .A1(n29275), .A2(n44), .Z(n5965) );
  XOR2_X1 U1997 ( .A1(n24773), .A2(n24476), .Z(n44) );
  NAND2_X2 U2014 ( .A1(n18400), .A2(n46), .ZN(n19294) );
  XOR2_X1 U2024 ( .A1(n4986), .A2(n702), .Z(n4984) );
  XOR2_X1 U2034 ( .A1(n52), .A2(n14809), .Z(n15733) );
  XOR2_X1 U2041 ( .A1(n23463), .A2(n54), .Z(n14783) );
  XOR2_X1 U2042 ( .A1(n23299), .A2(n23489), .Z(n54) );
  XOR2_X1 U2070 ( .A1(n23136), .A2(n62), .Z(n17591) );
  XOR2_X1 U2071 ( .A1(n26101), .A2(n14818), .Z(n62) );
  NAND2_X2 U2076 ( .A1(n2677), .A2(n16084), .ZN(n20529) );
  NAND2_X2 U2082 ( .A1(n16669), .A2(n31324), .ZN(n17239) );
  NAND2_X1 U2101 ( .A1(n18462), .A2(n18463), .ZN(n94) );
  AOI21_X2 U2102 ( .A1(n4879), .A2(n4643), .B(n8091), .ZN(n4878) );
  INV_X2 U2116 ( .I(n11562), .ZN(n22139) );
  NAND2_X2 U2150 ( .A1(n28904), .A2(n3157), .ZN(n20334) );
  XOR2_X1 U2151 ( .A1(n81), .A2(n23132), .Z(n23263) );
  NAND2_X2 U2157 ( .A1(n21559), .A2(n6489), .ZN(n21821) );
  XOR2_X1 U2162 ( .A1(n10399), .A2(n6571), .Z(n86) );
  INV_X2 U2165 ( .I(n87), .ZN(n563) );
  INV_X2 U2168 ( .I(n14980), .ZN(n13759) );
  OR2_X1 U2179 ( .A1(n14212), .A2(n28891), .Z(n4611) );
  NAND2_X1 U2185 ( .A1(n11419), .A2(n15835), .ZN(n92) );
  NAND2_X1 U2211 ( .A1(n33583), .A2(n31807), .ZN(n97) );
  OAI21_X1 U2243 ( .A1(n25278), .A2(n12431), .B(n25284), .ZN(n16290) );
  INV_X4 U2247 ( .I(n4746), .ZN(n15179) );
  INV_X2 U2251 ( .I(n11833), .ZN(n22926) );
  NAND2_X1 U2252 ( .A1(n107), .A2(n16347), .ZN(n25255) );
  OAI21_X2 U2265 ( .A1(n21298), .A2(n15807), .B(n21299), .ZN(n21721) );
  BUF_X4 U2292 ( .I(n9125), .Z(n9127) );
  NAND2_X2 U2294 ( .A1(n7144), .A2(n17888), .ZN(n21877) );
  XOR2_X1 U2302 ( .A1(n20746), .A2(n3209), .Z(n11689) );
  XOR2_X1 U2308 ( .A1(n16917), .A2(n6973), .Z(n119) );
  AOI21_X2 U2330 ( .A1(n11709), .A2(n9854), .B(n124), .ZN(n20727) );
  XOR2_X1 U2341 ( .A1(n34160), .A2(n22072), .Z(n22307) );
  XOR2_X1 U2343 ( .A1(n19554), .A2(n26032), .Z(n128) );
  NOR2_X1 U2348 ( .A1(n4953), .A2(n17927), .ZN(n4952) );
  OAI21_X1 U2367 ( .A1(n25526), .A2(n15295), .B(n15155), .ZN(n25527) );
  INV_X2 U2377 ( .I(n10371), .ZN(n8778) );
  NOR2_X2 U2379 ( .A1(n1352), .A2(n14545), .ZN(n10323) );
  XOR2_X1 U2381 ( .A1(n15353), .A2(n136), .Z(n10558) );
  XOR2_X1 U2382 ( .A1(n15352), .A2(n20962), .Z(n136) );
  OAI21_X1 U2386 ( .A1(n25488), .A2(n25487), .B(n25486), .ZN(n138) );
  XOR2_X1 U2388 ( .A1(n16693), .A2(n25190), .Z(n139) );
  NAND2_X2 U2390 ( .A1(n7278), .A2(n7277), .ZN(n12491) );
  INV_X2 U2394 ( .I(n23949), .ZN(n23947) );
  INV_X2 U2407 ( .I(n3340), .ZN(n19236) );
  INV_X2 U2419 ( .I(n4113), .ZN(n18241) );
  OAI22_X1 U2426 ( .A1(n25668), .A2(n9365), .B1(n25645), .B2(n25651), .ZN(
        n25642) );
  INV_X2 U2432 ( .I(n18884), .ZN(n18662) );
  BUF_X4 U2436 ( .I(n14702), .Z(n1337) );
  INV_X2 U2438 ( .I(n10146), .ZN(n24811) );
  NOR2_X2 U2449 ( .A1(n11759), .A2(n152), .ZN(n17927) );
  XOR2_X1 U2456 ( .A1(n153), .A2(n25195), .Z(Ciphertext[71]) );
  NAND3_X1 U2457 ( .A1(n4767), .A2(n4768), .A3(n4769), .ZN(n153) );
  INV_X2 U2459 ( .I(n12811), .ZN(n12992) );
  NAND2_X2 U2462 ( .A1(n7492), .A2(n5455), .ZN(n11074) );
  NAND2_X2 U2488 ( .A1(n4337), .A2(n28701), .ZN(n20940) );
  OAI21_X2 U2491 ( .A1(n16712), .A2(n10778), .B(n28240), .ZN(n10777) );
  XOR2_X1 U2497 ( .A1(n21035), .A2(n1993), .Z(n11424) );
  NAND2_X2 U2498 ( .A1(n11617), .A2(n11618), .ZN(n21035) );
  NAND2_X2 U2503 ( .A1(n21812), .A2(n18184), .ZN(n11848) );
  OR2_X2 U2511 ( .A1(n1850), .A2(n28591), .Z(n12247) );
  XOR2_X1 U2523 ( .A1(n1454), .A2(n168), .Z(n652) );
  XOR2_X1 U2524 ( .A1(n23199), .A2(n169), .Z(n168) );
  XOR2_X1 U2528 ( .A1(n170), .A2(n29108), .Z(n17535) );
  XOR2_X1 U2529 ( .A1(n6417), .A2(n15334), .Z(n170) );
  XOR2_X1 U2538 ( .A1(n175), .A2(n12062), .Z(n18037) );
  NAND2_X2 U2540 ( .A1(n15166), .A2(n15165), .ZN(n18997) );
  XOR2_X1 U2553 ( .A1(n3504), .A2(n5051), .Z(n24549) );
  XOR2_X1 U2558 ( .A1(n5231), .A2(n5229), .Z(n25112) );
  AOI22_X2 U2564 ( .A1(n11815), .A2(n18556), .B1(n16564), .B2(n18328), .ZN(
        n5892) );
  NAND3_X2 U2565 ( .A1(n5890), .A2(n5892), .A3(n5891), .ZN(n5545) );
  OR2_X1 U2575 ( .A1(n21733), .A2(n13872), .Z(n187) );
  INV_X2 U2579 ( .I(n10327), .ZN(n17814) );
  INV_X2 U2594 ( .I(n193), .ZN(n502) );
  XOR2_X1 U2595 ( .A1(n5151), .A2(n5152), .Z(n193) );
  INV_X2 U2596 ( .I(n29814), .ZN(n1353) );
  INV_X2 U2627 ( .I(n3967), .ZN(n19907) );
  XOR2_X1 U2631 ( .A1(n21990), .A2(n29259), .Z(n13704) );
  OAI21_X2 U2632 ( .A1(n6117), .A2(n15697), .B(n6116), .ZN(n7134) );
  XOR2_X1 U2634 ( .A1(n7674), .A2(n26085), .Z(n15309) );
  XOR2_X1 U2651 ( .A1(n2330), .A2(n19467), .Z(n2335) );
  NAND3_X1 U2653 ( .A1(n20361), .A2(n27887), .A3(n10939), .ZN(n5349) );
  INV_X4 U2659 ( .I(n17408), .ZN(n22705) );
  OR2_X1 U2661 ( .A1(n9719), .A2(n20375), .Z(n204) );
  NAND2_X1 U2672 ( .A1(n2209), .A2(n6288), .ZN(n13023) );
  INV_X2 U2674 ( .I(n625), .ZN(n5440) );
  OAI21_X2 U2709 ( .A1(n18956), .A2(n784), .B(n13009), .ZN(n13482) );
  XOR2_X1 U2717 ( .A1(n23254), .A2(n22841), .Z(n225) );
  XOR2_X1 U2726 ( .A1(n29194), .A2(n6923), .Z(n227) );
  XOR2_X1 U2734 ( .A1(n22230), .A2(n233), .Z(n17284) );
  XOR2_X1 U2735 ( .A1(n32084), .A2(n22092), .Z(n233) );
  NAND2_X2 U2751 ( .A1(n19283), .A2(n19285), .ZN(n19080) );
  NOR2_X2 U2756 ( .A1(n1864), .A2(n6073), .ZN(n10717) );
  INV_X4 U2786 ( .I(n5610), .ZN(n1378) );
  INV_X2 U2827 ( .I(n23143), .ZN(n23211) );
  NAND2_X1 U2856 ( .A1(n20573), .A2(n20572), .ZN(n258) );
  AOI21_X1 U2859 ( .A1(n7680), .A2(n16274), .B(n259), .ZN(n19250) );
  XOR2_X1 U2868 ( .A1(n30443), .A2(n19494), .Z(n19431) );
  OAI21_X2 U2869 ( .A1(n1451), .A2(n1453), .B(n1450), .ZN(n19494) );
  NAND2_X2 U2872 ( .A1(n9967), .A2(n11452), .ZN(n21651) );
  NAND2_X1 U2885 ( .A1(n5948), .A2(n12654), .ZN(n262) );
  OAI21_X2 U2896 ( .A1(n22774), .A2(n15718), .B(n22759), .ZN(n7625) );
  XOR2_X1 U2901 ( .A1(Plaintext[70]), .A2(Key[70]), .Z(n270) );
  XOR2_X1 U2917 ( .A1(n12011), .A2(n24441), .Z(n16877) );
  XOR2_X1 U2918 ( .A1(n24475), .A2(n9386), .Z(n24441) );
  NAND3_X2 U2924 ( .A1(n273), .A2(n2922), .A3(n23991), .ZN(n24664) );
  INV_X2 U2926 ( .I(n2236), .ZN(n694) );
  XOR2_X1 U2929 ( .A1(n24596), .A2(n24576), .Z(n17097) );
  INV_X2 U2936 ( .I(n23904), .ZN(n11050) );
  XOR2_X1 U2958 ( .A1(n6706), .A2(n15761), .Z(n281) );
  XOR2_X1 U2970 ( .A1(n9644), .A2(n13888), .Z(n16030) );
  INV_X2 U2983 ( .I(n292), .ZN(n547) );
  XOR2_X1 U2986 ( .A1(n16429), .A2(n293), .Z(n476) );
  NAND2_X2 U2992 ( .A1(n11961), .A2(n294), .ZN(n19951) );
  INV_X4 U2993 ( .I(n16681), .ZN(n2694) );
  NOR2_X2 U3004 ( .A1(n14659), .A2(n14658), .ZN(n14657) );
  XOR2_X1 U3008 ( .A1(n7387), .A2(n13863), .Z(n17126) );
  NAND2_X2 U3009 ( .A1(n13478), .A2(n13479), .ZN(n7387) );
  INV_X2 U3029 ( .I(n15057), .ZN(n16009) );
  INV_X4 U3032 ( .I(n17598), .ZN(n18761) );
  AND2_X1 U3044 ( .A1(n24138), .A2(n24141), .Z(n11832) );
  XOR2_X1 U3050 ( .A1(n5381), .A2(n30319), .Z(n23313) );
  XOR2_X1 U3052 ( .A1(n308), .A2(n19539), .Z(n7193) );
  XOR2_X1 U3053 ( .A1(n31568), .A2(n16301), .Z(n308) );
  INV_X4 U3065 ( .I(n21056), .ZN(n9191) );
  NAND2_X2 U3079 ( .A1(n5969), .A2(n5968), .ZN(n5970) );
  NAND2_X2 U3082 ( .A1(n10513), .A2(n24207), .ZN(n24062) );
  BUF_X2 U3100 ( .I(n24852), .Z(n322) );
  NOR2_X2 U3105 ( .A1(n14951), .A2(n16844), .ZN(n13800) );
  XOR2_X1 U3117 ( .A1(n15093), .A2(n15934), .Z(n16778) );
  XOR2_X1 U3118 ( .A1(n22114), .A2(n29851), .Z(n3101) );
  BUF_X4 U3127 ( .I(n13531), .Z(n13548) );
  NAND2_X1 U3135 ( .A1(n8305), .A2(n5595), .ZN(n329) );
  NAND2_X2 U3138 ( .A1(n10615), .A2(n10614), .ZN(n20412) );
  INV_X2 U3141 ( .I(n25228), .ZN(n25306) );
  NOR2_X2 U3144 ( .A1(n24036), .A2(n24035), .ZN(n24796) );
  OR2_X1 U3161 ( .A1(n11827), .A2(n11826), .Z(n337) );
  INV_X2 U3178 ( .I(n25711), .ZN(n1077) );
  XOR2_X1 U3183 ( .A1(n19626), .A2(n4942), .Z(n19577) );
  XOR2_X1 U3189 ( .A1(n22235), .A2(n22152), .Z(n2696) );
  XOR2_X1 U3190 ( .A1(n16210), .A2(n22017), .Z(n22235) );
  OAI22_X1 U3192 ( .A1(n18777), .A2(n28686), .B1(n954), .B2(n16585), .ZN(
        n12877) );
  INV_X1 U3200 ( .I(n8243), .ZN(n13730) );
  NAND2_X2 U3210 ( .A1(n2905), .A2(n15285), .ZN(n20632) );
  INV_X2 U3215 ( .I(n18048), .ZN(n349) );
  XOR2_X1 U3233 ( .A1(n15630), .A2(n26075), .Z(n5133) );
  NOR2_X2 U3235 ( .A1(n6943), .A2(n642), .ZN(n6874) );
  OR2_X1 U3237 ( .A1(n28338), .A2(n11899), .Z(n13819) );
  INV_X2 U3257 ( .I(n18654), .ZN(n18798) );
  INV_X2 U3264 ( .I(n5441), .ZN(n22585) );
  OAI21_X2 U3265 ( .A1(n18327), .A2(n180), .B(n9840), .ZN(n2581) );
  NAND3_X2 U3274 ( .A1(n365), .A2(n5990), .A3(n5989), .ZN(n5988) );
  OAI21_X2 U3280 ( .A1(n7330), .A2(n10460), .B(n7332), .ZN(n14522) );
  XOR2_X1 U3283 ( .A1(n10809), .A2(n367), .Z(n11969) );
  INV_X2 U3294 ( .I(n24204), .ZN(n24061) );
  INV_X4 U3297 ( .I(n8832), .ZN(n18515) );
  NOR2_X2 U3304 ( .A1(n5121), .A2(n5122), .ZN(n6846) );
  XOR2_X1 U3315 ( .A1(n1941), .A2(n1942), .Z(n7573) );
  NAND2_X2 U3321 ( .A1(n4130), .A2(n8144), .ZN(n3929) );
  XOR2_X1 U3345 ( .A1(n15367), .A2(n26057), .Z(n380) );
  INV_X2 U3351 ( .I(n627), .ZN(n1284) );
  XOR2_X1 U3361 ( .A1(n19611), .A2(n9599), .Z(n2672) );
  XOR2_X1 U3369 ( .A1(n16877), .A2(n385), .Z(n2315) );
  XOR2_X1 U3370 ( .A1(n18174), .A2(n18173), .Z(n385) );
  INV_X2 U3400 ( .I(n18037), .ZN(n17147) );
  NAND2_X2 U3405 ( .A1(n25402), .A2(n25401), .ZN(n25440) );
  AOI21_X2 U3423 ( .A1(n12026), .A2(n27455), .B(n6363), .ZN(n12434) );
  OR2_X1 U3442 ( .A1(n22439), .A2(n8409), .Z(n17008) );
  NAND2_X2 U3446 ( .A1(n25391), .A2(n17717), .ZN(n25346) );
  NAND2_X2 U3450 ( .A1(n3554), .A2(n3552), .ZN(n4746) );
  NAND3_X1 U3455 ( .A1(n12682), .A2(n20040), .A3(n20138), .ZN(n410) );
  NAND3_X1 U3463 ( .A1(n6072), .A2(n8409), .A3(n1125), .ZN(n413) );
  BUF_X2 U3467 ( .I(n26049), .Z(n414) );
  XOR2_X1 U3474 ( .A1(n10205), .A2(n10979), .Z(n5847) );
  INV_X4 U3477 ( .I(n18720), .ZN(n18855) );
  OR2_X1 U3481 ( .A1(n25366), .A2(n30400), .Z(n25371) );
  XOR2_X1 U3483 ( .A1(n3493), .A2(n416), .Z(n17932) );
  INV_X2 U3508 ( .I(n4798), .ZN(n424) );
  XOR2_X1 U3509 ( .A1(n17384), .A2(n425), .Z(n5340) );
  XOR2_X1 U3510 ( .A1(n30327), .A2(n24516), .Z(n425) );
  XOR2_X1 U3514 ( .A1(n22311), .A2(n22233), .Z(n9432) );
  XOR2_X1 U3515 ( .A1(n27130), .A2(n2863), .Z(n22311) );
  XOR2_X1 U3518 ( .A1(n19585), .A2(n10434), .Z(n2064) );
  XOR2_X1 U3526 ( .A1(n5244), .A2(n30311), .Z(n3584) );
  AOI21_X2 U3551 ( .A1(n19889), .A2(n11475), .B(n19949), .ZN(n7245) );
  XOR2_X1 U3563 ( .A1(n439), .A2(n16381), .Z(Ciphertext[7]) );
  INV_X2 U3569 ( .I(n12906), .ZN(n17373) );
  XOR2_X1 U3570 ( .A1(n12962), .A2(n440), .Z(n12960) );
  XOR2_X1 U3571 ( .A1(n11784), .A2(n26100), .Z(n440) );
  OR2_X1 U3583 ( .A1(n20376), .A2(n20361), .Z(n5351) );
  INV_X1 U3593 ( .I(n22677), .ZN(n22403) );
  XNOR2_X1 U3624 ( .A1(n19540), .A2(n1364), .ZN(n444) );
  XNOR2_X1 U3625 ( .A1(n19539), .A2(n16578), .ZN(n445) );
  XNOR2_X1 U3628 ( .A1(n20730), .A2(n25735), .ZN(n447) );
  XNOR2_X1 U3633 ( .A1(n30532), .A2(n16696), .ZN(n452) );
  XNOR2_X1 U3635 ( .A1(n34150), .A2(n16698), .ZN(n454) );
  XNOR2_X1 U3637 ( .A1(n19473), .A2(n25195), .ZN(n456) );
  XNOR2_X1 U3638 ( .A1(n31229), .A2(n1403), .ZN(n457) );
  XNOR2_X1 U3639 ( .A1(n283), .A2(n1409), .ZN(n458) );
  XNOR2_X1 U3642 ( .A1(n19691), .A2(n25108), .ZN(n461) );
  XNOR2_X1 U3644 ( .A1(n19463), .A2(n25182), .ZN(n463) );
  XNOR2_X1 U3646 ( .A1(n23475), .A2(n23474), .ZN(n465) );
  XNOR2_X1 U3652 ( .A1(n19651), .A2(n25465), .ZN(n467) );
  XNOR2_X1 U3660 ( .A1(n14132), .A2(n16674), .ZN(n474) );
  XNOR2_X1 U3661 ( .A1(n23535), .A2(n16679), .ZN(n475) );
  XNOR2_X1 U3662 ( .A1(n15517), .A2(n25098), .ZN(n477) );
  XNOR2_X1 U3663 ( .A1(n30212), .A2(n24386), .ZN(n478) );
  XNOR2_X1 U3665 ( .A1(n10294), .A2(n1197), .ZN(n480) );
  XNOR2_X1 U3666 ( .A1(n34100), .A2(n16619), .ZN(n481) );
  AND2_X2 U3670 ( .A1(n17558), .A2(n4869), .Z(n485) );
  XNOR2_X1 U3672 ( .A1(n15236), .A2(n25319), .ZN(n487) );
  XOR2_X1 U3673 ( .A1(Plaintext[34]), .A2(Key[34]), .Z(n488) );
  XOR2_X1 U3678 ( .A1(Plaintext[97]), .A2(Key[97]), .Z(n493) );
  XNOR2_X1 U3679 ( .A1(Plaintext[115]), .A2(Key[115]), .ZN(n494) );
  XOR2_X1 U3680 ( .A1(Plaintext[190]), .A2(Key[190]), .Z(n495) );
  XNOR2_X1 U3681 ( .A1(n10180), .A2(n8685), .ZN(n496) );
  XOR2_X1 U3683 ( .A1(Plaintext[96]), .A2(Key[96]), .Z(n498) );
  XNOR2_X1 U3685 ( .A1(n20963), .A2(n24065), .ZN(n500) );
  XNOR2_X1 U3689 ( .A1(n17010), .A2(n17009), .ZN(n503) );
  XNOR2_X1 U3692 ( .A1(n20813), .A2(n25693), .ZN(n506) );
  XNOR2_X1 U3693 ( .A1(n20921), .A2(n29707), .ZN(n507) );
  XNOR2_X1 U3694 ( .A1(n5414), .A2(n16654), .ZN(n508) );
  XNOR2_X1 U3697 ( .A1(n16634), .A2(n16448), .ZN(n511) );
  XNOR2_X1 U3699 ( .A1(n28762), .A2(n25001), .ZN(n513) );
  XNOR2_X1 U3700 ( .A1(n8269), .A2(n1427), .ZN(n514) );
  XNOR2_X1 U3704 ( .A1(n4285), .A2(n32130), .ZN(n518) );
  XNOR2_X1 U3707 ( .A1(n30309), .A2(n25506), .ZN(n521) );
  XNOR2_X1 U3710 ( .A1(n23475), .A2(n17400), .ZN(n524) );
  XNOR2_X1 U3713 ( .A1(n32050), .A2(n27176), .ZN(n528) );
  XNOR2_X1 U3714 ( .A1(n23196), .A2(n25648), .ZN(n529) );
  XNOR2_X1 U3715 ( .A1(n23200), .A2(n23291), .ZN(n530) );
  XNOR2_X1 U3716 ( .A1(n10535), .A2(n16504), .ZN(n531) );
  XNOR2_X1 U3717 ( .A1(n29217), .A2(n25716), .ZN(n532) );
  XNOR2_X1 U3718 ( .A1(n7046), .A2(n18019), .ZN(n533) );
  XOR2_X1 U3720 ( .A1(n10659), .A2(n11148), .Z(n535) );
  XNOR2_X1 U3721 ( .A1(n22056), .A2(n25457), .ZN(n536) );
  XNOR2_X1 U3722 ( .A1(n13844), .A2(n16381), .ZN(n537) );
  XNOR2_X1 U3723 ( .A1(n16160), .A2(n25001), .ZN(n538) );
  INV_X1 U3725 ( .I(n23931), .ZN(n23527) );
  XNOR2_X1 U3726 ( .A1(n6262), .A2(n23295), .ZN(n540) );
  XNOR2_X1 U3727 ( .A1(n22113), .A2(n3704), .ZN(n541) );
  XNOR2_X1 U3728 ( .A1(n22113), .A2(n22173), .ZN(n542) );
  XNOR2_X1 U3729 ( .A1(n25751), .A2(n27801), .ZN(n543) );
  XNOR2_X1 U3730 ( .A1(n24738), .A2(n24632), .ZN(n544) );
  XNOR2_X1 U3731 ( .A1(n24790), .A2(n25040), .ZN(n545) );
  XNOR2_X1 U3732 ( .A1(n24787), .A2(n25493), .ZN(n546) );
  XNOR2_X1 U3734 ( .A1(n14789), .A2(n25879), .ZN(n549) );
  XNOR2_X1 U3735 ( .A1(n24816), .A2(n24895), .ZN(n550) );
  XNOR2_X1 U3736 ( .A1(n23467), .A2(n13033), .ZN(n551) );
  XNOR2_X1 U3738 ( .A1(n24545), .A2(n25104), .ZN(n553) );
  XNOR2_X1 U3739 ( .A1(n25428), .A2(n24512), .ZN(n554) );
  XNOR2_X1 U3742 ( .A1(n12821), .A2(n25578), .ZN(n556) );
  XNOR2_X1 U3755 ( .A1(n9044), .A2(n6254), .ZN(n567) );
  XNOR2_X1 U3759 ( .A1(n10663), .A2(n10661), .ZN(n571) );
  XOR2_X1 U3764 ( .A1(n7636), .A2(n7634), .Z(n576) );
  BUF_X2 U3769 ( .I(n11910), .Z(n11350) );
  INV_X2 U3775 ( .I(n20117), .ZN(n20045) );
  XOR2_X1 U3782 ( .A1(n32478), .A2(n16705), .Z(n586) );
  XNOR2_X1 U3789 ( .A1(n20242), .A2(n20241), .ZN(n590) );
  XNOR2_X1 U3790 ( .A1(n20873), .A2(n25878), .ZN(n591) );
  XNOR2_X1 U3795 ( .A1(n18095), .A2(n16820), .ZN(n595) );
  XNOR2_X1 U3800 ( .A1(n8827), .A2(n8826), .ZN(n598) );
  INV_X2 U3803 ( .I(n8632), .ZN(n21149) );
  XNOR2_X1 U3804 ( .A1(n20699), .A2(n20698), .ZN(n600) );
  XOR2_X1 U3805 ( .A1(n1487), .A2(n2009), .Z(n601) );
  XNOR2_X1 U3807 ( .A1(n10164), .A2(n20390), .ZN(n603) );
  INV_X2 U3810 ( .I(n20468), .ZN(n3462) );
  NAND2_X2 U3817 ( .A1(n4785), .A2(n4784), .ZN(n21466) );
  XNOR2_X1 U3819 ( .A1(n15268), .A2(n20644), .ZN(n609) );
  NAND3_X2 U3826 ( .A1(n1651), .A2(n1649), .A3(n1648), .ZN(n22012) );
  XNOR2_X1 U3827 ( .A1(n22145), .A2(n25167), .ZN(n612) );
  XNOR2_X1 U3828 ( .A1(n18189), .A2(n24999), .ZN(n613) );
  XNOR2_X1 U3834 ( .A1(n22047), .A2(n22013), .ZN(n618) );
  XNOR2_X1 U3837 ( .A1(n22140), .A2(n22142), .ZN(n620) );
  XNOR2_X1 U3840 ( .A1(n22029), .A2(n22021), .ZN(n623) );
  XNOR2_X1 U3841 ( .A1(n5476), .A2(n31094), .ZN(n624) );
  NAND2_X2 U3852 ( .A1(n12845), .A2(n14878), .ZN(n12594) );
  NOR2_X2 U3858 ( .A1(n14044), .A2(n14765), .ZN(n22957) );
  NAND2_X2 U3867 ( .A1(n15608), .A2(n15607), .ZN(n12729) );
  XNOR2_X1 U3874 ( .A1(n14036), .A2(n9228), .ZN(n647) );
  XOR2_X1 U3884 ( .A1(n23304), .A2(n10129), .Z(n657) );
  XNOR2_X1 U3890 ( .A1(n11551), .A2(n23468), .ZN(n660) );
  XOR2_X1 U3891 ( .A1(n11039), .A2(n23077), .Z(n661) );
  NAND2_X2 U3900 ( .A1(n9343), .A2(n23671), .ZN(n9342) );
  OAI21_X2 U3904 ( .A1(n17730), .A2(n11975), .B(n13603), .ZN(n24275) );
  INV_X2 U3919 ( .I(n4951), .ZN(n17861) );
  INV_X4 U3923 ( .I(n25871), .ZN(n883) );
  INV_X2 U3942 ( .I(n17476), .ZN(n25903) );
  INV_X2 U3944 ( .I(n8044), .ZN(n25892) );
  OR2_X1 U3947 ( .A1(n25067), .A2(n1951), .Z(n693) );
  OR2_X1 U3949 ( .A1(n24922), .A2(n15799), .Z(n698) );
  NAND2_X2 U3965 ( .A1(n4420), .A2(n15350), .ZN(n20450) );
  AOI21_X2 U3970 ( .A1(n28395), .A2(n28838), .B(n2551), .ZN(n1771) );
  INV_X1 U3978 ( .I(n19583), .ZN(n16110) );
  NAND3_X2 U3988 ( .A1(n17511), .A2(n20490), .A3(n17513), .ZN(n20726) );
  OAI21_X2 U3997 ( .A1(n10167), .A2(n17269), .B(n10166), .ZN(n23053) );
  INV_X1 U4012 ( .I(n22390), .ZN(n22549) );
  AOI21_X2 U4021 ( .A1(n5473), .A2(n5053), .B(n5052), .ZN(n16047) );
  AOI21_X2 U4034 ( .A1(n12634), .A2(n20135), .B(n19964), .ZN(n2905) );
  NAND2_X1 U4039 ( .A1(n6288), .A2(n7842), .ZN(n25679) );
  OR2_X1 U4043 ( .A1(n24910), .A2(n10755), .Z(n8304) );
  NAND2_X2 U4050 ( .A1(n25765), .A2(n25704), .ZN(n9804) );
  AOI21_X2 U4051 ( .A1(n17475), .A2(n25904), .B(n8299), .ZN(n10285) );
  INV_X2 U4074 ( .I(n14142), .ZN(n25563) );
  INV_X2 U4101 ( .I(n7825), .ZN(n15423) );
  INV_X2 U4109 ( .I(n2200), .ZN(n23201) );
  INV_X2 U4144 ( .I(n9753), .ZN(n10622) );
  INV_X2 U4146 ( .I(n9750), .ZN(n10568) );
  INV_X2 U4154 ( .I(n8964), .ZN(n8965) );
  INV_X1 U4179 ( .I(n28429), .ZN(n12278) );
  NAND2_X2 U4213 ( .A1(n11141), .A2(n5910), .ZN(n17544) );
  NAND2_X2 U4214 ( .A1(n9099), .A2(n9098), .ZN(n12563) );
  INV_X2 U4221 ( .I(n29252), .ZN(n821) );
  BUF_X4 U4226 ( .I(n19455), .Z(n16694) );
  INV_X2 U4229 ( .I(n12467), .ZN(n20067) );
  AND2_X1 U4237 ( .A1(n13252), .A2(n1452), .Z(n1451) );
  AND2_X1 U4255 ( .A1(n15873), .A2(n5834), .Z(n15870) );
  INV_X2 U4262 ( .I(n3954), .ZN(n5225) );
  CLKBUF_X2 U4270 ( .I(n18823), .Z(n4868) );
  BUF_X1 U4272 ( .I(Key[133]), .Z(n25156) );
  BUF_X1 U4275 ( .I(Key[105]), .Z(n16506) );
  BUF_X1 U4286 ( .I(Key[189]), .Z(n24527) );
  BUF_X1 U4291 ( .I(Key[168]), .Z(n25086) );
  BUF_X1 U4293 ( .I(Key[161]), .Z(n25288) );
  BUF_X1 U4299 ( .I(Key[59]), .Z(n24231) );
  BUF_X1 U4304 ( .I(Key[135]), .Z(n24417) );
  BUF_X1 U4308 ( .I(Key[9]), .Z(n25570) );
  BUF_X1 U4312 ( .I(Key[165]), .Z(n16597) );
  BUF_X1 U4314 ( .I(Key[125]), .Z(n25108) );
  BUF_X1 U4315 ( .I(Key[104]), .Z(n24514) );
  BUF_X1 U4320 ( .I(Key[131]), .Z(n24426) );
  NAND3_X1 U4333 ( .A1(n25575), .A2(n25571), .A3(n30285), .ZN(n6730) );
  NAND3_X1 U4339 ( .A1(n25916), .A2(n25915), .A3(n25925), .ZN(n25917) );
  NAND2_X1 U4341 ( .A1(n25851), .A2(n13049), .ZN(n13953) );
  NAND2_X1 U4344 ( .A1(n24904), .A2(n24915), .ZN(n3820) );
  AOI21_X1 U4347 ( .A1(n15054), .A2(n25258), .B(n2191), .ZN(n25246) );
  INV_X1 U4359 ( .I(n25687), .ZN(n7843) );
  INV_X1 U4361 ( .I(n3229), .ZN(n3230) );
  NAND3_X1 U4363 ( .A1(n27113), .A2(n5926), .A3(n25571), .ZN(n25573) );
  NAND2_X1 U4366 ( .A1(n31178), .A2(n25313), .ZN(n25314) );
  AOI22_X1 U4384 ( .A1(n700), .A2(n14104), .B1(n10136), .B2(n25900), .ZN(
        n17195) );
  NAND2_X1 U4398 ( .A1(n12856), .A2(n25591), .ZN(n1751) );
  NAND2_X1 U4404 ( .A1(n24725), .A2(n25871), .ZN(n9110) );
  OAI21_X1 U4408 ( .A1(n12359), .A2(n12358), .B(n3828), .ZN(n5763) );
  AND2_X1 U4411 ( .A1(n18219), .A2(n10062), .Z(n10221) );
  NAND2_X1 U4431 ( .A1(n28096), .A2(n15295), .ZN(n9718) );
  INV_X1 U4445 ( .I(n25111), .ZN(n9506) );
  NAND4_X1 U4463 ( .A1(n1816), .A2(n1818), .A3(n1819), .A4(n23594), .ZN(n7962)
         );
  NAND2_X1 U4486 ( .A1(n23581), .A2(n29068), .ZN(n23582) );
  NAND3_X2 U4499 ( .A1(n22410), .A2(n9747), .A3(n17481), .ZN(n6386) );
  NAND2_X1 U4532 ( .A1(n22550), .A2(n22551), .ZN(n6366) );
  NAND2_X1 U4536 ( .A1(n22025), .A2(n628), .ZN(n11378) );
  INV_X2 U4538 ( .I(n8167), .ZN(n9737) );
  INV_X2 U4542 ( .I(n16136), .ZN(n996) );
  NOR3_X1 U4551 ( .A1(n14949), .A2(n11755), .A3(n11229), .ZN(n11228) );
  AND2_X1 U4552 ( .A1(n11755), .A2(n6442), .Z(n21676) );
  NAND2_X2 U4562 ( .A1(n6014), .A2(n6013), .ZN(n16077) );
  NOR2_X1 U4572 ( .A1(n5822), .A2(n16633), .ZN(n21311) );
  NAND3_X1 U4578 ( .A1(n14682), .A2(n10523), .A3(n20173), .ZN(n2647) );
  NOR2_X1 U4580 ( .A1(n20547), .A2(n30130), .ZN(n1961) );
  NOR2_X1 U4585 ( .A1(n20548), .A2(n710), .ZN(n6134) );
  NAND2_X1 U4591 ( .A1(n1964), .A2(n26182), .ZN(n1963) );
  INV_X1 U4595 ( .I(n20503), .ZN(n16146) );
  INV_X2 U4611 ( .I(n8373), .ZN(n8857) );
  INV_X2 U4612 ( .I(n11507), .ZN(n14761) );
  INV_X1 U4615 ( .I(n7575), .ZN(n7008) );
  INV_X2 U4643 ( .I(n15216), .ZN(n18307) );
  INV_X2 U4646 ( .I(n6265), .ZN(n15216) );
  BUF_X1 U4648 ( .I(Key[103]), .Z(n16701) );
  NAND3_X1 U4659 ( .A1(n1208), .A2(n24969), .A3(n24970), .ZN(n1934) );
  NAND2_X1 U4664 ( .A1(n10755), .A2(n24910), .ZN(n9991) );
  INV_X1 U4670 ( .I(n3843), .ZN(n12783) );
  INV_X1 U4677 ( .I(n32855), .ZN(n25613) );
  INV_X1 U4681 ( .I(n27173), .ZN(n2049) );
  NAND2_X1 U4700 ( .A1(n14267), .A2(n25890), .ZN(n12678) );
  NAND2_X1 U4704 ( .A1(n25233), .A2(n25232), .ZN(n17925) );
  NOR2_X1 U4720 ( .A1(n17535), .A2(n31920), .ZN(n4491) );
  AOI21_X1 U4726 ( .A1(n25229), .A2(n25306), .B(n18059), .ZN(n9428) );
  INV_X1 U4732 ( .I(n2378), .ZN(n25526) );
  INV_X2 U4736 ( .I(n686), .ZN(n13763) );
  INV_X2 U4741 ( .I(n30277), .ZN(n837) );
  INV_X1 U4749 ( .I(n10048), .ZN(n7602) );
  NAND2_X1 U4760 ( .A1(n9178), .A2(n10687), .ZN(n11788) );
  AOI21_X1 U4766 ( .A1(n27159), .A2(n26750), .B(n24106), .ZN(n13237) );
  NAND2_X1 U4769 ( .A1(n10687), .A2(n32737), .ZN(n15158) );
  NOR2_X1 U4787 ( .A1(n6474), .A2(n14078), .ZN(n9812) );
  INV_X1 U4803 ( .I(n17285), .ZN(n23708) );
  INV_X1 U4811 ( .I(n17857), .ZN(n23857) );
  INV_X1 U4812 ( .I(n23287), .ZN(n23242) );
  INV_X1 U4815 ( .I(n3600), .ZN(n4777) );
  NAND2_X1 U4819 ( .A1(n3773), .A2(n22977), .ZN(n2624) );
  INV_X1 U4833 ( .I(n9335), .ZN(n9334) );
  INV_X1 U4865 ( .I(n19894), .ZN(n20417) );
  INV_X1 U4867 ( .I(n20595), .ZN(n20499) );
  INV_X2 U4879 ( .I(n571), .ZN(n14559) );
  AOI21_X1 U4894 ( .A1(n18835), .A2(n13846), .B(n18832), .ZN(n14393) );
  AOI22_X1 U4917 ( .A1(n12783), .A2(n24969), .B1(n8622), .B2(n27134), .ZN(
        n3136) );
  AOI21_X1 U4953 ( .A1(n25637), .A2(n9718), .B(n27188), .ZN(n9717) );
  OR2_X1 U4954 ( .A1(n25876), .A2(n1211), .Z(n3955) );
  NAND3_X1 U4959 ( .A1(n14630), .A2(n17595), .A3(n14629), .ZN(n14628) );
  AOI21_X1 U4963 ( .A1(n17169), .A2(n24606), .B(n9941), .ZN(n24025) );
  NOR2_X1 U4977 ( .A1(n1083), .A2(n34115), .ZN(n8840) );
  AOI21_X1 U4995 ( .A1(n9202), .A2(n970), .B(n9275), .ZN(n9366) );
  NAND2_X1 U5022 ( .A1(n23715), .A2(n707), .ZN(n6248) );
  INV_X1 U5045 ( .I(n11621), .ZN(n4111) );
  NAND2_X1 U5076 ( .A1(n2418), .A2(n22567), .ZN(n22444) );
  NAND2_X1 U5095 ( .A1(n12794), .A2(n34046), .ZN(n21576) );
  INV_X1 U5102 ( .I(n7753), .ZN(n21752) );
  INV_X1 U5122 ( .I(n20650), .ZN(n20270) );
  NOR2_X1 U5161 ( .A1(n12316), .A2(n18993), .ZN(n1453) );
  NAND2_X1 U5175 ( .A1(n5328), .A2(n5327), .ZN(n4053) );
  NAND3_X1 U5180 ( .A1(n17073), .A2(n10786), .A3(n29659), .ZN(n10785) );
  INV_X1 U5181 ( .I(n5328), .ZN(n4178) );
  NOR2_X1 U5186 ( .A1(n493), .A2(n16450), .ZN(n5753) );
  NAND4_X1 U5194 ( .A1(n5622), .A2(n25206), .A3(n5621), .A4(n7304), .ZN(n7302)
         );
  NAND3_X1 U5195 ( .A1(n4770), .A2(n4781), .A3(n10858), .ZN(n4769) );
  NOR2_X1 U5200 ( .A1(n4781), .A2(n9247), .ZN(n3988) );
  NOR2_X1 U5221 ( .A1(n24484), .A2(n17684), .ZN(n6365) );
  INV_X1 U5230 ( .I(n11409), .ZN(n25263) );
  NAND2_X1 U5234 ( .A1(n15555), .A2(n25870), .ZN(n15670) );
  INV_X2 U5236 ( .I(n17861), .ZN(n25292) );
  INV_X2 U5240 ( .I(n15295), .ZN(n13032) );
  INV_X1 U5241 ( .I(n1786), .ZN(n25203) );
  INV_X1 U5242 ( .I(n17092), .ZN(n15355) );
  NOR2_X1 U5249 ( .A1(n25564), .A2(n25582), .ZN(n25634) );
  NAND2_X1 U5290 ( .A1(n707), .A2(n8370), .ZN(n7190) );
  NAND2_X1 U5295 ( .A1(n23816), .A2(n17616), .ZN(n17816) );
  NAND2_X1 U5301 ( .A1(n23949), .A2(n11621), .ZN(n9894) );
  NAND2_X1 U5303 ( .A1(n15865), .A2(n27136), .ZN(n23555) );
  OAI21_X1 U5304 ( .A1(n3553), .A2(n11621), .B(n30360), .ZN(n3552) );
  INV_X1 U5309 ( .I(n16536), .ZN(n23713) );
  AND2_X1 U5311 ( .A1(n34009), .A2(n28914), .Z(n8850) );
  OAI21_X1 U5315 ( .A1(n847), .A2(n8760), .B(n23721), .ZN(n23115) );
  INV_X1 U5324 ( .I(n11887), .ZN(n7088) );
  INV_X2 U5328 ( .I(n17591), .ZN(n23888) );
  INV_X1 U5329 ( .I(n26114), .ZN(n16097) );
  INV_X2 U5331 ( .I(n9798), .ZN(n11943) );
  INV_X2 U5335 ( .I(n23286), .ZN(n770) );
  NAND3_X1 U5337 ( .A1(n10528), .A2(n28891), .A3(n1271), .ZN(n17774) );
  NOR2_X1 U5375 ( .A1(n22608), .A2(n32512), .ZN(n7426) );
  NAND2_X1 U5378 ( .A1(n22535), .A2(n22428), .ZN(n22540) );
  INV_X1 U5433 ( .I(n17746), .ZN(n15468) );
  NAND3_X1 U5443 ( .A1(n6405), .A2(n13451), .A3(n32746), .ZN(n13301) );
  INV_X1 U5471 ( .I(n13450), .ZN(n19051) );
  OAI21_X1 U5476 ( .A1(n12707), .A2(n19048), .B(n28705), .ZN(n12600) );
  NAND2_X1 U5482 ( .A1(n5545), .A2(n5889), .ZN(n5907) );
  NAND2_X1 U5508 ( .A1(n13360), .A2(n8208), .ZN(n17073) );
  INV_X1 U5509 ( .I(n3344), .ZN(n18311) );
  INV_X1 U5516 ( .I(n13531), .ZN(n1063) );
  NAND2_X1 U5536 ( .A1(n830), .A2(n27123), .ZN(n3706) );
  NAND3_X1 U5542 ( .A1(n715), .A2(n25220), .A3(n25210), .ZN(n7304) );
  INV_X1 U5545 ( .I(n31236), .ZN(n25550) );
  INV_X1 U5555 ( .I(n25746), .ZN(n832) );
  AOI22_X1 U5559 ( .A1(n4492), .A2(n31920), .B1(n4407), .B2(n4491), .ZN(n5886)
         );
  AND2_X1 U5566 ( .A1(n833), .A2(n24667), .Z(n25537) );
  NAND2_X1 U5573 ( .A1(n13985), .A2(n25261), .ZN(n24581) );
  AND2_X1 U5576 ( .A1(n25334), .A2(n25536), .Z(n12088) );
  NOR2_X1 U5578 ( .A1(n317), .A2(n6551), .ZN(n6640) );
  AOI21_X1 U5580 ( .A1(n15235), .A2(n33393), .B(n765), .ZN(n5929) );
  NAND3_X1 U5581 ( .A1(n10497), .A2(n15295), .A3(n2378), .ZN(n25715) );
  AOI22_X1 U5582 ( .A1(n15235), .A2(n25561), .B1(n765), .B2(n16704), .ZN(n5930) );
  AND2_X1 U5591 ( .A1(n25586), .A2(n25590), .Z(n12423) );
  NAND2_X1 U5592 ( .A1(n678), .A2(n25409), .ZN(n25326) );
  INV_X1 U5599 ( .I(n25115), .ZN(n16025) );
  INV_X1 U5613 ( .I(n24763), .ZN(n1225) );
  NAND2_X1 U5625 ( .A1(n24156), .A2(n10513), .ZN(n9283) );
  NAND3_X1 U5627 ( .A1(n7150), .A2(n16868), .A3(n24253), .ZN(n3546) );
  AND2_X1 U5640 ( .A1(n24061), .A2(n24156), .Z(n2463) );
  NAND3_X1 U5641 ( .A1(n767), .A2(n29566), .A3(n2847), .ZN(n7094) );
  NAND3_X1 U5700 ( .A1(n23867), .A2(n17895), .A3(n23868), .ZN(n23821) );
  NAND3_X1 U5701 ( .A1(n8408), .A2(n23868), .A3(n1257), .ZN(n10132) );
  NAND2_X1 U5717 ( .A1(n23947), .A2(n4111), .ZN(n1525) );
  INV_X1 U5735 ( .I(n23346), .ZN(n23132) );
  AND3_X1 U5746 ( .A1(n4067), .A2(n22826), .A3(n30437), .Z(n22652) );
  OAI21_X1 U5766 ( .A1(n6593), .A2(n17720), .B(n22955), .ZN(n2002) );
  INV_X1 U5777 ( .I(n17890), .ZN(n22389) );
  NAND3_X1 U5788 ( .A1(n902), .A2(n22330), .A3(n14376), .ZN(n11008) );
  INV_X1 U5795 ( .I(n29451), .ZN(n14008) );
  INV_X1 U5801 ( .I(n22576), .ZN(n16148) );
  OAI21_X1 U5815 ( .A1(n21123), .A2(n31910), .B(n31260), .ZN(n21126) );
  INV_X2 U5838 ( .I(n21432), .ZN(n5049) );
  AOI21_X1 U5840 ( .A1(n21453), .A2(n9186), .B(n780), .ZN(n9393) );
  NOR2_X1 U5841 ( .A1(n11966), .A2(n21367), .ZN(n2605) );
  INV_X1 U5847 ( .I(n8398), .ZN(n3931) );
  OAI21_X1 U5862 ( .A1(n26182), .A2(n20545), .B(n3157), .ZN(n13631) );
  OAI21_X1 U5870 ( .A1(n2566), .A2(n17497), .B(n8293), .ZN(n19955) );
  NAND4_X1 U5875 ( .A1(n1678), .A2(n1680), .A3(n1677), .A4(n1679), .ZN(n20306)
         );
  OAI21_X1 U5886 ( .A1(n10286), .A2(n18142), .B(n14306), .ZN(n3945) );
  NOR2_X1 U5901 ( .A1(n13605), .A2(n20088), .ZN(n11501) );
  INV_X2 U5907 ( .I(n4881), .ZN(n6275) );
  AND2_X1 U5908 ( .A1(n16489), .A2(n20052), .Z(n16675) );
  INV_X1 U5916 ( .I(n11910), .ZN(n19863) );
  NAND2_X1 U5944 ( .A1(n27726), .A2(n3388), .ZN(n3390) );
  OAI21_X1 U5959 ( .A1(n15495), .A2(n9937), .B(n16538), .ZN(n15576) );
  OR2_X2 U5962 ( .A1(n18709), .A2(n17625), .Z(n10700) );
  NOR2_X1 U5964 ( .A1(n15902), .A2(n1709), .ZN(n9937) );
  NOR2_X1 U5974 ( .A1(n13548), .A2(n15146), .ZN(n13526) );
  INV_X1 U5997 ( .I(n17189), .ZN(n881) );
  INV_X2 U5999 ( .I(n18559), .ZN(n828) );
  CLKBUF_X2 U6002 ( .I(Key[58]), .Z(n16691) );
  CLKBUF_X2 U6004 ( .I(Key[187]), .Z(n16655) );
  CLKBUF_X2 U6006 ( .I(Key[91]), .Z(n24869) );
  CLKBUF_X2 U6007 ( .I(Key[79]), .Z(n16555) );
  CLKBUF_X2 U6010 ( .I(Key[151]), .Z(n16654) );
  NOR2_X1 U6015 ( .A1(n17927), .A2(n27123), .ZN(n9703) );
  AOI21_X1 U6020 ( .A1(n714), .A2(n25007), .B(n3232), .ZN(n3231) );
  OAI21_X1 U6021 ( .A1(n1076), .A2(n10376), .B(n25724), .ZN(n4253) );
  AND2_X1 U6022 ( .A1(n27123), .A2(n786), .Z(n12060) );
  NOR2_X1 U6023 ( .A1(n27123), .A2(n9247), .ZN(n3435) );
  OR2_X1 U6025 ( .A1(n4415), .A2(n25744), .Z(n24432) );
  INV_X1 U6027 ( .I(n32859), .ZN(n25105) );
  NAND2_X1 U6029 ( .A1(n28358), .A2(n16509), .ZN(n25216) );
  NOR2_X1 U6030 ( .A1(n5926), .A2(n5942), .ZN(n5918) );
  INV_X2 U6042 ( .I(n16509), .ZN(n15340) );
  INV_X1 U6053 ( .I(n25200), .ZN(n17005) );
  NOR2_X1 U6055 ( .A1(n27651), .A2(n16025), .ZN(n12165) );
  OAI21_X1 U6056 ( .A1(n25134), .A2(n5611), .B(n16589), .ZN(n25135) );
  NOR2_X1 U6057 ( .A1(n25117), .A2(n14495), .ZN(n9956) );
  INV_X1 U6058 ( .I(n24724), .ZN(n7963) );
  NOR2_X1 U6059 ( .A1(n14495), .A2(n27651), .ZN(n8608) );
  AND2_X1 U6065 ( .A1(n25884), .A2(n15152), .Z(n25886) );
  NOR2_X1 U6068 ( .A1(n25229), .A2(n13985), .ZN(n9427) );
  INV_X1 U6080 ( .I(n25977), .ZN(n1224) );
  NAND2_X1 U6104 ( .A1(n7361), .A2(n8399), .ZN(n13632) );
  AND2_X1 U6112 ( .A1(n7060), .A2(n16643), .Z(n7059) );
  NOR2_X1 U6128 ( .A1(n17178), .A2(n17180), .ZN(n16663) );
  NAND2_X1 U6129 ( .A1(n24177), .A2(n4897), .ZN(n5041) );
  NOR2_X1 U6153 ( .A1(n28222), .A2(n23754), .ZN(n23347) );
  OAI21_X1 U6160 ( .A1(n6869), .A2(n23917), .B(n8372), .ZN(n23116) );
  AND2_X1 U6181 ( .A1(n29272), .A2(n756), .Z(n7710) );
  NAND2_X1 U6198 ( .A1(n17895), .A2(n657), .ZN(n3650) );
  NOR2_X1 U6207 ( .A1(n16431), .A2(n29270), .ZN(n23643) );
  NAND2_X1 U6209 ( .A1(n1099), .A2(n29323), .ZN(n12817) );
  INV_X2 U6216 ( .I(n17506), .ZN(n843) );
  OR2_X1 U6238 ( .A1(n22868), .A2(n25994), .Z(n7103) );
  NAND2_X1 U6253 ( .A1(n12729), .A2(n16458), .ZN(n12726) );
  INV_X1 U6256 ( .I(n27719), .ZN(n11565) );
  NAND3_X1 U6263 ( .A1(n23066), .A2(n4734), .A3(n13807), .ZN(n10411) );
  NAND3_X1 U6265 ( .A1(n805), .A2(n2479), .A3(n31795), .ZN(n7582) );
  NAND3_X1 U6266 ( .A1(n1109), .A2(n31129), .A3(n22798), .ZN(n17481) );
  AND2_X1 U6308 ( .A1(n22430), .A2(n2538), .Z(n2537) );
  AND2_X1 U6309 ( .A1(n16529), .A2(n9515), .Z(n9516) );
  NAND3_X1 U6310 ( .A1(n14008), .A2(n809), .A3(n16483), .ZN(n14066) );
  NAND2_X1 U6324 ( .A1(n22575), .A2(n5743), .ZN(n5744) );
  OAI21_X1 U6330 ( .A1(n14251), .A2(n32830), .B(n14253), .ZN(n1663) );
  NAND2_X1 U6351 ( .A1(n11629), .A2(n22486), .ZN(n8318) );
  INV_X1 U6354 ( .I(n29868), .ZN(n22359) );
  NOR2_X1 U6370 ( .A1(n13167), .A2(n2801), .ZN(n7017) );
  NOR2_X1 U6428 ( .A1(n21074), .A2(n21434), .ZN(n14951) );
  OR2_X1 U6438 ( .A1(n12441), .A2(n21353), .Z(n12465) );
  NOR2_X1 U6441 ( .A1(n11272), .A2(n21095), .ZN(n7512) );
  AND3_X1 U6455 ( .A1(n10599), .A2(n21239), .A3(n5822), .Z(n13100) );
  INV_X1 U6470 ( .I(n20730), .ZN(n20824) );
  OR3_X1 U6501 ( .A1(n6679), .A2(n1357), .A3(n20635), .Z(n6616) );
  OR2_X1 U6506 ( .A1(n13282), .A2(n28836), .Z(n12115) );
  INV_X1 U6513 ( .I(n20605), .ZN(n20130) );
  OAI21_X1 U6517 ( .A1(n8100), .A2(n29253), .B(n19850), .ZN(n19234) );
  NAND3_X1 U6520 ( .A1(n12253), .A2(n18119), .A3(n1168), .ZN(n4854) );
  NOR2_X1 U6533 ( .A1(n1172), .A2(n31161), .ZN(n3311) );
  NAND2_X1 U6535 ( .A1(n16848), .A2(n29153), .ZN(n6960) );
  NAND3_X1 U6537 ( .A1(n15665), .A2(n4180), .A3(n20056), .ZN(n15313) );
  OR2_X1 U6539 ( .A1(n19456), .A2(n28293), .Z(n19994) );
  NAND3_X1 U6543 ( .A1(n4215), .A2(n33419), .A3(n20156), .ZN(n8589) );
  INV_X1 U6548 ( .I(n19936), .ZN(n14172) );
  INV_X2 U6551 ( .I(n29254), .ZN(n1168) );
  INV_X1 U6570 ( .I(n15786), .ZN(n19524) );
  NAND3_X1 U6580 ( .A1(n3822), .A2(n19016), .A3(n19017), .ZN(n4985) );
  AOI21_X1 U6585 ( .A1(n16669), .A2(n18838), .B(n13925), .ZN(n18839) );
  AND2_X1 U6589 ( .A1(n19183), .A2(n2612), .Z(n7568) );
  NAND3_X1 U6598 ( .A1(n28379), .A2(n16740), .A3(n19140), .ZN(n5333) );
  AND2_X1 U6611 ( .A1(n10423), .A2(n29781), .Z(n2149) );
  OAI21_X1 U6633 ( .A1(n15018), .A2(n8376), .B(n9886), .ZN(n3023) );
  NAND3_X1 U6637 ( .A1(n952), .A2(n711), .A3(n29315), .ZN(n10306) );
  NAND2_X1 U6647 ( .A1(n15902), .A2(n11459), .ZN(n10133) );
  NAND2_X1 U6653 ( .A1(n18480), .A2(n18605), .ZN(n16763) );
  NOR2_X1 U6657 ( .A1(n6783), .A2(n11389), .ZN(n14843) );
  NOR2_X1 U6661 ( .A1(n18682), .A2(n1659), .ZN(n12051) );
  NAND2_X1 U6677 ( .A1(n4677), .A2(n33621), .ZN(n6777) );
  NAND2_X1 U6680 ( .A1(n4808), .A2(n962), .ZN(n11389) );
  OR2_X2 U6697 ( .A1(n16855), .A2(n7216), .Z(n3779) );
  NAND2_X1 U6699 ( .A1(n6783), .A2(n14926), .ZN(n6887) );
  NAND2_X1 U6702 ( .A1(n493), .A2(n498), .ZN(n17557) );
  NOR2_X1 U6704 ( .A1(n9766), .A2(n16420), .ZN(n15697) );
  NAND2_X1 U6708 ( .A1(n16855), .A2(n7216), .ZN(n14906) );
  AND2_X1 U6714 ( .A1(n17223), .A2(n16948), .Z(n8948) );
  BUF_X2 U6719 ( .I(n16450), .Z(n5473) );
  INV_X1 U6720 ( .I(n25578), .ZN(n960) );
  CLKBUF_X2 U6723 ( .I(Key[82]), .Z(n16642) );
  CLKBUF_X2 U6725 ( .I(Key[87]), .Z(n25465) );
  CLKBUF_X2 U6726 ( .I(Key[80]), .Z(n25720) );
  INV_X2 U6728 ( .I(n18085), .ZN(n882) );
  CLKBUF_X2 U6729 ( .I(Key[14]), .Z(n25880) );
  NOR2_X1 U6736 ( .A1(n12431), .A2(n25271), .ZN(n10605) );
  NAND2_X1 U6737 ( .A1(n25571), .A2(n5942), .ZN(n3638) );
  AND2_X1 U6739 ( .A1(n5043), .A2(n15340), .Z(n4613) );
  NAND2_X1 U6740 ( .A1(n3646), .A2(n2191), .ZN(n25256) );
  NOR2_X1 U6743 ( .A1(n28736), .A2(n25128), .ZN(n6828) );
  NOR2_X1 U6745 ( .A1(n31456), .A2(n30241), .ZN(n14873) );
  NOR2_X1 U6758 ( .A1(n10097), .A2(n967), .ZN(n8247) );
  OAI21_X1 U6763 ( .A1(n25202), .A2(n16632), .B(n25203), .ZN(n3385) );
  INV_X1 U6770 ( .I(n16783), .ZN(n6641) );
  OR2_X1 U6772 ( .A1(n15425), .A2(n29063), .Z(n14925) );
  AND2_X1 U6775 ( .A1(n12039), .A2(n6034), .Z(n6825) );
  NAND2_X1 U6783 ( .A1(n11049), .A2(n16066), .ZN(n3212) );
  NAND2_X1 U6790 ( .A1(n8058), .A2(n24094), .ZN(n23382) );
  NOR2_X1 U6794 ( .A1(n7097), .A2(n7361), .ZN(n7100) );
  OAI21_X1 U6801 ( .A1(n32520), .A2(n23995), .B(n15175), .ZN(n9659) );
  AOI21_X1 U6804 ( .A1(n10987), .A2(n24328), .B(n24245), .ZN(n7097) );
  OAI21_X1 U6811 ( .A1(n24210), .A2(n24212), .B(n24211), .ZN(n6840) );
  NAND2_X1 U6815 ( .A1(n24132), .A2(n32102), .ZN(n8336) );
  NOR2_X1 U6816 ( .A1(n4024), .A2(n7503), .ZN(n24202) );
  NAND3_X1 U6817 ( .A1(n24097), .A2(n840), .A3(n26516), .ZN(n24038) );
  NAND2_X1 U6820 ( .A1(n24092), .A2(n17261), .ZN(n5914) );
  NAND2_X1 U6833 ( .A1(n23347), .A2(n28297), .ZN(n14118) );
  INV_X1 U6841 ( .I(n31096), .ZN(n14891) );
  NOR2_X1 U6871 ( .A1(n23848), .A2(n15423), .ZN(n6132) );
  NOR2_X1 U6885 ( .A1(n23872), .A2(n23695), .ZN(n23577) );
  NOR2_X1 U6892 ( .A1(n13308), .A2(n23949), .ZN(n3553) );
  NAND2_X1 U6910 ( .A1(n2623), .A2(n30573), .ZN(n11669) );
  NOR2_X1 U6931 ( .A1(n8954), .A2(n13751), .ZN(n8953) );
  INV_X1 U6934 ( .I(n22862), .ZN(n9435) );
  OAI21_X1 U6935 ( .A1(n10644), .A2(n849), .B(n10411), .ZN(n10410) );
  OR2_X1 U6938 ( .A1(n28314), .A2(n22810), .Z(n15730) );
  NOR2_X1 U6953 ( .A1(n12727), .A2(n851), .ZN(n5982) );
  AND2_X1 U6954 ( .A1(n23096), .A2(n25979), .Z(n3173) );
  NAND2_X1 U6966 ( .A1(n13694), .A2(n5915), .ZN(n4182) );
  INV_X1 U6967 ( .I(n23111), .ZN(n17099) );
  OAI21_X1 U6969 ( .A1(n13008), .A2(n29335), .B(n12688), .ZN(n12687) );
  NAND2_X1 U6977 ( .A1(n10388), .A2(n22681), .ZN(n10387) );
  NOR2_X1 U6986 ( .A1(n15260), .A2(n30668), .ZN(n7659) );
  INV_X1 U7001 ( .I(n22393), .ZN(n7490) );
  NOR2_X1 U7007 ( .A1(n27402), .A2(n22550), .ZN(n8098) );
  NOR2_X1 U7009 ( .A1(n26878), .A2(n29078), .ZN(n1519) );
  AOI21_X1 U7014 ( .A1(n628), .A2(n9234), .B(n9757), .ZN(n15643) );
  NOR2_X1 U7036 ( .A1(n22595), .A2(n22599), .ZN(n4055) );
  INV_X1 U7037 ( .I(n1289), .ZN(n11244) );
  INV_X2 U7046 ( .I(n17899), .ZN(n907) );
  INV_X1 U7047 ( .I(n22078), .ZN(n11859) );
  AOI22_X1 U7064 ( .A1(n534), .A2(n31765), .B1(n28450), .B2(n3821), .ZN(n10874) );
  NOR2_X1 U7081 ( .A1(n21856), .A2(n21), .ZN(n1595) );
  NOR2_X1 U7082 ( .A1(n30885), .A2(n1013), .ZN(n4435) );
  NOR2_X1 U7085 ( .A1(n27178), .A2(n21719), .ZN(n21720) );
  AND2_X1 U7106 ( .A1(n16386), .A2(n21842), .Z(n1535) );
  OAI22_X1 U7115 ( .A1(n17078), .A2(n14640), .B1(n1652), .B2(n14577), .ZN(
        n1769) );
  INV_X1 U7118 ( .I(n21350), .ZN(n1012) );
  NOR2_X1 U7119 ( .A1(n10720), .A2(n12561), .ZN(n15747) );
  NAND2_X1 U7124 ( .A1(n14577), .A2(n1652), .ZN(n21723) );
  INV_X2 U7128 ( .I(n8313), .ZN(n915) );
  INV_X1 U7135 ( .I(n8140), .ZN(n1139) );
  INV_X1 U7142 ( .I(n18213), .ZN(n6471) );
  AOI21_X1 U7157 ( .A1(n28642), .A2(n1017), .B(n20676), .ZN(n20677) );
  NAND2_X1 U7172 ( .A1(n6451), .A2(n26167), .ZN(n1784) );
  INV_X1 U7204 ( .I(n20657), .ZN(n21249) );
  AOI21_X1 U7207 ( .A1(n9405), .A2(n21452), .B(n21237), .ZN(n9406) );
  INV_X1 U7210 ( .I(n30727), .ZN(n8393) );
  INV_X1 U7240 ( .I(n20836), .ZN(n1592) );
  NOR2_X1 U7259 ( .A1(n16146), .A2(n14719), .ZN(n4857) );
  NOR2_X1 U7263 ( .A1(n28390), .A2(n20549), .ZN(n10834) );
  NAND3_X1 U7264 ( .A1(n20575), .A2(n420), .A3(n20571), .ZN(n4816) );
  INV_X1 U7273 ( .I(n20430), .ZN(n11017) );
  NAND2_X1 U7287 ( .A1(n13631), .A2(n28261), .ZN(n13630) );
  NOR2_X1 U7301 ( .A1(n20267), .A2(n26585), .ZN(n8293) );
  INV_X1 U7304 ( .I(n10939), .ZN(n20452) );
  NAND3_X1 U7313 ( .A1(n20256), .A2(n13380), .A3(n20404), .ZN(n13379) );
  BUF_X2 U7321 ( .I(n16452), .Z(n10057) );
  NAND2_X1 U7332 ( .A1(n13611), .A2(n12078), .ZN(n13608) );
  NAND2_X1 U7339 ( .A1(n5642), .A2(n17456), .ZN(n5641) );
  AOI21_X1 U7346 ( .A1(n29357), .A2(n29013), .B(n10340), .ZN(n19822) );
  NAND2_X1 U7347 ( .A1(n19876), .A2(n31103), .ZN(n20289) );
  INV_X1 U7380 ( .I(n11593), .ZN(n13841) );
  NAND2_X1 U7386 ( .A1(n1039), .A2(n14281), .ZN(n2291) );
  NAND2_X1 U7389 ( .A1(n13912), .A2(n5073), .ZN(n4051) );
  AND2_X1 U7394 ( .A1(n9748), .A2(n3526), .Z(n3525) );
  AND2_X1 U7401 ( .A1(n8301), .A2(n20008), .Z(n9875) );
  INV_X1 U7418 ( .I(n10696), .ZN(n20157) );
  INV_X1 U7429 ( .I(n8808), .ZN(n12100) );
  INV_X1 U7432 ( .I(n20088), .ZN(n16493) );
  NOR3_X1 U7439 ( .A1(n19174), .A2(n19134), .A3(n3535), .ZN(n19135) );
  NAND2_X1 U7455 ( .A1(n17370), .A2(n16699), .ZN(n1450) );
  NOR2_X1 U7458 ( .A1(n19313), .A2(n19152), .ZN(n11075) );
  NAND2_X1 U7468 ( .A1(n19604), .A2(n2799), .ZN(n3391) );
  NAND2_X1 U7474 ( .A1(n19176), .A2(n19253), .ZN(n2123) );
  NOR2_X1 U7476 ( .A1(n18994), .A2(n14892), .ZN(n5655) );
  AOI22_X1 U7478 ( .A1(n19287), .A2(n3388), .B1(n6059), .B2(n27726), .ZN(n1869) );
  NOR2_X1 U7479 ( .A1(n16916), .A2(n18979), .ZN(n2390) );
  NOR2_X1 U7486 ( .A1(n8606), .A2(n19229), .ZN(n9424) );
  AND2_X1 U7504 ( .A1(n19313), .A2(n763), .Z(n18969) );
  AND2_X1 U7508 ( .A1(n12707), .A2(n30682), .Z(n12131) );
  NOR2_X1 U7510 ( .A1(n16274), .A2(n9553), .ZN(n3244) );
  OR2_X1 U7511 ( .A1(n27726), .A2(n17817), .Z(n3365) );
  NOR2_X1 U7512 ( .A1(n19107), .A2(n19108), .ZN(n10054) );
  INV_X2 U7524 ( .I(n19123), .ZN(n8233) );
  AND2_X1 U7526 ( .A1(n25985), .A2(n1056), .Z(n9710) );
  OR2_X2 U7537 ( .A1(n10365), .A2(n4659), .Z(n4656) );
  OAI21_X1 U7565 ( .A1(n31579), .A2(n4259), .B(n18768), .ZN(n18765) );
  AOI21_X1 U7581 ( .A1(n13514), .A2(n8376), .B(n7454), .ZN(n11555) );
  NAND2_X1 U7584 ( .A1(n18795), .A2(n6119), .ZN(n7682) );
  AOI21_X1 U7585 ( .A1(n3601), .A2(n11941), .B(n26717), .ZN(n3111) );
  NAND2_X1 U7586 ( .A1(n17359), .A2(n18737), .ZN(n7733) );
  NOR2_X1 U7590 ( .A1(n17687), .A2(n18863), .ZN(n4506) );
  NAND2_X1 U7595 ( .A1(n18511), .A2(n16855), .ZN(n14453) );
  OAI21_X1 U7596 ( .A1(n13254), .A2(n34141), .B(n4677), .ZN(n12173) );
  NOR2_X1 U7598 ( .A1(n17477), .A2(n1060), .ZN(n6890) );
  OAI21_X1 U7599 ( .A1(n18785), .A2(n18801), .B(n8395), .ZN(n18628) );
  NAND3_X1 U7600 ( .A1(n3601), .A2(n10095), .A3(n732), .ZN(n3149) );
  NAND2_X1 U7603 ( .A1(n9766), .A2(n31724), .ZN(n11693) );
  NOR2_X1 U7607 ( .A1(n18815), .A2(n11918), .ZN(n8043) );
  NAND2_X1 U7611 ( .A1(n18797), .A2(n16420), .ZN(n7713) );
  NOR2_X1 U7613 ( .A1(n18706), .A2(n18707), .ZN(n18745) );
  INV_X1 U7621 ( .I(n10182), .ZN(n1189) );
  AND2_X1 U7626 ( .A1(n9909), .A2(n11459), .Z(n15495) );
  NAND2_X1 U7628 ( .A1(n16766), .A2(n31579), .ZN(n18764) );
  INV_X1 U7630 ( .I(n25832), .ZN(n1064) );
  INV_X1 U7631 ( .I(n25493), .ZN(n1065) );
  INV_X1 U7636 ( .I(n18335), .ZN(n18481) );
  INV_X2 U7638 ( .I(n32034), .ZN(n13254) );
  INV_X1 U7642 ( .I(n16464), .ZN(n1070) );
  BUF_X2 U7643 ( .I(n9909), .Z(n1709) );
  INV_X1 U7644 ( .I(n11905), .ZN(n8208) );
  INV_X1 U7646 ( .I(n16548), .ZN(n1419) );
  INV_X1 U7647 ( .I(n25108), .ZN(n1067) );
  INV_X1 U7653 ( .I(n16701), .ZN(n1069) );
  CLKBUF_X2 U7654 ( .I(Key[102]), .Z(n16548) );
  CLKBUF_X2 U7656 ( .I(Key[93]), .Z(n24968) );
  CLKBUF_X2 U7657 ( .I(Key[65]), .Z(n24386) );
  CLKBUF_X2 U7664 ( .I(Key[132]), .Z(n24943) );
  INV_X2 U7665 ( .I(n16914), .ZN(n962) );
  CLKBUF_X2 U7667 ( .I(Key[101]), .Z(n16423) );
  OAI21_X1 U7676 ( .A1(n25746), .A2(n27189), .B(n1979), .ZN(n4417) );
  NAND3_X1 U7679 ( .A1(n11003), .A2(n25816), .A3(n25804), .ZN(n11004) );
  NAND2_X1 U7683 ( .A1(n6111), .A2(n13624), .ZN(n5917) );
  NAND2_X1 U7684 ( .A1(n7929), .A2(n14511), .ZN(n11133) );
  INV_X1 U7685 ( .I(n25223), .ZN(n4188) );
  NAND2_X1 U7688 ( .A1(n25247), .A2(n2191), .ZN(n11135) );
  NAND2_X1 U7690 ( .A1(n25743), .A2(n32863), .ZN(n9414) );
  NAND2_X1 U7692 ( .A1(n25006), .A2(n3232), .ZN(n3155) );
  NAND2_X1 U7693 ( .A1(n715), .A2(n25214), .ZN(n4614) );
  AND2_X1 U7697 ( .A1(n7273), .A2(n1395), .Z(n7270) );
  INV_X1 U7699 ( .I(n11571), .ZN(n8035) );
  NAND2_X1 U7701 ( .A1(n25220), .A2(n7515), .ZN(n25222) );
  INV_X4 U7706 ( .I(n24896), .ZN(n965) );
  INV_X1 U7707 ( .I(n2983), .ZN(n2876) );
  NAND2_X1 U7710 ( .A1(n885), .A2(n17684), .ZN(n4101) );
  NAND2_X1 U7712 ( .A1(n10570), .A2(n25289), .ZN(n5535) );
  NOR2_X1 U7717 ( .A1(n24884), .A2(n25020), .ZN(n6473) );
  INV_X1 U7721 ( .I(n7081), .ZN(n10748) );
  NOR3_X1 U7725 ( .A1(n14454), .A2(n24780), .A3(n15719), .ZN(n2996) );
  OAI21_X1 U7730 ( .A1(n13042), .A2(n25885), .B(n25871), .ZN(n8541) );
  NAND2_X1 U7731 ( .A1(n15318), .A2(n4885), .ZN(n5659) );
  NOR2_X1 U7740 ( .A1(n5202), .A2(n25119), .ZN(n5203) );
  INV_X4 U7741 ( .I(n25382), .ZN(n16783) );
  OAI21_X1 U7743 ( .A1(n2158), .A2(n2156), .B(n10924), .ZN(n1645) );
  NAND2_X1 U7760 ( .A1(n24051), .A2(n15720), .ZN(n15790) );
  NOR2_X1 U7767 ( .A1(n9202), .A2(n796), .ZN(n17601) );
  AOI21_X1 U7786 ( .A1(n9323), .A2(n6286), .B(n16651), .ZN(n3548) );
  NAND2_X1 U7791 ( .A1(n2558), .A2(n14399), .ZN(n14995) );
  OAI21_X1 U7792 ( .A1(n13175), .A2(n24110), .B(n10530), .ZN(n10529) );
  OAI21_X1 U7793 ( .A1(n28945), .A2(n11200), .B(n13356), .ZN(n24178) );
  OR3_X1 U7796 ( .A1(n1087), .A2(n13343), .A3(n17068), .Z(n24115) );
  INV_X2 U7803 ( .I(n14123), .ZN(n1088) );
  OAI21_X1 U7805 ( .A1(n26158), .A2(n1775), .B(n27931), .ZN(n5045) );
  OR2_X1 U7811 ( .A1(n16643), .A2(n3718), .Z(n2686) );
  INV_X1 U7812 ( .I(n7581), .ZN(n24236) );
  NOR2_X1 U7831 ( .A1(n15660), .A2(n4408), .ZN(n3995) );
  NAND2_X1 U7832 ( .A1(n17980), .A2(n14664), .ZN(n14166) );
  NOR2_X1 U7849 ( .A1(n13521), .A2(n895), .ZN(n5954) );
  NAND2_X1 U7851 ( .A1(n15623), .A2(n23910), .ZN(n3449) );
  NAND3_X1 U7861 ( .A1(n4177), .A2(n28347), .A3(n23857), .ZN(n23801) );
  OR2_X1 U7869 ( .A1(n23778), .A2(n11392), .Z(n11391) );
  NAND2_X1 U7882 ( .A1(n29294), .A2(n11676), .ZN(n9893) );
  NOR2_X1 U7890 ( .A1(n10193), .A2(n34008), .ZN(n12070) );
  NOR2_X1 U7914 ( .A1(n22400), .A2(n33007), .ZN(n11411) );
  NAND2_X1 U7934 ( .A1(n1104), .A2(n10528), .ZN(n2342) );
  OAI21_X1 U7935 ( .A1(n1106), .A2(n7463), .B(n3668), .ZN(n3783) );
  NAND2_X1 U7944 ( .A1(n22944), .A2(n3657), .ZN(n9259) );
  NAND2_X1 U7948 ( .A1(n1484), .A2(n23104), .ZN(n10790) );
  NAND3_X1 U7950 ( .A1(n31531), .A2(n22981), .A3(n32935), .ZN(n17411) );
  NOR2_X1 U7951 ( .A1(n23109), .A2(n853), .ZN(n5895) );
  NOR2_X1 U7957 ( .A1(n6453), .A2(n16022), .ZN(n4937) );
  OAI21_X1 U7960 ( .A1(n29242), .A2(n31798), .B(n22828), .ZN(n8200) );
  INV_X1 U7982 ( .I(n32531), .ZN(n23032) );
  NAND2_X1 U7994 ( .A1(n1286), .A2(n8801), .ZN(n6712) );
  NOR2_X1 U7996 ( .A1(n31561), .A2(n22637), .ZN(n4511) );
  NAND2_X1 U8001 ( .A1(n1842), .A2(n7659), .ZN(n7658) );
  NOR2_X1 U8006 ( .A1(n22025), .A2(n8131), .ZN(n8349) );
  NAND2_X1 U8025 ( .A1(n21957), .A2(n10724), .ZN(n9547) );
  NAND2_X1 U8033 ( .A1(n12488), .A2(n639), .ZN(n10216) );
  NOR2_X1 U8038 ( .A1(n3063), .A2(n22503), .ZN(n3328) );
  AND2_X1 U8041 ( .A1(n14251), .A2(n1294), .Z(n1664) );
  NOR2_X1 U8048 ( .A1(n22690), .A2(n22689), .ZN(n3454) );
  OAI21_X1 U8055 ( .A1(n26878), .A2(n27378), .B(n12213), .ZN(n7541) );
  INV_X1 U8057 ( .I(n16375), .ZN(n22604) );
  NAND2_X1 U8059 ( .A1(n901), .A2(n22524), .ZN(n1727) );
  NOR2_X1 U8067 ( .A1(n22645), .A2(n16166), .ZN(n8595) );
  NAND2_X1 U8069 ( .A1(n10282), .A2(n10354), .ZN(n10355) );
  NOR2_X1 U8073 ( .A1(n22625), .A2(n634), .ZN(n7559) );
  INV_X1 U8076 ( .I(n11986), .ZN(n9155) );
  BUF_X2 U8078 ( .I(n22504), .Z(n3063) );
  INV_X1 U8104 ( .I(n22231), .ZN(n10429) );
  INV_X2 U8110 ( .I(n21910), .ZN(n1003) );
  AOI21_X1 U8128 ( .A1(n32073), .A2(n1134), .B(n13133), .ZN(n21599) );
  NAND3_X1 U8130 ( .A1(n1650), .A2(n21723), .A3(n28838), .ZN(n1649) );
  NOR2_X1 U8151 ( .A1(n727), .A2(n16441), .ZN(n2443) );
  NOR2_X1 U8158 ( .A1(n3043), .A2(n31197), .ZN(n3042) );
  NOR2_X1 U8161 ( .A1(n28581), .A2(n15302), .ZN(n21657) );
  NOR2_X1 U8168 ( .A1(n21489), .A2(n6718), .ZN(n3418) );
  NOR2_X1 U8175 ( .A1(n21738), .A2(n21866), .ZN(n2625) );
  NAND2_X1 U8178 ( .A1(n21235), .A2(n8029), .ZN(n11381) );
  NOR2_X1 U8182 ( .A1(n1136), .A2(n21581), .ZN(n21164) );
  NAND2_X1 U8186 ( .A1(n21461), .A2(n14640), .ZN(n1650) );
  INV_X1 U8227 ( .I(n15022), .ZN(n12587) );
  OAI22_X1 U8255 ( .A1(n1784), .A2(n1632), .B1(n925), .B2(n1783), .ZN(n1457)
         );
  NOR2_X1 U8262 ( .A1(n21451), .A2(n33498), .ZN(n1968) );
  OR2_X1 U8267 ( .A1(n21080), .A2(n17467), .Z(n13968) );
  NAND2_X1 U8268 ( .A1(n34131), .A2(n3236), .ZN(n20941) );
  NAND2_X1 U8274 ( .A1(n21393), .A2(n21367), .ZN(n16311) );
  AOI22_X1 U8280 ( .A1(n16505), .A2(n16473), .B1(n21152), .B2(n31835), .ZN(
        n12689) );
  NOR2_X1 U8292 ( .A1(n921), .A2(n21259), .ZN(n3867) );
  NOR2_X1 U8308 ( .A1(n21085), .A2(n26861), .ZN(n1867) );
  NOR2_X1 U8321 ( .A1(n1335), .A2(n14290), .ZN(n20790) );
  OR3_X1 U8328 ( .A1(n151), .A2(n21200), .A3(n17455), .Z(n9794) );
  INV_X1 U8329 ( .I(n7007), .ZN(n2277) );
  INV_X1 U8365 ( .I(n20885), .ZN(n5558) );
  OR2_X1 U8367 ( .A1(n20954), .A2(n6158), .Z(n6157) );
  NAND3_X1 U8385 ( .A1(n20601), .A2(n28288), .A3(n12583), .ZN(n2753) );
  OAI21_X1 U8416 ( .A1(n28390), .A2(n20549), .B(n12563), .ZN(n11827) );
  OR2_X1 U8418 ( .A1(n20487), .A2(n9808), .Z(n11139) );
  NOR2_X1 U8431 ( .A1(n31390), .A2(n13693), .ZN(n11826) );
  NOR2_X1 U8449 ( .A1(n1155), .A2(n30637), .ZN(n11055) );
  NOR2_X1 U8456 ( .A1(n32240), .A2(n20534), .ZN(n11839) );
  OR2_X1 U8465 ( .A1(n17947), .A2(n20485), .Z(n5878) );
  AND2_X1 U8470 ( .A1(n9688), .A2(n26881), .Z(n9689) );
  NAND2_X1 U8471 ( .A1(n8454), .A2(n4807), .ZN(n20572) );
  NOR2_X1 U8472 ( .A1(n15230), .A2(n28288), .ZN(n5030) );
  AND2_X1 U8476 ( .A1(n20570), .A2(n17236), .Z(n12999) );
  NAND2_X1 U8480 ( .A1(n1156), .A2(n20635), .ZN(n2904) );
  NOR2_X1 U8495 ( .A1(n33117), .A2(n30763), .ZN(n3442) );
  INV_X1 U8496 ( .I(n11557), .ZN(n12142) );
  NAND2_X1 U8497 ( .A1(n5641), .A2(n32296), .ZN(n5910) );
  NOR2_X1 U8498 ( .A1(n17237), .A2(n17236), .ZN(n5592) );
  NOR2_X1 U8505 ( .A1(n937), .A2(n13077), .ZN(n15849) );
  AND2_X1 U8506 ( .A1(n19952), .A2(n14927), .Z(n19953) );
  NAND2_X1 U8510 ( .A1(n3197), .A2(n729), .ZN(n1679) );
  NAND2_X1 U8523 ( .A1(n2291), .A2(n2289), .ZN(n2292) );
  NAND3_X1 U8536 ( .A1(n13771), .A2(n12100), .A3(n9876), .ZN(n1815) );
  NAND2_X1 U8539 ( .A1(n821), .A2(n19884), .ZN(n8382) );
  AOI21_X1 U8540 ( .A1(n13605), .A2(n16493), .B(n1161), .ZN(n5693) );
  NAND2_X1 U8542 ( .A1(n6263), .A2(n4674), .ZN(n14011) );
  NOR2_X1 U8545 ( .A1(n12179), .A2(n20156), .ZN(n12178) );
  NAND2_X1 U8553 ( .A1(n1438), .A2(n3790), .ZN(n12351) );
  INV_X1 U8555 ( .I(n19935), .ZN(n14171) );
  OAI21_X1 U8556 ( .A1(n20128), .A2(n875), .B(n431), .ZN(n7893) );
  NAND2_X1 U8570 ( .A1(n26551), .A2(n19456), .ZN(n5827) );
  NOR2_X1 U8571 ( .A1(n12075), .A2(n20052), .ZN(n7244) );
  NOR2_X1 U8585 ( .A1(n11959), .A2(n9724), .ZN(n9027) );
  NOR3_X1 U8587 ( .A1(n20052), .A2(n584), .A3(n17495), .ZN(n3769) );
  AND2_X1 U8588 ( .A1(n17243), .A2(n4215), .Z(n16029) );
  NOR2_X1 U8593 ( .A1(n15189), .A2(n9724), .ZN(n14793) );
  INV_X1 U8609 ( .I(n11219), .ZN(n9263) );
  INV_X1 U8610 ( .I(n7108), .ZN(n5606) );
  INV_X1 U8613 ( .I(n19589), .ZN(n13095) );
  NAND2_X1 U8614 ( .A1(n4592), .A2(n7810), .ZN(n10073) );
  NAND2_X1 U8617 ( .A1(n4405), .A2(n7680), .ZN(n4592) );
  NAND2_X1 U8635 ( .A1(n10943), .A2(n19284), .ZN(n9383) );
  AND2_X1 U8656 ( .A1(n14597), .A2(n8742), .Z(n19336) );
  INV_X1 U8657 ( .I(n26600), .ZN(n19202) );
  NOR2_X1 U8659 ( .A1(n1386), .A2(n2935), .ZN(n7201) );
  NOR2_X1 U8663 ( .A1(n13806), .A2(n947), .ZN(n6009) );
  NAND2_X1 U8665 ( .A1(n2612), .A2(n19325), .ZN(n16872) );
  NOR2_X1 U8669 ( .A1(n877), .A2(n4202), .ZN(n4218) );
  NAND2_X1 U8671 ( .A1(n2101), .A2(n19269), .ZN(n2100) );
  AND2_X1 U8678 ( .A1(n34018), .A2(n3340), .Z(n18935) );
  NOR2_X1 U8686 ( .A1(n31108), .A2(n10017), .ZN(n18908) );
  NAND2_X1 U8687 ( .A1(n19252), .A2(n29757), .ZN(n19176) );
  NOR2_X1 U8689 ( .A1(n18983), .A2(n8233), .ZN(n5636) );
  INV_X1 U8693 ( .I(n4436), .ZN(n19175) );
  NOR2_X1 U8695 ( .A1(n950), .A2(n19116), .ZN(n19117) );
  INV_X1 U8699 ( .I(n19020), .ZN(n13426) );
  NAND2_X1 U8702 ( .A1(n4053), .A2(n5646), .ZN(n5645) );
  INV_X1 U8703 ( .I(n25960), .ZN(n19121) );
  INV_X1 U8707 ( .I(n13796), .ZN(n19036) );
  NAND2_X1 U8709 ( .A1(n30958), .A2(n31949), .ZN(n4364) );
  INV_X1 U8715 ( .I(n19143), .ZN(n19253) );
  AND2_X1 U8718 ( .A1(n11203), .A2(n4016), .Z(n10453) );
  NAND2_X1 U8721 ( .A1(n8395), .A2(n6399), .ZN(n12174) );
  NOR2_X1 U8738 ( .A1(n11555), .A2(n18892), .ZN(n6794) );
  NOR2_X1 U8739 ( .A1(n28548), .A2(n12290), .ZN(n15695) );
  INV_X1 U8742 ( .I(n18653), .ZN(n9264) );
  OAI21_X1 U8745 ( .A1(n18737), .A2(n6429), .B(n6428), .ZN(n18740) );
  OAI22_X1 U8761 ( .A1(n6597), .A2(n18511), .B1(n956), .B2(n11380), .ZN(n18513) );
  NOR2_X1 U8762 ( .A1(n2733), .A2(n18893), .ZN(n2732) );
  NAND2_X1 U8765 ( .A1(n13548), .A2(n13514), .ZN(n7518) );
  NAND2_X1 U8766 ( .A1(n16403), .A2(n8395), .ZN(n18366) );
  OAI21_X1 U8768 ( .A1(n16435), .A2(n18602), .B(n15115), .ZN(n18292) );
  NAND2_X1 U8771 ( .A1(n15406), .A2(n1184), .ZN(n6173) );
  NAND2_X1 U8780 ( .A1(n18739), .A2(n18863), .ZN(n6428) );
  NOR2_X1 U8783 ( .A1(n29315), .A2(n31971), .ZN(n2596) );
  NAND2_X1 U8784 ( .A1(n18101), .A2(n1189), .ZN(n1571) );
  NOR2_X1 U8785 ( .A1(n16181), .A2(n8208), .ZN(n13243) );
  AOI21_X1 U8789 ( .A1(n28344), .A2(n18808), .B(n16474), .ZN(n2432) );
  INV_X1 U8790 ( .I(n18812), .ZN(n3180) );
  NOR2_X1 U8794 ( .A1(n7899), .A2(n18797), .ZN(n7681) );
  INV_X1 U8796 ( .I(n18569), .ZN(n15070) );
  INV_X2 U8797 ( .I(n16766), .ZN(n18642) );
  NAND2_X1 U8799 ( .A1(n16487), .A2(n497), .ZN(n6037) );
  OAI21_X1 U8808 ( .A1(n29087), .A2(n171), .B(n5473), .ZN(n17737) );
  INV_X1 U8810 ( .I(n493), .ZN(n1190) );
  NOR2_X1 U8814 ( .A1(n12290), .A2(n962), .ZN(n2964) );
  INV_X1 U8818 ( .I(n18548), .ZN(n18808) );
  AND2_X1 U8826 ( .A1(n1709), .A2(n961), .Z(n8184) );
  CLKBUF_X2 U8827 ( .I(n18707), .Z(n16487) );
  INV_X2 U8828 ( .I(n18888), .ZN(n1060) );
  INV_X1 U8831 ( .I(n18823), .ZN(n4869) );
  BUF_X2 U8832 ( .I(n18402), .Z(n18849) );
  INV_X2 U8833 ( .I(n15240), .ZN(n16855) );
  INV_X1 U8834 ( .I(n14926), .ZN(n16370) );
  INV_X1 U8836 ( .I(n16355), .ZN(n1191) );
  INV_X1 U8839 ( .I(n25190), .ZN(n1197) );
  INV_X1 U8840 ( .I(n16575), .ZN(n1196) );
  INV_X1 U8841 ( .I(n16685), .ZN(n1194) );
  INV_X1 U8842 ( .I(n16612), .ZN(n1192) );
  INV_X1 U8843 ( .I(n25373), .ZN(n1193) );
  CLKBUF_X2 U8846 ( .I(Key[140]), .Z(n24966) );
  CLKBUF_X2 U8847 ( .I(Key[41]), .Z(n25751) );
  CLKBUF_X2 U8848 ( .I(Key[68]), .Z(n25648) );
  CLKBUF_X2 U8849 ( .I(Key[77]), .Z(n24917) );
  CLKBUF_X2 U8851 ( .I(Key[127]), .Z(n16685) );
  CLKBUF_X2 U8854 ( .I(Key[38]), .Z(n24953) );
  CLKBUF_X2 U8856 ( .I(Key[188]), .Z(n25191) );
  CLKBUF_X2 U8865 ( .I(Key[176]), .Z(n25126) );
  CLKBUF_X2 U8868 ( .I(Key[86]), .Z(n25161) );
  CLKBUF_X2 U8870 ( .I(Key[95]), .Z(n25519) );
  NOR2_X1 U8872 ( .A1(n13624), .A2(n30557), .ZN(n10012) );
  NAND3_X1 U8873 ( .A1(n11005), .A2(n25819), .A3(n11004), .ZN(n15959) );
  AOI22_X1 U8876 ( .A1(n7270), .A2(n7271), .B1(n7274), .B2(n1395), .ZN(n7266)
         );
  OAI21_X1 U8881 ( .A1(n25510), .A2(n749), .B(n1946), .ZN(n1945) );
  OAI21_X1 U8885 ( .A1(n16833), .A2(n16973), .B(n963), .ZN(n6047) );
  OAI21_X1 U8889 ( .A1(n25812), .A2(n25803), .B(n25826), .ZN(n11005) );
  AOI22_X1 U8891 ( .A1(n10959), .A2(n25569), .B1(n5918), .B2(n5917), .ZN(n5916) );
  NAND2_X1 U8892 ( .A1(n7271), .A2(n7273), .ZN(n7269) );
  NOR2_X1 U8893 ( .A1(n3435), .A2(n786), .ZN(n3434) );
  AOI22_X1 U8899 ( .A1(n30318), .A2(n30288), .B1(n14737), .B2(n32059), .ZN(
        n5303) );
  NAND2_X1 U8900 ( .A1(n25193), .A2(n786), .ZN(n13245) );
  NOR2_X1 U8902 ( .A1(n32059), .A2(n2536), .ZN(n7339) );
  NAND2_X1 U8905 ( .A1(n25100), .A2(n1203), .ZN(n7335) );
  OAI21_X1 U8906 ( .A1(n9495), .A2(n13640), .B(n6915), .ZN(n9552) );
  OAI21_X1 U8907 ( .A1(n6092), .A2(n25575), .B(n25571), .ZN(n3639) );
  NAND2_X1 U8909 ( .A1(n11571), .A2(n25247), .ZN(n11569) );
  NAND2_X1 U8911 ( .A1(n25906), .A2(n1206), .ZN(n7716) );
  NAND2_X1 U8914 ( .A1(n10941), .A2(n15359), .ZN(n10940) );
  NAND2_X1 U8915 ( .A1(n27149), .A2(n4781), .ZN(n25189) );
  INV_X1 U8918 ( .I(n17637), .ZN(n8902) );
  NOR2_X1 U8919 ( .A1(n25665), .A2(n25657), .ZN(n6299) );
  NAND2_X1 U8935 ( .A1(n25391), .A2(n11556), .ZN(n6909) );
  NAND2_X1 U8944 ( .A1(n13323), .A2(n11306), .ZN(n5989) );
  NAND2_X1 U8945 ( .A1(n24734), .A2(n24733), .ZN(n24735) );
  AOI21_X1 U8951 ( .A1(n16442), .A2(n9127), .B(n11718), .ZN(n24364) );
  NOR2_X1 U8954 ( .A1(n25872), .A2(n25884), .ZN(n9111) );
  NOR2_X1 U8958 ( .A1(n9195), .A2(n24713), .ZN(n24714) );
  NAND2_X1 U8959 ( .A1(n5203), .A2(n25116), .ZN(n3794) );
  NOR2_X1 U8961 ( .A1(n3033), .A2(n17787), .ZN(n2998) );
  NAND2_X1 U8962 ( .A1(n24875), .A2(n14959), .ZN(n5624) );
  NOR2_X1 U8965 ( .A1(n5468), .A2(n25232), .ZN(n5467) );
  INV_X1 U8966 ( .I(n11752), .ZN(n25868) );
  NOR2_X1 U8969 ( .A1(n18219), .A2(n25900), .ZN(n14104) );
  NOR2_X1 U8973 ( .A1(n25388), .A2(n25590), .ZN(n10042) );
  NOR2_X1 U8976 ( .A1(n790), .A2(n1223), .ZN(n10548) );
  NAND2_X1 U8979 ( .A1(n24729), .A2(n754), .ZN(n8195) );
  NOR2_X1 U8980 ( .A1(n25566), .A2(n16648), .ZN(n10396) );
  OAI21_X1 U8983 ( .A1(n16025), .A2(n25116), .B(n25119), .ZN(n24981) );
  NAND2_X1 U8989 ( .A1(n25867), .A2(n1223), .ZN(n17489) );
  INV_X1 U8990 ( .I(n25117), .ZN(n12164) );
  NAND2_X1 U8993 ( .A1(n6034), .A2(n12039), .ZN(n25204) );
  AOI21_X1 U8994 ( .A1(n4407), .A2(n17120), .B(n25760), .ZN(n2872) );
  AOI21_X1 U8996 ( .A1(n25114), .A2(n560), .B(n18154), .ZN(n9957) );
  AND2_X1 U8998 ( .A1(n25760), .A2(n754), .Z(n13258) );
  AND2_X1 U9002 ( .A1(n5254), .A2(n28455), .Z(n12113) );
  NAND2_X1 U9004 ( .A1(n837), .A2(n12042), .ZN(n9859) );
  INV_X2 U9008 ( .I(n17867), .ZN(n25382) );
  INV_X1 U9012 ( .I(n24770), .ZN(n6862) );
  INV_X1 U9013 ( .I(n9681), .ZN(n8215) );
  INV_X1 U9016 ( .I(n18028), .ZN(n4244) );
  INV_X1 U9017 ( .I(n24622), .ZN(n3294) );
  INV_X1 U9018 ( .I(n12313), .ZN(n3305) );
  INV_X2 U9021 ( .I(n24548), .ZN(n1084) );
  NAND2_X1 U9039 ( .A1(n24140), .A2(n7203), .ZN(n6166) );
  NOR2_X1 U9047 ( .A1(n31862), .A2(n3181), .ZN(n24129) );
  NAND2_X1 U9052 ( .A1(n33680), .A2(n24242), .ZN(n2325) );
  OAI21_X1 U9054 ( .A1(n1237), .A2(n30061), .B(n3548), .ZN(n3547) );
  NAND3_X1 U9058 ( .A1(n14530), .A2(n24223), .A3(n24042), .ZN(n9965) );
  NOR2_X1 U9061 ( .A1(n24236), .A2(n32102), .ZN(n15271) );
  NOR2_X1 U9067 ( .A1(n24159), .A2(n29748), .ZN(n11435) );
  OR2_X1 U9071 ( .A1(n719), .A2(n24073), .Z(n11387) );
  NAND2_X1 U9073 ( .A1(n1240), .A2(n13412), .ZN(n7019) );
  OAI21_X1 U9084 ( .A1(n24237), .A2(n14542), .B(n32862), .ZN(n15270) );
  AOI21_X1 U9085 ( .A1(n2686), .A2(n13458), .B(n24209), .ZN(n6819) );
  OAI21_X1 U9090 ( .A1(n26750), .A2(n8058), .B(n23665), .ZN(n23666) );
  INV_X1 U9093 ( .I(n24228), .ZN(n13733) );
  NOR2_X1 U9103 ( .A1(n15065), .A2(n24177), .ZN(n13356) );
  NOR2_X1 U9106 ( .A1(n24251), .A2(n28553), .ZN(n3221) );
  NOR2_X1 U9112 ( .A1(n14399), .A2(n16868), .ZN(n3632) );
  AOI22_X1 U9118 ( .A1(n23895), .A2(n23894), .B1(n28265), .B2(n707), .ZN(n5754) );
  NAND2_X1 U9127 ( .A1(n15207), .A2(n13720), .ZN(n15206) );
  NAND2_X1 U9153 ( .A1(n23632), .A2(n33337), .ZN(n6467) );
  NOR2_X1 U9157 ( .A1(n8145), .A2(n23912), .ZN(n3446) );
  NAND2_X1 U9159 ( .A1(n16271), .A2(n8547), .ZN(n14038) );
  NAND2_X1 U9167 ( .A1(n31435), .A2(n23847), .ZN(n9329) );
  NAND2_X1 U9168 ( .A1(n7077), .A2(n1253), .ZN(n7076) );
  NOR2_X1 U9183 ( .A1(n23860), .A2(n17661), .ZN(n8865) );
  NAND2_X1 U9184 ( .A1(n4891), .A2(n8525), .ZN(n23952) );
  NOR2_X1 U9200 ( .A1(n23857), .A2(n4177), .ZN(n15186) );
  NOR2_X1 U9201 ( .A1(n31890), .A2(n13521), .ZN(n14496) );
  NOR2_X1 U9204 ( .A1(n17694), .A2(n29246), .ZN(n12031) );
  NAND2_X1 U9207 ( .A1(n10955), .A2(n29246), .ZN(n9740) );
  NAND3_X1 U9226 ( .A1(n12823), .A2(n16587), .A3(n22874), .ZN(n1671) );
  AOI21_X1 U9227 ( .A1(n12823), .A2(n22874), .B(n16587), .ZN(n1673) );
  AOI21_X1 U9234 ( .A1(n22893), .A2(n22894), .B(n23034), .ZN(n8150) );
  AOI21_X1 U9248 ( .A1(n31861), .A2(n4113), .B(n22915), .ZN(n15717) );
  NAND2_X1 U9259 ( .A1(n22972), .A2(n14420), .ZN(n2639) );
  NOR2_X1 U9263 ( .A1(n22862), .A2(n6800), .ZN(n4609) );
  INV_X1 U9264 ( .I(n11018), .ZN(n3348) );
  NAND2_X1 U9270 ( .A1(n1112), .A2(n1267), .ZN(n15831) );
  AOI21_X1 U9272 ( .A1(n897), .A2(n15704), .B(n15301), .ZN(n2029) );
  OAI21_X1 U9274 ( .A1(n11268), .A2(n641), .B(n10031), .ZN(n2032) );
  INV_X1 U9276 ( .I(n1267), .ZN(n2773) );
  NAND3_X1 U9278 ( .A1(n724), .A2(n13751), .A3(n23073), .ZN(n3162) );
  NAND2_X1 U9279 ( .A1(n10884), .A2(n723), .ZN(n10883) );
  OAI21_X1 U9280 ( .A1(n22962), .A2(n13592), .B(n8334), .ZN(n8127) );
  AND2_X1 U9297 ( .A1(n15718), .A2(n27090), .Z(n1719) );
  NAND2_X1 U9300 ( .A1(n27798), .A2(n31867), .ZN(n8201) );
  NOR2_X1 U9302 ( .A1(n27719), .A2(n31325), .ZN(n11828) );
  AND2_X1 U9312 ( .A1(n22834), .A2(n10360), .Z(n9384) );
  INV_X1 U9314 ( .I(n12687), .ZN(n12686) );
  INV_X1 U9315 ( .I(n22871), .ZN(n15389) );
  INV_X2 U9326 ( .I(n15243), .ZN(n1109) );
  OAI21_X1 U9328 ( .A1(n3502), .A2(n8260), .B(n16483), .ZN(n3501) );
  NAND3_X1 U9331 ( .A1(n15204), .A2(n12530), .A3(n13710), .ZN(n21883) );
  OAI21_X1 U9335 ( .A1(n3329), .A2(n3328), .B(n1287), .ZN(n3327) );
  AOI21_X1 U9348 ( .A1(n22449), .A2(n2381), .B(n22557), .ZN(n2380) );
  OAI21_X1 U9349 ( .A1(n11895), .A2(n28473), .B(n14591), .ZN(n14590) );
  NAND2_X1 U9358 ( .A1(n16367), .A2(n22461), .ZN(n16366) );
  AOI21_X1 U9360 ( .A1(n22404), .A2(n12496), .B(n3325), .ZN(n3324) );
  NAND2_X1 U9363 ( .A1(n11866), .A2(n29232), .ZN(n11865) );
  NAND2_X1 U9366 ( .A1(n22434), .A2(n28472), .ZN(n13008) );
  INV_X1 U9371 ( .I(n22430), .ZN(n22431) );
  NOR2_X1 U9373 ( .A1(n22329), .A2(n10354), .ZN(n9653) );
  NOR2_X1 U9374 ( .A1(n31701), .A2(n10355), .ZN(n6401) );
  NAND2_X1 U9376 ( .A1(n8594), .A2(n4315), .ZN(n8593) );
  NOR2_X1 U9387 ( .A1(n907), .A2(n10206), .ZN(n1820) );
  NOR2_X1 U9394 ( .A1(n22544), .A2(n10288), .ZN(n7237) );
  NAND2_X1 U9401 ( .A1(n13485), .A2(n8318), .ZN(n1658) );
  AOI21_X1 U9403 ( .A1(n15195), .A2(n1296), .B(n13169), .ZN(n13168) );
  NOR2_X1 U9404 ( .A1(n14376), .A2(n22672), .ZN(n4810) );
  NAND2_X1 U9407 ( .A1(n14307), .A2(n22576), .ZN(n4547) );
  NOR2_X1 U9422 ( .A1(n3063), .A2(n9370), .ZN(n3332) );
  AND2_X1 U9425 ( .A1(n17916), .A2(n1291), .Z(n15740) );
  NAND3_X1 U9427 ( .A1(n11244), .A2(n11629), .A3(n1296), .ZN(n11243) );
  NAND2_X1 U9431 ( .A1(n22540), .A2(n12844), .ZN(n4504) );
  AND2_X1 U9439 ( .A1(n12496), .A2(n3063), .Z(n3329) );
  NOR2_X1 U9443 ( .A1(n8318), .A2(n11244), .ZN(n2137) );
  AND2_X1 U9450 ( .A1(n16166), .A2(n22642), .Z(n22643) );
  AOI21_X1 U9452 ( .A1(n16166), .A2(n30641), .B(n22645), .ZN(n17191) );
  AND2_X1 U9453 ( .A1(n16432), .A2(n8527), .Z(n8529) );
  AND3_X1 U9458 ( .A1(n22452), .A2(n16567), .A3(n22576), .Z(n14219) );
  INV_X1 U9476 ( .I(n34160), .ZN(n1970) );
  NOR2_X1 U9490 ( .A1(n11796), .A2(n1647), .ZN(n7326) );
  NAND3_X1 U9495 ( .A1(n2551), .A2(n1647), .A3(n32282), .ZN(n1651) );
  NAND2_X1 U9504 ( .A1(n31910), .A2(n913), .ZN(n7323) );
  NAND2_X1 U9525 ( .A1(n21653), .A2(n21592), .ZN(n21154) );
  NAND2_X1 U9529 ( .A1(n11890), .A2(n21832), .ZN(n2300) );
  NOR2_X1 U9532 ( .A1(n21840), .A2(n4234), .ZN(n21610) );
  INV_X1 U9533 ( .I(n21823), .ZN(n8006) );
  NAND3_X1 U9546 ( .A1(n21663), .A2(n777), .A3(n31197), .ZN(n7949) );
  NAND2_X1 U9549 ( .A1(n21664), .A2(n21662), .ZN(n3049) );
  OR2_X1 U9551 ( .A1(n27619), .A2(n15026), .Z(n12448) );
  AND2_X1 U9559 ( .A1(n21737), .A2(n30152), .Z(n16371) );
  NAND2_X1 U9560 ( .A1(n11683), .A2(n11215), .ZN(n11682) );
  OAI21_X1 U9564 ( .A1(n1328), .A2(n28181), .B(n21460), .ZN(n9284) );
  NAND2_X1 U9567 ( .A1(n32642), .A2(n6489), .ZN(n16735) );
  INV_X1 U9570 ( .I(n21697), .ZN(n21656) );
  NAND2_X1 U9573 ( .A1(n432), .A2(n16194), .ZN(n6935) );
  NAND2_X1 U9588 ( .A1(n11684), .A2(n29460), .ZN(n11683) );
  NAND2_X1 U9591 ( .A1(n26407), .A2(n28642), .ZN(n11684) );
  NAND2_X1 U9610 ( .A1(n29256), .A2(n16933), .ZN(n17984) );
  INV_X1 U9625 ( .I(n21387), .ZN(n6182) );
  NAND2_X1 U9626 ( .A1(n12195), .A2(n20677), .ZN(n1559) );
  AND2_X1 U9635 ( .A1(n15506), .A2(n151), .Z(n2724) );
  NOR2_X1 U9636 ( .A1(n8657), .A2(n33454), .ZN(n5730) );
  NAND2_X1 U9645 ( .A1(n28257), .A2(n1022), .ZN(n4088) );
  NOR2_X1 U9656 ( .A1(n21269), .A2(n1017), .ZN(n12865) );
  AND2_X1 U9659 ( .A1(n21259), .A2(n21257), .Z(n10096) );
  NAND2_X1 U9667 ( .A1(n21149), .A2(n2738), .ZN(n2716) );
  NAND2_X1 U9668 ( .A1(n21389), .A2(n29901), .ZN(n6181) );
  NAND2_X1 U9675 ( .A1(n1332), .A2(n14483), .ZN(n14482) );
  INV_X1 U9679 ( .I(n349), .ZN(n21217) );
  OAI21_X1 U9683 ( .A1(n11272), .A2(n510), .B(n17455), .ZN(n12091) );
  NAND2_X1 U9684 ( .A1(n28737), .A2(n398), .ZN(n5683) );
  NAND3_X1 U9687 ( .A1(n927), .A2(n21441), .A3(n926), .ZN(n2664) );
  NAND2_X1 U9692 ( .A1(n8605), .A2(n10558), .ZN(n8604) );
  NAND2_X1 U9695 ( .A1(n21215), .A2(n12525), .ZN(n21216) );
  INV_X1 U9696 ( .I(n21263), .ZN(n21057) );
  NAND2_X1 U9706 ( .A1(n21448), .A2(n5822), .ZN(n21449) );
  INV_X1 U9709 ( .I(n30313), .ZN(n21084) );
  AOI22_X1 U9722 ( .A1(n4618), .A2(n1398), .B1(n4617), .B2(n4616), .ZN(n10110)
         );
  INV_X1 U9725 ( .I(n20711), .ZN(n8343) );
  NOR2_X1 U9726 ( .A1(n18265), .A2(n1398), .ZN(n4617) );
  NOR2_X1 U9737 ( .A1(n13572), .A2(n11634), .ZN(n8579) );
  NOR2_X1 U9752 ( .A1(n20338), .A2(n20590), .ZN(n20592) );
  INV_X1 U9755 ( .I(n14858), .ZN(n1828) );
  NAND2_X1 U9756 ( .A1(n5496), .A2(n8268), .ZN(n5350) );
  NAND2_X1 U9760 ( .A1(n4807), .A2(n816), .ZN(n8820) );
  AND2_X1 U9783 ( .A1(n9783), .A2(n31873), .Z(n10488) );
  NAND2_X1 U9787 ( .A1(n26041), .A2(n20523), .ZN(n15257) );
  NOR2_X1 U9789 ( .A1(n3443), .A2(n3442), .ZN(n3441) );
  NAND3_X1 U9790 ( .A1(n20313), .A2(n20314), .A3(n20481), .ZN(n20315) );
  NAND2_X1 U9795 ( .A1(n20525), .A2(n12169), .ZN(n9485) );
  NAND2_X1 U9799 ( .A1(n16190), .A2(n16144), .ZN(n2621) );
  NAND2_X1 U9801 ( .A1(n20377), .A2(n14179), .ZN(n5497) );
  NAND2_X1 U9808 ( .A1(n1350), .A2(n14545), .ZN(n3425) );
  OAI21_X1 U9809 ( .A1(n16518), .A2(n20533), .B(n15027), .ZN(n11038) );
  NOR2_X1 U9817 ( .A1(n20570), .A2(n31968), .ZN(n12793) );
  NOR2_X1 U9832 ( .A1(n819), .A2(n11988), .ZN(n5026) );
  NOR2_X1 U9848 ( .A1(n6864), .A2(n10752), .ZN(n7308) );
  NAND2_X1 U9849 ( .A1(n8382), .A2(n11593), .ZN(n2147) );
  NOR2_X1 U9850 ( .A1(n19921), .A2(n33525), .ZN(n7631) );
  OAI21_X1 U9853 ( .A1(n29003), .A2(n31742), .B(n15135), .ZN(n7551) );
  OR2_X1 U9868 ( .A1(n19883), .A2(n19794), .Z(n17944) );
  NOR2_X1 U9869 ( .A1(n28600), .A2(n19975), .ZN(n1898) );
  NOR2_X1 U9879 ( .A1(n10752), .A2(n19921), .ZN(n19922) );
  NOR2_X1 U9888 ( .A1(n19459), .A2(n7609), .ZN(n7607) );
  INV_X1 U9893 ( .I(n13859), .ZN(n9221) );
  NOR2_X1 U9895 ( .A1(n12168), .A2(n16848), .ZN(n5718) );
  NAND2_X1 U9901 ( .A1(n20120), .A2(n14815), .ZN(n6221) );
  AOI21_X1 U9909 ( .A1(n9563), .A2(n8100), .B(n17967), .ZN(n3270) );
  OR3_X1 U9917 ( .A1(n17260), .A2(n28600), .A3(n873), .Z(n15176) );
  INV_X1 U9923 ( .I(n13605), .ZN(n11119) );
  NAND2_X1 U9924 ( .A1(n34154), .A2(n29153), .ZN(n15602) );
  NOR2_X1 U9927 ( .A1(n12038), .A2(n11913), .ZN(n10804) );
  AND2_X1 U9929 ( .A1(n942), .A2(n15110), .Z(n9302) );
  INV_X1 U9931 ( .I(n15237), .ZN(n20138) );
  OR2_X1 U9935 ( .A1(n397), .A2(n14210), .Z(n6409) );
  INV_X1 U9939 ( .I(n20119), .ZN(n20018) );
  INV_X1 U9947 ( .I(n20098), .ZN(n19891) );
  INV_X1 U9956 ( .I(n15236), .ZN(n4976) );
  INV_X1 U9958 ( .I(n3652), .ZN(n3194) );
  INV_X1 U9963 ( .I(n11102), .ZN(n1365) );
  INV_X1 U9964 ( .I(n17430), .ZN(n5484) );
  NAND2_X1 U9974 ( .A1(n9383), .A2(n1376), .ZN(n3206) );
  OAI21_X1 U9979 ( .A1(n18935), .A2(n1386), .B(n7133), .ZN(n1655) );
  NAND2_X1 U9981 ( .A1(n8437), .A2(n33672), .ZN(n5222) );
  NOR2_X1 U9983 ( .A1(n2100), .A2(n2098), .ZN(n19073) );
  NAND2_X1 U9996 ( .A1(n14331), .A2(n4436), .ZN(n2587) );
  AOI21_X1 U10004 ( .A1(n19334), .A2(n8212), .B(n12815), .ZN(n6440) );
  NAND2_X1 U10007 ( .A1(n12502), .A2(n7557), .ZN(n6577) );
  NOR2_X1 U10008 ( .A1(n25999), .A2(n5636), .ZN(n5635) );
  AOI22_X1 U10011 ( .A1(n19182), .A2(n19181), .B1(n33078), .B2(n29769), .ZN(
        n2125) );
  NOR2_X1 U10013 ( .A1(n2283), .A2(n3340), .ZN(n6779) );
  AND2_X1 U10016 ( .A1(n19186), .A2(n947), .Z(n15675) );
  OAI22_X1 U10018 ( .A1(n17386), .A2(n19096), .B1(n29093), .B2(n10203), .ZN(
        n3115) );
  NAND2_X1 U10019 ( .A1(n31451), .A2(n5889), .ZN(n7187) );
  OR2_X1 U10020 ( .A1(n33845), .A2(n10260), .Z(n14113) );
  AND2_X1 U10021 ( .A1(n1386), .A2(n31139), .Z(n7200) );
  NAND2_X1 U10022 ( .A1(n15021), .A2(n1384), .ZN(n7901) );
  NAND2_X1 U10024 ( .A1(n13568), .A2(n824), .ZN(n9177) );
  NAND2_X1 U10026 ( .A1(n19110), .A2(n17725), .ZN(n6563) );
  OAI21_X1 U10028 ( .A1(n19334), .A2(n9538), .B(n8742), .ZN(n6282) );
  INV_X1 U10030 ( .I(n18454), .ZN(n18285) );
  NAND2_X1 U10032 ( .A1(n17817), .A2(n10124), .ZN(n3360) );
  INV_X1 U10034 ( .I(n16790), .ZN(n2871) );
  NAND2_X1 U10039 ( .A1(n27807), .A2(n6290), .ZN(n11262) );
  OAI21_X1 U10042 ( .A1(n9423), .A2(n19229), .B(n34107), .ZN(n18440) );
  OAI22_X1 U10046 ( .A1(n5877), .A2(n19199), .B1(n29047), .B2(n5876), .ZN(
        n18789) );
  INV_X1 U10047 ( .I(n5789), .ZN(n19209) );
  NOR2_X1 U10048 ( .A1(n9423), .A2(n19357), .ZN(n16769) );
  AND2_X1 U10049 ( .A1(n19262), .A2(n25971), .Z(n18751) );
  AOI21_X1 U10051 ( .A1(n25985), .A2(n33822), .B(n19146), .ZN(n10259) );
  NAND2_X1 U10054 ( .A1(n7134), .A2(n19002), .ZN(n5033) );
  NAND3_X1 U10060 ( .A1(n4365), .A2(n4364), .A3(n5789), .ZN(n4363) );
  NAND2_X1 U10064 ( .A1(n5545), .A2(n19360), .ZN(n18931) );
  AOI21_X1 U10067 ( .A1(n1053), .A2(n19109), .B(n19107), .ZN(n19111) );
  NAND2_X1 U10068 ( .A1(n19088), .A2(n19087), .ZN(n7435) );
  AND3_X1 U10069 ( .A1(n19216), .A2(n32805), .A3(n827), .Z(n6575) );
  AOI21_X1 U10072 ( .A1(n1054), .A2(n13796), .B(n11940), .ZN(n1836) );
  INV_X1 U10073 ( .I(n32788), .ZN(n18474) );
  NAND2_X1 U10074 ( .A1(n2901), .A2(n2902), .ZN(n19214) );
  NOR2_X1 U10081 ( .A1(n19257), .A2(n25971), .ZN(n4596) );
  INV_X1 U10082 ( .I(n4835), .ZN(n14806) );
  NAND2_X1 U10097 ( .A1(n8376), .A2(n7454), .ZN(n3364) );
  NAND2_X1 U10099 ( .A1(n18682), .A2(n746), .ZN(n7275) );
  NOR2_X1 U10100 ( .A1(n14614), .A2(n18407), .ZN(n10207) );
  NAND2_X1 U10101 ( .A1(n18653), .A2(n9266), .ZN(n9265) );
  NAND2_X1 U10105 ( .A1(n16854), .A2(n16855), .ZN(n3437) );
  NOR2_X1 U10108 ( .A1(n7163), .A2(n7216), .ZN(n7162) );
  NAND2_X1 U10109 ( .A1(n18311), .A2(n6173), .ZN(n6172) );
  NAND2_X1 U10115 ( .A1(n15211), .A2(n18854), .ZN(n3928) );
  NOR2_X1 U10118 ( .A1(n1571), .A2(n16538), .ZN(n14659) );
  NAND2_X1 U10124 ( .A1(n9437), .A2(n2936), .ZN(n14654) );
  NOR2_X1 U10134 ( .A1(n14695), .A2(n18875), .ZN(n14694) );
  NAND2_X1 U10135 ( .A1(n18881), .A2(n18880), .ZN(n9266) );
  NAND2_X1 U10136 ( .A1(n16995), .A2(n18539), .ZN(n14326) );
  OAI21_X1 U10146 ( .A1(n1709), .A2(n10181), .B(n11460), .ZN(n18686) );
  NOR2_X1 U10148 ( .A1(n14093), .A2(n18761), .ZN(n18336) );
  OR2_X1 U10149 ( .A1(n14906), .A2(n18511), .Z(n6918) );
  OR2_X1 U10150 ( .A1(n18566), .A2(n18492), .Z(n14678) );
  NAND2_X1 U10152 ( .A1(n18406), .A2(n18875), .ZN(n9401) );
  NAND3_X1 U10155 ( .A1(n3251), .A2(n18822), .A3(n29514), .ZN(n15957) );
  OR2_X1 U10156 ( .A1(n18463), .A2(n16915), .Z(n11954) );
  AOI21_X1 U10157 ( .A1(n18708), .A2(n18742), .B(n10665), .ZN(n17625) );
  NAND2_X1 U10159 ( .A1(n18854), .A2(n18307), .ZN(n18718) );
  NAND2_X1 U10160 ( .A1(n18856), .A2(n18853), .ZN(n3927) );
  NOR2_X1 U10161 ( .A1(n11097), .A2(n18085), .ZN(n11098) );
  NAND2_X1 U10163 ( .A1(n8739), .A2(n30371), .ZN(n6587) );
  AND2_X1 U10164 ( .A1(n34139), .A2(n18492), .Z(n18460) );
  OR2_X1 U10167 ( .A1(n18539), .A2(n14651), .Z(n2936) );
  BUF_X2 U10174 ( .I(n15265), .Z(n7454) );
  AND2_X1 U10175 ( .A1(n18770), .A2(n18774), .Z(n18274) );
  NOR2_X1 U10181 ( .A1(n18637), .A2(n18537), .ZN(n13381) );
  INV_X1 U10186 ( .I(n17419), .ZN(n11122) );
  INV_X1 U10188 ( .I(n16462), .ZN(n9729) );
  INV_X1 U10191 ( .I(n25879), .ZN(n1395) );
  INV_X1 U10193 ( .I(n16657), .ZN(n1427) );
  INV_X2 U10196 ( .I(n12166), .ZN(n18588) );
  INV_X1 U10197 ( .I(n25036), .ZN(n1398) );
  INV_X1 U10199 ( .I(n24999), .ZN(n1415) );
  INV_X1 U10200 ( .I(n25252), .ZN(n1424) );
  CLKBUF_X2 U10201 ( .I(n32034), .Z(n1446) );
  INV_X1 U10206 ( .I(n25156), .ZN(n1393) );
  INV_X1 U10207 ( .I(n16497), .ZN(n1396) );
  INV_X1 U10209 ( .I(n24707), .ZN(n1407) );
  INV_X1 U10210 ( .I(n25167), .ZN(n1413) );
  INV_X1 U10211 ( .I(n25772), .ZN(n1431) );
  INV_X1 U10212 ( .I(n24992), .ZN(n1406) );
  CLKBUF_X2 U10217 ( .I(Key[155]), .Z(n24738) );
  CLKBUF_X2 U10219 ( .I(Key[153]), .Z(n16666) );
  CLKBUF_X2 U10220 ( .I(Key[171]), .Z(n16622) );
  CLKBUF_X2 U10221 ( .I(Key[146]), .Z(n25549) );
  CLKBUF_X2 U10224 ( .I(Key[118]), .Z(n25319) );
  CLKBUF_X2 U10225 ( .I(Key[150]), .Z(n16520) );
  CLKBUF_X2 U10226 ( .I(Key[119]), .Z(n25669) );
  CLKBUF_X2 U10227 ( .I(Key[83]), .Z(n25457) );
  CLKBUF_X2 U10228 ( .I(Key[56]), .Z(n24374) );
  CLKBUF_X2 U10230 ( .I(Key[152]), .Z(n25001) );
  CLKBUF_X2 U10233 ( .I(Key[5]), .Z(n25560) );
  CLKBUF_X2 U10234 ( .I(Key[117]), .Z(n25079) );
  CLKBUF_X2 U10236 ( .I(Key[44]), .Z(n25506) );
  CLKBUF_X2 U10237 ( .I(Key[23]), .Z(n24895) );
  CLKBUF_X2 U10238 ( .I(Key[128]), .Z(n24923) );
  CLKBUF_X2 U10239 ( .I(Key[53]), .Z(n25827) );
  CLKBUF_X2 U10241 ( .I(Key[74]), .Z(n25098) );
  CLKBUF_X2 U10242 ( .I(Key[50]), .Z(n24992) );
  CLKBUF_X2 U10243 ( .I(Key[25]), .Z(n16687) );
  CLKBUF_X2 U10245 ( .I(Key[8]), .Z(n25252) );
  INV_X1 U10246 ( .I(n25641), .ZN(n1198) );
  CLKBUF_X2 U10249 ( .I(Key[71]), .Z(n25324) );
  CLKBUF_X2 U10250 ( .I(Key[62]), .Z(n25040) );
  CLKBUF_X2 U10255 ( .I(Key[149]), .Z(n25224) );
  AOI21_X1 U10267 ( .A1(n3706), .A2(n3434), .B(n3432), .ZN(n3431) );
  INV_X1 U10268 ( .I(n7303), .ZN(n5622) );
  OAI22_X1 U10278 ( .A1(n4642), .A2(n832), .B1(n25743), .B2(n1979), .ZN(n24434) );
  NAND2_X1 U10279 ( .A1(n25173), .A2(n25174), .ZN(n8339) );
  OAI21_X1 U10281 ( .A1(n5113), .A2(n7831), .B(n14321), .ZN(n14320) );
  NAND2_X1 U10285 ( .A1(n2129), .A2(n13935), .ZN(n2128) );
  NAND2_X1 U10287 ( .A1(n24934), .A2(n24925), .ZN(n5773) );
  OAI21_X1 U10292 ( .A1(n24967), .A2(n24970), .B(n3843), .ZN(n3135) );
  NAND2_X1 U10294 ( .A1(n25681), .A2(n26447), .ZN(n1757) );
  NAND2_X1 U10296 ( .A1(n25691), .A2(n25689), .ZN(n1758) );
  INV_X1 U10298 ( .I(n24972), .ZN(n2103) );
  NAND2_X1 U10299 ( .A1(n3376), .A2(n14208), .ZN(n5900) );
  NAND2_X1 U10301 ( .A1(n25650), .A2(n6299), .ZN(n7084) );
  NAND2_X1 U10302 ( .A1(n11428), .A2(n965), .ZN(n15250) );
  NAND2_X1 U10304 ( .A1(n24967), .A2(n33434), .ZN(n3846) );
  INV_X1 U10310 ( .I(n24913), .ZN(n10214) );
  NAND2_X1 U10312 ( .A1(n32859), .A2(n5712), .ZN(n5520) );
  INV_X1 U10318 ( .I(n25067), .ZN(n5865) );
  OAI21_X1 U10324 ( .A1(n3123), .A2(n3122), .B(n31640), .ZN(n6424) );
  OR3_X1 U10325 ( .A1(n25670), .A2(n25687), .A3(n25686), .Z(n24860) );
  NAND2_X1 U10328 ( .A1(n25222), .A2(n28651), .ZN(n5638) );
  NOR2_X1 U10332 ( .A1(n27183), .A2(n1074), .ZN(n9732) );
  NAND2_X1 U10335 ( .A1(n13023), .A2(n29243), .ZN(n12217) );
  INV_X1 U10336 ( .I(n25851), .ZN(n25860) );
  NOR2_X1 U10338 ( .A1(n25171), .A2(n18227), .ZN(n8930) );
  NOR2_X1 U10340 ( .A1(n2049), .A2(n25686), .ZN(n8156) );
  NOR2_X1 U10341 ( .A1(n25059), .A2(n25060), .ZN(n8257) );
  INV_X1 U10342 ( .I(n14732), .ZN(n2017) );
  INV_X1 U10349 ( .I(n27162), .ZN(n18022) );
  NAND2_X1 U10352 ( .A1(n2536), .A2(n10469), .ZN(n5408) );
  INV_X2 U10355 ( .I(n3019), .ZN(n3232) );
  INV_X1 U10358 ( .I(n17488), .ZN(n11247) );
  INV_X1 U10359 ( .I(n2191), .ZN(n25257) );
  OAI21_X1 U10361 ( .A1(n28136), .A2(n25391), .B(n6909), .ZN(n24587) );
  INV_X1 U10363 ( .I(n25172), .ZN(n18227) );
  INV_X1 U10370 ( .I(n28736), .ZN(n8073) );
  NAND2_X1 U10373 ( .A1(n15894), .A2(n11703), .ZN(n15771) );
  AND2_X1 U10393 ( .A1(n15964), .A2(n25590), .Z(n12025) );
  NAND2_X1 U10399 ( .A1(n29476), .A2(n13322), .ZN(n5990) );
  NAND2_X1 U10400 ( .A1(n5467), .A2(n17110), .ZN(n2214) );
  NOR2_X1 U10402 ( .A1(n25839), .A2(n7143), .ZN(n25840) );
  NOR2_X1 U10403 ( .A1(n10396), .A2(n10395), .ZN(n13422) );
  NAND2_X1 U10404 ( .A1(n15770), .A2(n32798), .ZN(n15894) );
  INV_X1 U10408 ( .I(n24718), .ZN(n12369) );
  NOR2_X1 U10417 ( .A1(n25761), .A2(n4407), .ZN(n4531) );
  NAND2_X1 U10420 ( .A1(n24448), .A2(n27127), .ZN(n11697) );
  OAI21_X1 U10423 ( .A1(n7064), .A2(n24714), .B(n25763), .ZN(n24717) );
  NAND2_X1 U10430 ( .A1(n1081), .A2(n13429), .ZN(n25010) );
  OR2_X1 U10432 ( .A1(n1786), .A2(n13709), .Z(n7855) );
  NOR2_X1 U10434 ( .A1(n752), .A2(n25299), .ZN(n10251) );
  NAND2_X1 U10441 ( .A1(n24981), .A2(n25114), .ZN(n3378) );
  NAND2_X1 U10442 ( .A1(n25326), .A2(n15528), .ZN(n6144) );
  INV_X1 U10447 ( .I(n4491), .ZN(n25761) );
  NAND2_X1 U10455 ( .A1(n24732), .A2(n13349), .ZN(n12968) );
  OAI21_X1 U10462 ( .A1(n17120), .A2(n25712), .B(n2872), .ZN(n2961) );
  AND2_X1 U10469 ( .A1(n13709), .A2(n25201), .Z(n25202) );
  OR2_X1 U10471 ( .A1(n25891), .A2(n25892), .Z(n12359) );
  OR2_X1 U10472 ( .A1(n25584), .A2(n718), .Z(n25585) );
  NOR2_X1 U10473 ( .A1(n886), .A2(n15528), .ZN(n10252) );
  NAND2_X1 U10475 ( .A1(n31945), .A2(n25590), .ZN(n11992) );
  NAND2_X1 U10480 ( .A1(n754), .A2(n24729), .ZN(n4452) );
  AND2_X1 U10481 ( .A1(n13050), .A2(n13042), .Z(n11976) );
  INV_X1 U10486 ( .I(n11973), .ZN(n25709) );
  INV_X2 U10488 ( .I(n675), .ZN(n1218) );
  INV_X4 U10492 ( .I(n24466), .ZN(n1221) );
  INV_X1 U10498 ( .I(n24575), .ZN(n17153) );
  INV_X1 U10499 ( .I(n17448), .ZN(n24845) );
  INV_X1 U10500 ( .I(n24518), .ZN(n13145) );
  INV_X1 U10507 ( .I(n24544), .ZN(n4566) );
  INV_X1 U10511 ( .I(n24773), .ZN(n17865) );
  INV_X1 U10512 ( .I(n24813), .ZN(n11537) );
  INV_X1 U10516 ( .I(n15508), .ZN(n8507) );
  INV_X1 U10518 ( .I(n24545), .ZN(n10257) );
  AND2_X1 U10524 ( .A1(n24166), .A2(n24165), .Z(n6051) );
  NAND2_X1 U10528 ( .A1(n3767), .A2(n3506), .ZN(n6268) );
  INV_X1 U10533 ( .I(n4728), .ZN(n8895) );
  NAND2_X1 U10534 ( .A1(n23994), .A2(n28691), .ZN(n11440) );
  INV_X2 U10541 ( .I(n283), .ZN(n1228) );
  NAND2_X1 U10549 ( .A1(n12068), .A2(n16090), .ZN(n18128) );
  NOR2_X1 U10569 ( .A1(n13047), .A2(n15253), .ZN(n7101) );
  NAND2_X1 U10573 ( .A1(n24336), .A2(n33680), .ZN(n2400) );
  OR2_X1 U10577 ( .A1(n24005), .A2(n1089), .Z(n5424) );
  INV_X1 U10578 ( .I(n17112), .ZN(n12353) );
  INV_X1 U10581 ( .I(n14530), .ZN(n13082) );
  NAND2_X1 U10583 ( .A1(n13748), .A2(n11346), .ZN(n10450) );
  NAND2_X1 U10594 ( .A1(n23666), .A2(n32459), .ZN(n7883) );
  NAND2_X1 U10601 ( .A1(n16574), .A2(n9323), .ZN(n3549) );
  NOR2_X1 U10607 ( .A1(n15271), .A2(n15270), .ZN(n24238) );
  NOR2_X1 U10608 ( .A1(n1096), .A2(n1800), .ZN(n14411) );
  INV_X1 U10610 ( .I(n6819), .ZN(n6818) );
  AND2_X1 U10613 ( .A1(n24138), .A2(n3880), .Z(n24140) );
  NOR2_X1 U10614 ( .A1(n10342), .A2(n1093), .ZN(n8399) );
  NAND2_X1 U10619 ( .A1(n2944), .A2(n13268), .ZN(n2943) );
  AND3_X1 U10620 ( .A1(n24305), .A2(n12903), .A3(n24304), .Z(n24306) );
  INV_X1 U10623 ( .I(n2686), .ZN(n2945) );
  NAND2_X1 U10636 ( .A1(n32041), .A2(n795), .ZN(n11725) );
  NAND2_X1 U10639 ( .A1(n24321), .A2(n8), .ZN(n6841) );
  NAND3_X1 U10645 ( .A1(n793), .A2(n27168), .A3(n13334), .ZN(n1838) );
  NAND2_X1 U10646 ( .A1(n15011), .A2(n24084), .ZN(n24085) );
  OR2_X1 U10654 ( .A1(n24210), .A2(n13530), .Z(n11963) );
  INV_X1 U10658 ( .I(n1090), .ZN(n1238) );
  INV_X1 U10659 ( .I(n24148), .ZN(n24121) );
  NAND4_X1 U10662 ( .A1(n4822), .A2(n4824), .A3(n4823), .A4(n4821), .ZN(n24256) );
  AND2_X1 U10663 ( .A1(n12997), .A2(n14907), .Z(n4775) );
  NAND2_X1 U10687 ( .A1(n5116), .A2(n13666), .ZN(n11079) );
  NAND2_X1 U10691 ( .A1(n13906), .A2(n13904), .ZN(n12237) );
  INV_X1 U10700 ( .I(n15474), .ZN(n5633) );
  AND2_X1 U10705 ( .A1(n16786), .A2(n23692), .Z(n8613) );
  NAND2_X1 U10708 ( .A1(n23875), .A2(n26882), .ZN(n16326) );
  NAND2_X1 U10710 ( .A1(n662), .A2(n23938), .ZN(n12080) );
  INV_X1 U10712 ( .I(n10069), .ZN(n2447) );
  NAND2_X1 U10715 ( .A1(n14164), .A2(n11095), .ZN(n12884) );
  NAND2_X1 U10729 ( .A1(n3873), .A2(n29839), .ZN(n3744) );
  NAND2_X1 U10733 ( .A1(n14088), .A2(n842), .ZN(n8344) );
  NAND2_X1 U10734 ( .A1(n12069), .A2(n14207), .ZN(n11310) );
  NAND2_X1 U10737 ( .A1(n23642), .A2(n4891), .ZN(n3757) );
  NAND2_X1 U10738 ( .A1(n12031), .A2(n548), .ZN(n3708) );
  NOR2_X1 U10740 ( .A1(n13103), .A2(n15446), .ZN(n8064) );
  NAND2_X1 U10765 ( .A1(n8865), .A2(n11904), .ZN(n2003) );
  NAND2_X1 U10767 ( .A1(n10140), .A2(n844), .ZN(n9931) );
  NAND2_X1 U10770 ( .A1(n33345), .A2(n844), .ZN(n8655) );
  NOR2_X1 U10771 ( .A1(n23637), .A2(n3650), .ZN(n11653) );
  NOR2_X1 U10776 ( .A1(n23868), .A2(n17895), .ZN(n13137) );
  OR2_X1 U10781 ( .A1(n23862), .A2(n23527), .Z(n4079) );
  INV_X1 U10783 ( .I(n16033), .ZN(n11157) );
  AND2_X1 U10785 ( .A1(n16320), .A2(n977), .Z(n12069) );
  INV_X1 U10794 ( .I(n23738), .ZN(n14155) );
  AND2_X1 U10798 ( .A1(n15682), .A2(n14325), .Z(n11975) );
  NAND3_X1 U10800 ( .A1(n1489), .A2(n23763), .A3(n23736), .ZN(n23737) );
  NOR2_X1 U10806 ( .A1(n757), .A2(n11887), .ZN(n10068) );
  INV_X1 U10808 ( .I(n13342), .ZN(n9444) );
  NAND2_X1 U10811 ( .A1(n23902), .A2(n27474), .ZN(n23176) );
  AND2_X1 U10814 ( .A1(n23848), .A2(n23807), .Z(n13544) );
  INV_X1 U10821 ( .I(n9391), .ZN(n3375) );
  NAND2_X1 U10830 ( .A1(n14585), .A2(n23763), .ZN(n23723) );
  CLKBUF_X2 U10837 ( .I(n23435), .Z(n8298) );
  INV_X1 U10842 ( .I(n12538), .ZN(n23298) );
  INV_X1 U10843 ( .I(n23386), .ZN(n9671) );
  INV_X1 U10848 ( .I(n10535), .ZN(n4409) );
  INV_X1 U10850 ( .I(n1673), .ZN(n1672) );
  INV_X1 U10856 ( .I(n23294), .ZN(n7520) );
  INV_X1 U10858 ( .I(n30321), .ZN(n23320) );
  INV_X1 U10861 ( .I(n23387), .ZN(n5514) );
  INV_X1 U10863 ( .I(n12491), .ZN(n11426) );
  INV_X1 U10868 ( .I(n4399), .ZN(n22811) );
  NAND2_X1 U10894 ( .A1(n12135), .A2(n4731), .ZN(n4730) );
  NAND2_X1 U10900 ( .A1(n2639), .A2(n2638), .ZN(n2637) );
  INV_X1 U10909 ( .I(n5971), .ZN(n2633) );
  NAND2_X1 U10912 ( .A1(n23030), .A2(n13066), .ZN(n14617) );
  NAND2_X1 U10915 ( .A1(n2624), .A2(n23103), .ZN(n2623) );
  NAND2_X1 U10921 ( .A1(n22399), .A2(n12375), .ZN(n3770) );
  AND2_X1 U10929 ( .A1(n12417), .A2(n12418), .Z(n12099) );
  OAI21_X1 U10931 ( .A1(n12016), .A2(n14114), .B(n31784), .ZN(n3513) );
  NOR2_X1 U10932 ( .A1(n23015), .A2(n27652), .ZN(n13288) );
  NAND2_X1 U10944 ( .A1(n11829), .A2(n11828), .ZN(n11837) );
  NOR2_X1 U10947 ( .A1(n22897), .A2(n27984), .ZN(n16142) );
  NAND2_X1 U10958 ( .A1(n13838), .A2(n4833), .ZN(n13837) );
  INV_X1 U10965 ( .I(n22961), .ZN(n5260) );
  AND2_X1 U10976 ( .A1(n23003), .A2(n23000), .Z(n12135) );
  AND2_X1 U10982 ( .A1(n32119), .A2(n33675), .Z(n23090) );
  NAND2_X1 U10984 ( .A1(n12218), .A2(n990), .ZN(n12180) );
  AND2_X1 U10989 ( .A1(n3891), .A2(n22836), .Z(n12033) );
  INV_X1 U10990 ( .I(n3614), .ZN(n5981) );
  INV_X1 U10992 ( .I(n22800), .ZN(n22801) );
  NAND2_X1 U10994 ( .A1(n852), .A2(n8967), .ZN(n8966) );
  INV_X1 U10998 ( .I(n9184), .ZN(n6098) );
  AOI21_X1 U11004 ( .A1(n17503), .A2(n31943), .B(n22753), .ZN(n17502) );
  NAND2_X1 U11012 ( .A1(n22592), .A2(n22705), .ZN(n11829) );
  NOR2_X1 U11013 ( .A1(n990), .A2(n30297), .ZN(n7747) );
  NAND3_X1 U11015 ( .A1(n23079), .A2(n23082), .A3(n22885), .ZN(n12646) );
  INV_X1 U11024 ( .I(n11330), .ZN(n7745) );
  INV_X1 U11029 ( .I(n3566), .ZN(n10166) );
  INV_X2 U11030 ( .I(n3668), .ZN(n23026) );
  AND2_X1 U11031 ( .A1(n23009), .A2(n23008), .Z(n23010) );
  NAND2_X1 U11033 ( .A1(n22900), .A2(n17211), .ZN(n11048) );
  AND4_X1 U11037 ( .A1(n22358), .A2(n17627), .A3(n12697), .A4(n22357), .Z(
        n9584) );
  NAND2_X1 U11038 ( .A1(n1274), .A2(n33591), .ZN(n13977) );
  INV_X1 U11049 ( .I(n17631), .ZN(n13746) );
  NAND2_X1 U11057 ( .A1(n1113), .A2(n10121), .ZN(n11853) );
  INV_X1 U11067 ( .I(n17569), .ZN(n11615) );
  AOI21_X1 U11070 ( .A1(n6384), .A2(n22678), .B(n32172), .ZN(n9738) );
  NOR2_X1 U11076 ( .A1(n30066), .A2(n22600), .ZN(n7649) );
  NAND2_X1 U11084 ( .A1(n22498), .A2(n5769), .ZN(n22499) );
  INV_X1 U11085 ( .I(n22409), .ZN(n1749) );
  NAND2_X1 U11089 ( .A1(n14830), .A2(n22639), .ZN(n15607) );
  NAND2_X1 U11091 ( .A1(n8529), .A2(n30066), .ZN(n7648) );
  NAND2_X1 U11092 ( .A1(n14830), .A2(n16240), .ZN(n11746) );
  OAI21_X1 U11097 ( .A1(n14221), .A2(n14220), .B(n22666), .ZN(n4628) );
  NAND2_X1 U11099 ( .A1(n1728), .A2(n1727), .ZN(n1726) );
  NAND2_X1 U11109 ( .A1(n9789), .A2(n1124), .ZN(n22254) );
  NOR2_X1 U11111 ( .A1(n22402), .A2(n16556), .ZN(n16232) );
  OR2_X1 U11114 ( .A1(n22544), .A2(n252), .Z(n10137) );
  INV_X1 U11116 ( .I(n22369), .ZN(n3522) );
  NAND2_X1 U11118 ( .A1(n14713), .A2(n701), .ZN(n3382) );
  NAND2_X1 U11120 ( .A1(n11575), .A2(n9603), .ZN(n3594) );
  INV_X1 U11121 ( .I(n22437), .ZN(n16414) );
  NAND2_X1 U11123 ( .A1(n4810), .A2(n905), .ZN(n4809) );
  NAND2_X1 U11137 ( .A1(n11011), .A2(n22673), .ZN(n11010) );
  INV_X2 U11139 ( .I(n12488), .ZN(n3567) );
  NOR2_X1 U11140 ( .A1(n22510), .A2(n8527), .ZN(n14765) );
  INV_X1 U11146 ( .I(n11378), .ZN(n3325) );
  NOR2_X1 U11149 ( .A1(n22536), .A2(n17626), .ZN(n17146) );
  NAND2_X1 U11156 ( .A1(n29158), .A2(n9737), .ZN(n8287) );
  INV_X1 U11158 ( .I(n22522), .ZN(n9654) );
  NOR2_X1 U11164 ( .A1(n7964), .A2(n22558), .ZN(n2844) );
  INV_X1 U11174 ( .I(n22455), .ZN(n13665) );
  NAND2_X1 U11175 ( .A1(n28865), .A2(n10622), .ZN(n11147) );
  NAND2_X1 U11178 ( .A1(n22639), .A2(n22640), .ZN(n13881) );
  AND2_X1 U11180 ( .A1(n1116), .A2(n28865), .Z(n22112) );
  NOR2_X1 U11183 ( .A1(n22537), .A2(n909), .ZN(n3188) );
  NOR2_X1 U11186 ( .A1(n22491), .A2(n26305), .ZN(n12931) );
  INV_X1 U11187 ( .I(n22669), .ZN(n15650) );
  NAND2_X1 U11199 ( .A1(n17394), .A2(n907), .ZN(n7897) );
  INV_X1 U11208 ( .I(n22504), .ZN(n22025) );
  INV_X2 U11210 ( .I(n22414), .ZN(n2066) );
  CLKBUF_X2 U11213 ( .I(n22677), .Z(n16556) );
  INV_X1 U11217 ( .I(n22289), .ZN(n16027) );
  INV_X1 U11225 ( .I(n10186), .ZN(n21874) );
  NOR2_X1 U11230 ( .A1(n14151), .A2(n14150), .ZN(n15698) );
  NAND2_X1 U11233 ( .A1(n15798), .A2(n22126), .ZN(n15797) );
  INV_X1 U11240 ( .I(n15606), .ZN(n4789) );
  INV_X1 U11242 ( .I(n13651), .ZN(n4187) );
  INV_X1 U11244 ( .I(n17362), .ZN(n4788) );
  NAND2_X1 U11250 ( .A1(n15840), .A2(n6176), .ZN(n10671) );
  OAI21_X1 U11251 ( .A1(n21562), .A2(n21561), .B(n22220), .ZN(n13370) );
  OR2_X1 U11252 ( .A1(n31930), .A2(n29180), .Z(n9961) );
  INV_X1 U11257 ( .I(n22196), .ZN(n9531) );
  NAND2_X1 U11260 ( .A1(n21756), .A2(n33403), .ZN(n15410) );
  INV_X1 U11268 ( .I(n21126), .ZN(n9312) );
  NAND2_X1 U11273 ( .A1(n21521), .A2(n21520), .ZN(n11590) );
  NAND2_X1 U11284 ( .A1(n21542), .A2(n30677), .ZN(n15129) );
  NAND2_X1 U11288 ( .A1(n5788), .A2(n5787), .ZN(n7792) );
  INV_X1 U11295 ( .I(n21754), .ZN(n21756) );
  OAI21_X1 U11299 ( .A1(n12041), .A2(n21610), .B(n27937), .ZN(n3050) );
  INV_X1 U11301 ( .I(n26113), .ZN(n2949) );
  OR2_X1 U11303 ( .A1(n2441), .A2(n7592), .Z(n2440) );
  INV_X1 U11313 ( .I(n21527), .ZN(n8459) );
  NAND2_X1 U11319 ( .A1(n21641), .A2(n21640), .ZN(n4688) );
  NAND2_X1 U11327 ( .A1(n21766), .A2(n28395), .ZN(n5997) );
  NOR2_X1 U11328 ( .A1(n21647), .A2(n26573), .ZN(n11633) );
  INV_X1 U11329 ( .I(n21818), .ZN(n21819) );
  AOI21_X1 U11340 ( .A1(n10357), .A2(n21864), .B(n15465), .ZN(n21527) );
  AND2_X1 U11343 ( .A1(n14738), .A2(n14739), .Z(n9299) );
  INV_X1 U11346 ( .I(n21491), .ZN(n11582) );
  NOR2_X1 U11347 ( .A1(n33325), .A2(n15302), .ZN(n9811) );
  NAND2_X1 U11348 ( .A1(n777), .A2(n3497), .ZN(n10346) );
  NOR2_X1 U11349 ( .A1(n16441), .A2(n25975), .ZN(n21479) );
  NOR2_X1 U11352 ( .A1(n1138), .A2(n16735), .ZN(n17164) );
  NAND2_X1 U11356 ( .A1(n21496), .A2(n21601), .ZN(n6237) );
  INV_X1 U11358 ( .I(n21797), .ZN(n21800) );
  INV_X1 U11371 ( .I(n21842), .ZN(n21750) );
  INV_X1 U11373 ( .I(n21643), .ZN(n8733) );
  INV_X1 U11375 ( .I(n21740), .ZN(n18055) );
  AND2_X1 U11377 ( .A1(n29864), .A2(n21460), .Z(n7388) );
  NOR2_X1 U11378 ( .A1(n1139), .A2(n9205), .ZN(n9204) );
  AND2_X1 U11381 ( .A1(n29980), .A2(n15302), .Z(n2202) );
  NAND2_X1 U11382 ( .A1(n13213), .A2(n28099), .ZN(n7947) );
  NOR2_X1 U11386 ( .A1(n14397), .A2(n7182), .ZN(n13869) );
  NAND2_X1 U11387 ( .A1(n6181), .A2(n21387), .ZN(n6179) );
  NOR2_X1 U11388 ( .A1(n31197), .A2(n28099), .ZN(n4098) );
  INV_X1 U11392 ( .I(n21510), .ZN(n9059) );
  INV_X1 U11397 ( .I(n10357), .ZN(n21587) );
  AND2_X1 U11398 ( .A1(n2575), .A2(n2576), .Z(n11362) );
  INV_X1 U11399 ( .I(n21723), .ZN(n13187) );
  NAND2_X1 U11401 ( .A1(n31042), .A2(n12827), .ZN(n7365) );
  NOR2_X1 U11407 ( .A1(n7182), .A2(n196), .ZN(n15827) );
  INV_X1 U11410 ( .I(n13800), .ZN(n11229) );
  INV_X1 U11412 ( .I(n21559), .ZN(n12229) );
  INV_X1 U11413 ( .I(n12792), .ZN(n1323) );
  NAND2_X1 U11414 ( .A1(n8267), .A2(n6182), .ZN(n6178) );
  INV_X1 U11416 ( .I(n12587), .ZN(n6751) );
  INV_X1 U11421 ( .I(n11266), .ZN(n21616) );
  NOR2_X1 U11429 ( .A1(n21084), .A2(n10573), .ZN(n10572) );
  OR2_X1 U11430 ( .A1(n26635), .A2(n20940), .Z(n12133) );
  INV_X1 U11433 ( .I(n13130), .ZN(n21107) );
  NAND2_X1 U11437 ( .A1(n7673), .A2(n17341), .ZN(n11315) );
  NAND2_X1 U11438 ( .A1(n21110), .A2(n21222), .ZN(n8468) );
  NOR2_X1 U11445 ( .A1(n21423), .A2(n32347), .ZN(n6881) );
  INV_X1 U11450 ( .I(n6199), .ZN(n6198) );
  NAND2_X1 U11452 ( .A1(n21413), .A2(n8657), .ZN(n3916) );
  OAI21_X1 U11456 ( .A1(n28257), .A2(n921), .B(n4088), .ZN(n21051) );
  NAND2_X1 U11460 ( .A1(n21115), .A2(n21114), .ZN(n6743) );
  NAND2_X1 U11463 ( .A1(n3105), .A2(n505), .ZN(n3104) );
  AND2_X1 U11469 ( .A1(n21209), .A2(n20874), .Z(n9095) );
  NAND2_X1 U11472 ( .A1(n11285), .A2(n21163), .ZN(n12536) );
  NAND2_X1 U11479 ( .A1(n21260), .A2(n921), .ZN(n10655) );
  NAND2_X1 U11481 ( .A1(n12492), .A2(n21270), .ZN(n10339) );
  INV_X1 U11482 ( .I(n21074), .ZN(n7147) );
  INV_X1 U11485 ( .I(n3937), .ZN(n3936) );
  INV_X1 U11492 ( .I(n6303), .ZN(n21361) );
  OAI21_X1 U11494 ( .A1(n5684), .A2(n17341), .B(n5683), .ZN(n3937) );
  INV_X1 U11495 ( .I(n1783), .ZN(n21127) );
  NAND2_X1 U11501 ( .A1(n32242), .A2(n27382), .ZN(n12340) );
  NAND2_X1 U11502 ( .A1(n21357), .A2(n6307), .ZN(n9462) );
  NOR2_X1 U11509 ( .A1(n398), .A2(n7673), .ZN(n1911) );
  INV_X1 U11512 ( .I(n21302), .ZN(n21447) );
  NAND2_X1 U11513 ( .A1(n21096), .A2(n15024), .ZN(n15023) );
  OAI21_X1 U11516 ( .A1(n4683), .A2(n320), .B(n29255), .ZN(n16545) );
  NAND2_X1 U11517 ( .A1(n1146), .A2(n320), .ZN(n21073) );
  NAND3_X1 U11518 ( .A1(n11292), .A2(n9186), .A3(n1143), .ZN(n11291) );
  NAND2_X1 U11522 ( .A1(n13101), .A2(n21311), .ZN(n11452) );
  NOR2_X1 U11524 ( .A1(n12091), .A2(n15506), .ZN(n2725) );
  OAI21_X1 U11525 ( .A1(n21131), .A2(n21307), .B(n31729), .ZN(n6199) );
  NOR2_X1 U11534 ( .A1(n8792), .A2(n8924), .ZN(n7343) );
  NOR2_X1 U11535 ( .A1(n599), .A2(n15015), .ZN(n21415) );
  NOR2_X1 U11536 ( .A1(n11513), .A2(n13367), .ZN(n14489) );
  AND2_X1 U11539 ( .A1(n21139), .A2(n21374), .Z(n11979) );
  INV_X1 U11541 ( .I(n21081), .ZN(n1868) );
  AND2_X1 U11544 ( .A1(n21295), .A2(n9721), .Z(n12111) );
  OAI21_X1 U11552 ( .A1(n15874), .A2(n21398), .B(n32625), .ZN(n15112) );
  INV_X1 U11561 ( .I(n21053), .ZN(n21054) );
  CLKBUF_X2 U11564 ( .I(n21053), .Z(n16308) );
  INV_X2 U11565 ( .I(n7738), .ZN(n21259) );
  INV_X1 U11566 ( .I(n20931), .ZN(n21182) );
  AND2_X1 U11570 ( .A1(n10533), .A2(n33566), .Z(n3032) );
  INV_X1 U11571 ( .I(n21184), .ZN(n21363) );
  INV_X1 U11573 ( .I(n27711), .ZN(n16905) );
  INV_X1 U11574 ( .I(n21136), .ZN(n21269) );
  INV_X2 U11578 ( .I(n9744), .ZN(n17985) );
  INV_X1 U11583 ( .I(n10110), .ZN(n9908) );
  INV_X1 U11585 ( .I(n8581), .ZN(n11512) );
  NAND2_X1 U11594 ( .A1(n7253), .A2(n7252), .ZN(n6158) );
  INV_X1 U11603 ( .I(n18266), .ZN(n4616) );
  INV_X1 U11612 ( .I(n20769), .ZN(n17592) );
  NAND2_X1 U11614 ( .A1(n20380), .A2(n20442), .ZN(n4913) );
  NOR2_X1 U11615 ( .A1(n20270), .A2(n28575), .ZN(n20271) );
  INV_X1 U11618 ( .I(n20861), .ZN(n7888) );
  NAND2_X1 U11625 ( .A1(n3441), .A2(n3462), .ZN(n3440) );
  NAND2_X1 U11628 ( .A1(n33902), .A2(n12224), .ZN(n6083) );
  NOR2_X1 U11629 ( .A1(n12757), .A2(n12759), .ZN(n5804) );
  INV_X1 U11630 ( .I(n20736), .ZN(n20816) );
  INV_X1 U11640 ( .I(n15168), .ZN(n3308) );
  INV_X1 U11641 ( .I(n20219), .ZN(n17003) );
  NAND2_X1 U11649 ( .A1(n20194), .A2(n32941), .ZN(n11216) );
  NOR2_X1 U11662 ( .A1(n5878), .A2(n20221), .ZN(n7478) );
  NAND2_X1 U11673 ( .A1(n9693), .A2(n1151), .ZN(n4130) );
  NOR2_X1 U11674 ( .A1(n20400), .A2(n819), .ZN(n8354) );
  NAND2_X1 U11675 ( .A1(n5498), .A2(n5497), .ZN(n5496) );
  INV_X1 U11676 ( .I(n26424), .ZN(n8868) );
  NAND2_X1 U11680 ( .A1(n34013), .A2(n1863), .ZN(n9419) );
  NAND2_X1 U11681 ( .A1(n5275), .A2(n20345), .ZN(n10716) );
  INV_X1 U11684 ( .I(n26041), .ZN(n17791) );
  NAND2_X1 U11689 ( .A1(n6925), .A2(n27771), .ZN(n5835) );
  NAND2_X1 U11692 ( .A1(n11038), .A2(n1153), .ZN(n11037) );
  INV_X1 U11693 ( .I(n20197), .ZN(n3069) );
  NAND2_X1 U11694 ( .A1(n10351), .A2(n20515), .ZN(n7254) );
  NAND2_X1 U11697 ( .A1(n12583), .A2(n5415), .ZN(n12582) );
  INV_X1 U11704 ( .I(n20405), .ZN(n11445) );
  NAND2_X1 U11712 ( .A1(n32940), .A2(n16190), .ZN(n10623) );
  OAI21_X1 U11713 ( .A1(n15553), .A2(n9774), .B(n20563), .ZN(n9773) );
  NAND3_X1 U11715 ( .A1(n14719), .A2(n12966), .A3(n28376), .ZN(n20501) );
  AND2_X1 U11724 ( .A1(n20284), .A2(n20527), .Z(n8582) );
  INV_X1 U11730 ( .I(n15225), .ZN(n20319) );
  NAND2_X1 U11731 ( .A1(n20227), .A2(n29938), .ZN(n11666) );
  NAND2_X1 U11733 ( .A1(n20304), .A2(n1028), .ZN(n7698) );
  INV_X1 U11740 ( .I(n9719), .ZN(n20199) );
  NOR2_X1 U11741 ( .A1(n1811), .A2(n1032), .ZN(n7033) );
  INV_X1 U11743 ( .I(n20304), .ZN(n5217) );
  INV_X1 U11744 ( .I(n20306), .ZN(n2134) );
  INV_X1 U11748 ( .I(n27600), .ZN(n20300) );
  OR2_X1 U11749 ( .A1(n5879), .A2(n5909), .Z(n5908) );
  AND2_X1 U11752 ( .A1(n16132), .A2(n933), .Z(n20230) );
  NAND2_X1 U11753 ( .A1(n819), .A2(n11988), .ZN(n10431) );
  AND2_X1 U11754 ( .A1(n20460), .A2(n20395), .Z(n20366) );
  NAND2_X1 U11755 ( .A1(n16606), .A2(n6531), .ZN(n17393) );
  NAND2_X1 U11768 ( .A1(n13538), .A2(n26881), .ZN(n20181) );
  NAND2_X1 U11769 ( .A1(n16146), .A2(n12421), .ZN(n20502) );
  NAND2_X1 U11770 ( .A1(n9688), .A2(n20310), .ZN(n20179) );
  OAI21_X1 U11778 ( .A1(n11502), .A2(n11501), .B(n11500), .ZN(n19816) );
  AND2_X1 U11783 ( .A1(n20290), .A2(n20289), .Z(n20291) );
  NAND2_X1 U11788 ( .A1(n19534), .A2(n20037), .ZN(n19535) );
  NAND2_X1 U11796 ( .A1(n11501), .A2(n28644), .ZN(n11500) );
  NAND2_X1 U11800 ( .A1(n11350), .A2(n568), .ZN(n19861) );
  NAND2_X1 U11805 ( .A1(n14989), .A2(n4841), .ZN(n5888) );
  INV_X1 U11810 ( .I(n6963), .ZN(n7001) );
  NAND2_X1 U11811 ( .A1(n14033), .A2(n31683), .ZN(n14032) );
  INV_X1 U11815 ( .I(n13058), .ZN(n19913) );
  NAND2_X1 U11818 ( .A1(n3271), .A2(n3270), .ZN(n3269) );
  NAND2_X1 U11819 ( .A1(n8148), .A2(n20061), .ZN(n19892) );
  NAND2_X1 U11822 ( .A1(n19869), .A2(n8137), .ZN(n19872) );
  OAI21_X1 U11825 ( .A1(n16193), .A2(n20088), .B(n1161), .ZN(n6963) );
  INV_X1 U11827 ( .I(n14801), .ZN(n3096) );
  NAND2_X1 U11828 ( .A1(n1955), .A2(n10750), .ZN(n1954) );
  OR2_X1 U11833 ( .A1(n13425), .A2(n19991), .Z(n13423) );
  NAND2_X1 U11836 ( .A1(n10683), .A2(n16346), .ZN(n8592) );
  NAND2_X1 U11837 ( .A1(n7153), .A2(n20045), .ZN(n6663) );
  NAND2_X1 U11841 ( .A1(n20055), .A2(n9379), .ZN(n11871) );
  AOI21_X1 U11846 ( .A1(n579), .A2(n16491), .B(n7460), .ZN(n15906) );
  AND2_X1 U11847 ( .A1(n1165), .A2(n5433), .Z(n6951) );
  NAND2_X1 U11853 ( .A1(n19818), .A2(n6961), .ZN(n14107) );
  INV_X1 U11855 ( .I(n10484), .ZN(n14173) );
  NAND2_X1 U11856 ( .A1(n5718), .A2(n13583), .ZN(n5717) );
  NAND2_X1 U11870 ( .A1(n29187), .A2(n25980), .ZN(n1799) );
  AND2_X1 U11875 ( .A1(n28183), .A2(n33848), .Z(n4308) );
  INV_X1 U11878 ( .I(n7525), .ZN(n1974) );
  INV_X1 U11880 ( .I(n13346), .ZN(n20077) );
  INV_X1 U11881 ( .I(n20118), .ZN(n7153) );
  INV_X1 U11884 ( .I(n34153), .ZN(n13425) );
  NOR2_X1 U11889 ( .A1(n17711), .A2(n20068), .ZN(n16516) );
  NOR2_X1 U11891 ( .A1(n19965), .A2(n8371), .ZN(n9105) );
  OAI21_X1 U11899 ( .A1(n19891), .A2(n20096), .B(n30692), .ZN(n8148) );
  NAND2_X1 U11904 ( .A1(n1040), .A2(n19456), .ZN(n5828) );
  NOR2_X1 U11909 ( .A1(n17060), .A2(n16694), .ZN(n8216) );
  NAND2_X1 U11910 ( .A1(n27097), .A2(n20152), .ZN(n19979) );
  INV_X1 U11911 ( .I(n12085), .ZN(n2290) );
  NAND2_X1 U11915 ( .A1(n1043), .A2(n16579), .ZN(n7737) );
  AND2_X1 U11916 ( .A1(n13852), .A2(n19942), .Z(n12061) );
  INV_X1 U11917 ( .I(n17060), .ZN(n11142) );
  INV_X1 U11921 ( .I(n20106), .ZN(n17696) );
  NAND3_X1 U11923 ( .A1(n20106), .A2(n20107), .A3(n16243), .ZN(n7579) );
  AND2_X1 U11924 ( .A1(n19874), .A2(n149), .Z(n11909) );
  INV_X2 U11932 ( .I(n5287), .ZN(n13605) );
  NAND2_X1 U11934 ( .A1(n577), .A2(n20096), .ZN(n17441) );
  INV_X1 U11940 ( .I(n19469), .ZN(n7191) );
  INV_X1 U11942 ( .I(n19433), .ZN(n4894) );
  INV_X1 U11945 ( .I(n19462), .ZN(n5190) );
  OAI21_X1 U11948 ( .A1(n17293), .A2(n17291), .B(n17290), .ZN(n19633) );
  INV_X1 U11949 ( .I(n19682), .ZN(n2469) );
  INV_X1 U11950 ( .I(n19545), .ZN(n6680) );
  INV_X1 U11953 ( .I(n18125), .ZN(n8266) );
  INV_X1 U11954 ( .I(n15188), .ZN(n19757) );
  INV_X1 U11962 ( .I(n19461), .ZN(n19696) );
  INV_X1 U11963 ( .I(n2282), .ZN(n2281) );
  INV_X1 U11965 ( .I(n26683), .ZN(n19570) );
  INV_X1 U11967 ( .I(n19352), .ZN(n3073) );
  INV_X1 U11969 ( .I(n32697), .ZN(n19448) );
  INV_X1 U11972 ( .I(n19445), .ZN(n19587) );
  INV_X1 U11975 ( .I(n7109), .ZN(n5608) );
  NAND2_X1 U11988 ( .A1(n15930), .A2(n11262), .ZN(n11261) );
  NOR2_X1 U11993 ( .A1(n7575), .A2(n32802), .ZN(n5332) );
  NAND2_X1 U11995 ( .A1(n10828), .A2(n19164), .ZN(n11278) );
  NAND2_X1 U11997 ( .A1(n6282), .A2(n13252), .ZN(n12894) );
  NAND2_X1 U12000 ( .A1(n10856), .A2(n10855), .ZN(n10854) );
  OAI21_X1 U12004 ( .A1(n8233), .A2(n19128), .B(n5635), .ZN(n5637) );
  INV_X1 U12007 ( .I(n6440), .ZN(n6029) );
  NAND2_X1 U12010 ( .A1(n11263), .A2(n30817), .ZN(n2518) );
  NAND2_X1 U12019 ( .A1(n3115), .A2(n15910), .ZN(n3114) );
  AND2_X1 U12021 ( .A1(n18987), .A2(n19033), .Z(n3116) );
  INV_X1 U12024 ( .I(n8092), .ZN(n4879) );
  INV_X2 U12027 ( .I(n19370), .ZN(n1372) );
  NAND2_X1 U12029 ( .A1(n1766), .A2(n19219), .ZN(n6795) );
  AOI21_X1 U12034 ( .A1(n19093), .A2(n5813), .B(n17386), .ZN(n5946) );
  OAI22_X1 U12035 ( .A1(n12034), .A2(n17725), .B1(n19107), .B2(n5907), .ZN(
        n18457) );
  NAND2_X1 U12036 ( .A1(n19209), .A2(n31948), .ZN(n9318) );
  NOR2_X1 U12038 ( .A1(n16444), .A2(n31451), .ZN(n18455) );
  NAND2_X1 U12042 ( .A1(n4363), .A2(n4202), .ZN(n4360) );
  INV_X1 U12043 ( .I(n19243), .ZN(n4217) );
  NAND2_X1 U12050 ( .A1(n3022), .A2(n14597), .ZN(n5221) );
  NAND2_X1 U12057 ( .A1(n19128), .A2(n7967), .ZN(n7966) );
  NOR2_X1 U12059 ( .A1(n14806), .A2(n10828), .ZN(n17527) );
  NAND2_X1 U12060 ( .A1(n19215), .A2(n1836), .ZN(n6603) );
  OAI21_X1 U12064 ( .A1(n13389), .A2(n11807), .B(n13390), .ZN(n13391) );
  INV_X1 U12075 ( .I(n9508), .ZN(n8671) );
  INV_X1 U12086 ( .I(n9887), .ZN(n3024) );
  INV_X1 U12087 ( .I(n3516), .ZN(n3499) );
  NOR2_X1 U12089 ( .A1(n19293), .A2(n7275), .ZN(n19297) );
  NAND2_X1 U12090 ( .A1(n15928), .A2(n15927), .ZN(n10910) );
  NOR2_X1 U12093 ( .A1(n7517), .A2(n13526), .ZN(n7516) );
  NAND2_X1 U12097 ( .A1(n14327), .A2(n14328), .ZN(n8489) );
  OAI21_X1 U12111 ( .A1(n18659), .A2(n12199), .B(n12198), .ZN(n10693) );
  NOR2_X1 U12117 ( .A1(n7454), .A2(n7518), .ZN(n7517) );
  INV_X1 U12120 ( .I(n18896), .ZN(n7714) );
  NOR2_X1 U12121 ( .A1(n12799), .A2(n18339), .ZN(n18996) );
  NAND2_X1 U12122 ( .A1(n18686), .A2(n15575), .ZN(n15574) );
  NAND2_X1 U12123 ( .A1(n5587), .A2(n1060), .ZN(n5561) );
  NAND2_X1 U12125 ( .A1(n5586), .A2(n18680), .ZN(n4717) );
  NAND2_X1 U12128 ( .A1(n18803), .A2(n18785), .ZN(n6399) );
  AOI21_X1 U12135 ( .A1(n10367), .A2(n10366), .B(n18678), .ZN(n10365) );
  NAND2_X1 U12136 ( .A1(n18336), .A2(n18755), .ZN(n9835) );
  NOR2_X1 U12138 ( .A1(n18499), .A2(n18605), .ZN(n16328) );
  NAND2_X1 U12140 ( .A1(n4868), .A2(n1190), .ZN(n8570) );
  OAI21_X1 U12143 ( .A1(n17926), .A2(n18894), .B(n18795), .ZN(n12814) );
  NOR2_X1 U12150 ( .A1(n18870), .A2(n18871), .ZN(n10305) );
  NOR2_X1 U12153 ( .A1(n3218), .A2(n18891), .ZN(n14544) );
  NAND3_X1 U12158 ( .A1(n15348), .A2(n18579), .A3(n18856), .ZN(n5124) );
  NAND2_X1 U12159 ( .A1(n11410), .A2(n6891), .ZN(n6889) );
  INV_X1 U12162 ( .I(n18410), .ZN(n18522) );
  NAND2_X1 U12163 ( .A1(n6612), .A2(n16614), .ZN(n18309) );
  AND2_X1 U12166 ( .A1(n18702), .A2(n16352), .Z(n12132) );
  NOR2_X1 U12169 ( .A1(n18130), .A2(n13738), .ZN(n18333) );
  NAND2_X1 U12172 ( .A1(n33205), .A2(n16287), .ZN(n6429) );
  INV_X1 U12174 ( .I(n18659), .ZN(n11517) );
  NAND2_X1 U12175 ( .A1(n18881), .A2(n28578), .ZN(n10639) );
  AND2_X1 U12177 ( .A1(n16474), .A2(n18349), .Z(n16120) );
  INV_X1 U12180 ( .I(n18576), .ZN(n10565) );
  INV_X1 U12182 ( .I(n15265), .ZN(n18792) );
  CLKBUF_X2 U12186 ( .I(n18654), .Z(n18446) );
  CLKBUF_X2 U12189 ( .I(n18756), .Z(n14093) );
  INV_X1 U12191 ( .I(n25693), .ZN(n25694) );
  INV_X1 U12192 ( .I(n25126), .ZN(n11034) );
  AND2_X1 U12193 ( .A1(n12006), .A2(n22), .Z(n12130) );
  INV_X1 U12194 ( .I(n25319), .ZN(n24507) );
  INV_X1 U12196 ( .I(n16479), .ZN(n3259) );
  INV_X1 U12197 ( .I(n16654), .ZN(n10308) );
  INV_X1 U12198 ( .I(n25815), .ZN(n10584) );
  INV_X1 U12199 ( .I(n25751), .ZN(n13033) );
  INV_X1 U12203 ( .I(n16502), .ZN(n15409) );
  INV_X1 U12204 ( .I(n24426), .ZN(n12754) );
  INV_X1 U12206 ( .I(n16423), .ZN(n9874) );
  INV_X1 U12208 ( .I(n25598), .ZN(n1546) );
  INV_X1 U12212 ( .I(n24943), .ZN(n24944) );
  INV_X1 U12218 ( .I(n25131), .ZN(n1653) );
  INV_X1 U12219 ( .I(n25288), .ZN(n14526) );
  INV_X1 U12220 ( .I(n25191), .ZN(n25192) );
  INV_X1 U12222 ( .I(n24738), .ZN(n5101) );
  INV_X1 U12223 ( .I(n16679), .ZN(n14300) );
  INV_X1 U12224 ( .I(n25465), .ZN(n25466) );
  INV_X1 U12225 ( .I(n25074), .ZN(n15742) );
  INV_X1 U12226 ( .I(n25506), .ZN(n25507) );
  INV_X1 U12227 ( .I(n24917), .ZN(n24918) );
  INV_X1 U12230 ( .I(n16454), .ZN(n15779) );
  INV_X1 U12232 ( .I(n24748), .ZN(n9527) );
  INV_X1 U12233 ( .I(n24907), .ZN(n13438) );
  INV_X1 U12237 ( .I(n25457), .ZN(n3027) );
  CLKBUF_X2 U12238 ( .I(n18335), .Z(n18755) );
  INV_X1 U12240 ( .I(n25560), .ZN(n8500) );
  INV_X1 U12241 ( .I(n16613), .ZN(n14885) );
  INV_X1 U12243 ( .I(n16671), .ZN(n17063) );
  INV_X1 U12244 ( .I(n16482), .ZN(n8139) );
  INV_X1 U12245 ( .I(n16602), .ZN(n10553) );
  INV_X1 U12246 ( .I(n16696), .ZN(n12719) );
  INV_X1 U12248 ( .I(n25001), .ZN(n12695) );
  INV_X1 U12249 ( .I(n16680), .ZN(n15147) );
  INV_X1 U12250 ( .I(n16642), .ZN(n1390) );
  CLKBUF_X2 U12254 ( .I(Key[89]), .Z(n24962) );
  INV_X1 U12255 ( .I(n16322), .ZN(n1397) );
  INV_X1 U12257 ( .I(n25722), .ZN(n1402) );
  INV_X1 U12259 ( .I(n16690), .ZN(n1403) );
  INV_X1 U12260 ( .I(n16631), .ZN(n1405) );
  INV_X1 U12262 ( .I(n25554), .ZN(n1409) );
  INV_X1 U12263 ( .I(n16390), .ZN(n1411) );
  CLKBUF_X2 U12266 ( .I(Key[137]), .Z(n25182) );
  INV_X1 U12268 ( .I(n25218), .ZN(n1414) );
  INV_X1 U12270 ( .I(n25049), .ZN(n1416) );
  INV_X1 U12271 ( .I(n25908), .ZN(n1417) );
  INV_X1 U12273 ( .I(n16578), .ZN(n1420) );
  INV_X1 U12274 ( .I(n25716), .ZN(n1421) );
  INV_X1 U12276 ( .I(n25038), .ZN(n1423) );
  CLKBUF_X2 U12277 ( .I(Key[21]), .Z(n16698) );
  CLKBUF_X2 U12278 ( .I(Key[63]), .Z(n25282) );
  INV_X1 U12280 ( .I(n16584), .ZN(n1425) );
  INV_X1 U12282 ( .I(n16506), .ZN(n1426) );
  INV_X1 U12283 ( .I(n16301), .ZN(n1429) );
  CLKBUF_X2 U12284 ( .I(Key[164]), .Z(n25074) );
  INV_X1 U12285 ( .I(n16666), .ZN(n1432) );
  INV_X1 U12286 ( .I(n25009), .ZN(n1433) );
  INV_X1 U12287 ( .I(n16622), .ZN(n1434) );
  XOR2_X1 U12289 ( .A1(n31491), .A2(n10776), .Z(n1436) );
  NAND3_X1 U12293 ( .A1(n1438), .A2(n3790), .A3(n1163), .ZN(n19934) );
  XOR2_X1 U12294 ( .A1(Plaintext[129]), .A2(Key[129]), .Z(n17189) );
  XOR2_X1 U12304 ( .A1(n22235), .A2(n13740), .Z(n1445) );
  NOR2_X1 U12305 ( .A1(n32787), .A2(n12317), .ZN(n18802) );
  INV_X2 U12306 ( .I(n6776), .ZN(n12317) );
  INV_X1 U12320 ( .I(n1464), .ZN(n19485) );
  XOR2_X1 U12321 ( .A1(n1464), .A2(n16654), .Z(n2980) );
  XOR2_X1 U12323 ( .A1(n1464), .A2(n3568), .Z(n19648) );
  XOR2_X1 U12324 ( .A1(n1464), .A2(n2469), .Z(n1541) );
  NOR2_X1 U12326 ( .A1(n1465), .A2(n31907), .ZN(n3746) );
  XOR2_X1 U12332 ( .A1(n24758), .A2(n24757), .Z(n1468) );
  XOR2_X1 U12337 ( .A1(n23277), .A2(n1470), .Z(n2164) );
  XOR2_X1 U12338 ( .A1(n23299), .A2(n25500), .Z(n1470) );
  OAI21_X2 U12339 ( .A1(n23080), .A2(n18129), .B(n3786), .ZN(n23299) );
  NAND2_X2 U12343 ( .A1(n1474), .A2(n1473), .ZN(n16798) );
  XOR2_X1 U12346 ( .A1(n17385), .A2(n3550), .Z(n2436) );
  XOR2_X1 U12348 ( .A1(n17385), .A2(n25554), .Z(n17564) );
  XOR2_X1 U12349 ( .A1(n22120), .A2(n17385), .Z(n4397) );
  XOR2_X1 U12350 ( .A1(n1481), .A2(n1483), .Z(n10287) );
  XOR2_X1 U12352 ( .A1(n27174), .A2(n24968), .Z(n1482) );
  XOR2_X1 U12355 ( .A1(n21014), .A2(n21015), .Z(n1483) );
  XOR2_X1 U12356 ( .A1(n20818), .A2(n20801), .Z(n21015) );
  XOR2_X1 U12359 ( .A1(n20819), .A2(n20717), .Z(n21014) );
  NOR2_X2 U12362 ( .A1(n10905), .A2(n10904), .ZN(n1485) );
  NOR2_X1 U12368 ( .A1(n23763), .A2(n1489), .ZN(n17537) );
  NAND2_X2 U12379 ( .A1(n1497), .A2(n1496), .ZN(n5268) );
  AOI22_X2 U12383 ( .A1(n1506), .A2(n23869), .B1(n13224), .B2(n23867), .ZN(
        n13223) );
  OAI21_X2 U12398 ( .A1(n1524), .A2(n1523), .B(n17357), .ZN(n22909) );
  XOR2_X1 U12405 ( .A1(n23166), .A2(n1537), .Z(n1536) );
  XOR2_X1 U12406 ( .A1(n23183), .A2(n23218), .Z(n23166) );
  XOR2_X1 U12407 ( .A1(n51), .A2(n1391), .Z(n1537) );
  NAND3_X2 U12412 ( .A1(n9950), .A2(n23054), .A3(n9949), .ZN(n23267) );
  NAND2_X2 U12417 ( .A1(n2281), .A2(n2279), .ZN(n3568) );
  XOR2_X1 U12418 ( .A1(n2470), .A2(n1541), .Z(n1540) );
  XOR2_X1 U12424 ( .A1(n32861), .A2(n27252), .Z(n4467) );
  XOR2_X1 U12427 ( .A1(n20670), .A2(n1546), .Z(n1545) );
  XOR2_X1 U12436 ( .A1(n24356), .A2(n1560), .Z(n18091) );
  XOR2_X1 U12438 ( .A1(n1560), .A2(n16655), .Z(n24391) );
  XOR2_X1 U12439 ( .A1(n14789), .A2(n1560), .Z(n7259) );
  XOR2_X1 U12440 ( .A1(n1560), .A2(n1230), .Z(n10089) );
  NAND2_X2 U12448 ( .A1(n1565), .A2(n1564), .ZN(n23293) );
  NOR2_X2 U12455 ( .A1(n32878), .A2(n4885), .ZN(n1573) );
  XOR2_X1 U12467 ( .A1(n3550), .A2(n21952), .Z(n1590) );
  XOR2_X1 U12468 ( .A1(n5482), .A2(n14289), .Z(n1587) );
  XOR2_X1 U12470 ( .A1(n22217), .A2(n454), .Z(n1588) );
  XOR2_X1 U12471 ( .A1(n11736), .A2(n22098), .Z(n22217) );
  NOR2_X1 U12481 ( .A1(n15110), .A2(n823), .ZN(n1596) );
  XOR2_X1 U12482 ( .A1(n31843), .A2(n16551), .Z(n17858) );
  XOR2_X1 U12497 ( .A1(n20443), .A2(n20669), .Z(n1612) );
  XOR2_X1 U12498 ( .A1(n8568), .A2(n20917), .Z(n20669) );
  XOR2_X1 U12504 ( .A1(n12121), .A2(n19519), .Z(n1616) );
  XOR2_X1 U12513 ( .A1(n4554), .A2(n23440), .Z(n1621) );
  XOR2_X1 U12517 ( .A1(n23334), .A2(n452), .Z(n1622) );
  XOR2_X1 U12522 ( .A1(n27114), .A2(n13545), .Z(n24538) );
  XOR2_X1 U12523 ( .A1(n27114), .A2(n7574), .Z(n18174) );
  OAI21_X1 U12528 ( .A1(n4150), .A2(n5872), .B(n25693), .ZN(n1627) );
  OR2_X1 U12529 ( .A1(n5872), .A2(n25693), .Z(n1628) );
  XOR2_X1 U12530 ( .A1(n19746), .A2(n9880), .Z(n19766) );
  AOI21_X2 U12532 ( .A1(n1631), .A2(n19254), .B(n1629), .ZN(n19746) );
  OAI21_X1 U12535 ( .A1(n20523), .A2(n1150), .B(n1635), .ZN(n20231) );
  NAND2_X2 U12537 ( .A1(n17786), .A2(n17784), .ZN(n1636) );
  XOR2_X1 U12543 ( .A1(n17384), .A2(n2155), .Z(n1644) );
  NAND2_X2 U12544 ( .A1(n1646), .A2(n1645), .ZN(n17384) );
  XOR2_X1 U12545 ( .A1(n22012), .A2(n25908), .Z(n21889) );
  INV_X2 U12549 ( .I(n11238), .ZN(n22487) );
  NAND2_X2 U12552 ( .A1(n12823), .A2(n22874), .ZN(n23331) );
  XOR2_X1 U12554 ( .A1(n10201), .A2(n23507), .Z(n1676) );
  NAND2_X2 U12555 ( .A1(n2112), .A2(n2111), .ZN(n23507) );
  AOI22_X2 U12559 ( .A1(n4255), .A2(n18784), .B1(n18787), .B2(n18786), .ZN(
        n4392) );
  NAND2_X1 U12560 ( .A1(n4392), .A2(n2150), .ZN(n5876) );
  XOR2_X1 U12561 ( .A1(n1686), .A2(n1682), .Z(n17271) );
  XOR2_X1 U12562 ( .A1(n1685), .A2(n1683), .Z(n1682) );
  XOR2_X1 U12563 ( .A1(n20970), .A2(n25001), .Z(n1683) );
  XOR2_X1 U12565 ( .A1(n20891), .A2(n20892), .Z(n1685) );
  NAND2_X2 U12567 ( .A1(n20385), .A2(n20386), .ZN(n20891) );
  XOR2_X1 U12569 ( .A1(n3705), .A2(n20839), .Z(n20890) );
  NAND2_X2 U12571 ( .A1(n20351), .A2(n20350), .ZN(n20982) );
  INV_X2 U12572 ( .I(n20727), .ZN(n20822) );
  XOR2_X1 U12578 ( .A1(n14789), .A2(n24403), .Z(n24556) );
  XOR2_X1 U12584 ( .A1(n9577), .A2(n2122), .Z(n1695) );
  XOR2_X1 U12592 ( .A1(n24567), .A2(n10163), .Z(n5530) );
  XOR2_X1 U12598 ( .A1(n20782), .A2(n3119), .Z(n1704) );
  INV_X2 U12599 ( .I(n15865), .ZN(n17661) );
  XOR2_X1 U12605 ( .A1(Plaintext[179]), .A2(Key[179]), .Z(n18874) );
  INV_X2 U12606 ( .I(n10181), .ZN(n18101) );
  XOR2_X1 U12607 ( .A1(Plaintext[178]), .A2(Key[178]), .Z(n9909) );
  XOR2_X1 U12609 ( .A1(n13477), .A2(n29312), .Z(n3178) );
  NAND2_X2 U12610 ( .A1(n2037), .A2(n12368), .ZN(n2041) );
  XOR2_X1 U12613 ( .A1(n28239), .A2(n24804), .Z(n1712) );
  NAND2_X2 U12618 ( .A1(n7325), .A2(n11590), .ZN(n10979) );
  INV_X1 U12623 ( .I(n23858), .ZN(n1732) );
  XOR2_X1 U12628 ( .A1(n11349), .A2(n25969), .Z(n1741) );
  XOR2_X1 U12634 ( .A1(n12124), .A2(n541), .Z(n1742) );
  INV_X2 U12639 ( .I(n6288), .ZN(n25687) );
  NOR2_X1 U12645 ( .A1(n25675), .A2(n14732), .ZN(n1756) );
  XOR2_X1 U12648 ( .A1(n9189), .A2(n1760), .Z(n1761) );
  XOR2_X1 U12649 ( .A1(n16693), .A2(n1069), .Z(n1760) );
  INV_X2 U12658 ( .I(n11628), .ZN(n6474) );
  XOR2_X1 U12679 ( .A1(n1780), .A2(n1779), .Z(n1778) );
  XOR2_X1 U12680 ( .A1(n14789), .A2(n13419), .Z(n1779) );
  XOR2_X1 U12681 ( .A1(n24761), .A2(n8306), .Z(n1780) );
  XOR2_X1 U12682 ( .A1(n24472), .A2(n14967), .Z(n1781) );
  NAND2_X2 U12683 ( .A1(n7660), .A2(n7658), .ZN(n4124) );
  XOR2_X1 U12685 ( .A1(n1791), .A2(n1794), .Z(n15365) );
  XOR2_X1 U12686 ( .A1(n1793), .A2(n1792), .Z(n1791) );
  XOR2_X1 U12687 ( .A1(n23336), .A2(n24374), .Z(n1792) );
  XOR2_X1 U12689 ( .A1(n1796), .A2(n1795), .Z(n1794) );
  OAI21_X1 U12693 ( .A1(n25980), .A2(n1362), .B(n1799), .ZN(n3925) );
  NAND2_X2 U12694 ( .A1(n1818), .A2(n23594), .ZN(n9964) );
  NAND4_X1 U12696 ( .A1(n14548), .A2(n1818), .A3(n14550), .A4(n23594), .ZN(
        n1800) );
  NAND2_X1 U12697 ( .A1(n3779), .A2(n32005), .ZN(n3856) );
  XOR2_X1 U12700 ( .A1(n20886), .A2(n5024), .Z(n1801) );
  NAND2_X1 U12704 ( .A1(n1803), .A2(n16041), .ZN(n17089) );
  OAI21_X1 U12706 ( .A1(n9732), .A2(n31178), .B(n32867), .ZN(n9731) );
  XOR2_X1 U12714 ( .A1(n1825), .A2(n23425), .Z(n23426) );
  XOR2_X1 U12716 ( .A1(n17775), .A2(n1825), .Z(n23062) );
  XOR2_X1 U12717 ( .A1(n23529), .A2(n1825), .Z(n23182) );
  XOR2_X1 U12721 ( .A1(n20593), .A2(n20997), .Z(n2009) );
  NOR3_X2 U12723 ( .A1(n7478), .A2(n19957), .A3(n7479), .ZN(n20699) );
  OAI21_X1 U12725 ( .A1(n7555), .A2(n28736), .B(n15323), .ZN(n1832) );
  NAND2_X1 U12726 ( .A1(n1834), .A2(n25124), .ZN(n1833) );
  NAND2_X1 U12727 ( .A1(n7554), .A2(n15323), .ZN(n1834) );
  NOR2_X1 U12729 ( .A1(n881), .A2(n32337), .ZN(n15429) );
  OAI21_X1 U12738 ( .A1(n5628), .A2(n30033), .B(n17644), .ZN(n20877) );
  XOR2_X1 U12741 ( .A1(n3929), .A2(n24748), .Z(n1844) );
  XOR2_X1 U12742 ( .A1(n20776), .A2(n7294), .Z(n1845) );
  NAND2_X2 U12762 ( .A1(n1862), .A2(n3385), .ZN(n25221) );
  XOR2_X1 U12767 ( .A1(n32822), .A2(n2388), .Z(n3357) );
  NAND2_X2 U12775 ( .A1(n9195), .A2(n25701), .ZN(n1874) );
  XOR2_X1 U12780 ( .A1(n1881), .A2(n3176), .Z(n3816) );
  XOR2_X1 U12781 ( .A1(n12413), .A2(n19441), .Z(n1881) );
  INV_X1 U12788 ( .I(n33621), .ZN(n18803) );
  XOR2_X1 U12790 ( .A1(n28730), .A2(n24923), .Z(n1884) );
  XOR2_X1 U12794 ( .A1(n20838), .A2(n20748), .Z(n1886) );
  XOR2_X1 U12795 ( .A1(n20747), .A2(n21043), .Z(n20838) );
  NAND2_X1 U12798 ( .A1(n19837), .A2(n20037), .ZN(n19838) );
  OR2_X1 U12808 ( .A1(n19976), .A2(n32746), .Z(n1900) );
  XOR2_X1 U12811 ( .A1(n859), .A2(n1903), .Z(n1902) );
  XOR2_X1 U12814 ( .A1(n10824), .A2(n1970), .Z(n1905) );
  INV_X1 U12817 ( .I(n11617), .ZN(n1909) );
  AOI21_X1 U12824 ( .A1(n28737), .A2(n17341), .B(n16184), .ZN(n1914) );
  XOR2_X1 U12827 ( .A1(n31616), .A2(n24962), .Z(n5012) );
  XOR2_X1 U12828 ( .A1(n31616), .A2(n25182), .Z(n21947) );
  XOR2_X1 U12829 ( .A1(n22055), .A2(n31616), .Z(n16912) );
  AOI21_X1 U12835 ( .A1(n25234), .A2(n16589), .B(n8219), .ZN(n8121) );
  XOR2_X1 U12837 ( .A1(n1928), .A2(n1927), .Z(n10436) );
  XOR2_X1 U12838 ( .A1(n20679), .A2(n25476), .Z(n1927) );
  XOR2_X1 U12839 ( .A1(n3929), .A2(n21016), .Z(n1928) );
  XOR2_X1 U12842 ( .A1(n14897), .A2(n11170), .Z(n11169) );
  XOR2_X1 U12844 ( .A1(n2362), .A2(n12141), .Z(n12260) );
  XOR2_X1 U12849 ( .A1(n4295), .A2(n32981), .Z(n1936) );
  XOR2_X1 U12864 ( .A1(n27167), .A2(n1191), .Z(n1948) );
  XOR2_X1 U12865 ( .A1(n13470), .A2(n14665), .Z(n24774) );
  NAND2_X1 U12868 ( .A1(n30330), .A2(n1951), .ZN(n25069) );
  NOR2_X1 U12869 ( .A1(n25076), .A2(n1951), .ZN(n12304) );
  NAND3_X1 U12870 ( .A1(n25076), .A2(n25066), .A3(n1951), .ZN(n25068) );
  OAI21_X1 U12874 ( .A1(n12329), .A2(n25066), .B(n1951), .ZN(n1950) );
  MUX2_X1 U12879 ( .I0(n10086), .I1(n19921), .S(n10752), .Z(n1955) );
  INV_X1 U12889 ( .I(n1982), .ZN(n13149) );
  XOR2_X1 U12891 ( .A1(n19672), .A2(n1984), .Z(n11627) );
  XOR2_X1 U12892 ( .A1(n1984), .A2(n16598), .Z(n17538) );
  NAND2_X1 U12894 ( .A1(n24076), .A2(n1233), .ZN(n24077) );
  XOR2_X1 U12899 ( .A1(n4134), .A2(n6966), .Z(n1988) );
  XOR2_X1 U12903 ( .A1(n34078), .A2(n22198), .Z(n1990) );
  XOR2_X1 U12905 ( .A1(n14851), .A2(n22240), .Z(n1992) );
  INV_X2 U12908 ( .I(n6462), .ZN(n13612) );
  XOR2_X1 U12913 ( .A1(n20852), .A2(n1993), .Z(n14668) );
  NAND2_X1 U12918 ( .A1(n219), .A2(n1040), .ZN(n19995) );
  XOR2_X1 U12929 ( .A1(n24812), .A2(n24554), .Z(n2012) );
  XOR2_X1 U12934 ( .A1(n24664), .A2(n25071), .Z(n2015) );
  AOI22_X2 U12937 ( .A1(n2018), .A2(n11497), .B1(n27947), .B2(n24460), .ZN(
        n25686) );
  XOR2_X1 U12947 ( .A1(n24486), .A2(n2048), .Z(n2043) );
  XOR2_X1 U12948 ( .A1(n24770), .A2(n2864), .Z(n24486) );
  XOR2_X1 U12949 ( .A1(n16917), .A2(n13810), .Z(n2044) );
  XOR2_X1 U12951 ( .A1(n1228), .A2(n14762), .Z(n13810) );
  NAND2_X1 U12955 ( .A1(n26447), .A2(n2049), .ZN(n25673) );
  XOR2_X1 U12959 ( .A1(n16608), .A2(n19767), .Z(n2053) );
  XOR2_X1 U12960 ( .A1(n3357), .A2(n3358), .Z(n2054) );
  XOR2_X1 U12968 ( .A1(n23233), .A2(n23536), .Z(n15497) );
  XOR2_X1 U12969 ( .A1(n1258), .A2(n721), .Z(n14122) );
  NOR2_X1 U12976 ( .A1(n22487), .A2(n2066), .ZN(n13169) );
  NAND2_X1 U12977 ( .A1(n31964), .A2(n2066), .ZN(n16963) );
  MUX2_X1 U12978 ( .I0(n2066), .I1(n31964), .S(n33046), .Z(n11246) );
  AOI22_X2 U12981 ( .A1(n13364), .A2(n17398), .B1(n8145), .B2(n13936), .ZN(
        n24240) );
  NAND2_X1 U12990 ( .A1(n1098), .A2(n34009), .ZN(n8852) );
  NAND3_X1 U12991 ( .A1(n763), .A2(n7197), .A3(n2081), .ZN(n18905) );
  OAI21_X1 U12992 ( .A1(n825), .A2(n31970), .B(n2081), .ZN(n16908) );
  XOR2_X1 U12996 ( .A1(n2082), .A2(n22155), .Z(n8341) );
  NOR2_X1 U12999 ( .A1(n23046), .A2(n808), .ZN(n2084) );
  NOR2_X1 U13000 ( .A1(n13121), .A2(n13120), .ZN(n2085) );
  XOR2_X1 U13018 ( .A1(n2095), .A2(n2097), .Z(n8099) );
  XOR2_X1 U13021 ( .A1(n22309), .A2(n22310), .Z(n2097) );
  XOR2_X1 U13022 ( .A1(n11736), .A2(n13564), .Z(n22310) );
  AOI21_X2 U13023 ( .A1(n4688), .A2(n21643), .B(n4687), .ZN(n13564) );
  NAND2_X2 U13029 ( .A1(n11396), .A2(n14844), .ZN(n15502) );
  INV_X2 U13040 ( .I(n2108), .ZN(n5897) );
  XOR2_X1 U13042 ( .A1(n3599), .A2(n19632), .Z(n19636) );
  XOR2_X1 U13043 ( .A1(n3599), .A2(n19072), .Z(n10224) );
  NAND2_X1 U13051 ( .A1(n11153), .A2(n2118), .ZN(n11152) );
  XOR2_X1 U13054 ( .A1(n2331), .A2(n25669), .Z(n2122) );
  XOR2_X1 U13068 ( .A1(n30749), .A2(n20729), .Z(n15936) );
  XOR2_X1 U13073 ( .A1(n22150), .A2(n5352), .Z(n2144) );
  NOR2_X1 U13079 ( .A1(n10203), .A2(n26417), .ZN(n19092) );
  NAND3_X1 U13080 ( .A1(n10203), .A2(n31658), .A3(n26417), .ZN(n18987) );
  AOI21_X1 U13081 ( .A1(n31658), .A2(n8141), .B(n26417), .ZN(n18790) );
  OAI21_X1 U13082 ( .A1(n5813), .A2(n8141), .B(n26417), .ZN(n5812) );
  NAND2_X1 U13087 ( .A1(n9521), .A2(n4019), .ZN(n2154) );
  XOR2_X1 U13089 ( .A1(n33700), .A2(n15000), .Z(n2155) );
  XOR2_X1 U13092 ( .A1(n13020), .A2(n5031), .Z(n2161) );
  INV_X2 U13093 ( .I(n2163), .ZN(n13297) );
  AND2_X1 U13095 ( .A1(n31916), .A2(n13297), .Z(n23562) );
  XOR2_X1 U13099 ( .A1(n582), .A2(n16678), .Z(n9201) );
  XOR2_X1 U13101 ( .A1(Plaintext[191]), .A2(Key[191]), .Z(n10891) );
  AOI21_X1 U13108 ( .A1(n24924), .A2(n2180), .B(n15799), .ZN(n24931) );
  XOR2_X1 U13115 ( .A1(n23454), .A2(n27243), .Z(n2190) );
  NOR2_X1 U13116 ( .A1(n5568), .A2(n2191), .ZN(n16348) );
  NAND3_X1 U13117 ( .A1(n3646), .A2(n7929), .A3(n2191), .ZN(n16583) );
  OAI21_X1 U13118 ( .A1(n25247), .A2(n34109), .B(n2191), .ZN(n8036) );
  NAND2_X2 U13119 ( .A1(n4552), .A2(n25245), .ZN(n2191) );
  NAND3_X2 U13123 ( .A1(n2197), .A2(n13563), .A3(n13562), .ZN(n16331) );
  NAND2_X1 U13128 ( .A1(n20379), .A2(n2205), .ZN(n2204) );
  NOR2_X1 U13129 ( .A1(n6679), .A2(n20635), .ZN(n2205) );
  NAND2_X1 U13132 ( .A1(n2209), .A2(n25687), .ZN(n25680) );
  OAI22_X1 U13134 ( .A1(n26447), .A2(n27173), .B1(n25687), .B2(n2209), .ZN(
        n2208) );
  XOR2_X1 U13136 ( .A1(n24370), .A2(n16733), .Z(n9681) );
  XOR2_X1 U13140 ( .A1(n2212), .A2(n24541), .Z(n2211) );
  XOR2_X1 U13141 ( .A1(n705), .A2(n26002), .Z(n2212) );
  OAI21_X2 U13143 ( .A1(n12919), .A2(n2219), .B(n2215), .ZN(n21910) );
  NAND2_X1 U13149 ( .A1(n3007), .A2(n1274), .ZN(n2226) );
  XOR2_X1 U13151 ( .A1(n11641), .A2(n620), .Z(n2547) );
  NOR2_X1 U13154 ( .A1(n31046), .A2(n2229), .ZN(n19817) );
  NAND3_X1 U13158 ( .A1(n28734), .A2(n25322), .A3(n16041), .ZN(n25323) );
  NAND2_X1 U13161 ( .A1(n25320), .A2(n28734), .ZN(n9733) );
  NOR2_X1 U13162 ( .A1(n8770), .A2(n2237), .ZN(n12917) );
  NAND3_X1 U13164 ( .A1(n1028), .A2(n1151), .A3(n2237), .ZN(n7252) );
  XOR2_X1 U13181 ( .A1(n22036), .A2(n16523), .Z(n2261) );
  XOR2_X1 U13182 ( .A1(n2262), .A2(n12695), .Z(Ciphertext[32]) );
  OAI21_X1 U13186 ( .A1(n3019), .A2(n30279), .B(n2266), .ZN(n2265) );
  XOR2_X1 U13189 ( .A1(n21023), .A2(n2268), .Z(n2267) );
  XOR2_X1 U13190 ( .A1(n7717), .A2(n25545), .Z(n2268) );
  XOR2_X1 U13195 ( .A1(n19701), .A2(n19697), .Z(n18166) );
  XNOR2_X1 U13196 ( .A1(n16349), .A2(n19661), .ZN(n19701) );
  NAND2_X1 U13198 ( .A1(n2271), .A2(n7001), .ZN(n6995) );
  NAND2_X1 U13199 ( .A1(n26088), .A2(n2271), .ZN(n6994) );
  XOR2_X1 U13202 ( .A1(Plaintext[54]), .A2(Key[54]), .Z(n16849) );
  XOR2_X1 U13207 ( .A1(n24747), .A2(n2278), .Z(n2699) );
  OAI21_X2 U13209 ( .A1(n11042), .A2(n24199), .B(n24020), .ZN(n2278) );
  AOI21_X1 U13210 ( .A1(n19038), .A2(n19039), .B(n28157), .ZN(n2282) );
  NAND2_X1 U13214 ( .A1(n2290), .A2(n10845), .ZN(n2289) );
  NAND2_X1 U13220 ( .A1(n12147), .A2(n12148), .ZN(n2302) );
  XOR2_X1 U13225 ( .A1(n21020), .A2(n2306), .Z(n2305) );
  XOR2_X1 U13226 ( .A1(n21019), .A2(n1923), .Z(n2306) );
  INV_X2 U13235 ( .I(n2312), .ZN(n2450) );
  INV_X2 U13236 ( .I(n2315), .ZN(n2378) );
  MUX2_X1 U13237 ( .I0(n15295), .I1(n18151), .S(n2378), .Z(n9198) );
  OAI21_X2 U13240 ( .A1(n20360), .A2(n2320), .B(n2319), .ZN(n20813) );
  INV_X2 U13243 ( .I(n14934), .ZN(n21438) );
  XOR2_X1 U13247 ( .A1(n19772), .A2(n24426), .Z(n2333) );
  XOR2_X1 U13248 ( .A1(n13106), .A2(n31731), .Z(n2334) );
  XOR2_X1 U13264 ( .A1(n7256), .A2(n24763), .Z(n24472) );
  XOR2_X1 U13268 ( .A1(n26623), .A2(n358), .Z(n2365) );
  XOR2_X1 U13270 ( .A1(n2367), .A2(n23151), .Z(n2968) );
  XOR2_X1 U13271 ( .A1(n2367), .A2(n23236), .Z(n15374) );
  OAI21_X1 U13279 ( .A1(n3032), .A2(n6520), .B(n2369), .ZN(n2371) );
  NOR2_X1 U13281 ( .A1(n33566), .A2(n30813), .ZN(n12027) );
  XNOR2_X1 U13288 ( .A1(n10979), .A2(n22028), .ZN(n22070) );
  OR2_X1 U13290 ( .A1(n6798), .A2(n22949), .Z(n6675) );
  XOR2_X1 U13298 ( .A1(n31950), .A2(n1413), .Z(n2384) );
  XOR2_X1 U13305 ( .A1(n19168), .A2(n2389), .Z(n5402) );
  XOR2_X1 U13306 ( .A1(n19484), .A2(n2388), .Z(n2389) );
  NOR2_X1 U13317 ( .A1(n2479), .A2(n22949), .ZN(n2405) );
  XOR2_X1 U13324 ( .A1(n11869), .A2(n14784), .Z(n2414) );
  XOR2_X1 U13325 ( .A1(n20958), .A2(n14785), .Z(n2415) );
  NAND3_X1 U13330 ( .A1(n10046), .A2(n24675), .A3(n23964), .ZN(n2420) );
  XOR2_X1 U13340 ( .A1(n5875), .A2(n2436), .Z(n2435) );
  NAND2_X2 U13344 ( .A1(n2442), .A2(n2440), .ZN(n17385) );
  AOI21_X1 U13345 ( .A1(n21715), .A2(n21601), .B(n21496), .ZN(n2441) );
  NAND2_X1 U13351 ( .A1(n2449), .A2(n28942), .ZN(n10496) );
  NOR2_X1 U13352 ( .A1(n9224), .A2(n2449), .ZN(n9003) );
  XOR2_X1 U13358 ( .A1(n2045), .A2(n16253), .Z(n2452) );
  XNOR2_X1 U13359 ( .A1(n24810), .A2(n91), .ZN(n16002) );
  INV_X2 U13370 ( .I(n2455), .ZN(n6976) );
  NAND2_X2 U13371 ( .A1(n1083), .A2(n18080), .ZN(n2456) );
  XOR2_X1 U13375 ( .A1(n2221), .A2(n6386), .Z(n2458) );
  INV_X2 U13376 ( .I(n12617), .ZN(n24308) );
  NAND2_X2 U13379 ( .A1(n2466), .A2(n2464), .ZN(n15716) );
  XOR2_X1 U13381 ( .A1(n4321), .A2(n1069), .Z(n2470) );
  XOR2_X1 U13382 ( .A1(n17830), .A2(n2472), .Z(n2473) );
  XOR2_X1 U13383 ( .A1(n20905), .A2(n25815), .Z(n2472) );
  XOR2_X1 U13388 ( .A1(n20928), .A2(n15), .Z(n2476) );
  INV_X1 U13389 ( .I(n22274), .ZN(n18058) );
  NAND2_X1 U13394 ( .A1(n1204), .A2(n6595), .ZN(n18215) );
  NAND2_X1 U13401 ( .A1(n25146), .A2(n5020), .ZN(n17525) );
  XOR2_X1 U13402 ( .A1(n24829), .A2(n5021), .Z(n2489) );
  OAI21_X2 U13403 ( .A1(n17385), .A2(n22099), .B(n2490), .ZN(n16971) );
  NAND2_X2 U13404 ( .A1(n2491), .A2(n21126), .ZN(n22099) );
  NOR2_X2 U13408 ( .A1(n23565), .A2(n23564), .ZN(n24150) );
  NAND2_X1 U13409 ( .A1(n4065), .A2(n25119), .ZN(n2498) );
  NAND2_X1 U13410 ( .A1(n1205), .A2(n254), .ZN(n15016) );
  NAND2_X2 U13411 ( .A1(n2498), .A2(n2497), .ZN(n25007) );
  AND2_X1 U13412 ( .A1(n24885), .A2(n24886), .Z(n2497) );
  XOR2_X1 U13415 ( .A1(n4028), .A2(n19681), .Z(n2500) );
  XOR2_X1 U13417 ( .A1(n19726), .A2(n5081), .Z(n2501) );
  NAND3_X1 U13419 ( .A1(n31074), .A2(n19252), .A3(n1180), .ZN(n2867) );
  AOI21_X2 U13420 ( .A1(n2794), .A2(n22071), .B(n2502), .ZN(n15123) );
  OAI21_X2 U13432 ( .A1(n911), .A2(n21602), .B(n2513), .ZN(n8533) );
  NAND3_X2 U13438 ( .A1(n11261), .A2(n2519), .A3(n2518), .ZN(n15786) );
  NAND2_X1 U13441 ( .A1(n8756), .A2(n29309), .ZN(n2523) );
  XOR2_X1 U13445 ( .A1(n1024), .A2(n28864), .Z(n2525) );
  XOR2_X1 U13446 ( .A1(n3351), .A2(n507), .Z(n2526) );
  NAND2_X2 U13456 ( .A1(n2535), .A2(n16951), .ZN(n9320) );
  NOR2_X1 U13457 ( .A1(n10752), .A2(n1826), .ZN(n2534) );
  INV_X2 U13460 ( .I(n2978), .ZN(n6200) );
  NAND2_X2 U13461 ( .A1(n5270), .A2(n5271), .ZN(n2536) );
  NAND2_X2 U13468 ( .A1(n29258), .A2(n21462), .ZN(n6599) );
  XOR2_X1 U13470 ( .A1(n2556), .A2(n26124), .Z(n3782) );
  XOR2_X1 U13471 ( .A1(n2557), .A2(n11681), .Z(n2556) );
  XOR2_X1 U13474 ( .A1(n23293), .A2(n1194), .Z(n2564) );
  NOR2_X1 U13477 ( .A1(n7287), .A2(n23057), .ZN(n2580) );
  XOR2_X1 U13479 ( .A1(n15960), .A2(n16657), .Z(n11726) );
  OAI21_X2 U13480 ( .A1(n18841), .A2(n12052), .B(n2583), .ZN(n15960) );
  XOR2_X1 U13488 ( .A1(n20786), .A2(n5414), .Z(n2590) );
  XOR2_X1 U13489 ( .A1(n4681), .A2(n13491), .Z(n2591) );
  NOR2_X1 U13495 ( .A1(n29330), .A2(n13684), .ZN(n2960) );
  NOR2_X1 U13496 ( .A1(n29331), .A2(n13640), .ZN(n12885) );
  OAI22_X1 U13499 ( .A1(n25717), .A2(n29331), .B1(n1076), .B2(n6915), .ZN(
        n5784) );
  XOR2_X1 U13504 ( .A1(n17931), .A2(n19719), .Z(n2607) );
  XOR2_X1 U13506 ( .A1(n17430), .A2(n1370), .Z(n19719) );
  XOR2_X1 U13507 ( .A1(n19701), .A2(n467), .Z(n2608) );
  XOR2_X1 U13508 ( .A1(n28822), .A2(n2616), .Z(n12673) );
  OR2_X1 U13511 ( .A1(n31156), .A2(n7394), .Z(n2610) );
  XOR2_X1 U13519 ( .A1(n14588), .A2(n2611), .Z(n19519) );
  NAND2_X1 U13521 ( .A1(n18648), .A2(n18373), .ZN(n2613) );
  NAND2_X1 U13522 ( .A1(n18650), .A2(n2614), .ZN(n18549) );
  XOR2_X1 U13530 ( .A1(n31477), .A2(n16698), .Z(n13725) );
  XOR2_X1 U13531 ( .A1(n31477), .A2(n1416), .Z(n9762) );
  XOR2_X1 U13535 ( .A1(n31908), .A2(n478), .Z(n2626) );
  NAND4_X1 U13544 ( .A1(n5973), .A2(n5971), .A3(n22654), .A4(n11669), .ZN(
        n2632) );
  INV_X1 U13545 ( .I(n11669), .ZN(n2634) );
  OAI21_X2 U13556 ( .A1(n2646), .A2(n730), .B(n26600), .ZN(n3051) );
  XOR2_X1 U13558 ( .A1(n10522), .A2(n21017), .Z(n10437) );
  NAND2_X2 U13559 ( .A1(n2648), .A2(n2647), .ZN(n10522) );
  XOR2_X1 U13564 ( .A1(n23231), .A2(n540), .Z(n2651) );
  XOR2_X1 U13571 ( .A1(n11636), .A2(n7717), .Z(n2661) );
  XOR2_X1 U13581 ( .A1(n3694), .A2(n7603), .Z(n2666) );
  XOR2_X1 U13583 ( .A1(n7562), .A2(n24769), .Z(n2668) );
  XOR2_X1 U13585 ( .A1(n19712), .A2(n876), .Z(n2671) );
  OAI21_X2 U13589 ( .A1(n19339), .A2(n20000), .B(n7327), .ZN(n15005) );
  NAND2_X1 U13590 ( .A1(n20196), .A2(n2675), .ZN(n5103) );
  OAI21_X1 U13598 ( .A1(n31753), .A2(n18893), .B(n11941), .ZN(n2682) );
  OAI21_X1 U13607 ( .A1(n4045), .A2(n2694), .B(n2693), .ZN(n19847) );
  XOR2_X1 U13609 ( .A1(n2696), .A2(n2695), .Z(n8396) );
  XOR2_X1 U13610 ( .A1(n22268), .A2(n22057), .Z(n2695) );
  XOR2_X1 U13612 ( .A1(n24790), .A2(n1391), .Z(n2698) );
  XOR2_X1 U13620 ( .A1(n22289), .A2(n2707), .Z(n2917) );
  XOR2_X1 U13621 ( .A1(n343), .A2(n1390), .Z(n2707) );
  XOR2_X1 U13625 ( .A1(n2483), .A2(n12719), .Z(n12718) );
  XOR2_X1 U13626 ( .A1(n32822), .A2(n1415), .Z(n19427) );
  OAI21_X2 U13648 ( .A1(n18555), .A2(n3429), .B(n2731), .ZN(n9553) );
  XOR2_X1 U13657 ( .A1(Plaintext[28]), .A2(Key[28]), .Z(n11605) );
  XOR2_X1 U13659 ( .A1(n4134), .A2(n14668), .Z(n2739) );
  NAND2_X2 U13666 ( .A1(n10710), .A2(n13173), .ZN(n13232) );
  XOR2_X1 U13669 ( .A1(n31755), .A2(n19763), .Z(n2747) );
  NAND2_X2 U13675 ( .A1(n2754), .A2(n2753), .ZN(n20921) );
  XOR2_X1 U13683 ( .A1(n2759), .A2(n2757), .Z(n20054) );
  XOR2_X1 U13684 ( .A1(n19742), .A2(n2758), .Z(n2757) );
  XOR2_X1 U13685 ( .A1(n19768), .A2(n16525), .Z(n2758) );
  XOR2_X1 U13701 ( .A1(n15560), .A2(n624), .Z(n10076) );
  XOR2_X1 U13710 ( .A1(n2786), .A2(n2784), .Z(n20882) );
  XOR2_X1 U13716 ( .A1(n17837), .A2(n24527), .Z(n2788) );
  NAND2_X2 U13717 ( .A1(n2790), .A2(n12536), .ZN(n12535) );
  XOR2_X1 U13721 ( .A1(n19431), .A2(n17104), .Z(n19687) );
  XOR2_X1 U13722 ( .A1(n17835), .A2(n17834), .Z(n2796) );
  XOR2_X1 U13723 ( .A1(n28460), .A2(n16701), .Z(n23113) );
  AOI21_X2 U13726 ( .A1(n24385), .A2(n24384), .B(n24383), .ZN(n6484) );
  NAND2_X1 U13729 ( .A1(n31228), .A2(n27104), .ZN(n24384) );
  XOR2_X1 U13739 ( .A1(n9018), .A2(n23470), .Z(n2808) );
  NOR2_X2 U13748 ( .A1(n2813), .A2(n2844), .ZN(n23057) );
  XOR2_X1 U13754 ( .A1(n9629), .A2(n16551), .Z(n2818) );
  XOR2_X1 U13755 ( .A1(n4134), .A2(n20989), .Z(n2819) );
  NAND3_X2 U13760 ( .A1(n3461), .A2(n3465), .A3(n6536), .ZN(n2989) );
  AOI21_X1 U13764 ( .A1(n12966), .A2(n28376), .B(n2821), .ZN(n20505) );
  NOR2_X1 U13765 ( .A1(n2822), .A2(n1145), .ZN(n21418) );
  NAND2_X1 U13767 ( .A1(n28017), .A2(n2822), .ZN(n7121) );
  XOR2_X1 U13773 ( .A1(n22126), .A2(n25274), .Z(n2825) );
  XOR2_X1 U13784 ( .A1(n32467), .A2(n25274), .Z(n2838) );
  XOR2_X1 U13786 ( .A1(n2842), .A2(n2840), .Z(n16563) );
  XOR2_X1 U13787 ( .A1(n15055), .A2(n2841), .Z(n2840) );
  NAND3_X1 U13791 ( .A1(n14054), .A2(n15005), .A3(n2843), .ZN(n14546) );
  XOR2_X1 U13794 ( .A1(n2331), .A2(n34082), .Z(n3654) );
  XOR2_X1 U13796 ( .A1(n34082), .A2(n25619), .Z(n19391) );
  XOR2_X1 U13797 ( .A1(n3653), .A2(n3651), .Z(n9469) );
  NAND2_X1 U13815 ( .A1(n19143), .A2(n2869), .ZN(n2868) );
  NAND3_X1 U13819 ( .A1(n2876), .A2(n25007), .A3(n254), .ZN(n25004) );
  NAND2_X2 U13823 ( .A1(n3293), .A2(n3292), .ZN(n8374) );
  XOR2_X1 U13824 ( .A1(n2881), .A2(n2880), .Z(n2946) );
  XOR2_X1 U13825 ( .A1(n9569), .A2(n20837), .Z(n2880) );
  XOR2_X1 U13826 ( .A1(n21007), .A2(n21043), .Z(n9569) );
  XOR2_X1 U13831 ( .A1(n20813), .A2(n1193), .Z(n2883) );
  XOR2_X1 U13837 ( .A1(n2891), .A2(n2890), .Z(n2889) );
  XOR2_X1 U13838 ( .A1(n29652), .A2(n24964), .Z(n2890) );
  XOR2_X1 U13839 ( .A1(n9303), .A2(n20926), .Z(n2891) );
  XOR2_X1 U13848 ( .A1(n22158), .A2(n1067), .Z(n2898) );
  XOR2_X1 U13849 ( .A1(n2894), .A2(n4285), .Z(n2899) );
  NOR2_X1 U13858 ( .A1(n2901), .A2(n2902), .ZN(n10808) );
  OAI22_X1 U13859 ( .A1(n26640), .A2(n32253), .B1(n11940), .B2(n2902), .ZN(
        n19037) );
  INV_X1 U13863 ( .I(n2909), .ZN(n25026) );
  INV_X2 U13868 ( .I(n2915), .ZN(n13998) );
  XOR2_X1 U13871 ( .A1(n22118), .A2(n22115), .Z(n2918) );
  XOR2_X1 U13874 ( .A1(n2920), .A2(n16697), .Z(n19442) );
  XOR2_X1 U13879 ( .A1(n20974), .A2(n2925), .Z(n2924) );
  XOR2_X1 U13882 ( .A1(n20743), .A2(n8774), .Z(n2926) );
  INV_X2 U13891 ( .I(n2946), .ZN(n21237) );
  XOR2_X1 U13898 ( .A1(n13908), .A2(n13909), .Z(n2952) );
  NAND2_X1 U13907 ( .A1(n868), .A2(n2958), .ZN(n15951) );
  AOI21_X1 U13911 ( .A1(n25732), .A2(n6915), .B(n2959), .ZN(n5838) );
  NOR2_X1 U13912 ( .A1(n13124), .A2(n2960), .ZN(n2959) );
  NOR2_X2 U13915 ( .A1(n13637), .A2(n13636), .ZN(n13640) );
  XOR2_X1 U13926 ( .A1(n2972), .A2(n2975), .Z(n8634) );
  XOR2_X1 U13930 ( .A1(n30041), .A2(n23387), .Z(n23522) );
  XOR2_X1 U13931 ( .A1(n13190), .A2(n17704), .Z(n2975) );
  NAND2_X2 U13933 ( .A1(n3658), .A2(n4982), .ZN(n23441) );
  OAI21_X2 U13939 ( .A1(n8867), .A2(n8864), .B(n8863), .ZN(n19484) );
  NAND2_X2 U13941 ( .A1(n18717), .A2(n17617), .ZN(n19470) );
  OAI22_X1 U13943 ( .A1(n25006), .A2(n3019), .B1(n2983), .B2(n14865), .ZN(
        n25008) );
  NOR2_X1 U13952 ( .A1(n9090), .A2(n27142), .ZN(n2986) );
  XOR2_X1 U13953 ( .A1(n2989), .A2(n25722), .Z(n20644) );
  INV_X2 U13956 ( .I(n11599), .ZN(n11941) );
  NAND2_X1 U13968 ( .A1(n11680), .A2(n1331), .ZN(n3003) );
  XOR2_X1 U13978 ( .A1(n6484), .A2(n7256), .Z(n17571) );
  INV_X2 U13979 ( .I(n3012), .ZN(n8370) );
  NAND4_X1 U13980 ( .A1(n24333), .A2(n24334), .A3(n24332), .A4(n3014), .ZN(
        n24336) );
  NAND2_X2 U13984 ( .A1(n24880), .A2(n24879), .ZN(n3019) );
  NOR2_X2 U13990 ( .A1(n24083), .A2(n24082), .ZN(n24753) );
  NOR2_X2 U13993 ( .A1(n3024), .A2(n3023), .ZN(n9885) );
  XOR2_X1 U13995 ( .A1(n33293), .A2(n3027), .Z(n3026) );
  XOR2_X1 U13996 ( .A1(n7229), .A2(n30320), .Z(n3028) );
  INV_X1 U13999 ( .I(n3033), .ZN(n15013) );
  NAND2_X1 U14008 ( .A1(n3049), .A2(n3048), .ZN(n3047) );
  NOR2_X1 U14018 ( .A1(n20196), .A2(n295), .ZN(n3068) );
  XOR2_X1 U14020 ( .A1(n19549), .A2(n3071), .Z(n3070) );
  XOR2_X1 U14021 ( .A1(n19550), .A2(n25049), .Z(n3071) );
  XOR2_X1 U14023 ( .A1(n19699), .A2(n7971), .Z(n19549) );
  NAND2_X2 U14028 ( .A1(n16363), .A2(n19131), .ZN(n16727) );
  XOR2_X1 U14029 ( .A1(n19661), .A2(n19580), .Z(n19551) );
  XOR2_X1 U14038 ( .A1(n3081), .A2(n3082), .Z(n23586) );
  XOR2_X1 U14043 ( .A1(n1262), .A2(n27186), .Z(n3083) );
  XOR2_X1 U14050 ( .A1(n20984), .A2(n20986), .Z(n3099) );
  XOR2_X1 U14051 ( .A1(n17377), .A2(n3101), .Z(n3100) );
  XOR2_X1 U14052 ( .A1(n12495), .A2(n21985), .Z(n3102) );
  OAI21_X1 U14059 ( .A1(n17640), .A2(n26677), .B(n4971), .ZN(n3105) );
  XOR2_X1 U14068 ( .A1(n10443), .A2(n32880), .Z(n3109) );
  INV_X1 U14074 ( .I(n20781), .ZN(n20867) );
  XOR2_X1 U14078 ( .A1(n17517), .A2(n16390), .Z(n3118) );
  XOR2_X1 U14079 ( .A1(n21019), .A2(n15275), .Z(n3119) );
  XOR2_X1 U14081 ( .A1(n22203), .A2(n10165), .Z(n3120) );
  XNOR2_X1 U14091 ( .A1(n23200), .A2(n7772), .ZN(n23165) );
  XOR2_X1 U14092 ( .A1(n33465), .A2(n14435), .Z(n3126) );
  INV_X2 U14096 ( .I(n19222), .ZN(n15137) );
  XOR2_X1 U14102 ( .A1(n3134), .A2(n24964), .Z(Ciphertext[18]) );
  XOR2_X1 U14107 ( .A1(n22030), .A2(n22031), .Z(n3142) );
  XOR2_X1 U14108 ( .A1(n16321), .A2(n16472), .Z(n24595) );
  XOR2_X1 U14109 ( .A1(n16321), .A2(n1417), .Z(n24357) );
  XOR2_X1 U14111 ( .A1(n15308), .A2(n17384), .Z(n3143) );
  NAND3_X1 U14116 ( .A1(n3148), .A2(n24268), .A3(n31228), .ZN(n23996) );
  XOR2_X1 U14119 ( .A1(n20772), .A2(n3158), .Z(n4246) );
  XOR2_X1 U14120 ( .A1(n32399), .A2(n20992), .Z(n3158) );
  XOR2_X1 U14126 ( .A1(n17519), .A2(n3164), .Z(n14494) );
  XOR2_X1 U14127 ( .A1(n29011), .A2(n8356), .Z(n3164) );
  NAND2_X1 U14128 ( .A1(n29043), .A2(n3165), .ZN(n17588) );
  XOR2_X1 U14137 ( .A1(n7987), .A2(n6464), .Z(n10791) );
  NAND2_X1 U14140 ( .A1(n24780), .A2(n24874), .ZN(n24604) );
  XOR2_X1 U14141 ( .A1(n32467), .A2(n21037), .Z(n12171) );
  XOR2_X1 U14143 ( .A1(n22143), .A2(n21984), .Z(n3175) );
  XOR2_X1 U14145 ( .A1(n27240), .A2(n13091), .Z(n3177) );
  NAND2_X1 U14147 ( .A1(n8125), .A2(n3181), .ZN(n17589) );
  AND2_X1 U14149 ( .A1(n22537), .A2(n28170), .Z(n3189) );
  XOR2_X1 U14151 ( .A1(n21038), .A2(n6872), .Z(n3190) );
  XOR2_X1 U14152 ( .A1(n21039), .A2(n586), .Z(n3191) );
  XOR2_X1 U14155 ( .A1(n3194), .A2(n19413), .Z(n19414) );
  XOR2_X1 U14157 ( .A1(n11422), .A2(n22194), .Z(n11421) );
  NOR2_X1 U14161 ( .A1(n10831), .A2(n19856), .ZN(n3197) );
  XOR2_X1 U14162 ( .A1(n3199), .A2(n3198), .Z(n13298) );
  XOR2_X1 U14163 ( .A1(n13236), .A2(n1420), .Z(n3198) );
  XOR2_X1 U14164 ( .A1(n28579), .A2(n28939), .Z(n3199) );
  NAND2_X1 U14168 ( .A1(n30678), .A2(n3203), .ZN(n21536) );
  NAND2_X1 U14172 ( .A1(n24260), .A2(n30280), .ZN(n16573) );
  AOI21_X1 U14188 ( .A1(n18891), .A2(n18676), .B(n3218), .ZN(n12198) );
  NOR2_X1 U14189 ( .A1(n11398), .A2(n3218), .ZN(n11397) );
  AOI21_X1 U14190 ( .A1(n3586), .A2(n14874), .B(n3218), .ZN(n3516) );
  NOR2_X1 U14194 ( .A1(n9162), .A2(n9164), .ZN(n3224) );
  OAI21_X2 U14200 ( .A1(n17906), .A2(n3240), .B(n3239), .ZN(n24242) );
  NAND2_X2 U14202 ( .A1(n5083), .A2(n3242), .ZN(n6387) );
  NAND3_X2 U14203 ( .A1(n3245), .A2(n19173), .A3(n19172), .ZN(n19473) );
  NAND2_X1 U14208 ( .A1(n12508), .A2(n6111), .ZN(n25572) );
  XOR2_X1 U14213 ( .A1(n1363), .A2(n3258), .Z(n3358) );
  XOR2_X1 U14214 ( .A1(n3260), .A2(n3259), .Z(n3258) );
  XOR2_X1 U14217 ( .A1(n23399), .A2(n23398), .Z(n3267) );
  NAND2_X1 U14220 ( .A1(n4663), .A2(n31742), .ZN(n3271) );
  XOR2_X1 U14238 ( .A1(n11604), .A2(n34082), .Z(n19591) );
  XOR2_X1 U14242 ( .A1(n17912), .A2(n1084), .Z(n24401) );
  INV_X2 U14247 ( .I(n23853), .ZN(n8614) );
  OAI21_X2 U14251 ( .A1(n2537), .A2(n1300), .B(n6685), .ZN(n22856) );
  NAND3_X2 U14254 ( .A1(n25342), .A2(n25341), .A3(n25340), .ZN(n3300) );
  NOR2_X1 U14255 ( .A1(n3300), .A2(n25367), .ZN(n25362) );
  AOI21_X1 U14256 ( .A1(n25367), .A2(n25368), .B(n3300), .ZN(n25350) );
  NOR2_X1 U14257 ( .A1(n18711), .A2(n27142), .ZN(n11269) );
  XOR2_X1 U14262 ( .A1(n3350), .A2(n1407), .Z(n20621) );
  XOR2_X1 U14263 ( .A1(n3350), .A2(n7705), .Z(n20798) );
  XOR2_X1 U14264 ( .A1(n3350), .A2(n30543), .Z(n13093) );
  INV_X2 U14266 ( .I(n13189), .ZN(n15522) );
  XOR2_X1 U14272 ( .A1(n438), .A2(n32796), .Z(n3319) );
  OAI21_X2 U14276 ( .A1(n3324), .A2(n29232), .B(n11865), .ZN(n15243) );
  XOR2_X1 U14279 ( .A1(n30041), .A2(n14613), .Z(n13777) );
  NAND2_X1 U14288 ( .A1(n18538), .A2(n3344), .ZN(n14327) );
  XOR2_X1 U14291 ( .A1(n3345), .A2(n31416), .Z(n24552) );
  XOR2_X1 U14292 ( .A1(n33700), .A2(n24804), .Z(n14532) );
  NAND2_X2 U14296 ( .A1(n4234), .A2(n13113), .ZN(n21839) );
  XOR2_X1 U14298 ( .A1(n3355), .A2(n3354), .Z(n3353) );
  XOR2_X1 U14299 ( .A1(n29121), .A2(n1421), .Z(n3354) );
  XOR2_X1 U14300 ( .A1(n12789), .A2(n7808), .Z(n3355) );
  OAI21_X2 U14302 ( .A1(n7516), .A2(n10125), .B(n3361), .ZN(n10124) );
  XOR2_X1 U14305 ( .A1(n22187), .A2(n3369), .Z(n3368) );
  XOR2_X1 U14306 ( .A1(n16060), .A2(n25910), .Z(n3369) );
  NAND3_X2 U14309 ( .A1(n3384), .A2(n32031), .A3(n3382), .ZN(n6798) );
  INV_X2 U14314 ( .I(n3392), .ZN(n4396) );
  XOR2_X1 U14316 ( .A1(n30571), .A2(n27920), .Z(n3396) );
  XOR2_X1 U14319 ( .A1(n19716), .A2(n10123), .Z(n3399) );
  XOR2_X1 U14324 ( .A1(n21045), .A2(n20967), .Z(n4260) );
  NOR2_X1 U14327 ( .A1(n3405), .A2(n25564), .ZN(n24460) );
  OAI21_X2 U14332 ( .A1(n1260), .A2(n9843), .B(n3408), .ZN(n4955) );
  XOR2_X1 U14336 ( .A1(n4955), .A2(n23386), .Z(n3410) );
  XOR2_X1 U14337 ( .A1(n3412), .A2(n537), .Z(n3411) );
  XOR2_X1 U14338 ( .A1(n27220), .A2(n5514), .Z(n3412) );
  XOR2_X1 U14342 ( .A1(n26623), .A2(n25218), .Z(n3415) );
  XOR2_X1 U14346 ( .A1(n13477), .A2(n3417), .Z(n19705) );
  XOR2_X1 U14348 ( .A1(n22119), .A2(n30993), .Z(n22120) );
  AND2_X1 U14355 ( .A1(n20419), .A2(n15005), .Z(n3428) );
  INV_X1 U14356 ( .I(n3430), .ZN(n10745) );
  XOR2_X1 U14357 ( .A1(n3431), .A2(n25192), .Z(Ciphertext[68]) );
  OAI21_X1 U14358 ( .A1(n10574), .A2(n27149), .B(n3433), .ZN(n3432) );
  NOR2_X1 U14372 ( .A1(n632), .A2(n14339), .ZN(n3502) );
  MUX2_X1 U14374 ( .I0(n809), .I1(n30065), .S(n14227), .Z(n22448) );
  XOR2_X1 U14376 ( .A1(n24749), .A2(n3477), .Z(n3476) );
  XOR2_X1 U14377 ( .A1(n24839), .A2(n25864), .Z(n3477) );
  NOR2_X1 U14389 ( .A1(n30318), .A2(n3489), .ZN(n5301) );
  NAND2_X1 U14390 ( .A1(n5408), .A2(n3489), .ZN(n5407) );
  XOR2_X1 U14394 ( .A1(n16998), .A2(n18015), .Z(n3493) );
  NAND2_X1 U14396 ( .A1(n26292), .A2(n3495), .ZN(n11420) );
  NAND2_X1 U14399 ( .A1(n31197), .A2(n32898), .ZN(n3497) );
  XOR2_X1 U14404 ( .A1(n10422), .A2(n10421), .Z(n16710) );
  XOR2_X1 U14410 ( .A1(n3514), .A2(n23535), .Z(n9983) );
  XOR2_X1 U14418 ( .A1(n23183), .A2(n26656), .Z(n23494) );
  NAND3_X1 U14435 ( .A1(n21781), .A2(n31220), .A3(n3539), .ZN(n21746) );
  XOR2_X1 U14439 ( .A1(n11217), .A2(n3541), .Z(n3540) );
  XOR2_X1 U14440 ( .A1(n17301), .A2(n8139), .Z(n3541) );
  XOR2_X1 U14442 ( .A1(n5932), .A2(n24652), .Z(n24824) );
  XOR2_X1 U14449 ( .A1(n20747), .A2(n1191), .Z(n3559) );
  NAND2_X1 U14454 ( .A1(n3567), .A2(n31019), .ZN(n17631) );
  NOR2_X1 U14456 ( .A1(n22406), .A2(n3567), .ZN(n3566) );
  INV_X1 U14457 ( .I(n3569), .ZN(n12159) );
  NAND3_X1 U14458 ( .A1(n3570), .A2(n22982), .A3(n22983), .ZN(n22984) );
  NOR2_X1 U14460 ( .A1(n22800), .A2(n3570), .ZN(n13045) );
  XOR2_X1 U14465 ( .A1(n23375), .A2(n23294), .Z(n23240) );
  NAND2_X2 U14466 ( .A1(n16993), .A2(n11837), .ZN(n23294) );
  NAND2_X2 U14468 ( .A1(n15208), .A2(n17175), .ZN(n16373) );
  XOR2_X1 U14470 ( .A1(n23343), .A2(n3575), .Z(n3574) );
  XOR2_X1 U14471 ( .A1(n15183), .A2(n16602), .Z(n3575) );
  XOR2_X1 U14483 ( .A1(n22139), .A2(n16390), .Z(n3583) );
  XOR2_X1 U14487 ( .A1(n27186), .A2(n12797), .Z(n10776) );
  XOR2_X1 U14488 ( .A1(n27186), .A2(n9223), .Z(n7131) );
  AOI21_X2 U14491 ( .A1(n19074), .A2(n29398), .B(n19073), .ZN(n3599) );
  XOR2_X1 U14497 ( .A1(n17918), .A2(n3606), .Z(n3605) );
  XOR2_X1 U14498 ( .A1(n8617), .A2(n16525), .Z(n3606) );
  XOR2_X1 U14500 ( .A1(n33468), .A2(n16598), .Z(n12624) );
  INV_X2 U14508 ( .I(n20788), .ZN(n20907) );
  XOR2_X1 U14511 ( .A1(n3621), .A2(n3622), .Z(n3618) );
  XOR2_X1 U14514 ( .A1(n23461), .A2(n23321), .Z(n3620) );
  XOR2_X1 U14516 ( .A1(n30322), .A2(n15114), .Z(n3622) );
  XOR2_X1 U14520 ( .A1(n3628), .A2(n20894), .Z(n3627) );
  XOR2_X1 U14521 ( .A1(n20992), .A2(n1069), .Z(n3628) );
  XOR2_X1 U14527 ( .A1(n3634), .A2(n25541), .Z(n9269) );
  XOR2_X1 U14543 ( .A1(n11762), .A2(n10278), .Z(n3648) );
  XOR2_X1 U14544 ( .A1(n3652), .A2(n18031), .Z(n3651) );
  XOR2_X1 U14545 ( .A1(n3815), .A2(n3654), .Z(n3653) );
  AOI21_X1 U14546 ( .A1(n17055), .A2(n15475), .B(n25996), .ZN(n15474) );
  MUX2_X1 U14549 ( .I0(n30769), .I1(n30885), .S(n21697), .Z(n3656) );
  NAND2_X2 U14550 ( .A1(n18136), .A2(n12133), .ZN(n21697) );
  AND2_X1 U14553 ( .A1(n33627), .A2(n29446), .Z(n4301) );
  XOR2_X1 U14555 ( .A1(n19620), .A2(n5919), .Z(n3665) );
  NAND2_X1 U14561 ( .A1(n5821), .A2(n3668), .ZN(n22750) );
  XOR2_X1 U14571 ( .A1(n24552), .A2(n3677), .Z(n4302) );
  XOR2_X1 U14572 ( .A1(n8949), .A2(n5268), .Z(n3677) );
  XOR2_X1 U14576 ( .A1(n21945), .A2(n3682), .Z(n3683) );
  INV_X2 U14577 ( .I(n3686), .ZN(n9172) );
  NOR2_X1 U14578 ( .A1(n17694), .A2(n3687), .ZN(n13879) );
  NAND2_X2 U14579 ( .A1(n22496), .A2(n22495), .ZN(n14686) );
  XOR2_X1 U14585 ( .A1(n3694), .A2(n2864), .Z(n9093) );
  XOR2_X1 U14591 ( .A1(n3704), .A2(n17555), .Z(n22300) );
  XOR2_X1 U14594 ( .A1(n9536), .A2(n3704), .Z(n9532) );
  XOR2_X1 U14597 ( .A1(n12342), .A2(n3705), .Z(n20242) );
  XOR2_X1 U14598 ( .A1(n20726), .A2(n3705), .Z(n21027) );
  NAND2_X2 U14599 ( .A1(n15142), .A2(n20237), .ZN(n3705) );
  OAI21_X2 U14609 ( .A1(n11991), .A2(n918), .B(n11856), .ZN(n3723) );
  XOR2_X1 U14617 ( .A1(n3727), .A2(n19679), .Z(n9819) );
  NAND2_X1 U14618 ( .A1(n5433), .A2(n502), .ZN(n4841) );
  NAND2_X2 U14620 ( .A1(n3730), .A2(n3728), .ZN(n6402) );
  INV_X2 U14621 ( .I(n18080), .ZN(n25236) );
  XOR2_X1 U14623 ( .A1(n30219), .A2(n24231), .Z(n3735) );
  XOR2_X1 U14624 ( .A1(n14858), .A2(n16173), .Z(n12618) );
  XOR2_X1 U14625 ( .A1(n20870), .A2(n3737), .Z(n3736) );
  XOR2_X1 U14626 ( .A1(n21040), .A2(n5772), .Z(n3737) );
  XOR2_X1 U14634 ( .A1(n24469), .A2(n17753), .Z(n17752) );
  AOI22_X2 U14639 ( .A1(n24378), .A2(n14547), .B1(n25753), .B2(n25581), .ZN(
        n25746) );
  NOR2_X1 U14643 ( .A1(n12906), .A2(n12948), .ZN(n9391) );
  NAND2_X2 U14647 ( .A1(n23792), .A2(n23791), .ZN(n12493) );
  INV_X2 U14654 ( .I(n3755), .ZN(n10182) );
  XOR2_X1 U14655 ( .A1(Plaintext[174]), .A2(Key[174]), .Z(n3755) );
  XOR2_X1 U14657 ( .A1(n4240), .A2(n16642), .Z(n24794) );
  NOR3_X2 U14663 ( .A1(n26025), .A2(n15466), .A3(n14098), .ZN(n8530) );
  XOR2_X1 U14667 ( .A1(n17524), .A2(n20514), .Z(n21442) );
  NAND2_X2 U14673 ( .A1(n20651), .A2(n20650), .ZN(n20769) );
  AOI21_X2 U14674 ( .A1(n2565), .A2(n20438), .B(n17424), .ZN(n20651) );
  NAND2_X1 U14679 ( .A1(n20501), .A2(n20502), .ZN(n16758) );
  OAI21_X1 U14682 ( .A1(n25349), .A2(n25360), .B(n25379), .ZN(n3771) );
  OR2_X1 U14683 ( .A1(n25350), .A2(n25361), .Z(n3772) );
  XOR2_X1 U14686 ( .A1(n24848), .A2(n17448), .Z(n5022) );
  XOR2_X1 U14693 ( .A1(n4915), .A2(n23245), .Z(n3777) );
  NAND2_X1 U14694 ( .A1(n4066), .A2(n14811), .ZN(n16007) );
  OAI21_X2 U14695 ( .A1(n4178), .A2(n5752), .B(n5751), .ZN(n4066) );
  XNOR2_X1 U14696 ( .A1(n13309), .A2(n11803), .ZN(n4004) );
  INV_X2 U14705 ( .I(n3782), .ZN(n11820) );
  AND2_X1 U14707 ( .A1(n25174), .A2(n25175), .Z(n8931) );
  NAND2_X2 U14708 ( .A1(n25172), .A2(n25169), .ZN(n25174) );
  NAND2_X1 U14718 ( .A1(n3788), .A2(n1425), .ZN(n14295) );
  XOR2_X1 U14730 ( .A1(Plaintext[116]), .A2(Key[116]), .Z(n18131) );
  XOR2_X1 U14731 ( .A1(n23220), .A2(n23198), .Z(n11144) );
  OAI21_X1 U14736 ( .A1(n14830), .A2(n22636), .B(n12043), .ZN(n22495) );
  XOR2_X1 U14748 ( .A1(n8656), .A2(n24050), .Z(n9968) );
  XOR2_X1 U14757 ( .A1(n9200), .A2(n660), .Z(n9199) );
  XOR2_X1 U14759 ( .A1(n23189), .A2(n4409), .Z(n23465) );
  XOR2_X1 U14761 ( .A1(n24533), .A2(n27950), .Z(n16891) );
  AND2_X1 U14762 ( .A1(n23660), .A2(n30252), .Z(n4350) );
  NAND2_X1 U14766 ( .A1(n32884), .A2(n32798), .ZN(n15867) );
  XOR2_X1 U14771 ( .A1(n24439), .A2(n3809), .Z(n11527) );
  XOR2_X1 U14772 ( .A1(n24592), .A2(n25364), .Z(n3809) );
  INV_X2 U14780 ( .I(n3816), .ZN(n11333) );
  NAND2_X1 U14783 ( .A1(n9469), .A2(n563), .ZN(n12119) );
  XOR2_X1 U14784 ( .A1(n3819), .A2(n12672), .Z(n8545) );
  XOR2_X1 U14785 ( .A1(n20796), .A2(n20797), .Z(n3819) );
  XOR2_X1 U14786 ( .A1(n21025), .A2(n6561), .Z(n6560) );
  NAND2_X2 U14789 ( .A1(n9237), .A2(n9238), .ZN(n14293) );
  AOI21_X1 U14794 ( .A1(n832), .A2(n27189), .B(n7038), .ZN(n7037) );
  OAI21_X2 U14797 ( .A1(n14693), .A2(n19889), .B(n3827), .ZN(n20485) );
  XNOR2_X1 U14801 ( .A1(n11481), .A2(n5848), .ZN(n9673) );
  XOR2_X1 U14803 ( .A1(n15708), .A2(n19552), .Z(n19555) );
  XOR2_X1 U14823 ( .A1(n23370), .A2(n16300), .Z(n6152) );
  XOR2_X1 U14824 ( .A1(n8630), .A2(n22301), .Z(n12828) );
  XOR2_X1 U14825 ( .A1(n4723), .A2(n15825), .Z(n22301) );
  NAND2_X1 U14826 ( .A1(n21594), .A2(n21145), .ZN(n21156) );
  NOR2_X1 U14828 ( .A1(n6778), .A2(n33621), .ZN(n6579) );
  OAI21_X2 U14837 ( .A1(n15675), .A2(n6009), .B(n3920), .ZN(n19778) );
  NOR2_X1 U14863 ( .A1(n13733), .A2(n24229), .ZN(n13732) );
  XOR2_X1 U14864 ( .A1(n23315), .A2(n13812), .Z(n11416) );
  XOR2_X1 U14866 ( .A1(n20600), .A2(n5209), .Z(n16239) );
  NAND2_X2 U14869 ( .A1(n414), .A2(n5834), .ZN(n18682) );
  XOR2_X1 U14887 ( .A1(n23385), .A2(n17188), .Z(n23284) );
  NAND2_X2 U14893 ( .A1(n6206), .A2(n6570), .ZN(n6571) );
  XOR2_X1 U14897 ( .A1(n14908), .A2(n26623), .Z(n3870) );
  OR2_X1 U14900 ( .A1(n24712), .A2(n4490), .Z(n4451) );
  XOR2_X1 U14904 ( .A1(n11221), .A2(n11220), .Z(n19958) );
  NAND2_X2 U14905 ( .A1(n21827), .A2(n21824), .ZN(n5170) );
  XNOR2_X1 U14912 ( .A1(n23203), .A2(n24917), .ZN(n4466) );
  NAND2_X1 U14913 ( .A1(n23690), .A2(n23856), .ZN(n17056) );
  XOR2_X1 U14921 ( .A1(n3884), .A2(n14206), .Z(n14296) );
  NAND2_X1 U14922 ( .A1(n14295), .A2(n14294), .ZN(n3884) );
  XOR2_X1 U14924 ( .A1(n12491), .A2(n30320), .Z(n9012) );
  INV_X1 U14928 ( .I(n4342), .ZN(n22188) );
  AOI21_X2 U14932 ( .A1(n18334), .A2(n3893), .B(n18333), .ZN(n16847) );
  XOR2_X1 U14933 ( .A1(n7184), .A2(n446), .Z(n16105) );
  XOR2_X1 U14943 ( .A1(n17565), .A2(n23320), .Z(n23194) );
  XOR2_X1 U14946 ( .A1(n10200), .A2(n3896), .Z(n17779) );
  XOR2_X1 U14947 ( .A1(n14779), .A2(n24098), .Z(n3896) );
  NAND2_X2 U14948 ( .A1(n7770), .A2(n7768), .ZN(n25107) );
  NAND3_X2 U14955 ( .A1(n3900), .A2(n5333), .A3(n19136), .ZN(n19773) );
  INV_X1 U14956 ( .I(n23446), .ZN(n17350) );
  AND2_X1 U14959 ( .A1(n4405), .A2(n7810), .Z(n19174) );
  XOR2_X1 U14961 ( .A1(n3905), .A2(n17457), .Z(n8834) );
  AND2_X1 U14963 ( .A1(n6483), .A2(n3467), .Z(n8970) );
  NAND2_X2 U14971 ( .A1(n3908), .A2(n12939), .ZN(n22291) );
  NAND2_X1 U14973 ( .A1(n19863), .A2(n10335), .ZN(n7922) );
  XOR2_X1 U14974 ( .A1(n9326), .A2(n9325), .Z(n10335) );
  INV_X1 U14979 ( .I(n25882), .ZN(n7274) );
  AND2_X1 U14980 ( .A1(n25882), .A2(n25879), .Z(n7268) );
  XNOR2_X1 U14985 ( .A1(n21281), .A2(n21280), .ZN(n9593) );
  NOR2_X1 U14992 ( .A1(n19799), .A2(n16625), .ZN(n19800) );
  INV_X2 U14995 ( .I(n9992), .ZN(n11887) );
  NAND2_X2 U14998 ( .A1(n13461), .A2(n13462), .ZN(n23066) );
  XOR2_X1 U15004 ( .A1(n23220), .A2(n3923), .Z(n8488) );
  XOR2_X1 U15005 ( .A1(n27252), .A2(n31354), .Z(n3923) );
  XNOR2_X1 U15006 ( .A1(n15341), .A2(n27763), .ZN(n14733) );
  NOR2_X1 U15010 ( .A1(n21066), .A2(n31965), .ZN(n6213) );
  XNOR2_X1 U15012 ( .A1(n28262), .A2(n16551), .ZN(n10878) );
  NAND2_X1 U15018 ( .A1(n8966), .A2(n3926), .ZN(n14465) );
  AOI21_X1 U15019 ( .A1(n5035), .A2(n6593), .B(n22957), .ZN(n3926) );
  NAND2_X2 U15021 ( .A1(n23989), .A2(n13144), .ZN(n7511) );
  NOR2_X1 U15025 ( .A1(n5842), .A2(n18945), .ZN(n18946) );
  NAND2_X2 U15027 ( .A1(n24217), .A2(n29010), .ZN(n23964) );
  NAND2_X2 U15028 ( .A1(n14966), .A2(n14965), .ZN(n6906) );
  XOR2_X1 U15035 ( .A1(n5881), .A2(n3938), .Z(n5880) );
  XOR2_X1 U15036 ( .A1(n5882), .A2(n524), .Z(n3938) );
  NAND2_X1 U15067 ( .A1(n6234), .A2(n694), .ZN(n16661) );
  XOR2_X1 U15071 ( .A1(Plaintext[9]), .A2(Key[9]), .Z(n3954) );
  AOI21_X1 U15072 ( .A1(n5113), .A2(n24994), .B(n9901), .ZN(n9903) );
  INV_X2 U15074 ( .I(n10725), .ZN(n16166) );
  XOR2_X1 U15078 ( .A1(n24846), .A2(n7256), .Z(n24849) );
  XOR2_X1 U15082 ( .A1(n20757), .A2(n20712), .Z(n20713) );
  XOR2_X1 U15085 ( .A1(n10109), .A2(n15562), .Z(n3957) );
  XOR2_X1 U15086 ( .A1(n3958), .A2(n9487), .Z(n9486) );
  XOR2_X1 U15087 ( .A1(n24778), .A2(n550), .Z(n3958) );
  XOR2_X1 U15088 ( .A1(n20852), .A2(n10159), .Z(n15630) );
  OAI22_X2 U15090 ( .A1(n21602), .A2(n21716), .B1(n21710), .B2(n21712), .ZN(
        n6462) );
  XOR2_X1 U15093 ( .A1(n6169), .A2(n15653), .Z(n16300) );
  OAI22_X2 U15104 ( .A1(n3963), .A2(n21298), .B1(n4989), .B2(n21199), .ZN(
        n21870) );
  XOR2_X1 U15106 ( .A1(n24634), .A2(n24494), .Z(n10945) );
  XOR2_X1 U15108 ( .A1(n20899), .A2(n9706), .Z(n10951) );
  NAND2_X2 U15114 ( .A1(n964), .A2(n5072), .ZN(n9481) );
  OAI22_X2 U15124 ( .A1(n19060), .A2(n1179), .B1(n4366), .B2(n16185), .ZN(
        n4150) );
  NAND2_X1 U15137 ( .A1(n22832), .A2(n13635), .ZN(n12156) );
  XOR2_X1 U15140 ( .A1(n16259), .A2(n23433), .Z(n17285) );
  XOR2_X1 U15146 ( .A1(n9528), .A2(n3980), .Z(n10934) );
  XOR2_X1 U15148 ( .A1(n3981), .A2(n444), .Z(n5074) );
  XOR2_X1 U15149 ( .A1(n4984), .A2(n15788), .Z(n3981) );
  INV_X1 U15150 ( .I(n19523), .ZN(n20141) );
  NAND2_X1 U15151 ( .A1(n27110), .A2(n15237), .ZN(n19523) );
  AND2_X1 U15157 ( .A1(n10182), .A2(n11460), .Z(n18877) );
  OR2_X1 U15159 ( .A1(n7465), .A2(n13334), .Z(n5490) );
  NAND2_X2 U15165 ( .A1(n3985), .A2(n12814), .ZN(n16699) );
  XOR2_X1 U15169 ( .A1(n20752), .A2(n3990), .Z(n18050) );
  XOR2_X1 U15170 ( .A1(n4618), .A2(n24804), .Z(n3990) );
  OAI21_X2 U15180 ( .A1(n3996), .A2(n3995), .B(n4675), .ZN(n24002) );
  OR2_X1 U15181 ( .A1(n4734), .A2(n23065), .Z(n3997) );
  XOR2_X1 U15186 ( .A1(n20759), .A2(n16191), .Z(n4000) );
  AND2_X1 U15197 ( .A1(n1278), .A2(n15633), .Z(n12218) );
  OR2_X1 U15209 ( .A1(n1430), .A2(n10080), .Z(n4008) );
  XOR2_X1 U15212 ( .A1(n4013), .A2(n13067), .Z(n10186) );
  INV_X1 U15216 ( .I(n24870), .ZN(n16607) );
  XOR2_X1 U15217 ( .A1(n4015), .A2(n9607), .Z(n9606) );
  XOR2_X1 U15218 ( .A1(n9608), .A2(n21007), .Z(n4015) );
  XOR2_X1 U15229 ( .A1(n5939), .A2(n14122), .Z(n4020) );
  XOR2_X1 U15238 ( .A1(n30327), .A2(n5539), .Z(n14779) );
  NAND2_X2 U15240 ( .A1(n4628), .A2(n4629), .ZN(n4599) );
  XOR2_X1 U15249 ( .A1(n4035), .A2(n16423), .Z(Ciphertext[29]) );
  AOI22_X1 U15259 ( .A1(n17165), .A2(n17687), .B1(n17166), .B2(n18863), .ZN(
        n12193) );
  NOR2_X2 U15261 ( .A1(n19816), .A2(n19817), .ZN(n20595) );
  OR2_X1 U15262 ( .A1(n10413), .A2(n19891), .Z(n17443) );
  XOR2_X1 U15268 ( .A1(n19695), .A2(n4042), .Z(n20088) );
  XOR2_X1 U15269 ( .A1(n19693), .A2(n19694), .Z(n4042) );
  XOR2_X1 U15286 ( .A1(n4052), .A2(n496), .Z(n8684) );
  XOR2_X1 U15294 ( .A1(n21035), .A2(n1409), .Z(n20929) );
  XOR2_X1 U15299 ( .A1(n23124), .A2(n481), .Z(n4059) );
  OR2_X1 U15303 ( .A1(n21707), .A2(n230), .Z(n14461) );
  NAND2_X2 U15309 ( .A1(n5801), .A2(n4062), .ZN(n4646) );
  XOR2_X1 U15311 ( .A1(n4063), .A2(n27126), .Z(n7381) );
  NAND2_X1 U15315 ( .A1(n24882), .A2(n25117), .ZN(n4065) );
  NOR2_X1 U15337 ( .A1(n14544), .A2(n14543), .ZN(n10128) );
  NAND2_X1 U15339 ( .A1(n4177), .A2(n23855), .ZN(n23800) );
  OAI21_X2 U15340 ( .A1(n8800), .A2(n18925), .B(n18924), .ZN(n19632) );
  AND2_X1 U15342 ( .A1(n23949), .A2(n11676), .Z(n9002) );
  NAND2_X1 U15343 ( .A1(n11623), .A2(n2635), .ZN(n5233) );
  XOR2_X1 U15347 ( .A1(n15308), .A2(n24387), .Z(n4419) );
  AND2_X1 U15351 ( .A1(n25867), .A2(n25897), .Z(n8780) );
  XOR2_X1 U15354 ( .A1(Plaintext[189]), .A2(Key[189]), .Z(n5594) );
  INV_X1 U15356 ( .I(n23705), .ZN(n4086) );
  OAI21_X1 U15360 ( .A1(n25375), .A2(n30276), .B(n4089), .ZN(n25357) );
  XOR2_X1 U15363 ( .A1(n11836), .A2(n11835), .Z(n11834) );
  XOR2_X1 U15365 ( .A1(n24593), .A2(n4091), .Z(n5429) );
  XOR2_X1 U15366 ( .A1(n24645), .A2(n28898), .Z(n4091) );
  NAND2_X1 U15375 ( .A1(n28825), .A2(n8846), .ZN(n5814) );
  INV_X1 U15379 ( .I(n16596), .ZN(n18779) );
  NAND2_X2 U15395 ( .A1(n1337), .A2(n9678), .ZN(n8041) );
  XOR2_X1 U15396 ( .A1(n1227), .A2(n4112), .Z(n15484) );
  XOR2_X1 U15397 ( .A1(n27151), .A2(n25856), .Z(n4112) );
  XOR2_X1 U15407 ( .A1(n24424), .A2(n24425), .Z(n6726) );
  XOR2_X1 U15408 ( .A1(n24416), .A2(n24796), .Z(n24425) );
  BUF_X2 U15410 ( .I(n8190), .Z(n4119) );
  OAI21_X1 U15420 ( .A1(n27619), .A2(n27336), .B(n12028), .ZN(n21549) );
  XOR2_X1 U15436 ( .A1(n23441), .A2(n17871), .Z(n4559) );
  INV_X2 U15440 ( .I(n4133), .ZN(n20156) );
  INV_X1 U15451 ( .I(n6259), .ZN(n12570) );
  NAND2_X1 U15452 ( .A1(n12570), .A2(n25197), .ZN(n4533) );
  XOR2_X1 U15457 ( .A1(n7731), .A2(n30540), .Z(n24629) );
  AOI22_X2 U15461 ( .A1(n8461), .A2(n18422), .B1(n18616), .B2(n17224), .ZN(
        n14811) );
  XOR2_X1 U15478 ( .A1(n22799), .A2(n4154), .Z(n14381) );
  XOR2_X1 U15479 ( .A1(n13347), .A2(n15941), .Z(n4154) );
  NOR2_X1 U15485 ( .A1(n12930), .A2(n12931), .ZN(n9502) );
  OAI21_X1 U15486 ( .A1(n917), .A2(n916), .B(n9898), .ZN(n9897) );
  NAND2_X1 U15487 ( .A1(n9897), .A2(n9896), .ZN(n9895) );
  OAI22_X2 U15488 ( .A1(n18647), .A2(n5456), .B1(n10125), .B2(n17792), .ZN(
        n5455) );
  XOR2_X1 U15490 ( .A1(n11860), .A2(n11859), .Z(n4158) );
  XNOR2_X1 U15491 ( .A1(n22273), .A2(n21931), .ZN(n6543) );
  INV_X1 U15493 ( .I(n10404), .ZN(n4456) );
  NAND2_X1 U15512 ( .A1(n15043), .A2(n15169), .ZN(n20341) );
  INV_X1 U15515 ( .I(n18002), .ZN(n4168) );
  NOR2_X1 U15525 ( .A1(n8207), .A2(n25179), .ZN(n8932) );
  NAND2_X2 U15528 ( .A1(n21867), .A2(n13652), .ZN(n21863) );
  INV_X1 U15530 ( .I(n20015), .ZN(n4893) );
  XOR2_X1 U15532 ( .A1(n8921), .A2(n19702), .Z(n7184) );
  XOR2_X1 U15533 ( .A1(n18911), .A2(n19743), .Z(n19702) );
  XOR2_X1 U15534 ( .A1(n14743), .A2(n14744), .Z(n17821) );
  XOR2_X1 U15536 ( .A1(n5702), .A2(n533), .Z(n4173) );
  AOI21_X2 U15539 ( .A1(n23818), .A2(n23819), .B(n23817), .ZN(n24327) );
  XOR2_X1 U15547 ( .A1(n4176), .A2(n19512), .Z(n16646) );
  XOR2_X1 U15548 ( .A1(n12801), .A2(n12683), .Z(n4176) );
  INV_X2 U15553 ( .I(n4180), .ZN(n11958) );
  XNOR2_X1 U15554 ( .A1(n17356), .A2(n17355), .ZN(n4180) );
  XOR2_X1 U15557 ( .A1(n6316), .A2(n10901), .Z(n10900) );
  XOR2_X1 U15559 ( .A1(n14833), .A2(n4187), .Z(n4186) );
  XOR2_X1 U15573 ( .A1(n8682), .A2(n4196), .Z(n8681) );
  XOR2_X1 U15574 ( .A1(n11783), .A2(n15936), .Z(n4196) );
  NAND3_X2 U15578 ( .A1(n24856), .A2(n7853), .A3(n7854), .ZN(n25082) );
  INV_X2 U15583 ( .I(n4200), .ZN(n18349) );
  XOR2_X1 U15587 ( .A1(n20723), .A2(n20859), .Z(n16803) );
  NAND2_X1 U15590 ( .A1(n4447), .A2(n9181), .ZN(n25814) );
  NAND2_X2 U15604 ( .A1(n6010), .A2(n8667), .ZN(n23111) );
  XOR2_X1 U15609 ( .A1(n19594), .A2(n463), .Z(n5138) );
  XNOR2_X1 U15613 ( .A1(n23249), .A2(n23450), .ZN(n5263) );
  INV_X2 U15614 ( .I(n4224), .ZN(n4373) );
  XOR2_X1 U15616 ( .A1(n21044), .A2(n27169), .Z(n9607) );
  NOR2_X1 U15619 ( .A1(n16440), .A2(n21338), .ZN(n7115) );
  AOI21_X2 U15633 ( .A1(n18084), .A2(n4232), .B(n24364), .ZN(n24910) );
  INV_X1 U15636 ( .I(n21146), .ZN(n4865) );
  NAND2_X1 U15639 ( .A1(n22645), .A2(n10724), .ZN(n13973) );
  INV_X2 U15641 ( .I(n4243), .ZN(n11045) );
  AOI21_X2 U15645 ( .A1(n24301), .A2(n24302), .B(n24306), .ZN(n24645) );
  OR2_X1 U15649 ( .A1(n18800), .A2(n8395), .Z(n4255) );
  XOR2_X1 U15650 ( .A1(n24281), .A2(n24280), .Z(n11717) );
  NAND3_X1 U15663 ( .A1(n7855), .A2(n16632), .A3(n15254), .ZN(n7853) );
  AOI21_X1 U15664 ( .A1(n5908), .A2(n12194), .B(n1346), .ZN(n4261) );
  XOR2_X1 U15668 ( .A1(n20762), .A2(n26058), .Z(n4263) );
  XOR2_X1 U15678 ( .A1(n8488), .A2(n9993), .Z(n9992) );
  XOR2_X1 U15685 ( .A1(n23441), .A2(n23368), .Z(n4273) );
  XOR2_X1 U15687 ( .A1(n24416), .A2(n30540), .Z(n12067) );
  OR2_X1 U15694 ( .A1(n10335), .A2(n568), .Z(n17060) );
  XOR2_X1 U15696 ( .A1(n8214), .A2(n4280), .Z(n9239) );
  XOR2_X1 U15697 ( .A1(n24371), .A2(n9241), .Z(n4280) );
  XOR2_X1 U15704 ( .A1(n32860), .A2(n12491), .Z(n11551) );
  XOR2_X1 U15705 ( .A1(n24847), .A2(n10084), .Z(n24541) );
  OR2_X1 U15712 ( .A1(n20575), .A2(n20574), .Z(n4290) );
  OAI21_X2 U15721 ( .A1(n4370), .A2(n4368), .B(n4367), .ZN(n20627) );
  NAND2_X2 U15722 ( .A1(n8332), .A2(n4299), .ZN(n17408) );
  XOR2_X1 U15725 ( .A1(Plaintext[102]), .A2(Key[102]), .Z(n6634) );
  OR2_X1 U15727 ( .A1(n5753), .A2(n5327), .Z(n5752) );
  AND2_X1 U15730 ( .A1(n7161), .A2(n27021), .Z(n7967) );
  AND2_X1 U15734 ( .A1(n21621), .A2(n21620), .Z(n4310) );
  XOR2_X1 U15745 ( .A1(n24549), .A2(n9694), .Z(n5231) );
  INV_X2 U15747 ( .I(n4330), .ZN(n8420) );
  XOR2_X1 U15749 ( .A1(n4332), .A2(n24646), .Z(n6417) );
  NAND2_X1 U15752 ( .A1(n8156), .A2(n7843), .ZN(n25671) );
  OAI21_X2 U15756 ( .A1(n5804), .A2(n26778), .B(n4335), .ZN(n17793) );
  XOR2_X1 U15758 ( .A1(n4338), .A2(n23377), .Z(n10936) );
  XOR2_X1 U15759 ( .A1(n3723), .A2(n25040), .Z(n7999) );
  XOR2_X1 U15760 ( .A1(n32881), .A2(n3723), .Z(n21900) );
  XOR2_X1 U15769 ( .A1(n24764), .A2(n24620), .Z(n4352) );
  XOR2_X1 U15770 ( .A1(n5268), .A2(n13060), .Z(n4353) );
  OAI21_X2 U15771 ( .A1(n12985), .A2(n14913), .B(n12983), .ZN(n13060) );
  XOR2_X1 U15772 ( .A1(n4355), .A2(n24354), .Z(n4354) );
  XOR2_X1 U15773 ( .A1(n5539), .A2(n1231), .Z(n4355) );
  INV_X2 U15777 ( .I(n4362), .ZN(n19630) );
  NAND2_X1 U15778 ( .A1(n18876), .A2(n31948), .ZN(n4365) );
  XOR2_X1 U15788 ( .A1(n28823), .A2(n25224), .Z(n15025) );
  XOR2_X1 U15789 ( .A1(n28823), .A2(n21018), .Z(n5068) );
  XOR2_X1 U15793 ( .A1(n22043), .A2(n22266), .Z(n4379) );
  XOR2_X1 U15794 ( .A1(n12627), .A2(n22045), .Z(n4380) );
  NOR2_X2 U15797 ( .A1(n4387), .A2(n4386), .ZN(n15028) );
  XOR2_X1 U15804 ( .A1(n7363), .A2(n29299), .Z(n7107) );
  XOR2_X1 U15807 ( .A1(n19537), .A2(n4403), .Z(n4401) );
  XOR2_X1 U15809 ( .A1(n19597), .A2(n25001), .Z(n4403) );
  XOR2_X1 U15814 ( .A1(n4413), .A2(n4412), .Z(n4411) );
  XOR2_X1 U15815 ( .A1(n29235), .A2(n26000), .Z(n4412) );
  XOR2_X1 U15816 ( .A1(n23383), .A2(n23465), .Z(n4414) );
  XOR2_X1 U15826 ( .A1(n21993), .A2(n514), .Z(n4427) );
  NAND3_X1 U15832 ( .A1(n23031), .A2(n22945), .A3(n773), .ZN(n7277) );
  INV_X2 U15834 ( .I(n16272), .ZN(n22681) );
  XOR2_X1 U15836 ( .A1(n22182), .A2(n22148), .Z(n4437) );
  XOR2_X1 U15840 ( .A1(n4446), .A2(n4444), .Z(n17150) );
  XOR2_X1 U15841 ( .A1(n4955), .A2(n4445), .Z(n4444) );
  XOR2_X1 U15842 ( .A1(n30321), .A2(n15147), .Z(n4445) );
  MUX2_X1 U15845 ( .I0(n25820), .I1(n25804), .S(n4450), .Z(n4447) );
  XOR2_X1 U15847 ( .A1(n20907), .A2(n28864), .Z(n4448) );
  INV_X2 U15848 ( .I(n4449), .ZN(n4490) );
  INV_X2 U15849 ( .I(n4450), .ZN(n25823) );
  XOR2_X1 U15850 ( .A1(n3682), .A2(n24374), .Z(n22081) );
  XOR2_X1 U15851 ( .A1(n3682), .A2(n25126), .Z(n21899) );
  XOR2_X1 U15854 ( .A1(n12419), .A2(n3682), .Z(n10815) );
  XOR2_X1 U15868 ( .A1(n6156), .A2(n5964), .Z(n4464) );
  XOR2_X1 U15870 ( .A1(n4792), .A2(n4466), .Z(n13932) );
  NOR2_X2 U15875 ( .A1(n6672), .A2(n6377), .ZN(n14564) );
  OAI21_X2 U15877 ( .A1(n24338), .A2(n767), .B(n2847), .ZN(n24165) );
  NAND2_X2 U15878 ( .A1(n16859), .A2(n33990), .ZN(n24166) );
  NAND2_X1 U15883 ( .A1(n15243), .A2(n31129), .ZN(n4486) );
  INV_X2 U15885 ( .I(n31920), .ZN(n25712) );
  OR2_X1 U15890 ( .A1(n10858), .A2(n4770), .Z(n9248) );
  OAI21_X2 U15891 ( .A1(n5532), .A2(n9428), .B(n9426), .ZN(n10858) );
  XOR2_X1 U15898 ( .A1(n4236), .A2(n1424), .Z(n6376) );
  NAND2_X1 U15903 ( .A1(n17767), .A2(n17971), .ZN(n16266) );
  MUX2_X1 U15909 ( .I0(n21536), .I1(n17274), .S(n21569), .Z(n21537) );
  NOR2_X1 U15910 ( .A1(n3376), .A2(n4525), .ZN(n14322) );
  NOR2_X1 U15911 ( .A1(n5113), .A2(n4525), .ZN(n17838) );
  OAI21_X1 U15912 ( .A1(n9481), .A2(n4525), .B(n4524), .ZN(n9480) );
  XOR2_X1 U15920 ( .A1(n28926), .A2(n1395), .Z(n4530) );
  XOR2_X1 U15921 ( .A1(n29918), .A2(n17723), .Z(n17722) );
  OR2_X1 U15925 ( .A1(n17662), .A2(n397), .Z(n12077) );
  XOR2_X1 U15928 ( .A1(n4557), .A2(n4556), .Z(n4555) );
  XOR2_X1 U15929 ( .A1(n26915), .A2(n16555), .Z(n4556) );
  XOR2_X1 U15930 ( .A1(n32899), .A2(n6905), .Z(n4557) );
  XOR2_X1 U15942 ( .A1(n13596), .A2(n4565), .Z(n9164) );
  XOR2_X1 U15943 ( .A1(n7173), .A2(n13595), .Z(n4565) );
  XOR2_X1 U15944 ( .A1(n5970), .A2(n24475), .Z(n7173) );
  XOR2_X1 U15946 ( .A1(n30314), .A2(n30329), .Z(n5600) );
  XOR2_X1 U15955 ( .A1(n26084), .A2(n5169), .Z(n4579) );
  XOR2_X1 U15959 ( .A1(n22153), .A2(n17187), .Z(n4583) );
  NAND2_X1 U15960 ( .A1(n20447), .A2(n31454), .ZN(n4585) );
  XOR2_X1 U15965 ( .A1(n6650), .A2(n22151), .Z(n4590) );
  NAND2_X1 U15966 ( .A1(n1271), .A2(n4599), .ZN(n23015) );
  NAND2_X1 U15967 ( .A1(n14540), .A2(n4599), .ZN(n17399) );
  INV_X2 U15969 ( .I(n29061), .ZN(n18891) );
  NOR2_X1 U15970 ( .A1(n29061), .A2(n14926), .ZN(n11410) );
  INV_X1 U15971 ( .I(Plaintext[16]), .ZN(n4601) );
  XOR2_X1 U15978 ( .A1(n15183), .A2(n27126), .Z(n4610) );
  OR2_X1 U15980 ( .A1(n18266), .A2(n18265), .Z(n4618) );
  XOR2_X1 U15983 ( .A1(n14382), .A2(n14381), .Z(n8523) );
  NOR2_X1 U15984 ( .A1(n32127), .A2(n18643), .ZN(n4624) );
  AOI21_X1 U15986 ( .A1(n17266), .A2(n4626), .B(n28238), .ZN(n18378) );
  AOI21_X1 U16000 ( .A1(n11893), .A2(n565), .B(n16317), .ZN(n4636) );
  AOI21_X1 U16002 ( .A1(n7039), .A2(n4642), .B(n7037), .ZN(n10157) );
  XOR2_X1 U16003 ( .A1(n2045), .A2(n25167), .Z(n10163) );
  OAI21_X1 U16011 ( .A1(n19301), .A2(n1052), .B(n4658), .ZN(n14736) );
  XOR2_X1 U16012 ( .A1(n23182), .A2(n538), .Z(n4660) );
  XOR2_X1 U16014 ( .A1(n23138), .A2(n529), .Z(n4662) );
  XOR2_X1 U16015 ( .A1(n23267), .A2(n31727), .Z(n23138) );
  INV_X1 U16016 ( .I(n31161), .ZN(n4663) );
  XNOR2_X1 U16025 ( .A1(Plaintext[182]), .A2(Key[182]), .ZN(n4669) );
  XOR2_X1 U16028 ( .A1(n32648), .A2(n16506), .Z(n4671) );
  NAND2_X1 U16035 ( .A1(n7802), .A2(n4834), .ZN(n4678) );
  XOR2_X1 U16039 ( .A1(n29918), .A2(n16525), .Z(n4681) );
  AOI21_X1 U16041 ( .A1(n25265), .A2(n25264), .B(n4685), .ZN(n25267) );
  OAI22_X1 U16042 ( .A1(n1207), .A2(n4686), .B1(n12431), .B2(n25284), .ZN(
        n4685) );
  OR2_X1 U16044 ( .A1(n25285), .A2(n25277), .Z(n4686) );
  AOI21_X1 U16048 ( .A1(n20635), .A2(n4693), .B(n26278), .ZN(n20322) );
  NOR2_X1 U16054 ( .A1(n21721), .A2(n3467), .ZN(n4699) );
  XOR2_X1 U16059 ( .A1(n4704), .A2(n16705), .Z(n8718) );
  XOR2_X1 U16060 ( .A1(n4704), .A2(n19570), .Z(n11354) );
  NAND2_X2 U16065 ( .A1(n18694), .A2(n18693), .ZN(n10714) );
  NAND2_X1 U16066 ( .A1(n7687), .A2(n11477), .ZN(n4716) );
  NAND2_X2 U16067 ( .A1(n15576), .A2(n15574), .ZN(n11477) );
  XOR2_X1 U16073 ( .A1(n8306), .A2(n16555), .Z(n4720) );
  XOR2_X1 U16080 ( .A1(n4727), .A2(n4724), .Z(n10337) );
  XOR2_X1 U16081 ( .A1(n4726), .A2(n4725), .Z(n4724) );
  XOR2_X1 U16082 ( .A1(n1923), .A2(n25669), .Z(n4725) );
  XOR2_X1 U16083 ( .A1(n20783), .A2(n20955), .Z(n4726) );
  XOR2_X1 U16088 ( .A1(n4783), .A2(n15707), .Z(n17498) );
  XOR2_X1 U16089 ( .A1(n4729), .A2(n13825), .Z(n4783) );
  NAND3_X2 U16091 ( .A1(n5130), .A2(n5129), .A3(n668), .ZN(n14855) );
  NAND2_X2 U16092 ( .A1(n10313), .A2(n9462), .ZN(n5016) );
  XOR2_X1 U16104 ( .A1(n22017), .A2(n22033), .Z(n4739) );
  XOR2_X1 U16106 ( .A1(n12376), .A2(n22108), .Z(n22016) );
  NOR2_X1 U16112 ( .A1(n8270), .A2(n9172), .ZN(n4743) );
  XOR2_X1 U16124 ( .A1(n20897), .A2(n11066), .Z(n4759) );
  NOR2_X1 U16125 ( .A1(n21604), .A2(n17098), .ZN(n11081) );
  XOR2_X1 U16126 ( .A1(n4763), .A2(n4762), .Z(n4761) );
  XOR2_X1 U16127 ( .A1(n10292), .A2(n25086), .Z(n4762) );
  NOR2_X2 U16128 ( .A1(n6266), .A2(n4765), .ZN(n10953) );
  NAND3_X2 U16129 ( .A1(n4772), .A2(n14546), .A3(n13933), .ZN(n6857) );
  XOR2_X1 U16132 ( .A1(Plaintext[15]), .A2(Key[15]), .Z(n4808) );
  XOR2_X1 U16133 ( .A1(n4783), .A2(n13824), .Z(n10617) );
  XOR2_X1 U16134 ( .A1(n15606), .A2(n25190), .Z(n5031) );
  XOR2_X1 U16135 ( .A1(n31597), .A2(n3977), .Z(n22320) );
  XOR2_X1 U16136 ( .A1(n3977), .A2(n4788), .Z(n22002) );
  XOR2_X1 U16137 ( .A1(n11750), .A2(n4789), .Z(n11748) );
  XOR2_X1 U16142 ( .A1(n23358), .A2(n25801), .Z(n4794) );
  XOR2_X1 U16149 ( .A1(n13970), .A2(n32310), .Z(n10799) );
  XOR2_X1 U16154 ( .A1(n27130), .A2(n30495), .Z(n22111) );
  INV_X2 U16159 ( .I(n4808), .ZN(n11390) );
  NAND2_X2 U16160 ( .A1(n4811), .A2(n4809), .ZN(n23056) );
  NAND2_X2 U16163 ( .A1(n7253), .A2(n7252), .ZN(n20899) );
  AOI21_X2 U16165 ( .A1(n23952), .A2(n16281), .B(n17664), .ZN(n4821) );
  XOR2_X1 U16174 ( .A1(n22264), .A2(n27120), .Z(n15367) );
  XOR2_X1 U16176 ( .A1(n22214), .A2(n16530), .Z(n4831) );
  NAND2_X2 U16181 ( .A1(n10693), .A2(n10694), .ZN(n4835) );
  NOR2_X1 U16183 ( .A1(n4835), .A2(n11444), .ZN(n11263) );
  NOR2_X1 U16186 ( .A1(n11085), .A2(n4835), .ZN(n11688) );
  XOR2_X1 U16191 ( .A1(n15674), .A2(n24267), .Z(n4840) );
  NAND2_X2 U16194 ( .A1(n24259), .A2(n17800), .ZN(n6547) );
  XOR2_X1 U16195 ( .A1(n4849), .A2(n598), .Z(n11733) );
  NOR2_X1 U16197 ( .A1(n29495), .A2(n4396), .ZN(n11195) );
  NOR2_X1 U16198 ( .A1(n22558), .A2(n22671), .ZN(n4850) );
  XOR2_X1 U16207 ( .A1(n21926), .A2(n8979), .Z(n4861) );
  NAND2_X1 U16208 ( .A1(n8079), .A2(n27543), .ZN(n21790) );
  AOI21_X2 U16209 ( .A1(n4865), .A2(n27842), .B(n4863), .ZN(n21789) );
  NAND2_X1 U16211 ( .A1(n171), .A2(n4869), .ZN(n18384) );
  NOR2_X1 U16212 ( .A1(n18571), .A2(n4869), .ZN(n18385) );
  OAI21_X1 U16213 ( .A1(n1190), .A2(n4869), .B(n29087), .ZN(n5053) );
  XOR2_X1 U16214 ( .A1(Plaintext[99]), .A2(Key[99]), .Z(n18823) );
  XOR2_X1 U16218 ( .A1(n19584), .A2(n8089), .Z(n4884) );
  XOR2_X1 U16219 ( .A1(n27733), .A2(n25911), .Z(n14407) );
  XOR2_X1 U16221 ( .A1(n27733), .A2(n24968), .Z(n24404) );
  XOR2_X1 U16222 ( .A1(n1604), .A2(n1394), .Z(n17041) );
  XOR2_X1 U16223 ( .A1(n10006), .A2(n27185), .Z(n10005) );
  INV_X2 U16224 ( .I(n11888), .ZN(n4891) );
  NAND2_X1 U16225 ( .A1(n23919), .A2(n4892), .ZN(n15095) );
  NAND2_X1 U16226 ( .A1(n16620), .A2(n33221), .ZN(n23349) );
  NAND3_X1 U16234 ( .A1(n24903), .A2(n27248), .A3(n10099), .ZN(n4899) );
  NAND2_X2 U16235 ( .A1(n4903), .A2(n4900), .ZN(n24915) );
  INV_X1 U16236 ( .I(n5763), .ZN(n4903) );
  XOR2_X1 U16242 ( .A1(n34047), .A2(n25319), .Z(n4915) );
  XOR2_X1 U16243 ( .A1(n18180), .A2(n20816), .Z(n20956) );
  NAND2_X2 U16247 ( .A1(n4919), .A2(n6501), .ZN(n16023) );
  OR2_X1 U16248 ( .A1(n1335), .A2(n11915), .Z(n4922) );
  NAND2_X2 U16263 ( .A1(n5534), .A2(n5533), .ZN(n5128) );
  OR2_X1 U16266 ( .A1(n13601), .A2(n30191), .Z(n4960) );
  XOR2_X1 U16269 ( .A1(n31229), .A2(n29121), .Z(n17042) );
  NAND2_X1 U16272 ( .A1(n3657), .A2(n32531), .ZN(n4982) );
  NOR2_X1 U16276 ( .A1(n19855), .A2(n3989), .ZN(n5909) );
  MUX2_X1 U16280 ( .I0(n5073), .I1(n20155), .S(n9724), .Z(n12322) );
  XOR2_X1 U16284 ( .A1(n4992), .A2(n26076), .Z(n11351) );
  XOR2_X1 U16296 ( .A1(n5013), .A2(n5011), .Z(n9757) );
  XOR2_X1 U16297 ( .A1(n5012), .A2(n9758), .Z(n5011) );
  XOR2_X1 U16301 ( .A1(n24830), .A2(n11297), .Z(n5021) );
  XNOR2_X1 U16304 ( .A1(n5022), .A2(n5023), .ZN(n5019) );
  NAND2_X2 U16306 ( .A1(n5027), .A2(n5025), .ZN(n20968) );
  XOR2_X1 U16307 ( .A1(n20968), .A2(n16612), .Z(n5431) );
  NOR2_X1 U16308 ( .A1(n16789), .A2(n20096), .ZN(n18041) );
  XOR2_X1 U16309 ( .A1(n7375), .A2(n7374), .Z(n10414) );
  XOR2_X1 U16311 ( .A1(n22012), .A2(n13067), .Z(n22168) );
  NAND2_X1 U16314 ( .A1(n15601), .A2(n5035), .ZN(n22959) );
  XOR2_X1 U16316 ( .A1(n23261), .A2(n556), .Z(n5038) );
  INV_X1 U16322 ( .I(n24132), .ZN(n5066) );
  XOR2_X1 U16324 ( .A1(n5070), .A2(n5069), .Z(n11515) );
  XOR2_X1 U16325 ( .A1(n20721), .A2(n5071), .Z(n5069) );
  XOR2_X1 U16326 ( .A1(n5772), .A2(n1067), .Z(n5071) );
  INV_X2 U16327 ( .I(n7940), .ZN(n7941) );
  INV_X2 U16331 ( .I(n5074), .ZN(n9724) );
  XOR2_X1 U16336 ( .A1(n2073), .A2(n16613), .Z(n5081) );
  OAI22_X2 U16337 ( .A1(n7438), .A2(n12532), .B1(n7437), .B2(n7436), .ZN(
        n19426) );
  INV_X1 U16343 ( .I(n5089), .ZN(n24656) );
  XOR2_X1 U16344 ( .A1(n5090), .A2(n16402), .Z(n9694) );
  XOR2_X1 U16345 ( .A1(n5090), .A2(n16605), .Z(n24379) );
  NAND2_X1 U16347 ( .A1(n979), .A2(n5097), .ZN(n6694) );
  XOR2_X1 U16350 ( .A1(n28709), .A2(n22248), .Z(n5099) );
  XOR2_X1 U16353 ( .A1(n5106), .A2(n5104), .Z(n22579) );
  XOR2_X1 U16354 ( .A1(n5105), .A2(n13371), .Z(n5104) );
  XOR2_X1 U16357 ( .A1(n22296), .A2(n22147), .Z(n5107) );
  XOR2_X1 U16359 ( .A1(n22149), .A2(n16613), .Z(n5109) );
  XOR2_X1 U16368 ( .A1(n22004), .A2(n21658), .Z(n5126) );
  XOR2_X1 U16372 ( .A1(n5133), .A2(n20661), .Z(n9980) );
  NOR2_X2 U16374 ( .A1(n12181), .A2(n15317), .ZN(n5380) );
  INV_X1 U16381 ( .I(n5140), .ZN(n9800) );
  XOR2_X1 U16385 ( .A1(n5146), .A2(n5147), .Z(n5145) );
  XOR2_X1 U16386 ( .A1(n16733), .A2(n29954), .Z(n5147) );
  NAND2_X2 U16388 ( .A1(n9314), .A2(n9317), .ZN(n17430) );
  XOR2_X1 U16389 ( .A1(n19551), .A2(n19465), .Z(n5152) );
  XOR2_X1 U16395 ( .A1(n23502), .A2(n7994), .Z(n5159) );
  XOR2_X1 U16409 ( .A1(n32255), .A2(n13438), .Z(n13437) );
  XOR2_X1 U16410 ( .A1(n32255), .A2(n25208), .Z(n13453) );
  XOR2_X1 U16411 ( .A1(n16429), .A2(n24907), .Z(n5169) );
  XOR2_X1 U16421 ( .A1(n30303), .A2(n20784), .Z(n21011) );
  INV_X2 U16422 ( .I(n5188), .ZN(n8443) );
  XOR2_X1 U16433 ( .A1(n5197), .A2(n10004), .Z(n16392) );
  XOR2_X1 U16434 ( .A1(n7288), .A2(n21457), .Z(n5197) );
  XOR2_X1 U16440 ( .A1(n13198), .A2(n26103), .Z(n5207) );
  XOR2_X1 U16442 ( .A1(n5462), .A2(n25450), .Z(n18902) );
  XOR2_X1 U16443 ( .A1(n24785), .A2(n25832), .Z(n24537) );
  XOR2_X1 U16444 ( .A1(n24785), .A2(n16520), .Z(n6053) );
  XOR2_X1 U16446 ( .A1(n20899), .A2(n24937), .Z(n5210) );
  XOR2_X1 U16451 ( .A1(n23502), .A2(n23406), .Z(n5215) );
  NAND2_X2 U16454 ( .A1(n5218), .A2(n5216), .ZN(n20885) );
  NOR2_X1 U16457 ( .A1(n21801), .A2(n5228), .ZN(n15639) );
  NAND2_X2 U16460 ( .A1(n10811), .A2(n24119), .ZN(n24573) );
  XNOR2_X1 U16461 ( .A1(n10631), .A2(n5790), .ZN(n10729) );
  XOR2_X1 U16465 ( .A1(n5237), .A2(n1045), .Z(n5236) );
  XOR2_X1 U16466 ( .A1(n19772), .A2(n1065), .Z(n5237) );
  NAND2_X1 U16467 ( .A1(n17640), .A2(n5239), .ZN(n9558) );
  XOR2_X1 U16472 ( .A1(n5724), .A2(n9908), .Z(n5240) );
  XOR2_X1 U16475 ( .A1(n20873), .A2(n20872), .Z(n20902) );
  XOR2_X1 U16477 ( .A1(n5243), .A2(n25225), .Z(Ciphertext[77]) );
  XOR2_X1 U16480 ( .A1(n5256), .A2(n5255), .Z(n6552) );
  XOR2_X1 U16481 ( .A1(n24415), .A2(n554), .Z(n5255) );
  XOR2_X1 U16487 ( .A1(Plaintext[140]), .A2(Key[140]), .Z(n10664) );
  INV_X1 U16488 ( .I(n5273), .ZN(n5272) );
  XOR2_X1 U16492 ( .A1(n23209), .A2(n16464), .Z(n5277) );
  XOR2_X1 U16495 ( .A1(n6156), .A2(n19707), .Z(n5279) );
  XOR2_X1 U16496 ( .A1(n14337), .A2(n11219), .Z(n19707) );
  XOR2_X1 U16497 ( .A1(n19709), .A2(n18082), .Z(n5280) );
  MUX2_X1 U16504 ( .I0(n16493), .I1(n20012), .S(n13605), .Z(n19880) );
  XOR2_X1 U16507 ( .A1(n29885), .A2(n26915), .Z(n15690) );
  XOR2_X1 U16515 ( .A1(n12414), .A2(n1070), .Z(n5297) );
  AOI22_X2 U16516 ( .A1(n21748), .A2(n21750), .B1(n13815), .B2(n30346), .ZN(
        n11458) );
  NOR2_X1 U16518 ( .A1(n23081), .A2(n1577), .ZN(n8126) );
  MUX2_X1 U16519 ( .I0(n6985), .I1(n23082), .S(n1577), .Z(n23080) );
  NOR2_X1 U16520 ( .A1(n12869), .A2(n1124), .ZN(n5305) );
  XOR2_X1 U16526 ( .A1(n5316), .A2(n29344), .Z(n5315) );
  XOR2_X1 U16531 ( .A1(n15527), .A2(n12998), .Z(n5322) );
  NAND3_X1 U16534 ( .A1(n25410), .A2(n752), .A3(n25405), .ZN(n24702) );
  XOR2_X1 U16536 ( .A1(n17548), .A2(Key[101]), .Z(n17558) );
  XOR2_X1 U16541 ( .A1(n20710), .A2(n5337), .Z(n5336) );
  XOR2_X1 U16545 ( .A1(n5340), .A2(n5338), .Z(n6143) );
  XOR2_X1 U16546 ( .A1(n24568), .A2(n5339), .Z(n5338) );
  XOR2_X1 U16547 ( .A1(n12454), .A2(n24943), .Z(n5339) );
  XOR2_X1 U16550 ( .A1(n15114), .A2(n17871), .Z(n12659) );
  XOR2_X1 U16555 ( .A1(n4295), .A2(n25358), .Z(n5352) );
  INV_X2 U16570 ( .I(n5361), .ZN(n6855) );
  NAND2_X1 U16571 ( .A1(n22462), .A2(n22343), .ZN(n23011) );
  MUX2_X1 U16580 ( .I0(n23902), .I1(n23629), .S(n1254), .Z(n23631) );
  INV_X2 U16583 ( .I(n11988), .ZN(n7116) );
  INV_X2 U16588 ( .I(n5392), .ZN(n11915) );
  XOR2_X1 U16589 ( .A1(Plaintext[133]), .A2(Key[133]), .Z(n14156) );
  INV_X2 U16590 ( .I(n5401), .ZN(n17967) );
  XOR2_X1 U16599 ( .A1(n11762), .A2(n5422), .Z(n5421) );
  XOR2_X1 U16600 ( .A1(n14125), .A2(n25598), .Z(n5422) );
  XOR2_X1 U16603 ( .A1(n29318), .A2(n24750), .Z(n5425) );
  NAND2_X1 U16609 ( .A1(n886), .A2(n752), .ZN(n24701) );
  INV_X2 U16614 ( .I(n5432), .ZN(n24975) );
  XOR2_X1 U16616 ( .A1(n19742), .A2(n5435), .Z(n5434) );
  XOR2_X1 U16617 ( .A1(n19466), .A2(n27995), .Z(n5435) );
  XOR2_X1 U16622 ( .A1(Key[136]), .A2(Plaintext[136]), .Z(n16995) );
  XOR2_X1 U16625 ( .A1(n23402), .A2(n23226), .Z(n5445) );
  XOR2_X1 U16636 ( .A1(n15844), .A2(n19641), .Z(n19467) );
  NAND2_X2 U16641 ( .A1(n5460), .A2(n9352), .ZN(n20554) );
  NAND2_X1 U16642 ( .A1(n20169), .A2(n5460), .ZN(n20172) );
  INV_X2 U16643 ( .I(n20521), .ZN(n5460) );
  XOR2_X1 U16644 ( .A1(n5472), .A2(n3929), .Z(n9605) );
  XOR2_X1 U16645 ( .A1(n5472), .A2(n16530), .Z(n10424) );
  XOR2_X1 U16646 ( .A1(Plaintext[98]), .A2(Key[98]), .Z(n16450) );
  INV_X2 U16649 ( .I(n7348), .ZN(n5476) );
  OAI21_X2 U16651 ( .A1(n18824), .A2(n17735), .B(n5478), .ZN(n19128) );
  NOR2_X1 U16653 ( .A1(n16093), .A2(n26600), .ZN(n13957) );
  NOR2_X1 U16654 ( .A1(n4656), .A2(n26600), .ZN(n19084) );
  INV_X2 U16656 ( .I(n6854), .ZN(n5480) );
  XOR2_X1 U16657 ( .A1(n5483), .A2(n19481), .Z(n19482) );
  XOR2_X1 U16658 ( .A1(n7971), .A2(n5484), .Z(n5483) );
  XOR2_X1 U16668 ( .A1(n5513), .A2(n21650), .Z(n5501) );
  XOR2_X1 U16670 ( .A1(n859), .A2(n22099), .Z(n5503) );
  INV_X2 U16671 ( .I(n5504), .ZN(n15746) );
  AOI21_X2 U16672 ( .A1(n23404), .A2(n5742), .B(n5505), .ZN(n11326) );
  XOR2_X1 U16675 ( .A1(n26582), .A2(n27179), .Z(n5508) );
  XOR2_X1 U16680 ( .A1(n14289), .A2(n4057), .Z(n5513) );
  XOR2_X1 U16681 ( .A1(n27148), .A2(n5399), .Z(n23386) );
  XOR2_X1 U16682 ( .A1(n5518), .A2(n5515), .Z(n21168) );
  XOR2_X1 U16683 ( .A1(n5517), .A2(n5516), .Z(n5515) );
  XOR2_X1 U16684 ( .A1(n20860), .A2(n16502), .Z(n5516) );
  XOR2_X1 U16685 ( .A1(n17554), .A2(n21016), .Z(n5517) );
  XOR2_X1 U16693 ( .A1(n31508), .A2(n24748), .Z(n5522) );
  XOR2_X1 U16696 ( .A1(n6156), .A2(n19343), .Z(n5526) );
  INV_X2 U16697 ( .I(n5527), .ZN(n23765) );
  NOR2_X1 U16701 ( .A1(n33714), .A2(n820), .ZN(n5582) );
  AOI21_X1 U16709 ( .A1(n17725), .A2(n19063), .B(n1053), .ZN(n7186) );
  NOR3_X1 U16711 ( .A1(n21560), .A2(n14236), .A3(n5546), .ZN(n15319) );
  NOR2_X1 U16713 ( .A1(n3657), .A2(n850), .ZN(n6696) );
  INV_X1 U16714 ( .I(n21636), .ZN(n21638) );
  NOR2_X2 U16715 ( .A1(n9186), .A2(n780), .ZN(n5575) );
  XOR2_X1 U16720 ( .A1(n19564), .A2(n456), .Z(n5562) );
  NAND2_X1 U16723 ( .A1(n5575), .A2(n21453), .ZN(n20436) );
  AOI21_X1 U16724 ( .A1(n25217), .A2(n5043), .B(n5577), .ZN(n25219) );
  INV_X2 U16732 ( .I(n22535), .ZN(n22537) );
  OAI21_X2 U16739 ( .A1(n31923), .A2(n12610), .B(n5602), .ZN(n19556) );
  NOR2_X2 U16742 ( .A1(n17556), .A2(n12744), .ZN(n19424) );
  XOR2_X1 U16744 ( .A1(n9955), .A2(n16824), .Z(n5609) );
  OAI21_X2 U16751 ( .A1(n5656), .A2(n5655), .B(n4643), .ZN(n15073) );
  XOR2_X1 U16756 ( .A1(n16708), .A2(n25355), .Z(n5629) );
  NAND2_X2 U16760 ( .A1(n18986), .A2(n5637), .ZN(n19589) );
  XNOR2_X1 U16770 ( .A1(n22144), .A2(n21920), .ZN(n5658) );
  XOR2_X1 U16771 ( .A1(n21726), .A2(n22100), .Z(n21920) );
  XOR2_X1 U16775 ( .A1(n9848), .A2(n5666), .Z(n5663) );
  XOR2_X1 U16779 ( .A1(n24532), .A2(n16301), .Z(n5666) );
  INV_X2 U16788 ( .I(n5675), .ZN(n16625) );
  NOR2_X1 U16790 ( .A1(n5677), .A2(n18493), .ZN(n18424) );
  NOR2_X1 U16791 ( .A1(n18326), .A2(n5677), .ZN(n5676) );
  NAND2_X2 U16792 ( .A1(n5682), .A2(n8786), .ZN(n23485) );
  NAND4_X2 U16795 ( .A1(n11725), .A2(n11724), .A3(n15781), .A4(n5690), .ZN(
        n11722) );
  XOR2_X1 U16797 ( .A1(n5692), .A2(n5691), .Z(n17812) );
  XOR2_X1 U16798 ( .A1(n23249), .A2(n23251), .Z(n5691) );
  OAI22_X1 U16804 ( .A1(n32868), .A2(n803), .B1(n724), .B2(n3163), .ZN(n22693)
         );
  XOR2_X1 U16805 ( .A1(n5699), .A2(n5697), .Z(n15009) );
  XOR2_X1 U16806 ( .A1(n5698), .A2(n14415), .Z(n5697) );
  XOR2_X1 U16807 ( .A1(n4400), .A2(n25098), .Z(n5698) );
  XOR2_X1 U16813 ( .A1(n34056), .A2(n23224), .Z(n5702) );
  NOR2_X1 U16818 ( .A1(n5707), .A2(n31017), .ZN(n13649) );
  NAND2_X1 U16822 ( .A1(n7334), .A2(n5713), .ZN(n25083) );
  NAND2_X1 U16823 ( .A1(n5713), .A2(n25106), .ZN(n5712) );
  XOR2_X1 U16827 ( .A1(n546), .A2(n24817), .Z(n5714) );
  XOR2_X1 U16832 ( .A1(n511), .A2(n13901), .Z(n5722) );
  INV_X2 U16834 ( .I(n6894), .ZN(n16668) );
  XOR2_X1 U16837 ( .A1(n26084), .A2(n18011), .Z(n5726) );
  XOR2_X1 U16842 ( .A1(n20977), .A2(n5733), .Z(n5732) );
  XOR2_X1 U16843 ( .A1(n16708), .A2(n16381), .Z(n5733) );
  NOR2_X1 U16851 ( .A1(n978), .A2(n28222), .ZN(n5745) );
  NAND2_X2 U16853 ( .A1(n7538), .A2(n5754), .ZN(n14147) );
  XOR2_X1 U16855 ( .A1(n22021), .A2(n21886), .Z(n21903) );
  XOR2_X1 U16857 ( .A1(n30069), .A2(n31308), .Z(n10923) );
  NAND2_X1 U16859 ( .A1(n1384), .A2(n5760), .ZN(n7434) );
  XOR2_X1 U16862 ( .A1(n24643), .A2(n30104), .Z(n24376) );
  XOR2_X1 U16866 ( .A1(n7135), .A2(n7606), .Z(n5767) );
  NAND2_X1 U16868 ( .A1(n16205), .A2(n1122), .ZN(n5771) );
  NAND3_X1 U16869 ( .A1(n30328), .A2(n24922), .A3(n15569), .ZN(n5774) );
  MUX2_X1 U16870 ( .I0(n32571), .I1(n1211), .S(n33585), .Z(n25786) );
  XOR2_X1 U16872 ( .A1(n5775), .A2(n6324), .Z(n15994) );
  INV_X1 U16879 ( .I(n5792), .ZN(n5791) );
  XOR2_X1 U16883 ( .A1(n8232), .A2(n17793), .Z(n13899) );
  NAND2_X1 U16884 ( .A1(n5805), .A2(n28987), .ZN(n5890) );
  NOR2_X2 U16893 ( .A1(n7464), .A2(n21929), .ZN(n7463) );
  XOR2_X1 U16896 ( .A1(n24785), .A2(n1421), .Z(n13793) );
  XOR2_X1 U16899 ( .A1(n22085), .A2(n22096), .Z(n21921) );
  XOR2_X1 U16903 ( .A1(n5838), .A2(n1194), .Z(Ciphertext[151]) );
  NAND3_X1 U16905 ( .A1(n30346), .A2(n13816), .A3(n21840), .ZN(n14739) );
  NAND2_X1 U16906 ( .A1(n16987), .A2(n5843), .ZN(n21685) );
  NAND2_X1 U16907 ( .A1(n16386), .A2(n30346), .ZN(n21841) );
  XOR2_X1 U16909 ( .A1(n5844), .A2(n11766), .Z(n11765) );
  XOR2_X1 U16912 ( .A1(n23474), .A2(n16597), .Z(n5846) );
  AOI21_X1 U16915 ( .A1(n18492), .A2(n17813), .B(n17316), .ZN(n5852) );
  NAND2_X1 U16922 ( .A1(n6493), .A2(n780), .ZN(n9273) );
  NAND2_X1 U16923 ( .A1(n17437), .A2(n1337), .ZN(n5857) );
  XOR2_X1 U16924 ( .A1(n5862), .A2(n5859), .Z(n5870) );
  XOR2_X1 U16925 ( .A1(n5861), .A2(n5860), .Z(n5859) );
  XOR2_X1 U16926 ( .A1(n14588), .A2(n16655), .Z(n5860) );
  INV_X1 U16933 ( .I(n22336), .ZN(n22413) );
  INV_X2 U16944 ( .I(n5870), .ZN(n16154) );
  XOR2_X1 U16946 ( .A1(n9160), .A2(n16734), .Z(n15077) );
  XOR2_X1 U16947 ( .A1(n23324), .A2(n12200), .Z(n5881) );
  INV_X1 U16948 ( .I(n23213), .ZN(n5882) );
  XOR2_X1 U16950 ( .A1(n21911), .A2(n6183), .Z(n5885) );
  NAND2_X1 U16952 ( .A1(n18274), .A2(n27129), .ZN(n5891) );
  XOR2_X1 U16960 ( .A1(n5904), .A2(n26701), .Z(n14036) );
  NOR2_X1 U16963 ( .A1(n6899), .A2(n17947), .ZN(n5911) );
  XOR2_X1 U16966 ( .A1(n5916), .A2(n1069), .Z(Ciphertext[127]) );
  XOR2_X1 U16968 ( .A1(n19649), .A2(n16506), .Z(n5919) );
  XOR2_X1 U16970 ( .A1(n19721), .A2(n5921), .Z(n5920) );
  NAND3_X2 U16981 ( .A1(n19904), .A2(n19905), .A3(n5931), .ZN(n20561) );
  XOR2_X1 U16983 ( .A1(n5940), .A2(n23535), .Z(n5939) );
  XOR2_X1 U16984 ( .A1(n23534), .A2(n16634), .Z(n5940) );
  XOR2_X1 U16985 ( .A1(n7933), .A2(n5941), .Z(n8167) );
  XOR2_X1 U16986 ( .A1(n22293), .A2(n610), .Z(n5941) );
  NAND2_X1 U16989 ( .A1(n19033), .A2(n5946), .ZN(n5945) );
  NAND2_X1 U16990 ( .A1(n21404), .A2(n596), .ZN(n5948) );
  INV_X2 U16992 ( .I(n5962), .ZN(n10871) );
  NAND2_X1 U16994 ( .A1(n2858), .A2(n5991), .ZN(n5963) );
  INV_X2 U16995 ( .I(n19230), .ZN(n19783) );
  XOR2_X1 U16996 ( .A1(n19230), .A2(n1406), .Z(n5964) );
  INV_X2 U16997 ( .I(n5965), .ZN(n17240) );
  NAND2_X1 U16998 ( .A1(n885), .A2(n25012), .ZN(n24477) );
  XOR2_X1 U17003 ( .A1(n22130), .A2(n22192), .Z(n22293) );
  NAND2_X2 U17008 ( .A1(n13707), .A2(n13708), .ZN(n19384) );
  INV_X2 U17010 ( .I(n9203), .ZN(n11912) );
  OAI21_X1 U17013 ( .A1(n15456), .A2(n5981), .B(n15457), .ZN(n5983) );
  XOR2_X1 U17016 ( .A1(n11332), .A2(n24442), .Z(n24795) );
  NAND2_X1 U17018 ( .A1(n22606), .A2(n5991), .ZN(n6186) );
  NAND2_X1 U17019 ( .A1(n4066), .A2(n19156), .ZN(n15120) );
  NOR2_X1 U17020 ( .A1(n18426), .A2(n4066), .ZN(n18979) );
  XOR2_X1 U17021 ( .A1(n3799), .A2(n25801), .Z(n20647) );
  XOR2_X1 U17022 ( .A1(n5994), .A2(n22005), .Z(n21916) );
  XOR2_X1 U17024 ( .A1(n28082), .A2(n31308), .Z(n8755) );
  NAND2_X1 U17027 ( .A1(n6003), .A2(n30146), .ZN(n12692) );
  XOR2_X1 U17031 ( .A1(n6008), .A2(n6005), .Z(n24459) );
  XOR2_X1 U17032 ( .A1(n6007), .A2(n6006), .Z(n6005) );
  XOR2_X1 U17033 ( .A1(n24526), .A2(n25722), .Z(n6006) );
  XOR2_X1 U17034 ( .A1(n24799), .A2(n24809), .Z(n6007) );
  NAND2_X2 U17039 ( .A1(n6322), .A2(n7648), .ZN(n23109) );
  XOR2_X1 U17044 ( .A1(n22130), .A2(n25545), .Z(n6018) );
  XOR2_X1 U17046 ( .A1(n13020), .A2(n22049), .Z(n6020) );
  INV_X1 U17048 ( .I(n6673), .ZN(n10011) );
  XOR2_X1 U17054 ( .A1(n24478), .A2(n25206), .Z(n12032) );
  XOR2_X1 U17057 ( .A1(n19763), .A2(n19649), .Z(n6028) );
  OAI21_X2 U17058 ( .A1(n6030), .A2(n6029), .B(n9134), .ZN(n19763) );
  XOR2_X1 U17059 ( .A1(n6033), .A2(n6032), .Z(n6031) );
  XOR2_X1 U17060 ( .A1(n19764), .A2(n25783), .Z(n6032) );
  XOR2_X1 U17066 ( .A1(n31229), .A2(n24833), .Z(n14217) );
  XOR2_X1 U17067 ( .A1(n7046), .A2(n25728), .Z(n7994) );
  XOR2_X1 U17068 ( .A1(n7046), .A2(n15409), .Z(n15408) );
  XOR2_X1 U17075 ( .A1(n13471), .A2(n6053), .Z(n6052) );
  XOR2_X1 U17080 ( .A1(n22213), .A2(n6056), .Z(n6055) );
  XOR2_X1 U17081 ( .A1(n15825), .A2(n16527), .Z(n6056) );
  XOR2_X1 U17089 ( .A1(n26683), .A2(n27101), .Z(n16824) );
  XOR2_X1 U17090 ( .A1(n26683), .A2(n16671), .Z(n7875) );
  XOR2_X1 U17091 ( .A1(n26683), .A2(n25506), .Z(n14315) );
  XOR2_X1 U17092 ( .A1(n26530), .A2(n20747), .Z(n6078) );
  XOR2_X1 U17101 ( .A1(n6088), .A2(n6087), .Z(n6086) );
  XOR2_X1 U17102 ( .A1(n20825), .A2(n25880), .Z(n6087) );
  XOR2_X1 U17103 ( .A1(n23181), .A2(n10218), .Z(n10219) );
  XOR2_X1 U17112 ( .A1(n6095), .A2(n25466), .Z(Ciphertext[111]) );
  MUX2_X1 U17114 ( .I0(n25462), .I1(n25473), .S(n6310), .Z(n6097) );
  AOI21_X2 U17115 ( .A1(n13249), .A2(n16490), .B(n9738), .ZN(n23051) );
  XOR2_X1 U17116 ( .A1(n6103), .A2(n24643), .Z(n9943) );
  NAND3_X1 U17119 ( .A1(n9625), .A2(n33597), .A3(n5308), .ZN(n6104) );
  XOR2_X1 U17122 ( .A1(n19385), .A2(n6115), .Z(n19387) );
  XOR2_X1 U17127 ( .A1(n2896), .A2(n13579), .Z(n6318) );
  XOR2_X1 U17132 ( .A1(n27922), .A2(n1192), .Z(n6127) );
  NAND2_X1 U17134 ( .A1(n14652), .A2(n6138), .ZN(n13686) );
  XOR2_X1 U17137 ( .A1(n16897), .A2(n22242), .Z(n9790) );
  NOR2_X1 U17141 ( .A1(n22963), .A2(n6149), .ZN(n6150) );
  XOR2_X1 U17144 ( .A1(n23449), .A2(n23288), .Z(n6151) );
  NAND2_X1 U17147 ( .A1(n8304), .A2(n24908), .ZN(n6155) );
  XOR2_X1 U17148 ( .A1(n6159), .A2(n6160), .Z(n13304) );
  NAND2_X2 U17152 ( .A1(n7255), .A2(n7254), .ZN(n20954) );
  INV_X2 U17153 ( .I(n9627), .ZN(n9706) );
  XOR2_X1 U17154 ( .A1(n20833), .A2(n6161), .Z(n6160) );
  XOR2_X1 U17155 ( .A1(n9627), .A2(n6162), .Z(n6161) );
  INV_X1 U17156 ( .I(n25324), .ZN(n6162) );
  XNOR2_X1 U17157 ( .A1(n17517), .A2(n6906), .ZN(n20833) );
  XOR2_X1 U17162 ( .A1(n11206), .A2(n16597), .Z(n6183) );
  XOR2_X1 U17163 ( .A1(n9809), .A2(n27837), .Z(n22042) );
  XOR2_X1 U17165 ( .A1(n24809), .A2(n25465), .Z(n6185) );
  NAND2_X1 U17167 ( .A1(n21256), .A2(n6192), .ZN(n21261) );
  OAI21_X1 U17170 ( .A1(n18979), .A2(n18425), .B(n18978), .ZN(n6193) );
  NOR2_X1 U17172 ( .A1(n14810), .A2(n6402), .ZN(n9227) );
  AND2_X1 U17173 ( .A1(n25312), .A2(n694), .Z(n17709) );
  NOR2_X1 U17175 ( .A1(n24121), .A2(n1775), .ZN(n13748) );
  NAND2_X1 U17176 ( .A1(n8932), .A2(n16273), .ZN(n8340) );
  XOR2_X1 U17179 ( .A1(Plaintext[22]), .A2(Key[22]), .Z(n8317) );
  OR2_X1 U17192 ( .A1(n19967), .A2(n14576), .Z(n20022) );
  XOR2_X1 U17193 ( .A1(n20669), .A2(n20667), .Z(n6205) );
  AND2_X1 U17196 ( .A1(n15528), .A2(n16528), .Z(n15530) );
  XOR2_X1 U17197 ( .A1(n18903), .A2(n6209), .Z(n6281) );
  XOR2_X1 U17200 ( .A1(n24768), .A2(n6211), .Z(n7042) );
  XOR2_X1 U17201 ( .A1(n13060), .A2(n16561), .Z(n6211) );
  NAND2_X1 U17204 ( .A1(n24084), .A2(n24087), .ZN(n14912) );
  OAI21_X2 U17207 ( .A1(n11788), .A2(n10119), .B(n10116), .ZN(n24819) );
  XOR2_X1 U17213 ( .A1(Plaintext[60]), .A2(Key[60]), .Z(n6215) );
  XOR2_X1 U17228 ( .A1(n31450), .A2(n11889), .Z(n6229) );
  NAND3_X1 U17229 ( .A1(n11517), .A2(n12197), .A3(n12196), .ZN(n10694) );
  XNOR2_X1 U17237 ( .A1(n24537), .A2(n24835), .ZN(n6341) );
  XOR2_X1 U17243 ( .A1(n22044), .A2(n9129), .Z(n6245) );
  XNOR2_X1 U17245 ( .A1(n19620), .A2(n15621), .ZN(n6867) );
  CLKBUF_X2 U17246 ( .I(Key[29]), .Z(n24861) );
  NAND2_X2 U17251 ( .A1(n6252), .A2(n16763), .ZN(n19348) );
  XOR2_X1 U17253 ( .A1(n10902), .A2(n19721), .Z(n6254) );
  NAND2_X1 U17254 ( .A1(n22156), .A2(n17151), .ZN(n22665) );
  XOR2_X1 U17264 ( .A1(Plaintext[158]), .A2(Key[158]), .Z(n6265) );
  XOR2_X1 U17268 ( .A1(n24654), .A2(n1226), .Z(n6267) );
  XOR2_X1 U17269 ( .A1(n21912), .A2(n6318), .Z(n6811) );
  NAND3_X2 U17271 ( .A1(n6268), .A2(n9542), .A3(n11534), .ZN(n10146) );
  XOR2_X1 U17277 ( .A1(n20957), .A2(n474), .Z(n6273) );
  AND2_X1 U17279 ( .A1(n25628), .A2(n4146), .Z(n16096) );
  NOR2_X2 U17286 ( .A1(n8064), .A2(n8063), .ZN(n24177) );
  INV_X1 U17289 ( .I(n16828), .ZN(n16827) );
  NOR2_X2 U17297 ( .A1(n13295), .A2(n34107), .ZN(n19356) );
  AND2_X1 U17298 ( .A1(n9692), .A2(n20576), .Z(n8144) );
  OR2_X1 U17299 ( .A1(n12042), .A2(n32875), .Z(n7974) );
  INV_X2 U17300 ( .I(n6281), .ZN(n11913) );
  OAI21_X2 U17303 ( .A1(n4245), .A2(n6283), .B(n24893), .ZN(n14954) );
  XOR2_X1 U17306 ( .A1(n14239), .A2(n8575), .Z(n14238) );
  XNOR2_X1 U17309 ( .A1(n12785), .A2(n13553), .ZN(n22256) );
  XOR2_X1 U17313 ( .A1(n24823), .A2(n24548), .Z(n18042) );
  NAND3_X2 U17314 ( .A1(n11830), .A2(n16950), .A3(n29292), .ZN(n24823) );
  XOR2_X1 U17323 ( .A1(n10869), .A2(n24574), .Z(n8747) );
  NOR2_X1 U17334 ( .A1(n15302), .A2(n21530), .ZN(n12095) );
  XOR2_X1 U17341 ( .A1(n18315), .A2(Key[130]), .Z(n16462) );
  XOR2_X1 U17347 ( .A1(n20977), .A2(n14522), .Z(n9635) );
  XOR2_X1 U17353 ( .A1(n10277), .A2(n10276), .Z(n9301) );
  XOR2_X1 U17354 ( .A1(n12971), .A2(n543), .Z(n6316) );
  NAND2_X1 U17362 ( .A1(n14258), .A2(n14257), .ZN(n10783) );
  XOR2_X1 U17367 ( .A1(n14428), .A2(n20871), .Z(n6324) );
  XOR2_X1 U17372 ( .A1(n17004), .A2(n22091), .Z(n6327) );
  XOR2_X1 U17373 ( .A1(n10813), .A2(n10816), .Z(n14514) );
  XNOR2_X1 U17376 ( .A1(n24814), .A2(n11537), .ZN(n8537) );
  XOR2_X1 U17387 ( .A1(n13163), .A2(n6341), .Z(n7080) );
  XOR2_X1 U17392 ( .A1(n15743), .A2(n17938), .Z(n15754) );
  NOR2_X1 U17394 ( .A1(n16534), .A2(n10937), .ZN(n11067) );
  NAND2_X1 U17398 ( .A1(n30308), .A2(n25345), .ZN(n6345) );
  INV_X2 U17399 ( .I(n6346), .ZN(n7216) );
  XOR2_X1 U17400 ( .A1(Plaintext[104]), .A2(Key[104]), .Z(n6346) );
  XOR2_X1 U17403 ( .A1(n18109), .A2(n11604), .Z(n19690) );
  XNOR2_X1 U17410 ( .A1(n23200), .A2(n16527), .ZN(n9228) );
  XOR2_X1 U17417 ( .A1(n16080), .A2(n19673), .Z(n6721) );
  NAND2_X2 U17421 ( .A1(n12547), .A2(n12546), .ZN(n23540) );
  NOR2_X1 U17424 ( .A1(n23067), .A2(n29070), .ZN(n6677) );
  XOR2_X1 U17426 ( .A1(n23152), .A2(n23240), .Z(n22518) );
  XOR2_X1 U17427 ( .A1(n20757), .A2(n15025), .Z(n7908) );
  XOR2_X1 U17433 ( .A1(n7452), .A2(n600), .Z(n7234) );
  XOR2_X1 U17434 ( .A1(n33380), .A2(n13638), .Z(n9131) );
  NAND2_X1 U17447 ( .A1(n7897), .A2(n13318), .ZN(n6710) );
  INV_X1 U17449 ( .I(n8951), .ZN(n8950) );
  XNOR2_X1 U17452 ( .A1(n19468), .A2(n19394), .ZN(n8401) );
  XOR2_X1 U17455 ( .A1(n24116), .A2(n24375), .Z(n6397) );
  NAND2_X2 U17459 ( .A1(n1356), .A2(n7577), .ZN(n20604) );
  XOR2_X1 U17460 ( .A1(n19731), .A2(n19732), .Z(n10576) );
  NAND2_X1 U17463 ( .A1(n2471), .A2(n10310), .ZN(n22806) );
  XOR2_X1 U17465 ( .A1(n20887), .A2(n10557), .Z(n7126) );
  XOR2_X1 U17468 ( .A1(n28983), .A2(n26530), .Z(n7565) );
  OR2_X1 U17470 ( .A1(n19899), .A2(n17688), .Z(n20106) );
  AND2_X1 U17489 ( .A1(n1786), .A2(n11987), .Z(n7656) );
  INV_X1 U17491 ( .I(n25020), .ZN(n9052) );
  NOR2_X1 U17493 ( .A1(n884), .A2(n14832), .ZN(n6425) );
  OR2_X1 U17498 ( .A1(n20755), .A2(n6431), .Z(n7952) );
  INV_X2 U17501 ( .I(n6434), .ZN(n17306) );
  INV_X1 U17509 ( .I(n15581), .ZN(n15195) );
  OR2_X1 U17510 ( .A1(n15581), .A2(n22487), .Z(n11245) );
  XOR2_X1 U17513 ( .A1(n7772), .A2(n1404), .Z(n17546) );
  XOR2_X1 U17516 ( .A1(n5381), .A2(n31491), .Z(n6445) );
  XOR2_X1 U17519 ( .A1(Plaintext[19]), .A2(Key[19]), .Z(n7712) );
  XOR2_X1 U17526 ( .A1(n16717), .A2(n16718), .Z(n6452) );
  OR2_X1 U17527 ( .A1(n10435), .A2(n579), .Z(n7525) );
  XOR2_X1 U17531 ( .A1(n22132), .A2(n31105), .Z(n22134) );
  OR2_X1 U17535 ( .A1(n21374), .A2(n4145), .Z(n12110) );
  XOR2_X1 U17547 ( .A1(n16949), .A2(n6465), .Z(n6464) );
  INV_X2 U17549 ( .I(n15721), .ZN(n16568) );
  XOR2_X1 U17551 ( .A1(n24474), .A2(n24421), .Z(n24373) );
  XOR2_X1 U17552 ( .A1(n17682), .A2(n458), .Z(n24678) );
  XOR2_X1 U17554 ( .A1(n6469), .A2(n1410), .Z(Ciphertext[144]) );
  NAND3_X1 U17556 ( .A1(n28767), .A2(n16154), .A3(n29840), .ZN(n18147) );
  OR2_X1 U17563 ( .A1(n11255), .A2(n24327), .Z(n7099) );
  NOR2_X1 U17569 ( .A1(n12937), .A2(n18842), .ZN(n10451) );
  OAI21_X1 U17570 ( .A1(n24432), .A2(n27164), .B(n6477), .ZN(n24433) );
  NAND2_X1 U17571 ( .A1(n24431), .A2(n27164), .ZN(n6477) );
  NAND2_X1 U17572 ( .A1(n22588), .A2(n16562), .ZN(n22590) );
  XOR2_X1 U17573 ( .A1(n22173), .A2(n28490), .Z(n22175) );
  XOR2_X1 U17576 ( .A1(n1345), .A2(n13970), .Z(n7030) );
  XOR2_X1 U17579 ( .A1(n17549), .A2(n9764), .Z(n6485) );
  OR2_X1 U17584 ( .A1(n13059), .A2(n16916), .Z(n16788) );
  NOR2_X1 U17596 ( .A1(n18609), .A2(n18485), .ZN(n18276) );
  XOR2_X1 U17598 ( .A1(n6720), .A2(n6885), .Z(n6719) );
  NOR2_X2 U17605 ( .A1(n6504), .A2(n10128), .ZN(n17820) );
  XOR2_X1 U17606 ( .A1(n6507), .A2(n348), .Z(n8485) );
  NOR2_X2 U17609 ( .A1(n18502), .A2(n18503), .ZN(n19089) );
  XOR2_X1 U17612 ( .A1(n24389), .A2(n24600), .Z(n6513) );
  XOR2_X1 U17613 ( .A1(n21965), .A2(n6515), .Z(n15229) );
  XOR2_X1 U17617 ( .A1(n23258), .A2(n23476), .Z(n23520) );
  AND2_X1 U17622 ( .A1(n24063), .A2(n9946), .Z(n9945) );
  XOR2_X1 U17629 ( .A1(n21037), .A2(n20389), .Z(n20390) );
  AOI21_X1 U17633 ( .A1(n25742), .A2(n25741), .B(n6524), .ZN(n10082) );
  AND2_X1 U17637 ( .A1(n33078), .A2(n13200), .Z(n8662) );
  OR2_X1 U17640 ( .A1(n21666), .A2(n28618), .Z(n11584) );
  XOR2_X1 U17643 ( .A1(n6526), .A2(n16454), .Z(Ciphertext[184]) );
  XOR2_X1 U17653 ( .A1(n19574), .A2(n10866), .Z(n10865) );
  NAND3_X2 U17663 ( .A1(n22356), .A2(n22511), .A3(n13078), .ZN(n22357) );
  XOR2_X1 U17669 ( .A1(n24796), .A2(n16525), .Z(n14689) );
  NAND3_X1 U17675 ( .A1(n9148), .A2(n32186), .A3(n31862), .ZN(n9147) );
  XOR2_X1 U17676 ( .A1(n2142), .A2(n12580), .Z(n12579) );
  XOR2_X1 U17683 ( .A1(n31277), .A2(n14206), .Z(n6561) );
  XOR2_X1 U17684 ( .A1(n20863), .A2(n508), .Z(n6562) );
  OR2_X1 U17687 ( .A1(n18931), .A2(n17725), .Z(n6567) );
  XOR2_X1 U17688 ( .A1(n9018), .A2(n11586), .Z(n6572) );
  XOR2_X1 U17690 ( .A1(n7861), .A2(n7860), .Z(n6574) );
  OAI21_X1 U17691 ( .A1(n12175), .A2(n6579), .B(n13254), .ZN(n7027) );
  XOR2_X1 U17692 ( .A1(Plaintext[51]), .A2(Key[51]), .Z(n6776) );
  XOR2_X1 U17701 ( .A1(n14401), .A2(n6601), .Z(n20049) );
  XOR2_X1 U17702 ( .A1(n28822), .A2(n20836), .Z(n6601) );
  XOR2_X1 U17703 ( .A1(n14132), .A2(n2616), .Z(n14401) );
  XOR2_X1 U17704 ( .A1(Plaintext[73]), .A2(Key[73]), .Z(n18557) );
  NAND2_X1 U17707 ( .A1(n15119), .A2(n29626), .ZN(n15326) );
  NAND2_X1 U17714 ( .A1(n23033), .A2(n6605), .ZN(n22893) );
  XOR2_X1 U17719 ( .A1(n51), .A2(n25161), .Z(n6607) );
  XOR2_X1 U17722 ( .A1(n2330), .A2(n6680), .Z(n6609) );
  OAI22_X1 U17727 ( .A1(n18853), .A2(n6860), .B1(n15216), .B2(n15211), .ZN(
        n6612) );
  INV_X2 U17728 ( .I(n8400), .ZN(n15211) );
  XOR2_X1 U17731 ( .A1(n11691), .A2(n28687), .Z(n6614) );
  XOR2_X1 U17737 ( .A1(n20987), .A2(n6618), .Z(n8160) );
  XOR2_X1 U17738 ( .A1(n20754), .A2(n16666), .Z(n6618) );
  XOR2_X1 U17740 ( .A1(n24783), .A2(n6621), .Z(n6620) );
  XOR2_X1 U17741 ( .A1(n30307), .A2(n16657), .Z(n6621) );
  XOR2_X1 U17746 ( .A1(n6627), .A2(n6628), .Z(n8632) );
  XOR2_X1 U17747 ( .A1(n587), .A2(n9984), .Z(n6628) );
  NAND2_X1 U17748 ( .A1(n33702), .A2(n7555), .ZN(n12251) );
  INV_X2 U17750 ( .I(n6634), .ZN(n16854) );
  NAND2_X2 U17753 ( .A1(n6919), .A2(n6918), .ZN(n19156) );
  INV_X2 U17755 ( .I(n33393), .ZN(n25562) );
  XOR2_X1 U17758 ( .A1(n24683), .A2(n6647), .Z(n6646) );
  XOR2_X1 U17759 ( .A1(n24474), .A2(n24789), .Z(n24683) );
  XOR2_X1 U17762 ( .A1(n25191), .A2(n27385), .Z(n6647) );
  XOR2_X1 U17765 ( .A1(n1129), .A2(n28005), .Z(n6650) );
  OAI21_X2 U17767 ( .A1(n22770), .A2(n32960), .B(n15914), .ZN(n23183) );
  NOR2_X1 U17774 ( .A1(n16418), .A2(n15108), .ZN(n6668) );
  MUX2_X1 U17777 ( .I0(n14729), .I1(n19959), .S(n20112), .Z(n6672) );
  NAND3_X1 U17778 ( .A1(n6673), .A2(n13624), .A3(n30557), .ZN(n10007) );
  NAND2_X2 U17781 ( .A1(n16085), .A2(n13580), .ZN(n21665) );
  XNOR2_X1 U17782 ( .A1(n15539), .A2(n6682), .ZN(n6681) );
  XOR2_X1 U17783 ( .A1(n6683), .A2(n15538), .Z(n6682) );
  XOR2_X1 U17786 ( .A1(n6687), .A2(n6688), .Z(n6686) );
  XOR2_X1 U17792 ( .A1(n6701), .A2(n6700), .Z(n21228) );
  XOR2_X1 U17796 ( .A1(n31950), .A2(n17600), .Z(n6702) );
  INV_X2 U17798 ( .I(n14834), .ZN(n19874) );
  INV_X2 U17799 ( .I(n6705), .ZN(n11922) );
  XOR2_X1 U17800 ( .A1(n6706), .A2(n6708), .Z(n6707) );
  XOR2_X1 U17801 ( .A1(n23300), .A2(n23535), .Z(n6708) );
  XOR2_X1 U17802 ( .A1(n23301), .A2(n10201), .Z(n23124) );
  NOR2_X1 U17807 ( .A1(n29757), .A2(n19143), .ZN(n7882) );
  INV_X2 U17810 ( .I(n6725), .ZN(n25697) );
  AOI21_X2 U17811 ( .A1(n13662), .A2(n1327), .B(n6728), .ZN(n8291) );
  NAND3_X2 U17813 ( .A1(n15023), .A2(n21097), .A3(n21098), .ZN(n15022) );
  XOR2_X1 U17819 ( .A1(n20926), .A2(n25832), .Z(n6737) );
  XOR2_X1 U17822 ( .A1(n16958), .A2(n20715), .Z(n6739) );
  XOR2_X1 U17825 ( .A1(n23256), .A2(n475), .Z(n6746) );
  XOR2_X1 U17830 ( .A1(n6756), .A2(n6755), .Z(n6893) );
  XOR2_X1 U17831 ( .A1(n21033), .A2(n31950), .Z(n6755) );
  XOR2_X1 U17834 ( .A1(n6757), .A2(n4771), .Z(n6756) );
  XOR2_X1 U17837 ( .A1(n6761), .A2(n23524), .Z(n6760) );
  XOR2_X1 U17838 ( .A1(n32899), .A2(n10773), .Z(n6761) );
  XOR2_X1 U17839 ( .A1(n23367), .A2(n2520), .Z(n23524) );
  XOR2_X1 U17840 ( .A1(n8882), .A2(n23248), .Z(n6762) );
  NAND2_X1 U17844 ( .A1(n3909), .A2(n31402), .ZN(n22654) );
  AOI21_X1 U17846 ( .A1(n747), .A2(n14737), .B(n32059), .ZN(n7373) );
  XOR2_X1 U17847 ( .A1(n22285), .A2(n16344), .Z(n10422) );
  XOR2_X1 U17848 ( .A1(n24492), .A2(n7132), .Z(n15427) );
  NAND3_X2 U17849 ( .A1(n6773), .A2(n7729), .A3(n7727), .ZN(n15671) );
  INV_X1 U17854 ( .I(n12317), .ZN(n6778) );
  OAI21_X2 U17858 ( .A1(n6786), .A2(n16473), .B(n6784), .ZN(n9472) );
  XOR2_X1 U17862 ( .A1(n20978), .A2(n10424), .Z(n6790) );
  INV_X1 U17863 ( .I(Plaintext[32]), .ZN(n6791) );
  XOR2_X1 U17864 ( .A1(n6791), .A2(Key[32]), .Z(n7194) );
  INV_X2 U17865 ( .I(n7368), .ZN(n7195) );
  OR2_X1 U17866 ( .A1(n22950), .A2(n6798), .Z(n6801) );
  XOR2_X1 U17872 ( .A1(n6808), .A2(n7138), .Z(n7137) );
  XOR2_X1 U17875 ( .A1(n12614), .A2(n6810), .Z(n6809) );
  XOR2_X1 U17876 ( .A1(n9412), .A2(n24386), .Z(n6810) );
  INV_X2 U17879 ( .I(n6820), .ZN(n9162) );
  XOR2_X1 U17884 ( .A1(n6827), .A2(n16584), .Z(Ciphertext[55]) );
  NAND3_X1 U17885 ( .A1(n1075), .A2(n28736), .A3(n7555), .ZN(n6829) );
  XOR2_X1 U17895 ( .A1(n11869), .A2(n13393), .Z(n6843) );
  NOR2_X1 U17901 ( .A1(n1214), .A2(n25889), .ZN(n24718) );
  INV_X1 U17902 ( .I(n13622), .ZN(n12231) );
  NOR2_X2 U17903 ( .A1(n22326), .A2(n22325), .ZN(n16267) );
  XNOR2_X1 U17906 ( .A1(n15309), .A2(n6856), .ZN(n6854) );
  XOR2_X1 U17907 ( .A1(n29285), .A2(n20998), .Z(n6856) );
  XOR2_X1 U17908 ( .A1(n15), .A2(n25436), .Z(n11374) );
  NAND3_X1 U17915 ( .A1(n6200), .A2(n6263), .A3(n4674), .ZN(n6866) );
  XOR2_X1 U17920 ( .A1(n21036), .A2(n21037), .Z(n6872) );
  NOR2_X1 U17921 ( .A1(n580), .A2(n1158), .ZN(n20616) );
  NAND2_X1 U17923 ( .A1(n14559), .A2(n16489), .ZN(n6930) );
  XOR2_X1 U17924 ( .A1(n19741), .A2(n25880), .Z(n6885) );
  XOR2_X1 U17925 ( .A1(n27156), .A2(n19424), .Z(n19673) );
  INV_X2 U17929 ( .I(n6893), .ZN(n12044) );
  XOR2_X1 U17935 ( .A1(n24638), .A2(n16581), .Z(n6897) );
  XOR2_X1 U17936 ( .A1(n9145), .A2(n24394), .Z(n24505) );
  XOR2_X1 U17938 ( .A1(n15886), .A2(n11194), .Z(n6903) );
  XOR2_X1 U17939 ( .A1(n21019), .A2(n6906), .Z(n20700) );
  NAND2_X1 U17942 ( .A1(n27501), .A2(n30586), .ZN(n9846) );
  NAND2_X1 U17943 ( .A1(n27501), .A2(n24158), .ZN(n24313) );
  XOR2_X1 U17945 ( .A1(n19705), .A2(n487), .Z(n6914) );
  AOI21_X1 U17946 ( .A1(n16854), .A2(n18459), .B(n7216), .ZN(n6921) );
  XOR2_X1 U17949 ( .A1(n32880), .A2(n23474), .Z(n6923) );
  XOR2_X1 U17952 ( .A1(n3322), .A2(n12059), .Z(n6924) );
  NAND2_X1 U17955 ( .A1(n21612), .A2(n17472), .ZN(n6937) );
  INV_X2 U17956 ( .I(n6938), .ZN(n6939) );
  XOR2_X1 U17958 ( .A1(n24377), .A2(n6941), .Z(n6940) );
  XOR2_X1 U17959 ( .A1(n24559), .A2(n1411), .Z(n6941) );
  INV_X2 U17964 ( .I(n6955), .ZN(n12076) );
  INV_X2 U17966 ( .I(n6957), .ZN(n21165) );
  XOR2_X1 U17970 ( .A1(n10159), .A2(n16301), .Z(n6966) );
  AOI21_X1 U17972 ( .A1(n19915), .A2(n19914), .B(n6970), .ZN(n19916) );
  XOR2_X1 U17974 ( .A1(n24771), .A2(n25610), .Z(n6973) );
  NAND2_X1 U17977 ( .A1(n18041), .A2(n2606), .ZN(n6999) );
  INV_X2 U17988 ( .I(n7020), .ZN(n16650) );
  INV_X2 U17990 ( .I(n7022), .ZN(n13905) );
  INV_X2 U17992 ( .I(n21970), .ZN(n7023) );
  XOR2_X1 U17994 ( .A1(n22167), .A2(n11027), .Z(n7025) );
  XOR2_X1 U17995 ( .A1(n7030), .A2(n7031), .Z(n7029) );
  NAND2_X1 U18000 ( .A1(n8820), .A2(n31968), .ZN(n8819) );
  NOR2_X1 U18003 ( .A1(n9985), .A2(n27901), .ZN(n11635) );
  XOR2_X1 U18004 ( .A1(n9467), .A2(n7042), .Z(n7043) );
  INV_X2 U18005 ( .I(n7043), .ZN(n25700) );
  OAI21_X1 U18010 ( .A1(n468), .A2(n2417), .B(n11250), .ZN(n7052) );
  AOI22_X2 U18013 ( .A1(n7055), .A2(n7116), .B1(n8353), .B2(n7054), .ZN(n20776) );
  XOR2_X1 U18014 ( .A1(n7057), .A2(n30305), .Z(n14415) );
  XOR2_X1 U18017 ( .A1(n29137), .A2(n25560), .Z(n13435) );
  XOR2_X1 U18024 ( .A1(n23362), .A2(n7823), .Z(n7071) );
  NOR2_X1 U18028 ( .A1(n7073), .A2(n12906), .ZN(n7077) );
  XOR2_X1 U18029 ( .A1(n3739), .A2(n24895), .Z(n9867) );
  XOR2_X1 U18030 ( .A1(n7078), .A2(n24836), .Z(n18138) );
  INV_X2 U18031 ( .I(n7080), .ZN(n25232) );
  INV_X2 U18032 ( .I(n17214), .ZN(n7081) );
  NOR2_X1 U18038 ( .A1(n10018), .A2(n7088), .ZN(n23221) );
  NAND2_X1 U18042 ( .A1(n11255), .A2(n24245), .ZN(n24128) );
  NOR2_X1 U18046 ( .A1(n22868), .A2(n28555), .ZN(n22869) );
  NAND2_X1 U18047 ( .A1(n23050), .A2(n28555), .ZN(n9950) );
  XOR2_X1 U18048 ( .A1(n23224), .A2(n1414), .Z(n11586) );
  XOR2_X1 U18049 ( .A1(n17929), .A2(n23224), .Z(n12387) );
  XOR2_X1 U18053 ( .A1(n20839), .A2(n20892), .Z(n7113) );
  INV_X2 U18056 ( .I(n21971), .ZN(n22411) );
  XOR2_X1 U18057 ( .A1(n7114), .A2(n21901), .Z(n21971) );
  INV_X2 U18061 ( .I(n7250), .ZN(n10205) );
  INV_X2 U18062 ( .I(n7124), .ZN(n8490) );
  XNOR2_X1 U18063 ( .A1(n7126), .A2(n7125), .ZN(n7124) );
  XOR2_X1 U18064 ( .A1(n15823), .A2(n20671), .Z(n7125) );
  XOR2_X1 U18066 ( .A1(n9222), .A2(n13739), .Z(n7129) );
  XOR2_X1 U18069 ( .A1(n10331), .A2(n16703), .Z(n7132) );
  XOR2_X1 U18072 ( .A1(n20837), .A2(n20860), .Z(n20978) );
  NAND2_X2 U18073 ( .A1(n20425), .A2(n20424), .ZN(n20837) );
  NAND2_X1 U18075 ( .A1(n7140), .A2(n13281), .ZN(n7139) );
  XOR2_X1 U18076 ( .A1(n22105), .A2(n12127), .Z(n7152) );
  XOR2_X1 U18079 ( .A1(n22318), .A2(n22295), .Z(n22273) );
  NAND2_X1 U18080 ( .A1(n16811), .A2(n19907), .ZN(n20118) );
  AOI21_X2 U18084 ( .A1(n18577), .A2(n33941), .B(n7162), .ZN(n7161) );
  OR2_X1 U18085 ( .A1(n16854), .A2(n11379), .Z(n7164) );
  NAND3_X1 U18090 ( .A1(n26232), .A2(n6230), .A3(n26471), .ZN(n20583) );
  XOR2_X1 U18102 ( .A1(n16005), .A2(n19763), .Z(n19469) );
  INV_X2 U18104 ( .I(n7194), .ZN(n15146) );
  NOR2_X1 U18108 ( .A1(n14940), .A2(n25995), .ZN(n7369) );
  NAND3_X1 U18115 ( .A1(n10511), .A2(n24991), .A3(n10510), .ZN(n7212) );
  NAND3_X1 U18117 ( .A1(n9320), .A2(n14436), .A3(n7218), .ZN(n9692) );
  XOR2_X1 U18120 ( .A1(n4157), .A2(n16527), .Z(n7222) );
  NOR2_X1 U18121 ( .A1(n17640), .A2(n4971), .ZN(n7224) );
  INV_X2 U18122 ( .I(n18197), .ZN(n21170) );
  XOR2_X1 U18125 ( .A1(n19699), .A2(n5150), .Z(n7938) );
  XOR2_X1 U18129 ( .A1(n16053), .A2(n7229), .Z(n23342) );
  NOR3_X1 U18133 ( .A1(n7776), .A2(n7775), .A3(n7232), .ZN(n7774) );
  XOR2_X1 U18135 ( .A1(n21041), .A2(n18010), .Z(n7235) );
  NAND2_X1 U18138 ( .A1(n21517), .A2(n21847), .ZN(n7241) );
  XOR2_X1 U18144 ( .A1(n7259), .A2(n7258), .Z(n7257) );
  XOR2_X1 U18145 ( .A1(n24796), .A2(n16696), .Z(n7258) );
  XOR2_X1 U18153 ( .A1(n31523), .A2(n24065), .Z(n23452) );
  XOR2_X1 U18160 ( .A1(n7294), .A2(n1405), .Z(n9608) );
  XOR2_X1 U18161 ( .A1(n21044), .A2(n28983), .Z(n14785) );
  NAND2_X2 U18163 ( .A1(n20368), .A2(n20367), .ZN(n7294) );
  XOR2_X1 U18165 ( .A1(n19733), .A2(n7296), .Z(n7295) );
  XOR2_X1 U18166 ( .A1(n15117), .A2(n16703), .Z(n7296) );
  NAND2_X1 U18168 ( .A1(n7303), .A2(n27920), .ZN(n7298) );
  NOR2_X1 U18169 ( .A1(n7301), .A2(n7300), .ZN(n7299) );
  NOR3_X1 U18170 ( .A1(n7305), .A2(n15359), .A3(n25206), .ZN(n7300) );
  NOR2_X1 U18171 ( .A1(n7304), .A2(n25206), .ZN(n7301) );
  NOR2_X1 U18173 ( .A1(n10750), .A2(n7308), .ZN(n7307) );
  NAND3_X1 U18179 ( .A1(n5834), .A2(n18683), .A3(n30116), .ZN(n7318) );
  NOR2_X1 U18180 ( .A1(n26049), .A2(n18683), .ZN(n9476) );
  XOR2_X1 U18182 ( .A1(n20688), .A2(n7331), .Z(n7328) );
  XOR2_X1 U18184 ( .A1(n32749), .A2(n16687), .Z(n7331) );
  XOR2_X1 U18186 ( .A1(n7336), .A2(n25881), .Z(Ciphertext[183]) );
  XOR2_X1 U18191 ( .A1(n16693), .A2(n7352), .Z(n24798) );
  XOR2_X1 U18192 ( .A1(n16128), .A2(n24741), .Z(n7352) );
  XOR2_X1 U18204 ( .A1(n7381), .A2(n14748), .Z(n7380) );
  XOR2_X1 U18205 ( .A1(n23511), .A2(n16482), .Z(n7382) );
  XOR2_X1 U18207 ( .A1(n24603), .A2(n15573), .Z(n12935) );
  XOR2_X1 U18208 ( .A1(n7387), .A2(n2363), .Z(n14391) );
  OR2_X1 U18214 ( .A1(n20387), .A2(n53), .Z(n7395) );
  OR2_X1 U18215 ( .A1(n18899), .A2(n878), .Z(n7402) );
  XOR2_X1 U18221 ( .A1(n23230), .A2(n12252), .Z(n15055) );
  AND2_X1 U18223 ( .A1(n22716), .A2(n22808), .Z(n7412) );
  INV_X1 U18225 ( .I(n7413), .ZN(n10567) );
  NAND2_X1 U18226 ( .A1(n16274), .A2(n9553), .ZN(n7417) );
  NOR2_X1 U18227 ( .A1(n28707), .A2(n7496), .ZN(n17368) );
  XOR2_X1 U18229 ( .A1(n7431), .A2(n7432), .Z(n11942) );
  XOR2_X1 U18230 ( .A1(n21045), .A2(n8526), .Z(n7432) );
  XOR2_X1 U18235 ( .A1(n25991), .A2(n1405), .Z(n7450) );
  NOR2_X1 U18237 ( .A1(n1063), .A2(n18792), .ZN(n18794) );
  XOR2_X1 U18238 ( .A1(n18350), .A2(Key[30]), .Z(n15265) );
  XOR2_X1 U18248 ( .A1(n7471), .A2(n7470), .Z(n7469) );
  XOR2_X1 U18249 ( .A1(n4997), .A2(n16604), .Z(n7470) );
  XOR2_X1 U18251 ( .A1(n10869), .A2(n24774), .Z(n7472) );
  NAND2_X1 U18252 ( .A1(n9025), .A2(n11312), .ZN(n11311) );
  OAI21_X2 U18258 ( .A1(n20299), .A2(n14835), .B(n20554), .ZN(n20698) );
  NOR2_X1 U18262 ( .A1(n4024), .A2(n24201), .ZN(n7485) );
  NAND2_X1 U18269 ( .A1(n470), .A2(n7496), .ZN(n7495) );
  NOR2_X1 U18270 ( .A1(n31407), .A2(n25317), .ZN(n11998) );
  NAND2_X1 U18281 ( .A1(n15906), .A2(n7525), .ZN(n9381) );
  XOR2_X1 U18283 ( .A1(n28953), .A2(n5024), .Z(n13209) );
  XOR2_X1 U18284 ( .A1(n400), .A2(n7530), .Z(n9373) );
  XOR2_X1 U18285 ( .A1(n27275), .A2(n7530), .Z(n8053) );
  INV_X2 U18291 ( .I(n10770), .ZN(n24780) );
  XOR2_X1 U18292 ( .A1(n4240), .A2(n1404), .Z(n7537) );
  INV_X1 U18303 ( .I(n12609), .ZN(n21042) );
  XOR2_X1 U18306 ( .A1(n31277), .A2(n33693), .Z(n7569) );
  INV_X2 U18308 ( .I(n7573), .ZN(n18089) );
  OAI21_X1 U18309 ( .A1(n24657), .A2(n24656), .B(n7576), .ZN(n24659) );
  NAND2_X1 U18310 ( .A1(n31428), .A2(n10325), .ZN(n18889) );
  XOR2_X1 U18317 ( .A1(n8785), .A2(n1365), .Z(n7589) );
  XOR2_X1 U18318 ( .A1(n33749), .A2(n19675), .Z(n7590) );
  NAND2_X1 U18320 ( .A1(n25115), .A2(n18156), .ZN(n25020) );
  XOR2_X1 U18324 ( .A1(n7595), .A2(n5024), .Z(n7594) );
  XOR2_X1 U18328 ( .A1(n17395), .A2(n7598), .Z(n7597) );
  XOR2_X1 U18329 ( .A1(n30331), .A2(n30906), .Z(n7598) );
  XOR2_X1 U18330 ( .A1(n12760), .A2(n16974), .Z(n7599) );
  NOR2_X1 U18331 ( .A1(n7600), .A2(n19255), .ZN(n15040) );
  AOI21_X2 U18332 ( .A1(n24676), .A2(n24799), .B(n7604), .ZN(n17811) );
  XOR2_X1 U18333 ( .A1(n17811), .A2(n16972), .Z(n7605) );
  XOR2_X1 U18334 ( .A1(n13236), .A2(n1432), .Z(n7606) );
  NOR2_X1 U18335 ( .A1(n7609), .A2(n12038), .ZN(n19997) );
  XOR2_X1 U18337 ( .A1(n7611), .A2(n9641), .Z(n9640) );
  XOR2_X1 U18338 ( .A1(n9006), .A2(n10210), .Z(n7611) );
  XOR2_X1 U18340 ( .A1(n23245), .A2(n7615), .Z(n7614) );
  XOR2_X1 U18341 ( .A1(n23186), .A2(n16605), .Z(n7615) );
  XOR2_X1 U18343 ( .A1(n32930), .A2(n19582), .Z(n7619) );
  XOR2_X1 U18346 ( .A1(n20904), .A2(n25610), .Z(n7622) );
  XOR2_X1 U18347 ( .A1(n8795), .A2(n20905), .Z(n7623) );
  INV_X1 U18348 ( .I(n32051), .ZN(n18518) );
  INV_X2 U18350 ( .I(n7624), .ZN(n25889) );
  XOR2_X1 U18352 ( .A1(n20736), .A2(n1923), .Z(n7628) );
  AOI22_X2 U18353 ( .A1(n9852), .A2(n16050), .B1(n7631), .B2(n14011), .ZN(
        n20614) );
  XOR2_X1 U18354 ( .A1(n19588), .A2(n7635), .Z(n7634) );
  XOR2_X1 U18355 ( .A1(n29890), .A2(n207), .Z(n7635) );
  XOR2_X1 U18360 ( .A1(n29011), .A2(n16464), .Z(n7638) );
  XOR2_X1 U18363 ( .A1(n21910), .A2(n21958), .Z(n22046) );
  XOR2_X1 U18368 ( .A1(n20648), .A2(n7645), .Z(n7644) );
  XOR2_X1 U18369 ( .A1(n20996), .A2(n12957), .Z(n7645) );
  XOR2_X1 U18370 ( .A1(n20698), .A2(n20954), .Z(n20648) );
  XOR2_X1 U18371 ( .A1(n19703), .A2(n27281), .Z(n7652) );
  XOR2_X1 U18372 ( .A1(n32581), .A2(n25465), .Z(n20858) );
  INV_X2 U18378 ( .I(n7657), .ZN(n21070) );
  NOR2_X1 U18379 ( .A1(n4202), .A2(n30010), .ZN(n9315) );
  NOR2_X1 U18381 ( .A1(n8408), .A2(n23867), .ZN(n7663) );
  INV_X2 U18382 ( .I(n15356), .ZN(n19938) );
  XOR2_X1 U18384 ( .A1(n2894), .A2(n24917), .Z(n7664) );
  XOR2_X1 U18386 ( .A1(n8997), .A2(n25131), .Z(n7675) );
  XOR2_X1 U18388 ( .A1(n19632), .A2(n1196), .Z(n7676) );
  XOR2_X1 U18394 ( .A1(n22076), .A2(n22158), .Z(n21919) );
  NAND2_X1 U18396 ( .A1(n12358), .A2(n7689), .ZN(n7688) );
  XOR2_X1 U18399 ( .A1(n29318), .A2(n1397), .Z(n7693) );
  XOR2_X1 U18400 ( .A1(n356), .A2(n25990), .Z(n7694) );
  INV_X2 U18404 ( .I(n7700), .ZN(n8408) );
  NAND2_X2 U18406 ( .A1(n17022), .A2(n17023), .ZN(n7702) );
  NOR2_X1 U18407 ( .A1(n25916), .A2(n7701), .ZN(n25907) );
  NOR2_X1 U18409 ( .A1(n31476), .A2(n1018), .ZN(n21272) );
  INV_X2 U18413 ( .I(n7712), .ZN(n16420) );
  NAND2_X1 U18414 ( .A1(n9272), .A2(n1287), .ZN(n11866) );
  MUX2_X1 U18418 ( .I0(n26950), .I1(n9323), .S(n7809), .Z(n7730) );
  XOR2_X1 U18420 ( .A1(n7731), .A2(n16687), .Z(n11484) );
  NOR2_X1 U18421 ( .A1(n8862), .A2(n7732), .ZN(n8867) );
  NAND2_X1 U18425 ( .A1(n2444), .A2(n1244), .ZN(n23621) );
  NAND2_X1 U18426 ( .A1(n24111), .A2(n1244), .ZN(n24112) );
  NOR2_X1 U18427 ( .A1(n15977), .A2(n1244), .ZN(n10177) );
  INV_X2 U18431 ( .I(n7912), .ZN(n10187) );
  XOR2_X1 U18435 ( .A1(n9904), .A2(n33749), .Z(n7741) );
  AOI22_X2 U18440 ( .A1(n7745), .A2(n22864), .B1(n7744), .B2(n14978), .ZN(
        n23262) );
  NAND2_X1 U18442 ( .A1(n31019), .A2(n12488), .ZN(n17268) );
  XOR2_X1 U18447 ( .A1(n7838), .A2(n17296), .Z(n7761) );
  OAI21_X1 U18449 ( .A1(n25154), .A2(n7765), .B(n25175), .ZN(n16098) );
  XOR2_X1 U18452 ( .A1(n7772), .A2(n16355), .Z(n23472) );
  AOI21_X1 U18457 ( .A1(n3994), .A2(n24936), .B(n15799), .ZN(n7785) );
  XOR2_X1 U18462 ( .A1(n7794), .A2(n7793), .Z(n24870) );
  XOR2_X1 U18463 ( .A1(n28258), .A2(n7795), .Z(n7793) );
  XOR2_X1 U18465 ( .A1(n30301), .A2(n7511), .Z(n7795) );
  INV_X1 U18467 ( .I(n14201), .ZN(n22855) );
  NAND2_X1 U18470 ( .A1(n29253), .A2(n27345), .ZN(n7803) );
  XOR2_X1 U18473 ( .A1(n7808), .A2(n14300), .Z(n14299) );
  XOR2_X1 U18477 ( .A1(n31950), .A2(n16038), .Z(n16754) );
  XOR2_X1 U18478 ( .A1(n27708), .A2(n25036), .Z(n7823) );
  XOR2_X1 U18484 ( .A1(n7828), .A2(n16530), .Z(n7829) );
  NOR2_X1 U18487 ( .A1(n24995), .A2(n7831), .ZN(n14450) );
  OR2_X1 U18492 ( .A1(n25677), .A2(n25678), .Z(n7842) );
  XOR2_X1 U18494 ( .A1(n22139), .A2(n30332), .Z(n16837) );
  XOR2_X1 U18498 ( .A1(n7859), .A2(n18231), .Z(n11220) );
  XOR2_X1 U18499 ( .A1(n24826), .A2(n1426), .Z(n7860) );
  XOR2_X1 U18500 ( .A1(n28579), .A2(n12313), .Z(n7861) );
  INV_X2 U18503 ( .I(n7865), .ZN(n13969) );
  XOR2_X1 U18504 ( .A1(n15357), .A2(n15819), .Z(n7866) );
  XOR2_X1 U18505 ( .A1(n1341), .A2(n7960), .Z(n7870) );
  XOR2_X1 U18508 ( .A1(n16080), .A2(n7875), .Z(n7874) );
  XOR2_X1 U18519 ( .A1(n13457), .A2(n7888), .Z(n13491) );
  XOR2_X1 U18521 ( .A1(n20906), .A2(n447), .Z(n7890) );
  NAND2_X1 U18524 ( .A1(n7895), .A2(n1099), .ZN(n23649) );
  NAND2_X1 U18525 ( .A1(n7895), .A2(n27455), .ZN(n23348) );
  NOR2_X1 U18529 ( .A1(n6215), .A2(n1430), .ZN(n7900) );
  XOR2_X1 U18530 ( .A1(Plaintext[65]), .A2(Key[65]), .Z(n18186) );
  XOR2_X1 U18533 ( .A1(n24686), .A2(n10924), .Z(n24524) );
  AOI21_X2 U18534 ( .A1(n11121), .A2(n28120), .B(n24169), .ZN(n24686) );
  XOR2_X1 U18537 ( .A1(n7910), .A2(n7909), .Z(n14307) );
  XOR2_X1 U18538 ( .A1(n16896), .A2(n15778), .Z(n7909) );
  XOR2_X1 U18539 ( .A1(n12495), .A2(n7911), .Z(n7910) );
  XOR2_X1 U18543 ( .A1(n23121), .A2(n22948), .Z(n7916) );
  XOR2_X1 U18544 ( .A1(n23184), .A2(n22954), .Z(n7917) );
  NAND2_X1 U18545 ( .A1(n8467), .A2(n17439), .ZN(n8466) );
  INV_X2 U18546 ( .I(n7918), .ZN(n17439) );
  XOR2_X1 U18548 ( .A1(n17766), .A2(n15121), .Z(n7931) );
  NAND2_X2 U18550 ( .A1(n21742), .A2(n14041), .ZN(n9960) );
  XOR2_X1 U18551 ( .A1(n11784), .A2(n7934), .Z(n7933) );
  XOR2_X1 U18552 ( .A1(n22294), .A2(n22295), .Z(n7934) );
  XOR2_X1 U18555 ( .A1(n7939), .A2(n7936), .Z(n12241) );
  XOR2_X1 U18556 ( .A1(n7937), .A2(n7938), .Z(n7936) );
  NAND2_X1 U18559 ( .A1(n713), .A2(n7941), .ZN(n14451) );
  NAND2_X2 U18560 ( .A1(n13940), .A2(n9422), .ZN(n19230) );
  OAI21_X2 U18561 ( .A1(n21310), .A2(n21447), .B(n21309), .ZN(n21662) );
  XOR2_X1 U18566 ( .A1(n22168), .A2(n28926), .Z(n22247) );
  AND2_X1 U18571 ( .A1(n19130), .A2(n7966), .Z(n16363) );
  INV_X2 U18572 ( .I(n11379), .ZN(n18459) );
  XOR2_X1 U18579 ( .A1(n19546), .A2(n19690), .Z(n7988) );
  XOR2_X1 U18581 ( .A1(n19734), .A2(n19401), .Z(n7989) );
  INV_X2 U18583 ( .I(n7993), .ZN(n23795) );
  XOR2_X1 U18585 ( .A1(n7999), .A2(n22250), .Z(n7998) );
  XOR2_X1 U18590 ( .A1(n8701), .A2(n17999), .Z(n8700) );
  XOR2_X1 U18593 ( .A1(n23393), .A2(n16454), .Z(n8018) );
  XOR2_X1 U18595 ( .A1(n8021), .A2(n23403), .Z(n8020) );
  XOR2_X1 U18596 ( .A1(n11193), .A2(n27613), .Z(n8021) );
  NAND2_X1 U18601 ( .A1(n12827), .A2(n8029), .ZN(n8030) );
  XOR2_X1 U18602 ( .A1(n27169), .A2(n3929), .Z(n20695) );
  INV_X2 U18604 ( .I(n14788), .ZN(n17110) );
  XOR2_X1 U18605 ( .A1(n10617), .A2(n10616), .Z(n14788) );
  NAND2_X2 U18607 ( .A1(n17959), .A2(n22527), .ZN(n22983) );
  INV_X2 U18609 ( .I(n8042), .ZN(n23742) );
  XOR2_X1 U18619 ( .A1(n8050), .A2(n24646), .Z(n24411) );
  XOR2_X1 U18622 ( .A1(n13339), .A2(n1024), .Z(n13338) );
  INV_X1 U18624 ( .I(n9481), .ZN(n9479) );
  NAND2_X2 U18631 ( .A1(n19241), .A2(n19240), .ZN(n19676) );
  NOR2_X2 U18632 ( .A1(n19239), .A2(n19238), .ZN(n19779) );
  NOR2_X1 U18633 ( .A1(n8058), .A2(n24106), .ZN(n14375) );
  NOR2_X1 U18634 ( .A1(n17310), .A2(n8058), .ZN(n12098) );
  XOR2_X1 U18636 ( .A1(n8060), .A2(n8059), .Z(n8721) );
  XOR2_X1 U18638 ( .A1(n27130), .A2(n16060), .Z(n8061) );
  NOR2_X1 U18641 ( .A1(n13102), .A2(n23930), .ZN(n8063) );
  XOR2_X1 U18643 ( .A1(n32895), .A2(n8066), .Z(n8065) );
  XOR2_X1 U18644 ( .A1(n23519), .A2(n25465), .Z(n8066) );
  XOR2_X1 U18645 ( .A1(n23518), .A2(n23520), .Z(n8067) );
  XOR2_X1 U18648 ( .A1(n23125), .A2(n15049), .Z(n8070) );
  AOI21_X1 U18651 ( .A1(n712), .A2(n14810), .B(n6402), .ZN(n25125) );
  XOR2_X1 U18655 ( .A1(n22296), .A2(n16381), .Z(n21878) );
  XOR2_X1 U18657 ( .A1(n16138), .A2(n16110), .Z(n8089) );
  NOR2_X2 U18667 ( .A1(n21306), .A2(n21305), .ZN(n8106) );
  XOR2_X1 U18673 ( .A1(n13695), .A2(n25009), .Z(n8112) );
  XOR2_X1 U18674 ( .A1(n14899), .A2(n20318), .Z(n8116) );
  XOR2_X1 U18676 ( .A1(n23387), .A2(n25772), .Z(n8129) );
  XOR2_X1 U18677 ( .A1(n10205), .A2(n1064), .Z(n22194) );
  XOR2_X1 U18678 ( .A1(n8133), .A2(n8132), .Z(n9871) );
  XOR2_X1 U18679 ( .A1(n21927), .A2(n10429), .Z(n8132) );
  XOR2_X1 U18683 ( .A1(n30729), .A2(n8139), .Z(n12103) );
  XOR2_X1 U18684 ( .A1(n30729), .A2(n16631), .Z(n19316) );
  NAND2_X2 U18686 ( .A1(n18769), .A2(n17905), .ZN(n8141) );
  NAND2_X2 U18694 ( .A1(n12371), .A2(n12373), .ZN(n8313) );
  NAND2_X2 U18697 ( .A1(n21609), .A2(n21608), .ZN(n22021) );
  NAND2_X1 U18702 ( .A1(n32605), .A2(n22608), .ZN(n12112) );
  OAI21_X1 U18706 ( .A1(n18583), .A2(n12190), .B(n18582), .ZN(n12191) );
  NOR2_X1 U18715 ( .A1(n22690), .A2(n16205), .ZN(n9603) );
  OAI21_X1 U18716 ( .A1(n17709), .A2(n17708), .B(n8629), .ZN(n11558) );
  OAI21_X1 U18718 ( .A1(n15858), .A2(n32867), .B(n25312), .ZN(n15857) );
  XOR2_X1 U18725 ( .A1(n11434), .A2(n11432), .Z(n16904) );
  NAND2_X2 U18727 ( .A1(n8481), .A2(n11347), .ZN(n9247) );
  INV_X1 U18730 ( .I(n12498), .ZN(n12497) );
  XOR2_X1 U18736 ( .A1(Plaintext[170]), .A2(Key[170]), .Z(n18411) );
  XOR2_X1 U18738 ( .A1(n19587), .A2(n32844), .Z(n15044) );
  NAND2_X1 U18748 ( .A1(n21653), .A2(n21595), .ZN(n21596) );
  OR2_X1 U18749 ( .A1(n29658), .A2(n8208), .Z(n10786) );
  NOR2_X1 U18756 ( .A1(n24328), .A2(n10987), .ZN(n10342) );
  INV_X2 U18757 ( .I(n18182), .ZN(n10213) );
  INV_X2 U18760 ( .I(n8213), .ZN(n18880) );
  XOR2_X1 U18762 ( .A1(n24845), .A2(n8215), .Z(n8214) );
  NAND2_X1 U18764 ( .A1(n23105), .A2(n22971), .ZN(n11623) );
  OAI22_X1 U18772 ( .A1(n19022), .A2(n19023), .B1(n19021), .B2(n19290), .ZN(
        n8227) );
  AOI21_X1 U18773 ( .A1(n17850), .A2(n25463), .B(n25470), .ZN(n17849) );
  INV_X2 U18774 ( .I(n8228), .ZN(n9133) );
  XOR2_X1 U18778 ( .A1(n1341), .A2(n11636), .Z(n8232) );
  XOR2_X1 U18785 ( .A1(n8236), .A2(n31094), .Z(Ciphertext[122]) );
  NAND3_X1 U18786 ( .A1(n25548), .A2(n17401), .A3(n25547), .ZN(n8236) );
  XOR2_X1 U18787 ( .A1(n24578), .A2(n14250), .Z(n17504) );
  XOR2_X1 U18792 ( .A1(n8241), .A2(n30275), .Z(n11271) );
  INV_X1 U18793 ( .I(n9536), .ZN(n8241) );
  NAND2_X1 U18803 ( .A1(n7144), .A2(n21876), .ZN(n8253) );
  XNOR2_X1 U18806 ( .A1(n32255), .A2(n22078), .ZN(n9208) );
  NOR2_X1 U18812 ( .A1(n881), .A2(n6295), .ZN(n18318) );
  OR2_X1 U18813 ( .A1(n15397), .A2(n19330), .Z(n19155) );
  XOR2_X1 U18814 ( .A1(n8556), .A2(n14429), .Z(n14534) );
  XOR2_X1 U18821 ( .A1(n11574), .A2(n8266), .Z(n8265) );
  NOR2_X1 U18824 ( .A1(n4373), .A2(n16848), .ZN(n19818) );
  NAND2_X1 U18825 ( .A1(n17670), .A2(n33561), .ZN(n12253) );
  AOI21_X1 U18830 ( .A1(n23108), .A2(n6453), .B(n23111), .ZN(n9042) );
  XOR2_X1 U18837 ( .A1(n22099), .A2(n22031), .Z(n8282) );
  OAI21_X1 U18844 ( .A1(n17877), .A2(n298), .B(n11257), .ZN(n17876) );
  INV_X1 U18849 ( .I(n21160), .ZN(n21139) );
  XOR2_X1 U18855 ( .A1(n20710), .A2(n20709), .Z(n11542) );
  OR2_X1 U18859 ( .A1(n17403), .A2(n13483), .Z(n25548) );
  NAND2_X1 U18860 ( .A1(n11646), .A2(n28203), .ZN(n11645) );
  AND2_X1 U18864 ( .A1(n1099), .A2(n29323), .Z(n12026) );
  OR3_X1 U18869 ( .A1(n17156), .A2(n17155), .A3(n4587), .Z(n10850) );
  XOR2_X1 U18870 ( .A1(n12342), .A2(n20921), .Z(n20758) );
  INV_X1 U18872 ( .I(n9612), .ZN(n9611) );
  AND2_X1 U18885 ( .A1(n10574), .A2(n27149), .Z(n9676) );
  NOR2_X1 U18890 ( .A1(n10549), .A2(n18219), .ZN(n8470) );
  NOR2_X1 U18893 ( .A1(n23670), .A2(n29198), .ZN(n9344) );
  XOR2_X1 U18895 ( .A1(n12681), .A2(n22221), .Z(n8324) );
  XOR2_X1 U18900 ( .A1(n8557), .A2(n8987), .Z(n10372) );
  NOR2_X2 U18907 ( .A1(n11983), .A2(n31854), .ZN(n22781) );
  AND2_X1 U18910 ( .A1(n21676), .A2(n15595), .Z(n8331) );
  OR2_X1 U18911 ( .A1(n18955), .A2(n18983), .Z(n18964) );
  AND3_X1 U18915 ( .A1(n14321), .A2(n24995), .A3(n24996), .Z(n9901) );
  XOR2_X1 U18919 ( .A1(n21892), .A2(n30332), .Z(n10963) );
  XOR2_X1 U18928 ( .A1(n8341), .A2(n14216), .Z(n22156) );
  NAND2_X1 U18929 ( .A1(n9273), .A2(n6908), .ZN(n8958) );
  XOR2_X1 U18934 ( .A1(n8345), .A2(n16402), .Z(Ciphertext[172]) );
  XOR2_X1 U18941 ( .A1(n22018), .A2(n521), .Z(n8352) );
  XOR2_X1 U18946 ( .A1(n8361), .A2(n11600), .Z(n9753) );
  XOR2_X1 U18948 ( .A1(n21885), .A2(n16439), .Z(n17109) );
  XOR2_X1 U18953 ( .A1(n14400), .A2(n8364), .Z(n12670) );
  XOR2_X1 U18954 ( .A1(n14647), .A2(n14646), .Z(n8364) );
  XOR2_X1 U18956 ( .A1(n11282), .A2(n8366), .Z(n11281) );
  NAND3_X1 U18965 ( .A1(n10897), .A2(n27162), .A3(n25851), .ZN(n18021) );
  XOR2_X1 U18968 ( .A1(n19406), .A2(n445), .Z(n8383) );
  AND2_X1 U18977 ( .A1(n11987), .A2(n28591), .Z(n14895) );
  XOR2_X1 U18984 ( .A1(n8394), .A2(n25910), .Z(Ciphertext[188]) );
  NAND2_X2 U18986 ( .A1(n12690), .A2(n12689), .ZN(n8457) );
  XOR2_X1 U18987 ( .A1(n10916), .A2(n10914), .Z(n14834) );
  NOR2_X1 U18988 ( .A1(n8397), .A2(n25416), .ZN(n25417) );
  AOI21_X1 U18989 ( .A1(n25415), .A2(n25418), .B(n25452), .ZN(n8397) );
  XOR2_X1 U18994 ( .A1(Key[159]), .A2(Plaintext[159]), .Z(n8400) );
  INV_X4 U18995 ( .I(n9162), .ZN(n14922) );
  INV_X2 U18997 ( .I(n20091), .ZN(n19936) );
  XOR2_X1 U18998 ( .A1(n14222), .A2(n8401), .Z(n20091) );
  INV_X1 U18999 ( .I(n16007), .ZN(n14611) );
  AND2_X1 U19000 ( .A1(n16275), .A2(n599), .Z(n12743) );
  NOR2_X1 U19001 ( .A1(n21590), .A2(n7144), .ZN(n8402) );
  XOR2_X1 U19003 ( .A1(n10076), .A2(n8405), .Z(n22390) );
  XOR2_X1 U19008 ( .A1(n27852), .A2(n322), .Z(n8413) );
  NAND2_X2 U19012 ( .A1(n985), .A2(n9280), .ZN(n8786) );
  INV_X2 U19014 ( .I(n10860), .ZN(n11198) );
  XOR2_X1 U19015 ( .A1(n10861), .A2(n8416), .Z(n10860) );
  XOR2_X1 U19021 ( .A1(Plaintext[94]), .A2(Key[94]), .Z(n16782) );
  INV_X2 U19023 ( .I(n8422), .ZN(n10080) );
  XOR2_X1 U19026 ( .A1(n11320), .A2(n15565), .Z(n8424) );
  XNOR2_X1 U19029 ( .A1(n22014), .A2(n16587), .ZN(n8979) );
  INV_X2 U19038 ( .I(n8435), .ZN(n19947) );
  XOR2_X1 U19043 ( .A1(n8440), .A2(n1426), .Z(Ciphertext[33]) );
  INV_X1 U19045 ( .I(n17578), .ZN(n23870) );
  NOR2_X1 U19047 ( .A1(n29294), .A2(n10187), .ZN(n10753) );
  INV_X2 U19050 ( .I(n8444), .ZN(n11945) );
  XOR2_X1 U19051 ( .A1(n14886), .A2(n14883), .Z(n8444) );
  XNOR2_X1 U19065 ( .A1(n19773), .A2(n13826), .ZN(n15188) );
  OR2_X1 U19072 ( .A1(n21490), .A2(n21489), .Z(n8463) );
  NAND2_X1 U19077 ( .A1(n34097), .A2(n15976), .ZN(n11740) );
  INV_X2 U19078 ( .I(n8469), .ZN(n21109) );
  INV_X2 U19080 ( .I(n10372), .ZN(n25867) );
  XOR2_X1 U19082 ( .A1(n6569), .A2(n16701), .Z(n8475) );
  OR2_X1 U19084 ( .A1(n17879), .A2(n22580), .Z(n22348) );
  NAND2_X1 U19099 ( .A1(n31549), .A2(n23103), .ZN(n8494) );
  XOR2_X1 U19101 ( .A1(n10391), .A2(n8496), .Z(n10390) );
  XOR2_X1 U19103 ( .A1(n3722), .A2(n22078), .Z(n8497) );
  XOR2_X1 U19108 ( .A1(n8997), .A2(n8500), .Z(n11066) );
  INV_X1 U19111 ( .I(n9839), .ZN(n10886) );
  INV_X2 U19114 ( .I(n8505), .ZN(n11920) );
  XOR2_X1 U19115 ( .A1(n14298), .A2(n14301), .Z(n8505) );
  XOR2_X1 U19116 ( .A1(n24777), .A2(n24778), .Z(n16719) );
  XOR2_X1 U19117 ( .A1(n8507), .A2(n24643), .Z(n24777) );
  NAND2_X1 U19120 ( .A1(n25804), .A2(n25818), .ZN(n25819) );
  NOR2_X2 U19123 ( .A1(n8515), .A2(n9956), .ZN(n25072) );
  XNOR2_X1 U19125 ( .A1(n19544), .A2(n19446), .ZN(n16678) );
  XOR2_X1 U19128 ( .A1(n24679), .A2(n24678), .Z(n24680) );
  XOR2_X1 U19132 ( .A1(n8949), .A2(n25878), .Z(n8531) );
  XOR2_X1 U19133 ( .A1(n19742), .A2(n13222), .Z(n8532) );
  NAND2_X1 U19134 ( .A1(n23822), .A2(n11887), .ZN(n18152) );
  XOR2_X1 U19135 ( .A1(n8536), .A2(n16587), .Z(Ciphertext[60]) );
  NAND2_X1 U19137 ( .A1(n14531), .A2(n25140), .ZN(n15228) );
  XOR2_X1 U19142 ( .A1(n23196), .A2(n16160), .Z(n23373) );
  NAND2_X1 U19145 ( .A1(n8542), .A2(n8541), .ZN(n10100) );
  NOR2_X1 U19148 ( .A1(n21478), .A2(n32904), .ZN(n9590) );
  AND2_X1 U19150 ( .A1(n23882), .A2(n8544), .Z(n10621) );
  INV_X2 U19153 ( .I(n8545), .ZN(n11966) );
  AOI22_X1 U19157 ( .A1(n25153), .A2(n25179), .B1(n14531), .B2(n25174), .ZN(
        n17635) );
  NAND2_X2 U19161 ( .A1(n8551), .A2(n8550), .ZN(n19104) );
  XOR2_X1 U19162 ( .A1(n24762), .A2(n24541), .Z(n14886) );
  OAI21_X2 U19166 ( .A1(n11318), .A2(n11319), .B(n8554), .ZN(n18257) );
  XOR2_X1 U19169 ( .A1(n24793), .A2(n17858), .Z(n8557) );
  XOR2_X1 U19172 ( .A1(n19698), .A2(n23239), .Z(n8561) );
  XOR2_X1 U19174 ( .A1(n19527), .A2(n19526), .Z(n20137) );
  NAND2_X1 U19176 ( .A1(n8664), .A2(n24276), .ZN(n8663) );
  NAND2_X1 U19186 ( .A1(n19233), .A2(n19274), .ZN(n9407) );
  OAI21_X2 U19190 ( .A1(n8581), .A2(n11636), .B(n8578), .ZN(n12539) );
  XOR2_X1 U19192 ( .A1(n1340), .A2(n11349), .Z(n8583) );
  NAND2_X1 U19194 ( .A1(n32857), .A2(n28228), .ZN(n25089) );
  XOR2_X1 U19200 ( .A1(n19503), .A2(n13829), .Z(n10060) );
  NOR2_X1 U19211 ( .A1(n19229), .A2(n8606), .ZN(n11807) );
  INV_X2 U19218 ( .I(n18541), .ZN(n13279) );
  XOR2_X1 U19222 ( .A1(n8633), .A2(n16679), .Z(n13951) );
  XOR2_X1 U19223 ( .A1(n8633), .A2(n12998), .Z(n12519) );
  INV_X2 U19224 ( .I(n8634), .ZN(n17895) );
  XOR2_X1 U19226 ( .A1(n8480), .A2(n25827), .Z(n8635) );
  INV_X2 U19228 ( .I(n24947), .ZN(n24958) );
  XOR2_X1 U19232 ( .A1(n32243), .A2(n8659), .Z(n23390) );
  INV_X1 U19233 ( .I(Plaintext[33]), .ZN(n8666) );
  XOR2_X1 U19234 ( .A1(n8666), .A2(Key[33]), .Z(n10058) );
  NOR2_X1 U19237 ( .A1(n25787), .A2(n8678), .ZN(n16670) );
  OAI21_X1 U19239 ( .A1(n25798), .A2(n26753), .B(n12611), .ZN(n25799) );
  NAND2_X1 U19240 ( .A1(n25782), .A2(n26753), .ZN(n17222) );
  INV_X2 U19243 ( .I(n8681), .ZN(n21253) );
  XOR2_X1 U19245 ( .A1(n31491), .A2(n25619), .Z(n23307) );
  XOR2_X1 U19247 ( .A1(n19589), .A2(n13826), .Z(n8685) );
  XOR2_X1 U19249 ( .A1(n19644), .A2(n19368), .Z(n19446) );
  INV_X1 U19252 ( .I(n29130), .ZN(n19337) );
  XOR2_X1 U19253 ( .A1(n29130), .A2(n25167), .Z(n13843) );
  XOR2_X1 U19255 ( .A1(n31279), .A2(n1432), .Z(n13854) );
  INV_X2 U19259 ( .I(n8694), .ZN(n23695) );
  XOR2_X1 U19261 ( .A1(Plaintext[166]), .A2(Key[166]), .Z(n18860) );
  NAND2_X1 U19262 ( .A1(n4683), .A2(n8010), .ZN(n16543) );
  XOR2_X1 U19263 ( .A1(n24539), .A2(n24454), .Z(n24398) );
  XOR2_X1 U19268 ( .A1(n8707), .A2(n24869), .Z(Ciphertext[115]) );
  OAI21_X1 U19269 ( .A1(n8766), .A2(n25515), .B(n25509), .ZN(n8708) );
  NOR2_X1 U19270 ( .A1(n8766), .A2(n25516), .ZN(n8709) );
  XOR2_X1 U19272 ( .A1(n8718), .A2(n9263), .Z(n8715) );
  AOI21_X1 U19274 ( .A1(n28736), .A2(n7555), .B(n25129), .ZN(n8722) );
  INV_X1 U19277 ( .I(n19164), .ZN(n9652) );
  INV_X1 U19278 ( .I(n8237), .ZN(n15029) );
  XOR2_X1 U19279 ( .A1(n28889), .A2(n11490), .Z(n19785) );
  XOR2_X1 U19281 ( .A1(n29838), .A2(n16696), .Z(n16949) );
  XOR2_X1 U19282 ( .A1(n29838), .A2(n25091), .Z(n20709) );
  AOI21_X1 U19283 ( .A1(n17814), .A2(n33480), .B(n25902), .ZN(n17621) );
  NOR2_X1 U19284 ( .A1(n11754), .A2(n1090), .ZN(n8731) );
  NAND2_X2 U19285 ( .A1(n21597), .A2(n21596), .ZN(n22210) );
  NAND2_X1 U19287 ( .A1(n13663), .A2(n11918), .ZN(n8737) );
  AOI21_X1 U19290 ( .A1(n8212), .A2(n8742), .B(n33672), .ZN(n14500) );
  XOR2_X1 U19295 ( .A1(n8747), .A2(n8745), .Z(n10171) );
  XOR2_X1 U19296 ( .A1(n10729), .A2(n8746), .Z(n8745) );
  XOR2_X1 U19297 ( .A1(n11332), .A2(n1193), .Z(n8746) );
  XOR2_X1 U19300 ( .A1(n11166), .A2(n22210), .Z(n8750) );
  XOR2_X1 U19307 ( .A1(n19677), .A2(n8755), .Z(n8754) );
  XOR2_X1 U19313 ( .A1(n8765), .A2(n8763), .Z(n10463) );
  XOR2_X1 U19314 ( .A1(n23190), .A2(n8764), .Z(n8763) );
  XOR2_X1 U19315 ( .A1(n29235), .A2(n1064), .Z(n8764) );
  XOR2_X1 U19316 ( .A1(n29217), .A2(n29299), .Z(n23190) );
  NAND2_X1 U19317 ( .A1(n8770), .A2(n31522), .ZN(n8769) );
  XOR2_X1 U19318 ( .A1(n19739), .A2(n19211), .Z(n8771) );
  XOR2_X1 U19320 ( .A1(n31755), .A2(n12620), .Z(n8772) );
  NAND2_X1 U19322 ( .A1(n17655), .A2(n30316), .ZN(n8773) );
  XOR2_X1 U19323 ( .A1(n32894), .A2(n1427), .Z(n8774) );
  NAND2_X1 U19326 ( .A1(n31161), .A2(n1172), .ZN(n8782) );
  XOR2_X1 U19327 ( .A1(n8791), .A2(n12355), .Z(n10350) );
  XOR2_X1 U19335 ( .A1(n12958), .A2(n8806), .Z(n8808) );
  XOR2_X1 U19338 ( .A1(n23163), .A2(n8812), .Z(n8811) );
  XOR2_X1 U19339 ( .A1(n23260), .A2(n16533), .Z(n8812) );
  XOR2_X1 U19342 ( .A1(Plaintext[79]), .A2(Key[79]), .Z(n16881) );
  XOR2_X1 U19346 ( .A1(n14858), .A2(n1065), .Z(n8826) );
  XNOR2_X1 U19348 ( .A1(Plaintext[119]), .A2(Key[119]), .ZN(n8832) );
  XOR2_X1 U19350 ( .A1(n8845), .A2(n8843), .Z(n17641) );
  XOR2_X1 U19352 ( .A1(n32870), .A2(n24618), .Z(n8844) );
  NAND2_X1 U19363 ( .A1(n8860), .A2(n18738), .ZN(n18124) );
  NAND2_X1 U19364 ( .A1(n25744), .A2(n1597), .ZN(n25740) );
  NAND2_X1 U19365 ( .A1(n25737), .A2(n25748), .ZN(n25742) );
  XOR2_X1 U19366 ( .A1(n30314), .A2(n22274), .Z(n8861) );
  NOR3_X1 U19369 ( .A1(n18261), .A2(n30365), .A3(n25979), .ZN(n8876) );
  XOR2_X1 U19375 ( .A1(n23247), .A2(n8883), .Z(n8882) );
  INV_X2 U19379 ( .I(n34169), .ZN(n25590) );
  OR2_X1 U19380 ( .A1(n34169), .A2(n8892), .Z(n25529) );
  XOR2_X1 U19383 ( .A1(n24624), .A2(n8895), .Z(n8894) );
  XOR2_X1 U19384 ( .A1(n24625), .A2(n13556), .Z(n8896) );
  XOR2_X1 U19385 ( .A1(n9217), .A2(n609), .Z(n8899) );
  INV_X2 U19386 ( .I(n8899), .ZN(n21056) );
  NOR2_X1 U19387 ( .A1(n8901), .A2(n25587), .ZN(n10395) );
  MUX2_X1 U19388 ( .I0(n24075), .I1(n24127), .S(n1235), .Z(n24078) );
  XOR2_X1 U19391 ( .A1(n24689), .A2(n25065), .Z(n17325) );
  XOR2_X1 U19392 ( .A1(n24689), .A2(n24964), .Z(n10195) );
  XOR2_X1 U19393 ( .A1(n23209), .A2(n1196), .Z(n8916) );
  XOR2_X1 U19394 ( .A1(n23257), .A2(n15497), .Z(n8917) );
  XOR2_X1 U19395 ( .A1(n24764), .A2(n25036), .Z(n8920) );
  XOR2_X1 U19396 ( .A1(n4028), .A2(n480), .Z(n8922) );
  NAND2_X1 U19397 ( .A1(n8207), .A2(n28196), .ZN(n16279) );
  NAND2_X1 U19398 ( .A1(n25154), .A2(n8926), .ZN(n25140) );
  OAI21_X1 U19400 ( .A1(n16273), .A2(n8207), .B(n8925), .ZN(n25160) );
  INV_X2 U19402 ( .I(n8933), .ZN(n12168) );
  NAND2_X1 U19403 ( .A1(n5966), .A2(n12168), .ZN(n8934) );
  NOR2_X1 U19406 ( .A1(n8944), .A2(n32193), .ZN(n22529) );
  INV_X2 U19408 ( .I(n9626), .ZN(n21452) );
  NAND2_X2 U19414 ( .A1(n14773), .A2(n14772), .ZN(n22871) );
  XOR2_X1 U19416 ( .A1(n15114), .A2(n1197), .Z(n8974) );
  XOR2_X1 U19417 ( .A1(n8976), .A2(n13190), .Z(n8975) );
  XOR2_X1 U19418 ( .A1(n23503), .A2(n28927), .Z(n8976) );
  XOR2_X1 U19421 ( .A1(n21964), .A2(n1065), .Z(n8992) );
  XOR2_X1 U19424 ( .A1(n22036), .A2(n17723), .Z(n9000) );
  INV_X1 U19425 ( .I(n20515), .ZN(n20174) );
  XOR2_X1 U19426 ( .A1(n9005), .A2(n9004), .Z(n11051) );
  INV_X2 U19429 ( .I(n11051), .ZN(n15110) );
  XOR2_X1 U19432 ( .A1(n23419), .A2(n24861), .Z(n9011) );
  XOR2_X1 U19433 ( .A1(n23359), .A2(n15897), .Z(n9013) );
  XOR2_X1 U19435 ( .A1(n11836), .A2(n9021), .Z(n9020) );
  XOR2_X1 U19436 ( .A1(n11897), .A2(n16301), .Z(n9021) );
  XOR2_X1 U19443 ( .A1(n8347), .A2(n14557), .Z(n9038) );
  NAND2_X1 U19445 ( .A1(n936), .A2(n26566), .ZN(n20313) );
  MUX2_X1 U19446 ( .I0(n20578), .I1(n20579), .S(n8528), .Z(n20585) );
  XOR2_X1 U19447 ( .A1(n19719), .A2(n9045), .Z(n9044) );
  XOR2_X1 U19448 ( .A1(n19763), .A2(n25104), .Z(n9045) );
  INV_X2 U19452 ( .I(n9064), .ZN(n12952) );
  NAND2_X1 U19454 ( .A1(n24308), .A2(n11041), .ZN(n12575) );
  XOR2_X1 U19458 ( .A1(n9907), .A2(n24953), .Z(n9087) );
  XOR2_X1 U19459 ( .A1(n16237), .A2(n25319), .Z(n12084) );
  XOR2_X1 U19460 ( .A1(n22114), .A2(n1307), .Z(n22115) );
  XOR2_X1 U19463 ( .A1(n19616), .A2(n18902), .Z(n18903) );
  XOR2_X1 U19465 ( .A1(n13586), .A2(n16672), .Z(n9092) );
  NAND2_X1 U19467 ( .A1(n19997), .A2(n19986), .ZN(n9098) );
  XOR2_X1 U19469 ( .A1(n19641), .A2(n25224), .Z(n9101) );
  XOR2_X1 U19470 ( .A1(n19686), .A2(n15117), .Z(n9102) );
  XOR2_X1 U19476 ( .A1(n16351), .A2(n19787), .Z(n9116) );
  XNOR2_X1 U19479 ( .A1(Plaintext[114]), .A2(Key[114]), .ZN(n9118) );
  XOR2_X1 U19487 ( .A1(n343), .A2(n22173), .Z(n21961) );
  AOI22_X1 U19492 ( .A1(n19336), .A2(n12815), .B1(n12316), .B2(n16699), .ZN(
        n9134) );
  XOR2_X1 U19495 ( .A1(n21926), .A2(n13303), .Z(n9136) );
  XOR2_X1 U19496 ( .A1(n19530), .A2(n32981), .Z(n9138) );
  XOR2_X1 U19497 ( .A1(n9141), .A2(n16402), .Z(n13856) );
  NOR2_X1 U19499 ( .A1(n31969), .A2(n27600), .ZN(n20359) );
  NAND2_X1 U19500 ( .A1(n10312), .A2(n31969), .ZN(n20239) );
  NAND2_X1 U19501 ( .A1(n19865), .A2(n31969), .ZN(n13246) );
  XOR2_X1 U19502 ( .A1(n23206), .A2(n23207), .Z(n9154) );
  AOI21_X2 U19509 ( .A1(n11470), .A2(n9174), .B(n18651), .ZN(n11085) );
  NAND2_X1 U19513 ( .A1(n11754), .A2(n31155), .ZN(n16090) );
  NAND2_X1 U19514 ( .A1(n1238), .A2(n24118), .ZN(n9178) );
  INV_X1 U19515 ( .I(n25818), .ZN(n25822) );
  NOR2_X1 U19517 ( .A1(n9182), .A2(n9181), .ZN(n9180) );
  NAND2_X2 U19518 ( .A1(n18491), .A2(n9183), .ZN(n18990) );
  XOR2_X1 U19520 ( .A1(n9185), .A2(n16390), .Z(n12580) );
  INV_X2 U19521 ( .I(n19255), .ZN(n19256) );
  NAND2_X1 U19531 ( .A1(n12143), .A2(n9219), .ZN(n12430) );
  XOR2_X1 U19533 ( .A1(n26562), .A2(n32881), .Z(n14902) );
  XOR2_X1 U19536 ( .A1(n9231), .A2(n9988), .Z(n9230) );
  OAI21_X1 U19538 ( .A1(n14503), .A2(n21662), .B(n32898), .ZN(n13803) );
  INV_X2 U19543 ( .I(n9239), .ZN(n11944) );
  XOR2_X1 U19545 ( .A1(n16693), .A2(n15147), .Z(n9241) );
  NAND2_X1 U19547 ( .A1(n830), .A2(n4770), .ZN(n9249) );
  NOR2_X2 U19549 ( .A1(n9014), .A2(n14005), .ZN(n9255) );
  XOR2_X1 U19553 ( .A1(n16586), .A2(n4975), .Z(n19522) );
  XOR2_X1 U19555 ( .A1(n24787), .A2(n25131), .Z(n9281) );
  NAND2_X2 U19557 ( .A1(n14161), .A2(n14005), .ZN(n20219) );
  XOR2_X1 U19560 ( .A1(n9290), .A2(n22099), .Z(n22165) );
  INV_X1 U19561 ( .I(n8386), .ZN(n9305) );
  INV_X1 U19566 ( .I(n10325), .ZN(n9296) );
  XOR2_X1 U19568 ( .A1(n26931), .A2(n22273), .Z(n9298) );
  NAND2_X1 U19574 ( .A1(n11264), .A2(n9302), .ZN(n19882) );
  XOR2_X1 U19576 ( .A1(n9303), .A2(n16662), .Z(n10557) );
  XOR2_X1 U19577 ( .A1(n9303), .A2(n1343), .Z(n20702) );
  XOR2_X1 U19578 ( .A1(n9308), .A2(n7603), .Z(n9307) );
  XOR2_X1 U19579 ( .A1(n9309), .A2(n9310), .Z(n11238) );
  XOR2_X1 U19580 ( .A1(n9311), .A2(n22310), .Z(n9309) );
  XOR2_X1 U19581 ( .A1(n16971), .A2(n21887), .Z(n9310) );
  XOR2_X1 U19584 ( .A1(n19464), .A2(n11361), .Z(n9325) );
  AND3_X1 U19588 ( .A1(n23950), .A2(n10187), .A3(n33659), .Z(n9345) );
  XOR2_X1 U19589 ( .A1(n23234), .A2(n9349), .Z(n9347) );
  XOR2_X1 U19591 ( .A1(n23438), .A2(n30557), .Z(n9349) );
  XOR2_X1 U19595 ( .A1(n14211), .A2(n9362), .Z(n9361) );
  XOR2_X1 U19596 ( .A1(n19682), .A2(n16680), .Z(n9362) );
  AOI21_X2 U19607 ( .A1(n13112), .A2(n13111), .B(n13110), .ZN(n19283) );
  XOR2_X1 U19609 ( .A1(n24441), .A2(n24505), .Z(n9385) );
  NAND3_X2 U19610 ( .A1(n24278), .A2(n14288), .A3(n24279), .ZN(n24475) );
  XOR2_X1 U19611 ( .A1(n21949), .A2(n9388), .Z(n9387) );
  XOR2_X1 U19612 ( .A1(n22033), .A2(n25669), .Z(n9388) );
  XOR2_X1 U19616 ( .A1(n16838), .A2(n544), .Z(n11995) );
  XOR2_X1 U19619 ( .A1(n9412), .A2(n17679), .Z(n21949) );
  XOR2_X1 U19620 ( .A1(n9412), .A2(n25751), .Z(n22142) );
  XOR2_X1 U19625 ( .A1(Plaintext[132]), .A2(Key[132]), .Z(n9437) );
  INV_X2 U19628 ( .I(n9920), .ZN(n23862) );
  INV_X2 U19633 ( .I(n9437), .ZN(n18537) );
  NAND2_X1 U19639 ( .A1(n9446), .A2(n22946), .ZN(n16921) );
  XOR2_X1 U19640 ( .A1(n22182), .A2(n9447), .Z(n16617) );
  XOR2_X1 U19641 ( .A1(n9960), .A2(n27281), .Z(n9447) );
  XOR2_X1 U19657 ( .A1(n11751), .A2(n1403), .Z(n9475) );
  INV_X2 U19662 ( .I(n9486), .ZN(n25763) );
  XOR2_X1 U19663 ( .A1(n16838), .A2(n9488), .Z(n9487) );
  XOR2_X1 U19664 ( .A1(n24533), .A2(n27157), .Z(n9488) );
  NAND2_X2 U19668 ( .A1(n21089), .A2(n21090), .ZN(n21687) );
  XOR2_X1 U19670 ( .A1(n9504), .A2(n27137), .Z(n9503) );
  XOR2_X1 U19671 ( .A1(n18453), .A2(n25881), .Z(n9504) );
  XOR2_X1 U19672 ( .A1(n1305), .A2(n27180), .Z(n9505) );
  XOR2_X1 U19673 ( .A1(n20736), .A2(n20996), .Z(n20738) );
  XOR2_X1 U19674 ( .A1(n9507), .A2(n20542), .Z(n10788) );
  NOR2_X1 U19675 ( .A1(n13548), .A2(n13514), .ZN(n9513) );
  XOR2_X1 U19678 ( .A1(n29312), .A2(n9527), .Z(n9526) );
  XOR2_X1 U19680 ( .A1(n9533), .A2(n9529), .Z(n9535) );
  XOR2_X1 U19681 ( .A1(n9532), .A2(n9530), .Z(n9529) );
  XOR2_X1 U19682 ( .A1(n22210), .A2(n9531), .Z(n9530) );
  NAND2_X2 U19685 ( .A1(n9540), .A2(n9539), .ZN(n19335) );
  AOI21_X1 U19687 ( .A1(n33594), .A2(n22641), .B(n22645), .ZN(n9544) );
  XOR2_X1 U19690 ( .A1(n23397), .A2(n9551), .Z(n9550) );
  XOR2_X1 U19691 ( .A1(n15183), .A2(n25693), .Z(n9551) );
  INV_X2 U19692 ( .I(n9564), .ZN(n11957) );
  XOR2_X1 U19694 ( .A1(n27015), .A2(n9568), .Z(n9567) );
  XOR2_X1 U19696 ( .A1(n9209), .A2(n24809), .Z(n9573) );
  XOR2_X1 U19697 ( .A1(n24808), .A2(n10583), .Z(n9574) );
  XOR2_X1 U19705 ( .A1(n29718), .A2(n1192), .Z(n9599) );
  XOR2_X1 U19709 ( .A1(n9606), .A2(n9604), .Z(n17218) );
  XOR2_X1 U19710 ( .A1(n27375), .A2(n9605), .Z(n9604) );
  NOR2_X1 U19711 ( .A1(n9612), .A2(n25235), .ZN(n9609) );
  NAND2_X1 U19715 ( .A1(n22414), .A2(n9617), .ZN(n15581) );
  XOR2_X1 U19716 ( .A1(n9623), .A2(n9621), .Z(n22394) );
  XOR2_X1 U19717 ( .A1(n9622), .A2(n21967), .Z(n9621) );
  XOR2_X1 U19718 ( .A1(n31457), .A2(n13651), .Z(n9622) );
  XOR2_X1 U19719 ( .A1(n22183), .A2(n14994), .Z(n9623) );
  XOR2_X1 U19721 ( .A1(n10169), .A2(n453), .Z(n9634) );
  INV_X2 U19726 ( .I(n9640), .ZN(n19998) );
  XOR2_X1 U19727 ( .A1(n19168), .A2(n18915), .Z(n9641) );
  NAND2_X1 U19729 ( .A1(n25193), .A2(n27149), .ZN(n13266) );
  AOI21_X1 U19730 ( .A1(n830), .A2(n25194), .B(n27149), .ZN(n9675) );
  XOR2_X1 U19733 ( .A1(n6484), .A2(n25156), .Z(n9650) );
  AND2_X1 U19736 ( .A1(n3148), .A2(n23995), .Z(n9658) );
  NAND3_X1 U19737 ( .A1(n31960), .A2(n7182), .A3(n27954), .ZN(n9896) );
  XOR2_X1 U19740 ( .A1(n9665), .A2(n16472), .Z(n10986) );
  XOR2_X1 U19743 ( .A1(n13777), .A2(n23232), .Z(n9672) );
  NOR2_X1 U19745 ( .A1(n25985), .A2(n9677), .ZN(n10853) );
  XOR2_X1 U19747 ( .A1(n11860), .A2(n21582), .Z(n9679) );
  NOR2_X1 U19749 ( .A1(n1358), .A2(n13327), .ZN(n11013) );
  NOR2_X1 U19750 ( .A1(n29338), .A2(n1358), .ZN(n14693) );
  AOI22_X1 U19753 ( .A1(n9696), .A2(n29085), .B1(n27123), .B2(n9247), .ZN(
        n9695) );
  NAND3_X1 U19754 ( .A1(n13266), .A2(n4781), .A3(n9698), .ZN(n9697) );
  NAND2_X1 U19755 ( .A1(n10858), .A2(n4953), .ZN(n9698) );
  NAND2_X1 U19759 ( .A1(n13245), .A2(n9703), .ZN(n9705) );
  NAND3_X1 U19760 ( .A1(n29085), .A2(n786), .A3(n9247), .ZN(n9704) );
  XOR2_X1 U19761 ( .A1(n646), .A2(n27171), .Z(n14818) );
  XOR2_X1 U19762 ( .A1(n12821), .A2(n646), .Z(n23075) );
  XOR2_X1 U19763 ( .A1(n1262), .A2(n646), .Z(n23469) );
  INV_X1 U19765 ( .I(n14179), .ZN(n15661) );
  NOR2_X1 U19767 ( .A1(n9729), .A2(n18711), .ZN(n13566) );
  NOR2_X1 U19768 ( .A1(n1835), .A2(n9729), .ZN(n18317) );
  OAI21_X1 U19773 ( .A1(n22807), .A2(n3614), .B(n851), .ZN(n22809) );
  NAND2_X1 U19774 ( .A1(n15457), .A2(n3614), .ZN(n12782) );
  NAND2_X1 U19775 ( .A1(n22403), .A2(n22678), .ZN(n9739) );
  XOR2_X1 U19779 ( .A1(n22158), .A2(n22205), .Z(n10626) );
  XOR2_X1 U19783 ( .A1(n22137), .A2(n11863), .Z(n9758) );
  XOR2_X1 U19789 ( .A1(n11897), .A2(n16698), .Z(n9764) );
  XOR2_X1 U19791 ( .A1(n32660), .A2(n24923), .Z(n24578) );
  XOR2_X1 U19792 ( .A1(n32660), .A2(n15653), .Z(n24453) );
  XOR2_X1 U19793 ( .A1(Plaintext[23]), .A2(Key[23]), .Z(n9930) );
  NOR2_X1 U19795 ( .A1(n11943), .A2(n16320), .ZN(n9768) );
  XOR2_X1 U19799 ( .A1(n9782), .A2(n9780), .Z(n9798) );
  XOR2_X1 U19800 ( .A1(n9781), .A2(n15963), .Z(n9780) );
  XOR2_X1 U19801 ( .A1(n23450), .A2(n16160), .Z(n9781) );
  NOR2_X2 U19803 ( .A1(n13384), .A2(n14552), .ZN(n23196) );
  NOR2_X1 U19808 ( .A1(n28581), .A2(n9793), .ZN(n11658) );
  OAI22_X1 U19810 ( .A1(n9811), .A2(n8886), .B1(n21585), .B2(n9793), .ZN(
        n10825) );
  NAND2_X1 U19811 ( .A1(n12095), .A2(n9793), .ZN(n11656) );
  NOR2_X1 U19813 ( .A1(n953), .A2(n4868), .ZN(n18573) );
  XOR2_X1 U19817 ( .A1(n9819), .A2(n9820), .Z(n9818) );
  XOR2_X1 U19818 ( .A1(n32286), .A2(n19703), .Z(n9820) );
  XOR2_X1 U19819 ( .A1(n19426), .A2(n16381), .Z(n9822) );
  XOR2_X1 U19826 ( .A1(n9843), .A2(n17986), .Z(n23248) );
  NAND2_X1 U19827 ( .A1(n9847), .A2(n9846), .ZN(n9933) );
  NAND2_X1 U19830 ( .A1(n31155), .A2(n24117), .ZN(n10118) );
  NAND2_X1 U19831 ( .A1(n1238), .A2(n24225), .ZN(n12068) );
  XOR2_X1 U19834 ( .A1(n20727), .A2(n1428), .Z(n13339) );
  XOR2_X1 U19838 ( .A1(n9863), .A2(n23242), .Z(n23447) );
  XOR2_X1 U19841 ( .A1(n23255), .A2(n9867), .Z(n9866) );
  INV_X2 U19853 ( .I(n14676), .ZN(n15089) );
  NOR2_X1 U19856 ( .A1(n16908), .A2(n12144), .ZN(n16907) );
  OR2_X1 U19859 ( .A1(n20556), .A2(n20236), .Z(n20170) );
  XOR2_X1 U19865 ( .A1(n11304), .A2(n9878), .Z(n9877) );
  XOR2_X1 U19866 ( .A1(n16708), .A2(n25038), .Z(n9878) );
  XOR2_X1 U19869 ( .A1(n24846), .A2(n25772), .Z(n17296) );
  INV_X2 U19872 ( .I(n11413), .ZN(n11676) );
  XOR2_X1 U19874 ( .A1(n9904), .A2(n19513), .Z(n19514) );
  XOR2_X1 U19878 ( .A1(n9907), .A2(n11370), .Z(n24546) );
  XOR2_X1 U19887 ( .A1(n16081), .A2(n24374), .Z(n9928) );
  INV_X2 U19888 ( .I(n9929), .ZN(n19857) );
  NAND3_X1 U19890 ( .A1(n25867), .A2(n700), .A3(n10062), .ZN(n11253) );
  NOR2_X2 U19902 ( .A1(n13071), .A2(n13070), .ZN(n9951) );
  XOR2_X1 U19903 ( .A1(n30943), .A2(n19479), .Z(n9955) );
  XOR2_X1 U19906 ( .A1(n356), .A2(n25054), .Z(n12918) );
  XOR2_X1 U19907 ( .A1(n24750), .A2(n356), .Z(n13824) );
  INV_X2 U19909 ( .I(n9968), .ZN(n11898) );
  XOR2_X1 U19910 ( .A1(n9969), .A2(n13438), .Z(Ciphertext[2]) );
  INV_X1 U19913 ( .I(n19322), .ZN(n19324) );
  OAI21_X2 U19916 ( .A1(n29282), .A2(n14004), .B(n9978), .ZN(n20630) );
  OAI21_X1 U19918 ( .A1(n25613), .A2(n9982), .B(n9981), .ZN(n10265) );
  XOR2_X1 U19920 ( .A1(n15275), .A2(n20996), .Z(n9984) );
  INV_X1 U19921 ( .I(n20479), .ZN(n9985) );
  XOR2_X1 U19923 ( .A1(n17040), .A2(n13388), .Z(n9993) );
  NOR2_X1 U19924 ( .A1(n21825), .A2(n9994), .ZN(n21829) );
  NAND2_X1 U19926 ( .A1(n30878), .A2(n28288), .ZN(n10764) );
  NAND3_X1 U19930 ( .A1(n10011), .A2(n10385), .A3(n16520), .ZN(n10010) );
  XOR2_X1 U19936 ( .A1(Plaintext[148]), .A2(Key[148]), .Z(n15519) );
  INV_X1 U19939 ( .I(Plaintext[83]), .ZN(n10044) );
  XOR2_X1 U19940 ( .A1(n10044), .A2(Key[83]), .Z(n18575) );
  AOI21_X2 U19943 ( .A1(n12837), .A2(n14537), .B(n10055), .ZN(n19108) );
  INV_X2 U19946 ( .I(n10058), .ZN(n13514) );
  XOR2_X1 U19947 ( .A1(Plaintext[35]), .A2(Key[35]), .Z(n13531) );
  AOI21_X1 U19951 ( .A1(n17489), .A2(n14108), .B(n10062), .ZN(n17488) );
  XOR2_X1 U19952 ( .A1(n770), .A2(n16263), .Z(n10064) );
  INV_X2 U19957 ( .I(n21228), .ZN(n21443) );
  XOR2_X1 U19959 ( .A1(n19517), .A2(n26005), .Z(n10077) );
  NAND2_X1 U19961 ( .A1(n23868), .A2(n844), .ZN(n12603) );
  XOR2_X1 U19963 ( .A1(n10082), .A2(n1405), .Z(Ciphertext[160]) );
  XOR2_X1 U19965 ( .A1(n10084), .A2(n32814), .Z(n24698) );
  XOR2_X1 U19967 ( .A1(n10088), .A2(n10090), .Z(n25710) );
  XOR2_X1 U19968 ( .A1(n24597), .A2(n10089), .Z(n10088) );
  XOR2_X1 U19969 ( .A1(n24556), .A2(n24382), .Z(n10090) );
  NAND2_X1 U19972 ( .A1(n11046), .A2(n10097), .ZN(n24864) );
  INV_X1 U19973 ( .I(n10099), .ZN(n10098) );
  NAND2_X2 U19975 ( .A1(n20316), .A2(n20315), .ZN(n20872) );
  XOR2_X1 U19977 ( .A1(n15710), .A2(n23453), .Z(n23180) );
  NOR2_X1 U19978 ( .A1(n28344), .A2(n18349), .ZN(n12013) );
  XNOR2_X1 U19979 ( .A1(Plaintext[40]), .A2(Key[40]), .ZN(n10114) );
  NOR2_X1 U19980 ( .A1(n24225), .A2(n24118), .ZN(n10119) );
  XOR2_X1 U19983 ( .A1(n32791), .A2(n24917), .Z(n10122) );
  XOR2_X1 U19985 ( .A1(n19634), .A2(n24623), .Z(n10123) );
  INV_X2 U19986 ( .I(n17820), .ZN(n19290) );
  XOR2_X1 U19987 ( .A1(n10130), .A2(n13517), .Z(n10129) );
  INV_X2 U19992 ( .I(n657), .ZN(n23868) );
  NOR2_X1 U19993 ( .A1(n29246), .A2(n10145), .ZN(n10542) );
  XOR2_X1 U19995 ( .A1(n23521), .A2(n12122), .Z(n10150) );
  XOR2_X1 U19999 ( .A1(n22198), .A2(n25054), .Z(n10155) );
  OAI21_X2 U20000 ( .A1(n21607), .A2(n21776), .B(n18163), .ZN(n22198) );
  XOR2_X1 U20002 ( .A1(n10157), .A2(n25735), .Z(Ciphertext[158]) );
  XOR2_X1 U20004 ( .A1(n20819), .A2(n10159), .Z(n15338) );
  XOR2_X1 U20008 ( .A1(n27180), .A2(n25570), .Z(n10165) );
  INV_X2 U20009 ( .I(n10171), .ZN(n25628) );
  XOR2_X1 U20012 ( .A1(n22157), .A2(n16237), .Z(n10370) );
  NAND3_X1 U20013 ( .A1(n11931), .A2(n27262), .A3(n10174), .ZN(n10268) );
  XOR2_X1 U20017 ( .A1(n19341), .A2(n25009), .Z(n10180) );
  NOR2_X1 U20018 ( .A1(n10182), .A2(n10181), .ZN(n18590) );
  XOR2_X1 U20021 ( .A1(n21924), .A2(n21577), .Z(n10184) );
  XOR2_X1 U20027 ( .A1(n24428), .A2(n10195), .Z(n10194) );
  NAND2_X2 U20029 ( .A1(n17118), .A2(n24610), .ZN(n10199) );
  XOR2_X1 U20031 ( .A1(n9706), .A2(n24895), .Z(n20712) );
  XOR2_X1 U20032 ( .A1(n10201), .A2(n16657), .Z(n14656) );
  AND2_X1 U20033 ( .A1(n629), .A2(n10206), .Z(n10908) );
  AOI21_X2 U20034 ( .A1(n10208), .A2(n18403), .B(n10207), .ZN(n16354) );
  INV_X2 U20035 ( .I(n10209), .ZN(n18219) );
  OAI21_X1 U20036 ( .A1(n4289), .A2(n816), .B(n20570), .ZN(n20573) );
  XOR2_X1 U20041 ( .A1(n29320), .A2(n11603), .Z(n10237) );
  XOR2_X1 U20042 ( .A1(n29320), .A2(n25728), .Z(n24443) );
  XOR2_X1 U20043 ( .A1(n29320), .A2(n24507), .Z(n24508) );
  AOI21_X1 U20044 ( .A1(n824), .A2(n10227), .B(n13568), .ZN(n17981) );
  XOR2_X1 U20052 ( .A1(n10087), .A2(n13075), .Z(n10249) );
  NOR2_X1 U20053 ( .A1(n974), .A2(n10281), .ZN(n24131) );
  NAND2_X1 U20054 ( .A1(n2575), .A2(n10254), .ZN(n14870) );
  XOR2_X1 U20058 ( .A1(n19710), .A2(n25086), .Z(n10262) );
  NAND3_X1 U20059 ( .A1(n29659), .A2(n28010), .A3(n15519), .ZN(n18438) );
  OAI22_X1 U20060 ( .A1(n10843), .A2(n29659), .B1(n17321), .B2(n959), .ZN(
        n10842) );
  XOR2_X1 U20062 ( .A1(n22079), .A2(n10270), .Z(n22082) );
  XOR2_X1 U20063 ( .A1(n32881), .A2(n2353), .Z(n10270) );
  XOR2_X1 U20068 ( .A1(n24624), .A2(n11699), .Z(n10276) );
  XOR2_X1 U20069 ( .A1(n22014), .A2(n1392), .Z(n10278) );
  XNOR2_X1 U20071 ( .A1(Plaintext[180]), .A2(Key[180]), .ZN(n10284) );
  INV_X2 U20072 ( .I(n10287), .ZN(n10533) );
  NAND2_X1 U20077 ( .A1(n12487), .A2(n10301), .ZN(n12486) );
  OAI22_X1 U20078 ( .A1(n16836), .A2(n14954), .B1(n28658), .B2(n10301), .ZN(
        n12302) );
  NOR2_X1 U20079 ( .A1(n1322), .A2(n21832), .ZN(n21835) );
  XOR2_X1 U20080 ( .A1(n12828), .A2(n10304), .Z(n16332) );
  XOR2_X1 U20081 ( .A1(n22300), .A2(n12084), .Z(n10304) );
  XOR2_X1 U20082 ( .A1(n23368), .A2(n10308), .Z(n23127) );
  MUX2_X1 U20083 ( .I0(n20360), .I1(n27600), .S(n29553), .Z(n20240) );
  XOR2_X1 U20088 ( .A1(n572), .A2(n14916), .Z(n10320) );
  NOR2_X1 U20092 ( .A1(n30558), .A2(n10325), .ZN(n18885) );
  XOR2_X1 U20094 ( .A1(n8356), .A2(n24964), .Z(n10328) );
  XOR2_X1 U20096 ( .A1(n27801), .A2(n27950), .Z(n24445) );
  XOR2_X1 U20101 ( .A1(n9145), .A2(n14727), .Z(n15588) );
  XOR2_X1 U20103 ( .A1(n15293), .A2(n15408), .Z(n10347) );
  INV_X2 U20104 ( .I(n10350), .ZN(n15318) );
  OR2_X1 U20105 ( .A1(n12691), .A2(n11608), .Z(n10358) );
  XOR2_X1 U20118 ( .A1(n30571), .A2(n16634), .Z(n21457) );
  XOR2_X1 U20119 ( .A1(n156), .A2(n1194), .Z(n10399) );
  XOR2_X1 U20121 ( .A1(n33219), .A2(n25213), .Z(n10412) );
  AND2_X1 U20123 ( .A1(n11346), .A2(n1775), .Z(n10416) );
  XOR2_X1 U20127 ( .A1(n22284), .A2(n22283), .Z(n10421) );
  INV_X2 U20129 ( .I(n10426), .ZN(n19724) );
  INV_X2 U20130 ( .I(n10430), .ZN(n11900) );
  XOR2_X1 U20132 ( .A1(n25993), .A2(n1431), .Z(n10434) );
  NAND2_X1 U20134 ( .A1(n17368), .A2(n14213), .ZN(n10485) );
  NAND2_X1 U20135 ( .A1(n12877), .A2(n14213), .ZN(n12533) );
  OAI21_X1 U20136 ( .A1(n16443), .A2(n26158), .B(n10449), .ZN(n10448) );
  XOR2_X1 U20139 ( .A1(n848), .A2(n29155), .Z(n10459) );
  XOR2_X1 U20141 ( .A1(n11762), .A2(n22083), .Z(n10461) );
  XOR2_X1 U20147 ( .A1(n19731), .A2(n10467), .Z(n10466) );
  XOR2_X1 U20148 ( .A1(n19375), .A2(n1369), .Z(n10467) );
  NOR2_X1 U20150 ( .A1(n5455), .A2(n7492), .ZN(n12144) );
  XOR2_X1 U20153 ( .A1(n12414), .A2(n1198), .Z(n10474) );
  NOR2_X2 U20157 ( .A1(n10491), .A2(n10490), .ZN(n22130) );
  INV_X2 U20161 ( .I(n10505), .ZN(n21398) );
  XOR2_X1 U20163 ( .A1(n20893), .A2(n10508), .Z(n10507) );
  XOR2_X1 U20164 ( .A1(n20970), .A2(n1338), .Z(n10508) );
  INV_X2 U20165 ( .I(n10514), .ZN(n19991) );
  XOR2_X1 U20167 ( .A1(n24429), .A2(n15473), .Z(n10515) );
  XOR2_X1 U20168 ( .A1(n30795), .A2(n7879), .Z(n24429) );
  XOR2_X1 U20169 ( .A1(n10585), .A2(n15815), .Z(n10516) );
  XOR2_X1 U20173 ( .A1(n10525), .A2(n22712), .Z(n15116) );
  NOR2_X1 U20177 ( .A1(n71), .A2(n20103), .ZN(n16980) );
  NAND2_X1 U20178 ( .A1(n15551), .A2(n71), .ZN(n20105) );
  XOR2_X1 U20179 ( .A1(n10539), .A2(n13419), .Z(n24529) );
  XOR2_X1 U20180 ( .A1(n24635), .A2(n10539), .Z(n16394) );
  OAI21_X2 U20182 ( .A1(n10548), .A2(n10756), .B(n10547), .ZN(n10755) );
  XOR2_X1 U20185 ( .A1(n29312), .A2(n10553), .Z(n10552) );
  INV_X2 U20189 ( .I(n16881), .ZN(n16948) );
  NAND2_X2 U20190 ( .A1(n11247), .A2(n10566), .ZN(n24970) );
  NAND2_X1 U20191 ( .A1(n18035), .A2(n12323), .ZN(n10571) );
  NAND2_X1 U20193 ( .A1(n20580), .A2(n26566), .ZN(n20584) );
  XOR2_X1 U20195 ( .A1(n32399), .A2(n16685), .Z(n10581) );
  XOR2_X1 U20197 ( .A1(n2864), .A2(n10584), .Z(n10583) );
  XOR2_X1 U20198 ( .A1(n10587), .A2(n16533), .Z(Ciphertext[69]) );
  AND2_X1 U20200 ( .A1(n30234), .A2(n8365), .Z(n10589) );
  NOR2_X1 U20205 ( .A1(n24590), .A2(n30018), .ZN(n10600) );
  INV_X1 U20206 ( .I(n24590), .ZN(n10603) );
  NOR2_X1 U20207 ( .A1(n10606), .A2(n10605), .ZN(n10604) );
  XOR2_X1 U20213 ( .A1(n22056), .A2(n17679), .Z(n22268) );
  XOR2_X1 U20215 ( .A1(n11694), .A2(n1309), .Z(n11884) );
  XOR2_X1 U20216 ( .A1(n31105), .A2(n9960), .Z(n21879) );
  XOR2_X1 U20217 ( .A1(n7828), .A2(n15775), .Z(n10616) );
  XOR2_X1 U20220 ( .A1(n10626), .A2(n13956), .Z(n11600) );
  XOR2_X1 U20225 ( .A1(n16076), .A2(n10773), .Z(n17915) );
  XOR2_X1 U20227 ( .A1(n9536), .A2(n10650), .Z(n10649) );
  NOR2_X1 U20229 ( .A1(n13509), .A2(n7007), .ZN(n10658) );
  NAND2_X1 U20231 ( .A1(n21424), .A2(n6855), .ZN(n15564) );
  NOR2_X1 U20232 ( .A1(n30854), .A2(n21424), .ZN(n21337) );
  OAI21_X1 U20233 ( .A1(n21243), .A2(n30854), .B(n11912), .ZN(n17803) );
  MUX2_X1 U20234 ( .I0(n20071), .I1(n31080), .S(n729), .Z(n20072) );
  XOR2_X1 U20235 ( .A1(n19666), .A2(n10662), .Z(n10661) );
  XOR2_X1 U20236 ( .A1(n29312), .A2(n1193), .Z(n10662) );
  NAND2_X1 U20239 ( .A1(n18747), .A2(n10665), .ZN(n17874) );
  NAND2_X1 U20240 ( .A1(n16487), .A2(n10665), .ZN(n14706) );
  NOR2_X1 U20241 ( .A1(n12575), .A2(n12574), .ZN(n10666) );
  XOR2_X1 U20244 ( .A1(n22211), .A2(n22226), .Z(n22242) );
  XNOR2_X1 U20245 ( .A1(n10675), .A2(n10674), .ZN(n10673) );
  XOR2_X1 U20263 ( .A1(n10704), .A2(n10701), .Z(n10725) );
  XOR2_X1 U20264 ( .A1(n10703), .A2(n10702), .Z(n10701) );
  XOR2_X1 U20265 ( .A1(n17362), .A2(n25038), .Z(n10702) );
  OAI21_X2 U20272 ( .A1(n6303), .A2(n14955), .B(n10721), .ZN(n12561) );
  XOR2_X1 U20273 ( .A1(n17213), .A2(n15708), .Z(n10722) );
  XOR2_X1 U20274 ( .A1(n19586), .A2(n461), .Z(n10723) );
  XOR2_X1 U20275 ( .A1(n10727), .A2(n17205), .Z(n17203) );
  XOR2_X1 U20276 ( .A1(n10728), .A2(n34160), .Z(n10727) );
  XOR2_X1 U20277 ( .A1(n17697), .A2(n1429), .Z(n10728) );
  XOR2_X1 U20284 ( .A1(n20857), .A2(n20905), .Z(n10737) );
  XOR2_X1 U20285 ( .A1(n19626), .A2(n19708), .Z(n10738) );
  NOR2_X1 U20288 ( .A1(n17110), .A2(n25292), .ZN(n10744) );
  NOR2_X1 U20289 ( .A1(n10748), .A2(n17110), .ZN(n10747) );
  AOI22_X2 U20291 ( .A1(n10763), .A2(n23850), .B1(n14664), .B2(n10762), .ZN(
        n24299) );
  XOR2_X1 U20302 ( .A1(n2353), .A2(n22248), .Z(n17219) );
  NOR2_X2 U20303 ( .A1(n11493), .A2(n19953), .ZN(n11984) );
  XOR2_X1 U20307 ( .A1(n10800), .A2(n10797), .Z(n17144) );
  XOR2_X1 U20308 ( .A1(n10799), .A2(n10798), .Z(n10797) );
  XOR2_X1 U20309 ( .A1(n20848), .A2(n16679), .Z(n10798) );
  XOR2_X1 U20313 ( .A1(n10810), .A2(n19591), .Z(n10809) );
  XOR2_X1 U20315 ( .A1(n28848), .A2(n25191), .Z(n10814) );
  AND2_X1 U20316 ( .A1(n25066), .A2(n10822), .Z(n10821) );
  NOR2_X1 U20322 ( .A1(n13304), .A2(n18048), .ZN(n21387) );
  XOR2_X1 U20335 ( .A1(n19763), .A2(n17091), .Z(n10866) );
  XOR2_X1 U20337 ( .A1(n10873), .A2(n14979), .Z(n10872) );
  XOR2_X1 U20341 ( .A1(n20916), .A2(n10878), .Z(n10877) );
  XOR2_X1 U20344 ( .A1(n2353), .A2(n24953), .Z(n10887) );
  XOR2_X1 U20345 ( .A1(n10889), .A2(n18190), .Z(n10888) );
  XOR2_X1 U20346 ( .A1(n30212), .A2(n25801), .Z(n19340) );
  NAND3_X1 U20347 ( .A1(n20569), .A2(n29069), .A3(n4289), .ZN(n11761) );
  INV_X2 U20351 ( .I(n10900), .ZN(n16442) );
  NAND2_X2 U20353 ( .A1(n10910), .A2(n10909), .ZN(n19199) );
  XOR2_X1 U20354 ( .A1(n10915), .A2(n15029), .Z(n10914) );
  XOR2_X1 U20356 ( .A1(n15031), .A2(n4400), .Z(n10917) );
  INV_X1 U20357 ( .I(n24004), .ZN(n13984) );
  NAND2_X1 U20358 ( .A1(n31096), .A2(n24004), .ZN(n14889) );
  INV_X2 U20361 ( .I(n10932), .ZN(n16633) );
  INV_X2 U20362 ( .I(n10936), .ZN(n16534) );
  XOR2_X1 U20364 ( .A1(n10945), .A2(n10944), .Z(n25308) );
  XOR2_X1 U20366 ( .A1(n10946), .A2(n24895), .Z(n12779) );
  XOR2_X1 U20367 ( .A1(n10946), .A2(n22056), .Z(n21948) );
  OAI22_X2 U20369 ( .A1(n17581), .A2(n3219), .B1(n15086), .B2(n15085), .ZN(
        n24636) );
  MUX2_X1 U20373 ( .I0(n802), .I1(n22766), .S(n9293), .Z(n22767) );
  XOR2_X1 U20379 ( .A1(n12614), .A2(n10961), .Z(n10960) );
  XOR2_X1 U20380 ( .A1(n14952), .A2(n960), .Z(n10961) );
  XOR2_X1 U20385 ( .A1(n10979), .A2(n24943), .Z(n21661) );
  XOR2_X1 U20386 ( .A1(n22303), .A2(n10979), .Z(n22155) );
  XOR2_X1 U20391 ( .A1(n19517), .A2(n10986), .Z(n10985) );
  NAND2_X1 U20392 ( .A1(n26830), .A2(n19229), .ZN(n15845) );
  XOR2_X1 U20395 ( .A1(n22244), .A2(n10990), .Z(n10989) );
  XOR2_X1 U20396 ( .A1(n22291), .A2(n10991), .Z(n10990) );
  INV_X1 U20397 ( .I(n24968), .ZN(n10991) );
  NAND2_X2 U20398 ( .A1(n16364), .A2(n19810), .ZN(n20429) );
  XOR2_X1 U20400 ( .A1(n23526), .A2(n23525), .Z(n23931) );
  INV_X2 U20409 ( .I(n11006), .ZN(n12657) );
  XOR2_X1 U20410 ( .A1(n27138), .A2(n32918), .Z(n19700) );
  XOR2_X1 U20411 ( .A1(n32889), .A2(n21016), .Z(n11012) );
  XOR2_X1 U20417 ( .A1(n22085), .A2(n11028), .Z(n11027) );
  INV_X1 U20418 ( .I(n16636), .ZN(n11028) );
  XOR2_X1 U20422 ( .A1(n400), .A2(n25036), .Z(n19638) );
  NAND2_X1 U20425 ( .A1(n16291), .A2(n25276), .ZN(n25280) );
  XOR2_X1 U20427 ( .A1(n10870), .A2(n16438), .Z(n15775) );
  NAND3_X1 U20431 ( .A1(n32941), .A2(n13499), .A3(n33721), .ZN(n20051) );
  XOR2_X1 U20433 ( .A1(n20985), .A2(n12957), .Z(n20896) );
  XOR2_X1 U20434 ( .A1(n7256), .A2(n16685), .Z(n24628) );
  NOR2_X1 U20441 ( .A1(n23578), .A2(n12287), .ZN(n11095) );
  NAND3_X1 U20442 ( .A1(n14232), .A2(n23958), .A3(n11096), .ZN(n23959) );
  MUX2_X1 U20443 ( .I0(n21252), .I1(n17437), .S(n1337), .Z(n21254) );
  AOI22_X1 U20444 ( .A1(n16017), .A2(n30283), .B1(n14677), .B2(n11107), .ZN(
        n24036) );
  XOR2_X1 U20449 ( .A1(n20982), .A2(n25648), .Z(n11118) );
  XOR2_X1 U20451 ( .A1(n11128), .A2(n15460), .Z(n11124) );
  XOR2_X1 U20453 ( .A1(n22128), .A2(n2353), .Z(n11126) );
  XOR2_X1 U20455 ( .A1(n11130), .A2(n11129), .Z(n13080) );
  XOR2_X1 U20456 ( .A1(n19441), .A2(n19442), .Z(n11129) );
  XOR2_X1 U20457 ( .A1(n13829), .A2(n12453), .Z(n11130) );
  INV_X1 U20460 ( .I(n17110), .ZN(n14509) );
  NOR2_X1 U20461 ( .A1(n34109), .A2(n25247), .ZN(n11136) );
  NOR2_X1 U20466 ( .A1(n14376), .A2(n11147), .ZN(n11146) );
  XOR2_X1 U20467 ( .A1(n23190), .A2(n12123), .Z(n11148) );
  XOR2_X1 U20468 ( .A1(n23363), .A2(n23189), .Z(n23276) );
  NAND2_X1 U20470 ( .A1(n17661), .A2(n23806), .ZN(n11159) );
  XOR2_X1 U20472 ( .A1(n25969), .A2(n25908), .Z(n20482) );
  INV_X1 U20474 ( .I(n21811), .ZN(n14917) );
  AOI21_X2 U20475 ( .A1(n21809), .A2(n2801), .B(n11167), .ZN(n11166) );
  XOR2_X1 U20476 ( .A1(n24638), .A2(n25252), .Z(n11170) );
  XOR2_X1 U20477 ( .A1(n24455), .A2(n24600), .Z(n11171) );
  INV_X2 U20480 ( .I(n11175), .ZN(n22640) );
  XOR2_X1 U20484 ( .A1(n23393), .A2(n26701), .Z(n11194) );
  XOR2_X1 U20491 ( .A1(n11206), .A2(n21886), .Z(n21997) );
  AND3_X1 U20497 ( .A1(n26026), .A2(n17828), .A3(n23104), .Z(n17585) );
  XOR2_X1 U20498 ( .A1(n11225), .A2(n11223), .Z(n12906) );
  XOR2_X1 U20503 ( .A1(n23453), .A2(n1402), .Z(n11227) );
  INV_X1 U20511 ( .I(n25285), .ZN(n25279) );
  NAND2_X1 U20512 ( .A1(n18483), .A2(n9549), .ZN(n15165) );
  INV_X2 U20513 ( .I(n24565), .ZN(n25295) );
  INV_X2 U20520 ( .I(n11281), .ZN(n11916) );
  XOR2_X1 U20523 ( .A1(n23532), .A2(n25735), .Z(n16263) );
  NOR2_X1 U20526 ( .A1(n11734), .A2(n11966), .ZN(n11285) );
  XOR2_X1 U20527 ( .A1(n11290), .A2(n14481), .Z(n11289) );
  XOR2_X1 U20532 ( .A1(n11297), .A2(n29707), .Z(n14079) );
  XOR2_X1 U20534 ( .A1(n11297), .A2(n31687), .Z(n24423) );
  XOR2_X1 U20535 ( .A1(n11297), .A2(n16671), .Z(n24048) );
  NAND2_X1 U20536 ( .A1(n11302), .A2(n743), .ZN(n19219) );
  XOR2_X1 U20542 ( .A1(Plaintext[156]), .A2(Key[156]), .Z(n14159) );
  OR2_X1 U20543 ( .A1(n18543), .A2(n18858), .Z(n11318) );
  XOR2_X1 U20548 ( .A1(n24642), .A2(n24861), .Z(n24517) );
  INV_X2 U20549 ( .I(n15401), .ZN(n23755) );
  XOR2_X1 U20550 ( .A1(n22616), .A2(n11326), .Z(n13132) );
  NAND3_X2 U20551 ( .A1(n21757), .A2(n11719), .A3(n15410), .ZN(n22096) );
  XOR2_X1 U20552 ( .A1(n20989), .A2(n11339), .Z(n11338) );
  XOR2_X1 U20553 ( .A1(n20904), .A2(n16672), .Z(n11339) );
  INV_X2 U20555 ( .I(n11348), .ZN(n14290) );
  XOR2_X1 U20556 ( .A1(n11353), .A2(n11351), .Z(n11910) );
  XOR2_X1 U20558 ( .A1(n11354), .A2(n19707), .Z(n11353) );
  XOR2_X1 U20560 ( .A1(n11357), .A2(n11356), .Z(n11355) );
  XOR2_X1 U20561 ( .A1(n22189), .A2(n30954), .Z(n11356) );
  XOR2_X1 U20562 ( .A1(n2896), .A2(n4342), .Z(n11357) );
  NOR2_X1 U20566 ( .A1(n25082), .A2(n11360), .ZN(n25094) );
  XOR2_X1 U20568 ( .A1(n19494), .A2(n25288), .Z(n11361) );
  NAND3_X1 U20569 ( .A1(n15434), .A2(n15005), .A3(n14545), .ZN(n13933) );
  INV_X2 U20570 ( .I(n11364), .ZN(n16317) );
  XOR2_X1 U20574 ( .A1(n11722), .A2(n25720), .Z(n24639) );
  XOR2_X1 U20580 ( .A1(Plaintext[26]), .A2(Key[26]), .Z(n11599) );
  XNOR2_X1 U20581 ( .A1(Plaintext[103]), .A2(Key[103]), .ZN(n11379) );
  NOR2_X1 U20583 ( .A1(n27188), .A2(n18151), .ZN(n12235) );
  NAND2_X1 U20585 ( .A1(n962), .A2(n11390), .ZN(n14543) );
  XOR2_X1 U20588 ( .A1(n11568), .A2(n22728), .Z(n23745) );
  NOR2_X2 U20589 ( .A1(n6783), .A2(n12290), .ZN(n12238) );
  OAI21_X2 U20595 ( .A1(n24485), .A2(n29629), .B(n11429), .ZN(n24960) );
  XOR2_X1 U20596 ( .A1(n19564), .A2(n11433), .Z(n11432) );
  XOR2_X1 U20597 ( .A1(n15117), .A2(n25324), .Z(n11433) );
  NOR2_X1 U20601 ( .A1(n16627), .A2(n22435), .ZN(n11443) );
  XOR2_X1 U20602 ( .A1(n14214), .A2(n17551), .Z(n11450) );
  XNOR2_X1 U20603 ( .A1(n19408), .A2(n19398), .ZN(n18072) );
  INV_X2 U20604 ( .I(n11451), .ZN(n16627) );
  XOR2_X1 U20608 ( .A1(n26562), .A2(n20389), .Z(n18113) );
  NAND2_X1 U20609 ( .A1(n10181), .A2(n11459), .ZN(n14695) );
  XOR2_X1 U20611 ( .A1(Plaintext[177]), .A2(Key[177]), .Z(n18873) );
  NOR2_X1 U20613 ( .A1(n10673), .A2(n499), .ZN(n23633) );
  OAI21_X1 U20614 ( .A1(n17947), .A2(n4254), .B(n20486), .ZN(n11465) );
  INV_X1 U20615 ( .I(n11468), .ZN(n25153) );
  OAI22_X1 U20616 ( .A1(n25166), .A2(n25174), .B1(n25179), .B2(n11468), .ZN(
        n12457) );
  OAI21_X2 U20617 ( .A1(n14971), .A2(n33904), .B(n24463), .ZN(n24956) );
  XOR2_X1 U20618 ( .A1(n30628), .A2(n1196), .Z(n11476) );
  XOR2_X1 U20620 ( .A1(n11485), .A2(n11484), .Z(n11483) );
  XOR2_X1 U20622 ( .A1(n16693), .A2(n705), .Z(n11485) );
  INV_X1 U20624 ( .I(n21258), .ZN(n21255) );
  XOR2_X1 U20626 ( .A1(n19541), .A2(n17072), .Z(n11488) );
  XOR2_X1 U20630 ( .A1(n1045), .A2(n13826), .Z(n17213) );
  XOR2_X1 U20632 ( .A1(n11504), .A2(n25506), .Z(n23167) );
  NAND2_X2 U20635 ( .A1(n19040), .A2(n19042), .ZN(n13925) );
  XOR2_X1 U20638 ( .A1(n19495), .A2(n11523), .Z(n11522) );
  XOR2_X1 U20639 ( .A1(n30193), .A2(n1419), .Z(n11523) );
  XOR2_X1 U20640 ( .A1(n17552), .A2(n15983), .Z(n11524) );
  XOR2_X1 U20641 ( .A1(n13810), .A2(n11526), .Z(n11525) );
  XOR2_X1 U20642 ( .A1(n24675), .A2(n7603), .Z(n11526) );
  XOR2_X1 U20643 ( .A1(n11529), .A2(n11528), .Z(n22486) );
  XOR2_X1 U20645 ( .A1(n16457), .A2(n17174), .Z(n11529) );
  XOR2_X1 U20646 ( .A1(n11532), .A2(n11531), .Z(n11530) );
  XOR2_X1 U20647 ( .A1(n13970), .A2(n13331), .Z(n11531) );
  XOR2_X1 U20651 ( .A1(n16513), .A2(n11544), .Z(n11543) );
  XOR2_X1 U20652 ( .A1(n16349), .A2(n19649), .Z(n11544) );
  NOR2_X1 U20655 ( .A1(n25391), .A2(n32884), .ZN(n25392) );
  XOR2_X1 U20657 ( .A1(n11558), .A2(n16649), .Z(Ciphertext[91]) );
  XOR2_X1 U20659 ( .A1(n22032), .A2(n16703), .Z(n11819) );
  NOR2_X1 U20662 ( .A1(n11567), .A2(n30089), .ZN(n23597) );
  XOR2_X1 U20664 ( .A1(n9434), .A2(n30943), .Z(n11574) );
  XOR2_X1 U20665 ( .A1(n11578), .A2(n516), .Z(n11577) );
  XOR2_X1 U20668 ( .A1(n18401), .A2(Key[172]), .Z(n18847) );
  AND2_X1 U20673 ( .A1(n11601), .A2(n21070), .Z(n12933) );
  INV_X1 U20676 ( .I(n16674), .ZN(n11603) );
  XOR2_X1 U20677 ( .A1(n19772), .A2(n11604), .Z(n19775) );
  XOR2_X1 U20678 ( .A1(n22790), .A2(n11611), .Z(n11610) );
  XOR2_X1 U20679 ( .A1(n10773), .A2(n1393), .Z(n11611) );
  XOR2_X1 U20680 ( .A1(n23318), .A2(n23273), .Z(n22790) );
  XOR2_X1 U20681 ( .A1(n23173), .A2(n23460), .Z(n11612) );
  NOR2_X1 U20682 ( .A1(n13175), .A2(n24110), .ZN(n11613) );
  INV_X2 U20684 ( .I(n11620), .ZN(n22476) );
  XNOR2_X1 U20686 ( .A1(n471), .A2(n11631), .ZN(n11630) );
  XOR2_X1 U20687 ( .A1(n17840), .A2(n19536), .Z(n11631) );
  XOR2_X1 U20689 ( .A1(Plaintext[74]), .A2(Key[74]), .Z(n11773) );
  XOR2_X1 U20692 ( .A1(n33453), .A2(n15816), .Z(n17095) );
  XOR2_X1 U20693 ( .A1(n33453), .A2(n23191), .Z(n14967) );
  NAND2_X1 U20698 ( .A1(n24250), .A2(n28553), .ZN(n17409) );
  XOR2_X1 U20702 ( .A1(n19780), .A2(n24964), .Z(n11661) );
  XOR2_X1 U20705 ( .A1(n1369), .A2(n876), .Z(n11663) );
  NAND2_X2 U20709 ( .A1(n11675), .A2(n12187), .ZN(n24393) );
  XOR2_X1 U20710 ( .A1(n18356), .A2(Key[18]), .Z(n18654) );
  NOR2_X1 U20712 ( .A1(n1334), .A2(n11814), .ZN(n11680) );
  XOR2_X1 U20713 ( .A1(n24676), .A2(n16533), .Z(n11681) );
  NAND2_X2 U20714 ( .A1(n11686), .A2(n11682), .ZN(n15296) );
  XOR2_X1 U20715 ( .A1(n11689), .A2(n11690), .Z(n16784) );
  XOR2_X1 U20716 ( .A1(n20894), .A2(n15652), .Z(n11690) );
  XOR2_X1 U20719 ( .A1(n24652), .A2(n15779), .Z(n11699) );
  XOR2_X1 U20726 ( .A1(n5932), .A2(n25990), .Z(n14363) );
  XOR2_X1 U20727 ( .A1(n31508), .A2(n25991), .Z(n24651) );
  XOR2_X1 U20733 ( .A1(n22063), .A2(n16479), .Z(n11750) );
  INV_X1 U20736 ( .I(n23263), .ZN(n11766) );
  XOR2_X1 U20739 ( .A1(n17091), .A2(n33918), .Z(n19481) );
  XNOR2_X1 U20740 ( .A1(n17091), .A2(n19337), .ZN(n15157) );
  INV_X2 U20741 ( .I(n11773), .ZN(n18559) );
  XOR2_X1 U20743 ( .A1(n14656), .A2(n11776), .Z(n11775) );
  XOR2_X1 U20744 ( .A1(n24836), .A2(n14533), .Z(n11782) );
  XOR2_X1 U20745 ( .A1(n32310), .A2(n27920), .Z(n11783) );
  XOR2_X1 U20747 ( .A1(n17301), .A2(n16507), .Z(n11803) );
  XOR2_X1 U20749 ( .A1(n27252), .A2(n15415), .Z(n13739) );
  XOR2_X1 U20751 ( .A1(n20954), .A2(n20955), .Z(n14854) );
  XOR2_X1 U20752 ( .A1(n19445), .A2(n33587), .Z(n11817) );
  XOR2_X1 U20756 ( .A1(n11841), .A2(n11843), .Z(n11844) );
  XOR2_X1 U20757 ( .A1(n11842), .A2(n24637), .Z(n11841) );
  INV_X2 U20759 ( .I(n11844), .ZN(n12042) );
  XNOR2_X1 U20761 ( .A1(n15047), .A2(n15048), .ZN(n11847) );
  NAND3_X2 U20763 ( .A1(n11854), .A2(n22458), .A3(n11853), .ZN(n23086) );
  NAND2_X1 U20764 ( .A1(n17670), .A2(n11855), .ZN(n19547) );
  NAND2_X1 U20767 ( .A1(n15797), .A2(n15796), .ZN(n11860) );
  NAND3_X2 U20768 ( .A1(n17101), .A2(n16048), .A3(n20373), .ZN(n12424) );
  XOR2_X1 U20772 ( .A1(n11869), .A2(n14401), .Z(n14400) );
  XOR2_X1 U20773 ( .A1(n24805), .A2(n5268), .Z(n24668) );
  OAI21_X1 U20777 ( .A1(n694), .A2(n25322), .B(n16041), .ZN(n15854) );
  NAND3_X1 U20778 ( .A1(n32867), .A2(n16041), .A3(n694), .ZN(n25309) );
  INV_X2 U20779 ( .I(n11877), .ZN(n18035) );
  XOR2_X1 U20781 ( .A1(n18348), .A2(Key[37]), .Z(n18548) );
  INV_X1 U20787 ( .I(n33848), .ZN(n20034) );
  NAND4_X1 U20788 ( .A1(n11214), .A2(n12642), .A3(n12640), .A4(n12641), .ZN(
        n21546) );
  NOR2_X1 U20789 ( .A1(n20944), .A2(n21181), .ZN(n15321) );
  AOI22_X1 U20790 ( .A1(n24780), .A2(n24874), .B1(n10770), .B2(n15719), .ZN(
        n15234) );
  NOR2_X1 U20792 ( .A1(n1205), .A2(n24998), .ZN(n14837) );
  NAND3_X1 U20793 ( .A1(n1291), .A2(n29336), .A3(n855), .ZN(n14772) );
  NAND2_X1 U20794 ( .A1(n13962), .A2(n31161), .ZN(n15135) );
  INV_X1 U20797 ( .I(n12257), .ZN(n15062) );
  NAND2_X1 U20798 ( .A1(n18437), .A2(n958), .ZN(n16207) );
  NOR2_X1 U20799 ( .A1(n18007), .A2(n18427), .ZN(n18428) );
  INV_X1 U20802 ( .I(n19412), .ZN(n19592) );
  NOR2_X1 U20804 ( .A1(n12244), .A2(n20338), .ZN(n12843) );
  INV_X1 U20805 ( .I(n20574), .ZN(n12812) );
  INV_X1 U20818 ( .I(n18623), .ZN(n18771) );
  INV_X1 U20821 ( .I(n18423), .ZN(n17102) );
  NAND2_X1 U20824 ( .A1(n14828), .A2(n13738), .ZN(n17231) );
  INV_X1 U20834 ( .I(n20842), .ZN(n17759) );
  NAND4_X1 U20839 ( .A1(n13285), .A2(n13284), .A3(n19892), .A4(n13283), .ZN(
        n13282) );
  INV_X1 U20844 ( .I(n17672), .ZN(n20266) );
  INV_X1 U20847 ( .I(n20351), .ZN(n12367) );
  NAND2_X1 U20850 ( .A1(n14156), .A2(n9437), .ZN(n13788) );
  NOR2_X1 U20852 ( .A1(n962), .A2(n14926), .ZN(n12291) );
  NAND2_X1 U20854 ( .A1(n16226), .A2(n29256), .ZN(n14174) );
  NAND2_X1 U20855 ( .A1(n21365), .A2(n20945), .ZN(n20705) );
  NAND2_X1 U20858 ( .A1(n19258), .A2(n19257), .ZN(n19259) );
  NAND2_X1 U20865 ( .A1(n957), .A2(n12956), .ZN(n18519) );
  NAND2_X1 U20874 ( .A1(n18439), .A2(n19355), .ZN(n17996) );
  NOR2_X1 U20875 ( .A1(n13390), .A2(n28386), .ZN(n18439) );
  NAND2_X1 U20878 ( .A1(n18825), .A2(n17553), .ZN(n14859) );
  NAND3_X1 U20880 ( .A1(n15417), .A2(n1048), .A3(n15780), .ZN(n18452) );
  NAND2_X1 U20881 ( .A1(n19271), .A2(n19265), .ZN(n15780) );
  INV_X1 U20882 ( .I(n21379), .ZN(n21178) );
  OAI21_X1 U20883 ( .A1(n16905), .A2(n13319), .B(n13581), .ZN(n13580) );
  NAND3_X1 U20885 ( .A1(n14384), .A2(n8029), .A3(n31042), .ZN(n21519) );
  OAI21_X1 U20886 ( .A1(n17078), .A2(n14640), .B(n15171), .ZN(n21521) );
  NOR2_X1 U20889 ( .A1(n14008), .A2(n15752), .ZN(n15635) );
  NAND2_X1 U20892 ( .A1(n22478), .A2(n22377), .ZN(n13186) );
  NAND2_X1 U20898 ( .A1(n16493), .A2(n16105), .ZN(n16262) );
  INV_X1 U20899 ( .I(n19368), .ZN(n17104) );
  NOR2_X1 U20902 ( .A1(n13561), .A2(n14253), .ZN(n13587) );
  AOI21_X1 U20907 ( .A1(n23778), .A2(n8547), .B(n23776), .ZN(n13140) );
  NAND2_X1 U20908 ( .A1(n28367), .A2(n23871), .ZN(n23876) );
  INV_X1 U20917 ( .I(n12720), .ZN(n13825) );
  INV_X1 U20918 ( .I(n24356), .ZN(n24493) );
  NAND2_X1 U20919 ( .A1(n17047), .A2(n17037), .ZN(n17046) );
  INV_X1 U20922 ( .I(n20454), .ZN(n14086) );
  NAND2_X1 U20925 ( .A1(n868), .A2(n20525), .ZN(n20276) );
  INV_X1 U20927 ( .I(n20350), .ZN(n12366) );
  INV_X1 U20931 ( .I(n25856), .ZN(n14557) );
  INV_X1 U20934 ( .I(n18882), .ZN(n17478) );
  INV_X1 U20936 ( .I(n18695), .ZN(n18697) );
  NOR2_X1 U20937 ( .A1(n30271), .A2(n12006), .ZN(n15141) );
  AOI22_X1 U20938 ( .A1(n14271), .A2(n15589), .B1(n7690), .B2(n3931), .ZN(
        n14270) );
  NOR2_X1 U20939 ( .A1(n15261), .A2(n14721), .ZN(n14271) );
  NAND2_X1 U20943 ( .A1(n15874), .A2(n21398), .ZN(n16258) );
  INV_X1 U20946 ( .I(n17822), .ZN(n14305) );
  NAND2_X1 U20947 ( .A1(n14290), .A2(n1335), .ZN(n15160) );
  NOR2_X1 U20950 ( .A1(n21073), .A2(n29255), .ZN(n16844) );
  INV_X1 U20951 ( .I(n16545), .ZN(n16544) );
  INV_X1 U20958 ( .I(n21362), .ZN(n14903) );
  AOI21_X1 U20963 ( .A1(n16403), .A2(n18801), .B(n18785), .ZN(n18629) );
  NAND2_X1 U20964 ( .A1(n828), .A2(n18775), .ZN(n18624) );
  NOR2_X1 U20966 ( .A1(n13254), .A2(n12317), .ZN(n13408) );
  NOR2_X1 U20970 ( .A1(n1048), .A2(n31726), .ZN(n18975) );
  NOR2_X1 U20972 ( .A1(n19097), .A2(n19098), .ZN(n14030) );
  NAND2_X1 U20973 ( .A1(n21095), .A2(n8190), .ZN(n21295) );
  AOI21_X1 U20975 ( .A1(n26782), .A2(n15838), .B(n21793), .ZN(n21791) );
  NOR2_X1 U20977 ( .A1(n14488), .A2(n29497), .ZN(n14487) );
  NOR2_X1 U20978 ( .A1(n14489), .A2(n21412), .ZN(n14488) );
  NAND3_X1 U20981 ( .A1(n21084), .A2(n28406), .A3(n17985), .ZN(n13315) );
  NAND3_X1 U20987 ( .A1(n9), .A2(n15956), .A3(n18829), .ZN(n17135) );
  NAND2_X1 U20993 ( .A1(n16624), .A2(n16417), .ZN(n12799) );
  AOI21_X1 U20995 ( .A1(n10828), .A2(n19165), .B(n19308), .ZN(n15930) );
  NAND2_X1 U20997 ( .A1(n17737), .A2(n17736), .ZN(n17735) );
  NAND2_X1 U21009 ( .A1(n19037), .A2(n2901), .ZN(n14455) );
  NAND2_X1 U21010 ( .A1(n16916), .A2(n27587), .ZN(n12645) );
  INV_X1 U21013 ( .I(n33698), .ZN(n19767) );
  NAND3_X1 U21014 ( .A1(n19255), .A2(n19143), .A3(n1180), .ZN(n18528) );
  NOR2_X1 U21018 ( .A1(n30205), .A2(n137), .ZN(n13485) );
  INV_X1 U21022 ( .I(n22536), .ZN(n12844) );
  NAND2_X1 U21031 ( .A1(n20255), .A2(n16951), .ZN(n13380) );
  INV_X1 U21040 ( .I(n22619), .ZN(n15349) );
  NAND2_X1 U21042 ( .A1(n7957), .A2(n708), .ZN(n22253) );
  INV_X1 U21044 ( .I(n23218), .ZN(n23250) );
  NAND2_X1 U21046 ( .A1(n19947), .A2(n15110), .ZN(n15109) );
  OAI21_X1 U21047 ( .A1(n11958), .A2(n20056), .B(n14099), .ZN(n17945) );
  NAND2_X1 U21051 ( .A1(n23637), .A2(n13137), .ZN(n13136) );
  NOR2_X1 U21054 ( .A1(n23797), .A2(n14193), .ZN(n15187) );
  INV_X1 U21057 ( .I(n23490), .ZN(n17194) );
  INV_X1 U21058 ( .I(n23583), .ZN(n14523) );
  OAI21_X1 U21061 ( .A1(n23653), .A2(n8547), .B(n13140), .ZN(n13139) );
  NAND2_X1 U21066 ( .A1(n13905), .A2(n23759), .ZN(n13904) );
  INV_X1 U21068 ( .I(n23958), .ZN(n23957) );
  INV_X1 U21073 ( .I(n16634), .ZN(n15000) );
  INV_X1 U21074 ( .I(n13698), .ZN(n16826) );
  INV_X1 U21075 ( .I(n13060), .ZN(n12513) );
  INV_X1 U21077 ( .I(n11974), .ZN(n14020) );
  NOR2_X1 U21081 ( .A1(n24975), .A2(n25012), .ZN(n14992) );
  NAND2_X1 U21084 ( .A1(n13349), .A2(n4993), .ZN(n24733) );
  NOR2_X1 U21089 ( .A1(n15756), .A2(n16451), .ZN(n15755) );
  NOR2_X1 U21091 ( .A1(n15770), .A2(n28136), .ZN(n15757) );
  INV_X2 U21092 ( .I(n17044), .ZN(n25536) );
  NOR2_X1 U21093 ( .A1(n11900), .A2(n11090), .ZN(n13323) );
  NAND2_X1 U21097 ( .A1(n965), .A2(n24960), .ZN(n14933) );
  OAI21_X1 U21099 ( .A1(n12783), .A2(n33434), .B(n12204), .ZN(n12203) );
  NAND2_X1 U21100 ( .A1(n24972), .A2(n8622), .ZN(n12204) );
  NAND2_X1 U21101 ( .A1(n24969), .A2(n24970), .ZN(n13737) );
  INV_X1 U21103 ( .I(n14638), .ZN(n14637) );
  NAND2_X1 U21104 ( .A1(n1074), .A2(n72), .ZN(n15858) );
  INV_X1 U21109 ( .I(n20953), .ZN(n20997) );
  NAND3_X1 U21110 ( .A1(n20498), .A2(n20497), .A3(n30869), .ZN(n16759) );
  NAND2_X1 U21115 ( .A1(n20461), .A2(n20462), .ZN(n13546) );
  INV_X1 U21116 ( .I(n20773), .ZN(n12732) );
  NAND2_X1 U21117 ( .A1(n13700), .A2(n21182), .ZN(n12913) );
  NAND3_X1 U21119 ( .A1(n14486), .A2(n14485), .A3(n16584), .ZN(n14294) );
  NAND2_X1 U21120 ( .A1(n10182), .A2(n11459), .ZN(n15575) );
  NOR2_X1 U21125 ( .A1(n18797), .A2(n16420), .ZN(n17926) );
  NOR2_X1 U21128 ( .A1(n1017), .A2(n21267), .ZN(n21064) );
  INV_X1 U21134 ( .I(n12654), .ZN(n14860) );
  OAI21_X1 U21136 ( .A1(n14802), .A2(n21379), .B(n7007), .ZN(n21179) );
  NAND2_X1 U21139 ( .A1(n13506), .A2(n21424), .ZN(n17666) );
  NOR2_X1 U21141 ( .A1(n13149), .A2(n21634), .ZN(n13148) );
  NOR2_X1 U21143 ( .A1(n21366), .A2(n21365), .ZN(n12348) );
  AOI21_X1 U21146 ( .A1(n6783), .A2(n962), .B(n12290), .ZN(n12197) );
  NOR2_X1 U21148 ( .A1(n9423), .A2(n19355), .ZN(n16750) );
  AOI21_X1 U21152 ( .A1(n13787), .A2(n9437), .B(n18638), .ZN(n13201) );
  NAND2_X1 U21155 ( .A1(n19268), .A2(n18974), .ZN(n18449) );
  NAND2_X1 U21158 ( .A1(n16487), .A2(n18706), .ZN(n18708) );
  NOR2_X1 U21159 ( .A1(n33078), .A2(n19178), .ZN(n14426) );
  NOR2_X1 U21160 ( .A1(n4016), .A2(n19348), .ZN(n19218) );
  AOI21_X1 U21164 ( .A1(n15874), .A2(n27955), .B(n21143), .ZN(n15024) );
  NAND3_X1 U21165 ( .A1(n29552), .A2(n6176), .A3(n21772), .ZN(n14868) );
  NAND2_X1 U21169 ( .A1(n31826), .A2(n26021), .ZN(n12507) );
  NOR2_X1 U21171 ( .A1(n21052), .A2(n21257), .ZN(n14643) );
  NAND2_X1 U21172 ( .A1(n8631), .A2(n2738), .ZN(n14853) );
  INV_X1 U21175 ( .I(n22021), .ZN(n22162) );
  NAND2_X1 U21178 ( .A1(n15774), .A2(n21812), .ZN(n13167) );
  AOI21_X1 U21182 ( .A1(n19323), .A2(n19317), .B(n19324), .ZN(n12384) );
  AND2_X1 U21183 ( .A1(n6416), .A2(n16538), .Z(n14696) );
  INV_X1 U21184 ( .I(n17165), .ZN(n18865) );
  AOI21_X1 U21188 ( .A1(n18432), .A2(n18433), .B(n18743), .ZN(n13501) );
  INV_X1 U21191 ( .I(n18135), .ZN(n12928) );
  NAND2_X1 U21193 ( .A1(n19114), .A2(n19115), .ZN(n13227) );
  NOR2_X1 U21196 ( .A1(n17455), .A2(n9721), .ZN(n14999) );
  NAND2_X1 U21204 ( .A1(n16447), .A2(n22403), .ZN(n15204) );
  NAND2_X1 U21205 ( .A1(n22678), .A2(n22562), .ZN(n13710) );
  INV_X1 U21206 ( .I(n19878), .ZN(n13987) );
  NAND2_X1 U21209 ( .A1(n33561), .A2(n29013), .ZN(n15737) );
  NOR2_X1 U21211 ( .A1(n18803), .A2(n16403), .ZN(n12175) );
  NOR2_X1 U21214 ( .A1(n3626), .A2(n3790), .ZN(n12590) );
  NOR2_X1 U21218 ( .A1(n6275), .A2(n33264), .ZN(n15267) );
  INV_X1 U21220 ( .I(n28638), .ZN(n17293) );
  INV_X1 U21221 ( .I(n32057), .ZN(n17291) );
  NOR2_X1 U21222 ( .A1(n20059), .A2(n17608), .ZN(n19420) );
  NOR2_X1 U21227 ( .A1(n12112), .A2(n22610), .ZN(n14157) );
  NOR2_X1 U21229 ( .A1(n15008), .A2(n22570), .ZN(n14081) );
  NAND2_X1 U21233 ( .A1(n22503), .A2(n34125), .ZN(n12254) );
  AOI21_X1 U21234 ( .A1(n15322), .A2(n701), .B(n22434), .ZN(n14591) );
  NAND2_X1 U21237 ( .A1(n873), .A2(n19819), .ZN(n13451) );
  INV_X1 U21239 ( .I(n20133), .ZN(n20025) );
  OAI21_X1 U21240 ( .A1(n19987), .A2(n16623), .B(n14440), .ZN(n19339) );
  NOR2_X1 U21241 ( .A1(n19986), .A2(n19998), .ZN(n14622) );
  NOR2_X1 U21242 ( .A1(n19308), .A2(n19165), .ZN(n17526) );
  INV_X1 U21248 ( .I(n20079), .ZN(n19803) );
  NOR2_X1 U21261 ( .A1(n137), .A2(n31964), .ZN(n14160) );
  NAND2_X1 U21271 ( .A1(n15230), .A2(n6996), .ZN(n20400) );
  NAND2_X1 U21274 ( .A1(n13499), .A2(n16144), .ZN(n14265) );
  NAND2_X1 U21276 ( .A1(n22490), .A2(n22489), .ZN(n12930) );
  AND2_X1 U21279 ( .A1(n16078), .A2(n23003), .Z(n11929) );
  NAND2_X1 U21280 ( .A1(n23848), .A2(n23847), .ZN(n13576) );
  NOR2_X1 U21282 ( .A1(n20239), .A2(n20238), .ZN(n17317) );
  NAND2_X1 U21283 ( .A1(n1255), .A2(n14164), .ZN(n13982) );
  OAI22_X1 U21287 ( .A1(n17665), .A2(n13125), .B1(n16431), .B2(n23951), .ZN(
        n17664) );
  NAND3_X1 U21298 ( .A1(n23528), .A2(n23933), .A3(n23681), .ZN(n12546) );
  NAND2_X1 U21299 ( .A1(n23698), .A2(n23867), .ZN(n13138) );
  NOR2_X1 U21301 ( .A1(n13048), .A2(n24276), .ZN(n13047) );
  NAND3_X1 U21304 ( .A1(n16343), .A2(n16496), .A3(n29965), .ZN(n23131) );
  NOR2_X1 U21308 ( .A1(n24150), .A2(n797), .ZN(n12189) );
  NAND2_X1 U21312 ( .A1(n23718), .A2(n13031), .ZN(n14924) );
  NAND3_X1 U21317 ( .A1(n23770), .A2(n11567), .A3(n23769), .ZN(n15402) );
  INV_X1 U21318 ( .I(n12775), .ZN(n12774) );
  NOR2_X1 U21329 ( .A1(n24153), .A2(n1245), .ZN(n16983) );
  NOR2_X1 U21331 ( .A1(n25013), .A2(n31274), .ZN(n14021) );
  NAND2_X1 U21333 ( .A1(n17110), .A2(n7081), .ZN(n25197) );
  AOI21_X1 U21336 ( .A1(n17038), .A2(n25539), .B(n24667), .ZN(n16828) );
  INV_X1 U21337 ( .I(n25876), .ZN(n17762) );
  OAI21_X1 U21340 ( .A1(n25398), .A2(n25403), .B(n25397), .ZN(n15882) );
  NOR2_X1 U21342 ( .A1(n31783), .A2(n25198), .ZN(n15705) );
  NOR2_X1 U21350 ( .A1(n11090), .A2(n25582), .ZN(n15598) );
  OAI21_X1 U21351 ( .A1(n11945), .A2(n17118), .B(n15046), .ZN(n24462) );
  NAND2_X1 U21354 ( .A1(n24955), .A2(n24956), .ZN(n14932) );
  NAND2_X1 U21357 ( .A1(n30302), .A2(n25375), .ZN(n15478) );
  OAI21_X1 U21361 ( .A1(n14454), .A2(n15084), .B(n15223), .ZN(n17771) );
  NOR2_X1 U21365 ( .A1(n27118), .A2(n1223), .ZN(n15673) );
  INV_X1 U21371 ( .I(n17594), .ZN(n15332) );
  NAND3_X1 U21372 ( .A1(n14627), .A2(n15641), .A3(n25145), .ZN(n14631) );
  NOR2_X1 U21373 ( .A1(n25199), .A2(n12476), .ZN(n25147) );
  NAND2_X1 U21374 ( .A1(n966), .A2(n25214), .ZN(n25215) );
  NAND2_X1 U21375 ( .A1(n25231), .A2(n25398), .ZN(n17924) );
  NOR2_X1 U21376 ( .A1(n15770), .A2(n17717), .ZN(n15896) );
  NAND2_X1 U21379 ( .A1(n25369), .A2(n25376), .ZN(n16246) );
  NAND2_X1 U21380 ( .A1(n24863), .A2(n9858), .ZN(n16187) );
  AOI21_X1 U21381 ( .A1(n25564), .A2(n17655), .B(n25582), .ZN(n13322) );
  NAND3_X1 U21382 ( .A1(n25752), .A2(n25707), .A3(n25620), .ZN(n25580) );
  NAND2_X1 U21385 ( .A1(n13768), .A2(n20236), .ZN(n12224) );
  NAND2_X1 U21391 ( .A1(n15006), .A2(n20417), .ZN(n20274) );
  NOR2_X1 U21398 ( .A1(n33515), .A2(n13759), .ZN(n13786) );
  NAND2_X1 U21399 ( .A1(n13880), .A2(n20524), .ZN(n12345) );
  INV_X1 U21402 ( .I(n20498), .ZN(n16762) );
  NOR2_X1 U21404 ( .A1(n2618), .A2(n30987), .ZN(n17758) );
  NOR2_X1 U21405 ( .A1(n31835), .A2(n865), .ZN(n16505) );
  NAND3_X1 U21406 ( .A1(n17971), .A2(n28502), .A3(n21251), .ZN(n20935) );
  NAND3_X1 U21407 ( .A1(n779), .A2(n16933), .A3(n21249), .ZN(n20936) );
  INV_X1 U21413 ( .I(n17984), .ZN(n16780) );
  NOR2_X1 U21415 ( .A1(n21473), .A2(n27532), .ZN(n12275) );
  INV_X1 U21418 ( .I(n13872), .ZN(n21458) );
  NAND2_X1 U21424 ( .A1(n17687), .A2(n18738), .ZN(n18531) );
  NAND2_X1 U21425 ( .A1(n28171), .A2(n878), .ZN(n12807) );
  NAND2_X1 U21426 ( .A1(n882), .A2(n28707), .ZN(n15927) );
  OAI21_X1 U21429 ( .A1(n18843), .A2(n746), .B(n25981), .ZN(n16713) );
  NAND2_X1 U21430 ( .A1(n19321), .A2(n19322), .ZN(n19232) );
  AOI22_X1 U21436 ( .A1(n12130), .A2(n30271), .B1(n13846), .B2(n18699), .ZN(
        n15196) );
  NOR2_X1 U21438 ( .A1(n13200), .A2(n19180), .ZN(n19182) );
  INV_X1 U21440 ( .I(n19507), .ZN(n12683) );
  NAND2_X1 U21443 ( .A1(n21668), .A2(n918), .ZN(n14673) );
  NAND2_X1 U21445 ( .A1(n17547), .A2(n7553), .ZN(n12786) );
  INV_X1 U21446 ( .I(n14950), .ZN(n14949) );
  NAND2_X1 U21449 ( .A1(n16519), .A2(n16165), .ZN(n12712) );
  NAND2_X1 U21450 ( .A1(n27336), .A2(n432), .ZN(n16863) );
  INV_X1 U21455 ( .I(n34040), .ZN(n19263) );
  NAND2_X1 U21456 ( .A1(n19269), .A2(n19265), .ZN(n15505) );
  NOR2_X1 U21459 ( .A1(n18581), .A2(n17419), .ZN(n13036) );
  NOR2_X1 U21460 ( .A1(n16403), .A2(n18785), .ZN(n18786) );
  NAND2_X1 U21461 ( .A1(n4677), .A2(n18801), .ZN(n18787) );
  NAND2_X1 U21462 ( .A1(n746), .A2(n15873), .ZN(n16867) );
  NAND2_X1 U21463 ( .A1(n16370), .A2(n6783), .ZN(n12196) );
  NAND2_X1 U21471 ( .A1(n19181), .A2(n19118), .ZN(n13012) );
  OAI21_X1 U21475 ( .A1(n18467), .A2(n18468), .B(n945), .ZN(n13708) );
  NAND2_X1 U21477 ( .A1(n18532), .A2(n17166), .ZN(n15583) );
  AOI21_X1 U21479 ( .A1(n15685), .A2(n18254), .B(n18434), .ZN(n18709) );
  INV_X1 U21480 ( .I(n18704), .ZN(n15685) );
  NOR2_X1 U21481 ( .A1(n33205), .A2(n16287), .ZN(n17359) );
  NOR2_X1 U21495 ( .A1(n919), .A2(n21687), .ZN(n12332) );
  NOR2_X1 U21497 ( .A1(n13500), .A2(n21641), .ZN(n13613) );
  NOR2_X1 U21500 ( .A1(n16519), .A2(n16165), .ZN(n14503) );
  OAI21_X1 U21501 ( .A1(n21840), .A2(n16987), .B(n26163), .ZN(n13815) );
  NOR2_X1 U21504 ( .A1(n29854), .A2(n9076), .ZN(n15680) );
  INV_X1 U21509 ( .I(n22160), .ZN(n17968) );
  NAND2_X1 U21512 ( .A1(n21731), .A2(n15655), .ZN(n12939) );
  NOR2_X1 U21516 ( .A1(n14976), .A2(n14172), .ZN(n20093) );
  INV_X1 U21523 ( .I(n22220), .ZN(n12681) );
  NOR2_X1 U21528 ( .A1(n31017), .A2(n34103), .ZN(n13655) );
  AOI21_X1 U21529 ( .A1(n19862), .A2(n16579), .B(n19863), .ZN(n18002) );
  NOR3_X1 U21530 ( .A1(n34103), .A2(n14458), .A3(n31017), .ZN(n14282) );
  NAND3_X1 U21534 ( .A1(n14747), .A2(n11959), .A3(n3486), .ZN(n13570) );
  NOR3_X1 U21535 ( .A1(n20142), .A2(n11911), .A3(n11248), .ZN(n12851) );
  INV_X1 U21540 ( .I(n19984), .ZN(n12397) );
  AOI21_X1 U21541 ( .A1(n22803), .A2(n22983), .B(n16140), .ZN(n12596) );
  NOR2_X1 U21546 ( .A1(n22805), .A2(n14420), .ZN(n14419) );
  NAND2_X1 U21549 ( .A1(n22798), .A2(n23053), .ZN(n22868) );
  INV_X1 U21551 ( .I(n23336), .ZN(n14583) );
  NAND3_X1 U21552 ( .A1(n11980), .A2(n13892), .A3(n16486), .ZN(n15577) );
  NAND2_X1 U21554 ( .A1(n13575), .A2(n22780), .ZN(n13574) );
  OAI21_X1 U21558 ( .A1(n3184), .A2(n3183), .B(n22781), .ZN(n16716) );
  NOR2_X1 U21559 ( .A1(n28948), .A2(n17084), .ZN(n14603) );
  AOI21_X1 U21562 ( .A1(n31684), .A2(n13061), .B(n29013), .ZN(n14989) );
  NAND2_X1 U21564 ( .A1(n26232), .A2(n20577), .ZN(n20579) );
  OAI21_X1 U21565 ( .A1(n20153), .A2(n11199), .B(n20150), .ZN(n15350) );
  NAND2_X1 U21568 ( .A1(n19812), .A2(n20018), .ZN(n19814) );
  NAND2_X1 U21575 ( .A1(n22952), .A2(n2479), .ZN(n13004) );
  NAND2_X1 U21578 ( .A1(n28277), .A2(n25994), .ZN(n13251) );
  AOI21_X1 U21582 ( .A1(n13995), .A2(n23106), .B(n14131), .ZN(n14552) );
  INV_X1 U21588 ( .I(n23375), .ZN(n23260) );
  INV_X1 U21596 ( .I(n23507), .ZN(n13287) );
  NAND2_X1 U21605 ( .A1(n16167), .A2(n20510), .ZN(n14366) );
  NOR2_X1 U21607 ( .A1(n20228), .A2(n7242), .ZN(n20516) );
  NOR2_X1 U21609 ( .A1(n20337), .A2(n20531), .ZN(n14261) );
  OAI21_X1 U21611 ( .A1(n15806), .A2(n22865), .B(n989), .ZN(n22707) );
  INV_X1 U21614 ( .I(n16076), .ZN(n23321) );
  NAND2_X1 U21616 ( .A1(n20240), .A2(n27386), .ZN(n16857) );
  INV_X1 U21619 ( .I(n24226), .ZN(n24042) );
  NAND3_X1 U21621 ( .A1(n24325), .A2(n7361), .A3(n24245), .ZN(n24079) );
  INV_X1 U21622 ( .I(n24276), .ZN(n24195) );
  OR3_X1 U21625 ( .A1(n27430), .A2(n24304), .A3(n12904), .Z(n11937) );
  NAND2_X1 U21628 ( .A1(n13082), .A2(n32737), .ZN(n12629) );
  AOI21_X1 U21639 ( .A1(n12189), .A2(n2913), .B(n12188), .ZN(n12187) );
  OAI21_X1 U21643 ( .A1(n791), .A2(n26916), .B(n12357), .ZN(n23626) );
  NOR2_X1 U21645 ( .A1(n24270), .A2(n11768), .ZN(n14502) );
  INV_X1 U21646 ( .I(n3935), .ZN(n14938) );
  NAND3_X1 U21650 ( .A1(n14889), .A2(n28694), .A3(n16621), .ZN(n14888) );
  OAI21_X1 U21651 ( .A1(n28694), .A2(n17261), .B(n13260), .ZN(n24229) );
  NAND2_X1 U21652 ( .A1(n1786), .A2(n1850), .ZN(n15254) );
  INV_X1 U21654 ( .I(n24816), .ZN(n18217) );
  INV_X1 U21656 ( .I(n24403), .ZN(n12240) );
  NAND2_X1 U21657 ( .A1(n317), .A2(n15880), .ZN(n14139) );
  INV_X1 U21659 ( .I(n25584), .ZN(n18196) );
  NOR2_X1 U21661 ( .A1(n10755), .A2(n14752), .ZN(n24912) );
  NAND2_X1 U21662 ( .A1(n25258), .A2(n17273), .ZN(n14511) );
  NOR2_X1 U21663 ( .A1(n14960), .A2(n8622), .ZN(n16383) );
  NAND2_X1 U21665 ( .A1(n18151), .A2(n28096), .ZN(n15185) );
  NOR2_X1 U21666 ( .A1(n1209), .A2(n32897), .ZN(n25496) );
  INV_X1 U21667 ( .I(n25058), .ZN(n25050) );
  NAND2_X1 U21673 ( .A1(n25705), .A2(n11944), .ZN(n13359) );
  AOI21_X1 U21675 ( .A1(n32856), .A2(n25615), .B(n9982), .ZN(n25618) );
  INV_X1 U21677 ( .I(n25224), .ZN(n25225) );
  NAND2_X1 U21679 ( .A1(n14780), .A2(n26447), .ZN(n12215) );
  NAND2_X1 U21681 ( .A1(n25605), .A2(n831), .ZN(n13996) );
  OAI21_X1 U21685 ( .A1(n24911), .A2(n10755), .B(n14752), .ZN(n24906) );
  NAND2_X1 U21688 ( .A1(n25861), .A2(n18022), .ZN(n18020) );
  OAI21_X1 U21689 ( .A1(n25052), .A2(n28070), .B(n17744), .ZN(n17743) );
  NAND2_X1 U21690 ( .A1(n15479), .A2(n15478), .ZN(n25356) );
  AOI21_X1 U21693 ( .A1(n3843), .A2(n24965), .B(n13627), .ZN(n12202) );
  AOI21_X1 U21694 ( .A1(n28736), .A2(n14810), .B(n28200), .ZN(n12250) );
  OAI21_X1 U21695 ( .A1(n14634), .A2(n14638), .B(n1420), .ZN(n14633) );
  NAND2_X1 U21696 ( .A1(n27183), .A2(n1074), .ZN(n17708) );
  NAND2_X1 U21699 ( .A1(n25516), .A2(n32897), .ZN(n16468) );
  INV_X1 U21702 ( .I(n24447), .ZN(n25705) );
  XOR2_X1 U21704 ( .A1(Plaintext[145]), .A2(Key[145]), .Z(n11905) );
  INV_X1 U21706 ( .I(n21305), .ZN(n21131) );
  AND2_X1 U21708 ( .A1(n22664), .A2(n14307), .Z(n11928) );
  AND2_X1 U21711 ( .A1(n3843), .A2(n24965), .Z(n11939) );
  AND2_X1 U21714 ( .A1(n25705), .A2(n25707), .Z(n11951) );
  OR2_X1 U21715 ( .A1(n20039), .A2(n20040), .Z(n11952) );
  OR2_X1 U21719 ( .A1(n20411), .A2(n28261), .Z(n11964) );
  NOR2_X1 U21721 ( .A1(n13894), .A2(n13893), .ZN(n11980) );
  XNOR2_X1 U21723 ( .A1(n20822), .A2(n13093), .ZN(n11982) );
  INV_X1 U21724 ( .I(n19355), .ZN(n15842) );
  OR2_X1 U21727 ( .A1(n24610), .A2(n680), .Z(n11994) );
  XNOR2_X1 U21728 ( .A1(n33293), .A2(n25827), .ZN(n11996) );
  AND2_X1 U21729 ( .A1(n25884), .A2(n25872), .Z(n11999) );
  NOR2_X1 U21733 ( .A1(n24112), .A2(n24289), .ZN(n12002) );
  XNOR2_X1 U21737 ( .A1(n23430), .A2(n25224), .ZN(n12014) );
  AND2_X1 U21738 ( .A1(n27166), .A2(n13622), .Z(n12016) );
  AND2_X1 U21739 ( .A1(n781), .A2(n1351), .Z(n12021) );
  AND2_X1 U21740 ( .A1(n969), .A2(n24194), .Z(n12022) );
  AND2_X1 U21741 ( .A1(n16933), .A2(n21249), .Z(n12029) );
  AND2_X1 U21742 ( .A1(n16413), .A2(n11944), .Z(n12030) );
  NAND3_X1 U21743 ( .A1(n16688), .A2(n1096), .A3(n24218), .ZN(n24043) );
  OR2_X2 U21747 ( .A1(n12384), .A2(n12382), .Z(n12048) );
  OR2_X1 U21750 ( .A1(n14458), .A2(n31017), .Z(n12053) );
  XNOR2_X1 U21756 ( .A1(n31499), .A2(n24417), .ZN(n12059) );
  XNOR2_X1 U21757 ( .A1(n17145), .A2(n22041), .ZN(n12062) );
  AND2_X1 U21758 ( .A1(n15909), .A2(n18757), .Z(n12065) );
  INV_X1 U21759 ( .I(n25916), .ZN(n25926) );
  INV_X1 U21761 ( .I(n16778), .ZN(n25400) );
  INV_X1 U21765 ( .I(n22412), .ZN(n22639) );
  XNOR2_X1 U21766 ( .A1(n22029), .A2(n25722), .ZN(n12082) );
  INV_X1 U21770 ( .I(n11944), .ZN(n25706) );
  INV_X1 U21775 ( .I(n24168), .ZN(n24194) );
  XNOR2_X1 U21777 ( .A1(n22034), .A2(n22035), .ZN(n12101) );
  INV_X1 U21778 ( .I(n23639), .ZN(n23873) );
  XNOR2_X1 U21779 ( .A1(n8298), .A2(n23436), .ZN(n12104) );
  INV_X1 U21784 ( .I(n23132), .ZN(n14464) );
  AND2_X1 U21789 ( .A1(n23487), .A2(n23486), .Z(n12122) );
  INV_X1 U21790 ( .I(n18973), .ZN(n19271) );
  XNOR2_X1 U21791 ( .A1(n15130), .A2(n25086), .ZN(n12123) );
  XNOR2_X1 U21792 ( .A1(n34078), .A2(n16551), .ZN(n12124) );
  XNOR2_X1 U21795 ( .A1(n22130), .A2(n24869), .ZN(n12127) );
  XNOR2_X1 U21798 ( .A1(n19736), .A2(n24968), .ZN(n12136) );
  XNOR2_X1 U21799 ( .A1(n19566), .A2(n16523), .ZN(n12137) );
  AND2_X1 U21802 ( .A1(n20456), .A2(n14086), .Z(n12139) );
  INV_X1 U21804 ( .I(n13401), .ZN(n21059) );
  XNOR2_X1 U21805 ( .A1(n19630), .A2(n25476), .ZN(n12141) );
  INV_X1 U21806 ( .I(n27698), .ZN(n19808) );
  INV_X2 U21809 ( .I(n16682), .ZN(n22634) );
  INV_X1 U21810 ( .I(n16587), .ZN(n15566) );
  INV_X1 U21811 ( .I(n8548), .ZN(n17723) );
  INV_X1 U21813 ( .I(n25545), .ZN(n15816) );
  INV_X1 U21815 ( .I(n16687), .ZN(n17986) );
  INV_X1 U21816 ( .I(n25864), .ZN(n18019) );
  INV_X1 U21817 ( .I(n16550), .ZN(n13394) );
  INV_X1 U21818 ( .I(n8487), .ZN(n16438) );
  INV_X1 U21821 ( .I(n16698), .ZN(n14648) );
  INV_X1 U21822 ( .I(n16507), .ZN(n13091) );
  INV_X1 U21824 ( .I(n16597), .ZN(n16038) );
  INV_X1 U21826 ( .I(n25086), .ZN(n13331) );
  INV_X1 U21827 ( .I(n24962), .ZN(n15415) );
  INV_X1 U21828 ( .I(n16533), .ZN(n18102) );
  INV_X2 U21829 ( .I(n13567), .ZN(n15255) );
  INV_X2 U21834 ( .I(n16310), .ZN(n17813) );
  NAND2_X1 U21835 ( .A1(n27651), .A2(n25119), .ZN(n12163) );
  XNOR2_X1 U21836 ( .A1(Plaintext[164]), .A2(Key[164]), .ZN(n12166) );
  XOR2_X1 U21837 ( .A1(n20983), .A2(n12171), .Z(n12170) );
  XOR2_X1 U21838 ( .A1(n20758), .A2(n20621), .Z(n12172) );
  XNOR2_X1 U21839 ( .A1(n18083), .A2(n19374), .ZN(n12182) );
  XOR2_X1 U21840 ( .A1(n4975), .A2(n32367), .Z(n19751) );
  NAND2_X1 U21841 ( .A1(n17525), .A2(n1850), .ZN(n18132) );
  XOR2_X1 U21843 ( .A1(n14841), .A2(n14136), .Z(n12185) );
  XOR2_X1 U21846 ( .A1(n23391), .A2(n25911), .Z(n12200) );
  NAND2_X1 U21850 ( .A1(n28263), .A2(n28669), .ZN(n12209) );
  XOR2_X1 U21852 ( .A1(n12223), .A2(n12410), .Z(n12409) );
  NOR2_X1 U21854 ( .A1(n22590), .A2(n12236), .ZN(n17584) );
  XOR2_X1 U21855 ( .A1(n22028), .A2(n16548), .Z(n16816) );
  XOR2_X1 U21857 ( .A1(n24741), .A2(n12240), .Z(n12239) );
  NAND2_X2 U21858 ( .A1(n14674), .A2(n14673), .ZN(n21726) );
  XOR2_X1 U21860 ( .A1(n12252), .A2(n25252), .Z(n18108) );
  XOR2_X1 U21861 ( .A1(n12252), .A2(n14583), .Z(n14582) );
  XOR2_X1 U21872 ( .A1(n19764), .A2(n17600), .Z(n12283) );
  XOR2_X1 U21873 ( .A1(n12286), .A2(n12285), .Z(n12284) );
  XOR2_X1 U21874 ( .A1(n5348), .A2(n24953), .Z(n12285) );
  XOR2_X1 U21875 ( .A1(n28813), .A2(n12494), .Z(n12286) );
  XOR2_X1 U21877 ( .A1(n23279), .A2(n23278), .Z(n12288) );
  NAND2_X1 U21879 ( .A1(n28450), .A2(n15864), .ZN(n14524) );
  NAND2_X1 U21880 ( .A1(n534), .A2(n28450), .ZN(n21873) );
  AND2_X1 U21882 ( .A1(n12085), .A2(n15057), .Z(n12300) );
  NAND3_X2 U21884 ( .A1(n19955), .A2(n19956), .A3(n19954), .ZN(n14858) );
  NAND2_X2 U21885 ( .A1(n12616), .A2(n12553), .ZN(n16173) );
  XOR2_X1 U21887 ( .A1(n12313), .A2(n27125), .Z(n16972) );
  NOR2_X1 U21888 ( .A1(n25676), .A2(n12314), .ZN(n25677) );
  NOR2_X1 U21891 ( .A1(n12315), .A2(n15456), .ZN(n15729) );
  NAND3_X1 U21892 ( .A1(n12727), .A2(n22715), .A3(n12315), .ZN(n22717) );
  OAI21_X1 U21893 ( .A1(n18727), .A2(n11123), .B(n18726), .ZN(n18729) );
  NAND2_X1 U21897 ( .A1(n12325), .A2(n21400), .ZN(n21096) );
  MUX2_X1 U21901 ( .I0(n32900), .I1(n12329), .S(n10822), .Z(n25081) );
  XOR2_X1 U21904 ( .A1(n11324), .A2(n12387), .Z(n12331) );
  INV_X2 U21905 ( .I(n12960), .ZN(n16375) );
  XOR2_X1 U21913 ( .A1(n21007), .A2(n27169), .Z(n13395) );
  NAND2_X2 U21916 ( .A1(n14990), .A2(n22833), .ZN(n16799) );
  XOR2_X1 U21917 ( .A1(n24422), .A2(n24215), .Z(n12355) );
  XNOR2_X1 U21918 ( .A1(n24522), .A2(n24618), .ZN(n24422) );
  NAND2_X1 U21920 ( .A1(n26516), .A2(n30146), .ZN(n23659) );
  INV_X2 U21921 ( .I(n15518), .ZN(n25891) );
  XOR2_X1 U21924 ( .A1(n12376), .A2(n25131), .Z(n21050) );
  XOR2_X1 U21927 ( .A1(n19723), .A2(n19667), .Z(n12380) );
  XOR2_X1 U21928 ( .A1(n19584), .A2(n13682), .Z(n12381) );
  AOI21_X1 U21929 ( .A1(n27131), .A2(n12383), .B(n19274), .ZN(n12382) );
  NAND2_X1 U21930 ( .A1(n19318), .A2(n19275), .ZN(n12383) );
  INV_X1 U21932 ( .I(n12390), .ZN(n12392) );
  NOR2_X1 U21934 ( .A1(n20105), .A2(n12398), .ZN(n20454) );
  NOR2_X1 U21936 ( .A1(n14913), .A2(n33295), .ZN(n12402) );
  MUX2_X1 U21937 ( .I0(n24086), .I1(n24085), .S(n14913), .Z(n12403) );
  XOR2_X1 U21940 ( .A1(n19577), .A2(n19380), .Z(n12411) );
  XOR2_X1 U21949 ( .A1(n12456), .A2(n1413), .Z(Ciphertext[63]) );
  XOR2_X1 U21951 ( .A1(n12462), .A2(n612), .Z(n12461) );
  XOR2_X1 U21952 ( .A1(n4057), .A2(n32695), .Z(n12462) );
  XOR2_X1 U21953 ( .A1(n30489), .A2(n4295), .Z(n21898) );
  XOR2_X1 U21961 ( .A1(n13814), .A2(n1198), .Z(n12475) );
  XOR2_X1 U21962 ( .A1(n12944), .A2(n12942), .Z(n25188) );
  INV_X2 U21963 ( .I(n22638), .ZN(n22636) );
  XOR2_X1 U21965 ( .A1(n5381), .A2(n12491), .Z(n22948) );
  XOR2_X1 U21967 ( .A1(n12493), .A2(n24966), .Z(n24389) );
  XOR2_X1 U21968 ( .A1(n12494), .A2(n25098), .Z(n20684) );
  XOR2_X1 U21969 ( .A1(n12494), .A2(n25549), .Z(n20971) );
  AOI21_X1 U21972 ( .A1(n827), .A2(n32485), .B(n12502), .ZN(n19346) );
  INV_X2 U21976 ( .I(n17074), .ZN(n24466) );
  XOR2_X1 U21977 ( .A1(n13849), .A2(n12513), .Z(n12512) );
  NAND2_X1 U21985 ( .A1(n12169), .A2(n12541), .ZN(n12540) );
  NOR2_X2 U21987 ( .A1(n24114), .A2(n16356), .ZN(n23608) );
  XOR2_X1 U21990 ( .A1(n348), .A2(n24386), .Z(n12552) );
  MUX2_X1 U21996 ( .I0(n32397), .I1(n12561), .S(n21646), .Z(n15748) );
  XOR2_X1 U22002 ( .A1(n12573), .A2(n13932), .Z(n13931) );
  INV_X2 U22006 ( .I(n12584), .ZN(n21305) );
  NAND2_X1 U22008 ( .A1(n1175), .A2(n12585), .ZN(n16591) );
  NOR2_X1 U22009 ( .A1(n25961), .A2(n12585), .ZN(n16361) );
  XOR2_X1 U22017 ( .A1(n12610), .A2(n25191), .Z(n19380) );
  NAND2_X1 U22021 ( .A1(n16603), .A2(n23886), .ZN(n12615) );
  OAI21_X1 U22025 ( .A1(n4016), .A2(n14194), .B(n19348), .ZN(n19000) );
  XOR2_X1 U22026 ( .A1(n702), .A2(n17430), .Z(n12620) );
  XOR2_X1 U22029 ( .A1(n24836), .A2(n24764), .Z(n12628) );
  XOR2_X1 U22033 ( .A1(n24750), .A2(n16602), .Z(n12636) );
  OAI21_X2 U22036 ( .A1(n13891), .A2(n13890), .B(n13889), .ZN(n19408) );
  NOR2_X1 U22040 ( .A1(n13210), .A2(n949), .ZN(n12649) );
  XOR2_X1 U22048 ( .A1(n17912), .A2(n12665), .Z(n24625) );
  XOR2_X1 U22050 ( .A1(n20959), .A2(n12673), .Z(n12672) );
  XOR2_X1 U22051 ( .A1(n12675), .A2(n27423), .Z(n13519) );
  INV_X1 U22054 ( .I(n23905), .ZN(n16238) );
  OR2_X1 U22055 ( .A1(n14974), .A2(n12680), .Z(n15943) );
  NAND2_X2 U22058 ( .A1(n25871), .A2(n25885), .ZN(n12699) );
  NAND3_X1 U22059 ( .A1(n941), .A2(n821), .A3(n17608), .ZN(n12704) );
  NOR2_X2 U22061 ( .A1(n18920), .A2(n18921), .ZN(n12707) );
  XOR2_X1 U22063 ( .A1(n13844), .A2(n26002), .Z(n12717) );
  XOR2_X1 U22064 ( .A1(n12721), .A2(n16482), .Z(n20797) );
  XOR2_X1 U22065 ( .A1(n12721), .A2(n16507), .Z(n20915) );
  NAND3_X1 U22066 ( .A1(n22715), .A2(n851), .A3(n12729), .ZN(n22716) );
  OAI21_X1 U22067 ( .A1(n22807), .A2(n12729), .B(n16458), .ZN(n15101) );
  XOR2_X1 U22068 ( .A1(n12731), .A2(n20774), .Z(n21375) );
  XOR2_X1 U22069 ( .A1(n20772), .A2(n12732), .Z(n12731) );
  NOR2_X2 U22073 ( .A1(n21386), .A2(n21385), .ZN(n21630) );
  XOR2_X1 U22075 ( .A1(n9145), .A2(n31687), .Z(n24792) );
  INV_X2 U22076 ( .I(n12735), .ZN(n18110) );
  XOR2_X1 U22078 ( .A1(n23155), .A2(n23414), .Z(n23537) );
  NAND2_X1 U22079 ( .A1(n6842), .A2(n12747), .ZN(n21069) );
  XOR2_X1 U22081 ( .A1(n20995), .A2(n17793), .Z(n12749) );
  XOR2_X1 U22082 ( .A1(n4728), .A2(n16527), .Z(n15573) );
  NAND3_X1 U22083 ( .A1(n16699), .A2(n19335), .A3(n14597), .ZN(n12755) );
  XOR2_X1 U22085 ( .A1(n22189), .A2(n22056), .Z(n12760) );
  XOR2_X1 U22087 ( .A1(n34120), .A2(n23425), .Z(n12765) );
  NOR2_X2 U22094 ( .A1(n17378), .A2(n17379), .ZN(n13627) );
  NAND2_X1 U22095 ( .A1(n21642), .A2(n29234), .ZN(n21473) );
  XOR2_X1 U22096 ( .A1(n12800), .A2(n16548), .Z(n24354) );
  XOR2_X1 U22097 ( .A1(n12795), .A2(n12057), .Z(n15237) );
  XOR2_X1 U22100 ( .A1(Plaintext[169]), .A2(Key[169]), .Z(n15966) );
  XOR2_X1 U22101 ( .A1(n15913), .A2(n19514), .Z(n12803) );
  NAND2_X1 U22103 ( .A1(n12812), .A2(n29069), .ZN(n18270) );
  OAI21_X2 U22106 ( .A1(n12432), .A2(n12816), .B(n14942), .ZN(n24164) );
  NAND2_X2 U22107 ( .A1(n6072), .A2(n1125), .ZN(n22439) );
  XOR2_X1 U22108 ( .A1(n12821), .A2(n25131), .Z(n17500) );
  NOR2_X1 U22115 ( .A1(n12587), .A2(n30291), .ZN(n21606) );
  NOR2_X1 U22116 ( .A1(n2575), .A2(n30291), .ZN(n21759) );
  XOR2_X1 U22119 ( .A1(n30171), .A2(n24943), .Z(n15993) );
  OR2_X1 U22120 ( .A1(n15022), .A2(n21761), .Z(n12853) );
  AOI21_X2 U22121 ( .A1(n12855), .A2(n26386), .B(n21606), .ZN(n21952) );
  INV_X2 U22122 ( .I(n23579), .ZN(n23833) );
  OR2_X1 U22123 ( .A1(n24219), .A2(n16554), .Z(n12861) );
  XOR2_X1 U22124 ( .A1(Plaintext[45]), .A2(Key[45]), .Z(n18777) );
  XOR2_X1 U22125 ( .A1(n28977), .A2(n27125), .Z(n13741) );
  XOR2_X1 U22126 ( .A1(n20730), .A2(n20842), .Z(n20732) );
  XOR2_X1 U22131 ( .A1(n14215), .A2(n19559), .Z(n12896) );
  XOR2_X1 U22136 ( .A1(n24761), .A2(n16584), .Z(n12905) );
  XOR2_X1 U22137 ( .A1(n23517), .A2(n12955), .Z(n12954) );
  INV_X1 U22138 ( .I(n12907), .ZN(n12908) );
  XOR2_X1 U22141 ( .A1(n12915), .A2(n13529), .Z(n21965) );
  XOR2_X1 U22142 ( .A1(n20704), .A2(n12916), .Z(n20931) );
  XOR2_X1 U22143 ( .A1(n20768), .A2(n20703), .Z(n12916) );
  XOR2_X1 U22145 ( .A1(Plaintext[121]), .A2(Key[121]), .Z(n14409) );
  XOR2_X1 U22146 ( .A1(n24793), .A2(n12918), .Z(n14065) );
  OAI21_X1 U22147 ( .A1(n16600), .A2(n2217), .B(n6660), .ZN(n12919) );
  XOR2_X1 U22150 ( .A1(n23529), .A2(n12922), .Z(n12921) );
  XOR2_X1 U22154 ( .A1(n24473), .A2(n18042), .Z(n12936) );
  XOR2_X1 U22157 ( .A1(n24838), .A2(n12943), .Z(n12942) );
  XOR2_X1 U22159 ( .A1(n24835), .A2(n24834), .Z(n12944) );
  XOR2_X1 U22160 ( .A1(n11751), .A2(n12945), .Z(n24835) );
  NAND3_X1 U22163 ( .A1(n30375), .A2(n20028), .A3(n28423), .ZN(n19905) );
  MUX2_X1 U22164 ( .I0(n19805), .I1(n19806), .S(n19724), .Z(n19807) );
  AOI21_X1 U22165 ( .A1(n30271), .A2(n13846), .B(n27687), .ZN(n18390) );
  XOR2_X1 U22167 ( .A1(n23262), .A2(n23444), .Z(n12955) );
  NOR2_X1 U22168 ( .A1(n12956), .A2(n18848), .ZN(n18593) );
  NOR2_X1 U22169 ( .A1(n12956), .A2(n17184), .ZN(n18594) );
  OAI21_X1 U22170 ( .A1(n15967), .A2(n12956), .B(n18846), .ZN(n18734) );
  NAND2_X1 U22171 ( .A1(n31972), .A2(n10283), .ZN(n18870) );
  XOR2_X1 U22173 ( .A1(n12957), .A2(n24426), .Z(n13404) );
  XOR2_X1 U22174 ( .A1(n20720), .A2(n12957), .Z(n20721) );
  XOR2_X1 U22175 ( .A1(n23438), .A2(n12934), .Z(n23283) );
  XOR2_X1 U22177 ( .A1(n12959), .A2(n18072), .Z(n12958) );
  XOR2_X1 U22178 ( .A1(n28908), .A2(n25541), .Z(n12959) );
  XOR2_X1 U22179 ( .A1(n22000), .A2(n22002), .Z(n12962) );
  XOR2_X1 U22182 ( .A1(n32648), .A2(n20905), .Z(n13179) );
  XOR2_X1 U22184 ( .A1(n27211), .A2(n12969), .Z(n12971) );
  NOR2_X1 U22186 ( .A1(n12973), .A2(n28869), .ZN(n21121) );
  AOI21_X1 U22188 ( .A1(n7203), .A2(n33295), .B(n24139), .ZN(n12985) );
  INV_X2 U22191 ( .I(n13177), .ZN(n21095) );
  NAND3_X1 U22192 ( .A1(n19255), .A2(n19143), .A3(n19252), .ZN(n12993) );
  NOR2_X2 U22193 ( .A1(n19791), .A2(n19790), .ZN(n20582) );
  NOR2_X1 U22196 ( .A1(n9484), .A2(n868), .ZN(n13880) );
  XOR2_X1 U22198 ( .A1(n19676), .A2(n29515), .Z(n19677) );
  XOR2_X1 U22199 ( .A1(n33749), .A2(n29515), .Z(n19377) );
  INV_X2 U22201 ( .I(n13022), .ZN(n17731) );
  NAND2_X1 U22203 ( .A1(n18738), .A2(n18737), .ZN(n13024) );
  NOR2_X1 U22204 ( .A1(n2378), .A2(n13032), .ZN(n24446) );
  NAND2_X1 U22205 ( .A1(n15155), .A2(n13032), .ZN(n25714) );
  XOR2_X1 U22208 ( .A1(n20820), .A2(n13041), .Z(n17576) );
  XOR2_X1 U22209 ( .A1(n13041), .A2(n25079), .Z(n20988) );
  XOR2_X1 U22214 ( .A1(n13065), .A2(n16662), .Z(Ciphertext[66]) );
  INV_X1 U22215 ( .I(n13067), .ZN(n15795) );
  NOR2_X1 U22216 ( .A1(n3880), .A2(n24084), .ZN(n16100) );
  AND2_X1 U22217 ( .A1(n3880), .A2(n16286), .Z(n15010) );
  INV_X1 U22220 ( .I(n22303), .ZN(n13075) );
  NOR2_X1 U22221 ( .A1(n18781), .A2(n10080), .ZN(n13076) );
  INV_X2 U22223 ( .I(n13080), .ZN(n17711) );
  XOR2_X1 U22226 ( .A1(n24524), .A2(n13086), .Z(n13085) );
  NOR2_X1 U22228 ( .A1(n20439), .A2(n14863), .ZN(n13090) );
  XOR2_X1 U22229 ( .A1(n13106), .A2(n13095), .Z(n19554) );
  XOR2_X1 U22232 ( .A1(n19379), .A2(n24065), .Z(n13099) );
  NAND2_X1 U22233 ( .A1(n8412), .A2(n24271), .ZN(n15899) );
  NOR2_X1 U22234 ( .A1(n23555), .A2(n23806), .ZN(n17701) );
  NAND2_X1 U22237 ( .A1(n32874), .A2(n25795), .ZN(n15304) );
  NAND2_X1 U22238 ( .A1(n15242), .A2(n1009), .ZN(n15676) );
  NAND2_X1 U22239 ( .A1(n17467), .A2(n27382), .ZN(n20932) );
  OAI21_X1 U22244 ( .A1(n14312), .A2(n10700), .B(n15143), .ZN(n17617) );
  NOR2_X1 U22250 ( .A1(n19874), .A2(n20092), .ZN(n15383) );
  NAND2_X1 U22251 ( .A1(n16957), .A2(n28763), .ZN(n17038) );
  OAI21_X1 U22252 ( .A1(n20065), .A2(n16630), .B(n10413), .ZN(n15311) );
  NOR3_X1 U22255 ( .A1(n834), .A2(n25865), .A3(n29063), .ZN(n14872) );
  NAND2_X1 U22258 ( .A1(n23889), .A2(n23888), .ZN(n17257) );
  BUF_X2 U22267 ( .I(n19618), .Z(n20154) );
  OAI21_X1 U22271 ( .A1(n16694), .A2(n13852), .B(n19863), .ZN(n17061) );
  NAND2_X1 U22272 ( .A1(n14960), .A2(n13627), .ZN(n13935) );
  NAND2_X1 U22273 ( .A1(n8919), .A2(n14845), .ZN(n15699) );
  NAND2_X1 U22275 ( .A1(n953), .A2(n17649), .ZN(n17736) );
  NAND2_X1 U22276 ( .A1(n21713), .A2(n727), .ZN(n21478) );
  NOR2_X1 U22283 ( .A1(n22468), .A2(n15089), .ZN(n15939) );
  NAND2_X1 U22286 ( .A1(n23822), .A2(n23942), .ZN(n13668) );
  INV_X1 U22289 ( .I(n23933), .ZN(n13102) );
  OAI21_X1 U22290 ( .A1(n28010), .A2(n4194), .B(n16181), .ZN(n13111) );
  NAND2_X1 U22291 ( .A1(n338), .A2(n16987), .ZN(n21844) );
  NOR2_X2 U22292 ( .A1(n13265), .A2(n20934), .ZN(n13114) );
  OAI21_X1 U22293 ( .A1(n17644), .A2(n29523), .B(n13115), .ZN(n21591) );
  XOR2_X1 U22298 ( .A1(n600), .A2(n20700), .Z(n13122) );
  XNOR2_X1 U22299 ( .A1(n17871), .A2(n30322), .ZN(n13123) );
  NAND2_X1 U22300 ( .A1(n29270), .A2(n13125), .ZN(n23642) );
  AOI21_X1 U22301 ( .A1(n16431), .A2(n13125), .B(n354), .ZN(n16281) );
  NAND2_X1 U22306 ( .A1(n12871), .A2(n17074), .ZN(n24606) );
  NOR2_X2 U22309 ( .A1(n17935), .A2(n16818), .ZN(n23003) );
  XOR2_X1 U22317 ( .A1(n20753), .A2(n13179), .Z(n13178) );
  XOR2_X1 U22320 ( .A1(n20786), .A2(n16655), .Z(n13181) );
  MUX2_X1 U22324 ( .I0(n13186), .I1(n13185), .S(n900), .Z(n17249) );
  XOR2_X1 U22330 ( .A1(n30273), .A2(n13209), .Z(n13208) );
  XOR2_X1 U22331 ( .A1(n23464), .A2(n23414), .Z(n13214) );
  XOR2_X1 U22334 ( .A1(n2073), .A2(n16555), .Z(n13222) );
  XOR2_X1 U22338 ( .A1(n23497), .A2(n23180), .Z(n13234) );
  XOR2_X1 U22340 ( .A1(n23181), .A2(n17934), .Z(n13235) );
  MUX2_X1 U22346 ( .I0(n14756), .I1(n842), .S(n299), .Z(n13261) );
  XOR2_X1 U22358 ( .A1(n16175), .A2(n17998), .Z(n13293) );
  XOR2_X1 U22359 ( .A1(n20972), .A2(n20971), .Z(n13294) );
  NAND2_X2 U22361 ( .A1(n14521), .A2(n23959), .ZN(n16868) );
  XOR2_X1 U22362 ( .A1(n27151), .A2(n2864), .Z(n13299) );
  NAND2_X2 U22363 ( .A1(n13302), .A2(n13301), .ZN(n14980) );
  XOR2_X1 U22364 ( .A1(n33150), .A2(n16612), .Z(n13303) );
  NOR2_X1 U22369 ( .A1(n9191), .A2(n30313), .ZN(n13312) );
  NAND3_X1 U22370 ( .A1(n17985), .A2(n30313), .A3(n18035), .ZN(n13313) );
  INV_X2 U22372 ( .I(n18110), .ZN(n13319) );
  NAND2_X1 U22374 ( .A1(n10700), .A2(n25968), .ZN(n17510) );
  NAND2_X1 U22376 ( .A1(n13329), .A2(n8787), .ZN(n13328) );
  NAND3_X1 U22377 ( .A1(n16066), .A2(n27500), .A3(n794), .ZN(n23609) );
  XOR2_X1 U22380 ( .A1(n13336), .A2(n21028), .Z(n17440) );
  AOI21_X2 U22384 ( .A1(n23222), .A2(n23223), .B(n23221), .ZN(n24276) );
  XOR2_X1 U22391 ( .A1(n19445), .A2(n15117), .Z(n19373) );
  XOR2_X1 U22393 ( .A1(n20960), .A2(n13357), .Z(n14930) );
  XOR2_X1 U22403 ( .A1(n6462), .A2(n15779), .Z(n15778) );
  XOR2_X1 U22404 ( .A1(n13375), .A2(n13372), .Z(n17768) );
  XOR2_X1 U22405 ( .A1(n13373), .A2(n13374), .Z(n13372) );
  XOR2_X1 U22406 ( .A1(n15183), .A2(n16674), .Z(n13373) );
  XOR2_X1 U22407 ( .A1(n13638), .A2(n27613), .Z(n13374) );
  XOR2_X1 U22409 ( .A1(n16053), .A2(n25195), .Z(n13388) );
  XOR2_X1 U22410 ( .A1(n28262), .A2(n13394), .Z(n13393) );
  XOR2_X1 U22412 ( .A1(n13405), .A2(n13404), .Z(n13403) );
  XOR2_X1 U22413 ( .A1(n20996), .A2(n14858), .Z(n13405) );
  INV_X1 U22414 ( .I(n13407), .ZN(n21416) );
  INV_X2 U22415 ( .I(n12317), .ZN(n18785) );
  XOR2_X1 U22419 ( .A1(n24403), .A2(n13419), .Z(n23551) );
  NOR2_X1 U22420 ( .A1(n17339), .A2(n27033), .ZN(n19126) );
  NOR2_X1 U22421 ( .A1(n17339), .A2(n32414), .ZN(n18985) );
  NOR2_X1 U22423 ( .A1(n17382), .A2(n15719), .ZN(n17770) );
  NOR2_X1 U22424 ( .A1(n17382), .A2(n14454), .ZN(n13429) );
  XOR2_X1 U22426 ( .A1(n13439), .A2(n13441), .Z(n16777) );
  XOR2_X1 U22427 ( .A1(n19546), .A2(n13440), .Z(n13439) );
  XOR2_X1 U22428 ( .A1(n13826), .A2(n25064), .Z(n13440) );
  XOR2_X1 U22430 ( .A1(n19463), .A2(n19772), .Z(n19545) );
  XOR2_X1 U22439 ( .A1(n13454), .A2(n13453), .Z(n13452) );
  XOR2_X1 U22440 ( .A1(n33468), .A2(n4295), .Z(n13454) );
  OR2_X1 U22442 ( .A1(n23975), .A2(n23976), .Z(n13459) );
  NOR2_X1 U22444 ( .A1(n8320), .A2(n13483), .ZN(n25544) );
  NAND3_X1 U22446 ( .A1(n24059), .A2(n14501), .A3(n13394), .ZN(n13467) );
  INV_X1 U22447 ( .I(n13469), .ZN(n13468) );
  AOI21_X1 U22448 ( .A1(n14501), .A2(n24059), .B(n13394), .ZN(n13469) );
  XOR2_X1 U22452 ( .A1(n16060), .A2(n25648), .Z(n21938) );
  NAND2_X1 U22457 ( .A1(n950), .A2(n19116), .ZN(n13494) );
  XOR2_X1 U22458 ( .A1(n13498), .A2(n23450), .Z(n13497) );
  XOR2_X1 U22462 ( .A1(n22264), .A2(n25218), .Z(n22265) );
  XOR2_X1 U22463 ( .A1(n22264), .A2(n25693), .Z(n14979) );
  XOR2_X1 U22470 ( .A1(n23300), .A2(n23299), .Z(n13517) );
  NAND2_X2 U22471 ( .A1(n22054), .A2(n22053), .ZN(n23300) );
  XOR2_X1 U22474 ( .A1(n13527), .A2(n13394), .Z(Ciphertext[124]) );
  AOI21_X1 U22475 ( .A1(n25556), .A2(n33414), .B(n16853), .ZN(n13528) );
  INV_X1 U22476 ( .I(n25542), .ZN(n25556) );
  XOR2_X1 U22477 ( .A1(n30331), .A2(n14526), .Z(n13529) );
  XOR2_X1 U22479 ( .A1(n32871), .A2(n13545), .Z(n24637) );
  XOR2_X1 U22480 ( .A1(n24421), .A2(n13545), .Z(n24415) );
  NOR2_X1 U22483 ( .A1(n17328), .A2(n20563), .ZN(n20564) );
  NAND2_X1 U22487 ( .A1(n13558), .A2(n22971), .ZN(n22972) );
  OAI21_X1 U22489 ( .A1(n2635), .A2(n13558), .B(n13191), .ZN(n15753) );
  NAND2_X1 U22490 ( .A1(n23106), .A2(n13558), .ZN(n22804) );
  XOR2_X1 U22493 ( .A1(n32084), .A2(n13564), .Z(n22178) );
  XOR2_X1 U22495 ( .A1(n13586), .A2(n24532), .Z(n17309) );
  XOR2_X1 U22496 ( .A1(n30795), .A2(n13586), .Z(n24828) );
  XOR2_X1 U22497 ( .A1(n25969), .A2(n24869), .Z(n13590) );
  NOR2_X1 U22498 ( .A1(n11198), .A2(n13591), .ZN(n17155) );
  XOR2_X1 U22500 ( .A1(n24830), .A2(n25506), .Z(n13595) );
  XOR2_X1 U22501 ( .A1(n15588), .A2(n24815), .Z(n13596) );
  XOR2_X1 U22502 ( .A1(n24513), .A2(n24512), .Z(n24815) );
  XOR2_X1 U22506 ( .A1(n13606), .A2(n16613), .Z(n20864) );
  XOR2_X1 U22507 ( .A1(n13606), .A2(n1431), .Z(n15652) );
  NAND2_X2 U22508 ( .A1(n13609), .A2(n13608), .ZN(n20158) );
  NOR2_X1 U22511 ( .A1(n24965), .A2(n13627), .ZN(n17331) );
  INV_X2 U22512 ( .I(n15514), .ZN(n14133) );
  NAND2_X1 U22514 ( .A1(n19824), .A2(n1165), .ZN(n19825) );
  XOR2_X1 U22519 ( .A1(Plaintext[117]), .A2(Key[117]), .Z(n13719) );
  NOR2_X1 U22522 ( .A1(n13319), .A2(n21167), .ZN(n13680) );
  XOR2_X1 U22523 ( .A1(n13681), .A2(n1434), .Z(n15793) );
  XOR2_X1 U22524 ( .A1(n32367), .A2(n25864), .Z(n13682) );
  XOR2_X1 U22529 ( .A1(n19384), .A2(n17091), .Z(n13689) );
  NAND2_X1 U22542 ( .A1(n30682), .A2(n19048), .ZN(n19016) );
  AOI21_X1 U22544 ( .A1(n13736), .A2(n24970), .B(n13934), .ZN(n13735) );
  NAND2_X1 U22545 ( .A1(n32493), .A2(n992), .ZN(n22436) );
  XOR2_X1 U22546 ( .A1(n11862), .A2(n25619), .Z(n13740) );
  XOR2_X1 U22547 ( .A1(n968), .A2(n15161), .Z(n13742) );
  XOR2_X1 U22550 ( .A1(n24770), .A2(n24993), .Z(n13745) );
  OAI21_X1 U22556 ( .A1(n31921), .A2(n29539), .B(n13763), .ZN(n16188) );
  NAND3_X1 U22557 ( .A1(n17177), .A2(n19866), .A3(n1395), .ZN(n13765) );
  INV_X1 U22558 ( .I(n13767), .ZN(n13766) );
  AOI21_X1 U22559 ( .A1(n17177), .A2(n19866), .B(n1395), .ZN(n13767) );
  AND2_X1 U22562 ( .A1(n13785), .A2(n13537), .Z(n13784) );
  XOR2_X1 U22566 ( .A1(n24783), .A2(n24668), .Z(n13794) );
  INV_X2 U22568 ( .I(n17047), .ZN(n25334) );
  MUX2_X1 U22569 ( .I0(n33110), .I1(n33583), .S(n31807), .Z(n23222) );
  NOR2_X1 U22571 ( .A1(n31716), .A2(n17189), .ZN(n13809) );
  XOR2_X1 U22572 ( .A1(n32753), .A2(n26931), .Z(n22131) );
  MUX2_X1 U22573 ( .I0(n23624), .I1(n23625), .S(n791), .Z(n23627) );
  XOR2_X1 U22574 ( .A1(n17188), .A2(n24964), .Z(n13812) );
  XOR2_X1 U22575 ( .A1(n8347), .A2(n19718), .Z(n15557) );
  XOR2_X1 U22576 ( .A1(n13817), .A2(n19411), .Z(n15679) );
  XOR2_X1 U22577 ( .A1(n32271), .A2(n13826), .Z(n19430) );
  INV_X1 U22586 ( .I(n15139), .ZN(n13845) );
  XOR2_X1 U22589 ( .A1(n19405), .A2(n13854), .Z(n13853) );
  XNOR2_X1 U22590 ( .A1(n19658), .A2(n19461), .ZN(n19405) );
  XOR2_X1 U22591 ( .A1(n19574), .A2(n19480), .Z(n13855) );
  XOR2_X1 U22592 ( .A1(n16727), .A2(n19353), .Z(n19480) );
  OR2_X1 U22596 ( .A1(n22721), .A2(n28849), .Z(n13861) );
  OAI22_X1 U22599 ( .A1(n15655), .A2(n920), .B1(n27024), .B2(n13872), .ZN(
        n21275) );
  XOR2_X1 U22601 ( .A1(n16891), .A2(n13877), .Z(n13876) );
  XOR2_X1 U22602 ( .A1(n27423), .A2(n25929), .Z(n13877) );
  AND2_X1 U22604 ( .A1(n25542), .A2(n31236), .Z(n13883) );
  XOR2_X1 U22607 ( .A1(n5348), .A2(n20825), .Z(n20799) );
  XOR2_X1 U22608 ( .A1(n20764), .A2(n13887), .Z(n13886) );
  XOR2_X1 U22609 ( .A1(n20843), .A2(n25074), .Z(n13887) );
  XOR2_X1 U22610 ( .A1(Plaintext[63]), .A2(Key[63]), .Z(n16596) );
  INV_X1 U22611 ( .I(n13895), .ZN(n13893) );
  XOR2_X1 U22613 ( .A1(n28687), .A2(n25190), .Z(n13898) );
  XOR2_X1 U22615 ( .A1(n21009), .A2(n20924), .Z(n13901) );
  XOR2_X1 U22616 ( .A1(n13902), .A2(n12797), .Z(Ciphertext[185]) );
  XOR2_X1 U22618 ( .A1(n27252), .A2(n25182), .Z(n13907) );
  XOR2_X1 U22619 ( .A1(n14908), .A2(n4157), .Z(n13909) );
  XOR2_X1 U22623 ( .A1(n27481), .A2(n16322), .Z(n13927) );
  XOR2_X1 U22624 ( .A1(n23271), .A2(n23291), .Z(n13928) );
  INV_X2 U22627 ( .I(n13931), .ZN(n23855) );
  INV_X1 U22631 ( .I(n13944), .ZN(n15946) );
  XOR2_X1 U22633 ( .A1(n22108), .A2(n25224), .Z(n13956) );
  NAND2_X1 U22634 ( .A1(n8371), .A2(n14334), .ZN(n19811) );
  NOR2_X1 U22639 ( .A1(n14392), .A2(n22791), .ZN(n22759) );
  NOR3_X1 U22644 ( .A1(n17066), .A2(n17065), .A3(n17068), .ZN(n17067) );
  NAND3_X1 U22646 ( .A1(n25613), .A2(n11931), .A3(n9982), .ZN(n25609) );
  NAND3_X1 U22650 ( .A1(n16783), .A2(n25561), .A3(n16704), .ZN(n13979) );
  XOR2_X1 U22655 ( .A1(n22202), .A2(n22146), .Z(n15686) );
  XOR2_X1 U22656 ( .A1(n22284), .A2(n18113), .Z(n15548) );
  NOR2_X1 U22659 ( .A1(n25254), .A2(n17273), .ZN(n15094) );
  NAND2_X1 U22664 ( .A1(n21866), .A2(n21736), .ZN(n16235) );
  OAI21_X1 U22665 ( .A1(n21189), .A2(n21321), .B(n14023), .ZN(n14022) );
  OAI21_X1 U22666 ( .A1(n25808), .A2(n25811), .B(n14009), .ZN(n25810) );
  OR2_X1 U22674 ( .A1(n20099), .A2(n19990), .Z(n14019) );
  XOR2_X1 U22675 ( .A1(n19596), .A2(n19595), .Z(n19601) );
  NAND2_X2 U22678 ( .A1(n21191), .A2(n14022), .ZN(n21872) );
  XOR2_X1 U22680 ( .A1(n14908), .A2(n16110), .Z(n14916) );
  XOR2_X1 U22688 ( .A1(n22169), .A2(n21924), .Z(n17919) );
  NAND3_X1 U22691 ( .A1(n25773), .A2(n25788), .A3(n25796), .ZN(n25768) );
  NOR2_X1 U22693 ( .A1(n10364), .A2(n18662), .ZN(n17910) );
  XOR2_X1 U22696 ( .A1(n14043), .A2(n14494), .Z(n17518) );
  XOR2_X1 U22697 ( .A1(n618), .A2(n21661), .Z(n14043) );
  OR2_X1 U22699 ( .A1(n30949), .A2(n23938), .Z(n15238) );
  XOR2_X1 U22700 ( .A1(n15612), .A2(n23374), .Z(n23936) );
  INV_X2 U22701 ( .I(n15613), .ZN(n23533) );
  NAND2_X1 U22703 ( .A1(n20609), .A2(n20608), .ZN(n14050) );
  NAND2_X1 U22704 ( .A1(n20610), .A2(n33397), .ZN(n14051) );
  XOR2_X1 U22705 ( .A1(n28262), .A2(n2616), .Z(n20639) );
  XOR2_X1 U22706 ( .A1(n14053), .A2(n4047), .Z(n15099) );
  NAND2_X1 U22708 ( .A1(n828), .A2(n18774), .ZN(n14056) );
  XOR2_X1 U22713 ( .A1(n14070), .A2(n25274), .Z(Ciphertext[86]) );
  AND2_X1 U22721 ( .A1(n19243), .A2(n877), .Z(n14699) );
  NAND2_X1 U22723 ( .A1(n16156), .A2(n11774), .ZN(n14100) );
  XOR2_X1 U22725 ( .A1(n16128), .A2(n24696), .Z(n24697) );
  INV_X2 U22729 ( .I(n18090), .ZN(n20113) );
  XNOR2_X1 U22733 ( .A1(n15787), .A2(n19654), .ZN(n18051) );
  OAI21_X1 U22738 ( .A1(n29815), .A2(n16872), .B(n16871), .ZN(n16870) );
  OR3_X1 U22739 ( .A1(n20335), .A2(n30130), .A3(n20158), .Z(n20159) );
  XOR2_X1 U22741 ( .A1(n14391), .A2(n19617), .Z(n19618) );
  XOR2_X1 U22742 ( .A1(n22137), .A2(n22138), .Z(n22140) );
  AOI21_X1 U22744 ( .A1(n22338), .A2(n906), .B(n22645), .ZN(n14145) );
  XOR2_X1 U22746 ( .A1(n29876), .A2(n3727), .Z(n14146) );
  NAND2_X1 U22748 ( .A1(n1385), .A2(n18990), .ZN(n14148) );
  NAND2_X1 U22749 ( .A1(n25471), .A2(n25472), .ZN(n14149) );
  INV_X1 U22750 ( .I(n25057), .ZN(n25045) );
  OR2_X1 U22751 ( .A1(n25058), .A2(n25057), .Z(n25043) );
  AND2_X1 U22753 ( .A1(n2061), .A2(n6533), .Z(n14150) );
  XOR2_X1 U22754 ( .A1(n17309), .A2(n24355), .Z(n17308) );
  XOR2_X1 U22756 ( .A1(n14370), .A2(n14154), .Z(n23352) );
  NAND2_X2 U22760 ( .A1(n14657), .A2(n14660), .ZN(n19255) );
  NAND2_X1 U22762 ( .A1(n28070), .A2(n25062), .ZN(n17741) );
  XOR2_X1 U22764 ( .A1(n20912), .A2(n20914), .Z(n15035) );
  OR2_X1 U22766 ( .A1(n5394), .A2(n20940), .Z(n15925) );
  NAND3_X1 U22769 ( .A1(n17403), .A2(n15134), .A3(n17402), .ZN(n17401) );
  NOR2_X2 U22771 ( .A1(n19912), .A2(n19913), .ZN(n14187) );
  INV_X2 U22774 ( .I(n14190), .ZN(n23871) );
  NAND2_X1 U22776 ( .A1(n23876), .A2(n801), .ZN(n16325) );
  NOR2_X1 U22777 ( .A1(n24137), .A2(n15011), .ZN(n14196) );
  XOR2_X1 U22782 ( .A1(n24806), .A2(n14203), .Z(n14202) );
  XOR2_X1 U22783 ( .A1(n24764), .A2(n26000), .Z(n14203) );
  XOR2_X1 U22786 ( .A1(n19561), .A2(n25993), .Z(n14211) );
  INV_X2 U22795 ( .I(n18763), .ZN(n18768) );
  XOR2_X1 U22797 ( .A1(n24648), .A2(n14578), .Z(n14239) );
  XOR2_X1 U22798 ( .A1(n29190), .A2(n19718), .Z(n14242) );
  XOR2_X1 U22799 ( .A1(n23376), .A2(n16373), .Z(n23289) );
  NOR2_X1 U22804 ( .A1(n14438), .A2(n32253), .ZN(n14437) );
  XOR2_X1 U22807 ( .A1(n28864), .A2(n20892), .Z(n15525) );
  NAND3_X1 U22808 ( .A1(n15073), .A2(n15074), .A3(n17986), .ZN(n14257) );
  INV_X1 U22809 ( .I(n14259), .ZN(n14258) );
  AND2_X1 U22813 ( .A1(n1218), .A2(n25183), .Z(n14276) );
  XOR2_X1 U22814 ( .A1(n24762), .A2(n14279), .Z(n14277) );
  XOR2_X1 U22816 ( .A1(n33447), .A2(n24759), .Z(n14279) );
  XOR2_X1 U22818 ( .A1(n22180), .A2(n14299), .Z(n14298) );
  XOR2_X1 U22820 ( .A1(n14316), .A2(n14315), .Z(n19532) );
  NAND2_X1 U22824 ( .A1(n19078), .A2(n31254), .ZN(n19079) );
  XOR2_X1 U22825 ( .A1(n5772), .A2(n24962), .Z(n21022) );
  XOR2_X1 U22826 ( .A1(n5772), .A2(n25519), .Z(n20914) );
  XOR2_X1 U22827 ( .A1(n5772), .A2(n25827), .Z(n20166) );
  XOR2_X1 U22833 ( .A1(n14349), .A2(n23185), .Z(n14348) );
  XOR2_X1 U22834 ( .A1(n29462), .A2(n33293), .Z(n14349) );
  XOR2_X1 U22839 ( .A1(n14364), .A2(n14361), .Z(n15294) );
  XOR2_X1 U22840 ( .A1(n14362), .A2(n14363), .Z(n14361) );
  XOR2_X1 U22842 ( .A1(n24685), .A2(n24443), .Z(n14364) );
  OR2_X1 U22843 ( .A1(n20434), .A2(n20432), .Z(n14368) );
  XOR2_X1 U22844 ( .A1(n19624), .A2(n25549), .Z(n17009) );
  XOR2_X1 U22848 ( .A1(n33574), .A2(n17301), .Z(n14385) );
  NAND2_X1 U22849 ( .A1(n16554), .A2(n24219), .ZN(n14444) );
  NAND2_X1 U22850 ( .A1(n16554), .A2(n24218), .ZN(n23602) );
  INV_X2 U22854 ( .I(n14409), .ZN(n16249) );
  INV_X2 U22856 ( .I(n18429), .ZN(n18822) );
  NOR2_X1 U22857 ( .A1(n1245), .A2(n29634), .ZN(n16800) );
  XOR2_X1 U22858 ( .A1(n21726), .A2(n25079), .Z(n14416) );
  XOR2_X1 U22859 ( .A1(n22294), .A2(n22064), .Z(n14422) );
  XOR2_X1 U22860 ( .A1(n20225), .A2(n20226), .Z(n14429) );
  XOR2_X1 U22864 ( .A1(n27126), .A2(n13091), .Z(n14435) );
  XOR2_X1 U22867 ( .A1(n23488), .A2(n29299), .Z(n14442) );
  NAND3_X1 U22869 ( .A1(n30279), .A2(n714), .A3(n3232), .ZN(n14607) );
  NAND2_X1 U22875 ( .A1(n14451), .A2(n14450), .ZN(n14449) );
  NAND2_X2 U22877 ( .A1(n23571), .A2(n23572), .ZN(n15663) );
  NAND3_X2 U22882 ( .A1(n14472), .A2(n14471), .A3(n14470), .ZN(n14682) );
  OR2_X1 U22884 ( .A1(n14683), .A2(n1355), .Z(n14472) );
  NAND2_X1 U22885 ( .A1(n23643), .A2(n3760), .ZN(n23644) );
  NAND2_X1 U22886 ( .A1(n14478), .A2(n17163), .ZN(n21979) );
  XOR2_X1 U22890 ( .A1(n1261), .A2(n23203), .Z(n14481) );
  XOR2_X1 U22891 ( .A1(n23503), .A2(n16523), .Z(n14492) );
  XOR2_X1 U22893 ( .A1(n22197), .A2(n22239), .Z(n21813) );
  XOR2_X1 U22895 ( .A1(n14506), .A2(n14504), .Z(n21869) );
  XOR2_X1 U22896 ( .A1(n21838), .A2(n14505), .Z(n14504) );
  XOR2_X1 U22897 ( .A1(n22243), .A2(n27180), .Z(n14505) );
  XOR2_X1 U22898 ( .A1(n33969), .A2(n31513), .Z(n14507) );
  NAND2_X1 U22900 ( .A1(n25338), .A2(n14509), .ZN(n25341) );
  XOR2_X1 U22903 ( .A1(n14517), .A2(n14519), .Z(n16845) );
  XOR2_X1 U22904 ( .A1(n20827), .A2(n14930), .Z(n14519) );
  INV_X2 U22910 ( .I(n14534), .ZN(n14556) );
  XOR2_X1 U22912 ( .A1(n29235), .A2(n24943), .Z(n23316) );
  XOR2_X1 U22918 ( .A1(n24809), .A2(n24417), .Z(n14578) );
  XOR2_X1 U22920 ( .A1(n23219), .A2(n14586), .Z(n14580) );
  XOR2_X1 U22921 ( .A1(n14584), .A2(n14582), .Z(n14581) );
  XOR2_X1 U22922 ( .A1(n23266), .A2(n25880), .Z(n14586) );
  XOR2_X1 U22923 ( .A1(n15374), .A2(n15372), .Z(n15399) );
  XOR2_X1 U22926 ( .A1(n28730), .A2(n1407), .Z(n15900) );
  INV_X1 U22927 ( .I(n14717), .ZN(n17225) );
  NAND2_X1 U22929 ( .A1(n24154), .A2(n31883), .ZN(n23117) );
  XOR2_X1 U22931 ( .A1(n20917), .A2(n16642), .Z(n14646) );
  AND2_X1 U22933 ( .A1(n18638), .A2(n18539), .Z(n14653) );
  INV_X2 U22934 ( .I(n14661), .ZN(n16489) );
  NAND2_X1 U22937 ( .A1(n31907), .A2(n14365), .ZN(n20508) );
  XOR2_X1 U22944 ( .A1(n14682), .A2(n16454), .Z(n20810) );
  XOR2_X1 U22945 ( .A1(n22123), .A2(n21952), .Z(n14684) );
  XOR2_X1 U22947 ( .A1(n21998), .A2(n21953), .Z(n14685) );
  XOR2_X1 U22954 ( .A1(n20794), .A2(n20793), .Z(n14701) );
  NAND2_X2 U22955 ( .A1(n18225), .A2(n18224), .ZN(n16093) );
  NOR2_X1 U22961 ( .A1(n16627), .A2(n11895), .ZN(n14713) );
  XOR2_X1 U22962 ( .A1(n12459), .A2(n7717), .Z(n14716) );
  XOR2_X1 U22965 ( .A1(n8491), .A2(n1396), .Z(n15368) );
  OAI21_X1 U22966 ( .A1(n20112), .A2(n20045), .B(n16812), .ZN(n17609) );
  XOR2_X1 U22967 ( .A1(n23179), .A2(n24763), .Z(n24634) );
  XOR2_X1 U22968 ( .A1(n19537), .A2(n32046), .Z(n14744) );
  XOR2_X1 U22970 ( .A1(n23355), .A2(n7045), .Z(n14748) );
  XOR2_X1 U22973 ( .A1(n22196), .A2(n16631), .Z(n14754) );
  XOR2_X1 U22979 ( .A1(n23330), .A2(n14782), .Z(n14781) );
  XOR2_X1 U22980 ( .A1(n29299), .A2(n1410), .Z(n14782) );
  XOR2_X1 U22981 ( .A1(n23507), .A2(n23209), .Z(n23330) );
  XOR2_X1 U22982 ( .A1(n20776), .A2(n25319), .Z(n14784) );
  XOR2_X1 U22984 ( .A1(n22201), .A2(n16578), .Z(n14787) );
  XOR2_X1 U22985 ( .A1(n23437), .A2(n23329), .Z(n14791) );
  NOR2_X1 U22989 ( .A1(n32590), .A2(n14805), .ZN(n16532) );
  XOR2_X1 U22991 ( .A1(n21017), .A2(n20915), .Z(n14809) );
  INV_X2 U22992 ( .I(n14814), .ZN(n14815) );
  XOR2_X1 U22995 ( .A1(n22139), .A2(n4342), .Z(n16036) );
  XOR2_X1 U22996 ( .A1(n14820), .A2(n15702), .Z(n15701) );
  NAND2_X1 U22998 ( .A1(n7486), .A2(n20555), .ZN(n20297) );
  XOR2_X1 U23002 ( .A1(Plaintext[95]), .A2(Key[95]), .Z(n15955) );
  XOR2_X1 U23005 ( .A1(n21913), .A2(n910), .Z(n14833) );
  AND2_X1 U23007 ( .A1(n19936), .A2(n14834), .Z(n15382) );
  NAND3_X1 U23010 ( .A1(n2551), .A2(n28395), .A3(n1647), .ZN(n21724) );
  XOR2_X1 U23012 ( .A1(n24504), .A2(n477), .Z(n14842) );
  XOR2_X1 U23014 ( .A1(n22238), .A2(n1404), .Z(n21930) );
  XOR2_X1 U23015 ( .A1(n22238), .A2(n16438), .Z(n22041) );
  NOR2_X1 U23016 ( .A1(n14863), .A2(n20494), .ZN(n19804) );
  NOR2_X1 U23018 ( .A1(n26585), .A2(n14863), .ZN(n20437) );
  NOR2_X2 U23020 ( .A1(n14866), .A2(n16469), .ZN(n14865) );
  XOR2_X1 U23022 ( .A1(n27179), .A2(n16550), .Z(n15049) );
  XOR2_X1 U23027 ( .A1(n24425), .A2(n14884), .Z(n14883) );
  XOR2_X1 U23028 ( .A1(n24813), .A2(n14885), .Z(n14884) );
  XOR2_X1 U23029 ( .A1(n14887), .A2(n17643), .Z(n16938) );
  XOR2_X1 U23030 ( .A1(n11668), .A2(n25126), .Z(n23495) );
  OAI21_X1 U23032 ( .A1(n14893), .A2(n14892), .B(n100), .ZN(n17810) );
  OR2_X1 U23033 ( .A1(n21440), .A2(n8115), .Z(n14896) );
  XOR2_X1 U23034 ( .A1(Key[105]), .A2(Plaintext[105]), .Z(n14898) );
  INV_X2 U23035 ( .I(n14898), .ZN(n16732) );
  XOR2_X1 U23036 ( .A1(n14902), .A2(n21112), .Z(n14901) );
  NOR2_X1 U23038 ( .A1(n25863), .A2(n14915), .ZN(n25861) );
  XOR2_X1 U23044 ( .A1(n24790), .A2(n25161), .Z(n14920) );
  XOR2_X1 U23046 ( .A1(n24816), .A2(n28898), .Z(n24818) );
  XOR2_X1 U23049 ( .A1(n24473), .A2(n15674), .Z(n14935) );
  XOR2_X1 U23050 ( .A1(n17301), .A2(n14938), .Z(n14937) );
  XOR2_X1 U23051 ( .A1(n2896), .A2(n25324), .Z(n17187) );
  NOR2_X1 U23060 ( .A1(n19874), .A2(n14976), .ZN(n16065) );
  NAND2_X1 U23065 ( .A1(n13300), .A2(n1154), .ZN(n20178) );
  XOR2_X1 U23069 ( .A1(n19733), .A2(n19467), .Z(n14985) );
  XOR2_X1 U23071 ( .A1(n12594), .A2(n17063), .Z(n16344) );
  XOR2_X1 U23072 ( .A1(n12594), .A2(n25161), .Z(n22233) );
  XOR2_X1 U23073 ( .A1(n22251), .A2(n12594), .Z(n22018) );
  XOR2_X1 U23074 ( .A1(n23506), .A2(n23407), .Z(n22387) );
  XOR2_X1 U23075 ( .A1(n11370), .A2(n25126), .Z(n24476) );
  XOR2_X1 U23076 ( .A1(n156), .A2(n28411), .Z(n14994) );
  NAND2_X1 U23078 ( .A1(n1350), .A2(n15005), .ZN(n20420) );
  NAND2_X1 U23079 ( .A1(n20419), .A2(n1352), .ZN(n15006) );
  NOR2_X1 U23083 ( .A1(n15027), .A2(n20463), .ZN(n20352) );
  XOR2_X1 U23086 ( .A1(n19423), .A2(n24953), .Z(n15031) );
  XOR2_X1 U23088 ( .A1(n20911), .A2(n15037), .Z(n15036) );
  XOR2_X1 U23089 ( .A1(n3799), .A2(n348), .Z(n15037) );
  XOR2_X1 U23090 ( .A1(n20925), .A2(n591), .Z(n15048) );
  XOR2_X1 U23094 ( .A1(n29644), .A2(n16674), .Z(n19669) );
  XOR2_X1 U23099 ( .A1(n31584), .A2(n20872), .Z(n15083) );
  XOR2_X1 U23102 ( .A1(n19634), .A2(n19633), .Z(n19635) );
  XOR2_X1 U23104 ( .A1(n23138), .A2(n15099), .Z(n16283) );
  OR2_X1 U23105 ( .A1(n21963), .A2(n15103), .Z(n22418) );
  XOR2_X1 U23107 ( .A1(n15106), .A2(n16730), .Z(n16711) );
  OR2_X1 U23109 ( .A1(n19947), .A2(n19857), .Z(n15111) );
  INV_X2 U23110 ( .I(n15115), .ZN(n17598) );
  XOR2_X1 U23111 ( .A1(Key[71]), .A2(Plaintext[71]), .Z(n15115) );
  XOR2_X1 U23113 ( .A1(n438), .A2(n16373), .Z(n15121) );
  INV_X1 U23115 ( .I(n16676), .ZN(n23612) );
  NAND2_X1 U23117 ( .A1(n15124), .A2(n25251), .ZN(n16582) );
  NAND2_X1 U23119 ( .A1(n21719), .A2(n17227), .ZN(n15127) );
  INV_X1 U23124 ( .I(Plaintext[101]), .ZN(n17548) );
  NAND2_X2 U23128 ( .A1(n15140), .A2(n15196), .ZN(n19115) );
  XOR2_X1 U23136 ( .A1(n15153), .A2(n16753), .Z(n16756) );
  NAND2_X1 U23138 ( .A1(n25527), .A2(n28096), .ZN(n15156) );
  NAND2_X1 U23142 ( .A1(n20626), .A2(n14005), .ZN(n15173) );
  NAND2_X1 U23147 ( .A1(n21707), .A2(n21512), .ZN(n21482) );
  INV_X1 U23150 ( .I(n21071), .ZN(n21427) );
  INV_X1 U23151 ( .I(n16558), .ZN(n22635) );
  XOR2_X1 U23154 ( .A1(n1130), .A2(n21938), .Z(n21940) );
  NAND2_X2 U23156 ( .A1(n18143), .A2(n22499), .ZN(n22955) );
  XOR2_X1 U23158 ( .A1(Plaintext[87]), .A2(Key[87]), .Z(n15194) );
  BUF_X4 U23163 ( .I(n24459), .Z(n25582) );
  XOR2_X1 U23164 ( .A1(n15205), .A2(n15701), .Z(n20015) );
  XOR2_X1 U23166 ( .A1(Plaintext[13]), .A2(Key[13]), .Z(n16914) );
  AND2_X1 U23167 ( .A1(n22984), .A2(n22985), .Z(n15208) );
  XOR2_X1 U23169 ( .A1(n16586), .A2(n11889), .Z(n19502) );
  INV_X1 U23173 ( .I(Key[118]), .ZN(n16378) );
  NAND2_X1 U23175 ( .A1(n20205), .A2(n8206), .ZN(n18171) );
  INV_X2 U23177 ( .I(n15229), .ZN(n18098) );
  NOR3_X1 U23178 ( .A1(n26350), .A2(n10700), .A3(n14312), .ZN(n18716) );
  NAND2_X1 U23179 ( .A1(n21791), .A2(n21790), .ZN(n21796) );
  NOR2_X1 U23181 ( .A1(n24610), .A2(n680), .ZN(n15231) );
  XOR2_X1 U23182 ( .A1(Plaintext[161]), .A2(Key[161]), .Z(n15347) );
  NAND2_X2 U23183 ( .A1(n17196), .A2(n17195), .ZN(n25916) );
  INV_X2 U23189 ( .I(n15235), .ZN(n16704) );
  NOR2_X1 U23190 ( .A1(n15722), .A2(n15238), .ZN(n17180) );
  MUX2_X1 U23191 ( .I0(n23549), .I1(n23548), .S(n16066), .Z(n23550) );
  XOR2_X1 U23192 ( .A1(n23512), .A2(n6901), .Z(n15307) );
  XOR2_X1 U23193 ( .A1(Key[107]), .A2(Plaintext[107]), .Z(n15240) );
  AND3_X1 U23199 ( .A1(n21181), .A2(n21182), .A3(n4076), .Z(n16282) );
  XOR2_X1 U23201 ( .A1(n17141), .A2(n12101), .Z(n17140) );
  INV_X1 U23203 ( .I(Plaintext[124]), .ZN(n17622) );
  XOR2_X1 U23204 ( .A1(n19580), .A2(n27137), .Z(n19582) );
  OAI21_X2 U23207 ( .A1(n19623), .A2(n19622), .B(n19621), .ZN(n20310) );
  NAND3_X1 U23208 ( .A1(n24878), .A2(n24877), .A3(n24876), .ZN(n24880) );
  INV_X1 U23210 ( .I(n17525), .ZN(n15274) );
  AND3_X1 U23211 ( .A1(n24316), .A2(n16305), .A3(n26938), .Z(n16304) );
  NAND2_X1 U23214 ( .A1(n15413), .A2(n15412), .ZN(n21483) );
  XNOR2_X1 U23219 ( .A1(n31374), .A2(n25364), .ZN(n17106) );
  XOR2_X1 U23221 ( .A1(n15292), .A2(n25560), .Z(Ciphertext[125]) );
  INV_X2 U23222 ( .I(n15294), .ZN(n15295) );
  INV_X1 U23224 ( .I(n23282), .ZN(n15305) );
  NOR2_X1 U23228 ( .A1(n832), .A2(n27189), .ZN(n25733) );
  XOR2_X1 U23232 ( .A1(n24691), .A2(n12969), .Z(n15334) );
  INV_X1 U23236 ( .I(n20851), .ZN(n15337) );
  XOR2_X1 U23238 ( .A1(n29190), .A2(n25364), .Z(n23207) );
  XOR2_X1 U23240 ( .A1(n23168), .A2(n15370), .Z(n15346) );
  INV_X2 U23241 ( .I(n15347), .ZN(n18720) );
  OR2_X1 U23242 ( .A1(n18720), .A2(n16614), .Z(n15348) );
  XOR2_X1 U23244 ( .A1(n8491), .A2(n32813), .Z(n15744) );
  XOR2_X1 U23245 ( .A1(n11481), .A2(n30309), .Z(n18190) );
  XOR2_X1 U23246 ( .A1(n20183), .A2(n24991), .Z(n15352) );
  INV_X1 U23249 ( .I(n15364), .ZN(n22803) );
  XOR2_X1 U23251 ( .A1(n23297), .A2(n16581), .Z(n15370) );
  XOR2_X1 U23252 ( .A1(n23150), .A2(n25669), .Z(n15373) );
  XOR2_X1 U23254 ( .A1(n17407), .A2(n24855), .Z(n25201) );
  INV_X2 U23257 ( .I(n15384), .ZN(n21923) );
  XOR2_X1 U23259 ( .A1(n17918), .A2(n15386), .Z(n17917) );
  XOR2_X1 U23260 ( .A1(n22130), .A2(n25772), .Z(n15386) );
  XOR2_X1 U23266 ( .A1(n207), .A2(n15415), .Z(n18105) );
  INV_X2 U23268 ( .I(n25710), .ZN(n25760) );
  XOR2_X1 U23269 ( .A1(n14428), .A2(n25500), .Z(n21010) );
  XOR2_X1 U23270 ( .A1(n5149), .A2(n15420), .Z(n15419) );
  XOR2_X1 U23271 ( .A1(n702), .A2(n16597), .Z(n15420) );
  XOR2_X1 U23272 ( .A1(n5482), .A2(n24527), .Z(n21905) );
  INV_X1 U23273 ( .I(n15421), .ZN(n22754) );
  MUX2_X1 U23274 ( .I0(n23000), .I1(n13159), .S(n15421), .Z(n23006) );
  XOR2_X1 U23279 ( .A1(n15432), .A2(n15431), .Z(n15430) );
  XOR2_X1 U23280 ( .A1(n16076), .A2(n16584), .Z(n15431) );
  NAND2_X1 U23284 ( .A1(n15442), .A2(n21239), .ZN(n15441) );
  XOR2_X1 U23286 ( .A1(n27151), .A2(n24809), .Z(n15452) );
  XOR2_X1 U23287 ( .A1(n21945), .A2(n25880), .Z(n15460) );
  XOR2_X1 U23292 ( .A1(n15329), .A2(n22970), .Z(n23153) );
  XOR2_X1 U23293 ( .A1(n23152), .A2(n23154), .Z(n15470) );
  XOR2_X1 U23294 ( .A1(n460), .A2(n15471), .Z(n15472) );
  NAND2_X1 U23296 ( .A1(n23855), .A2(n4177), .ZN(n15475) );
  NAND2_X2 U23298 ( .A1(n25336), .A2(n15480), .ZN(n25368) );
  XOR2_X1 U23301 ( .A1(n23399), .A2(n23217), .Z(n15489) );
  INV_X2 U23303 ( .I(n15496), .ZN(n15528) );
  XOR2_X1 U23310 ( .A1(n23284), .A2(n23283), .Z(n15515) );
  XOR2_X1 U23311 ( .A1(n15517), .A2(n11370), .Z(n15987) );
  XOR2_X1 U23313 ( .A1(n15526), .A2(n15523), .Z(n21233) );
  XOR2_X1 U23314 ( .A1(n15525), .A2(n15524), .Z(n15523) );
  XOR2_X1 U23315 ( .A1(n20733), .A2(n25208), .Z(n15524) );
  XOR2_X1 U23318 ( .A1(n20975), .A2(n1070), .Z(n15538) );
  XOR2_X1 U23319 ( .A1(n15875), .A2(n15540), .Z(n15539) );
  XOR2_X1 U23320 ( .A1(n20821), .A2(n30303), .Z(n15540) );
  XOR2_X1 U23324 ( .A1(n24515), .A2(n24815), .Z(n15543) );
  INV_X2 U23328 ( .I(n23352), .ZN(n23764) );
  XOR2_X1 U23331 ( .A1(n22062), .A2(n22060), .Z(n15561) );
  XOR2_X1 U23332 ( .A1(n21048), .A2(n31584), .Z(n15562) );
  XOR2_X1 U23333 ( .A1(n19513), .A2(n15566), .Z(n15565) );
  NAND3_X2 U23338 ( .A1(n15579), .A2(n21983), .A3(n15578), .ZN(n23209) );
  XOR2_X1 U23339 ( .A1(Plaintext[165]), .A2(Key[165]), .Z(n17167) );
  NOR2_X1 U23340 ( .A1(n31533), .A2(n2928), .ZN(n15590) );
  NAND2_X2 U23341 ( .A1(n15594), .A2(n15592), .ZN(n20395) );
  NOR2_X1 U23342 ( .A1(n6842), .A2(n5480), .ZN(n21244) );
  NAND2_X1 U23343 ( .A1(n13506), .A2(n6842), .ZN(n21633) );
  NAND2_X1 U23348 ( .A1(n10183), .A2(n9234), .ZN(n15644) );
  XOR2_X1 U23351 ( .A1(n15668), .A2(n15667), .Z(n15666) );
  XOR2_X1 U23352 ( .A1(n20869), .A2(n21018), .Z(n15667) );
  XOR2_X1 U23354 ( .A1(n24816), .A2(n15671), .Z(n24452) );
  INV_X2 U23356 ( .I(n16939), .ZN(n16451) );
  INV_X2 U23360 ( .I(n18071), .ZN(n18743) );
  XOR2_X1 U23361 ( .A1(n15788), .A2(n19447), .Z(n19449) );
  XOR2_X1 U23363 ( .A1(n23210), .A2(n23212), .Z(n15691) );
  XOR2_X1 U23365 ( .A1(n15978), .A2(n25054), .Z(n15702) );
  XOR2_X1 U23367 ( .A1(n30183), .A2(n24839), .Z(n15707) );
  XOR2_X1 U23370 ( .A1(Plaintext[171]), .A2(Key[171]), .Z(n17029) );
  XOR2_X1 U23374 ( .A1(n21994), .A2(n1398), .Z(n15725) );
  INV_X2 U23382 ( .I(n15754), .ZN(n25238) );
  XOR2_X1 U23385 ( .A1(n32893), .A2(n1394), .Z(n15761) );
  INV_X1 U23386 ( .I(n24823), .ZN(n15765) );
  OAI21_X2 U23387 ( .A1(n15896), .A2(n15771), .B(n15769), .ZN(n25258) );
  XOR2_X1 U23392 ( .A1(n15792), .A2(n7511), .Z(n15791) );
  XOR2_X1 U23395 ( .A1(n10522), .A2(n15802), .Z(n15801) );
  XOR2_X1 U23398 ( .A1(n19703), .A2(n15816), .Z(n15815) );
  XOR2_X1 U23399 ( .A1(n15817), .A2(n20357), .Z(n21225) );
  XOR2_X1 U23402 ( .A1(n19483), .A2(n25879), .Z(n15819) );
  XOR2_X1 U23405 ( .A1(n22164), .A2(n15822), .Z(n15821) );
  OR2_X1 U23407 ( .A1(n21603), .A2(n31960), .Z(n15828) );
  NOR2_X1 U23408 ( .A1(n21629), .A2(n21630), .ZN(n15840) );
  XOR2_X1 U23409 ( .A1(n15861), .A2(n24644), .Z(n15860) );
  XOR2_X1 U23410 ( .A1(n25182), .A2(n12969), .Z(n15861) );
  MUX2_X1 U23419 ( .I0(n24256), .I1(n24255), .S(n15876), .Z(n24259) );
  XOR2_X1 U23424 ( .A1(n15183), .A2(n16636), .Z(n15886) );
  XNOR2_X1 U23425 ( .A1(n5932), .A2(n6547), .ZN(n15887) );
  XOR2_X1 U23426 ( .A1(n21027), .A2(n15890), .Z(n15889) );
  XOR2_X1 U23427 ( .A1(n20641), .A2(n20921), .Z(n15890) );
  XOR2_X1 U23428 ( .A1(n20919), .A2(n20922), .Z(n15891) );
  XOR2_X1 U23429 ( .A1(n646), .A2(n23430), .Z(n15897) );
  NAND3_X1 U23431 ( .A1(n22754), .A2(n806), .A3(n13159), .ZN(n22755) );
  XOR2_X1 U23433 ( .A1(n19378), .A2(n27672), .Z(n15904) );
  INV_X1 U23434 ( .I(n15909), .ZN(n18762) );
  AOI21_X1 U23435 ( .A1(n15909), .A2(n18499), .B(n33472), .ZN(n18503) );
  XOR2_X1 U23436 ( .A1(Plaintext[69]), .A2(Key[69]), .Z(n18498) );
  XOR2_X1 U23437 ( .A1(n15913), .A2(n19602), .Z(n19613) );
  INV_X1 U23440 ( .I(n15929), .ZN(n17318) );
  XOR2_X1 U23443 ( .A1(n24546), .A2(n545), .Z(n15934) );
  NOR2_X1 U23445 ( .A1(n19124), .A2(n8233), .ZN(n19125) );
  NAND3_X1 U23450 ( .A1(n25845), .A2(n25844), .A3(n25846), .ZN(n15947) );
  XOR2_X1 U23451 ( .A1(n24777), .A2(n15949), .Z(n15948) );
  XOR2_X1 U23452 ( .A1(n12969), .A2(n7511), .Z(n15949) );
  XOR2_X1 U23454 ( .A1(n15959), .A2(n16657), .Z(Ciphertext[168]) );
  XOR2_X1 U23455 ( .A1(n400), .A2(n25716), .Z(n19376) );
  XOR2_X1 U23456 ( .A1(n11891), .A2(n25208), .Z(n15963) );
  XOR2_X1 U23457 ( .A1(Plaintext[125]), .A2(Key[125]), .Z(n17143) );
  NOR2_X1 U23458 ( .A1(n17184), .A2(n18845), .ZN(n15967) );
  INV_X2 U23459 ( .I(n17029), .ZN(n17184) );
  XOR2_X1 U23461 ( .A1(n9327), .A2(n19507), .Z(n19415) );
  XOR2_X1 U23462 ( .A1(n22072), .A2(n34150), .Z(n15969) );
  NAND2_X1 U23463 ( .A1(n15976), .A2(n3183), .ZN(n22051) );
  XOR2_X1 U23466 ( .A1(n19408), .A2(n17551), .Z(n15983) );
  XOR2_X1 U23468 ( .A1(n15992), .A2(n15994), .Z(n16129) );
  XOR2_X1 U23469 ( .A1(n15993), .A2(n20902), .Z(n15992) );
  XOR2_X1 U23470 ( .A1(n21997), .A2(n15998), .Z(n16000) );
  XOR2_X1 U23471 ( .A1(n22030), .A2(n22305), .Z(n15998) );
  XOR2_X1 U23472 ( .A1(n21998), .A2(n21999), .Z(n15999) );
  XOR2_X1 U23473 ( .A1(n19378), .A2(n30411), .Z(n16005) );
  XOR2_X1 U23474 ( .A1(n23367), .A2(n23368), .Z(n16010) );
  AOI22_X1 U23477 ( .A1(n24615), .A2(n33434), .B1(n16383), .B2(n1208), .ZN(
        n16021) );
  XOR2_X1 U23478 ( .A1(n16302), .A2(n16997), .Z(n16996) );
  XOR2_X1 U23481 ( .A1(n16036), .A2(n17529), .Z(n16035) );
  OAI21_X1 U23482 ( .A1(n20608), .A2(n20606), .B(n16481), .ZN(n20368) );
  NAND2_X1 U23487 ( .A1(n24912), .A2(n24911), .ZN(n17883) );
  INV_X1 U23489 ( .I(n24144), .ZN(n16039) );
  NAND2_X1 U23491 ( .A1(n23815), .A2(n354), .ZN(n23818) );
  XOR2_X1 U23494 ( .A1(n322), .A2(n25669), .Z(n17991) );
  AND2_X1 U23497 ( .A1(n19614), .A2(n4587), .Z(n19622) );
  INV_X2 U23498 ( .I(n16062), .ZN(n25701) );
  XOR2_X1 U23501 ( .A1(n19533), .A2(n19532), .Z(n19833) );
  XOR2_X1 U23512 ( .A1(n16104), .A2(n16697), .Z(Ciphertext[46]) );
  AOI21_X2 U23518 ( .A1(n21156), .A2(n27543), .B(n21155), .ZN(n22072) );
  XNOR2_X1 U23519 ( .A1(n19708), .A2(n24514), .ZN(n18082) );
  NAND2_X1 U23523 ( .A1(n11892), .A2(n11804), .ZN(n17076) );
  XOR2_X1 U23524 ( .A1(n28813), .A2(n25161), .Z(n16773) );
  XOR2_X1 U23526 ( .A1(n24695), .A2(n24357), .Z(n16416) );
  OR2_X1 U23530 ( .A1(n25912), .A2(n25922), .Z(n25920) );
  OAI22_X1 U23535 ( .A1(n18624), .A2(n16522), .B1(n828), .B2(n18623), .ZN(
        n16156) );
  XOR2_X1 U23539 ( .A1(n23363), .A2(n23535), .Z(n16162) );
  AOI21_X1 U23541 ( .A1(n25281), .A2(n733), .B(n17876), .ZN(n17875) );
  XOR2_X1 U23544 ( .A1(n20907), .A2(n21036), .Z(n16191) );
  INV_X1 U23545 ( .I(n15116), .ZN(n23595) );
  XOR2_X1 U23546 ( .A1(n21900), .A2(n21899), .Z(n21901) );
  NAND2_X1 U23553 ( .A1(n18785), .A2(n32108), .ZN(n18367) );
  XOR2_X1 U23555 ( .A1(n21923), .A2(n22012), .Z(n21281) );
  INV_X2 U23556 ( .I(n16220), .ZN(n16766) );
  XOR2_X1 U23557 ( .A1(Plaintext[56]), .A2(Key[56]), .Z(n16220) );
  XOR2_X1 U23559 ( .A1(Plaintext[143]), .A2(Key[143]), .Z(n18071) );
  NAND2_X2 U23561 ( .A1(n24709), .A2(n24708), .ZN(n25820) );
  XOR2_X1 U23563 ( .A1(n20930), .A2(n17106), .Z(n17957) );
  XOR2_X1 U23564 ( .A1(n16237), .A2(n30275), .Z(n18149) );
  NAND2_X1 U23565 ( .A1(n19089), .A2(n5760), .ZN(n19090) );
  INV_X1 U23572 ( .I(n1053), .ZN(n19361) );
  XOR2_X1 U23574 ( .A1(n19689), .A2(n19690), .Z(n19695) );
  INV_X2 U23578 ( .I(n16277), .ZN(n22433) );
  XOR2_X1 U23581 ( .A1(n16284), .A2(n16581), .Z(Ciphertext[92]) );
  INV_X1 U23586 ( .I(n22873), .ZN(n22916) );
  XOR2_X1 U23590 ( .A1(Plaintext[89]), .A2(Key[89]), .Z(n16310) );
  OAI21_X1 U23591 ( .A1(n25745), .A2(n25746), .B(n25744), .ZN(n25747) );
  XOR2_X1 U23597 ( .A1(Key[81]), .A2(Plaintext[81]), .Z(n18613) );
  NAND2_X1 U23603 ( .A1(n21760), .A2(n21759), .ZN(n21765) );
  INV_X1 U23604 ( .I(n19108), .ZN(n18930) );
  INV_X1 U23613 ( .I(n29269), .ZN(n23932) );
  XOR2_X1 U23615 ( .A1(n16378), .A2(n18382), .Z(n18818) );
  INV_X1 U23616 ( .I(n32874), .ZN(n25773) );
  XOR2_X1 U23617 ( .A1(n4400), .A2(n16081), .Z(n19787) );
  XOR2_X1 U23618 ( .A1(n17042), .A2(n17041), .Z(n17119) );
  NAND2_X1 U23625 ( .A1(n16412), .A2(n16411), .ZN(n18169) );
  XOR2_X1 U23630 ( .A1(n19628), .A2(n16437), .Z(n19631) );
  XOR2_X1 U23631 ( .A1(n29030), .A2(n16438), .Z(n16437) );
  XOR2_X1 U23632 ( .A1(n22154), .A2(n21884), .Z(n16439) );
  XOR2_X1 U23633 ( .A1(n7879), .A2(n25282), .Z(n24769) );
  XOR2_X1 U23634 ( .A1(n20984), .A2(n20593), .Z(n20600) );
  XOR2_X1 U23638 ( .A1(n16242), .A2(n21889), .Z(n16457) );
  XOR2_X1 U23642 ( .A1(n17434), .A2(n17435), .Z(n20064) );
  OR2_X1 U23644 ( .A1(n23753), .A2(n11922), .Z(n23727) );
  BUF_X2 U23650 ( .I(n20015), .Z(n16491) );
  NOR2_X1 U23655 ( .A1(n18196), .A2(n18195), .ZN(n18194) );
  XOR2_X1 U23657 ( .A1(n26794), .A2(n16672), .Z(n16513) );
  OR3_X1 U23661 ( .A1(n1141), .A2(n29497), .A3(n929), .Z(n17171) );
  XOR2_X1 U23665 ( .A1(n16541), .A2(n30993), .Z(Ciphertext[147]) );
  AOI22_X1 U23669 ( .A1(n21065), .A2(n29460), .B1(n21064), .B2(n28642), .ZN(
        n16553) );
  XOR2_X1 U23671 ( .A1(Plaintext[17]), .A2(Key[17]), .Z(n18198) );
  NAND3_X1 U23681 ( .A1(n25365), .A2(n750), .A3(n25366), .ZN(n25372) );
  NAND2_X1 U23692 ( .A1(n16937), .A2(n25322), .ZN(n16660) );
  XOR2_X1 U23699 ( .A1(n21997), .A2(n21920), .Z(n17452) );
  XOR2_X1 U23701 ( .A1(n16689), .A2(n22179), .Z(n22589) );
  XOR2_X1 U23703 ( .A1(n21951), .A2(n21949), .Z(n16692) );
  INV_X2 U23704 ( .I(n16695), .ZN(n18064) );
  XOR2_X1 U23707 ( .A1(Plaintext[55]), .A2(Key[55]), .Z(n16819) );
  BUF_X2 U23708 ( .I(Key[191]), .Z(n16703) );
  XOR2_X1 U23709 ( .A1(n24768), .A2(n29274), .Z(n16730) );
  INV_X2 U23710 ( .I(n16711), .ZN(n25145) );
  XOR2_X1 U23713 ( .A1(n12), .A2(n30301), .Z(n16718) );
  NOR2_X1 U23714 ( .A1(n11930), .A2(n16432), .ZN(n16724) );
  XOR2_X1 U23715 ( .A1(n19502), .A2(n19501), .Z(n16734) );
  XOR2_X1 U23717 ( .A1(n8109), .A2(n16738), .Z(n16737) );
  XOR2_X1 U23718 ( .A1(n18216), .A2(n24671), .Z(n16739) );
  XOR2_X1 U23724 ( .A1(n16754), .A2(n17576), .Z(n16753) );
  INV_X2 U23725 ( .I(n16756), .ZN(n21203) );
  XOR2_X1 U23727 ( .A1(n17555), .A2(n16604), .Z(n16767) );
  INV_X2 U23733 ( .I(n16776), .ZN(n23575) );
  NAND2_X1 U23734 ( .A1(n17079), .A2(n16780), .ZN(n17982) );
  NAND2_X1 U23735 ( .A1(n17079), .A2(n13401), .ZN(n17983) );
  OAI21_X1 U23739 ( .A1(n21259), .A2(n16652), .B(n21257), .ZN(n21260) );
  AND2_X1 U23741 ( .A1(n16819), .A2(n16766), .Z(n18486) );
  XOR2_X1 U23742 ( .A1(n13602), .A2(n10766), .Z(n16823) );
  XOR2_X1 U23744 ( .A1(n28163), .A2(n16649), .Z(n20827) );
  NAND2_X1 U23745 ( .A1(n20325), .A2(n28011), .ZN(n17514) );
  XOR2_X1 U23748 ( .A1(n19550), .A2(n27137), .Z(n16841) );
  XOR2_X1 U23750 ( .A1(n19474), .A2(n16690), .Z(n19475) );
  INV_X1 U23751 ( .I(n16448), .ZN(n20821) );
  MUX2_X1 U23753 ( .I0(n18943), .I1(n18944), .S(n18995), .Z(n18947) );
  XOR2_X1 U23756 ( .A1(n11166), .A2(n22198), .Z(n17258) );
  XOR2_X1 U23757 ( .A1(n16869), .A2(n25545), .Z(Ciphertext[121]) );
  NAND3_X1 U23758 ( .A1(n1049), .A2(n29815), .A3(n19326), .ZN(n16871) );
  AOI21_X1 U23759 ( .A1(n20627), .A2(n7280), .B(n14005), .ZN(n16883) );
  INV_X2 U23760 ( .I(n16885), .ZN(n22435) );
  XOR2_X1 U23762 ( .A1(n17913), .A2(n17915), .Z(n16887) );
  XOR2_X1 U23765 ( .A1(Plaintext[75]), .A2(Key[75]), .Z(n16899) );
  INV_X2 U23766 ( .I(n16899), .ZN(n18774) );
  XOR2_X1 U23768 ( .A1(n22015), .A2(n16911), .Z(n16910) );
  INV_X2 U23769 ( .I(n16913), .ZN(n18151) );
  NAND2_X2 U23770 ( .A1(n16926), .A2(n16928), .ZN(n23453) );
  XOR2_X1 U23773 ( .A1(n26701), .A2(n24748), .Z(n23279) );
  XOR2_X1 U23776 ( .A1(n22013), .A2(n26000), .Z(n16945) );
  XOR2_X1 U23777 ( .A1(n22303), .A2(n21994), .Z(n16946) );
  XOR2_X1 U23783 ( .A1(n22141), .A2(n24231), .Z(n16974) );
  INV_X2 U23784 ( .I(n16996), .ZN(n20103) );
  XOR2_X1 U23785 ( .A1(n19567), .A2(n12137), .Z(n16997) );
  XOR2_X1 U23787 ( .A1(n23440), .A2(n17013), .Z(n17012) );
  XOR2_X1 U23788 ( .A1(n10773), .A2(n16613), .Z(n17013) );
  XOR2_X1 U23791 ( .A1(n20722), .A2(n20724), .Z(n17026) );
  XOR2_X1 U23796 ( .A1(n24666), .A2(n17049), .Z(n17048) );
  XOR2_X1 U23797 ( .A1(n16128), .A2(n705), .Z(n17049) );
  INV_X2 U23798 ( .I(n17050), .ZN(n23735) );
  MUX2_X1 U23802 ( .I0(n27143), .I1(n13896), .S(n16072), .Z(n21199) );
  XOR2_X1 U23803 ( .A1(n29312), .A2(n16636), .Z(n17072) );
  XOR2_X1 U23804 ( .A1(Plaintext[88]), .A2(Key[88]), .Z(n18569) );
  AOI21_X1 U23806 ( .A1(n16337), .A2(n23763), .B(n17087), .ZN(n17086) );
  XOR2_X1 U23807 ( .A1(n19698), .A2(n17091), .Z(n17090) );
  OR2_X1 U23812 ( .A1(n751), .A2(n25627), .Z(n17108) );
  XOR2_X1 U23814 ( .A1(n17115), .A2(n8139), .Z(Ciphertext[16]) );
  XOR2_X1 U23818 ( .A1(n19766), .A2(n12103), .Z(n17125) );
  INV_X2 U23819 ( .I(n17127), .ZN(n19867) );
  XOR2_X1 U23821 ( .A1(n5380), .A2(n1433), .Z(n23340) );
  NAND2_X1 U23822 ( .A1(n17134), .A2(n31959), .ZN(n23542) );
  INV_X2 U23823 ( .I(n24726), .ZN(n25885) );
  XOR2_X1 U23828 ( .A1(n22067), .A2(n22198), .Z(n17145) );
  NOR2_X1 U23830 ( .A1(n27597), .A2(n10831), .ZN(n17363) );
  MUX2_X1 U23831 ( .I0(n19856), .I1(n17365), .S(n10831), .Z(n17364) );
  NAND2_X2 U23832 ( .A1(n20189), .A2(n20191), .ZN(n20531) );
  XOR2_X1 U23833 ( .A1(n24518), .A2(n24444), .Z(n17159) );
  NAND2_X1 U23835 ( .A1(n6638), .A2(n12548), .ZN(n17162) );
  OR2_X1 U23836 ( .A1(n22636), .A2(n22637), .Z(n17163) );
  XNOR2_X1 U23838 ( .A1(Plaintext[90]), .A2(Key[90]), .ZN(n17168) );
  NAND3_X1 U23839 ( .A1(n33972), .A2(n29497), .A3(n21414), .ZN(n17172) );
  XOR2_X1 U23841 ( .A1(n33572), .A2(n29951), .Z(n17174) );
  XOR2_X1 U23843 ( .A1(n22108), .A2(n22055), .Z(n22152) );
  XOR2_X1 U23844 ( .A1(n17188), .A2(n23413), .Z(n23415) );
  XOR2_X1 U23845 ( .A1(n17193), .A2(n17192), .Z(n20133) );
  XOR2_X1 U23847 ( .A1(n30305), .A2(n28806), .Z(n19729) );
  NAND2_X1 U23848 ( .A1(n25899), .A2(n18219), .ZN(n17196) );
  XOR2_X1 U23851 ( .A1(n30284), .A2(n17206), .Z(n17205) );
  INV_X1 U23852 ( .I(n22029), .ZN(n17206) );
  XOR2_X1 U23853 ( .A1(n17207), .A2(n17258), .Z(n22090) );
  OAI21_X2 U23857 ( .A1(n21390), .A2(n17217), .B(n17215), .ZN(n21849) );
  XOR2_X1 U23859 ( .A1(n4554), .A2(n23478), .Z(n17235) );
  NAND2_X1 U23860 ( .A1(n17237), .A2(n20401), .ZN(n20574) );
  XOR2_X1 U23861 ( .A1(n1004), .A2(n1306), .Z(n17244) );
  INV_X2 U23865 ( .I(n17255), .ZN(n17582) );
  XOR2_X1 U23866 ( .A1(n21961), .A2(n21962), .Z(n17259) );
  XOR2_X1 U23872 ( .A1(n20668), .A2(n17282), .Z(n17281) );
  XOR2_X1 U23873 ( .A1(n21044), .A2(n20586), .Z(n17282) );
  INV_X1 U23875 ( .I(n17289), .ZN(n17290) );
  NAND2_X1 U23876 ( .A1(n32063), .A2(n24955), .ZN(n24957) );
  XOR2_X1 U23881 ( .A1(n24674), .A2(n24429), .Z(n17307) );
  NAND2_X1 U23882 ( .A1(n24103), .A2(n17310), .ZN(n23664) );
  XOR2_X1 U23885 ( .A1(n24526), .A2(n16038), .Z(n24542) );
  XOR2_X1 U23886 ( .A1(n24526), .A2(n14648), .Z(n24752) );
  AND2_X1 U23887 ( .A1(n18965), .A2(n18955), .Z(n17320) );
  NOR2_X2 U23888 ( .A1(n19273), .A2(n19272), .ZN(n19772) );
  XOR2_X1 U23890 ( .A1(n30443), .A2(n17324), .Z(n17323) );
  INV_X1 U23891 ( .I(n25827), .ZN(n17324) );
  NOR2_X1 U23894 ( .A1(n14312), .A2(n947), .ZN(n18982) );
  XOR2_X1 U23895 ( .A1(n29312), .A2(n16402), .Z(n19750) );
  XNOR2_X1 U23896 ( .A1(n23336), .A2(n23335), .ZN(n23446) );
  XOR2_X1 U23897 ( .A1(n17353), .A2(n23445), .Z(n17351) );
  XOR2_X1 U23899 ( .A1(n31908), .A2(n19342), .Z(n17355) );
  XOR2_X1 U23900 ( .A1(n19588), .A2(n19340), .Z(n17356) );
  NOR2_X1 U23902 ( .A1(n25590), .A2(n26912), .ZN(n17367) );
  XOR2_X1 U23904 ( .A1(n17380), .A2(n17381), .Z(n20117) );
  XOR2_X1 U23905 ( .A1(n19739), .A2(n12136), .Z(n17381) );
  OR2_X1 U23906 ( .A1(n25316), .A2(n1074), .Z(n17383) );
  XOR2_X1 U23907 ( .A1(n26582), .A2(n16642), .Z(n18015) );
  NAND2_X1 U23909 ( .A1(n25546), .A2(n25542), .ZN(n17402) );
  AND2_X1 U23915 ( .A1(n21349), .A2(n21348), .Z(n17418) );
  NOR2_X1 U23916 ( .A1(n17419), .A2(n18722), .ZN(n18301) );
  XOR2_X1 U23920 ( .A1(n17436), .A2(n19706), .Z(n17435) );
  XOR2_X1 U23921 ( .A1(n31450), .A2(n1191), .Z(n17436) );
  INV_X4 U23923 ( .I(n18923), .ZN(n17445) );
  MUX2_X1 U23924 ( .I0(n18719), .I1(n18718), .S(n18855), .Z(n17446) );
  NAND2_X2 U23925 ( .A1(n18734), .A2(n18735), .ZN(n18980) );
  INV_X2 U23926 ( .I(n17450), .ZN(n22332) );
  XOR2_X1 U23928 ( .A1(n23168), .A2(n23167), .Z(n17457) );
  XOR2_X1 U23933 ( .A1(Key[0]), .A2(Plaintext[0]), .Z(n18882) );
  XOR2_X1 U23938 ( .A1(n6547), .A2(n16697), .Z(n24375) );
  XOR2_X1 U23939 ( .A1(n6547), .A2(n24839), .Z(n24840) );
  XOR2_X1 U23944 ( .A1(n22033), .A2(n22205), .Z(n17529) );
  NAND2_X1 U23953 ( .A1(n17630), .A2(n22472), .ZN(n17567) );
  NAND3_X1 U23954 ( .A1(n13746), .A2(n17569), .A3(n22472), .ZN(n17568) );
  XOR2_X1 U23955 ( .A1(n24597), .A2(n17571), .Z(n17570) );
  XOR2_X1 U23956 ( .A1(n24596), .A2(n24595), .Z(n17572) );
  XOR2_X1 U23960 ( .A1(Plaintext[44]), .A2(Key[44]), .Z(n18076) );
  INV_X1 U23961 ( .I(n25911), .ZN(n17600) );
  XOR2_X1 U23962 ( .A1(n16319), .A2(n25519), .Z(n18144) );
  XOR2_X1 U23963 ( .A1(n16319), .A2(n30954), .Z(n24451) );
  XOR2_X1 U23964 ( .A1(n16319), .A2(n25324), .Z(n24671) );
  XOR2_X1 U23966 ( .A1(n12), .A2(n16423), .Z(n24481) );
  XOR2_X1 U23968 ( .A1(n19463), .A2(n19412), .Z(n17613) );
  NOR2_X2 U23972 ( .A1(n18741), .A2(n18740), .ZN(n19262) );
  XOR2_X1 U23976 ( .A1(n34120), .A2(n16671), .Z(n17628) );
  NOR2_X1 U23978 ( .A1(n25495), .A2(n30935), .ZN(n25498) );
  OAI21_X1 U23979 ( .A1(n25496), .A2(n30935), .B(n17636), .ZN(n25497) );
  XOR2_X1 U23982 ( .A1(n20868), .A2(n20867), .Z(n17643) );
  XNOR2_X1 U23984 ( .A1(Plaintext[100]), .A2(Key[100]), .ZN(n17649) );
  XOR2_X1 U23985 ( .A1(n19730), .A2(n17651), .Z(n17650) );
  XOR2_X1 U23986 ( .A1(n19779), .A2(n25832), .Z(n17651) );
  OR2_X1 U23988 ( .A1(n20651), .A2(n23191), .Z(n17658) );
  NOR2_X1 U23989 ( .A1(n25057), .A2(n25058), .ZN(n17744) );
  NOR2_X1 U23992 ( .A1(n17675), .A2(n19794), .ZN(n20209) );
  XOR2_X1 U23993 ( .A1(n25249), .A2(n16548), .Z(Ciphertext[78]) );
  XOR2_X1 U23994 ( .A1(n17679), .A2(n22032), .Z(n22035) );
  INV_X2 U23996 ( .I(n17683), .ZN(n25012) );
  XOR2_X1 U23999 ( .A1(n27148), .A2(n27995), .Z(n17704) );
  XOR2_X1 U24001 ( .A1(n24646), .A2(n25457), .Z(n17705) );
  NAND3_X1 U24004 ( .A1(n6072), .A2(n32483), .A3(n22584), .ZN(n17718) );
  XNOR2_X1 U24007 ( .A1(n33373), .A2(n20699), .ZN(n20868) );
  XOR2_X1 U24009 ( .A1(n17738), .A2(n20675), .Z(n21136) );
  OR2_X1 U24012 ( .A1(n25059), .A2(n28070), .Z(n17742) );
  XOR2_X1 U24013 ( .A1(n17752), .A2(n17754), .Z(n24368) );
  XOR2_X1 U24014 ( .A1(n24673), .A2(n17755), .Z(n17754) );
  XOR2_X1 U24015 ( .A1(n24531), .A2(n24801), .Z(n17755) );
  XOR2_X1 U24016 ( .A1(n22165), .A2(n22163), .Z(n17765) );
  INV_X2 U24017 ( .I(n17768), .ZN(n23942) );
  NAND2_X1 U24018 ( .A1(n17781), .A2(n15046), .ZN(n17778) );
  NAND2_X1 U24020 ( .A1(n17810), .A2(n945), .ZN(n18897) );
  NAND2_X1 U24026 ( .A1(n31533), .A2(n2928), .ZN(n17809) );
  XOR2_X1 U24027 ( .A1(n19637), .A2(n1366), .Z(n19639) );
  NAND2_X1 U24029 ( .A1(n28528), .A2(n17817), .ZN(n18359) );
  XOR2_X1 U24032 ( .A1(n15844), .A2(n29728), .Z(n17834) );
  XOR2_X1 U24033 ( .A1(n17837), .A2(n21035), .Z(n20660) );
  XOR2_X1 U24035 ( .A1(n17844), .A2(n25619), .Z(Ciphertext[137]) );
  OR2_X1 U24037 ( .A1(n25488), .A2(n25478), .Z(n17850) );
  XOR2_X1 U24043 ( .A1(n24687), .A2(n24688), .Z(n17869) );
  XOR2_X1 U24044 ( .A1(n17875), .A2(n27672), .Z(Ciphertext[87]) );
  NAND2_X1 U24045 ( .A1(n23899), .A2(n4069), .ZN(n17881) );
  OR2_X1 U24046 ( .A1(n24908), .A2(n6154), .Z(n17884) );
  INV_X2 U24047 ( .I(n17886), .ZN(n24610) );
  INV_X2 U24049 ( .I(n17903), .ZN(n25755) );
  XOR2_X1 U24050 ( .A1(n24825), .A2(n24401), .Z(n17904) );
  XNOR2_X1 U24052 ( .A1(n17919), .A2(n17917), .ZN(n17916) );
  XOR2_X1 U24054 ( .A1(n17933), .A2(n293), .Z(Ciphertext[74]) );
  XOR2_X1 U24055 ( .A1(n23259), .A2(n25856), .Z(n17934) );
  XOR2_X1 U24057 ( .A1(n24491), .A2(n18138), .Z(n17938) );
  NOR2_X1 U24061 ( .A1(n17948), .A2(n25446), .ZN(n25424) );
  NAND2_X1 U24065 ( .A1(n739), .A2(n23889), .ZN(n17949) );
  XOR2_X1 U24069 ( .A1(n14337), .A2(n26751), .Z(n17958) );
  XOR2_X1 U24072 ( .A1(Plaintext[134]), .A2(Key[134]), .Z(n17970) );
  AOI21_X1 U24074 ( .A1(n31435), .A2(n3241), .B(n28365), .ZN(n17977) );
  NAND2_X1 U24075 ( .A1(n23807), .A2(n23848), .ZN(n17978) );
  XOR2_X1 U24076 ( .A1(n25181), .A2(n25182), .Z(Ciphertext[65]) );
  XOR2_X1 U24082 ( .A1(n20970), .A2(n32052), .Z(n17998) );
  XOR2_X1 U24083 ( .A1(n21040), .A2(n25009), .Z(n18010) );
  XOR2_X1 U24084 ( .A1(n28806), .A2(n24966), .Z(n18011) );
  AND2_X1 U24086 ( .A1(n22610), .A2(n22634), .Z(n18013) );
  XOR2_X1 U24089 ( .A1(n20957), .A2(n20682), .Z(n18024) );
  XOR2_X1 U24092 ( .A1(n19445), .A2(n24917), .Z(n18031) );
  NAND2_X1 U24093 ( .A1(n16345), .A2(n21463), .ZN(n18034) );
  NOR2_X1 U24095 ( .A1(n21812), .A2(n21811), .ZN(n18043) );
  INV_X2 U24103 ( .I(n18075), .ZN(n25198) );
  XNOR2_X1 U24105 ( .A1(Plaintext[46]), .A2(Key[46]), .ZN(n18085) );
  XOR2_X1 U24111 ( .A1(n18096), .A2(n20959), .Z(n18095) );
  XOR2_X1 U24112 ( .A1(n30163), .A2(n31233), .Z(n18096) );
  XOR2_X1 U24113 ( .A1(n23166), .A2(n18108), .Z(n18107) );
  NAND2_X1 U24115 ( .A1(n842), .A2(n667), .ZN(n23629) );
  INV_X1 U24117 ( .I(n23079), .ZN(n18129) );
  NAND2_X1 U24118 ( .A1(n18827), .A2(n18489), .ZN(n18130) );
  NOR2_X1 U24119 ( .A1(n18146), .A2(n24197), .ZN(n18145) );
  XOR2_X1 U24120 ( .A1(n18149), .A2(n18148), .Z(n21815) );
  XOR2_X1 U24121 ( .A1(n22240), .A2(n16602), .Z(n18148) );
  INV_X2 U24122 ( .I(n18155), .ZN(n25119) );
  XOR2_X1 U24124 ( .A1(n19619), .A2(n112), .Z(n18165) );
  XOR2_X1 U24125 ( .A1(n24513), .A2(n15742), .Z(n18173) );
  OAI21_X1 U24128 ( .A1(n4146), .A2(n25697), .B(n25699), .ZN(n18195) );
  XOR2_X1 U24132 ( .A1(n322), .A2(n18217), .Z(n18216) );
  INV_X2 U24133 ( .I(n18220), .ZN(n24436) );
  XOR2_X1 U24135 ( .A1(n29890), .A2(n19769), .Z(n19770) );
  XOR2_X1 U24137 ( .A1(n19741), .A2(n25161), .Z(n18231) );
  NAND2_X1 U24140 ( .A1(n19971), .A2(n18237), .ZN(n18236) );
  NAND2_X1 U24141 ( .A1(n19900), .A2(n19899), .ZN(n18237) );
  XOR2_X1 U24142 ( .A1(n18238), .A2(n19685), .Z(n20108) );
  XOR2_X1 U24143 ( .A1(n19681), .A2(n19680), .Z(n18238) );
  XOR2_X1 U24149 ( .A1(Plaintext[141]), .A2(Key[141]), .Z(n18314) );
  OAI22_X1 U24152 ( .A1(n25248), .A2(n27429), .B1(n25247), .B2(n25246), .ZN(
        n25249) );
  BUF_X2 U24156 ( .I(n18569), .Z(n18493) );
  INV_X1 U24158 ( .I(n20616), .ZN(n20363) );
  BUF_X2 U24161 ( .I(n21100), .Z(n21307) );
  NAND4_X1 U24163 ( .A1(n23998), .A2(n23997), .A3(n23922), .A4(n23921), .ZN(
        n23934) );
  XOR2_X1 U24166 ( .A1(Key[72]), .A2(Plaintext[72]), .Z(n18773) );
  INV_X1 U24167 ( .I(n18773), .ZN(n18770) );
  INV_X1 U24168 ( .I(Plaintext[59]), .ZN(n18275) );
  XOR2_X1 U24169 ( .A1(n18275), .A2(Key[59]), .Z(n18763) );
  INV_X1 U24171 ( .I(Plaintext[64]), .ZN(n18280) );
  INV_X1 U24172 ( .I(Plaintext[62]), .ZN(n18281) );
  XOR2_X1 U24173 ( .A1(n18281), .A2(Key[62]), .Z(n18780) );
  INV_X1 U24174 ( .I(Plaintext[80]), .ZN(n18282) );
  XOR2_X1 U24175 ( .A1(n18282), .A2(Key[80]), .Z(n18283) );
  INV_X1 U24176 ( .I(Plaintext[66]), .ZN(n18286) );
  XOR2_X1 U24177 ( .A1(n18286), .A2(Key[66]), .Z(n18756) );
  XOR2_X1 U24178 ( .A1(Key[67]), .A2(Plaintext[67]), .Z(n18335) );
  INV_X1 U24180 ( .I(Plaintext[68]), .ZN(n18287) );
  XOR2_X1 U24181 ( .A1(n18287), .A2(Key[68]), .Z(n18293) );
  NAND2_X1 U24182 ( .A1(n18338), .A2(n18605), .ZN(n18294) );
  NAND2_X1 U24183 ( .A1(n32437), .A2(n19108), .ZN(n18297) );
  XOR2_X1 U24186 ( .A1(Key[85]), .A2(Plaintext[85]), .Z(n18323) );
  XOR2_X1 U24189 ( .A1(Key[150]), .A2(Plaintext[150]), .Z(n18540) );
  XOR2_X1 U24190 ( .A1(Key[155]), .A2(Plaintext[155]), .Z(n18300) );
  XOR2_X1 U24191 ( .A1(Key[154]), .A2(Plaintext[154]), .Z(n18580) );
  XOR2_X1 U24192 ( .A1(Key[152]), .A2(Plaintext[152]), .Z(n18541) );
  INV_X1 U24193 ( .I(n18302), .ZN(n18304) );
  XOR2_X1 U24195 ( .A1(Key[137]), .A2(Plaintext[137]), .Z(n18310) );
  INV_X1 U24196 ( .I(n18314), .ZN(n18747) );
  INV_X1 U24197 ( .I(Plaintext[142]), .ZN(n18313) );
  XOR2_X1 U24198 ( .A1(n18313), .A2(Key[142]), .Z(n18434) );
  XOR2_X1 U24199 ( .A1(Key[139]), .A2(Plaintext[139]), .Z(n18707) );
  INV_X1 U24200 ( .I(Plaintext[130]), .ZN(n18315) );
  OAI21_X1 U24201 ( .A1(n1439), .A2(n18317), .B(n18316), .ZN(n18320) );
  XOR2_X1 U24202 ( .A1(Key[131]), .A2(Plaintext[131]), .Z(n18392) );
  MUX2_X1 U24203 ( .I0(n18492), .I1(n18566), .S(n18324), .Z(n18327) );
  NOR2_X1 U24205 ( .A1(n18328), .A2(n16564), .ZN(n18331) );
  AOI21_X1 U24208 ( .A1(n18840), .A2(n1181), .B(n30937), .ZN(n18347) );
  NAND2_X1 U24209 ( .A1(n26181), .A2(n19052), .ZN(n18346) );
  NAND3_X1 U24211 ( .A1(n18339), .A2(n18779), .A3(n10080), .ZN(n18341) );
  XOR2_X1 U24214 ( .A1(Key[39]), .A2(Plaintext[39]), .Z(n18649) );
  INV_X1 U24215 ( .I(Plaintext[37]), .ZN(n18348) );
  INV_X1 U24216 ( .I(Plaintext[30]), .ZN(n18350) );
  INV_X1 U24220 ( .I(Plaintext[8]), .ZN(n18354) );
  XOR2_X1 U24222 ( .A1(Key[11]), .A2(Plaintext[11]), .Z(n18674) );
  INV_X1 U24223 ( .I(Plaintext[18]), .ZN(n18356) );
  XOR2_X1 U24224 ( .A1(Key[21]), .A2(Plaintext[21]), .Z(n18357) );
  NAND2_X1 U24226 ( .A1(n18793), .A2(n26810), .ZN(n18361) );
  INV_X1 U24227 ( .I(Plaintext[48]), .ZN(n18364) );
  INV_X1 U24228 ( .I(Plaintext[49]), .ZN(n18365) );
  XOR2_X1 U24230 ( .A1(Key[42]), .A2(Plaintext[42]), .Z(n18811) );
  OAI21_X1 U24231 ( .A1(n8422), .A2(n18779), .B(n6215), .ZN(n18368) );
  NAND2_X1 U24232 ( .A1(n18368), .A2(n18618), .ZN(n18372) );
  NOR2_X1 U24235 ( .A1(n12074), .A2(n18642), .ZN(n18375) );
  NAND2_X1 U24236 ( .A1(n18378), .A2(n18377), .ZN(n18379) );
  INV_X1 U24237 ( .I(Plaintext[118]), .ZN(n18382) );
  NOR2_X1 U24238 ( .A1(n956), .A2(n18459), .ZN(n18387) );
  XOR2_X1 U24241 ( .A1(Key[113]), .A2(Plaintext[113]), .Z(n18696) );
  XOR2_X1 U24242 ( .A1(Key[108]), .A2(Plaintext[108]), .Z(n18831) );
  XOR2_X1 U24243 ( .A1(Key[109]), .A2(Plaintext[109]), .Z(n18700) );
  XOR2_X1 U24245 ( .A1(Key[123]), .A2(Plaintext[123]), .Z(n18429) );
  INV_X1 U24246 ( .I(Plaintext[120]), .ZN(n18393) );
  INV_X1 U24249 ( .I(Plaintext[3]), .ZN(n18395) );
  XOR2_X1 U24250 ( .A1(n18395), .A2(Key[3]), .Z(n18888) );
  XOR2_X1 U24251 ( .A1(Key[1]), .A2(Plaintext[1]), .Z(n18660) );
  INV_X1 U24252 ( .I(Plaintext[183]), .ZN(n18396) );
  XOR2_X1 U24254 ( .A1(Key[181]), .A2(Plaintext[181]), .Z(n18688) );
  INV_X1 U24255 ( .I(Plaintext[184]), .ZN(n18398) );
  XOR2_X1 U24256 ( .A1(Key[187]), .A2(Plaintext[187]), .Z(n18844) );
  INV_X2 U24257 ( .I(n18844), .ZN(n18681) );
  XOR2_X1 U24258 ( .A1(Key[173]), .A2(Plaintext[173]), .Z(n18402) );
  INV_X1 U24259 ( .I(Plaintext[172]), .ZN(n18401) );
  XOR2_X1 U24261 ( .A1(Key[167]), .A2(Plaintext[167]), .Z(n18861) );
  XOR2_X1 U24262 ( .A1(Key[162]), .A2(Plaintext[162]), .Z(n18862) );
  INV_X1 U24263 ( .I(Plaintext[163]), .ZN(n18404) );
  NAND2_X1 U24265 ( .A1(n10182), .A2(n18101), .ZN(n18406) );
  NAND2_X1 U24267 ( .A1(n31821), .A2(n18726), .ZN(n18408) );
  NAND3_X1 U24274 ( .A1(n18720), .A2(n16614), .A3(n8411), .ZN(n18416) );
  NAND2_X2 U24275 ( .A1(n18417), .A2(n18416), .ZN(n19318) );
  NAND2_X1 U24276 ( .A1(n33432), .A2(n19318), .ZN(n18418) );
  NAND3_X1 U24277 ( .A1(n19321), .A2(n18419), .A3(n18418), .ZN(n18420) );
  NOR2_X1 U24278 ( .A1(n19158), .A2(n14811), .ZN(n18425) );
  INV_X1 U24280 ( .I(n18831), .ZN(n18427) );
  INV_X1 U24281 ( .I(n18434), .ZN(n18746) );
  NAND2_X1 U24282 ( .A1(n8208), .A2(n6359), .ZN(n18437) );
  NOR2_X1 U24284 ( .A1(n18446), .A2(n18797), .ZN(n18444) );
  NAND2_X1 U24287 ( .A1(n18454), .A2(n17725), .ZN(n18456) );
  NOR2_X1 U24288 ( .A1(n18456), .A2(n18455), .ZN(n18458) );
  NOR2_X1 U24289 ( .A1(n18995), .A2(n18976), .ZN(n18468) );
  NOR2_X1 U24292 ( .A1(n18994), .A2(n100), .ZN(n18467) );
  NOR2_X1 U24294 ( .A1(n18006), .A2(n18699), .ZN(n18471) );
  NAND2_X1 U24298 ( .A1(n16585), .A2(n18811), .ZN(n18479) );
  NOR3_X1 U24300 ( .A1(n18481), .A2(n17597), .A3(n14093), .ZN(n18482) );
  NOR2_X1 U24301 ( .A1(n16417), .A2(n10080), .ZN(n18483) );
  NAND2_X1 U24302 ( .A1(n18601), .A2(n18755), .ZN(n18501) );
  NAND2_X1 U24303 ( .A1(n18761), .A2(n18605), .ZN(n18500) );
  AOI21_X1 U24304 ( .A1(n18501), .A2(n18500), .B(n27940), .ZN(n18502) );
  OR2_X1 U24305 ( .A1(n18899), .A2(n19088), .Z(n18504) );
  NOR2_X1 U24306 ( .A1(n17516), .A2(n15888), .ZN(n18507) );
  NAND2_X1 U24308 ( .A1(n16732), .A2(n33941), .ZN(n18512) );
  NOR2_X1 U24310 ( .A1(n18845), .A2(n18731), .ZN(n18520) );
  OAI21_X1 U24311 ( .A1(n957), .A2(n18520), .B(n18519), .ZN(n18524) );
  NOR2_X1 U24312 ( .A1(n17184), .A2(n18847), .ZN(n18521) );
  NAND2_X1 U24316 ( .A1(n18704), .A2(n18743), .ZN(n18536) );
  NAND2_X1 U24320 ( .A1(n18349), .A2(n18548), .ZN(n18550) );
  MUX2_X1 U24321 ( .I0(n18550), .I1(n18549), .S(n17114), .Z(n18551) );
  AOI21_X1 U24323 ( .A1(n18559), .A2(n18623), .B(n27129), .ZN(n18561) );
  NAND2_X1 U24324 ( .A1(n18774), .A2(n18771), .ZN(n18560) );
  NOR2_X1 U24329 ( .A1(n18848), .A2(n17030), .ZN(n18596) );
  NOR2_X1 U24330 ( .A1(n18402), .A2(n18846), .ZN(n18595) );
  INV_X1 U24332 ( .I(n19158), .ZN(n18599) );
  OAI21_X1 U24333 ( .A1(n18599), .A2(n14812), .B(n12548), .ZN(n18600) );
  NOR2_X1 U24335 ( .A1(n18618), .A2(n1430), .ZN(n18619) );
  NOR2_X1 U24336 ( .A1(n13254), .A2(n17937), .ZN(n18627) );
  INV_X1 U24337 ( .I(n18821), .ZN(n18632) );
  NOR2_X1 U24341 ( .A1(n18683), .A2(n5700), .ZN(n18651) );
  AOI22_X1 U24343 ( .A1(n18798), .A2(n31724), .B1(n18797), .B2(n18655), .ZN(
        n18656) );
  NOR2_X1 U24344 ( .A1(n18656), .A2(n16420), .ZN(n18657) );
  AOI21_X1 U24345 ( .A1(n31971), .A2(n28675), .B(n18687), .ZN(n18664) );
  NOR2_X1 U24346 ( .A1(n18866), .A2(n18871), .ZN(n18663) );
  NOR2_X1 U24347 ( .A1(n18664), .A2(n18663), .ZN(n18666) );
  NAND2_X1 U24351 ( .A1(n18692), .A2(n711), .ZN(n18693) );
  NAND2_X1 U24354 ( .A1(n18853), .A2(n15211), .ZN(n18719) );
  AOI21_X1 U24355 ( .A1(n18720), .A2(n16614), .B(n18307), .ZN(n18721) );
  NOR2_X1 U24358 ( .A1(n18736), .A2(n17687), .ZN(n18741) );
  NOR2_X1 U24359 ( .A1(n18747), .A2(n18742), .ZN(n18744) );
  NAND2_X1 U24360 ( .A1(n18747), .A2(n18746), .ZN(n18748) );
  NAND2_X1 U24362 ( .A1(n14093), .A2(n18755), .ZN(n18757) );
  NAND2_X1 U24364 ( .A1(n18762), .A2(n18761), .ZN(n19095) );
  NOR2_X1 U24365 ( .A1(n18775), .A2(n18770), .ZN(n18772) );
  NAND2_X1 U24367 ( .A1(n31095), .A2(n1430), .ZN(n18781) );
  NAND2_X1 U24369 ( .A1(n18798), .A2(n18797), .ZN(n18799) );
  XOR2_X1 U24371 ( .A1(n9665), .A2(n24869), .Z(n18814) );
  NOR2_X1 U24373 ( .A1(n785), .A2(n18515), .ZN(n18819) );
  NAND2_X1 U24374 ( .A1(n18819), .A2(n16393), .ZN(n19041) );
  NOR2_X1 U24375 ( .A1(n171), .A2(n4868), .ZN(n18825) );
  NAND2_X1 U24376 ( .A1(n18829), .A2(n18827), .ZN(n18828) );
  INV_X1 U24378 ( .I(n18921), .ZN(n18836) );
  NAND3_X1 U24379 ( .A1(n32784), .A2(n18836), .A3(n31324), .ZN(n18838) );
  NOR2_X1 U24380 ( .A1(n18848), .A2(n18847), .ZN(n18851) );
  XOR2_X1 U24385 ( .A1(n29030), .A2(n16454), .Z(n18898) );
  NAND2_X1 U24387 ( .A1(n19315), .A2(n825), .ZN(n18904) );
  XOR2_X1 U24388 ( .A1(n32262), .A2(n25038), .Z(n18915) );
  NOR2_X1 U24390 ( .A1(n28935), .A2(n18923), .ZN(n18925) );
  XOR2_X1 U24392 ( .A1(n28806), .A2(n25910), .Z(n18932) );
  NAND3_X1 U24394 ( .A1(n30959), .A2(n18939), .A3(n31949), .ZN(n18940) );
  XOR2_X1 U24396 ( .A1(n30443), .A2(n25519), .Z(n18948) );
  NOR2_X1 U24402 ( .A1(n31850), .A2(n16288), .ZN(n18984) );
  NOR2_X1 U24403 ( .A1(n14498), .A2(n18990), .ZN(n18989) );
  INV_X1 U24407 ( .I(n13925), .ZN(n19017) );
  NAND3_X1 U24411 ( .A1(n10124), .A2(n745), .A3(n19196), .ZN(n19024) );
  NAND2_X1 U24413 ( .A1(n14130), .A2(n19202), .ZN(n19028) );
  NAND2_X1 U24414 ( .A1(n19301), .A2(n26600), .ZN(n19027) );
  NAND3_X1 U24415 ( .A1(n19028), .A2(n730), .A3(n19027), .ZN(n19031) );
  NOR2_X1 U24416 ( .A1(n16354), .A2(n16093), .ZN(n19029) );
  INV_X1 U24417 ( .I(n19040), .ZN(n19045) );
  INV_X1 U24418 ( .I(n19041), .ZN(n19044) );
  INV_X1 U24419 ( .I(n19042), .ZN(n19043) );
  NOR3_X1 U24420 ( .A1(n19045), .A2(n19044), .A3(n19043), .ZN(n19047) );
  NOR3_X1 U24422 ( .A1(n1053), .A2(n19109), .A3(n19063), .ZN(n19064) );
  NOR2_X1 U24424 ( .A1(n19318), .A2(n19275), .ZN(n19068) );
  NOR2_X1 U24425 ( .A1(n19317), .A2(n30894), .ZN(n19067) );
  INV_X1 U24426 ( .I(n19356), .ZN(n19069) );
  NAND2_X1 U24427 ( .A1(n19069), .A2(n6516), .ZN(n19071) );
  NAND2_X1 U24428 ( .A1(n15842), .A2(n6516), .ZN(n19070) );
  AOI22_X1 U24429 ( .A1(n19071), .A2(n19281), .B1(n19070), .B2(n19354), .ZN(
        n19072) );
  INV_X1 U24432 ( .I(n19094), .ZN(n19098) );
  AOI22_X1 U24433 ( .A1(n19126), .A2(n31850), .B1(n19125), .B2(n7968), .ZN(
        n19131) );
  XOR2_X1 U24434 ( .A1(n19651), .A2(n16727), .Z(n19447) );
  NOR2_X1 U24435 ( .A1(n7810), .A2(n1379), .ZN(n19134) );
  OAI21_X1 U24437 ( .A1(n19137), .A2(n744), .B(n25971), .ZN(n19141) );
  NOR2_X1 U24438 ( .A1(n19257), .A2(n19258), .ZN(n19139) );
  NOR2_X1 U24439 ( .A1(n19255), .A2(n19143), .ZN(n19144) );
  NAND2_X1 U24440 ( .A1(n4747), .A2(n25961), .ZN(n19150) );
  NAND2_X1 U24442 ( .A1(n16007), .A2(n19160), .ZN(n19161) );
  XOR2_X1 U24445 ( .A1(n19474), .A2(n16561), .Z(n19193) );
  XOR2_X1 U24446 ( .A1(n19384), .A2(n25815), .Z(n19211) );
  MUX2_X1 U24448 ( .I0(n19275), .I1(n30894), .S(n19318), .Z(n19233) );
  NAND2_X1 U24449 ( .A1(n11940), .A2(n26603), .ZN(n19240) );
  NAND3_X1 U24450 ( .A1(n19243), .A2(n19242), .A3(n877), .ZN(n19246) );
  MUX2_X1 U24455 ( .I0(n19318), .I1(n27132), .S(n19275), .Z(n19277) );
  NAND2_X1 U24456 ( .A1(n19322), .A2(n19320), .ZN(n19276) );
  OAI21_X2 U24457 ( .A1(n19278), .A2(n19277), .B(n19276), .ZN(n19641) );
  INV_X1 U24459 ( .I(n19292), .ZN(n19293) );
  OAI21_X1 U24460 ( .A1(n746), .A2(n19295), .B(n19294), .ZN(n19296) );
  NOR2_X1 U24462 ( .A1(n19302), .A2(n19301), .ZN(n19303) );
  XOR2_X1 U24466 ( .A1(n19412), .A2(n15117), .Z(n19342) );
  XOR2_X1 U24467 ( .A1(n19625), .A2(n25074), .Z(n19344) );
  XOR2_X1 U24468 ( .A1(n11218), .A2(n19344), .Z(n19345) );
  INV_X1 U24470 ( .I(n19349), .ZN(n19347) );
  NAND2_X1 U24471 ( .A1(n19347), .A2(n19346), .ZN(n19351) );
  NAND2_X1 U24472 ( .A1(n19349), .A2(n27941), .ZN(n19350) );
  NAND2_X1 U24474 ( .A1(n19361), .A2(n16444), .ZN(n19362) );
  NAND2_X1 U24475 ( .A1(n19363), .A2(n19362), .ZN(n19366) );
  XOR2_X1 U24477 ( .A1(n30212), .A2(n25929), .Z(n19372) );
  XOR2_X1 U24478 ( .A1(n19373), .A2(n19372), .Z(n19374) );
  XOR2_X1 U24483 ( .A1(n19630), .A2(n16550), .Z(n19390) );
  XOR2_X1 U24484 ( .A1(n19755), .A2(n16619), .Z(n19394) );
  XOR2_X1 U24486 ( .A1(n15028), .A2(n25720), .Z(n19397) );
  XOR2_X1 U24487 ( .A1(n19644), .A2(n24231), .Z(n19401) );
  XOR2_X1 U24488 ( .A1(n19405), .A2(n19549), .Z(n19407) );
  XOR2_X1 U24489 ( .A1(n19409), .A2(n19754), .Z(n19411) );
  XOR2_X1 U24491 ( .A1(n19412), .A2(n19589), .Z(n19507) );
  XOR2_X1 U24492 ( .A1(n29890), .A2(n16423), .Z(n19413) );
  XOR2_X1 U24493 ( .A1(n19414), .A2(n19415), .Z(n19419) );
  NAND3_X1 U24494 ( .A1(n29156), .A2(n19799), .A3(n19886), .ZN(n19422) );
  XOR2_X1 U24495 ( .A1(n19416), .A2(n25358), .Z(n19417) );
  XOR2_X1 U24497 ( .A1(n19684), .A2(n19427), .Z(n19428) );
  XOR2_X1 U24498 ( .A1(n19429), .A2(n19428), .Z(n19796) );
  XOR2_X1 U24500 ( .A1(n19711), .A2(n19434), .Z(n19435) );
  NAND3_X1 U24504 ( .A1(n25997), .A2(n12038), .A3(n11913), .ZN(n19460) );
  XOR2_X1 U24505 ( .A1(n19649), .A2(n25722), .Z(n19465) );
  XOR2_X1 U24506 ( .A1(n16138), .A2(n16604), .Z(n19471) );
  XOR2_X1 U24508 ( .A1(n15787), .A2(n25079), .Z(n19487) );
  XOR2_X1 U24509 ( .A1(n19509), .A2(n16390), .Z(n19496) );
  XOR2_X1 U24510 ( .A1(n19498), .A2(n19524), .Z(n19500) );
  XOR2_X1 U24511 ( .A1(n28399), .A2(n16653), .Z(n19501) );
  INV_X1 U24512 ( .I(Key[2]), .ZN(n24831) );
  XOR2_X1 U24514 ( .A1(n19508), .A2(n34077), .Z(n19511) );
  XOR2_X1 U24515 ( .A1(n19509), .A2(n24895), .Z(n19510) );
  XOR2_X1 U24516 ( .A1(n19511), .A2(n19510), .Z(n19512) );
  XOR2_X1 U24517 ( .A1(n19755), .A2(n24833), .Z(n19516) );
  XOR2_X1 U24519 ( .A1(n19764), .A2(n19524), .Z(n19525) );
  XOR2_X1 U24520 ( .A1(n19699), .A2(n19525), .Z(n19526) );
  INV_X1 U24521 ( .I(n19530), .ZN(n19531) );
  INV_X1 U24522 ( .I(n19833), .ZN(n20040) );
  OAI21_X1 U24523 ( .A1(n20040), .A2(n1169), .B(n19834), .ZN(n19534) );
  XOR2_X1 U24524 ( .A1(n19736), .A2(n19539), .Z(n19540) );
  XOR2_X1 U24527 ( .A1(n19754), .A2(n16634), .Z(n19559) );
  XOR2_X1 U24528 ( .A1(n30766), .A2(n25554), .Z(n19573) );
  XOR2_X1 U24529 ( .A1(n19589), .A2(n24738), .Z(n19590) );
  XOR2_X1 U24530 ( .A1(n19591), .A2(n19590), .Z(n19596) );
  XOR2_X1 U24531 ( .A1(n15844), .A2(n19592), .Z(n19593) );
  XOR2_X1 U24532 ( .A1(n19594), .A2(n19593), .Z(n19595) );
  XOR2_X1 U24534 ( .A1(n19676), .A2(n25641), .Z(n19602) );
  INV_X1 U24535 ( .I(n19603), .ZN(n19607) );
  AOI22_X1 U24536 ( .A1(n19607), .A2(n19606), .B1(n19605), .B2(n19604), .ZN(
        n19609) );
  XOR2_X1 U24537 ( .A1(n29718), .A2(n19609), .Z(n19610) );
  XOR2_X1 U24538 ( .A1(n19611), .A2(n19610), .Z(n19612) );
  XOR2_X1 U24539 ( .A1(n19612), .A2(n19613), .Z(n19829) );
  XOR2_X1 U24540 ( .A1(n12048), .A2(n16530), .Z(n19615) );
  XOR2_X1 U24543 ( .A1(n30411), .A2(n19649), .Z(n19653) );
  XOR2_X1 U24545 ( .A1(n32697), .A2(n25436), .Z(n19655) );
  XOR2_X1 U24549 ( .A1(n19661), .A2(n24417), .Z(n19663) );
  NAND2_X1 U24554 ( .A1(n18199), .A2(n19899), .ZN(n20107) );
  XOR2_X1 U24556 ( .A1(n19682), .A2(n25091), .Z(n19683) );
  XOR2_X1 U24557 ( .A1(n19684), .A2(n19683), .Z(n19685) );
  XOR2_X1 U24558 ( .A1(n32271), .A2(n19691), .Z(n19694) );
  XOR2_X1 U24560 ( .A1(n19696), .A2(n25610), .Z(n19697) );
  XOR2_X1 U24562 ( .A1(n19712), .A2(n16662), .Z(n19713) );
  INV_X1 U24563 ( .I(Key[27]), .ZN(n19718) );
  XOR2_X1 U24569 ( .A1(n19751), .A2(n19750), .Z(n19752) );
  OAI21_X1 U24570 ( .A1(n31683), .A2(n26368), .B(n20112), .ZN(n19761) );
  XOR2_X1 U24573 ( .A1(n19771), .A2(n19770), .Z(n19777) );
  XOR2_X1 U24574 ( .A1(n19773), .A2(n25751), .Z(n19774) );
  XOR2_X1 U24575 ( .A1(n19775), .A2(n19774), .Z(n19776) );
  XOR2_X1 U24576 ( .A1(n19777), .A2(n19776), .Z(n20083) );
  XOR2_X1 U24577 ( .A1(n8571), .A2(n25040), .Z(n19786) );
  AOI21_X1 U24578 ( .A1(n19789), .A2(n20085), .B(n16664), .ZN(n19790) );
  NAND3_X1 U24580 ( .A1(n20034), .A2(n20032), .A3(n19971), .ZN(n19810) );
  INV_X1 U24582 ( .I(n20083), .ZN(n20007) );
  NOR2_X1 U24585 ( .A1(n15394), .A2(n17299), .ZN(n19831) );
  NAND2_X1 U24594 ( .A1(n27600), .A2(n11453), .ZN(n19865) );
  AOI21_X2 U24597 ( .A1(n19872), .A2(n821), .B(n19871), .ZN(n20521) );
  NAND2_X1 U24598 ( .A1(n29339), .A2(n16491), .ZN(n19875) );
  INV_X1 U24599 ( .I(n19933), .ZN(n19876) );
  NAND3_X1 U24601 ( .A1(n2606), .A2(n20096), .A3(n3915), .ZN(n20293) );
  MUX2_X1 U24605 ( .I0(n19896), .I1(n12682), .S(n20136), .Z(n20229) );
  NAND2_X1 U24606 ( .A1(n16595), .A2(n20021), .ZN(n19897) );
  NOR3_X1 U24609 ( .A1(n19912), .A2(n19913), .A3(n12142), .ZN(n19911) );
  INV_X1 U24611 ( .I(n8259), .ZN(n19917) );
  NOR2_X1 U24617 ( .A1(n4254), .A2(n20486), .ZN(n19957) );
  INV_X1 U24619 ( .I(n20631), .ZN(n19972) );
  NAND2_X1 U24620 ( .A1(n19965), .A2(n20018), .ZN(n19968) );
  AOI21_X1 U24621 ( .A1(n20033), .A2(n2795), .B(n16243), .ZN(n19970) );
  NAND2_X1 U24623 ( .A1(n19819), .A2(n32745), .ZN(n19975) );
  XOR2_X1 U24629 ( .A1(n20693), .A2(n16602), .Z(n20005) );
  XOR2_X1 U24630 ( .A1(n20722), .A2(n20005), .Z(n20050) );
  OAI21_X1 U24631 ( .A1(n20020), .A2(n20019), .B(n20119), .ZN(n20024) );
  INV_X1 U24638 ( .I(n20060), .ZN(n20063) );
  INV_X1 U24640 ( .I(n20070), .ZN(n20073) );
  MUX2_X1 U24644 ( .I0(n20122), .I1(n20121), .S(n14334), .Z(n20127) );
  NOR2_X2 U24645 ( .A1(n20127), .A2(n20126), .ZN(n20460) );
  NAND2_X1 U24650 ( .A1(n20266), .A2(n28376), .ZN(n20163) );
  XOR2_X1 U24651 ( .A1(n20868), .A2(n20166), .Z(n20167) );
  XOR2_X1 U24652 ( .A1(n20168), .A2(n20167), .Z(n21258) );
  MUX2_X1 U24653 ( .I0(n13768), .I1(n16374), .S(n20556), .Z(n20169) );
  NAND2_X1 U24656 ( .A1(n28414), .A2(n20499), .ZN(n20175) );
  INV_X1 U24659 ( .I(n20188), .ZN(n20193) );
  INV_X1 U24660 ( .I(n20190), .ZN(n20192) );
  INV_X1 U24663 ( .I(n20209), .ZN(n20210) );
  NAND2_X1 U24666 ( .A1(n4254), .A2(n20221), .ZN(n20222) );
  XOR2_X1 U24667 ( .A1(n20729), .A2(n20784), .Z(n20226) );
  XOR2_X1 U24668 ( .A1(n20715), .A2(n16548), .Z(n20225) );
  NAND3_X1 U24669 ( .A1(n20520), .A2(n16218), .A3(n20556), .ZN(n20237) );
  XOR2_X1 U24670 ( .A1(n20733), .A2(n25252), .Z(n20241) );
  INV_X1 U24672 ( .I(n16050), .ZN(n20255) );
  NAND2_X1 U24673 ( .A1(n16951), .A2(n11182), .ZN(n20256) );
  AOI22_X1 U24675 ( .A1(n20651), .A2(n20271), .B1(n28575), .B2(n20270), .ZN(
        n20272) );
  MUX2_X1 U24676 ( .I0(n20273), .I1(n1157), .S(n15434), .Z(n20275) );
  INV_X1 U24679 ( .I(n20280), .ZN(n20281) );
  INV_X1 U24681 ( .I(n16515), .ZN(n20284) );
  NAND4_X1 U24682 ( .A1(n20294), .A2(n20291), .A3(n20292), .A4(n20293), .ZN(
        n20296) );
  NAND2_X1 U24685 ( .A1(n12872), .A2(n6230), .ZN(n20314) );
  XOR2_X1 U24686 ( .A1(n3009), .A2(n16619), .Z(n20318) );
  NAND3_X1 U24687 ( .A1(n818), .A2(n710), .A3(n20335), .ZN(n20336) );
  XOR2_X1 U24690 ( .A1(n33969), .A2(n25358), .Z(n20356) );
  XOR2_X1 U24691 ( .A1(n21038), .A2(n20356), .Z(n20357) );
  INV_X1 U24695 ( .I(n25428), .ZN(n20389) );
  AOI21_X1 U24703 ( .A1(n20562), .A2(n30931), .B(n20523), .ZN(n20415) );
  OAI21_X2 U24706 ( .A1(n20422), .A2(n20421), .B(n20420), .ZN(n21043) );
  NAND2_X1 U24707 ( .A1(n17329), .A2(n4647), .ZN(n20424) );
  INV_X1 U24708 ( .I(n20431), .ZN(n20432) );
  INV_X1 U24709 ( .I(n20433), .ZN(n20434) );
  INV_X1 U24710 ( .I(n20495), .ZN(n20440) );
  NAND2_X1 U24712 ( .A1(n4468), .A2(n31768), .ZN(n20446) );
  INV_X1 U24714 ( .I(n20453), .ZN(n20456) );
  NAND3_X1 U24716 ( .A1(n29695), .A2(n20489), .A3(n28812), .ZN(n20490) );
  NOR2_X1 U24717 ( .A1(n20495), .A2(n20494), .ZN(n20496) );
  XOR2_X1 U24719 ( .A1(n20920), .A2(n7705), .Z(n20513) );
  XOR2_X1 U24720 ( .A1(n20824), .A2(n16581), .Z(n20512) );
  XOR2_X1 U24721 ( .A1(n20512), .A2(n20513), .Z(n20514) );
  XOR2_X1 U24724 ( .A1(n21046), .A2(n16497), .Z(n20542) );
  XOR2_X1 U24725 ( .A1(n20586), .A2(n2616), .Z(n20588) );
  NAND4_X1 U24732 ( .A1(n20625), .A2(n20624), .A3(n20623), .A4(n20622), .ZN(
        n20626) );
  XOR2_X1 U24735 ( .A1(n32162), .A2(n25126), .Z(n20640) );
  XOR2_X1 U24736 ( .A1(n20690), .A2(n16504), .Z(n20642) );
  XOR2_X1 U24737 ( .A1(n32791), .A2(n24861), .Z(n20645) );
  XOR2_X1 U24738 ( .A1(n20984), .A2(n20647), .Z(n20649) );
  XOR2_X1 U24741 ( .A1(n20658), .A2(n24417), .Z(n20659) );
  XOR2_X1 U24742 ( .A1(n20660), .A2(n20659), .Z(n20661) );
  XOR2_X1 U24743 ( .A1(n20857), .A2(n25783), .Z(n20663) );
  XOR2_X1 U24746 ( .A1(n20747), .A2(n8487), .Z(n20667) );
  XOR2_X1 U24748 ( .A1(n5348), .A2(n25191), .Z(n20672) );
  XOR2_X1 U24749 ( .A1(n20673), .A2(n20672), .Z(n20675) );
  XOR2_X1 U24751 ( .A1(n21016), .A2(n16697), .Z(n20682) );
  XOR2_X1 U24753 ( .A1(n20775), .A2(n25054), .Z(n20694) );
  XOR2_X1 U24754 ( .A1(n20695), .A2(n20694), .Z(n20696) );
  XOR2_X1 U24755 ( .A1(n25619), .A2(n20720), .Z(n20697) );
  XOR2_X1 U24757 ( .A1(n20743), .A2(n20702), .Z(n20704) );
  XOR2_X1 U24758 ( .A1(n20848), .A2(n24623), .Z(n20703) );
  XOR2_X1 U24759 ( .A1(n20837), .A2(n16604), .Z(n20706) );
  XOR2_X1 U24761 ( .A1(n10522), .A2(n20756), .Z(n20707) );
  XOR2_X1 U24762 ( .A1(n20851), .A2(n16578), .Z(n20719) );
  XOR2_X1 U24763 ( .A1(n20917), .A2(n20836), .Z(n20724) );
  XOR2_X1 U24764 ( .A1(n21029), .A2(n16671), .Z(n20731) );
  XOR2_X1 U24766 ( .A1(n21019), .A2(n25182), .Z(n20737) );
  INV_X1 U24768 ( .I(n23239), .ZN(n25213) );
  XOR2_X1 U24769 ( .A1(n32749), .A2(n16680), .Z(n20744) );
  XOR2_X1 U24770 ( .A1(n14132), .A2(n25728), .Z(n20749) );
  XOR2_X1 U24772 ( .A1(n21001), .A2(n24514), .Z(n20759) );
  XOR2_X1 U24775 ( .A1(n1342), .A2(n16555), .Z(n20770) );
  XOR2_X1 U24776 ( .A1(n20771), .A2(n20770), .Z(n20774) );
  INV_X1 U24778 ( .I(n21402), .ZN(n20795) );
  XOR2_X1 U24779 ( .A1(n29241), .A2(n18019), .Z(n20793) );
  XOR2_X1 U24784 ( .A1(n30219), .A2(n25288), .Z(n20815) );
  XOR2_X1 U24789 ( .A1(n28864), .A2(n20839), .Z(n20840) );
  XOR2_X1 U24790 ( .A1(n20841), .A2(n20840), .Z(n20846) );
  XOR2_X1 U24791 ( .A1(n20843), .A2(n24907), .Z(n20844) );
  XOR2_X1 U24792 ( .A1(n20919), .A2(n20844), .Z(n20845) );
  XOR2_X1 U24793 ( .A1(n20845), .A2(n20846), .Z(n21389) );
  XOR2_X1 U24795 ( .A1(n21024), .A2(n20183), .Z(n20865) );
  XOR2_X1 U24796 ( .A1(n20865), .A2(n20864), .Z(n20866) );
  NAND2_X1 U24797 ( .A1(n20880), .A2(n6408), .ZN(n20875) );
  XOR2_X1 U24800 ( .A1(n1023), .A2(n25040), .Z(n20908) );
  NOR2_X1 U24802 ( .A1(n20909), .A2(n31760), .ZN(n20910) );
  XOR2_X1 U24803 ( .A1(n32478), .A2(n24992), .Z(n20922) );
  XOR2_X1 U24804 ( .A1(n20926), .A2(n16575), .Z(n20927) );
  AOI21_X1 U24805 ( .A1(n21363), .A2(n20932), .B(n21182), .ZN(n20934) );
  NAND2_X1 U24806 ( .A1(n21363), .A2(n27382), .ZN(n20933) );
  NOR2_X1 U24808 ( .A1(n27773), .A2(n20945), .ZN(n20944) );
  XOR2_X1 U24812 ( .A1(n20975), .A2(n25641), .Z(n20976) );
  XOR2_X1 U24813 ( .A1(n20985), .A2(n25064), .Z(n20986) );
  XOR2_X1 U24814 ( .A1(n28687), .A2(n24999), .Z(n20995) );
  XOR2_X1 U24815 ( .A1(n20996), .A2(n20997), .Z(n20998) );
  XOR2_X1 U24817 ( .A1(n21001), .A2(n24374), .Z(n21002) );
  XOR2_X1 U24818 ( .A1(n21003), .A2(n21002), .Z(n21004) );
  XOR2_X1 U24819 ( .A1(n21005), .A2(n21004), .Z(n21068) );
  INV_X1 U24820 ( .I(n21068), .ZN(n21424) );
  XOR2_X1 U24821 ( .A1(n21029), .A2(n25506), .Z(n21030) );
  XOR2_X1 U24822 ( .A1(n21031), .A2(n21030), .Z(n21032) );
  NOR2_X1 U24825 ( .A1(n16034), .A2(n8490), .ZN(n21066) );
  NOR2_X1 U24827 ( .A1(n5480), .A2(n21075), .ZN(n21076) );
  NAND2_X1 U24828 ( .A1(n21160), .A2(n4145), .ZN(n21088) );
  MUX2_X1 U24829 ( .I0(n21088), .I1(n32452), .S(n26777), .Z(n21090) );
  NAND2_X1 U24831 ( .A1(n21206), .A2(n15874), .ZN(n21098) );
  NAND3_X1 U24832 ( .A1(n21289), .A2(n21143), .A3(n21396), .ZN(n21097) );
  INV_X1 U24833 ( .I(n21100), .ZN(n21303) );
  NAND2_X1 U24837 ( .A1(n925), .A2(n6451), .ZN(n21110) );
  INV_X1 U24838 ( .I(n24514), .ZN(n25849) );
  XOR2_X1 U24839 ( .A1(n8291), .A2(n25849), .Z(n21112) );
  NAND2_X1 U24841 ( .A1(n11187), .A2(n4381), .ZN(n21118) );
  NAND2_X1 U24842 ( .A1(n21306), .A2(n21307), .ZN(n21129) );
  NAND3_X1 U24845 ( .A1(n16034), .A2(n28642), .A3(n31965), .ZN(n21137) );
  NAND2_X1 U24846 ( .A1(n16222), .A2(n21592), .ZN(n21594) );
  NOR2_X1 U24849 ( .A1(n28190), .A2(n21379), .ZN(n21159) );
  NAND2_X1 U24854 ( .A1(n21439), .A2(n17832), .ZN(n21226) );
  NOR2_X1 U24857 ( .A1(n9186), .A2(n21237), .ZN(n21634) );
  XOR2_X1 U24861 ( .A1(n22147), .A2(n16680), .Z(n21280) );
  NAND2_X1 U24862 ( .A1(n1312), .A2(n1136), .ZN(n21282) );
  MUX2_X1 U24866 ( .I0(n21305), .I1(n21304), .S(n21306), .Z(n21310) );
  NAND2_X1 U24875 ( .A1(n1328), .A2(n17416), .ZN(n21346) );
  NAND3_X1 U24877 ( .A1(n21340), .A2(n26542), .A3(n21339), .ZN(n21345) );
  NOR2_X1 U24880 ( .A1(n21369), .A2(n11966), .ZN(n21370) );
  NOR3_X1 U24883 ( .A1(n27711), .A2(n922), .A3(n6408), .ZN(n21385) );
  NAND2_X1 U24884 ( .A1(n21392), .A2(n21391), .ZN(n21393) );
  NAND2_X1 U24885 ( .A1(n8587), .A2(n812), .ZN(n21394) );
  MUX2_X1 U24890 ( .I0(n21469), .I1(n21467), .S(n21793), .Z(n21472) );
  NAND3_X1 U24892 ( .A1(n21470), .A2(n21469), .A3(n8079), .ZN(n21471) );
  NAND2_X1 U24893 ( .A1(n21933), .A2(n21932), .ZN(n21477) );
  NOR2_X1 U24895 ( .A1(n21934), .A2(n28895), .ZN(n21475) );
  MUX2_X1 U24899 ( .I0(n21613), .I1(n21482), .S(n21755), .Z(n21485) );
  INV_X1 U24900 ( .I(n31765), .ZN(n21487) );
  INV_X1 U24902 ( .I(n21497), .ZN(n21502) );
  INV_X1 U24903 ( .I(n21498), .ZN(n21501) );
  INV_X1 U24904 ( .I(n21499), .ZN(n21500) );
  NOR3_X1 U24905 ( .A1(n21502), .A2(n21501), .A3(n21500), .ZN(n21503) );
  NOR2_X1 U24912 ( .A1(n30677), .A2(n21532), .ZN(n21534) );
  NAND2_X1 U24914 ( .A1(n21539), .A2(n21857), .ZN(n21540) );
  XOR2_X1 U24917 ( .A1(n30495), .A2(n16705), .Z(n21582) );
  OAI21_X1 U24918 ( .A1(n31978), .A2(n21628), .B(n2217), .ZN(n21608) );
  INV_X1 U24919 ( .I(n21614), .ZN(n21615) );
  NOR2_X1 U24920 ( .A1(n21616), .A2(n21615), .ZN(n21621) );
  INV_X1 U24921 ( .I(n21617), .ZN(n21618) );
  NOR2_X1 U24922 ( .A1(n21619), .A2(n21618), .ZN(n21620) );
  INV_X1 U24924 ( .I(n21633), .ZN(n21635) );
  NOR2_X1 U24925 ( .A1(n21635), .A2(n21634), .ZN(n21639) );
  NAND4_X1 U24926 ( .A1(n31511), .A2(n21639), .A3(n21637), .A4(n21638), .ZN(
        n21640) );
  NAND2_X1 U24927 ( .A1(n30506), .A2(n15864), .ZN(n21648) );
  XOR2_X1 U24928 ( .A1(n3550), .A2(n25282), .Z(n21650) );
  XOR2_X1 U24929 ( .A1(n8291), .A2(n24992), .Z(n21658) );
  NAND3_X1 U24930 ( .A1(n21850), .A2(n21763), .A3(n15022), .ZN(n21684) );
  OAI21_X1 U24932 ( .A1(n26474), .A2(n21730), .B(n920), .ZN(n21731) );
  NAND2_X1 U24936 ( .A1(n27649), .A2(n21755), .ZN(n21753) );
  NAND2_X1 U24938 ( .A1(n12587), .A2(n21763), .ZN(n21760) );
  XOR2_X1 U24939 ( .A1(n22086), .A2(n16550), .Z(n21768) );
  NAND2_X1 U24942 ( .A1(n21811), .A2(n21808), .ZN(n21809) );
  XOR2_X1 U24943 ( .A1(n21916), .A2(n21813), .Z(n21814) );
  XOR2_X1 U24944 ( .A1(n21815), .A2(n21814), .Z(n22677) );
  INV_X1 U24945 ( .I(n21824), .ZN(n21825) );
  INV_X1 U24946 ( .I(n21826), .ZN(n21828) );
  INV_X1 U24947 ( .I(n21831), .ZN(n21836) );
  NOR2_X1 U24948 ( .A1(n11890), .A2(n25815), .ZN(n21833) );
  OAI21_X1 U24949 ( .A1(n1009), .A2(n15242), .B(n21833), .ZN(n21834) );
  OAI22_X1 U24950 ( .A1(n21836), .A2(n25815), .B1(n21835), .B2(n21834), .ZN(
        n21837) );
  AOI21_X1 U24951 ( .A1(n25815), .A2(n34016), .B(n21837), .ZN(n21838) );
  INV_X1 U24952 ( .I(n21857), .ZN(n21861) );
  XOR2_X1 U24955 ( .A1(n21875), .A2(n21874), .Z(n21881) );
  XOR2_X1 U24956 ( .A1(n21878), .A2(n21879), .Z(n21880) );
  XOR2_X1 U24959 ( .A1(n22188), .A2(n25827), .Z(n21884) );
  INV_X1 U24960 ( .I(n24417), .ZN(n24435) );
  XOR2_X1 U24961 ( .A1(n30306), .A2(n24435), .Z(n21887) );
  XOR2_X1 U24962 ( .A1(n16355), .A2(n22197), .Z(n21888) );
  XOR2_X1 U24963 ( .A1(n21923), .A2(n16687), .Z(n21893) );
  INV_X1 U24964 ( .I(n12785), .ZN(n21894) );
  XOR2_X1 U24969 ( .A1(n21906), .A2(n21905), .Z(n21907) );
  XOR2_X1 U24970 ( .A1(n22044), .A2(n24748), .Z(n21915) );
  XOR2_X1 U24975 ( .A1(n22111), .A2(n22018), .Z(n21939) );
  XOR2_X1 U24976 ( .A1(n21940), .A2(n21939), .Z(n21941) );
  XOR2_X1 U24978 ( .A1(n21948), .A2(n21947), .Z(n21950) );
  XOR2_X1 U24979 ( .A1(n27180), .A2(n25104), .Z(n21953) );
  NAND2_X1 U24980 ( .A1(n22641), .A2(n33594), .ZN(n21957) );
  XOR2_X1 U24981 ( .A1(n21959), .A2(n22123), .Z(n21960) );
  XOR2_X1 U24982 ( .A1(n22226), .A2(n18019), .Z(n21962) );
  XOR2_X1 U24983 ( .A1(n22295), .A2(n16555), .Z(n21967) );
  NAND2_X1 U24985 ( .A1(n28124), .A2(n22489), .ZN(n21972) );
  NAND2_X1 U24990 ( .A1(n21979), .A2(n16240), .ZN(n21980) );
  NAND3_X1 U24991 ( .A1(n33007), .A2(n33115), .A3(n17930), .ZN(n21983) );
  XOR2_X1 U24993 ( .A1(n30495), .A2(n25735), .Z(n21988) );
  XOR2_X1 U24994 ( .A1(n22291), .A2(n25465), .Z(n21999) );
  XOR2_X1 U24997 ( .A1(n22239), .A2(n16507), .Z(n22006) );
  XOR2_X1 U25002 ( .A1(n22145), .A2(n25856), .Z(n22022) );
  XOR2_X1 U25005 ( .A1(n22251), .A2(n16581), .Z(n22038) );
  XOR2_X1 U25006 ( .A1(n22039), .A2(n22038), .Z(n22040) );
  XOR2_X1 U25007 ( .A1(n26957), .A2(n16402), .Z(n22045) );
  NAND2_X1 U25009 ( .A1(n22741), .A2(n22780), .ZN(n22053) );
  XOR2_X1 U25010 ( .A1(n7477), .A2(n25519), .Z(n22057) );
  INV_X1 U25011 ( .I(n22185), .ZN(n22058) );
  XOR2_X1 U25012 ( .A1(n32885), .A2(n22058), .Z(n22060) );
  XOR2_X1 U25013 ( .A1(n28848), .A2(n25074), .Z(n22062) );
  XOR2_X1 U25019 ( .A1(n29011), .A2(n25500), .Z(n22083) );
  XOR2_X1 U25020 ( .A1(n32404), .A2(n22086), .Z(n22088) );
  XOR2_X1 U25021 ( .A1(n17555), .A2(n25373), .Z(n22087) );
  XOR2_X1 U25022 ( .A1(n22088), .A2(n22087), .Z(n22089) );
  XOR2_X1 U25023 ( .A1(n22090), .A2(n22089), .Z(n22662) );
  XOR2_X1 U25024 ( .A1(n22201), .A2(n25911), .Z(n22093) );
  XOR2_X1 U25025 ( .A1(n22093), .A2(n22259), .Z(n22094) );
  XOR2_X1 U25026 ( .A1(n16649), .A2(n27850), .Z(n22103) );
  XOR2_X1 U25027 ( .A1(n22104), .A2(n22103), .Z(n22107) );
  XOR2_X1 U25031 ( .A1(n22295), .A2(n16654), .Z(n22133) );
  XOR2_X1 U25034 ( .A1(n3550), .A2(n16666), .Z(n22146) );
  INV_X1 U25035 ( .I(n22579), .ZN(n22452) );
  XOR2_X1 U25036 ( .A1(n28848), .A2(n24966), .Z(n22151) );
  XOR2_X1 U25037 ( .A1(n22162), .A2(n25049), .Z(n22163) );
  XOR2_X1 U25038 ( .A1(n17555), .A2(n16674), .Z(n22174) );
  XOR2_X1 U25039 ( .A1(n22175), .A2(n22174), .Z(n22176) );
  XOR2_X1 U25042 ( .A1(n22318), .A2(n25071), .Z(n22181) );
  XOR2_X1 U25049 ( .A1(n22238), .A2(n16502), .Z(n22241) );
  MUX2_X1 U25051 ( .I0(n22254), .I1(n22253), .S(n28424), .Z(n22258) );
  XOR2_X1 U25052 ( .A1(n22260), .A2(n25783), .Z(n22261) );
  NOR2_X1 U25054 ( .A1(n28924), .A2(n32078), .ZN(n22297) );
  XOR2_X1 U25055 ( .A1(n22308), .A2(n25881), .Z(n22309) );
  XOR2_X1 U25056 ( .A1(n32154), .A2(n16655), .Z(n22319) );
  NOR2_X1 U25060 ( .A1(n22745), .A2(n27166), .ZN(n22328) );
  NAND2_X1 U25068 ( .A1(n11930), .A2(n22599), .ZN(n22356) );
  XOR2_X1 U25074 ( .A1(n23367), .A2(n25091), .Z(n22384) );
  XOR2_X1 U25075 ( .A1(n22385), .A2(n22384), .Z(n22386) );
  XOR2_X1 U25076 ( .A1(n22387), .A2(n22386), .Z(n22617) );
  AOI21_X1 U25079 ( .A1(n22408), .A2(n22534), .B(n909), .ZN(n22409) );
  NAND2_X1 U25081 ( .A1(n22644), .A2(n33594), .ZN(n22422) );
  NAND3_X1 U25084 ( .A1(n22604), .A2(n17960), .A3(n14728), .ZN(n22426) );
  NAND2_X1 U25085 ( .A1(n16503), .A2(n22923), .ZN(n22458) );
  NAND2_X1 U25086 ( .A1(n22460), .A2(n5379), .ZN(n22461) );
  NOR2_X1 U25090 ( .A1(n22681), .A2(n11926), .ZN(n22471) );
  NAND2_X1 U25092 ( .A1(n22546), .A2(n1282), .ZN(n22480) );
  OAI21_X1 U25094 ( .A1(n14493), .A2(n22689), .B(n15746), .ZN(n22498) );
  XOR2_X1 U25100 ( .A1(n9153), .A2(n25079), .Z(n22515) );
  XOR2_X1 U25101 ( .A1(n22516), .A2(n22515), .Z(n22517) );
  NAND2_X1 U25105 ( .A1(n22562), .A2(n16447), .ZN(n22561) );
  NAND2_X1 U25109 ( .A1(n22659), .A2(n22658), .ZN(n22575) );
  INV_X1 U25110 ( .I(n22806), .ZN(n22581) );
  NOR3_X1 U25111 ( .A1(n22724), .A2(n22581), .A3(n22723), .ZN(n22582) );
  XOR2_X1 U25114 ( .A1(n23393), .A2(n16551), .Z(n22616) );
  OAI21_X1 U25119 ( .A1(n14183), .A2(n23072), .B(n28970), .ZN(n22692) );
  INV_X1 U25121 ( .I(n22697), .ZN(n22698) );
  OAI21_X1 U25122 ( .A1(n7181), .A2(n7881), .B(n22827), .ZN(n22706) );
  XOR2_X1 U25123 ( .A1(n23328), .A2(n23363), .Z(n22711) );
  MUX2_X1 U25124 ( .I0(n30365), .I1(n26667), .S(n23100), .Z(n22710) );
  XOR2_X1 U25125 ( .A1(n22711), .A2(n8298), .Z(n22712) );
  XOR2_X1 U25126 ( .A1(n23230), .A2(n25428), .Z(n22719) );
  XOR2_X1 U25127 ( .A1(n23373), .A2(n22719), .Z(n22728) );
  NAND2_X1 U25128 ( .A1(n6012), .A2(n23109), .ZN(n22726) );
  MUX2_X1 U25134 ( .I0(n22740), .I1(n22739), .S(n3184), .Z(n22743) );
  MUX2_X1 U25136 ( .I0(n23583), .I1(n23745), .S(n23770), .Z(n22765) );
  NAND3_X1 U25138 ( .A1(n22757), .A2(n23042), .A3(n13474), .ZN(n22758) );
  XOR2_X1 U25143 ( .A1(n23274), .A2(n25038), .Z(n22799) );
  XOR2_X1 U25149 ( .A1(n23467), .A2(n25064), .Z(n22841) );
  INV_X1 U25152 ( .I(n3183), .ZN(n22888) );
  OAI21_X1 U25153 ( .A1(n29175), .A2(n3183), .B(n22849), .ZN(n22851) );
  XOR2_X1 U25157 ( .A1(n23258), .A2(n25610), .Z(n22867) );
  XOR2_X1 U25158 ( .A1(n23439), .A2(n23189), .Z(n22875) );
  XOR2_X1 U25159 ( .A1(n23331), .A2(n22875), .Z(n22877) );
  XOR2_X1 U25161 ( .A1(n23274), .A2(n16472), .Z(n22896) );
  NAND2_X1 U25165 ( .A1(n22921), .A2(n22920), .ZN(n22929) );
  INV_X1 U25166 ( .I(n22922), .ZN(n22928) );
  INV_X1 U25167 ( .I(n22923), .ZN(n22925) );
  OAI21_X1 U25168 ( .A1(n31267), .A2(n22925), .B(n22924), .ZN(n22927) );
  NOR3_X1 U25169 ( .A1(n22929), .A2(n22928), .A3(n22927), .ZN(n22931) );
  XOR2_X1 U25171 ( .A1(n23511), .A2(n23125), .Z(n22934) );
  XOR2_X1 U25172 ( .A1(n22935), .A2(n22934), .Z(n22936) );
  NAND2_X1 U25173 ( .A1(n22940), .A2(n27694), .ZN(n22942) );
  INV_X2 U25174 ( .I(n32860), .ZN(n23203) );
  XOR2_X1 U25175 ( .A1(n23203), .A2(n1067), .Z(n22954) );
  NOR2_X1 U25177 ( .A1(n14129), .A2(n22965), .ZN(n22966) );
  NAND2_X1 U25178 ( .A1(n31935), .A2(n28680), .ZN(n22996) );
  INV_X1 U25179 ( .I(n23007), .ZN(n23008) );
  INV_X1 U25180 ( .I(n23011), .ZN(n23012) );
  NOR2_X1 U25181 ( .A1(n23013), .A2(n23012), .ZN(n23014) );
  XOR2_X1 U25182 ( .A1(n7070), .A2(n721), .Z(n23023) );
  XOR2_X1 U25184 ( .A1(n29217), .A2(n24833), .Z(n23022) );
  XOR2_X1 U25185 ( .A1(n23023), .A2(n23022), .Z(n23024) );
  XOR2_X1 U25187 ( .A1(n8659), .A2(n23376), .Z(n23039) );
  XOR2_X1 U25188 ( .A1(n27875), .A2(n25554), .Z(n23038) );
  XOR2_X1 U25189 ( .A1(n23038), .A2(n23039), .Z(n23040) );
  NAND3_X1 U25190 ( .A1(n27612), .A2(n1108), .A3(n28277), .ZN(n23054) );
  NAND2_X1 U25191 ( .A1(n1269), .A2(n26231), .ZN(n23060) );
  XOR2_X1 U25194 ( .A1(n23420), .A2(n16423), .Z(n23076) );
  XOR2_X1 U25195 ( .A1(n23075), .A2(n23076), .Z(n23077) );
  NAND2_X1 U25197 ( .A1(n14602), .A2(n17639), .ZN(n23089) );
  XOR2_X1 U25200 ( .A1(n24992), .A2(n11891), .Z(n23118) );
  XOR2_X1 U25201 ( .A1(n23122), .A2(n32893), .Z(n23123) );
  XOR2_X1 U25204 ( .A1(n13321), .A2(n16697), .Z(n23139) );
  XOR2_X1 U25205 ( .A1(n23344), .A2(n23139), .Z(n23140) );
  XOR2_X1 U25207 ( .A1(n24953), .A2(n3519), .Z(n23146) );
  XOR2_X1 U25210 ( .A1(n27763), .A2(n16666), .Z(n23154) );
  INV_X1 U25211 ( .I(n23530), .ZN(n23162) );
  XOR2_X1 U25212 ( .A1(n32050), .A2(n23474), .Z(n23163) );
  NAND2_X1 U25216 ( .A1(n12658), .A2(n31796), .ZN(n23177) );
  OAI21_X1 U25217 ( .A1(n24385), .A2(n24383), .B(n24384), .ZN(n23179) );
  XOR2_X1 U25218 ( .A1(n23420), .A2(n24231), .Z(n23185) );
  XOR2_X1 U25222 ( .A1(n3868), .A2(n25324), .Z(n23198) );
  XOR2_X1 U25223 ( .A1(n23454), .A2(n23346), .Z(n23205) );
  XOR2_X1 U25225 ( .A1(n24759), .A2(n23211), .Z(n23212) );
  OAI21_X1 U25226 ( .A1(n757), .A2(n32998), .B(n23823), .ZN(n23223) );
  XOR2_X1 U25227 ( .A1(n23216), .A2(n24966), .Z(n23217) );
  XOR2_X1 U25228 ( .A1(n7045), .A2(n30315), .Z(n23226) );
  XOR2_X1 U25229 ( .A1(n23385), .A2(n23227), .Z(n23228) );
  XOR2_X1 U25230 ( .A1(n27875), .A2(n25282), .Z(n23231) );
  XOR2_X1 U25231 ( .A1(n32899), .A2(n16479), .Z(n23232) );
  XOR2_X1 U25233 ( .A1(n848), .A2(n25549), .Z(n23243) );
  XOR2_X1 U25234 ( .A1(n23250), .A2(n25910), .Z(n23251) );
  XOR2_X1 U25236 ( .A1(n24707), .A2(n11891), .Z(n23268) );
  XOR2_X1 U25237 ( .A1(n23298), .A2(n23268), .Z(n23269) );
  XOR2_X1 U25238 ( .A1(n5512), .A2(n5211), .Z(n23278) );
  XOR2_X1 U25239 ( .A1(n26656), .A2(n23287), .Z(n23288) );
  XOR2_X1 U25240 ( .A1(n27708), .A2(n23413), .Z(n23303) );
  XOR2_X1 U25241 ( .A1(n7363), .A2(n25311), .Z(n23302) );
  XOR2_X1 U25242 ( .A1(n23303), .A2(n23302), .Z(n23304) );
  XOR2_X1 U25243 ( .A1(n26656), .A2(n31513), .Z(n23310) );
  XOR2_X1 U25248 ( .A1(n23328), .A2(n25878), .Z(n23329) );
  XOR2_X1 U25249 ( .A1(n16160), .A2(n24514), .Z(n23338) );
  NAND2_X1 U25250 ( .A1(n23871), .A2(n27163), .ZN(n24186) );
  NOR2_X1 U25252 ( .A1(n23726), .A2(n23348), .ZN(n23971) );
  NOR2_X1 U25253 ( .A1(n23510), .A2(n23721), .ZN(n23350) );
  NAND2_X1 U25254 ( .A1(n23351), .A2(n16337), .ZN(n23353) );
  XOR2_X1 U25256 ( .A1(n16530), .A2(n23405), .Z(n23356) );
  XOR2_X1 U25258 ( .A1(n15130), .A2(n25206), .Z(n23364) );
  XOR2_X1 U25259 ( .A1(n23371), .A2(n25191), .Z(n23372) );
  XOR2_X1 U25260 ( .A1(n23373), .A2(n23372), .Z(n23374) );
  INV_X1 U25265 ( .I(n23395), .ZN(n23396) );
  XOR2_X1 U25266 ( .A1(n33971), .A2(n23396), .Z(n23397) );
  XOR2_X1 U25267 ( .A1(n16631), .A2(n23405), .Z(n23406) );
  XOR2_X1 U25269 ( .A1(n23420), .A2(n25493), .Z(n23421) );
  XOR2_X1 U25272 ( .A1(n23429), .A2(n23430), .Z(n23432) );
  XOR2_X1 U25273 ( .A1(n33293), .A2(n24937), .Z(n23431) );
  XOR2_X1 U25274 ( .A1(n23431), .A2(n23432), .Z(n23433) );
  XOR2_X1 U25275 ( .A1(n27708), .A2(n16612), .Z(n23436) );
  XOR2_X1 U25276 ( .A1(n23467), .A2(n25560), .Z(n23468) );
  INV_X1 U25277 ( .I(n23485), .ZN(n23481) );
  INV_X1 U25278 ( .I(n23479), .ZN(n23483) );
  NOR2_X1 U25279 ( .A1(n23483), .A2(n25545), .ZN(n23480) );
  OAI21_X1 U25280 ( .A1(n23481), .A2(n23482), .B(n23480), .ZN(n23487) );
  NOR2_X1 U25281 ( .A1(n23482), .A2(n15816), .ZN(n23484) );
  AOI22_X1 U25282 ( .A1(n23485), .A2(n23484), .B1(n23483), .B2(n25545), .ZN(
        n23486) );
  XOR2_X1 U25283 ( .A1(n982), .A2(n23511), .Z(n23512) );
  XOR2_X1 U25284 ( .A1(n31554), .A2(n8487), .Z(n23513) );
  XOR2_X1 U25287 ( .A1(n10773), .A2(n24869), .Z(n23523) );
  XOR2_X1 U25288 ( .A1(n23524), .A2(n23523), .Z(n23525) );
  NAND2_X1 U25289 ( .A1(n26290), .A2(n23527), .ZN(n23528) );
  NAND2_X1 U25293 ( .A1(n23540), .A2(n13343), .ZN(n23548) );
  XOR2_X1 U25294 ( .A1(n23552), .A2(n23551), .Z(n23553) );
  XOR2_X1 U25295 ( .A1(n23554), .A2(n23553), .Z(n24359) );
  NAND2_X1 U25301 ( .A1(n16186), .A2(n23917), .ZN(n23573) );
  NOR2_X1 U25307 ( .A1(n23770), .A2(n23768), .ZN(n23598) );
  AOI21_X1 U25308 ( .A1(n23778), .A2(n11392), .B(n23775), .ZN(n23604) );
  NAND3_X1 U25309 ( .A1(n24220), .A2(n1096), .A3(n24218), .ZN(n23606) );
  NAND2_X1 U25310 ( .A1(n791), .A2(n24219), .ZN(n23605) );
  NOR2_X1 U25312 ( .A1(n24289), .A2(n24110), .ZN(n23618) );
  NAND3_X1 U25317 ( .A1(n16388), .A2(n29272), .A3(n28510), .ZN(n23636) );
  INV_X1 U25322 ( .I(n23655), .ZN(n23656) );
  NAND2_X1 U25324 ( .A1(n13308), .A2(n11621), .ZN(n23670) );
  MUX2_X1 U25325 ( .I0(n24142), .I1(n24144), .S(n319), .Z(n23680) );
  NAND2_X1 U25329 ( .A1(n13549), .A2(n1253), .ZN(n23676) );
  OAI21_X1 U25338 ( .A1(n29269), .A2(n23527), .B(n23717), .ZN(n23718) );
  NAND3_X1 U25339 ( .A1(n23765), .A2(n1101), .A3(n23352), .ZN(n23724) );
  INV_X1 U25340 ( .I(n23728), .ZN(n23731) );
  MUX2_X1 U25343 ( .I0(n23735), .I1(n29865), .S(n23736), .Z(n23740) );
  AOI21_X2 U25344 ( .A1(n23740), .A2(n28676), .B(n23739), .ZN(n24072) );
  NAND3_X1 U25347 ( .A1(n23776), .A2(n8547), .A3(n23775), .ZN(n23780) );
  XOR2_X1 U25348 ( .A1(n24638), .A2(n16705), .Z(n23790) );
  NOR2_X1 U25350 ( .A1(n14975), .A2(n16238), .ZN(n23784) );
  NAND2_X1 U25353 ( .A1(n23797), .A2(n23857), .ZN(n23799) );
  INV_X1 U25357 ( .I(n23868), .ZN(n23869) );
  NAND2_X1 U25358 ( .A1(n23870), .A2(n31179), .ZN(n23978) );
  INV_X1 U25360 ( .I(n23929), .ZN(n23922) );
  INV_X1 U25361 ( .I(n23928), .ZN(n23921) );
  INV_X1 U25364 ( .I(n23966), .ZN(n23969) );
  INV_X1 U25365 ( .I(n23967), .ZN(n23968) );
  INV_X1 U25366 ( .I(n23971), .ZN(n23972) );
  NAND3_X1 U25367 ( .A1(n23974), .A2(n23973), .A3(n23972), .ZN(n23975) );
  INV_X1 U25370 ( .I(n24183), .ZN(n23994) );
  XOR2_X1 U25374 ( .A1(n24992), .A2(n24520), .Z(n24021) );
  NOR2_X1 U25379 ( .A1(n24305), .A2(n14252), .ZN(n24032) );
  NAND2_X1 U25380 ( .A1(n24114), .A2(n24040), .ZN(n24041) );
  XOR2_X1 U25381 ( .A1(n24513), .A2(n31687), .Z(n24049) );
  XOR2_X1 U25382 ( .A1(n24049), .A2(n24048), .Z(n24050) );
  INV_X1 U25384 ( .I(n24065), .ZN(n24993) );
  MUX2_X1 U25388 ( .I0(n33540), .I1(n33680), .S(n24243), .Z(n24076) );
  NAND3_X1 U25389 ( .A1(n890), .A2(n10987), .A3(n24326), .ZN(n24081) );
  NOR2_X1 U25390 ( .A1(n890), .A2(n24128), .ZN(n24082) );
  XOR2_X1 U25392 ( .A1(n24786), .A2(n12969), .Z(n24089) );
  XOR2_X1 U25395 ( .A1(n16679), .A2(n24622), .Z(n24098) );
  NOR2_X1 U25396 ( .A1(n24878), .A2(n24974), .ZN(n24099) );
  INV_X1 U25399 ( .I(n24174), .ZN(n24607) );
  NAND4_X1 U25402 ( .A1(n24189), .A2(n24188), .A3(n24187), .A4(n24186), .ZN(
        n24190) );
  NAND2_X1 U25403 ( .A1(n9368), .A2(n32349), .ZN(n24208) );
  XOR2_X1 U25405 ( .A1(n24474), .A2(n24707), .Z(n24215) );
  NAND2_X1 U25406 ( .A1(n32737), .A2(n24225), .ZN(n24227) );
  INV_X1 U25407 ( .I(n24231), .ZN(n25259) );
  XOR2_X1 U25408 ( .A1(n4728), .A2(n16636), .Z(n24241) );
  NAND3_X1 U25411 ( .A1(n24265), .A2(n31096), .A3(n16621), .ZN(n24266) );
  XOR2_X1 U25412 ( .A1(n25450), .A2(n11332), .Z(n24267) );
  XOR2_X1 U25413 ( .A1(n24394), .A2(n31687), .Z(n24281) );
  XOR2_X1 U25414 ( .A1(n24475), .A2(n25910), .Z(n24280) );
  NAND2_X1 U25417 ( .A1(n28240), .A2(n319), .ZN(n24300) );
  NAND2_X1 U25418 ( .A1(n24300), .A2(n1241), .ZN(n24301) );
  INV_X1 U25420 ( .I(n24330), .ZN(n24333) );
  INV_X1 U25421 ( .I(n24331), .ZN(n24332) );
  XOR2_X1 U25425 ( .A1(n25436), .A2(n24592), .Z(n24355) );
  XOR2_X1 U25431 ( .A1(n24761), .A2(n30540), .Z(n24371) );
  INV_X1 U25432 ( .I(n24374), .ZN(n25567) );
  NOR2_X1 U25433 ( .A1(n25620), .A2(n25752), .ZN(n24378) );
  XOR2_X1 U25436 ( .A1(n24686), .A2(n25086), .Z(n24387) );
  XOR2_X1 U25437 ( .A1(n24814), .A2(n24391), .Z(n24392) );
  XOR2_X1 U25441 ( .A1(n25218), .A2(n11868), .Z(n24402) );
  XOR2_X1 U25443 ( .A1(n24786), .A2(n25578), .Z(n24410) );
  XOR2_X1 U25444 ( .A1(n24411), .A2(n24410), .Z(n24412) );
  XOR2_X1 U25446 ( .A1(n887), .A2(n24620), .Z(n24428) );
  XOR2_X1 U25449 ( .A1(n24962), .A2(n24753), .Z(n24444) );
  XOR2_X1 U25451 ( .A1(n24453), .A2(n24547), .Z(n24457) );
  INV_X1 U25453 ( .I(n16757), .ZN(n25564) );
  OAI21_X1 U25456 ( .A1(n18264), .A2(n8758), .B(n32012), .ZN(n24485) );
  XOR2_X1 U25458 ( .A1(n24781), .A2(n24622), .Z(n24491) );
  NAND2_X1 U25459 ( .A1(n24498), .A2(n15409), .ZN(n24501) );
  NAND2_X1 U25460 ( .A1(n24499), .A2(n15409), .ZN(n24500) );
  NAND2_X1 U25462 ( .A1(n32798), .A2(n28136), .ZN(n24506) );
  XOR2_X1 U25464 ( .A1(n24660), .A2(n24514), .Z(n24515) );
  XOR2_X1 U25465 ( .A1(n24518), .A2(n24517), .Z(n24519) );
  XOR2_X1 U25467 ( .A1(n24522), .A2(n27385), .Z(n24523) );
  OAI21_X1 U25469 ( .A1(n16650), .A2(n25397), .B(n25343), .ZN(n24557) );
  XOR2_X1 U25470 ( .A1(n24937), .A2(n24559), .Z(n24560) );
  NOR2_X1 U25475 ( .A1(n11409), .A2(n24570), .ZN(n24584) );
  INV_X1 U25476 ( .I(n24572), .ZN(n24583) );
  NAND2_X1 U25477 ( .A1(n33761), .A2(n25229), .ZN(n24580) );
  MUX2_X1 U25478 ( .I0(n24581), .I1(n24580), .S(n32864), .Z(n24582) );
  NOR2_X1 U25482 ( .A1(n24969), .A2(n24970), .ZN(n24615) );
  INV_X1 U25485 ( .I(n24623), .ZN(n25065) );
  INV_X1 U25488 ( .I(n24655), .ZN(n24657) );
  XOR2_X1 U25489 ( .A1(n24658), .A2(n24659), .Z(n24662) );
  INV_X1 U25491 ( .I(n24664), .ZN(n24665) );
  XOR2_X1 U25492 ( .A1(n31713), .A2(n24665), .Z(n24666) );
  INV_X1 U25499 ( .I(Key[10]), .ZN(n25864) );
  XOR2_X1 U25500 ( .A1(n24836), .A2(n24686), .Z(n24688) );
  INV_X1 U25502 ( .I(n16523), .ZN(n24696) );
  XOR2_X1 U25503 ( .A1(n24698), .A2(n24697), .Z(n24699) );
  NAND3_X2 U25505 ( .A1(n24704), .A2(n24703), .A3(n24702), .ZN(n25478) );
  NOR2_X1 U25506 ( .A1(n25403), .A2(n25400), .ZN(n24705) );
  INV_X1 U25507 ( .I(n25701), .ZN(n24713) );
  NOR2_X1 U25509 ( .A1(n25816), .A2(n11003), .ZN(n24721) );
  INV_X1 U25510 ( .I(n25804), .ZN(n25805) );
  NAND2_X1 U25511 ( .A1(n25805), .A2(n4450), .ZN(n24720) );
  XOR2_X1 U25514 ( .A1(n24741), .A2(n24999), .Z(n24742) );
  XOR2_X1 U25515 ( .A1(n24743), .A2(n24742), .Z(n24744) );
  XOR2_X1 U25516 ( .A1(n24745), .A2(n24744), .Z(n25022) );
  XOR2_X1 U25518 ( .A1(n30307), .A2(n25500), .Z(n24757) );
  XOR2_X1 U25521 ( .A1(n24801), .A2(n16622), .Z(n24802) );
  XOR2_X1 U25522 ( .A1(n24817), .A2(n24818), .Z(n24822) );
  XOR2_X1 U25523 ( .A1(n24819), .A2(n25288), .Z(n24820) );
  XOR2_X1 U25524 ( .A1(n12800), .A2(n24833), .Z(n24834) );
  XOR2_X1 U25526 ( .A1(n31713), .A2(n24869), .Z(n24848) );
  NAND2_X1 U25527 ( .A1(n25148), .A2(n17005), .ZN(n24856) );
  XOR2_X1 U25529 ( .A1(n24862), .A2(n24861), .Z(Ciphertext[149]) );
  INV_X1 U25531 ( .I(n25529), .ZN(n24865) );
  NAND2_X1 U25533 ( .A1(n15046), .A2(n11898), .ZN(n24876) );
  NAND2_X1 U25534 ( .A1(n15046), .A2(n24973), .ZN(n24879) );
  OR2_X1 U25536 ( .A1(n27651), .A2(n25019), .Z(n24882) );
  NAND3_X1 U25537 ( .A1(n25019), .A2(n5202), .A3(n560), .ZN(n24886) );
  NAND3_X1 U25539 ( .A1(n24884), .A2(n25114), .A3(n16025), .ZN(n24885) );
  NAND3_X1 U25542 ( .A1(n1201), .A2(n24938), .A3(n965), .ZN(n24897) );
  NOR3_X1 U25544 ( .A1(n24905), .A2(n10755), .A3(n24902), .ZN(n24899) );
  AOI21_X1 U25545 ( .A1(n24916), .A2(n24908), .B(n24899), .ZN(n24901) );
  XOR2_X1 U25546 ( .A1(n24901), .A2(n28575), .Z(Ciphertext[1]) );
  OAI22_X1 U25547 ( .A1(n24928), .A2(n24927), .B1(n24936), .B2(n24926), .ZN(
        n24929) );
  AOI21_X1 U25548 ( .A1(n24931), .A2(n24930), .B(n24929), .ZN(n24932) );
  XOR2_X1 U25549 ( .A1(n24932), .A2(n15409), .Z(Ciphertext[10]) );
  NAND2_X1 U25550 ( .A1(n24939), .A2(n24938), .ZN(n24942) );
  INV_X1 U25551 ( .I(n28662), .ZN(n24940) );
  AOI22_X1 U25552 ( .A1(n24942), .A2(n24955), .B1(n24941), .B2(n24940), .ZN(
        n24945) );
  XOR2_X1 U25553 ( .A1(n24945), .A2(n24944), .Z(Ciphertext[12]) );
  OAI21_X1 U25554 ( .A1(n24948), .A2(n24947), .B(n24946), .ZN(n24949) );
  OAI21_X1 U25557 ( .A1(n24958), .A2(n965), .B(n24954), .ZN(n24961) );
  NAND2_X1 U25558 ( .A1(n24957), .A2(n24956), .ZN(n24959) );
  XOR2_X1 U25562 ( .A1(n25000), .A2(n1415), .Z(Ciphertext[31]) );
  NOR2_X1 U25564 ( .A1(n25050), .A2(n25057), .ZN(n25029) );
  NOR2_X1 U25565 ( .A1(n25121), .A2(n8210), .ZN(n25024) );
  NAND3_X1 U25566 ( .A1(n25025), .A2(n25120), .A3(n25152), .ZN(n25028) );
  NAND2_X1 U25567 ( .A1(n25026), .A2(n16293), .ZN(n25027) );
  NOR2_X1 U25569 ( .A1(n32760), .A2(n32106), .ZN(n25031) );
  OAI21_X1 U25571 ( .A1(n25063), .A2(n25044), .B(n25057), .ZN(n25034) );
  NAND2_X1 U25572 ( .A1(n25035), .A2(n25034), .ZN(n25037) );
  XOR2_X1 U25573 ( .A1(n25037), .A2(n25036), .Z(Ciphertext[36]) );
  NAND2_X1 U25576 ( .A1(n25058), .A2(n25051), .ZN(n25042) );
  MUX2_X1 U25579 ( .I0(n25062), .I1(n31640), .S(n25057), .Z(n25053) );
  XOR2_X1 U25580 ( .A1(n25055), .A2(n25054), .Z(Ciphertext[40]) );
  NAND2_X1 U25582 ( .A1(n25078), .A2(n16809), .ZN(n25070) );
  AOI21_X1 U25585 ( .A1(n25105), .A2(n25100), .B(n32857), .ZN(n25084) );
  XOR2_X1 U25587 ( .A1(n25087), .A2(n13331), .Z(Ciphertext[48]) );
  INV_X1 U25588 ( .I(n25088), .ZN(n25090) );
  INV_X1 U25590 ( .I(n25094), .ZN(n25095) );
  INV_X1 U25591 ( .I(n25185), .ZN(n25183) );
  NAND2_X1 U25593 ( .A1(n25187), .A2(n8219), .ZN(n25132) );
  NOR2_X1 U25596 ( .A1(n14627), .A2(n15641), .ZN(n25143) );
  NAND2_X1 U25597 ( .A1(n7765), .A2(n25175), .ZN(n25155) );
  OAI22_X1 U25598 ( .A1(n25180), .A2(n25153), .B1(n25158), .B2(n25155), .ZN(
        n25157) );
  XOR2_X1 U25599 ( .A1(n25157), .A2(n25156), .Z(Ciphertext[61]) );
  INV_X1 U25600 ( .I(n25161), .ZN(n25162) );
  XOR2_X1 U25601 ( .A1(n25163), .A2(n25162), .Z(Ciphertext[62]) );
  NAND2_X1 U25602 ( .A1(n25165), .A2(n25175), .ZN(n25166) );
  NAND3_X1 U25603 ( .A1(n25170), .A2(n25169), .A3(n25168), .ZN(n25171) );
  NOR2_X1 U25607 ( .A1(n25339), .A2(n25232), .ZN(n25196) );
  XOR2_X1 U25608 ( .A1(n25219), .A2(n1414), .Z(Ciphertext[76]) );
  OAI21_X1 U25609 ( .A1(n16650), .A2(n25400), .B(n14246), .ZN(n25231) );
  NOR2_X1 U25610 ( .A1(n25253), .A2(n25237), .ZN(n25248) );
  OAI21_X1 U25611 ( .A1(n25977), .A2(n32601), .B(n9162), .ZN(n25243) );
  NAND3_X1 U25612 ( .A1(n31268), .A2(n1224), .A3(n33493), .ZN(n25245) );
  XOR2_X1 U25613 ( .A1(n25255), .A2(n16602), .Z(Ciphertext[82]) );
  AOI21_X1 U25614 ( .A1(n733), .A2(n25279), .B(n25278), .ZN(n25265) );
  NAND2_X1 U25615 ( .A1(n25284), .A2(n28532), .ZN(n25264) );
  NAND3_X1 U25616 ( .A1(n13985), .A2(n25302), .A3(n25261), .ZN(n25262) );
  XOR2_X1 U25617 ( .A1(n25267), .A2(n26000), .Z(Ciphertext[84]) );
  NAND2_X1 U25619 ( .A1(n25279), .A2(n25278), .ZN(n25268) );
  NAND2_X1 U25622 ( .A1(n16291), .A2(n25278), .ZN(n25272) );
  OAI21_X1 U25626 ( .A1(n7081), .A2(n11132), .B(n25290), .ZN(n25294) );
  NAND2_X1 U25627 ( .A1(n11132), .A2(n25339), .ZN(n25291) );
  NAND3_X1 U25628 ( .A1(n17110), .A2(n25292), .A3(n25291), .ZN(n25293) );
  NAND3_X1 U25634 ( .A1(n17110), .A2(n32659), .A3(n25339), .ZN(n25340) );
  NOR2_X1 U25636 ( .A1(n25352), .A2(n25375), .ZN(n25349) );
  INV_X1 U25637 ( .I(n25368), .ZN(n25379) );
  NOR2_X1 U25639 ( .A1(n25367), .A2(n25368), .ZN(n25354) );
  NAND2_X1 U25640 ( .A1(n25352), .A2(n25361), .ZN(n25353) );
  NAND2_X1 U25644 ( .A1(n30276), .A2(n25376), .ZN(n25365) );
  NAND3_X1 U25645 ( .A1(n30400), .A2(n30302), .A3(n25368), .ZN(n25370) );
  AOI21_X1 U25647 ( .A1(n25376), .A2(n25375), .B(n30276), .ZN(n25377) );
  NAND2_X1 U25651 ( .A1(n25331), .A2(n25562), .ZN(n25383) );
  OAI21_X1 U25656 ( .A1(n25430), .A2(n25425), .B(n25445), .ZN(n25416) );
  NAND2_X1 U25658 ( .A1(n16650), .A2(n25400), .ZN(n25401) );
  XOR2_X1 U25664 ( .A1(n25417), .A2(n1394), .Z(Ciphertext[102]) );
  NAND2_X1 U25667 ( .A1(n25425), .A2(n25429), .ZN(n25419) );
  AOI22_X1 U25671 ( .A1(n29280), .A2(n25453), .B1(n25424), .B2(n25437), .ZN(
        n25427) );
  NAND2_X1 U25674 ( .A1(n29280), .A2(n25437), .ZN(n25449) );
  NAND3_X1 U25677 ( .A1(n25452), .A2(n25446), .A3(n25455), .ZN(n25447) );
  NOR2_X1 U25681 ( .A1(n25462), .A2(n6310), .ZN(n25459) );
  XOR2_X1 U25684 ( .A1(n25467), .A2(n1404), .Z(n25468) );
  NAND3_X1 U25685 ( .A1(n25468), .A2(n25470), .A3(n25475), .ZN(n25485) );
  INV_X1 U25686 ( .I(n25482), .ZN(n25472) );
  NAND3_X1 U25692 ( .A1(n25477), .A2(n4183), .A3(n25476), .ZN(n25481) );
  NAND3_X1 U25693 ( .A1(n25479), .A2(n1404), .A3(n6310), .ZN(n25480) );
  XOR2_X1 U25695 ( .A1(n25494), .A2(n1065), .Z(Ciphertext[113]) );
  OAI21_X1 U25696 ( .A1(n2480), .A2(n32897), .B(n8766), .ZN(n25499) );
  INV_X1 U25697 ( .I(n32897), .ZN(n25495) );
  OAI21_X1 U25698 ( .A1(n25499), .A2(n25498), .B(n25497), .ZN(n25501) );
  XOR2_X1 U25699 ( .A1(n25501), .A2(n25500), .Z(Ciphertext[114]) );
  NAND2_X1 U25701 ( .A1(n749), .A2(n32897), .ZN(n25514) );
  NAND2_X1 U25702 ( .A1(n25561), .A2(n16783), .ZN(n25522) );
  NAND2_X1 U25706 ( .A1(n25550), .A2(n15134), .ZN(n25543) );
  NAND3_X1 U25707 ( .A1(n25550), .A2(n31647), .A3(n8320), .ZN(n25547) );
  NAND2_X1 U25709 ( .A1(n25707), .A2(n11944), .ZN(n25579) );
  NAND3_X1 U25711 ( .A1(n25593), .A2(n12042), .A3(n837), .ZN(n25594) );
  NAND2_X1 U25719 ( .A1(n11931), .A2(n25615), .ZN(n25608) );
  XOR2_X1 U25723 ( .A1(n25642), .A2(n16472), .Z(Ciphertext[139]) );
  AOI21_X1 U25731 ( .A1(n34094), .A2(n3883), .B(n26322), .ZN(n25667) );
  NAND3_X1 U25732 ( .A1(n25691), .A2(n25687), .A3(n32879), .ZN(n25672) );
  AOI21_X1 U25735 ( .A1(n17120), .A2(n33976), .B(n25760), .ZN(n25676) );
  NAND3_X1 U25736 ( .A1(n25680), .A2(n26447), .A3(n25679), .ZN(n25683) );
  NAND3_X1 U25738 ( .A1(n33386), .A2(n10376), .A3(n25731), .ZN(n25718) );
  NAND2_X1 U25739 ( .A1(n25719), .A2(n25718), .ZN(n25721) );
  XOR2_X1 U25740 ( .A1(n25721), .A2(n25720), .Z(Ciphertext[152]) );
  NAND3_X1 U25742 ( .A1(n25731), .A2(n16494), .A3(n25729), .ZN(n25726) );
  OAI21_X1 U25744 ( .A1(n13640), .A2(n16494), .B(n25729), .ZN(n25730) );
  NAND2_X1 U25745 ( .A1(n25746), .A2(n32863), .ZN(n25737) );
  OAI21_X1 U25746 ( .A1(n25743), .A2(n27164), .B(n25738), .ZN(n25741) );
  INV_X1 U25747 ( .I(n25743), .ZN(n25749) );
  NAND3_X1 U25749 ( .A1(n25788), .A2(n25781), .A3(n12611), .ZN(n25770) );
  NAND2_X1 U25750 ( .A1(n25763), .A2(n146), .ZN(n25764) );
  NOR2_X1 U25751 ( .A1(n32874), .A2(n25795), .ZN(n25798) );
  AOI21_X1 U25752 ( .A1(n25775), .A2(n12611), .B(n25774), .ZN(n25776) );
  OAI21_X1 U25753 ( .A1(n25798), .A2(n25777), .B(n25776), .ZN(n25778) );
  XOR2_X1 U25754 ( .A1(n25778), .A2(n17063), .Z(Ciphertext[164]) );
  INV_X1 U25755 ( .I(n25780), .ZN(n25782) );
  INV_X1 U25756 ( .I(n25784), .ZN(n25785) );
  OAI21_X1 U25757 ( .A1(n11899), .A2(n25786), .B(n25785), .ZN(n25787) );
  NAND2_X1 U25758 ( .A1(n25789), .A2(n25788), .ZN(n25792) );
  XOR2_X1 U25763 ( .A1(n25802), .A2(n25801), .Z(Ciphertext[167]) );
  NOR2_X1 U25764 ( .A1(n4450), .A2(n25804), .ZN(n25803) );
  OAI21_X1 U25765 ( .A1(n25823), .A2(n25805), .B(n11003), .ZN(n25808) );
  XOR2_X1 U25766 ( .A1(n25810), .A2(n32981), .Z(Ciphertext[170]) );
  NAND2_X1 U25767 ( .A1(n25817), .A2(n25816), .ZN(n25821) );
  AOI21_X1 U25768 ( .A1(n25823), .A2(n25804), .B(n25822), .ZN(n25824) );
  OAI22_X1 U25769 ( .A1(n25826), .A2(n25825), .B1(n9181), .B2(n25824), .ZN(
        n25828) );
  XOR2_X1 U25770 ( .A1(n25828), .A2(n25827), .Z(Ciphertext[173]) );
  OAI21_X1 U25771 ( .A1(n25834), .A2(n25851), .B(n14199), .ZN(n25830) );
  NOR3_X1 U25772 ( .A1(n16673), .A2(n10897), .A3(n25851), .ZN(n25829) );
  XOR2_X1 U25774 ( .A1(n25833), .A2(n1064), .Z(Ciphertext[174]) );
  NOR2_X1 U25775 ( .A1(n25851), .A2(n13049), .ZN(n25835) );
  OAI22_X1 U25776 ( .A1(n25836), .A2(n25852), .B1(n25835), .B2(n25853), .ZN(
        n25837) );
  XOR2_X1 U25777 ( .A1(n25837), .A2(n16654), .Z(Ciphertext[175]) );
  NOR2_X1 U25779 ( .A1(n25838), .A2(n25901), .ZN(n25841) );
  NOR4_X1 U25780 ( .A1(n25843), .A2(n31979), .A3(n25841), .A4(n25840), .ZN(
        n25847) );
  INV_X1 U25784 ( .I(n25923), .ZN(n25906) );
  MUX2_X1 U25785 ( .I0(n25922), .I1(n25925), .S(n25915), .Z(n25909) );
  AOI21_X1 U25787 ( .A1(n25923), .A2(n14359), .B(n25922), .ZN(n25924) );
  INV_X2 U6220 ( .I(n23944), .ZN(n1256) );
  INV_X2 U322 ( .I(n23275), .ZN(n721) );
  INV_X4 U5017 ( .I(n10302), .ZN(n6003) );
  INV_X4 U20459 ( .I(n25232), .ZN(n11132) );
  INV_X2 U923 ( .I(n19300), .ZN(n730) );
  BUF_X2 U1607 ( .I(n22390), .Z(n15260) );
  INV_X4 U6339 ( .I(n17394), .ZN(n992) );
  INV_X4 U7806 ( .I(n28202), .ZN(n24335) );
  NAND2_X2 U944 ( .A1(n5119), .A2(n5118), .ZN(n19103) );
  NAND2_X2 U5101 ( .A1(n27619), .A2(n26445), .ZN(n21550) );
  NAND2_X2 U668 ( .A1(n21095), .A2(n9322), .ZN(n12811) );
  NAND2_X2 U1745 ( .A1(n725), .A2(n14540), .ZN(n7746) );
  NAND2_X2 U2920 ( .A1(n24120), .A2(n1775), .ZN(n23791) );
  INV_X2 U799 ( .I(n20228), .ZN(n20325) );
  NOR2_X2 U6586 ( .A1(n19269), .A2(n19265), .ZN(n19226) );
  INV_X4 U203 ( .I(n23540), .ZN(n24114) );
  AOI21_X2 U5929 ( .A1(n17239), .A2(n18922), .B(n17238), .ZN(n15991) );
  INV_X2 U10570 ( .I(n24198), .ZN(n16712) );
  INV_X4 U287 ( .I(n13297), .ZN(n23828) );
  BUF_X2 U4738 ( .I(n24360), .Z(n25884) );
  OAI21_X2 U4497 ( .A1(n2633), .A2(n2634), .B(n23137), .ZN(n2631) );
  AOI22_X2 U8397 ( .A1(n20506), .A2(n14367), .B1(n10057), .B2(n20435), .ZN(
        n6775) );
  INV_X2 U107 ( .I(n18156), .ZN(n18154) );
  INV_X2 U4429 ( .I(n17535), .ZN(n25711) );
  INV_X2 U4446 ( .I(n25962), .ZN(n15770) );
  AOI22_X2 U4784 ( .A1(n9813), .A2(n801), .B1(n9812), .B2(n27163), .ZN(n5258)
         );
  NAND2_X2 U990 ( .A1(n12327), .A2(n7164), .ZN(n18577) );
  AOI21_X2 U751 ( .A1(n11809), .A2(n125), .B(n11808), .ZN(n12147) );
  NAND2_X2 U1673 ( .A1(n24925), .A2(n24927), .ZN(n24922) );
  INV_X2 U5851 ( .I(n15733), .ZN(n21379) );
  OAI22_X2 U553 ( .A1(n11981), .A2(n21876), .B1(n13345), .B2(n8602), .ZN(
        n21702) );
  INV_X2 U208 ( .I(n24234), .ZN(n24130) );
  INV_X2 U5996 ( .I(n33094), .ZN(n18006) );
  NOR2_X2 U7575 ( .A1(n18005), .A2(n18470), .ZN(n17253) );
  NAND2_X2 U793 ( .A1(n15310), .A2(n15311), .ZN(n20463) );
  INV_X2 U23623 ( .I(n16401), .ZN(n17405) );
  OAI21_X2 U803 ( .A1(n937), .A2(n28876), .B(n27343), .ZN(n19931) );
  NAND2_X2 U4485 ( .A1(n8614), .A2(n23852), .ZN(n12722) );
  INV_X2 U859 ( .I(n12517), .ZN(n16298) );
  INV_X2 U983 ( .I(n18588), .ZN(n17687) );
  INV_X2 U304 ( .I(n9199), .ZN(n13773) );
  INV_X2 U1001 ( .I(n17030), .ZN(n12956) );
  AOI22_X2 U9851 ( .A1(n29423), .A2(n17495), .B1(n20052), .B2(n1358), .ZN(
        n3827) );
  BUF_X2 U8103 ( .I(n9170), .Z(n1842) );
  NAND2_X2 U5052 ( .A1(n22997), .A2(n22996), .ZN(n23489) );
  INV_X2 U12247 ( .I(n6215), .ZN(n9549) );
  BUF_X4 U922 ( .I(n14233), .Z(n29) );
  AOI21_X2 U8115 ( .A1(n15315), .A2(n32076), .B(n14822), .ZN(n15314) );
  NOR2_X2 U6685 ( .A1(n18798), .A2(n18797), .ZN(n18896) );
  NAND2_X2 U363 ( .A1(n31937), .A2(n4084), .ZN(n23067) );
  INV_X2 U118 ( .I(n3339), .ZN(n16589) );
  NAND2_X2 U7276 ( .A1(n1355), .A2(n15282), .ZN(n20506) );
  NOR2_X2 U206 ( .A1(n15179), .A2(n24254), .ZN(n17801) );
  INV_X2 U9205 ( .I(n14726), .ZN(n23843) );
  NOR2_X2 U8727 ( .A1(n9631), .A2(n8309), .ZN(n10784) );
  OAI21_X2 U9747 ( .A1(n5589), .A2(n5592), .B(n27785), .ZN(n5588) );
  NAND2_X2 U1566 ( .A1(n2141), .A2(n24243), .ZN(n24127) );
  NAND2_X2 U4948 ( .A1(n15051), .A2(n1573), .ZN(n2270) );
  OAI21_X2 U5772 ( .A1(n15464), .A2(n3567), .B(n10282), .ZN(n10386) );
  NOR2_X2 U529 ( .A1(n7641), .A2(n14541), .ZN(n22047) );
  NOR2_X2 U4575 ( .A1(n16512), .A2(n31874), .ZN(n20880) );
  AOI21_X2 U1907 ( .A1(n32064), .A2(n17162), .B(n12549), .ZN(n1871) );
  OAI21_X2 U399 ( .A1(n11614), .A2(n17630), .B(n22472), .ZN(n23079) );
  NAND2_X2 U9838 ( .A1(n13986), .A2(n8549), .ZN(n20294) );
  INV_X4 U6679 ( .I(n5327), .ZN(n951) );
  BUF_X2 U8704 ( .I(n10423), .Z(n4017) );
  INV_X2 U3581 ( .I(n10414), .ZN(n16789) );
  NAND2_X2 U4253 ( .A1(n4645), .A2(n4644), .ZN(n5625) );
  INV_X2 U959 ( .I(n10228), .ZN(n10229) );
  INV_X2 U569 ( .I(n21767), .ZN(n914) );
  INV_X2 U403 ( .I(n7881), .ZN(n1275) );
  NOR2_X2 U17706 ( .A1(n828), .A2(n28987), .ZN(n11815) );
  INV_X2 U4535 ( .I(n10258), .ZN(n16529) );
  NAND2_X2 U1007 ( .A1(n829), .A2(n1188), .ZN(n8788) );
  INV_X4 U209 ( .I(n9964), .ZN(n16688) );
  INV_X2 U839 ( .I(n9724), .ZN(n9748) );
  INV_X2 U103 ( .I(n17523), .ZN(n25699) );
  BUF_X2 U6466 ( .I(n21375), .Z(n16421) );
  NAND2_X2 U747 ( .A1(n1351), .A2(n9025), .ZN(n20406) );
  AOI21_X2 U9357 ( .A1(n22431), .A2(n22626), .B(n17123), .ZN(n17122) );
  INV_X2 U666 ( .I(n11847), .ZN(n12654) );
  OAI21_X2 U11620 ( .A1(n12582), .A2(n12407), .B(n10000), .ZN(n14966) );
  BUF_X2 U8844 ( .I(Key[147]), .Z(n25815) );
  NOR2_X2 U13130 ( .A1(n8212), .A2(n17370), .ZN(n12892) );
  NAND2_X2 U5370 ( .A1(n12338), .A2(n901), .ZN(n22523) );
  INV_X2 U1003 ( .I(n16849), .ZN(n4259) );
  INV_X2 U4576 ( .I(n21389), .ZN(n21147) );
  INV_X1 U2783 ( .I(n21224), .ZN(n8115) );
  INV_X2 U5523 ( .I(n18643), .ZN(n4626) );
  OAI21_X2 U5390 ( .A1(n9312), .A2(n9313), .B(n17385), .ZN(n2490) );
  INV_X2 U565 ( .I(n21122), .ZN(n913) );
  INV_X1 U117 ( .I(n12358), .ZN(n716) );
  OAI21_X2 U241 ( .A1(n144), .A2(n10068), .B(n23940), .ZN(n2448) );
  NAND2_X2 U3422 ( .A1(n14280), .A2(n13379), .ZN(n7228) );
  INV_X4 U4804 ( .I(n23806), .ZN(n1100) );
  INV_X2 U493 ( .I(n31932), .ZN(n11917) );
  INV_X2 U232 ( .I(n5317), .ZN(n5318) );
  NAND2_X2 U22011 ( .A1(n3891), .A2(n12586), .ZN(n22834) );
  OAI21_X2 U6492 ( .A1(n16174), .A2(n20515), .B(n20517), .ZN(n10731) );
  INV_X2 U1170 ( .I(n7746), .ZN(n17149) );
  INV_X4 U865 ( .I(n16317), .ZN(n15665) );
  AOI21_X2 U9771 ( .A1(n12089), .A2(n20333), .B(n12880), .ZN(n12879) );
  OAI21_X2 U730 ( .A1(n29444), .A2(n16070), .B(n1157), .ZN(n4772) );
  AOI22_X2 U8662 ( .A1(n13806), .A2(n26350), .B1(n10700), .B2(n14312), .ZN(
        n3920) );
  INV_X2 U5401 ( .I(n29523), .ZN(n21859) );
  NAND2_X2 U7302 ( .A1(n33091), .A2(n20158), .ZN(n20333) );
  INV_X2 U704 ( .I(n6684), .ZN(n21085) );
  NAND2_X2 U13709 ( .A1(n11947), .A2(n9436), .ZN(n25205) );
  OAI21_X2 U7053 ( .A1(n8274), .A2(n21607), .B(n21775), .ZN(n21609) );
  AOI21_X2 U353 ( .A1(n1274), .A2(n2580), .B(n2579), .ZN(n4543) );
  OR2_X2 U5609 ( .A1(n17499), .A2(n24447), .Z(n17092) );
  NAND2_X2 U8434 ( .A1(n1153), .A2(n28028), .ZN(n14177) );
  NOR2_X2 U236 ( .A1(n23170), .A2(n23169), .ZN(n24060) );
  INV_X4 U6618 ( .I(n2080), .ZN(n19315) );
  INV_X2 U5657 ( .I(n11041), .ZN(n23714) );
  INV_X2 U211 ( .I(n18077), .ZN(n17310) );
  INV_X2 U4543 ( .I(n22363), .ZN(n22588) );
  OAI21_X2 U1658 ( .A1(n23758), .A2(n23757), .B(n28671), .ZN(n11418) );
  INV_X2 U4352 ( .I(n27134), .ZN(n1208) );
  INV_X2 U491 ( .I(n17140), .ZN(n22428) );
  OAI21_X2 U9729 ( .A1(n12010), .A2(n20321), .B(n18078), .ZN(n13851) );
  INV_X4 U5805 ( .I(n32082), .ZN(n22576) );
  INV_X2 U3614 ( .I(n24002), .ZN(n767) );
  NAND2_X2 U10547 ( .A1(n6632), .A2(n6633), .ZN(n3380) );
  NOR2_X2 U6149 ( .A1(n3222), .A2(n24248), .ZN(n14972) );
  INV_X2 U698 ( .I(n13921), .ZN(n12747) );
  INV_X2 U4989 ( .I(n9163), .ZN(n12039) );
  NAND2_X2 U46 ( .A1(n9754), .A2(n1462), .ZN(n25513) );
  AOI21_X2 U7949 ( .A1(n23085), .A2(n22884), .B(n17668), .ZN(n8455) );
  INV_X4 U8469 ( .I(n32240), .ZN(n1153) );
  NAND2_X2 U342 ( .A1(n8226), .A2(n11467), .ZN(n12181) );
  INV_X2 U5184 ( .I(n18139), .ZN(n8376) );
  OAI21_X2 U6593 ( .A1(n15050), .A2(n19248), .B(n4591), .ZN(n14757) );
  INV_X4 U6564 ( .I(n4577), .ZN(n17670) );
  INV_X1 U1623 ( .I(n8558), .ZN(n1617) );
  BUF_X2 U7660 ( .I(Key[113]), .Z(n25064) );
  INV_X1 U11202 ( .I(n22656), .ZN(n1286) );
  INV_X4 U4508 ( .I(n1485), .ZN(n22977) );
  INV_X2 U5083 ( .I(n632), .ZN(n15752) );
  BUF_X4 U4627 ( .I(n5545), .Z(n1053) );
  BUF_X4 U8705 ( .I(n19222), .Z(n16185) );
  NAND2_X2 U4849 ( .A1(n18210), .A2(n18209), .ZN(n21646) );
  NAND2_X2 U11253 ( .A1(n21276), .A2(n21277), .ZN(n15385) );
  NAND2_X2 U6485 ( .A1(n14731), .A2(n11086), .ZN(n19826) );
  INV_X2 U545 ( .I(n21821), .ZN(n1317) );
  OAI21_X2 U10111 ( .A1(n18772), .A2(n5805), .B(n18771), .ZN(n5311) );
  OAI22_X2 U5426 ( .A1(n20475), .A2(n33288), .B1(n7394), .B2(n12758), .ZN(
        n12757) );
  NAND2_X2 U9992 ( .A1(n19085), .A2(n1046), .ZN(n18405) );
  INV_X1 U8181 ( .I(n8602), .ZN(n8569) );
  NAND2_X2 U571 ( .A1(n27532), .A2(n11401), .ZN(n21643) );
  OAI22_X2 U5264 ( .A1(n12054), .A2(n29866), .B1(n24153), .B2(n26314), .ZN(
        n3918) );
  NOR2_X2 U6665 ( .A1(n6295), .A2(n328), .ZN(n9090) );
  INV_X4 U3434 ( .I(n17306), .ZN(n834) );
  INV_X1 U1283 ( .I(n13020), .ZN(n9346) );
  AOI21_X2 U5923 ( .A1(n3391), .A2(n19603), .B(n19195), .ZN(n19780) );
  NAND2_X2 U6584 ( .A1(n3390), .A2(n3389), .ZN(n19603) );
  AOI21_X2 U9483 ( .A1(n13188), .A2(n33322), .B(n13187), .ZN(n21725) );
  INV_X2 U7493 ( .I(n14624), .ZN(n9423) );
  INV_X2 U5153 ( .I(n4632), .ZN(n10831) );
  INV_X2 U2517 ( .I(n11966), .ZN(n812) );
  NOR2_X2 U8755 ( .A1(n18445), .A2(n18444), .ZN(n2099) );
  OAI21_X2 U7567 ( .A1(n18798), .A2(n7899), .B(n17843), .ZN(n18445) );
  INV_X2 U7179 ( .I(n11601), .ZN(n12363) );
  OAI21_X2 U15105 ( .A1(n12367), .A2(n12366), .B(n1023), .ZN(n12365) );
  NAND2_X2 U5931 ( .A1(n13011), .A2(n13012), .ZN(n13481) );
  NOR2_X2 U1714 ( .A1(n6219), .A2(n21359), .ZN(n10313) );
  INV_X4 U7265 ( .I(n31522), .ZN(n1026) );
  INV_X2 U769 ( .I(n20445), .ZN(n20381) );
  NAND2_X2 U4236 ( .A1(n4361), .A2(n4360), .ZN(n4362) );
  BUF_X2 U10216 ( .I(Key[182]), .Z(n25735) );
  OAI21_X2 U961 ( .A1(n18766), .A2(n14284), .B(n18765), .ZN(n18769) );
  NAND2_X2 U4639 ( .A1(n1183), .A2(n7216), .ZN(n12327) );
  NAND2_X2 U9749 ( .A1(n1026), .A2(n20257), .ZN(n3556) );
  BUF_X4 U6621 ( .I(n16960), .Z(n8862) );
  OR2_X2 U7609 ( .A1(n17558), .A2(n16450), .Z(n12989) );
  INV_X2 U947 ( .I(n16960), .ZN(n19116) );
  INV_X2 U5128 ( .I(n20526), .ZN(n868) );
  INV_X2 U6414 ( .I(n21581), .ZN(n16127) );
  INV_X4 U22830 ( .I(n14339), .ZN(n18073) );
  AOI21_X2 U12115 ( .A1(n17422), .A2(n28707), .B(n3018), .ZN(n10909) );
  BUF_X4 U5062 ( .I(n13679), .Z(n803) );
  OAI21_X2 U6622 ( .A1(n12065), .A2(n18759), .B(n15281), .ZN(n19094) );
  INV_X2 U5733 ( .I(n23267), .ZN(n14077) );
  INV_X2 U5461 ( .I(n19418), .ZN(n20059) );
  INV_X2 U9266 ( .I(n985), .ZN(n7047) );
  INV_X2 U5079 ( .I(n1299), .ZN(n22388) );
  OAI21_X2 U4614 ( .A1(n26081), .A2(n26518), .B(n8211), .ZN(n18668) );
  AOI21_X2 U9046 ( .A1(n12353), .A2(n24152), .B(n3903), .ZN(n3902) );
  NAND3_X2 U5820 ( .A1(n17983), .A2(n17982), .A3(n1652), .ZN(n14642) );
  INV_X2 U4744 ( .I(n9164), .ZN(n17824) );
  INV_X4 U11568 ( .I(n17971), .ZN(n4518) );
  NAND2_X2 U1700 ( .A1(n14244), .A2(n14247), .ZN(n14243) );
  INV_X2 U388 ( .I(n6874), .ZN(n9954) );
  INV_X2 U465 ( .I(n17518), .ZN(n22690) );
  AOI22_X2 U4898 ( .A1(n18877), .A2(n961), .B1(n14658), .B2(n18101), .ZN(
        n18939) );
  INV_X2 U225 ( .I(n31155), .ZN(n24225) );
  INV_X2 U3574 ( .I(n10284), .ZN(n18871) );
  NAND2_X2 U4076 ( .A1(n16982), .A2(n23117), .ZN(n24763) );
  INV_X2 U9945 ( .I(n17662), .ZN(n20142) );
  NOR2_X2 U5173 ( .A1(n13202), .A2(n13201), .ZN(n13673) );
  INV_X2 U6083 ( .I(n25118), .ZN(n25116) );
  NAND2_X1 U1823 ( .A1(n14344), .A2(n15406), .ZN(n10) );
  INV_X2 U4442 ( .I(n11622), .ZN(n11947) );
  INV_X2 U4243 ( .I(n9553), .ZN(n15050) );
  AOI21_X2 U6231 ( .A1(n4155), .A2(n27612), .B(n6099), .ZN(n5593) );
  OR2_X2 U4058 ( .A1(n9120), .A2(n23668), .Z(n15550) );
  INV_X2 U7234 ( .I(n32648), .ZN(n2789) );
  NAND2_X2 U6979 ( .A1(n5453), .A2(n5744), .ZN(n5448) );
  NAND2_X2 U896 ( .A1(n379), .A2(n9787), .ZN(n7438) );
  NAND2_X2 U953 ( .A1(n2684), .A2(n2683), .ZN(n19020) );
  BUF_X2 U4651 ( .I(Key[0]), .Z(n25206) );
  INV_X2 U511 ( .I(n22047), .ZN(n21996) );
  INV_X4 U5943 ( .I(n10700), .ZN(n947) );
  INV_X2 U10213 ( .I(n10664), .ZN(n10665) );
  AOI22_X2 U6681 ( .A1(n12238), .A2(n6891), .B1(n18553), .B2(n18891), .ZN(
        n14844) );
  NAND4_X1 U1491 ( .A1(n24497), .A2(n16502), .A3(n24495), .A4(n24496), .ZN(
        n24502) );
  INV_X4 U3620 ( .I(n676), .ZN(n11306) );
  NOR2_X2 U5791 ( .A1(n22537), .A2(n22428), .ZN(n22407) );
  AOI21_X2 U8401 ( .A1(n12139), .A2(n33154), .B(n20455), .ZN(n20458) );
  NOR2_X2 U9303 ( .A1(n772), .A2(n25994), .ZN(n22760) );
  CLKBUF_X4 U4905 ( .I(n12282), .Z(n6783) );
  INV_X2 U3905 ( .I(n24117), .ZN(n24223) );
  NAND2_X2 U24874 ( .A1(n13921), .A2(n27193), .ZN(n21336) );
  INV_X2 U4382 ( .I(n2536), .ZN(n7273) );
  OAI21_X2 U6540 ( .A1(n822), .A2(n3626), .B(n13346), .ZN(n20006) );
  BUF_X2 U5792 ( .I(n22589), .Z(n16562) );
  NAND3_X2 U7365 ( .A1(n6644), .A2(n14172), .A3(n20066), .ZN(n6643) );
  NAND2_X1 U14244 ( .A1(n22572), .A2(n1298), .ZN(n14775) );
  OAI21_X2 U7270 ( .A1(n8353), .A2(n16182), .B(n7056), .ZN(n7055) );
  NAND2_X2 U5858 ( .A1(n4648), .A2(n4266), .ZN(n20423) );
  AOI21_X2 U18858 ( .A1(n16221), .A2(n28404), .B(n8303), .ZN(n16106) );
  INV_X2 U4478 ( .I(n5306), .ZN(n9625) );
  INV_X2 U5035 ( .I(n23576), .ZN(n14207) );
  INV_X2 U843 ( .I(n12182), .ZN(n822) );
  NAND2_X2 U897 ( .A1(n28386), .A2(n13390), .ZN(n19281) );
  NAND2_X2 U607 ( .A1(n14397), .A2(n7182), .ZN(n21846) );
  NOR2_X2 U3598 ( .A1(n7310), .A2(n3909), .ZN(n8084) );
  BUF_X2 U6724 ( .I(Key[70]), .Z(n16697) );
  OR2_X1 U4023 ( .A1(n893), .A2(n23834), .Z(n12020) );
  INV_X2 U4189 ( .I(n7119), .ZN(n21322) );
  INV_X1 U2340 ( .I(n22307), .ZN(n16700) );
  AOI21_X2 U6419 ( .A1(n1142), .A2(n5049), .B(n5047), .ZN(n9396) );
  AOI21_X2 U6573 ( .A1(n16336), .A2(n16335), .B(n15239), .ZN(n18937) );
  BUF_X4 U795 ( .I(n20305), .Z(n15434) );
  INV_X2 U1733 ( .I(n19788), .ZN(n20009) );
  NOR2_X2 U6581 ( .A1(n19004), .A2(n7176), .ZN(n7283) );
  INV_X1 U18831 ( .I(n8277), .ZN(n23717) );
  INV_X4 U855 ( .I(n20009), .ZN(n9876) );
  NAND3_X2 U4185 ( .A1(n7667), .A2(n21429), .A3(n7430), .ZN(n21614) );
  NAND2_X2 U1629 ( .A1(n13872), .A2(n16327), .ZN(n12626) );
  NAND2_X2 U6139 ( .A1(n24154), .A2(n16799), .ZN(n17112) );
  NOR2_X2 U5261 ( .A1(n5632), .A2(n7778), .ZN(n10104) );
  BUF_X4 U5428 ( .I(n14980), .Z(n13300) );
  AOI21_X2 U25416 ( .A1(n33444), .A2(n15520), .B(n24010), .ZN(n24296) );
  INV_X4 U6650 ( .I(n19330), .ZN(n880) );
  INV_X2 U4126 ( .I(n3773), .ZN(n17161) );
  INV_X2 U659 ( .I(n9663), .ZN(n21441) );
  AOI21_X2 U7952 ( .A1(n15915), .A2(n899), .B(n22769), .ZN(n15914) );
  NOR2_X2 U24701 ( .A1(n420), .A2(n29069), .ZN(n20403) );
  INV_X2 U111 ( .I(n6143), .ZN(n25409) );
  AOI22_X2 U4696 ( .A1(n25328), .A2(n25406), .B1(n25329), .B2(n25410), .ZN(
        n6411) );
  NAND2_X1 U18918 ( .A1(n13917), .A2(n10293), .ZN(n13916) );
  INV_X2 U5190 ( .I(n18498), .ZN(n18601) );
  INV_X1 U4988 ( .I(n25628), .ZN(n755) );
  INV_X2 U6706 ( .I(n18293), .ZN(n18605) );
  BUF_X2 U4193 ( .I(n26448), .Z(n8757) );
  NOR2_X1 U10790 ( .A1(n13068), .A2(n10993), .ZN(n23539) );
  NAND2_X1 U14983 ( .A1(n21261), .A2(n21054), .ZN(n10656) );
  INV_X4 U9585 ( .I(n9076), .ZN(n21730) );
  INV_X2 U6568 ( .I(n19375), .ZN(n12998) );
  NAND2_X1 U24604 ( .A1(n8558), .A2(n15593), .ZN(n19896) );
  INV_X1 U3797 ( .I(n3933), .ZN(n21143) );
  INV_X4 U7139 ( .I(n17416), .ZN(n21812) );
  OAI21_X2 U17871 ( .A1(n8735), .A2(n829), .B(n8737), .ZN(n8734) );
  INV_X2 U6412 ( .I(n16327), .ZN(n920) );
  NAND2_X2 U6313 ( .A1(n12613), .A2(n7964), .ZN(n11161) );
  INV_X2 U4844 ( .I(n16222), .ZN(n15838) );
  INV_X2 U466 ( .I(n5975), .ZN(n8409) );
  OAI21_X2 U18231 ( .A1(n16185), .A2(n28147), .B(n4), .ZN(n7436) );
  AOI22_X2 U5217 ( .A1(n31974), .A2(n25633), .B1(n25582), .B2(n25632), .ZN(
        n15599) );
  INV_X2 U946 ( .I(n19360), .ZN(n19109) );
  INV_X1 U20868 ( .I(n21353), .ZN(n21172) );
  AND2_X2 U13467 ( .A1(n13272), .A2(n11720), .Z(n12337) );
  NAND3_X2 U5054 ( .A1(n22937), .A2(n27694), .A3(n30925), .ZN(n22852) );
  BUF_X4 U1155 ( .I(n9159), .Z(n7144) );
  AOI22_X2 U9785 ( .A1(n5029), .A2(n16182), .B1(n32035), .B2(n20603), .ZN(
        n5027) );
  INV_X4 U14381 ( .I(n3483), .ZN(n5741) );
  INV_X1 U3036 ( .I(n24561), .ZN(n304) );
  INV_X4 U4847 ( .I(n16278), .ZN(n5546) );
  INV_X4 U9323 ( .I(n22785), .ZN(n7310) );
  NAND2_X1 U11601 ( .A1(n14266), .A2(n20531), .ZN(n14262) );
  NAND2_X2 U828 ( .A1(n10831), .A2(n563), .ZN(n19855) );
  INV_X4 U9690 ( .I(n11915), .ZN(n7830) );
  NAND3_X2 U24170 ( .A1(n34140), .A2(n28757), .A3(n18642), .ZN(n18278) );
  OAI21_X2 U6251 ( .A1(n5972), .A2(n5252), .B(n17161), .ZN(n5971) );
  NAND2_X2 U4178 ( .A1(n2569), .A2(n2568), .ZN(n9999) );
  INV_X2 U5125 ( .I(n14720), .ZN(n14719) );
  NOR2_X2 U4388 ( .A1(n25639), .A2(n25638), .ZN(n25640) );
  INV_X2 U6219 ( .I(n3874), .ZN(n846) );
  NAND2_X2 U6386 ( .A1(n1137), .A2(n21816), .ZN(n21820) );
  INV_X2 U4850 ( .I(n21225), .ZN(n15261) );
  NOR2_X2 U6431 ( .A1(n164), .A2(n7430), .ZN(n21120) );
  AOI21_X2 U5358 ( .A1(n22605), .A2(n22604), .B(n22603), .ZN(n14045) );
  AOI22_X2 U8626 ( .A1(n13377), .A2(n28386), .B1(n19359), .B2(n19229), .ZN(
        n13940) );
  AOI21_X2 U22241 ( .A1(n6511), .A2(n28935), .B(n18912), .ZN(n18914) );
  INV_X4 U5464 ( .I(n10059), .ZN(n11959) );
  NAND2_X2 U6187 ( .A1(n23756), .A2(n26115), .ZN(n7885) );
  BUF_X2 U4197 ( .I(n21136), .Z(n16034) );
  NAND2_X2 U9907 ( .A1(n7804), .A2(n19450), .ZN(n3309) );
  INV_X4 U5675 ( .I(n12841), .ZN(n24052) );
  NAND2_X2 U775 ( .A1(n20213), .A2(n14564), .ZN(n20631) );
  BUF_X2 U5480 ( .I(n9319), .Z(n4714) );
  NAND2_X2 U16652 ( .A1(n26600), .A2(n16093), .ZN(n19302) );
  AOI22_X2 U7470 ( .A1(n12052), .A2(n26181), .B1(n19007), .B2(n19052), .ZN(
        n19008) );
  INV_X2 U7230 ( .I(n26448), .ZN(n1022) );
  INV_X4 U7889 ( .I(n667), .ZN(n23901) );
  INV_X1 U3525 ( .I(n3994), .ZN(n24924) );
  OAI21_X2 U13316 ( .A1(n2479), .A2(n28853), .B(n805), .ZN(n2404) );
  NOR2_X2 U1354 ( .A1(n2734), .A2(n2732), .ZN(n2731) );
  NAND2_X2 U5981 ( .A1(n13548), .A2(n13514), .ZN(n15018) );
  OR2_X2 U4254 ( .A1(n18585), .A2(n12191), .Z(n11970) );
  INV_X2 U3626 ( .I(n27154), .ZN(n6263) );
  NAND2_X2 U47 ( .A1(n25151), .A2(n34057), .ZN(n25172) );
  NOR2_X2 U21608 ( .A1(n28836), .A2(n34052), .ZN(n17228) );
  BUF_X2 U10187 ( .I(n16462), .Z(n6295) );
  INV_X4 U8464 ( .I(n1636), .ZN(n20523) );
  INV_X2 U7605 ( .I(n11918), .ZN(n18714) );
  INV_X2 U11939 ( .I(n16777), .ZN(n3486) );
  BUF_X4 U2928 ( .I(n18300), .Z(n18722) );
  INV_X2 U929 ( .I(n18980), .ZN(n19257) );
  NAND3_X2 U8598 ( .A1(n761), .A2(n11959), .A3(n9724), .ZN(n4050) );
  BUF_X2 U4265 ( .I(n11605), .Z(n2990) );
  INV_X2 U12972 ( .I(n8741), .ZN(n9665) );
  OR2_X2 U11537 ( .A1(n16938), .A2(n16743), .Z(n21087) );
  BUF_X2 U6008 ( .I(Key[126]), .Z(n16561) );
  INV_X4 U7859 ( .I(n23843), .ZN(n5373) );
  NAND2_X2 U17098 ( .A1(n7830), .A2(n6082), .ZN(n8256) );
  INV_X4 U9215 ( .I(n5191), .ZN(n6661) );
  NOR2_X2 U8653 ( .A1(n8051), .A2(n16485), .ZN(n8831) );
  NAND2_X2 U6997 ( .A1(n8131), .A2(n3063), .ZN(n22531) );
  AOI21_X2 U10910 ( .A1(n17149), .A2(n17148), .B(n4652), .ZN(n4651) );
  INV_X4 U3538 ( .I(n22641), .ZN(n906) );
  AOI21_X2 U15433 ( .A1(n14478), .A2(n29360), .B(n29626), .ZN(n15328) );
  NAND2_X2 U13792 ( .A1(n1350), .A2(n2843), .ZN(n11838) );
  INV_X2 U7154 ( .I(n17956), .ZN(n7238) );
  INV_X2 U10041 ( .I(n19280), .ZN(n13377) );
  NAND2_X2 U3275 ( .A1(n6071), .A2(n27947), .ZN(n365) );
  OAI22_X2 U8218 ( .A1(n5048), .A2(n16779), .B1(n1142), .B2(n5049), .ZN(n13292) );
  INV_X2 U63 ( .I(n25397), .ZN(n14247) );
  OAI21_X2 U9143 ( .A1(n16540), .A2(n33103), .B(n16539), .ZN(n1819) );
  INV_X4 U6644 ( .I(n8802), .ZN(n879) );
  INV_X2 U9296 ( .I(n11626), .ZN(n8479) );
  OR3_X2 U4407 ( .A1(n1224), .A2(n33493), .A3(n31268), .Z(n25109) );
  AOI21_X2 U10762 ( .A1(n13342), .A2(n23510), .B(n23918), .ZN(n8983) );
  OR2_X2 U7737 ( .A1(n24870), .A2(n8492), .Z(n25149) );
  OAI21_X2 U24482 ( .A1(n20078), .A2(n1163), .B(n19381), .ZN(n19382) );
  NOR3_X2 U4893 ( .A1(n9511), .A2(n29683), .A3(n9514), .ZN(n9509) );
  NAND2_X1 U18961 ( .A1(n15129), .A2(n16228), .ZN(n21545) );
  NAND3_X1 U151 ( .A1(n11963), .A2(n24212), .A3(n24211), .ZN(n17420) );
  INV_X2 U22628 ( .I(n23855), .ZN(n23797) );
  INV_X2 U3609 ( .I(n23860), .ZN(n2752) );
  INV_X1 U6352 ( .I(n11629), .ZN(n10931) );
  INV_X2 U9066 ( .I(n24244), .ZN(n1233) );
  NAND3_X1 U5096 ( .A1(n8584), .A2(n8360), .A3(n17472), .ZN(n1772) );
  NAND2_X2 U10086 ( .A1(n24), .A2(n8335), .ZN(n19328) );
  AOI21_X2 U7765 ( .A1(n9257), .A2(n7203), .B(n15010), .ZN(n9256) );
  INV_X2 U564 ( .I(n14691), .ZN(n17139) );
  OAI21_X2 U8646 ( .A1(n4218), .A2(n4217), .B(n27818), .ZN(n4361) );
  NAND2_X2 U11986 ( .A1(n13938), .A2(n29437), .ZN(n13937) );
  NAND2_X2 U894 ( .A1(n8862), .A2(n24), .ZN(n15397) );
  INV_X2 U14002 ( .I(n5035), .ZN(n8967) );
  INV_X2 U6698 ( .I(n16420), .ZN(n7899) );
  OR2_X2 U15307 ( .A1(n21330), .A2(n7453), .Z(n21429) );
  OAI21_X2 U20976 ( .A1(n16016), .A2(n21781), .B(n17021), .ZN(n16014) );
  INV_X2 U7573 ( .I(n13514), .ZN(n18793) );
  NOR2_X2 U9409 ( .A1(n239), .A2(n904), .ZN(n2794) );
  INV_X2 U5245 ( .I(n25385), .ZN(n25331) );
  INV_X2 U2658 ( .I(n3629), .ZN(n11691) );
  NAND2_X2 U7013 ( .A1(n16884), .A2(n1296), .ZN(n7817) );
  INV_X1 U5272 ( .I(n7778), .ZN(n24012) );
  BUF_X2 U10253 ( .I(Key[134]), .Z(n24707) );
  INV_X2 U5434 ( .I(n4693), .ZN(n1156) );
  NAND3_X2 U9614 ( .A1(n8256), .A2(n27230), .A3(n1335), .ZN(n1882) );
  NAND2_X2 U4432 ( .A1(n24723), .A2(n25905), .ZN(n25838) );
  AOI21_X2 U5137 ( .A1(n19918), .A2(n19917), .B(n19916), .ZN(n20526) );
  INV_X2 U20250 ( .I(n10681), .ZN(n17201) );
  INV_X2 U14432 ( .I(n276), .ZN(n21522) );
  NAND2_X1 U14547 ( .A1(n17056), .A2(n25996), .ZN(n5634) );
  INV_X2 U4258 ( .I(n18631), .ZN(n16352) );
  INV_X2 U5515 ( .I(n5473), .ZN(n953) );
  AOI21_X2 U5740 ( .A1(n12107), .A2(n27865), .B(n6591), .ZN(n14466) );
  INV_X2 U7632 ( .I(n16585), .ZN(n18228) );
  NAND2_X2 U11698 ( .A1(n11838), .A2(n15434), .ZN(n10321) );
  INV_X2 U5492 ( .I(n5455), .ZN(n825) );
  NAND2_X2 U5134 ( .A1(n1815), .A2(n13772), .ZN(n4693) );
  INV_X2 U6509 ( .I(n14564), .ZN(n9062) );
  AOI22_X2 U7280 ( .A1(n20323), .A2(n5471), .B1(n8268), .B2(n15661), .ZN(
        n13850) );
  NAND2_X2 U5206 ( .A1(n11019), .A2(n25915), .ZN(n14170) );
  INV_X4 U7898 ( .I(n11821), .ZN(n1257) );
  INV_X2 U4238 ( .I(n11302), .ZN(n946) );
  NAND2_X2 U7143 ( .A1(n21120), .A2(n21429), .ZN(n21499) );
  NAND2_X2 U11293 ( .A1(n8006), .A2(n34087), .ZN(n1543) );
  NOR2_X2 U21194 ( .A1(n19883), .A2(n8616), .ZN(n17574) );
  OAI21_X2 U7781 ( .A1(n15179), .A2(n27436), .B(n24253), .ZN(n3604) );
  INV_X2 U16330 ( .I(n9690), .ZN(n5073) );
  AOI21_X2 U9999 ( .A1(n19034), .A2(n19088), .B(n10867), .ZN(n7316) );
  INV_X2 U4218 ( .I(n20110), .ZN(n19971) );
  INV_X2 U3197 ( .I(n25473), .ZN(n25470) );
  INV_X2 U7174 ( .I(n13304), .ZN(n17956) );
  NAND2_X1 U995 ( .A1(n6890), .A2(n10669), .ZN(n5560) );
  NOR2_X2 U5742 ( .A1(n30960), .A2(n15851), .ZN(n3689) );
  INV_X2 U850 ( .I(n20142), .ZN(n20036) );
  OAI21_X2 U10963 ( .A1(n11925), .A2(n16919), .B(n32766), .ZN(n16918) );
  BUF_X2 U8853 ( .I(Key[129]), .Z(n16578) );
  INV_X2 U9577 ( .I(n12452), .ZN(n21673) );
  OAI22_X2 U4756 ( .A1(n11064), .A2(n8731), .B1(n10687), .B2(n24223), .ZN(
        n9966) );
  AOI22_X2 U7147 ( .A1(n11487), .A2(n21255), .B1(n8757), .B2(n4633), .ZN(n7754) );
  INV_X2 U36 ( .I(n7702), .ZN(n25915) );
  AND2_X2 U19164 ( .A1(n10058), .A2(n18139), .Z(n9514) );
  INV_X2 U830 ( .I(n33264), .ZN(n6961) );
  INV_X2 U9694 ( .I(n18049), .ZN(n21428) );
  NOR2_X2 U4399 ( .A1(n13052), .A2(n6425), .ZN(n13051) );
  BUF_X4 U4979 ( .I(n25885), .Z(n4318) );
  OR2_X1 U19124 ( .A1(n20029), .A2(n19961), .Z(n16923) );
  INV_X1 U8092 ( .I(n22662), .ZN(n22660) );
  INV_X2 U4907 ( .I(n16782), .ZN(n13738) );
  OAI21_X2 U8972 ( .A1(n14922), .A2(n1213), .B(n16169), .ZN(n11786) );
  INV_X2 U25538 ( .I(n24883), .ZN(n25114) );
  INV_X2 U16068 ( .I(n4718), .ZN(n15038) );
  AOI21_X2 U7166 ( .A1(n21369), .A2(n1148), .B(n17522), .ZN(n4786) );
  AOI21_X2 U12107 ( .A1(n4043), .A2(n17874), .B(n16358), .ZN(n13502) );
  BUF_X2 U8345 ( .I(n6556), .Z(n3236) );
  NAND2_X2 U6932 ( .A1(n22814), .A2(n4678), .ZN(n9844) );
  NOR3_X1 U16468 ( .A1(n7224), .A2(n7225), .A3(n5239), .ZN(n18137) );
  NOR2_X2 U5983 ( .A1(n18676), .A2(n12290), .ZN(n18553) );
  INV_X2 U13028 ( .I(n15502), .ZN(n19269) );
  AND2_X2 U323 ( .A1(n5971), .A2(n11669), .Z(n11668) );
  INV_X4 U18570 ( .I(n7965), .ZN(n17764) );
  BUF_X2 U4295 ( .I(Key[170]), .Z(n16598) );
  BUF_X4 U4502 ( .I(n13415), .Z(n5381) );
  AOI21_X2 U22012 ( .A1(n29435), .A2(n21763), .B(n21762), .ZN(n21764) );
  INV_X2 U716 ( .I(n28813), .ZN(n1023) );
  INV_X4 U1854 ( .I(n6416), .ZN(n15902) );
  AND2_X2 U7407 ( .A1(n10863), .A2(n571), .Z(n12075) );
  OAI21_X2 U3589 ( .A1(n29435), .A2(n21762), .B(n6751), .ZN(n12845) );
  INV_X1 U16150 ( .I(n22110), .ZN(n13802) );
  NAND2_X1 U10970 ( .A1(n3826), .A2(n27984), .ZN(n10970) );
  AOI22_X2 U23233 ( .A1(n15335), .A2(n16072), .B1(n4989), .B2(n21406), .ZN(
        n21299) );
  INV_X4 U7423 ( .I(n20156), .ZN(n940) );
  INV_X2 U11267 ( .I(n8291), .ZN(n1310) );
  INV_X2 U4688 ( .I(n5412), .ZN(n25922) );
  INV_X4 U9003 ( .I(n9127), .ZN(n5387) );
  NAND2_X2 U7582 ( .A1(n15108), .A2(n18018), .ZN(n18574) );
  INV_X4 U16901 ( .I(n25981), .ZN(n5834) );
  INV_X2 U18746 ( .I(n15009), .ZN(n14457) );
  AOI21_X2 U16955 ( .A1(n5896), .A2(n22606), .B(n2858), .ZN(n5958) );
  INV_X4 U23056 ( .I(n22427), .ZN(n22534) );
  INV_X2 U696 ( .I(n17731), .ZN(n1332) );
  INV_X4 U3424 ( .I(n19942), .ZN(n1164) );
  OAI21_X1 U19059 ( .A1(n8710), .A2(n8709), .B(n8708), .ZN(n8707) );
  NAND2_X1 U22888 ( .A1(n29216), .A2(n28876), .ZN(n14479) );
  INV_X1 U8083 ( .I(n645), .ZN(n22368) );
  BUF_X2 U6893 ( .I(n14398), .Z(n8525) );
  OR2_X2 U15560 ( .A1(n10390), .A2(n8469), .Z(n21061) );
  NOR2_X2 U9891 ( .A1(n10072), .A2(n20149), .ZN(n5550) );
  INV_X4 U4687 ( .I(n15483), .ZN(n16041) );
  INV_X2 U4715 ( .I(n9941), .ZN(n2886) );
  NAND2_X1 U8634 ( .A1(n2599), .A2(n2935), .ZN(n2598) );
  BUF_X2 U4173 ( .I(n21630), .Z(n16601) );
  BUF_X2 U8852 ( .I(Key[108]), .Z(n25878) );
  CLKBUF_X2 U4652 ( .I(Key[39]), .Z(n25167) );
  BUF_X2 U12251 ( .I(Key[22]), .Z(n16551) );
  BUF_X2 U12265 ( .I(Key[112]), .Z(n16454) );
  CLKBUF_X2 U4654 ( .I(Key[84]), .Z(n16612) );
  BUF_X2 U7662 ( .I(Key[154]), .Z(n16605) );
  BUF_X2 U8869 ( .I(Key[109]), .Z(n25038) );
  BUF_X2 U6000 ( .I(Key[130]), .Z(n25450) );
  CLKBUF_X2 U4290 ( .I(Key[123]), .Z(n24487) );
  CLKBUF_X2 U4276 ( .I(Key[88]), .Z(n16631) );
  BUF_X2 U8866 ( .I(Key[114]), .Z(n25311) );
  BUF_X2 U8864 ( .I(Key[142]), .Z(n16674) );
  BUF_X2 U8845 ( .I(Key[48]), .Z(n25541) );
  BUF_X2 U6001 ( .I(Key[169]), .Z(n25355) );
  BUF_X2 U10252 ( .I(Key[76]), .Z(n25693) );
  CLKBUF_X2 U4306 ( .I(Key[34]), .Z(n16502) );
  CLKBUF_X2 U4294 ( .I(Key[184]), .Z(n8487) );
  BUF_X2 U5532 ( .I(Key[85]), .Z(n16523) );
  BUF_X2 U10223 ( .I(Key[31]), .Z(n16584) );
  CLKBUF_X2 U4323 ( .I(Key[52]), .Z(n16550) );
  BUF_X2 U7673 ( .I(Key[24]), .Z(n16619) );
  CLKBUF_X2 U4301 ( .I(Key[94]), .Z(n16355) );
  BUF_X2 U7674 ( .I(Key[90]), .Z(n16662) );
  BUF_X2 U5531 ( .I(Key[166]), .Z(n16604) );
  BUF_X2 U8862 ( .I(Key[138]), .Z(n25500) );
  BUF_X2 U12258 ( .I(Key[148]), .Z(n16636) );
  BUF_X2 U10232 ( .I(Key[61]), .Z(n25879) );
  CLKBUF_X2 U2766 ( .I(Key[173]), .Z(n16390) );
  BUF_X2 U8863 ( .I(Key[64]), .Z(n16322) );
  BUF_X2 U6012 ( .I(Key[49]), .Z(n24759) );
  BUF_X2 U10235 ( .I(Key[30]), .Z(n24833) );
  CLKBUF_X2 U4319 ( .I(Key[162]), .Z(n25641) );
  BUF_X2 U7669 ( .I(Key[172]), .Z(n16527) );
  CLKBUF_X2 U4302 ( .I(Key[3]), .Z(n24065) );
  BUF_X2 U4902 ( .I(n18882), .Z(n17477) );
  INV_X1 U2900 ( .I(n270), .ZN(n17597) );
  CLKBUF_X4 U6717 ( .I(n17189), .Z(n1439) );
  CLKBUF_X2 U4267 ( .I(n11905), .Z(n4194) );
  INV_X1 U12253 ( .I(n16504), .ZN(n1392) );
  INV_X1 U12252 ( .I(n25274), .ZN(n1391) );
  INV_X2 U979 ( .I(n18485), .ZN(n18767) );
  CLKBUF_X1 U12179 ( .I(n12120), .Z(n16426) );
  INV_X1 U12118 ( .I(n13466), .ZN(n18749) );
  INV_X2 U10080 ( .I(n4392), .ZN(n5813) );
  CLKBUF_X4 U1929 ( .I(n8802), .Z(n24) );
  INV_X2 U5176 ( .I(n33986), .ZN(n764) );
  NAND2_X1 U21483 ( .A1(n19354), .A2(n19355), .ZN(n14708) );
  NAND2_X1 U23965 ( .A1(n18904), .A2(n32932), .ZN(n17606) );
  NAND2_X1 U10005 ( .A1(n824), .A2(n10229), .ZN(n10855) );
  NAND2_X1 U21154 ( .A1(n15869), .A2(n18449), .ZN(n15418) );
  AOI21_X1 U1531 ( .A1(n19366), .A2(n19365), .B(n19364), .ZN(n19367) );
  CLKBUF_X2 U11931 ( .I(n10696), .Z(n4233) );
  INV_X1 U11885 ( .I(n5267), .ZN(n5405) );
  NAND2_X1 U8558 ( .A1(n20111), .A2(n32408), .ZN(n7580) );
  INV_X1 U11742 ( .I(n20576), .ZN(n7706) );
  INV_X2 U788 ( .I(n15043), .ZN(n20338) );
  CLKBUF_X4 U1243 ( .I(n20339), .Z(n384) );
  NAND2_X1 U8386 ( .A1(n20554), .A2(n20553), .ZN(n20557) );
  NAND2_X1 U24702 ( .A1(n20540), .A2(n782), .ZN(n20408) );
  NOR2_X1 U4579 ( .A1(n1961), .A2(n6134), .ZN(n1960) );
  AOI21_X1 U2571 ( .A1(n5835), .A2(n15898), .B(n184), .ZN(n183) );
  BUF_X4 U4581 ( .I(n20968), .Z(n5024) );
  BUF_X2 U7228 ( .I(n20931), .Z(n21365) );
  INV_X2 U23648 ( .I(n21189), .ZN(n21419) );
  NOR2_X1 U23736 ( .A1(n28642), .A2(n1017), .ZN(n21065) );
  NAND2_X1 U8200 ( .A1(n8457), .A2(n21736), .ZN(n21737) );
  NAND2_X1 U11317 ( .A1(n9350), .A2(n27532), .ZN(n9448) );
  NAND3_X1 U9489 ( .A1(n21753), .A2(n1316), .A3(n21752), .ZN(n21757) );
  NAND2_X1 U11270 ( .A1(n6937), .A2(n6935), .ZN(n6600) );
  INV_X1 U5091 ( .I(n22100), .ZN(n9290) );
  INV_X1 U16077 ( .I(n15825), .ZN(n22214) );
  CLKBUF_X2 U4160 ( .I(n15606), .Z(n3977) );
  BUF_X2 U4545 ( .I(n22662), .Z(n16483) );
  BUF_X2 U8095 ( .I(n22412), .Z(n16240) );
  CLKBUF_X2 U4152 ( .I(n21869), .Z(n16447) );
  BUF_X2 U4137 ( .I(n22565), .Z(n16490) );
  BUF_X2 U11173 ( .I(n11986), .Z(n4100) );
  INV_X1 U9442 ( .I(n15805), .ZN(n22663) );
  NOR2_X1 U11197 ( .A1(n12530), .A2(n22403), .ZN(n22333) );
  INV_X2 U4539 ( .I(n16166), .ZN(n22484) );
  NOR2_X1 U8043 ( .A1(n8098), .A2(n1842), .ZN(n7662) );
  CLKBUF_X4 U4121 ( .I(n14600), .Z(n897) );
  INV_X2 U1887 ( .I(n23103), .ZN(n11399) );
  INV_X1 U25186 ( .I(n23027), .ZN(n23029) );
  NAND2_X1 U9246 ( .A1(n10790), .A2(n30573), .ZN(n4780) );
  CLKBUF_X2 U1109 ( .I(n14612), .Z(n6461) );
  BUF_X2 U7910 ( .I(n11205), .Z(n8659) );
  INV_X1 U1307 ( .I(n23246), .ZN(n5316) );
  INV_X1 U5048 ( .I(n13216), .ZN(n11776) );
  CLKBUF_X2 U4106 ( .I(n23925), .Z(n16121) );
  NAND2_X1 U25290 ( .A1(n23691), .A2(n23857), .ZN(n23543) );
  BUF_X2 U10827 ( .I(n17245), .Z(n13549) );
  INV_X1 U10719 ( .I(n7524), .ZN(n9137) );
  INV_X2 U196 ( .I(n4821), .ZN(n14399) );
  INV_X2 U17285 ( .I(n24177), .ZN(n8062) );
  INV_X2 U5678 ( .I(n24060), .ZN(n792) );
  NAND2_X1 U25391 ( .A1(n24139), .A2(n24141), .ZN(n24086) );
  NAND2_X1 U194 ( .A1(n17277), .A2(n24288), .ZN(n3767) );
  NOR2_X1 U10609 ( .A1(n794), .A2(n16356), .ZN(n17066) );
  INV_X1 U13127 ( .I(n13306), .ZN(n24277) );
  INV_X1 U10508 ( .I(n24842), .ZN(n3544) );
  BUF_X2 U5594 ( .I(n11973), .Z(n8307) );
  CLKBUF_X4 U3559 ( .I(n12871), .Z(n12358) );
  INV_X2 U18573 ( .I(n13763), .ZN(n9858) );
  NAND2_X1 U6766 ( .A1(n4407), .A2(n33976), .ZN(n8194) );
  NAND2_X1 U8934 ( .A1(n7678), .A2(n8608), .ZN(n7647) );
  OAI21_X1 U1508 ( .A1(n3922), .A2(n15598), .B(n25630), .ZN(n15597) );
  NAND2_X1 U8950 ( .A1(n25027), .A2(n25028), .ZN(n1549) );
  OR2_X1 U10394 ( .A1(n17782), .A2(n17778), .Z(n14309) );
  CLKBUF_X4 U8927 ( .I(n25478), .Z(n6310) );
  CLKBUF_X4 U4689 ( .I(n5412), .Z(n5411) );
  NAND2_X1 U25691 ( .A1(n25479), .A2(n6310), .ZN(n25477) );
  INV_X1 U10263 ( .I(n10385), .ZN(n10009) );
  CLKBUF_X2 U10248 ( .I(Key[55]), .Z(n16479) );
  BUF_X2 U4322 ( .I(Key[136]), .Z(n16482) );
  BUF_X2 U4318 ( .I(Key[139]), .Z(n25772) );
  BUF_X2 U4303 ( .I(Key[181]), .Z(n16613) );
  BUF_X2 U7672 ( .I(Key[73]), .Z(n23191) );
  BUF_X2 U4284 ( .I(Key[4]), .Z(n25218) );
  BUF_X2 U4307 ( .I(Key[16]), .Z(n16653) );
  BUF_X2 U8857 ( .I(Key[67]), .Z(n16649) );
  BUF_X2 U12269 ( .I(Key[186]), .Z(n16634) );
  BUF_X2 U4297 ( .I(Key[163]), .Z(n25908) );
  CLKBUF_X2 U4908 ( .I(Key[12]), .Z(n25266) );
  CLKBUF_X2 U4277 ( .I(Key[26]), .Z(n24907) );
  CLKBUF_X2 U4282 ( .I(Key[11]), .Z(n25009) );
  OAI21_X1 U24366 ( .A1(n18775), .A2(n18774), .B(n18773), .ZN(n18776) );
  INV_X1 U1367 ( .I(n21662), .ZN(n10345) );
  AOI21_X1 U8056 ( .A1(n22503), .A2(n628), .B(n3063), .ZN(n11737) );
  INV_X1 U1496 ( .I(n22897), .ZN(n10885) );
  INV_X1 U10750 ( .I(n23930), .ZN(n9262) );
  NOR2_X1 U9208 ( .A1(n7073), .A2(n17373), .ZN(n3873) );
  NAND2_X2 U134 ( .A1(n3547), .A2(n2361), .ZN(n24370) );
  BUF_X4 U935 ( .I(n16047), .Z(n5760) );
  INV_X2 U11576 ( .I(n8028), .ZN(n5394) );
  OAI21_X2 U11426 ( .A1(n21382), .A2(n21383), .B(n15985), .ZN(n21386) );
  OAI21_X2 U7592 ( .A1(n18755), .A2(n18605), .B(n18761), .ZN(n18607) );
  INV_X2 U22408 ( .I(n17970), .ZN(n18638) );
  OAI21_X2 U11312 ( .A1(n8706), .A2(n8705), .B(n34087), .ZN(n2355) );
  INV_X4 U21769 ( .I(n26891), .ZN(n16485) );
  OAI21_X2 U9724 ( .A1(n12809), .A2(n28085), .B(n12808), .ZN(n20287) );
  AOI22_X2 U17395 ( .A1(n14573), .A2(n14334), .B1(n16092), .B2(n14575), .ZN(
        n14084) );
  OAI21_X2 U21015 ( .A1(n20019), .A2(n16595), .B(n14083), .ZN(n14573) );
  NAND2_X1 U5514 ( .A1(n16450), .A2(n17649), .ZN(n5328) );
  INV_X2 U22855 ( .I(n31012), .ZN(n18702) );
  NAND2_X1 U8821 ( .A1(n18706), .A2(n18535), .ZN(n18432) );
  INV_X2 U22396 ( .I(n13360), .ZN(n16181) );
  INV_X1 U2642 ( .I(n18811), .ZN(n7496) );
  INV_X2 U1052 ( .I(n18638), .ZN(n955) );
  INV_X1 U5192 ( .I(n17649), .ZN(n18572) );
  AOI21_X1 U24268 ( .A1(n18848), .A2(n18845), .B(n18730), .ZN(n18409) );
  OAI21_X1 U21441 ( .A1(n16995), .A2(n955), .B(n14651), .ZN(n14328) );
  AOI21_X1 U12170 ( .A1(n28731), .A2(n4194), .B(n27958), .ZN(n10843) );
  NAND2_X1 U6684 ( .A1(n18891), .A2(n6783), .ZN(n14874) );
  NOR2_X1 U10145 ( .A1(n18679), .A2(n10669), .ZN(n5586) );
  INV_X1 U20800 ( .I(n12006), .ZN(n18698) );
  NOR2_X1 U5512 ( .A1(n10283), .A2(n10284), .ZN(n18692) );
  NOR2_X1 U5187 ( .A1(n32901), .A2(n12951), .ZN(n18832) );
  AOI21_X1 U7589 ( .A1(n16352), .A2(n31012), .B(n18701), .ZN(n13949) );
  NOR2_X1 U13035 ( .A1(n2107), .A2(n962), .ZN(n15694) );
  NOR2_X1 U5972 ( .A1(n13466), .A2(n29659), .ZN(n13110) );
  AOI21_X1 U976 ( .A1(n18804), .A2(n17114), .B(n11880), .ZN(n18810) );
  NAND2_X1 U14843 ( .A1(n18409), .A2(n18410), .ZN(n3844) );
  OAI21_X1 U7536 ( .A1(n14666), .A2(n15902), .B(n10133), .ZN(n10208) );
  OAI21_X1 U5988 ( .A1(n14651), .A2(n18637), .B(n18638), .ZN(n5459) );
  OAI21_X1 U20823 ( .A1(n18616), .A2(n12837), .B(n10043), .ZN(n18422) );
  NAND2_X1 U5969 ( .A1(n7682), .A2(n7681), .ZN(n18074) );
  INV_X1 U7563 ( .I(n12989), .ZN(n18824) );
  INV_X1 U12084 ( .I(n19224), .ZN(n1380) );
  INV_X2 U8701 ( .I(n4016), .ZN(n12502) );
  INV_X2 U924 ( .I(n34107), .ZN(n19228) );
  INV_X1 U6625 ( .I(n2150), .ZN(n19096) );
  INV_X1 U13321 ( .I(n12468), .ZN(n2412) );
  NAND3_X1 U3309 ( .A1(n2150), .A2(n18769), .A3(n17905), .ZN(n19200) );
  INV_X1 U6608 ( .I(n14597), .ZN(n18993) );
  INV_X1 U5493 ( .I(n19348), .ZN(n19217) );
  OAI22_X1 U24430 ( .A1(n19076), .A2(n19196), .B1(n19075), .B2(n27726), .ZN(
        n19077) );
  OAI21_X1 U16522 ( .A1(n5813), .A2(n10203), .B(n19200), .ZN(n13890) );
  OAI21_X1 U7520 ( .A1(n880), .A2(n19116), .B(n879), .ZN(n8864) );
  NAND2_X1 U22024 ( .A1(n4016), .A2(n19348), .ZN(n16335) );
  NOR2_X1 U1467 ( .A1(n19364), .A2(n19064), .ZN(n19065) );
  NAND2_X1 U18070 ( .A1(n1386), .A2(n11302), .ZN(n7133) );
  INV_X1 U9993 ( .I(n18123), .ZN(n3059) );
  NAND3_X1 U9995 ( .A1(n9318), .A2(n19210), .A3(n4202), .ZN(n9317) );
  BUF_X2 U4274 ( .I(Key[15]), .Z(n25049) );
  AOI21_X1 U24295 ( .A1(n18474), .A2(n28147), .B(n1378), .ZN(n18478) );
  INV_X1 U875 ( .I(n4704), .ZN(n8571) );
  CLKBUF_X2 U11961 ( .I(n19520), .Z(n16586) );
  INV_X1 U9959 ( .I(n5127), .ZN(n9988) );
  NAND2_X1 U22449 ( .A1(n13477), .A2(n13480), .ZN(n13479) );
  BUF_X2 U6003 ( .I(Key[190]), .Z(n16530) );
  INV_X1 U1304 ( .I(n19763), .ZN(n1364) );
  NOR2_X1 U13705 ( .A1(n2780), .A2(n20155), .ZN(n13912) );
  NOR2_X1 U7333 ( .A1(n5188), .A2(n19921), .ZN(n1957) );
  BUF_X2 U2738 ( .I(n16646), .Z(n12682) );
  INV_X1 U2452 ( .I(n6200), .ZN(n10750) );
  NOR3_X1 U22451 ( .A1(n19799), .A2(n19867), .A3(n19886), .ZN(n13489) );
  INV_X1 U5899 ( .I(n18142), .ZN(n20143) );
  NAND3_X1 U7383 ( .A1(n1167), .A2(n20080), .A3(n1359), .ZN(n2052) );
  INV_X1 U5903 ( .I(n565), .ZN(n19794) );
  NOR2_X1 U2873 ( .A1(n27655), .A2(n19900), .ZN(n20111) );
  INV_X1 U4220 ( .I(n16105), .ZN(n20013) );
  INV_X1 U821 ( .I(n8816), .ZN(n1166) );
  NOR2_X1 U14421 ( .A1(n11959), .A2(n5073), .ZN(n3526) );
  AOI21_X1 U1030 ( .A1(n20095), .A2(n579), .B(n10439), .ZN(n10394) );
  NAND3_X1 U21027 ( .A1(n761), .A2(n3530), .A3(n15189), .ZN(n13569) );
  NAND2_X1 U11791 ( .A1(n20124), .A2(n20018), .ZN(n17542) );
  OAI21_X1 U9943 ( .A1(n14644), .A2(n19987), .B(n5707), .ZN(n20622) );
  INV_X1 U21106 ( .I(n20507), .ZN(n17975) );
  NOR2_X1 U9804 ( .A1(n1350), .A2(n2843), .ZN(n20418) );
  NAND2_X1 U24729 ( .A1(n7291), .A2(n20607), .ZN(n20609) );
  NAND2_X1 U21397 ( .A1(n20554), .A2(n7486), .ZN(n13433) );
  INV_X1 U4863 ( .I(n20345), .ZN(n760) );
  NOR2_X1 U7272 ( .A1(n20517), .A2(n28011), .ZN(n17297) );
  NOR2_X1 U11707 ( .A1(n26424), .A2(n9025), .ZN(n8869) );
  NOR2_X1 U21403 ( .A1(n20334), .A2(n710), .ZN(n12880) );
  OAI21_X1 U11657 ( .A1(n782), .A2(n1863), .B(n20342), .ZN(n20349) );
  AOI22_X1 U8417 ( .A1(n20531), .A2(n33721), .B1(n11055), .B2(n930), .ZN(
        n11412) );
  NAND3_X1 U24665 ( .A1(n111), .A2(n8998), .A3(n4468), .ZN(n20217) );
  NAND3_X1 U24718 ( .A1(n14731), .A2(n14719), .A3(n32747), .ZN(n20504) );
  NAND2_X1 U7282 ( .A1(n8868), .A2(n29628), .ZN(n20350) );
  INV_X1 U3031 ( .I(n7330), .ZN(n7960) );
  NAND2_X1 U9682 ( .A1(n11733), .A2(n21391), .ZN(n11732) );
  NOR2_X1 U13593 ( .A1(n925), .A2(n1329), .ZN(n2676) );
  NAND2_X1 U5117 ( .A1(n601), .A2(n21221), .ZN(n21060) );
  NAND3_X1 U24848 ( .A1(n21147), .A2(n29901), .A3(n21218), .ZN(n21148) );
  NOR3_X1 U6426 ( .A1(n10837), .A2(n31614), .A3(n21387), .ZN(n8560) );
  NOR2_X1 U1500 ( .A1(n4274), .A2(n28668), .ZN(n9816) );
  NAND2_X1 U24801 ( .A1(n8028), .A2(n5395), .ZN(n20909) );
  INV_X1 U7195 ( .I(n15874), .ZN(n21289) );
  NAND3_X1 U8253 ( .A1(n26971), .A2(n31614), .A3(n17956), .ZN(n8170) );
  NAND2_X1 U8249 ( .A1(n14853), .A2(n21151), .ZN(n9378) );
  NOR2_X1 U7199 ( .A1(n15002), .A2(n510), .ZN(n9454) );
  NAND2_X1 U630 ( .A1(n8170), .A2(n21148), .ZN(n4863) );
  INV_X2 U9572 ( .I(n21789), .ZN(n21653) );
  NAND2_X1 U8228 ( .A1(n8457), .A2(n13652), .ZN(n10357) );
  NAND2_X1 U21419 ( .A1(n15838), .A2(n21653), .ZN(n21467) );
  INV_X1 U6407 ( .I(n12827), .ZN(n11394) );
  NAND2_X1 U6404 ( .A1(n196), .A2(n27954), .ZN(n21603) );
  OAI21_X1 U4549 ( .A1(n11362), .A2(n10254), .B(n26443), .ZN(n14878) );
  AOI21_X1 U9540 ( .A1(n16222), .A2(n21653), .B(n21592), .ZN(n3807) );
  INV_X1 U9563 ( .I(n21462), .ZN(n21520) );
  OAI21_X1 U9544 ( .A1(n3703), .A2(n17347), .B(n1013), .ZN(n3702) );
  NOR2_X1 U8212 ( .A1(n14577), .A2(n14640), .ZN(n21766) );
  NOR2_X1 U7107 ( .A1(n1009), .A2(n2296), .ZN(n15241) );
  OAI21_X1 U1632 ( .A1(n17734), .A2(n29864), .B(n28181), .ZN(n21728) );
  NAND2_X1 U11285 ( .A1(n27686), .A2(n13162), .ZN(n13161) );
  AOI21_X1 U9498 ( .A1(n21154), .A2(n21468), .B(n21705), .ZN(n21155) );
  INV_X1 U11236 ( .I(n9960), .ZN(n11694) );
  INV_X2 U8097 ( .I(n4581), .ZN(n16567) );
  INV_X1 U21725 ( .I(n22457), .ZN(n22659) );
  INV_X1 U6326 ( .I(n8919), .ZN(n4500) );
  NOR2_X1 U21228 ( .A1(n9910), .A2(n26292), .ZN(n18181) );
  INV_X1 U463 ( .I(n9592), .ZN(n16745) );
  INV_X1 U21801 ( .I(n22428), .ZN(n17626) );
  INV_X1 U5782 ( .I(n1125), .ZN(n12236) );
  INV_X1 U4834 ( .I(n22610), .ZN(n855) );
  INV_X1 U17763 ( .I(n16334), .ZN(n17473) );
  AOI21_X1 U5784 ( .A1(n22454), .A2(n22578), .B(n15020), .ZN(n15019) );
  NOR2_X1 U9433 ( .A1(n468), .A2(n12733), .ZN(n4560) );
  NAND2_X1 U25095 ( .A1(n27638), .A2(n30014), .ZN(n22502) );
  NAND3_X1 U22129 ( .A1(n2471), .A2(n22574), .A3(n22657), .ZN(n12887) );
  NOR2_X1 U25059 ( .A1(n1842), .A2(n25947), .ZN(n22325) );
  NOR2_X1 U11195 ( .A1(n1001), .A2(n2132), .ZN(n1523) );
  NAND2_X1 U18985 ( .A1(n22650), .A2(n22651), .ZN(n10928) );
  NOR2_X1 U10938 ( .A1(n32766), .A2(n28313), .ZN(n5096) );
  INV_X1 U17711 ( .I(n6605), .ZN(n17327) );
  NAND2_X1 U25137 ( .A1(n23043), .A2(n896), .ZN(n22757) );
  INV_X1 U7988 ( .I(n3898), .ZN(n17148) );
  INV_X1 U391 ( .I(n22655), .ZN(n22895) );
  OAI21_X1 U4816 ( .A1(n17161), .A2(n22977), .B(n28227), .ZN(n2078) );
  INV_X1 U4505 ( .I(n23262), .ZN(n23443) );
  AOI21_X1 U25120 ( .A1(n23158), .A2(n22693), .B(n22692), .ZN(n23425) );
  INV_X1 U3610 ( .I(n666), .ZN(n23847) );
  NOR2_X1 U22212 ( .A1(n14297), .A2(n23813), .ZN(n13056) );
  INV_X1 U6213 ( .I(n4408), .ZN(n16099) );
  INV_X2 U3193 ( .I(n23940), .ZN(n23823) );
  INV_X1 U22042 ( .I(n28765), .ZN(n23822) );
  NAND2_X1 U7856 ( .A1(n895), .A2(n31890), .ZN(n16211) );
  NAND2_X1 U21286 ( .A1(n14164), .A2(n23578), .ZN(n15642) );
  NAND2_X1 U21285 ( .A1(n23824), .A2(n23825), .ZN(n15615) );
  INV_X1 U6898 ( .I(n11922), .ZN(n7895) );
  NOR2_X1 U21320 ( .A1(n16496), .A2(n16343), .ZN(n13364) );
  NAND3_X1 U21291 ( .A1(n3241), .A2(n23848), .A3(n28365), .ZN(n13173) );
  NOR2_X1 U9186 ( .A1(n26641), .A2(n976), .ZN(n14939) );
  OAI21_X1 U12453 ( .A1(n1920), .A2(n15912), .B(n26416), .ZN(n5679) );
  INV_X1 U21315 ( .I(n24094), .ZN(n24103) );
  INV_X2 U181 ( .I(n29977), .ZN(n1237) );
  INV_X1 U4473 ( .I(n12904), .ZN(n12903) );
  NAND2_X1 U6830 ( .A1(n24315), .A2(n13232), .ZN(n14336) );
  INV_X1 U10579 ( .I(n17801), .ZN(n6632) );
  NAND3_X1 U9096 ( .A1(n15179), .A2(n14399), .A3(n16868), .ZN(n6633) );
  NAND2_X1 U13663 ( .A1(n14663), .A2(n24316), .ZN(n2745) );
  NAND2_X1 U6121 ( .A1(n9581), .A2(n34137), .ZN(n24059) );
  NAND3_X1 U14790 ( .A1(n28120), .A2(n7068), .A3(n28784), .ZN(n23989) );
  INV_X1 U4750 ( .I(n6484), .ZN(n1230) );
  NAND2_X1 U21085 ( .A1(n25897), .A2(n24607), .ZN(n14108) );
  NAND2_X1 U18574 ( .A1(n12042), .A2(n16397), .ZN(n7973) );
  NAND2_X1 U25737 ( .A1(n25701), .A2(n146), .ZN(n25702) );
  INV_X1 U21785 ( .I(n17117), .ZN(n24611) );
  NAND2_X1 U6051 ( .A1(n25708), .A2(n16413), .ZN(n13643) );
  OAI21_X1 U1261 ( .A1(n25147), .A2(n25148), .B(n25203), .ZN(n9028) );
  INV_X1 U21355 ( .I(n25329), .ZN(n24703) );
  NAND2_X1 U5224 ( .A1(n25630), .A2(n8773), .ZN(n11497) );
  NOR2_X1 U8920 ( .A1(n27113), .A2(n5926), .ZN(n10038) );
  NAND2_X1 U21943 ( .A1(n25278), .A2(n12431), .ZN(n17877) );
  INV_X1 U2759 ( .I(n7941), .ZN(n5901) );
  NAND3_X1 U8 ( .A1(n27113), .A2(n25577), .A3(n25575), .ZN(n10039) );
  NAND2_X1 U62 ( .A1(n13273), .A2(n14922), .ZN(n3792) );
  AND2_X1 U100 ( .A1(n1083), .A2(n25235), .Z(n25134) );
  AND2_X1 U101 ( .A1(n25695), .A2(n25628), .Z(n6468) );
  BUF_X2 U119 ( .I(n25325), .Z(n11366) );
  NOR2_X1 U132 ( .A1(n3565), .A2(n9195), .ZN(n26466) );
  NAND2_X1 U136 ( .A1(n14495), .A2(n25119), .ZN(n27625) );
  INV_X1 U168 ( .I(n24533), .ZN(n7796) );
  NAND3_X1 U182 ( .A1(n15876), .A2(n7150), .A3(n28296), .ZN(n3545) );
  NAND2_X1 U195 ( .A1(n23964), .A2(n10046), .ZN(n27961) );
  INV_X1 U245 ( .I(n24072), .ZN(n7891) );
  BUF_X2 U250 ( .I(n24014), .Z(n16535) );
  NOR2_X1 U259 ( .A1(n12904), .A2(n27430), .ZN(n10778) );
  OR2_X1 U267 ( .A1(n11041), .A2(n3421), .Z(n11997) );
  INV_X2 U297 ( .I(n3880), .ZN(n15011) );
  OR2_X1 U328 ( .A1(n23918), .A2(n6869), .Z(n26073) );
  NAND2_X1 U339 ( .A1(n26716), .A2(n23675), .ZN(n26211) );
  OR2_X1 U376 ( .A1(n32998), .A2(n3004), .Z(n26070) );
  AOI22_X1 U382 ( .A1(n23902), .A2(n23843), .B1(n28034), .B2(n11067), .ZN(
        n29081) );
  OAI21_X1 U394 ( .A1(n23892), .A2(n32657), .B(n26801), .ZN(n23581) );
  OR2_X1 U398 ( .A1(n16620), .A2(n4892), .Z(n26074) );
  NAND2_X1 U414 ( .A1(n28266), .A2(n29498), .ZN(n26801) );
  AOI21_X1 U441 ( .A1(n16343), .A2(n23832), .B(n7005), .ZN(n3448) );
  CLKBUF_X2 U479 ( .I(n29323), .Z(n28297) );
  NAND2_X1 U517 ( .A1(n4542), .A2(n4543), .ZN(n29160) );
  NAND2_X1 U540 ( .A1(n806), .A2(n4110), .ZN(n26422) );
  NOR2_X1 U547 ( .A1(n5982), .A2(n4399), .ZN(n26994) );
  NOR2_X1 U559 ( .A1(n22848), .A2(n31854), .ZN(n22940) );
  NAND2_X1 U572 ( .A1(n28680), .A2(n27752), .ZN(n28327) );
  OAI21_X1 U583 ( .A1(n29242), .A2(n27752), .B(n22992), .ZN(n9582) );
  INV_X2 U618 ( .I(n15704), .ZN(n802) );
  NAND2_X1 U683 ( .A1(n21972), .A2(n22277), .ZN(n21975) );
  AOI22_X1 U693 ( .A1(n22688), .A2(n2417), .B1(n6232), .B2(n2418), .ZN(n28205)
         );
  OR2_X1 U703 ( .A1(n22449), .A2(n16137), .Z(n22973) );
  OAI21_X1 U736 ( .A1(n10206), .A2(n28669), .B(n32493), .ZN(n1702) );
  OR2_X1 U754 ( .A1(n6976), .A2(n1284), .Z(n22449) );
  NOR2_X1 U761 ( .A1(n27122), .A2(n22476), .ZN(n27207) );
  OAI21_X1 U789 ( .A1(n22670), .A2(n1127), .B(n22558), .ZN(n27357) );
  NOR2_X1 U797 ( .A1(n22665), .A2(n22576), .ZN(n15020) );
  NAND2_X1 U824 ( .A1(n28924), .A2(n32078), .ZN(n22420) );
  OAI21_X1 U914 ( .A1(n3742), .A2(n26572), .B(n13490), .ZN(n5004) );
  NAND3_X1 U915 ( .A1(n27707), .A2(n4331), .A3(n27706), .ZN(n5075) );
  NOR2_X1 U921 ( .A1(n26438), .A2(n21673), .ZN(n26282) );
  INV_X1 U962 ( .I(n16194), .ZN(n1325) );
  NOR2_X1 U964 ( .A1(n21872), .A2(n7813), .ZN(n13162) );
  NOR2_X1 U982 ( .A1(n21865), .A2(n21738), .ZN(n28068) );
  NAND2_X1 U991 ( .A1(n27454), .A2(n17098), .ZN(n11856) );
  AND2_X1 U1029 ( .A1(n4234), .A2(n26163), .Z(n12036) );
  NOR2_X1 U1043 ( .A1(n1533), .A2(n21842), .ZN(n27816) );
  NAND2_X1 U1046 ( .A1(n14640), .A2(n29258), .ZN(n15171) );
  INV_X1 U1056 ( .I(n15414), .ZN(n1319) );
  NOR2_X1 U1065 ( .A1(n21370), .A2(n26506), .ZN(n26505) );
  NOR2_X1 U1077 ( .A1(n13593), .A2(n21368), .ZN(n26506) );
  AND2_X1 U1093 ( .A1(n28668), .A2(n17341), .Z(n11138) );
  NAND2_X1 U1105 ( .A1(n17466), .A2(n27382), .ZN(n27658) );
  NAND2_X1 U1111 ( .A1(n9191), .A2(n15522), .ZN(n26993) );
  NOR2_X1 U1113 ( .A1(n4755), .A2(n17271), .ZN(n2173) );
  NOR2_X1 U1123 ( .A1(n5239), .A2(n8028), .ZN(n26142) );
  NOR2_X1 U1125 ( .A1(n6082), .A2(n21202), .ZN(n14292) );
  NOR2_X1 U1136 ( .A1(n29256), .A2(n4518), .ZN(n26736) );
  NOR2_X1 U1143 ( .A1(n21402), .A2(n12654), .ZN(n28425) );
  AOI21_X1 U1148 ( .A1(n17305), .A2(n4145), .B(n17590), .ZN(n12232) );
  NAND2_X1 U1154 ( .A1(n21325), .A2(n21326), .ZN(n27684) );
  NOR2_X1 U1164 ( .A1(n2468), .A2(n5883), .ZN(n26412) );
  INV_X1 U1169 ( .I(n21168), .ZN(n27711) );
  NOR2_X1 U1173 ( .A1(n21136), .A2(n31965), .ZN(n28375) );
  NOR3_X1 U1198 ( .A1(n6255), .A2(n6230), .A3(n26232), .ZN(n19792) );
  NAND2_X1 U1204 ( .A1(n20352), .A2(n1153), .ZN(n26722) );
  NOR2_X1 U1210 ( .A1(n17329), .A2(n17328), .ZN(n12809) );
  AOI21_X1 U1236 ( .A1(n20410), .A2(n20332), .B(n6475), .ZN(n7953) );
  AND2_X1 U1240 ( .A1(n20345), .A2(n10717), .Z(n20540) );
  AND2_X1 U1244 ( .A1(n15230), .A2(n25966), .Z(n5029) );
  NAND2_X1 U1247 ( .A1(n2843), .A2(n14054), .ZN(n20273) );
  OR2_X1 U1279 ( .A1(n5781), .A2(n6610), .Z(n27876) );
  OR2_X1 U1292 ( .A1(n14179), .A2(n20450), .Z(n5498) );
  BUF_X2 U1305 ( .I(n17236), .Z(n29069) );
  NOR2_X1 U1320 ( .A1(n28199), .A2(n27374), .ZN(n27373) );
  NAND2_X1 U1331 ( .A1(n28001), .A2(n875), .ZN(n27569) );
  NAND3_X1 U1332 ( .A1(n20043), .A2(n20157), .A3(n20156), .ZN(n29225) );
  OR2_X1 U1339 ( .A1(n28645), .A2(n26547), .Z(n26007) );
  NAND2_X1 U1346 ( .A1(n20068), .A2(n15110), .ZN(n27716) );
  NAND3_X1 U1349 ( .A1(n761), .A2(n20155), .A3(n3486), .ZN(n19925) );
  NAND2_X1 U1352 ( .A1(n729), .A2(n18126), .ZN(n29034) );
  NAND2_X1 U1356 ( .A1(n14589), .A2(n11959), .ZN(n6067) );
  NAND2_X1 U1363 ( .A1(n20147), .A2(n783), .ZN(n27374) );
  NAND2_X1 U1376 ( .A1(n15189), .A2(n20155), .ZN(n9026) );
  AND2_X1 U1379 ( .A1(n12179), .A2(n2391), .Z(n26006) );
  NOR2_X1 U1380 ( .A1(n8576), .A2(n27491), .ZN(n9149) );
  NAND2_X1 U1391 ( .A1(n12077), .A2(n14306), .ZN(n9173) );
  NAND3_X1 U1404 ( .A1(n19990), .A2(n12895), .A3(n28876), .ZN(n3087) );
  NAND2_X1 U1409 ( .A1(n579), .A2(n570), .ZN(n28154) );
  NAND2_X1 U1430 ( .A1(n11333), .A2(n575), .ZN(n6859) );
  NOR2_X1 U1434 ( .A1(n16193), .A2(n1161), .ZN(n19939) );
  INV_X1 U1437 ( .I(n25997), .ZN(n10805) );
  INV_X1 U1449 ( .I(n19399), .ZN(n3195) );
  INV_X1 U1453 ( .I(n16349), .ZN(n27825) );
  OAI21_X1 U1463 ( .A1(n19260), .A2(n25971), .B(n19257), .ZN(n7419) );
  NOR2_X1 U1480 ( .A1(n19261), .A2(n33206), .ZN(n6343) );
  OAI22_X1 U1483 ( .A1(n32932), .A2(n11000), .B1(n7492), .B2(n825), .ZN(n26918) );
  OAI21_X1 U1514 ( .A1(n28528), .A2(n10124), .B(n3388), .ZN(n19604) );
  BUF_X4 U1567 ( .I(n2150), .Z(n26417) );
  OAI21_X1 U1574 ( .A1(n26717), .A2(n18893), .B(n13087), .ZN(n18555) );
  OAI21_X1 U1578 ( .A1(n13408), .A2(n4474), .B(n4677), .ZN(n28172) );
  NAND2_X1 U1580 ( .A1(n18893), .A2(n10579), .ZN(n28573) );
  NAND2_X1 U1583 ( .A1(n7345), .A2(n14892), .ZN(n1603) );
  OAI21_X1 U1584 ( .A1(n18778), .A2(n18619), .B(n16624), .ZN(n15004) );
  AOI21_X1 U1585 ( .A1(n12863), .A2(n10903), .B(n7496), .ZN(n18554) );
  AND2_X1 U1586 ( .A1(n18805), .A2(n18806), .Z(n26035) );
  OAI21_X1 U1590 ( .A1(n18805), .A2(n18650), .B(n27908), .ZN(n9786) );
  NAND2_X1 U1592 ( .A1(n3601), .A2(n27690), .ZN(n9539) );
  OAI21_X1 U1598 ( .A1(n18805), .A2(n17114), .B(n17465), .ZN(n27238) );
  NAND2_X1 U1599 ( .A1(n27384), .A2(n6118), .ZN(n6117) );
  NAND2_X1 U1609 ( .A1(n25981), .A2(n18683), .ZN(n19292) );
  NAND2_X1 U1612 ( .A1(n18895), .A2(n16420), .ZN(n27384) );
  NAND2_X1 U1613 ( .A1(n26444), .A2(n6887), .ZN(n4765) );
  NOR2_X1 U1634 ( .A1(n18808), .A2(n16474), .ZN(n27908) );
  NAND2_X1 U1637 ( .A1(n18742), .A2(n18706), .ZN(n18635) );
  NOR2_X1 U1640 ( .A1(n12951), .A2(n12006), .ZN(n13016) );
  BUF_X2 U1652 ( .I(n18780), .Z(n16417) );
  OAI22_X2 U1661 ( .A1(n30375), .A2(n20028), .B1(n16461), .B2(n16637), .ZN(
        n19940) );
  INV_X2 U1668 ( .I(n4066), .ZN(n6638) );
  NAND2_X2 U1674 ( .A1(n18623), .A2(n27129), .ZN(n11864) );
  NOR2_X1 U1676 ( .A1(n18900), .A2(n28171), .ZN(n28993) );
  INV_X2 U1679 ( .I(n19618), .ZN(n20150) );
  INV_X2 U1702 ( .I(n22667), .ZN(n13664) );
  INV_X2 U1703 ( .I(n22330), .ZN(n22672) );
  OAI22_X2 U1783 ( .A1(n20940), .A2(n3236), .B1(n5395), .B2(n7990), .ZN(n5396)
         );
  AOI22_X2 U1799 ( .A1(n1026), .A2(n7707), .B1(n7706), .B2(n26587), .ZN(n7709)
         );
  NAND2_X1 U1801 ( .A1(n3883), .A2(n734), .ZN(n11213) );
  NAND2_X1 U1835 ( .A1(n24585), .A2(n24588), .ZN(n26217) );
  INV_X2 U1839 ( .I(n21992), .ZN(n1714) );
  INV_X2 U1856 ( .I(n16267), .ZN(n722) );
  BUF_X2 U1862 ( .I(n22679), .Z(n16570) );
  AOI21_X2 U1864 ( .A1(n5832), .A2(n31402), .B(n722), .ZN(n27451) );
  INV_X2 U1865 ( .I(n23866), .ZN(n9741) );
  NAND3_X1 U1871 ( .A1(n17333), .A2(n21712), .A3(n32904), .ZN(n28995) );
  OAI21_X2 U1917 ( .A1(n13170), .A2(n32298), .B(n32299), .ZN(n11675) );
  NAND2_X1 U1935 ( .A1(n16955), .A2(n29180), .ZN(n26370) );
  CLKBUF_X2 U1939 ( .I(n4908), .Z(n27622) );
  NAND2_X1 U1995 ( .A1(n9365), .A2(n25653), .ZN(n7085) );
  OAI21_X1 U2003 ( .A1(n10745), .A2(n10744), .B(n25232), .ZN(n10743) );
  BUF_X2 U2025 ( .I(n25723), .Z(n9495) );
  INV_X1 U2026 ( .I(n27117), .ZN(n17453) );
  CLKBUF_X2 U2029 ( .I(n27117), .Z(n28784) );
  CLKBUF_X2 U2033 ( .I(n5544), .Z(n5466) );
  NOR2_X1 U2043 ( .A1(n4381), .A2(n28017), .ZN(n21420) );
  OAI21_X1 U2056 ( .A1(n5926), .A2(n6092), .B(n25569), .ZN(n6673) );
  NAND2_X1 U2075 ( .A1(n14443), .A2(n6003), .ZN(n17492) );
  CLKBUF_X2 U2081 ( .I(n2236), .Z(n28734) );
  INV_X1 U2090 ( .I(n26848), .ZN(n12643) );
  NOR2_X1 U2123 ( .A1(n22619), .A2(n29314), .ZN(n28320) );
  NOR2_X1 U2140 ( .A1(n15011), .A2(n24141), .ZN(n15052) );
  NOR2_X1 U2143 ( .A1(n13627), .A2(n14960), .ZN(n24967) );
  AND2_X1 U2149 ( .A1(n12329), .A2(n32900), .Z(n5867) );
  BUF_X2 U2174 ( .I(n24275), .Z(n28120) );
  NAND2_X1 U2176 ( .A1(n24277), .A2(n26247), .ZN(n24278) );
  INV_X2 U2178 ( .I(n691), .ZN(n13624) );
  AOI21_X1 U2183 ( .A1(n24587), .A2(n753), .B(n26217), .ZN(n10609) );
  NAND2_X1 U2184 ( .A1(n123), .A2(n17764), .ZN(n13417) );
  AND2_X1 U2186 ( .A1(n25062), .A2(n25057), .Z(n3123) );
  AND2_X1 U2187 ( .A1(n25063), .A2(n25062), .Z(n16377) );
  OR2_X1 U2193 ( .A1(n7915), .A2(n28343), .Z(n23655) );
  OR3_X1 U2205 ( .A1(n767), .A2(n24340), .A3(n24163), .Z(n7091) );
  NAND2_X1 U2299 ( .A1(n25250), .A2(n7929), .ZN(n15124) );
  NOR2_X1 U2300 ( .A1(n25250), .A2(n7929), .ZN(n5543) );
  NAND2_X1 U2301 ( .A1(n7929), .A2(n25258), .ZN(n25254) );
  OAI22_X1 U2305 ( .A1(n25569), .A2(n13624), .B1(n25568), .B2(n6092), .ZN(
        n6114) );
  NAND2_X1 U2307 ( .A1(n9616), .A2(n5226), .ZN(n24288) );
  NOR2_X1 U2315 ( .A1(n8307), .A2(n25756), .ZN(n26270) );
  OR2_X1 U2317 ( .A1(n25709), .A2(n25756), .Z(n26056) );
  NAND2_X1 U2327 ( .A1(n25082), .A2(n11360), .ZN(n25100) );
  NAND2_X1 U2329 ( .A1(n25057), .A2(n25058), .ZN(n27609) );
  NAND2_X1 U2339 ( .A1(n3569), .A2(n547), .ZN(n17023) );
  NOR2_X1 U2363 ( .A1(n10097), .A2(n31921), .ZN(n11181) );
  INV_X2 U2364 ( .I(n31921), .ZN(n9862) );
  AOI21_X1 U2370 ( .A1(n22626), .A2(n16170), .B(n17955), .ZN(n22627) );
  NOR2_X1 U2374 ( .A1(n22982), .A2(n12586), .ZN(n28318) );
  OR2_X1 U2385 ( .A1(n29317), .A2(n13694), .Z(n10293) );
  OR2_X1 U2396 ( .A1(n10724), .A2(n17638), .Z(n250) );
  NOR2_X1 U2428 ( .A1(n13343), .A2(n4151), .ZN(n17065) );
  NOR2_X1 U2440 ( .A1(n23566), .A2(n769), .ZN(n26464) );
  NOR2_X1 U2443 ( .A1(n17373), .A2(n3874), .ZN(n23675) );
  NOR2_X1 U2447 ( .A1(n25900), .A2(n25867), .ZN(n6981) );
  OAI21_X1 U2453 ( .A1(n7935), .A2(n24157), .B(n796), .ZN(n17602) );
  NOR2_X1 U2467 ( .A1(n1567), .A2(n2092), .ZN(n27514) );
  INV_X1 U2485 ( .I(n25060), .ZN(n25052) );
  AND2_X1 U2512 ( .A1(n25699), .A2(n25696), .Z(n12086) );
  OR2_X1 U2546 ( .A1(n22816), .A2(n16315), .Z(n15167) );
  INV_X1 U2547 ( .I(n24682), .ZN(n9386) );
  NAND2_X1 U2567 ( .A1(n5226), .A2(n11503), .ZN(n17232) );
  NAND3_X1 U2587 ( .A1(n9917), .A2(n25390), .A3(n24667), .ZN(n14062) );
  OAI21_X1 U2597 ( .A1(n17110), .A2(n25232), .B(n5468), .ZN(n6259) );
  BUF_X2 U2608 ( .I(n19624), .Z(n27395) );
  OR2_X1 U2609 ( .A1(n1511), .A2(n25973), .Z(n1508) );
  NOR2_X1 U2618 ( .A1(n21766), .A2(n6599), .ZN(n3796) );
  NAND2_X1 U2624 ( .A1(n12058), .A2(n1218), .ZN(n24894) );
  NAND2_X1 U2637 ( .A1(n15255), .A2(n17641), .ZN(n8901) );
  INV_X2 U2650 ( .I(n31894), .ZN(n23482) );
  NAND2_X1 U2655 ( .A1(n7093), .A2(n24163), .ZN(n2852) );
  INV_X1 U2671 ( .I(n25375), .ZN(n25361) );
  NOR2_X1 U2678 ( .A1(n20507), .A2(n16452), .ZN(n17760) );
  BUF_X2 U2681 ( .I(n16831), .Z(n28163) );
  INV_X1 U2690 ( .I(n12593), .ZN(n24010) );
  CLKBUF_X4 U2694 ( .I(n22125), .Z(n8356) );
  NAND3_X1 U2700 ( .A1(n12005), .A2(n16152), .A3(n32298), .ZN(n16409) );
  INV_X2 U2715 ( .I(n20819), .ZN(n20658) );
  AND2_X1 U2716 ( .A1(n19911), .A2(n12770), .Z(n25941) );
  INV_X1 U2732 ( .I(n9159), .ZN(n13345) );
  XOR2_X1 U2733 ( .A1(n22121), .A2(n16622), .Z(n25945) );
  INV_X2 U2737 ( .I(n10824), .ZN(n22030) );
  INV_X2 U2754 ( .I(n14002), .ZN(n23017) );
  INV_X1 U2755 ( .I(n22580), .ZN(n9913) );
  NOR3_X2 U2767 ( .A1(n12445), .A2(n17740), .A3(n12444), .ZN(n27176) );
  INV_X2 U2772 ( .I(n23945), .ZN(n1253) );
  NAND2_X2 U2793 ( .A1(n27660), .A2(n27439), .ZN(n27125) );
  INV_X2 U2794 ( .I(n24299), .ZN(n24304) );
  INV_X1 U2796 ( .I(n25325), .ZN(n25410) );
  INV_X2 U2801 ( .I(n25051), .ZN(n28070) );
  INV_X2 U2803 ( .I(n31939), .ZN(n27127) );
  NAND2_X2 U2805 ( .A1(n11786), .A2(n13267), .ZN(n27149) );
  NAND2_X1 U2815 ( .A1(n802), .A2(n22876), .ZN(n2028) );
  AND2_X1 U2825 ( .A1(n14864), .A2(n13345), .Z(n5078) );
  NAND2_X1 U2846 ( .A1(n10717), .A2(n10106), .ZN(n20342) );
  NOR2_X1 U2853 ( .A1(n1718), .A2(n25628), .ZN(n26563) );
  AND2_X1 U2864 ( .A1(n25795), .A2(n8678), .Z(n8676) );
  NAND2_X1 U2880 ( .A1(n6544), .A2(n5546), .ZN(n4358) );
  INV_X1 U2898 ( .I(n8533), .ZN(n26493) );
  NOR2_X1 U2906 ( .A1(n7811), .A2(n21872), .ZN(n10492) );
  NAND2_X1 U2909 ( .A1(n18727), .A2(n13279), .ZN(n26398) );
  AND2_X2 U2910 ( .A1(n18548), .A2(n18649), .Z(n18804) );
  NAND2_X1 U2939 ( .A1(n16194), .A2(n5016), .ZN(n8360) );
  NAND2_X1 U2951 ( .A1(n26244), .A2(n26242), .ZN(n17083) );
  NAND2_X1 U2955 ( .A1(n24251), .A2(n28553), .ZN(n12551) );
  INV_X2 U2977 ( .I(n13614), .ZN(n24421) );
  NAND3_X1 U2987 ( .A1(n125), .A2(n12563), .A3(n20329), .ZN(n12564) );
  NAND2_X1 U2988 ( .A1(n15571), .A2(n24031), .ZN(n15570) );
  NOR2_X1 U3013 ( .A1(n15278), .A2(n20095), .ZN(n15907) );
  CLKBUF_X1 U3020 ( .I(n19149), .Z(n25959) );
  CLKBUF_X12 U3022 ( .I(n23944), .Z(n16677) );
  INV_X1 U3028 ( .I(n15275), .ZN(n26715) );
  NOR3_X1 U3045 ( .A1(n32642), .A2(n21559), .A3(n6489), .ZN(n8007) );
  NOR2_X1 U3083 ( .A1(n12982), .A2(n3421), .ZN(n27863) );
  NAND2_X1 U3115 ( .A1(n17084), .A2(n23087), .ZN(n26244) );
  NAND3_X1 U3120 ( .A1(n26070), .A2(n31807), .A3(n33583), .ZN(n2992) );
  NOR2_X1 U3126 ( .A1(n19178), .A2(n29769), .ZN(n27273) );
  AOI21_X1 U3139 ( .A1(n12038), .A2(n25997), .B(n19998), .ZN(n26823) );
  AOI21_X2 U3149 ( .A1(n17268), .A2(n11202), .B(n34074), .ZN(n10167) );
  NAND2_X1 U3172 ( .A1(n12535), .A2(n28580), .ZN(n12140) );
  NAND2_X1 U3184 ( .A1(n3203), .A2(n21532), .ZN(n12347) );
  AOI21_X1 U3195 ( .A1(n14619), .A2(n16799), .B(n839), .ZN(n10112) );
  AND2_X2 U3253 ( .A1(n15216), .A2(n15347), .Z(n18543) );
  INV_X1 U3259 ( .I(n22970), .ZN(n23259) );
  INV_X1 U3279 ( .I(n26750), .ZN(n14373) );
  AND2_X2 U3290 ( .A1(n21224), .A2(n14934), .Z(n21317) );
  INV_X1 U3307 ( .I(n7810), .ZN(n1050) );
  NAND3_X1 U3308 ( .A1(n16274), .A2(n7810), .A3(n7680), .ZN(n2585) );
  NAND2_X1 U3312 ( .A1(n26806), .A2(n24244), .ZN(n2324) );
  NAND2_X1 U3319 ( .A1(n27685), .A2(n30832), .ZN(n26283) );
  OR2_X2 U3322 ( .A1(n10932), .A2(n14439), .Z(n21451) );
  BUF_X4 U3328 ( .I(n22856), .Z(n25979) );
  NAND2_X1 U3342 ( .A1(n15829), .A2(n22990), .ZN(n22619) );
  INV_X1 U3343 ( .I(n22990), .ZN(n14977) );
  INV_X1 U3373 ( .I(n21232), .ZN(n21132) );
  OR2_X2 U3376 ( .A1(n21232), .A2(n21228), .Z(n21302) );
  NAND2_X1 U3377 ( .A1(n1289), .A2(n9617), .ZN(n22336) );
  OAI21_X1 U3380 ( .A1(n18146), .A2(n27430), .B(n12903), .ZN(n15571) );
  OAI21_X1 U3396 ( .A1(n28157), .A2(n3340), .B(n3515), .ZN(n19003) );
  NAND2_X1 U3428 ( .A1(n9630), .A2(n29288), .ZN(n12613) );
  AND2_X2 U3451 ( .A1(n10891), .A2(n495), .Z(n18843) );
  INV_X1 U3454 ( .I(n495), .ZN(n1389) );
  NAND2_X1 U3457 ( .A1(n1318), .A2(n26439), .ZN(n26438) );
  OAI22_X1 U3475 ( .A1(n7219), .A2(n985), .B1(n7221), .B2(n9280), .ZN(n28402)
         );
  NAND3_X1 U3487 ( .A1(n21284), .A2(n33889), .A3(n33147), .ZN(n8866) );
  NOR2_X1 U3490 ( .A1(n7068), .A2(n31461), .ZN(n8665) );
  INV_X1 U3493 ( .I(n18076), .ZN(n16372) );
  AOI22_X2 U3494 ( .A1(n3522), .A2(n32021), .B1(n31551), .B2(n3521), .ZN(n3520) );
  NAND3_X1 U3512 ( .A1(n4071), .A2(n34013), .A3(n5275), .ZN(n10290) );
  NAND3_X1 U3517 ( .A1(n10106), .A2(n20344), .A3(n20345), .ZN(n27225) );
  BUF_X2 U3519 ( .I(n7811), .Z(n5383) );
  NAND2_X1 U3529 ( .A1(n24276), .A2(n24168), .ZN(n24167) );
  NAND2_X1 U3532 ( .A1(n25066), .A2(n12329), .ZN(n12487) );
  OAI21_X1 U3533 ( .A1(n24139), .A2(n24138), .B(n3880), .ZN(n6978) );
  INV_X1 U3539 ( .I(n2643), .ZN(n21468) );
  INV_X1 U3566 ( .I(n11217), .ZN(n26540) );
  BUF_X4 U3567 ( .I(n10260), .Z(n25985) );
  OAI21_X1 U3602 ( .A1(n28659), .A2(n30904), .B(n28318), .ZN(n17175) );
  NAND2_X1 U3605 ( .A1(n10360), .A2(n28697), .ZN(n22985) );
  NAND2_X1 U3634 ( .A1(n21070), .A2(n3192), .ZN(n21328) );
  AND3_X2 U3641 ( .A1(n21630), .A2(n21573), .A3(n21628), .Z(n3798) );
  NOR2_X1 U3647 ( .A1(n1327), .A2(n21707), .ZN(n27648) );
  BUF_X2 U3768 ( .I(n10772), .Z(n17906) );
  AND2_X2 U3772 ( .A1(n33531), .A2(n15393), .Z(n20148) );
  NAND2_X1 U3814 ( .A1(n4755), .A2(n26345), .ZN(n21081) );
  AOI21_X1 U3832 ( .A1(n25410), .A2(n16528), .B(n25411), .ZN(n26892) );
  CLKBUF_X1 U3843 ( .I(n24276), .Z(n26247) );
  AOI21_X1 U3847 ( .A1(n27734), .A2(n23943), .B(n13549), .ZN(n23326) );
  NAND2_X1 U3849 ( .A1(n23562), .A2(n33260), .ZN(n7141) );
  NOR2_X1 U3855 ( .A1(n23634), .A2(n28510), .ZN(n28509) );
  CLKBUF_X1 U3857 ( .I(n9490), .Z(n26290) );
  BUF_X2 U3872 ( .I(n31566), .Z(n26231) );
  CLKBUF_X2 U3875 ( .I(n6593), .Z(n27865) );
  BUF_X4 U3876 ( .I(n23051), .Z(n25994) );
  CLKBUF_X2 U3887 ( .I(n10402), .Z(n26292) );
  CLKBUF_X2 U3897 ( .I(n22036), .Z(n28411) );
  CLKBUF_X1 U3909 ( .I(n14730), .Z(n26899) );
  NAND2_X1 U3911 ( .A1(n21850), .A2(n13490), .ZN(n27005) );
  OAI21_X1 U3918 ( .A1(n16147), .A2(n31958), .B(n33766), .ZN(n2720) );
  BUF_X2 U3922 ( .I(n16147), .Z(n26904) );
  OAI21_X1 U3937 ( .A1(n5026), .A2(n5030), .B(n1160), .ZN(n5025) );
  NAND2_X1 U3946 ( .A1(n17882), .A2(n1170), .ZN(n4045) );
  CLKBUF_X2 U3956 ( .I(n6974), .Z(n28889) );
  INV_X1 U3981 ( .I(n16649), .ZN(n26002) );
  OAI22_X1 U3990 ( .A1(n11134), .A2(n11136), .B1(n14510), .B2(n11133), .ZN(
        n27047) );
  NAND3_X1 U3992 ( .A1(n24946), .A2(n26199), .A3(n26197), .ZN(n15249) );
  INV_X2 U4001 ( .I(n25723), .ZN(n16494) );
  NAND2_X1 U4014 ( .A1(n28738), .A2(n26892), .ZN(n695) );
  BUF_X4 U4015 ( .I(n7198), .Z(n25995) );
  NAND2_X1 U4020 ( .A1(n30269), .A2(n26390), .ZN(n28888) );
  NAND2_X1 U4024 ( .A1(n11254), .A2(n11253), .ZN(n17295) );
  NAND2_X1 U4025 ( .A1(n26281), .A2(n31822), .ZN(n14267) );
  NAND2_X1 U4035 ( .A1(n25760), .A2(n24729), .ZN(n12265) );
  INV_X1 U4036 ( .I(n28223), .ZN(n24734) );
  CLKBUF_X1 U4044 ( .I(n15528), .Z(n28634) );
  NOR2_X1 U4066 ( .A1(n32017), .A2(n27982), .ZN(n9398) );
  INV_X1 U4070 ( .I(n7511), .ZN(n27791) );
  NAND2_X1 U4072 ( .A1(n17069), .A2(n794), .ZN(n27267) );
  NOR2_X1 U4078 ( .A1(n7019), .A2(n1086), .ZN(n7018) );
  NAND2_X1 U4093 ( .A1(n31772), .A2(n27591), .ZN(n6767) );
  NOR2_X1 U4104 ( .A1(n6286), .A2(n1931), .ZN(n27854) );
  CLKBUF_X2 U4105 ( .I(n24308), .Z(n28590) );
  CLKBUF_X2 U4119 ( .I(n4821), .Z(n27436) );
  CLKBUF_X2 U4123 ( .I(n24110), .Z(n29010) );
  NAND2_X1 U4128 ( .A1(n28509), .A2(n28507), .ZN(n10383) );
  NAND2_X1 U4129 ( .A1(n17086), .A2(n23766), .ZN(n14587) );
  NAND2_X1 U4134 ( .A1(n27078), .A2(n1253), .ZN(n57) );
  NAND2_X1 U4163 ( .A1(n23116), .A2(n23115), .ZN(n26150) );
  CLKBUF_X2 U4168 ( .I(n23157), .Z(n29068) );
  INV_X1 U4174 ( .I(n8674), .ZN(n27321) );
  NAND2_X1 U4187 ( .A1(n23917), .A2(n6869), .ZN(n26533) );
  INV_X1 U4331 ( .I(n23458), .ZN(n29220) );
  INV_X1 U4335 ( .I(n23494), .ZN(n26924) );
  INV_X1 U4342 ( .I(n33265), .ZN(n28492) );
  INV_X1 U4348 ( .I(n28402), .ZN(n28401) );
  NOR2_X1 U4349 ( .A1(n26026), .A2(n28227), .ZN(n28862) );
  NAND2_X1 U4353 ( .A1(n2028), .A2(n2029), .ZN(n26336) );
  NAND2_X1 U4362 ( .A1(n27191), .A2(n29176), .ZN(n22054) );
  INV_X1 U4365 ( .I(n11084), .ZN(n2031) );
  OAI21_X1 U4379 ( .A1(n28778), .A2(n28777), .B(n23055), .ZN(n17458) );
  OAI21_X1 U4381 ( .A1(n26106), .A2(n29174), .B(n29173), .ZN(n27191) );
  NAND2_X1 U4383 ( .A1(n22051), .A2(n31824), .ZN(n29176) );
  NAND2_X1 U4391 ( .A1(n23029), .A2(n23028), .ZN(n27079) );
  INV_X1 U4392 ( .I(n17707), .ZN(n27969) );
  CLKBUF_X2 U4397 ( .I(n15633), .Z(n28891) );
  OR2_X1 U4418 ( .A1(n1271), .A2(n10528), .Z(n26104) );
  AND2_X1 U4423 ( .A1(n22780), .A2(n30925), .Z(n26106) );
  CLKBUF_X2 U4455 ( .I(n3670), .Z(n26169) );
  CLKBUF_X2 U4466 ( .I(n12700), .Z(n27389) );
  CLKBUF_X8 U4475 ( .I(n15829), .Z(n27752) );
  CLKBUF_X2 U4481 ( .I(n8040), .Z(n26868) );
  CLKBUF_X2 U4531 ( .I(n14307), .Z(n28635) );
  INV_X1 U4570 ( .I(n22217), .ZN(n26845) );
  CLKBUF_X2 U4590 ( .I(n22172), .Z(n28490) );
  INV_X1 U4597 ( .I(n22149), .ZN(n28465) );
  AND2_X1 U4604 ( .A1(n21597), .A2(n21596), .Z(n27120) );
  NAND2_X1 U4608 ( .A1(n26265), .A2(n26625), .ZN(n13539) );
  NAND2_X1 U4631 ( .A1(n26522), .A2(n27005), .ZN(n7240) );
  NAND2_X1 U4634 ( .A1(n3807), .A2(n15837), .ZN(n15836) );
  NOR2_X1 U4635 ( .A1(n26386), .A2(n13490), .ZN(n14871) );
  OAI21_X1 U4662 ( .A1(n21682), .A2(n2575), .B(n26341), .ZN(n21517) );
  NOR2_X1 U4673 ( .A1(n21682), .A2(n2575), .ZN(n3742) );
  NAND2_X1 U4680 ( .A1(n21509), .A2(n21510), .ZN(n26451) );
  NOR2_X1 U4682 ( .A1(n16327), .A2(n12866), .ZN(n17429) );
  CLKBUF_X2 U4691 ( .I(n21462), .Z(n28838) );
  NAND2_X1 U4707 ( .A1(n27720), .A2(n13313), .ZN(n13310) );
  NAND2_X1 U4708 ( .A1(n21255), .A2(n21259), .ZN(n28255) );
  NAND2_X1 U4710 ( .A1(n21255), .A2(n21257), .ZN(n21256) );
  INV_X1 U4711 ( .I(n27198), .ZN(n21292) );
  NAND2_X1 U4718 ( .A1(n20935), .A2(n20938), .ZN(n28298) );
  NAND2_X1 U4724 ( .A1(n28501), .A2(n32357), .ZN(n16934) );
  NOR2_X1 U4725 ( .A1(n21325), .A2(n1146), .ZN(n8012) );
  OR2_X1 U4739 ( .A1(n10546), .A2(n16034), .Z(n11700) );
  NAND2_X1 U4742 ( .A1(n17455), .A2(n21295), .ZN(n27305) );
  CLKBUF_X2 U4763 ( .I(n15226), .Z(n26407) );
  NOR2_X1 U4771 ( .A1(n7822), .A2(n510), .ZN(n9879) );
  CLKBUF_X2 U4778 ( .I(n14029), .Z(n26798) );
  CLKBUF_X2 U4788 ( .I(n6854), .Z(n27193) );
  CLKBUF_X4 U4796 ( .I(n20946), .Z(n29062) );
  INV_X1 U4799 ( .I(n8972), .ZN(n27200) );
  INV_X1 U4800 ( .I(n10508), .ZN(n20823) );
  NAND2_X1 U4806 ( .A1(n20272), .A2(n17658), .ZN(n27923) );
  CLKBUF_X2 U4807 ( .I(n20953), .Z(n28823) );
  NAND2_X1 U4831 ( .A1(n442), .A2(n1863), .ZN(n26296) );
  INV_X1 U4845 ( .I(n20601), .ZN(n27621) );
  NAND2_X1 U4848 ( .A1(n1160), .A2(n10431), .ZN(n27620) );
  NAND2_X1 U4857 ( .A1(n20383), .A2(n15162), .ZN(n26986) );
  NAND2_X1 U4861 ( .A1(n20419), .A2(n14054), .ZN(n19893) );
  NOR2_X1 U4869 ( .A1(n27105), .A2(n5748), .ZN(n443) );
  OR2_X1 U4871 ( .A1(n710), .A2(n28261), .Z(n12149) );
  NOR2_X1 U4911 ( .A1(n27301), .A2(n19842), .ZN(n27300) );
  NAND2_X1 U4915 ( .A1(n26825), .A2(n26823), .ZN(n28454) );
  OAI21_X1 U4916 ( .A1(n12682), .A2(n20136), .B(n28012), .ZN(n19837) );
  NAND2_X1 U4918 ( .A1(n3486), .A2(n27398), .ZN(n7473) );
  NOR2_X1 U4934 ( .A1(n31046), .A2(n16108), .ZN(n27019) );
  NOR2_X1 U4935 ( .A1(n29339), .A2(n1166), .ZN(n20017) );
  NOR2_X1 U4936 ( .A1(n6859), .A2(n17882), .ZN(n27301) );
  AND2_X1 U4943 ( .A1(n13488), .A2(n821), .Z(n26093) );
  INV_X2 U4965 ( .I(n11969), .ZN(n25997) );
  NAND2_X1 U4973 ( .A1(n29135), .A2(n29134), .ZN(n29133) );
  AOI21_X1 U4987 ( .A1(n12649), .A2(n16669), .B(n26043), .ZN(n50) );
  INV_X1 U4990 ( .I(n10398), .ZN(n29135) );
  NAND2_X1 U4991 ( .A1(n28498), .A2(n18297), .ZN(n18298) );
  NAND2_X1 U4994 ( .A1(n14611), .A2(n12549), .ZN(n28371) );
  NOR2_X1 U4997 ( .A1(n19214), .A2(n29963), .ZN(n28133) );
  NAND2_X1 U5000 ( .A1(n19092), .A2(n19093), .ZN(n27929) );
  INV_X2 U5006 ( .I(n2207), .ZN(n5491) );
  OAI21_X1 U5011 ( .A1(n13444), .A2(n958), .B(n16207), .ZN(n27857) );
  NAND2_X1 U5016 ( .A1(n18851), .A2(n18730), .ZN(n27762) );
  NAND2_X1 U5030 ( .A1(n18850), .A2(n18849), .ZN(n27761) );
  NAND2_X1 U5033 ( .A1(n18662), .A2(n17477), .ZN(n29239) );
  INV_X1 U5034 ( .I(n18858), .ZN(n28102) );
  CLKBUF_X2 U5041 ( .I(n954), .Z(n28707) );
  INV_X1 U5047 ( .I(n16691), .ZN(n28422) );
  CLKBUF_X2 U5050 ( .I(n488), .Z(n26810) );
  CLKBUF_X2 U5053 ( .I(n270), .Z(n27940) );
  CLKBUF_X2 U5056 ( .I(n18811), .Z(n28686) );
  INV_X1 U5059 ( .I(n25728), .ZN(n28711) );
  CLKBUF_X2 U5060 ( .I(n10114), .Z(n28344) );
  INV_X1 U5061 ( .I(n16527), .ZN(n28462) );
  INV_X1 U5063 ( .I(n25282), .ZN(n27672) );
  INV_X1 U5068 ( .I(n25079), .ZN(n26001) );
  NAND2_X1 U5069 ( .A1(n18662), .A2(n17478), .ZN(n11406) );
  CLKBUF_X1 U5092 ( .I(n8386), .Z(n28578) );
  AOI21_X1 U5104 ( .A1(n15956), .A2(n18487), .B(n9), .ZN(n18488) );
  NOR2_X1 U5105 ( .A1(n18635), .A2(n18743), .ZN(n16359) );
  AOI21_X1 U5123 ( .A1(n10669), .A2(n18679), .B(n10537), .ZN(n10829) );
  NOR2_X1 U5130 ( .A1(n4868), .A2(n5327), .ZN(n5644) );
  NOR2_X1 U5135 ( .A1(n18648), .A2(n18650), .ZN(n2430) );
  NAND2_X1 U5157 ( .A1(n2614), .A2(n16474), .ZN(n26594) );
  NAND2_X1 U5172 ( .A1(n31821), .A2(n18722), .ZN(n18724) );
  AOI22_X1 U5178 ( .A1(n16181), .A2(n28010), .B1(n29659), .B2(n13360), .ZN(
        n13444) );
  INV_X1 U5202 ( .I(n5032), .ZN(n3341) );
  NAND3_X1 U5203 ( .A1(n7714), .A2(n9766), .A3(n7713), .ZN(n12826) );
  NOR2_X1 U5222 ( .A1(n745), .A2(n19021), .ZN(n6059) );
  NOR2_X1 U5223 ( .A1(n6846), .A2(n7995), .ZN(n28929) );
  AND3_X1 U5235 ( .A1(n27743), .A2(n13925), .A3(n949), .Z(n26043) );
  NAND2_X1 U5256 ( .A1(n14354), .A2(n13475), .ZN(n274) );
  CLKBUF_X1 U5283 ( .I(n4632), .Z(n294) );
  NOR2_X1 U5316 ( .A1(n3790), .A2(n27805), .ZN(n28419) );
  CLKBUF_X2 U5327 ( .I(n567), .Z(n28423) );
  AND3_X1 U5339 ( .A1(n16108), .A2(n1161), .A3(n13605), .Z(n6073) );
  NAND2_X1 U5340 ( .A1(n19456), .A2(n16681), .ZN(n19846) );
  NOR2_X1 U5374 ( .A1(n10613), .A2(n28904), .ZN(n28269) );
  NAND2_X1 U5405 ( .A1(n19906), .A2(n17790), .ZN(n15256) );
  NOR2_X1 U5412 ( .A1(n8031), .A2(n7577), .ZN(n3750) );
  NAND2_X1 U5423 ( .A1(n20564), .A2(n12263), .ZN(n20568) );
  NOR2_X1 U5435 ( .A1(n20418), .A2(n20417), .ZN(n20422) );
  INV_X1 U5444 ( .I(n20917), .ZN(n20809) );
  INV_X1 U5447 ( .I(n5724), .ZN(n10109) );
  NOR2_X1 U5486 ( .A1(n8190), .A2(n21095), .ZN(n17841) );
  NOR2_X1 U5504 ( .A1(n26677), .A2(n26635), .ZN(n7225) );
  NAND2_X1 U5513 ( .A1(n17832), .A2(n21317), .ZN(n20373) );
  NAND2_X1 U5521 ( .A1(n4683), .A2(n27684), .ZN(n28549) );
  NAND2_X1 U5537 ( .A1(n21752), .A2(n15414), .ZN(n15412) );
  AOI21_X1 U5538 ( .A1(n9699), .A2(n28037), .B(n8197), .ZN(n15905) );
  NAND3_X1 U5546 ( .A1(n28737), .A2(n18218), .A3(n1019), .ZN(n10555) );
  NAND2_X1 U5563 ( .A1(n26993), .A2(n12643), .ZN(n12641) );
  NAND2_X1 U5569 ( .A1(n16544), .A2(n16543), .ZN(n14950) );
  AND2_X1 U5587 ( .A1(n32506), .A2(n21568), .Z(n3315) );
  INV_X1 U5588 ( .I(n22291), .ZN(n1903) );
  NOR2_X1 U5595 ( .A1(n21736), .A2(n21867), .ZN(n26298) );
  OAI22_X1 U5600 ( .A1(n11848), .A2(n14917), .B1(n21346), .B2(n8140), .ZN(
        n21347) );
  NAND3_X1 U5605 ( .A1(n15127), .A2(n31954), .A3(n21741), .ZN(n14041) );
  INV_X1 U5607 ( .I(n22005), .ZN(n22086) );
  INV_X1 U5614 ( .I(n21937), .ZN(n28941) );
  NAND2_X1 U5623 ( .A1(n22484), .A2(n6297), .ZN(n8594) );
  NOR2_X1 U5637 ( .A1(n6297), .A2(n22641), .ZN(n4300) );
  NAND3_X1 U5674 ( .A1(n11250), .A2(n16334), .A3(n27959), .ZN(n14069) );
  NOR2_X1 U5681 ( .A1(n22664), .A2(n27415), .ZN(n22437) );
  NOR2_X1 U5684 ( .A1(n898), .A2(n32595), .ZN(n10645) );
  NAND2_X1 U5690 ( .A1(n7819), .A2(n28131), .ZN(n135) );
  INV_X1 U5706 ( .I(n23051), .ZN(n28555) );
  INV_X1 U5710 ( .I(n30234), .ZN(n1267) );
  NAND2_X1 U5719 ( .A1(n2937), .A2(n8308), .ZN(n26590) );
  AOI21_X1 U5725 ( .A1(n17707), .A2(n23026), .B(n6190), .ZN(n6189) );
  INV_X2 U5743 ( .I(n13694), .ZN(n23158) );
  INV_X1 U5748 ( .I(n23196), .ZN(n23216) );
  INV_X1 U5757 ( .I(n11897), .ZN(n10218) );
  INV_X1 U5761 ( .I(n528), .ZN(n26888) );
  INV_X1 U5763 ( .I(n23447), .ZN(n27080) );
  INV_X1 U5773 ( .I(n29178), .ZN(n15971) );
  NAND2_X1 U5797 ( .A1(n23855), .A2(n29178), .ZN(n9167) );
  INV_X1 U5808 ( .I(n9490), .ZN(n10967) );
  INV_X1 U5810 ( .I(n23851), .ZN(n8615) );
  NOR2_X1 U5816 ( .A1(n27455), .A2(n1099), .ZN(n14119) );
  INV_X1 U5825 ( .I(n14350), .ZN(n300) );
  NOR2_X1 U5837 ( .A1(n23940), .A2(n31807), .ZN(n2563) );
  AND2_X1 U5845 ( .A1(n6394), .A2(n30282), .Z(n15017) );
  INV_X1 U5846 ( .I(n14193), .ZN(n23544) );
  NAND2_X1 U5866 ( .A1(n13260), .A2(n24004), .ZN(n2865) );
  NOR3_X1 U5885 ( .A1(n15011), .A2(n24084), .A3(n14913), .ZN(n24035) );
  NOR2_X1 U5896 ( .A1(n24288), .A2(n9625), .ZN(n24108) );
  OAI21_X1 U5898 ( .A1(n12402), .A2(n24140), .B(n24087), .ZN(n29184) );
  INV_X1 U5920 ( .I(n25115), .ZN(n27650) );
  OR2_X1 U5946 ( .A1(n10170), .A2(n27181), .Z(n15459) );
  NOR2_X1 U5958 ( .A1(n9198), .A2(n28096), .ZN(n7806) );
  NOR2_X1 U5963 ( .A1(n25900), .A2(n18219), .ZN(n6325) );
  NAND2_X1 U5975 ( .A1(n33919), .A2(n33915), .ZN(n28562) );
  NOR2_X1 U6014 ( .A1(n9611), .A2(n25234), .ZN(n9610) );
  NOR2_X1 U6038 ( .A1(n25390), .A2(n24867), .ZN(n24672) );
  NAND2_X1 U6052 ( .A1(n25316), .A2(n2236), .ZN(n17028) );
  CLKBUF_X1 U6054 ( .I(n24909), .Z(n14075) );
  INV_X1 U6087 ( .I(n25206), .ZN(n27920) );
  NAND2_X1 U6088 ( .A1(n25362), .A2(n25361), .ZN(n28517) );
  AOI21_X1 U6091 ( .A1(n7701), .A2(n25916), .B(n5411), .ZN(n11155) );
  INV_X1 U6096 ( .I(n25064), .ZN(n16911) );
  XNOR2_X1 U6103 ( .A1(n19518), .A2(n2980), .ZN(n26004) );
  XNOR2_X1 U6105 ( .A1(n19599), .A2(n25355), .ZN(n26005) );
  OR2_X1 U6107 ( .A1(n31721), .A2(n9831), .Z(n26008) );
  AND2_X1 U6120 ( .A1(n9329), .A2(n6129), .Z(n26012) );
  AND2_X1 U6123 ( .A1(n21400), .A2(n21398), .Z(n26013) );
  AND2_X1 U6125 ( .A1(n924), .A2(n1337), .Z(n26014) );
  XNOR2_X1 U6127 ( .A1(n16349), .A2(n702), .ZN(n26016) );
  OR3_X1 U6135 ( .A1(n11306), .A2(n11090), .A3(n25633), .Z(n26022) );
  AND2_X1 U6138 ( .A1(n11366), .A2(n25412), .Z(n26023) );
  XNOR2_X1 U6143 ( .A1(n6906), .A2(n25751), .ZN(n26028) );
  XOR2_X1 U6144 ( .A1(n33835), .A2(n23191), .Z(n26029) );
  XNOR2_X1 U6145 ( .A1(n20692), .A2(n16523), .ZN(n26030) );
  XNOR2_X1 U6148 ( .A1(n34016), .A2(n16506), .ZN(n26031) );
  XNOR2_X1 U6154 ( .A1(n19773), .A2(n24937), .ZN(n26032) );
  AND2_X1 U6155 ( .A1(n1672), .A2(n1671), .Z(n26033) );
  INV_X1 U6158 ( .I(n8376), .ZN(n18791) );
  AND2_X1 U6162 ( .A1(n23754), .A2(n22617), .Z(n26036) );
  AND2_X1 U6169 ( .A1(n28958), .A2(n15528), .Z(n26038) );
  CLKBUF_X2 U6173 ( .I(n5748), .Z(n26730) );
  OR2_X1 U6182 ( .A1(n20413), .A2(n20414), .Z(n26041) );
  XNOR2_X1 U6186 ( .A1(n356), .A2(n24573), .ZN(n26045) );
  INV_X1 U6192 ( .I(n18557), .ZN(n18775) );
  XOR2_X1 U6211 ( .A1(n33835), .A2(n25908), .Z(n26053) );
  XOR2_X1 U6212 ( .A1(n12376), .A2(n24738), .Z(n26054) );
  XNOR2_X1 U6214 ( .A1(n19712), .A2(n24943), .ZN(n26055) );
  XNOR2_X1 U6215 ( .A1(n22226), .A2(n16691), .ZN(n26057) );
  XNOR2_X1 U6221 ( .A1(n20861), .A2(n16479), .ZN(n26058) );
  XNOR2_X1 U6222 ( .A1(n23476), .A2(n25167), .ZN(n26059) );
  NAND2_X1 U6225 ( .A1(n23842), .A2(n23887), .ZN(n26060) );
  AND2_X1 U6226 ( .A1(n25278), .A2(n16291), .Z(n26061) );
  AND2_X1 U6232 ( .A1(n16170), .A2(n16306), .Z(n26065) );
  AND2_X1 U6234 ( .A1(n12500), .A2(n13925), .Z(n26067) );
  NAND2_X1 U6235 ( .A1(n31915), .A2(n976), .ZN(n26069) );
  OR2_X1 U6239 ( .A1(n10724), .A2(n16166), .Z(n26072) );
  XNOR2_X1 U6245 ( .A1(n7653), .A2(n20820), .ZN(n26075) );
  XNOR2_X1 U6250 ( .A1(n27156), .A2(n25735), .ZN(n26076) );
  AND3_X1 U6259 ( .A1(n791), .A2(n9964), .A3(n24220), .Z(n26079) );
  CLKBUF_X4 U6262 ( .I(n1484), .Z(n28227) );
  INV_X1 U6267 ( .I(n1484), .ZN(n26160) );
  NOR2_X1 U6279 ( .A1(n11051), .A2(n13080), .ZN(n26083) );
  XNOR2_X1 U6284 ( .A1(n12957), .A2(n9874), .ZN(n26085) );
  XNOR2_X1 U6293 ( .A1(n20732), .A2(n20731), .ZN(n26087) );
  AND2_X2 U6294 ( .A1(n19938), .A2(n16105), .Z(n26088) );
  XNOR2_X1 U6311 ( .A1(n17385), .A2(n25436), .ZN(n26094) );
  XNOR2_X1 U6316 ( .A1(n21994), .A2(n24623), .ZN(n26096) );
  XNOR2_X1 U6323 ( .A1(n22031), .A2(n25610), .ZN(n26097) );
  XNOR2_X1 U6333 ( .A1(n22130), .A2(n16472), .ZN(n26100) );
  XNOR2_X1 U6337 ( .A1(n4732), .A2(n25929), .ZN(n26101) );
  XNOR2_X1 U6341 ( .A1(n7477), .A2(n16423), .ZN(n26103) );
  XNOR2_X1 U6347 ( .A1(n7229), .A2(n12754), .ZN(n26108) );
  INV_X1 U6355 ( .I(n11983), .ZN(n29175) );
  XNOR2_X1 U6359 ( .A1(n24629), .A2(n24628), .ZN(n26111) );
  AND2_X2 U6369 ( .A1(n31957), .A2(n4646), .Z(n26113) );
  XNOR2_X1 U6372 ( .A1(n227), .A2(n6924), .ZN(n26115) );
  XNOR2_X1 U6374 ( .A1(n16162), .A2(n23364), .ZN(n26116) );
  XNOR2_X1 U6382 ( .A1(n23467), .A2(n14526), .ZN(n26118) );
  INV_X1 U6385 ( .I(n13308), .ZN(n23559) );
  INV_X1 U6389 ( .I(n24327), .ZN(n1093) );
  XOR2_X1 U6390 ( .A1(n14645), .A2(n25693), .Z(n26121) );
  XNOR2_X1 U6394 ( .A1(n33971), .A2(n25450), .ZN(n26123) );
  XNOR2_X1 U6397 ( .A1(n32623), .A2(n13858), .ZN(n26124) );
  OR2_X1 U6403 ( .A1(n25659), .A2(n25657), .Z(n26127) );
  XNOR2_X1 U6418 ( .A1(n8269), .A2(n7808), .ZN(n3393) );
  INV_X2 U6421 ( .I(n31451), .ZN(n19107) );
  NAND2_X1 U6422 ( .A1(n19063), .A2(n31451), .ZN(n19062) );
  AND2_X1 U6448 ( .A1(n32855), .A2(n10948), .Z(n25611) );
  XOR2_X1 U6463 ( .A1(n4397), .A2(n9505), .Z(n4395) );
  XOR2_X1 U6467 ( .A1(n22147), .A2(n28465), .Z(n6396) );
  NAND2_X2 U6475 ( .A1(n18032), .A2(n21279), .ZN(n22147) );
  NAND2_X1 U6488 ( .A1(n31654), .A2(n21777), .ZN(n4211) );
  XOR2_X1 U6489 ( .A1(n12422), .A2(n12032), .Z(n13084) );
  NOR2_X2 U6508 ( .A1(n29027), .A2(n29026), .ZN(n987) );
  XOR2_X1 U6542 ( .A1(n20779), .A2(n11374), .Z(n26140) );
  AOI21_X1 U6559 ( .A1(n24283), .A2(n16356), .B(n4151), .ZN(n3862) );
  XOR2_X1 U6575 ( .A1(n10289), .A2(n23498), .Z(n26145) );
  NOR2_X2 U6576 ( .A1(n12358), .A2(n24466), .ZN(n26334) );
  NAND2_X2 U6607 ( .A1(n26150), .A2(n26073), .ZN(n839) );
  INV_X2 U6624 ( .I(n26153), .ZN(n19942) );
  XOR2_X1 U6626 ( .A1(n9821), .A2(n9818), .Z(n26153) );
  XOR2_X1 U6630 ( .A1(n16035), .A2(n26154), .Z(n16682) );
  XOR2_X1 U6632 ( .A1(n21918), .A2(n21919), .Z(n26154) );
  XOR2_X1 U6645 ( .A1(n24394), .A2(n9907), .Z(n24395) );
  NOR2_X2 U6662 ( .A1(n11608), .A2(n12691), .ZN(n12313) );
  INV_X2 U6666 ( .I(n15393), .ZN(n27748) );
  XOR2_X1 U6669 ( .A1(n11092), .A2(n11093), .Z(n15393) );
  AOI21_X2 U6676 ( .A1(n4926), .A2(n5700), .B(n26156), .ZN(n4508) );
  INV_X2 U6759 ( .I(n26162), .ZN(n13989) );
  NAND2_X2 U6773 ( .A1(n17960), .A2(n16375), .ZN(n22505) );
  INV_X2 U6774 ( .I(n15053), .ZN(n26633) );
  NAND2_X2 U6802 ( .A1(n2902), .A2(n2692), .ZN(n19212) );
  NAND2_X2 U6803 ( .A1(n18309), .A2(n18308), .ZN(n2692) );
  NAND3_X1 U6809 ( .A1(n17373), .A2(n26775), .A3(n23945), .ZN(n23677) );
  NAND2_X2 U6821 ( .A1(n2771), .A2(n26165), .ZN(n20926) );
  XOR2_X1 U6824 ( .A1(n9790), .A2(n26168), .Z(n11100) );
  XOR2_X1 U6827 ( .A1(n22241), .A2(n12898), .Z(n26168) );
  XOR2_X1 U6829 ( .A1(n24512), .A2(n31866), .Z(n26502) );
  INV_X2 U6836 ( .I(n26170), .ZN(n5736) );
  NAND2_X2 U6842 ( .A1(n9806), .A2(n9804), .ZN(n25654) );
  XOR2_X1 U6868 ( .A1(n9761), .A2(n26172), .Z(n7657) );
  XOR2_X1 U6870 ( .A1(n21034), .A2(n11424), .Z(n26172) );
  XOR2_X1 U6873 ( .A1(n23343), .A2(n27041), .Z(n5314) );
  OAI21_X2 U6917 ( .A1(n27802), .A2(n822), .B(n16059), .ZN(n3962) );
  XNOR2_X1 U6926 ( .A1(n33699), .A2(n13519), .ZN(n29108) );
  OR2_X1 U6957 ( .A1(n20158), .A2(n26182), .Z(n10615) );
  XOR2_X1 U6958 ( .A1(n20893), .A2(n20890), .Z(n1686) );
  XOR2_X1 U6959 ( .A1(n20982), .A2(n20822), .Z(n20893) );
  XOR2_X1 U6960 ( .A1(n1944), .A2(n9880), .Z(n11062) );
  NAND2_X1 U7021 ( .A1(n6102), .A2(n23052), .ZN(n6101) );
  INV_X2 U7050 ( .I(n24158), .ZN(n9934) );
  OAI21_X2 U7054 ( .A1(n7377), .A2(n7378), .B(n16629), .ZN(n7376) );
  XOR2_X1 U7066 ( .A1(n5241), .A2(n5240), .Z(n26194) );
  NAND2_X1 U7076 ( .A1(n26198), .A2(n24955), .ZN(n26197) );
  OR2_X1 U7077 ( .A1(n24955), .A2(n24956), .Z(n26199) );
  OAI22_X1 U7080 ( .A1(n8073), .A2(n1075), .B1(n7554), .B2(n28736), .ZN(n14764) );
  NAND2_X1 U7090 ( .A1(n24244), .A2(n28374), .ZN(n24075) );
  NOR2_X2 U7095 ( .A1(n24330), .A2(n24331), .ZN(n24244) );
  NAND2_X2 U7102 ( .A1(n7447), .A2(n26202), .ZN(n14864) );
  XOR2_X1 U7105 ( .A1(n22203), .A2(n14787), .Z(n14786) );
  XOR2_X1 U7109 ( .A1(n32084), .A2(n22031), .Z(n22203) );
  NAND3_X2 U7123 ( .A1(n26204), .A2(n9147), .A3(n23981), .ZN(n9145) );
  NOR2_X1 U7141 ( .A1(n15070), .A2(n180), .ZN(n28773) );
  OR2_X2 U7159 ( .A1(n7918), .A2(n10390), .Z(n1783) );
  XOR2_X1 U7170 ( .A1(n7574), .A2(n26208), .Z(n681) );
  INV_X1 U7171 ( .I(n25880), .ZN(n26208) );
  XOR2_X1 U7182 ( .A1(n12473), .A2(n17194), .Z(n663) );
  XOR2_X1 U7197 ( .A1(n3619), .A2(n3618), .Z(n16961) );
  XOR2_X1 U7217 ( .A1(n26215), .A2(n19388), .Z(n15476) );
  XOR2_X1 U7219 ( .A1(n19387), .A2(n19567), .Z(n26215) );
  XOR2_X1 U7220 ( .A1(n24654), .A2(n24683), .Z(n16930) );
  NAND2_X1 U7274 ( .A1(n16954), .A2(n15296), .ZN(n28) );
  XOR2_X1 U7303 ( .A1(n23457), .A2(n23404), .Z(n23314) );
  NAND2_X2 U7309 ( .A1(n14610), .A2(n22738), .ZN(n23457) );
  AOI22_X2 U7320 ( .A1(n26228), .A2(n20877), .B1(n21691), .B2(n5628), .ZN(
        n22056) );
  NAND3_X2 U7323 ( .A1(n31927), .A2(n21), .A3(n13115), .ZN(n26228) );
  XOR2_X1 U7349 ( .A1(n5856), .A2(n26233), .Z(n11068) );
  XOR2_X1 U7350 ( .A1(n4975), .A2(n3870), .Z(n26233) );
  XOR2_X1 U7395 ( .A1(n5563), .A2(n5562), .Z(n26237) );
  NOR2_X2 U7399 ( .A1(n26239), .A2(n26238), .ZN(n2285) );
  NOR2_X2 U7400 ( .A1(n5825), .A2(n17882), .ZN(n26239) );
  NAND2_X1 U7405 ( .A1(n27934), .A2(n8125), .ZN(n5079) );
  OAI21_X2 U7409 ( .A1(n26241), .A2(n23946), .B(n23950), .ZN(n3554) );
  NOR2_X2 U7422 ( .A1(n154), .A2(n1337), .ZN(n21099) );
  OAI22_X2 U7457 ( .A1(n1857), .A2(n28784), .B1(n13324), .B2(n17453), .ZN(
        n13586) );
  XOR2_X1 U7480 ( .A1(Plaintext[82]), .A2(Key[82]), .Z(n26249) );
  AOI21_X2 U7490 ( .A1(n18970), .A2(n12645), .B(n26250), .ZN(n19710) );
  NAND2_X1 U7533 ( .A1(n20481), .A2(n26566), .ZN(n8171) );
  XOR2_X1 U7542 ( .A1(n21946), .A2(n6245), .Z(n26256) );
  NAND2_X2 U7559 ( .A1(n27741), .A2(n32594), .ZN(n13867) );
  NAND2_X1 U7610 ( .A1(n18150), .A2(n18151), .ZN(n12230) );
  XOR2_X1 U7625 ( .A1(n26262), .A2(n15987), .Z(n8522) );
  XOR2_X1 U7633 ( .A1(n15986), .A2(n24373), .Z(n26262) );
  XOR2_X1 U7714 ( .A1(n11527), .A2(n11525), .Z(n18150) );
  NAND2_X2 U7727 ( .A1(n6432), .A2(n3894), .ZN(n28942) );
  NAND3_X2 U7728 ( .A1(n7961), .A2(n27627), .A3(n17992), .ZN(n7330) );
  AOI21_X2 U7733 ( .A1(n26268), .A2(n21430), .B(n7666), .ZN(n21617) );
  XOR2_X1 U7761 ( .A1(n15787), .A2(n6488), .Z(n6033) );
  XOR2_X1 U7770 ( .A1(n16792), .A2(n6028), .Z(n26272) );
  NAND2_X1 U7778 ( .A1(n29048), .A2(n29050), .ZN(n26275) );
  XOR2_X1 U7783 ( .A1(n26276), .A2(n7328), .Z(n20939) );
  XOR2_X1 U7784 ( .A1(n14522), .A2(n20687), .Z(n26276) );
  XOR2_X1 U7795 ( .A1(n16080), .A2(n14404), .Z(n5699) );
  XOR2_X1 U7800 ( .A1(n19626), .A2(n14293), .Z(n14404) );
  AOI21_X2 U7808 ( .A1(n17272), .A2(n21171), .B(n27424), .ZN(n27379) );
  NAND2_X2 U7813 ( .A1(n10232), .A2(n10233), .ZN(n22014) );
  INV_X4 U7825 ( .I(n26640), .ZN(n11940) );
  XOR2_X1 U7829 ( .A1(n28411), .A2(n27850), .Z(n4529) );
  INV_X2 U7839 ( .I(n26284), .ZN(n22429) );
  OR2_X1 U7854 ( .A1(n8044), .A2(n15518), .Z(n24605) );
  INV_X1 U7865 ( .I(n26439), .ZN(n21669) );
  AOI21_X2 U7878 ( .A1(n3128), .A2(n12178), .B(n26006), .ZN(n26291) );
  XOR2_X1 U7884 ( .A1(n26294), .A2(n24089), .Z(n24090) );
  XOR2_X1 U7885 ( .A1(n28258), .A2(n25619), .Z(n26294) );
  XOR2_X1 U7886 ( .A1(n26295), .A2(n16038), .Z(Ciphertext[93]) );
  NAND3_X2 U7902 ( .A1(n17420), .A2(n24214), .A3(n17676), .ZN(n24474) );
  OR2_X1 U7906 ( .A1(n28199), .A2(n16568), .Z(n9233) );
  XOR2_X1 U7908 ( .A1(n30319), .A2(n3589), .Z(n4003) );
  NAND2_X1 U7913 ( .A1(n31636), .A2(n29335), .ZN(n22573) );
  XOR2_X1 U7923 ( .A1(n26300), .A2(n2363), .Z(n3511) );
  AND2_X1 U7939 ( .A1(n27378), .A2(n7965), .Z(n26301) );
  OAI22_X1 U7942 ( .A1(n25667), .A2(n25666), .B1(n734), .B2(n25668), .ZN(
        n28052) );
  NOR2_X1 U7945 ( .A1(n11981), .A2(n7144), .ZN(n15215) );
  NAND3_X2 U7965 ( .A1(n26304), .A2(n27761), .A3(n27762), .ZN(n19206) );
  NAND3_X1 U7966 ( .A1(n6312), .A2(n6313), .A3(n957), .ZN(n26304) );
  NOR2_X2 U7976 ( .A1(n4856), .A2(n4857), .ZN(n18266) );
  XOR2_X1 U7983 ( .A1(n29030), .A2(n4157), .Z(n19491) );
  BUF_X2 U7995 ( .I(n7024), .Z(n26305) );
  AOI21_X2 U8004 ( .A1(n11436), .A2(n11437), .B(n26307), .ZN(n11439) );
  XOR2_X1 U8018 ( .A1(n23266), .A2(n30272), .Z(n6608) );
  XOR2_X1 U8061 ( .A1(n27290), .A2(n3476), .Z(n14142) );
  XOR2_X1 U8065 ( .A1(n21033), .A2(n9762), .Z(n9761) );
  OAI21_X2 U8075 ( .A1(n26318), .A2(n18573), .B(n29087), .ZN(n5478) );
  NAND2_X2 U8079 ( .A1(n951), .A2(n4868), .ZN(n12490) );
  NAND2_X2 U8084 ( .A1(n3181), .A2(n6555), .ZN(n24347) );
  NAND2_X2 U8106 ( .A1(n9917), .A2(n8105), .ZN(n24867) );
  NAND3_X2 U8107 ( .A1(n26362), .A2(n12215), .A3(n24860), .ZN(n24862) );
  NAND2_X2 U8112 ( .A1(n24436), .A2(n25696), .ZN(n25627) );
  NAND2_X2 U8123 ( .A1(n4075), .A2(n10056), .ZN(n11988) );
  OAI21_X2 U8126 ( .A1(n25539), .A2(n25536), .B(n17046), .ZN(n25297) );
  XOR2_X1 U8134 ( .A1(n6548), .A2(n16958), .Z(n20767) );
  AND2_X1 U8160 ( .A1(n15968), .A2(n20676), .Z(n26328) );
  XOR2_X1 U8185 ( .A1(n30628), .A2(n22014), .Z(n22027) );
  INV_X2 U8189 ( .I(n26330), .ZN(n522) );
  XOR2_X1 U8191 ( .A1(n5796), .A2(n13452), .Z(n26330) );
  INV_X2 U8216 ( .I(n26334), .ZN(n13326) );
  AND2_X1 U8225 ( .A1(n30978), .A2(n13114), .Z(n4433) );
  XOR2_X1 U8237 ( .A1(n26338), .A2(n10052), .Z(n10051) );
  OR2_X1 U8242 ( .A1(n20344), .A2(n10717), .Z(n20538) );
  NOR2_X1 U8243 ( .A1(n26445), .A2(n432), .ZN(n3168) );
  INV_X2 U8271 ( .I(n26340), .ZN(n11762) );
  NAND2_X2 U8279 ( .A1(n30995), .A2(n19224), .ZN(n19060) );
  OAI22_X2 U8337 ( .A1(n26355), .A2(n33635), .B1(n32951), .B2(n19185), .ZN(
        n11385) );
  NAND2_X2 U8347 ( .A1(n2612), .A2(n7687), .ZN(n13219) );
  AOI21_X2 U8350 ( .A1(n26357), .A2(n19868), .B(n941), .ZN(n19871) );
  NOR2_X2 U8360 ( .A1(n4633), .A2(n8757), .ZN(n5111) );
  NOR2_X2 U8362 ( .A1(n14556), .A2(n21053), .ZN(n4633) );
  XOR2_X1 U8380 ( .A1(n5436), .A2(n5434), .Z(n4060) );
  INV_X2 U8391 ( .I(n20555), .ZN(n28166) );
  OAI22_X2 U8392 ( .A1(n19881), .A2(n19880), .B1(n31046), .B2(n11119), .ZN(
        n20555) );
  XOR2_X1 U8410 ( .A1(n24440), .A2(n24664), .Z(n24596) );
  OAI21_X2 U8411 ( .A1(n2921), .A2(n7101), .B(n13046), .ZN(n24440) );
  NAND2_X1 U8421 ( .A1(n12217), .A2(n25689), .ZN(n26362) );
  NAND2_X2 U8428 ( .A1(n11795), .A2(n7457), .ZN(n22013) );
  XOR2_X1 U8436 ( .A1(n23282), .A2(n2520), .Z(n23408) );
  XOR2_X1 U8453 ( .A1(n26365), .A2(n8537), .Z(n9163) );
  BUF_X2 U8458 ( .I(n20117), .Z(n26368) );
  OAI22_X2 U8460 ( .A1(n26909), .A2(n2430), .B1(n2432), .B2(n16120), .ZN(
        n11203) );
  INV_X2 U8516 ( .I(n15839), .ZN(n28714) );
  XOR2_X1 U8519 ( .A1(n7032), .A2(n7029), .Z(n15839) );
  NOR2_X2 U8525 ( .A1(n23754), .A2(n1099), .ZN(n12432) );
  XOR2_X1 U8530 ( .A1(n32581), .A2(n31374), .Z(n20779) );
  INV_X1 U8543 ( .I(n19188), .ZN(n26376) );
  NOR2_X1 U8554 ( .A1(n18802), .A2(n33621), .ZN(n26378) );
  AOI21_X2 U8574 ( .A1(n20349), .A2(n760), .B(n27227), .ZN(n28813) );
  NAND2_X1 U8583 ( .A1(n28366), .A2(n5288), .ZN(n1864) );
  XOR2_X1 U8589 ( .A1(n8071), .A2(n26423), .Z(n23130) );
  XOR2_X1 U8616 ( .A1(n3411), .A2(n3410), .Z(n26385) );
  XOR2_X1 U8618 ( .A1(n24479), .A2(n12969), .Z(n24778) );
  NAND2_X2 U8619 ( .A1(n12403), .A2(n29184), .ZN(n12969) );
  NOR2_X2 U8625 ( .A1(n8984), .A2(n8983), .ZN(n26387) );
  NAND2_X1 U8638 ( .A1(n25144), .A2(n17595), .ZN(n16729) );
  NOR2_X2 U8647 ( .A1(n3698), .A2(n3695), .ZN(n14396) );
  AOI21_X2 U8654 ( .A1(n2176), .A2(n21172), .B(n2174), .ZN(n15172) );
  XOR2_X1 U8676 ( .A1(n10482), .A2(n9673), .Z(n26388) );
  NAND2_X2 U8710 ( .A1(n727), .A2(n7592), .ZN(n21712) );
  NOR2_X2 U8711 ( .A1(n1456), .A2(n1457), .ZN(n7592) );
  NAND2_X2 U8722 ( .A1(n26393), .A2(n22629), .ZN(n4734) );
  NOR2_X1 U8801 ( .A1(n6433), .A2(n31531), .ZN(n13835) );
  AOI22_X2 U8875 ( .A1(n26400), .A2(n28815), .B1(n24462), .B2(n8648), .ZN(
        n14931) );
  XOR2_X1 U8894 ( .A1(n32537), .A2(n22148), .Z(n5105) );
  NAND3_X2 U8904 ( .A1(n21505), .A2(n21510), .A3(n21506), .ZN(n21706) );
  NOR2_X2 U8910 ( .A1(n26772), .A2(n26408), .ZN(n17720) );
  INV_X1 U8921 ( .I(n15786), .ZN(n27098) );
  INV_X1 U8931 ( .I(n26585), .ZN(n20439) );
  INV_X2 U8941 ( .I(n12948), .ZN(n3874) );
  NAND2_X1 U8946 ( .A1(n26775), .A2(n12948), .ZN(n23943) );
  XOR2_X1 U8952 ( .A1(n6539), .A2(n12950), .Z(n12948) );
  AND2_X1 U8956 ( .A1(n16811), .A2(n20117), .Z(n19959) );
  INV_X2 U8964 ( .I(n11774), .ZN(n5805) );
  INV_X2 U8978 ( .I(n2022), .ZN(n26415) );
  AOI21_X2 U8992 ( .A1(n1563), .A2(n26373), .B(n27451), .ZN(n23387) );
  INV_X2 U8997 ( .I(n26418), .ZN(n18373) );
  XNOR2_X1 U8999 ( .A1(Key[41]), .A2(Plaintext[41]), .ZN(n26418) );
  XOR2_X1 U9009 ( .A1(n32537), .A2(n21923), .Z(n21577) );
  NOR2_X1 U9020 ( .A1(n8742), .A2(n9885), .ZN(n3022) );
  XOR2_X1 U9051 ( .A1(n23128), .A2(n23127), .Z(n26423) );
  XOR2_X1 U9104 ( .A1(n15161), .A2(n27125), .Z(n26429) );
  XOR2_X1 U9105 ( .A1(n12413), .A2(n19748), .Z(n4701) );
  XOR2_X1 U9128 ( .A1(n1259), .A2(n15130), .Z(n6706) );
  INV_X1 U9137 ( .I(n32917), .ZN(n840) );
  NAND2_X2 U9142 ( .A1(n990), .A2(n30297), .ZN(n11626) );
  INV_X4 U9145 ( .I(n10528), .ZN(n990) );
  INV_X2 U9150 ( .I(n26433), .ZN(n22427) );
  INV_X2 U9163 ( .I(n12701), .ZN(n22982) );
  OAI21_X2 U9164 ( .A1(n4503), .A2(n4504), .B(n4502), .ZN(n12701) );
  NAND3_X2 U9169 ( .A1(n6251), .A2(n6250), .A3(n26916), .ZN(n27439) );
  XOR2_X1 U9174 ( .A1(n26435), .A2(n17991), .Z(n17407) );
  NOR2_X1 U9192 ( .A1(n7867), .A2(n25941), .ZN(n8264) );
  XOR2_X1 U9197 ( .A1(n19505), .A2(n9138), .Z(n26436) );
  XOR2_X1 U9198 ( .A1(n11884), .A2(n6396), .Z(n6395) );
  NOR2_X2 U9203 ( .A1(n18941), .A2(n18942), .ZN(n19509) );
  NAND2_X1 U9209 ( .A1(n11390), .A2(n14926), .ZN(n11398) );
  NAND2_X1 U9210 ( .A1(n7941), .A2(n26440), .ZN(n434) );
  XOR2_X1 U9222 ( .A1(n8762), .A2(n25598), .Z(n10697) );
  NAND2_X1 U9245 ( .A1(n2105), .A2(n6891), .ZN(n26444) );
  NAND2_X1 U9250 ( .A1(n8373), .A2(n26774), .ZN(n20029) );
  XOR2_X1 U9292 ( .A1(n23370), .A2(n26452), .Z(n15612) );
  XOR2_X1 U9293 ( .A1(n32975), .A2(n6169), .Z(n26452) );
  NAND2_X1 U9294 ( .A1(n22665), .A2(n22576), .ZN(n26453) );
  XOR2_X1 U9298 ( .A1(n28460), .A2(n8548), .Z(n3621) );
  NAND2_X2 U9308 ( .A1(n14272), .A2(n14270), .ZN(n27954) );
  NOR2_X1 U9310 ( .A1(n26455), .A2(n27648), .ZN(n26690) );
  OAI21_X1 U9311 ( .A1(n27649), .A2(n230), .B(n32441), .ZN(n26455) );
  XOR2_X1 U9319 ( .A1(n3285), .A2(n3283), .Z(n26774) );
  NAND2_X2 U9327 ( .A1(n2593), .A2(n2595), .ZN(n26600) );
  XOR2_X1 U9330 ( .A1(n19490), .A2(n3415), .Z(n26456) );
  NOR2_X1 U9340 ( .A1(n1360), .A2(n1043), .ZN(n10273) );
  NAND2_X2 U9343 ( .A1(n18598), .A2(n26458), .ZN(n19330) );
  XNOR2_X1 U9353 ( .A1(n20801), .A2(n25881), .ZN(n29054) );
  XOR2_X1 U9400 ( .A1(n24390), .A2(n24472), .Z(n17653) );
  NAND2_X2 U9418 ( .A1(n13831), .A2(n26469), .ZN(n19074) );
  OAI21_X2 U9434 ( .A1(n15870), .A2(n9476), .B(n1389), .ZN(n26627) );
  AOI21_X2 U9457 ( .A1(n18809), .A2(n18650), .B(n26472), .ZN(n28944) );
  AND2_X1 U9459 ( .A1(n18648), .A2(n18349), .Z(n26472) );
  NOR2_X2 U9460 ( .A1(n2614), .A2(n18648), .ZN(n18809) );
  OR2_X1 U9494 ( .A1(n20393), .A2(n15468), .Z(n26478) );
  NAND2_X2 U9501 ( .A1(n24334), .A2(n3014), .ZN(n28202) );
  NOR2_X2 U9502 ( .A1(n1876), .A2(n1875), .ZN(n24334) );
  XOR2_X1 U9516 ( .A1(n20755), .A2(n26530), .Z(n13857) );
  INV_X1 U9521 ( .I(n8121), .ZN(n27768) );
  INV_X4 U9522 ( .I(n13412), .ZN(n791) );
  XOR2_X1 U9547 ( .A1(n8109), .A2(n24525), .Z(n8113) );
  XOR2_X1 U9562 ( .A1(n26484), .A2(n22247), .Z(n8471) );
  XOR2_X1 U9576 ( .A1(n13602), .A2(n27147), .Z(n13727) );
  NAND2_X2 U9578 ( .A1(n26485), .A2(n11037), .ZN(n20849) );
  XOR2_X1 U9592 ( .A1(n14682), .A2(n12671), .Z(n20796) );
  AND2_X1 U9595 ( .A1(n691), .A2(n8168), .Z(n12508) );
  XOR2_X1 U9604 ( .A1(n15726), .A2(n15725), .Z(n26487) );
  XOR2_X1 U9611 ( .A1(n5976), .A2(n29170), .Z(n5975) );
  XOR2_X1 U9630 ( .A1(n26490), .A2(n7652), .Z(n446) );
  XOR2_X1 U9634 ( .A1(n9665), .A2(n4314), .Z(n26490) );
  XOR2_X1 U9639 ( .A1(n26492), .A2(n21988), .Z(n29259) );
  XOR2_X1 U9641 ( .A1(n3723), .A2(n26493), .Z(n26492) );
  AOI22_X2 U9730 ( .A1(n16549), .A2(n22534), .B1(n12698), .B2(n17146), .ZN(
        n12697) );
  OR2_X1 U9731 ( .A1(n22655), .A2(n22951), .Z(n22862) );
  XOR2_X1 U9733 ( .A1(n26502), .A2(n7173), .Z(n29275) );
  NAND2_X2 U9748 ( .A1(n26505), .A2(n26504), .ZN(n16194) );
  BUF_X2 U9810 ( .I(n20137), .Z(n8558) );
  XOR2_X1 U9828 ( .A1(n26511), .A2(n11542), .Z(n8625) );
  INV_X2 U9847 ( .I(n26515), .ZN(n16333) );
  BUF_X2 U9859 ( .I(n12356), .Z(n26516) );
  AOI22_X2 U9861 ( .A1(n27696), .A2(n14734), .B1(n29223), .B2(n19203), .ZN(
        n8692) );
  XOR2_X1 U9862 ( .A1(n22295), .A2(n18189), .Z(n21944) );
  NAND2_X2 U9886 ( .A1(n26520), .A2(n16915), .ZN(n14831) );
  NAND2_X2 U9896 ( .A1(n25033), .A2(n26521), .ZN(n25044) );
  OAI21_X1 U9902 ( .A1(n25031), .A2(n14055), .B(n29334), .ZN(n26521) );
  NAND2_X2 U9922 ( .A1(n26524), .A2(n9453), .ZN(n13652) );
  INV_X2 U9936 ( .I(n26525), .ZN(n11513) );
  XNOR2_X1 U9940 ( .A1(n11514), .A2(n26977), .ZN(n26525) );
  NAND2_X2 U9965 ( .A1(n12515), .A2(n31470), .ZN(n20385) );
  AOI22_X2 U9968 ( .A1(n3571), .A2(n3401), .B1(n32004), .B2(n23577), .ZN(
        n24201) );
  NAND2_X2 U10063 ( .A1(n6332), .A2(n18810), .ZN(n2207) );
  XOR2_X1 U10077 ( .A1(n25998), .A2(n28479), .Z(n26534) );
  INV_X2 U10095 ( .I(n26537), .ZN(n7965) );
  OR2_X1 U10153 ( .A1(n14290), .A2(n21403), .Z(n4920) );
  XOR2_X1 U10154 ( .A1(n20848), .A2(n30304), .Z(n20671) );
  XOR2_X1 U10259 ( .A1(n12474), .A2(n23228), .Z(n12473) );
  XOR2_X1 U10261 ( .A1(n13864), .A2(n20715), .Z(n5184) );
  NAND2_X2 U10269 ( .A1(n9158), .A2(n9156), .ZN(n849) );
  NAND2_X1 U10290 ( .A1(n16111), .A2(n25790), .ZN(n12308) );
  XOR2_X1 U10323 ( .A1(n26552), .A2(n12552), .Z(n5166) );
  XOR2_X1 U10326 ( .A1(n20736), .A2(n31043), .Z(n26552) );
  XOR2_X1 U10327 ( .A1(n19449), .A2(n27824), .Z(n8435) );
  AOI22_X2 U10344 ( .A1(n3463), .A2(n3462), .B1(n26555), .B2(n28316), .ZN(
        n3461) );
  XOR2_X1 U10350 ( .A1(n3177), .A2(n3178), .Z(n3176) );
  XOR2_X1 U10360 ( .A1(n26556), .A2(n119), .Z(n24174) );
  XOR2_X1 U10362 ( .A1(n24405), .A2(n24649), .Z(n26556) );
  OR2_X1 U10364 ( .A1(n4632), .A2(n9469), .Z(n18126) );
  XOR2_X1 U10369 ( .A1(n4631), .A2(n29039), .Z(n4632) );
  OAI21_X2 U10379 ( .A1(n26557), .A2(n15849), .B(n15850), .ZN(n20329) );
  NOR2_X2 U10385 ( .A1(n15614), .A2(n14014), .ZN(n12904) );
  XOR2_X1 U10407 ( .A1(n21006), .A2(n16636), .Z(n27573) );
  OAI21_X2 U10410 ( .A1(n4469), .A2(n4471), .B(n20446), .ZN(n21006) );
  XOR2_X1 U10431 ( .A1(n23272), .A2(n25355), .Z(n643) );
  AND2_X1 U10433 ( .A1(n10599), .A2(n5822), .Z(n4248) );
  OAI21_X2 U10437 ( .A1(n26563), .A2(n6468), .B(n33120), .ZN(n6722) );
  AOI21_X2 U10445 ( .A1(n14163), .A2(n33787), .B(n14162), .ZN(n8726) );
  XOR2_X1 U10464 ( .A1(n23369), .A2(n27201), .Z(n16776) );
  OAI22_X1 U10478 ( .A1(n15167), .A2(n776), .B1(n22964), .B2(n15852), .ZN(
        n22820) );
  OAI22_X2 U10479 ( .A1(n26569), .A2(n17621), .B1(n7143), .B2(n25905), .ZN(
        n5412) );
  XOR2_X1 U10489 ( .A1(n5315), .A2(n5314), .Z(n5527) );
  AOI22_X2 U10494 ( .A1(n18807), .A2(n17465), .B1(n18809), .B2(n27909), .ZN(
        n6332) );
  XOR2_X1 U10496 ( .A1(n26571), .A2(n16634), .Z(Ciphertext[162]) );
  AND2_X1 U10501 ( .A1(n17370), .A2(n16699), .Z(n6030) );
  NOR2_X1 U10513 ( .A1(n16023), .A2(n30291), .ZN(n26572) );
  NAND2_X2 U10555 ( .A1(n26022), .A2(n26581), .ZN(n25664) );
  XOR2_X1 U10560 ( .A1(n2365), .A2(n7222), .Z(n2364) );
  OAI21_X1 U10567 ( .A1(n26290), .A2(n23862), .B(n13068), .ZN(n6235) );
  INV_X2 U10584 ( .I(n26583), .ZN(n13829) );
  XOR2_X1 U10591 ( .A1(n19520), .A2(n4157), .Z(n26583) );
  AOI21_X2 U10629 ( .A1(n15397), .A2(n13072), .B(n15395), .ZN(n19754) );
  AOI21_X2 U10649 ( .A1(n26589), .A2(n26588), .B(n10480), .ZN(n24004) );
  NAND2_X1 U10650 ( .A1(n17881), .A2(n32308), .ZN(n26588) );
  NAND2_X2 U10661 ( .A1(n3994), .A2(n14001), .ZN(n24926) );
  AOI21_X2 U10668 ( .A1(n28242), .A2(n13641), .B(n718), .ZN(n13636) );
  NAND2_X1 U10682 ( .A1(n26829), .A2(n5141), .ZN(n15422) );
  NOR2_X2 U10685 ( .A1(n11861), .A2(n31317), .ZN(n16016) );
  INV_X2 U10692 ( .I(n26593), .ZN(n29279) );
  XOR2_X1 U10693 ( .A1(n391), .A2(n13358), .Z(n26593) );
  NAND2_X2 U10694 ( .A1(n11199), .A2(n11198), .ZN(n10072) );
  AOI22_X1 U10713 ( .A1(n25812), .A2(n25816), .B1(n17642), .B2(n25811), .ZN(
        n25813) );
  INV_X2 U10731 ( .I(n26597), .ZN(n5961) );
  NOR2_X1 U10755 ( .A1(n26611), .A2(n16115), .ZN(n17115) );
  AOI21_X2 U10757 ( .A1(n25951), .A2(n28347), .B(n23796), .ZN(n2234) );
  INV_X2 U10795 ( .I(n18373), .ZN(n2614) );
  AND2_X1 U10832 ( .A1(n32253), .A2(n26640), .Z(n3643) );
  NAND2_X1 U10888 ( .A1(n16187), .A2(n16188), .ZN(n26614) );
  NAND2_X1 U10896 ( .A1(n2728), .A2(n15038), .ZN(n27064) );
  NOR2_X2 U10905 ( .A1(n15376), .A2(n5160), .ZN(n28525) );
  NOR2_X1 U10917 ( .A1(n16954), .A2(n29980), .ZN(n16953) );
  XOR2_X1 U10924 ( .A1(n3599), .A2(n16504), .Z(n26617) );
  NAND2_X2 U10934 ( .A1(n14758), .A2(n9256), .ZN(n24520) );
  NOR2_X2 U10951 ( .A1(n29224), .A2(n25678), .ZN(n25675) );
  XOR2_X1 U10997 ( .A1(n23041), .A2(n23040), .Z(n23720) );
  XOR2_X1 U11006 ( .A1(n22237), .A2(n21931), .Z(n10704) );
  OAI21_X1 U11010 ( .A1(n22641), .A2(n22484), .B(n9544), .ZN(n27445) );
  OAI21_X1 U11018 ( .A1(n9026), .A2(n9027), .B(n19974), .ZN(n26644) );
  INV_X1 U11021 ( .I(n26644), .ZN(n7474) );
  AOI21_X1 U11026 ( .A1(n3468), .A2(n17077), .B(n1135), .ZN(n26625) );
  INV_X4 U11053 ( .I(n25488), .ZN(n25462) );
  NAND2_X1 U11054 ( .A1(n4151), .A2(n13343), .ZN(n28275) );
  INV_X2 U11061 ( .I(n26630), .ZN(n3004) );
  NOR2_X2 U11068 ( .A1(n27446), .A2(n26631), .ZN(n24014) );
  XOR2_X1 U11081 ( .A1(n20808), .A2(n20807), .Z(n4849) );
  XOR2_X1 U11086 ( .A1(n30219), .A2(n20869), .Z(n20807) );
  NAND2_X2 U11087 ( .A1(n3499), .A2(n28380), .ZN(n3515) );
  AOI21_X1 U11104 ( .A1(n17120), .A2(n754), .B(n4407), .ZN(n26637) );
  NAND2_X2 U11130 ( .A1(n12650), .A2(n10100), .ZN(n10099) );
  NOR2_X2 U11133 ( .A1(n13502), .A2(n13501), .ZN(n26640) );
  XOR2_X1 U11152 ( .A1(n23471), .A2(n23472), .Z(n26642) );
  XOR2_X1 U11155 ( .A1(n26643), .A2(n17723), .Z(Ciphertext[157]) );
  AOI22_X1 U11163 ( .A1(n25750), .A2(n1979), .B1(n25734), .B2(n25733), .ZN(
        n26643) );
  XOR2_X1 U11181 ( .A1(n2875), .A2(n438), .Z(n26646) );
  NAND3_X2 U11198 ( .A1(n26648), .A2(n18536), .A3(n32530), .ZN(n19284) );
  NAND2_X1 U11203 ( .A1(n18256), .A2(n18745), .ZN(n26648) );
  XOR2_X1 U11218 ( .A1(n7452), .A2(n12805), .Z(n7646) );
  AOI22_X2 U11235 ( .A1(n28638), .A2(n29715), .B1(n3206), .B2(n13475), .ZN(
        n19197) );
  XOR2_X1 U11263 ( .A1(n26655), .A2(n22039), .Z(n10816) );
  XOR2_X1 U11272 ( .A1(n28730), .A2(n16060), .Z(n26655) );
  NAND2_X2 U11279 ( .A1(n4050), .A2(n4051), .ZN(n13911) );
  NAND2_X2 U11294 ( .A1(n9786), .A2(n9785), .ZN(n19224) );
  NAND2_X2 U11300 ( .A1(n5004), .A2(n10968), .ZN(n4342) );
  XOR2_X1 U11308 ( .A1(n24838), .A2(n24552), .Z(n18188) );
  AOI21_X2 U11360 ( .A1(n26007), .A2(n26741), .B(n942), .ZN(n26663) );
  XOR2_X1 U11370 ( .A1(n12736), .A2(n26665), .Z(n12735) );
  XOR2_X1 U11372 ( .A1(n20858), .A2(n10737), .Z(n26665) );
  NAND2_X1 U11394 ( .A1(n17467), .A2(n34089), .ZN(n12911) );
  INV_X1 U11395 ( .I(n26666), .ZN(n27862) );
  NAND3_X1 U11400 ( .A1(n25621), .A2(n11944), .A3(n25707), .ZN(n26666) );
  XOR2_X1 U11402 ( .A1(n27733), .A2(n23239), .Z(n2048) );
  NAND2_X1 U11406 ( .A1(n2107), .A2(n18676), .ZN(n3586) );
  XOR2_X1 U11424 ( .A1(n12495), .A2(n21921), .Z(n6329) );
  XOR2_X1 U11435 ( .A1(n29285), .A2(n7458), .Z(n3237) );
  NAND2_X2 U11458 ( .A1(n11560), .A2(n15836), .ZN(n22032) );
  INV_X2 U11462 ( .I(n10791), .ZN(n26677) );
  NAND2_X2 U11464 ( .A1(n26635), .A2(n26677), .ZN(n7990) );
  NOR2_X2 U11465 ( .A1(n1156), .A2(n26278), .ZN(n20321) );
  NOR2_X2 U11466 ( .A1(n28381), .A2(n28382), .ZN(n28380) );
  XOR2_X1 U11467 ( .A1(n29072), .A2(n27823), .Z(n7020) );
  OAI21_X2 U11476 ( .A1(n31975), .A2(n20480), .B(n26471), .ZN(n20316) );
  AOI21_X2 U11483 ( .A1(n1184), .A2(n13381), .B(n26680), .ZN(n6170) );
  NAND2_X2 U11484 ( .A1(n14651), .A2(n18638), .ZN(n6138) );
  NAND2_X2 U11486 ( .A1(n1214), .A2(n25889), .ZN(n7350) );
  XNOR2_X1 U11540 ( .A1(n20680), .A2(n20693), .ZN(n20859) );
  NAND2_X2 U11575 ( .A1(n25995), .A2(n30288), .ZN(n25882) );
  XOR2_X1 U11589 ( .A1(n3143), .A2(n3144), .Z(n15012) );
  NOR2_X1 U11592 ( .A1(n2902), .A2(n2692), .ZN(n14438) );
  NOR2_X1 U11593 ( .A1(n22674), .A2(n22467), .ZN(n8252) );
  XOR2_X1 U11609 ( .A1(n26692), .A2(n8312), .Z(n26691) );
  XOR2_X1 U11616 ( .A1(n3175), .A2(n26693), .Z(n22504) );
  XOR2_X1 U11617 ( .A1(n21906), .A2(n25945), .Z(n26693) );
  NAND2_X2 U11632 ( .A1(n26696), .A2(n19882), .ZN(n20515) );
  XOR2_X1 U11664 ( .A1(n3399), .A2(n26702), .Z(n577) );
  BUF_X2 U11695 ( .I(n709), .Z(n26710) );
  XOR2_X1 U11745 ( .A1(n26711), .A2(n16523), .Z(Ciphertext[13]) );
  OAI21_X2 U11774 ( .A1(n10686), .A2(n15002), .B(n151), .ZN(n14996) );
  OR2_X1 U11801 ( .A1(n13297), .A2(n5736), .Z(n7386) );
  OR2_X1 U11821 ( .A1(n26040), .A2(n26717), .Z(n3179) );
  XOR2_X1 U11840 ( .A1(n14215), .A2(n26055), .Z(n4895) );
  XOR2_X1 U11860 ( .A1(n10201), .A2(n16662), .Z(n23412) );
  NAND2_X2 U11888 ( .A1(n19298), .A2(n27831), .ZN(n14606) );
  INV_X2 U11895 ( .I(n11570), .ZN(n7929) );
  NAND2_X2 U11902 ( .A1(n15768), .A2(n17924), .ZN(n11570) );
  NOR2_X1 U11906 ( .A1(n15094), .A2(n16348), .ZN(n16347) );
  NAND2_X2 U11907 ( .A1(n19006), .A2(n18939), .ZN(n27077) );
  BUF_X2 U11922 ( .I(n24883), .Z(n25019) );
  INV_X4 U11930 ( .I(n3004), .ZN(n23940) );
  XOR2_X1 U11947 ( .A1(n12595), .A2(n14901), .Z(n15343) );
  NOR2_X1 U11977 ( .A1(n21646), .A2(n28580), .ZN(n21647) );
  XOR2_X1 U11998 ( .A1(n29652), .A2(n15566), .Z(n27643) );
  XOR2_X1 U12015 ( .A1(n30306), .A2(n22243), .Z(n28835) );
  INV_X2 U12018 ( .I(n26738), .ZN(n17688) );
  XOR2_X1 U12025 ( .A1(n26740), .A2(n17663), .Z(n25115) );
  XOR2_X1 U12026 ( .A1(n24788), .A2(n1226), .Z(n26740) );
  NAND3_X2 U12037 ( .A1(n12876), .A2(n12875), .A3(n1182), .ZN(n26742) );
  NAND2_X1 U12045 ( .A1(n10359), .A2(n25995), .ZN(n26744) );
  NOR2_X1 U12058 ( .A1(n20067), .A2(n13080), .ZN(n27542) );
  OAI21_X1 U12069 ( .A1(n12904), .A2(n24305), .B(n26747), .ZN(n24302) );
  AOI21_X1 U12070 ( .A1(n27430), .A2(n12904), .B(n1241), .ZN(n26747) );
  NAND2_X1 U12081 ( .A1(n867), .A2(n18078), .ZN(n2512) );
  XOR2_X1 U12094 ( .A1(n4955), .A2(n22790), .Z(n14382) );
  INV_X2 U12129 ( .I(n19597), .ZN(n26751) );
  AND2_X1 U12132 ( .A1(n15149), .A2(n21147), .Z(n11151) );
  NAND2_X1 U12142 ( .A1(n3646), .A2(n7929), .ZN(n7926) );
  XOR2_X1 U12147 ( .A1(n26755), .A2(n15904), .Z(n27824) );
  XOR2_X1 U12149 ( .A1(n27825), .A2(n19448), .Z(n26755) );
  NOR2_X2 U12178 ( .A1(n2395), .A2(n7986), .ZN(n2394) );
  INV_X1 U12185 ( .I(n2380), .ZN(n26758) );
  NAND2_X2 U12239 ( .A1(n4909), .A2(n4913), .ZN(n5348) );
  XOR2_X1 U12275 ( .A1(n13145), .A2(n24409), .Z(n27951) );
  NOR2_X1 U12295 ( .A1(n15456), .A2(n12315), .ZN(n12118) );
  INV_X2 U12301 ( .I(n26761), .ZN(n579) );
  XOR2_X1 U12303 ( .A1(n5768), .A2(n503), .Z(n26761) );
  NAND2_X2 U12307 ( .A1(n26762), .A2(n3594), .ZN(n16297) );
  NAND2_X2 U12310 ( .A1(n3597), .A2(n3598), .ZN(n22500) );
  XOR2_X1 U12311 ( .A1(n10631), .A2(n13470), .Z(n13309) );
  XOR2_X1 U12315 ( .A1(n26765), .A2(n22102), .Z(n4161) );
  OAI21_X1 U12322 ( .A1(n2536), .A2(n14940), .B(n25995), .ZN(n5300) );
  NOR2_X2 U12329 ( .A1(n7732), .A2(n11970), .ZN(n13495) );
  NAND2_X2 U12372 ( .A1(n25670), .A2(n25675), .ZN(n25691) );
  OAI22_X2 U12376 ( .A1(n9083), .A2(n17370), .B1(n18993), .B2(n13252), .ZN(
        n26768) );
  XOR2_X1 U12378 ( .A1(n110), .A2(n7025), .Z(n7024) );
  AND2_X1 U12382 ( .A1(n19857), .A2(n20067), .Z(n27541) );
  INV_X1 U12394 ( .I(n28504), .ZN(n15824) );
  OR2_X1 U12395 ( .A1(n28504), .A2(n31967), .Z(n16251) );
  OR2_X1 U12402 ( .A1(n5410), .A2(n25995), .Z(n7425) );
  AND3_X1 U12404 ( .A1(n22505), .A2(n22524), .A3(n8314), .Z(n29026) );
  INV_X2 U12408 ( .I(n23144), .ZN(n23841) );
  NAND2_X2 U12421 ( .A1(n15137), .A2(n30995), .ZN(n18477) );
  INV_X1 U12422 ( .I(n21214), .ZN(n21215) );
  XOR2_X1 U12441 ( .A1(n23241), .A2(n23533), .Z(n9863) );
  AND2_X1 U12450 ( .A1(n8083), .A2(n12231), .Z(n26780) );
  OR2_X1 U12456 ( .A1(n23843), .A2(n31796), .Z(n14350) );
  NOR2_X1 U12475 ( .A1(n4006), .A2(n1109), .ZN(n16927) );
  XOR2_X1 U12492 ( .A1(n9843), .A2(n28927), .Z(n23210) );
  NAND2_X2 U12493 ( .A1(n4542), .A2(n4543), .ZN(n9843) );
  NOR2_X2 U12499 ( .A1(n10373), .A2(n1384), .ZN(n12744) );
  XNOR2_X1 U12510 ( .A1(Key[93]), .A2(Plaintext[93]), .ZN(n26791) );
  OAI21_X2 U12521 ( .A1(n17320), .A2(n15378), .B(n17319), .ZN(n19436) );
  NAND2_X2 U12526 ( .A1(n8286), .A2(n14551), .ZN(n24218) );
  AND2_X1 U12548 ( .A1(n20334), .A2(n28261), .Z(n12089) );
  XNOR2_X1 U12557 ( .A1(n10075), .A2(n22080), .ZN(n26822) );
  NAND2_X2 U12576 ( .A1(n26799), .A2(n16414), .ZN(n22919) );
  INV_X1 U12590 ( .I(n5373), .ZN(n28740) );
  NAND2_X1 U12617 ( .A1(n7040), .A2(n25734), .ZN(n7039) );
  INV_X2 U12620 ( .I(n27105), .ZN(n20541) );
  XOR2_X1 U12625 ( .A1(n15618), .A2(n26807), .Z(n15617) );
  XOR2_X1 U12626 ( .A1(n2477), .A2(n371), .Z(n26807) );
  OAI21_X2 U12630 ( .A1(n28347), .A2(n4177), .B(n25996), .ZN(n26808) );
  NOR2_X1 U12632 ( .A1(n6816), .A2(n25128), .ZN(n27518) );
  INV_X2 U12661 ( .I(n20305), .ZN(n20419) );
  AOI21_X1 U12664 ( .A1(n31821), .A2(n11123), .B(n13279), .ZN(n18303) );
  INV_X2 U12668 ( .I(n26812), .ZN(n13496) );
  XOR2_X1 U12676 ( .A1(n9636), .A2(n26815), .Z(n20102) );
  XOR2_X1 U12705 ( .A1(n5279), .A2(n5280), .Z(n5287) );
  XOR2_X1 U12712 ( .A1(n26821), .A2(n22082), .Z(n10681) );
  XOR2_X1 U12718 ( .A1(n22081), .A2(n26822), .Z(n26821) );
  NOR2_X2 U12730 ( .A1(n24498), .A2(n24499), .ZN(n24750) );
  NAND2_X1 U12732 ( .A1(n13747), .A2(n10805), .ZN(n26825) );
  OAI22_X2 U12745 ( .A1(n31079), .A2(n11637), .B1(n29077), .B2(n8454), .ZN(
        n11634) );
  XOR2_X1 U12750 ( .A1(n23426), .A2(n23427), .Z(n10674) );
  NOR3_X1 U12757 ( .A1(n28704), .A2(n1168), .A3(n17670), .ZN(n26827) );
  XOR2_X1 U12765 ( .A1(n21006), .A2(n6431), .Z(n20748) );
  INV_X2 U12770 ( .I(n19284), .ZN(n28721) );
  NAND2_X2 U12776 ( .A1(n1680), .A2(n1679), .ZN(n20467) );
  XOR2_X1 U12782 ( .A1(n3195), .A2(n19691), .Z(n3652) );
  NAND2_X1 U12796 ( .A1(n16265), .A2(n16266), .ZN(n21104) );
  AOI21_X2 U12800 ( .A1(n14867), .A2(n25123), .B(n16607), .ZN(n14866) );
  NAND2_X2 U12807 ( .A1(n7310), .A2(n13622), .ZN(n22890) );
  OR2_X1 U12810 ( .A1(n9406), .A2(n6908), .Z(n6013) );
  OAI22_X2 U12813 ( .A1(n26078), .A2(n9146), .B1(n24347), .B2(n29043), .ZN(
        n29143) );
  XOR2_X1 U12852 ( .A1(n21896), .A2(n26096), .Z(n26842) );
  XOR2_X1 U12858 ( .A1(n26844), .A2(n12461), .Z(n27004) );
  XOR2_X1 U12861 ( .A1(n22165), .A2(n26845), .Z(n26844) );
  INV_X2 U12872 ( .I(n26846), .ZN(n17971) );
  OAI21_X2 U12877 ( .A1(n11106), .A2(n7656), .B(n26432), .ZN(n1862) );
  NAND2_X2 U12881 ( .A1(n27765), .A2(n21140), .ZN(n21592) );
  XOR2_X1 U12884 ( .A1(n27613), .A2(n26582), .Z(n23514) );
  NAND3_X1 U12910 ( .A1(n33750), .A2(n630), .A3(n26305), .ZN(n21909) );
  AOI22_X2 U12911 ( .A1(n26855), .A2(n1773), .B1(n22375), .B2(n1282), .ZN(
        n9575) );
  OAI21_X1 U12915 ( .A1(n23026), .A2(n26169), .B(n16280), .ZN(n26856) );
  XOR2_X1 U12924 ( .A1(n32861), .A2(n24738), .Z(n23151) );
  INV_X1 U12925 ( .I(n5826), .ZN(n27302) );
  NOR2_X1 U12953 ( .A1(n14102), .A2(n750), .ZN(n14101) );
  XOR2_X1 U12956 ( .A1(n29220), .A2(n7382), .Z(n26865) );
  AOI22_X2 U12961 ( .A1(n19992), .A2(n16681), .B1(n19993), .B2(n19943), .ZN(
        n28786) );
  AOI22_X1 U12963 ( .A1(n25492), .A2(n30047), .B1(n138), .B2(n4183), .ZN(
        n25494) );
  XOR2_X1 U12964 ( .A1(n23417), .A2(n23444), .Z(n23497) );
  OAI21_X2 U12974 ( .A1(n26023), .A2(n28634), .B(n6144), .ZN(n25330) );
  XOR2_X1 U12993 ( .A1(n9269), .A2(n30314), .Z(n27055) );
  XOR2_X1 U13007 ( .A1(n11324), .A2(n26869), .Z(n6502) );
  XOR2_X1 U13009 ( .A1(n23457), .A2(n16402), .Z(n26869) );
  OAI21_X1 U13017 ( .A1(n28166), .A2(n16374), .B(n16218), .ZN(n14876) );
  XOR2_X1 U13036 ( .A1(n9006), .A2(n462), .Z(n26872) );
  NAND3_X2 U13047 ( .A1(n27437), .A2(n29404), .A3(n9055), .ZN(n26875) );
  XOR2_X1 U13050 ( .A1(n26877), .A2(n16479), .Z(Ciphertext[79]) );
  NOR2_X2 U13064 ( .A1(n27683), .A2(n18435), .ZN(n8606) );
  NAND2_X2 U13069 ( .A1(n26885), .A2(n16028), .ZN(n23189) );
  NOR2_X1 U13072 ( .A1(n22808), .A2(n11308), .ZN(n26886) );
  INV_X1 U13074 ( .I(n22809), .ZN(n26887) );
  XOR2_X1 U13137 ( .A1(n10087), .A2(n22046), .Z(n7640) );
  NAND2_X1 U13146 ( .A1(n8544), .A2(n9375), .ZN(n5116) );
  AND2_X1 U13155 ( .A1(n15704), .A2(n28077), .Z(n28613) );
  INV_X2 U13156 ( .I(n26896), .ZN(n29256) );
  XOR2_X1 U13157 ( .A1(n16770), .A2(n11982), .Z(n26896) );
  XOR2_X1 U13169 ( .A1(n9038), .A2(n26897), .Z(n9037) );
  XOR2_X1 U13170 ( .A1(n15877), .A2(n15), .Z(n26897) );
  AND2_X1 U13193 ( .A1(n30506), .A2(n15863), .Z(n27326) );
  NOR3_X2 U13241 ( .A1(n13475), .A2(n17311), .A3(n948), .ZN(n28175) );
  INV_X1 U13250 ( .I(n27561), .ZN(n28913) );
  NAND3_X2 U13251 ( .A1(n258), .A2(n4290), .A3(n8143), .ZN(n9141) );
  NOR2_X1 U13252 ( .A1(n21529), .A2(n21697), .ZN(n26913) );
  NAND2_X1 U13266 ( .A1(n26724), .A2(n758), .ZN(n5481) );
  NAND2_X1 U13274 ( .A1(n6910), .A2(n25394), .ZN(n26917) );
  INV_X1 U13286 ( .I(n22401), .ZN(n4983) );
  NAND2_X1 U13291 ( .A1(n17477), .A2(n10325), .ZN(n10366) );
  NAND2_X2 U13323 ( .A1(n22965), .A2(n14129), .ZN(n22814) );
  XOR2_X1 U13336 ( .A1(n1971), .A2(n859), .Z(n22292) );
  AOI22_X2 U13338 ( .A1(n26921), .A2(n33460), .B1(n25297), .B2(n28763), .ZN(
        n15483) );
  XOR2_X1 U13347 ( .A1(n22193), .A2(n26922), .Z(n17487) );
  XOR2_X1 U13348 ( .A1(n16619), .A2(n30314), .Z(n26922) );
  XOR2_X1 U13350 ( .A1(n6396), .A2(n32154), .Z(n11528) );
  NAND2_X2 U13356 ( .A1(n22615), .A2(n11308), .ZN(n4399) );
  XOR2_X1 U13361 ( .A1(n4660), .A2(n26923), .Z(n666) );
  XOR2_X1 U13362 ( .A1(n26924), .A2(n23249), .Z(n26923) );
  OAI21_X1 U13385 ( .A1(n26051), .A2(n1318), .B(n26927), .ZN(n14674) );
  INV_X2 U13399 ( .I(n26930), .ZN(n13308) );
  INV_X2 U13414 ( .I(n22048), .ZN(n26931) );
  OAI22_X2 U13422 ( .A1(n5694), .A2(n13605), .B1(n11120), .B2(n5693), .ZN(
        n20634) );
  XOR2_X1 U13426 ( .A1(n26934), .A2(n26933), .Z(n27880) );
  XOR2_X1 U13436 ( .A1(n5742), .A2(n26936), .Z(n1708) );
  INV_X1 U13437 ( .I(n16604), .ZN(n26936) );
  NAND2_X2 U13442 ( .A1(n11873), .A2(n14623), .ZN(n5742) );
  XOR2_X1 U13448 ( .A1(n2981), .A2(n26004), .Z(n2978) );
  NOR3_X2 U13449 ( .A1(n34131), .A2(n3236), .A3(n31760), .ZN(n6958) );
  OAI21_X2 U13450 ( .A1(n6101), .A2(n4489), .B(n26937), .ZN(n22870) );
  INV_X2 U13452 ( .I(n9890), .ZN(n26938) );
  AOI22_X2 U13464 ( .A1(n6858), .A2(n6859), .B1(n16681), .B2(n19944), .ZN(
        n8118) );
  XOR2_X1 U13466 ( .A1(n12878), .A2(n17929), .Z(n23245) );
  OAI22_X2 U13469 ( .A1(n6964), .A2(n896), .B1(n13142), .B2(n6965), .ZN(n17929) );
  OAI21_X2 U13487 ( .A1(n14653), .A2(n14654), .B(n13686), .ZN(n27242) );
  AOI21_X2 U13490 ( .A1(n21274), .A2(n21273), .B(n21272), .ZN(n16327) );
  AOI21_X2 U13491 ( .A1(n22892), .A2(n23037), .B(n899), .ZN(n8149) );
  NAND2_X2 U13512 ( .A1(n16663), .A2(n23542), .ZN(n16066) );
  OR2_X1 U13513 ( .A1(n4274), .A2(n27838), .Z(n5684) );
  XOR2_X1 U13517 ( .A1(n15560), .A2(n26941), .Z(n12595) );
  XOR2_X1 U13518 ( .A1(n26942), .A2(n22248), .Z(n26941) );
  NAND2_X2 U13527 ( .A1(n1602), .A2(n18977), .ZN(n15074) );
  XOR2_X1 U13529 ( .A1(n29162), .A2(n26945), .Z(n28373) );
  XOR2_X1 U13536 ( .A1(n17128), .A2(n32024), .Z(n26945) );
  XOR2_X1 U13539 ( .A1(n26947), .A2(n11289), .Z(n29273) );
  XOR2_X1 U13543 ( .A1(n5382), .A2(n26118), .Z(n26947) );
  NAND3_X1 U13546 ( .A1(n25788), .A2(n25796), .A3(n12611), .ZN(n26948) );
  NAND2_X2 U13547 ( .A1(n9323), .A2(n26950), .ZN(n26949) );
  OAI21_X2 U13563 ( .A1(n23722), .A2(n23349), .B(n9443), .ZN(n18077) );
  NOR2_X1 U13565 ( .A1(n2512), .A2(n31873), .ZN(n26953) );
  XOR2_X1 U13575 ( .A1(n2388), .A2(n3727), .Z(n2982) );
  NOR2_X2 U13588 ( .A1(n772), .A2(n31129), .ZN(n4489) );
  XOR2_X1 U13592 ( .A1(n19709), .A2(n19397), .Z(n17953) );
  XOR2_X1 U13595 ( .A1(n22085), .A2(n26957), .Z(n10873) );
  NAND2_X2 U13611 ( .A1(n26958), .A2(n4854), .ZN(n20374) );
  OAI21_X1 U13617 ( .A1(n25556), .A2(n28760), .B(n28759), .ZN(n28758) );
  AOI21_X2 U13619 ( .A1(n30502), .A2(n22706), .B(n26960), .ZN(n13814) );
  XOR2_X1 U13631 ( .A1(n26426), .A2(n32893), .Z(n27548) );
  NAND2_X2 U13644 ( .A1(n25914), .A2(n25913), .ZN(n25923) );
  XOR2_X1 U13651 ( .A1(n23275), .A2(n24623), .Z(n23174) );
  NOR2_X2 U13652 ( .A1(n13289), .A2(n13288), .ZN(n23275) );
  XOR2_X1 U13665 ( .A1(n8893), .A2(n26111), .Z(n8892) );
  NAND2_X2 U13670 ( .A1(n13918), .A2(n11057), .ZN(n27763) );
  XOR2_X1 U13686 ( .A1(n24682), .A2(n13614), .Z(n14897) );
  XOR2_X1 U13689 ( .A1(n20736), .A2(n20953), .Z(n20808) );
  OAI21_X2 U13690 ( .A1(n5879), .A2(n5909), .B(n12194), .ZN(n17947) );
  NOR2_X2 U13695 ( .A1(n27460), .A2(n19014), .ZN(n19699) );
  NAND2_X1 U13697 ( .A1(n12777), .A2(n23912), .ZN(n26967) );
  XOR2_X1 U13698 ( .A1(n9459), .A2(n21993), .Z(n1713) );
  OR2_X1 U13731 ( .A1(n3157), .A2(n30130), .Z(n10613) );
  NOR2_X1 U13740 ( .A1(n9690), .A2(n5074), .ZN(n14589) );
  NAND2_X1 U13741 ( .A1(n15228), .A2(n16098), .ZN(n13971) );
  NAND2_X1 U13746 ( .A1(n13766), .A2(n13765), .ZN(n26974) );
  NAND2_X2 U13752 ( .A1(n7474), .A2(n7473), .ZN(n9025) );
  XOR2_X1 U13756 ( .A1(n14296), .A2(n21023), .Z(n26977) );
  INV_X2 U13761 ( .I(n26978), .ZN(n700) );
  XOR2_X1 U13763 ( .A1(n11171), .A2(n11169), .Z(n26978) );
  NAND2_X1 U13776 ( .A1(n21285), .A2(n29303), .ZN(n27431) );
  INV_X2 U13790 ( .I(n26980), .ZN(n1835) );
  XOR2_X1 U13798 ( .A1(Plaintext[127]), .A2(Key[127]), .Z(n26980) );
  AND2_X1 U13814 ( .A1(n5741), .A2(n24190), .Z(n6770) );
  XOR2_X1 U13828 ( .A1(n26983), .A2(n31912), .Z(n616) );
  XOR2_X1 U13829 ( .A1(n28490), .A2(n13612), .Z(n26983) );
  XOR2_X1 U13830 ( .A1(n28177), .A2(n2458), .Z(n17826) );
  INV_X2 U13853 ( .I(n8040), .ZN(n10360) );
  XOR2_X1 U13872 ( .A1(n589), .A2(n3237), .Z(n6556) );
  XOR2_X1 U13887 ( .A1(n20449), .A2(n20748), .Z(n1613) );
  NOR2_X2 U13892 ( .A1(n11447), .A2(n11446), .ZN(n6500) );
  NAND2_X1 U13899 ( .A1(n24335), .A2(n24242), .ZN(n11563) );
  OAI21_X2 U13902 ( .A1(n26991), .A2(n27889), .B(n904), .ZN(n6836) );
  NAND3_X1 U13903 ( .A1(n1896), .A2(n25717), .A3(n26992), .ZN(n25719) );
  INV_X2 U13905 ( .I(n1102), .ZN(n23393) );
  NOR2_X2 U13909 ( .A1(n26995), .A2(n26994), .ZN(n1102) );
  XOR2_X1 U13914 ( .A1(n20049), .A2(n20050), .Z(n21221) );
  AND2_X1 U13920 ( .A1(n23944), .A2(n16961), .Z(n16676) );
  NAND3_X2 U13928 ( .A1(n7777), .A2(n5776), .A3(n664), .ZN(n9220) );
  XOR2_X1 U13929 ( .A1(n16303), .A2(n19682), .Z(n19486) );
  XOR2_X1 U13934 ( .A1(n19744), .A2(n3568), .Z(n16303) );
  NAND3_X2 U13936 ( .A1(n4212), .A2(n4211), .A3(n17021), .ZN(n26998) );
  NAND2_X2 U13942 ( .A1(n27752), .A2(n29314), .ZN(n14978) );
  OAI21_X2 U13951 ( .A1(n27865), .A2(n22904), .B(n18177), .ZN(n23247) );
  INV_X4 U13957 ( .I(n5073), .ZN(n761) );
  NAND2_X2 U13961 ( .A1(n14627), .A2(n15641), .ZN(n2726) );
  NOR2_X2 U13967 ( .A1(n777), .A2(n32898), .ZN(n11756) );
  NOR2_X2 U13973 ( .A1(n3312), .A2(n10572), .ZN(n21350) );
  NAND2_X2 U13975 ( .A1(n14719), .A2(n2821), .ZN(n20428) );
  NOR2_X2 U13977 ( .A1(n3527), .A2(n3525), .ZN(n2821) );
  XOR2_X1 U13997 ( .A1(n7535), .A2(n28144), .Z(n10770) );
  OAI21_X2 U13998 ( .A1(n27010), .A2(n11187), .B(n21421), .ZN(n14236) );
  XOR2_X1 U14001 ( .A1(n27011), .A2(n721), .Z(n23490) );
  INV_X2 U14004 ( .I(n27012), .ZN(n599) );
  NOR2_X1 U14006 ( .A1(n8270), .A2(n28847), .ZN(n29080) );
  XOR2_X1 U14011 ( .A1(n12924), .A2(n14077), .Z(n12923) );
  XOR2_X1 U14022 ( .A1(n27169), .A2(n27015), .Z(n27014) );
  OR2_X1 U14025 ( .A1(n579), .A2(n29250), .Z(n10484) );
  INV_X4 U14031 ( .I(n9280), .ZN(n5178) );
  XOR2_X1 U14033 ( .A1(n3568), .A2(n14588), .Z(n19726) );
  NAND2_X2 U14035 ( .A1(n25440), .A2(n25441), .ZN(n25429) );
  XOR2_X1 U14040 ( .A1(n21992), .A2(n22013), .Z(n13873) );
  XOR2_X1 U14054 ( .A1(n20907), .A2(n21028), .Z(n3617) );
  NOR2_X2 U14075 ( .A1(n2705), .A2(n2706), .ZN(n8506) );
  XOR2_X1 U14082 ( .A1(n23507), .A2(n27708), .Z(n4413) );
  AND2_X1 U14086 ( .A1(n23968), .A2(n23969), .Z(n27026) );
  NAND4_X1 U14097 ( .A1(n25440), .A2(n25442), .A3(n25439), .A4(n25441), .ZN(
        n25443) );
  NAND2_X2 U14112 ( .A1(n13800), .A2(n14950), .ZN(n6442) );
  NAND2_X2 U14115 ( .A1(n5973), .A2(n22654), .ZN(n23137) );
  OR2_X1 U14125 ( .A1(n25675), .A2(n25686), .Z(n25685) );
  NAND3_X1 U14166 ( .A1(n17087), .A2(n23723), .A3(n23738), .ZN(n28506) );
  XOR2_X1 U14167 ( .A1(n6168), .A2(n24809), .Z(n24405) );
  NAND2_X2 U14169 ( .A1(n6167), .A2(n6166), .ZN(n24809) );
  XOR2_X1 U14170 ( .A1(n27613), .A2(n27126), .Z(n27041) );
  XOR2_X1 U14173 ( .A1(n27190), .A2(n22131), .Z(n22136) );
  XOR2_X1 U14174 ( .A1(n22192), .A2(n22130), .Z(n27190) );
  XOR2_X1 U14181 ( .A1(n3280), .A2(n27042), .Z(n17799) );
  AOI22_X2 U14183 ( .A1(n12886), .A2(n2990), .B1(n16318), .B2(n11323), .ZN(
        n11322) );
  NAND2_X1 U14195 ( .A1(n5327), .A2(n17649), .ZN(n17553) );
  NAND2_X2 U14204 ( .A1(n27044), .A2(n2992), .ZN(n24315) );
  NAND2_X1 U14212 ( .A1(n24168), .A2(n5454), .ZN(n3984) );
  XOR2_X1 U14219 ( .A1(n27047), .A2(n1424), .Z(Ciphertext[80]) );
  AOI22_X2 U14224 ( .A1(n3297), .A2(n28649), .B1(n3296), .B2(n33132), .ZN(
        n1565) );
  INV_X2 U14228 ( .I(n27050), .ZN(n4577) );
  XOR2_X1 U14229 ( .A1(n4578), .A2(n4579), .Z(n27050) );
  XOR2_X1 U14231 ( .A1(n16998), .A2(n23165), .Z(n27052) );
  XOR2_X1 U14232 ( .A1(n24621), .A2(n17325), .Z(n13513) );
  XOR2_X1 U14243 ( .A1(n20815), .A2(n21018), .Z(n27054) );
  XOR2_X1 U14252 ( .A1(n11836), .A2(n23295), .Z(n11822) );
  XOR2_X1 U14253 ( .A1(n23519), .A2(n23294), .Z(n11836) );
  INV_X2 U14283 ( .I(n27058), .ZN(n14083) );
  OR2_X1 U14307 ( .A1(n7425), .A2(n25879), .Z(n7265) );
  XOR2_X1 U14315 ( .A1(n27063), .A2(n25319), .Z(Ciphertext[94]) );
  XOR2_X1 U14318 ( .A1(n19483), .A2(n26002), .Z(n19305) );
  AOI21_X2 U14325 ( .A1(n27066), .A2(n11376), .B(n22280), .ZN(n22785) );
  OAI21_X2 U14329 ( .A1(n8479), .A2(n29115), .B(n27652), .ZN(n27067) );
  XOR2_X1 U14341 ( .A1(n22970), .A2(n30993), .Z(n7011) );
  AOI21_X2 U14344 ( .A1(n15730), .A2(n15729), .B(n14680), .ZN(n22970) );
  XOR2_X1 U14350 ( .A1(n24456), .A2(n24457), .Z(n27072) );
  INV_X2 U14364 ( .I(n7453), .ZN(n21241) );
  NAND2_X2 U14383 ( .A1(n27392), .A2(n29131), .ZN(n24138) );
  XOR2_X1 U14385 ( .A1(n27081), .A2(n27080), .Z(n28151) );
  XOR2_X1 U14387 ( .A1(n8432), .A2(n23243), .Z(n27081) );
  XOR2_X1 U14391 ( .A1(n3491), .A2(n27082), .Z(n416) );
  XOR2_X1 U14392 ( .A1(n33971), .A2(n26701), .Z(n27082) );
  AND2_X1 U14393 ( .A1(n28123), .A2(n15038), .Z(n9734) );
  XOR2_X1 U14414 ( .A1(n6151), .A2(n6152), .Z(n14255) );
  XOR2_X1 U14423 ( .A1(n30193), .A2(n9904), .Z(n19575) );
  XOR2_X1 U14431 ( .A1(n23313), .A2(n17500), .Z(n12950) );
  INV_X1 U14452 ( .I(n22933), .ZN(n27088) );
  XOR2_X1 U14462 ( .A1(n1302), .A2(n22027), .Z(n8680) );
  BUF_X2 U14475 ( .I(n11622), .Z(n6034) );
  XOR2_X1 U14492 ( .A1(n22043), .A2(n10155), .Z(n10154) );
  XOR2_X1 U14494 ( .A1(n22173), .A2(n22196), .Z(n22043) );
  NAND2_X2 U14502 ( .A1(n4167), .A2(n4168), .ZN(n15043) );
  XOR2_X1 U14507 ( .A1(n4448), .A2(n20908), .Z(n27091) );
  OAI22_X1 U14530 ( .A1(n10009), .A2(n10012), .B1(n10385), .B2(n30557), .ZN(
        n27092) );
  NAND2_X2 U14531 ( .A1(n17364), .A2(n14), .ZN(n2843) );
  INV_X2 U14534 ( .I(n1696), .ZN(n8100) );
  XOR2_X1 U14537 ( .A1(n1698), .A2(n29079), .Z(n1696) );
  NOR2_X1 U14539 ( .A1(n14881), .A2(n22522), .ZN(n27094) );
  XNOR2_X1 U14542 ( .A1(n12789), .A2(n21994), .ZN(n22193) );
  AOI21_X1 U14563 ( .A1(n28973), .A2(n28972), .B(n27532), .ZN(n28494) );
  NOR2_X2 U14580 ( .A1(n28455), .A2(n25902), .ZN(n10085) );
  NAND3_X2 U14582 ( .A1(n20290), .A2(n20289), .A3(n20292), .ZN(n14821) );
  AOI21_X2 U14586 ( .A1(n28167), .A2(n28166), .B(n34132), .ZN(n15749) );
  XOR2_X1 U14590 ( .A1(n22311), .A2(n12621), .Z(n8405) );
  XOR2_X1 U14592 ( .A1(Key[47]), .A2(Plaintext[47]), .Z(n28946) );
  XOR2_X1 U14600 ( .A1(n15489), .A2(n15487), .Z(n28765) );
  NOR2_X2 U14607 ( .A1(n19135), .A2(n15126), .ZN(n19654) );
  NAND2_X2 U14619 ( .A1(n4801), .A2(n4804), .ZN(n11193) );
  XOR2_X1 U14629 ( .A1(n24792), .A2(n27100), .Z(n17663) );
  XOR2_X1 U14630 ( .A1(n24790), .A2(n27101), .Z(n27100) );
  INV_X1 U14631 ( .I(n25648), .ZN(n27101) );
  XOR2_X1 U14645 ( .A1(n10172), .A2(n8562), .Z(n10170) );
  XOR2_X1 U14651 ( .A1(n12675), .A2(n24786), .Z(n24817) );
  OAI21_X2 U14653 ( .A1(n9658), .A2(n9659), .B(n23996), .ZN(n24786) );
  XOR2_X1 U14658 ( .A1(n32880), .A2(n25436), .Z(n15923) );
  XOR2_X1 U14662 ( .A1(n24821), .A2(n24822), .Z(n25242) );
  AOI21_X2 U14670 ( .A1(n2726), .A2(n1218), .B(n16276), .ZN(n1547) );
  OAI21_X2 U14678 ( .A1(n7147), .A2(n6427), .B(n8603), .ZN(n8602) );
  NAND2_X1 U14687 ( .A1(n17273), .A2(n7925), .ZN(n5568) );
  OAI22_X2 U14689 ( .A1(n3529), .A2(n27111), .B1(n761), .B2(n2089), .ZN(n3527)
         );
  NOR2_X2 U14697 ( .A1(n4871), .A2(n28449), .ZN(n23430) );
  OR2_X1 U14703 ( .A1(n17239), .A2(n28705), .Z(n12565) );
  INV_X4 U14712 ( .I(n27214), .ZN(n7492) );
  INV_X2 U14721 ( .I(n11934), .ZN(n16397) );
  OAI21_X1 U14726 ( .A1(n25559), .A2(n14944), .B(n28758), .ZN(n15292) );
  NOR3_X1 U14742 ( .A1(n24311), .A2(n7503), .A3(n9962), .ZN(n27982) );
  NAND3_X2 U14746 ( .A1(n24017), .A2(n24016), .A3(n24018), .ZN(n27115) );
  NAND3_X1 U14747 ( .A1(n24017), .A2(n24016), .A3(n24018), .ZN(n24832) );
  INV_X1 U14758 ( .I(n28761), .ZN(n28760) );
  NAND2_X1 U14760 ( .A1(n16092), .A2(n16595), .ZN(n29020) );
  NAND2_X1 U14767 ( .A1(n28244), .A2(n28243), .ZN(n25471) );
  NAND3_X1 U14773 ( .A1(n4183), .A2(n25476), .A3(n25470), .ZN(n28244) );
  NAND2_X1 U14777 ( .A1(n25405), .A2(n25412), .ZN(n28738) );
  NOR2_X1 U14781 ( .A1(n15665), .A2(n8616), .ZN(n29098) );
  NAND2_X1 U14800 ( .A1(n16684), .A2(n20561), .ZN(n19906) );
  AND2_X1 U14809 ( .A1(n8238), .A2(n14195), .Z(n5376) );
  NOR2_X1 U14817 ( .A1(n25302), .A2(n25229), .ZN(n1858) );
  OAI21_X1 U14820 ( .A1(n14959), .A2(n4245), .B(n26020), .ZN(n25017) );
  INV_X1 U14829 ( .I(n23043), .ZN(n28356) );
  OR2_X1 U14834 ( .A1(n16425), .A2(n25570), .Z(n11852) );
  INV_X2 U14835 ( .I(n30783), .ZN(n2088) );
  AND2_X1 U14845 ( .A1(n1218), .A2(n15641), .Z(n25186) );
  NAND2_X1 U14849 ( .A1(n25611), .A2(n25612), .ZN(n10266) );
  INV_X1 U14850 ( .I(n9982), .ZN(n25612) );
  NAND2_X1 U14851 ( .A1(n750), .A2(n25368), .ZN(n15479) );
  NAND3_X1 U14852 ( .A1(n9731), .A2(n9733), .A3(n25323), .ZN(n27330) );
  AOI22_X1 U14855 ( .A1(n25539), .A2(n12088), .B1(n9917), .B2(n15481), .ZN(
        n15480) );
  NAND2_X1 U14856 ( .A1(n14454), .A2(n17382), .ZN(n3033) );
  NOR2_X1 U14865 ( .A1(n27926), .A2(n14454), .ZN(n689) );
  AND2_X1 U14895 ( .A1(n8555), .A2(n4415), .Z(n4416) );
  NOR2_X1 U14896 ( .A1(n17336), .A2(n32092), .ZN(n17335) );
  NAND3_X1 U14907 ( .A1(n25651), .A2(n25666), .A3(n7087), .ZN(n7086) );
  INV_X1 U14918 ( .I(n24181), .ZN(n14111) );
  NOR2_X1 U14919 ( .A1(n25378), .A2(n25369), .ZN(n25360) );
  NOR2_X1 U14949 ( .A1(n27162), .A2(n25858), .ZN(n405) );
  OR2_X1 U14951 ( .A1(n15496), .A2(n25409), .Z(n27119) );
  AND2_X1 U14952 ( .A1(n5343), .A2(n17873), .Z(n27121) );
  NAND2_X1 U14957 ( .A1(n25394), .A2(n25238), .ZN(n15756) );
  INV_X1 U14958 ( .I(n19122), .ZN(n1055) );
  XOR2_X1 U14962 ( .A1(n9623), .A2(n9621), .Z(n27122) );
  NAND2_X1 U14964 ( .A1(n31236), .A2(n25557), .ZN(n28761) );
  OAI22_X1 U14965 ( .A1(n25559), .A2(n25552), .B1(n25544), .B2(n25543), .ZN(
        n16869) );
  INV_X1 U14989 ( .I(n11781), .ZN(n5206) );
  NOR2_X1 U14997 ( .A1(n4041), .A2(n3673), .ZN(n14802) );
  NAND2_X2 U15000 ( .A1(n3724), .A2(n3725), .ZN(n27123) );
  AOI21_X1 U15002 ( .A1(n24996), .A2(n7941), .B(n5113), .ZN(n12035) );
  CLKBUF_X4 U15003 ( .I(n25110), .Z(n8219) );
  AOI21_X1 U15011 ( .A1(n8248), .A2(n7809), .B(n8178), .ZN(n15973) );
  NAND2_X2 U15037 ( .A1(n803), .A2(n29317), .ZN(n22914) );
  NAND3_X1 U15045 ( .A1(n25105), .A2(n787), .A3(n32857), .ZN(n3824) );
  INV_X1 U15046 ( .I(n23403), .ZN(n27552) );
  INV_X1 U15048 ( .I(n25617), .ZN(n25602) );
  OR2_X1 U15062 ( .A1(n8277), .A2(n9920), .Z(n13068) );
  NAND2_X1 U15063 ( .A1(n28904), .A2(n20545), .ZN(n20548) );
  NAND2_X1 U15080 ( .A1(n24780), .A2(n17382), .ZN(n28520) );
  OAI21_X1 U15081 ( .A1(n18648), .A2(n16474), .B(n4200), .ZN(n27561) );
  XNOR2_X1 U15107 ( .A1(Plaintext[77]), .A2(Key[77]), .ZN(n27129) );
  NAND2_X1 U15116 ( .A1(n13037), .A2(n13035), .ZN(n27132) );
  AOI21_X1 U15133 ( .A1(n21306), .A2(n21305), .B(n21303), .ZN(n21101) );
  NAND2_X2 U15144 ( .A1(n9166), .A2(n9167), .ZN(n28350) );
  OR2_X2 U15152 ( .A1(n17378), .A2(n17379), .Z(n27134) );
  NOR2_X1 U15161 ( .A1(n29180), .A2(n33325), .ZN(n13230) );
  NAND2_X2 U15162 ( .A1(n723), .A2(n27719), .ZN(n22897) );
  CLKBUF_X1 U15168 ( .I(n6552), .Z(n5254) );
  AOI21_X1 U15175 ( .A1(n17068), .A2(n24283), .B(n16356), .ZN(n24284) );
  NAND2_X1 U15191 ( .A1(n24436), .A2(n25699), .ZN(n17863) );
  OR2_X1 U15196 ( .A1(n24919), .A2(n15569), .Z(n17480) );
  INV_X1 U15198 ( .I(n24919), .ZN(n1200) );
  XOR2_X1 U15199 ( .A1(n10659), .A2(n11148), .Z(n27136) );
  NAND2_X2 U15201 ( .A1(n12597), .A2(n12596), .ZN(n23332) );
  NAND3_X2 U15204 ( .A1(n2870), .A2(n2868), .A3(n2867), .ZN(n27137) );
  NAND3_X2 U15207 ( .A1(n2870), .A2(n2868), .A3(n2867), .ZN(n27138) );
  INV_X1 U15228 ( .I(n29121), .ZN(n27277) );
  OR2_X2 U15230 ( .A1(n495), .A2(n10891), .Z(n9651) );
  NAND2_X1 U15246 ( .A1(n6068), .A2(n6067), .ZN(n27139) );
  OAI21_X1 U15251 ( .A1(n29222), .A2(n10680), .B(n14339), .ZN(n3475) );
  NAND2_X1 U15253 ( .A1(n10680), .A2(n809), .ZN(n15812) );
  OR2_X2 U15267 ( .A1(n11605), .A2(n4036), .Z(n10578) );
  INV_X1 U15276 ( .I(n19335), .ZN(n9538) );
  AOI21_X1 U15278 ( .A1(n5491), .A2(n19335), .B(n14597), .ZN(n1452) );
  XOR2_X1 U15289 ( .A1(n20740), .A2(n20739), .Z(n27143) );
  NAND2_X1 U15304 ( .A1(n25360), .A2(n25368), .ZN(n28516) );
  XOR2_X1 U15308 ( .A1(Key[92]), .A2(Plaintext[92]), .Z(n27146) );
  NAND3_X2 U15313 ( .A1(n8797), .A2(n10765), .A3(n10764), .ZN(n27147) );
  OR2_X2 U15314 ( .A1(n10000), .A2(n7116), .Z(n10765) );
  INV_X2 U15321 ( .I(n16568), .ZN(n20147) );
  INV_X1 U15326 ( .I(n22940), .ZN(n22938) );
  OR2_X2 U15330 ( .A1(n13862), .A2(n636), .Z(n14231) );
  OAI21_X1 U15335 ( .A1(n7361), .A2(n24327), .B(n24245), .ZN(n5286) );
  INV_X1 U15341 ( .I(n16053), .ZN(n17051) );
  NOR2_X2 U15355 ( .A1(n4665), .A2(n4664), .ZN(n27151) );
  NAND2_X1 U15371 ( .A1(n28801), .A2(n16280), .ZN(n11494) );
  NAND2_X2 U15374 ( .A1(n20364), .A2(n20363), .ZN(n4225) );
  NAND2_X1 U15378 ( .A1(n27188), .A2(n18151), .ZN(n9197) );
  XOR2_X1 U15389 ( .A1(n2366), .A2(n2364), .Z(n27154) );
  NAND2_X1 U15394 ( .A1(n16008), .A2(n19156), .ZN(n28372) );
  XOR2_X1 U15398 ( .A1(n15982), .A2(n27155), .Z(n265) );
  XNOR2_X1 U15399 ( .A1(n27115), .A2(n32981), .ZN(n27155) );
  AOI21_X1 U15402 ( .A1(n14813), .A2(n15437), .B(n7188), .ZN(n28403) );
  NAND2_X1 U15403 ( .A1(n32898), .A2(n28099), .ZN(n3043) );
  NAND2_X1 U15404 ( .A1(n27127), .A2(n33681), .ZN(n1890) );
  BUF_X4 U15411 ( .I(n20054), .Z(n8616) );
  OAI21_X1 U15424 ( .A1(n19051), .A2(n19000), .B(n27877), .ZN(n27156) );
  INV_X2 U15435 ( .I(n8721), .ZN(n22599) );
  INV_X2 U15437 ( .I(n25145), .ZN(n17595) );
  OAI21_X1 U15442 ( .A1(n15376), .A2(n888), .B(n33544), .ZN(n15375) );
  NOR3_X1 U15443 ( .A1(n12304), .A2(n25072), .A3(n25078), .ZN(n27925) );
  AND2_X2 U15449 ( .A1(n11063), .A2(n11272), .Z(n15506) );
  INV_X2 U15453 ( .I(n33117), .ZN(n741) );
  OR3_X2 U15460 ( .A1(n1052), .A2(n26600), .A3(n7251), .Z(n18123) );
  NOR2_X1 U15466 ( .A1(n4405), .A2(n1379), .ZN(n3243) );
  INV_X2 U15467 ( .I(n4405), .ZN(n7415) );
  OAI21_X1 U15484 ( .A1(n19058), .A2(n7345), .B(n5625), .ZN(n4914) );
  INV_X1 U15501 ( .I(n25789), .ZN(n29168) );
  NOR2_X1 U15507 ( .A1(n24969), .A2(n3843), .ZN(n2129) );
  NOR2_X1 U15523 ( .A1(n25221), .A2(n7515), .ZN(n10941) );
  CLKBUF_X4 U15526 ( .I(n16045), .Z(n28898) );
  NAND2_X1 U15545 ( .A1(n20401), .A2(n20569), .ZN(n27904) );
  NAND2_X1 U15546 ( .A1(n6765), .A2(n21876), .ZN(n27706) );
  OR2_X1 U15571 ( .A1(n4019), .A2(n24148), .Z(n8963) );
  NOR2_X1 U15579 ( .A1(n11571), .A2(n7929), .ZN(n25253) );
  INV_X2 U15580 ( .I(n6402), .ZN(n1075) );
  OR2_X1 U15591 ( .A1(n22781), .A2(n11383), .Z(n11382) );
  AOI21_X1 U15600 ( .A1(n28659), .A2(n28697), .B(n8040), .ZN(n8038) );
  XOR2_X1 U15627 ( .A1(n11349), .A2(n7717), .Z(n27165) );
  AND2_X2 U15628 ( .A1(n28083), .A2(n4221), .Z(n27166) );
  NAND3_X1 U15676 ( .A1(n6997), .A2(n6995), .A3(n6994), .ZN(n5415) );
  NAND2_X1 U15683 ( .A1(n6431), .A2(n20755), .ZN(n7951) );
  INV_X1 U15692 ( .I(n7093), .ZN(n28715) );
  NAND2_X1 U15701 ( .A1(n20045), .A2(n19907), .ZN(n4143) );
  NAND2_X2 U15706 ( .A1(n10486), .A2(n10489), .ZN(n27169) );
  XOR2_X1 U15709 ( .A1(n3819), .A2(n12672), .Z(n27170) );
  OAI21_X1 U15713 ( .A1(n5274), .A2(n22919), .B(n32967), .ZN(n11539) );
  NAND2_X1 U15726 ( .A1(n6555), .A2(n29043), .ZN(n15437) );
  AND2_X1 U15729 ( .A1(n19724), .A2(n14082), .Z(n19902) );
  NAND3_X2 U15735 ( .A1(n60), .A2(n22943), .A3(n22942), .ZN(n27171) );
  NOR2_X1 U15737 ( .A1(n24164), .A2(n2826), .ZN(n27525) );
  NOR2_X1 U15739 ( .A1(n19249), .A2(n7810), .ZN(n14332) );
  INV_X1 U15751 ( .I(n31394), .ZN(n23442) );
  OAI22_X1 U15755 ( .A1(n27719), .A2(n17211), .B1(n31325), .B2(n723), .ZN(
        n3826) );
  NOR2_X1 U15763 ( .A1(n23066), .A2(n23065), .ZN(n10643) );
  INV_X1 U15774 ( .I(n23066), .ZN(n1281) );
  INV_X2 U15779 ( .I(n12446), .ZN(n12445) );
  INV_X2 U15781 ( .I(n14029), .ZN(n4041) );
  NOR3_X1 U15783 ( .A1(n7232), .A2(n7776), .A3(n7775), .ZN(n27177) );
  AOI21_X2 U15802 ( .A1(n5055), .A2(n5619), .B(n5054), .ZN(n27179) );
  NAND2_X2 U15803 ( .A1(n21537), .A2(n8196), .ZN(n27180) );
  NAND3_X1 U15817 ( .A1(n25199), .A2(n32873), .A3(n9294), .ZN(n7854) );
  INV_X2 U15818 ( .I(n32877), .ZN(n15068) );
  NOR2_X1 U15828 ( .A1(n12482), .A2(n17928), .ZN(n152) );
  NAND2_X1 U15829 ( .A1(n1161), .A2(n9759), .ZN(n20014) );
  XOR2_X1 U15833 ( .A1(n8747), .A2(n8745), .Z(n27181) );
  NAND2_X2 U15839 ( .A1(n27811), .A2(n4800), .ZN(n27184) );
  INV_X1 U15855 ( .I(n25973), .ZN(n12520) );
  OR2_X2 U15864 ( .A1(n16778), .A2(n24565), .Z(n25296) );
  OAI21_X1 U15867 ( .A1(n1071), .A2(n27123), .B(n9247), .ZN(n11365) );
  NAND2_X1 U15869 ( .A1(n27650), .A2(n24883), .ZN(n27461) );
  NAND2_X1 U15899 ( .A1(n10038), .A2(n32876), .ZN(n37) );
  AOI21_X1 U15902 ( .A1(n742), .A2(n741), .B(n31961), .ZN(n20161) );
  OR2_X1 U15905 ( .A1(n31939), .A2(n25700), .Z(n9805) );
  XNOR2_X1 U15906 ( .A1(n7984), .A2(n28746), .ZN(n27188) );
  NAND3_X2 U15914 ( .A1(n8194), .A2(n8195), .A3(n12314), .ZN(n1600) );
  AOI21_X1 U15916 ( .A1(n7287), .A2(n23057), .B(n3007), .ZN(n2911) );
  NAND3_X2 U15918 ( .A1(n26231), .A2(n31437), .A3(n28974), .ZN(n8308) );
  AND2_X2 U15923 ( .A1(n7043), .A2(n31939), .Z(n7064) );
  INV_X1 U15933 ( .I(n18777), .ZN(n954) );
  INV_X1 U15937 ( .I(n14899), .ZN(n5980) );
  INV_X2 U15951 ( .I(n25023), .ZN(n2092) );
  XOR2_X1 U15952 ( .A1(n8939), .A2(n28663), .Z(n25023) );
  MUX2_X1 U15954 ( .I0(n33115), .I1(n22795), .S(n13473), .Z(n6964) );
  OAI21_X2 U15975 ( .A1(n11091), .A2(n12743), .B(n15015), .ZN(n7146) );
  NOR2_X2 U15988 ( .A1(n16165), .A2(n21662), .ZN(n3379) );
  AOI21_X1 U15991 ( .A1(n17595), .A2(n675), .B(n25185), .ZN(n17594) );
  INV_X2 U15992 ( .I(n27202), .ZN(n2499) );
  XOR2_X1 U15993 ( .A1(n2500), .A2(n2501), .Z(n27202) );
  INV_X2 U15995 ( .I(n27203), .ZN(n16792) );
  XOR2_X1 U15996 ( .A1(n19651), .A2(n19384), .Z(n27203) );
  OAI21_X2 U16006 ( .A1(n27402), .A2(n22547), .B(n22393), .ZN(n22375) );
  AOI21_X1 U16017 ( .A1(n25854), .A2(n14199), .B(n10897), .ZN(n25848) );
  NAND3_X1 U16033 ( .A1(n25781), .A2(n16111), .A3(n32874), .ZN(n25769) );
  NOR2_X1 U16043 ( .A1(n10031), .A2(n15704), .ZN(n27212) );
  NOR2_X2 U16056 ( .A1(n7493), .A2(n27215), .ZN(n27214) );
  NAND2_X2 U16063 ( .A1(n27218), .A2(n11291), .ZN(n196) );
  XOR2_X1 U16064 ( .A1(n14250), .A2(n681), .Z(n8562) );
  XOR2_X1 U16069 ( .A1(n24617), .A2(n24421), .Z(n14250) );
  XOR2_X1 U16078 ( .A1(n27220), .A2(n17871), .Z(n23319) );
  XOR2_X1 U16102 ( .A1(n14796), .A2(n518), .Z(n3812) );
  XOR2_X1 U16118 ( .A1(n1902), .A2(n26031), .Z(n27226) );
  BUF_X2 U16119 ( .I(n15455), .Z(n27228) );
  NOR2_X2 U16139 ( .A1(n24064), .A2(n16425), .ZN(n24770) );
  XOR2_X1 U16143 ( .A1(n27234), .A2(n23024), .Z(n23746) );
  OR2_X2 U16147 ( .A1(n9125), .A2(n27894), .Z(n11752) );
  BUF_X2 U16148 ( .I(n16704), .Z(n27236) );
  OAI21_X2 U16161 ( .A1(n26035), .A2(n27238), .B(n27237), .ZN(n2080) );
  AND2_X1 U16169 ( .A1(n6149), .A2(n31637), .Z(n27590) );
  XOR2_X1 U16172 ( .A1(n24372), .A2(n15982), .Z(n28916) );
  AOI21_X1 U16178 ( .A1(n1299), .A2(n16647), .B(n857), .ZN(n6064) );
  INV_X2 U16190 ( .I(n27244), .ZN(n9234) );
  XOR2_X1 U16196 ( .A1(n9235), .A2(n9679), .Z(n27244) );
  AND2_X1 U16210 ( .A1(n19315), .A2(n7197), .Z(n28025) );
  NAND2_X1 U16220 ( .A1(n11135), .A2(n15054), .ZN(n11134) );
  NAND2_X2 U16249 ( .A1(n18408), .A2(n27253), .ZN(n13037) );
  NOR2_X1 U16252 ( .A1(n17605), .A2(n27719), .ZN(n17604) );
  AOI21_X1 U16254 ( .A1(n21859), .A2(n21858), .B(n21860), .ZN(n18251) );
  INV_X2 U16255 ( .I(n27257), .ZN(n11734) );
  NAND2_X1 U16268 ( .A1(n5219), .A2(n27605), .ZN(n5218) );
  NAND2_X1 U16270 ( .A1(n17191), .A2(n26072), .ZN(n13462) );
  NAND2_X2 U16274 ( .A1(n15693), .A2(n15151), .ZN(n7810) );
  NAND2_X2 U16282 ( .A1(n27261), .A2(n18748), .ZN(n19258) );
  XOR2_X1 U16286 ( .A1(n10515), .A2(n15472), .Z(n17523) );
  XOR2_X1 U16300 ( .A1(n29415), .A2(n22042), .Z(n27268) );
  NAND2_X1 U16313 ( .A1(n17637), .A2(n1204), .ZN(n17636) );
  XOR2_X1 U16317 ( .A1(n9087), .A2(n8844), .Z(n8843) );
  NAND2_X2 U16321 ( .A1(n27271), .A2(n13422), .ZN(n5942) );
  NAND2_X1 U16328 ( .A1(n13421), .A2(n25588), .ZN(n27271) );
  NAND2_X2 U16335 ( .A1(n14425), .A2(n14423), .ZN(n29130) );
  XOR2_X1 U16339 ( .A1(n10815), .A2(n10814), .Z(n10813) );
  XOR2_X1 U16342 ( .A1(n19468), .A2(n27275), .Z(n471) );
  XOR2_X1 U16349 ( .A1(n28107), .A2(n27276), .Z(n5640) );
  XOR2_X1 U16352 ( .A1(n5847), .A2(n27277), .Z(n27276) );
  NAND2_X1 U16361 ( .A1(n27282), .A2(n27281), .ZN(n7213) );
  INV_X1 U16362 ( .I(n24991), .ZN(n27281) );
  XOR2_X1 U16364 ( .A1(n28797), .A2(n1225), .Z(n27283) );
  OAI22_X2 U16369 ( .A1(n32095), .A2(n24304), .B1(n16039), .B2(n27284), .ZN(
        n283) );
  OR2_X1 U16373 ( .A1(n18145), .A2(n319), .Z(n27284) );
  XOR2_X1 U16387 ( .A1(n7131), .A2(n23516), .Z(n27289) );
  NAND2_X2 U16392 ( .A1(n15665), .A2(n8616), .ZN(n17675) );
  NOR2_X2 U16393 ( .A1(n19909), .A2(n870), .ZN(n16132) );
  NOR2_X2 U16397 ( .A1(n23560), .A2(n23561), .ZN(n16305) );
  NAND2_X1 U16407 ( .A1(n10435), .A2(n871), .ZN(n10439) );
  NAND2_X2 U16427 ( .A1(n27297), .A2(n21202), .ZN(n5944) );
  NAND2_X2 U16432 ( .A1(n7830), .A2(n21401), .ZN(n27297) );
  OAI22_X2 U16437 ( .A1(n1359), .A2(n20010), .B1(n16664), .B2(n12100), .ZN(
        n3366) );
  AOI22_X2 U16439 ( .A1(n12432), .A2(n28222), .B1(n23646), .B2(n23726), .ZN(
        n27551) );
  NOR2_X1 U16458 ( .A1(n18801), .A2(n32034), .ZN(n4474) );
  INV_X2 U16462 ( .I(n17937), .ZN(n18801) );
  XOR2_X1 U16469 ( .A1(Plaintext[52]), .A2(Key[52]), .Z(n17937) );
  NAND2_X2 U16471 ( .A1(n28789), .A2(n14234), .ZN(n28616) );
  NAND2_X2 U16482 ( .A1(n27302), .A2(n27300), .ZN(n20339) );
  NAND2_X2 U16485 ( .A1(n5906), .A2(n21226), .ZN(n2386) );
  XOR2_X1 U16498 ( .A1(n29140), .A2(n8531), .Z(n6689) );
  XOR2_X1 U16508 ( .A1(n32809), .A2(n19716), .Z(n8283) );
  XOR2_X1 U16509 ( .A1(n19780), .A2(n8785), .Z(n19716) );
  XOR2_X1 U16513 ( .A1(n27308), .A2(n16696), .Z(Ciphertext[133]) );
  OAI21_X1 U16523 ( .A1(n27309), .A2(n24129), .B(n24346), .ZN(n3334) );
  INV_X2 U16529 ( .I(n27311), .ZN(n6416) );
  XNOR2_X1 U16532 ( .A1(Plaintext[176]), .A2(Key[176]), .ZN(n27311) );
  XOR2_X1 U16533 ( .A1(n27312), .A2(n22176), .Z(n22363) );
  INV_X1 U16553 ( .I(n1533), .ZN(n12041) );
  INV_X2 U16554 ( .I(n27315), .ZN(n29116) );
  INV_X2 U16558 ( .I(n25473), .ZN(n27315) );
  NAND2_X1 U16568 ( .A1(n23853), .A2(n23852), .ZN(n27320) );
  NOR2_X2 U16582 ( .A1(n27334), .A2(n27662), .ZN(n27660) );
  INV_X2 U16587 ( .I(n27324), .ZN(n3601) );
  XOR2_X1 U16591 ( .A1(Plaintext[27]), .A2(Key[27]), .Z(n27324) );
  OAI22_X1 U16592 ( .A1(n14564), .A2(n20630), .B1(n9062), .B2(n31471), .ZN(
        n20216) );
  NOR2_X1 U16607 ( .A1(n10217), .A2(n14080), .ZN(n12528) );
  XOR2_X1 U16615 ( .A1(n27330), .A2(n25324), .Z(Ciphertext[95]) );
  NAND2_X1 U16627 ( .A1(n27332), .A2(n25977), .ZN(n3225) );
  AND2_X2 U16630 ( .A1(n24257), .A2(n4746), .Z(n24232) );
  NOR3_X2 U16639 ( .A1(n18805), .A2(n18349), .A3(n16122), .ZN(n18374) );
  AOI21_X2 U16688 ( .A1(n23669), .A2(n1250), .B(n23953), .ZN(n16842) );
  NAND2_X2 U16689 ( .A1(n27731), .A2(n25021), .ZN(n25057) );
  OAI21_X2 U16702 ( .A1(n4422), .A2(n21367), .B(n16311), .ZN(n27337) );
  XOR2_X1 U16725 ( .A1(n14613), .A2(n17914), .Z(n17913) );
  XOR2_X1 U16752 ( .A1(n4562), .A2(n4563), .Z(n7022) );
  NAND3_X2 U16758 ( .A1(n28672), .A2(n28670), .A3(n23651), .ZN(n27341) );
  NAND2_X2 U16769 ( .A1(n14890), .A2(n14888), .ZN(n24790) );
  OR2_X1 U16773 ( .A1(n33684), .A2(n21259), .Z(n28256) );
  XOR2_X1 U16777 ( .A1(n16002), .A2(n2452), .Z(n27344) );
  XOR2_X1 U16793 ( .A1(n6560), .A2(n6562), .Z(n7738) );
  XNOR2_X1 U16794 ( .A1(n28493), .A2(n28492), .ZN(n27881) );
  NOR2_X2 U16821 ( .A1(n24572), .A2(n24570), .ZN(n12431) );
  NAND2_X2 U16824 ( .A1(n16398), .A2(n16400), .ZN(n24572) );
  INV_X1 U16825 ( .I(n4551), .ZN(n27769) );
  OAI21_X1 U16828 ( .A1(n11852), .A2(n24064), .B(n27354), .ZN(n9585) );
  XOR2_X1 U16839 ( .A1(n20985), .A2(n15275), .Z(n15668) );
  XOR2_X1 U16877 ( .A1(n19734), .A2(n10810), .Z(n7297) );
  XOR2_X1 U16878 ( .A1(n19473), .A2(n13106), .Z(n19734) );
  NAND2_X1 U16887 ( .A1(n9663), .A2(n8243), .ZN(n27358) );
  NAND2_X2 U16890 ( .A1(n20441), .A2(n2650), .ZN(n20917) );
  INV_X2 U16898 ( .I(n10835), .ZN(n18059) );
  XOR2_X1 U16900 ( .A1(n5529), .A2(n5530), .Z(n10835) );
  XOR2_X1 U16904 ( .A1(n10766), .A2(n31526), .Z(n27361) );
  AND2_X1 U16919 ( .A1(n23084), .A2(n23088), .Z(n14192) );
  AND2_X1 U16920 ( .A1(n667), .A2(n23843), .Z(n13263) );
  NAND2_X2 U16921 ( .A1(n27363), .A2(n20436), .ZN(n3539) );
  XOR2_X1 U16929 ( .A1(n16303), .A2(n19565), .Z(n16302) );
  XOR2_X1 U16935 ( .A1(n2750), .A2(n26016), .Z(n27365) );
  AND2_X1 U16945 ( .A1(n22955), .A2(n5035), .Z(n22508) );
  NAND2_X1 U16962 ( .A1(n25375), .A2(n25376), .ZN(n4089) );
  XOR2_X1 U16977 ( .A1(n28632), .A2(n21925), .Z(n9267) );
  XOR2_X1 U16993 ( .A1(n11143), .A2(n11144), .Z(n11559) );
  XOR2_X1 U17026 ( .A1(n3868), .A2(n2221), .Z(n2367) );
  OAI21_X2 U17041 ( .A1(n3604), .A2(n3603), .B(n27381), .ZN(n4665) );
  XNOR2_X1 U17042 ( .A1(n1044), .A2(n8785), .ZN(n28458) );
  NAND2_X1 U17050 ( .A1(n22627), .A2(n22628), .ZN(n22629) );
  NAND2_X2 U17053 ( .A1(n2283), .A2(n11302), .ZN(n19038) );
  OR2_X1 U17064 ( .A1(n16868), .A2(n24257), .Z(n9889) );
  INV_X4 U17072 ( .I(n29196), .ZN(n10773) );
  XOR2_X1 U17079 ( .A1(n23246), .A2(n27388), .Z(n8069) );
  XOR2_X1 U17083 ( .A1(n5904), .A2(n13638), .Z(n27388) );
  AOI22_X2 U17088 ( .A1(n15017), .A2(n976), .B1(n9734), .B2(n1249), .ZN(n27392) );
  NOR2_X1 U17108 ( .A1(n15189), .A2(n11959), .ZN(n27398) );
  INV_X2 U17130 ( .I(n27401), .ZN(n2019) );
  XOR2_X1 U17131 ( .A1(Plaintext[149]), .A2(Key[149]), .Z(n27401) );
  NAND2_X2 U17136 ( .A1(n27403), .A2(n18591), .ZN(n8802) );
  AOI22_X2 U17139 ( .A1(n1710), .A2(n11459), .B1(n1709), .B2(n14658), .ZN(
        n27403) );
  NAND2_X1 U17146 ( .A1(n27408), .A2(n32898), .ZN(n9601) );
  NAND2_X1 U17149 ( .A1(n21662), .A2(n4097), .ZN(n27408) );
  AOI22_X2 U17178 ( .A1(n18875), .A2(n10182), .B1(n1709), .B2(n18590), .ZN(
        n18591) );
  NOR2_X2 U17190 ( .A1(n28124), .A2(n17302), .ZN(n12929) );
  XOR2_X1 U17199 ( .A1(n8055), .A2(n29515), .Z(n8054) );
  XOR2_X1 U17234 ( .A1(Plaintext[112]), .A2(Key[112]), .Z(n27428) );
  OAI22_X2 U17247 ( .A1(n2099), .A2(n18447), .B1(n18446), .B2(n18796), .ZN(
        n19268) );
  XOR2_X1 U17259 ( .A1(n23391), .A2(n16622), .Z(n11835) );
  NAND2_X1 U17262 ( .A1(n18844), .A2(n27747), .ZN(n4925) );
  INV_X2 U17273 ( .I(n27435), .ZN(n692) );
  NAND2_X2 U17278 ( .A1(n8081), .A2(n6519), .ZN(n23420) );
  NAND2_X2 U17295 ( .A1(n6068), .A2(n6067), .ZN(n20615) );
  INV_X2 U17301 ( .I(n27441), .ZN(n13413) );
  OAI21_X1 U17302 ( .A1(n16176), .A2(n27442), .B(n782), .ZN(n2771) );
  XOR2_X1 U17312 ( .A1(n14337), .A2(n25428), .Z(n27444) );
  INV_X2 U17321 ( .I(n27453), .ZN(n3933) );
  AOI22_X1 U17322 ( .A1(n15939), .A2(n12530), .B1(n14034), .B2(n22333), .ZN(
        n14750) );
  XOR2_X1 U17324 ( .A1(n4732), .A2(n18122), .Z(n11427) );
  NOR2_X1 U17326 ( .A1(n27456), .A2(n11201), .ZN(n5002) );
  NAND2_X1 U17328 ( .A1(n4999), .A2(n33425), .ZN(n27456) );
  INV_X2 U17344 ( .I(n14577), .ZN(n17078) );
  NAND2_X2 U17348 ( .A1(n3924), .A2(n21067), .ZN(n14577) );
  NOR2_X2 U17351 ( .A1(n12341), .A2(n3380), .ZN(n24682) );
  NAND2_X2 U17374 ( .A1(n13390), .A2(n19355), .ZN(n19280) );
  AND2_X1 U17380 ( .A1(n28865), .A2(n22330), .Z(n28456) );
  INV_X2 U17390 ( .I(n27471), .ZN(n628) );
  XOR2_X1 U17391 ( .A1(n3102), .A2(n3100), .Z(n27471) );
  INV_X2 U17419 ( .I(n27475), .ZN(n10059) );
  XOR2_X1 U17420 ( .A1(n10060), .A2(n11488), .Z(n27475) );
  INV_X4 U17444 ( .I(n29658), .ZN(n28010) );
  XOR2_X1 U17448 ( .A1(n10235), .A2(n10237), .Z(n10236) );
  NAND2_X1 U17473 ( .A1(n8336), .A2(n32862), .ZN(n27480) );
  NOR2_X1 U17482 ( .A1(n21170), .A2(n6957), .ZN(n27482) );
  XOR2_X1 U17484 ( .A1(n24616), .A2(n11722), .Z(n15982) );
  NOR2_X2 U17485 ( .A1(n11723), .A2(n11767), .ZN(n24616) );
  INV_X2 U17497 ( .I(n27485), .ZN(n9430) );
  XOR2_X1 U17515 ( .A1(n27487), .A2(n16390), .Z(Ciphertext[101]) );
  INV_X2 U17520 ( .I(n27490), .ZN(n25339) );
  INV_X2 U17525 ( .I(n31468), .ZN(n27491) );
  AOI21_X2 U17529 ( .A1(n2878), .A2(n1610), .B(n17396), .ZN(n23967) );
  AND3_X1 U17537 ( .A1(n15699), .A2(n29903), .A3(n32080), .Z(n27993) );
  NAND2_X2 U17541 ( .A1(n25999), .A2(n27033), .ZN(n18753) );
  XOR2_X1 U17543 ( .A1(n2331), .A2(n8456), .Z(n10810) );
  XOR2_X1 U17550 ( .A1(n9866), .A2(n9865), .Z(n23696) );
  XOR2_X1 U17583 ( .A1(n27505), .A2(n16636), .Z(Ciphertext[28]) );
  OAI22_X1 U17587 ( .A1(n14318), .A2(n12035), .B1(n14320), .B2(n14322), .ZN(
        n27505) );
  OR2_X1 U17603 ( .A1(n23855), .A2(n9152), .Z(n23690) );
  INV_X2 U17616 ( .I(n27147), .ZN(n20857) );
  OAI21_X2 U17618 ( .A1(n18472), .A2(n18471), .B(n13846), .ZN(n15148) );
  NAND2_X1 U17621 ( .A1(n29376), .A2(n24069), .ZN(n27735) );
  NAND2_X1 U17625 ( .A1(n19053), .A2(n2581), .ZN(n29102) );
  OAI22_X2 U17634 ( .A1(n18622), .A2(n18331), .B1(n18330), .B2(n18329), .ZN(
        n19053) );
  OAI21_X2 U17635 ( .A1(n23798), .A2(n23570), .B(n23797), .ZN(n23571) );
  NOR2_X2 U17636 ( .A1(n13963), .A2(n27509), .ZN(n19222) );
  XNOR2_X1 U17657 ( .A1(n19673), .A2(n11627), .ZN(n29032) );
  XOR2_X1 U17679 ( .A1(n24603), .A2(n24647), .Z(n27516) );
  NAND2_X2 U17680 ( .A1(n2929), .A2(n27517), .ZN(n2928) );
  XNOR2_X1 U17689 ( .A1(n32052), .A2(n20842), .ZN(n20919) );
  INV_X2 U17696 ( .I(n7576), .ZN(n27520) );
  NAND2_X2 U17697 ( .A1(n10198), .A2(n16535), .ZN(n7576) );
  NAND2_X1 U17700 ( .A1(n21568), .A2(n3203), .ZN(n21542) );
  NAND2_X1 U17716 ( .A1(n27525), .A2(n7093), .ZN(n7095) );
  INV_X2 U17730 ( .I(n14794), .ZN(n27529) );
  XOR2_X1 U17735 ( .A1(n24764), .A2(n13060), .Z(n24687) );
  AND2_X1 U17742 ( .A1(n25443), .A2(n25444), .Z(n27531) );
  NOR2_X1 U17751 ( .A1(n14912), .A2(n24141), .ZN(n27534) );
  NAND2_X2 U17756 ( .A1(n28944), .A2(n2680), .ZN(n19289) );
  AND2_X1 U17760 ( .A1(n7195), .A2(n30813), .Z(n15632) );
  NOR2_X1 U17771 ( .A1(n31894), .A2(n985), .ZN(n5177) );
  XOR2_X1 U17785 ( .A1(n27538), .A2(n2473), .Z(n17829) );
  XOR2_X1 U17788 ( .A1(n2476), .A2(n28513), .Z(n27538) );
  XOR2_X1 U17814 ( .A1(n9468), .A2(n24622), .Z(n24768) );
  XOR2_X1 U17826 ( .A1(n28940), .A2(n9387), .Z(n622) );
  NAND2_X2 U17853 ( .A1(n25739), .A2(n1597), .ZN(n1979) );
  AOI21_X2 U17855 ( .A1(n12989), .A2(n17557), .B(n17649), .ZN(n5052) );
  XOR2_X1 U17892 ( .A1(n5149), .A2(n5148), .Z(n5151) );
  XOR2_X1 U17893 ( .A1(n19461), .A2(n17430), .Z(n5149) );
  INV_X4 U17894 ( .I(n25116), .ZN(n27651) );
  NOR2_X1 U17897 ( .A1(n502), .A2(n5433), .ZN(n6954) );
  AOI22_X2 U17898 ( .A1(n28105), .A2(n28104), .B1(n9648), .B2(n7415), .ZN(
        n27553) );
  OAI22_X1 U17909 ( .A1(n10364), .A2(n18884), .B1(n18677), .B2(n17477), .ZN(
        n4659) );
  XOR2_X1 U17931 ( .A1(n5284), .A2(n10111), .Z(n24803) );
  INV_X2 U17948 ( .I(n27563), .ZN(n21505) );
  NOR2_X2 U17950 ( .A1(n21265), .A2(n28375), .ZN(n27563) );
  NAND2_X2 U17976 ( .A1(n7942), .A2(n7943), .ZN(n27566) );
  AOI21_X1 U18012 ( .A1(n13200), .A2(n19178), .B(n19181), .ZN(n8906) );
  OR2_X1 U18026 ( .A1(n24149), .A2(n32178), .Z(n10446) );
  INV_X2 U18027 ( .I(n27570), .ZN(n11821) );
  OAI21_X2 U18035 ( .A1(n6511), .A2(n5119), .B(n17445), .ZN(n18912) );
  XOR2_X1 U18036 ( .A1(n27571), .A2(n18269), .Z(n15721) );
  XOR2_X1 U18052 ( .A1(n27573), .A2(n29241), .Z(n6079) );
  OAI21_X2 U18088 ( .A1(n18749), .A2(n17073), .B(n27582), .ZN(n13160) );
  XNOR2_X1 U18114 ( .A1(n22102), .A2(n25641), .ZN(n27943) );
  XOR2_X1 U18119 ( .A1(n28977), .A2(n26001), .Z(n460) );
  XOR2_X1 U18127 ( .A1(n19630), .A2(n4157), .Z(n14817) );
  OAI21_X2 U18130 ( .A1(n15629), .A2(n15842), .B(n15627), .ZN(n4157) );
  OAI21_X2 U18131 ( .A1(n16318), .A2(n10579), .B(n3179), .ZN(n12886) );
  OR2_X2 U18172 ( .A1(n29334), .A2(n15318), .Z(n15051) );
  XOR2_X1 U18175 ( .A1(n4287), .A2(n24810), .Z(n29236) );
  OAI21_X2 U18181 ( .A1(n27590), .A2(n27589), .B(n27588), .ZN(n13276) );
  INV_X4 U18183 ( .I(n33382), .ZN(n27589) );
  NOR2_X2 U18185 ( .A1(n31973), .A2(n8831), .ZN(n8829) );
  NOR2_X1 U18196 ( .A1(n5741), .A2(n24193), .ZN(n27591) );
  XOR2_X1 U18198 ( .A1(n27593), .A2(n9459), .Z(n13833) );
  XOR2_X1 U18199 ( .A1(n14237), .A2(n3030), .Z(n27593) );
  NOR2_X2 U18200 ( .A1(n10833), .A2(n16359), .ZN(n16357) );
  NOR3_X2 U18201 ( .A1(n32041), .A2(n24273), .A3(n13040), .ZN(n24499) );
  AND2_X2 U18206 ( .A1(n13960), .A2(n7702), .Z(n690) );
  NAND2_X1 U18210 ( .A1(n21663), .A2(n13828), .ZN(n27594) );
  XOR2_X1 U18218 ( .A1(n19784), .A2(n19783), .Z(n16351) );
  INV_X2 U18219 ( .I(n29446), .ZN(n27597) );
  AND2_X2 U18246 ( .A1(n13391), .A2(n27745), .Z(n14094) );
  OAI22_X2 U18247 ( .A1(n16358), .A2(n18433), .B1(n18432), .B2(n5269), .ZN(
        n27683) );
  INV_X2 U18255 ( .I(n25654), .ZN(n25650) );
  NOR2_X2 U18261 ( .A1(n13911), .A2(n27604), .ZN(n9831) );
  XOR2_X1 U18267 ( .A1(n12370), .A2(n21768), .Z(n21769) );
  NAND2_X1 U18277 ( .A1(n18184), .A2(n17416), .ZN(n2802) );
  XOR2_X1 U18295 ( .A1(n14094), .A2(n27607), .Z(n15357) );
  NOR2_X1 U18321 ( .A1(n8051), .A2(n947), .ZN(n18715) );
  NAND2_X1 U18358 ( .A1(n3181), .A2(n31862), .ZN(n14813) );
  XOR2_X1 U18389 ( .A1(n1714), .A2(n10979), .Z(n9459) );
  NAND2_X2 U18408 ( .A1(n28683), .A2(n14134), .ZN(n20404) );
  INV_X1 U18416 ( .I(n17061), .ZN(n28685) );
  NAND3_X1 U18429 ( .A1(n19893), .A2(n14545), .A3(n19894), .ZN(n27627) );
  OAI21_X2 U18437 ( .A1(n31987), .A2(n18692), .B(n952), .ZN(n27628) );
  NOR2_X1 U18438 ( .A1(n7418), .A2(n27629), .ZN(n7420) );
  NOR2_X1 U18441 ( .A1(n7417), .A2(n7415), .ZN(n27629) );
  AOI22_X2 U18488 ( .A1(n19902), .A2(n16637), .B1(n19903), .B2(n27938), .ZN(
        n19904) );
  INV_X4 U18491 ( .I(n692), .ZN(n25229) );
  BUF_X2 U18496 ( .I(n9592), .Z(n27638) );
  AOI21_X2 U18506 ( .A1(n2147), .A2(n19867), .B(n2146), .ZN(n14138) );
  NAND2_X1 U18509 ( .A1(n18798), .A2(n7712), .ZN(n7898) );
  NOR2_X1 U18517 ( .A1(n18803), .A2(n12317), .ZN(n27641) );
  XOR2_X1 U18522 ( .A1(Plaintext[24]), .A2(Key[24]), .Z(n15455) );
  INV_X2 U18523 ( .I(n27642), .ZN(n632) );
  XOR2_X1 U18526 ( .A1(n10461), .A2(n10462), .Z(n27642) );
  XOR2_X1 U18531 ( .A1(n27645), .A2(n32759), .Z(n24855) );
  XOR2_X1 U18535 ( .A1(n24645), .A2(n15671), .Z(n27645) );
  BUF_X2 U18554 ( .I(n725), .Z(n27652) );
  NAND2_X2 U18564 ( .A1(n20619), .A2(n20620), .ZN(n21029) );
  AOI21_X2 U18569 ( .A1(n17542), .A2(n20024), .B(n27654), .ZN(n20345) );
  OAI22_X1 U18575 ( .A1(n20123), .A2(n16595), .B1(n20022), .B2(n20021), .ZN(
        n27654) );
  OR2_X2 U18576 ( .A1(n22617), .A2(n15401), .Z(n23753) );
  OR2_X1 U18611 ( .A1(n25923), .A2(n14359), .Z(n27659) );
  OAI22_X2 U18613 ( .A1(n25348), .A2(n31941), .B1(n25347), .B2(n25346), .ZN(
        n25376) );
  XOR2_X1 U18616 ( .A1(n27664), .A2(n25131), .Z(Ciphertext[59]) );
  XOR2_X1 U18618 ( .A1(n16200), .A2(n13907), .Z(n4562) );
  AND2_X2 U18626 ( .A1(n19053), .A2(n30663), .Z(n12052) );
  OAI21_X2 U18635 ( .A1(n7904), .A2(n7905), .B(n22552), .ZN(n27719) );
  NAND2_X2 U18649 ( .A1(n15820), .A2(n21740), .ZN(n22031) );
  OR2_X1 U18654 ( .A1(n22641), .A2(n10725), .Z(n5648) );
  XOR2_X1 U18682 ( .A1(n17659), .A2(n27672), .Z(n449) );
  AOI21_X2 U18689 ( .A1(n13659), .A2(n15520), .B(n29473), .ZN(n13658) );
  NOR2_X1 U18709 ( .A1(n298), .A2(n30281), .ZN(n27680) );
  XOR2_X1 U18733 ( .A1(n20958), .A2(n20959), .Z(n8076) );
  BUF_X2 U18741 ( .I(n12951), .Z(n27687) );
  NOR2_X2 U18742 ( .A1(n10113), .A2(n865), .ZN(n27688) );
  NAND2_X1 U18752 ( .A1(n1279), .A2(n23017), .ZN(n22963) );
  OR2_X1 U18753 ( .A1(n22791), .A2(n14392), .Z(n15391) );
  NAND3_X2 U18755 ( .A1(n28442), .A2(n19024), .A3(n19026), .ZN(n19658) );
  NAND2_X2 U18767 ( .A1(n19302), .A2(n730), .ZN(n27696) );
  NAND2_X2 U18770 ( .A1(n23658), .A2(n23657), .ZN(n12356) );
  NAND3_X1 U18777 ( .A1(n867), .A2(n1156), .A3(n6679), .ZN(n8996) );
  XOR2_X1 U18784 ( .A1(n22195), .A2(n22193), .Z(n11423) );
  XOR2_X1 U18791 ( .A1(n27703), .A2(n1067), .Z(Ciphertext[53]) );
  AOI22_X1 U18794 ( .A1(n3208), .A2(n25082), .B1(n1203), .B2(n5520), .ZN(
        n27703) );
  NAND2_X2 U18800 ( .A1(n16747), .A2(n19717), .ZN(n6255) );
  XOR2_X1 U18804 ( .A1(n702), .A2(n19539), .Z(n17931) );
  NOR2_X2 U18816 ( .A1(n18816), .A2(n18714), .ZN(n27709) );
  XOR2_X1 U18823 ( .A1(n28262), .A2(n20775), .Z(n1848) );
  INV_X2 U18828 ( .I(n23157), .ZN(n707) );
  INV_X2 U18834 ( .I(n20569), .ZN(n816) );
  XOR2_X1 U18843 ( .A1(n10685), .A2(n321), .Z(n11172) );
  XOR2_X1 U18850 ( .A1(n5402), .A2(n27717), .Z(n5401) );
  OAI22_X2 U18857 ( .A1(n19606), .A2(n3388), .B1(n9356), .B2(n826), .ZN(n27718) );
  NAND2_X1 U18862 ( .A1(n13312), .A2(n12323), .ZN(n27720) );
  OR3_X1 U18873 ( .A1(n4066), .A2(n19156), .A3(n18599), .Z(n19160) );
  XOR2_X1 U18878 ( .A1(n27721), .A2(n9475), .Z(n3144) );
  XOR2_X1 U18882 ( .A1(n3146), .A2(n24781), .Z(n27721) );
  NAND2_X2 U18892 ( .A1(n2903), .A2(n19934), .ZN(n18078) );
  NAND2_X2 U18906 ( .A1(n24179), .A2(n24178), .ZN(n24512) );
  XOR2_X1 U18913 ( .A1(n1612), .A2(n1613), .Z(n21100) );
  NAND2_X2 U18917 ( .A1(n7826), .A2(n27724), .ZN(n13478) );
  OR2_X1 U18920 ( .A1(n13481), .A2(n13482), .Z(n27724) );
  XOR2_X1 U18926 ( .A1(n26255), .A2(n11349), .Z(n28541) );
  INV_X1 U18936 ( .I(n32052), .ZN(n27729) );
  INV_X1 U18944 ( .I(n20674), .ZN(n28803) );
  XOR2_X1 U18952 ( .A1(n12801), .A2(n27728), .Z(n5137) );
  NAND2_X2 U18958 ( .A1(n6864), .A2(n19921), .ZN(n19844) );
  NAND2_X2 U18962 ( .A1(n12879), .A2(n20336), .ZN(n20842) );
  INV_X2 U18967 ( .I(n27732), .ZN(n10787) );
  XOR2_X1 U18976 ( .A1(n15308), .A2(n24783), .Z(n24173) );
  NAND3_X1 U18980 ( .A1(n14795), .A2(n25222), .A3(n15340), .ZN(n5174) );
  INV_X2 U18983 ( .I(n27736), .ZN(n17305) );
  XOR2_X1 U18992 ( .A1(n21992), .A2(n10205), .Z(n7639) );
  XOR2_X1 U19006 ( .A1(n16893), .A2(n30007), .Z(n21986) );
  OAI21_X1 U19011 ( .A1(n16749), .A2(n16750), .B(n6516), .ZN(n27745) );
  INV_X2 U19017 ( .I(n27747), .ZN(n469) );
  XOR2_X1 U19018 ( .A1(Plaintext[186]), .A2(Key[186]), .Z(n27747) );
  NAND2_X2 U19025 ( .A1(n21956), .A2(n8853), .ZN(n23301) );
  NAND2_X2 U19033 ( .A1(n27756), .A2(n14924), .ZN(n24087) );
  NOR2_X1 U19034 ( .A1(n15330), .A2(n16276), .ZN(n27758) );
  XOR2_X1 U19035 ( .A1(n11337), .A2(n11338), .Z(n13195) );
  NAND2_X2 U19044 ( .A1(n1351), .A2(n20447), .ZN(n20224) );
  XOR2_X1 U19060 ( .A1(n23319), .A2(n3620), .Z(n3619) );
  AOI22_X2 U19068 ( .A1(n27769), .A2(n27768), .B1(n9506), .B2(n8120), .ZN(
        n7925) );
  OAI22_X1 U19085 ( .A1(n13568), .A2(n8450), .B1(n25985), .B2(n10227), .ZN(
        n2517) );
  AOI21_X2 U19086 ( .A1(n27775), .A2(n29329), .B(n13835), .ZN(n13834) );
  NAND2_X2 U19094 ( .A1(n27776), .A2(n28084), .ZN(n2902) );
  NAND2_X1 U19097 ( .A1(n18303), .A2(n18304), .ZN(n27776) );
  NAND2_X1 U19100 ( .A1(n13953), .A2(n13952), .ZN(n29095) );
  NOR2_X2 U19102 ( .A1(n5704), .A2(n25975), .ZN(n21716) );
  XOR2_X1 U19126 ( .A1(n27375), .A2(n1592), .Z(n27778) );
  AOI21_X1 U19136 ( .A1(n7361), .A2(n24327), .B(n28030), .ZN(n28029) );
  AOI22_X2 U19141 ( .A1(n23982), .A2(n28538), .B1(n5286), .B2(n24325), .ZN(
        n24785) );
  AOI22_X2 U19151 ( .A1(n12105), .A2(n28436), .B1(n14891), .B2(n5913), .ZN(
        n14890) );
  NAND2_X2 U19184 ( .A1(n10523), .A2(n20173), .ZN(n17554) );
  INV_X2 U19201 ( .I(n27797), .ZN(n18648) );
  XNOR2_X1 U19202 ( .A1(Key[38]), .A2(Plaintext[38]), .ZN(n27797) );
  AND2_X1 U19209 ( .A1(n18648), .A2(n18649), .Z(n17113) );
  XOR2_X1 U19214 ( .A1(n27243), .A2(n11897), .Z(n22516) );
  XOR2_X1 U19236 ( .A1(n5212), .A2(n27179), .Z(n3491) );
  XOR2_X1 U19242 ( .A1(n2362), .A2(n2363), .Z(n2366) );
  XOR2_X1 U19264 ( .A1(n412), .A2(n27804), .Z(n2022) );
  XOR2_X1 U19271 ( .A1(n1676), .A2(n26033), .Z(n27804) );
  NAND2_X1 U19273 ( .A1(n822), .A2(n13348), .ZN(n27805) );
  XOR2_X1 U19276 ( .A1(n11490), .A2(n19740), .Z(n11222) );
  OAI22_X2 U19302 ( .A1(n11050), .A2(n12680), .B1(n23786), .B2(n23785), .ZN(
        n15692) );
  INV_X2 U19328 ( .I(n1266), .ZN(n22953) );
  XOR2_X1 U19333 ( .A1(n4291), .A2(n13298), .Z(n14605) );
  INV_X2 U19351 ( .I(n27819), .ZN(n16205) );
  OAI21_X1 U19362 ( .A1(n3136), .A2(n24972), .B(n3135), .ZN(n3134) );
  XOR2_X1 U19371 ( .A1(n15887), .A2(n24549), .Z(n27823) );
  NOR2_X1 U19376 ( .A1(n28954), .A2(n13735), .ZN(n29004) );
  OR2_X1 U19399 ( .A1(n8558), .A2(n20136), .Z(n27829) );
  NAND2_X1 U19413 ( .A1(n10501), .A2(n25608), .ZN(n27833) );
  OAI22_X1 U19427 ( .A1(n1376), .A2(n30501), .B1(n31254), .B2(n10943), .ZN(
        n14354) );
  XOR2_X1 U19438 ( .A1(n29262), .A2(n14684), .Z(n335) );
  INV_X2 U19449 ( .I(n27838), .ZN(n28668) );
  XNOR2_X1 U19450 ( .A1(n7890), .A2(n28748), .ZN(n27838) );
  OR2_X1 U19482 ( .A1(n32747), .A2(n11086), .Z(n28857) );
  XOR2_X1 U19490 ( .A1(Plaintext[5]), .A2(Key[5]), .Z(n27936) );
  XOR2_X1 U19503 ( .A1(n28239), .A2(n21894), .Z(n21896) );
  OAI22_X2 U19522 ( .A1(n27845), .A2(n24285), .B1(n27500), .B2(n24284), .ZN(
        n24478) );
  AND2_X1 U19523 ( .A1(n28275), .A2(n4604), .Z(n27845) );
  NAND2_X2 U19526 ( .A1(n15965), .A2(n7736), .ZN(n16144) );
  XOR2_X1 U19530 ( .A1(n23366), .A2(n26116), .Z(n28811) );
  XOR2_X1 U19546 ( .A1(n227), .A2(n6924), .Z(n2839) );
  XOR2_X1 U19572 ( .A1(n22161), .A2(n22110), .Z(n22019) );
  NAND2_X2 U19575 ( .A1(n27857), .A2(n18438), .ZN(n19355) );
  INV_X2 U19597 ( .I(n6168), .ZN(n24526) );
  NAND2_X2 U19598 ( .A1(n2939), .A2(n27998), .ZN(n6168) );
  BUF_X2 U19599 ( .I(n23508), .Z(n27860) );
  NOR2_X2 U19600 ( .A1(n21), .A2(n21857), .ZN(n21691) );
  NOR3_X1 U19614 ( .A1(n6939), .A2(n25707), .A3(n25705), .ZN(n27861) );
  XOR2_X1 U19624 ( .A1(n17659), .A2(n20904), .Z(n5282) );
  NAND2_X1 U19626 ( .A1(n19287), .A2(n19021), .ZN(n19026) );
  XNOR2_X1 U19660 ( .A1(n8568), .A2(n16691), .ZN(n29205) );
  NAND2_X2 U19665 ( .A1(n27867), .A2(n13973), .ZN(n13972) );
  NAND2_X2 U19686 ( .A1(n580), .A2(n20614), .ZN(n20455) );
  INV_X2 U19720 ( .I(n15734), .ZN(n28190) );
  NOR2_X1 U19724 ( .A1(n3495), .A2(n29158), .ZN(n3494) );
  XOR2_X1 U19735 ( .A1(n16590), .A2(n28457), .Z(n578) );
  AND2_X1 U19738 ( .A1(n21392), .A2(n27170), .Z(n2602) );
  XOR2_X1 U19752 ( .A1(n20982), .A2(n20891), .Z(n20673) );
  NAND2_X1 U19757 ( .A1(n27873), .A2(n27872), .ZN(n25281) );
  NAND2_X1 U19758 ( .A1(n30281), .A2(n25276), .ZN(n27872) );
  OAI21_X2 U19781 ( .A1(n12111), .A2(n16546), .B(n14692), .ZN(n28450) );
  XOR2_X1 U19784 ( .A1(n22231), .A2(n29121), .Z(n4763) );
  AND2_X1 U19790 ( .A1(n14650), .A2(n14954), .Z(n16810) );
  NOR2_X2 U19807 ( .A1(n19301), .A2(n16354), .ZN(n19085) );
  INV_X2 U19809 ( .I(n27883), .ZN(n5191) );
  XOR2_X1 U19815 ( .A1(n19558), .A2(n25998), .Z(n27884) );
  NAND2_X1 U19821 ( .A1(n28704), .A2(n4577), .ZN(n18119) );
  NAND2_X2 U19824 ( .A1(n1297), .A2(n22660), .ZN(n22446) );
  XOR2_X1 U19835 ( .A1(n16733), .A2(n32683), .Z(n673) );
  AOI21_X2 U19837 ( .A1(n24034), .A2(n24033), .B(n24032), .ZN(n16733) );
  AND2_X1 U19849 ( .A1(n2180), .A2(n3994), .Z(n24934) );
  NAND2_X2 U19855 ( .A1(n14355), .A2(n274), .ZN(n19698) );
  XOR2_X1 U19875 ( .A1(n4944), .A2(n9434), .Z(n27895) );
  MUX2_X1 U19880 ( .I0(n27430), .I1(n12904), .S(n24305), .Z(n24034) );
  INV_X2 U19883 ( .I(n18146), .ZN(n24305) );
  XOR2_X1 U19884 ( .A1(n16989), .A2(n27896), .Z(n11934) );
  XOR2_X1 U19885 ( .A1(n673), .A2(n16394), .Z(n27896) );
  NAND2_X2 U19892 ( .A1(n8024), .A2(n30010), .ZN(n19004) );
  NAND2_X2 U19895 ( .A1(n10307), .A2(n10306), .ZN(n8024) );
  NOR3_X2 U19908 ( .A1(n10687), .A2(n13), .A3(n24042), .ZN(n27899) );
  NAND2_X2 U19929 ( .A1(n21617), .A2(n21614), .ZN(n6489) );
  XOR2_X1 U19933 ( .A1(n6373), .A2(n13844), .Z(n23460) );
  INV_X2 U19938 ( .I(n27907), .ZN(n29255) );
  XOR2_X1 U19942 ( .A1(n6273), .A2(n8076), .Z(n27907) );
  OAI21_X2 U19948 ( .A1(n8222), .A2(n14081), .B(n12472), .ZN(n22968) );
  AOI21_X2 U19962 ( .A1(n18478), .A2(n18477), .B(n18476), .ZN(n19461) );
  XOR2_X1 U19964 ( .A1(n22037), .A2(n10887), .Z(n8328) );
  NAND3_X2 U19974 ( .A1(n15004), .A2(n437), .A3(n436), .ZN(n19122) );
  NAND2_X2 U19976 ( .A1(n27914), .A2(n26060), .ZN(n14770) );
  NAND3_X1 U19984 ( .A1(n53), .A2(n32481), .A3(n29774), .ZN(n7834) );
  INV_X2 U19994 ( .I(n31324), .ZN(n12500) );
  XOR2_X1 U19997 ( .A1(n19433), .A2(n27919), .Z(n3932) );
  XOR2_X1 U19998 ( .A1(n33749), .A2(n27920), .Z(n27919) );
  NAND2_X2 U20003 ( .A1(n28309), .A2(n29667), .ZN(n20283) );
  XOR2_X1 U20015 ( .A1(n12048), .A2(n14908), .Z(n19541) );
  NAND2_X2 U20016 ( .A1(n13706), .A2(n13705), .ZN(n19651) );
  XOR2_X1 U20020 ( .A1(n14716), .A2(n27923), .Z(n8249) );
  OR2_X1 U20048 ( .A1(n20037), .A2(n27911), .Z(n19835) );
  NAND2_X1 U20049 ( .A1(n21204), .A2(n27955), .ZN(n16197) );
  OAI21_X2 U20051 ( .A1(n4539), .A2(n4538), .B(n4536), .ZN(n3421) );
  INV_X1 U20057 ( .I(n19460), .ZN(n28453) );
  XOR2_X1 U20070 ( .A1(n15028), .A2(n19424), .Z(n19443) );
  NOR2_X1 U20085 ( .A1(n18662), .A2(n18678), .ZN(n18450) );
  NAND2_X2 U20098 ( .A1(n27930), .A2(n27929), .ZN(n4387) );
  INV_X2 U20138 ( .I(n27936), .ZN(n18884) );
  BUF_X2 U20142 ( .I(n21842), .Z(n27937) );
  INV_X2 U20155 ( .I(n21429), .ZN(n27939) );
  XNOR2_X1 U20156 ( .A1(n22211), .A2(n22210), .ZN(n28873) );
  XOR2_X1 U20186 ( .A1(n27946), .A2(n6328), .Z(n6820) );
  NOR2_X1 U20210 ( .A1(n6300), .A2(n22956), .ZN(n16203) );
  XOR2_X1 U20243 ( .A1(n14733), .A2(n15923), .Z(n27952) );
  OAI21_X2 U20246 ( .A1(n18407), .A2(n9401), .B(n27953), .ZN(n19322) );
  NOR3_X1 U20266 ( .A1(n11845), .A2(n24315), .A3(n13232), .ZN(n12188) );
  OAI21_X1 U20270 ( .A1(n33721), .A2(n13499), .B(n17878), .ZN(n14266) );
  INV_X2 U20279 ( .I(n27957), .ZN(n572) );
  INV_X2 U20292 ( .I(n27960), .ZN(n29268) );
  NAND2_X1 U20296 ( .A1(n27962), .A2(n27961), .ZN(n2421) );
  INV_X1 U20300 ( .I(n24675), .ZN(n27962) );
  XOR2_X1 U20314 ( .A1(n7686), .A2(n7684), .Z(n17450) );
  NOR2_X1 U20320 ( .A1(n27963), .A2(n14490), .ZN(n15818) );
  OAI21_X2 U20332 ( .A1(n15841), .A2(n33783), .B(n2778), .ZN(n17515) );
  XOR2_X1 U20343 ( .A1(n27968), .A2(n24993), .Z(Ciphertext[27]) );
  NAND3_X1 U20360 ( .A1(n27969), .A2(n23027), .A3(n16976), .ZN(n22749) );
  NAND2_X2 U20375 ( .A1(n27972), .A2(n11448), .ZN(n13553) );
  XOR2_X1 U20390 ( .A1(n32286), .A2(n8548), .Z(n12121) );
  OR2_X1 U20404 ( .A1(n469), .A2(n26049), .Z(n4927) );
  XOR2_X1 U20415 ( .A1(n8053), .A2(n8054), .Z(n27976) );
  NOR2_X1 U20435 ( .A1(n676), .A2(n25564), .ZN(n3922) );
  XOR2_X1 U20446 ( .A1(n304), .A2(n24560), .Z(n27977) );
  NAND2_X1 U20447 ( .A1(n23825), .A2(n14164), .ZN(n13721) );
  NOR2_X1 U20452 ( .A1(n16849), .A2(n31579), .ZN(n27980) );
  NAND2_X2 U20473 ( .A1(n8962), .A2(n8963), .ZN(n10510) );
  NOR2_X2 U20489 ( .A1(n9500), .A2(n9502), .ZN(n16458) );
  INV_X4 U20493 ( .I(n12700), .ZN(n12586) );
  NAND2_X1 U20494 ( .A1(n22983), .A2(n12700), .ZN(n22800) );
  NOR2_X2 U20495 ( .A1(n27994), .A2(n27993), .ZN(n12700) );
  XOR2_X1 U20501 ( .A1(n28163), .A2(n27995), .Z(n453) );
  XOR2_X1 U20505 ( .A1(n5472), .A2(n20836), .Z(n20916) );
  NOR2_X1 U20510 ( .A1(n23842), .A2(n23887), .ZN(n28016) );
  XOR2_X1 U20515 ( .A1(n12478), .A2(n16958), .Z(n8526) );
  XOR2_X1 U20524 ( .A1(n22023), .A2(n28000), .Z(n110) );
  XOR2_X1 U20533 ( .A1(n19515), .A2(n28004), .Z(n16590) );
  XOR2_X1 U20539 ( .A1(n28908), .A2(n26000), .Z(n28004) );
  BUF_X2 U20544 ( .I(n22185), .Z(n28005) );
  NAND2_X2 U20557 ( .A1(n19839), .A2(n19838), .ZN(n20507) );
  INV_X2 U20565 ( .I(n28014), .ZN(n28865) );
  NOR2_X1 U20572 ( .A1(n4182), .A2(n724), .ZN(n6382) );
  OAI22_X1 U20576 ( .A1(n9438), .A2(n14156), .B1(n955), .B2(n15406), .ZN(
        n14652) );
  XOR2_X1 U20623 ( .A1(n18050), .A2(n28027), .Z(n18049) );
  XOR2_X1 U20688 ( .A1(n3630), .A2(n3627), .Z(n18197) );
  INV_X2 U20695 ( .I(n28034), .ZN(n667) );
  NAND2_X2 U20704 ( .A1(n13284), .A2(n13283), .ZN(n20519) );
  OAI21_X2 U20721 ( .A1(n7051), .A2(n21178), .B(n28038), .ZN(n21581) );
  XOR2_X1 U20723 ( .A1(n2333), .A2(n2334), .Z(n28039) );
  NAND2_X1 U20775 ( .A1(n4425), .A2(n31914), .ZN(n6244) );
  OR2_X1 U20796 ( .A1(n11072), .A2(n19315), .Z(n11070) );
  OAI21_X1 U20816 ( .A1(n18587), .A2(n18532), .B(n33205), .ZN(n18530) );
  XOR2_X1 U20826 ( .A1(n28052), .A2(n25669), .Z(Ciphertext[143]) );
  INV_X2 U20830 ( .I(n21454), .ZN(n6493) );
  NAND2_X1 U20833 ( .A1(n780), .A2(n27912), .ZN(n11292) );
  XOR2_X1 U20840 ( .A1(n17804), .A2(n603), .Z(n21454) );
  XNOR2_X1 U20863 ( .A1(n12609), .A2(n6789), .ZN(n28086) );
  XOR2_X1 U20897 ( .A1(n28057), .A2(n18065), .Z(n16695) );
  XOR2_X1 U20903 ( .A1(n17958), .A2(n6376), .Z(n28057) );
  NOR2_X2 U20915 ( .A1(n11596), .A2(n14864), .ZN(n28059) );
  XOR2_X1 U20920 ( .A1(n22178), .A2(n22177), .Z(n22179) );
  XOR2_X1 U20960 ( .A1(n23496), .A2(n23118), .Z(n28062) );
  NAND2_X2 U20986 ( .A1(n14539), .A2(n12004), .ZN(n12329) );
  XOR2_X1 U21001 ( .A1(n6454), .A2(n22056), .Z(n22312) );
  NAND2_X1 U21029 ( .A1(n17673), .A2(n24565), .ZN(n25344) );
  INV_X4 U21039 ( .I(n17855), .ZN(n10031) );
  XOR2_X1 U21052 ( .A1(n7411), .A2(n51), .Z(n28072) );
  OAI21_X1 U21090 ( .A1(n14331), .A2(n9553), .B(n19249), .ZN(n8672) );
  INV_X2 U21095 ( .I(n28078), .ZN(n6860) );
  XOR2_X1 U21096 ( .A1(Plaintext[160]), .A2(Key[160]), .Z(n28078) );
  XOR2_X1 U21102 ( .A1(n17423), .A2(n14206), .Z(n20773) );
  XNOR2_X1 U21130 ( .A1(n9517), .A2(n19516), .ZN(n28174) );
  AOI22_X1 U21157 ( .A1(n18301), .A2(n13279), .B1(n18302), .B2(n18722), .ZN(
        n28084) );
  INV_X2 U21189 ( .I(n12895), .ZN(n20099) );
  XOR2_X1 U21212 ( .A1(n24684), .A2(n6646), .Z(n28093) );
  AND2_X1 U21230 ( .A1(n15216), .A2(n6860), .Z(n18858) );
  OAI21_X1 U21231 ( .A1(n27719), .A2(n27007), .B(n17408), .ZN(n22825) );
  NOR2_X1 U21235 ( .A1(n25760), .A2(n17120), .ZN(n24437) );
  INV_X2 U21243 ( .I(n18150), .ZN(n28096) );
  OR2_X1 U21253 ( .A1(n18638), .A2(n9437), .Z(n9438) );
  XOR2_X1 U21255 ( .A1(n23233), .A2(n29231), .Z(n28100) );
  NAND2_X2 U21262 ( .A1(n11086), .A2(n12966), .ZN(n20426) );
  NAND3_X1 U21265 ( .A1(n28102), .A2(n18855), .A3(n26068), .ZN(n5154) );
  XOR2_X1 U21269 ( .A1(n23358), .A2(n23306), .Z(n23236) );
  XOR2_X1 U21277 ( .A1(n16128), .A2(n8548), .Z(n24382) );
  NOR2_X2 U21278 ( .A1(n7098), .A2(n7100), .ZN(n16128) );
  INV_X2 U21294 ( .I(n3535), .ZN(n28104) );
  INV_X2 U21295 ( .I(n19133), .ZN(n28105) );
  INV_X2 U21300 ( .I(n30281), .ZN(n1207) );
  AOI22_X1 U21324 ( .A1(n20617), .A2(n32594), .B1(n7873), .B2(n20616), .ZN(
        n20620) );
  XOR2_X1 U21328 ( .A1(n28109), .A2(n8596), .Z(n17638) );
  AOI21_X2 U21335 ( .A1(n21672), .A2(n21673), .B(n28111), .ZN(n7641) );
  INV_X1 U21343 ( .I(n28114), .ZN(n28113) );
  OAI21_X1 U21344 ( .A1(n888), .A2(n23665), .B(n23382), .ZN(n28114) );
  XOR2_X1 U21356 ( .A1(n28116), .A2(n16598), .Z(Ciphertext[146]) );
  XOR2_X1 U21363 ( .A1(n23244), .A2(n530), .Z(n13131) );
  XOR2_X1 U21368 ( .A1(n28118), .A2(n23276), .Z(n10659) );
  INV_X1 U21369 ( .I(n23383), .ZN(n28118) );
  NAND2_X2 U21388 ( .A1(n7376), .A2(n3104), .ZN(n10720) );
  XOR2_X1 U21390 ( .A1(n9569), .A2(n9567), .Z(n28121) );
  XOR2_X1 U21408 ( .A1(n4414), .A2(n4411), .Z(n28123) );
  OR2_X1 U21412 ( .A1(n20527), .A2(n20566), .Z(n28126) );
  XNOR2_X1 U21414 ( .A1(n16946), .A2(n16945), .ZN(n28751) );
  NAND2_X2 U21439 ( .A1(n10234), .A2(n15640), .ZN(n22255) );
  XOR2_X1 U21464 ( .A1(n20983), .A2(n11118), .Z(n28134) );
  NAND2_X2 U21487 ( .A1(n14233), .A2(n14194), .ZN(n19050) );
  INV_X2 U21505 ( .I(n28142), .ZN(n2967) );
  NAND2_X2 U21513 ( .A1(n3885), .A2(n6722), .ZN(n25689) );
  NAND2_X1 U21527 ( .A1(n24921), .A2(n24933), .ZN(n24348) );
  XOR2_X1 U21553 ( .A1(n10255), .A2(n28150), .Z(n15496) );
  XOR2_X1 U21555 ( .A1(n9307), .A2(n15452), .Z(n28150) );
  INV_X2 U21556 ( .I(n28151), .ZN(n11621) );
  INV_X2 U21566 ( .I(n16291), .ZN(n733) );
  XOR2_X1 U21580 ( .A1(n17775), .A2(n28152), .Z(n8432) );
  XOR2_X1 U21581 ( .A1(n23286), .A2(n23297), .Z(n28152) );
  NAND3_X1 U21589 ( .A1(n12952), .A2(n8527), .A3(n9580), .ZN(n22513) );
  NAND2_X1 U21592 ( .A1(n224), .A2(n19868), .ZN(n19869) );
  OR2_X1 U21593 ( .A1(n17971), .A2(n12670), .Z(n4517) );
  NOR2_X1 U21602 ( .A1(n24874), .A2(n28520), .ZN(n28519) );
  AOI21_X1 U21613 ( .A1(n28471), .A2(n20306), .B(n28316), .ZN(n20162) );
  XOR2_X1 U21615 ( .A1(n28156), .A2(n25610), .Z(Ciphertext[135]) );
  NAND2_X1 U21632 ( .A1(n18251), .A2(n21740), .ZN(n28158) );
  XOR2_X1 U21633 ( .A1(n20686), .A2(n2976), .Z(n2756) );
  XOR2_X1 U21634 ( .A1(n20766), .A2(n20921), .Z(n20686) );
  NAND2_X1 U21638 ( .A1(n11406), .A2(n10670), .ZN(n6380) );
  XOR2_X1 U21669 ( .A1(n3739), .A2(n27171), .Z(n13702) );
  NAND2_X2 U21680 ( .A1(n7462), .A2(n882), .ZN(n9555) );
  NAND2_X2 U21682 ( .A1(n9805), .A2(n9363), .ZN(n25765) );
  NAND2_X2 U21683 ( .A1(n25701), .A2(n25703), .ZN(n9363) );
  BUF_X2 U21684 ( .I(n22428), .Z(n28170) );
  NAND2_X2 U21691 ( .A1(n4472), .A2(n28172), .ZN(n4016) );
  XOR2_X1 U21698 ( .A1(n22023), .A2(n1992), .Z(n1991) );
  NAND2_X1 U21700 ( .A1(n17624), .A2(n21341), .ZN(n10468) );
  OAI22_X2 U21703 ( .A1(n5978), .A2(n21076), .B1(n9842), .B2(n21243), .ZN(
        n5830) );
  XOR2_X1 U21709 ( .A1(n28174), .A2(n12803), .Z(n562) );
  XOR2_X1 U21731 ( .A1(n20825), .A2(n25910), .Z(n16775) );
  NAND2_X2 U21732 ( .A1(n20233), .A2(n285), .ZN(n20825) );
  XOR2_X1 U21762 ( .A1(n28179), .A2(n10507), .Z(n10505) );
  NOR2_X2 U21776 ( .A1(n23749), .A2(n23757), .ZN(n8330) );
  XOR2_X1 U21780 ( .A1(n22229), .A2(n16971), .Z(n5196) );
  XOR2_X1 U21833 ( .A1(n24761), .A2(n1225), .Z(n28188) );
  NAND2_X1 U21853 ( .A1(n9858), .A2(n837), .ZN(n11046) );
  NOR2_X2 U21868 ( .A1(n18997), .A2(n18996), .ZN(n28197) );
  NAND2_X2 U21869 ( .A1(n3915), .A2(n20097), .ZN(n19878) );
  XOR2_X1 U21886 ( .A1(n5148), .A2(n16841), .Z(n12750) );
  NAND2_X1 U21889 ( .A1(n30937), .A2(n29102), .ZN(n3091) );
  NAND2_X1 U21945 ( .A1(n14795), .A2(n25215), .ZN(n25217) );
  XOR2_X1 U21950 ( .A1(n17126), .A2(n17125), .Z(n17127) );
  OR2_X1 U21958 ( .A1(n295), .A2(n16144), .Z(n2622) );
  XOR2_X1 U21964 ( .A1(n28216), .A2(n19492), .Z(n6693) );
  NOR2_X2 U21995 ( .A1(n10397), .A2(n8543), .ZN(n10511) );
  OAI21_X2 U21997 ( .A1(n9242), .A2(n32037), .B(n32858), .ZN(n9243) );
  INV_X1 U22000 ( .I(n5713), .ZN(n28228) );
  XNOR2_X1 U22014 ( .A1(n17400), .A2(n23519), .ZN(n29194) );
  INV_X4 U22015 ( .I(n701), .ZN(n28473) );
  AOI21_X2 U22022 ( .A1(n11078), .A2(n977), .B(n11077), .ZN(n28235) );
  OAI21_X1 U22030 ( .A1(n3915), .A2(n27832), .B(n30692), .ZN(n8549) );
  XOR2_X1 U22034 ( .A1(n32052), .A2(n21028), .Z(n2976) );
  INV_X2 U22041 ( .I(n28236), .ZN(n9678) );
  NAND2_X2 U22057 ( .A1(n17907), .A2(n12116), .ZN(n19252) );
  BUF_X2 U22080 ( .I(n9342), .Z(n28240) );
  OR2_X1 U22090 ( .A1(n25470), .A2(n25476), .Z(n28243) );
  XNOR2_X1 U22098 ( .A1(Plaintext[146]), .A2(Key[146]), .ZN(n28245) );
  NAND2_X2 U22118 ( .A1(n10387), .A2(n10386), .ZN(n28697) );
  XOR2_X1 U22130 ( .A1(n19574), .A2(n16792), .Z(n13780) );
  XOR2_X1 U22134 ( .A1(n28251), .A2(n16698), .Z(Ciphertext[141]) );
  NAND3_X1 U22139 ( .A1(n28252), .A2(n15185), .A3(n15295), .ZN(n15184) );
  INV_X1 U22144 ( .I(n12235), .ZN(n28252) );
  OAI21_X2 U22151 ( .A1(n23752), .A2(n7895), .B(n31984), .ZN(n6716) );
  BUF_X2 U22156 ( .I(n24755), .Z(n28258) );
  INV_X2 U22195 ( .I(n15092), .ZN(n28266) );
  NOR2_X1 U22206 ( .A1(n25093), .A2(n32857), .ZN(n28270) );
  XOR2_X1 U22213 ( .A1(n21044), .A2(n16322), .Z(n7138) );
  XOR2_X1 U22227 ( .A1(n23337), .A2(n23338), .Z(n14103) );
  NAND2_X2 U22243 ( .A1(n10481), .A2(n10485), .ZN(n14597) );
  NAND2_X2 U22263 ( .A1(n16050), .A2(n34108), .ZN(n2535) );
  NAND2_X1 U22268 ( .A1(n27188), .A2(n28096), .ZN(n28283) );
  AND2_X1 U22278 ( .A1(n19451), .A2(n4180), .Z(n3593) );
  NAND2_X2 U22279 ( .A1(n7952), .A2(n7951), .ZN(n20959) );
  BUF_X2 U22311 ( .I(n10001), .Z(n28288) );
  XOR2_X1 U22321 ( .A1(n28289), .A2(n12957), .Z(n4021) );
  NAND2_X2 U22322 ( .A1(n20275), .A2(n20274), .ZN(n12957) );
  XOR2_X1 U22342 ( .A1(n31043), .A2(n31966), .Z(n8827) );
  NAND2_X1 U22357 ( .A1(n19224), .A2(n5610), .ZN(n4366) );
  AND2_X1 U22387 ( .A1(n6474), .A2(n23872), .Z(n9813) );
  AOI21_X1 U22388 ( .A1(n6097), .A2(n25475), .B(n28302), .ZN(n6095) );
  OR2_X1 U22397 ( .A1(n17151), .A2(n32082), .Z(n29021) );
  NAND2_X2 U22401 ( .A1(n17404), .A2(n32917), .ZN(n24039) );
  OAI21_X2 U22417 ( .A1(n8841), .A2(n8840), .B(n28304), .ZN(n5578) );
  OAI21_X2 U22433 ( .A1(n5163), .A2(n1249), .B(n9736), .ZN(n28307) );
  OAI21_X2 U22437 ( .A1(n933), .A2(n1636), .B(n15213), .ZN(n28309) );
  XOR2_X1 U22450 ( .A1(n23290), .A2(n28311), .Z(n29203) );
  XOR2_X1 U22453 ( .A1(n14242), .A2(n23289), .Z(n28311) );
  AOI21_X2 U22460 ( .A1(n5851), .A2(n31102), .B(n5849), .ZN(n5848) );
  INV_X2 U22467 ( .I(n28312), .ZN(n635) );
  OR2_X1 U22482 ( .A1(n8457), .A2(n13652), .Z(n12725) );
  NOR2_X1 U22531 ( .A1(n11454), .A2(n2387), .ZN(n28451) );
  XOR2_X1 U22538 ( .A1(n29876), .A2(n16685), .Z(n462) );
  XOR2_X1 U22553 ( .A1(Plaintext[12]), .A2(Key[12]), .Z(n28321) );
  AND2_X1 U22555 ( .A1(n5191), .A2(n13413), .Z(n23758) );
  NAND2_X1 U22585 ( .A1(n25666), .A2(n25650), .ZN(n25643) );
  NAND2_X2 U22588 ( .A1(n25640), .A2(n15184), .ZN(n25666) );
  XOR2_X1 U22593 ( .A1(n28331), .A2(n16464), .Z(Ciphertext[186]) );
  OR2_X1 U22600 ( .A1(n9831), .A2(n14980), .Z(n9833) );
  NAND2_X2 U22603 ( .A1(n17405), .A2(n32745), .ZN(n19820) );
  NAND2_X2 U22614 ( .A1(n28332), .A2(n13865), .ZN(n13864) );
  NAND2_X2 U22637 ( .A1(n12586), .A2(n28697), .ZN(n15364) );
  NAND2_X2 U22640 ( .A1(n15696), .A2(n18074), .ZN(n7680) );
  NOR2_X2 U22641 ( .A1(n7726), .A2(n28796), .ZN(n15696) );
  XOR2_X1 U22654 ( .A1(n528), .A2(n23205), .Z(n6294) );
  NAND2_X2 U22660 ( .A1(n12863), .A2(n28686), .ZN(n9667) );
  XOR2_X1 U22662 ( .A1(n28903), .A2(n3635), .Z(n2163) );
  NAND2_X2 U22668 ( .A1(n4508), .A2(n4507), .ZN(n28885) );
  NOR2_X1 U22670 ( .A1(n19822), .A2(n9619), .ZN(n28856) );
  NOR2_X1 U22671 ( .A1(n18650), .A2(n18373), .ZN(n16196) );
  NAND3_X1 U22707 ( .A1(n1247), .A2(n27136), .A3(n23860), .ZN(n5685) );
  XOR2_X1 U22719 ( .A1(n9274), .A2(n5558), .Z(n28354) );
  OR2_X1 U22720 ( .A1(n7305), .A2(n15359), .Z(n5621) );
  XOR2_X1 U22727 ( .A1(n10865), .A2(n26003), .Z(n10863) );
  XOR2_X1 U22735 ( .A1(n20987), .A2(n20988), .Z(n2820) );
  OR2_X1 U22759 ( .A1(n22674), .A2(n10568), .Z(n13105) );
  NOR2_X1 U22773 ( .A1(n23847), .A2(n26114), .ZN(n17980) );
  OAI21_X1 U22775 ( .A1(n18775), .A2(n18556), .B(n29074), .ZN(n29073) );
  NAND3_X1 U22779 ( .A1(n20014), .A2(n20013), .A3(n5267), .ZN(n28366) );
  OR2_X1 U22792 ( .A1(n627), .A2(n5379), .Z(n2793) );
  INV_X2 U22853 ( .I(n28373), .ZN(n1926) );
  NAND2_X2 U22871 ( .A1(n11464), .A2(n20222), .ZN(n20729) );
  NAND2_X2 U22872 ( .A1(n16785), .A2(n21267), .ZN(n21265) );
  OAI22_X2 U22879 ( .A1(n1534), .A2(n21748), .B1(n1532), .B2(n1533), .ZN(
        n22211) );
  XOR2_X1 U22880 ( .A1(n28399), .A2(n16322), .Z(n28859) );
  AND2_X1 U22902 ( .A1(n2964), .A2(n2107), .Z(n28381) );
  NOR2_X1 U22905 ( .A1(n28383), .A2(n2107), .ZN(n28382) );
  AOI21_X2 U22950 ( .A1(n9686), .A2(n28838), .B(n28393), .ZN(n9691) );
  NAND2_X2 U22975 ( .A1(n28397), .A2(n3794), .ZN(n8515) );
  NAND2_X1 U22976 ( .A1(n9957), .A2(n9402), .ZN(n28397) );
  BUF_X2 U22978 ( .I(n19197), .Z(n28399) );
  OAI21_X2 U22986 ( .A1(n3797), .A2(n3796), .B(n5997), .ZN(n22005) );
  OAI22_X2 U23013 ( .A1(n25767), .A2(n25766), .B1(n25764), .B2(n25765), .ZN(
        n25795) );
  OR2_X1 U23019 ( .A1(n14780), .A2(n29243), .Z(n11518) );
  OAI22_X1 U23043 ( .A1(n25207), .A2(n5173), .B1(n5043), .B2(n715), .ZN(n5172)
         );
  INV_X2 U23045 ( .I(n28407), .ZN(n29269) );
  INV_X2 U23055 ( .I(n9625), .ZN(n28410) );
  XOR2_X1 U23101 ( .A1(n22206), .A2(n28416), .Z(n29162) );
  XOR2_X1 U23103 ( .A1(n1308), .A2(n22205), .Z(n28416) );
  NOR2_X1 U23118 ( .A1(n3663), .A2(n12408), .ZN(n28418) );
  AOI21_X2 U23122 ( .A1(n12232), .A2(n12110), .B(n28420), .ZN(n206) );
  XOR2_X1 U23125 ( .A1(n19522), .A2(n28421), .Z(n12057) );
  XOR2_X1 U23126 ( .A1(n28601), .A2(n28422), .Z(n28421) );
  NOR2_X2 U23129 ( .A1(n28426), .A2(n28425), .ZN(n263) );
  XOR2_X1 U23140 ( .A1(n22288), .A2(n22289), .Z(n9911) );
  INV_X2 U23143 ( .I(n28430), .ZN(n20080) );
  NAND3_X2 U23155 ( .A1(n28437), .A2(n13867), .A3(n29676), .ZN(n13865) );
  NAND3_X1 U23160 ( .A1(n28438), .A2(n18855), .A3(n8411), .ZN(n8554) );
  XNOR2_X1 U23170 ( .A1(n22048), .A2(n22148), .ZN(n21931) );
  XOR2_X1 U23172 ( .A1(n9000), .A2(n1128), .Z(n28441) );
  NAND2_X1 U23187 ( .A1(n13426), .A2(n19021), .ZN(n19022) );
  NAND2_X1 U23188 ( .A1(n8227), .A2(n17817), .ZN(n28442) );
  XOR2_X1 U23195 ( .A1(n19579), .A2(n19480), .Z(n17300) );
  XOR2_X1 U23197 ( .A1(n28443), .A2(n5663), .Z(n17214) );
  NAND2_X2 U23216 ( .A1(n28444), .A2(n18452), .ZN(n19764) );
  XOR2_X1 U23239 ( .A1(n7160), .A2(n11476), .Z(n28446) );
  NAND2_X1 U23248 ( .A1(n28447), .A2(n18973), .ZN(n16725) );
  XOR2_X1 U23255 ( .A1(n9154), .A2(n6294), .Z(n9152) );
  XOR2_X1 U23261 ( .A1(n12422), .A2(n13496), .Z(n28448) );
  NOR2_X1 U23263 ( .A1(n18088), .A2(n15753), .ZN(n28449) );
  XOR2_X1 U23302 ( .A1(n15527), .A2(n28458), .Z(n28457) );
  BUF_X2 U23312 ( .I(n23318), .Z(n28460) );
  XOR2_X1 U23317 ( .A1(n20639), .A2(n28461), .Z(n16820) );
  XOR2_X1 U23325 ( .A1(n29241), .A2(n28462), .Z(n28461) );
  XOR2_X1 U23334 ( .A1(n24455), .A2(n24454), .Z(n24456) );
  XOR2_X1 U23335 ( .A1(n8703), .A2(n14727), .Z(n24454) );
  XOR2_X1 U23337 ( .A1(n2483), .A2(n25993), .Z(n15485) );
  NAND2_X2 U23345 ( .A1(n14734), .A2(n28466), .ZN(n19298) );
  OR2_X1 U23346 ( .A1(n19296), .A2(n19297), .Z(n28466) );
  XOR2_X1 U23350 ( .A1(n27165), .A2(n12539), .Z(n10582) );
  INV_X1 U23353 ( .I(n8519), .ZN(n22553) );
  NAND2_X1 U23357 ( .A1(n11451), .A2(n34161), .ZN(n8519) );
  NAND2_X1 U23373 ( .A1(n16627), .A2(n32532), .ZN(n10244) );
  OR2_X1 U23381 ( .A1(n701), .A2(n32532), .Z(n22572) );
  NAND2_X1 U23390 ( .A1(n25357), .A2(n25367), .ZN(n28469) );
  NAND2_X1 U23393 ( .A1(n25356), .A2(n30400), .ZN(n28470) );
  XOR2_X1 U23397 ( .A1(n19711), .A2(n7530), .Z(n15527) );
  NAND2_X2 U23400 ( .A1(n4914), .A2(n19059), .ZN(n7530) );
  XOR2_X1 U23401 ( .A1(n8715), .A2(n12212), .Z(n8714) );
  NAND2_X2 U23404 ( .A1(n5633), .A2(n5634), .ZN(n16052) );
  NAND2_X2 U23406 ( .A1(n28475), .A2(n28474), .ZN(n22848) );
  OR2_X1 U23412 ( .A1(n11737), .A2(n34125), .Z(n28474) );
  NOR2_X2 U23414 ( .A1(n22026), .A2(n3186), .ZN(n28475) );
  NOR2_X2 U23423 ( .A1(n23976), .A2(n23971), .ZN(n888) );
  NAND2_X2 U23430 ( .A1(n5371), .A2(n375), .ZN(n6704) );
  XOR2_X1 U23432 ( .A1(n7530), .A2(n16464), .Z(n28479) );
  INV_X2 U23438 ( .I(n28480), .ZN(n497) );
  XOR2_X1 U23442 ( .A1(Plaintext[138]), .A2(Key[138]), .Z(n28480) );
  NOR2_X1 U23444 ( .A1(n824), .A2(n9677), .ZN(n12128) );
  NAND2_X2 U23447 ( .A1(n16357), .A2(n18636), .ZN(n19167) );
  XOR2_X1 U23453 ( .A1(n24551), .A2(n6050), .Z(n6054) );
  NAND2_X2 U23467 ( .A1(n8203), .A2(n18534), .ZN(n19285) );
  XOR2_X1 U23476 ( .A1(n28482), .A2(n12185), .Z(n14031) );
  XOR2_X1 U23479 ( .A1(n23451), .A2(n13497), .Z(n28482) );
  AOI21_X2 U23480 ( .A1(n6482), .A2(n7090), .B(n28483), .ZN(n6835) );
  NOR2_X1 U23483 ( .A1(n1284), .A2(n7090), .ZN(n28483) );
  AOI21_X2 U23493 ( .A1(n14696), .A2(n1709), .B(n14694), .ZN(n19006) );
  XOR2_X1 U23496 ( .A1(n28486), .A2(n16911), .Z(Ciphertext[41]) );
  XOR2_X1 U23510 ( .A1(n8691), .A2(n24412), .Z(n11973) );
  NAND2_X1 U23525 ( .A1(n5172), .A2(n5174), .ZN(n17933) );
  AOI21_X2 U23527 ( .A1(n11712), .A2(n10848), .B(n8869), .ZN(n9803) );
  NOR2_X2 U23537 ( .A1(n25650), .A2(n25666), .ZN(n9365) );
  OAI21_X1 U23538 ( .A1(n22338), .A2(n16166), .B(n22337), .ZN(n22339) );
  INV_X2 U23540 ( .I(n28496), .ZN(n561) );
  NAND2_X1 U23547 ( .A1(n23833), .A2(n30252), .ZN(n28497) );
  OAI22_X1 U23558 ( .A1(n5043), .A2(n25216), .B1(n15359), .B2(n15462), .ZN(
        n5577) );
  AOI22_X2 U23582 ( .A1(n13238), .A2(n15376), .B1(n13237), .B2(n13459), .ZN(
        n13236) );
  XNOR2_X1 U23583 ( .A1(n23464), .A2(n23463), .ZN(n287) );
  NAND2_X1 U23592 ( .A1(n5438), .A2(n23655), .ZN(n28503) );
  XOR2_X1 U23593 ( .A1(n3781), .A2(n542), .Z(n17703) );
  XOR2_X1 U23610 ( .A1(n8795), .A2(n27174), .Z(n28513) );
  INV_X2 U23611 ( .I(n28514), .ZN(n11985) );
  NAND2_X2 U23621 ( .A1(n13409), .A2(n13249), .ZN(n22470) );
  XOR2_X1 U23635 ( .A1(n19598), .A2(n2982), .Z(n2981) );
  OAI21_X2 U23654 ( .A1(n29123), .A2(n28525), .B(n28524), .ZN(n24789) );
  NAND2_X2 U23656 ( .A1(n1869), .A2(n1870), .ZN(n2483) );
  XOR2_X1 U23662 ( .A1(n31499), .A2(n23180), .Z(n23377) );
  AOI21_X2 U23673 ( .A1(n3482), .A2(n3481), .B(n28534), .ZN(n3483) );
  NAND2_X2 U23678 ( .A1(n1751), .A2(n28536), .ZN(n6288) );
  NAND2_X1 U23679 ( .A1(n25636), .A2(n24446), .ZN(n28536) );
  NAND2_X2 U23682 ( .A1(n22664), .A2(n22578), .ZN(n5452) );
  NAND3_X1 U23700 ( .A1(n28781), .A2(n4151), .A3(n28779), .ZN(n3213) );
  INV_X2 U23719 ( .I(n562), .ZN(n1169) );
  INV_X2 U23720 ( .I(n7677), .ZN(n19474) );
  NAND2_X2 U23722 ( .A1(n28540), .A2(n28539), .ZN(n7677) );
  OAI21_X2 U23730 ( .A1(n10259), .A2(n17981), .B(n14113), .ZN(n13826) );
  XOR2_X1 U23732 ( .A1(n6624), .A2(n28542), .Z(n17662) );
  XOR2_X1 U23738 ( .A1(n19757), .A2(n18105), .Z(n28542) );
  INV_X2 U23755 ( .I(n28545), .ZN(n22606) );
  XOR2_X1 U23774 ( .A1(n23335), .A2(n11891), .Z(n23400) );
  OAI22_X2 U23778 ( .A1(n5458), .A2(n5457), .B1(n18311), .B2(n5459), .ZN(
        n10260) );
  XOR2_X1 U23781 ( .A1(n21992), .A2(n30628), .Z(n21891) );
  XOR2_X1 U23799 ( .A1(n4601), .A2(Key[16]), .Z(n29061) );
  OAI22_X2 U23801 ( .A1(n844), .A2(n23867), .B1(n33345), .B2(n11821), .ZN(
        n1506) );
  XOR2_X1 U23805 ( .A1(n23286), .A2(n24907), .Z(n28552) );
  INV_X2 U23810 ( .I(n28554), .ZN(n9953) );
  INV_X2 U23834 ( .I(n28560), .ZN(n16528) );
  XOR2_X1 U23840 ( .A1(n17097), .A2(n17094), .Z(n28560) );
  NAND2_X1 U23846 ( .A1(n32911), .A2(n5202), .ZN(n7678) );
  XOR2_X1 U23849 ( .A1(n17377), .A2(n14755), .Z(n14753) );
  XOR2_X1 U23854 ( .A1(n19662), .A2(n19663), .Z(n19664) );
  NAND2_X1 U23858 ( .A1(n16280), .A2(n3668), .ZN(n3669) );
  NAND2_X1 U23863 ( .A1(n24705), .A2(n16650), .ZN(n28564) );
  OR2_X1 U23864 ( .A1(n13194), .A2(n21313), .Z(n28565) );
  XOR2_X1 U23868 ( .A1(n28566), .A2(n17452), .Z(n28979) );
  XOR2_X1 U23880 ( .A1(n3041), .A2(n26097), .Z(n28566) );
  NAND2_X2 U23910 ( .A1(n3336), .A2(n3334), .ZN(n24741) );
  OAI21_X2 U23927 ( .A1(n1594), .A2(n857), .B(n1001), .ZN(n28567) );
  XOR2_X1 U23936 ( .A1(n8921), .A2(n28571), .Z(n2759) );
  XOR2_X1 U23937 ( .A1(n3568), .A2(n2761), .Z(n28571) );
  INV_X1 U23958 ( .I(n23191), .ZN(n28575) );
  XOR2_X1 U23990 ( .A1(n8680), .A2(n17119), .Z(n22625) );
  XOR2_X1 U23997 ( .A1(n32124), .A2(n18100), .Z(n17141) );
  NOR2_X1 U24030 ( .A1(n443), .A2(n30139), .ZN(n442) );
  NAND2_X2 U24034 ( .A1(n11957), .A2(n25710), .ZN(n24712) );
  NOR2_X2 U24040 ( .A1(n28586), .A2(n29221), .ZN(n16309) );
  XNOR2_X1 U24051 ( .A1(n9517), .A2(n7676), .ZN(n29007) );
  XOR2_X1 U24053 ( .A1(Plaintext[7]), .A2(Key[7]), .Z(n8386) );
  NOR2_X1 U24064 ( .A1(n4040), .A2(n14903), .ZN(n4906) );
  INV_X2 U24067 ( .I(n28589), .ZN(n639) );
  XOR2_X1 U24071 ( .A1(n27145), .A2(n24836), .Z(n12943) );
  XOR2_X1 U24090 ( .A1(n19729), .A2(n28593), .Z(n17192) );
  XOR2_X1 U24091 ( .A1(n4400), .A2(n16581), .Z(n28593) );
  XNOR2_X1 U24102 ( .A1(n20707), .A2(n20708), .ZN(n28594) );
  INV_X2 U24106 ( .I(n8088), .ZN(n1333) );
  XOR2_X1 U24107 ( .A1(n9815), .A2(n28595), .Z(n8088) );
  OR2_X1 U24130 ( .A1(n21490), .A2(n423), .Z(n6146) );
  NAND2_X2 U24139 ( .A1(n28602), .A2(n3378), .ZN(n7940) );
  OAI21_X1 U24146 ( .A1(n9252), .A2(n1158), .B(n28603), .ZN(n20617) );
  INV_X2 U24148 ( .I(n28605), .ZN(n21403) );
  XOR2_X1 U24160 ( .A1(n1306), .A2(n27185), .Z(n28606) );
  OAI21_X2 U24204 ( .A1(n5590), .A2(n12793), .B(n5588), .ZN(n20924) );
  INV_X2 U24212 ( .I(n28607), .ZN(n21392) );
  INV_X2 U24233 ( .I(n28608), .ZN(n651) );
  XOR2_X1 U24285 ( .A1(n16242), .A2(n15795), .Z(n28612) );
  OAI21_X2 U24296 ( .A1(n4398), .A2(n14187), .B(n8794), .ZN(n8795) );
  XOR2_X1 U24322 ( .A1(n24808), .A2(n553), .Z(n2809) );
  AND2_X1 U24327 ( .A1(n15021), .A2(n19088), .Z(n28614) );
  OR2_X1 U24331 ( .A1(n32883), .A2(n29215), .Z(n21423) );
  INV_X2 U24339 ( .I(n28617), .ZN(n12074) );
  XOR2_X1 U24340 ( .A1(Plaintext[58]), .A2(Key[58]), .Z(n28617) );
  NOR2_X1 U24381 ( .A1(n7004), .A2(n13558), .ZN(n7003) );
  NAND2_X1 U24401 ( .A1(n14745), .A2(n16799), .ZN(n28623) );
  INV_X2 U24405 ( .I(n28624), .ZN(n14339) );
  XOR2_X1 U24408 ( .A1(n6615), .A2(n28627), .Z(n8228) );
  XOR2_X1 U24409 ( .A1(n6614), .A2(n20744), .Z(n28627) );
  XOR2_X1 U24423 ( .A1(n4161), .A2(n618), .Z(n28633) );
  XOR2_X1 U24441 ( .A1(Plaintext[106]), .A2(Key[106]), .Z(n13445) );
  XOR2_X1 U24461 ( .A1(n28636), .A2(n2045), .Z(n10255) );
  XOR2_X1 U24464 ( .A1(n10257), .A2(n24807), .Z(n28636) );
  BUF_X2 U24546 ( .I(n8398), .Z(n28641) );
  XOR2_X1 U24566 ( .A1(n13419), .A2(n24553), .Z(n24626) );
  INV_X2 U24593 ( .I(n15324), .ZN(n28649) );
  NAND2_X1 U24632 ( .A1(n28658), .A2(n25072), .ZN(n28657) );
  XOR2_X1 U24648 ( .A1(n23388), .A2(n27171), .Z(n23255) );
  XOR2_X1 U24649 ( .A1(n20788), .A2(n3705), .Z(n6088) );
  NAND2_X2 U24664 ( .A1(n10048), .A2(n18120), .ZN(n24799) );
  XOR2_X1 U24694 ( .A1(n2698), .A2(n2699), .Z(n28663) );
  NAND2_X2 U24698 ( .A1(n974), .A2(n10281), .ZN(n6319) );
  NAND2_X2 U24734 ( .A1(n33731), .A2(n1133), .ZN(n7502) );
  INV_X1 U24740 ( .I(n17167), .ZN(n28964) );
  XOR2_X1 U24771 ( .A1(n28673), .A2(n3599), .Z(n5324) );
  XOR2_X1 U24773 ( .A1(n19408), .A2(n16520), .Z(n28673) );
  AOI22_X1 U24774 ( .A1(n5543), .A2(n17273), .B1(n7928), .B2(n25247), .ZN(
        n4226) );
  NOR2_X1 U24782 ( .A1(n19183), .A2(n19105), .ZN(n15291) );
  NAND2_X2 U24785 ( .A1(n28674), .A2(n18905), .ZN(n16349) );
  XOR2_X1 U24807 ( .A1(n7630), .A2(n26028), .Z(n15669) );
  XOR2_X1 U24852 ( .A1(n1085), .A2(n24689), .Z(n5358) );
  NOR3_X2 U24867 ( .A1(n29211), .A2(n26093), .A3(n13489), .ZN(n20518) );
  NOR2_X2 U24886 ( .A1(n28696), .A2(n11769), .ZN(n14161) );
  OAI21_X2 U24891 ( .A1(n8037), .A2(n8038), .B(n12702), .ZN(n13844) );
  NAND2_X2 U24897 ( .A1(n28698), .A2(n1730), .ZN(n6286) );
  XOR2_X1 U24907 ( .A1(n5925), .A2(n26029), .Z(n7374) );
  AND2_X1 U24915 ( .A1(n9953), .A2(n639), .Z(n15464) );
  XOR2_X1 U24940 ( .A1(n15787), .A2(n15786), .Z(n15788) );
  OR2_X1 U24992 ( .A1(n11006), .A2(n19936), .Z(n28852) );
  XOR2_X1 U24999 ( .A1(n28708), .A2(n4158), .Z(n14676) );
  XOR2_X1 U25000 ( .A1(n22187), .A2(n15900), .Z(n28708) );
  NAND2_X2 U25001 ( .A1(n12599), .A2(n12598), .ZN(n15230) );
  XOR2_X1 U25015 ( .A1(n253), .A2(n28711), .Z(n28710) );
  NAND3_X2 U25028 ( .A1(n607), .A2(n28712), .A3(n10671), .ZN(n11562) );
  XOR2_X1 U25053 ( .A1(n10331), .A2(n24755), .Z(n8109) );
  NAND2_X2 U25067 ( .A1(n15058), .A2(n2270), .ZN(n25006) );
  NAND2_X2 U25078 ( .A1(n18910), .A2(n18909), .ZN(n14120) );
  OAI21_X2 U25083 ( .A1(n15486), .A2(n17311), .B(n17819), .ZN(n19599) );
  INV_X2 U25117 ( .I(n28723), .ZN(n676) );
  XOR2_X1 U25145 ( .A1(n2012), .A2(n2013), .Z(n28723) );
  NAND2_X1 U25147 ( .A1(n25664), .A2(n25650), .ZN(n7087) );
  XOR2_X1 U25148 ( .A1(n17219), .A2(n28724), .Z(n11806) );
  XOR2_X1 U25162 ( .A1(n1310), .A2(n6435), .Z(n28724) );
  NAND3_X1 U25203 ( .A1(n19597), .A2(n18668), .A3(n18669), .ZN(n8716) );
  INV_X2 U25209 ( .I(n28731), .ZN(n13360) );
  XOR2_X1 U25213 ( .A1(Plaintext[147]), .A2(Key[147]), .Z(n28731) );
  AOI22_X2 U25261 ( .A1(n2709), .A2(n4359), .B1(n2710), .B2(n21823), .ZN(
        n22196) );
  XOR2_X1 U25264 ( .A1(n28735), .A2(n25311), .Z(Ciphertext[90]) );
  XOR2_X1 U25300 ( .A1(n14000), .A2(n24686), .Z(n24783) );
  NOR2_X2 U25305 ( .A1(n3256), .A2(n3257), .ZN(n14000) );
  XOR2_X1 U25356 ( .A1(n20787), .A2(n7113), .Z(n28748) );
  INV_X2 U25375 ( .I(n28750), .ZN(n25014) );
  AOI22_X2 U25377 ( .A1(n18577), .A2(n3779), .B1(n14453), .B2(n18387), .ZN(
        n7995) );
  XOR2_X1 U25387 ( .A1(n9193), .A2(n28751), .Z(n22414) );
  XOR2_X1 U25423 ( .A1(n29190), .A2(n29206), .Z(n28753) );
  OR2_X2 U25430 ( .A1(n8251), .A2(n2450), .Z(n23885) );
  OAI22_X2 U25452 ( .A1(n28755), .A2(n8271), .B1(n414), .B2(n9651), .ZN(n7233)
         );
  OAI21_X2 U25454 ( .A1(n1059), .A2(n5834), .B(n1659), .ZN(n28755) );
  XNOR2_X1 U25494 ( .A1(n19193), .A2(n11450), .ZN(n29079) );
  INV_X2 U25497 ( .I(n10937), .ZN(n14756) );
  INV_X2 U25528 ( .I(n28763), .ZN(n8105) );
  XOR2_X1 U25535 ( .A1(n16737), .A2(n16739), .Z(n28763) );
  XOR2_X1 U25570 ( .A1(n19495), .A2(n28769), .Z(n11321) );
  XOR2_X1 U25574 ( .A1(n19637), .A2(n28908), .Z(n28769) );
  NAND2_X2 U25586 ( .A1(n28770), .A2(n14100), .ZN(n18626) );
  XOR2_X1 U25595 ( .A1(n28771), .A2(n19551), .Z(n3074) );
  XOR2_X1 U25604 ( .A1(n1370), .A2(n3076), .Z(n28771) );
  NAND2_X1 U25643 ( .A1(n24283), .A2(n26387), .ZN(n28779) );
  NOR2_X1 U25654 ( .A1(n22577), .A2(n28635), .ZN(n14220) );
  OAI21_X1 U25659 ( .A1(n1200), .A2(n24934), .B(n24933), .ZN(n7787) );
  NAND2_X2 U25660 ( .A1(n8778), .A2(n14001), .ZN(n24919) );
  XOR2_X1 U25662 ( .A1(n20733), .A2(n20891), .Z(n20765) );
  XOR2_X1 U25668 ( .A1(n12442), .A2(n15978), .Z(n19666) );
  NAND2_X2 U25670 ( .A1(n11777), .A2(n11778), .ZN(n12442) );
  INV_X1 U25675 ( .I(n24283), .ZN(n24040) );
  XNOR2_X1 U25687 ( .A1(n22182), .A2(n22181), .ZN(n29170) );
  XOR2_X1 U25708 ( .A1(n28788), .A2(n4000), .Z(n8190) );
  XOR2_X1 U25710 ( .A1(n20758), .A2(n29832), .Z(n28788) );
  OAI21_X2 U25712 ( .A1(n18486), .A2(n14284), .B(n18768), .ZN(n28789) );
  NAND2_X2 U25713 ( .A1(n7708), .A2(n7709), .ZN(n7705) );
  OAI21_X1 U25715 ( .A1(n32856), .A2(n9982), .B(n28791), .ZN(n25605) );
  AOI21_X1 U25718 ( .A1(n1034), .A2(n27177), .B(n9320), .ZN(n5219) );
  OR2_X1 U25724 ( .A1(n14331), .A2(n15050), .Z(n259) );
  NAND2_X1 U25727 ( .A1(n12195), .A2(n6213), .ZN(n6212) );
  NAND2_X1 U25729 ( .A1(n16785), .A2(n8490), .ZN(n12195) );
  XOR2_X1 U25730 ( .A1(n20806), .A2(n13590), .Z(n13456) );
  NOR2_X1 U25743 ( .A1(n7898), .A2(n9766), .ZN(n28796) );
  NAND2_X1 U25760 ( .A1(n7213), .A2(n7212), .ZN(n28797) );
  INV_X2 U25761 ( .I(n9240), .ZN(n25621) );
  XOR2_X1 U25773 ( .A1(n8522), .A2(n17833), .Z(n9240) );
  OR2_X1 U25786 ( .A1(n20605), .A2(n7892), .Z(n28799) );
  NAND2_X1 U25790 ( .A1(n28800), .A2(n28580), .ZN(n4123) );
  NOR2_X1 U25791 ( .A1(n12535), .A2(n10720), .ZN(n28800) );
  OAI21_X1 U25798 ( .A1(n16193), .A2(n16493), .B(n16105), .ZN(n11502) );
  NAND2_X2 U25799 ( .A1(n22773), .A2(n9075), .ZN(n11891) );
  XOR2_X1 U25803 ( .A1(n19629), .A2(n15978), .Z(n19441) );
  XOR2_X1 U25806 ( .A1(n8635), .A2(n16319), .Z(n28807) );
  NAND2_X2 U25813 ( .A1(n18514), .A2(n14393), .ZN(n19178) );
  XOR2_X1 U25816 ( .A1(n3190), .A2(n3191), .Z(n3192) );
  XOR2_X1 U25817 ( .A1(n20767), .A2(n21046), .Z(n28814) );
  INV_X2 U25821 ( .I(n28816), .ZN(n680) );
  XOR2_X1 U25822 ( .A1(n28817), .A2(n23522), .Z(n2972) );
  XOR2_X1 U25823 ( .A1(n9843), .A2(n2974), .Z(n28817) );
  AND2_X1 U25824 ( .A1(n29207), .A2(n11966), .Z(n4423) );
  NAND3_X1 U25826 ( .A1(n24069), .A2(n1092), .A3(n25973), .ZN(n3021) );
  XOR2_X1 U25827 ( .A1(n28818), .A2(n2190), .Z(n4338) );
  NAND2_X1 U25828 ( .A1(n12291), .A2(n12290), .ZN(n10127) );
  OAI21_X2 U25835 ( .A1(n6051), .A2(n30307), .B(n28830), .ZN(n6050) );
  XOR2_X1 U25842 ( .A1(n22202), .A2(n28835), .Z(n4140) );
  XOR2_X1 U25843 ( .A1(n28837), .A2(n24759), .Z(Ciphertext[169]) );
  OAI22_X1 U25844 ( .A1(n25825), .A2(n25812), .B1(n24721), .B2(n24720), .ZN(
        n28837) );
  AND2_X1 U25850 ( .A1(n20180), .A2(n20181), .Z(n28844) );
  XOR2_X1 U25861 ( .A1(n24562), .A2(n8112), .Z(n8110) );
  NOR2_X1 U25868 ( .A1(n25775), .A2(n15304), .ZN(n28854) );
  NOR2_X2 U25870 ( .A1(n3161), .A2(n3159), .ZN(n23328) );
  NAND2_X2 U25872 ( .A1(n415), .A2(n4595), .ZN(n253) );
  NAND2_X2 U25874 ( .A1(n13539), .A2(n13540), .ZN(n22294) );
  INV_X2 U25878 ( .I(n16275), .ZN(n21189) );
  XOR2_X1 U25881 ( .A1(n24824), .A2(n28861), .Z(n6328) );
  XOR2_X1 U25882 ( .A1(n24839), .A2(n28422), .Z(n28861) );
  NAND2_X2 U25883 ( .A1(n15381), .A2(n11006), .ZN(n6027) );
  NAND2_X2 U25890 ( .A1(n15521), .A2(n23689), .ZN(n4286) );
  XOR2_X1 U25893 ( .A1(n28870), .A2(n8917), .Z(n28975) );
  XOR2_X1 U25898 ( .A1(n6058), .A2(n28873), .Z(n28872) );
  XOR2_X1 U25909 ( .A1(n28887), .A2(n24738), .Z(Ciphertext[179]) );
  NAND2_X2 U25911 ( .A1(n12686), .A2(n14590), .ZN(n15704) );
  NAND2_X1 U25912 ( .A1(n24920), .A2(n3994), .ZN(n24930) );
  NAND2_X2 U25917 ( .A1(n16807), .A2(n16806), .ZN(n5889) );
  AOI22_X2 U25918 ( .A1(n22784), .A2(n7746), .B1(n14212), .B2(n7747), .ZN(
        n23444) );
  XOR2_X1 U25922 ( .A1(n23456), .A2(n25373), .Z(n22932) );
  XOR2_X1 U25927 ( .A1(n23430), .A2(n3589), .Z(n23254) );
  XOR2_X1 U25935 ( .A1(n23263), .A2(n26059), .Z(n28903) );
  XOR2_X1 U25938 ( .A1(n20953), .A2(n16703), .Z(n6507) );
  OAI22_X2 U25939 ( .A1(n17002), .A2(n17003), .B1(n9255), .B2(n10978), .ZN(
        n20953) );
  XOR2_X1 U25940 ( .A1(n20956), .A2(n28909), .Z(n8605) );
  XOR2_X1 U25941 ( .A1(n8485), .A2(n14854), .Z(n28909) );
  NOR2_X1 U25942 ( .A1(n32877), .A2(n24060), .ZN(n13600) );
  XOR2_X1 U25946 ( .A1(n30443), .A2(n19508), .Z(n19564) );
  NOR2_X2 U25948 ( .A1(n13279), .A2(n18580), .ZN(n29182) );
  XOR2_X1 U25951 ( .A1(n28916), .A2(n11717), .Z(n15777) );
  XOR2_X1 U25956 ( .A1(n9141), .A2(n3929), .Z(n6808) );
  NAND2_X1 U25957 ( .A1(n25606), .A2(n27262), .ZN(n28917) );
  XOR2_X1 U25958 ( .A1(n27841), .A2(n6127), .Z(n28918) );
  NAND2_X2 U25961 ( .A1(n28921), .A2(n21265), .ZN(n11214) );
  OAI21_X1 U25972 ( .A1(n25685), .A2(n32879), .B(n28931), .ZN(n25692) );
  INV_X2 U25973 ( .I(n28932), .ZN(n701) );
  XOR2_X1 U25974 ( .A1(n14786), .A2(n4140), .Z(n28932) );
  NOR2_X2 U25975 ( .A1(n28933), .A2(n17910), .ZN(n17907) );
  XOR2_X1 U25976 ( .A1(n1761), .A2(n6726), .Z(n6725) );
  INV_X2 U25982 ( .I(n4192), .ZN(n9515) );
  OAI21_X2 U25983 ( .A1(n28938), .A2(n28937), .B(n16375), .ZN(n17959) );
  NOR2_X1 U25984 ( .A1(n22524), .A2(n16665), .ZN(n28937) );
  NOR3_X1 U25985 ( .A1(n16915), .A2(n18827), .A3(n18489), .ZN(n18490) );
  XOR2_X1 U25986 ( .A1(n13198), .A2(n28941), .Z(n28940) );
  INV_X2 U25991 ( .I(n28946), .ZN(n470) );
  NAND2_X2 U25992 ( .A1(n14601), .A2(n28947), .ZN(n23450) );
  OAI21_X1 U25993 ( .A1(n22967), .A2(n22966), .B(n28948), .ZN(n28947) );
  NAND2_X1 U25998 ( .A1(n23664), .A2(n14373), .ZN(n15377) );
  XOR2_X1 U25999 ( .A1(n28953), .A2(n20803), .Z(n6683) );
  AOI21_X1 U26001 ( .A1(n3006), .A2(n13737), .B(n2103), .ZN(n28954) );
  XOR2_X1 U26002 ( .A1(n24632), .A2(n24853), .Z(n24377) );
  NOR2_X1 U26005 ( .A1(n5869), .A2(n8576), .ZN(n14004) );
  OAI21_X2 U26010 ( .A1(n8472), .A2(n8473), .B(n1256), .ZN(n28956) );
  XOR2_X1 U26017 ( .A1(n18404), .A2(Key[163]), .Z(n18586) );
  XOR2_X1 U26018 ( .A1(n24813), .A2(n8306), .Z(n17096) );
  AND2_X1 U26021 ( .A1(n22577), .A2(n22664), .Z(n14221) );
  NAND2_X2 U26024 ( .A1(n1897), .A2(n1900), .ZN(n8903) );
  OAI21_X2 U26025 ( .A1(n12021), .A2(n10848), .B(n28967), .ZN(n20351) );
  OAI22_X1 U26027 ( .A1(n14933), .A2(n24958), .B1(n965), .B2(n14932), .ZN(
        n16115) );
  NAND2_X1 U26030 ( .A1(n11401), .A2(n21651), .ZN(n28972) );
  XOR2_X1 U26034 ( .A1(n28978), .A2(n30435), .Z(n18269) );
  INV_X2 U26036 ( .I(n28979), .ZN(n11932) );
  OAI22_X2 U26037 ( .A1(n29147), .A2(n18381), .B1(n1179), .B2(n15137), .ZN(
        n19399) );
  XOR2_X1 U26048 ( .A1(n19371), .A2(n19426), .Z(n4028) );
  NAND2_X1 U26050 ( .A1(n5582), .A2(n20147), .ZN(n28982) );
  NAND2_X1 U26051 ( .A1(n981), .A2(n16431), .ZN(n17665) );
  AOI21_X1 U26052 ( .A1(n20606), .A2(n20130), .B(n7292), .ZN(n16481) );
  AOI21_X2 U26056 ( .A1(n4477), .A2(n1275), .B(n4476), .ZN(n5904) );
  NAND2_X2 U26059 ( .A1(n6025), .A2(n6026), .ZN(n18988) );
  NOR2_X1 U26060 ( .A1(n18978), .A2(n14812), .ZN(n16008) );
  NAND2_X1 U26066 ( .A1(n25666), .A2(n25653), .ZN(n28992) );
  NAND2_X2 U26070 ( .A1(n16274), .A2(n4436), .ZN(n19133) );
  INV_X2 U26071 ( .I(n3815), .ZN(n19594) );
  NAND2_X2 U26072 ( .A1(n3055), .A2(n3056), .ZN(n3815) );
  OR2_X1 U26074 ( .A1(n22937), .A2(n31824), .Z(n22943) );
  XOR2_X1 U26078 ( .A1(n5378), .A2(n5539), .Z(n28999) );
  XOR2_X1 U26079 ( .A1(n23328), .A2(n10625), .Z(n23464) );
  XOR2_X1 U26080 ( .A1(n24841), .A2(n29000), .Z(n6421) );
  OAI21_X2 U26085 ( .A1(n29002), .A2(n29001), .B(n21406), .ZN(n5801) );
  XOR2_X1 U26090 ( .A1(n5512), .A2(n27481), .Z(n11325) );
  XOR2_X1 U26091 ( .A1(n29004), .A2(n18122), .Z(Ciphertext[23]) );
  NAND3_X1 U26092 ( .A1(n25314), .A2(n25315), .A3(n32867), .ZN(n25318) );
  XOR2_X1 U26098 ( .A1(n12764), .A2(n15346), .Z(n12763) );
  XOR2_X1 U26101 ( .A1(n8491), .A2(n12454), .Z(n29009) );
  XOR2_X1 U26103 ( .A1(n8129), .A2(n15305), .Z(n29012) );
  XOR2_X1 U26114 ( .A1(n12067), .A2(n12905), .Z(n321) );
  XOR2_X1 U26115 ( .A1(n26053), .A2(n19647), .Z(n14060) );
  XOR2_X1 U26116 ( .A1(n19371), .A2(n17342), .Z(n19647) );
  XOR2_X1 U26119 ( .A1(n29320), .A2(n30183), .Z(n7471) );
  XOR2_X1 U26120 ( .A1(n29028), .A2(n9822), .Z(n9821) );
  XOR2_X1 U26121 ( .A1(n12381), .A2(n12380), .Z(n29029) );
  NAND3_X2 U26122 ( .A1(n9728), .A2(n3269), .A3(n3272), .ZN(n14049) );
  XOR2_X1 U26125 ( .A1(n18200), .A2(n29032), .Z(n18199) );
  NOR2_X1 U26128 ( .A1(n14321), .A2(n7940), .ZN(n8202) );
  XOR2_X1 U26130 ( .A1(n24794), .A2(n24795), .Z(n29033) );
  XOR2_X1 U26131 ( .A1(n20687), .A2(n20834), .Z(n7570) );
  XOR2_X1 U26132 ( .A1(n8728), .A2(n12459), .Z(n20834) );
  INV_X2 U26134 ( .I(n19951), .ZN(n29035) );
  XOR2_X1 U26137 ( .A1(n10738), .A2(n476), .Z(n29039) );
  XOR2_X1 U26146 ( .A1(n4236), .A2(n29046), .Z(n7859) );
  AOI21_X1 U26149 ( .A1(n3843), .A2(n13627), .B(n29049), .ZN(n29048) );
  NAND2_X1 U26151 ( .A1(n29051), .A2(n7503), .ZN(n7481) );
  NAND2_X1 U26152 ( .A1(n17635), .A2(n13971), .ZN(n8536) );
  NAND2_X2 U26153 ( .A1(n10062), .A2(n25897), .ZN(n7413) );
  XOR2_X1 U26157 ( .A1(n20966), .A2(n29054), .Z(n8496) );
  OAI21_X1 U26159 ( .A1(n1207), .A2(n25284), .B(n32882), .ZN(n11294) );
  OR2_X1 U26162 ( .A1(n29255), .A2(n10558), .Z(n7148) );
  XOR2_X1 U26166 ( .A1(n8630), .A2(n22066), .Z(n29057) );
  INV_X2 U26171 ( .I(n29064), .ZN(n9959) );
  NOR2_X1 U26177 ( .A1(n28987), .A2(n18556), .ZN(n10374) );
  NAND3_X2 U26182 ( .A1(n6659), .A2(n14906), .A3(n16732), .ZN(n29071) );
  OAI21_X2 U26185 ( .A1(n29073), .A2(n18561), .B(n18560), .ZN(n19123) );
  NAND2_X1 U26186 ( .A1(n18556), .A2(n16522), .ZN(n29074) );
  INV_X2 U26187 ( .I(n29075), .ZN(n23949) );
  OAI21_X1 U26190 ( .A1(n25093), .A2(n25106), .B(n18175), .ZN(n29076) );
  NAND2_X1 U26195 ( .A1(n828), .A2(n18776), .ZN(n29149) );
  BUF_X2 U26200 ( .I(n498), .Z(n29087) );
  XOR2_X1 U26201 ( .A1(n29090), .A2(n5150), .Z(n15621) );
  NOR2_X1 U26207 ( .A1(n27637), .A2(n676), .ZN(n29094) );
  AOI21_X1 U26208 ( .A1(n29095), .A2(n25830), .B(n25829), .ZN(n25833) );
  INV_X1 U26211 ( .I(n3005), .ZN(n29099) );
  OAI21_X1 U26214 ( .A1(n11939), .A2(n17331), .B(n13934), .ZN(n17330) );
  NAND3_X1 U26215 ( .A1(n24039), .A2(n23659), .A3(n14195), .ZN(n23663) );
  XOR2_X1 U26225 ( .A1(n19571), .A2(n31361), .Z(n19492) );
  NOR2_X1 U26226 ( .A1(n25005), .A2(n2876), .ZN(n29110) );
  NAND2_X1 U26228 ( .A1(n23715), .A2(n29498), .ZN(n29111) );
  XOR2_X1 U26235 ( .A1(n12212), .A2(n29119), .Z(n8416) );
  XOR2_X1 U26236 ( .A1(n14293), .A2(n11034), .Z(n29119) );
  XOR2_X1 U26238 ( .A1(n24024), .A2(n26126), .Z(n15518) );
  XOR2_X1 U26240 ( .A1(n2591), .A2(n2589), .Z(n11348) );
  NAND2_X1 U26241 ( .A1(n1951), .A2(n16809), .ZN(n12485) );
  XOR2_X1 U26243 ( .A1(n5380), .A2(n5381), .Z(n5382) );
  NAND2_X2 U26244 ( .A1(n29124), .A2(n14587), .ZN(n8058) );
  AOI21_X1 U26248 ( .A1(n5827), .A2(n5828), .B(n575), .ZN(n5826) );
  NAND3_X1 U26252 ( .A1(n30285), .A2(n25577), .A3(n6092), .ZN(n4056) );
  INV_X1 U26253 ( .I(n13541), .ZN(n29134) );
  XOR2_X1 U26259 ( .A1(n3517), .A2(n3518), .Z(n29139) );
  XOR2_X1 U26262 ( .A1(n7759), .A2(n7761), .Z(n8044) );
  XOR2_X1 U26267 ( .A1(n29236), .A2(n6545), .Z(n24470) );
  NAND2_X2 U26268 ( .A1(n5311), .A2(n29149), .ZN(n2150) );
  INV_X2 U26269 ( .I(n2971), .ZN(n8787) );
  NAND2_X1 U26272 ( .A1(n193), .A2(n13922), .ZN(n29152) );
  BUF_X2 U26274 ( .I(n23530), .Z(n29155) );
  INV_X2 U26276 ( .I(n32078), .ZN(n29158) );
  XOR2_X1 U26277 ( .A1(n29159), .A2(n8302), .Z(n12517) );
  XOR2_X1 U26278 ( .A1(n15527), .A2(n12519), .Z(n29159) );
  NOR2_X2 U26283 ( .A1(n3998), .A2(n13076), .ZN(n10974) );
  XOR2_X1 U26285 ( .A1(n7452), .A2(n29285), .Z(n20740) );
  XOR2_X1 U26287 ( .A1(n4419), .A2(n4418), .Z(n4449) );
  XOR2_X1 U26289 ( .A1(Plaintext[36]), .A2(Key[36]), .Z(n4200) );
  OAI21_X2 U26293 ( .A1(n1702), .A2(n10908), .B(n1486), .ZN(n1484) );
  XOR2_X1 U26302 ( .A1(n28939), .A2(n24801), .Z(n15471) );
  NAND2_X1 U26303 ( .A1(n29172), .A2(n32441), .ZN(n7789) );
  OAI21_X1 U26304 ( .A1(n1319), .A2(n230), .B(n6351), .ZN(n29172) );
  XOR2_X1 U26306 ( .A1(n12675), .A2(n24479), .Z(n24644) );
  XOR2_X1 U26312 ( .A1(n19634), .A2(n19675), .Z(n19444) );
  NAND2_X2 U26313 ( .A1(n19065), .A2(n7591), .ZN(n19675) );
  XOR2_X1 U26318 ( .A1(n29189), .A2(n25126), .Z(Ciphertext[56]) );
  AOI22_X1 U26319 ( .A1(n25125), .A2(n25127), .B1(n12250), .B2(n12251), .ZN(
        n29189) );
  AOI21_X2 U26326 ( .A1(n13460), .A2(n30437), .B(n10410), .ZN(n29196) );
  NAND2_X2 U26329 ( .A1(n252), .A2(n22397), .ZN(n22396) );
  NAND2_X2 U26334 ( .A1(n29634), .A2(n5317), .ZN(n24005) );
  NAND2_X1 U26340 ( .A1(n15115), .A2(n270), .ZN(n18499) );
  NAND2_X1 U26341 ( .A1(n24117), .A2(n30505), .ZN(n9374) );
  INV_X2 U26344 ( .I(n29203), .ZN(n16981) );
  XOR2_X1 U26346 ( .A1(n23444), .A2(n25213), .Z(n29206) );
  XOR2_X1 U26349 ( .A1(n2484), .A2(n9361), .Z(n4133) );
  AOI21_X1 U26351 ( .A1(n1439), .A2(n18710), .B(n328), .ZN(n18509) );
  XOR2_X1 U26352 ( .A1(Plaintext[128]), .A2(Key[128]), .Z(n11707) );
  XOR2_X1 U26357 ( .A1(n30193), .A2(n19675), .Z(n19432) );
  NAND2_X1 U26359 ( .A1(n21538), .A2(n18235), .ZN(n29212) );
  OAI21_X2 U26362 ( .A1(n29214), .A2(n9095), .B(n20875), .ZN(n21857) );
  NAND3_X2 U26366 ( .A1(n6564), .A2(n6567), .A3(n6563), .ZN(n6974) );
  INV_X2 U26374 ( .I(n21193), .ZN(n16440) );
  XOR2_X1 U26375 ( .A1(n2524), .A2(n2526), .Z(n21193) );
  XOR2_X1 U26380 ( .A1(n9013), .A2(n9010), .Z(n15917) );
  NOR2_X1 U26381 ( .A1(n25130), .A2(n25124), .ZN(n29227) );
  INV_X2 U26382 ( .I(n29228), .ZN(n1850) );
  INV_X2 U26385 ( .I(n29230), .ZN(n510) );
  NAND2_X2 U26389 ( .A1(n25136), .A2(n25135), .ZN(n25154) );
  BUF_X2 U26395 ( .I(n12792), .Z(n29234) );
  OAI21_X2 U26400 ( .A1(n15040), .A2(n8909), .B(n8908), .ZN(n19624) );
  NAND2_X2 U26401 ( .A1(n20171), .A2(n20172), .ZN(n20680) );
  XOR2_X1 U26405 ( .A1(n6079), .A2(n6078), .Z(n29244) );
  NOR2_X1 U26406 ( .A1(n19257), .A2(n19137), .ZN(n29245) );
  XOR2_X1 U26413 ( .A1(n13645), .A2(n14293), .Z(n12410) );
  INV_X2 U26415 ( .I(n12379), .ZN(n13348) );
  INV_X2 U26420 ( .I(n2956), .ZN(n3030) );
  XNOR2_X1 U26421 ( .A1(n22206), .A2(n3583), .ZN(n29260) );
  INV_X2 U26423 ( .I(n17109), .ZN(n1289) );
  AOI21_X2 U26425 ( .A1(n22020), .A2(n1117), .B(n2257), .ZN(n2256) );
  OR2_X1 U26428 ( .A1(n22707), .A2(n32089), .Z(n29266) );
  INV_X2 U26431 ( .I(n5880), .ZN(n23860) );
  XNOR2_X1 U26438 ( .A1(n1231), .A2(n16587), .ZN(n29274) );
  INV_X1 U26441 ( .I(n25150), .ZN(n25120) );
  INV_X2 U26444 ( .I(n5019), .ZN(n16632) );
  AOI21_X2 U1504 ( .A1(n18488), .A2(n14831), .B(n18490), .ZN(n9183) );
  INV_X2 U1964 ( .I(n19206), .ZN(n7176) );
  AOI21_X2 U6752 ( .A1(n6850), .A2(n31456), .B(n6849), .ZN(n2001) );
  NOR2_X2 U8793 ( .A1(n17843), .A2(n18895), .ZN(n14091) );
  INV_X2 U12023 ( .I(n26969), .ZN(n1630) );
  OR2_X1 U3103 ( .A1(n4378), .A2(n9064), .Z(n12572) );
  OAI21_X2 U8729 ( .A1(n15695), .A2(n18659), .B(n2107), .ZN(n15151) );
  INV_X2 U15014 ( .I(n14864), .ZN(n17887) );
  INV_X2 U7211 ( .I(n3192), .ZN(n11601) );
  INV_X2 U22246 ( .I(n21671), .ZN(n21668) );
  INV_X2 U11943 ( .I(n15343), .ZN(n8919) );
  NOR2_X2 U2415 ( .A1(n4835), .A2(n30817), .ZN(n11280) );
  BUF_X2 U4768 ( .I(n606), .Z(n28869) );
  INV_X2 U23141 ( .I(n32532), .ZN(n28472) );
  NAND2_X2 U2323 ( .A1(n25756), .A2(n2967), .ZN(n4708) );
  BUF_X2 U4471 ( .I(n9624), .Z(n7546) );
  INV_X4 U14451 ( .I(n9678), .ZN(n8197) );
  AOI22_X2 U7067 ( .A1(n6447), .A2(n27178), .B1(n21720), .B2(n1007), .ZN(n2393) );
  NAND2_X2 U1274 ( .A1(n14049), .A2(n17544), .ZN(n9808) );
  NOR2_X2 U1357 ( .A1(n161), .A2(n29003), .ZN(n12625) );
  NAND2_X2 U18501 ( .A1(n14010), .A2(n13168), .ZN(n18261) );
  NOR2_X2 U1131 ( .A1(n26412), .A2(n26411), .ZN(n2466) );
  AOI21_X2 U9119 ( .A1(n2023), .A2(n1732), .B(n1731), .ZN(n1730) );
  NAND2_X2 U1053 ( .A1(n20302), .A2(n20075), .ZN(n9588) );
  NOR2_X2 U1036 ( .A1(n27529), .A2(n17716), .ZN(n2395) );
  INV_X2 U20028 ( .I(n10197), .ZN(n16136) );
  NAND3_X1 U26110 ( .A1(n29020), .A2(n20022), .A3(n20021), .ZN(n19657) );
  NOR2_X2 U2707 ( .A1(n13969), .A2(n17299), .ZN(n28199) );
  INV_X4 U23943 ( .I(n17522), .ZN(n21367) );
  NOR2_X2 U3486 ( .A1(n16569), .A2(n18007), .ZN(n18835) );
  NAND3_X1 U16423 ( .A1(n27296), .A2(n22913), .A3(n29317), .ZN(n4711) );
  INV_X2 U10180 ( .I(n18101), .ZN(n1572) );
  AOI22_X2 U515 ( .A1(n22775), .A2(n15718), .B1(n18241), .B2(n31861), .ZN(
        n22777) );
  OR2_X1 U20600 ( .A1(n14329), .A2(n11443), .Z(n11442) );
  INV_X2 U1022 ( .I(n21707), .ZN(n27649) );
  INV_X2 U15785 ( .I(n19197), .ZN(n9880) );
  BUF_X4 U6937 ( .I(n23003), .Z(n13159) );
  NAND2_X2 U11034 ( .A1(n18094), .A2(n14017), .ZN(n16818) );
  NAND2_X2 U8775 ( .A1(n18705), .A2(n18743), .ZN(n18256) );
  INV_X2 U718 ( .I(n20652), .ZN(n1340) );
  NOR2_X2 U3578 ( .A1(n11460), .A2(n10182), .ZN(n18407) );
  BUF_X4 U2337 ( .I(n21350), .Z(n21566) );
  NOR2_X2 U898 ( .A1(n19325), .A2(n9646), .ZN(n19185) );
  OAI21_X2 U5425 ( .A1(n20631), .A2(n20381), .B(n8998), .ZN(n8994) );
  NOR2_X1 U1631 ( .A1(n14197), .A2(n14196), .ZN(n14311) );
  OAI21_X2 U1355 ( .A1(n3311), .A2(n9563), .B(n7804), .ZN(n1677) );
  OR2_X1 U8307 ( .A1(n22425), .A2(n22602), .Z(n12334) );
  NOR2_X2 U21451 ( .A1(n21781), .A2(n517), .ZN(n12545) );
  OAI21_X2 U12314 ( .A1(n1458), .A2(n17662), .B(n14210), .ZN(n11730) );
  INV_X2 U1006 ( .I(n17167), .ZN(n18737) );
  INV_X2 U15126 ( .I(n20565), .ZN(n20527) );
  OAI21_X2 U1474 ( .A1(n13495), .A2(n5162), .B(n24), .ZN(n8863) );
  NAND2_X2 U7538 ( .A1(n12490), .A2(n18572), .ZN(n18386) );
  INV_X2 U10190 ( .I(n18402), .ZN(n18730) );
  NAND2_X2 U6648 ( .A1(n9838), .A2(n18337), .ZN(n9837) );
  NAND2_X2 U1000 ( .A1(n18759), .A2(n18761), .ZN(n9838) );
  INV_X1 U1237 ( .I(n16847), .ZN(n10017) );
  NAND2_X2 U1059 ( .A1(n5843), .A2(n13113), .ZN(n1533) );
  NOR2_X2 U827 ( .A1(n15381), .A2(n20066), .ZN(n19935) );
  OAI21_X1 U11996 ( .A1(n6779), .A2(n6780), .B(n31139), .ZN(n1654) );
  OAI21_X2 U2615 ( .A1(n1647), .A2(n14641), .B(n6599), .ZN(n13188) );
  OAI21_X2 U2673 ( .A1(n6133), .A2(n1125), .B(n3970), .ZN(n2407) );
  NAND2_X2 U4694 ( .A1(n883), .A2(n3800), .ZN(n8542) );
  INV_X2 U22865 ( .I(n14439), .ZN(n21239) );
  NAND2_X2 U17993 ( .A1(n13657), .A2(n1039), .ZN(n13656) );
  AOI21_X2 U15431 ( .A1(n9654), .A2(n22353), .B(n8918), .ZN(n9224) );
  NAND2_X2 U2720 ( .A1(n29173), .A2(n3184), .ZN(n11383) );
  NOR2_X2 U1135 ( .A1(n1889), .A2(n26997), .ZN(n20751) );
  BUF_X2 U6350 ( .I(n8471), .Z(n7957) );
  NAND2_X2 U1494 ( .A1(n16740), .A2(n25971), .ZN(n19261) );
  INV_X4 U852 ( .I(n14210), .ZN(n1362) );
  INV_X2 U1267 ( .I(n30099), .ZN(n2566) );
  INV_X2 U23643 ( .I(n16845), .ZN(n21395) );
  INV_X2 U393 ( .I(n22983), .ZN(n22836) );
  AOI21_X2 U9338 ( .A1(n18013), .A2(n15853), .B(n18012), .ZN(n14856) );
  INV_X4 U3359 ( .I(n11985), .ZN(n13985) );
  INV_X2 U7224 ( .I(n8700), .ZN(n16639) );
  NOR2_X2 U3964 ( .A1(n20377), .A2(n20450), .ZN(n20202) );
  INV_X2 U5992 ( .I(n18459), .ZN(n11380) );
  OR2_X2 U10892 ( .A1(n15955), .A2(n28231), .Z(n18563) );
  OAI22_X2 U7398 ( .A1(n19960), .A2(n6748), .B1(n31906), .B2(n19961), .ZN(
        n6733) );
  INV_X2 U5500 ( .I(n10423), .ZN(n10015) );
  INV_X2 U5809 ( .I(n21726), .ZN(n22201) );
  AOI21_X2 U16885 ( .A1(n10374), .A2(n11864), .B(n5805), .ZN(n6025) );
  INV_X2 U9919 ( .I(n20150), .ZN(n4587) );
  INV_X2 U1303 ( .I(n20374), .ZN(n8268) );
  INV_X2 U552 ( .I(n21877), .ZN(n1315) );
  INV_X4 U7523 ( .I(n7161), .ZN(n18983) );
  INV_X1 U10928 ( .I(n30832), .ZN(n27686) );
  NAND2_X2 U5663 ( .A1(n10757), .A2(n10288), .ZN(n28160) );
  OAI21_X2 U8731 ( .A1(n31986), .A2(n2509), .B(n711), .ZN(n2508) );
  INV_X2 U6675 ( .I(n17638), .ZN(n22641) );
  INV_X2 U810 ( .I(n29101), .ZN(n29261) );
  INV_X2 U6741 ( .I(n25107), .ZN(n1203) );
  OAI21_X2 U6046 ( .A1(n32038), .A2(n7771), .B(n34057), .ZN(n7770) );
  NAND2_X2 U2522 ( .A1(n23017), .A2(n9377), .ZN(n22882) );
  AOI21_X2 U1990 ( .A1(n17112), .A2(n24005), .B(n1245), .ZN(n4521) );
  INV_X2 U945 ( .I(n11085), .ZN(n19310) );
  NOR2_X2 U2870 ( .A1(n8616), .A2(n20056), .ZN(n17713) );
  INV_X4 U1008 ( .I(n29309), .ZN(n711) );
  NAND2_X2 U2493 ( .A1(n8657), .A2(n1141), .ZN(n9906) );
  BUF_X4 U4210 ( .I(n20605), .Z(n7577) );
  AOI21_X1 U17914 ( .A1(n636), .A2(n1805), .B(n28568), .ZN(n13965) );
  OAI21_X2 U21021 ( .A1(n17764), .A2(n996), .B(n13664), .ZN(n13414) );
  CLKBUF_X4 U3889 ( .I(n23130), .Z(n23832) );
  NOR2_X2 U9380 ( .A1(n15589), .A2(n5595), .ZN(n21439) );
  BUF_X2 U3326 ( .I(n14834), .Z(n375) );
  NOR2_X2 U2202 ( .A1(n21763), .A2(n21761), .ZN(n21762) );
  INV_X2 U499 ( .I(n27799), .ZN(n23754) );
  INV_X2 U5897 ( .I(n11958), .ZN(n20055) );
  INV_X2 U3252 ( .I(n20460), .ZN(n20606) );
  NAND2_X2 U6673 ( .A1(n12238), .A2(n18891), .ZN(n6888) );
  NAND2_X2 U4818 ( .A1(n18240), .A2(n1719), .ZN(n22874) );
  NAND2_X2 U21431 ( .A1(n31726), .A2(n18973), .ZN(n15417) );
  NAND2_X2 U2473 ( .A1(n1087), .A2(n24283), .ZN(n4604) );
  INV_X2 U3548 ( .I(n16356), .ZN(n1087) );
  INV_X2 U10055 ( .I(n27921), .ZN(n17725) );
  NAND2_X1 U9881 ( .A1(n16298), .A2(n20044), .ZN(n14033) );
  INV_X1 U8022 ( .I(n1284), .ZN(n16367) );
  INV_X4 U5727 ( .I(n13998), .ZN(n23953) );
  AOI21_X2 U951 ( .A1(n11719), .A2(n21754), .B(n27649), .ZN(n6728) );
  INV_X2 U16351 ( .I(n11515), .ZN(n13367) );
  INV_X2 U12674 ( .I(n16297), .ZN(n23101) );
  NAND2_X2 U5284 ( .A1(n31982), .A2(n7190), .ZN(n4375) );
  OR2_X1 U2961 ( .A1(n4177), .A2(n28615), .Z(n17055) );
  INV_X2 U13296 ( .I(n621), .ZN(n22462) );
  NAND2_X2 U506 ( .A1(n9243), .A2(n9244), .ZN(n27126) );
  OAI22_X1 U15176 ( .A1(n25320), .A2(n16041), .B1(n25312), .B2(n25322), .ZN(
        n8629) );
  AOI22_X2 U10703 ( .A1(n33104), .A2(n4069), .B1(n23705), .B2(n23897), .ZN(
        n4536) );
  NAND2_X2 U3839 ( .A1(n27377), .A2(n14118), .ZN(n23976) );
  NAND2_X2 U6672 ( .A1(n18759), .A2(n18601), .ZN(n18289) );
  NAND2_X2 U8623 ( .A1(n29378), .A2(n12502), .ZN(n12798) );
  INV_X2 U2959 ( .I(n31095), .ZN(n18618) );
  INV_X2 U8077 ( .I(n12490), .ZN(n26318) );
  INV_X1 U5191 ( .I(n18540), .ZN(n18723) );
  NOR2_X2 U9075 ( .A1(n24139), .A2(n30969), .ZN(n9257) );
  INV_X2 U12491 ( .I(n31671), .ZN(n27097) );
  INV_X4 U6075 ( .I(n29063), .ZN(n1214) );
  NOR2_X2 U1201 ( .A1(n20406), .A2(n1349), .ZN(n15714) );
  INV_X2 U1017 ( .I(n14640), .ZN(n14641) );
  NOR2_X2 U3148 ( .A1(n7317), .A2(n6473), .ZN(n6494) );
  OAI21_X2 U21488 ( .A1(n8683), .A2(n803), .B(n8577), .ZN(n28138) );
  NAND2_X2 U5713 ( .A1(n8990), .A2(n22908), .ZN(n16898) );
  INV_X2 U1444 ( .I(n28082), .ZN(n1366) );
  NAND2_X2 U12546 ( .A1(n1655), .A2(n1654), .ZN(n11604) );
  NOR2_X2 U10001 ( .A1(n18284), .A2(n18285), .ZN(n18299) );
  INV_X4 U5859 ( .I(n5548), .ZN(n12966) );
  NOR2_X2 U2036 ( .A1(n11848), .A2(n21811), .ZN(n9206) );
  OAI21_X2 U4600 ( .A1(n12562), .A2(n861), .B(n4123), .ZN(n10491) );
  INV_X2 U15643 ( .I(n24645), .ZN(n24559) );
  INV_X2 U412 ( .I(n29294), .ZN(n23950) );
  INV_X2 U907 ( .I(n16354), .ZN(n14734) );
  NAND2_X2 U13465 ( .A1(n28831), .A2(n803), .ZN(n8577) );
  AOI21_X2 U4169 ( .A1(n23815), .A2(n6694), .B(n8525), .ZN(n26631) );
  NOR2_X2 U10725 ( .A1(n9444), .A2(n23350), .ZN(n9443) );
  BUF_X4 U6331 ( .I(n11208), .Z(n10699) );
  INV_X2 U2677 ( .I(n17641), .ZN(n25586) );
  INV_X4 U285 ( .I(n25987), .ZN(n23938) );
  INV_X4 U10835 ( .I(n26606), .ZN(n2858) );
  NAND2_X2 U8942 ( .A1(n13643), .A2(n13359), .ZN(n5810) );
  AND2_X2 U812 ( .A1(n9630), .A2(n3392), .Z(n26098) );
  NAND2_X2 U3703 ( .A1(n15149), .A2(n31614), .ZN(n2118) );
  NAND2_X1 U2460 ( .A1(n14032), .A2(n17609), .ZN(n27992) );
  BUF_X4 U1311 ( .I(n6997), .Z(n25966) );
  OAI21_X2 U5665 ( .A1(n14227), .A2(n18073), .B(n16260), .ZN(n15636) );
  AOI21_X2 U3060 ( .A1(n23074), .A2(n23073), .B(n8953), .ZN(n13690) );
  NAND2_X2 U4713 ( .A1(n13042), .A2(n14832), .ZN(n3800) );
  INV_X2 U4748 ( .I(n5051), .ZN(n12665) );
  BUF_X4 U13106 ( .I(n15144), .Z(n26891) );
  OAI21_X2 U5922 ( .A1(n32952), .A2(n4210), .B(n4714), .ZN(n5329) );
  NOR2_X2 U715 ( .A1(n22343), .A2(n7090), .ZN(n26991) );
  INV_X2 U5422 ( .I(n8795), .ZN(n10766) );
  OAI21_X2 U2699 ( .A1(n19144), .A2(n2871), .B(n19254), .ZN(n2870) );
  INV_X2 U4599 ( .I(n25966), .ZN(n1160) );
  INV_X2 U9206 ( .I(n17373), .ZN(n23826) );
  NAND3_X2 U20627 ( .A1(n20038), .A2(n20039), .A3(n20135), .ZN(n20042) );
  NOR2_X2 U1373 ( .A1(n19451), .A2(n20056), .ZN(n20053) );
  INV_X4 U2519 ( .I(n19724), .ZN(n20028) );
  AOI21_X2 U22284 ( .A1(n10273), .A2(n11350), .B(n10271), .ZN(n28285) );
  NAND2_X2 U12832 ( .A1(n16842), .A2(n29372), .ZN(n26834) );
  NOR3_X2 U2840 ( .A1(n30692), .A2(n20097), .A3(n16630), .ZN(n10241) );
  INV_X2 U1193 ( .I(n20837), .ZN(n27015) );
  INV_X2 U176 ( .I(n30795), .ZN(n968) );
  NOR2_X2 U22939 ( .A1(n24062), .A2(n24156), .ZN(n28391) );
  AOI21_X2 U8047 ( .A1(n22689), .A2(n14493), .B(n5769), .ZN(n5770) );
  AND3_X1 U3124 ( .A1(n22990), .A2(n29313), .A3(n15829), .Z(n13430) );
  BUF_X2 U8867 ( .I(Key[116]), .Z(n25910) );
  NAND2_X2 U12446 ( .A1(n27279), .A2(n16923), .ZN(n6398) );
  INV_X2 U3921 ( .I(n920), .ZN(n27024) );
  INV_X2 U15897 ( .I(n4236), .ZN(n19784) );
  AND2_X1 U2883 ( .A1(n6489), .A2(n6544), .Z(n21855) );
  INV_X2 U4033 ( .I(n16442), .ZN(n26390) );
  INV_X2 U504 ( .I(n23120), .ZN(n1262) );
  INV_X2 U5437 ( .I(n7852), .ZN(n20608) );
  INV_X4 U7033 ( .I(n22433), .ZN(n22651) );
  BUF_X2 U10229 ( .I(Key[167]), .Z(n25929) );
  INV_X2 U16428 ( .I(n16392), .ZN(n10862) );
  NOR2_X2 U1402 ( .A1(n19820), .A2(n28600), .ZN(n15246) );
  NAND2_X2 U8774 ( .A1(n18764), .A2(n27981), .ZN(n18766) );
  NAND2_X2 U1179 ( .A1(n10280), .A2(n23030), .ZN(n22738) );
  INV_X2 U302 ( .I(n5097), .ZN(n11888) );
  INV_X2 U3582 ( .I(n13348), .ZN(n1163) );
  INV_X4 U13030 ( .I(n11322), .ZN(n19267) );
  AOI21_X2 U24404 ( .A1(n18989), .A2(n18988), .B(n19034), .ZN(n18992) );
  NOR2_X2 U8690 ( .A1(n1385), .A2(n19089), .ZN(n19034) );
  INV_X2 U1259 ( .I(n9403), .ZN(n1159) );
  INV_X2 U5796 ( .I(n14297), .ZN(n3860) );
  INV_X1 U17438 ( .I(n13176), .ZN(n24217) );
  AOI21_X2 U931 ( .A1(n12545), .A2(n11861), .B(n29434), .ZN(n28155) );
  AOI21_X2 U3101 ( .A1(n9192), .A2(n16751), .B(n25186), .ZN(n8481) );
  NAND2_X2 U10536 ( .A1(n24296), .A2(n24297), .ZN(n3780) );
  BUF_X4 U5668 ( .I(n9890), .Z(n2913) );
  INV_X2 U6223 ( .I(n12821), .ZN(n1980) );
  BUF_X4 U4245 ( .I(n19285), .Z(n17311) );
  BUF_X2 U822 ( .I(n34162), .Z(n28568) );
  CLKBUF_X4 U8344 ( .I(n8605), .Z(n1146) );
  NAND2_X2 U1503 ( .A1(n784), .A2(n13200), .ZN(n27274) );
  OAI21_X2 U14671 ( .A1(n27941), .A2(n15239), .B(n10740), .ZN(n10739) );
  NAND2_X1 U13439 ( .A1(n14775), .A2(n2522), .ZN(n14774) );
  INV_X2 U4022 ( .I(n16384), .ZN(n16781) );
  OR2_X1 U2855 ( .A1(n4146), .A2(n25628), .Z(n277) );
  INV_X2 U8093 ( .I(n15617), .ZN(n22658) );
  NAND3_X2 U9615 ( .A1(n3852), .A2(n23021), .A3(n3851), .ZN(n23202) );
  INV_X2 U457 ( .I(n28123), .ZN(n4408) );
  INV_X2 U1366 ( .I(n567), .ZN(n13994) );
  INV_X2 U12825 ( .I(n398), .ZN(n16184) );
  INV_X2 U2799 ( .I(n23018), .ZN(n1279) );
  INV_X4 U7122 ( .I(n21665), .ZN(n1134) );
  NAND2_X2 U3341 ( .A1(n28328), .A2(n31798), .ZN(n15830) );
  INV_X2 U10955 ( .I(n2130), .ZN(n22722) );
  AOI21_X2 U2669 ( .A1(n21692), .A2(n21857), .B(n2797), .ZN(n15847) );
  NAND2_X2 U9230 ( .A1(n3770), .A2(n896), .ZN(n6965) );
  NOR2_X2 U5598 ( .A1(n13030), .A2(n12036), .ZN(n13029) );
  NAND2_X2 U537 ( .A1(n9844), .A2(n6236), .ZN(n26796) );
  INV_X2 U6024 ( .I(n25755), .ZN(n1212) );
  AOI21_X2 U1094 ( .A1(n7226), .A2(n21354), .B(n2088), .ZN(n3698) );
  AOI21_X2 U7820 ( .A1(n8850), .A2(n27615), .B(n8849), .ZN(n8848) );
  NAND2_X2 U1287 ( .A1(n16488), .A2(n12345), .ZN(n12344) );
  NAND3_X1 U7708 ( .A1(n4451), .A2(n24711), .A3(n4452), .ZN(n3835) );
  NOR2_X2 U5664 ( .A1(n14972), .A2(n24251), .ZN(n17581) );
  NAND2_X2 U10974 ( .A1(n12762), .A2(n23068), .ZN(n14914) );
  NOR2_X2 U6799 ( .A1(n16620), .A2(n23721), .ZN(n11812) );
  INV_X4 U123 ( .I(n4490), .ZN(n4407) );
  NAND3_X2 U1994 ( .A1(n7086), .A2(n7085), .A3(n7084), .ZN(n28251) );
  INV_X2 U1005 ( .I(n16819), .ZN(n18485) );
  NAND2_X2 U3277 ( .A1(n26750), .A2(n24106), .ZN(n24093) );
  AOI21_X2 U19409 ( .A1(n26600), .A2(n16354), .B(n4656), .ZN(n27831) );
  INV_X4 U606 ( .I(n34163), .ZN(n22981) );
  INV_X2 U4647 ( .I(n18688), .ZN(n10283) );
  BUF_X2 U7093 ( .I(n21626), .Z(n6176) );
  OAI22_X2 U26265 ( .A1(n1179), .A2(n9787), .B1(n1380), .B2(n15137), .ZN(
        n29147) );
  AOI21_X2 U1506 ( .A1(n15814), .A2(n15428), .B(n21162), .ZN(n7049) );
  INV_X2 U6264 ( .I(n6975), .ZN(n1104) );
  BUF_X4 U4247 ( .I(n19283), .Z(n13475) );
  OAI22_X2 U4372 ( .A1(n26104), .A2(n29115), .B1(n23016), .B2(n28891), .ZN(
        n13289) );
  NAND2_X2 U7016 ( .A1(n2177), .A2(n16790), .ZN(n26289) );
  INV_X2 U17035 ( .I(n29767), .ZN(n14195) );
  INV_X4 U6594 ( .I(n4747), .ZN(n1175) );
  INV_X2 U6329 ( .I(n11208), .ZN(n21799) );
  INV_X2 U41 ( .I(n14960), .ZN(n24972) );
  INV_X1 U8717 ( .I(n2902), .ZN(n19035) );
  INV_X4 U17631 ( .I(n6899), .ZN(n20489) );
  INV_X2 U885 ( .I(n5848), .ZN(n22248) );
  NAND2_X2 U6380 ( .A1(n3539), .A2(n21780), .ZN(n21583) );
  NAND2_X2 U12472 ( .A1(n10441), .A2(n10442), .ZN(n22098) );
  INV_X1 U15273 ( .I(n31960), .ZN(n15595) );
  OAI21_X2 U9865 ( .A1(n20071), .A2(n729), .B(n19888), .ZN(n18036) );
  OR2_X2 U205 ( .A1(n16552), .A2(n7171), .Z(n24342) );
  AND2_X1 U3440 ( .A1(n27921), .A2(n5889), .Z(n6566) );
  NAND2_X1 U26343 ( .A1(n20170), .A2(n20298), .ZN(n29202) );
  NOR2_X2 U10089 ( .A1(n10638), .A2(n10637), .ZN(n7286) );
  INV_X2 U5915 ( .I(n13272), .ZN(n18142) );
  BUF_X2 U5326 ( .I(n31906), .Z(n28767) );
  OAI21_X2 U24357 ( .A1(n18733), .A2(n18732), .B(n18731), .ZN(n18735) );
  INV_X2 U5615 ( .I(n17697), .ZN(n22305) );
  NAND2_X2 U1454 ( .A1(n1491), .A2(n26293), .ZN(n19682) );
  NAND2_X2 U6792 ( .A1(n23965), .A2(n13), .ZN(n18120) );
  NAND2_X2 U7186 ( .A1(n865), .A2(n2738), .ZN(n21284) );
  INV_X2 U8692 ( .I(n27242), .ZN(n13685) );
  OAI21_X2 U5639 ( .A1(n22657), .A2(n22658), .B(n16503), .ZN(n5766) );
  NOR2_X2 U2241 ( .A1(n28914), .A2(n654), .ZN(n4538) );
  CLKBUF_X2 U4287 ( .I(Key[78]), .Z(n16504) );
  INV_X4 U9064 ( .I(n24335), .ZN(n1235) );
  NOR2_X2 U8433 ( .A1(n3317), .A2(n21572), .ZN(n3316) );
  BUF_X4 U4030 ( .I(n18613), .Z(n17223) );
  NAND2_X2 U2201 ( .A1(n15022), .A2(n21761), .ZN(n21850) );
  INV_X2 U3820 ( .I(n21095), .ZN(n21408) );
  OAI21_X2 U11605 ( .A1(n13915), .A2(n33902), .B(n6083), .ZN(n15142) );
  OR3_X1 U3989 ( .A1(n18186), .A2(n1430), .A3(n6215), .Z(n10975) );
  OAI21_X2 U1398 ( .A1(n11052), .A2(n26083), .B(n11264), .ZN(n29008) );
  OAI22_X2 U6472 ( .A1(n10718), .A2(n9419), .B1(n5275), .B2(n20541), .ZN(n9418) );
  NOR2_X2 U8373 ( .A1(n26358), .A2(n17758), .ZN(n7392) );
  OR2_X2 U5369 ( .A1(n29395), .A2(n3567), .Z(n9801) );
  INV_X1 U7448 ( .I(n4386), .ZN(n4385) );
  INV_X2 U8331 ( .I(n13367), .ZN(n1141) );
  NAND2_X2 U5935 ( .A1(n12937), .A2(n4016), .ZN(n13450) );
  INV_X2 U24496 ( .I(n19419), .ZN(n19868) );
  BUF_X2 U9944 ( .I(n31671), .Z(n11199) );
  OAI21_X2 U21362 ( .A1(n27236), .A2(n16783), .B(n25520), .ZN(n25521) );
  NAND2_X2 U1189 ( .A1(n10460), .A2(n7330), .ZN(n7332) );
  INV_X2 U12423 ( .I(n16421), .ZN(n26777) );
  INV_X1 U26417 ( .I(n21375), .ZN(n21374) );
  AOI22_X2 U895 ( .A1(n17428), .A2(n17773), .B1(n21459), .B2(n21458), .ZN(
        n11795) );
  NAND2_X2 U21138 ( .A1(n17699), .A2(n29062), .ZN(n20947) );
  BUF_X4 U9928 ( .I(n15237), .Z(n20135) );
  NOR2_X2 U3554 ( .A1(n22705), .A2(n27007), .ZN(n16236) );
  BUF_X4 U26192 ( .I(n16136), .Z(n29078) );
  INV_X2 U13001 ( .I(n3084), .ZN(n20589) );
  OAI21_X2 U10117 ( .A1(n18517), .A2(n18878), .B(n18112), .ZN(n2704) );
  OAI21_X2 U7354 ( .A1(n8421), .A2(n16243), .B(n32408), .ZN(n3825) );
  OAI21_X2 U5097 ( .A1(n2443), .A2(n21716), .B(n911), .ZN(n2442) );
  NOR2_X2 U21201 ( .A1(n15872), .A2(n15506), .ZN(n14692) );
  INV_X2 U2848 ( .I(n10717), .ZN(n5275) );
  OR2_X2 U7226 ( .A1(n21184), .A2(n13989), .Z(n12756) );
  OAI21_X2 U24283 ( .A1(n16466), .A2(n18672), .B(n18441), .ZN(n18443) );
  AOI21_X2 U4842 ( .A1(n6121), .A2(n29938), .B(n3972), .ZN(n4965) );
  INV_X4 U1431 ( .I(n15110), .ZN(n27715) );
  INV_X1 U21005 ( .I(n22490), .ZN(n14671) );
  NOR2_X1 U4632 ( .A1(n1014), .A2(n12028), .ZN(n2743) );
  NOR2_X2 U13097 ( .A1(n6446), .A2(n13685), .ZN(n26890) );
  INV_X2 U5611 ( .I(n16896), .ZN(n12370) );
  NOR2_X2 U5572 ( .A1(n31927), .A2(n21), .ZN(n2797) );
  AOI22_X2 U2391 ( .A1(n11802), .A2(n1377), .B1(n26518), .B2(n10828), .ZN(
        n11801) );
  INV_X2 U5491 ( .I(n19053), .ZN(n1181) );
  OAI21_X2 U5692 ( .A1(n983), .A2(n12259), .B(n12910), .ZN(n12909) );
  INV_X2 U24023 ( .I(n17799), .ZN(n23813) );
  NOR2_X2 U2824 ( .A1(n897), .A2(n22876), .ZN(n12910) );
  INV_X2 U11490 ( .I(n5111), .ZN(n3866) );
  INV_X2 U1522 ( .I(n18626), .ZN(n19147) );
  INV_X1 U15419 ( .I(n18186), .ZN(n16624) );
  AND2_X2 U18887 ( .A1(n10303), .A2(n16332), .Z(n22479) );
  NAND2_X2 U21571 ( .A1(n4468), .A2(n15162), .ZN(n12516) );
  INV_X4 U5526 ( .I(n18815), .ZN(n785) );
  AOI21_X2 U8735 ( .A1(n4843), .A2(n1188), .B(n8043), .ZN(n4644) );
  INV_X2 U19478 ( .I(n9118), .ZN(n11918) );
  NAND2_X1 U15441 ( .A1(n10134), .A2(n33972), .ZN(n7815) );
  OAI21_X2 U5145 ( .A1(n18370), .A2(n18369), .B(n12120), .ZN(n18371) );
  NOR2_X1 U4821 ( .A1(n26953), .A2(n12010), .ZN(n8995) );
  OAI21_X2 U1742 ( .A1(n10977), .A2(n18778), .B(n10975), .ZN(n3998) );
  INV_X1 U19862 ( .I(n16202), .ZN(n28878) );
  INV_X1 U23003 ( .I(n24359), .ZN(n14832) );
  NAND2_X2 U5910 ( .A1(n23606), .A2(n23605), .ZN(n16815) );
  AOI21_X1 U12965 ( .A1(n864), .A2(n33139), .B(n2061), .ZN(n2060) );
  INV_X2 U23628 ( .I(n23696), .ZN(n16431) );
  INV_X4 U3439 ( .I(n31967), .ZN(n1347) );
  AOI21_X2 U12943 ( .A1(n12865), .A2(n11215), .B(n27608), .ZN(n12642) );
  BUF_X4 U2424 ( .I(n31448), .Z(n149) );
  INV_X2 U1441 ( .I(n29029), .ZN(n12379) );
  AND2_X2 U1501 ( .A1(n17201), .A2(n8452), .Z(n22570) );
  INV_X4 U2028 ( .I(n20092), .ZN(n15192) );
  AOI22_X2 U10106 ( .A1(n18894), .A2(n31724), .B1(n18896), .B2(n6119), .ZN(
        n6116) );
  INV_X2 U10078 ( .I(n17821), .ZN(n20155) );
  NAND2_X2 U5107 ( .A1(n497), .A2(n18747), .ZN(n18433) );
  BUF_X2 U2464 ( .I(n519), .Z(n154) );
  INV_X4 U5638 ( .I(n17960), .ZN(n12338) );
  NOR2_X2 U16864 ( .A1(n6699), .A2(n6698), .ZN(n10946) );
  BUF_X2 U10833 ( .I(n23905), .Z(n12680) );
  INV_X2 U13667 ( .I(n20080), .ZN(n20084) );
  NAND2_X1 U22425 ( .A1(n15191), .A2(n15190), .ZN(n28776) );
  INV_X4 U12317 ( .I(n25980), .ZN(n1458) );
  INV_X4 U7044 ( .I(n16124), .ZN(n17960) );
  NAND2_X2 U9101 ( .A1(n28296), .A2(n6476), .ZN(n7151) );
  INV_X4 U661 ( .I(n27752), .ZN(n28328) );
  BUF_X2 U4244 ( .I(n19360), .Z(n16444) );
  OAI21_X2 U1971 ( .A1(n26113), .A2(n16229), .B(n21817), .ZN(n5757) );
  BUF_X2 U1432 ( .I(n13510), .Z(n29208) );
  AOI21_X2 U12101 ( .A1(n18878), .A2(n18881), .B(n6754), .ZN(n6753) );
  NOR2_X2 U17829 ( .A1(n18672), .A2(n18881), .ZN(n6754) );
  OAI21_X2 U1462 ( .A1(n19170), .A2(n19171), .B(n948), .ZN(n3245) );
  NOR2_X2 U22400 ( .A1(n34005), .A2(n28721), .ZN(n19170) );
  NOR2_X2 U22728 ( .A1(n25974), .A2(n24251), .ZN(n15086) );
  NAND2_X2 U22647 ( .A1(n20139), .A2(n32141), .ZN(n15594) );
  NOR3_X1 U5166 ( .A1(n1053), .A2(n5889), .A3(n31451), .ZN(n6565) );
  NAND2_X2 U2908 ( .A1(n18722), .A2(n13279), .ZN(n18582) );
  BUF_X4 U1326 ( .I(n1736), .Z(n1632) );
  NAND2_X2 U24810 ( .A1(n21451), .A2(n20950), .ZN(n20951) );
  INV_X4 U22817 ( .I(n14458), .ZN(n20000) );
  INV_X4 U17258 ( .I(n33740), .ZN(n10757) );
  OR2_X1 U3811 ( .A1(n31970), .A2(n3093), .Z(n15284) );
  INV_X4 U13638 ( .I(n8924), .ZN(n16473) );
  AOI22_X2 U1981 ( .A1(n13210), .A2(n13925), .B1(n19046), .B2(n19047), .ZN(
        n12601) );
  BUF_X2 U2676 ( .I(n23827), .Z(n16467) );
  NAND3_X2 U25782 ( .A1(n14925), .A2(n34149), .A3(n32590), .ZN(n25913) );
  INV_X1 U11206 ( .I(n3911), .ZN(n22552) );
  OAI21_X2 U1233 ( .A1(n30602), .A2(n19256), .B(n2703), .ZN(n2124) );
  BUF_X2 U4695 ( .I(n14396), .Z(n26337) );
  OAI21_X2 U5814 ( .A1(n4668), .A2(n18043), .B(n21808), .ZN(n21727) );
  OR2_X1 U6142 ( .A1(n3773), .A2(n22977), .Z(n26026) );
  NAND2_X2 U2148 ( .A1(n5481), .A2(n11399), .ZN(n27975) );
  INV_X2 U4858 ( .I(n4740), .ZN(n4755) );
  INV_X1 U1680 ( .I(n5511), .ZN(n6901) );
  BUF_X4 U2996 ( .I(n11984), .Z(n295) );
  NAND2_X2 U7539 ( .A1(n9837), .A2(n9836), .ZN(n4571) );
  OAI22_X2 U725 ( .A1(n20416), .A2(n20415), .B1(n30931), .B2(n20414), .ZN(
        n20860) );
  INV_X2 U5057 ( .I(n32595), .ZN(n11059) );
  NAND2_X2 U451 ( .A1(n22488), .A2(n31551), .ZN(n75) );
  NOR3_X2 U1302 ( .A1(n8619), .A2(n2625), .A3(n30152), .ZN(n8618) );
  OR2_X1 U5392 ( .A1(n15713), .A2(n16167), .Z(n27299) );
  INV_X2 U12749 ( .I(n1850), .ZN(n9294) );
  NAND2_X2 U1412 ( .A1(n19884), .A2(n224), .ZN(n26357) );
  OR2_X2 U15510 ( .A1(n12654), .A2(n14290), .Z(n7205) );
  BUF_X2 U4298 ( .I(Key[96]), .Z(n16657) );
  BUF_X2 U2518 ( .I(n19698), .Z(n112) );
  BUF_X2 U2740 ( .I(n22625), .Z(n16170) );
  BUF_X2 U5507 ( .I(n11272), .Z(n6584) );
  NAND2_X2 U11440 ( .A1(n18213), .A2(n29369), .ZN(n18210) );
  OR2_X1 U2857 ( .A1(n5736), .A2(n2163), .Z(n3480) );
  INV_X1 U21925 ( .I(n16440), .ZN(n28211) );
  INV_X2 U129 ( .I(n6545), .ZN(n24771) );
  OAI21_X2 U10689 ( .A1(n23682), .A2(n23681), .B(n14124), .ZN(n23685) );
  NOR2_X2 U16763 ( .A1(n11730), .A2(n8775), .ZN(n6631) );
  NAND2_X1 U17263 ( .A1(n11213), .A2(n25658), .ZN(n11212) );
  NOR2_X1 U21252 ( .A1(n12377), .A2(n23034), .ZN(n15191) );
  INV_X2 U879 ( .I(n18453), .ZN(n1370) );
  INV_X4 U389 ( .I(n33115), .ZN(n23045) );
  BUF_X2 U2808 ( .I(n14000), .Z(n27841) );
  NAND2_X1 U5 ( .A1(n11211), .A2(n34094), .ZN(n28631) );
  NAND3_X1 U17453 ( .A1(n18361), .A2(n17792), .A3(n18362), .ZN(n18162) );
  INV_X2 U6196 ( .I(n893), .ZN(n8835) );
  AOI22_X2 U6982 ( .A1(n1669), .A2(n9580), .B1(n13079), .B2(n22599), .ZN(n1668) );
  OAI21_X2 U7162 ( .A1(n11405), .A2(n28869), .B(n21431), .ZN(n13150) );
  INV_X2 U5067 ( .I(n23000), .ZN(n16078) );
  NOR2_X2 U11161 ( .A1(n630), .A2(n28124), .ZN(n3521) );
  INV_X1 U6197 ( .I(n14398), .ZN(n13125) );
  NOR2_X2 U14822 ( .A1(n18374), .A2(n18809), .ZN(n9785) );
  INV_X4 U3108 ( .I(n635), .ZN(n16137) );
  OAI22_X2 U11717 ( .A1(n26008), .A2(n13537), .B1(n13759), .B2(n13538), .ZN(
        n13783) );
  OR2_X2 U23824 ( .A1(n5097), .A2(n29270), .Z(n23819) );
  OAI21_X2 U908 ( .A1(n27326), .A2(n864), .B(n1), .ZN(n3685) );
  OAI21_X2 U9262 ( .A1(n32595), .A2(n1275), .B(n30502), .ZN(n13460) );
  NAND2_X1 U10879 ( .A1(n8494), .A2(n17828), .ZN(n4779) );
  INV_X2 U5113 ( .I(n606), .ZN(n12925) );
  OAI21_X2 U7345 ( .A1(n15737), .A2(n10340), .B(n15735), .ZN(n19912) );
  INV_X2 U12921 ( .I(n16510), .ZN(n17717) );
  AOI22_X2 U5535 ( .A1(n12992), .A2(n10686), .B1(n15002), .B2(n7512), .ZN(
        n28664) );
  INV_X2 U5452 ( .I(n7014), .ZN(n20071) );
  BUF_X2 U7659 ( .I(Key[13]), .Z(n16696) );
  AOI21_X2 U18598 ( .A1(n18940), .A2(n19244), .B(n27818), .ZN(n18941) );
  NOR2_X2 U7295 ( .A1(n13589), .A2(n17328), .ZN(n20234) );
  INV_X2 U18458 ( .I(n10371), .ZN(n15799) );
  OAI22_X2 U2053 ( .A1(n25591), .A2(n10497), .B1(n9197), .B2(n13032), .ZN(
        n28557) );
  NAND2_X2 U8172 ( .A1(n21805), .A2(n3467), .ZN(n7501) );
  OAI21_X2 U899 ( .A1(n1766), .A2(n2283), .B(n2280), .ZN(n2279) );
  INV_X2 U5086 ( .I(n15455), .ZN(n26717) );
  CLKBUF_X4 U1539 ( .I(n19348), .Z(n27941) );
  OR2_X1 U21250 ( .A1(n22680), .A2(n32172), .Z(n12531) );
  NAND2_X2 U2052 ( .A1(n10497), .A2(n18151), .ZN(n25636) );
  INV_X4 U15707 ( .I(n30885), .ZN(n17348) );
  INV_X2 U11812 ( .I(n26278), .ZN(n1357) );
  INV_X2 U1906 ( .I(n16781), .ZN(n28671) );
  NAND2_X2 U6658 ( .A1(n6888), .A2(n6889), .ZN(n6266) );
  BUF_X4 U3406 ( .I(n8506), .Z(n29118) );
  INV_X2 U476 ( .I(n6882), .ZN(n5769) );
  NOR2_X2 U7361 ( .A1(n19884), .A2(n19868), .ZN(n20057) );
  NAND2_X2 U11451 ( .A1(n1915), .A2(n1914), .ZN(n1913) );
  NAND2_X2 U5913 ( .A1(n7730), .A2(n1237), .ZN(n6773) );
  INV_X1 U13802 ( .I(n18151), .ZN(n28097) );
  INV_X2 U3395 ( .I(n24104), .ZN(n15376) );
  OR2_X1 U3462 ( .A1(n12452), .A2(n26439), .Z(n28654) );
  NOR2_X2 U22510 ( .A1(n31402), .A2(n7310), .ZN(n14114) );
  OAI21_X2 U5393 ( .A1(n31996), .A2(n13869), .B(n26727), .ZN(n10441) );
  INV_X2 U3371 ( .I(n31074), .ZN(n19254) );
  OAI21_X1 U11072 ( .A1(n6187), .A2(n28825), .B(n5814), .ZN(n2861) );
  NOR2_X1 U11307 ( .A1(n11582), .A2(n3580), .ZN(n3579) );
  INV_X2 U18158 ( .I(n20395), .ZN(n7291) );
  INV_X4 U13502 ( .I(n11734), .ZN(n21369) );
  NAND2_X1 U11746 ( .A1(n24950), .A2(n24949), .ZN(n26711) );
  INV_X4 U14982 ( .I(n12145), .ZN(n16681) );
  NAND2_X1 U2138 ( .A1(n25256), .A2(n7871), .ZN(n26497) );
  AND2_X1 U3404 ( .A1(n19252), .A2(n8506), .Z(n18525) );
  NAND3_X1 U2566 ( .A1(n25530), .A2(n25588), .A3(n25529), .ZN(n25535) );
  OAI22_X2 U904 ( .A1(n3468), .A2(n21660), .B1(n3467), .B2(n21659), .ZN(n11053) );
  BUF_X2 U7670 ( .I(Key[17]), .Z(n25619) );
  INV_X2 U5873 ( .I(n20582), .ZN(n12872) );
  NOR2_X2 U8928 ( .A1(n9114), .A2(n23960), .ZN(n9113) );
  INV_X2 U6090 ( .I(n16321), .ZN(n7837) );
  NOR2_X1 U20872 ( .A1(n15215), .A2(n8602), .ZN(n12751) );
  NAND2_X1 U15799 ( .A1(n17172), .A2(n17171), .ZN(n4390) );
  INV_X2 U9587 ( .I(n21872), .ZN(n21871) );
  INV_X4 U3762 ( .I(n10465), .ZN(n3626) );
  NAND3_X1 U17210 ( .A1(n20487), .A2(n20252), .A3(n5878), .ZN(n11140) );
  OAI21_X2 U21533 ( .A1(n9876), .A2(n12100), .B(n20007), .ZN(n17785) );
  NAND2_X1 U22256 ( .A1(n15417), .A2(n19267), .ZN(n15416) );
  INV_X4 U2919 ( .I(n11390), .ZN(n2107) );
  NOR2_X1 U2429 ( .A1(n27971), .A2(n5936), .ZN(n5933) );
  INV_X1 U2482 ( .I(n32998), .ZN(n10018) );
  NAND2_X2 U4367 ( .A1(n27537), .A2(n26222), .ZN(n6519) );
  AOI22_X2 U15561 ( .A1(n21534), .A2(n21566), .B1(n29806), .B2(n21568), .ZN(
        n8196) );
  NAND2_X1 U16881 ( .A1(n27358), .A2(n6520), .ZN(n2369) );
  BUF_X2 U10257 ( .I(Key[107]), .Z(n25578) );
  INV_X2 U6093 ( .I(n32317), .ZN(n1232) );
  NOR2_X2 U3659 ( .A1(n7176), .A2(n30010), .ZN(n1494) );
  INV_X1 U3179 ( .I(n18874), .ZN(n961) );
  NOR2_X2 U3334 ( .A1(n30355), .A2(n2679), .ZN(n2678) );
  OAI21_X2 U21437 ( .A1(n15141), .A2(n18697), .B(n33098), .ZN(n15140) );
  INV_X2 U20675 ( .I(n20102), .ZN(n12038) );
  NOR2_X2 U15051 ( .A1(n5205), .A2(n30573), .ZN(n28863) );
  OAI21_X2 U3682 ( .A1(n10947), .A2(n11521), .B(n25997), .ZN(n18949) );
  BUF_X2 U10166 ( .I(n18434), .Z(n18705) );
  INV_X2 U12217 ( .I(n10891), .ZN(n18683) );
  NAND2_X1 U8660 ( .A1(n28157), .A2(n19236), .ZN(n2599) );
  AOI22_X2 U5672 ( .A1(n7560), .A2(n16170), .B1(n17955), .B2(n7559), .ZN(
        n27916) );
  AOI21_X2 U25895 ( .A1(n17392), .A2(n17393), .B(n3562), .ZN(n8425) );
  INV_X1 U5468 ( .I(n14340), .ZN(n27412) );
  NAND2_X1 U11408 ( .A1(n11687), .A2(n16034), .ZN(n11686) );
  NAND4_X2 U4550 ( .A1(n21829), .A2(n21828), .A3(n21827), .A4(n21832), .ZN(
        n17406) );
  NAND3_X2 U1322 ( .A1(n13994), .A2(n20028), .A3(n16461), .ZN(n12947) );
  INV_X4 U18707 ( .I(n8408), .ZN(n27678) );
  OAI21_X2 U8760 ( .A1(n18399), .A2(n2596), .B(n29309), .ZN(n2595) );
  INV_X4 U23330 ( .I(n15559), .ZN(n17624) );
  INV_X1 U6566 ( .I(n16904), .ZN(n873) );
  NAND2_X1 U24080 ( .A1(n12572), .A2(n9065), .ZN(n28592) );
  BUF_X4 U8091 ( .I(n29451), .Z(n1297) );
  NAND2_X2 U12104 ( .A1(n16338), .A2(n18576), .ZN(n8461) );
  OAI21_X2 U4912 ( .A1(n8931), .A2(n8930), .B(n8929), .ZN(n8928) );
  NAND2_X2 U11824 ( .A1(n3366), .A2(n32780), .ZN(n17786) );
  NAND3_X1 U14633 ( .A1(n9903), .A2(n24997), .A3(n9902), .ZN(n4035) );
  OR2_X1 U17288 ( .A1(n16777), .A2(n15189), .Z(n4163) );
  BUF_X2 U8153 ( .I(n21860), .Z(n3756) );
  INV_X2 U4640 ( .I(n497), .ZN(n18742) );
  NAND2_X2 U17538 ( .A1(n27981), .A2(n27980), .ZN(n14234) );
  CLKBUF_X8 U14489 ( .I(n16051), .Z(n27090) );
  INV_X2 U637 ( .I(n1104), .ZN(n29115) );
  AOI21_X2 U2640 ( .A1(n10199), .A2(n24361), .B(n680), .ZN(n15150) );
  NOR2_X1 U23026 ( .A1(n8919), .A2(n16745), .ZN(n14881) );
  INV_X4 U1647 ( .I(n18768), .ZN(n27981) );
  INV_X2 U276 ( .I(n8125), .ZN(n3165) );
  INV_X4 U5042 ( .I(n2450), .ZN(n756) );
  AOI21_X2 U6635 ( .A1(n6921), .A2(n32005), .B(n6920), .ZN(n6919) );
  INV_X1 U1811 ( .I(n14083), .ZN(n20123) );
  NOR2_X2 U11799 ( .A1(n15259), .A2(n15258), .ZN(n14711) );
  INV_X2 U12669 ( .I(n9170), .ZN(n1773) );
  NAND2_X2 U20989 ( .A1(n19196), .A2(n3388), .ZN(n19075) );
  AND2_X1 U3616 ( .A1(n32595), .A2(n7881), .Z(n10646) );
  NAND2_X1 U12695 ( .A1(n32253), .A2(n19212), .ZN(n26818) );
  NAND3_X1 U2324 ( .A1(n28531), .A2(n25309), .A3(n25315), .ZN(n28735) );
  INV_X2 U21179 ( .I(n15261), .ZN(n17832) );
  BUF_X4 U1851 ( .I(n11513), .Z(n8657) );
  INV_X4 U11389 ( .I(n1137), .ZN(n2368) );
  NOR2_X2 U23297 ( .A1(n28453), .A2(n7607), .ZN(n28452) );
  NOR2_X1 U21293 ( .A1(n13056), .A2(n23611), .ZN(n13055) );
  INV_X2 U15277 ( .I(n25198), .ZN(n25302) );
  INV_X2 U7005 ( .I(n8553), .ZN(n10206) );
  NOR2_X2 U5353 ( .A1(n10846), .A2(n14282), .ZN(n7549) );
  AOI21_X2 U2087 ( .A1(n11158), .A2(n11159), .B(n11157), .ZN(n4164) );
  INV_X1 U167 ( .I(n24499), .ZN(n24497) );
  AOI22_X2 U17441 ( .A1(n20285), .A2(n20284), .B1(n12263), .B2(n13589), .ZN(
        n27478) );
  OAI22_X2 U20507 ( .A1(n10317), .A2(n902), .B1(n10316), .B2(n1116), .ZN(
        n10315) );
  NOR3_X2 U2111 ( .A1(n15152), .A2(n883), .A3(n13050), .ZN(n9114) );
  INV_X1 U5802 ( .I(n13704), .ZN(n14253) );
  NOR2_X2 U20056 ( .A1(n22658), .A2(n9515), .ZN(n22923) );
  NOR2_X2 U12622 ( .A1(n2023), .A2(n23859), .ZN(n1731) );
  INV_X1 U18652 ( .I(n8074), .ZN(n21300) );
  NAND2_X1 U26358 ( .A1(n29212), .A2(n21540), .ZN(n15820) );
  NOR2_X2 U22432 ( .A1(n2678), .A2(n26083), .ZN(n2677) );
  BUF_X2 U6011 ( .I(Key[81]), .Z(n16301) );
  NOR2_X1 U21454 ( .A1(n28133), .A2(n28132), .ZN(n6602) );
  BUF_X4 U5171 ( .I(n13673), .Z(n13200) );
  OAI21_X2 U18897 ( .A1(n22823), .A2(n10972), .B(n22705), .ZN(n10971) );
  NAND2_X2 U19529 ( .A1(n9213), .A2(n9212), .ZN(n14882) );
  NAND2_X2 U9906 ( .A1(n12398), .A2(n19819), .ZN(n12396) );
  NAND2_X1 U18905 ( .A1(n8913), .A2(n8911), .ZN(n10003) );
  AOI21_X1 U15892 ( .A1(n27638), .A2(n29142), .B(n4500), .ZN(n8913) );
  OAI21_X2 U8293 ( .A1(n21081), .A2(n21353), .B(n3696), .ZN(n3695) );
  INV_X2 U3116 ( .I(n15966), .ZN(n18845) );
  INV_X2 U1682 ( .I(n219), .ZN(n19993) );
  OAI21_X1 U1947 ( .A1(n16954), .A2(n9793), .B(n27338), .ZN(n16955) );
  NAND3_X2 U13354 ( .A1(n2621), .A2(n2622), .A3(n27755), .ZN(n2620) );
  AOI22_X2 U22210 ( .A1(n4318), .A2(n883), .B1(n25872), .B2(n13042), .ZN(
        n14971) );
  BUF_X2 U4938 ( .I(n31161), .Z(n29003) );
  NAND2_X2 U12105 ( .A1(n9513), .A2(n7454), .ZN(n9512) );
  AOI21_X2 U5342 ( .A1(n22913), .A2(n5915), .B(n803), .ZN(n8943) );
  BUF_X2 U21781 ( .I(n15144), .Z(n14312) );
  NAND2_X2 U230 ( .A1(n13974), .A2(n33557), .ZN(n18127) );
  INV_X2 U17790 ( .I(n6693), .ZN(n19456) );
  NAND2_X2 U4403 ( .A1(n12856), .A2(n10392), .ZN(n13555) );
  NAND2_X2 U6906 ( .A1(n23047), .A2(n33007), .ZN(n23048) );
  BUF_X2 U4102 ( .I(n16799), .Z(n26314) );
  BUF_X2 U3787 ( .I(n5612), .Z(n25990) );
  NOR2_X1 U9632 ( .A1(n13692), .A2(n21357), .ZN(n11678) );
  OAI21_X2 U10122 ( .A1(n33098), .A2(n18698), .B(n18833), .ZN(n18514) );
  NAND2_X2 U7178 ( .A1(n1145), .A2(n599), .ZN(n13407) );
  NAND2_X2 U9701 ( .A1(n30813), .A2(n926), .ZN(n5469) );
  INV_X4 U6627 ( .I(n30010), .ZN(n877) );
  NAND2_X2 U15634 ( .A1(n12872), .A2(n6255), .ZN(n7978) );
  CLKBUF_X4 U4235 ( .I(n7748), .Z(n4236) );
  AOI21_X2 U8384 ( .A1(n31975), .A2(n936), .B(n12873), .ZN(n18205) );
  OAI22_X2 U5685 ( .A1(n9894), .A2(n33659), .B1(n29198), .B2(n9893), .ZN(
        n23561) );
  NAND2_X2 U7922 ( .A1(n27583), .A2(n10264), .ZN(n27582) );
  NAND2_X2 U18089 ( .A1(n10844), .A2(n17321), .ZN(n27583) );
  INV_X2 U8494 ( .I(n26374), .ZN(n24338) );
  INV_X2 U7425 ( .I(n27597), .ZN(n19853) );
  NAND3_X1 U631 ( .A1(n21449), .A2(n9518), .A3(n21451), .ZN(n1965) );
  INV_X4 U14814 ( .I(n14931), .ZN(n24955) );
  INV_X4 U8591 ( .I(n20103), .ZN(n12398) );
  NOR2_X2 U8180 ( .A1(n26955), .A2(n17701), .ZN(n13603) );
  BUF_X2 U4283 ( .I(Key[156]), .Z(n25036) );
  NAND2_X1 U10542 ( .A1(n13055), .A2(n8674), .ZN(n26579) );
  BUF_X2 U4279 ( .I(Key[40]), .Z(n25476) );
  CLKBUF_X2 U4321 ( .I(Key[174]), .Z(n25716) );
  BUF_X2 U12281 ( .I(Key[46]), .Z(n16507) );
  BUF_X2 U12272 ( .I(Key[1]), .Z(n25545) );
  BUF_X2 U4316 ( .I(Key[141]), .Z(n16533) );
  CLKBUF_X2 U4313 ( .I(Key[120]), .Z(n16679) );
  BUF_X2 U4305 ( .I(Key[37]), .Z(n8548) );
  BUF_X2 U10256 ( .I(Key[100]), .Z(n16402) );
  BUF_X2 U8850 ( .I(Key[28]), .Z(n25373) );
  BUF_X2 U10218 ( .I(Key[42]), .Z(n24964) );
  BUF_X2 U7661 ( .I(Key[178]), .Z(n25728) );
  BUF_X2 U4310 ( .I(Key[180]), .Z(n16587) );
  BUF_X2 U6727 ( .I(Key[124]), .Z(n24748) );
  INV_X1 U10205 ( .I(n25720), .ZN(n1428) );
  CLKBUF_X1 U4268 ( .I(n14159), .Z(n8411) );
  CLKBUF_X4 U3362 ( .I(n5594), .Z(n25981) );
  INV_X1 U13955 ( .I(n11605), .ZN(n10095) );
  CLKBUF_X2 U10215 ( .I(n18314), .Z(n18706) );
  BUF_X2 U6270 ( .I(n18674), .Z(n16572) );
  INV_X1 U21819 ( .I(n25358), .ZN(n15653) );
  INV_X2 U6204 ( .I(n27146), .ZN(n16915) );
  CLKBUF_X2 U3982 ( .I(n18688), .Z(n28675) );
  INV_X1 U5724 ( .I(n25071), .ZN(n27995) );
  CLKBUF_X4 U7606 ( .I(n18293), .Z(n18759) );
  NOR2_X1 U18747 ( .A1(n732), .A2(n27691), .ZN(n27690) );
  NOR2_X1 U6686 ( .A1(n16417), .A2(n16624), .ZN(n18340) );
  NOR2_X1 U8740 ( .A1(n16328), .A2(n18482), .ZN(n6252) );
  NAND2_X1 U25592 ( .A1(n18625), .A2(n16522), .ZN(n28770) );
  INV_X2 U13211 ( .I(n7134), .ZN(n2283) );
  INV_X2 U7532 ( .I(n18257), .ZN(n948) );
  INV_X2 U12473 ( .I(n8506), .ZN(n7600) );
  OR2_X1 U10083 ( .A1(n3388), .A2(n28528), .Z(n3389) );
  NOR2_X1 U1466 ( .A1(n16444), .A2(n19062), .ZN(n19364) );
  OAI21_X1 U7440 ( .A1(n3244), .A2(n3243), .B(n19175), .ZN(n3242) );
  INV_X1 U11952 ( .I(n19504), .ZN(n8504) );
  CLKBUF_X2 U3240 ( .I(n19436), .Z(n358) );
  INV_X1 U14367 ( .I(n33339), .ZN(n16852) );
  CLKBUF_X1 U3771 ( .I(n20088), .Z(n16108) );
  CLKBUF_X4 U9948 ( .I(n20102), .Z(n10947) );
  INV_X1 U11918 ( .I(n4893), .ZN(n8816) );
  NOR2_X1 U14063 ( .A1(n20013), .A2(n13605), .ZN(n27018) );
  BUF_X2 U11920 ( .I(n20083), .Z(n16664) );
  INV_X1 U5317 ( .I(n4602), .ZN(n11757) );
  NAND2_X1 U19401 ( .A1(n28826), .A2(n8558), .ZN(n27830) );
  NAND2_X1 U11874 ( .A1(n12784), .A2(n11911), .ZN(n6630) );
  NAND2_X1 U24602 ( .A1(n30794), .A2(n28644), .ZN(n19879) );
  OAI21_X1 U14062 ( .A1(n27019), .A2(n27018), .B(n20012), .ZN(n19717) );
  AOI21_X1 U5307 ( .A1(n10465), .A2(n822), .B(n20076), .ZN(n27846) );
  CLKBUF_X2 U24406 ( .I(n8057), .Z(n28625) );
  INV_X2 U2714 ( .I(n9115), .ZN(n20602) );
  NOR2_X1 U1213 ( .A1(n32903), .A2(n14265), .ZN(n14264) );
  INV_X1 U22325 ( .I(n10949), .ZN(n28289) );
  NAND3_X1 U19359 ( .A1(n26255), .A2(n13766), .A3(n13765), .ZN(n1733) );
  CLKBUF_X2 U3935 ( .I(n7124), .Z(n27285) );
  BUF_X2 U14827 ( .I(n21068), .Z(n21243) );
  INV_X2 U9712 ( .I(n3879), .ZN(n6520) );
  BUF_X2 U2448 ( .I(n21095), .Z(n151) );
  INV_X1 U1141 ( .I(n26829), .ZN(n21343) );
  OR2_X1 U19054 ( .A1(n21141), .A2(n21373), .Z(n27765) );
  INV_X2 U2530 ( .I(n21338), .ZN(n14168) );
  INV_X2 U5562 ( .I(n12221), .ZN(n17227) );
  CLKBUF_X4 U1060 ( .I(n16077), .Z(n423) );
  INV_X2 U5564 ( .I(n15172), .ZN(n6074) );
  INV_X2 U3111 ( .I(n29302), .ZN(n15026) );
  CLKBUF_X4 U12758 ( .I(n21779), .Z(n29084) );
  INV_X2 U13059 ( .I(n15863), .ZN(n15864) );
  INV_X1 U23949 ( .I(n17547), .ZN(n21785) );
  INV_X1 U9530 ( .I(n6231), .ZN(n11924) );
  INV_X1 U20683 ( .I(n27560), .ZN(n21732) );
  BUF_X2 U2903 ( .I(n8533), .Z(n28848) );
  BUF_X2 U770 ( .I(n1289), .Z(n28131) );
  BUF_X2 U4523 ( .I(n22597), .Z(n8527) );
  CLKBUF_X2 U796 ( .I(n22362), .Z(n28424) );
  NAND2_X1 U4546 ( .A1(n9752), .A2(n9751), .ZN(n10316) );
  CLKBUF_X4 U18975 ( .I(n7023), .Z(n28124) );
  INV_X2 U5082 ( .I(n22645), .ZN(n1292) );
  OAI21_X1 U25071 ( .A1(n22368), .A2(n16225), .B(n7023), .ZN(n22369) );
  INV_X2 U14138 ( .I(n11916), .ZN(n856) );
  NAND2_X1 U25103 ( .A1(n22526), .A2(n16665), .ZN(n22527) );
  NOR2_X1 U15310 ( .A1(n27298), .A2(n5035), .ZN(n9242) );
  OAI21_X1 U1257 ( .A1(n11494), .A2(n22748), .B(n3669), .ZN(n4453) );
  INV_X1 U10946 ( .I(n22860), .ZN(n14163) );
  NAND2_X1 U6735 ( .A1(n26161), .A2(n26160), .ZN(n2076) );
  INV_X1 U10838 ( .I(n23257), .ZN(n6745) );
  INV_X2 U4100 ( .I(n9152), .ZN(n14193) );
  CLKBUF_X2 U4227 ( .I(n29273), .Z(n299) );
  CLKBUF_X2 U22698 ( .I(n28615), .Z(n28347) );
  BUF_X4 U1760 ( .I(n8523), .Z(n976) );
  BUF_X2 U4207 ( .I(n10954), .Z(n29246) );
  BUF_X2 U4219 ( .I(n28765), .Z(n26965) );
  AOI21_X1 U10058 ( .A1(n26533), .A2(n23919), .B(n29185), .ZN(n8984) );
  NAND2_X1 U7835 ( .A1(n23612), .A2(n16467), .ZN(n23613) );
  NAND2_X1 U10684 ( .A1(n15615), .A2(n15642), .ZN(n15614) );
  NOR2_X1 U21907 ( .A1(n23768), .A2(n27910), .ZN(n12336) );
  NOR2_X1 U26227 ( .A1(n32434), .A2(n29111), .ZN(n4099) );
  NAND2_X1 U17413 ( .A1(n10560), .A2(n8852), .ZN(n8851) );
  NAND2_X1 U2180 ( .A1(n23752), .A2(n23726), .ZN(n26790) );
  CLKBUF_X4 U1882 ( .I(n13530), .Z(n13268) );
  INV_X2 U6693 ( .I(n15663), .ZN(n26158) );
  OAI22_X1 U9029 ( .A1(n12022), .A2(n26247), .B1(n8665), .B2(n8663), .ZN(
        n13144) );
  BUF_X2 U2000 ( .I(n10331), .Z(n27950) );
  CLKBUF_X2 U19559 ( .I(n24753), .Z(n27852) );
  CLKBUF_X4 U1694 ( .I(n91), .Z(n28939) );
  INV_X1 U4942 ( .I(n25260), .ZN(n11112) );
  NAND2_X1 U4728 ( .A1(n24605), .A2(n24606), .ZN(n3569) );
  INV_X1 U4702 ( .I(n12295), .ZN(n25148) );
  NAND2_X1 U10391 ( .A1(n24892), .A2(n31274), .ZN(n24893) );
  NAND2_X1 U15731 ( .A1(n14269), .A2(n14268), .ZN(n12679) );
  NAND3_X1 U14199 ( .A1(n28722), .A2(n26127), .A3(n25660), .ZN(n16094) );
  INV_X2 U10331 ( .I(n2180), .ZN(n15569) );
  INV_X1 U8880 ( .I(n24954), .ZN(n11469) );
  BUF_X2 U5728 ( .I(n23476), .Z(n29082) );
  NAND2_X2 U16699 ( .A1(n26612), .A2(n31549), .ZN(n4339) );
  INV_X2 U1672 ( .I(n26049), .ZN(n5700) );
  BUF_X2 U10214 ( .I(n18873), .Z(n11459) );
  BUF_X2 U13720 ( .I(n18397), .Z(n18866) );
  OAI21_X1 U6640 ( .A1(n18866), .A2(n29309), .B(n18871), .ZN(n18867) );
  NAND2_X1 U24210 ( .A1(n18481), .A2(n18601), .ZN(n18337) );
  INV_X1 U24187 ( .I(n18323), .ZN(n18567) );
  INV_X1 U6721 ( .I(n18660), .ZN(n18678) );
  BUF_X2 U5995 ( .I(n9930), .Z(n9766) );
  INV_X2 U22010 ( .I(n28231), .ZN(n18827) );
  INV_X1 U4641 ( .I(n469), .ZN(n746) );
  INV_X2 U5193 ( .I(n4677), .ZN(n8395) );
  INV_X1 U23837 ( .I(n17168), .ZN(n18489) );
  INV_X1 U4644 ( .I(n10114), .ZN(n18650) );
  INV_X1 U2607 ( .I(n18349), .ZN(n18806) );
  NAND2_X1 U10144 ( .A1(n34139), .A2(n18567), .ZN(n4550) );
  INV_X1 U4645 ( .I(n8317), .ZN(n18795) );
  NOR2_X1 U6683 ( .A1(n1389), .A2(n4925), .ZN(n26156) );
  INV_X1 U18750 ( .I(n10578), .ZN(n27691) );
  NOR2_X1 U6667 ( .A1(n16417), .A2(n12120), .ZN(n18778) );
  INV_X1 U8822 ( .I(n4259), .ZN(n17266) );
  NAND2_X1 U13643 ( .A1(n16522), .A2(n18774), .ZN(n26962) );
  NAND2_X1 U10104 ( .A1(n10669), .A2(n9296), .ZN(n10326) );
  INV_X1 U3688 ( .I(n17223), .ZN(n17224) );
  INV_X1 U985 ( .I(n18860), .ZN(n18532) );
  NAND2_X1 U24372 ( .A1(n30371), .A2(n785), .ZN(n18817) );
  INV_X1 U6712 ( .I(n18357), .ZN(n18895) );
  NAND2_X1 U8777 ( .A1(n10579), .A2(n2990), .ZN(n6457) );
  OAI21_X1 U24299 ( .A1(n18481), .A2(n18601), .B(n18602), .ZN(n18480) );
  AOI21_X1 U13783 ( .A1(n955), .A2(n16995), .B(n1184), .ZN(n5458) );
  NAND3_X1 U2233 ( .A1(n18332), .A2(n18489), .A3(n6256), .ZN(n18334) );
  NAND2_X1 U21122 ( .A1(n16249), .A2(n18822), .ZN(n13946) );
  NOR2_X1 U24356 ( .A1(n18730), .A2(n18846), .ZN(n18732) );
  NOR2_X1 U8787 ( .A1(n18759), .A2(n27940), .ZN(n18606) );
  NAND2_X1 U5189 ( .A1(n18532), .A2(n18588), .ZN(n17599) );
  NAND3_X1 U2237 ( .A1(n1659), .A2(n5700), .A3(n46), .ZN(n7319) );
  AOI22_X1 U16162 ( .A1(n16196), .A2(n18648), .B1(n18373), .B2(n18804), .ZN(
        n27237) );
  NOR2_X1 U10098 ( .A1(n14843), .A2(n11397), .ZN(n11396) );
  OAI21_X1 U10140 ( .A1(n28010), .A2(n959), .B(n27958), .ZN(n16018) );
  NOR2_X1 U5174 ( .A1(n18532), .A2(n18588), .ZN(n18739) );
  INV_X1 U10183 ( .I(n12120), .ZN(n18339) );
  INV_X1 U2682 ( .I(n10264), .ZN(n18750) );
  NAND2_X1 U9648 ( .A1(n18846), .A2(n18847), .ZN(n18410) );
  OAI21_X1 U8737 ( .A1(n6579), .A2(n18802), .B(n8395), .ZN(n4472) );
  AOI22_X1 U6899 ( .A1(n18340), .A2(n18339), .B1(n1430), .B2(n6215), .ZN(
        n26176) );
  OAI21_X1 U24206 ( .A1(n27129), .A2(n28987), .B(n18556), .ZN(n18329) );
  NOR2_X1 U7552 ( .A1(n11864), .A2(n18559), .ZN(n18330) );
  OAI21_X1 U2620 ( .A1(n17113), .A2(n12013), .B(n18808), .ZN(n2680) );
  NAND2_X1 U7562 ( .A1(n18812), .A2(n2990), .ZN(n2683) );
  NOR2_X1 U15208 ( .A1(n15136), .A2(n4008), .ZN(n18260) );
  BUF_X2 U1314 ( .I(n10579), .Z(n3429) );
  BUF_X2 U8491 ( .I(n19049), .Z(n28705) );
  AOI21_X1 U6670 ( .A1(n17360), .A2(n18587), .B(n18863), .ZN(n13025) );
  INV_X2 U3971 ( .I(n9677), .ZN(n13568) );
  NOR2_X1 U18050 ( .A1(n19011), .A2(n5119), .ZN(n7110) );
  INV_X1 U21515 ( .I(n14811), .ZN(n18426) );
  NAND2_X1 U19805 ( .A1(n9787), .A2(n19224), .ZN(n12505) );
  NAND2_X1 U5484 ( .A1(n1053), .A2(n31451), .ZN(n18454) );
  INV_X2 U22187 ( .I(n19048), .ZN(n16669) );
  INV_X1 U7495 ( .I(n16699), .ZN(n19334) );
  NAND2_X1 U15115 ( .A1(n13037), .A2(n13035), .ZN(n27131) );
  NOR2_X1 U21485 ( .A1(n13200), .A2(n19118), .ZN(n14424) );
  INV_X1 U22712 ( .I(n19033), .ZN(n4102) );
  NAND3_X1 U7477 ( .A1(n7435), .A2(n7434), .A3(n1047), .ZN(n7439) );
  AOI22_X1 U7450 ( .A1(n9424), .A2(n9423), .B1(n18068), .B2(n26830), .ZN(n9422) );
  BUF_X2 U5501 ( .I(n18980), .Z(n16740) );
  NOR3_X1 U16708 ( .A1(n18930), .A2(n16444), .A3(n1053), .ZN(n18284) );
  BUF_X2 U3973 ( .I(n2581), .Z(n26181) );
  AOI21_X1 U13526 ( .A1(n15074), .A2(n15073), .B(n17986), .ZN(n14259) );
  NAND3_X1 U5233 ( .A1(n19087), .A2(n19089), .A3(n1384), .ZN(n10868) );
  NOR2_X1 U21457 ( .A1(n19215), .A2(n2901), .ZN(n28132) );
  OAI21_X1 U900 ( .A1(n10013), .A2(n11080), .B(n4017), .ZN(n18910) );
  NOR2_X1 U5481 ( .A1(n19332), .A2(n8335), .ZN(n5162) );
  NOR2_X1 U7999 ( .A1(n19359), .A2(n19356), .ZN(n15629) );
  NAND2_X1 U19389 ( .A1(n1180), .A2(n19255), .ZN(n8910) );
  INV_X1 U5490 ( .I(n19080), .ZN(n19171) );
  NOR2_X1 U7509 ( .A1(n19116), .A2(n19330), .ZN(n3784) );
  INV_X1 U10330 ( .I(n19148), .ZN(n26554) );
  NAND3_X1 U12769 ( .A1(n3365), .A2(n745), .A3(n3360), .ZN(n1870) );
  AOI21_X1 U7489 ( .A1(n32064), .A2(n15120), .B(n16916), .ZN(n19162) );
  INV_X1 U9991 ( .I(n12996), .ZN(n5710) );
  INV_X1 U21998 ( .I(n12830), .ZN(n12567) );
  INV_X1 U5252 ( .I(n19128), .ZN(n15378) );
  INV_X1 U12039 ( .I(n11074), .ZN(n17678) );
  NAND2_X1 U5941 ( .A1(n12707), .A2(n16669), .ZN(n3822) );
  NAND2_X1 U21514 ( .A1(n16592), .A2(n16591), .ZN(n18268) );
  NAND3_X1 U5924 ( .A1(n18967), .A2(n11085), .A3(n19165), .ZN(n11800) );
  AOI21_X1 U20394 ( .A1(n19280), .A2(n32908), .B(n26830), .ZN(n19282) );
  NAND3_X1 U2876 ( .A1(n34005), .A2(n29715), .A3(n17311), .ZN(n19173) );
  OAI21_X1 U12044 ( .A1(n18983), .A2(n19128), .B(n18963), .ZN(n18966) );
  OAI21_X1 U15672 ( .A1(n764), .A2(n25985), .B(n9677), .ZN(n9709) );
  NOR2_X1 U15974 ( .A1(n1378), .A2(n29146), .ZN(n12532) );
  INV_X1 U6188 ( .I(n1180), .ZN(n26288) );
  OAI21_X1 U8621 ( .A1(n1382), .A2(n19004), .B(n19210), .ZN(n18942) );
  AOI22_X1 U12330 ( .A1(n13495), .A2(n19116), .B1(n879), .B2(n5162), .ZN(
        n28003) );
  INV_X1 U19512 ( .I(n19151), .ZN(n9176) );
  NAND3_X1 U18141 ( .A1(n16354), .A2(n19291), .A3(n7251), .ZN(n19204) );
  BUF_X2 U7668 ( .I(Key[160]), .Z(n25054) );
  INV_X1 U9966 ( .I(n16727), .ZN(n3076) );
  INV_X1 U2889 ( .I(n2073), .ZN(n2761) );
  INV_X1 U878 ( .I(n2483), .ZN(n6115) );
  BUF_X2 U4273 ( .I(Key[122]), .Z(n25358) );
  INV_X1 U11959 ( .I(n19644), .ZN(n1916) );
  BUF_X2 U6100 ( .I(Key[45]), .Z(n25783) );
  BUF_X2 U4278 ( .I(Key[99]), .Z(n25554) );
  INV_X1 U847 ( .I(n20067), .ZN(n823) );
  NAND2_X1 U4925 ( .A1(n823), .A2(n19947), .ZN(n28021) );
  INV_X2 U19508 ( .I(n10934), .ZN(n14210) );
  INV_X2 U8377 ( .I(n4060), .ZN(n5433) );
  INV_X1 U3238 ( .I(n577), .ZN(n1041) );
  INV_X2 U825 ( .I(n17688), .ZN(n20110) );
  INV_X1 U24625 ( .I(n29981), .ZN(n19976) );
  INV_X2 U5892 ( .I(n1164), .ZN(n7920) );
  INV_X2 U2496 ( .I(n16811), .ZN(n16812) );
  INV_X2 U837 ( .I(n29253), .ZN(n1036) );
  INV_X1 U863 ( .I(n26774), .ZN(n875) );
  OAI22_X1 U5347 ( .A1(n12038), .A2(n25997), .B1(n13747), .B2(n10947), .ZN(
        n17371) );
  INV_X1 U833 ( .I(n20109), .ZN(n20035) );
  INV_X1 U9941 ( .I(n16193), .ZN(n20012) );
  NAND2_X1 U16819 ( .A1(n5707), .A2(n19987), .ZN(n14440) );
  NAND2_X1 U7388 ( .A1(n3626), .A2(n20076), .ZN(n3663) );
  NAND2_X1 U5277 ( .A1(n12008), .A2(n10086), .ZN(n8946) );
  AOI21_X1 U11780 ( .A1(n19861), .A2(n7923), .B(n1164), .ZN(n7921) );
  INV_X2 U21988 ( .I(n19986), .ZN(n28219) );
  INV_X1 U20149 ( .I(n20134), .ZN(n20132) );
  INV_X1 U7424 ( .I(n3486), .ZN(n3530) );
  NAND2_X1 U11848 ( .A1(n16346), .A2(n17243), .ZN(n3128) );
  NOR2_X1 U8504 ( .A1(n9876), .A2(n8301), .ZN(n2933) );
  NOR3_X1 U13885 ( .A1(n20007), .A2(n20008), .A3(n20009), .ZN(n2930) );
  NAND2_X1 U5299 ( .A1(n1036), .A2(n31161), .ZN(n8033) );
  OAI21_X1 U8550 ( .A1(n5871), .A2(n5869), .B(n31468), .ZN(n3292) );
  INV_X1 U9937 ( .I(n4215), .ZN(n17389) );
  NAND2_X1 U20249 ( .A1(n584), .A2(n14559), .ZN(n11475) );
  NAND2_X1 U11804 ( .A1(n26088), .A2(n30794), .ZN(n5288) );
  NAND2_X1 U14929 ( .A1(n20132), .A2(n16461), .ZN(n5931) );
  NOR2_X1 U19858 ( .A1(n13987), .A2(n10241), .ZN(n13986) );
  NAND2_X1 U7385 ( .A1(n15278), .A2(n1166), .ZN(n20292) );
  AND2_X1 U5338 ( .A1(n10831), .A2(n33627), .Z(n19952) );
  NOR2_X1 U9898 ( .A1(n20154), .A2(n27097), .ZN(n16307) );
  NOR2_X1 U6528 ( .A1(n4215), .A2(n17243), .ZN(n12078) );
  AOI21_X1 U19422 ( .A1(n17243), .A2(n4233), .B(n4215), .ZN(n9139) );
  NAND3_X1 U14805 ( .A1(n20100), .A2(n12895), .A3(n19990), .ZN(n17035) );
  OAI21_X1 U819 ( .A1(n29281), .A2(n25997), .B(n12038), .ZN(n13954) );
  NAND2_X1 U5357 ( .A1(n19952), .A2(n19856), .ZN(n12194) );
  OAI21_X1 U11802 ( .A1(n32559), .A2(n13058), .B(n19823), .ZN(n10478) );
  NOR2_X1 U8529 ( .A1(n19884), .A2(n19886), .ZN(n19421) );
  NOR2_X1 U1348 ( .A1(n12408), .A2(n3626), .ZN(n27802) );
  NAND2_X1 U21532 ( .A1(n17785), .A2(n20010), .ZN(n17784) );
  INV_X1 U2404 ( .I(n20485), .ZN(n1346) );
  NAND2_X1 U806 ( .A1(n20006), .A2(n20078), .ZN(n13107) );
  NAND2_X1 U15780 ( .A1(n19998), .A2(n28219), .ZN(n4367) );
  NAND3_X1 U13038 ( .A1(n20100), .A2(n29216), .A3(n29944), .ZN(n20623) );
  AOI21_X1 U1310 ( .A1(n19986), .A2(n25997), .B(n11521), .ZN(n4368) );
  INV_X1 U21264 ( .I(n20312), .ZN(n20578) );
  INV_X2 U4594 ( .I(n20492), .ZN(n20494) );
  INV_X1 U1298 ( .I(n8374), .ZN(n20525) );
  INV_X2 U771 ( .I(n31504), .ZN(n12169) );
  NAND2_X1 U22617 ( .A1(n17947), .A2(n20485), .ZN(n17532) );
  NOR2_X1 U23017 ( .A1(n20268), .A2(n14863), .ZN(n20269) );
  INV_X1 U3325 ( .I(n9320), .ZN(n1028) );
  INV_X2 U1242 ( .I(n15027), .ZN(n27771) );
  NOR2_X1 U8444 ( .A1(n935), .A2(n29628), .ZN(n17414) );
  NAND2_X1 U19867 ( .A1(n27105), .A2(n30643), .ZN(n20347) );
  NAND2_X1 U3199 ( .A1(n20268), .A2(n5781), .ZN(n5670) );
  BUF_X2 U2892 ( .I(n20267), .Z(n266) );
  NAND2_X1 U6503 ( .A1(n9320), .A2(n14436), .ZN(n20257) );
  BUF_X2 U22722 ( .I(n14049), .Z(n28357) );
  INV_X2 U14587 ( .I(n5748), .ZN(n782) );
  NAND2_X1 U6504 ( .A1(n20268), .A2(n20210), .ZN(n5782) );
  NAND2_X1 U4830 ( .A1(n15169), .A2(n20590), .ZN(n28893) );
  INV_X2 U23091 ( .I(n2928), .ZN(n28414) );
  NOR2_X1 U11727 ( .A1(n12771), .A2(n9484), .ZN(n5061) );
  AOI21_X1 U16049 ( .A1(n30971), .A2(n31873), .B(n20379), .ZN(n20380) );
  NAND3_X1 U23485 ( .A1(n28893), .A2(n31967), .A3(n15824), .ZN(n28485) );
  NOR2_X1 U8414 ( .A1(n7978), .A2(n936), .ZN(n12873) );
  OAI21_X1 U16113 ( .A1(n20347), .A2(n26730), .B(n27225), .ZN(n27227) );
  INV_X1 U26129 ( .I(n17947), .ZN(n17896) );
  NAND2_X1 U24715 ( .A1(n1159), .A2(n30987), .ZN(n20475) );
  NOR2_X1 U13112 ( .A1(n31804), .A2(n31533), .ZN(n5993) );
  INV_X1 U9953 ( .I(n31471), .ZN(n1354) );
  INV_X1 U14535 ( .I(n3644), .ZN(n12407) );
  AOI21_X1 U22901 ( .A1(n15042), .A2(n15043), .B(n28840), .ZN(n15041) );
  OAI22_X1 U8390 ( .A1(n29972), .A2(n20426), .B1(n16146), .B2(n20427), .ZN(
        n1930) );
  NOR2_X1 U15874 ( .A1(n1354), .A2(n4468), .ZN(n4471) );
  NAND2_X1 U23867 ( .A1(n817), .A2(n31804), .ZN(n17270) );
  NAND3_X1 U12457 ( .A1(n1351), .A2(n11312), .A3(n1349), .ZN(n20407) );
  OAI21_X1 U24661 ( .A1(n20202), .A2(n20201), .B(n27887), .ZN(n20203) );
  NOR2_X1 U3535 ( .A1(n5003), .A2(n32504), .ZN(n20164) );
  NOR2_X1 U11737 ( .A1(n2965), .A2(n1159), .ZN(n2764) );
  INV_X1 U24658 ( .I(n20462), .ZN(n20187) );
  INV_X1 U9719 ( .I(n9303), .ZN(n20871) );
  INV_X1 U19160 ( .I(n20755), .ZN(n12674) );
  INV_X1 U2704 ( .I(n20939), .ZN(n21270) );
  NOR2_X1 U19708 ( .A1(n7007), .A2(n28190), .ZN(n6303) );
  INV_X2 U5115 ( .I(n21170), .ZN(n14803) );
  INV_X1 U9718 ( .I(n11733), .ZN(n1148) );
  INV_X1 U4754 ( .I(n34157), .ZN(n21167) );
  NOR2_X1 U8306 ( .A1(n21398), .A2(n32625), .ZN(n21206) );
  NOR2_X1 U6435 ( .A1(n5049), .A2(n29255), .ZN(n5047) );
  NOR2_X1 U21135 ( .A1(n21165), .A2(n14803), .ZN(n21086) );
  INV_X2 U7165 ( .I(n21428), .ZN(n21341) );
  INV_X1 U2645 ( .I(n2118), .ZN(n8267) );
  INV_X1 U11538 ( .I(n28190), .ZN(n13509) );
  NOR2_X1 U20930 ( .A1(n1334), .A2(n21270), .ZN(n12243) );
  NAND2_X1 U9698 ( .A1(n5141), .A2(n14168), .ZN(n21340) );
  NAND3_X1 U15904 ( .A1(n28502), .A2(n21079), .A3(n4518), .ZN(n20938) );
  INV_X1 U11542 ( .I(n15751), .ZN(n17093) );
  NOR2_X1 U7185 ( .A1(n17640), .A2(n3106), .ZN(n7378) );
  NOR2_X1 U8254 ( .A1(n6451), .A2(n1736), .ZN(n4569) );
  OAI21_X1 U14558 ( .A1(n11151), .A2(n27842), .B(n21217), .ZN(n11150) );
  NAND2_X1 U13282 ( .A1(n7196), .A2(n6520), .ZN(n2568) );
  NOR2_X1 U8383 ( .A1(n28502), .A2(n16933), .ZN(n16484) );
  CLKBUF_X2 U4751 ( .I(n21170), .Z(n26861) );
  NOR2_X1 U8287 ( .A1(n21212), .A2(n6408), .ZN(n18213) );
  INV_X1 U24830 ( .I(n31909), .ZN(n21093) );
  NAND2_X1 U5413 ( .A1(n21405), .A2(n4989), .ZN(n4988) );
  OAI22_X1 U8246 ( .A1(n20933), .A2(n21080), .B1(n21365), .B2(n21183), .ZN(
        n13265) );
  OAI21_X1 U632 ( .A1(n9454), .A2(n7822), .B(n17455), .ZN(n9453) );
  NAND2_X1 U16203 ( .A1(n8175), .A2(n21434), .ZN(n27249) );
  NOR2_X1 U9642 ( .A1(n20662), .A2(n4518), .ZN(n4283) );
  OAI21_X1 U7129 ( .A1(n8012), .A2(n16639), .B(n7526), .ZN(n21437) );
  NAND2_X1 U15029 ( .A1(n7123), .A2(n7120), .ZN(n5843) );
  NAND2_X1 U3913 ( .A1(n2575), .A2(n21849), .ZN(n26341) );
  NOR3_X1 U23415 ( .A1(n21408), .A2(n4119), .A3(n30755), .ZN(n15872) );
  AOI21_X1 U9593 ( .A1(n7148), .A2(n8604), .B(n8010), .ZN(n6427) );
  NOR2_X1 U1032 ( .A1(n13133), .A2(n1136), .ZN(n26175) );
  BUF_X2 U24342 ( .I(n21665), .Z(n28618) );
  NAND3_X1 U6368 ( .A1(n16577), .A2(n13133), .A3(n1312), .ZN(n21667) );
  INV_X2 U6399 ( .I(n21463), .ZN(n918) );
  AOI21_X1 U14233 ( .A1(n15813), .A2(n10401), .B(n11890), .ZN(n27053) );
  INV_X1 U597 ( .I(n28232), .ZN(n1328) );
  AOI21_X1 U24913 ( .A1(n21690), .A2(n21859), .B(n21857), .ZN(n21538) );
  NAND3_X1 U1016 ( .A1(n1328), .A2(n15772), .A3(n21811), .ZN(n8174) );
  NOR2_X1 U11968 ( .A1(n21709), .A2(n30441), .ZN(n27383) );
  NAND2_X1 U3649 ( .A1(n8276), .A2(n21707), .ZN(n9055) );
  NOR2_X1 U23200 ( .A1(n30885), .A2(n27635), .ZN(n17347) );
  NOR2_X1 U1015 ( .A1(n21629), .A2(n21628), .ZN(n27991) );
  NOR2_X1 U11957 ( .A1(n31954), .A2(n27178), .ZN(n26731) );
  BUF_X2 U8183 ( .I(n8602), .Z(n4331) );
  INV_X2 U8196 ( .I(n21779), .ZN(n21781) );
  INV_X1 U3251 ( .I(n6489), .ZN(n21853) );
  NOR2_X1 U557 ( .A1(n21806), .A2(n6483), .ZN(n279) );
  NAND2_X1 U11404 ( .A1(n21690), .A2(n29523), .ZN(n2708) );
  NAND2_X1 U11337 ( .A1(n21164), .A2(n16577), .ZN(n12994) );
  INV_X1 U3590 ( .I(n21715), .ZN(n911) );
  INV_X1 U4165 ( .I(n14095), .ZN(n21775) );
  INV_X1 U4633 ( .I(n7502), .ZN(n28665) );
  NOR2_X1 U22789 ( .A1(n30440), .A2(n31309), .ZN(n21934) );
  NAND3_X1 U940 ( .A1(n17644), .A2(n3756), .A3(n21857), .ZN(n28159) );
  NAND3_X1 U9505 ( .A1(n21800), .A2(n21801), .A3(n21799), .ZN(n15640) );
  NAND2_X1 U18456 ( .A1(n21678), .A2(n28203), .ZN(n27630) );
  OAI21_X1 U23082 ( .A1(n17472), .A2(n15026), .B(n16194), .ZN(n21495) );
  AOI21_X1 U11322 ( .A1(n12102), .A2(n21686), .B(n26513), .ZN(n10490) );
  NAND2_X1 U3432 ( .A1(n9119), .A2(n21655), .ZN(n21936) );
  NAND2_X1 U21170 ( .A1(n15091), .A2(n31085), .ZN(n14012) );
  NOR2_X1 U5396 ( .A1(n21622), .A2(n28387), .ZN(n21561) );
  NAND2_X1 U13782 ( .A1(n10028), .A2(n27619), .ZN(n26979) );
  NOR2_X1 U11282 ( .A1(n17164), .A2(n15319), .ZN(n16164) );
  OAI21_X1 U13910 ( .A1(n12626), .A2(n9076), .B(n11619), .ZN(n9088) );
  NAND2_X1 U3902 ( .A1(n21819), .A2(n26904), .ZN(n27103) );
  AOI21_X1 U9515 ( .A1(n9666), .A2(n15091), .B(n28618), .ZN(n13804) );
  NAND2_X1 U22785 ( .A1(n21934), .A2(n915), .ZN(n21935) );
  INV_X1 U524 ( .I(n22172), .ZN(n4723) );
  INV_X1 U4839 ( .I(n32055), .ZN(n9065) );
  INV_X1 U6356 ( .I(n11100), .ZN(n22543) );
  NAND2_X1 U6318 ( .A1(n1122), .A2(n31931), .ZN(n11575) );
  INV_X2 U2572 ( .I(n22543), .ZN(n1124) );
  NAND2_X1 U23842 ( .A1(n28472), .A2(n16627), .ZN(n22571) );
  NAND2_X1 U21002 ( .A1(n15752), .A2(n29451), .ZN(n15008) );
  OAI21_X1 U8027 ( .A1(n4055), .A2(n4054), .B(n8527), .ZN(n7610) );
  NOR2_X1 U9350 ( .A1(n18098), .A2(n12076), .ZN(n17263) );
  NAND2_X1 U20086 ( .A1(n22330), .A2(n14376), .ZN(n10317) );
  NOR2_X1 U782 ( .A1(n998), .A2(n22330), .ZN(n17132) );
  INV_X2 U3597 ( .I(n22626), .ZN(n1117) );
  INV_X1 U4141 ( .I(n8409), .ZN(n22586) );
  INV_X1 U4132 ( .I(n30668), .ZN(n1282) );
  INV_X2 U492 ( .I(n16205), .ZN(n22689) );
  OAI21_X1 U25106 ( .A1(n22565), .A2(n22561), .B(n22560), .ZN(n22566) );
  NAND2_X1 U430 ( .A1(n15229), .A2(n22476), .ZN(n13534) );
  NAND3_X1 U724 ( .A1(n26878), .A2(n27378), .A3(n996), .ZN(n26178) );
  OAI21_X1 U17275 ( .A1(n22610), .A2(n29336), .B(n22631), .ZN(n22613) );
  NOR2_X1 U8005 ( .A1(n22531), .A2(n9234), .ZN(n9777) );
  NOR2_X1 U18681 ( .A1(n7957), .A2(n1124), .ZN(n8136) );
  OAI21_X1 U21232 ( .A1(n17960), .A2(n16375), .B(n1728), .ZN(n22526) );
  INV_X1 U9386 ( .I(n9272), .ZN(n8348) );
  NOR2_X1 U2334 ( .A1(n16170), .A2(n25), .ZN(n26862) );
  NAND2_X1 U11069 ( .A1(n1113), .A2(n22923), .ZN(n3854) );
  NAND2_X1 U21922 ( .A1(n1294), .A2(n26884), .ZN(n28206) );
  NAND2_X1 U9438 ( .A1(n9271), .A2(n9234), .ZN(n9270) );
  OAI22_X1 U19882 ( .A1(n13417), .A2(n9913), .B1(n22667), .B2(n29078), .ZN(
        n22723) );
  INV_X2 U14894 ( .I(n4908), .ZN(n724) );
  OAI21_X1 U6546 ( .A1(n26144), .A2(n26660), .B(n14728), .ZN(n26394) );
  AOI21_X1 U9367 ( .A1(n8595), .A2(n30641), .B(n4300), .ZN(n4299) );
  NAND2_X1 U4529 ( .A1(n22392), .A2(n22546), .ZN(n14024) );
  NAND2_X1 U1044 ( .A1(n22407), .A2(n22429), .ZN(n17627) );
  INV_X1 U15007 ( .I(n23072), .ZN(n8683) );
  NOR2_X1 U6949 ( .A1(n22878), .A2(n31437), .ZN(n2169) );
  NOR2_X1 U9236 ( .A1(n14131), .A2(n2635), .ZN(n6285) );
  INV_X1 U9322 ( .I(n6798), .ZN(n1107) );
  INV_X1 U590 ( .I(n31637), .ZN(n13778) );
  INV_X2 U7972 ( .I(n849), .ZN(n7181) );
  INV_X1 U6287 ( .I(n5915), .ZN(n23073) );
  INV_X1 U615 ( .I(n22968), .ZN(n23083) );
  NOR2_X1 U16802 ( .A1(n27622), .A2(n3163), .ZN(n13917) );
  NAND3_X1 U25193 ( .A1(n23070), .A2(n10641), .A3(n23069), .ZN(n23071) );
  NOR2_X1 U6261 ( .A1(n26724), .A2(n23104), .ZN(n5972) );
  OAI21_X1 U21545 ( .A1(n18241), .A2(n22916), .B(n27090), .ZN(n18047) );
  INV_X1 U4409 ( .I(n28214), .ZN(n27409) );
  NOR2_X1 U26084 ( .A1(n22798), .A2(n23053), .ZN(n23050) );
  NAND2_X1 U1427 ( .A1(n641), .A2(n11268), .ZN(n6227) );
  NAND2_X1 U16265 ( .A1(n32091), .A2(n10296), .ZN(n22441) );
  NAND3_X1 U19331 ( .A1(n15852), .A2(n15851), .A3(n30960), .ZN(n13598) );
  NOR2_X1 U22109 ( .A1(n22872), .A2(n31861), .ZN(n12824) );
  OAI22_X1 U14459 ( .A1(n10360), .A2(n3570), .B1(n3891), .B2(n12586), .ZN(
        n22714) );
  INV_X1 U10853 ( .I(n15941), .ZN(n2974) );
  INV_X1 U10860 ( .I(n12716), .ZN(n3282) );
  INV_X1 U312 ( .I(n23475), .ZN(n6262) );
  INV_X1 U458 ( .I(n28811), .ZN(n662) );
  OAI21_X1 U9134 ( .A1(n11887), .A2(n11933), .B(n3004), .ZN(n10069) );
  INV_X1 U7887 ( .I(n23719), .ZN(n23919) );
  INV_X1 U6218 ( .I(n23567), .ZN(n23849) );
  INV_X1 U8286 ( .I(n23683), .ZN(n23681) );
  NAND2_X1 U25891 ( .A1(n32998), .A2(n11933), .ZN(n15490) );
  NAND2_X1 U5789 ( .A1(n23491), .A2(n23712), .ZN(n17520) );
  INV_X1 U477 ( .I(n10954), .ZN(n11968) );
  OR2_X1 U2850 ( .A1(n28611), .A2(n8166), .Z(n8674) );
  NOR2_X1 U5695 ( .A1(n23713), .A2(n23889), .ZN(n23842) );
  INV_X2 U413 ( .I(n756), .ZN(n28510) );
  NAND2_X1 U10532 ( .A1(n23813), .A2(n663), .ZN(n23692) );
  INV_X2 U9216 ( .I(n27455), .ZN(n23752) );
  INV_X1 U9199 ( .I(n11567), .ZN(n8095) );
  INV_X1 U4113 ( .I(n9430), .ZN(n15912) );
  AND2_X1 U19075 ( .A1(n7022), .A2(n2839), .Z(n14092) );
  NOR2_X1 U20458 ( .A1(n23864), .A2(n23527), .ZN(n11131) );
  NAND2_X1 U7815 ( .A1(n23894), .A2(n29068), .ZN(n6249) );
  NAND2_X1 U9180 ( .A1(n7915), .A2(n23778), .ZN(n11393) );
  INV_X1 U25320 ( .I(n23646), .ZN(n23647) );
  NOR2_X1 U3881 ( .A1(n707), .A2(n8370), .ZN(n655) );
  AOI21_X1 U18362 ( .A1(n10193), .A2(n34008), .B(n23897), .ZN(n10560) );
  NAND2_X1 U5831 ( .A1(n17520), .A2(n17234), .ZN(n11491) );
  INV_X1 U5711 ( .I(n976), .ZN(n1249) );
  NOR2_X1 U10819 ( .A1(n13549), .A2(n27219), .ZN(n8473) );
  NOR2_X1 U6856 ( .A1(n8544), .A2(n14207), .ZN(n11309) );
  INV_X2 U404 ( .I(n15423), .ZN(n23850) );
  NAND2_X1 U9139 ( .A1(n978), .A2(n8273), .ZN(n15351) );
  INV_X1 U4790 ( .I(n14092), .ZN(n23651) );
  OAI21_X1 U2110 ( .A1(n13544), .A2(n13578), .B(n17906), .ZN(n7613) );
  NAND2_X1 U25328 ( .A1(n11192), .A2(n16337), .ZN(n28744) );
  NAND3_X1 U6895 ( .A1(n16467), .A2(n846), .A3(n27219), .ZN(n7075) );
  NAND3_X1 U16858 ( .A1(n847), .A2(n23573), .A3(n5759), .ZN(n23574) );
  NAND2_X1 U21319 ( .A1(n23832), .A2(n23912), .ZN(n17398) );
  NOR2_X1 U21050 ( .A1(n8408), .A2(n17895), .ZN(n17806) );
  NAND2_X1 U2242 ( .A1(n32711), .A2(n654), .ZN(n26384) );
  INV_X1 U21292 ( .I(n23923), .ZN(n16118) );
  INV_X1 U375 ( .I(n32308), .ZN(n26383) );
  INV_X1 U8694 ( .I(n26392), .ZN(n26391) );
  NOR2_X1 U348 ( .A1(n9797), .A2(n14207), .ZN(n9769) );
  NAND2_X1 U10741 ( .A1(n17618), .A2(n13503), .ZN(n3484) );
  NOR2_X1 U24025 ( .A1(n17807), .A2(n17806), .ZN(n17805) );
  INV_X1 U1627 ( .I(n9919), .ZN(n10530) );
  INV_X1 U218 ( .I(n6911), .ZN(n24312) );
  CLKBUF_X2 U3087 ( .I(n24299), .Z(n319) );
  BUF_X2 U26435 ( .I(n24314), .Z(n7503) );
  INV_X2 U6831 ( .I(n3205), .ZN(n9323) );
  INV_X1 U204 ( .I(n5199), .ZN(n24245) );
  INV_X1 U1655 ( .I(n9342), .ZN(n14252) );
  INV_X1 U9113 ( .I(n16799), .ZN(n1089) );
  NAND2_X1 U8289 ( .A1(n24243), .A2(n24242), .ZN(n1480) );
  NAND2_X1 U8049 ( .A1(n1089), .A2(n14619), .ZN(n5615) );
  AOI21_X1 U9049 ( .A1(n796), .A2(n10226), .B(n970), .ZN(n9282) );
  NOR2_X1 U20904 ( .A1(n24305), .A2(n24197), .ZN(n16901) );
  NAND2_X1 U2309 ( .A1(n27159), .A2(n24094), .ZN(n13239) );
  NOR2_X1 U9043 ( .A1(n16985), .A2(n1245), .ZN(n5616) );
  INV_X1 U4097 ( .I(n14725), .ZN(n27550) );
  INV_X1 U15179 ( .I(n3148), .ZN(n3038) );
  NAND2_X1 U9027 ( .A1(n24061), .A2(n10651), .ZN(n11342) );
  NOR2_X1 U4777 ( .A1(n3483), .A2(n24193), .ZN(n24057) );
  NAND2_X1 U3528 ( .A1(n27117), .A2(n24168), .ZN(n13306) );
  NOR2_X1 U4779 ( .A1(n10033), .A2(n24201), .ZN(n7669) );
  OAI21_X1 U14171 ( .A1(n7809), .A2(n30280), .B(n16651), .ZN(n5937) );
  NAND3_X1 U5263 ( .A1(n24211), .A2(n24213), .A3(n24209), .ZN(n6990) );
  NAND3_X1 U8171 ( .A1(n24322), .A2(n29785), .A3(n24209), .ZN(n6817) );
  NAND2_X1 U10544 ( .A1(n28120), .A2(n13048), .ZN(n13046) );
  INV_X1 U10615 ( .I(n11346), .ZN(n10428) );
  NOR2_X1 U15680 ( .A1(n24097), .A2(n24096), .ZN(n5377) );
  NOR2_X1 U7785 ( .A1(n14443), .A2(n17404), .ZN(n7105) );
  OAI21_X1 U2256 ( .A1(n32036), .A2(n7669), .B(n24008), .ZN(n7668) );
  NAND2_X1 U7810 ( .A1(n8058), .A2(n24106), .ZN(n23665) );
  NAND2_X1 U3284 ( .A1(n11342), .A2(n11341), .ZN(n11340) );
  NAND2_X1 U14084 ( .A1(n6001), .A2(n27026), .ZN(n12693) );
  NAND3_X1 U18424 ( .A1(n1244), .A2(n29010), .A3(n24216), .ZN(n10175) );
  NAND2_X1 U23247 ( .A1(n23748), .A2(n27184), .ZN(n24018) );
  NAND2_X1 U9069 ( .A1(n10188), .A2(n31355), .ZN(n8000) );
  NAND3_X1 U3711 ( .A1(n24322), .A2(n13268), .A3(n29785), .ZN(n24324) );
  NAND2_X1 U25404 ( .A1(n24213), .A2(n13268), .ZN(n24214) );
  NAND2_X1 U1058 ( .A1(n2852), .A2(n29567), .ZN(n2849) );
  AOI21_X1 U11550 ( .A1(n14336), .A2(n24317), .B(n32298), .ZN(n2156) );
  NAND3_X1 U22969 ( .A1(n1089), .A2(n12054), .A3(n14745), .ZN(n15224) );
  INV_X1 U10526 ( .I(n24442), .ZN(n10070) );
  OR2_X1 U173 ( .A1(n6877), .A2(n4207), .Z(n27153) );
  INV_X1 U9015 ( .I(n24839), .ZN(n3233) );
  INV_X1 U21655 ( .I(n24522), .ZN(n24658) );
  INV_X1 U6784 ( .I(n16319), .ZN(n7466) );
  INV_X1 U3744 ( .I(n13695), .ZN(n24642) );
  BUF_X2 U3027 ( .I(n25308), .Z(n25962) );
  NOR2_X1 U17370 ( .A1(n7413), .A2(n24607), .ZN(n6326) );
  NOR2_X1 U2117 ( .A1(n13532), .A2(n16397), .ZN(n6691) );
  NAND2_X1 U8419 ( .A1(n15719), .A2(n24874), .ZN(n27926) );
  INV_X2 U2261 ( .I(n12676), .ZN(n24725) );
  INV_X1 U19329 ( .I(n4885), .ZN(n18264) );
  INV_X1 U4424 ( .I(n25012), .ZN(n17684) );
  AOI21_X1 U16251 ( .A1(n13050), .A2(n25872), .B(n884), .ZN(n4931) );
  NAND2_X1 U4393 ( .A1(n16729), .A2(n16276), .ZN(n16728) );
  NAND2_X1 U26368 ( .A1(n4885), .A2(n32760), .ZN(n11953) );
  NOR2_X1 U25363 ( .A1(n4318), .A2(n25871), .ZN(n23960) );
  NOR2_X1 U4731 ( .A1(n13985), .A2(n18059), .ZN(n5793) );
  NOR2_X1 U2316 ( .A1(n717), .A2(n25756), .ZN(n3275) );
  OAI21_X1 U12928 ( .A1(n12086), .A2(n12926), .B(n718), .ZN(n3885) );
  INV_X1 U15073 ( .I(n1221), .ZN(n27128) );
  NAND2_X1 U7762 ( .A1(n2967), .A2(n26270), .ZN(n24413) );
  NOR2_X1 U19613 ( .A1(n27862), .A2(n27861), .ZN(n28875) );
  INV_X1 U52 ( .I(n25712), .ZN(n12314) );
  NAND2_X1 U10317 ( .A1(n2536), .A2(n30288), .ZN(n10359) );
  INV_X1 U5554 ( .I(n25664), .ZN(n25659) );
  INV_X1 U2146 ( .I(n24970), .ZN(n29049) );
  INV_X2 U9260 ( .I(n25689), .ZN(n26447) );
  INV_X1 U25541 ( .I(n24956), .ZN(n24938) );
  INV_X1 U25495 ( .I(n25490), .ZN(n25475) );
  INV_X1 U6035 ( .I(n12611), .ZN(n12309) );
  OAI21_X1 U23695 ( .A1(n8676), .A2(n16670), .B(n12611), .ZN(n25793) );
  OR2_X1 U1 ( .A1(n14208), .A2(n964), .Z(n9902) );
  NAND2_X1 U9 ( .A1(n25474), .A2(n25475), .ZN(n30118) );
  NAND3_X1 U11 ( .A1(n31647), .A2(n8320), .A3(n13483), .ZN(n30134) );
  NAND3_X1 U12 ( .A1(n14944), .A2(n15134), .A3(n31236), .ZN(n8804) );
  OR2_X1 U13 ( .A1(n27164), .A2(n1597), .Z(n7040) );
  OR2_X1 U15 ( .A1(n8515), .A2(n9956), .Z(n30330) );
  NOR2_X1 U34 ( .A1(n28070), .A2(n25060), .ZN(n17728) );
  INV_X1 U43 ( .I(n25214), .ZN(n25220) );
  INV_X1 U58 ( .I(n25665), .ZN(n25658) );
  OAI21_X1 U90 ( .A1(n31602), .A2(n31603), .B(n33278), .ZN(n29911) );
  NOR2_X1 U124 ( .A1(n32571), .A2(n1212), .ZN(n30876) );
  NOR2_X1 U127 ( .A1(n17781), .A2(n11945), .ZN(n31603) );
  INV_X1 U131 ( .I(n24471), .ZN(n30461) );
  NAND2_X1 U133 ( .A1(n14959), .A2(n25012), .ZN(n30145) );
  NOR2_X1 U135 ( .A1(n884), .A2(n13042), .ZN(n31463) );
  OR2_X1 U137 ( .A1(n25892), .A2(n25890), .Z(n14042) );
  NOR2_X1 U139 ( .A1(n883), .A2(n25885), .ZN(n4930) );
  NOR2_X1 U158 ( .A1(n24725), .A2(n13050), .ZN(n31464) );
  OAI21_X1 U163 ( .A1(n30998), .A2(n6691), .B(n837), .ZN(n30386) );
  INV_X2 U164 ( .I(n547), .ZN(n14268) );
  OR2_X1 U170 ( .A1(n5897), .A2(n14454), .Z(n29351) );
  NOR2_X1 U171 ( .A1(n14055), .A2(n15318), .ZN(n14484) );
  NAND2_X1 U213 ( .A1(n25900), .A2(n25897), .ZN(n24461) );
  INV_X1 U231 ( .I(n25700), .ZN(n3565) );
  CLKBUF_X2 U240 ( .I(n25023), .Z(n8210) );
  INV_X1 U268 ( .I(n24531), .ZN(n29589) );
  NAND3_X1 U295 ( .A1(n24124), .A2(n24182), .A3(n11463), .ZN(n13204) );
  NAND2_X1 U303 ( .A1(n12312), .A2(n6001), .ZN(n29502) );
  NAND2_X1 U316 ( .A1(n24162), .A2(n14592), .ZN(n16859) );
  CLKBUF_X1 U319 ( .I(n4151), .Z(n27500) );
  NAND3_X1 U329 ( .A1(n17588), .A2(n1232), .A3(n17589), .ZN(n17587) );
  NOR2_X1 U335 ( .A1(n24039), .A2(n6001), .ZN(n31016) );
  OR2_X1 U356 ( .A1(n2444), .A2(n13175), .Z(n10859) );
  NAND2_X1 U357 ( .A1(n26314), .A2(n839), .ZN(n5366) );
  CLKBUF_X2 U369 ( .I(n15536), .Z(n29306) );
  AND2_X1 U373 ( .A1(n1244), .A2(n24289), .Z(n29293) );
  NAND2_X1 U383 ( .A1(n14252), .A2(n319), .ZN(n29512) );
  INV_X1 U395 ( .I(n24314), .ZN(n10033) );
  NAND2_X1 U406 ( .A1(n28350), .A2(n9214), .ZN(n30280) );
  CLKBUF_X2 U407 ( .I(n14619), .Z(n31883) );
  CLKBUF_X1 U408 ( .I(n14335), .Z(n31271) );
  NAND2_X1 U411 ( .A1(n28210), .A2(n23880), .ZN(n23709) );
  NAND2_X1 U424 ( .A1(n7993), .A2(n30251), .ZN(n664) );
  OAI21_X1 U426 ( .A1(n11131), .A2(n15446), .B(n23932), .ZN(n30898) );
  OAI21_X1 U455 ( .A1(n27678), .A2(n23867), .B(n10142), .ZN(n17807) );
  OAI21_X1 U461 ( .A1(n14513), .A2(n29590), .B(n5417), .ZN(n14990) );
  AND2_X1 U490 ( .A1(n23904), .A2(n23905), .Z(n17287) );
  NAND3_X1 U496 ( .A1(n26074), .A2(n23721), .A3(n15095), .ZN(n28194) );
  NAND2_X1 U497 ( .A1(n31696), .A2(n739), .ZN(n25954) );
  INV_X1 U503 ( .I(n23590), .ZN(n14746) );
  NOR2_X1 U514 ( .A1(n14975), .A2(n12680), .ZN(n30620) );
  INV_X1 U521 ( .I(n17694), .ZN(n31175) );
  OAI21_X1 U523 ( .A1(n16786), .A2(n14297), .B(n23852), .ZN(n29682) );
  OR2_X1 U543 ( .A1(n23720), .A2(n23719), .Z(n23510) );
  NOR2_X1 U568 ( .A1(n23887), .A2(n23840), .ZN(n23632) );
  NOR2_X1 U570 ( .A1(n29240), .A2(n23713), .ZN(n31158) );
  INV_X1 U588 ( .I(n23720), .ZN(n23917) );
  AOI22_X1 U605 ( .A1(n3173), .A2(n23100), .B1(n3174), .B2(n986), .ZN(n3172)
         );
  AND2_X1 U622 ( .A1(n30231), .A2(n16280), .Z(n16975) );
  NAND2_X1 U629 ( .A1(n5874), .A2(n23111), .ZN(n30123) );
  AND2_X1 U638 ( .A1(n22832), .A2(n31943), .Z(n17064) );
  NOR2_X1 U646 ( .A1(n17828), .A2(n31549), .ZN(n31548) );
  NOR3_X1 U647 ( .A1(n28957), .A2(n28801), .A3(n22748), .ZN(n30247) );
  NAND2_X1 U651 ( .A1(n23083), .A2(n7802), .ZN(n23084) );
  NAND2_X1 U664 ( .A1(n16254), .A2(n30476), .ZN(n27834) );
  OAI21_X1 U675 ( .A1(n15039), .A2(n32119), .B(n33675), .ZN(n5619) );
  OAI22_X1 U700 ( .A1(n22761), .A2(n641), .B1(n15704), .B2(n15301), .ZN(n10404) );
  CLKBUF_X2 U719 ( .I(n26898), .Z(n30976) );
  NOR2_X1 U733 ( .A1(n3163), .A2(n29317), .ZN(n23074) );
  NAND2_X2 U786 ( .A1(n30762), .A2(n30349), .ZN(n31637) );
  OR2_X1 U790 ( .A1(n22587), .A2(n1125), .Z(n29406) );
  OR2_X1 U791 ( .A1(n13710), .A2(n15089), .Z(n12019) );
  NAND3_X1 U808 ( .A1(n31559), .A2(n22646), .A3(n4459), .ZN(n9156) );
  NAND3_X1 U844 ( .A1(n858), .A2(n22670), .A3(n29495), .ZN(n1516) );
  NAND2_X1 U860 ( .A1(n22681), .A2(n10354), .ZN(n17569) );
  NAND2_X1 U873 ( .A1(n22647), .A2(n5961), .ZN(n31559) );
  NOR2_X1 U887 ( .A1(n18062), .A2(n22651), .ZN(n29583) );
  NOR2_X1 U892 ( .A1(n17960), .A2(n22524), .ZN(n26144) );
  OR2_X1 U911 ( .A1(n11895), .A2(n32532), .Z(n22200) );
  NOR3_X1 U916 ( .A1(n5769), .A2(n355), .A3(n31931), .ZN(n28661) );
  AOI21_X1 U917 ( .A1(n1000), .A2(n22681), .B(n10282), .ZN(n17269) );
  OAI21_X1 U925 ( .A1(n6257), .A2(n28424), .B(n29342), .ZN(n31363) );
  OR2_X1 U928 ( .A1(n16277), .A2(n13704), .Z(n22648) );
  AND2_X1 U932 ( .A1(n22670), .A2(n1127), .Z(n29371) );
  AND2_X1 U933 ( .A1(n22636), .A2(n12043), .Z(n29355) );
  NAND2_X1 U937 ( .A1(n10725), .A2(n22645), .ZN(n29562) );
  NAND2_X1 U939 ( .A1(n31838), .A2(n11083), .ZN(n118) );
  AND2_X1 U941 ( .A1(n15089), .A2(n32172), .Z(n12556) );
  INV_X1 U949 ( .I(n22670), .ZN(n30106) );
  NOR2_X1 U957 ( .A1(n17960), .A2(n1728), .ZN(n15033) );
  NAND2_X1 U989 ( .A1(n10622), .A2(n10568), .ZN(n9752) );
  BUF_X2 U1020 ( .I(n11907), .Z(n29304) );
  INV_X1 U1037 ( .I(n22232), .ZN(n2863) );
  INV_X1 U1041 ( .I(n3704), .ZN(n30087) );
  INV_X1 U1045 ( .I(n3634), .ZN(n26863) );
  INV_X1 U1047 ( .I(n22227), .ZN(n30747) );
  OAI21_X1 U1068 ( .A1(n10215), .A2(n11081), .B(n21673), .ZN(n17681) );
  AND2_X1 U1071 ( .A1(n21465), .A2(n1134), .Z(n29455) );
  AOI21_X1 U1073 ( .A1(n31511), .A2(n21786), .B(n1323), .ZN(n4687) );
  NAND2_X1 U1078 ( .A1(n15091), .A2(n21581), .ZN(n31089) );
  AND2_X1 U1084 ( .A1(n2575), .A2(n16023), .Z(n29435) );
  AND2_X1 U1095 ( .A1(n32252), .A2(n27635), .Z(n29407) );
  AND2_X1 U1096 ( .A1(n17098), .A2(n21463), .Z(n10215) );
  NOR2_X1 U1098 ( .A1(n17472), .A2(n29302), .ZN(n10028) );
  NAND3_X1 U1114 ( .A1(n861), .A2(n21687), .A3(n21688), .ZN(n31121) );
  AND2_X1 U1116 ( .A1(n30506), .A2(n28429), .Z(n12279) );
  NOR2_X1 U1118 ( .A1(n21717), .A2(n26710), .ZN(n7986) );
  NOR2_X1 U1130 ( .A1(n21645), .A2(n21646), .ZN(n21091) );
  NAND2_X1 U1134 ( .A1(n11861), .A2(n21583), .ZN(n3588) );
  OR2_X1 U1137 ( .A1(n21687), .A2(n21688), .Z(n12102) );
  NOR2_X1 U1138 ( .A1(n28729), .A2(n12394), .ZN(n29796) );
  AOI22_X1 U1144 ( .A1(n1008), .A2(n8313), .B1(n21799), .B2(n21797), .ZN(
        n31026) );
  NAND2_X1 U1174 ( .A1(n30326), .A2(n21553), .ZN(n21678) );
  NAND2_X1 U1175 ( .A1(n21716), .A2(n21715), .ZN(n7276) );
  OR2_X1 U1186 ( .A1(n5170), .A2(n9999), .Z(n2337) );
  OR2_X1 U1200 ( .A1(n29258), .A2(n1652), .Z(n11796) );
  NOR3_X1 U1208 ( .A1(n27560), .A2(n29854), .A3(n21730), .ZN(n29943) );
  INV_X1 U1224 ( .I(n9666), .ZN(n11729) );
  NAND2_X1 U1226 ( .A1(n21755), .A2(n26451), .ZN(n30902) );
  OR2_X1 U1229 ( .A1(n26445), .A2(n27336), .Z(n16864) );
  NOR2_X1 U1232 ( .A1(n31511), .A2(n21786), .ZN(n11938) );
  NOR2_X1 U1278 ( .A1(n27563), .A2(n29777), .ZN(n21509) );
  NAND2_X1 U1289 ( .A1(n12340), .A2(n21183), .ZN(n30700) );
  NOR2_X1 U1290 ( .A1(n10921), .A2(n21127), .ZN(n31677) );
  OAI21_X1 U1306 ( .A1(n21396), .A2(n27955), .B(n3933), .ZN(n31815) );
  NOR2_X1 U1308 ( .A1(n21306), .A2(n21303), .ZN(n30544) );
  NAND2_X1 U1334 ( .A1(n3933), .A2(n29303), .ZN(n21286) );
  INV_X1 U1337 ( .I(n21506), .ZN(n29777) );
  INV_X1 U1340 ( .I(n4683), .ZN(n728) );
  NAND2_X1 U1341 ( .A1(n16639), .A2(n320), .ZN(n7526) );
  NOR2_X1 U1393 ( .A1(n28037), .A2(n21253), .ZN(n15932) );
  OR2_X1 U1399 ( .A1(n31614), .A2(n349), .Z(n31613) );
  NOR2_X1 U1400 ( .A1(n11734), .A2(n1148), .ZN(n30863) );
  AOI21_X1 U1406 ( .A1(n11187), .A2(n21189), .B(n2822), .ZN(n14023) );
  OR2_X1 U1407 ( .A1(n21442), .A2(n21100), .Z(n21304) );
  OAI21_X1 U1414 ( .A1(n21307), .A2(n21443), .B(n21306), .ZN(n21308) );
  INV_X1 U1428 ( .I(n21270), .ZN(n31476) );
  CLKBUF_X2 U1485 ( .I(n21356), .Z(n28701) );
  BUF_X2 U1486 ( .I(n21165), .Z(n27075) );
  OR2_X1 U1498 ( .A1(n9405), .A2(n9626), .Z(n31004) );
  BUF_X2 U1499 ( .I(n21432), .Z(n320) );
  INV_X1 U1515 ( .I(n13092), .ZN(n30543) );
  NAND3_X1 U1533 ( .A1(n10765), .A2(n8797), .A3(n10764), .ZN(n31608) );
  INV_X1 U1534 ( .I(n6500), .ZN(n30430) );
  OR2_X1 U1535 ( .A1(n14177), .A2(n32329), .Z(n7956) );
  NAND3_X1 U1560 ( .A1(n16004), .A2(n9688), .A3(n8087), .ZN(n30197) );
  NAND2_X1 U1561 ( .A1(n3644), .A2(n31047), .ZN(n5413) );
  NAND2_X1 U1563 ( .A1(n16132), .A2(n20523), .ZN(n30414) );
  INV_X1 U1600 ( .I(n31211), .ZN(n31210) );
  OR2_X1 U1626 ( .A1(n20471), .A2(n29337), .Z(n2766) );
  NAND2_X1 U1635 ( .A1(n30425), .A2(n32504), .ZN(n2767) );
  INV_X1 U1642 ( .I(n20537), .ZN(n31250) );
  OAI22_X1 U1645 ( .A1(n20528), .A2(n13499), .B1(n13599), .B2(n11984), .ZN(
        n31022) );
  NOR2_X1 U1646 ( .A1(n8206), .A2(n27771), .ZN(n30471) );
  NOR2_X1 U1650 ( .A1(n28626), .A2(n741), .ZN(n29724) );
  OAI21_X1 U1654 ( .A1(n2879), .A2(n14187), .B(n33530), .ZN(n7867) );
  NAND2_X1 U1684 ( .A1(n7242), .A2(n6530), .ZN(n15833) );
  CLKBUF_X2 U1687 ( .I(n2928), .Z(n31804) );
  NAND2_X1 U1691 ( .A1(n8770), .A2(n14436), .ZN(n3787) );
  NAND3_X1 U1693 ( .A1(n31721), .A2(n13759), .A3(n20310), .ZN(n29983) );
  BUF_X2 U1708 ( .I(n20384), .Z(n30594) );
  INV_X1 U1711 ( .I(n20345), .ZN(n30138) );
  NOR2_X1 U1715 ( .A1(n20463), .A2(n20371), .ZN(n20464) );
  BUF_X2 U1729 ( .I(n20581), .Z(n6230) );
  INV_X1 U1731 ( .I(n19909), .ZN(n29668) );
  NAND2_X1 U1744 ( .A1(n15286), .A2(n31766), .ZN(n15285) );
  OAI21_X1 U1759 ( .A1(n8421), .A2(n19971), .B(n31164), .ZN(n8759) );
  NOR3_X1 U1767 ( .A1(n20010), .A2(n20008), .A3(n9876), .ZN(n9341) );
  NAND3_X1 U1772 ( .A1(n20028), .A2(n20025), .A3(n1042), .ZN(n19735) );
  AOI22_X1 U1774 ( .A1(n1361), .A2(n11893), .B1(n3591), .B2(n19794), .ZN(n3590) );
  NOR2_X1 U1777 ( .A1(n34153), .A2(n20100), .ZN(n19562) );
  NOR2_X1 U1780 ( .A1(n30064), .A2(n16966), .ZN(n16979) );
  NOR2_X1 U1792 ( .A1(n20136), .A2(n20037), .ZN(n31766) );
  NAND2_X1 U1795 ( .A1(n10072), .A2(n19979), .ZN(n31443) );
  NAND3_X1 U1808 ( .A1(n18089), .A2(n7804), .A3(n31445), .ZN(n8015) );
  INV_X1 U1812 ( .I(n875), .ZN(n29840) );
  INV_X2 U1817 ( .I(n19867), .ZN(n17608) );
  AND2_X1 U1818 ( .A1(n29153), .A2(n4224), .Z(n29358) );
  INV_X1 U1829 ( .I(n10413), .ZN(n8147) );
  AND2_X1 U1845 ( .A1(n20113), .A2(n19907), .Z(n29373) );
  NOR2_X1 U1855 ( .A1(n27808), .A2(n16812), .ZN(n31697) );
  INV_X1 U1860 ( .I(n13650), .ZN(n30017) );
  NOR2_X1 U1869 ( .A1(n19901), .A2(n19900), .ZN(n5999) );
  CLKBUF_X2 U1875 ( .I(n12040), .Z(n6532) );
  INV_X1 U1878 ( .I(n1368), .ZN(n30819) );
  INV_X1 U1879 ( .I(n19764), .ZN(n31646) );
  INV_X1 U1886 ( .I(n27138), .ZN(n29689) );
  NAND2_X1 U1895 ( .A1(n5709), .A2(n5710), .ZN(n31573) );
  NAND2_X1 U1926 ( .A1(n16874), .A2(n30789), .ZN(n16873) );
  INV_X1 U1930 ( .I(n29781), .ZN(n31217) );
  NAND2_X1 U1932 ( .A1(n18977), .A2(n8092), .ZN(n30660) );
  AOI21_X1 U1933 ( .A1(n27743), .A2(n28705), .B(n16669), .ZN(n12498) );
  AND2_X1 U1945 ( .A1(n30663), .A2(n339), .Z(n10013) );
  CLKBUF_X2 U1962 ( .I(n19332), .Z(n28404) );
  NAND2_X1 U1968 ( .A1(n29815), .A2(n7687), .ZN(n30789) );
  NOR2_X1 U1972 ( .A1(n1384), .A2(n31352), .ZN(n31351) );
  NAND2_X1 U1975 ( .A1(n16960), .A2(n8335), .ZN(n19333) );
  BUF_X2 U1978 ( .I(n8606), .Z(n26830) );
  NAND3_X1 U1999 ( .A1(n29684), .A2(n3364), .A3(n29683), .ZN(n3361) );
  NAND3_X1 U2001 ( .A1(n26398), .A2(n18581), .A3(n18724), .ZN(n26591) );
  NOR2_X1 U2005 ( .A1(n18578), .A2(n30866), .ZN(n11319) );
  AOI22_X1 U2008 ( .A1(n485), .A2(n18571), .B1(n5753), .B2(n4868), .ZN(n5751)
         );
  NAND3_X1 U2011 ( .A1(n26717), .A2(n3601), .A3(n10579), .ZN(n2684) );
  NAND2_X1 U2018 ( .A1(n15956), .A2(n31519), .ZN(n18491) );
  NOR2_X1 U2020 ( .A1(n469), .A2(n25981), .ZN(n8271) );
  NOR2_X1 U2030 ( .A1(n1188), .A2(n8739), .ZN(n7977) );
  OAI22_X1 U2031 ( .A1(n16247), .A2(n16352), .B1(n18822), .B2(n18820), .ZN(
        n30001) );
  NAND3_X1 U2035 ( .A1(n18635), .A2(n5269), .A3(n6037), .ZN(n18636) );
  NAND2_X1 U2038 ( .A1(n17582), .A2(n16948), .ZN(n31339) );
  OR2_X1 U2044 ( .A1(n18574), .A2(n18617), .Z(n8821) );
  NOR2_X1 U2045 ( .A1(n6256), .A2(n13738), .ZN(n31519) );
  AND2_X1 U2048 ( .A1(n18586), .A2(n28964), .Z(n17165) );
  NOR2_X1 U2051 ( .A1(n18822), .A2(n16249), .ZN(n30698) );
  NOR2_X1 U2058 ( .A1(n18867), .A2(n31986), .ZN(n30908) );
  OAI21_X1 U2059 ( .A1(n3601), .A2(n26040), .B(n27228), .ZN(n11323) );
  NAND3_X1 U2060 ( .A1(n1188), .A2(n8739), .A3(n18639), .ZN(n18640) );
  NOR2_X1 U2061 ( .A1(n16569), .A2(n12006), .ZN(n18469) );
  CLKBUF_X1 U2064 ( .I(n15966), .Z(n26155) );
  BUF_X1 U2091 ( .I(n18186), .Z(n30744) );
  AOI21_X2 U2097 ( .A1(n18324), .A2(n34139), .B(n180), .ZN(n12214) );
  BUF_X4 U2099 ( .I(n24257), .Z(n6476) );
  OAI22_X2 U2106 ( .A1(n10731), .A2(n17228), .B1(n15832), .B2(n20516), .ZN(
        n30304) );
  OAI21_X2 U2107 ( .A1(n13300), .A2(n33301), .B(n13830), .ZN(n20311) );
  NOR2_X2 U2113 ( .A1(n18487), .A2(n18827), .ZN(n18462) );
  BUF_X2 U2114 ( .I(n15955), .Z(n14828) );
  NAND2_X2 U2121 ( .A1(n29398), .A2(n19225), .ZN(n13938) );
  BUF_X2 U2124 ( .I(n17237), .Z(n8454) );
  BUF_X4 U2125 ( .I(n2396), .Z(n2141) );
  AOI21_X2 U2127 ( .A1(n1373), .A2(n11940), .B(n1764), .ZN(n1763) );
  AND2_X1 U2129 ( .A1(n18768), .A2(n16849), .Z(n18376) );
  BUF_X4 U2142 ( .I(n18722), .Z(n29602) );
  OR2_X1 U2154 ( .A1(n10568), .A2(n28014), .Z(n22466) );
  OAI21_X2 U2161 ( .A1(n12590), .A2(n20079), .B(n6444), .ZN(n26961) );
  INV_X2 U2170 ( .I(n14789), .ZN(n27545) );
  NAND2_X1 U2171 ( .A1(n30976), .A2(n5374), .ZN(n29621) );
  INV_X2 U2177 ( .I(n26445), .ZN(n28435) );
  AOI21_X2 U2198 ( .A1(n1287), .A2(n30405), .B(n29232), .ZN(n27565) );
  NAND3_X2 U2200 ( .A1(n12053), .A2(n14283), .A3(n1039), .ZN(n31319) );
  AND2_X1 U2210 ( .A1(n21306), .A2(n21305), .Z(n29382) );
  NAND2_X2 U2218 ( .A1(n15830), .A2(n22992), .ZN(n30388) );
  INV_X2 U2230 ( .I(n23156), .ZN(n18133) );
  AOI21_X2 U2231 ( .A1(n1170), .A2(n19456), .B(n16681), .ZN(n6858) );
  BUF_X2 U2232 ( .I(n18696), .Z(n16569) );
  INV_X4 U2234 ( .I(n7287), .ZN(n23055) );
  OR2_X1 U2245 ( .A1(n18696), .A2(n18831), .Z(n13015) );
  OR2_X1 U2246 ( .A1(n23540), .A2(n24283), .Z(n28781) );
  INV_X2 U2254 ( .I(n28091), .ZN(n30737) );
  INV_X2 U2266 ( .I(n25201), .ZN(n25200) );
  INV_X4 U2268 ( .I(n16651), .ZN(n29056) );
  INV_X2 U2270 ( .I(n29153), .ZN(n6962) );
  OAI22_X1 U2274 ( .A1(n16254), .A2(n6360), .B1(n6012), .B2(n16022), .ZN(n5874) );
  OAI21_X1 U2275 ( .A1(n23708), .A2(n16238), .B(n14974), .ZN(n12509) );
  NAND2_X1 U2283 ( .A1(n12837), .A2(n17223), .ZN(n18029) );
  NAND2_X1 U2284 ( .A1(n17582), .A2(n17223), .ZN(n16338) );
  INV_X1 U2285 ( .I(n17223), .ZN(n29751) );
  CLKBUF_X2 U2286 ( .I(n10469), .Z(n7371) );
  NAND3_X1 U2291 ( .A1(n1290), .A2(n6478), .A3(n8409), .ZN(n22555) );
  INV_X1 U2293 ( .I(n25903), .ZN(n29771) );
  NAND2_X1 U2295 ( .A1(n31801), .A2(n7093), .ZN(n29584) );
  NAND2_X1 U2303 ( .A1(n5417), .A2(n15038), .ZN(n30515) );
  OAI21_X1 U2321 ( .A1(n29261), .A2(n900), .B(n22476), .ZN(n30383) );
  AOI21_X1 U2331 ( .A1(n15757), .A2(n11556), .B(n15755), .ZN(n15769) );
  NOR2_X1 U2336 ( .A1(n17120), .A2(n30221), .ZN(n31245) );
  AND2_X1 U2338 ( .A1(n33007), .A2(n22795), .Z(n29438) );
  INV_X1 U2345 ( .I(n10111), .ZN(n24781) );
  NAND2_X1 U2352 ( .A1(n29107), .A2(n23058), .ZN(n14418) );
  INV_X2 U2357 ( .I(n25736), .ZN(n25744) );
  NAND2_X1 U2358 ( .A1(n14721), .A2(n21223), .ZN(n21316) );
  NOR3_X1 U2360 ( .A1(n26868), .A2(n14188), .A3(n28697), .ZN(n16140) );
  NOR2_X1 U2395 ( .A1(n18764), .A2(n18767), .ZN(n31521) );
  NAND2_X1 U2397 ( .A1(n30369), .A2(n25211), .ZN(n10942) );
  NAND2_X1 U2406 ( .A1(n6483), .A2(n21721), .ZN(n14076) );
  CLKBUF_X2 U2416 ( .I(n24914), .Z(n27248) );
  OAI22_X1 U2417 ( .A1(n12615), .A2(n23144), .B1(n17257), .B2(n6479), .ZN(
        n26392) );
  INV_X1 U2431 ( .I(n12329), .ZN(n25076) );
  INV_X1 U2439 ( .I(n661), .ZN(n4892) );
  CLKBUF_X4 U2444 ( .I(n16141), .Z(n12) );
  NOR2_X1 U2454 ( .A1(n13985), .A2(n25198), .ZN(n1861) );
  AOI21_X1 U2463 ( .A1(n16117), .A2(n5056), .B(n13073), .ZN(n18221) );
  OAI21_X1 U2480 ( .A1(n7655), .A2(n1215), .B(n27342), .ZN(n1859) );
  NAND2_X1 U2495 ( .A1(n13268), .A2(n24210), .ZN(n24321) );
  OAI21_X1 U2521 ( .A1(n28473), .A2(n28472), .B(n22435), .ZN(n11441) );
  OAI21_X1 U2537 ( .A1(n15359), .A2(n25214), .B(n15339), .ZN(n30369) );
  AND2_X1 U2544 ( .A1(n29304), .A2(n8275), .Z(n4812) );
  NAND3_X1 U2545 ( .A1(n27123), .A2(n29085), .A3(n1071), .ZN(n4768) );
  OAI21_X1 U2548 ( .A1(n16097), .A2(n23848), .B(n23847), .ZN(n10762) );
  BUF_X2 U2554 ( .I(n23567), .Z(n23848) );
  INV_X1 U2574 ( .I(n9664), .ZN(n10483) );
  BUF_X2 U2584 ( .I(n4599), .Z(n3898) );
  NOR2_X1 U2593 ( .A1(n15054), .A2(n2191), .ZN(n7928) );
  BUF_X2 U2599 ( .I(n24147), .Z(n4019) );
  NAND2_X1 U2623 ( .A1(n2746), .A2(n2745), .ZN(n30110) );
  BUF_X2 U2626 ( .I(n5128), .Z(n4781) );
  NAND2_X1 U2628 ( .A1(n25132), .A2(n1083), .ZN(n31780) );
  INV_X1 U2630 ( .I(n1083), .ZN(n31779) );
  INV_X2 U2644 ( .I(n25867), .ZN(n790) );
  NOR3_X1 U2646 ( .A1(n29706), .A2(n13049), .A3(n25847), .ZN(n15944) );
  OAI21_X1 U2666 ( .A1(n24715), .A2(n16323), .B(n9195), .ZN(n24716) );
  NOR2_X1 U2670 ( .A1(n16323), .A2(n25701), .ZN(n24449) );
  OR2_X1 U2679 ( .A1(n9163), .A2(n9164), .Z(n27376) );
  NOR2_X1 U2687 ( .A1(n11575), .A2(n6882), .ZN(n642) );
  AND2_X1 U2702 ( .A1(n17927), .A2(n10858), .Z(n9655) );
  NOR2_X1 U2758 ( .A1(n19857), .A2(n17711), .ZN(n11903) );
  NAND2_X1 U2768 ( .A1(n31920), .A2(n4490), .ZN(n24711) );
  OAI21_X1 U2770 ( .A1(n16467), .A2(n9391), .B(n7073), .ZN(n7505) );
  NAND2_X1 U2771 ( .A1(n27479), .A2(n13709), .ZN(n12293) );
  NAND2_X1 U2780 ( .A1(n22422), .A2(n906), .ZN(n30639) );
  NOR2_X1 U2790 ( .A1(n11299), .A2(n12363), .ZN(n12372) );
  AND2_X1 U2810 ( .A1(n9199), .A2(n651), .Z(n13666) );
  NOR2_X1 U2817 ( .A1(n6910), .A2(n25394), .ZN(n25347) );
  NOR2_X1 U2822 ( .A1(n30139), .A2(n1863), .ZN(n31286) );
  NAND2_X1 U2823 ( .A1(n6668), .A2(n2042), .ZN(n6667) );
  INV_X1 U2826 ( .I(n19509), .ZN(n8456) );
  AND2_X1 U2838 ( .A1(n14335), .A2(n3860), .Z(n1978) );
  AND2_X1 U2841 ( .A1(n14335), .A2(n31294), .Z(n31293) );
  AND2_X1 U2842 ( .A1(n6595), .A2(n8766), .Z(n8710) );
  INV_X1 U2845 ( .I(n11334), .ZN(n6133) );
  NOR2_X1 U2849 ( .A1(n11334), .A2(n22584), .ZN(n17007) );
  NAND2_X1 U2879 ( .A1(n15550), .A2(n13050), .ZN(n12677) );
  BUF_X2 U2894 ( .I(n25221), .Z(n28651) );
  CLKBUF_X2 U2915 ( .I(n29157), .Z(n31722) );
  NAND3_X1 U2916 ( .A1(n30328), .A2(n24927), .A3(n2180), .ZN(n24350) );
  CLKBUF_X1 U2921 ( .I(n11931), .Z(n27057) );
  NOR2_X1 U2922 ( .A1(n11931), .A2(n10504), .ZN(n25617) );
  CLKBUF_X2 U2923 ( .I(n14865), .Z(n254) );
  INV_X1 U2925 ( .I(n14865), .ZN(n25003) );
  NAND2_X1 U2950 ( .A1(n29253), .A2(n8100), .ZN(n13962) );
  NAND2_X1 U2953 ( .A1(n12677), .A2(n25884), .ZN(n24463) );
  NAND2_X1 U2954 ( .A1(n25884), .A2(n14832), .ZN(n4932) );
  AND2_X1 U2965 ( .A1(n25973), .A2(n24251), .Z(n29376) );
  NOR2_X1 U2971 ( .A1(n25060), .A2(n25051), .ZN(n25063) );
  NAND3_X1 U2976 ( .A1(n12974), .A2(n842), .A3(n14756), .ZN(n16947) );
  NOR2_X1 U2979 ( .A1(n25980), .A2(n14210), .ZN(n12784) );
  AND2_X1 U2981 ( .A1(n7748), .A2(n1984), .Z(n1983) );
  AND3_X1 U2985 ( .A1(n5760), .A2(n18990), .A3(n18017), .Z(n10867) );
  BUF_X2 U2989 ( .I(n18017), .Z(n28171) );
  AOI21_X1 U3002 ( .A1(n21811), .A2(n28181), .B(n1328), .ZN(n21349) );
  AOI22_X1 U3017 ( .A1(n891), .A2(n3506), .B1(n29576), .B2(n28410), .ZN(n6106)
         );
  AOI22_X1 U3019 ( .A1(n10567), .A2(n790), .B1(n18219), .B2(n790), .ZN(n10566)
         );
  NOR2_X1 U3026 ( .A1(n16041), .A2(n72), .ZN(n16937) );
  INV_X2 U3030 ( .I(n16041), .ZN(n25312) );
  NAND2_X1 U3040 ( .A1(n31916), .A2(n29268), .ZN(n23616) );
  INV_X1 U3056 ( .I(n13159), .ZN(n16817) );
  OAI21_X1 U3077 ( .A1(n16149), .A2(n22576), .B(n16567), .ZN(n6657) );
  NOR3_X1 U3112 ( .A1(n1119), .A2(n1926), .A3(n1805), .ZN(n1887) );
  OAI21_X1 U3125 ( .A1(n1165), .A2(n13061), .B(n31684), .ZN(n14988) );
  NAND3_X1 U3131 ( .A1(n15736), .A2(n31684), .A3(n1165), .ZN(n15735) );
  NOR2_X1 U3132 ( .A1(n1165), .A2(n29152), .ZN(n15306) );
  OAI21_X1 U3152 ( .A1(n15189), .A2(n20155), .B(n3486), .ZN(n6069) );
  INV_X1 U3156 ( .I(n5988), .ZN(n25575) );
  AOI22_X1 U3157 ( .A1(n19117), .A2(n28404), .B1(n19154), .B2(n8862), .ZN(
        n12368) );
  OAI21_X1 U3162 ( .A1(n880), .A2(n879), .B(n19154), .ZN(n16221) );
  NOR2_X1 U3169 ( .A1(n11366), .A2(n16528), .ZN(n30372) );
  NOR2_X1 U3182 ( .A1(n17894), .A2(n25901), .ZN(n4205) );
  AND2_X1 U3186 ( .A1(n386), .A2(n30089), .Z(n15404) );
  NOR2_X1 U3191 ( .A1(n7195), .A2(n21441), .ZN(n2689) );
  OAI21_X1 U3196 ( .A1(n31195), .A2(n7195), .B(n21441), .ZN(n7196) );
  AOI21_X1 U3198 ( .A1(n796), .A2(n10226), .B(n7935), .ZN(n11341) );
  NOR2_X1 U3208 ( .A1(n21864), .A2(n21865), .ZN(n8619) );
  NAND4_X1 U3225 ( .A1(n3052), .A2(n3057), .A3(n3051), .A4(n18123), .ZN(n3056)
         );
  NAND2_X1 U3226 ( .A1(n15283), .A2(n30586), .ZN(n12319) );
  INV_X1 U3227 ( .I(n19754), .ZN(n26230) );
  OAI22_X1 U3243 ( .A1(n24988), .A2(n713), .B1(n24994), .B2(n4525), .ZN(n24989) );
  NAND2_X1 U3248 ( .A1(n6500), .A2(n11617), .ZN(n30551) );
  AOI21_X1 U3250 ( .A1(n21587), .A2(n26766), .B(n30806), .ZN(n21589) );
  NOR3_X1 U3267 ( .A1(n1211), .A2(n28338), .A3(n1212), .ZN(n13296) );
  AOI21_X1 U3271 ( .A1(n6763), .A2(n3340), .B(n7134), .ZN(n3343) );
  INV_X2 U3273 ( .I(n6763), .ZN(n31139) );
  BUF_X2 U3291 ( .I(n15255), .Z(n26912) );
  INV_X1 U3298 ( .I(n15255), .ZN(n25588) );
  NAND3_X1 U3299 ( .A1(n15255), .A2(n11820), .A3(n34169), .ZN(n25534) );
  OAI21_X1 U3305 ( .A1(n4281), .A2(n28265), .B(n30527), .ZN(n7538) );
  BUF_X2 U3311 ( .I(n32309), .Z(n4281) );
  NAND3_X1 U3313 ( .A1(n15278), .A2(n10484), .A3(n19933), .ZN(n1813) );
  NAND2_X1 U3332 ( .A1(n26447), .A2(n27173), .ZN(n28931) );
  NAND2_X1 U3336 ( .A1(n791), .A2(n16688), .ZN(n6250) );
  INV_X1 U3337 ( .I(n5932), .ZN(n15264) );
  NOR2_X1 U3344 ( .A1(n25637), .A2(n2378), .ZN(n25638) );
  CLKBUF_X2 U3346 ( .I(n21455), .Z(n29088) );
  CLKBUF_X2 U3347 ( .I(n3880), .Z(n30969) );
  NAND2_X1 U3348 ( .A1(n24084), .A2(n3880), .ZN(n14677) );
  NAND2_X1 U3354 ( .A1(n33722), .A2(n23813), .ZN(n31294) );
  INV_X1 U3363 ( .I(n25816), .ZN(n25826) );
  INV_X1 U3374 ( .I(n23924), .ZN(n23736) );
  OAI21_X1 U3386 ( .A1(n20437), .A2(n20438), .B(n30099), .ZN(n2650) );
  OAI22_X1 U3391 ( .A1(n26520), .A2(n18827), .B1(n18489), .B2(n18487), .ZN(
        n17251) );
  NAND2_X1 U3392 ( .A1(n18487), .A2(n18827), .ZN(n18332) );
  INV_X2 U3393 ( .I(n26791), .ZN(n18487) );
  AOI21_X1 U3394 ( .A1(n11888), .A2(n354), .B(n8217), .ZN(n13503) );
  NAND2_X1 U3402 ( .A1(n32063), .A2(n24956), .ZN(n24954) );
  NOR2_X1 U3403 ( .A1(n1201), .A2(n32063), .ZN(n8639) );
  INV_X1 U3416 ( .I(n23266), .ZN(n23445) );
  INV_X1 U3430 ( .I(n14031), .ZN(n1247) );
  AND2_X2 U3443 ( .A1(n11913), .A2(n16), .Z(n29281) );
  AND2_X1 U3445 ( .A1(n29022), .A2(n20100), .Z(n29283) );
  INV_X1 U3447 ( .I(n8713), .ZN(n19921) );
  BUF_X2 U3449 ( .I(n8713), .Z(n1826) );
  XNOR2_X1 U3461 ( .A1(n10949), .A2(n6906), .ZN(n29285) );
  NOR2_X2 U3465 ( .A1(n7954), .A2(n7955), .ZN(n6431) );
  INV_X1 U3470 ( .I(n20882), .ZN(n21391) );
  INV_X2 U3485 ( .I(n14045), .ZN(n853) );
  XNOR2_X1 U3497 ( .A1(n23224), .A2(n16691), .ZN(n29291) );
  INV_X2 U3502 ( .I(n6169), .ZN(n14136) );
  INV_X2 U3513 ( .I(n4286), .ZN(n15520) );
  INV_X2 U3520 ( .I(n23301), .ZN(n30380) );
  INV_X4 U3527 ( .I(n25756), .ZN(n1211) );
  BUF_X2 U3543 ( .I(n7242), .Z(n28836) );
  AND2_X2 U3550 ( .A1(n9490), .A2(n8277), .Z(n15446) );
  INV_X1 U3560 ( .I(n4110), .ZN(n22830) );
  NAND3_X1 U3572 ( .A1(n16835), .A2(n700), .A3(n25867), .ZN(n11254) );
  INV_X1 U3573 ( .I(n6255), .ZN(n20481) );
  BUF_X2 U3584 ( .I(n29471), .Z(n29294) );
  OAI21_X1 U3585 ( .A1(n5272), .A2(n836), .B(n25901), .ZN(n5271) );
  INV_X1 U3617 ( .I(n23808), .ZN(n31483) );
  AOI21_X1 U3627 ( .A1(n5670), .A2(n5779), .B(n26585), .ZN(n5669) );
  OR2_X2 U3629 ( .A1(n28545), .A2(n26606), .Z(n22646) );
  NAND2_X1 U3632 ( .A1(n20527), .A2(n16515), .ZN(n17392) );
  INV_X2 U3648 ( .I(n11372), .ZN(n13273) );
  NAND2_X1 U3650 ( .A1(n11372), .A2(n25977), .ZN(n3791) );
  AND2_X2 U3651 ( .A1(n9280), .A2(n9951), .Z(n22843) );
  NAND3_X1 U3654 ( .A1(n30902), .A2(n21512), .A3(n9057), .ZN(n27437) );
  NOR2_X1 U3657 ( .A1(n21755), .A2(n21512), .ZN(n8276) );
  INV_X2 U3674 ( .I(n6669), .ZN(n17077) );
  NAND2_X1 U3676 ( .A1(n31911), .A2(n31309), .ZN(n21801) );
  OAI22_X1 U3687 ( .A1(n17255), .A2(n18617), .B1(n17062), .B2(n16948), .ZN(
        n31333) );
  NAND2_X1 U3696 ( .A1(n15108), .A2(n18617), .ZN(n14536) );
  AND2_X1 U3701 ( .A1(n1119), .A2(n13862), .Z(n1594) );
  INV_X1 U3733 ( .I(n24621), .ZN(n31088) );
  NOR2_X1 U3741 ( .A1(n18546), .A2(n1185), .ZN(n9510) );
  INV_X1 U3743 ( .I(n18546), .ZN(n18647) );
  NOR2_X1 U3746 ( .A1(n18546), .A2(n26810), .ZN(n18363) );
  NOR2_X2 U3753 ( .A1(n21321), .A2(n21322), .ZN(n21190) );
  NOR2_X1 U3761 ( .A1(n18110), .A2(n16129), .ZN(n13582) );
  AOI21_X1 U3778 ( .A1(n1041), .A2(n20097), .B(n16789), .ZN(n17442) );
  INV_X1 U3794 ( .I(n13720), .ZN(n798) );
  BUF_X4 U3806 ( .I(n17278), .Z(n29299) );
  NAND2_X1 U3815 ( .A1(n12902), .A2(n20311), .ZN(n31188) );
  AOI21_X2 U3822 ( .A1(n17639), .A2(n14603), .B(n14602), .ZN(n14601) );
  NAND2_X2 U3823 ( .A1(n12836), .A2(n9439), .ZN(n27218) );
  NAND2_X1 U3833 ( .A1(n11368), .A2(n20423), .ZN(n26399) );
  INV_X1 U3853 ( .I(n19057), .ZN(n1387) );
  INV_X2 U3864 ( .I(n14954), .ZN(n10822) );
  NAND2_X1 U3865 ( .A1(n12329), .A2(n14954), .ZN(n25067) );
  NAND2_X1 U3880 ( .A1(n10883), .A2(n27007), .ZN(n39) );
  INV_X1 U3883 ( .I(n27007), .ZN(n29635) );
  NAND2_X1 U3885 ( .A1(n27007), .A2(n22824), .ZN(n17605) );
  AND2_X2 U3886 ( .A1(n27007), .A2(n22592), .Z(n22823) );
  OAI21_X1 U3899 ( .A1(n14168), .A2(n21072), .B(n5141), .ZN(n31025) );
  BUF_X2 U3914 ( .I(n10631), .Z(n31508) );
  NOR2_X1 U3933 ( .A1(n15864), .A2(n30506), .ZN(n12280) );
  BUF_X2 U3948 ( .I(n16710), .Z(n28378) );
  AND3_X1 U3962 ( .A1(n21568), .A2(n21569), .A3(n30389), .Z(n21570) );
  NOR4_X1 U3976 ( .A1(n22729), .A2(n22730), .A3(n22731), .A4(n22732), .ZN(
        n12055) );
  INV_X1 U3980 ( .I(n5454), .ZN(n13048) );
  AOI21_X1 U3983 ( .A1(n14620), .A2(n20261), .B(n32747), .ZN(n1929) );
  AOI21_X1 U4005 ( .A1(n16688), .A2(n16554), .B(n24219), .ZN(n12357) );
  CLKBUF_X12 U4006 ( .I(n16554), .Z(n26916) );
  NOR2_X1 U4029 ( .A1(n1323), .A2(n7868), .ZN(n17547) );
  OR2_X2 U4032 ( .A1(n10438), .A2(n4735), .Z(n7561) );
  OR3_X2 U4049 ( .A1(n11208), .A2(n12211), .A3(n8313), .Z(n5309) );
  NAND2_X1 U4077 ( .A1(n16018), .A2(n16181), .ZN(n5428) );
  NOR3_X1 U4079 ( .A1(n16181), .A2(n489), .A3(n29658), .ZN(n9631) );
  OAI22_X1 U4080 ( .A1(n19333), .A2(n28404), .B1(n19331), .B2(n8862), .ZN(
        n26503) );
  NAND2_X1 U4090 ( .A1(n1094), .A2(n13412), .ZN(n1640) );
  BUF_X4 U4120 ( .I(n15536), .Z(n29307) );
  INV_X1 U4122 ( .I(n23438), .ZN(n29231) );
  INV_X1 U4124 ( .I(n12652), .ZN(n5157) );
  INV_X1 U4136 ( .I(n18283), .ZN(n12837) );
  BUF_X2 U4139 ( .I(n18283), .Z(n18617) );
  AOI21_X2 U4140 ( .A1(n28278), .A2(n34046), .B(n11890), .ZN(n12794) );
  NAND2_X1 U4149 ( .A1(n16688), .A2(n24220), .ZN(n23624) );
  INV_X1 U4175 ( .I(n21551), .ZN(n30511) );
  OAI21_X2 U4182 ( .A1(n20057), .A2(n20058), .B(n19867), .ZN(n27840) );
  OAI22_X1 U4188 ( .A1(n11199), .A2(n20154), .B1(n11198), .B2(n19926), .ZN(
        n19918) );
  NOR2_X1 U4194 ( .A1(n20157), .A2(n20156), .ZN(n16795) );
  NAND3_X1 U4202 ( .A1(n30934), .A2(n33687), .A3(n34139), .ZN(n11919) );
  OAI21_X1 U4211 ( .A1(n18567), .A2(n34139), .B(n12154), .ZN(n12153) );
  NAND2_X1 U4225 ( .A1(n23956), .A2(n23955), .ZN(n14521) );
  OR3_X2 U4249 ( .A1(n25121), .A2(n1567), .A3(n16293), .Z(n24889) );
  OAI22_X1 U4288 ( .A1(n11311), .A2(n781), .B1(n20447), .B2(n26424), .ZN(n7955) );
  INV_X2 U4338 ( .I(n20756), .ZN(n6218) );
  INV_X1 U4345 ( .I(n27077), .ZN(n1382) );
  NAND3_X1 U4356 ( .A1(n15646), .A2(n24780), .A3(n24983), .ZN(n4216) );
  INV_X2 U4357 ( .I(n24780), .ZN(n15084) );
  CLKBUF_X4 U4371 ( .I(n25146), .Z(n1786) );
  NOR2_X1 U4385 ( .A1(n21832), .A2(n5170), .ZN(n12161) );
  NOR2_X1 U4413 ( .A1(n14839), .A2(n24163), .ZN(n29568) );
  INV_X1 U4415 ( .I(n23333), .ZN(n28323) );
  NAND2_X2 U4434 ( .A1(n583), .A2(n9288), .ZN(n30530) );
  NOR2_X2 U4450 ( .A1(n25985), .A2(n33335), .ZN(n19146) );
  NOR2_X1 U4462 ( .A1(n22361), .A2(n4135), .ZN(n26609) );
  AND2_X1 U4468 ( .A1(n31637), .A2(n22361), .Z(n29430) );
  INV_X2 U4472 ( .I(n20450), .ZN(n20378) );
  OR2_X2 U4479 ( .A1(n32055), .A2(n9064), .Z(n22600) );
  INV_X1 U4483 ( .I(n18184), .ZN(n21808) );
  INV_X1 U4487 ( .I(n18411), .ZN(n18848) );
  BUF_X2 U4488 ( .I(n18411), .Z(n18846) );
  INV_X1 U4491 ( .I(n18078), .ZN(n9783) );
  NAND2_X1 U4504 ( .A1(n23079), .A2(n22885), .ZN(n31712) );
  NOR2_X1 U4514 ( .A1(n20160), .A2(n14138), .ZN(n26555) );
  OAI22_X1 U4517 ( .A1(n4683), .A2(n1146), .B1(n8010), .B2(n5049), .ZN(n8175)
         );
  BUF_X4 U4522 ( .I(n31951), .Z(n19926) );
  NAND2_X1 U4525 ( .A1(n5889), .A2(n27921), .ZN(n19363) );
  AND2_X2 U4528 ( .A1(n15343), .A2(n22521), .Z(n22522) );
  INV_X1 U4540 ( .I(n21198), .ZN(n21405) );
  INV_X1 U4563 ( .I(n30637), .ZN(n16190) );
  NAND2_X1 U4565 ( .A1(n15692), .A2(n23877), .ZN(n9975) );
  NOR2_X1 U4573 ( .A1(n4820), .A2(n23742), .ZN(n30172) );
  NAND2_X1 U4582 ( .A1(n13759), .A2(n8087), .ZN(n13785) );
  AOI21_X1 U4583 ( .A1(n8087), .A2(n33515), .B(n9688), .ZN(n13830) );
  OAI21_X1 U4589 ( .A1(n13509), .A2(n17313), .B(n26133), .ZN(n14955) );
  NAND2_X1 U4601 ( .A1(n19057), .A2(n7345), .ZN(n8092) );
  AND2_X2 U4613 ( .A1(n25894), .A2(n9125), .Z(n28910) );
  AND2_X2 U4624 ( .A1(n8899), .A2(n595), .Z(n7721) );
  NAND2_X1 U4636 ( .A1(n20529), .A2(n30637), .ZN(n20528) );
  NOR2_X1 U4653 ( .A1(n20529), .A2(n30637), .ZN(n20196) );
  NAND2_X1 U4655 ( .A1(n19088), .A2(n18990), .ZN(n31352) );
  CLKBUF_X12 U4667 ( .I(n18869), .Z(n29308) );
  BUF_X4 U4668 ( .I(n18869), .Z(n29309) );
  INV_X1 U4685 ( .I(n5414), .ZN(n31059) );
  INV_X2 U4697 ( .I(n5440), .ZN(n6072) );
  NAND2_X1 U4699 ( .A1(n5440), .A2(n5441), .ZN(n11334) );
  NAND2_X1 U4705 ( .A1(n22586), .A2(n33320), .ZN(n22587) );
  NAND2_X1 U4709 ( .A1(n12421), .A2(n2821), .ZN(n19830) );
  INV_X1 U4735 ( .I(n27503), .ZN(n21080) );
  NAND2_X1 U4740 ( .A1(n29655), .A2(n27931), .ZN(n14460) );
  OR2_X2 U4743 ( .A1(n8469), .A2(n4568), .Z(n8467) );
  NAND2_X1 U4746 ( .A1(n5433), .A2(n1168), .ZN(n13058) );
  NAND2_X1 U4758 ( .A1(n5433), .A2(n17670), .ZN(n4744) );
  INV_X1 U4767 ( .I(n12040), .ZN(n19987) );
  BUF_X4 U4776 ( .I(n2041), .Z(n29312) );
  NAND2_X1 U4782 ( .A1(n16621), .A2(n24180), .ZN(n27786) );
  CLKBUF_X12 U4783 ( .I(n30410), .Z(n29313) );
  BUF_X4 U4789 ( .I(n30410), .Z(n29314) );
  CLKBUF_X4 U4795 ( .I(n4669), .Z(n29315) );
  CLKBUF_X12 U4798 ( .I(n16354), .Z(n14130) );
  AOI21_X1 U4817 ( .A1(n21357), .A2(n12037), .B(n21358), .ZN(n30226) );
  NOR2_X1 U4823 ( .A1(n12863), .A2(n10903), .ZN(n12663) );
  OAI22_X1 U4827 ( .A1(n7497), .A2(n10903), .B1(n7495), .B2(n12863), .ZN(
        n27215) );
  AOI22_X1 U4846 ( .A1(n18595), .A2(n18731), .B1(n18845), .B2(n18596), .ZN(
        n26458) );
  CLKBUF_X4 U4853 ( .I(n20064), .Z(n16630) );
  INV_X1 U4873 ( .I(n16022), .ZN(n6360) );
  NOR2_X1 U4914 ( .A1(n22865), .A2(n4084), .ZN(n12578) );
  INV_X2 U4919 ( .I(n4084), .ZN(n10641) );
  BUF_X4 U4920 ( .I(n29321), .Z(n29322) );
  NAND3_X1 U4921 ( .A1(n16490), .A2(n32172), .A3(n15089), .ZN(n21882) );
  OAI21_X1 U4923 ( .A1(n22678), .A2(n15089), .B(n16570), .ZN(n15911) );
  NOR2_X1 U4926 ( .A1(n16563), .A2(n2839), .ZN(n23757) );
  INV_X2 U4931 ( .I(n432), .ZN(n17472) );
  NOR2_X1 U4933 ( .A1(n432), .A2(n16194), .ZN(n31557) );
  NAND2_X1 U4955 ( .A1(n20630), .A2(n14564), .ZN(n30496) );
  NOR2_X1 U4958 ( .A1(n30326), .A2(n12827), .ZN(n13332) );
  OAI22_X1 U4974 ( .A1(n6671), .A2(n12517), .B1(n19908), .B2(n16298), .ZN(
        n6377) );
  CLKBUF_X4 U4975 ( .I(n7552), .Z(n53) );
  NOR2_X1 U4986 ( .A1(n29253), .A2(n17967), .ZN(n8108) );
  INV_X2 U4998 ( .I(n17967), .ZN(n7804) );
  BUF_X2 U5020 ( .I(n20152), .Z(n8259) );
  NAND2_X1 U5037 ( .A1(n29118), .A2(n26969), .ZN(n9441) );
  INV_X2 U5064 ( .I(n5696), .ZN(n14183) );
  NAND2_X1 U5070 ( .A1(n6453), .A2(n3103), .ZN(n14555) );
  INV_X2 U5078 ( .I(n21870), .ZN(n12394) );
  NOR2_X1 U5098 ( .A1(n18078), .A2(n6679), .ZN(n20223) );
  CLKBUF_X12 U5110 ( .I(n18586), .Z(n18587) );
  OR3_X2 U5121 ( .A1(n27619), .A2(n26445), .A3(n27336), .Z(n615) );
  INV_X2 U5129 ( .I(n27726), .ZN(n826) );
  NAND2_X1 U5131 ( .A1(n29302), .A2(n16194), .ZN(n21494) );
  NOR2_X1 U5147 ( .A1(n21211), .A2(n16906), .ZN(n12066) );
  NAND2_X1 U5149 ( .A1(n14402), .A2(n7287), .ZN(n31790) );
  BUF_X4 U5158 ( .I(n22909), .Z(n29329) );
  NOR2_X1 U5165 ( .A1(n16249), .A2(n18820), .ZN(n12976) );
  NOR2_X1 U5169 ( .A1(n9484), .A2(n2958), .ZN(n9483) );
  NAND2_X1 U5188 ( .A1(n31837), .A2(n11789), .ZN(n8279) );
  INV_X1 U5196 ( .I(n11789), .ZN(n24222) );
  BUF_X2 U5198 ( .I(n2600), .Z(n29331) );
  NAND3_X1 U5204 ( .A1(n13751), .A2(n5915), .A3(n14183), .ZN(n3160) );
  CLKBUF_X12 U5228 ( .I(n18763), .Z(n16559) );
  NAND2_X1 U5232 ( .A1(n28028), .A2(n20534), .ZN(n6925) );
  NAND2_X1 U5265 ( .A1(n1239), .A2(n24262), .ZN(n16574) );
  INV_X2 U5268 ( .I(n24262), .ZN(n26950) );
  INV_X1 U5278 ( .I(n17015), .ZN(n23785) );
  INV_X1 U5282 ( .I(n17927), .ZN(n830) );
  OAI22_X1 U5291 ( .A1(n15944), .A2(n25848), .B1(n25857), .B2(n14915), .ZN(
        n30808) );
  NAND2_X1 U5293 ( .A1(n27057), .A2(n12049), .ZN(n30831) );
  INV_X2 U5308 ( .I(n24965), .ZN(n24969) );
  NAND2_X1 U5325 ( .A1(n29593), .A2(n7688), .ZN(n4900) );
  INV_X1 U5334 ( .I(n29594), .ZN(n29593) );
  NAND2_X1 U5348 ( .A1(n9857), .A2(n9859), .ZN(n9856) );
  INV_X1 U5384 ( .I(n24878), .ZN(n31602) );
  BUF_X2 U5387 ( .I(n25762), .Z(n17120) );
  CLKBUF_X1 U5411 ( .I(n679), .Z(n30308) );
  INV_X1 U5415 ( .I(n24390), .ZN(n30883) );
  INV_X1 U5419 ( .I(n14727), .ZN(n24660) );
  NAND2_X1 U5431 ( .A1(n16901), .A2(n29512), .ZN(n13660) );
  AND2_X1 U5446 ( .A1(n24244), .A2(n1235), .Z(n29387) );
  NOR2_X1 U5451 ( .A1(n15996), .A2(n11200), .ZN(n31033) );
  AND3_X1 U5455 ( .A1(n6003), .A2(n33868), .A3(n24095), .Z(n29397) );
  OR2_X1 U5466 ( .A1(n30270), .A2(n31772), .Z(n273) );
  NOR2_X1 U5469 ( .A1(n27826), .A2(n9323), .ZN(n27971) );
  CLKBUF_X2 U5502 ( .I(n14770), .Z(n29985) );
  INV_X1 U5503 ( .I(n9368), .ZN(n31544) );
  CLKBUF_X2 U5506 ( .I(n4655), .Z(n31355) );
  CLKBUF_X2 U5511 ( .I(n15663), .Z(n29655) );
  AND2_X1 U5525 ( .A1(n27392), .A2(n29131), .Z(n30283) );
  INV_X1 U5540 ( .I(n27184), .ZN(n31615) );
  INV_X1 U5547 ( .I(n29590), .ZN(n12399) );
  NAND2_X1 U5550 ( .A1(n7475), .A2(n14133), .ZN(n30886) );
  OAI21_X1 U5553 ( .A1(n7088), .A2(n26965), .B(n2447), .ZN(n31247) );
  NAND2_X1 U5556 ( .A1(n18152), .A2(n23940), .ZN(n29708) );
  AND2_X1 U5565 ( .A1(n27474), .A2(n30408), .Z(n29368) );
  INV_X1 U5570 ( .I(n6309), .ZN(n23954) );
  NAND2_X1 U5583 ( .A1(n13291), .A2(n31916), .ZN(n31601) );
  INV_X1 U5586 ( .I(n299), .ZN(n30408) );
  CLKBUF_X4 U5619 ( .I(n27996), .Z(n31491) );
  NAND2_X1 U5621 ( .A1(n14417), .A2(n13977), .ZN(n29614) );
  NOR2_X1 U5629 ( .A1(n30868), .A2(n10296), .ZN(n17464) );
  NOR2_X1 U5632 ( .A1(n1277), .A2(n15577), .ZN(n30968) );
  AOI22_X1 U5633 ( .A1(n23104), .A2(n26724), .B1(n5448), .B2(n22582), .ZN(
        n22591) );
  NAND3_X1 U5634 ( .A1(n15391), .A2(n22873), .A3(n15390), .ZN(n393) );
  BUF_X2 U5647 ( .I(n849), .Z(n30437) );
  NAND2_X1 U5659 ( .A1(n31363), .A2(n10288), .ZN(n6540) );
  NAND2_X1 U5666 ( .A1(n31315), .A2(n22680), .ZN(n4156) );
  CLKBUF_X2 U5699 ( .I(n9953), .Z(n31019) );
  BUF_X2 U5705 ( .I(n27160), .Z(n22524) );
  CLKBUF_X4 U5712 ( .I(n11110), .Z(n29335) );
  INV_X1 U5720 ( .I(n22213), .ZN(n31331) );
  OAI21_X1 U5723 ( .A1(n29408), .A2(n21475), .B(n21936), .ZN(n21481) );
  AND2_X1 U5726 ( .A1(n21477), .A2(n28895), .Z(n29408) );
  NAND2_X1 U5729 ( .A1(n7813), .A2(n29796), .ZN(n30622) );
  NOR2_X1 U5732 ( .A1(n29433), .A2(n29943), .ZN(n3908) );
  NOR2_X1 U5734 ( .A1(n21785), .A2(n7553), .ZN(n30374) );
  CLKBUF_X4 U5741 ( .I(n1917), .Z(n31616) );
  NOR2_X1 U5758 ( .A1(n21282), .A2(n28618), .ZN(n31073) );
  NAND2_X1 U5759 ( .A1(n31557), .A2(n31458), .ZN(n31572) );
  NOR2_X1 U5760 ( .A1(n9601), .A2(n13213), .ZN(n13212) );
  NAND2_X1 U5764 ( .A1(n21278), .A2(n29827), .ZN(n21279) );
  INV_X2 U5767 ( .I(n5863), .ZN(n7813) );
  NAND2_X1 U5768 ( .A1(n21), .A2(n30033), .ZN(n21539) );
  CLKBUF_X2 U5774 ( .I(n12535), .Z(n30243) );
  NAND2_X1 U5776 ( .A1(n12725), .A2(n31334), .ZN(n12724) );
  CLKBUF_X4 U5779 ( .I(n6533), .Z(n31765) );
  INV_X1 U5819 ( .I(n31484), .ZN(n16925) );
  INV_X1 U5821 ( .I(n2802), .ZN(n29931) );
  AND3_X1 U5822 ( .A1(n21733), .A2(n26474), .A3(n13872), .Z(n29433) );
  NAND2_X1 U5824 ( .A1(n16257), .A2(n16258), .ZN(n29711) );
  INV_X1 U5836 ( .I(n21316), .ZN(n14230) );
  OAI21_X1 U5844 ( .A1(n12325), .A2(n3933), .B(n21400), .ZN(n15113) );
  NOR2_X1 U5852 ( .A1(n6277), .A2(n21302), .ZN(n18207) );
  NAND2_X1 U5853 ( .A1(n21167), .A2(n16905), .ZN(n30005) );
  INV_X1 U5854 ( .I(n20880), .ZN(n30006) );
  NAND2_X1 U5857 ( .A1(n1334), .A2(n31476), .ZN(n31475) );
  BUF_X2 U5871 ( .I(n3106), .Z(n26635) );
  NAND2_X1 U5874 ( .A1(n17439), .A2(n925), .ZN(n1785) );
  INV_X1 U5880 ( .I(n20972), .ZN(n29810) );
  BUF_X2 U5884 ( .I(n21220), .Z(n15149) );
  INV_X1 U5890 ( .I(n2756), .ZN(n29833) );
  INV_X1 U5891 ( .I(n20978), .ZN(n31235) );
  CLKBUF_X2 U5919 ( .I(n8728), .Z(n29838) );
  OR2_X1 U5926 ( .A1(n20247), .A2(n7394), .Z(n1684) );
  NOR2_X1 U5932 ( .A1(n30915), .A2(n20317), .ZN(n17732) );
  NOR2_X1 U5934 ( .A1(n30414), .A2(n30413), .ZN(n20282) );
  INV_X1 U5937 ( .I(n1354), .ZN(n31470) );
  INV_X1 U5938 ( .I(n931), .ZN(n30545) );
  CLKBUF_X2 U5945 ( .I(n6531), .Z(n31863) );
  CLKBUF_X2 U5947 ( .I(n9115), .Z(n30878) );
  CLKBUF_X2 U5951 ( .I(n4693), .Z(n31873) );
  INV_X2 U5952 ( .I(n6996), .ZN(n16182) );
  CLKBUF_X2 U5998 ( .I(n19849), .Z(n31742) );
  CLKBUF_X4 U6016 ( .I(n17711), .Z(n30355) );
  INV_X4 U6019 ( .I(n29882), .ZN(n20010) );
  CLKBUF_X2 U6041 ( .I(n19389), .Z(n31410) );
  NAND2_X1 U6043 ( .A1(n30710), .A2(n3341), .ZN(n19239) );
  NOR2_X1 U6044 ( .A1(n19011), .A2(n7995), .ZN(n30401) );
  INV_X1 U6045 ( .I(n19205), .ZN(n9316) );
  BUF_X2 U6061 ( .I(n11477), .Z(n4210) );
  BUF_X4 U6063 ( .I(n13320), .Z(n25968) );
  AOI21_X1 U6069 ( .A1(n12132), .A2(n18701), .B(n29366), .ZN(n8551) );
  INV_X1 U6071 ( .I(n18462), .ZN(n31903) );
  OAI21_X1 U6076 ( .A1(n17478), .A2(n31428), .B(n31427), .ZN(n12116) );
  OAI21_X1 U6082 ( .A1(n8411), .A2(n16614), .B(n18307), .ZN(n30866) );
  INV_X1 U6085 ( .I(n9836), .ZN(n18338) );
  NAND3_X1 U6092 ( .A1(n3152), .A2(n2990), .A3(n18893), .ZN(n30919) );
  CLKBUF_X2 U6095 ( .I(n18018), .Z(n31115) );
  INV_X1 U6102 ( .I(n24966), .ZN(n30881) );
  INV_X1 U6110 ( .I(n24923), .ZN(n31513) );
  BUF_X2 U6117 ( .I(n18557), .Z(n28987) );
  INV_X1 U6124 ( .I(n25450), .ZN(n29851) );
  INV_X1 U6130 ( .I(n16520), .ZN(n30557) );
  CLKBUF_X2 U6132 ( .I(n8317), .Z(n31724) );
  INV_X1 U6136 ( .I(n25195), .ZN(n30954) );
  INV_X1 U6137 ( .I(n16653), .ZN(n30018) );
  NAND2_X1 U6163 ( .A1(n18730), .A2(n18846), .ZN(n6313) );
  OAI21_X1 U6164 ( .A1(n16370), .A2(n962), .B(n6783), .ZN(n12199) );
  NAND2_X1 U6165 ( .A1(n1186), .A2(n18822), .ZN(n16247) );
  NOR2_X1 U6183 ( .A1(n18835), .A2(n32901), .ZN(n13013) );
  NOR2_X1 U6195 ( .A1(n10578), .A2(n11941), .ZN(n2734) );
  BUF_X2 U6201 ( .I(n16766), .Z(n28238) );
  INV_X1 U6205 ( .I(n7320), .ZN(n9174) );
  CLKBUF_X2 U6224 ( .I(n29061), .Z(n28548) );
  INV_X1 U6227 ( .I(n9514), .ZN(n17792) );
  NAND2_X1 U6228 ( .A1(n18792), .A2(n13514), .ZN(n29684) );
  NAND2_X1 U6240 ( .A1(n19315), .A2(n11000), .ZN(n10999) );
  NOR2_X1 U6241 ( .A1(n10857), .A2(n13568), .ZN(n10856) );
  INV_X2 U6246 ( .I(n19154), .ZN(n2040) );
  NAND2_X1 U6247 ( .A1(n7415), .A2(n14332), .ZN(n19247) );
  CLKBUF_X2 U6271 ( .I(n7134), .Z(n1386) );
  INV_X2 U6273 ( .I(n27807), .ZN(n26518) );
  NAND2_X1 U6274 ( .A1(n27077), .A2(n5789), .ZN(n19210) );
  INV_X1 U6277 ( .I(n6488), .ZN(n1367) );
  INV_X1 U6280 ( .I(n16429), .ZN(n31750) );
  NAND2_X1 U6281 ( .A1(n19190), .A2(n19261), .ZN(n28540) );
  NAND2_X1 U6289 ( .A1(n15239), .A2(n19218), .ZN(n19352) );
  OAI21_X1 U6297 ( .A1(n1630), .A2(n19176), .B(n12993), .ZN(n1629) );
  AOI21_X1 U6300 ( .A1(n18908), .A2(n26181), .B(n16353), .ZN(n18909) );
  INV_X1 U6304 ( .I(n2499), .ZN(n29727) );
  INV_X1 U6306 ( .I(n19343), .ZN(n30258) );
  INV_X1 U6307 ( .I(n15913), .ZN(n17220) );
  NAND2_X1 U6317 ( .A1(n20000), .A2(n14457), .ZN(n13654) );
  NAND2_X1 U6325 ( .A1(n1043), .A2(n11350), .ZN(n5642) );
  CLKBUF_X2 U6327 ( .I(n20011), .Z(n30794) );
  INV_X1 U6328 ( .I(n30600), .ZN(n8687) );
  OAI21_X1 U6336 ( .A1(n15192), .A2(n19874), .B(n149), .ZN(n12669) );
  NAND2_X1 U6357 ( .A1(n29373), .A2(n31694), .ZN(n31693) );
  NAND2_X1 U6358 ( .A1(n28021), .A2(n20068), .ZN(n28020) );
  NAND2_X1 U6371 ( .A1(n5999), .A2(n20033), .ZN(n4201) );
  NAND2_X1 U6379 ( .A1(n20017), .A2(n15278), .ZN(n30072) );
  INV_X1 U6388 ( .I(n20107), .ZN(n31164) );
  OAI21_X1 U6395 ( .A1(n19808), .A2(n15278), .B(n8816), .ZN(n10742) );
  NAND2_X1 U6396 ( .A1(n20090), .A2(n19879), .ZN(n19881) );
  INV_X2 U6398 ( .I(n34151), .ZN(n729) );
  NAND2_X1 U6423 ( .A1(n15953), .A2(n9484), .ZN(n30464) );
  CLKBUF_X2 U6429 ( .I(n10414), .Z(n3915) );
  NAND3_X1 U6432 ( .A1(n2879), .A2(n31504), .A3(n20524), .ZN(n31563) );
  AND2_X1 U6433 ( .A1(n17647), .A2(n6230), .Z(n29409) );
  NAND2_X1 U6437 ( .A1(n28288), .A2(n6997), .ZN(n7056) );
  INV_X1 U6440 ( .I(n20536), .ZN(n20535) );
  AOI21_X1 U6442 ( .A1(n33288), .A2(n20472), .B(n32504), .ZN(n20165) );
  INV_X2 U6446 ( .I(n8903), .ZN(n1349) );
  NAND2_X1 U6450 ( .A1(n9115), .A2(n6996), .ZN(n12583) );
  NAND2_X1 U6452 ( .A1(n8702), .A2(n9854), .ZN(n31496) );
  OAI21_X1 U6453 ( .A1(n818), .A2(n710), .B(n20334), .ZN(n20048) );
  NOR2_X1 U6454 ( .A1(n10718), .A2(n10716), .ZN(n10715) );
  NAND2_X1 U6456 ( .A1(n32068), .A2(n20452), .ZN(n15662) );
  OAI21_X1 U6468 ( .A1(n1160), .A2(n27621), .B(n27620), .ZN(n2754) );
  INV_X1 U6478 ( .I(n20863), .ZN(n29734) );
  NOR2_X1 U6490 ( .A1(n21060), .A2(n4568), .ZN(n10921) );
  NAND2_X1 U6491 ( .A1(n29255), .A2(n26712), .ZN(n6337) );
  NAND2_X1 U6493 ( .A1(n21203), .A2(n3933), .ZN(n21204) );
  INV_X1 U6495 ( .I(n29802), .ZN(n13700) );
  AND2_X1 U6496 ( .A1(n4145), .A2(n32452), .Z(n29361) );
  NAND2_X1 U6502 ( .A1(n8197), .A2(n924), .ZN(n1555) );
  INV_X1 U6505 ( .I(n31197), .ZN(n30816) );
  NOR2_X1 U6510 ( .A1(n21113), .A2(n1332), .ZN(n27539) );
  NOR2_X1 U6516 ( .A1(n18218), .A2(n31030), .ZN(n7845) );
  NAND2_X1 U6523 ( .A1(n14721), .A2(n8115), .ZN(n14087) );
  NAND3_X1 U6524 ( .A1(n20883), .A2(n21369), .A3(n1148), .ZN(n20884) );
  NOR2_X1 U6531 ( .A1(n21358), .A2(n11814), .ZN(n6307) );
  NAND2_X1 U6541 ( .A1(n21211), .A2(n13319), .ZN(n20874) );
  NAND2_X1 U6547 ( .A1(n30227), .A2(n30226), .ZN(n30225) );
  INV_X1 U6552 ( .I(n21147), .ZN(n17217) );
  NOR2_X1 U6561 ( .A1(n3140), .A2(n30885), .ZN(n27836) );
  AOI21_X1 U6562 ( .A1(n16755), .A2(n27955), .B(n21400), .ZN(n16257) );
  NAND2_X1 U6563 ( .A1(n4293), .A2(n31613), .ZN(n31612) );
  AOI21_X1 U6565 ( .A1(n30006), .A2(n30005), .B(n21209), .ZN(n29214) );
  INV_X1 U6572 ( .I(n11861), .ZN(n31653) );
  AOI21_X1 U6578 ( .A1(n10345), .A2(n16519), .B(n777), .ZN(n10344) );
  INV_X1 U6579 ( .I(n16605), .ZN(n30007) );
  INV_X1 U6597 ( .I(n2576), .ZN(n21682) );
  NAND2_X1 U6601 ( .A1(n31475), .A2(n31474), .ZN(n21274) );
  INV_X2 U6603 ( .I(n5795), .ZN(n1135) );
  NAND2_X1 U6617 ( .A1(n18055), .A2(n21), .ZN(n30608) );
  OAI21_X1 U6634 ( .A1(n21696), .A2(n30769), .B(n1013), .ZN(n21699) );
  NAND2_X1 U6651 ( .A1(n15748), .A2(n26513), .ZN(n10232) );
  INV_X1 U6663 ( .I(n10519), .ZN(n22244) );
  INV_X2 U6664 ( .I(n22092), .ZN(n14289) );
  INV_X1 U6671 ( .I(n1716), .ZN(n29896) );
  OAI21_X1 U6674 ( .A1(n13371), .A2(n22220), .B(n13370), .ZN(n22246) );
  INV_X1 U6695 ( .I(n22565), .ZN(n22468) );
  NOR3_X1 U6696 ( .A1(n22543), .A2(n10757), .A3(n252), .ZN(n7236) );
  CLKBUF_X4 U6716 ( .I(n632), .Z(n14227) );
  NOR2_X1 U6730 ( .A1(n22682), .A2(n9802), .ZN(n3455) );
  NAND3_X1 U6732 ( .A1(n900), .A2(n11920), .A3(n22476), .ZN(n14017) );
  NAND2_X1 U6744 ( .A1(n29335), .A2(n22435), .ZN(n31634) );
  NOR2_X1 U6748 ( .A1(n16986), .A2(n9370), .ZN(n22026) );
  OAI21_X1 U6750 ( .A1(n29461), .A2(n15635), .B(n29222), .ZN(n28894) );
  NOR2_X1 U6753 ( .A1(n29508), .A2(n22574), .ZN(n10121) );
  INV_X1 U6769 ( .I(n22560), .ZN(n31315) );
  AOI22_X1 U6781 ( .A1(n12281), .A2(n10288), .B1(n22542), .B2(n22397), .ZN(
        n22299) );
  NAND3_X1 U6791 ( .A1(n29222), .A2(n18073), .A3(n10680), .ZN(n12472) );
  NAND2_X1 U6793 ( .A1(n15033), .A2(n8314), .ZN(n15032) );
  INV_X2 U6797 ( .I(n7004), .ZN(n14131) );
  NAND2_X1 U6808 ( .A1(n2635), .A2(n13191), .ZN(n2638) );
  NAND2_X1 U6818 ( .A1(n14131), .A2(n23106), .ZN(n15280) );
  OAI22_X1 U6835 ( .A1(n22502), .A2(n32449), .B1(n13874), .B2(n30014), .ZN(
        n26772) );
  NAND3_X1 U6847 ( .A1(n29610), .A2(n4113), .A3(n22791), .ZN(n22776) );
  AOI21_X1 U6848 ( .A1(n3783), .A2(n28801), .B(n30247), .ZN(n9075) );
  INV_X1 U6852 ( .I(n9185), .ZN(n31056) );
  CLKBUF_X2 U6857 ( .I(n8762), .Z(n29235) );
  INV_X1 U6863 ( .I(n14464), .ZN(n29675) );
  INV_X1 U6864 ( .I(n23331), .ZN(n23509) );
  NAND2_X1 U6866 ( .A1(n23873), .A2(n23872), .ZN(n23874) );
  AOI21_X1 U6867 ( .A1(n27298), .A2(n8967), .B(n22957), .ZN(n22904) );
  INV_X1 U6869 ( .I(n23742), .ZN(n23768) );
  INV_X1 U6877 ( .I(n23778), .ZN(n975) );
  INV_X1 U6883 ( .I(n8045), .ZN(n11960) );
  NAND2_X1 U6884 ( .A1(n1252), .A2(n23603), .ZN(n14039) );
  NOR2_X1 U6886 ( .A1(n23611), .A2(n33144), .ZN(n1892) );
  NAND2_X1 U6887 ( .A1(n23647), .A2(n26790), .ZN(n28303) );
  INV_X1 U6891 ( .I(n28615), .ZN(n23691) );
  INV_X2 U6896 ( .I(n9828), .ZN(n16686) );
  CLKBUF_X2 U6900 ( .I(n23924), .Z(n1101) );
  OAI21_X1 U6903 ( .A1(n15187), .A2(n15186), .B(n23691), .ZN(n23572) );
  NAND3_X1 U6907 ( .A1(n23799), .A2(n23798), .A3(n23800), .ZN(n23802) );
  NAND2_X1 U6908 ( .A1(n23855), .A2(n652), .ZN(n23856) );
  INV_X2 U6912 ( .I(n23603), .ZN(n23776) );
  NAND2_X1 U6923 ( .A1(n793), .A2(n6713), .ZN(n5132) );
  AND2_X1 U6928 ( .A1(n11438), .A2(n29748), .Z(n29379) );
  NAND2_X1 U6936 ( .A1(n23707), .A2(n23786), .ZN(n23711) );
  NOR2_X1 U6947 ( .A1(n30283), .A2(n24087), .ZN(n11107) );
  OAI22_X1 U6964 ( .A1(n7068), .A2(n24196), .B1(n13048), .B2(n969), .ZN(n13324) );
  AND2_X1 U6972 ( .A1(n24234), .A2(n7581), .Z(n8004) );
  CLKBUF_X4 U6978 ( .I(n13508), .Z(n7828) );
  INV_X1 U6981 ( .I(n14897), .ZN(n1226) );
  INV_X1 U6988 ( .I(n24427), .ZN(n29639) );
  NAND2_X1 U6992 ( .A1(n16113), .A2(n25870), .ZN(n24732) );
  CLKBUF_X4 U7006 ( .I(n16757), .Z(n11090) );
  NAND2_X1 U7011 ( .A1(n26917), .A2(n15770), .ZN(n25396) );
  NAND2_X1 U7015 ( .A1(n25870), .A2(n4993), .ZN(n11718) );
  NAND2_X1 U7023 ( .A1(n419), .A2(n11366), .ZN(n16339) );
  AOI21_X1 U7027 ( .A1(n24955), .A2(n24956), .B(n24947), .ZN(n29664) );
  OAI21_X1 U7029 ( .A1(n25204), .A2(n32601), .B(n25205), .ZN(n18259) );
  CLKBUF_X1 U7031 ( .I(n11974), .Z(n4245) );
  INV_X1 U7034 ( .I(n29664), .ZN(n29663) );
  CLKBUF_X1 U7056 ( .I(n25258), .Z(n27429) );
  INV_X2 U7060 ( .I(n5128), .ZN(n786) );
  CLKBUF_X1 U7062 ( .I(Key[158]), .Z(n16705) );
  XNOR2_X1 U7071 ( .A1(n5150), .A2(n14648), .ZN(n29341) );
  XNOR2_X1 U7074 ( .A1(n19580), .A2(n32796), .ZN(n29343) );
  XNOR2_X1 U7075 ( .A1(n23271), .A2(n16653), .ZN(n29344) );
  XNOR2_X1 U7084 ( .A1(n27423), .A2(n25108), .ZN(n29345) );
  XNOR2_X1 U7086 ( .A1(n24635), .A2(n16654), .ZN(n29346) );
  XNOR2_X1 U7087 ( .A1(n16237), .A2(n28711), .ZN(n29347) );
  XNOR2_X1 U7088 ( .A1(n24617), .A2(n25735), .ZN(n29348) );
  OR2_X1 U7089 ( .A1(n32021), .A2(n31551), .Z(n29349) );
  AND2_X1 U7092 ( .A1(n24293), .A2(n5632), .Z(n29352) );
  AND2_X1 U7096 ( .A1(n14980), .A2(n31721), .Z(n29354) );
  OR2_X1 U7103 ( .A1(n28293), .A2(n1170), .Z(n29359) );
  AND2_X1 U7112 ( .A1(n20263), .A2(n16146), .Z(n29363) );
  AND2_X1 U7113 ( .A1(n3791), .A2(n6034), .Z(n29364) );
  OR2_X1 U7120 ( .A1(n17694), .A2(n11968), .Z(n29367) );
  OR2_X2 U7132 ( .A1(n28197), .A2(n33232), .Z(n29378) );
  OR2_X1 U7136 ( .A1(n28669), .A2(n10206), .Z(n29380) );
  AND2_X1 U7140 ( .A1(n21779), .A2(n31654), .Z(n29383) );
  OR2_X1 U7144 ( .A1(n26547), .A2(n1596), .Z(n29385) );
  XNOR2_X1 U7149 ( .A1(n24598), .A2(n29416), .ZN(n29386) );
  OR2_X1 U7153 ( .A1(n28833), .A2(n5615), .Z(n29389) );
  OR2_X1 U7155 ( .A1(n22659), .A2(n22658), .Z(n29390) );
  AND2_X1 U7160 ( .A1(n28801), .A2(n11235), .Z(n29391) );
  AND3_X1 U7161 ( .A1(n6012), .A2(n16254), .A3(n23110), .Z(n29392) );
  AND2_X1 U7163 ( .A1(n17077), .A2(n21579), .Z(n29393) );
  INV_X1 U7176 ( .I(n3106), .ZN(n4971) );
  XNOR2_X1 U7183 ( .A1(n17586), .A2(n12082), .ZN(n29400) );
  INV_X1 U7190 ( .I(n10124), .ZN(n29730) );
  AND2_X1 U7191 ( .A1(n24436), .A2(n25695), .Z(n29402) );
  OR3_X2 U7192 ( .A1(n7753), .A2(n26622), .A3(n15414), .Z(n29404) );
  AND2_X1 U7194 ( .A1(n15465), .A2(n21866), .Z(n29405) );
  INV_X1 U7196 ( .I(n19283), .ZN(n30932) );
  XNOR2_X1 U7201 ( .A1(n20885), .A2(n25716), .ZN(n29412) );
  XNOR2_X1 U7202 ( .A1(n21043), .A2(n30007), .ZN(n29413) );
  XNOR2_X1 U7212 ( .A1(n34150), .A2(n16533), .ZN(n29415) );
  XNOR2_X1 U7221 ( .A1(n24616), .A2(n24907), .ZN(n29416) );
  XNOR2_X1 U7222 ( .A1(n27167), .A2(n16653), .ZN(n29417) );
  XNOR2_X1 U7223 ( .A1(n34150), .A2(n24065), .ZN(n29418) );
  XNOR2_X1 U7225 ( .A1(n23153), .A2(n14464), .ZN(n29420) );
  AND2_X1 U7229 ( .A1(n17828), .A2(n26160), .Z(n29421) );
  XNOR2_X1 U7241 ( .A1(n19651), .A2(n19658), .ZN(n29426) );
  XNOR2_X1 U7242 ( .A1(n8497), .A2(n513), .ZN(n29428) );
  INV_X2 U7251 ( .I(n16132), .ZN(n15213) );
  XNOR2_X1 U7256 ( .A1(n19727), .A2(n18814), .ZN(n29441) );
  XNOR2_X1 U7257 ( .A1(n34082), .A2(n25560), .ZN(n29442) );
  INV_X1 U7261 ( .I(n18199), .ZN(n19900) );
  XNOR2_X1 U7267 ( .A1(n4107), .A2(n27361), .ZN(n29443) );
  XNOR2_X1 U7281 ( .A1(n9102), .A2(n9101), .ZN(n29445) );
  XNOR2_X1 U7288 ( .A1(n3665), .A2(n5920), .ZN(n29446) );
  XNOR2_X1 U7289 ( .A1(n10224), .A2(n1365), .ZN(n29447) );
  OR2_X1 U7290 ( .A1(n19226), .A2(n19227), .Z(n29448) );
  XOR2_X1 U7293 ( .A1(n21916), .A2(n21915), .Z(n29450) );
  XOR2_X1 U7294 ( .A1(n30070), .A2(n22094), .Z(n29451) );
  AND2_X2 U7300 ( .A1(n6357), .A2(n9999), .Z(n29454) );
  XNOR2_X1 U7306 ( .A1(n22076), .A2(n24937), .ZN(n29457) );
  XNOR2_X1 U7310 ( .A1(n22154), .A2(n22152), .ZN(n29458) );
  INV_X1 U7316 ( .I(n27160), .ZN(n28915) );
  NOR2_X1 U7318 ( .A1(n632), .A2(n22662), .ZN(n29461) );
  XNOR2_X1 U7324 ( .A1(n2899), .A2(n2898), .ZN(n29463) );
  OR2_X1 U7325 ( .A1(n8381), .A2(n5211), .Z(n29464) );
  XNOR2_X1 U7328 ( .A1(n11427), .A2(n11426), .ZN(n29467) );
  INV_X1 U7334 ( .I(n12375), .ZN(n808) );
  CLKBUF_X2 U7337 ( .I(n16536), .Z(n6479) );
  AND2_X1 U7340 ( .A1(n17394), .A2(n13318), .Z(n29469) );
  INV_X1 U7351 ( .I(n5736), .ZN(n13281) );
  XOR2_X1 U7352 ( .A1(n281), .A2(n15515), .Z(n29472) );
  NOR2_X1 U7363 ( .A1(n2855), .A2(n23767), .ZN(n29474) );
  XNOR2_X1 U7364 ( .A1(n24819), .A2(n24632), .ZN(n29475) );
  CLKBUF_X2 U7366 ( .I(n24975), .Z(n31274) );
  NAND2_X1 U7373 ( .A1(n10430), .A2(n27072), .ZN(n29476) );
  NAND2_X2 U7376 ( .A1(n2550), .A2(n6409), .ZN(n11557) );
  NOR2_X1 U7377 ( .A1(n4135), .A2(n29325), .ZN(n29477) );
  XOR2_X1 U7379 ( .A1(n19726), .A2(n12718), .Z(n29487) );
  INV_X2 U7387 ( .I(n28196), .ZN(n7765) );
  NAND2_X2 U7397 ( .A1(n25170), .A2(n25168), .ZN(n28196) );
  XOR2_X1 U7406 ( .A1(n11423), .A2(n11421), .Z(n11451) );
  NOR3_X1 U7408 ( .A1(n21865), .A2(n21738), .A3(n13652), .ZN(n30806) );
  OAI21_X2 U7414 ( .A1(n29358), .A2(n29480), .B(n8927), .ZN(n9097) );
  INV_X1 U7416 ( .I(n576), .ZN(n29480) );
  INV_X2 U7419 ( .I(n33373), .ZN(n29481) );
  NOR3_X1 U7430 ( .A1(n11516), .A2(n9430), .A3(n7993), .ZN(n5777) );
  XOR2_X1 U7435 ( .A1(n5431), .A2(n30171), .Z(n29482) );
  INV_X4 U7436 ( .I(n29483), .ZN(n9677) );
  NOR2_X2 U7437 ( .A1(n10842), .A2(n4267), .ZN(n29483) );
  NAND2_X1 U7443 ( .A1(n896), .A2(n23045), .ZN(n22400) );
  NAND3_X1 U7447 ( .A1(n9962), .A2(n10033), .A3(n24311), .ZN(n12318) );
  OAI21_X2 U7452 ( .A1(n29654), .A2(n30233), .B(n31960), .ZN(n6123) );
  NOR3_X2 U7460 ( .A1(n11411), .A2(n2085), .A3(n2084), .ZN(n23306) );
  XOR2_X1 U7462 ( .A1(n29485), .A2(n24486), .Z(n31005) );
  XOR2_X1 U7464 ( .A1(n24488), .A2(n24771), .Z(n29485) );
  XOR2_X1 U7465 ( .A1(n7537), .A2(n24603), .Z(n28144) );
  XOR2_X1 U7482 ( .A1(n27977), .A2(n24564), .Z(n17673) );
  OR2_X1 U7483 ( .A1(n23086), .A2(n4834), .Z(n4833) );
  XOR2_X1 U7488 ( .A1(n29486), .A2(n29487), .Z(n8327) );
  NAND2_X2 U7496 ( .A1(n29488), .A2(n28875), .ZN(n25653) );
  OAI21_X2 U7499 ( .A1(n15355), .A2(n15354), .B(n25706), .ZN(n29488) );
  XOR2_X1 U7506 ( .A1(n29489), .A2(n4761), .Z(n8553) );
  XOR2_X1 U7507 ( .A1(n10087), .A2(n28868), .Z(n29489) );
  XOR2_X1 U7514 ( .A1(n24635), .A2(n10146), .Z(n17448) );
  NOR2_X2 U7515 ( .A1(n7480), .A2(n7483), .ZN(n24635) );
  NAND2_X2 U7518 ( .A1(n13341), .A2(n28356), .ZN(n28355) );
  NAND2_X1 U7519 ( .A1(n26325), .A2(n1318), .ZN(n26927) );
  XOR2_X1 U7521 ( .A1(n7694), .A2(n7693), .Z(n29543) );
  XOR2_X1 U7531 ( .A1(n8714), .A2(n8265), .Z(n8713) );
  XOR2_X1 U7534 ( .A1(n6513), .A2(n9385), .Z(n9564) );
  NOR2_X1 U7549 ( .A1(n29792), .A2(n20549), .ZN(n31232) );
  NAND2_X2 U7557 ( .A1(n11466), .A2(n22783), .ZN(n8226) );
  OAI21_X1 U7569 ( .A1(n22558), .A2(n9630), .B(n29495), .ZN(n29494) );
  INV_X2 U7570 ( .I(n994), .ZN(n29495) );
  INV_X1 U7576 ( .I(n32957), .ZN(n29497) );
  INV_X2 U7577 ( .I(n15365), .ZN(n29498) );
  OR2_X1 U7579 ( .A1(n596), .A2(n14290), .Z(n14562) );
  XOR2_X1 U7583 ( .A1(n14727), .A2(n25549), .Z(n31093) );
  NAND2_X2 U7593 ( .A1(n13633), .A2(n13632), .ZN(n14727) );
  NAND2_X2 U7617 ( .A1(n2394), .A2(n2393), .ZN(n22102) );
  NAND2_X1 U7677 ( .A1(n14661), .A2(n29213), .ZN(n19889) );
  NAND2_X1 U7680 ( .A1(n12042), .A2(n32875), .ZN(n24863) );
  XOR2_X1 U7700 ( .A1(n16886), .A2(n16887), .Z(n23156) );
  OR2_X1 U7711 ( .A1(n9411), .A2(n30668), .Z(n7488) );
  NAND2_X2 U7722 ( .A1(n30856), .A2(n9803), .ZN(n20715) );
  NOR2_X2 U7739 ( .A1(n6533), .A2(n28429), .ZN(n16736) );
  NAND2_X2 U7744 ( .A1(n30483), .A2(n21216), .ZN(n6533) );
  NAND2_X2 U7745 ( .A1(n30139), .A2(n30138), .ZN(n20536) );
  NAND2_X2 U7749 ( .A1(n32075), .A2(n31734), .ZN(n21866) );
  NAND2_X2 U7756 ( .A1(n5743), .A2(n29508), .ZN(n29507) );
  NOR2_X1 U7759 ( .A1(n30666), .A2(n14803), .ZN(n29510) );
  OAI21_X2 U7763 ( .A1(n28510), .A2(n11240), .B(n29509), .ZN(n17580) );
  NAND2_X1 U7764 ( .A1(n10673), .A2(n499), .ZN(n29509) );
  NAND2_X2 U7787 ( .A1(n9123), .A2(n31573), .ZN(n4704) );
  XOR2_X1 U7821 ( .A1(n23504), .A2(n23164), .Z(n14370) );
  NAND2_X1 U7828 ( .A1(n31815), .A2(n21289), .ZN(n21291) );
  NOR2_X1 U7837 ( .A1(n5273), .A2(n17814), .ZN(n4204) );
  NAND2_X1 U7841 ( .A1(n27320), .A2(n27321), .ZN(n29517) );
  NAND2_X2 U7847 ( .A1(n17579), .A2(n16388), .ZN(n29518) );
  XOR2_X1 U7862 ( .A1(n22896), .A2(n23126), .Z(n14154) );
  NAND2_X2 U7867 ( .A1(n30705), .A2(n20163), .ZN(n20720) );
  OR2_X1 U7876 ( .A1(n17405), .A2(n16996), .Z(n11508) );
  OAI21_X2 U7877 ( .A1(n23158), .A2(n22914), .B(n29522), .ZN(n14613) );
  NOR2_X2 U7879 ( .A1(n8943), .A2(n6382), .ZN(n29522) );
  NOR2_X2 U7880 ( .A1(n1350), .A2(n15434), .ZN(n29586) );
  NOR2_X2 U7888 ( .A1(n9962), .A2(n27501), .ZN(n15283) );
  NOR2_X1 U7891 ( .A1(n29714), .A2(n8314), .ZN(n13770) );
  BUF_X2 U7895 ( .I(n19049), .Z(n29525) );
  NOR3_X2 U7896 ( .A1(n8378), .A2(n12925), .A3(n21430), .ZN(n7666) );
  NAND2_X2 U7899 ( .A1(n24461), .A2(n29526), .ZN(n31656) );
  NAND3_X2 U7901 ( .A1(n27118), .A2(n1223), .A3(n18219), .ZN(n29526) );
  NAND2_X2 U7903 ( .A1(n29527), .A2(n30938), .ZN(n16831) );
  XOR2_X1 U7911 ( .A1(n19476), .A2(n19575), .Z(n11093) );
  OR2_X1 U7915 ( .A1(n29213), .A2(n14661), .Z(n4938) );
  XOR2_X1 U7916 ( .A1(n24826), .A2(n7879), .Z(n29534) );
  XOR2_X1 U7920 ( .A1(n12413), .A2(n19490), .Z(n9528) );
  XOR2_X1 U7921 ( .A1(n19746), .A2(n12442), .Z(n19490) );
  XOR2_X1 U7936 ( .A1(n24090), .A2(n29531), .Z(n28816) );
  XOR2_X1 U7940 ( .A1(n24419), .A2(n29639), .Z(n29531) );
  OAI21_X2 U7943 ( .A1(n15673), .A2(n15672), .B(n29532), .ZN(n10371) );
  NAND2_X2 U7956 ( .A1(n30953), .A2(n25874), .ZN(n14737) );
  OAI22_X1 U7958 ( .A1(n790), .A2(n25900), .B1(n25867), .B2(n27118), .ZN(
        n25899) );
  XOR2_X1 U7970 ( .A1(n24807), .A2(n28939), .Z(n24439) );
  AOI22_X1 U7974 ( .A1(n4417), .A2(n25743), .B1(n9414), .B2(n4416), .ZN(n29572) );
  XOR2_X1 U7975 ( .A1(n29534), .A2(n33927), .Z(n26125) );
  XOR2_X1 U7986 ( .A1(n30767), .A2(n7071), .Z(n7825) );
  XOR2_X1 U7987 ( .A1(n29536), .A2(n22303), .Z(n21927) );
  NAND2_X2 U7989 ( .A1(n21589), .A2(n21588), .ZN(n22303) );
  INV_X2 U7990 ( .I(n13553), .ZN(n29536) );
  AOI22_X2 U7997 ( .A1(n23850), .A2(n32477), .B1(n23847), .B2(n23809), .ZN(
        n3239) );
  INV_X2 U7998 ( .I(n29537), .ZN(n10435) );
  XNOR2_X1 U8002 ( .A1(n26854), .A2(n2064), .ZN(n29537) );
  XOR2_X1 U8009 ( .A1(n29538), .A2(n24824), .Z(n31598) );
  CLKBUF_X12 U8019 ( .I(n10248), .Z(n29539) );
  NOR2_X2 U8030 ( .A1(n709), .A2(n31953), .ZN(n14794) );
  INV_X4 U8032 ( .I(n10435), .ZN(n15278) );
  OR2_X1 U8040 ( .A1(n33981), .A2(n21832), .Z(n10401) );
  NAND3_X1 U8063 ( .A1(n15146), .A2(n1063), .A3(n1185), .ZN(n9886) );
  OAI21_X1 U8064 ( .A1(n17497), .A2(n30099), .B(n5781), .ZN(n15929) );
  NOR2_X2 U8066 ( .A1(n6610), .A2(n20209), .ZN(n30099) );
  NOR2_X2 U8074 ( .A1(n12433), .A2(n23753), .ZN(n6363) );
  NAND3_X1 U8090 ( .A1(n31924), .A2(n29013), .A3(n4744), .ZN(n26958) );
  XOR2_X1 U8096 ( .A1(n2142), .A2(n17040), .Z(n2143) );
  XOR2_X1 U8098 ( .A1(n6386), .A2(n17052), .Z(n17040) );
  NAND2_X2 U8101 ( .A1(n8453), .A2(n164), .ZN(n7667) );
  XOR2_X1 U8133 ( .A1(n14136), .A2(n51), .Z(n3847) );
  XOR2_X1 U8140 ( .A1(n29545), .A2(n24699), .Z(n25385) );
  OAI21_X1 U8146 ( .A1(n13526), .A2(n18794), .B(n18793), .ZN(n9887) );
  NOR2_X2 U8152 ( .A1(n1898), .A2(n29548), .ZN(n1897) );
  XOR2_X1 U8169 ( .A1(n19568), .A2(n10552), .Z(n29550) );
  NAND3_X1 U8173 ( .A1(n4916), .A2(n22651), .A3(n14253), .ZN(n29551) );
  NAND2_X2 U8176 ( .A1(n30988), .A2(n11948), .ZN(n7226) );
  XOR2_X1 U8184 ( .A1(n27226), .A2(n29554), .Z(n10402) );
  XOR2_X1 U8188 ( .A1(n1971), .A2(n1905), .Z(n29554) );
  NOR2_X1 U8193 ( .A1(n20162), .A2(n20161), .ZN(n29725) );
  NOR2_X2 U8194 ( .A1(n18666), .A2(n29555), .ZN(n19308) );
  OAI22_X1 U8195 ( .A1(n2523), .A2(n18866), .B1(n18665), .B2(n711), .ZN(n29555) );
  NAND2_X2 U8199 ( .A1(n1008), .A2(n10699), .ZN(n21932) );
  AOI22_X2 U8202 ( .A1(n5252), .A2(n1265), .B1(n4777), .B2(n26612), .ZN(n4776)
         );
  NAND2_X2 U8204 ( .A1(n4780), .A2(n4779), .ZN(n4778) );
  NAND2_X2 U8205 ( .A1(n29557), .A2(n17718), .ZN(n30538) );
  XOR2_X1 U8223 ( .A1(n22109), .A2(n22111), .Z(n4797) );
  XOR2_X1 U8231 ( .A1(n29559), .A2(n27243), .Z(n31611) );
  XOR2_X1 U8232 ( .A1(n23262), .A2(n25049), .Z(n29559) );
  NOR2_X1 U8245 ( .A1(n19972), .A2(n20444), .ZN(n29560) );
  NAND2_X1 U8250 ( .A1(n10132), .A2(n23821), .ZN(n29561) );
  NAND2_X2 U8251 ( .A1(n29562), .A2(n30641), .ZN(n30640) );
  XOR2_X1 U8263 ( .A1(n20769), .A2(n1340), .Z(n20687) );
  NAND2_X2 U8269 ( .A1(n29563), .A2(n22436), .ZN(n8365) );
  XOR2_X1 U8276 ( .A1(n20839), .A2(n28813), .Z(n8855) );
  NAND3_X2 U8277 ( .A1(n29899), .A2(n20500), .A3(n16759), .ZN(n20839) );
  AOI22_X1 U8278 ( .A1(n10229), .A2(n19167), .B1(n25985), .B2(n10228), .ZN(
        n9711) );
  INV_X2 U8284 ( .I(n24339), .ZN(n24163) );
  NAND3_X2 U8285 ( .A1(n8720), .A2(n8719), .A3(n23780), .ZN(n24339) );
  XOR2_X1 U8323 ( .A1(n1044), .A2(n31138), .Z(n14223) );
  XOR2_X1 U8326 ( .A1(n29572), .A2(n1192), .Z(Ciphertext[156]) );
  NAND2_X2 U8327 ( .A1(n25846), .A2(n25844), .ZN(n27162) );
  NAND2_X2 U8332 ( .A1(n25838), .A2(n7143), .ZN(n25846) );
  NAND2_X1 U8342 ( .A1(n21132), .A2(n21442), .ZN(n29573) );
  XOR2_X1 U8370 ( .A1(n4949), .A2(n30463), .Z(n18048) );
  XOR2_X1 U8382 ( .A1(n2308), .A2(n22096), .Z(n22166) );
  OAI21_X1 U8393 ( .A1(n31144), .A2(n22377), .B(n31143), .ZN(n13535) );
  NAND3_X2 U8398 ( .A1(n11139), .A2(n11140), .A3(n20254), .ZN(n12459) );
  AOI21_X2 U8399 ( .A1(n25901), .A2(n25904), .B(n29578), .ZN(n26569) );
  NAND2_X2 U8400 ( .A1(n28455), .A2(n25902), .ZN(n29578) );
  XOR2_X1 U8402 ( .A1(n9781), .A2(n23264), .Z(n23311) );
  OAI22_X2 U8424 ( .A1(n18917), .A2(n18916), .B1(n13200), .B2(n19119), .ZN(
        n29581) );
  XOR2_X1 U8427 ( .A1(n9121), .A2(n29582), .Z(n9120) );
  XOR2_X1 U8429 ( .A1(n17705), .A2(n29475), .Z(n29582) );
  NOR2_X2 U8440 ( .A1(n29586), .A2(n16070), .ZN(n28802) );
  INV_X4 U8442 ( .I(n4834), .ZN(n23085) );
  NAND2_X1 U8446 ( .A1(n5673), .A2(n12593), .ZN(n5672) );
  INV_X4 U8447 ( .I(n23832), .ZN(n29965) );
  OAI21_X2 U8450 ( .A1(n22448), .A2(n1297), .B(n27886), .ZN(n14402) );
  XOR2_X1 U8455 ( .A1(n24492), .A2(n29588), .Z(n10841) );
  XOR2_X1 U8459 ( .A1(n28258), .A2(n12), .Z(n29588) );
  NOR2_X1 U8468 ( .A1(n11915), .A2(n8074), .ZN(n29743) );
  XOR2_X1 U8474 ( .A1(n19544), .A2(n19431), .Z(n18083) );
  NAND3_X1 U8477 ( .A1(n21316), .A2(n20330), .A3(n8115), .ZN(n16048) );
  INV_X2 U8524 ( .I(n10187), .ZN(n30360) );
  XOR2_X1 U8526 ( .A1(n29600), .A2(n15415), .Z(Ciphertext[17]) );
  AOI22_X1 U8528 ( .A1(n24961), .A2(n28662), .B1(n24958), .B2(n24959), .ZN(
        n29600) );
  OAI22_X2 U8532 ( .A1(n9842), .A2(n21335), .B1(n21337), .B2(n21336), .ZN(
        n8140) );
  BUF_X4 U8557 ( .I(n29268), .Z(n4991) );
  NOR2_X2 U8566 ( .A1(n9900), .A2(n9899), .ZN(n29606) );
  XOR2_X1 U8578 ( .A1(n23192), .A2(n23462), .Z(n29719) );
  NAND2_X2 U8579 ( .A1(n27008), .A2(n29607), .ZN(n9280) );
  OAI21_X2 U8582 ( .A1(n28456), .A2(n28019), .B(n905), .ZN(n29607) );
  NAND2_X1 U8590 ( .A1(n817), .A2(n20595), .ZN(n20598) );
  AOI22_X2 U8595 ( .A1(n1297), .A2(n15763), .B1(n22570), .B2(n18073), .ZN(
        n29608) );
  NOR2_X2 U8597 ( .A1(n17348), .A2(n27635), .ZN(n21696) );
  XOR2_X1 U8608 ( .A1(n4260), .A2(n8116), .Z(n21224) );
  NOR3_X1 U8620 ( .A1(n19322), .A2(n19274), .A3(n30894), .ZN(n6023) );
  INV_X1 U8622 ( .I(n10075), .ZN(n12419) );
  XOR2_X1 U8624 ( .A1(n10075), .A2(n29609), .Z(n22003) );
  INV_X1 U8629 ( .I(n25098), .ZN(n29609) );
  NAND2_X2 U8631 ( .A1(n6766), .A2(n6764), .ZN(n10075) );
  OR2_X2 U8643 ( .A1(n2019), .A2(n28245), .Z(n10264) );
  OAI22_X2 U8661 ( .A1(n21843), .A2(n338), .B1(n21841), .B2(n27937), .ZN(
        n14595) );
  NAND2_X1 U8674 ( .A1(n4259), .A2(n18767), .ZN(n18377) );
  INV_X2 U8683 ( .I(n29330), .ZN(n10376) );
  NAND2_X2 U8684 ( .A1(n4709), .A2(n4706), .ZN(n2600) );
  OAI21_X2 U8691 ( .A1(n19843), .A2(n7609), .B(n29615), .ZN(n15169) );
  XOR2_X1 U8720 ( .A1(n22078), .A2(n22059), .Z(n22284) );
  NAND2_X2 U8732 ( .A1(n9545), .A2(n27445), .ZN(n13473) );
  XOR2_X1 U8743 ( .A1(n29618), .A2(n19713), .Z(n9760) );
  XOR2_X1 U8744 ( .A1(n19711), .A2(n25998), .Z(n29618) );
  NOR2_X1 U8751 ( .A1(n27910), .A2(n386), .ZN(n15405) );
  OR2_X1 U8764 ( .A1(n9759), .A2(n5287), .Z(n5267) );
  NAND3_X1 U8772 ( .A1(n22670), .A2(n858), .A3(n994), .ZN(n29620) );
  NAND2_X1 U8779 ( .A1(n18089), .A2(n8100), .ZN(n8783) );
  INV_X2 U8792 ( .I(n16209), .ZN(n18976) );
  XOR2_X1 U8830 ( .A1(n29828), .A2(n20671), .Z(n29624) );
  XOR2_X1 U8877 ( .A1(n24116), .A2(n25990), .Z(n30774) );
  INV_X2 U8883 ( .I(n15633), .ZN(n725) );
  NAND2_X2 U8884 ( .A1(n15636), .A2(n28894), .ZN(n15633) );
  OR2_X1 U8898 ( .A1(n10899), .A2(n10900), .Z(n18118) );
  INV_X2 U8901 ( .I(n11172), .ZN(n29629) );
  BUF_X4 U8924 ( .I(n4646), .Z(n38) );
  INV_X2 U8930 ( .I(n29631), .ZN(n12974) );
  NAND2_X1 U8937 ( .A1(n3673), .A2(n4041), .ZN(n4040) );
  XOR2_X1 U8938 ( .A1(n14385), .A2(n24602), .Z(n8987) );
  NAND2_X2 U8939 ( .A1(n8989), .A2(n8988), .ZN(n24602) );
  NAND2_X2 U8940 ( .A1(n23046), .A2(n23045), .ZN(n23047) );
  XOR2_X1 U8949 ( .A1(n24755), .A2(n12754), .Z(n18001) );
  NAND2_X2 U8960 ( .A1(n17587), .A2(n8114), .ZN(n24755) );
  NAND2_X1 U8984 ( .A1(n25736), .A2(n10285), .ZN(n8555) );
  NOR2_X1 U8991 ( .A1(n31325), .A2(n27007), .ZN(n10972) );
  XOR2_X1 U9014 ( .A1(n13716), .A2(n29633), .Z(n20657) );
  XOR2_X1 U9019 ( .A1(n27643), .A2(n26647), .Z(n29633) );
  OAI22_X2 U9030 ( .A1(n834), .A2(n1214), .B1(n32590), .B2(n33155), .ZN(n1620)
         );
  BUF_X4 U9032 ( .I(n13646), .Z(n29769) );
  NOR2_X1 U9035 ( .A1(n22899), .A2(n31325), .ZN(n27410) );
  NOR2_X1 U9037 ( .A1(n15947), .A2(n15946), .ZN(n29706) );
  INV_X2 U9038 ( .I(n14238), .ZN(n18242) );
  NAND2_X2 U9042 ( .A1(n7049), .A2(n7050), .ZN(n31085) );
  XOR2_X1 U9050 ( .A1(n15083), .A2(n29636), .Z(n27766) );
  XOR2_X1 U9055 ( .A1(n3009), .A2(n24833), .Z(n29636) );
  NAND2_X1 U9063 ( .A1(n23984), .A2(n1233), .ZN(n31553) );
  XOR2_X1 U9086 ( .A1(n29638), .A2(n15427), .Z(n15425) );
  NOR2_X1 U9091 ( .A1(n29213), .A2(n14661), .ZN(n31442) );
  XOR2_X1 U9092 ( .A1(n22237), .A2(n1716), .Z(n85) );
  XOR2_X1 U9094 ( .A1(n22294), .A2(n18189), .Z(n22237) );
  XOR2_X1 U9100 ( .A1(n4400), .A2(n11219), .Z(n6720) );
  NAND2_X1 U9116 ( .A1(n24210), .A2(n29785), .ZN(n2944) );
  NAND2_X2 U9117 ( .A1(n7261), .A2(n23582), .ZN(n24210) );
  NAND2_X1 U9124 ( .A1(n3094), .A2(n3096), .ZN(n20189) );
  AND2_X2 U9125 ( .A1(n11333), .A2(n26551), .Z(n19845) );
  INV_X2 U9129 ( .I(n29642), .ZN(n596) );
  NAND2_X2 U9136 ( .A1(n31074), .A2(n8910), .ZN(n8909) );
  NOR2_X2 U9148 ( .A1(n21573), .A2(n33992), .ZN(n21627) );
  XOR2_X1 U9154 ( .A1(n12714), .A2(n29643), .Z(n16886) );
  XOR2_X1 U9160 ( .A1(n29042), .A2(n2616), .Z(n20794) );
  NAND2_X2 U9161 ( .A1(n30942), .A2(n2610), .ZN(n2616) );
  NOR2_X1 U9162 ( .A1(n28455), .A2(n11045), .ZN(n1522) );
  BUF_X2 U9165 ( .I(n19668), .Z(n29644) );
  AOI22_X2 U9166 ( .A1(n30854), .A2(n11912), .B1(n5480), .B2(n6842), .ZN(n9842) );
  XOR2_X1 U9175 ( .A1(n4884), .A2(n29645), .Z(n4881) );
  XOR2_X1 U9178 ( .A1(n4883), .A2(n28859), .Z(n29645) );
  XOR2_X1 U9179 ( .A1(n29646), .A2(n5207), .Z(n6039) );
  XOR2_X1 U9182 ( .A1(n14593), .A2(n5206), .Z(n29646) );
  XOR2_X1 U9185 ( .A1(n20920), .A2(n20892), .Z(n20972) );
  OAI22_X2 U9193 ( .A1(n9435), .A2(n6675), .B1(n17202), .B2(n22861), .ZN(
        n23519) );
  NAND2_X1 U9195 ( .A1(n30637), .A2(n28064), .ZN(n17878) );
  NAND2_X2 U9202 ( .A1(n20188), .A2(n20190), .ZN(n30637) );
  XOR2_X1 U9220 ( .A1(n9303), .A2(n4858), .Z(n20974) );
  INV_X2 U9232 ( .I(n29650), .ZN(n15467) );
  XOR2_X1 U9235 ( .A1(n27135), .A2(n1445), .Z(n29650) );
  NOR2_X2 U9239 ( .A1(n32800), .A2(n15371), .ZN(n21652) );
  XOR2_X1 U9241 ( .A1(n22269), .A2(n31913), .Z(n27106) );
  XOR2_X1 U9242 ( .A1(n21945), .A2(n26193), .Z(n22269) );
  XOR2_X1 U9243 ( .A1(n8571), .A2(n30943), .Z(n31857) );
  NOR2_X1 U9247 ( .A1(n20258), .A2(n29603), .ZN(n29651) );
  XOR2_X1 U9249 ( .A1(n6609), .A2(n29653), .Z(n30905) );
  XOR2_X1 U9255 ( .A1(n30540), .A2(n16479), .Z(n23552) );
  NAND2_X2 U9257 ( .A1(n28113), .A2(n4928), .ZN(n30540) );
  INV_X2 U9265 ( .I(n21846), .ZN(n29654) );
  NOR2_X1 U9267 ( .A1(n29118), .A2(n1180), .ZN(n2869) );
  XOR2_X1 U9281 ( .A1(n19664), .A2(n29657), .Z(n19901) );
  XOR2_X1 U9287 ( .A1(n19659), .A2(n19660), .Z(n29657) );
  XOR2_X1 U9295 ( .A1(n29660), .A2(n23264), .Z(n23265) );
  XOR2_X1 U9301 ( .A1(n29661), .A2(n19305), .Z(n19307) );
  AND2_X1 U9325 ( .A1(n11333), .A2(n6693), .Z(n15072) );
  NOR2_X1 U9332 ( .A1(n29663), .A2(n29662), .ZN(n26611) );
  NOR2_X1 U9333 ( .A1(n26198), .A2(n24956), .ZN(n29662) );
  INV_X2 U9352 ( .I(n29666), .ZN(n19418) );
  XNOR2_X1 U9354 ( .A1(n5487), .A2(n11591), .ZN(n29666) );
  INV_X2 U9355 ( .I(n10871), .ZN(n903) );
  INV_X2 U9359 ( .I(n8438), .ZN(n17590) );
  XOR2_X1 U9361 ( .A1(n10707), .A2(n27766), .Z(n8438) );
  OR2_X1 U9362 ( .A1(n20120), .A2(n16595), .Z(n6223) );
  INV_X2 U9364 ( .I(n29667), .ZN(n20278) );
  BUF_X4 U9375 ( .I(n20990), .Z(n31584) );
  XOR2_X1 U9377 ( .A1(n24747), .A2(n29670), .Z(n31849) );
  NAND2_X2 U9378 ( .A1(n3902), .A2(n15224), .ZN(n24747) );
  NOR2_X2 U9381 ( .A1(n4521), .A2(n4522), .ZN(n12414) );
  OAI22_X2 U9382 ( .A1(n3624), .A2(n1163), .B1(n29671), .B2(n13348), .ZN(n9352) );
  AOI22_X2 U9383 ( .A1(n12408), .A2(n822), .B1(n3626), .B2(n3790), .ZN(n29671)
         );
  NOR2_X2 U9392 ( .A1(n28862), .A2(n28863), .ZN(n14623) );
  XOR2_X1 U9397 ( .A1(n12330), .A2(n14518), .Z(n14517) );
  INV_X2 U9398 ( .I(n29673), .ZN(n12408) );
  XOR2_X1 U9402 ( .A1(n12411), .A2(n12409), .Z(n29673) );
  XOR2_X1 U9408 ( .A1(n3109), .A2(n29675), .Z(n29674) );
  NAND2_X2 U9415 ( .A1(n26291), .A2(n29225), .ZN(n31504) );
  NOR2_X2 U9420 ( .A1(n5966), .A2(n26615), .ZN(n6016) );
  AND2_X1 U9421 ( .A1(n12471), .A2(n23085), .Z(n13839) );
  NAND2_X2 U9426 ( .A1(n31139), .A2(n34018), .ZN(n5485) );
  NOR2_X2 U9428 ( .A1(n6794), .A2(n6793), .ZN(n6763) );
  INV_X4 U9448 ( .I(n29679), .ZN(n8178) );
  OAI22_X2 U9449 ( .A1(n155), .A2(n1933), .B1(n15681), .B2(n15683), .ZN(n29679) );
  XOR2_X1 U9451 ( .A1(n29680), .A2(n5421), .Z(n5441) );
  XOR2_X1 U9454 ( .A1(n22180), .A2(n2763), .Z(n29680) );
  NOR2_X2 U9456 ( .A1(n9510), .A2(n9509), .ZN(n9508) );
  XOR2_X1 U9462 ( .A1(n13606), .A2(n13457), .Z(n20806) );
  AOI22_X2 U9464 ( .A1(n12030), .A2(n8186), .B1(n11951), .B2(n1082), .ZN(
        n29681) );
  NAND2_X1 U9475 ( .A1(n29682), .A2(n23851), .ZN(n4106) );
  AOI21_X2 U9491 ( .A1(n12209), .A2(n29380), .B(n992), .ZN(n13894) );
  NAND2_X2 U9507 ( .A1(n30966), .A2(n4268), .ZN(n6169) );
  XOR2_X1 U9512 ( .A1(n1344), .A2(n20996), .Z(n20911) );
  AOI22_X2 U9518 ( .A1(n13548), .A2(n18892), .B1(n18792), .B2(n8376), .ZN(
        n5456) );
  XOR2_X1 U9534 ( .A1(n12258), .A2(n29687), .Z(n5500) );
  XOR2_X1 U9536 ( .A1(n30048), .A2(n5348), .Z(n12258) );
  INV_X2 U9537 ( .I(n29688), .ZN(n9390) );
  XOR2_X1 U9541 ( .A1(n7887), .A2(n29689), .Z(n30600) );
  XOR2_X1 U9542 ( .A1(n9629), .A2(n9292), .Z(n2363) );
  AOI22_X2 U9545 ( .A1(n1768), .A2(n19236), .B1(n1766), .B2(n1767), .ZN(n9292)
         );
  NAND2_X1 U9558 ( .A1(n21412), .A2(n11513), .ZN(n21113) );
  XOR2_X1 U9568 ( .A1(n29696), .A2(n29447), .Z(n575) );
  XOR2_X1 U9579 ( .A1(n19444), .A2(n26534), .Z(n29696) );
  NAND2_X2 U9606 ( .A1(n19928), .A2(n19929), .ZN(n16606) );
  INV_X2 U9624 ( .I(n4107), .ZN(n9218) );
  XOR2_X1 U9628 ( .A1(n13644), .A2(n17837), .Z(n4107) );
  NAND2_X2 U9637 ( .A1(n4456), .A2(n28364), .ZN(n23273) );
  XOR2_X1 U9653 ( .A1(n13347), .A2(n23333), .Z(n23440) );
  AOI22_X2 U9661 ( .A1(n22574), .A2(n9959), .B1(n16503), .B2(n22926), .ZN(
        n9647) );
  NAND2_X2 U9664 ( .A1(n29699), .A2(n26713), .ZN(n24328) );
  XOR2_X1 U9674 ( .A1(n6229), .A2(n14817), .Z(n29702) );
  OAI22_X2 U9677 ( .A1(n16013), .A2(n21488), .B1(n16736), .B2(n16012), .ZN(
        n22044) );
  XOR2_X1 U9686 ( .A1(n8810), .A2(n8811), .Z(n29704) );
  XOR2_X1 U9705 ( .A1(n23242), .A2(n29707), .Z(n450) );
  INV_X1 U9707 ( .I(n16598), .ZN(n29707) );
  XOR2_X1 U9734 ( .A1(n28552), .A2(n23264), .Z(n29709) );
  AND2_X1 U9740 ( .A1(n23840), .A2(n739), .Z(n23493) );
  XOR2_X1 U9742 ( .A1(n30057), .A2(n7874), .Z(n31248) );
  INV_X2 U9744 ( .I(n22251), .ZN(n6435) );
  NAND2_X2 U9751 ( .A1(n29711), .A2(n21399), .ZN(n21628) );
  XOR2_X1 U9758 ( .A1(n7796), .A2(n24632), .Z(n24754) );
  INV_X2 U9761 ( .I(n29712), .ZN(n11805) );
  XNOR2_X1 U9762 ( .A1(n7998), .A2(n11806), .ZN(n29712) );
  XOR2_X1 U9764 ( .A1(n33633), .A2(n16138), .Z(n29989) );
  NOR2_X2 U9772 ( .A1(n28915), .A2(n17960), .ZN(n29714) );
  OAI22_X2 U9779 ( .A1(n21343), .A2(n5141), .B1(n9073), .B2(n21341), .ZN(
        n29717) );
  OAI21_X2 U9782 ( .A1(n30681), .A2(n27574), .B(n15032), .ZN(n30410) );
  BUF_X2 U9792 ( .I(n28951), .Z(n29718) );
  XOR2_X1 U9803 ( .A1(n33492), .A2(n12454), .Z(n6687) );
  NOR2_X2 U9806 ( .A1(n31785), .A2(n15973), .ZN(n27922) );
  AND2_X1 U9807 ( .A1(n17963), .A2(n10327), .Z(n1521) );
  AND2_X1 U9813 ( .A1(n8857), .A2(n19960), .Z(n29841) );
  OAI22_X2 U9821 ( .A1(n9191), .A2(n17985), .B1(n30313), .B2(n18035), .ZN(
        n21264) );
  XOR2_X1 U9834 ( .A1(n29720), .A2(n12628), .Z(n10475) );
  OAI22_X2 U9842 ( .A1(n1008), .A2(n21708), .B1(n21709), .B2(n30440), .ZN(
        n29721) );
  NAND2_X2 U9852 ( .A1(n30688), .A2(n29722), .ZN(n9107) );
  NOR2_X1 U9857 ( .A1(n11916), .A2(n15467), .ZN(n29922) );
  XOR2_X1 U9867 ( .A1(n29723), .A2(n25071), .Z(Ciphertext[43]) );
  NOR2_X2 U9874 ( .A1(n29725), .A2(n29724), .ZN(n10949) );
  AND2_X1 U9876 ( .A1(n432), .A2(n5016), .Z(n5017) );
  NAND2_X2 U9878 ( .A1(n31136), .A2(n26431), .ZN(n432) );
  NAND2_X2 U9894 ( .A1(n29727), .A2(n12379), .ZN(n13346) );
  NOR2_X2 U9908 ( .A1(n12296), .A2(n12297), .ZN(n11454) );
  AOI21_X2 U9914 ( .A1(n6864), .A2(n1826), .B(n6263), .ZN(n29729) );
  NAND2_X2 U9915 ( .A1(n24152), .A2(n5317), .ZN(n27259) );
  NAND2_X1 U9925 ( .A1(n3204), .A2(n18359), .ZN(n29731) );
  XOR2_X1 U9926 ( .A1(n29732), .A2(n16507), .Z(Ciphertext[22]) );
  NAND2_X1 U9930 ( .A1(n16021), .A2(n26275), .ZN(n29732) );
  XOR2_X1 U9933 ( .A1(n29733), .A2(n4004), .Z(n4243) );
  XOR2_X1 U9934 ( .A1(n30774), .A2(n5425), .Z(n29733) );
  XOR2_X1 U9942 ( .A1(n1342), .A2(n20861), .Z(n6465) );
  NOR2_X2 U9978 ( .A1(n15991), .A2(n18839), .ZN(n19389) );
  NOR2_X2 U9986 ( .A1(n729), .A2(n19853), .ZN(n19854) );
  NAND3_X1 U9997 ( .A1(n16389), .A2(n16466), .A3(n16572), .ZN(n29738) );
  NAND2_X2 U10023 ( .A1(n2360), .A2(n30140), .ZN(n7256) );
  OR2_X1 U10031 ( .A1(n11814), .A2(n12037), .Z(n30227) );
  BUF_X4 U10043 ( .I(n28885), .Z(n30010) );
  NAND2_X1 U10045 ( .A1(n28736), .A2(n7554), .ZN(n6816) );
  XOR2_X1 U10087 ( .A1(n20717), .A2(n31526), .Z(n20785) );
  NAND2_X1 U10094 ( .A1(n15298), .A2(n26109), .ZN(n29741) );
  NAND3_X2 U10123 ( .A1(n2337), .A2(n8753), .A3(n396), .ZN(n31051) );
  NOR2_X2 U10131 ( .A1(n2795), .A2(n28183), .ZN(n31408) );
  NAND2_X2 U10151 ( .A1(n887), .A2(n24805), .ZN(n1646) );
  NAND2_X2 U10189 ( .A1(n29751), .A2(n16948), .ZN(n18576) );
  NAND2_X2 U10204 ( .A1(n29148), .A2(n31404), .ZN(n21945) );
  AOI21_X1 U10258 ( .A1(n1074), .A2(n27183), .B(n32867), .ZN(n15855) );
  NAND2_X2 U10266 ( .A1(n22974), .A2(n22973), .ZN(n7004) );
  NAND2_X1 U10273 ( .A1(n29755), .A2(n3931), .ZN(n8305) );
  NAND2_X1 U10274 ( .A1(n12804), .A2(n8813), .ZN(n29755) );
  NAND2_X2 U10275 ( .A1(n14176), .A2(n20466), .ZN(n21018) );
  INV_X2 U10280 ( .I(n16451), .ZN(n753) );
  OAI21_X1 U10309 ( .A1(n26753), .A2(n25773), .B(n25788), .ZN(n25777) );
  NAND2_X2 U10311 ( .A1(n14703), .A2(n11200), .ZN(n17566) );
  NAND2_X1 U10320 ( .A1(n21165), .A2(n4755), .ZN(n7063) );
  NOR2_X2 U10321 ( .A1(n3308), .A2(n3307), .ZN(n3350) );
  NAND2_X2 U10333 ( .A1(n29934), .A2(n29759), .ZN(n24094) );
  NAND3_X1 U10334 ( .A1(n15803), .A2(n23939), .A3(n12080), .ZN(n29759) );
  XOR2_X1 U10343 ( .A1(n19439), .A2(n19440), .Z(n9004) );
  XOR2_X1 U10365 ( .A1(n8283), .A2(n9760), .Z(n9759) );
  OAI21_X2 U10368 ( .A1(n8084), .A2(n7544), .B(n29761), .ZN(n7357) );
  NAND2_X2 U10371 ( .A1(n22890), .A2(n16501), .ZN(n29761) );
  XOR2_X1 U10374 ( .A1(n22157), .A2(n33437), .Z(n22213) );
  XOR2_X1 U10382 ( .A1(n24503), .A2(n29762), .Z(n16510) );
  NAND2_X2 U10396 ( .A1(n3556), .A2(n8769), .ZN(n30450) );
  XOR2_X1 U10397 ( .A1(n29765), .A2(n24833), .Z(Ciphertext[6]) );
  NAND4_X2 U10398 ( .A1(n24348), .A2(n24349), .A3(n24930), .A4(n24350), .ZN(
        n29765) );
  NAND2_X2 U10401 ( .A1(n14579), .A2(n26793), .ZN(n25796) );
  NOR2_X2 U10413 ( .A1(n31016), .A2(n29396), .ZN(n31015) );
  INV_X4 U10415 ( .I(n11904), .ZN(n15682) );
  AOI21_X2 U10416 ( .A1(n17566), .A2(n5041), .B(n28945), .ZN(n26874) );
  OAI21_X2 U10426 ( .A1(n21668), .A2(n11991), .B(n21674), .ZN(n5996) );
  OAI21_X2 U10438 ( .A1(n30512), .A2(n17963), .B(n17894), .ZN(n17475) );
  NAND2_X2 U10439 ( .A1(n29771), .A2(n33480), .ZN(n17894) );
  NOR2_X1 U10446 ( .A1(n16194), .A2(n31379), .ZN(n16195) );
  XOR2_X1 U10457 ( .A1(Plaintext[144]), .A2(Key[144]), .Z(n29776) );
  XOR2_X1 U10458 ( .A1(n6702), .A2(n29778), .Z(n6700) );
  XOR2_X1 U10459 ( .A1(n13644), .A2(n20801), .Z(n29778) );
  NOR3_X2 U10485 ( .A1(n2582), .A2(n4017), .A3(n1181), .ZN(n16353) );
  NOR2_X1 U10490 ( .A1(n30727), .A2(n29978), .ZN(n6786) );
  NAND2_X2 U10503 ( .A1(n21698), .A2(n21699), .ZN(n3704) );
  XOR2_X1 U10522 ( .A1(n24766), .A2(n29787), .Z(n13511) );
  XOR2_X1 U10523 ( .A1(n30290), .A2(n3294), .Z(n29787) );
  XOR2_X1 U10525 ( .A1(n24393), .A2(n12493), .Z(n24829) );
  NAND3_X2 U10529 ( .A1(n31208), .A2(n13576), .A3(n31209), .ZN(n29788) );
  XOR2_X1 U10531 ( .A1(n2489), .A2(n265), .Z(n5020) );
  OR2_X1 U10551 ( .A1(n12615), .A2(n23841), .Z(n31691) );
  OAI21_X2 U10552 ( .A1(n29791), .A2(n8990), .B(n2113), .ZN(n2112) );
  XOR2_X1 U10557 ( .A1(n23230), .A2(n16073), .Z(n23427) );
  NAND3_X2 U10559 ( .A1(n7412), .A2(n26705), .A3(n22717), .ZN(n23230) );
  XOR2_X1 U10568 ( .A1(n29536), .A2(n27185), .Z(n28868) );
  NAND2_X2 U10572 ( .A1(n1544), .A2(n1543), .ZN(n27185) );
  AOI21_X2 U10586 ( .A1(n18386), .A2(n3836), .B(n18385), .ZN(n5118) );
  NAND2_X2 U10598 ( .A1(n20624), .A2(n20622), .ZN(n29814) );
  XOR2_X1 U10599 ( .A1(n30997), .A2(n21958), .Z(n26340) );
  AND2_X1 U10612 ( .A1(n15394), .A2(n13969), .Z(n18172) );
  XOR2_X1 U10628 ( .A1(n29800), .A2(n23509), .Z(n28870) );
  XOR2_X1 U10630 ( .A1(n8916), .A2(n8915), .Z(n29800) );
  XOR2_X1 U10633 ( .A1(n2665), .A2(n2668), .Z(n25141) );
  OR2_X1 U10638 ( .A1(n28731), .A2(n27958), .Z(n28009) );
  INV_X2 U10642 ( .I(n29803), .ZN(n29270) );
  XOR2_X1 U10643 ( .A1(n6762), .A2(n6760), .Z(n29803) );
  NAND3_X2 U10652 ( .A1(n7580), .A2(n7579), .A3(n29804), .ZN(n20605) );
  OR2_X1 U10653 ( .A1(n16243), .A2(n20109), .Z(n29804) );
  NAND2_X1 U10664 ( .A1(n28263), .A2(n8553), .ZN(n26046) );
  XOR2_X1 U10666 ( .A1(n5462), .A2(n16642), .Z(n9231) );
  INV_X2 U10670 ( .I(n21356), .ZN(n5395) );
  NAND2_X1 U10672 ( .A1(n9106), .A2(n9151), .ZN(n28001) );
  XOR2_X1 U10673 ( .A1(n4465), .A2(n4464), .Z(n4224) );
  XOR2_X1 U10678 ( .A1(n6445), .A2(n29969), .Z(n29807) );
  NOR2_X2 U10679 ( .A1(n4279), .A2(n29808), .ZN(n19048) );
  XOR2_X1 U10681 ( .A1(n29809), .A2(n6185), .Z(n27352) );
  XOR2_X1 U10695 ( .A1(n20822), .A2(n20842), .Z(n21000) );
  XOR2_X1 U10704 ( .A1(n29813), .A2(n29812), .Z(n9929) );
  XOR2_X1 U10707 ( .A1(n14404), .A2(n19443), .Z(n29812) );
  XOR2_X1 U10709 ( .A1(n19538), .A2(n9928), .Z(n29813) );
  NAND2_X1 U10724 ( .A1(n17597), .A2(n17598), .ZN(n9836) );
  XOR2_X1 U10728 ( .A1(n4087), .A2(n18121), .Z(n22457) );
  AND2_X1 U10753 ( .A1(n10199), .A2(n3013), .Z(n30067) );
  NAND2_X2 U10754 ( .A1(n10970), .A2(n10971), .ZN(n23200) );
  XOR2_X1 U10763 ( .A1(n22021), .A2(n21952), .Z(n21984) );
  NOR2_X2 U10777 ( .A1(n23623), .A2(n23622), .ZN(n24816) );
  NAND2_X2 U10792 ( .A1(n29818), .A2(n29817), .ZN(n7363) );
  XOR2_X1 U10799 ( .A1(n29820), .A2(n960), .Z(Ciphertext[131]) );
  AOI22_X1 U10801 ( .A1(n10959), .A2(n691), .B1(n3639), .B2(n30285), .ZN(
        n29820) );
  AOI22_X1 U10804 ( .A1(n15429), .A2(n27142), .B1(n13809), .B2(n15888), .ZN(
        n29821) );
  NOR2_X2 U10813 ( .A1(n29070), .A2(n10641), .ZN(n12762) );
  OAI22_X2 U10823 ( .A1(n10321), .A2(n29444), .B1(n10322), .B2(n10323), .ZN(
        n10332) );
  NAND2_X1 U10836 ( .A1(n13561), .A2(n22648), .ZN(n8427) );
  XOR2_X1 U10849 ( .A1(n26842), .A2(n29825), .Z(n3536) );
  XOR2_X1 U10851 ( .A1(n9267), .A2(n28606), .Z(n29825) );
  OR2_X1 U10852 ( .A1(n30506), .A2(n28450), .Z(n14525) );
  OR2_X1 U10855 ( .A1(n21669), .A2(n21604), .Z(n29827) );
  XOR2_X1 U10859 ( .A1(n21881), .A2(n21880), .Z(n22565) );
  XOR2_X1 U10880 ( .A1(n22264), .A2(n13612), .Z(n22023) );
  NOR2_X2 U10881 ( .A1(n30965), .A2(n13613), .ZN(n22264) );
  NAND2_X2 U10884 ( .A1(n13355), .A2(n11295), .ZN(n15117) );
  INV_X2 U10891 ( .I(n29829), .ZN(n11983) );
  NOR2_X2 U10895 ( .A1(n27307), .A2(n13587), .ZN(n29829) );
  AND2_X1 U10902 ( .A1(n16249), .A2(n18510), .Z(n17623) );
  AND2_X1 U10908 ( .A1(n8758), .A2(n15318), .Z(n16406) );
  NOR2_X2 U10911 ( .A1(n25670), .A2(n27173), .ZN(n14780) );
  NOR2_X1 U10916 ( .A1(n9582), .A2(n9584), .ZN(n29830) );
  INV_X2 U10923 ( .I(n8189), .ZN(n29832) );
  NAND2_X2 U10926 ( .A1(n16606), .A2(n20565), .ZN(n13253) );
  NOR2_X1 U10930 ( .A1(n10409), .A2(n23768), .ZN(n29834) );
  AOI22_X2 U10935 ( .A1(n20234), .A2(n12263), .B1(n8942), .B2(n4647), .ZN(
        n29835) );
  NAND3_X2 U10940 ( .A1(n3546), .A2(n3545), .A3(n29836), .ZN(n7731) );
  NOR2_X2 U10943 ( .A1(n4164), .A2(n29837), .ZN(n16356) );
  OAI21_X2 U10945 ( .A1(n15682), .A2(n23804), .B(n12248), .ZN(n29837) );
  XOR2_X1 U10949 ( .A1(n23451), .A2(n23265), .Z(n23270) );
  OAI21_X2 U10952 ( .A1(n29841), .A2(n26774), .B(n16154), .ZN(n3293) );
  NAND2_X1 U10971 ( .A1(n29843), .A2(n26527), .ZN(n30054) );
  OAI21_X2 U10978 ( .A1(n7245), .A2(n7244), .B(n29844), .ZN(n7242) );
  NOR2_X2 U11000 ( .A1(n13525), .A2(n4916), .ZN(n4918) );
  NAND2_X2 U11002 ( .A1(n29847), .A2(n29846), .ZN(n5492) );
  NAND2_X2 U11005 ( .A1(n27294), .A2(n32106), .ZN(n29847) );
  NOR2_X1 U11019 ( .A1(n26635), .A2(n28701), .ZN(n29849) );
  XOR2_X1 U11022 ( .A1(n20693), .A2(n29851), .Z(n29850) );
  OR2_X1 U11043 ( .A1(n16781), .A2(n13905), .Z(n28670) );
  NOR2_X2 U11047 ( .A1(n4774), .A2(n12981), .ZN(n24133) );
  XOR2_X1 U11055 ( .A1(n31709), .A2(n9020), .Z(n27485) );
  XOR2_X1 U11059 ( .A1(n29855), .A2(n19440), .Z(n10780) );
  XOR2_X1 U11060 ( .A1(n34119), .A2(n11867), .Z(n19440) );
  XOR2_X1 U11062 ( .A1(n10783), .A2(n29856), .Z(n29855) );
  INV_X2 U11064 ( .I(n1372), .ZN(n29856) );
  NOR2_X1 U11071 ( .A1(n10680), .A2(n29451), .ZN(n8260) );
  NAND2_X1 U11108 ( .A1(n11898), .A2(n24611), .ZN(n24362) );
  INV_X2 U11117 ( .I(n5572), .ZN(n30048) );
  NAND3_X2 U11119 ( .A1(n5351), .A2(n5349), .A3(n5350), .ZN(n5572) );
  OAI22_X2 U11122 ( .A1(n10752), .A2(n8443), .B1(n6263), .B2(n6200), .ZN(
        n16050) );
  INV_X2 U11124 ( .I(n5187), .ZN(n10752) );
  XOR2_X1 U11131 ( .A1(n9573), .A2(n9571), .Z(n6458) );
  XOR2_X1 U11134 ( .A1(n14289), .A2(n1590), .Z(n29858) );
  XOR2_X1 U11160 ( .A1(n24543), .A2(n24542), .Z(n30029) );
  BUF_X2 U11168 ( .I(n28232), .Z(n29864) );
  NAND2_X1 U11169 ( .A1(n29865), .A2(n1101), .ZN(n30295) );
  XOR2_X1 U11170 ( .A1(n5278), .A2(n22877), .Z(n23924) );
  AND2_X1 U11172 ( .A1(n29296), .A2(n20569), .Z(n29867) );
  NAND2_X2 U11176 ( .A1(n7218), .A2(n2237), .ZN(n14280) );
  NAND2_X2 U11177 ( .A1(n7549), .A2(n31319), .ZN(n7218) );
  INV_X2 U11188 ( .I(n16603), .ZN(n23840) );
  NAND2_X1 U11189 ( .A1(n23887), .A2(n32611), .ZN(n23491) );
  BUF_X2 U11193 ( .I(n16332), .Z(n29868) );
  INV_X2 U11211 ( .I(n20992), .ZN(n29870) );
  XOR2_X1 U11222 ( .A1(n4861), .A2(n4859), .Z(n4862) );
  NAND2_X2 U11224 ( .A1(n7240), .A2(n7241), .ZN(n21958) );
  XOR2_X1 U11226 ( .A1(n4894), .A2(n29873), .Z(n4014) );
  XOR2_X1 U11227 ( .A1(n7530), .A2(n1366), .Z(n29873) );
  NOR2_X1 U11231 ( .A1(n12347), .A2(n14983), .ZN(n29875) );
  OAI21_X2 U11245 ( .A1(n5553), .A2(n16532), .B(n33196), .ZN(n29877) );
  NOR2_X2 U11255 ( .A1(n8337), .A2(n8164), .ZN(n29878) );
  XOR2_X1 U11274 ( .A1(n23256), .A2(n29880), .Z(n5278) );
  XOR2_X1 U11276 ( .A1(n5277), .A2(n23536), .Z(n29880) );
  OAI21_X2 U11280 ( .A1(n17289), .A2(n28638), .B(n32057), .ZN(n28951) );
  AND2_X1 U11281 ( .A1(n9170), .A2(n29868), .Z(n22391) );
  AND2_X1 U11296 ( .A1(n14083), .A2(n20120), .Z(n19965) );
  XNOR2_X1 U11302 ( .A1(n20723), .A2(n506), .ZN(n30265) );
  NAND2_X2 U11305 ( .A1(n29888), .A2(n3475), .ZN(n27886) );
  NAND2_X2 U11306 ( .A1(n22446), .A2(n18073), .ZN(n29888) );
  NOR2_X1 U11310 ( .A1(n18957), .A2(n29769), .ZN(n18114) );
  OAI21_X2 U11311 ( .A1(n13949), .A2(n30648), .B(n13945), .ZN(n13646) );
  NOR2_X2 U11341 ( .A1(n8270), .A2(n10955), .ZN(n23638) );
  XNOR2_X1 U11342 ( .A1(n10262), .A2(n19462), .ZN(n30137) );
  AOI21_X2 U11363 ( .A1(n20506), .A2(n17531), .B(n10057), .ZN(n20511) );
  AOI21_X1 U11364 ( .A1(n20392), .A2(n9252), .B(n1158), .ZN(n20393) );
  XOR2_X1 U11367 ( .A1(n29895), .A2(n9593), .Z(n9592) );
  XOR2_X1 U11374 ( .A1(n22322), .A2(n29896), .Z(n29895) );
  NAND2_X1 U11384 ( .A1(n15377), .A2(n15375), .ZN(n7884) );
  AOI22_X2 U11411 ( .A1(n7446), .A2(n33882), .B1(n7430), .B2(n12933), .ZN(
        n26202) );
  XOR2_X1 U11415 ( .A1(n16897), .A2(n8630), .Z(n9474) );
  NOR2_X2 U11418 ( .A1(n7144), .A2(n14864), .ZN(n21700) );
  INV_X2 U11419 ( .I(n27070), .ZN(n817) );
  OAI21_X2 U11420 ( .A1(n10440), .A2(n10394), .B(n19809), .ZN(n27070) );
  INV_X2 U11428 ( .I(n14845), .ZN(n26410) );
  NAND2_X2 U11436 ( .A1(n24094), .A2(n18077), .ZN(n5160) );
  AOI21_X2 U11447 ( .A1(n7238), .A2(n27842), .B(n29900), .ZN(n21390) );
  INV_X1 U11449 ( .I(n21220), .ZN(n29901) );
  NAND2_X2 U11454 ( .A1(n31021), .A2(n2770), .ZN(n3009) );
  BUF_X2 U11457 ( .I(n21248), .Z(n29903) );
  OAI21_X2 U11470 ( .A1(n13840), .A2(n13841), .B(n17608), .ZN(n29904) );
  XOR2_X1 U11488 ( .A1(n15862), .A2(n15860), .Z(n25394) );
  XOR2_X1 U11489 ( .A1(n22294), .A2(n28162), .Z(n22322) );
  XOR2_X1 U11503 ( .A1(n29907), .A2(n10877), .Z(n26971) );
  XOR2_X1 U11506 ( .A1(n20838), .A2(n27014), .Z(n29907) );
  AND2_X1 U11511 ( .A1(n7901), .A2(n10868), .Z(n29089) );
  NAND2_X2 U11519 ( .A1(n29909), .A2(n18524), .ZN(n19143) );
  OAI21_X2 U11521 ( .A1(n18521), .A2(n18522), .B(n18849), .ZN(n29909) );
  NAND2_X2 U11530 ( .A1(n31356), .A2(n18926), .ZN(n18928) );
  XOR2_X1 U11547 ( .A1(n4219), .A2(n11481), .Z(n22250) );
  XOR2_X1 U11553 ( .A1(n10923), .A2(n24524), .Z(n29912) );
  INV_X2 U11554 ( .I(n29913), .ZN(n19177) );
  NAND2_X2 U11556 ( .A1(n29769), .A2(n19120), .ZN(n29913) );
  INV_X4 U11562 ( .I(n29914), .ZN(n5781) );
  INV_X4 U11563 ( .I(n14248), .ZN(n31012) );
  INV_X2 U11581 ( .I(n26677), .ZN(n4337) );
  NAND2_X1 U11586 ( .A1(n30025), .A2(n14062), .ZN(n84) );
  XOR2_X1 U11595 ( .A1(n31005), .A2(n26125), .Z(n16939) );
  XOR2_X1 U11596 ( .A1(n12801), .A2(n29442), .Z(n30229) );
  XOR2_X1 U11597 ( .A1(n19473), .A2(n27781), .Z(n12801) );
  NAND2_X2 U11598 ( .A1(n29915), .A2(n8013), .ZN(n19749) );
  NAND2_X2 U11599 ( .A1(n28883), .A2(n30412), .ZN(n29915) );
  INV_X2 U11602 ( .I(n29916), .ZN(n28087) );
  INV_X2 U11611 ( .I(n29919), .ZN(n29278) );
  NAND2_X2 U11637 ( .A1(n9113), .A2(n29921), .ZN(n2180) );
  NAND2_X1 U11642 ( .A1(n9110), .A2(n9111), .ZN(n29921) );
  XOR2_X1 U11646 ( .A1(n24593), .A2(n24644), .Z(n9121) );
  AND2_X1 U11651 ( .A1(n4274), .A2(n28737), .Z(n9817) );
  INV_X4 U11661 ( .I(n28087), .ZN(n20100) );
  XOR2_X1 U11663 ( .A1(n30321), .A2(n23247), .Z(n23478) );
  INV_X2 U11668 ( .I(n7935), .ZN(n24156) );
  XOR2_X1 U11708 ( .A1(n24369), .A2(n29930), .Z(n24447) );
  XOR2_X1 U11709 ( .A1(n24687), .A2(n28918), .Z(n29930) );
  AOI22_X1 U11714 ( .A1(n12077), .A2(n1362), .B1(n14210), .B2(n10286), .ZN(
        n3946) );
  OAI21_X2 U11720 ( .A1(n29932), .A2(n29931), .B(n21811), .ZN(n16477) );
  NOR2_X2 U11721 ( .A1(n1132), .A2(n15772), .ZN(n29932) );
  NAND2_X1 U11722 ( .A1(n33474), .A2(n12358), .ZN(n17169) );
  NAND3_X2 U11723 ( .A1(n24011), .A2(n12143), .A3(n24012), .ZN(n15988) );
  NAND3_X1 U11732 ( .A1(n5901), .A2(n964), .A3(n314), .ZN(n24997) );
  XOR2_X1 U11756 ( .A1(n6731), .A2(n13951), .Z(n30093) );
  NOR2_X2 U11758 ( .A1(n5161), .A2(n5389), .ZN(n24622) );
  OAI21_X2 U11762 ( .A1(n33745), .A2(n179), .B(n7690), .ZN(n29933) );
  XOR2_X1 U11763 ( .A1(n23387), .A2(n23333), .Z(n23504) );
  OAI21_X2 U11765 ( .A1(n22888), .A2(n22889), .B(n1561), .ZN(n23333) );
  AND2_X1 U11767 ( .A1(n30763), .A2(n28471), .Z(n3443) );
  OAI21_X2 U11777 ( .A1(n29937), .A2(n5730), .B(n5758), .ZN(n14849) );
  BUF_X2 U11781 ( .I(n20519), .Z(n29938) );
  INV_X1 U11784 ( .I(n1357), .ZN(n30971) );
  NAND2_X1 U11786 ( .A1(n21664), .A2(n8323), .ZN(n3016) );
  AND2_X1 U11792 ( .A1(n13896), .A2(n27143), .Z(n29002) );
  NAND2_X1 U11826 ( .A1(n32081), .A2(n14676), .ZN(n22402) );
  XOR2_X1 U11835 ( .A1(n2073), .A2(n2075), .Z(n2072) );
  AOI21_X2 U11849 ( .A1(n14705), .A2(n14706), .B(n18743), .ZN(n18435) );
  AND2_X1 U11850 ( .A1(n3486), .A2(n20155), .Z(n3529) );
  XOR2_X1 U11851 ( .A1(n14132), .A2(n20813), .Z(n6081) );
  NOR2_X2 U11852 ( .A1(n9418), .A2(n10715), .ZN(n14132) );
  OAI22_X2 U11862 ( .A1(n890), .A2(n24325), .B1(n29141), .B2(n24327), .ZN(
        n23982) );
  NAND2_X1 U11865 ( .A1(n15907), .A2(n7460), .ZN(n30036) );
  NOR2_X2 U11869 ( .A1(n20951), .A2(n29946), .ZN(n21876) );
  OAI22_X2 U11871 ( .A1(n20947), .A2(n13194), .B1(n21313), .B2(n20949), .ZN(
        n29946) );
  OAI21_X2 U11883 ( .A1(n12276), .A2(n2741), .B(n12277), .ZN(n30628) );
  XOR2_X1 U11900 ( .A1(n10598), .A2(n29951), .Z(n26933) );
  OR3_X2 U11908 ( .A1(n27134), .A2(n24970), .A3(n3843), .Z(n699) );
  INV_X4 U11914 ( .I(n29952), .ZN(n6985) );
  XOR2_X1 U11925 ( .A1(n22246), .A2(n29953), .Z(n26214) );
  XOR2_X1 U11929 ( .A1(n21923), .A2(n29954), .Z(n29953) );
  INV_X1 U11936 ( .I(n25091), .ZN(n29954) );
  XOR2_X1 U11944 ( .A1(n13477), .A2(n2818), .Z(n29955) );
  NOR2_X2 U11951 ( .A1(n33675), .A2(n4208), .ZN(n22886) );
  XNOR2_X1 U11966 ( .A1(n14120), .A2(n19580), .ZN(n19406) );
  NAND2_X2 U11970 ( .A1(n6602), .A2(n6603), .ZN(n19580) );
  AND2_X1 U11973 ( .A1(n3147), .A2(n3077), .Z(n10938) );
  AND2_X1 U11978 ( .A1(n9285), .A2(n28203), .Z(n9286) );
  NAND2_X2 U11979 ( .A1(n7312), .A2(n10339), .ZN(n9285) );
  INV_X2 U11990 ( .I(n9313), .ZN(n2491) );
  NAND2_X2 U11991 ( .A1(n21125), .A2(n21678), .ZN(n9313) );
  INV_X2 U11999 ( .I(n29960), .ZN(n26114) );
  XOR2_X1 U12001 ( .A1(n13235), .A2(n13234), .Z(n29960) );
  AOI21_X2 U12005 ( .A1(n13109), .A2(n32459), .B(n33544), .ZN(n5389) );
  XOR2_X1 U12032 ( .A1(n12310), .A2(n29970), .Z(n29969) );
  NAND3_X2 U12033 ( .A1(n11991), .A2(n21673), .A3(n918), .ZN(n5995) );
  INV_X2 U12041 ( .I(n25859), .ZN(n10897) );
  NAND2_X2 U12047 ( .A1(n13051), .A2(n13053), .ZN(n25859) );
  XOR2_X1 U12051 ( .A1(n10535), .A2(n16690), .Z(n23122) );
  NAND2_X2 U12052 ( .A1(n1471), .A2(n4936), .ZN(n10535) );
  INV_X2 U12053 ( .I(n4378), .ZN(n9578) );
  AND2_X1 U12055 ( .A1(n19104), .A2(n18923), .Z(n27616) );
  XOR2_X1 U12056 ( .A1(n27352), .A2(n24470), .Z(n24471) );
  AOI22_X2 U12065 ( .A1(n8086), .A2(n8165), .B1(n13268), .B2(n24213), .ZN(
        n31086) );
  INV_X2 U12082 ( .I(n32747), .ZN(n29972) );
  NAND2_X2 U12099 ( .A1(n30088), .A2(n11919), .ZN(n14498) );
  OAI21_X2 U12108 ( .A1(n26067), .A2(n13210), .B(n29973), .ZN(n13001) );
  NAND2_X2 U12109 ( .A1(n13210), .A2(n12708), .ZN(n29973) );
  NAND2_X1 U12113 ( .A1(n4378), .A2(n9064), .ZN(n26333) );
  NAND2_X2 U12154 ( .A1(n349), .A2(n26971), .ZN(n21219) );
  AND2_X1 U12164 ( .A1(n1299), .A2(n16647), .Z(n15449) );
  NAND2_X2 U12176 ( .A1(n29975), .A2(n31612), .ZN(n21860) );
  NOR2_X1 U12187 ( .A1(n9133), .A2(n8632), .ZN(n29978) );
  XOR2_X1 U12216 ( .A1(n22249), .A2(n22160), .Z(n2349) );
  OAI22_X2 U12221 ( .A1(n2352), .A2(n21861), .B1(n2351), .B2(n3756), .ZN(
        n22160) );
  NAND2_X2 U12228 ( .A1(n6099), .A2(n1109), .ZN(n26937) );
  XOR2_X1 U12256 ( .A1(n13305), .A2(n471), .Z(n11507) );
  XOR2_X1 U12279 ( .A1(n22114), .A2(n22096), .Z(n22171) );
  NAND3_X2 U12288 ( .A1(n27569), .A2(n18147), .A3(n27764), .ZN(n4289) );
  NAND2_X1 U12292 ( .A1(n19035), .A2(n13796), .ZN(n26817) );
  NAND2_X2 U12296 ( .A1(n6170), .A2(n6172), .ZN(n13796) );
  XOR2_X1 U12299 ( .A1(n31373), .A2(n16128), .Z(n24528) );
  XOR2_X1 U12334 ( .A1(n29986), .A2(n19752), .Z(n3967) );
  INV_X2 U12336 ( .I(n29987), .ZN(n4677) );
  XOR2_X1 U12340 ( .A1(Plaintext[53]), .A2(Key[53]), .Z(n29987) );
  NAND2_X1 U12341 ( .A1(n31799), .A2(n26818), .ZN(n18322) );
  XOR2_X1 U12344 ( .A1(n34082), .A2(n19644), .Z(n29988) );
  XOR2_X1 U12357 ( .A1(n29989), .A2(n19669), .Z(n19671) );
  XOR2_X1 U12361 ( .A1(n27395), .A2(n19783), .Z(n19505) );
  OAI21_X2 U12365 ( .A1(n17242), .A2(n32618), .B(n17241), .ZN(n16452) );
  NAND2_X1 U12366 ( .A1(n30656), .A2(n10173), .ZN(n25604) );
  XOR2_X1 U12370 ( .A1(n5429), .A2(n24519), .Z(n678) );
  OR2_X1 U12391 ( .A1(n31360), .A2(n13483), .Z(n8805) );
  XNOR2_X1 U12393 ( .A1(n8785), .A2(n1410), .ZN(n31749) );
  AOI21_X1 U12403 ( .A1(n16648), .A2(n11820), .B(n26912), .ZN(n30568) );
  AOI22_X2 U12413 ( .A1(n19940), .A2(n13994), .B1(n19941), .B2(n16637), .ZN(
        n26278) );
  XOR2_X1 U12415 ( .A1(n17552), .A2(n11661), .Z(n11660) );
  XOR2_X1 U12431 ( .A1(n5324), .A2(n16852), .Z(n27192) );
  NAND2_X1 U12432 ( .A1(n20013), .A2(n31046), .ZN(n16261) );
  XOR2_X1 U12442 ( .A1(n2608), .A2(n2607), .Z(n20098) );
  OAI21_X2 U12443 ( .A1(n30004), .A2(n30003), .B(n1030), .ZN(n11617) );
  XOR2_X1 U12447 ( .A1(n19483), .A2(n19599), .Z(n19681) );
  OAI21_X2 U12452 ( .A1(n18391), .A2(n18390), .B(n18389), .ZN(n19101) );
  XOR2_X1 U12454 ( .A1(n26623), .A2(n30007), .Z(n7572) );
  NAND2_X2 U12458 ( .A1(n11336), .A2(n11489), .ZN(n26623) );
  NAND2_X2 U12463 ( .A1(n26543), .A2(n10850), .ZN(n10847) );
  XOR2_X1 U12469 ( .A1(n3030), .A2(n22274), .Z(n2477) );
  AND2_X1 U12478 ( .A1(n22364), .A2(n22588), .Z(n30507) );
  OAI21_X2 U12479 ( .A1(n26015), .A2(n25303), .B(n18059), .ZN(n11111) );
  XOR2_X1 U12480 ( .A1(n13743), .A2(n30011), .Z(n17886) );
  XOR2_X1 U12483 ( .A1(n13741), .A2(n13742), .Z(n30011) );
  AOI22_X1 U12484 ( .A1(n2130), .A2(n28849), .B1(n22981), .B2(n1280), .ZN(
        n17893) );
  XOR2_X1 U12485 ( .A1(n32623), .A2(n25881), .Z(n17753) );
  OR2_X1 U12489 ( .A1(n23777), .A2(n23778), .Z(n8720) );
  NAND2_X1 U12501 ( .A1(n16725), .A2(n1048), .ZN(n30012) );
  NOR2_X1 U12506 ( .A1(n5657), .A2(n26317), .ZN(n6232) );
  BUF_X2 U12509 ( .I(n8919), .Z(n30014) );
  INV_X2 U12512 ( .I(n5003), .ZN(n7394) );
  AND2_X1 U12515 ( .A1(n19422), .A2(n12704), .Z(n30015) );
  AOI22_X2 U12520 ( .A1(n21091), .A2(n21687), .B1(n29286), .B2(n26513), .ZN(
        n29148) );
  XOR2_X1 U12525 ( .A1(n31088), .A2(n29009), .Z(n31087) );
  BUF_X4 U12527 ( .I(n25700), .Z(n146) );
  XOR2_X1 U12538 ( .A1(n27976), .A2(n30016), .Z(n14456) );
  OR2_X1 U12551 ( .A1(n22332), .A2(n468), .Z(n13369) );
  XOR2_X1 U12556 ( .A1(n20792), .A2(n30018), .Z(n20449) );
  INV_X2 U12566 ( .I(n30020), .ZN(n10465) );
  XOR2_X1 U12568 ( .A1(n16324), .A2(n10466), .Z(n30020) );
  NAND2_X2 U12577 ( .A1(n31793), .A2(n30021), .ZN(n6595) );
  OAI22_X2 U12579 ( .A1(n30522), .A2(n30983), .B1(n765), .B2(n16783), .ZN(
        n30021) );
  OAI21_X2 U12583 ( .A1(n18618), .A2(n10080), .B(n10964), .ZN(n10977) );
  NOR2_X2 U12591 ( .A1(n9403), .A2(n20472), .ZN(n31532) );
  OAI22_X1 U12600 ( .A1(n25464), .A2(n25467), .B1(n25463), .B2(n25473), .ZN(
        n28302) );
  NAND2_X2 U12602 ( .A1(n19056), .A2(n6022), .ZN(n2075) );
  OAI21_X2 U12627 ( .A1(n26047), .A2(n28495), .B(n852), .ZN(n9244) );
  NAND2_X1 U12640 ( .A1(n25715), .A2(n25714), .ZN(n14352) );
  XOR2_X1 U12651 ( .A1(n23516), .A2(n16382), .Z(n16259) );
  INV_X2 U12654 ( .I(n30032), .ZN(n26049) );
  XOR2_X1 U12655 ( .A1(Plaintext[188]), .A2(Key[188]), .Z(n30032) );
  AND2_X1 U12656 ( .A1(n17298), .A2(n17514), .Z(n30222) );
  NAND2_X2 U12660 ( .A1(n12977), .A2(n12975), .ZN(n19049) );
  NAND3_X2 U12670 ( .A1(n30036), .A2(n30072), .A3(n9381), .ZN(n27105) );
  NAND2_X2 U12702 ( .A1(n26742), .A2(n12533), .ZN(n30039) );
  NAND2_X1 U12709 ( .A1(n20464), .A2(n30728), .ZN(n20466) );
  INV_X2 U12713 ( .I(n21860), .ZN(n5628) );
  INV_X2 U12719 ( .I(n30042), .ZN(n15623) );
  OAI22_X2 U12735 ( .A1(n27318), .A2(n8107), .B1(n8108), .B2(n18089), .ZN(
        n20188) );
  XOR2_X1 U12736 ( .A1(Plaintext[43]), .A2(Key[43]), .Z(n16585) );
  XNOR2_X1 U12744 ( .A1(n14819), .A2(n23419), .ZN(n30317) );
  OAI21_X2 U12753 ( .A1(n7429), .A2(n22342), .B(n26173), .ZN(n30044) );
  NAND2_X1 U12761 ( .A1(n20411), .A2(n29356), .ZN(n20047) );
  INV_X2 U12766 ( .I(n21049), .ZN(n30045) );
  OAI21_X2 U12774 ( .A1(n11444), .A2(n11280), .B(n11474), .ZN(n19312) );
  OAI21_X2 U12784 ( .A1(n3092), .A2(n3091), .B(n31226), .ZN(n6022) );
  NAND2_X1 U12785 ( .A1(n28913), .A2(n26594), .ZN(n30192) );
  NAND2_X1 U12792 ( .A1(n13905), .A2(n6662), .ZN(n28672) );
  XOR2_X1 U12793 ( .A1(n13817), .A2(n9373), .Z(n30049) );
  NAND2_X2 U12797 ( .A1(n12563), .A2(n13693), .ZN(n20328) );
  OR2_X1 U12799 ( .A1(n29629), .A2(n29334), .Z(n4968) );
  OAI21_X2 U12801 ( .A1(n11633), .A2(n12332), .B(n30054), .ZN(n17697) );
  NOR2_X1 U12805 ( .A1(n32055), .A2(n4378), .ZN(n4054) );
  NAND2_X2 U12809 ( .A1(n12542), .A2(n28155), .ZN(n22078) );
  INV_X2 U12815 ( .I(n24996), .ZN(n713) );
  INV_X1 U12819 ( .I(n19571), .ZN(n30058) );
  NAND3_X2 U12820 ( .A1(n10369), .A2(n20051), .A3(n11216), .ZN(n21047) );
  BUF_X2 U12831 ( .I(n23579), .Z(n30059) );
  OAI21_X2 U12834 ( .A1(n29375), .A2(n30060), .B(n8835), .ZN(n3166) );
  NAND2_X2 U12846 ( .A1(n30062), .A2(n7199), .ZN(n19661) );
  OAI21_X2 U12850 ( .A1(n16463), .A2(n13619), .B(n13618), .ZN(n23171) );
  XOR2_X1 U12851 ( .A1(n30063), .A2(n16691), .Z(Ciphertext[34]) );
  INV_X2 U12856 ( .I(n10303), .ZN(n22551) );
  NAND2_X2 U12867 ( .A1(n24187), .A2(n24188), .ZN(n15536) );
  OAI21_X2 U12871 ( .A1(n12326), .A2(n14529), .B(n798), .ZN(n24187) );
  XOR2_X1 U12880 ( .A1(n22269), .A2(n8061), .Z(n8060) );
  XOR2_X1 U12888 ( .A1(n19741), .A2(n19708), .Z(n17010) );
  BUF_X2 U12896 ( .I(n6407), .Z(n252) );
  NAND2_X2 U12909 ( .A1(n5627), .A2(n34008), .ZN(n23896) );
  XOR2_X1 U12944 ( .A1(n30074), .A2(n26436), .Z(n8373) );
  INV_X2 U12952 ( .I(n30076), .ZN(n15719) );
  XOR2_X1 U12958 ( .A1(n17570), .A2(n17572), .Z(n30076) );
  XOR2_X1 U12962 ( .A1(n23355), .A2(n23395), .Z(n11324) );
  XOR2_X1 U12971 ( .A1(n1044), .A2(n19780), .Z(n19495) );
  INV_X2 U12983 ( .I(n30078), .ZN(n11521) );
  XOR2_X1 U12984 ( .A1(n11522), .A2(n11524), .Z(n30078) );
  AOI21_X2 U12989 ( .A1(n14500), .A2(n32054), .B(n26768), .ZN(n17369) );
  NAND2_X2 U13012 ( .A1(n388), .A2(n387), .ZN(n25473) );
  NAND2_X2 U13014 ( .A1(n30080), .A2(n10329), .ZN(n4732) );
  XOR2_X1 U13015 ( .A1(n8762), .A2(n16497), .Z(n30596) );
  NAND2_X2 U13016 ( .A1(n7584), .A2(n30142), .ZN(n8762) );
  NAND2_X2 U13024 ( .A1(n21207), .A2(n30081), .ZN(n14691) );
  NAND2_X2 U13033 ( .A1(n30082), .A2(n9496), .ZN(n25723) );
  NAND3_X2 U13041 ( .A1(n27359), .A2(n25702), .A3(n27127), .ZN(n30082) );
  NAND2_X2 U13049 ( .A1(n10281), .A2(n24014), .ZN(n11883) );
  XOR2_X1 U13052 ( .A1(n13511), .A2(n13513), .Z(n13567) );
  NAND2_X2 U13055 ( .A1(n4734), .A2(n23065), .ZN(n10644) );
  OAI22_X2 U13067 ( .A1(n2152), .A2(n26918), .B1(n10472), .B2(n19152), .ZN(
        n19644) );
  XOR2_X1 U13070 ( .A1(n2330), .A2(n17213), .Z(n11434) );
  XOR2_X1 U13071 ( .A1(n2331), .A2(n1916), .Z(n2330) );
  XOR2_X1 U13075 ( .A1(n19493), .A2(n14223), .Z(n14222) );
  XOR2_X1 U13078 ( .A1(n19632), .A2(n33749), .Z(n19493) );
  XOR2_X1 U13083 ( .A1(n982), .A2(n5211), .Z(n23402) );
  OR2_X1 U13084 ( .A1(n23755), .A2(n6705), .Z(n15400) );
  XOR2_X1 U13088 ( .A1(n3932), .A2(n30188), .Z(n29213) );
  XOR2_X1 U13090 ( .A1(n30912), .A2(n3777), .Z(n5097) );
  AOI22_X2 U13096 ( .A1(n10627), .A2(n24237), .B1(n24131), .B2(n24130), .ZN(
        n30084) );
  OAI22_X2 U13100 ( .A1(n3866), .A2(n3867), .B1(n6568), .B2(n10096), .ZN(
        n25975) );
  NOR2_X1 U13120 ( .A1(n20630), .A2(n31471), .ZN(n20383) );
  OAI22_X2 U13121 ( .A1(n4230), .A2(n32618), .B1(n10695), .B2(n9139), .ZN(
        n31471) );
  NAND2_X2 U13125 ( .A1(n6580), .A2(n28459), .ZN(n5879) );
  INV_X4 U13135 ( .I(n16453), .ZN(n14233) );
  NOR2_X2 U13138 ( .A1(n32935), .A2(n29329), .ZN(n22840) );
  NAND2_X1 U13139 ( .A1(n30085), .A2(n11465), .ZN(n11464) );
  OAI21_X1 U13142 ( .A1(n5911), .A2(n4261), .B(n28812), .ZN(n30085) );
  INV_X2 U13144 ( .I(n30086), .ZN(n17316) );
  XNOR2_X1 U13145 ( .A1(Plaintext[86]), .A2(Key[86]), .ZN(n30086) );
  XOR2_X1 U13147 ( .A1(n13645), .A2(n28889), .Z(n30679) );
  AOI22_X2 U13152 ( .A1(n15716), .A2(n21496), .B1(n21601), .B2(n25975), .ZN(
        n21602) );
  XOR2_X1 U13159 ( .A1(n6462), .A2(n30087), .Z(n31660) );
  AOI22_X2 U13172 ( .A1(n5852), .A2(n4550), .B1(n14117), .B2(n18493), .ZN(
        n30088) );
  AOI21_X1 U13178 ( .A1(n14498), .A2(n18988), .B(n19089), .ZN(n18900) );
  XOR2_X1 U13185 ( .A1(n22195), .A2(n17244), .Z(n14301) );
  XOR2_X1 U13188 ( .A1(n22255), .A2(n22014), .Z(n22195) );
  NAND2_X2 U13191 ( .A1(n30090), .A2(n31814), .ZN(n3157) );
  INV_X2 U13201 ( .I(n29328), .ZN(n1280) );
  OAI22_X1 U13203 ( .A1(n12551), .A2(n12520), .B1(n3222), .B2(n24249), .ZN(
        n8204) );
  INV_X2 U13205 ( .I(n24250), .ZN(n3222) );
  NOR2_X1 U13217 ( .A1(n28183), .A2(n33848), .ZN(n16159) );
  XOR2_X1 U13221 ( .A1(n11251), .A2(n30093), .Z(n31128) );
  INV_X2 U13222 ( .I(n30094), .ZN(n15559) );
  XOR2_X1 U13223 ( .A1(n16178), .A2(n20691), .Z(n3010) );
  XOR2_X1 U13227 ( .A1(n20802), .A2(n20690), .Z(n16178) );
  NAND2_X2 U13229 ( .A1(n9460), .A2(n22774), .ZN(n22778) );
  OAI22_X2 U13232 ( .A1(n19078), .A2(n19283), .B1(n28721), .B2(n31254), .ZN(
        n28638) );
  AOI21_X2 U13245 ( .A1(n27023), .A2(n16327), .B(n27560), .ZN(n16796) );
  NOR3_X2 U13246 ( .A1(n3214), .A2(n30096), .A3(n24108), .ZN(n3504) );
  NAND2_X1 U13249 ( .A1(n4069), .A2(n29305), .ZN(n12568) );
  XOR2_X1 U13253 ( .A1(n20820), .A2(n20851), .Z(n20966) );
  XOR2_X1 U13255 ( .A1(n12610), .A2(n6974), .Z(n19343) );
  NOR2_X2 U13256 ( .A1(n30097), .A2(n2930), .ZN(n2929) );
  NOR2_X2 U13257 ( .A1(n13585), .A2(n20084), .ZN(n30097) );
  NAND2_X2 U13261 ( .A1(n12640), .A2(n12641), .ZN(n13872) );
  XOR2_X1 U13263 ( .A1(n22016), .A2(n10963), .Z(n30098) );
  XOR2_X1 U13265 ( .A1(n9468), .A2(n12800), .Z(n6688) );
  XOR2_X1 U13272 ( .A1(n12675), .A2(n25560), .Z(n6103) );
  OAI21_X2 U13273 ( .A1(n6105), .A2(n6106), .B(n6104), .ZN(n12675) );
  XOR2_X1 U13280 ( .A1(n10150), .A2(n27866), .Z(n10291) );
  XOR2_X1 U13292 ( .A1(n30137), .A2(n30102), .Z(n568) );
  XOR2_X1 U13294 ( .A1(n19476), .A2(n7741), .Z(n30102) );
  OAI21_X2 U13297 ( .A1(n29976), .A2(n16752), .B(n25143), .ZN(n25168) );
  NOR2_X2 U13304 ( .A1(n8760), .A2(n23721), .ZN(n23722) );
  XOR2_X1 U13308 ( .A1(n28730), .A2(n2825), .Z(n2824) );
  XOR2_X1 U13313 ( .A1(n30107), .A2(n5166), .Z(n12584) );
  NAND2_X1 U13320 ( .A1(n7515), .A2(n25214), .ZN(n15339) );
  XOR2_X1 U13322 ( .A1(n19579), .A2(n30109), .Z(n7939) );
  XOR2_X1 U13326 ( .A1(n19737), .A2(n1367), .Z(n30109) );
  XOR2_X1 U13331 ( .A1(n24399), .A2(n29348), .Z(n13358) );
  NAND2_X2 U13334 ( .A1(n30110), .A2(n24319), .ZN(n14789) );
  XOR2_X1 U13349 ( .A1(n22066), .A2(n21986), .Z(n61) );
  XOR2_X1 U13353 ( .A1(n22157), .A2(n22225), .Z(n22066) );
  XOR2_X1 U13357 ( .A1(n11660), .A2(n30111), .Z(n12467) );
  XOR2_X1 U13360 ( .A1(n19444), .A2(n11663), .Z(n30111) );
  NAND2_X1 U13368 ( .A1(n14016), .A2(n5820), .ZN(n30888) );
  XOR2_X1 U13372 ( .A1(n13436), .A2(n30644), .Z(n637) );
  NOR3_X2 U13378 ( .A1(n7857), .A2(n26667), .A3(n26739), .ZN(n30578) );
  NAND3_X2 U13386 ( .A1(n7488), .A2(n14024), .A3(n30112), .ZN(n14600) );
  OAI21_X1 U13391 ( .A1(n18843), .A2(n5700), .B(n4927), .ZN(n4507) );
  NAND2_X2 U13392 ( .A1(n30115), .A2(n30114), .ZN(n13579) );
  INV_X2 U13393 ( .I(n24110), .ZN(n889) );
  BUF_X2 U13405 ( .I(n469), .Z(n30116) );
  AND2_X1 U13427 ( .A1(n7320), .A2(n414), .Z(n2705) );
  AND2_X1 U13429 ( .A1(n25480), .A2(n25482), .Z(n30117) );
  NAND2_X1 U13435 ( .A1(n3181), .A2(n29043), .ZN(n27934) );
  NAND2_X2 U13472 ( .A1(n30122), .A2(n26568), .ZN(n4208) );
  NOR2_X2 U13497 ( .A1(n25229), .A2(n18059), .ZN(n11409) );
  AOI21_X1 U13500 ( .A1(n9832), .A2(n9833), .B(n8087), .ZN(n30236) );
  OAI22_X2 U13501 ( .A1(n18784), .A2(n34141), .B1(n6777), .B2(n18785), .ZN(
        n13963) );
  NAND2_X2 U13503 ( .A1(n8395), .A2(n13254), .ZN(n18784) );
  INV_X2 U13523 ( .I(n30125), .ZN(n11516) );
  XOR2_X1 U13528 ( .A1(n30127), .A2(n8920), .Z(n30126) );
  BUF_X2 U13537 ( .I(n21816), .Z(n30129) );
  NAND2_X2 U13551 ( .A1(n8378), .A2(n21430), .ZN(n11299) );
  OR2_X1 U13555 ( .A1(n11516), .A2(n29139), .Z(n23859) );
  XOR2_X1 U13568 ( .A1(n6904), .A2(n30135), .Z(n6886) );
  XOR2_X1 U13570 ( .A1(n22138), .A2(n30906), .Z(n30135) );
  XOR2_X1 U13572 ( .A1(n30136), .A2(n14885), .Z(Ciphertext[109]) );
  AOI22_X1 U13573 ( .A1(n25492), .A2(n25464), .B1(n25460), .B2(n25459), .ZN(
        n30136) );
  NAND2_X2 U13586 ( .A1(n13001), .A2(n13002), .ZN(n14337) );
  INV_X2 U13591 ( .I(n25557), .ZN(n15134) );
  XOR2_X1 U13599 ( .A1(n21003), .A2(n21038), .Z(n6895) );
  NAND2_X2 U13600 ( .A1(n12365), .A2(n12364), .ZN(n21038) );
  OR2_X1 U13603 ( .A1(n4054), .A2(n9580), .Z(n8199) );
  NAND3_X2 U13614 ( .A1(n24166), .A2(n31416), .A3(n24165), .ZN(n28830) );
  AOI22_X2 U13615 ( .A1(n25657), .A2(n25664), .B1(n7083), .B2(n25666), .ZN(
        n25668) );
  INV_X2 U13616 ( .I(n20344), .ZN(n30139) );
  XNOR2_X1 U13622 ( .A1(n24638), .A2(n25208), .ZN(n30607) );
  XOR2_X1 U13628 ( .A1(n28762), .A2(n17898), .Z(n22004) );
  NAND2_X1 U13630 ( .A1(n6841), .A2(n6840), .ZN(n30140) );
  NOR2_X2 U13635 ( .A1(n28361), .A2(n18994), .ZN(n19058) );
  NAND2_X2 U13636 ( .A1(n31856), .A2(n94), .ZN(n18994) );
  XOR2_X1 U13649 ( .A1(n24540), .A2(n9681), .Z(n2210) );
  AOI21_X2 U13653 ( .A1(n782), .A2(n20535), .B(n31250), .ZN(n26082) );
  NAND2_X2 U13672 ( .A1(n31244), .A2(n10825), .ZN(n3550) );
  INV_X2 U13674 ( .I(n30143), .ZN(n636) );
  XOR2_X1 U13676 ( .A1(n1589), .A2(n1588), .Z(n30143) );
  NAND2_X2 U13677 ( .A1(n29307), .A2(n24171), .ZN(n24191) );
  NOR2_X2 U13687 ( .A1(n29307), .A2(n24171), .ZN(n24273) );
  NAND2_X2 U13706 ( .A1(n4683), .A2(n320), .ZN(n6338) );
  NOR2_X2 U13711 ( .A1(n30148), .A2(n8354), .ZN(n8797) );
  XOR2_X1 U13714 ( .A1(n30149), .A2(n9116), .Z(n19788) );
  XOR2_X1 U13715 ( .A1(n19785), .A2(n19786), .Z(n30149) );
  OAI21_X2 U13719 ( .A1(n16096), .A2(n29402), .B(n751), .ZN(n30151) );
  XNOR2_X1 U13728 ( .A1(n32894), .A2(n25541), .ZN(n30722) );
  XOR2_X1 U13736 ( .A1(n9683), .A2(n5462), .Z(n27957) );
  NAND2_X2 U13742 ( .A1(n27159), .A2(n17310), .ZN(n26459) );
  NAND2_X2 U13751 ( .A1(n22845), .A2(n14882), .ZN(n23287) );
  OAI22_X2 U13759 ( .A1(n14232), .A2(n27577), .B1(n14133), .B2(n13720), .ZN(
        n23956) );
  INV_X2 U13762 ( .I(n25657), .ZN(n26322) );
  XOR2_X1 U13771 ( .A1(n27952), .A2(n12954), .Z(n23905) );
  NAND2_X2 U13777 ( .A1(n795), .A2(n29307), .ZN(n23991) );
  NAND2_X1 U13779 ( .A1(n11960), .A2(n33813), .ZN(n17562) );
  XOR2_X1 U13780 ( .A1(n23389), .A2(n23444), .Z(n23296) );
  XOR2_X1 U13795 ( .A1(n8154), .A2(n30559), .Z(n627) );
  XOR2_X1 U13799 ( .A1(n14499), .A2(n29345), .Z(n671) );
  XOR2_X1 U13811 ( .A1(n27882), .A2(n27881), .Z(n28343) );
  NAND2_X1 U13821 ( .A1(n30458), .A2(n30157), .ZN(n31065) );
  AOI22_X1 U13822 ( .A1(n17845), .A2(n25606), .B1(n25612), .B2(n32856), .ZN(
        n30157) );
  XOR2_X1 U13836 ( .A1(n20794), .A2(n20706), .Z(n20708) );
  XOR2_X1 U13842 ( .A1(n2672), .A2(n30159), .Z(n87) );
  XOR2_X1 U13846 ( .A1(n2671), .A2(n19732), .Z(n30159) );
  NAND2_X2 U13847 ( .A1(n32866), .A2(n2234), .ZN(n2654) );
  NAND3_X2 U13855 ( .A1(n24115), .A2(n3213), .A3(n3212), .ZN(n24116) );
  NOR2_X2 U13860 ( .A1(n22724), .A2(n22723), .ZN(n23103) );
  NAND2_X2 U13864 ( .A1(n26324), .A2(n26178), .ZN(n22724) );
  OR2_X1 U13865 ( .A1(n7941), .A2(n5492), .Z(n5112) );
  XOR2_X1 U13890 ( .A1(n19539), .A2(n19384), .Z(n19721) );
  NOR2_X2 U13893 ( .A1(n18457), .A2(n18458), .ZN(n19539) );
  NAND2_X2 U13894 ( .A1(n2729), .A2(n30169), .ZN(n13175) );
  OR2_X1 U13896 ( .A1(n5889), .A2(n19108), .Z(n12034) );
  NAND2_X2 U13904 ( .A1(n5632), .A2(n9219), .ZN(n24295) );
  XOR2_X1 U13937 ( .A1(n2356), .A2(n21009), .Z(n7016) );
  XOR2_X1 U13938 ( .A1(n30173), .A2(n31869), .Z(n686) );
  BUF_X4 U13940 ( .I(n17361), .Z(n3506) );
  BUF_X2 U13944 ( .I(n18879), .Z(n16588) );
  AOI21_X2 U13945 ( .A1(n15827), .A2(n26726), .B(n26725), .ZN(n27472) );
  NAND2_X2 U13946 ( .A1(n30174), .A2(n1763), .ZN(n9629) );
  XOR2_X1 U13949 ( .A1(n19376), .A2(n19377), .Z(n16324) );
  NAND2_X2 U13971 ( .A1(n30175), .A2(n18320), .ZN(n8379) );
  XOR2_X1 U13974 ( .A1(n30177), .A2(n30176), .Z(n21266) );
  XOR2_X1 U13976 ( .A1(n20889), .A2(n20850), .Z(n30176) );
  XOR2_X1 U13982 ( .A1(n20664), .A2(n20663), .Z(n30177) );
  NAND2_X1 U13983 ( .A1(n17543), .A2(n1101), .ZN(n30198) );
  AOI21_X2 U13985 ( .A1(n15286), .A2(n8558), .B(n20136), .ZN(n20139) );
  NOR2_X2 U14014 ( .A1(n17698), .A2(n30180), .ZN(n16519) );
  NOR3_X1 U14015 ( .A1(n4248), .A2(n9518), .A3(n21311), .ZN(n30180) );
  NAND2_X2 U14024 ( .A1(n16435), .A2(n18481), .ZN(n18604) );
  NAND2_X1 U14030 ( .A1(n13669), .A2(n13668), .ZN(n26713) );
  BUF_X2 U14045 ( .I(n3935), .Z(n30183) );
  XOR2_X1 U14058 ( .A1(n32255), .A2(n10075), .Z(n1937) );
  XOR2_X1 U14060 ( .A1(n1441), .A2(n29386), .Z(n31184) );
  NAND2_X2 U14061 ( .A1(n9954), .A2(n23031), .ZN(n30442) );
  NAND3_X2 U14065 ( .A1(n11700), .A2(n4082), .A3(n21137), .ZN(n21496) );
  XOR2_X1 U14069 ( .A1(n20552), .A2(n20752), .Z(n10789) );
  INV_X2 U14093 ( .I(n30187), .ZN(n31915) );
  NOR3_X2 U14094 ( .A1(n28037), .A2(n32644), .A3(n924), .ZN(n26411) );
  OAI21_X2 U14098 ( .A1(n951), .A2(n17557), .B(n12989), .ZN(n26203) );
  INV_X2 U14104 ( .I(n26203), .ZN(n13752) );
  NAND2_X2 U14105 ( .A1(n12567), .A2(n12565), .ZN(n30193) );
  XOR2_X1 U14113 ( .A1(n19432), .A2(n19435), .Z(n30188) );
  XOR2_X1 U14121 ( .A1(n23501), .A2(n30189), .Z(n5158) );
  XOR2_X1 U14122 ( .A1(n11193), .A2(n5157), .Z(n30189) );
  NAND2_X1 U14124 ( .A1(n17439), .A2(n1329), .ZN(n2833) );
  NOR2_X2 U14129 ( .A1(n11621), .A2(n13308), .ZN(n23946) );
  INV_X2 U14130 ( .I(n13764), .ZN(n16853) );
  XOR2_X1 U14133 ( .A1(n23505), .A2(n14492), .Z(n30190) );
  INV_X2 U14177 ( .I(n1787), .ZN(n2356) );
  NAND2_X2 U14179 ( .A1(n15662), .A2(n30195), .ZN(n20736) );
  OAI22_X2 U14184 ( .A1(n32068), .A2(n20451), .B1(n20450), .B2(n5471), .ZN(
        n30195) );
  XOR2_X1 U14196 ( .A1(n20737), .A2(n20738), .Z(n20739) );
  XOR2_X1 U14206 ( .A1(n20964), .A2(n500), .Z(n8701) );
  XOR2_X1 U14207 ( .A1(n31950), .A2(n2789), .Z(n20964) );
  OAI22_X2 U14222 ( .A1(n5653), .A2(n19121), .B1(n1051), .B2(n19148), .ZN(
        n31438) );
  OR2_X1 U14225 ( .A1(n25665), .A2(n25664), .Z(n25651) );
  AOI21_X2 U14236 ( .A1(n25292), .A2(n5468), .B(n7081), .ZN(n11069) );
  NAND2_X2 U14237 ( .A1(n30198), .A2(n23927), .ZN(n15227) );
  XOR2_X1 U14241 ( .A1(n19386), .A2(n1363), .Z(n19168) );
  XOR2_X1 U14245 ( .A1(n30199), .A2(n24991), .Z(Ciphertext[25]) );
  NAND2_X2 U14249 ( .A1(n6768), .A2(n6767), .ZN(n7879) );
  XOR2_X1 U14271 ( .A1(n30203), .A2(n16010), .Z(n27201) );
  XOR2_X1 U14273 ( .A1(n7211), .A2(n12715), .Z(n30203) );
  NOR2_X2 U14274 ( .A1(n2158), .A2(n2156), .ZN(n24805) );
  XOR2_X1 U14280 ( .A1(n24743), .A2(n7838), .Z(n7984) );
  NAND2_X2 U14284 ( .A1(n26120), .A2(n27184), .ZN(n24073) );
  NAND2_X1 U14287 ( .A1(n15528), .A2(n24511), .ZN(n30204) );
  OAI22_X2 U14289 ( .A1(n17906), .A2(n14664), .B1(n28365), .B2(n16097), .ZN(
        n10763) );
  OR2_X1 U14294 ( .A1(n24315), .A2(n13232), .Z(n16152) );
  NAND2_X2 U14304 ( .A1(n4730), .A2(n30207), .ZN(n9153) );
  INV_X2 U14326 ( .I(n32886), .ZN(n25620) );
  XOR2_X1 U14328 ( .A1(n17498), .A2(n6397), .Z(n17499) );
  BUF_X2 U14340 ( .I(n23587), .Z(n23588) );
  NOR2_X1 U14345 ( .A1(n12049), .A2(n25617), .ZN(n30497) );
  INV_X2 U14349 ( .I(n32887), .ZN(n789) );
  INV_X4 U14363 ( .I(n20414), .ZN(n1150) );
  OAI21_X2 U14365 ( .A1(n32746), .A2(n14761), .B(n873), .ZN(n11510) );
  XOR2_X1 U14371 ( .A1(n23218), .A2(n15742), .Z(n13498) );
  AOI22_X2 U14373 ( .A1(n10108), .A2(n26251), .B1(n10107), .B2(n850), .ZN(
        n23218) );
  AOI21_X2 U14379 ( .A1(n7361), .A2(n29141), .B(n890), .ZN(n9824) );
  OAI21_X2 U14380 ( .A1(n23035), .A2(n23034), .B(n13063), .ZN(n12446) );
  XOR2_X1 U14382 ( .A1(n30214), .A2(n7908), .Z(n29230) );
  BUF_X2 U14403 ( .I(n10469), .Z(n30318) );
  NAND2_X2 U14406 ( .A1(n18279), .A2(n18278), .ZN(n31451) );
  XOR2_X1 U14409 ( .A1(n30216), .A2(n671), .Z(n9932) );
  XOR2_X1 U14411 ( .A1(n24450), .A2(n16738), .Z(n30216) );
  NOR2_X2 U14415 ( .A1(n31459), .A2(n31333), .ZN(n30879) );
  XOR2_X1 U14417 ( .A1(n20896), .A2(n30218), .Z(n4756) );
  XOR2_X1 U14419 ( .A1(n15275), .A2(n4758), .Z(n30218) );
  XOR2_X1 U14420 ( .A1(n30220), .A2(n31405), .Z(n25762) );
  NAND3_X1 U14425 ( .A1(n932), .A2(n28011), .A3(n7242), .ZN(n17298) );
  NAND2_X2 U14429 ( .A1(n8854), .A2(n25594), .ZN(n25615) );
  XOR2_X1 U14433 ( .A1(n23171), .A2(n16672), .Z(n6091) );
  NOR2_X2 U14438 ( .A1(n8079), .A2(n21793), .ZN(n30223) );
  NOR2_X2 U14441 ( .A1(n932), .A2(n7242), .ZN(n10351) );
  NAND2_X2 U14444 ( .A1(n9408), .A2(n9407), .ZN(n30943) );
  XOR2_X1 U14445 ( .A1(n225), .A2(n30224), .Z(n17050) );
  XOR2_X1 U14446 ( .A1(n4792), .A2(n4467), .Z(n30224) );
  NAND3_X1 U14447 ( .A1(n14562), .A2(n15160), .A3(n11915), .ZN(n14561) );
  BUF_X2 U14448 ( .I(n33566), .Z(n16459) );
  NAND2_X2 U14464 ( .A1(n12849), .A2(n14455), .ZN(n19744) );
  OAI21_X2 U14467 ( .A1(n28385), .A2(n10093), .B(n30225), .ZN(n21463) );
  OAI21_X2 U14469 ( .A1(n24052), .A2(n30595), .B(n9973), .ZN(n5968) );
  INV_X2 U14478 ( .I(n3519), .ZN(n23532) );
  NAND2_X2 U14479 ( .A1(n32253), .A2(n8379), .ZN(n19215) );
  XOR2_X1 U14480 ( .A1(n10130), .A2(n8609), .Z(n412) );
  XOR2_X1 U14481 ( .A1(n30380), .A2(n23536), .Z(n10130) );
  INV_X2 U14484 ( .I(n17941), .ZN(n12105) );
  BUF_X2 U14490 ( .I(n24335), .Z(n30230) );
  XOR2_X1 U14504 ( .A1(n26256), .A2(n30815), .Z(n31467) );
  INV_X2 U14513 ( .I(n18994), .ZN(n14893) );
  NAND2_X2 U14515 ( .A1(n29330), .A2(n32887), .ZN(n6915) );
  INV_X2 U14517 ( .I(n15955), .ZN(n15956) );
  AOI21_X1 U14519 ( .A1(n13528), .A2(n25555), .B(n30232), .ZN(n13527) );
  OAI22_X1 U14522 ( .A1(n28759), .A2(n6391), .B1(n25555), .B2(n12864), .ZN(
        n30232) );
  NOR2_X2 U14526 ( .A1(n20087), .A2(n20086), .ZN(n9115) );
  NOR2_X2 U14528 ( .A1(n7182), .A2(n27954), .ZN(n30233) );
  OR2_X1 U14533 ( .A1(n24910), .A2(n24909), .Z(n10754) );
  XOR2_X1 U14536 ( .A1(n30235), .A2(n18019), .Z(Ciphertext[178]) );
  NAND3_X1 U14541 ( .A1(n27217), .A2(n18021), .A3(n18020), .ZN(n30235) );
  INV_X1 U14552 ( .I(n30236), .ZN(n2197) );
  XOR2_X1 U14554 ( .A1(n17745), .A2(n16816), .Z(n5601) );
  XOR2_X1 U14562 ( .A1(n30237), .A2(n20966), .Z(n17999) );
  XOR2_X1 U14564 ( .A1(n13681), .A2(n33219), .Z(n30237) );
  INV_X2 U14567 ( .I(n25855), .ZN(n25858) );
  NAND2_X2 U14569 ( .A1(n12697), .A2(n17627), .ZN(n30293) );
  NAND2_X2 U14595 ( .A1(n11899), .A2(n25756), .ZN(n5292) );
  XOR2_X1 U14596 ( .A1(n23166), .A2(n23199), .Z(n3905) );
  XOR2_X1 U14601 ( .A1(n23266), .A2(n11891), .Z(n23199) );
  NAND2_X2 U14635 ( .A1(n2045), .A2(n10358), .ZN(n30248) );
  INV_X1 U14636 ( .I(n31560), .ZN(n23601) );
  XOR2_X1 U14637 ( .A1(n17128), .A2(n5244), .Z(n8361) );
  XOR2_X1 U14641 ( .A1(n29137), .A2(n4285), .Z(n5244) );
  INV_X1 U14652 ( .I(n2861), .ZN(n31629) );
  NAND2_X2 U14659 ( .A1(n30779), .A2(n28754), .ZN(n30389) );
  NOR2_X2 U14660 ( .A1(n29224), .A2(n25678), .ZN(n27173) );
  NOR2_X2 U14661 ( .A1(n24438), .A2(n24437), .ZN(n29224) );
  XOR2_X1 U14665 ( .A1(n27868), .A2(n30250), .Z(n28624) );
  XOR2_X1 U14676 ( .A1(n19658), .A2(n27138), .Z(n19659) );
  NAND2_X1 U14691 ( .A1(n22455), .A2(n7965), .ZN(n30833) );
  NAND2_X2 U14699 ( .A1(n20429), .A2(n31533), .ZN(n20594) );
  XOR2_X1 U14700 ( .A1(n24762), .A2(n24626), .Z(n8893) );
  INV_X2 U14701 ( .I(n8834), .ZN(n30252) );
  AOI22_X2 U14714 ( .A1(n6660), .A2(n33992), .B1(n16600), .B2(n21628), .ZN(
        n21776) );
  INV_X2 U14715 ( .I(n21626), .ZN(n16600) );
  NOR2_X2 U14722 ( .A1(n31084), .A2(n31083), .ZN(n27914) );
  AND2_X1 U14737 ( .A1(n2317), .A2(n20376), .Z(n2316) );
  NAND2_X2 U14745 ( .A1(n9378), .A2(n8866), .ZN(n2575) );
  XOR2_X1 U14749 ( .A1(n30257), .A2(n5726), .Z(n5725) );
  XOR2_X1 U14755 ( .A1(n20693), .A2(n20776), .Z(n12609) );
  NAND2_X2 U14764 ( .A1(n20004), .A2(n20003), .ZN(n20693) );
  NAND2_X2 U14765 ( .A1(n24728), .A2(n30259), .ZN(n14915) );
  NOR2_X1 U14775 ( .A1(n146), .A2(n25763), .ZN(n24715) );
  BUF_X4 U14779 ( .I(n20483), .Z(n21306) );
  NAND2_X2 U14787 ( .A1(n30262), .A2(n7027), .ZN(n7197) );
  NAND2_X1 U14788 ( .A1(n12174), .A2(n12173), .ZN(n30262) );
  NOR2_X1 U14798 ( .A1(n25607), .A2(n10504), .ZN(n10501) );
  NAND2_X2 U14810 ( .A1(n24716), .A2(n24717), .ZN(n25818) );
  INV_X1 U14815 ( .I(n8243), .ZN(n28308) );
  XNOR2_X1 U14816 ( .A1(n2305), .A2(n30849), .ZN(n8243) );
  XOR2_X1 U14830 ( .A1(n17859), .A2(n12538), .Z(n1538) );
  OR2_X1 U14836 ( .A1(n23003), .A2(n23000), .Z(n31225) );
  NAND2_X2 U14840 ( .A1(n30342), .A2(n7815), .ZN(n5863) );
  NAND2_X2 U14848 ( .A1(n6369), .A2(n13043), .ZN(n13638) );
  XOR2_X1 U14859 ( .A1(n15776), .A2(n29441), .Z(n30387) );
  XOR2_X1 U14861 ( .A1(n17026), .A2(n30265), .Z(n30713) );
  NAND2_X2 U14871 ( .A1(n1882), .A2(n5944), .ZN(n30506) );
  OAI21_X2 U14876 ( .A1(n6661), .A2(n28671), .B(n4026), .ZN(n4025) );
  NAND2_X2 U14878 ( .A1(n27426), .A2(n13943), .ZN(n12616) );
  NAND2_X2 U14902 ( .A1(n951), .A2(n5473), .ZN(n31710) );
  NAND2_X2 U14903 ( .A1(n13764), .A2(n12864), .ZN(n17403) );
  OAI22_X2 U14914 ( .A1(n18118), .A2(n9127), .B1(n4993), .B2(n16113), .ZN(
        n9017) );
  INV_X2 U14930 ( .I(n19289), .ZN(n745) );
  OAI21_X1 U14935 ( .A1(n7397), .A2(n7836), .B(n20628), .ZN(n7396) );
  INV_X1 U14966 ( .I(n22598), .ZN(n22595) );
  AOI22_X1 U14969 ( .A1(n1521), .A2(n836), .B1(n1522), .B2(n25901), .ZN(n26793) );
  AOI21_X1 U14972 ( .A1(n24724), .A2(n29771), .B(n836), .ZN(n8299) );
  OR2_X1 U14977 ( .A1(n22336), .A2(n22486), .Z(n22416) );
  NAND2_X1 U14991 ( .A1(n24104), .A2(n18077), .ZN(n30459) );
  NAND3_X1 U14993 ( .A1(n15770), .A2(n17717), .A3(n28136), .ZN(n24585) );
  OAI22_X1 U15015 ( .A1(n18828), .A2(n16782), .B1(n17231), .B2(n16915), .ZN(
        n4279) );
  NAND3_X1 U15016 ( .A1(n17053), .A2(n21767), .A3(n21520), .ZN(n1648) );
  NOR2_X1 U15023 ( .A1(n9127), .A2(n4993), .ZN(n30269) );
  NOR2_X1 U15024 ( .A1(n757), .A2(n23940), .ZN(n13677) );
  INV_X1 U15032 ( .I(n24479), .ZN(n31762) );
  NAND2_X1 U15041 ( .A1(n24735), .A2(n9126), .ZN(n13944) );
  BUF_X4 U15042 ( .I(n16315), .Z(n13597) );
  INV_X1 U15047 ( .I(n19261), .ZN(n28544) );
  NAND2_X1 U15049 ( .A1(n21537), .A2(n8196), .ZN(n22308) );
  NAND2_X1 U15052 ( .A1(n5741), .A2(n29307), .ZN(n30270) );
  NAND3_X1 U15053 ( .A1(n24130), .A2(n32515), .A3(n974), .ZN(n8005) );
  OAI21_X1 U15054 ( .A1(n1858), .A2(n1861), .B(n25227), .ZN(n26380) );
  XOR2_X1 U15055 ( .A1(n18388), .A2(Key[111]), .Z(n30271) );
  AND2_X1 U15056 ( .A1(n4651), .A2(n4650), .Z(n30272) );
  INV_X2 U15058 ( .I(Plaintext[111]), .ZN(n18388) );
  INV_X1 U15064 ( .I(n1227), .ZN(n24648) );
  XNOR2_X1 U15068 ( .A1(n16448), .A2(n13864), .ZN(n30273) );
  INV_X2 U15069 ( .I(n31772), .ZN(n31918) );
  INV_X2 U15084 ( .I(n21455), .ZN(n780) );
  NAND2_X1 U15102 ( .A1(n115), .A2(n34084), .ZN(n22286) );
  CLKBUF_X12 U15112 ( .I(n23720), .Z(n16620) );
  AND3_X1 U15121 ( .A1(n17963), .A2(n11045), .A3(n25903), .Z(n10792) );
  INV_X1 U15125 ( .I(n18655), .ZN(n6118) );
  AND3_X2 U15128 ( .A1(n25342), .A2(n25341), .A3(n25340), .Z(n30276) );
  OAI21_X1 U15130 ( .A1(n25712), .A2(n25711), .B(n27208), .ZN(n31403) );
  NAND2_X1 U15134 ( .A1(n355), .A2(n6882), .ZN(n3597) );
  AOI22_X1 U15145 ( .A1(n11469), .A2(n965), .B1(n24960), .B2(n24948), .ZN(
        n24950) );
  NAND2_X1 U15147 ( .A1(n31564), .A2(n22871), .ZN(n30638) );
  NAND2_X1 U15155 ( .A1(n6338), .A2(n6337), .ZN(n21315) );
  NAND2_X1 U15160 ( .A1(n28037), .A2(n924), .ZN(n2468) );
  NOR2_X1 U15163 ( .A1(n924), .A2(n9678), .ZN(n1553) );
  NOR2_X1 U15164 ( .A1(n5883), .A2(n924), .ZN(n26369) );
  NOR3_X1 U15171 ( .A1(n21568), .A2(n30389), .A3(n21569), .ZN(n21351) );
  OAI21_X1 U15173 ( .A1(n14983), .A2(n21569), .B(n30389), .ZN(n3580) );
  NAND2_X1 U15189 ( .A1(n837), .A2(n967), .ZN(n13464) );
  NOR2_X1 U15195 ( .A1(n29269), .A2(n23681), .ZN(n8535) );
  NAND2_X1 U15202 ( .A1(n22314), .A2(n22549), .ZN(n22315) );
  XOR2_X1 U15213 ( .A1(n9868), .A2(n30278), .Z(n30277) );
  XNOR2_X1 U15214 ( .A1(n24774), .A2(n1948), .ZN(n30278) );
  NOR2_X1 U15220 ( .A1(n9127), .A2(n4993), .ZN(n28223) );
  INV_X2 U15222 ( .I(n25707), .ZN(n25708) );
  NAND2_X1 U15225 ( .A1(n27864), .A2(n27863), .ZN(n24020) );
  INV_X1 U15241 ( .I(n24133), .ZN(n27864) );
  AND2_X1 U15243 ( .A1(n24052), .A2(n29157), .Z(n31424) );
  INV_X2 U15244 ( .I(n17133), .ZN(n23872) );
  AND3_X2 U15245 ( .A1(n23695), .A2(n18182), .A3(n17133), .Z(n31396) );
  INV_X2 U15248 ( .I(n22824), .ZN(n723) );
  NAND2_X1 U15254 ( .A1(n24913), .A2(n27248), .ZN(n8278) );
  NOR2_X1 U15266 ( .A1(n14686), .A2(n15852), .ZN(n5689) );
  INV_X2 U15282 ( .I(n14686), .ZN(n15039) );
  OAI21_X1 U15283 ( .A1(n25760), .A2(n33976), .B(n25712), .ZN(n24438) );
  NAND3_X1 U15287 ( .A1(n8902), .A2(n749), .A3(n1204), .ZN(n1946) );
  NAND2_X2 U15297 ( .A1(n2997), .A2(n30855), .ZN(n30279) );
  NOR2_X2 U15298 ( .A1(n2999), .A2(n2998), .ZN(n2997) );
  NAND2_X1 U15312 ( .A1(n28691), .A2(n32176), .ZN(n11436) );
  INV_X2 U15316 ( .I(n21300), .ZN(n6082) );
  OAI21_X1 U15317 ( .A1(n20791), .A2(n20790), .B(n6082), .ZN(n3973) );
  NAND2_X1 U15320 ( .A1(n1808), .A2(n7581), .ZN(n24132) );
  NAND2_X1 U15331 ( .A1(n10135), .A2(n1332), .ZN(n30342) );
  NAND2_X1 U15332 ( .A1(n25343), .A2(n25344), .ZN(n14244) );
  CLKBUF_X4 U15348 ( .I(n25855), .Z(n14199) );
  NOR2_X1 U15349 ( .A1(n14681), .A2(n21704), .ZN(n21595) );
  INV_X2 U15353 ( .I(n14681), .ZN(n21705) );
  NOR2_X1 U15361 ( .A1(n21816), .A2(n1137), .ZN(n6626) );
  NAND2_X1 U15362 ( .A1(n21816), .A2(n31958), .ZN(n21818) );
  NAND2_X1 U15364 ( .A1(n254), .A2(n3019), .ZN(n24881) );
  NAND2_X1 U15372 ( .A1(n9953), .A2(n10354), .ZN(n22406) );
  INV_X1 U15373 ( .I(n10354), .ZN(n1000) );
  NAND2_X1 U15380 ( .A1(n25604), .A2(n27057), .ZN(n28775) );
  NAND2_X1 U15384 ( .A1(n16633), .A2(n16239), .ZN(n15442) );
  INV_X2 U15386 ( .I(n17721), .ZN(n23867) );
  INV_X1 U15390 ( .I(n23025), .ZN(n23653) );
  INV_X1 U15418 ( .I(n11931), .ZN(n831) );
  NAND2_X1 U15448 ( .A1(n22377), .A2(n17936), .ZN(n28225) );
  NOR2_X1 U15454 ( .A1(n11931), .A2(n10174), .ZN(n25606) );
  AOI21_X1 U15462 ( .A1(n10497), .A2(n25713), .B(n10393), .ZN(n11511) );
  NAND3_X2 U15470 ( .A1(n12399), .A2(n9736), .A3(n26069), .ZN(n29131) );
  NOR2_X1 U15473 ( .A1(n12541), .A2(n2958), .ZN(n10419) );
  NAND2_X1 U15474 ( .A1(n20525), .A2(n2958), .ZN(n2957) );
  CLKBUF_X4 U15494 ( .I(n5988), .Z(n5926) );
  AOI21_X1 U15498 ( .A1(n26887), .A2(n22808), .B(n26886), .ZN(n26885) );
  NAND2_X1 U15505 ( .A1(n34089), .A2(n13989), .ZN(n21181) );
  INV_X1 U15508 ( .I(n13989), .ZN(n17467) );
  INV_X2 U15517 ( .I(n8168), .ZN(n221) );
  NAND2_X1 U15518 ( .A1(n9342), .A2(n24031), .ZN(n24142) );
  NAND2_X1 U15522 ( .A1(n26479), .A2(n8079), .ZN(n6619) );
  OAI21_X1 U15527 ( .A1(n21479), .A2(n21711), .B(n21496), .ZN(n21480) );
  AOI21_X1 U15531 ( .A1(n28623), .A2(n16985), .B(n12374), .ZN(n16984) );
  NOR2_X1 U15537 ( .A1(n16984), .A2(n16983), .ZN(n16982) );
  NAND2_X1 U15538 ( .A1(n11943), .A2(n651), .ZN(n9772) );
  INV_X1 U15549 ( .I(n23916), .ZN(n23920) );
  NAND2_X1 U15550 ( .A1(n13326), .A2(n24985), .ZN(n14269) );
  NAND3_X1 U15555 ( .A1(n907), .A2(n10206), .A3(n856), .ZN(n13892) );
  INV_X1 U15556 ( .I(n907), .ZN(n10907) );
  INV_X1 U15558 ( .I(n14865), .ZN(n714) );
  NAND2_X2 U15569 ( .A1(n2000), .A2(n2001), .ZN(n30288) );
  INV_X1 U15572 ( .I(n2795), .ZN(n11587) );
  INV_X1 U15581 ( .I(n3718), .ZN(n24211) );
  NAND2_X1 U15582 ( .A1(n17426), .A2(n3718), .ZN(n7060) );
  OAI21_X1 U15585 ( .A1(n11132), .A2(n25339), .B(n10569), .ZN(n25338) );
  OR2_X2 U15586 ( .A1(n10569), .A2(n14788), .Z(n3430) );
  NOR2_X1 U15594 ( .A1(n16066), .A2(n4151), .ZN(n17069) );
  INV_X2 U15595 ( .I(n16066), .ZN(n24285) );
  NAND2_X1 U15597 ( .A1(n21805), .A2(n17077), .ZN(n10689) );
  NAND2_X1 U15601 ( .A1(n19220), .A2(n30995), .ZN(n18475) );
  NOR2_X1 U15602 ( .A1(n19220), .A2(n30995), .ZN(n31757) );
  AND2_X1 U15603 ( .A1(n4025), .A2(n27341), .Z(n30289) );
  AOI21_X1 U15610 ( .A1(n12485), .A2(n10822), .B(n25066), .ZN(n31206) );
  NAND2_X1 U15612 ( .A1(n13622), .A2(n30584), .ZN(n22745) );
  OAI21_X1 U15618 ( .A1(n5864), .A2(n5865), .B(n16809), .ZN(n30961) );
  NOR2_X2 U15620 ( .A1(n16815), .A2(n26966), .ZN(n30290) );
  NOR2_X1 U15624 ( .A1(n11298), .A2(n4184), .ZN(n18088) );
  OAI21_X1 U15625 ( .A1(n32652), .A2(n2092), .B(n25120), .ZN(n16611) );
  NAND2_X1 U15631 ( .A1(n25121), .A2(n2092), .ZN(n14867) );
  NAND2_X1 U15644 ( .A1(n25412), .A2(n25405), .ZN(n25299) );
  NAND3_X1 U15646 ( .A1(n32602), .A2(n10955), .A3(n843), .ZN(n9225) );
  INV_X2 U15647 ( .I(n10955), .ZN(n17694) );
  BUF_X2 U15648 ( .I(n23639), .Z(n14078) );
  NAND2_X1 U15651 ( .A1(n23735), .A2(n23765), .ZN(n30296) );
  NAND3_X1 U15652 ( .A1(n24213), .A2(n24210), .A3(n24209), .ZN(n23987) );
  NAND2_X1 U15656 ( .A1(n22622), .A2(n22497), .ZN(n22628) );
  NOR2_X1 U15681 ( .A1(n8576), .A2(n20029), .ZN(n30474) );
  OAI22_X1 U15686 ( .A1(n14793), .A2(n14747), .B1(n20155), .B2(n3486), .ZN(
        n5347) );
  NAND2_X1 U15693 ( .A1(n16812), .A2(n27808), .ZN(n6671) );
  OR2_X1 U15698 ( .A1(n25429), .A2(n17948), .Z(n25415) );
  INV_X1 U15703 ( .I(n27189), .ZN(n25745) );
  CLKBUF_X12 U15708 ( .I(Key[185]), .Z(n25493) );
  NAND2_X2 U15724 ( .A1(n11439), .A2(n11440), .ZN(n30301) );
  XNOR2_X1 U15738 ( .A1(n23371), .A2(n23530), .ZN(n23249) );
  OAI21_X2 U15743 ( .A1(n14247), .A2(n14245), .B(n14243), .ZN(n30302) );
  CLKBUF_X4 U15746 ( .I(n14577), .Z(n1647) );
  OAI21_X2 U15757 ( .A1(n18959), .A2(n4622), .B(n4619), .ZN(n30305) );
  NAND3_X1 U15775 ( .A1(n21433), .A2(n4683), .A3(n5049), .ZN(n8603) );
  NAND2_X1 U15786 ( .A1(n11438), .A2(n29157), .ZN(n11236) );
  NAND2_X1 U15805 ( .A1(n8057), .A2(n28451), .ZN(n20301) );
  INV_X1 U15806 ( .I(n20301), .ZN(n6559) );
  OAI22_X1 U15820 ( .A1(n24909), .A2(n10099), .B1(n24911), .B2(n24910), .ZN(
        n24916) );
  NAND2_X1 U15822 ( .A1(n30816), .A2(n4097), .ZN(n31202) );
  NAND2_X1 U15852 ( .A1(n21308), .A2(n16180), .ZN(n21309) );
  NOR3_X1 U15853 ( .A1(n21307), .A2(n21443), .A3(n21306), .ZN(n21230) );
  NAND2_X1 U15857 ( .A1(n19290), .A2(n27726), .ZN(n3204) );
  NAND2_X1 U15865 ( .A1(n4580), .A2(n16486), .ZN(n22905) );
  NAND2_X1 U15871 ( .A1(n9522), .A2(n24148), .ZN(n2153) );
  NOR2_X1 U15872 ( .A1(n24881), .A2(n30279), .ZN(n27062) );
  OAI21_X1 U15881 ( .A1(n5631), .A2(n9219), .B(n4286), .ZN(n10103) );
  INV_X1 U15884 ( .I(n19654), .ZN(n30766) );
  AOI22_X1 U15894 ( .A1(n7813), .A2(n7811), .B1(n5863), .B2(n21870), .ZN(
        n10493) );
  AOI22_X2 U15907 ( .A1(n31284), .A2(n34098), .B1(n21495), .B2(n1014), .ZN(
        n30309) );
  AOI22_X1 U15908 ( .A1(n31284), .A2(n34098), .B1(n21495), .B2(n1014), .ZN(
        n22080) );
  NAND2_X1 U15919 ( .A1(n10847), .A2(n29628), .ZN(n11616) );
  NOR2_X1 U15926 ( .A1(n14133), .A2(n12287), .ZN(n30991) );
  NAND2_X1 U15938 ( .A1(n21504), .A2(n21749), .ZN(n11585) );
  INV_X1 U15947 ( .I(n30033), .ZN(n21690) );
  INV_X2 U15949 ( .I(n16528), .ZN(n25405) );
  NOR2_X1 U15956 ( .A1(n10112), .A2(n29866), .ZN(n4522) );
  XOR2_X1 U15957 ( .A1(n4228), .A2(n7477), .Z(n30311) );
  NAND2_X1 U15958 ( .A1(n25277), .A2(n25276), .ZN(n25271) );
  NOR2_X1 U15976 ( .A1(n25780), .A2(n12611), .ZN(n25774) );
  XNOR2_X1 U15989 ( .A1(n18095), .A2(n16820), .ZN(n30313) );
  NAND3_X1 U15994 ( .A1(n6111), .A2(n13624), .A3(n30285), .ZN(n10035) );
  NOR2_X1 U15997 ( .A1(n7004), .A2(n13191), .ZN(n2712) );
  CLKBUF_X4 U15999 ( .I(n11722), .Z(n11370) );
  OAI21_X1 U16013 ( .A1(n17726), .A2(n8045), .B(n30252), .ZN(n9382) );
  NOR2_X1 U16020 ( .A1(n7083), .A2(n25653), .ZN(n25645) );
  NAND2_X1 U16021 ( .A1(n7083), .A2(n25659), .ZN(n25644) );
  AOI21_X1 U16029 ( .A1(n7083), .A2(n25653), .B(n25657), .ZN(n11211) );
  AND3_X1 U16045 ( .A1(n25403), .A2(n30308), .A3(n25295), .Z(n11259) );
  INV_X1 U16047 ( .I(n3405), .ZN(n30316) );
  INV_X1 U16052 ( .I(n10469), .ZN(n14940) );
  INV_X2 U16055 ( .I(n25334), .ZN(n25390) );
  OR2_X1 U16058 ( .A1(n17133), .A2(n8694), .Z(n23640) );
  OR2_X1 U16085 ( .A1(n29658), .A2(n15519), .Z(n13466) );
  NAND2_X1 U16086 ( .A1(n26322), .A2(n7083), .ZN(n6497) );
  INV_X1 U16087 ( .I(n9517), .ZN(n19515) );
  OAI22_X1 U16090 ( .A1(n8950), .A2(n7373), .B1(n7370), .B2(n7369), .ZN(n6526)
         );
  INV_X1 U16097 ( .I(n22063), .ZN(n1128) );
  NOR2_X1 U16103 ( .A1(n9041), .A2(n9042), .ZN(n30322) );
  INV_X2 U16122 ( .I(n23833), .ZN(n17726) );
  NAND2_X1 U16131 ( .A1(n25317), .A2(n31407), .ZN(n25315) );
  INV_X2 U16138 ( .I(n8606), .ZN(n19357) );
  NAND2_X1 U16151 ( .A1(n7312), .A2(n10339), .ZN(n30326) );
  NOR2_X1 U16152 ( .A1(n13279), .A2(n18581), .ZN(n8627) );
  NAND2_X1 U16153 ( .A1(n490), .A2(n18581), .ZN(n18583) );
  NAND2_X1 U16156 ( .A1(n18581), .A2(n31821), .ZN(n31820) );
  INV_X1 U16158 ( .I(n14770), .ZN(n24346) );
  NAND2_X1 U16170 ( .A1(n6075), .A2(n4755), .ZN(n30666) );
  INV_X2 U16171 ( .I(n4755), .ZN(n30784) );
  NOR2_X1 U16180 ( .A1(n30473), .A2(n24025), .ZN(n30328) );
  OAI21_X1 U16182 ( .A1(n16406), .A2(n1573), .B(n32760), .ZN(n25033) );
  NAND2_X2 U16184 ( .A1(n2394), .A2(n2393), .ZN(n30329) );
  INV_X1 U16206 ( .I(n25666), .ZN(n25660) );
  NOR2_X2 U16215 ( .A1(n22820), .A2(n22819), .ZN(n23120) );
  NOR2_X1 U16228 ( .A1(n7273), .A2(n7371), .ZN(n16833) );
  AOI22_X1 U16230 ( .A1(n7339), .A2(n7371), .B1(n14737), .B2(n16973), .ZN(
        n30740) );
  OAI21_X1 U16231 ( .A1(n7371), .A2(n32059), .B(n3489), .ZN(n7370) );
  INV_X2 U16232 ( .I(n28839), .ZN(n899) );
  AND2_X2 U16240 ( .A1(n23035), .A2(n28839), .Z(n17740) );
  NAND2_X1 U16241 ( .A1(n26261), .A2(n3469), .ZN(n30332) );
  NAND3_X1 U16253 ( .A1(n27785), .A2(n20575), .A3(n31968), .ZN(n8143) );
  AOI22_X1 U16259 ( .A1(n22509), .A2(n15601), .B1(n987), .B2(n22508), .ZN(
        n6503) );
  NOR2_X1 U16262 ( .A1(n987), .A2(n22955), .ZN(n6300) );
  AOI21_X1 U16267 ( .A1(n13532), .A2(n967), .B(n9858), .ZN(n9857) );
  NAND2_X1 U16273 ( .A1(n26566), .A2(n20577), .ZN(n20244) );
  INV_X2 U16290 ( .I(n27021), .ZN(n7968) );
  OR3_X2 U16291 ( .A1(n29306), .A2(n24171), .A3(n3483), .Z(n15781) );
  NOR2_X1 U16292 ( .A1(n1181), .A2(n339), .ZN(n11080) );
  OR2_X2 U16293 ( .A1(n30059), .A2(n28069), .Z(n23600) );
  INV_X1 U16295 ( .I(n15077), .ZN(n19961) );
  AND2_X1 U16298 ( .A1(n15077), .A2(n5870), .Z(n5871) );
  NAND2_X1 U16299 ( .A1(n8062), .A2(n4897), .ZN(n4999) );
  INV_X1 U16332 ( .I(n11707), .ZN(n328) );
  NOR2_X1 U16346 ( .A1(n10943), .A2(n31254), .ZN(n26037) );
  INV_X1 U16355 ( .I(n10943), .ZN(n11876) );
  NOR2_X1 U16358 ( .A1(n13129), .A2(n28942), .ZN(n13066) );
  INV_X1 U16376 ( .I(n10579), .ZN(n3152) );
  AND2_X2 U16377 ( .A1(n4036), .A2(n11599), .Z(n18812) );
  OR2_X2 U16383 ( .A1(n4036), .A2(n11599), .Z(n2733) );
  AOI22_X1 U16384 ( .A1(n18450), .A2(n17477), .B1(n18677), .B2(n18662), .ZN(
        n28943) );
  AOI21_X1 U16391 ( .A1(n17478), .A2(n18660), .B(n18677), .ZN(n31427) );
  NAND2_X1 U16396 ( .A1(n20635), .A2(n4693), .ZN(n30970) );
  AOI21_X1 U16398 ( .A1(n28408), .A2(n22949), .B(n805), .ZN(n6802) );
  NOR2_X1 U16400 ( .A1(n28555), .A2(n31129), .ZN(n17483) );
  NAND2_X2 U16403 ( .A1(n6950), .A2(n6952), .ZN(n8870) );
  AND2_X1 U16405 ( .A1(n31324), .A2(n19049), .Z(n12927) );
  NAND2_X2 U16406 ( .A1(n13752), .A2(n14859), .ZN(n31324) );
  INV_X2 U16408 ( .I(n13363), .ZN(n18581) );
  XOR2_X1 U16412 ( .A1(Plaintext[153]), .A2(Key[153]), .Z(n13363) );
  XOR2_X1 U16413 ( .A1(n5503), .A2(n5875), .Z(n31576) );
  XNOR2_X1 U16415 ( .A1(n22123), .A2(n13564), .ZN(n5875) );
  NAND2_X2 U16419 ( .A1(n14815), .A2(n14572), .ZN(n20124) );
  NAND2_X1 U16420 ( .A1(n31127), .A2(n31126), .ZN(n11706) );
  XNOR2_X1 U16424 ( .A1(n12868), .A2(n13236), .ZN(n1227) );
  XOR2_X1 U16445 ( .A1(n14682), .A2(n26575), .Z(n30338) );
  XOR2_X1 U16447 ( .A1(n32050), .A2(n30339), .Z(n6833) );
  XOR2_X1 U16448 ( .A1(n23294), .A2(n25815), .Z(n30339) );
  OAI21_X2 U16449 ( .A1(n17414), .A2(n30340), .B(n10848), .ZN(n28967) );
  NAND2_X2 U16453 ( .A1(n12449), .A2(n30341), .ZN(n23388) );
  AOI22_X1 U16455 ( .A1(n11210), .A2(n22961), .B1(n13396), .B2(n22962), .ZN(
        n30341) );
  XNOR2_X1 U16456 ( .A1(n21964), .A2(n2894), .ZN(n21951) );
  OAI21_X2 U16459 ( .A1(n26899), .A2(n10346), .B(n10343), .ZN(n2894) );
  AOI21_X2 U16473 ( .A1(n28306), .A2(n8760), .B(n30344), .ZN(n10500) );
  NOR2_X2 U16478 ( .A1(n5759), .A2(n23920), .ZN(n30344) );
  INV_X2 U16479 ( .I(n30345), .ZN(n30731) );
  XOR2_X1 U16483 ( .A1(n4136), .A2(n28446), .Z(n30345) );
  XOR2_X1 U16486 ( .A1(n20781), .A2(n20783), .Z(n3117) );
  NAND2_X1 U16494 ( .A1(n7485), .A2(n24312), .ZN(n30348) );
  XOR2_X1 U16499 ( .A1(n20746), .A2(n20993), .Z(n9815) );
  NAND3_X1 U16500 ( .A1(n10243), .A2(n10244), .A3(n11895), .ZN(n30349) );
  XOR2_X1 U16503 ( .A1(n22255), .A2(n30571), .Z(n7160) );
  NAND2_X1 U16525 ( .A1(n14174), .A2(n4518), .ZN(n16265) );
  NAND2_X2 U16537 ( .A1(n19450), .A2(n18089), .ZN(n3310) );
  OAI21_X1 U16543 ( .A1(n30353), .A2(n15746), .B(n22690), .ZN(n3451) );
  NOR2_X1 U16548 ( .A1(n1122), .A2(n31931), .ZN(n30353) );
  NAND2_X2 U16556 ( .A1(n1641), .A2(n26224), .ZN(n30354) );
  OAI21_X2 U16559 ( .A1(n30357), .A2(n30356), .B(n12947), .ZN(n20344) );
  OR2_X1 U16562 ( .A1(n18151), .A2(n15295), .Z(n25637) );
  XOR2_X1 U16563 ( .A1(n16158), .A2(n18109), .Z(n19552) );
  AOI22_X2 U16564 ( .A1(n2124), .A2(n28276), .B1(n30602), .B2(n2123), .ZN(
        n18109) );
  NOR2_X1 U16567 ( .A1(n515), .A2(n10433), .ZN(n4382) );
  NAND2_X2 U16573 ( .A1(n8897), .A2(n16797), .ZN(n14588) );
  AND2_X1 U16584 ( .A1(n31408), .A2(n19971), .Z(n31514) );
  NOR2_X1 U16586 ( .A1(n33809), .A2(n27491), .ZN(n30475) );
  NOR2_X2 U16597 ( .A1(n8062), .A2(n14490), .ZN(n24176) );
  AND2_X2 U16598 ( .A1(n18655), .A2(n32358), .Z(n18894) );
  BUF_X4 U16601 ( .I(n7600), .Z(n30602) );
  NAND2_X2 U16604 ( .A1(n21637), .A2(n21633), .ZN(n12792) );
  OAI21_X2 U16605 ( .A1(n5978), .A2(n21244), .B(n17803), .ZN(n21637) );
  BUF_X2 U16606 ( .I(n19991), .Z(n30366) );
  OAI21_X1 U16608 ( .A1(n29438), .A2(n23045), .B(n6553), .ZN(n29114) );
  XOR2_X1 U16611 ( .A1(n24551), .A2(n30367), .Z(n26754) );
  XOR2_X1 U16613 ( .A1(n24620), .A2(n16662), .Z(n30367) );
  INV_X1 U16621 ( .I(n8275), .ZN(n902) );
  XOR2_X1 U16623 ( .A1(n21927), .A2(n30368), .Z(n4859) );
  XOR2_X1 U16626 ( .A1(n10006), .A2(n8356), .Z(n30368) );
  XOR2_X1 U16634 ( .A1(n13661), .A2(n30370), .Z(n31098) );
  XOR2_X1 U16635 ( .A1(n14613), .A2(n24999), .Z(n30370) );
  NAND3_X1 U16648 ( .A1(n29958), .A2(n1577), .A3(n8334), .ZN(n14516) );
  AOI22_X2 U16659 ( .A1(n29383), .A2(n31653), .B1(n21744), .B2(n17021), .ZN(
        n17692) );
  INV_X2 U16690 ( .I(n17679), .ZN(n31493) );
  NAND2_X2 U16691 ( .A1(n17680), .A2(n17681), .ZN(n17679) );
  INV_X2 U16698 ( .I(n20818), .ZN(n31526) );
  NOR2_X2 U16703 ( .A1(n20246), .A2(n20245), .ZN(n20818) );
  NOR2_X2 U16704 ( .A1(n17685), .A2(n16282), .ZN(n21604) );
  XOR2_X1 U16716 ( .A1(n21937), .A2(n11819), .Z(n8596) );
  XOR2_X1 U16719 ( .A1(n22189), .A2(n22055), .Z(n21937) );
  OAI21_X1 U16726 ( .A1(n7197), .A2(n31970), .B(n825), .ZN(n17593) );
  NAND2_X2 U16728 ( .A1(n4025), .A2(n27341), .ZN(n13601) );
  AOI21_X2 U16730 ( .A1(n30379), .A2(n2574), .B(n32248), .ZN(n27973) );
  XOR2_X1 U16737 ( .A1(n8761), .A2(n30381), .Z(n29209) );
  XOR2_X1 U16738 ( .A1(n23536), .A2(n23189), .Z(n30381) );
  XOR2_X1 U16743 ( .A1(n30382), .A2(n31534), .Z(n14576) );
  XOR2_X1 U16747 ( .A1(n19653), .A2(n18051), .Z(n30382) );
  XOR2_X1 U16753 ( .A1(n30385), .A2(n8249), .Z(n8813) );
  XOR2_X1 U16754 ( .A1(n20654), .A2(n30045), .Z(n30385) );
  NAND2_X2 U16755 ( .A1(n3962), .A2(n13107), .ZN(n5748) );
  NOR2_X2 U16762 ( .A1(n30442), .A2(n773), .ZN(n31273) );
  XOR2_X1 U16765 ( .A1(n29244), .A2(n8972), .Z(n6957) );
  XOR2_X1 U16768 ( .A1(n6081), .A2(n30240), .Z(n8972) );
  NAND2_X2 U16781 ( .A1(n8245), .A2(n30386), .ZN(n8168) );
  INV_X2 U16783 ( .I(n30387), .ZN(n6344) );
  NAND2_X2 U16784 ( .A1(n15599), .A2(n15597), .ZN(n10174) );
  INV_X2 U16800 ( .I(n30390), .ZN(n15424) );
  INV_X2 U16808 ( .I(n7811), .ZN(n27685) );
  NAND2_X2 U16810 ( .A1(n4208), .A2(n12619), .ZN(n22964) );
  NAND2_X2 U16812 ( .A1(n7610), .A2(n28681), .ZN(n12619) );
  XOR2_X1 U16814 ( .A1(n10870), .A2(n24652), .Z(n24653) );
  OAI21_X2 U16826 ( .A1(n2604), .A2(n2605), .B(n30391), .ZN(n3286) );
  OAI21_X2 U16829 ( .A1(n2602), .A2(n2603), .B(n29207), .ZN(n30391) );
  OAI21_X2 U16833 ( .A1(n10735), .A2(n30441), .B(n11552), .ZN(n10935) );
  XOR2_X1 U16835 ( .A1(n23473), .A2(n770), .Z(n6094) );
  XOR2_X1 U16840 ( .A1(n1302), .A2(n22256), .Z(n4136) );
  XOR2_X1 U16844 ( .A1(n29898), .A2(n12459), .Z(n14875) );
  NAND2_X2 U16847 ( .A1(n30394), .A2(n10160), .ZN(n11789) );
  XOR2_X1 U16848 ( .A1(n28730), .A2(n30495), .Z(n11128) );
  XOR2_X1 U16856 ( .A1(n5127), .A2(n15236), .Z(n2362) );
  NAND2_X2 U16860 ( .A1(n8692), .A2(n19204), .ZN(n5127) );
  INV_X2 U16865 ( .I(n30047), .ZN(n25467) );
  INV_X2 U16874 ( .I(n25883), .ZN(n25872) );
  NOR3_X1 U16882 ( .A1(n30401), .A2(n19013), .A3(n19009), .ZN(n19014) );
  XOR2_X1 U16886 ( .A1(n24478), .A2(n24516), .Z(n24806) );
  NAND2_X2 U16888 ( .A1(n24166), .A2(n24165), .ZN(n24516) );
  NAND3_X1 U16895 ( .A1(n6497), .A2(n25643), .A3(n25658), .ZN(n26745) );
  XOR2_X1 U16908 ( .A1(n30402), .A2(n1604), .Z(n22224) );
  AOI22_X2 U16911 ( .A1(n5488), .A2(n67), .B1(n2574), .B2(n1632), .ZN(n30403)
         );
  NAND2_X2 U16939 ( .A1(n12746), .A2(n21423), .ZN(n5978) );
  XOR2_X1 U16940 ( .A1(n1338), .A2(n20843), .Z(n20674) );
  XOR2_X1 U16958 ( .A1(n8359), .A2(n28162), .Z(n8358) );
  INV_X1 U16973 ( .I(n7672), .ZN(n30973) );
  AOI22_X1 U16976 ( .A1(n12928), .A2(n27743), .B1(n13925), .B2(n12927), .ZN(
        n13002) );
  NAND2_X2 U16979 ( .A1(n19046), .A2(n19041), .ZN(n27743) );
  XOR2_X1 U16988 ( .A1(n16076), .A2(n30041), .Z(n23407) );
  XOR2_X1 U17002 ( .A1(n2592), .A2(n2590), .Z(n2589) );
  BUF_X2 U17005 ( .I(n31658), .Z(n30412) );
  NAND2_X2 U17030 ( .A1(n30417), .A2(n3508), .ZN(n7603) );
  XOR2_X1 U17037 ( .A1(n30418), .A2(n24937), .Z(Ciphertext[11]) );
  NAND2_X1 U17038 ( .A1(n7787), .A2(n31348), .ZN(n30418) );
  NOR2_X2 U17049 ( .A1(n7430), .A2(n12363), .ZN(n26268) );
  XOR2_X1 U17055 ( .A1(n23383), .A2(n30420), .Z(n27673) );
  XOR2_X1 U17056 ( .A1(n26426), .A2(n23536), .Z(n30420) );
  NOR2_X2 U17070 ( .A1(n30423), .A2(n25634), .ZN(n26581) );
  NOR2_X2 U17073 ( .A1(n11090), .A2(n3405), .ZN(n25632) );
  XOR2_X1 U17099 ( .A1(n30309), .A2(n32885), .Z(n22039) );
  OAI21_X1 U17100 ( .A1(n9472), .A2(n21870), .B(n5385), .ZN(n5384) );
  INV_X2 U17106 ( .I(n27655), .ZN(n2795) );
  XOR2_X1 U17107 ( .A1(n2796), .A2(n19687), .Z(n27655) );
  XOR2_X1 U17113 ( .A1(n7630), .A2(n7675), .Z(n30427) );
  NAND2_X2 U17117 ( .A1(n8995), .A2(n30428), .ZN(n8997) );
  AND2_X1 U17118 ( .A1(n10063), .A2(n8996), .Z(n30428) );
  NAND2_X2 U17123 ( .A1(n30429), .A2(n22822), .ZN(n9185) );
  NAND2_X1 U17125 ( .A1(n16203), .A2(n16202), .ZN(n30429) );
  NOR3_X1 U17126 ( .A1(n21872), .A2(n9472), .A3(n7811), .ZN(n4220) );
  AOI21_X2 U17143 ( .A1(n20247), .A2(n20248), .B(n17732), .ZN(n20717) );
  XOR2_X1 U17145 ( .A1(n1468), .A2(n1466), .Z(n25150) );
  XOR2_X1 U17180 ( .A1(n23419), .A2(n14819), .Z(n11290) );
  NAND2_X2 U17183 ( .A1(n31096), .A2(n14147), .ZN(n17941) );
  XOR2_X1 U17191 ( .A1(n30439), .A2(n16253), .Z(Ciphertext[117]) );
  NOR2_X1 U17194 ( .A1(n25511), .A2(n1945), .ZN(n30439) );
  INV_X2 U17195 ( .I(n21655), .ZN(n30441) );
  XOR2_X1 U17203 ( .A1(n27545), .A2(n8306), .Z(n24812) );
  INV_X2 U17216 ( .I(n30444), .ZN(n26606) );
  XOR2_X1 U17219 ( .A1(n3303), .A2(n3304), .Z(n30444) );
  INV_X2 U17220 ( .I(n30445), .ZN(n11272) );
  BUF_X2 U17226 ( .I(n15360), .Z(n31554) );
  NAND2_X2 U17227 ( .A1(n30446), .A2(n15745), .ZN(n9303) );
  NAND2_X2 U17236 ( .A1(n25581), .A2(n1082), .ZN(n15287) );
  OAI22_X2 U17238 ( .A1(n16413), .A2(n25707), .B1(n25621), .B2(n11944), .ZN(
        n25581) );
  AOI21_X2 U17239 ( .A1(n30641), .A2(n30448), .B(n22644), .ZN(n27867) );
  BUF_X4 U17241 ( .I(n3989), .Z(n31080) );
  NAND2_X2 U17249 ( .A1(n26990), .A2(n7360), .ZN(n7358) );
  XOR2_X1 U17284 ( .A1(n5509), .A2(n30453), .Z(n23157) );
  XOR2_X1 U17287 ( .A1(n5508), .A2(n29291), .Z(n30453) );
  AND2_X1 U17307 ( .A1(n16022), .A2(n14045), .Z(n28491) );
  XOR2_X1 U17317 ( .A1(n7234), .A2(n7235), .Z(n7453) );
  NAND2_X1 U17318 ( .A1(n5704), .A2(n15716), .ZN(n17333) );
  AOI21_X1 U17327 ( .A1(n25611), .A2(n27262), .B(n27528), .ZN(n30458) );
  OAI22_X1 U17331 ( .A1(n710), .A2(n3157), .B1(n28261), .B2(n30130), .ZN(n1964) );
  NOR2_X2 U17332 ( .A1(n6398), .A2(n16924), .ZN(n28261) );
  NAND2_X2 U17342 ( .A1(n28307), .A2(n30515), .ZN(n23974) );
  XOR2_X1 U17352 ( .A1(n14935), .A2(n30462), .Z(n5432) );
  XOR2_X1 U17355 ( .A1(n14937), .A2(n7829), .Z(n30462) );
  NOR2_X2 U17356 ( .A1(n1312), .A2(n21466), .ZN(n21465) );
  XOR2_X1 U17360 ( .A1(n5630), .A2(n5629), .Z(n30463) );
  XOR2_X1 U17364 ( .A1(n21026), .A2(n2525), .Z(n2524) );
  OR2_X2 U17365 ( .A1(n16440), .A2(n15559), .Z(n9073) );
  NAND2_X1 U17366 ( .A1(n31309), .A2(n11208), .ZN(n21708) );
  XOR2_X1 U17369 ( .A1(n30465), .A2(n12260), .Z(n29254) );
  XOR2_X1 U17371 ( .A1(n11062), .A2(n30466), .Z(n30465) );
  INV_X1 U17375 ( .I(n19748), .ZN(n30466) );
  OAI21_X2 U17382 ( .A1(n28757), .A2(n18609), .B(n18608), .ZN(n30467) );
  NOR2_X2 U17384 ( .A1(n31309), .A2(n21655), .ZN(n21797) );
  NAND2_X2 U17385 ( .A1(n30469), .A2(n7733), .ZN(n19332) );
  NAND2_X2 U17389 ( .A1(n2391), .A2(n20156), .ZN(n5470) );
  NAND2_X2 U17393 ( .A1(n31275), .A2(n5373), .ZN(n30470) );
  XOR2_X1 U17396 ( .A1(n1644), .A2(n1642), .Z(n23668) );
  NAND2_X2 U17406 ( .A1(n26956), .A2(n9046), .ZN(n14194) );
  XOR2_X1 U17409 ( .A1(n22150), .A2(n9208), .Z(n9207) );
  NAND2_X1 U17415 ( .A1(n30731), .A2(n11805), .ZN(n22544) );
  XOR2_X1 U17423 ( .A1(n24786), .A2(n24776), .Z(n24518) );
  NOR2_X2 U17425 ( .A1(n30475), .A2(n30474), .ZN(n20433) );
  NAND2_X2 U17428 ( .A1(n15074), .A2(n15073), .ZN(n19703) );
  NAND2_X1 U17437 ( .A1(n21847), .A2(n30291), .ZN(n30479) );
  NAND2_X2 U17439 ( .A1(n30480), .A2(n8459), .ZN(n9809) );
  OAI21_X2 U17440 ( .A1(n29405), .A2(n26298), .B(n1016), .ZN(n30480) );
  XOR2_X1 U17454 ( .A1(n20832), .A2(n8997), .Z(n18180) );
  OAI22_X1 U17461 ( .A1(n966), .A2(n25214), .B1(n5578), .B2(n16509), .ZN(
        n25223) );
  NOR2_X2 U17467 ( .A1(n26528), .A2(n18259), .ZN(n25214) );
  BUF_X2 U17469 ( .I(n5511), .Z(n30482) );
  NOR2_X1 U17472 ( .A1(n8334), .A2(n1577), .ZN(n11210) );
  XOR2_X1 U17474 ( .A1(n6052), .A2(n6054), .Z(n16757) );
  AOI22_X2 U17475 ( .A1(n8856), .A2(n21214), .B1(n15428), .B2(n21372), .ZN(
        n30483) );
  XOR2_X1 U17481 ( .A1(n30486), .A2(n2889), .Z(n30861) );
  BUF_X2 U17490 ( .I(n4219), .Z(n30489) );
  XOR2_X1 U17505 ( .A1(n23272), .A2(n5399), .Z(n23334) );
  AOI21_X2 U17508 ( .A1(n18073), .A2(n9456), .B(n29222), .ZN(n16260) );
  XOR2_X1 U17514 ( .A1(n30493), .A2(n30290), .Z(n24369) );
  OAI21_X2 U17517 ( .A1(n11637), .A2(n20575), .B(n20571), .ZN(n5590) );
  OR2_X1 U17518 ( .A1(n1877), .A2(n14436), .Z(n27605) );
  NAND2_X2 U17521 ( .A1(n28235), .A2(n11079), .ZN(n30505) );
  AOI21_X1 U17530 ( .A1(n25692), .A2(n25691), .B(n30494), .ZN(n30521) );
  AOI21_X1 U17534 ( .A1(n2017), .A2(n2016), .B(n26447), .ZN(n30494) );
  OAI22_X1 U17539 ( .A1(n30497), .A2(n17845), .B1(n25618), .B2(n10174), .ZN(
        n17844) );
  INV_X2 U17540 ( .I(n30498), .ZN(n490) );
  XOR2_X1 U17542 ( .A1(Plaintext[151]), .A2(Key[151]), .Z(n30498) );
  XOR2_X1 U17545 ( .A1(n19544), .A2(n19545), .Z(n13441) );
  BUF_X2 U17553 ( .I(n23066), .Z(n30502) );
  NAND2_X1 U17568 ( .A1(n10812), .A2(n30508), .ZN(n23965) );
  OR2_X1 U17575 ( .A1(n31155), .A2(n11754), .Z(n30508) );
  OAI21_X2 U17592 ( .A1(n30511), .A2(n21514), .B(n30243), .ZN(n31404) );
  XOR2_X1 U17593 ( .A1(n30513), .A2(n29082), .Z(n28640) );
  XOR2_X1 U17595 ( .A1(n27875), .A2(n11897), .Z(n30513) );
  XOR2_X1 U17608 ( .A1(n32564), .A2(n30306), .Z(n15822) );
  NAND2_X2 U17610 ( .A1(n21525), .A2(n21524), .ZN(n22306) );
  XOR2_X1 U17614 ( .A1(n20808), .A2(n20645), .Z(n30514) );
  XOR2_X1 U17630 ( .A1(n24756), .A2(n30517), .Z(n1466) );
  XOR2_X1 U17632 ( .A1(n30358), .A2(n30069), .Z(n30517) );
  NOR2_X1 U17641 ( .A1(n15283), .A2(n9934), .ZN(n9847) );
  NAND2_X1 U17648 ( .A1(n33928), .A2(n28934), .ZN(n28349) );
  XOR2_X1 U17650 ( .A1(n30521), .A2(n25694), .Z(Ciphertext[148]) );
  AOI22_X2 U17654 ( .A1(n27565), .A2(n12254), .B1(n29232), .B2(n12256), .ZN(
        n8040) );
  XOR2_X1 U17656 ( .A1(n17775), .A2(n23218), .Z(n23399) );
  INV_X1 U17660 ( .I(n7503), .ZN(n30586) );
  AND2_X1 U17664 ( .A1(n29270), .A2(n14398), .Z(n6759) );
  XOR2_X1 U17667 ( .A1(n15710), .A2(n16253), .Z(n30524) );
  AOI22_X1 U17686 ( .A1(n14434), .A2(n1206), .B1(n690), .B2(n25916), .ZN(
        n14433) );
  XOR2_X1 U17693 ( .A1(n27841), .A2(n30069), .Z(n24418) );
  INV_X2 U17708 ( .I(n30526), .ZN(n17963) );
  XOR2_X1 U17710 ( .A1(n17703), .A2(n29450), .Z(n26597) );
  INV_X2 U17721 ( .I(n1994), .ZN(n16138) );
  NOR2_X2 U17723 ( .A1(n11770), .A2(n13859), .ZN(n11769) );
  XOR2_X1 U17729 ( .A1(n16831), .A2(n3629), .Z(n20894) );
  XNOR2_X1 U17736 ( .A1(n21946), .A2(n10370), .ZN(n30575) );
  AOI21_X2 U17744 ( .A1(n16883), .A2(n20220), .B(n30530), .ZN(n14428) );
  XOR2_X1 U17770 ( .A1(n2854), .A2(n30317), .Z(n30535) );
  XOR2_X1 U17772 ( .A1(n30536), .A2(n4719), .Z(n17903) );
  XOR2_X1 U17773 ( .A1(n24797), .A2(n12239), .Z(n30536) );
  XOR2_X1 U17776 ( .A1(n18024), .A2(n18025), .Z(n11677) );
  NAND2_X2 U17789 ( .A1(n30537), .A2(n29406), .ZN(n3773) );
  NOR2_X2 U17793 ( .A1(n30538), .A2(n17584), .ZN(n30537) );
  AOI21_X2 U17795 ( .A1(n6876), .A2(n23032), .B(n31273), .ZN(n14610) );
  XOR2_X1 U17806 ( .A1(n14103), .A2(n30541), .Z(n23639) );
  XOR2_X1 U17815 ( .A1(n23446), .A2(n11667), .Z(n30541) );
  XOR2_X1 U17820 ( .A1(n4797), .A2(n30542), .Z(n9750) );
  XOR2_X1 U17823 ( .A1(n22110), .A2(n13437), .Z(n30542) );
  XOR2_X1 U17832 ( .A1(n20856), .A2(n20785), .Z(n9040) );
  INV_X1 U17833 ( .I(n29263), .ZN(n1122) );
  XOR2_X1 U17836 ( .A1(n27792), .A2(n5126), .Z(n29263) );
  XOR2_X1 U17850 ( .A1(n16893), .A2(n22264), .Z(n6058) );
  OAI21_X2 U17852 ( .A1(n30546), .A2(n28911), .B(n4602), .ZN(n20569) );
  XOR2_X1 U17859 ( .A1(n23113), .A2(n13123), .Z(n30547) );
  OAI21_X2 U17861 ( .A1(n276), .A2(n517), .B(n21777), .ZN(n30548) );
  XOR2_X1 U17868 ( .A1(n22198), .A2(n22197), .Z(n14755) );
  BUF_X2 U17870 ( .I(n21592), .Z(n30549) );
  XOR2_X1 U17878 ( .A1(n32881), .A2(n28005), .Z(n30550) );
  OAI22_X2 U17883 ( .A1(n1908), .A2(n31374), .B1(n30552), .B2(n30551), .ZN(
        n5647) );
  XOR2_X1 U17888 ( .A1(n13321), .A2(n5742), .Z(n23471) );
  NAND2_X2 U17890 ( .A1(n10849), .A2(n31454), .ZN(n30553) );
  BUF_X2 U17896 ( .I(n27097), .Z(n30554) );
  XOR2_X1 U17899 ( .A1(n30556), .A2(n5980), .Z(n5979) );
  XOR2_X1 U17910 ( .A1(n28315), .A2(n30557), .Z(n30556) );
  NAND2_X2 U17918 ( .A1(n14774), .A2(n14776), .ZN(n28934) );
  XOR2_X1 U17926 ( .A1(n26094), .A2(n16700), .Z(n30559) );
  NOR2_X2 U17927 ( .A1(n9133), .A2(n31040), .ZN(n21152) );
  INV_X2 U17934 ( .I(n30563), .ZN(n16738) );
  NAND2_X1 U17940 ( .A1(n5991), .A2(n28825), .ZN(n30564) );
  XOR2_X1 U17947 ( .A1(n23355), .A2(n31554), .Z(n30565) );
  XOR2_X1 U17953 ( .A1(n19473), .A2(n32267), .Z(n9577) );
  NAND2_X1 U17954 ( .A1(n29424), .A2(n26803), .ZN(n30658) );
  NAND2_X1 U17957 ( .A1(n9990), .A2(n10098), .ZN(n30587) );
  OAI21_X2 U17962 ( .A1(n30569), .A2(n30568), .B(n11992), .ZN(n9982) );
  AOI22_X1 U17963 ( .A1(n6825), .A2(n14922), .B1(n13273), .B2(n9162), .ZN(
        n6824) );
  NAND2_X2 U17973 ( .A1(n8743), .A2(n25109), .ZN(n25128) );
  NAND2_X2 U17980 ( .A1(n18205), .A2(n6228), .ZN(n20835) );
  NAND2_X1 U17984 ( .A1(n25944), .A2(n8253), .ZN(n11597) );
  INV_X2 U17985 ( .I(n30570), .ZN(n1736) );
  NAND2_X2 U17997 ( .A1(n7550), .A2(n7551), .ZN(n8770) );
  XOR2_X1 U17999 ( .A1(n19668), .A2(n253), .Z(n4883) );
  AOI21_X2 U18001 ( .A1(n10073), .A2(n28104), .B(n14757), .ZN(n19668) );
  XOR2_X1 U18008 ( .A1(n16727), .A2(n6488), .Z(n19660) );
  OR2_X1 U18018 ( .A1(n20109), .A2(n28183), .Z(n30614) );
  XOR2_X1 U18022 ( .A1(n10917), .A2(n30574), .Z(n10916) );
  XOR2_X1 U18023 ( .A1(n31750), .A2(n9434), .Z(n30574) );
  XOR2_X1 U18034 ( .A1(n10154), .A2(n30575), .Z(n28589) );
  NAND2_X1 U18040 ( .A1(n31306), .A2(n5477), .ZN(n15193) );
  INV_X1 U18044 ( .I(n9107), .ZN(n23096) );
  NOR2_X1 U18068 ( .A1(n12973), .A2(n21241), .ZN(n11405) );
  INV_X1 U18071 ( .I(n21330), .ZN(n12973) );
  XOR2_X1 U18082 ( .A1(n20778), .A2(n13725), .Z(n13724) );
  NOR2_X2 U18087 ( .A1(n19172), .A2(n19078), .ZN(n11875) );
  NAND2_X2 U18092 ( .A1(n1376), .A2(n10943), .ZN(n19172) );
  XOR2_X1 U18106 ( .A1(n20925), .A2(n20927), .Z(n7032) );
  XOR2_X1 U18112 ( .A1(n2520), .A2(n31394), .Z(n23126) );
  NAND2_X2 U18116 ( .A1(n18160), .A2(n18162), .ZN(n30995) );
  NOR3_X1 U18126 ( .A1(n25026), .A2(n25025), .A3(n25024), .ZN(n31320) );
  XOR2_X1 U18128 ( .A1(n24424), .A2(n4720), .Z(n4719) );
  XOR2_X1 U18134 ( .A1(n7731), .A2(n24440), .Z(n24424) );
  XOR2_X1 U18136 ( .A1(n30583), .A2(n25038), .Z(Ciphertext[37]) );
  NOR2_X2 U18142 ( .A1(n24008), .A2(n10033), .ZN(n26027) );
  NAND2_X2 U18147 ( .A1(n31163), .A2(n27679), .ZN(n27676) );
  NOR2_X1 U18149 ( .A1(n14133), .A2(n29203), .ZN(n14529) );
  NAND3_X1 U18150 ( .A1(n7302), .A2(n7299), .A3(n7298), .ZN(Ciphertext[72]) );
  NAND2_X2 U18157 ( .A1(n1172), .A2(n7573), .ZN(n19850) );
  OAI21_X2 U18176 ( .A1(n7001), .A2(n26088), .B(n2271), .ZN(n6996) );
  XOR2_X1 U18178 ( .A1(n13198), .A2(n29457), .Z(n27868) );
  OAI21_X2 U18187 ( .A1(n31938), .A2(n14513), .B(n16099), .ZN(n1776) );
  NOR2_X2 U18188 ( .A1(n15038), .A2(n976), .ZN(n14513) );
  OAI22_X1 U18211 ( .A1(n898), .A2(n23066), .B1(n849), .B2(n4067), .ZN(n4477)
         );
  INV_X2 U18222 ( .I(n30592), .ZN(n12120) );
  XOR2_X1 U18224 ( .A1(n18280), .A2(Key[64]), .Z(n30592) );
  INV_X2 U18232 ( .I(n30593), .ZN(n6444) );
  NAND2_X2 U18241 ( .A1(n5945), .A2(n29044), .ZN(n6488) );
  BUF_X2 U18242 ( .I(n14123), .Z(n30595) );
  XOR2_X1 U18245 ( .A1(n30596), .A2(n23507), .Z(n31429) );
  XOR2_X1 U18256 ( .A1(n30597), .A2(n4186), .Z(n11749) );
  XOR2_X1 U18257 ( .A1(n11748), .A2(n21944), .Z(n30597) );
  NAND2_X2 U18260 ( .A1(n23627), .A2(n23626), .ZN(n24479) );
  XOR2_X1 U18264 ( .A1(n22302), .A2(n10292), .Z(n7289) );
  NAND2_X2 U18271 ( .A1(n2338), .A2(n31051), .ZN(n10292) );
  XOR2_X1 U18272 ( .A1(n7363), .A2(n23332), .Z(n23383) );
  OAI22_X2 U18275 ( .A1(n30598), .A2(n9066), .B1(n24199), .B2(n12574), .ZN(
        n24764) );
  XOR2_X1 U18282 ( .A1(n30601), .A2(n30600), .Z(n26551) );
  XOR2_X1 U18286 ( .A1(n13842), .A2(n19447), .Z(n30601) );
  XOR2_X1 U18307 ( .A1(n23162), .A2(n6169), .Z(n1796) );
  NAND3_X2 U18314 ( .A1(n30608), .A2(n28158), .A3(n28159), .ZN(n22149) );
  XOR2_X1 U18326 ( .A1(n30610), .A2(n5107), .Z(n5106) );
  XOR2_X1 U18336 ( .A1(n33572), .A2(n5109), .Z(n30610) );
  INV_X1 U18344 ( .I(n16109), .ZN(n31167) );
  NOR2_X2 U18359 ( .A1(n5308), .A2(n7546), .ZN(n24046) );
  NAND2_X2 U18367 ( .A1(n30615), .A2(n25149), .ZN(n25151) );
  XOR2_X1 U18380 ( .A1(n5336), .A2(n6604), .Z(n10932) );
  NAND2_X1 U18383 ( .A1(n26237), .A2(n820), .ZN(n9232) );
  AND2_X2 U18385 ( .A1(n18186), .A2(n16417), .Z(n18370) );
  NOR2_X1 U18391 ( .A1(n31823), .A2(n20045), .ZN(n30617) );
  NAND2_X2 U18397 ( .A1(n30618), .A2(n39), .ZN(n23368) );
  OAI21_X2 U18398 ( .A1(n10885), .A2(n16236), .B(n22900), .ZN(n30618) );
  NAND3_X2 U18433 ( .A1(n29335), .A2(n28472), .A3(n28473), .ZN(n31181) );
  NAND3_X2 U18434 ( .A1(n30623), .A2(n13161), .A3(n30622), .ZN(n13651) );
  XOR2_X1 U18445 ( .A1(n19546), .A2(n19591), .Z(n3285) );
  NAND2_X1 U18450 ( .A1(n18184), .A2(n28232), .ZN(n9205) );
  NAND2_X2 U18451 ( .A1(n30624), .A2(n2908), .ZN(n20445) );
  OR2_X2 U18453 ( .A1(n4735), .A2(n31287), .Z(n2538) );
  NAND2_X2 U18454 ( .A1(n11069), .A2(n3430), .ZN(n5533) );
  NOR2_X2 U18455 ( .A1(n29353), .A2(n30625), .ZN(n10302) );
  NAND2_X1 U18460 ( .A1(n5640), .A2(n33594), .ZN(n22338) );
  NAND2_X2 U18464 ( .A1(n30626), .A2(n4872), .ZN(n24544) );
  OR3_X1 U18471 ( .A1(n2958), .A2(n868), .A3(n8374), .Z(n28353) );
  NOR2_X1 U18476 ( .A1(n15564), .A2(n11912), .ZN(n30627) );
  OAI22_X2 U18485 ( .A1(n31149), .A2(n25561), .B1(n25562), .B2(n25331), .ZN(
        n25523) );
  NAND3_X2 U18495 ( .A1(n6645), .A2(n6643), .A3(n14171), .ZN(n20267) );
  XOR2_X1 U18515 ( .A1(n13084), .A2(n13085), .Z(n16913) );
  XOR2_X1 U18528 ( .A1(n20924), .A2(n20885), .Z(n14899) );
  NAND2_X2 U18532 ( .A1(n28452), .A2(n28454), .ZN(n14436) );
  AOI21_X2 U18542 ( .A1(n14076), .A2(n4262), .B(n8784), .ZN(n30634) );
  XOR2_X1 U18547 ( .A1(n30635), .A2(n4401), .Z(n564) );
  INV_X2 U18553 ( .I(n10915), .ZN(n30636) );
  AND2_X1 U18558 ( .A1(n20479), .A2(n11637), .Z(n28226) );
  AOI21_X1 U18563 ( .A1(n22872), .A2(n15718), .B(n30638), .ZN(n30800) );
  XOR2_X1 U18568 ( .A1(n22218), .A2(n1131), .Z(n1716) );
  NAND2_X2 U18577 ( .A1(n21292), .A2(n21291), .ZN(n6669) );
  XOR2_X1 U18586 ( .A1(n16150), .A2(n13435), .Z(n30644) );
  NOR2_X2 U18588 ( .A1(n30645), .A2(n29084), .ZN(n8337) );
  NAND2_X2 U18589 ( .A1(n30940), .A2(n517), .ZN(n30645) );
  NAND2_X1 U18592 ( .A1(n3203), .A2(n30677), .ZN(n26207) );
  NAND2_X2 U18600 ( .A1(n3001), .A2(n3003), .ZN(n3203) );
  AOI22_X2 U18620 ( .A1(n31990), .A2(n31175), .B1(n23788), .B2(n15272), .ZN(
        n30649) );
  NAND2_X1 U18629 ( .A1(n1134), .A2(n30652), .ZN(n12995) );
  OAI21_X2 U18642 ( .A1(n31934), .A2(n13127), .B(n22444), .ZN(n22878) );
  XOR2_X1 U18646 ( .A1(n30653), .A2(n16030), .Z(n3686) );
  XOR2_X1 U18647 ( .A1(n6094), .A2(n17628), .Z(n30653) );
  XOR2_X1 U18656 ( .A1(n19636), .A2(n19635), .Z(n19640) );
  XOR2_X1 U18658 ( .A1(n22317), .A2(n156), .Z(n21924) );
  NOR2_X2 U18659 ( .A1(n21562), .A2(n21561), .ZN(n156) );
  XOR2_X1 U18668 ( .A1(n4574), .A2(n4572), .Z(n24726) );
  INV_X4 U18671 ( .I(n11521), .ZN(n13747) );
  INV_X1 U18675 ( .I(n27262), .ZN(n17845) );
  NAND2_X2 U18685 ( .A1(n18192), .A2(n25585), .ZN(n27262) );
  INV_X2 U18695 ( .I(n16847), .ZN(n30663) );
  OR2_X1 U18698 ( .A1(n30663), .A2(n2581), .Z(n30936) );
  INV_X1 U18699 ( .I(n22312), .ZN(n31203) );
  INV_X2 U18700 ( .I(n18397), .ZN(n18687) );
  XOR2_X1 U18703 ( .A1(n18396), .A2(Key[183]), .Z(n18397) );
  XOR2_X1 U18704 ( .A1(n19667), .A2(n19666), .Z(n17689) );
  XOR2_X1 U18710 ( .A1(n12048), .A2(n5462), .Z(n19667) );
  XOR2_X1 U18713 ( .A1(n26530), .A2(n21007), .Z(n30664) );
  NAND2_X2 U18719 ( .A1(n30824), .A2(n12465), .ZN(n28580) );
  INV_X2 U18729 ( .I(n14600), .ZN(n9293) );
  AOI22_X2 U18735 ( .A1(n22375), .A2(n9411), .B1(n25947), .B2(n22479), .ZN(
        n23000) );
  INV_X2 U18737 ( .I(n9168), .ZN(n30668) );
  NOR2_X1 U18740 ( .A1(n31150), .A2(n28949), .ZN(n30670) );
  XOR2_X1 U18744 ( .A1(n28086), .A2(n6790), .Z(n31040) );
  AOI21_X2 U18751 ( .A1(n24712), .A2(n24711), .B(n1077), .ZN(n25678) );
  OAI22_X1 U18765 ( .A1(n1028), .A2(n7774), .B1(n2237), .B2(n7218), .ZN(n9693)
         );
  INV_X2 U18766 ( .I(n11089), .ZN(n3405) );
  XOR2_X1 U18783 ( .A1(n24749), .A2(n5525), .Z(n30676) );
  NAND2_X2 U18797 ( .A1(n27232), .A2(n23547), .ZN(n24283) );
  INV_X4 U18799 ( .I(n31668), .ZN(n1351) );
  NAND2_X2 U18801 ( .A1(n7820), .A2(n28622), .ZN(n31668) );
  NAND2_X1 U18807 ( .A1(n30961), .A2(n5866), .ZN(n30777) );
  XOR2_X1 U18808 ( .A1(n30679), .A2(n18932), .Z(n26815) );
  NAND2_X2 U18810 ( .A1(n14084), .A2(n19968), .ZN(n20384) );
  NOR2_X2 U18811 ( .A1(n13770), .A2(n27878), .ZN(n30681) );
  BUF_X2 U18819 ( .I(n31324), .Z(n30682) );
  XOR2_X1 U18826 ( .A1(n15516), .A2(n20691), .Z(n8682) );
  OAI22_X1 U18832 ( .A1(n20332), .A2(n28390), .B1(n20549), .B2(n11710), .ZN(
        n11709) );
  XOR2_X1 U18833 ( .A1(n15329), .A2(n16506), .Z(n10443) );
  NAND2_X2 U18835 ( .A1(n12908), .A2(n12909), .ZN(n15329) );
  INV_X2 U18836 ( .I(n7012), .ZN(n14251) );
  XOR2_X1 U18840 ( .A1(n11889), .A2(n29312), .Z(n14820) );
  NAND2_X2 U18841 ( .A1(n19311), .A2(n19312), .ZN(n11889) );
  XOR2_X1 U18842 ( .A1(n15236), .A2(n19668), .Z(n13863) );
  AOI21_X2 U18845 ( .A1(n12798), .A2(n10452), .B(n10451), .ZN(n15236) );
  XOR2_X1 U18846 ( .A1(n28121), .A2(n30685), .Z(n3106) );
  XOR2_X1 U18851 ( .A1(n10081), .A2(n29205), .Z(n30685) );
  NOR2_X2 U18853 ( .A1(n10828), .A2(n1377), .ZN(n19309) );
  INV_X2 U18854 ( .I(n19308), .ZN(n1377) );
  NOR3_X1 U18866 ( .A1(n33722), .A2(n23813), .A3(n8166), .ZN(n30687) );
  XOR2_X1 U18898 ( .A1(n7677), .A2(n19712), .Z(n9517) );
  NAND3_X2 U18901 ( .A1(n2585), .A2(n8672), .A3(n2587), .ZN(n19712) );
  XOR2_X1 U18902 ( .A1(n23270), .A2(n23269), .Z(n31034) );
  INV_X2 U18904 ( .I(n12287), .ZN(n13720) );
  XOR2_X1 U18912 ( .A1(n47), .A2(n12288), .Z(n12287) );
  NAND2_X2 U18916 ( .A1(n21804), .A2(n11231), .ZN(n115) );
  NAND2_X2 U18922 ( .A1(n12711), .A2(n12712), .ZN(n21804) );
  INV_X2 U18923 ( .I(n30690), .ZN(n31911) );
  NAND3_X2 U18931 ( .A1(n21119), .A2(n7913), .A3(n21118), .ZN(n30690) );
  XOR2_X1 U18933 ( .A1(n30691), .A2(n9911), .Z(n31839) );
  XOR2_X1 U18935 ( .A1(n11271), .A2(n22287), .Z(n30691) );
  OAI21_X2 U18938 ( .A1(n30693), .A2(n30692), .B(n16789), .ZN(n30923) );
  XOR2_X1 U18940 ( .A1(n23297), .A2(n1825), .Z(n23119) );
  AND2_X1 U18950 ( .A1(n3251), .A2(n31012), .Z(n14314) );
  NAND2_X2 U18951 ( .A1(n2186), .A2(n30695), .ZN(n2864) );
  XOR2_X1 U18963 ( .A1(n7256), .A2(n30540), .Z(n24540) );
  OAI21_X2 U18970 ( .A1(n30698), .A2(n30697), .B(n31012), .ZN(n12977) );
  OAI21_X2 U18972 ( .A1(n30700), .A2(n30699), .B(n13968), .ZN(n14983) );
  NOR2_X1 U18979 ( .A1(n3042), .A2(n31201), .ZN(n3045) );
  XOR2_X1 U18981 ( .A1(n6792), .A2(n30702), .Z(n7368) );
  XOR2_X1 U18982 ( .A1(n7870), .A2(n13181), .Z(n30702) );
  NAND2_X2 U19002 ( .A1(n16552), .A2(n24056), .ZN(n26374) );
  NAND2_X2 U19004 ( .A1(n4483), .A2(n4481), .ZN(n24056) );
  NAND2_X2 U19009 ( .A1(n8482), .A2(n18294), .ZN(n27921) );
  XNOR2_X1 U19010 ( .A1(n2304), .A2(n21022), .ZN(n30849) );
  XOR2_X1 U19019 ( .A1(n23467), .A2(n9185), .Z(n16200) );
  XOR2_X1 U19020 ( .A1(n11862), .A2(n22205), .Z(n22153) );
  OAI22_X2 U19022 ( .A1(n10493), .A2(n28729), .B1(n5495), .B2(n10492), .ZN(
        n22205) );
  AOI21_X2 U19028 ( .A1(n6505), .A2(n30703), .B(n9777), .ZN(n5035) );
  NAND2_X2 U19036 ( .A1(n30748), .A2(n28857), .ZN(n30705) );
  XOR2_X1 U19042 ( .A1(n20810), .A2(n20809), .Z(n30706) );
  XOR2_X1 U19046 ( .A1(n29140), .A2(n30707), .Z(n1642) );
  XOR2_X1 U19049 ( .A1(n3295), .A2(n9468), .Z(n30707) );
  XOR2_X1 U19052 ( .A1(n22154), .A2(n7685), .Z(n7684) );
  NAND2_X1 U19061 ( .A1(n3343), .A2(n743), .ZN(n30710) );
  OR2_X2 U19062 ( .A1(n7), .A2(n21970), .Z(n22488) );
  XOR2_X1 U19064 ( .A1(n8809), .A2(n30711), .Z(n8806) );
  XOR2_X1 U19069 ( .A1(n31138), .A2(n30712), .Z(n30711) );
  INV_X2 U19071 ( .I(n30713), .ZN(n21412) );
  XOR2_X1 U19073 ( .A1(n22008), .A2(n30714), .Z(n27160) );
  XOR2_X1 U19076 ( .A1(n22288), .A2(n22006), .Z(n30714) );
  NOR2_X2 U19083 ( .A1(n30716), .A2(n17016), .ZN(n30732) );
  NAND2_X2 U19088 ( .A1(n24047), .A2(n8567), .ZN(n30716) );
  OR2_X1 U19089 ( .A1(n9073), .A2(n21428), .Z(n17415) );
  NOR3_X2 U19091 ( .A1(n6414), .A2(n14975), .A3(n14974), .ZN(n30717) );
  AOI21_X1 U19092 ( .A1(n1284), .A2(n6976), .B(n30718), .ZN(n2348) );
  INV_X2 U19096 ( .I(n980), .ZN(n30720) );
  XOR2_X1 U19104 ( .A1(n13208), .A2(n30721), .Z(n21432) );
  XOR2_X1 U19105 ( .A1(n20967), .A2(n30722), .Z(n30721) );
  AOI21_X2 U19106 ( .A1(n29398), .A2(n15505), .B(n30760), .ZN(n19273) );
  XOR2_X1 U19107 ( .A1(n30723), .A2(n19687), .Z(n5837) );
  XOR2_X1 U19109 ( .A1(n5236), .A2(n19430), .Z(n30723) );
  NOR3_X2 U19110 ( .A1(n17211), .A2(n28214), .A3(n22705), .ZN(n30724) );
  NAND2_X1 U19112 ( .A1(n23640), .A2(n14078), .ZN(n30725) );
  NAND2_X2 U19118 ( .A1(n30931), .A2(n16684), .ZN(n27317) );
  BUF_X2 U19121 ( .I(n31040), .Z(n30727) );
  OR2_X1 U19127 ( .A1(n32051), .A2(n5225), .Z(n18352) );
  OAI22_X2 U19146 ( .A1(n9741), .A2(n9740), .B1(n5764), .B2(n23788), .ZN(n7581) );
  NAND3_X2 U19158 ( .A1(n7324), .A2(n21519), .A3(n7323), .ZN(n22028) );
  XOR2_X1 U19168 ( .A1(n14742), .A2(n19503), .Z(n17434) );
  BUF_X2 U19177 ( .I(n31882), .Z(n30729) );
  NAND2_X2 U19181 ( .A1(n15123), .A2(n6605), .ZN(n22946) );
  OAI22_X2 U19185 ( .A1(n12601), .A2(n28705), .B1(n12131), .B2(n12600), .ZN(
        n19370) );
  INV_X1 U19187 ( .I(n30730), .ZN(n8631) );
  NAND2_X2 U19198 ( .A1(n31223), .A2(n6667), .ZN(n339) );
  OAI21_X2 U19199 ( .A1(n2409), .A2(n2408), .B(n2407), .ZN(n13762) );
  NAND2_X2 U19206 ( .A1(n7798), .A2(n14945), .ZN(n17837) );
  XOR2_X1 U19208 ( .A1(n22085), .A2(n6462), .Z(n17377) );
  AND2_X1 U19213 ( .A1(n632), .A2(n10681), .Z(n15763) );
  NAND3_X2 U19216 ( .A1(n31963), .A2(n29078), .A3(n123), .ZN(n26324) );
  AND2_X1 U19217 ( .A1(n23843), .A2(n299), .Z(n14088) );
  NAND2_X1 U19220 ( .A1(n20339), .A2(n15169), .ZN(n15042) );
  NAND2_X2 U19238 ( .A1(n11090), .A2(n3405), .ZN(n25565) );
  XOR2_X1 U19250 ( .A1(n23342), .A2(n30733), .Z(n23136) );
  NOR2_X1 U19251 ( .A1(n1348), .A2(n19402), .ZN(n26358) );
  XOR2_X1 U19256 ( .A1(n30734), .A2(n31321), .Z(n14726) );
  OAI21_X2 U19266 ( .A1(n30737), .A2(n30736), .B(n23864), .ZN(n17183) );
  NOR2_X2 U19288 ( .A1(n19023), .A2(n19020), .ZN(n27726) );
  AOI21_X2 U19292 ( .A1(n3429), .A2(n732), .B(n2682), .ZN(n19023) );
  XOR2_X1 U19293 ( .A1(n9848), .A2(n24567), .Z(n8575) );
  NOR2_X2 U19298 ( .A1(n23404), .A2(n30741), .ZN(n5505) );
  XOR2_X1 U19299 ( .A1(n30742), .A2(n25880), .Z(Ciphertext[182]) );
  OAI22_X1 U19303 ( .A1(n5303), .A2(n25995), .B1(n5301), .B2(n5300), .ZN(
        n30742) );
  XOR2_X1 U19311 ( .A1(n30746), .A2(n16555), .Z(Ciphertext[103]) );
  AND2_X1 U19321 ( .A1(n3911), .A2(n22420), .Z(n30758) );
  NAND3_X1 U19334 ( .A1(n17087), .A2(n23764), .A3(n1101), .ZN(n17088) );
  XOR2_X1 U19340 ( .A1(n11062), .A2(n15297), .Z(n1941) );
  NAND2_X1 U19341 ( .A1(n7486), .A2(n28166), .ZN(n20553) );
  AOI21_X2 U19344 ( .A1(n27372), .A2(n29317), .B(n30753), .ZN(n26656) );
  NAND2_X2 U19345 ( .A1(n30754), .A2(n28956), .ZN(n24289) );
  INV_X2 U19356 ( .I(n12945), .ZN(n1231) );
  NAND2_X2 U19358 ( .A1(n7246), .A2(n27480), .ZN(n12945) );
  XOR2_X1 U19367 ( .A1(n30757), .A2(n19417), .Z(n11591) );
  NOR2_X2 U19372 ( .A1(n29156), .A2(n19884), .ZN(n13840) );
  XOR2_X1 U19377 ( .A1(n11545), .A2(n11543), .Z(n20152) );
  BUF_X2 U19378 ( .I(n19268), .Z(n30760) );
  XOR2_X1 U19411 ( .A1(n112), .A2(n30766), .Z(n30765) );
  XOR2_X1 U19420 ( .A1(n15424), .A2(n23411), .Z(n30767) );
  XOR2_X1 U19428 ( .A1(n20753), .A2(n15557), .Z(n15556) );
  OAI22_X1 U19434 ( .A1(n19079), .A2(n34005), .B1(n19080), .B2(n948), .ZN(
        n30768) );
  NAND3_X1 U19437 ( .A1(n13286), .A2(n17624), .A3(n21338), .ZN(n2242) );
  NAND2_X2 U19441 ( .A1(n8489), .A2(n14326), .ZN(n31254) );
  INV_X2 U19444 ( .I(n30770), .ZN(n14458) );
  XOR2_X1 U19464 ( .A1(n19736), .A2(n19654), .Z(n7887) );
  NAND2_X2 U19468 ( .A1(n10532), .A2(n4098), .ZN(n11231) );
  XOR2_X1 U19472 ( .A1(n5146), .A2(n30776), .Z(n31747) );
  XOR2_X1 U19473 ( .A1(n24741), .A2(n16381), .Z(n30776) );
  XOR2_X1 U19474 ( .A1(n30777), .A2(n24895), .Z(Ciphertext[47]) );
  XOR2_X1 U19477 ( .A1(n1938), .A2(n1935), .Z(n9870) );
  OR2_X2 U19480 ( .A1(n26345), .A2(n4740), .Z(n21173) );
  NAND2_X2 U19483 ( .A1(n30780), .A2(n31694), .ZN(n16804) );
  OAI22_X2 U19485 ( .A1(n4142), .A2(n16812), .B1(n20044), .B2(n20045), .ZN(
        n30780) );
  XOR2_X1 U19510 ( .A1(n21996), .A2(n8356), .Z(n15726) );
  XOR2_X1 U19525 ( .A1(n11304), .A2(n20773), .Z(n28621) );
  INV_X2 U19528 ( .I(n14383), .ZN(n21358) );
  XOR2_X1 U19535 ( .A1(n3010), .A2(n11530), .Z(n14383) );
  NAND2_X2 U19540 ( .A1(n31036), .A2(n10297), .ZN(n19743) );
  NAND2_X1 U19542 ( .A1(n1734), .A2(n1733), .ZN(n30792) );
  XOR2_X1 U19548 ( .A1(n22252), .A2(n21919), .Z(n7686) );
  NAND2_X2 U19550 ( .A1(n20089), .A2(n5405), .ZN(n2271) );
  NAND2_X2 U19551 ( .A1(n31046), .A2(n1161), .ZN(n20089) );
  NAND4_X2 U19558 ( .A1(n17756), .A2(n12758), .A3(n2619), .A4(n2618), .ZN(
        n30942) );
  NAND3_X2 U19565 ( .A1(n5581), .A2(n9597), .A3(n20407), .ZN(n8728) );
  AND2_X1 U19570 ( .A1(n30293), .A2(n29313), .Z(n7529) );
  NAND2_X1 U19592 ( .A1(n654), .A2(n23899), .ZN(n23628) );
  NOR2_X2 U19594 ( .A1(n31399), .A2(n30800), .ZN(n1260) );
  XOR2_X1 U19617 ( .A1(n30532), .A2(n17871), .Z(n13661) );
  XOR2_X1 U19623 ( .A1(n30807), .A2(n16002), .Z(n4574) );
  XOR2_X1 U19627 ( .A1(n30808), .A2(n25849), .Z(Ciphertext[176]) );
  NAND2_X2 U19631 ( .A1(n8628), .A2(n30810), .ZN(n16748) );
  AOI22_X1 U19632 ( .A1(n8627), .A2(n11123), .B1(n18541), .B2(n31821), .ZN(
        n30810) );
  NOR2_X2 U19646 ( .A1(n743), .A2(n11302), .ZN(n5034) );
  INV_X1 U19652 ( .I(n31180), .ZN(n5056) );
  AOI21_X1 U19655 ( .A1(n12486), .A2(n28658), .B(n31206), .ZN(n31214) );
  XOR2_X1 U19656 ( .A1(n8750), .A2(n29347), .Z(n30815) );
  AND2_X1 U19658 ( .A1(n25429), .A2(n17948), .Z(n31142) );
  NAND2_X1 U19667 ( .A1(n28353), .A2(n31563), .ZN(n14394) );
  XOR2_X1 U19676 ( .A1(n33509), .A2(n23239), .Z(n31191) );
  NOR2_X1 U19679 ( .A1(n28915), .A2(n8314), .ZN(n26660) );
  INV_X2 U19684 ( .I(n22602), .ZN(n8314) );
  XOR2_X1 U19688 ( .A1(n15727), .A2(n26487), .Z(n22602) );
  XOR2_X1 U19701 ( .A1(n2375), .A2(n30818), .Z(n31495) );
  XOR2_X1 U19702 ( .A1(n30819), .A2(n11889), .Z(n30818) );
  INV_X2 U19706 ( .I(n30820), .ZN(n23807) );
  XOR2_X1 U19707 ( .A1(n7616), .A2(n7614), .Z(n30820) );
  OAI22_X2 U19725 ( .A1(n14678), .A2(n18424), .B1(n17102), .B2(n14117), .ZN(
        n19158) );
  XOR2_X1 U19728 ( .A1(n30822), .A2(n15765), .Z(n3987) );
  AND2_X1 U19746 ( .A1(n7251), .A2(n4656), .Z(n2646) );
  XOR2_X1 U19751 ( .A1(n21036), .A2(n20842), .Z(n11578) );
  NOR2_X2 U19756 ( .A1(n12514), .A2(n20742), .ZN(n21036) );
  AOI21_X1 U19766 ( .A1(n19128), .A2(n7968), .B(n31177), .ZN(n12268) );
  NAND2_X2 U19772 ( .A1(n79), .A2(n31942), .ZN(n22831) );
  NOR2_X2 U19776 ( .A1(n27455), .A2(n11922), .ZN(n23646) );
  AND3_X1 U19788 ( .A1(n23730), .A2(n23938), .A3(n12469), .Z(n31028) );
  AOI21_X1 U19794 ( .A1(n30828), .A2(n27265), .B(n17181), .ZN(n17178) );
  NOR2_X1 U19816 ( .A1(n30326), .A2(n11394), .ZN(n21123) );
  XOR2_X1 U19823 ( .A1(n30830), .A2(n15307), .Z(n23683) );
  XOR2_X1 U19825 ( .A1(n23513), .A2(n23514), .Z(n30830) );
  INV_X4 U19828 ( .I(n7552), .ZN(n14005) );
  INV_X2 U19832 ( .I(n14851), .ZN(n22238) );
  NAND2_X2 U19833 ( .A1(n21765), .A2(n21764), .ZN(n14851) );
  XOR2_X1 U19848 ( .A1(n30837), .A2(n16655), .Z(Ciphertext[19]) );
  XOR2_X1 U19857 ( .A1(n30840), .A2(n25648), .Z(Ciphertext[140]) );
  AOI22_X1 U19860 ( .A1(n26745), .A2(n25646), .B1(n25660), .B2(n25645), .ZN(
        n30840) );
  XOR2_X1 U19870 ( .A1(n24645), .A2(n4244), .Z(n24482) );
  NAND2_X1 U19886 ( .A1(n24977), .A2(n17684), .ZN(n24892) );
  NOR2_X2 U19891 ( .A1(n15169), .A2(n15043), .ZN(n28504) );
  XOR2_X1 U19894 ( .A1(n7772), .A2(n30843), .Z(n9018) );
  BUF_X4 U19899 ( .I(n14396), .Z(n30885) );
  AND2_X1 U19900 ( .A1(n27748), .A2(n29688), .Z(n13083) );
  XOR2_X1 U19912 ( .A1(n30844), .A2(n7570), .Z(n14702) );
  XOR2_X1 U19917 ( .A1(n10169), .A2(n7569), .Z(n30844) );
  XOR2_X1 U19928 ( .A1(n33492), .A2(n24620), .Z(n24766) );
  XOR2_X1 U19932 ( .A1(n20692), .A2(n20769), .Z(n11304) );
  XOR2_X1 U19945 ( .A1(n30850), .A2(n5067), .Z(n1487) );
  XOR2_X1 U19949 ( .A1(n5100), .A2(n8997), .Z(n30850) );
  NAND2_X2 U19982 ( .A1(n27391), .A2(n6716), .ZN(n6713) );
  XOR2_X1 U19989 ( .A1(n15630), .A2(n5647), .Z(n4672) );
  NAND2_X2 U20005 ( .A1(n2997), .A2(n30855), .ZN(n3229) );
  NOR2_X2 U20006 ( .A1(n2996), .A2(n28519), .ZN(n30855) );
  OAI21_X2 U20014 ( .A1(n13083), .A2(n33714), .B(n13157), .ZN(n30857) );
  XOR2_X1 U20038 ( .A1(n10539), .A2(n24846), .Z(n24597) );
  OAI21_X2 U20039 ( .A1(n2851), .A2(n2849), .B(n2848), .ZN(n24846) );
  XOR2_X1 U20065 ( .A1(n9526), .A2(n19491), .Z(n3980) );
  NAND2_X1 U20066 ( .A1(n12270), .A2(n18983), .ZN(n31177) );
  INV_X2 U20074 ( .I(n30861), .ZN(n17522) );
  OAI21_X1 U20075 ( .A1(n30863), .A2(n30862), .B(n21368), .ZN(n26504) );
  NOR2_X1 U20087 ( .A1(n21367), .A2(n21391), .ZN(n30862) );
  NAND2_X2 U20090 ( .A1(n30957), .A2(n30959), .ZN(n19245) );
  NAND3_X1 U20091 ( .A1(n25121), .A2(n2092), .A3(n25120), .ZN(n13667) );
  AOI22_X1 U20093 ( .A1(n11518), .A2(n2209), .B1(n2208), .B2(n25670), .ZN(
        n6469) );
  NAND2_X1 U20095 ( .A1(n146), .A2(n9195), .ZN(n30867) );
  NAND2_X1 U20097 ( .A1(n30933), .A2(n30932), .ZN(n31150) );
  NOR2_X2 U20112 ( .A1(n30869), .A2(n29603), .ZN(n15591) );
  NOR2_X2 U20113 ( .A1(n9560), .A2(n6958), .ZN(n31136) );
  NAND2_X2 U20117 ( .A1(n8015), .A2(n8016), .ZN(n2387) );
  XOR2_X1 U20120 ( .A1(n23471), .A2(n23356), .Z(n15712) );
  XOR2_X1 U20124 ( .A1(n6886), .A2(n30871), .Z(n16277) );
  XOR2_X1 U20125 ( .A1(n16912), .A2(n16910), .Z(n30871) );
  XOR2_X1 U20126 ( .A1(n1261), .A2(n12491), .Z(n9222) );
  NAND2_X1 U20133 ( .A1(n30872), .A2(n16699), .ZN(n8437) );
  NAND2_X1 U20137 ( .A1(n19335), .A2(n2207), .ZN(n30872) );
  OR2_X1 U20146 ( .A1(n31532), .A2(n20471), .Z(n30873) );
  NAND3_X2 U20154 ( .A1(n5222), .A2(n5221), .A3(n12755), .ZN(n19627) );
  INV_X2 U20158 ( .I(n13530), .ZN(n24209) );
  XOR2_X1 U20162 ( .A1(n15825), .A2(n22226), .Z(n12495) );
  XNOR2_X1 U20174 ( .A1(n10539), .A2(n24760), .ZN(n24576) );
  NOR2_X1 U20181 ( .A1(n10542), .A2(n30980), .ZN(n30979) );
  NAND2_X1 U20183 ( .A1(n29367), .A2(n30979), .ZN(n3840) );
  NAND2_X1 U20184 ( .A1(n20602), .A2(n15230), .ZN(n20601) );
  OAI22_X2 U20187 ( .A1(n21839), .A2(n21840), .B1(n13816), .B2(n21844), .ZN(
        n14594) );
  XOR2_X1 U20192 ( .A1(n14969), .A2(n22300), .Z(n22008) );
  XOR2_X1 U20201 ( .A1(n20799), .A2(n30880), .Z(n31841) );
  XOR2_X1 U20203 ( .A1(n20921), .A2(n30881), .Z(n30880) );
  XOR2_X1 U20204 ( .A1(n31043), .A2(n21018), .Z(n2304) );
  NAND2_X2 U20211 ( .A1(n27646), .A2(n5103), .ZN(n31043) );
  NAND2_X2 U20222 ( .A1(n31967), .A2(n28840), .ZN(n11103) );
  INV_X2 U20228 ( .I(n2347), .ZN(n5379) );
  XOR2_X1 U20230 ( .A1(n29057), .A2(n616), .Z(n2347) );
  XOR2_X1 U20261 ( .A1(n17546), .A2(n30887), .Z(n31875) );
  XOR2_X1 U20262 ( .A1(n5211), .A2(n27613), .Z(n30887) );
  AOI21_X2 U20269 ( .A1(n10468), .A2(n30889), .B(n32816), .ZN(n9071) );
  NAND2_X2 U20278 ( .A1(n327), .A2(n16334), .ZN(n6649) );
  INV_X1 U20280 ( .I(n1694), .ZN(n19771) );
  OR2_X1 U20294 ( .A1(n26040), .A2(n3601), .Z(n13087) );
  OR2_X1 U20298 ( .A1(n20322), .A2(n20379), .Z(n30892) );
  OR2_X1 U20311 ( .A1(n20008), .A2(n20080), .Z(n13771) );
  NAND2_X2 U20312 ( .A1(n17183), .A2(n30898), .ZN(n1931) );
  XOR2_X1 U20318 ( .A1(n19662), .A2(n13099), .Z(n30899) );
  XOR2_X1 U20321 ( .A1(n30900), .A2(n13689), .Z(n14621) );
  XOR2_X1 U20323 ( .A1(n26794), .A2(n30993), .Z(n30900) );
  XOR2_X1 U20325 ( .A1(n22016), .A2(n4739), .Z(n30901) );
  AOI21_X2 U20334 ( .A1(n867), .A2(n10488), .B(n31135), .ZN(n10486) );
  XOR2_X1 U20339 ( .A1(n2117), .A2(n25783), .Z(n4567) );
  NAND2_X2 U20340 ( .A1(n31297), .A2(n31872), .ZN(n2117) );
  XOR2_X1 U20363 ( .A1(n30749), .A2(n16690), .Z(n26929) );
  INV_X2 U20365 ( .I(n30905), .ZN(n20092) );
  BUF_X2 U20368 ( .I(n8392), .Z(n30906) );
  XOR2_X1 U20378 ( .A1(n13132), .A2(n13131), .Z(n15401) );
  OAI21_X2 U20399 ( .A1(n30914), .A2(n30913), .B(n728), .ZN(n28821) );
  INV_X2 U20405 ( .I(n21433), .ZN(n30914) );
  NOR2_X1 U20406 ( .A1(n31207), .A2(n25072), .ZN(n5864) );
  NAND2_X1 U20407 ( .A1(n33288), .A2(n5003), .ZN(n30915) );
  NAND2_X1 U20412 ( .A1(n11195), .A2(n858), .ZN(n30989) );
  OR2_X1 U20423 ( .A1(n25072), .A2(n32900), .Z(n28655) );
  AOI21_X2 U20437 ( .A1(n29394), .A2(n30727), .B(n2941), .ZN(n10769) );
  NAND3_X2 U20440 ( .A1(n30919), .A2(n27618), .A3(n3149), .ZN(n3093) );
  NAND2_X2 U20454 ( .A1(n25966), .A2(n11988), .ZN(n13353) );
  NAND3_X1 U20464 ( .A1(n28734), .A2(n25312), .A3(n25322), .ZN(n17105) );
  NAND2_X2 U20481 ( .A1(n23679), .A2(n23680), .ZN(n24652) );
  XOR2_X1 U20482 ( .A1(n3322), .A2(n3319), .Z(n3318) );
  XOR2_X1 U20483 ( .A1(n27176), .A2(n23295), .Z(n3322) );
  NOR2_X2 U20485 ( .A1(n2272), .A2(n31215), .ZN(n30978) );
  NAND2_X2 U20490 ( .A1(n10769), .A2(n2719), .ZN(n21816) );
  INV_X2 U20508 ( .I(n30926), .ZN(n22425) );
  XOR2_X1 U20509 ( .A1(n16000), .A2(n15999), .Z(n30926) );
  XNOR2_X1 U20521 ( .A1(n12442), .A2(n29030), .ZN(n19584) );
  AOI22_X2 U20529 ( .A1(n23962), .A2(n28410), .B1(n24046), .B2(n3506), .ZN(
        n3508) );
  NAND2_X2 U20538 ( .A1(n25442), .A2(n25439), .ZN(n25437) );
  OAI21_X2 U20563 ( .A1(n739), .A2(n23887), .B(n23841), .ZN(n8689) );
  NOR2_X2 U20575 ( .A1(n11742), .A2(n13732), .ZN(n16141) );
  NAND2_X2 U20587 ( .A1(n21532), .A2(n30389), .ZN(n17274) );
  XOR2_X1 U20592 ( .A1(n21951), .A2(n16036), .Z(n13436) );
  OR2_X1 U20606 ( .A1(n12974), .A2(n23843), .Z(n7524) );
  XOR2_X1 U20612 ( .A1(n30380), .A2(n23233), .Z(n23384) );
  NAND2_X2 U20619 ( .A1(n11162), .A2(n23089), .ZN(n23233) );
  NAND2_X2 U20629 ( .A1(n27793), .A2(n23550), .ZN(n24403) );
  NAND3_X1 U20631 ( .A1(n24325), .A2(n24327), .A3(n29141), .ZN(n24080) );
  AOI21_X2 U20650 ( .A1(n30948), .A2(n25121), .B(n25025), .ZN(n16469) );
  AOI22_X2 U20660 ( .A1(n15902), .A2(n8184), .B1(n16538), .B2(n18407), .ZN(
        n27953) );
  OAI21_X2 U20661 ( .A1(n13839), .A2(n22967), .B(n13837), .ZN(n23475) );
  NOR2_X2 U20667 ( .A1(n9959), .A2(n10258), .ZN(n9958) );
  XOR2_X1 U20670 ( .A1(n26054), .A2(n22268), .Z(n30951) );
  OR2_X1 U20690 ( .A1(n16226), .A2(n20657), .Z(n20662) );
  NAND2_X2 U20691 ( .A1(n5448), .A2(n22806), .ZN(n26724) );
  AOI22_X2 U20697 ( .A1(n4931), .A2(n4932), .B1(n4930), .B2(n33904), .ZN(
        n30953) );
  XOR2_X1 U20699 ( .A1(n20955), .A2(n30954), .Z(n587) );
  NAND2_X2 U20703 ( .A1(n13276), .A2(n13275), .ZN(n7229) );
  XOR2_X1 U20707 ( .A1(n17400), .A2(n30955), .Z(n28818) );
  NOR2_X2 U20720 ( .A1(n31949), .A2(n30958), .ZN(n30957) );
  INV_X2 U20722 ( .I(n18876), .ZN(n30959) );
  OR2_X2 U20724 ( .A1(n15721), .A2(n7865), .Z(n4602) );
  XOR2_X1 U20746 ( .A1(n12936), .A2(n12935), .Z(n24360) );
  XOR2_X1 U20750 ( .A1(n30964), .A2(n23188), .Z(n10772) );
  XOR2_X1 U20774 ( .A1(n24841), .A2(n26121), .Z(n29072) );
  XOR2_X1 U20782 ( .A1(n11651), .A2(n1084), .Z(n24841) );
  OAI21_X1 U20783 ( .A1(n30971), .A2(n20635), .B(n30970), .ZN(n1811) );
  NAND2_X1 U20785 ( .A1(n15569), .A2(n3994), .ZN(n7786) );
  OR2_X1 U20786 ( .A1(n28702), .A2(n30973), .Z(n5836) );
  INV_X2 U20814 ( .I(n843), .ZN(n30980) );
  XOR2_X1 U20815 ( .A1(n30981), .A2(n29467), .Z(n31140) );
  XOR2_X1 U20827 ( .A1(n16992), .A2(n13702), .Z(n30981) );
  NOR2_X2 U20831 ( .A1(n27555), .A2(n10030), .ZN(n30982) );
  XOR2_X1 U20832 ( .A1(n30985), .A2(n20719), .Z(n26401) );
  XOR2_X1 U20851 ( .A1(n5296), .A2(n6050), .Z(n30986) );
  NOR2_X1 U20860 ( .A1(n18098), .A2(n22394), .ZN(n31144) );
  XOR2_X1 U20861 ( .A1(n20757), .A2(n5210), .Z(n5209) );
  XOR2_X1 U20870 ( .A1(n23282), .A2(n32899), .Z(n15432) );
  NAND2_X2 U20871 ( .A1(n16630), .A2(n16789), .ZN(n10413) );
  XOR2_X1 U20877 ( .A1(n2192), .A2(n30992), .Z(n509) );
  XOR2_X1 U20887 ( .A1(n31477), .A2(n30993), .Z(n30992) );
  INV_X2 U20895 ( .I(n30994), .ZN(n9170) );
  NAND2_X2 U20906 ( .A1(n29525), .A2(n13925), .ZN(n18922) );
  XOR2_X1 U20932 ( .A1(n1781), .A2(n1778), .Z(n17683) );
  BUF_X2 U20940 ( .I(n22634), .Z(n31001) );
  XOR2_X1 U20941 ( .A1(n7646), .A2(n7644), .Z(n12804) );
  NAND2_X2 U20945 ( .A1(n29088), .A2(n424), .ZN(n9439) );
  NAND3_X1 U20948 ( .A1(n5494), .A2(n30832), .A3(n21872), .ZN(n12604) );
  AND2_X1 U20952 ( .A1(n22421), .A2(n22420), .Z(n31006) );
  AOI21_X1 U20967 ( .A1(n18822), .A2(n18701), .B(n31012), .ZN(n16395) );
  NAND2_X2 U20969 ( .A1(n23663), .A2(n31015), .ZN(n24632) );
  NOR2_X2 U20971 ( .A1(n16442), .A2(n10899), .ZN(n25893) );
  INV_X2 U20974 ( .I(n24096), .ZN(n17404) );
  OAI21_X2 U20979 ( .A1(n28303), .A2(n17490), .B(n23649), .ZN(n24096) );
  XOR2_X1 U20996 ( .A1(n4059), .A2(n6707), .Z(n6705) );
  INV_X4 U21004 ( .I(n26157), .ZN(n3748) );
  NOR2_X1 U21019 ( .A1(n19165), .A2(n4835), .ZN(n31029) );
  INV_X2 U21025 ( .I(n27933), .ZN(n468) );
  XOR2_X1 U21026 ( .A1(n19642), .A2(n19163), .Z(n6624) );
  AOI22_X2 U21032 ( .A1(n31781), .A2(n21846), .B1(n21518), .B2(n7969), .ZN(
        n31032) );
  XOR2_X1 U21033 ( .A1(n15433), .A2(n15430), .Z(n15514) );
  AND2_X1 U21041 ( .A1(n16686), .A2(n29268), .Z(n31524) );
  INV_X2 U21048 ( .I(n31034), .ZN(n9828) );
  XOR2_X1 U21049 ( .A1(n23516), .A2(n23254), .Z(n9865) );
  OAI21_X2 U21056 ( .A1(n12160), .A2(n2886), .B(n12159), .ZN(n31037) );
  NOR2_X2 U21063 ( .A1(n29397), .A2(n7105), .ZN(n31039) );
  OAI21_X1 U21065 ( .A1(n9285), .A2(n31042), .B(n31041), .ZN(n11646) );
  INV_X2 U21067 ( .I(n31044), .ZN(n20120) );
  XOR2_X1 U21069 ( .A1(n19640), .A2(n14574), .Z(n31044) );
  NOR2_X2 U21076 ( .A1(n18658), .A2(n18657), .ZN(n27807) );
  INV_X2 U21079 ( .I(n20011), .ZN(n31046) );
  AND2_X1 U21088 ( .A1(n5415), .A2(n819), .Z(n31047) );
  XOR2_X1 U21112 ( .A1(n7288), .A2(n34050), .Z(n27699) );
  OAI22_X2 U21114 ( .A1(n18344), .A2(n26181), .B1(n19052), .B2(n10015), .ZN(
        n18345) );
  XOR2_X1 U21147 ( .A1(n8113), .A2(n8110), .Z(n18080) );
  NAND2_X1 U21151 ( .A1(n17277), .A2(n13950), .ZN(n24107) );
  NAND2_X1 U21167 ( .A1(n25876), .A2(n25875), .ZN(n25877) );
  OAI22_X1 U21174 ( .A1(n22329), .A2(n1000), .B1(n22406), .B2(n30529), .ZN(
        n13071) );
  XOR2_X1 U21181 ( .A1(n5380), .A2(n31056), .Z(n31055) );
  NAND2_X2 U21187 ( .A1(n1146), .A2(n16639), .ZN(n21433) );
  OAI22_X2 U21195 ( .A1(n18841), .A2(n18840), .B1(n2148), .B2(n1181), .ZN(
        n31882) );
  NOR2_X1 U21198 ( .A1(n963), .A2(n14940), .ZN(n6043) );
  NOR2_X1 U21200 ( .A1(n18944), .A2(n7345), .ZN(n8573) );
  INV_X2 U21202 ( .I(n25313), .ZN(n1074) );
  NAND2_X2 U21217 ( .A1(n25293), .A2(n25294), .ZN(n25313) );
  AND2_X1 U21219 ( .A1(n22523), .A2(n22605), .Z(n29027) );
  XOR2_X1 U21223 ( .A1(n31059), .A2(n20835), .Z(n20895) );
  AOI21_X2 U21224 ( .A1(n5413), .A2(n5416), .B(n31976), .ZN(n5414) );
  XOR2_X1 U21236 ( .A1(n31731), .A2(n25457), .Z(n19693) );
  NAND2_X2 U21238 ( .A1(n16106), .A2(n19155), .ZN(n31731) );
  XNOR2_X1 U21246 ( .A1(n24646), .A2(n24231), .ZN(n31312) );
  NAND2_X2 U21254 ( .A1(n13985), .A2(n25302), .ZN(n31060) );
  NAND2_X2 U21260 ( .A1(n13768), .A2(n20556), .ZN(n20520) );
  XOR2_X1 U21263 ( .A1(n9135), .A2(n9136), .Z(n10197) );
  XOR2_X1 U21266 ( .A1(n8152), .A2(n24452), .Z(n28896) );
  XOR2_X1 U21267 ( .A1(n12283), .A2(n19737), .Z(n2750) );
  NAND2_X2 U21281 ( .A1(n21312), .A2(n21448), .ZN(n21314) );
  NOR2_X2 U21288 ( .A1(n17699), .A2(n16633), .ZN(n21312) );
  XOR2_X1 U21289 ( .A1(n18091), .A2(n31063), .Z(n10944) );
  XOR2_X1 U21290 ( .A1(n10084), .A2(n1423), .Z(n31063) );
  XOR2_X1 U21296 ( .A1(n31065), .A2(n25598), .Z(Ciphertext[132]) );
  NAND2_X2 U21297 ( .A1(n19031), .A2(n31066), .ZN(n7971) );
  XOR2_X1 U21305 ( .A1(n3235), .A2(n3233), .Z(n24503) );
  NAND2_X1 U21321 ( .A1(n26891), .A2(n27965), .ZN(n2970) );
  NAND2_X1 U21322 ( .A1(n23706), .A2(n499), .ZN(n15266) );
  XOR2_X1 U21326 ( .A1(n31070), .A2(n6086), .Z(n8074) );
  INV_X2 U21330 ( .I(n24091), .ZN(n10198) );
  NAND2_X2 U21338 ( .A1(n1035), .A2(n19990), .ZN(n13077) );
  XOR2_X1 U21339 ( .A1(n20850), .A2(n16823), .Z(n20853) );
  XOR2_X1 U21341 ( .A1(n20963), .A2(n20904), .Z(n20850) );
  NAND2_X2 U21359 ( .A1(n919), .A2(n21687), .ZN(n21686) );
  AOI22_X1 U21370 ( .A1(n6043), .A2(n25995), .B1(n30318), .B2(n3489), .ZN(
        n31075) );
  NAND2_X2 U21386 ( .A1(n31077), .A2(n9975), .ZN(n29157) );
  OAI21_X2 U21387 ( .A1(n28210), .A2(n14973), .B(n23784), .ZN(n31077) );
  NAND2_X1 U21400 ( .A1(n9485), .A2(n9483), .ZN(n31078) );
  XOR2_X1 U21410 ( .A1(n15438), .A2(n13793), .Z(n13792) );
  OAI21_X2 U21411 ( .A1(n24013), .A2(n10198), .B(n24130), .ZN(n7246) );
  XOR2_X1 U21420 ( .A1(n31151), .A2(n27812), .Z(n24883) );
  XOR2_X1 U21422 ( .A1(n11775), .A2(n14442), .Z(n31081) );
  XOR2_X1 U21434 ( .A1(n4792), .A2(n4790), .Z(n4791) );
  OAI22_X2 U21447 ( .A1(n31086), .A2(n24322), .B1(n7059), .B2(n24213), .ZN(
        n9468) );
  XOR2_X1 U21448 ( .A1(n20765), .A2(n20764), .Z(n3793) );
  XOR2_X1 U21452 ( .A1(n31087), .A2(n14202), .Z(n28750) );
  NAND2_X2 U21468 ( .A1(n31091), .A2(n16088), .ZN(n19046) );
  NAND2_X2 U21473 ( .A1(n27709), .A2(n16086), .ZN(n31091) );
  XOR2_X1 U21474 ( .A1(n24569), .A2(n5358), .Z(n31092) );
  INV_X1 U21476 ( .I(n23536), .ZN(n1258) );
  XOR2_X1 U21478 ( .A1(n20835), .A2(n17592), .Z(n20771) );
  XOR2_X1 U21490 ( .A1(n24662), .A2(n31093), .Z(n12083) );
  INV_X1 U21494 ( .I(n25549), .ZN(n31094) );
  NOR2_X2 U21502 ( .A1(n4017), .A2(n10017), .ZN(n19007) );
  BUF_X4 U21503 ( .I(n841), .Z(n31096) );
  NOR2_X1 U21507 ( .A1(n8946), .A2(n1826), .ZN(n31097) );
  XOR2_X1 U21510 ( .A1(n23384), .A2(n531), .Z(n12738) );
  XOR2_X1 U21511 ( .A1(n19463), .A2(n19445), .Z(n19642) );
  INV_X2 U21537 ( .I(n31099), .ZN(n18623) );
  AOI21_X1 U21544 ( .A1(n25306), .A2(n18059), .B(n692), .ZN(n5792) );
  XOR2_X1 U21567 ( .A1(n613), .A2(n10186), .Z(n31100) );
  NAND2_X2 U21570 ( .A1(n548), .A2(n32602), .ZN(n23866) );
  INV_X2 U21572 ( .I(n31101), .ZN(n515) );
  XOR2_X1 U21590 ( .A1(n31104), .A2(n4427), .Z(n31561) );
  XOR2_X1 U21594 ( .A1(n21995), .A2(n22275), .Z(n31104) );
  INV_X2 U21620 ( .I(n11248), .ZN(n397) );
  NOR2_X2 U21627 ( .A1(n31110), .A2(n31109), .ZN(n25743) );
  XOR2_X1 U21637 ( .A1(n19638), .A2(n19639), .Z(n14574) );
  XOR2_X1 U21644 ( .A1(n23286), .A2(n4047), .Z(n1795) );
  NAND2_X2 U21648 ( .A1(n13861), .A2(n17893), .ZN(n4047) );
  OAI21_X2 U21653 ( .A1(n3911), .A2(n18181), .B(n9737), .ZN(n28058) );
  NAND2_X2 U21658 ( .A1(n21799), .A2(n12211), .ZN(n21709) );
  XOR2_X1 U21660 ( .A1(n2747), .A2(n27365), .Z(n28430) );
  INV_X2 U21664 ( .I(n31114), .ZN(n31909) );
  XOR2_X1 U21668 ( .A1(n6895), .A2(n26087), .Z(n31114) );
  XOR2_X1 U21671 ( .A1(n1845), .A2(n1844), .Z(n31116) );
  XOR2_X1 U21672 ( .A1(n31117), .A2(n31756), .Z(n7672) );
  XOR2_X1 U21674 ( .A1(n20888), .A2(n5282), .Z(n31117) );
  NAND2_X1 U21676 ( .A1(n4714), .A2(n32619), .ZN(n4715) );
  NOR2_X1 U21686 ( .A1(n2720), .A2(n30129), .ZN(n2948) );
  NOR2_X2 U21687 ( .A1(n27406), .A2(n22479), .ZN(n31145) );
  NOR2_X2 U21707 ( .A1(n31118), .A2(n2178), .ZN(n22216) );
  INV_X1 U21726 ( .I(n23052), .ZN(n31120) );
  XOR2_X1 U21735 ( .A1(n26145), .A2(n3318), .Z(n31409) );
  XOR2_X1 U21752 ( .A1(n23530), .A2(n1428), .Z(n17353) );
  AOI21_X2 U21760 ( .A1(n11048), .A2(n10896), .B(n31758), .ZN(n23530) );
  XOR2_X1 U21772 ( .A1(n31123), .A2(n24820), .Z(n24821) );
  XOR2_X1 U21774 ( .A1(n27801), .A2(n24853), .Z(n31123) );
  OAI22_X1 U21787 ( .A1(n9655), .A2(n25194), .B1(n1071), .B2(n9247), .ZN(n4767) );
  INV_X2 U21788 ( .I(n4770), .ZN(n1071) );
  NAND2_X2 U21793 ( .A1(n13267), .A2(n11786), .ZN(n4770) );
  NAND2_X1 U21797 ( .A1(n10071), .A2(n11441), .ZN(n31124) );
  INV_X2 U21814 ( .I(n31128), .ZN(n15189) );
  NOR2_X2 U21823 ( .A1(n22870), .A2(n22869), .ZN(n23439) );
  XOR2_X1 U21844 ( .A1(n15543), .A2(n31132), .Z(n25325) );
  XOR2_X1 U21859 ( .A1(n14639), .A2(n25720), .Z(n31133) );
  OAI21_X2 U21864 ( .A1(n31784), .A2(n16501), .B(n22890), .ZN(n1563) );
  NAND3_X1 U21866 ( .A1(n24911), .A2(n10099), .A3(n24910), .ZN(n4898) );
  NOR3_X1 U21876 ( .A1(n1032), .A2(n20379), .A3(n18078), .ZN(n31135) );
  NAND2_X1 U21878 ( .A1(n31137), .A2(n29385), .ZN(n26696) );
  OAI21_X1 U21881 ( .A1(n17712), .A2(n16516), .B(n26547), .ZN(n31137) );
  NAND2_X2 U21883 ( .A1(n7281), .A2(n16009), .ZN(n20624) );
  BUF_X2 U21890 ( .I(n19779), .Z(n31138) );
  NAND3_X2 U21894 ( .A1(n7396), .A2(n7395), .A3(n7834), .ZN(n21037) );
  INV_X2 U21895 ( .I(n19002), .ZN(n743) );
  NAND2_X2 U21896 ( .A1(n6753), .A2(n9265), .ZN(n19002) );
  XOR2_X1 U21898 ( .A1(n27523), .A2(n26125), .Z(n28119) );
  INV_X2 U21899 ( .I(n31140), .ZN(n10955) );
  OAI21_X2 U21915 ( .A1(n31145), .A2(n22482), .B(n22480), .ZN(n22824) );
  NOR2_X2 U21931 ( .A1(n1353), .A2(n7280), .ZN(n7397) );
  NAND2_X1 U21933 ( .A1(n25877), .A2(n25709), .ZN(n31146) );
  INV_X2 U21939 ( .I(n31147), .ZN(n31579) );
  XNOR2_X1 U21942 ( .A1(Plaintext[57]), .A2(Key[57]), .ZN(n31147) );
  NAND2_X2 U21959 ( .A1(n11149), .A2(n11150), .ZN(n15091) );
  NOR2_X2 U21980 ( .A1(n6907), .A2(n9324), .ZN(n9994) );
  XOR2_X1 U21982 ( .A1(n24800), .A2(n26429), .Z(n31151) );
  NAND2_X2 U21983 ( .A1(n5119), .A2(n7995), .ZN(n8800) );
  XOR2_X1 U21984 ( .A1(n29728), .A2(n19769), .Z(n2628) );
  NOR2_X2 U21989 ( .A1(n3060), .A2(n3059), .ZN(n19769) );
  XOR2_X1 U22013 ( .A1(n8695), .A2(n27996), .Z(n23341) );
  NOR2_X2 U22016 ( .A1(n6676), .A2(n6677), .ZN(n8695) );
  OR3_X1 U22018 ( .A1(n11814), .A2(n14383), .A3(n3193), .Z(n31583) );
  AOI21_X2 U22019 ( .A1(n6108), .A2(n28423), .B(n31157), .ZN(n7292) );
  NOR2_X1 U22027 ( .A1(n18973), .A2(n15502), .ZN(n19227) );
  NAND2_X2 U22035 ( .A1(n26627), .A2(n16713), .ZN(n18973) );
  XOR2_X1 U22039 ( .A1(n16319), .A2(n7511), .Z(n24409) );
  NOR2_X2 U22043 ( .A1(n23992), .A2(n28725), .ZN(n16319) );
  BUF_X4 U22046 ( .I(n24789), .Z(n31687) );
  XOR2_X1 U22060 ( .A1(n31159), .A2(n14300), .Z(Ciphertext[0]) );
  AOI22_X1 U22062 ( .A1(n6155), .A2(n6154), .B1(n8980), .B2(n10755), .ZN(
        n31159) );
  OAI22_X2 U22071 ( .A1(n29448), .A2(n15869), .B1(n15759), .B2(n18975), .ZN(
        n19679) );
  XOR2_X1 U22072 ( .A1(n22319), .A2(n22320), .Z(n22324) );
  XOR2_X1 U22088 ( .A1(n31527), .A2(n1695), .Z(n13941) );
  INV_X2 U22089 ( .I(n5725), .ZN(n31161) );
  NAND2_X2 U22093 ( .A1(n3327), .A2(n31162), .ZN(n22990) );
  XOR2_X1 U22111 ( .A1(n3682), .A2(n22128), .Z(n10889) );
  OAI21_X2 U22112 ( .A1(n21487), .A2(n21488), .B(n3685), .ZN(n3682) );
  XOR2_X1 U22128 ( .A1(n23306), .A2(n27252), .Z(n2142) );
  XOR2_X1 U22133 ( .A1(n343), .A2(n16322), .Z(n22287) );
  XOR2_X1 U22135 ( .A1(n7477), .A2(n22205), .Z(n22313) );
  XOR2_X1 U22148 ( .A1(n31168), .A2(n18166), .Z(n20011) );
  XOR2_X1 U22153 ( .A1(n18165), .A2(n19700), .Z(n31168) );
  XOR2_X1 U22161 ( .A1(n19485), .A2(n31169), .Z(n19388) );
  XOR2_X1 U22176 ( .A1(n2611), .A2(n27144), .Z(n31169) );
  NAND2_X2 U22180 ( .A1(n11287), .A2(n11310), .ZN(n24158) );
  INV_X4 U22181 ( .I(n20375), .ZN(n20361) );
  XOR2_X1 U22194 ( .A1(n22259), .A2(n22261), .Z(n18121) );
  XOR2_X1 U22200 ( .A1(n22119), .A2(n22291), .Z(n22259) );
  INV_X2 U22202 ( .I(n16042), .ZN(n18539) );
  NAND2_X1 U22207 ( .A1(n14156), .A2(n16042), .ZN(n13787) );
  XOR2_X1 U22222 ( .A1(Plaintext[135]), .A2(Key[135]), .Z(n16042) );
  NAND3_X1 U22224 ( .A1(n15534), .A2(n28478), .A3(n33143), .ZN(n11778) );
  XOR2_X1 U22253 ( .A1(n19439), .A2(n15485), .Z(n14459) );
  XOR2_X1 U22257 ( .A1(n17554), .A2(n26530), .Z(n6789) );
  NAND2_X1 U22259 ( .A1(n18530), .A2(n18531), .ZN(n18534) );
  OR2_X1 U22277 ( .A1(n25316), .A2(n31178), .Z(n17058) );
  OAI21_X2 U22295 ( .A1(n22573), .A2(n1298), .B(n31181), .ZN(n10905) );
  OAI22_X2 U22296 ( .A1(n22524), .A2(n1728), .B1(n901), .B2(n17960), .ZN(
        n22605) );
  XOR2_X1 U22304 ( .A1(n31182), .A2(n16690), .Z(Ciphertext[30]) );
  AOI21_X1 U22308 ( .A1(n24250), .A2(n24251), .B(n28553), .ZN(n1513) );
  NAND2_X1 U22312 ( .A1(n32902), .A2(n21374), .ZN(n21377) );
  INV_X2 U22314 ( .I(n31184), .ZN(n24874) );
  XOR2_X1 U22319 ( .A1(n31186), .A2(n14754), .Z(n11327) );
  XOR2_X1 U22323 ( .A1(n22286), .A2(n11166), .Z(n31186) );
  INV_X2 U22329 ( .I(n20872), .ZN(n31189) );
  XOR2_X1 U22332 ( .A1(n6327), .A2(n31190), .Z(n6955) );
  XOR2_X1 U22333 ( .A1(n21960), .A2(n31191), .Z(n31190) );
  XOR2_X1 U22341 ( .A1(n3982), .A2(n31194), .Z(n14572) );
  XOR2_X1 U22343 ( .A1(n17540), .A2(n17541), .Z(n31194) );
  BUF_X2 U22347 ( .I(n8243), .Z(n31195) );
  AOI22_X1 U22351 ( .A1(n5638), .A2(n5043), .B1(n25223), .B2(n28358), .ZN(
        n5243) );
  AND2_X1 U22353 ( .A1(n16117), .A2(n1141), .Z(n4496) );
  XOR2_X1 U22367 ( .A1(n23341), .A2(n23340), .Z(n31200) );
  XOR2_X1 U22368 ( .A1(n17395), .A2(n31203), .Z(n2104) );
  NAND2_X2 U22371 ( .A1(n30744), .A2(n1430), .ZN(n18187) );
  NAND2_X2 U22373 ( .A1(n17900), .A2(n27067), .ZN(n16076) );
  XOR2_X1 U22382 ( .A1(n31205), .A2(n18898), .Z(n27599) );
  XOR2_X1 U22383 ( .A1(n19630), .A2(n4976), .Z(n31205) );
  INV_X2 U22386 ( .I(n17906), .ZN(n31208) );
  AOI22_X2 U22395 ( .A1(n27975), .A2(n26160), .B1(n5400), .B2(n1265), .ZN(
        n5399) );
  NAND2_X2 U22399 ( .A1(n22977), .A2(n1484), .ZN(n3600) );
  XOR2_X1 U22411 ( .A1(n20715), .A2(n20926), .Z(n20752) );
  NAND2_X2 U22418 ( .A1(n12504), .A2(n31213), .ZN(n12610) );
  XOR2_X1 U22435 ( .A1(n31214), .A2(n25065), .Z(Ciphertext[42]) );
  NAND3_X2 U22436 ( .A1(n22778), .A2(n22777), .A3(n22776), .ZN(n23335) );
  NAND2_X1 U22455 ( .A1(n24969), .A2(n3843), .ZN(n13736) );
  NAND2_X2 U22481 ( .A1(n10203), .A2(n19199), .ZN(n19033) );
  NAND2_X2 U22484 ( .A1(n22470), .A2(n4156), .ZN(n22885) );
  INV_X2 U22486 ( .I(n11438), .ZN(n24182) );
  AOI21_X1 U22494 ( .A1(n21286), .A2(n21285), .B(n21398), .ZN(n27198) );
  XOR2_X1 U22499 ( .A1(n14094), .A2(n19682), .Z(n8921) );
  XOR2_X1 U22504 ( .A1(n2261), .A2(n2554), .Z(n31221) );
  NAND2_X1 U22515 ( .A1(n21705), .A2(n21704), .ZN(n21145) );
  NAND3_X1 U22530 ( .A1(n24920), .A2(n15799), .A3(n15569), .ZN(n24353) );
  XOR2_X1 U22539 ( .A1(n29320), .A2(n24750), .Z(n5525) );
  XOR2_X1 U22541 ( .A1(n11562), .A2(n22189), .Z(n11781) );
  NAND2_X2 U22543 ( .A1(n12183), .A2(n16477), .ZN(n22189) );
  OAI21_X2 U22554 ( .A1(n7388), .A2(n21812), .B(n5474), .ZN(n11481) );
  XOR2_X1 U22563 ( .A1(n20979), .A2(n31235), .Z(n31234) );
  XOR2_X1 U22579 ( .A1(n6706), .A2(n31703), .Z(n31237) );
  XOR2_X1 U22580 ( .A1(n16861), .A2(n17259), .Z(n29101) );
  XOR2_X1 U22581 ( .A1(n24676), .A2(n15161), .Z(n15473) );
  NAND2_X2 U22584 ( .A1(n31238), .A2(n13021), .ZN(n20625) );
  OAI21_X2 U22595 ( .A1(n9855), .A2(n27343), .B(n19991), .ZN(n31238) );
  NAND2_X2 U22621 ( .A1(n31241), .A2(n13089), .ZN(n20820) );
  OAI21_X2 U22622 ( .A1(n10380), .A2(n19804), .B(n2565), .ZN(n31241) );
  NOR2_X2 U22625 ( .A1(n2149), .A2(n2584), .ZN(n18841) );
  NAND2_X1 U22630 ( .A1(n19984), .A2(n11508), .ZN(n31242) );
  XOR2_X1 U22632 ( .A1(n1690), .A2(n31243), .Z(n25345) );
  XOR2_X1 U22638 ( .A1(n24626), .A2(n29346), .Z(n31243) );
  XOR2_X1 U22642 ( .A1(n15941), .A2(n16076), .Z(n23505) );
  AOI21_X2 U22645 ( .A1(n7882), .A2(n29118), .B(n31246), .ZN(n8908) );
  NAND2_X2 U22651 ( .A1(n2448), .A2(n31247), .ZN(n9919) );
  INV_X2 U22652 ( .I(n31248), .ZN(n16966) );
  XOR2_X1 U22667 ( .A1(n4013), .A2(n1128), .Z(n31252) );
  XOR2_X1 U22673 ( .A1(n4013), .A2(n9960), .Z(n31253) );
  XOR2_X1 U22695 ( .A1(n21950), .A2(n16692), .Z(n22412) );
  XOR2_X1 U22702 ( .A1(n1886), .A2(n31258), .Z(n28260) );
  XOR2_X1 U22709 ( .A1(n11012), .A2(n20749), .Z(n31258) );
  XOR2_X1 U22710 ( .A1(n24598), .A2(n24523), .Z(n14918) );
  XOR2_X1 U22711 ( .A1(n7574), .A2(n31259), .Z(n24598) );
  INV_X2 U22714 ( .I(n24520), .ZN(n31259) );
  BUF_X2 U22718 ( .I(n21122), .Z(n31260) );
  OAI21_X2 U22730 ( .A1(n15154), .A2(n31262), .B(n12811), .ZN(n21704) );
  NAND3_X2 U22734 ( .A1(n21549), .A2(n21548), .A3(n21550), .ZN(n22067) );
  OAI21_X2 U22758 ( .A1(n17251), .A2(n15956), .B(n31265), .ZN(n31264) );
  NAND2_X2 U22768 ( .A1(n14831), .A2(n15956), .ZN(n31265) );
  OAI21_X1 U22778 ( .A1(n12033), .A2(n22801), .B(n26868), .ZN(n12597) );
  NAND2_X2 U22781 ( .A1(n20294), .A2(n20293), .ZN(n20556) );
  XOR2_X1 U22787 ( .A1(n12453), .A2(n19316), .Z(n31828) );
  XOR2_X1 U22788 ( .A1(n29030), .A2(n12048), .Z(n12453) );
  XOR2_X1 U22790 ( .A1(n20654), .A2(n28541), .Z(n17973) );
  BUF_X2 U22811 ( .I(n11947), .Z(n31268) );
  NAND2_X2 U22822 ( .A1(n25968), .A2(n19115), .ZN(n13330) );
  INV_X2 U22829 ( .I(n31272), .ZN(n13255) );
  OR2_X1 U22832 ( .A1(n22873), .A2(n22791), .Z(n22872) );
  OAI22_X2 U22835 ( .A1(n1664), .A2(n1663), .B1(n1661), .B2(n14253), .ZN(
        n22873) );
  NAND3_X1 U22866 ( .A1(n7924), .A2(n7926), .A3(n11571), .ZN(n31281) );
  NOR2_X2 U22870 ( .A1(n13482), .A2(n13481), .ZN(n13477) );
  NAND2_X2 U22894 ( .A1(n21550), .A2(n21494), .ZN(n31284) );
  INV_X2 U22906 ( .I(n25144), .ZN(n16751) );
  NAND2_X1 U22909 ( .A1(n25144), .A2(n25145), .ZN(n15330) );
  XOR2_X1 U22911 ( .A1(n16719), .A2(n6452), .Z(n25144) );
  NOR2_X2 U22913 ( .A1(n10495), .A2(n31285), .ZN(n10201) );
  AND2_X1 U22914 ( .A1(n6696), .A2(n22944), .Z(n31285) );
  OAI21_X2 U22917 ( .A1(n31286), .A2(n20540), .B(n26730), .ZN(n26165) );
  INV_X2 U22928 ( .I(n31287), .ZN(n634) );
  XNOR2_X1 U22930 ( .A1(n22019), .A2(n8352), .ZN(n31287) );
  OR2_X1 U22935 ( .A1(n19203), .A2(n19291), .Z(n31356) );
  NOR2_X2 U22936 ( .A1(n1052), .A2(n19300), .ZN(n19203) );
  XOR2_X1 U22946 ( .A1(n28983), .A2(n20792), .Z(n14647) );
  OAI21_X2 U22956 ( .A1(n1572), .A2(n33548), .B(n16538), .ZN(n18403) );
  NAND2_X2 U22957 ( .A1(n20625), .A2(n20623), .ZN(n7280) );
  NAND2_X2 U22959 ( .A1(n31292), .A2(n13397), .ZN(n6679) );
  OAI21_X2 U22963 ( .A1(n15477), .A2(n19935), .B(n5371), .ZN(n31292) );
  NAND2_X2 U22988 ( .A1(n23109), .A2(n853), .ZN(n23112) );
  XOR2_X1 U22993 ( .A1(n31296), .A2(n8687), .Z(n13272) );
  OR2_X1 U22997 ( .A1(n12535), .A2(n861), .Z(n21247) );
  NAND2_X1 U22999 ( .A1(n7785), .A2(n7786), .ZN(n31348) );
  XOR2_X1 U23004 ( .A1(n2785), .A2(n2788), .Z(n2784) );
  XOR2_X1 U23021 ( .A1(n26754), .A2(n18188), .Z(n679) );
  NOR2_X2 U23031 ( .A1(n10444), .A2(n502), .ZN(n9619) );
  XOR2_X1 U23041 ( .A1(n20975), .A2(n16958), .Z(n20887) );
  NAND2_X2 U23048 ( .A1(n20311), .A2(n12902), .ZN(n20975) );
  XOR2_X1 U23057 ( .A1(n11504), .A2(n32981), .Z(n14053) );
  NAND2_X2 U23058 ( .A1(n23049), .A2(n23048), .ZN(n11504) );
  XOR2_X1 U23061 ( .A1(n11816), .A2(n31301), .Z(n11833) );
  XOR2_X1 U23063 ( .A1(n15950), .A2(n22265), .Z(n31301) );
  NAND2_X2 U23067 ( .A1(n23009), .A2(n23011), .ZN(n6975) );
  AND2_X2 U23092 ( .A1(n9753), .A2(n9750), .Z(n22467) );
  XOR2_X1 U23097 ( .A1(n22167), .A2(n16767), .Z(n31303) );
  OR2_X1 U23098 ( .A1(n18879), .A2(n8213), .Z(n18441) );
  XNOR2_X1 U23106 ( .A1(n30329), .A2(n21994), .ZN(n21926) );
  NAND2_X2 U23112 ( .A1(n21796), .A2(n21795), .ZN(n21994) );
  NAND2_X2 U23114 ( .A1(n25738), .A2(n27189), .ZN(n4642) );
  OAI22_X2 U23131 ( .A1(n18047), .A2(n9460), .B1(n15717), .B2(n27090), .ZN(
        n12878) );
  OR2_X1 U23137 ( .A1(n31960), .A2(n6442), .Z(n26726) );
  OR2_X1 U23139 ( .A1(n11932), .A2(n32606), .Z(n16531) );
  OR2_X1 U23145 ( .A1(n32414), .A2(n19128), .Z(n31306) );
  NAND2_X2 U23148 ( .A1(n28660), .A2(n5573), .ZN(n28659) );
  XOR2_X1 U23159 ( .A1(n1604), .A2(n31308), .Z(n371) );
  INV_X1 U23161 ( .I(n25311), .ZN(n31308) );
  NAND2_X2 U23162 ( .A1(n1543), .A2(n1544), .ZN(n1604) );
  NAND2_X2 U23180 ( .A1(n27472), .A2(n15828), .ZN(n22226) );
  XOR2_X1 U23218 ( .A1(n24377), .A2(n31312), .Z(n6293) );
  NOR2_X2 U23223 ( .A1(n31798), .A2(n27752), .ZN(n11330) );
  XOR2_X1 U23225 ( .A1(n12980), .A2(n8992), .Z(n4251) );
  AOI21_X2 U23226 ( .A1(n21522), .A2(n21523), .B(n21744), .ZN(n21524) );
  INV_X4 U23235 ( .I(n31746), .ZN(n4747) );
  NAND2_X2 U23237 ( .A1(n3631), .A2(n3633), .ZN(n15508) );
  NAND2_X1 U23243 ( .A1(n23176), .A2(n28740), .ZN(n31314) );
  XOR2_X1 U23250 ( .A1(n31316), .A2(n17487), .Z(n22679) );
  XOR2_X1 U23253 ( .A1(n17486), .A2(n17485), .Z(n31316) );
  XOR2_X1 U23256 ( .A1(n32052), .A2(n21001), .Z(n13336) );
  INV_X1 U23264 ( .I(n18540), .ZN(n31821) );
  XOR2_X1 U23267 ( .A1(n6808), .A2(n20678), .Z(n7596) );
  XOR2_X1 U23275 ( .A1(n20776), .A2(n12721), .Z(n20678) );
  NOR2_X2 U23276 ( .A1(n12864), .A2(n13764), .ZN(n13811) );
  NAND2_X2 U23277 ( .A1(n13555), .A2(n15156), .ZN(n25546) );
  OR2_X1 U23278 ( .A1(n14236), .A2(n6489), .Z(n7476) );
  NAND2_X2 U23281 ( .A1(n13690), .A2(n28138), .ZN(n27996) );
  XNOR2_X1 U23285 ( .A1(n20680), .A2(n20679), .ZN(n31423) );
  OAI22_X2 U23288 ( .A1(n17897), .A2(n17896), .B1(n28357), .B2(n2609), .ZN(
        n20679) );
  INV_X2 U23289 ( .I(n6454), .ZN(n22017) );
  OAI22_X2 U23290 ( .A1(n28067), .A2(n28068), .B1(n4516), .B2(n28018), .ZN(
        n6454) );
  AND2_X1 U23299 ( .A1(n18540), .A2(n13363), .Z(n18302) );
  NAND3_X2 U23305 ( .A1(n4101), .A2(n24591), .A3(n25013), .ZN(n14964) );
  XOR2_X1 U23307 ( .A1(n3868), .A2(n23420), .Z(n23359) );
  INV_X2 U23316 ( .I(n31318), .ZN(n31920) );
  XOR2_X1 U23321 ( .A1(n2044), .A2(n2043), .Z(n31318) );
  NAND2_X1 U23322 ( .A1(n25022), .A2(n13427), .ZN(n2909) );
  NOR2_X2 U23326 ( .A1(n1549), .A2(n31320), .ZN(n25060) );
  XOR2_X1 U23327 ( .A1(n13927), .A2(n13928), .Z(n31321) );
  NOR2_X1 U23344 ( .A1(n15133), .A2(n15132), .ZN(n31323) );
  NAND2_X2 U23347 ( .A1(n13279), .A2(n490), .ZN(n12320) );
  NAND2_X1 U23359 ( .A1(n9284), .A2(n14917), .ZN(n12183) );
  OR2_X2 U23368 ( .A1(n26733), .A2(n14082), .Z(n20134) );
  NAND2_X1 U23369 ( .A1(n31811), .A2(n20460), .ZN(n20461) );
  INV_X2 U23371 ( .I(n17338), .ZN(n25999) );
  OAI21_X2 U23372 ( .A1(n17054), .A2(n18565), .B(n17135), .ZN(n17338) );
  NAND2_X2 U23391 ( .A1(n13546), .A2(n13547), .ZN(n17517) );
  NAND2_X1 U23411 ( .A1(n31932), .A2(n17879), .ZN(n31327) );
  XOR2_X1 U23418 ( .A1(n9574), .A2(n6458), .Z(n9436) );
  NAND2_X2 U23420 ( .A1(n13285), .A2(n19892), .ZN(n20228) );
  OAI21_X2 U23421 ( .A1(n8147), .A2(n8146), .B(n19891), .ZN(n13285) );
  XOR2_X1 U23441 ( .A1(n22172), .A2(n9129), .Z(n15950) );
  OAI22_X2 U23448 ( .A1(n28137), .A2(n21702), .B1(n11981), .B2(n32519), .ZN(
        n22172) );
  OAI21_X2 U23449 ( .A1(n31329), .A2(n11480), .B(n12925), .ZN(n7447) );
  XOR2_X1 U23464 ( .A1(n31330), .A2(n1742), .Z(n27819) );
  XOR2_X1 U23475 ( .A1(n31331), .A2(n31336), .Z(n31330) );
  INV_X1 U23488 ( .I(n15950), .ZN(n31336) );
  OAI21_X1 U23492 ( .A1(n17582), .A2(n17223), .B(n31339), .ZN(n14537) );
  XNOR2_X1 U23495 ( .A1(n17090), .A2(n19573), .ZN(n31387) );
  OAI21_X2 U23499 ( .A1(n10405), .A2(n28613), .B(n22876), .ZN(n28364) );
  XOR2_X1 U23508 ( .A1(n11636), .A2(n7889), .Z(n14518) );
  NOR2_X2 U23509 ( .A1(n28226), .A2(n11634), .ZN(n11636) );
  NAND2_X2 U23516 ( .A1(n31345), .A2(n31344), .ZN(n9399) );
  XOR2_X1 U23521 ( .A1(n31346), .A2(n9298), .Z(n10258) );
  XOR2_X1 U23528 ( .A1(n22271), .A2(n28575), .Z(n28574) );
  NAND3_X1 U23531 ( .A1(n16112), .A2(n12309), .A3(n25796), .ZN(n25791) );
  XOR2_X1 U23533 ( .A1(n7826), .A2(n31410), .Z(n31529) );
  OR2_X1 U23536 ( .A1(n26600), .A2(n19300), .Z(n31350) );
  BUF_X2 U23550 ( .I(n8695), .Z(n31354) );
  INV_X2 U23552 ( .I(n31357), .ZN(n7915) );
  XOR2_X1 U23560 ( .A1(n7916), .A2(n7917), .Z(n31357) );
  XOR2_X1 U23562 ( .A1(n13419), .A2(n24664), .Z(n24814) );
  AOI21_X2 U23566 ( .A1(n9367), .A2(n24061), .B(n9366), .ZN(n13419) );
  OAI21_X2 U23569 ( .A1(n27466), .A2(n21871), .B(n27596), .ZN(n31359) );
  NAND2_X1 U23571 ( .A1(n17255), .A2(n26249), .ZN(n17062) );
  OR2_X1 U23605 ( .A1(n15101), .A2(n12118), .Z(n31365) );
  NOR2_X1 U23607 ( .A1(n16453), .A2(n4016), .ZN(n31366) );
  INV_X2 U23608 ( .I(n9468), .ZN(n8491) );
  NAND2_X1 U23612 ( .A1(n4806), .A2(n22905), .ZN(n4805) );
  XOR2_X1 U23614 ( .A1(n4791), .A2(n31367), .Z(n23579) );
  XOR2_X1 U23619 ( .A1(n31588), .A2(n4794), .Z(n31367) );
  NAND2_X2 U23620 ( .A1(n21085), .A2(n21170), .ZN(n21354) );
  OAI21_X2 U23624 ( .A1(n31369), .A2(n31368), .B(n16819), .ZN(n28073) );
  NOR2_X2 U23626 ( .A1(n4259), .A2(n12074), .ZN(n31368) );
  XOR2_X1 U23627 ( .A1(n31370), .A2(n25519), .Z(Ciphertext[119]) );
  NAND4_X2 U23637 ( .A1(n4325), .A2(n16468), .A3(n18215), .A4(n25518), .ZN(
        n31370) );
  XOR2_X1 U23640 ( .A1(n17517), .A2(n5772), .Z(n20897) );
  NAND2_X2 U23645 ( .A1(n26082), .A2(n26296), .ZN(n5772) );
  XOR2_X1 U23649 ( .A1(n31371), .A2(n10024), .Z(n10426) );
  XOR2_X1 U23651 ( .A1(n19723), .A2(n15990), .Z(n31371) );
  AND2_X1 U23652 ( .A1(n9959), .A2(n11833), .Z(n10310) );
  XOR2_X1 U23660 ( .A1(n1259), .A2(n27708), .Z(n8609) );
  NAND2_X2 U23667 ( .A1(n31547), .A2(n5058), .ZN(n27708) );
  XOR2_X1 U23670 ( .A1(n20963), .A2(n20820), .Z(n20888) );
  NAND2_X2 U23672 ( .A1(n3835), .A2(n31372), .ZN(n4450) );
  XOR2_X1 U23676 ( .A1(n24528), .A2(n24529), .Z(n16125) );
  INV_X2 U23677 ( .I(n24440), .ZN(n31373) );
  BUF_X2 U23680 ( .I(n6500), .Z(n31374) );
  NOR2_X1 U23683 ( .A1(n16819), .A2(n31579), .ZN(n18608) );
  XOR2_X1 U23686 ( .A1(n17128), .A2(n17395), .Z(n27135) );
  XOR2_X1 U23689 ( .A1(n32537), .A2(n22192), .Z(n12882) );
  XOR2_X1 U23691 ( .A1(n6948), .A2(n29428), .Z(n6093) );
  NOR2_X1 U23702 ( .A1(n26445), .A2(n29302), .ZN(n31379) );
  INV_X1 U23721 ( .I(n31532), .ZN(n20476) );
  XOR2_X1 U23723 ( .A1(n31380), .A2(n21930), .Z(n9533) );
  NAND2_X1 U23728 ( .A1(n9180), .A2(n25819), .ZN(n31381) );
  NAND2_X2 U23737 ( .A1(n3792), .A2(n29364), .ZN(n13267) );
  AOI22_X2 U23752 ( .A1(n31385), .A2(n12394), .B1(n5383), .B2(n4689), .ZN(
        n22123) );
  NAND2_X1 U23761 ( .A1(n26283), .A2(n12354), .ZN(n31385) );
  XOR2_X1 U23767 ( .A1(n13780), .A2(n31387), .Z(n245) );
  NOR2_X1 U23782 ( .A1(n20329), .A2(n31390), .ZN(n31389) );
  NAND3_X1 U23786 ( .A1(n15304), .A2(n12308), .A3(n12309), .ZN(n28989) );
  INV_X2 U23789 ( .I(n5016), .ZN(n31458) );
  INV_X2 U23790 ( .I(n9285), .ZN(n14384) );
  XOR2_X1 U23792 ( .A1(n17014), .A2(n17012), .Z(n17015) );
  NAND2_X1 U23800 ( .A1(n10419), .A2(n31393), .ZN(n27738) );
  XOR2_X1 U23811 ( .A1(n31395), .A2(n7866), .Z(n7865) );
  NOR2_X2 U23816 ( .A1(n31397), .A2(n78), .ZN(n1471) );
  NOR2_X1 U23820 ( .A1(n4935), .A2(n23110), .ZN(n31397) );
  NOR2_X2 U23829 ( .A1(n8425), .A2(n31398), .ZN(n20425) );
  INV_X1 U23850 ( .I(n1260), .ZN(n6905) );
  AOI21_X2 U23869 ( .A1(n31400), .A2(n12140), .B(n32397), .ZN(n28439) );
  XOR2_X1 U23871 ( .A1(n9353), .A2(n5268), .Z(n12422) );
  BUF_X2 U23892 ( .I(n13622), .Z(n31402) );
  NAND2_X1 U23908 ( .A1(n26637), .A2(n12265), .ZN(n12264) );
  XOR2_X1 U23932 ( .A1(n12212), .A2(n19729), .Z(n4631) );
  NAND2_X2 U23934 ( .A1(n8717), .A2(n8716), .ZN(n12212) );
  XOR2_X1 U23935 ( .A1(n18042), .A2(n24379), .Z(n31405) );
  NAND2_X2 U23940 ( .A1(n10854), .A2(n31406), .ZN(n19597) );
  NAND3_X1 U23942 ( .A1(n25671), .A2(n25673), .A3(n25672), .ZN(n31478) );
  XOR2_X1 U23946 ( .A1(n16893), .A2(n14851), .Z(n16896) );
  NOR2_X2 U23947 ( .A1(n27753), .A2(n27754), .ZN(n16893) );
  INV_X2 U23952 ( .I(n31409), .ZN(n17133) );
  NAND2_X1 U23957 ( .A1(n1387), .A2(n18994), .ZN(n18943) );
  XOR2_X1 U23971 ( .A1(n22033), .A2(n25801), .Z(n22034) );
  NAND2_X2 U23977 ( .A1(n16888), .A2(n16889), .ZN(n22033) );
  AND2_X1 U23981 ( .A1(n13921), .A2(n5480), .Z(n11457) );
  XOR2_X1 U24000 ( .A1(n19345), .A2(n5526), .Z(n17575) );
  INV_X2 U24006 ( .I(n20371), .ZN(n20533) );
  XOR2_X1 U24010 ( .A1(n20853), .A2(n17957), .Z(n21220) );
  AOI21_X1 U24019 ( .A1(n2858), .A2(n5962), .B(n4459), .ZN(n3810) );
  NAND2_X2 U24036 ( .A1(n18928), .A2(n18927), .ZN(n31415) );
  NOR2_X1 U24056 ( .A1(n11596), .A2(n21876), .ZN(n14822) );
  NAND2_X1 U24063 ( .A1(n31922), .A2(n20133), .ZN(n19806) );
  NOR2_X1 U24073 ( .A1(n7802), .A2(n14129), .ZN(n13838) );
  NAND2_X2 U24087 ( .A1(n13878), .A2(n28850), .ZN(n24204) );
  NAND2_X2 U24088 ( .A1(n10848), .A2(n32953), .ZN(n31422) );
  XOR2_X1 U24097 ( .A1(n31423), .A2(n20678), .Z(n18025) );
  NAND3_X2 U24109 ( .A1(n4717), .A2(n5561), .A3(n5560), .ZN(n9319) );
  NOR3_X1 U24116 ( .A1(n18884), .A2(n18660), .A3(n18888), .ZN(n10537) );
  OAI21_X2 U24126 ( .A1(n29379), .A2(n31424), .B(n10381), .ZN(n13205) );
  XOR2_X1 U24145 ( .A1(n31426), .A2(n24795), .Z(n12637) );
  XOR2_X1 U24147 ( .A1(n10870), .A2(n4997), .Z(n31426) );
  NAND2_X2 U24150 ( .A1(n6362), .A2(n28943), .ZN(n19265) );
  XOR2_X1 U24151 ( .A1(n20899), .A2(n15275), .Z(n21041) );
  XOR2_X1 U24155 ( .A1(n23284), .A2(n31429), .Z(n10525) );
  NAND2_X2 U24159 ( .A1(n31689), .A2(n1668), .ZN(n14392) );
  XOR2_X1 U24207 ( .A1(n31432), .A2(n16551), .Z(Ciphertext[190]) );
  NAND4_X2 U24213 ( .A1(n25920), .A2(n25919), .A3(n25918), .A4(n25917), .ZN(
        n31432) );
  XOR2_X1 U24218 ( .A1(n28633), .A2(n22224), .Z(n8275) );
  NOR2_X2 U24240 ( .A1(n24265), .A2(n31096), .ZN(n24230) );
  NAND2_X2 U24253 ( .A1(n21405), .A2(n32069), .ZN(n15807) );
  NOR2_X2 U24279 ( .A1(n26220), .A2(n27329), .ZN(n24141) );
  XOR2_X1 U24290 ( .A1(n19550), .A2(n19661), .Z(n19739) );
  NAND2_X2 U24293 ( .A1(n3072), .A2(n6576), .ZN(n19550) );
  XOR2_X1 U24313 ( .A1(n14689), .A2(n1230), .Z(n31440) );
  INV_X2 U24314 ( .I(n8327), .ZN(n26733) );
  INV_X1 U24317 ( .I(n31564), .ZN(n22915) );
  XOR2_X1 U24338 ( .A1(n11868), .A2(n24442), .Z(n14362) );
  INV_X2 U24348 ( .I(n31445), .ZN(n29253) );
  XOR2_X1 U24349 ( .A1(n8772), .A2(n8771), .Z(n31445) );
  NAND2_X1 U24386 ( .A1(n26284), .A2(n17626), .ZN(n16411) );
  NAND3_X1 U24389 ( .A1(n547), .A2(n24466), .A3(n12358), .ZN(n3828) );
  BUF_X2 U24398 ( .I(n19629), .Z(n31450) );
  XOR2_X1 U24400 ( .A1(n24416), .A2(n7837), .Z(n5146) );
  NAND3_X2 U24410 ( .A1(n20406), .A2(n32061), .A3(n10849), .ZN(n9597) );
  NAND2_X2 U24421 ( .A1(n1913), .A2(n1910), .ZN(n21655) );
  OAI22_X2 U24451 ( .A1(n13262), .A2(n6392), .B1(n13261), .B2(n12658), .ZN(
        n24180) );
  INV_X2 U24463 ( .I(n26785), .ZN(n31457) );
  NAND2_X2 U24465 ( .A1(n21472), .A2(n21471), .ZN(n26785) );
  OAI21_X2 U24476 ( .A1(n4585), .A2(n10849), .B(n4586), .ZN(n7954) );
  AND2_X1 U24481 ( .A1(n564), .A2(n13510), .Z(n12179) );
  NOR2_X1 U24485 ( .A1(n2958), .A2(n31504), .ZN(n15953) );
  NAND2_X1 U24499 ( .A1(n28435), .A2(n31458), .ZN(n8584) );
  OAI22_X1 U24526 ( .A1(n23729), .A2(n23939), .B1(n23730), .B2(n23731), .ZN(
        n26220) );
  INV_X4 U24544 ( .I(n32040), .ZN(n21811) );
  NAND3_X1 U24548 ( .A1(n29351), .A2(n15084), .A3(n17787), .ZN(n12004) );
  XOR2_X1 U24550 ( .A1(n1344), .A2(n1923), .Z(n5067) );
  INV_X2 U24552 ( .I(n31467), .ZN(n31914) );
  NAND2_X2 U24555 ( .A1(n28350), .A2(n9214), .ZN(n3205) );
  OAI21_X1 U24559 ( .A1(n4415), .A2(n25736), .B(n25739), .ZN(n7038) );
  NAND2_X2 U24561 ( .A1(n1601), .A2(n1600), .ZN(n4415) );
  XOR2_X1 U24584 ( .A1(n30304), .A2(n20872), .Z(n26647) );
  INV_X2 U24587 ( .I(n15299), .ZN(n15301) );
  OAI22_X2 U24589 ( .A1(n15450), .A2(n13966), .B1(n15449), .B2(n15448), .ZN(
        n15299) );
  NOR2_X2 U24591 ( .A1(n31473), .A2(n28882), .ZN(n7312) );
  NAND2_X1 U24596 ( .A1(n21270), .A2(n11814), .ZN(n31474) );
  XOR2_X1 U24600 ( .A1(n24116), .A2(n17912), .Z(n24574) );
  AOI21_X1 U24603 ( .A1(n23940), .A2(n11933), .B(n757), .ZN(n98) );
  OAI21_X1 U24607 ( .A1(n16425), .A2(n24064), .B(n25570), .ZN(n27354) );
  NOR2_X2 U24608 ( .A1(n28488), .A2(n10428), .ZN(n16425) );
  XOR2_X1 U24610 ( .A1(n31478), .A2(n16687), .Z(Ciphertext[145]) );
  NAND2_X2 U24618 ( .A1(n5886), .A2(n12264), .ZN(n12611) );
  NAND2_X2 U24624 ( .A1(n21180), .A2(n21179), .ZN(n26439) );
  NOR2_X1 U24633 ( .A1(n24729), .A2(n4490), .ZN(n4492) );
  INV_X1 U24635 ( .I(n25762), .ZN(n24729) );
  NAND3_X2 U24636 ( .A1(n4713), .A2(n4710), .A3(n4711), .ZN(n23292) );
  NOR2_X1 U24637 ( .A1(n563), .A2(n9469), .ZN(n7014) );
  NOR2_X1 U24646 ( .A1(n18711), .A2(n11707), .ZN(n18506) );
  NAND3_X1 U24677 ( .A1(n6595), .A2(n17637), .A3(n33400), .ZN(n25518) );
  NAND2_X2 U24678 ( .A1(n13246), .A2(n13247), .ZN(n19866) );
  XOR2_X1 U24697 ( .A1(n210), .A2(n22231), .Z(n31486) );
  NAND2_X2 U24704 ( .A1(n31487), .A2(n13003), .ZN(n15613) );
  OAI21_X2 U24711 ( .A1(n13006), .A2(n22861), .B(n22895), .ZN(n31487) );
  NAND2_X1 U24713 ( .A1(n23943), .A2(n3375), .ZN(n27078) );
  NOR2_X2 U24739 ( .A1(n32076), .A2(n21700), .ZN(n28137) );
  XOR2_X1 U24744 ( .A1(n31488), .A2(n32796), .Z(Ciphertext[129]) );
  NOR2_X1 U24747 ( .A1(n31489), .A2(n6114), .ZN(n31488) );
  NAND2_X1 U24750 ( .A1(n25696), .A2(n25695), .ZN(n31490) );
  NOR2_X2 U24765 ( .A1(n28278), .A2(n5170), .ZN(n27704) );
  XOR2_X1 U24780 ( .A1(n128), .A2(n19555), .Z(n17559) );
  XNOR2_X1 U24783 ( .A1(n9189), .A2(n28188), .ZN(n31552) );
  XOR2_X1 U24787 ( .A1(n20754), .A2(n13041), .Z(n20889) );
  NAND2_X2 U24794 ( .A1(n20399), .A2(n26216), .ZN(n20754) );
  AND2_X1 U24824 ( .A1(n12932), .A2(n14770), .Z(n7767) );
  XOR2_X1 U24826 ( .A1(n23296), .A2(n23206), .Z(n8810) );
  AOI21_X2 U24834 ( .A1(n18124), .A2(n17360), .B(n31500), .ZN(n19300) );
  OAI22_X2 U24835 ( .A1(n17599), .A2(n18863), .B1(n15583), .B2(n17360), .ZN(
        n31500) );
  NAND2_X2 U24850 ( .A1(n13852), .A2(n16694), .ZN(n19862) );
  NOR2_X1 U24856 ( .A1(n11173), .A2(n14055), .ZN(n5662) );
  NAND3_X1 U24860 ( .A1(n5774), .A2(n5773), .A3(n24919), .ZN(n439) );
  AOI21_X2 U24864 ( .A1(n10808), .A2(n29963), .B(n31503), .ZN(n18321) );
  NOR2_X2 U24870 ( .A1(n10315), .A2(n11146), .ZN(n31505) );
  NAND2_X2 U24888 ( .A1(n31675), .A2(n17443), .ZN(n9403) );
  OAI21_X2 U24896 ( .A1(n22881), .A2(n33395), .B(n17463), .ZN(n23534) );
  XNOR2_X1 U24910 ( .A1(n19395), .A2(n17369), .ZN(n19709) );
  NAND2_X2 U24933 ( .A1(n13937), .A2(n13939), .ZN(n19395) );
  OAI21_X1 U24937 ( .A1(n406), .A2(n405), .B(n25863), .ZN(n27217) );
  NAND2_X2 U24941 ( .A1(n26778), .A2(n16641), .ZN(n4335) );
  XOR2_X1 U24953 ( .A1(n31509), .A2(n24828), .Z(n1851) );
  XOR2_X1 U24957 ( .A1(n11612), .A2(n11610), .Z(n8042) );
  INV_X4 U24977 ( .I(n22977), .ZN(n31549) );
  XOR2_X1 U24984 ( .A1(n14348), .A2(n31510), .Z(n23567) );
  XOR2_X1 U24989 ( .A1(n23184), .A2(n4003), .Z(n31510) );
  NAND2_X2 U24995 ( .A1(n9170), .A2(n22390), .ZN(n22393) );
  XOR2_X1 U24996 ( .A1(n12410), .A2(n31512), .Z(n18200) );
  XOR2_X1 U24998 ( .A1(n19740), .A2(n31513), .Z(n31512) );
  XOR2_X1 U25016 ( .A1(n14645), .A2(n31516), .Z(n13556) );
  NAND2_X1 U25017 ( .A1(n13468), .A2(n13467), .ZN(n31516) );
  INV_X2 U25046 ( .I(n6544), .ZN(n21854) );
  XOR2_X1 U25047 ( .A1(n19509), .A2(n15844), .Z(n19544) );
  INV_X2 U25048 ( .I(n4820), .ZN(n23741) );
  NOR2_X2 U25050 ( .A1(n28616), .A2(n31521), .ZN(n16453) );
  XOR2_X1 U25064 ( .A1(n23258), .A2(n29190), .Z(n17549) );
  XOR2_X1 U25082 ( .A1(n31525), .A2(n29400), .Z(n26433) );
  XOR2_X1 U25088 ( .A1(n1303), .A2(n3142), .Z(n31525) );
  XOR2_X1 U25089 ( .A1(n17551), .A2(n15064), .Z(n19468) );
  NAND2_X2 U25099 ( .A1(n18505), .A2(n18504), .ZN(n17551) );
  XOR2_X1 U25102 ( .A1(n1694), .A2(n19552), .Z(n31527) );
  INV_X2 U25116 ( .I(n13507), .ZN(n13921) );
  XOR2_X1 U25130 ( .A1(n13504), .A2(n12749), .Z(n13507) );
  NAND4_X2 U25131 ( .A1(n28728), .A2(n31528), .A3(n3401), .A4(n17578), .ZN(
        n24189) );
  XOR2_X1 U25132 ( .A1(n3009), .A2(n20926), .Z(n20691) );
  XOR2_X1 U25133 ( .A1(n10949), .A2(n9706), .Z(n8312) );
  XOR2_X1 U25139 ( .A1(n13829), .A2(n31529), .Z(n6209) );
  XOR2_X1 U25146 ( .A1(n19655), .A2(n29426), .Z(n31534) );
  XOR2_X1 U25156 ( .A1(n27951), .A2(n13876), .Z(n292) );
  INV_X2 U25199 ( .I(n19124), .ZN(n16288) );
  NAND2_X2 U25202 ( .A1(n26442), .A2(n10564), .ZN(n19124) );
  XOR2_X1 U25221 ( .A1(n8424), .A2(n11321), .Z(n31538) );
  INV_X2 U25247 ( .I(n16588), .ZN(n31542) );
  NAND2_X1 U25262 ( .A1(n25243), .A2(n31545), .ZN(n4552) );
  OAI21_X2 U25271 ( .A1(n29421), .A2(n31548), .B(n11399), .ZN(n31547) );
  NAND2_X2 U25285 ( .A1(n28205), .A2(n31902), .ZN(n5696) );
  NOR2_X1 U25291 ( .A1(n17338), .A2(n19124), .ZN(n18963) );
  AOI21_X2 U25297 ( .A1(n18106), .A2(n11745), .B(n21055), .ZN(n28396) );
  XOR2_X1 U25298 ( .A1(n22185), .A2(n11458), .Z(n22110) );
  NAND2_X2 U25302 ( .A1(n13034), .A2(n13803), .ZN(n22185) );
  XOR2_X1 U25311 ( .A1(n20960), .A2(n7717), .Z(n20962) );
  XOR2_X1 U25315 ( .A1(n1560), .A2(n16733), .Z(n24762) );
  OR2_X1 U25319 ( .A1(n13382), .A2(n2547), .Z(n7964) );
  NAND2_X2 U25331 ( .A1(n26835), .A2(n26834), .ZN(n10987) );
  NAND2_X2 U25332 ( .A1(n4135), .A2(n23018), .ZN(n22883) );
  XOR2_X1 U25337 ( .A1(n22084), .A2(n22195), .Z(n10462) );
  INV_X2 U25341 ( .I(n31561), .ZN(n4425) );
  INV_X2 U25342 ( .I(n31562), .ZN(n31921) );
  XOR2_X1 U25346 ( .A1(n4222), .A2(n24855), .Z(n31562) );
  NAND3_X2 U25351 ( .A1(n18966), .A2(n18964), .A3(n18965), .ZN(n19398) );
  NAND3_X2 U25354 ( .A1(n13653), .A2(n21863), .A3(n12724), .ZN(n9129) );
  NOR3_X2 U25383 ( .A1(n12280), .A2(n12279), .A3(n1), .ZN(n12276) );
  OAI21_X2 U25401 ( .A1(n12416), .A2(n9377), .B(n29325), .ZN(n12781) );
  NOR2_X1 U25409 ( .A1(n17462), .A2(n31566), .ZN(n28778) );
  XOR2_X1 U25415 ( .A1(n10077), .A2(n10079), .Z(n31671) );
  OAI21_X1 U25426 ( .A1(n25621), .A2(n25705), .B(n31570), .ZN(n31569) );
  XOR2_X1 U25427 ( .A1(n31571), .A2(n24707), .Z(Ciphertext[110]) );
  NOR2_X1 U25435 ( .A1(n21243), .A2(n11912), .ZN(n25942) );
  AOI21_X1 U25438 ( .A1(n31614), .A2(n21147), .B(n15149), .ZN(n4293) );
  XOR2_X1 U25439 ( .A1(n24746), .A2(n24681), .Z(n24684) );
  NOR2_X2 U25442 ( .A1(n6600), .A2(n16445), .ZN(n22121) );
  NAND2_X2 U25447 ( .A1(n17017), .A2(n26998), .ZN(n22138) );
  XOR2_X1 U25455 ( .A1(Plaintext[91]), .A2(Key[91]), .Z(n31574) );
  NOR2_X2 U25461 ( .A1(n28737), .A2(n398), .ZN(n1889) );
  XNOR2_X1 U25466 ( .A1(n7989), .A2(n7988), .ZN(n26699) );
  XOR2_X1 U25468 ( .A1(n3083), .A2(n12014), .Z(n3082) );
  XOR2_X1 U25472 ( .A1(n31575), .A2(n32025), .Z(n28595) );
  AND2_X1 U25479 ( .A1(n6593), .A2(n22955), .Z(n26507) );
  NAND2_X2 U25501 ( .A1(n28081), .A2(n32032), .ZN(n13617) );
  NAND2_X2 U25512 ( .A1(n1956), .A2(n1954), .ZN(n28390) );
  NAND2_X1 U25525 ( .A1(n25963), .A2(n22350), .ZN(n13561) );
  NAND2_X1 U25530 ( .A1(n3448), .A2(n3449), .ZN(n3447) );
  NAND2_X2 U25532 ( .A1(n31585), .A2(n20229), .ZN(n20413) );
  XOR2_X1 U25540 ( .A1(n19679), .A2(n19743), .Z(n19680) );
  NAND2_X1 U25560 ( .A1(n21414), .A2(n8657), .ZN(n5758) );
  XOR2_X1 U25561 ( .A1(n702), .A2(n24527), .Z(n7937) );
  NAND2_X2 U25577 ( .A1(n4985), .A2(n50), .ZN(n702) );
  XOR2_X1 U25584 ( .A1(n4732), .A2(n1262), .Z(n31588) );
  XOR2_X1 U25620 ( .A1(n4756), .A2(n4759), .Z(n6684) );
  XOR2_X1 U25621 ( .A1(n31590), .A2(n22147), .Z(n26462) );
  XOR2_X1 U25624 ( .A1(n19711), .A2(n19398), .Z(n19462) );
  AOI22_X2 U25625 ( .A1(n32028), .A2(n27127), .B1(n146), .B2(n7065), .ZN(
        n31591) );
  OAI21_X2 U25669 ( .A1(n15898), .A2(n1153), .B(n8206), .ZN(n10324) );
  XOR2_X1 U25672 ( .A1(n20804), .A2(n21047), .Z(n20552) );
  NAND2_X1 U25682 ( .A1(n8506), .A2(n19143), .ZN(n16790) );
  INV_X2 U25683 ( .I(n31594), .ZN(n31916) );
  XOR2_X1 U25688 ( .A1(n10536), .A2(n2164), .Z(n31594) );
  XOR2_X1 U25705 ( .A1(n31596), .A2(n23276), .Z(n10536) );
  XOR2_X1 U25714 ( .A1(n13287), .A2(n721), .Z(n31596) );
  XOR2_X1 U25716 ( .A1(n27633), .A2(n29350), .Z(n22223) );
  INV_X2 U25720 ( .I(n22317), .ZN(n31597) );
  XOR2_X1 U25722 ( .A1(n31598), .A2(n3540), .Z(n10430) );
  NAND3_X1 U25733 ( .A1(n27658), .A2(n21365), .A3(n12756), .ZN(n1688) );
  XOR2_X1 U25748 ( .A1(n31599), .A2(n13033), .Z(Ciphertext[161]) );
  XOR2_X1 U25794 ( .A1(n22260), .A2(n21959), .Z(n31606) );
  NAND3_X1 U25796 ( .A1(n29390), .A2(n29508), .A3(n31607), .ZN(n11854) );
  NAND2_X1 U25797 ( .A1(n22659), .A2(n22926), .ZN(n31607) );
  INV_X2 U25800 ( .I(n14983), .ZN(n21568) );
  XOR2_X1 U25808 ( .A1(n24596), .A2(n24634), .Z(n23554) );
  XOR2_X1 U25815 ( .A1(n24740), .A2(n12067), .Z(n24745) );
  XOR2_X1 U25818 ( .A1(n7731), .A2(n24370), .Z(n24740) );
  XOR2_X1 U25831 ( .A1(n8795), .A2(n31608), .Z(n4134) );
  NAND2_X1 U25838 ( .A1(n31617), .A2(n712), .ZN(n1830) );
  OR2_X1 U25847 ( .A1(n16421), .A2(n4145), .Z(n31619) );
  INV_X2 U25855 ( .I(n31622), .ZN(n23603) );
  XOR2_X1 U25857 ( .A1(n22969), .A2(n5263), .Z(n31622) );
  AOI22_X1 U25860 ( .A1(n23643), .A2(n15732), .B1(n6759), .B2(n11888), .ZN(
        n31623) );
  XOR2_X1 U25866 ( .A1(n7363), .A2(n10201), .Z(n23257) );
  XOR2_X1 U25871 ( .A1(n32604), .A2(n3682), .Z(n31626) );
  NAND3_X2 U25873 ( .A1(n21811), .A2(n29864), .A3(n8140), .ZN(n31627) );
  NAND2_X1 U25876 ( .A1(n18582), .A2(n18584), .ZN(n6207) );
  OR2_X1 U25877 ( .A1(n22640), .A2(n31914), .Z(n6242) );
  XOR2_X1 U25886 ( .A1(n31630), .A2(n14217), .Z(n14216) );
  XOR2_X1 U25887 ( .A1(n1004), .A2(n13146), .Z(n31630) );
  INV_X2 U25892 ( .I(n20635), .ZN(n867) );
  XOR2_X1 U25894 ( .A1(n13855), .A2(n13853), .Z(n27698) );
  NAND2_X1 U25901 ( .A1(n22816), .A2(n33675), .ZN(n22818) );
  OAI21_X1 U25914 ( .A1(n2576), .A2(n16023), .B(n21763), .ZN(n26522) );
  NAND2_X1 U25915 ( .A1(n31635), .A2(n31634), .ZN(n22360) );
  XOR2_X1 U25920 ( .A1(n19500), .A2(n29343), .Z(n31638) );
  NAND2_X1 U25921 ( .A1(n14840), .A2(n2826), .ZN(n14592) );
  XOR2_X1 U25925 ( .A1(n1937), .A2(n1936), .Z(n1935) );
  XOR2_X1 U25934 ( .A1(n6091), .A2(n23443), .Z(n6090) );
  NAND2_X2 U25936 ( .A1(n11643), .A2(n11645), .ZN(n22137) );
  XOR2_X1 U25943 ( .A1(n27395), .A2(n31361), .Z(n31642) );
  NAND3_X2 U25944 ( .A1(n2245), .A2(n2247), .A3(n16651), .ZN(n31643) );
  AOI21_X2 U25949 ( .A1(n19994), .A2(n19846), .B(n17882), .ZN(n31644) );
  AND2_X1 U25952 ( .A1(n16354), .A2(n19301), .Z(n19030) );
  INV_X2 U25953 ( .I(n7971), .ZN(n19737) );
  XOR2_X1 U25954 ( .A1(n7971), .A2(n31646), .Z(n101) );
  NAND2_X2 U25955 ( .A1(n19094), .A2(n19095), .ZN(n31658) );
  NAND2_X2 U25964 ( .A1(n27630), .A2(n27631), .ZN(n21681) );
  XOR2_X1 U25987 ( .A1(n9103), .A2(n29445), .Z(n27058) );
  XOR2_X1 U25997 ( .A1(n31655), .A2(n5714), .Z(n560) );
  AND2_X1 U26003 ( .A1(n17341), .A2(n4274), .Z(n31673) );
  OAI22_X1 U26006 ( .A1(n26198), .A2(n24955), .B1(n965), .B2(n24947), .ZN(
        n24941) );
  NOR2_X1 U26012 ( .A1(n27610), .A2(n25057), .ZN(n31661) );
  INV_X1 U26013 ( .I(n27609), .ZN(n31662) );
  NAND2_X1 U26016 ( .A1(n31663), .A2(n17409), .ZN(n11962) );
  NAND2_X2 U26033 ( .A1(n26851), .A2(n15158), .ZN(n10048) );
  XOR2_X1 U26043 ( .A1(n31666), .A2(n24802), .Z(n27812) );
  XOR2_X1 U26044 ( .A1(n24799), .A2(n2864), .Z(n31666) );
  OR2_X1 U26046 ( .A1(n28228), .A2(n7862), .Z(n25102) );
  AOI21_X1 U26047 ( .A1(n31667), .A2(n34167), .B(n23910), .ZN(n12775) );
  NAND2_X2 U26054 ( .A1(n10713), .A2(n18479), .ZN(n7462) );
  NAND2_X2 U26057 ( .A1(n31670), .A2(n31669), .ZN(n10713) );
  NAND2_X1 U26062 ( .A1(n16326), .A2(n16325), .ZN(n27900) );
  NAND2_X2 U26067 ( .A1(n25542), .A2(n25557), .ZN(n25555) );
  INV_X1 U26069 ( .I(n5587), .ZN(n18680) );
  NOR2_X1 U26073 ( .A1(n16805), .A2(n18660), .ZN(n5587) );
  AOI21_X2 U26075 ( .A1(n21169), .A2(n11678), .B(n31674), .ZN(n3001) );
  AOI21_X2 U26076 ( .A1(n15843), .A2(n15842), .B(n19282), .ZN(n15844) );
  NAND2_X2 U26082 ( .A1(n27900), .A2(n23978), .ZN(n25973) );
  AOI22_X2 U26083 ( .A1(n7997), .A2(n30692), .B1(n17442), .B2(n17441), .ZN(
        n31675) );
  NAND2_X2 U26087 ( .A1(n31676), .A2(n27992), .ZN(n20335) );
  XOR2_X1 U26094 ( .A1(n26279), .A2(n14791), .Z(n14190) );
  NOR2_X2 U26095 ( .A1(n19284), .A2(n10943), .ZN(n28949) );
  NAND2_X1 U26096 ( .A1(n19523), .A2(n31678), .ZN(n19528) );
  NAND2_X1 U26097 ( .A1(n15593), .A2(n19834), .ZN(n31678) );
  XOR2_X1 U26099 ( .A1(n2353), .A2(n17968), .Z(n26996) );
  NOR2_X1 U26102 ( .A1(n793), .A2(n719), .ZN(n31679) );
  XOR2_X1 U26107 ( .A1(n31043), .A2(n5101), .Z(n5100) );
  XOR2_X1 U26112 ( .A1(n24782), .A2(n27153), .Z(n13086) );
  NOR3_X1 U26113 ( .A1(n25546), .A2(n25557), .A3(n25542), .ZN(n15132) );
  XOR2_X1 U26117 ( .A1(n9327), .A2(n19689), .Z(n9326) );
  XOR2_X1 U26118 ( .A1(n19589), .A2(n19508), .Z(n19689) );
  NOR3_X1 U26124 ( .A1(n17306), .A2(n15425), .A3(n29063), .ZN(n6849) );
  INV_X2 U26126 ( .I(n14911), .ZN(n29063) );
  XNOR2_X1 U26136 ( .A1(n23498), .A2(n23497), .ZN(n31709) );
  OAI21_X2 U26142 ( .A1(n18813), .A2(n17370), .B(n31682), .ZN(n8741) );
  BUF_X2 U26147 ( .I(n16811), .Z(n31683) );
  OAI21_X2 U26154 ( .A1(n2060), .A2(n3821), .B(n31686), .ZN(n1917) );
  AOI22_X2 U26155 ( .A1(n534), .A2(n1326), .B1(n1), .B2(n16736), .ZN(n31686)
         );
  XOR2_X1 U26160 ( .A1(n24636), .A2(n24832), .Z(n24600) );
  OR2_X1 U26163 ( .A1(n27419), .A2(n33675), .Z(n22817) );
  NOR2_X1 U26167 ( .A1(n12329), .A2(n32900), .ZN(n25078) );
  OAI21_X2 U26168 ( .A1(n6204), .A2(n28706), .B(n24889), .ZN(n14650) );
  NAND2_X2 U26174 ( .A1(n31695), .A2(n31693), .ZN(n19909) );
  NAND3_X1 U26175 ( .A1(n4143), .A2(n16298), .A3(n4142), .ZN(n31695) );
  NOR2_X1 U26183 ( .A1(n8010), .A2(n8605), .ZN(n16779) );
  XOR2_X1 U26191 ( .A1(n19620), .A2(n31698), .Z(n11545) );
  XOR2_X1 U26193 ( .A1(n19619), .A2(n1173), .Z(n31698) );
  AOI21_X2 U26194 ( .A1(n26133), .A2(n2277), .B(n31699), .ZN(n2272) );
  OAI21_X2 U26196 ( .A1(n26798), .A2(n28714), .B(n3673), .ZN(n31699) );
  XOR2_X1 U26199 ( .A1(n10697), .A2(n23331), .Z(n31703) );
  AOI22_X2 U26202 ( .A1(n3113), .A2(n3112), .B1(n3111), .B2(n28573), .ZN(n3340) );
  XOR2_X1 U26205 ( .A1(n24521), .A2(n14920), .Z(n31704) );
  XOR2_X1 U26213 ( .A1(n31706), .A2(n31913), .Z(n27792) );
  NAND2_X2 U26220 ( .A1(n1256), .A2(n27219), .ZN(n26716) );
  XOR2_X1 U26221 ( .A1(n2900), .A2(n29463), .Z(n26537) );
  XOR2_X1 U26222 ( .A1(n22239), .A2(n22240), .Z(n12898) );
  XOR2_X1 U26229 ( .A1(n24489), .A2(n15744), .Z(n15743) );
  INV_X2 U26230 ( .I(n24197), .ZN(n27430) );
  NAND3_X2 U26231 ( .A1(n26211), .A2(n23676), .A3(n23677), .ZN(n24197) );
  OAI21_X1 U26247 ( .A1(n15912), .A2(n11516), .B(n29271), .ZN(n8914) );
  NAND3_X2 U26250 ( .A1(n31710), .A2(n18384), .A3(n17649), .ZN(n3836) );
  NAND2_X2 U26251 ( .A1(n18559), .A2(n18494), .ZN(n11774) );
  XOR2_X1 U26254 ( .A1(Plaintext[77]), .A2(Key[77]), .Z(n18494) );
  BUF_X2 U26255 ( .I(n24847), .Z(n31713) );
  NAND2_X2 U26261 ( .A1(n31834), .A2(n31714), .ZN(n20399) );
  NAND3_X1 U26275 ( .A1(n24051), .A2(n14490), .A3(n4897), .ZN(n305) );
  OAI22_X1 U26279 ( .A1(n15857), .A2(n11998), .B1(n15855), .B2(n15854), .ZN(
        n26295) );
  INV_X2 U26281 ( .I(n31716), .ZN(n17516) );
  XOR2_X1 U26284 ( .A1(Plaintext[126]), .A2(Key[126]), .Z(n31716) );
  NAND3_X2 U26288 ( .A1(n31718), .A2(n24038), .A3(n24039), .ZN(n24416) );
  XOR2_X1 U26291 ( .A1(n24758), .A2(n31719), .Z(n28968) );
  XOR2_X1 U26292 ( .A1(n5539), .A2(n31720), .Z(n31719) );
  INV_X1 U26294 ( .I(n16619), .ZN(n31720) );
  OAI22_X2 U26297 ( .A1(n19605), .A2(n29730), .B1(n2717), .B2(n19196), .ZN(
        n1944) );
  NOR2_X2 U26300 ( .A1(n3207), .A2(n19195), .ZN(n19605) );
  INV_X2 U26305 ( .I(n736), .ZN(n25539) );
  XOR2_X1 U26314 ( .A1(n8617), .A2(n25156), .Z(n610) );
  XOR2_X1 U26321 ( .A1(n15130), .A2(n8762), .Z(n27011) );
  NAND3_X2 U26324 ( .A1(n28846), .A2(n7582), .A3(n22276), .ZN(n15130) );
  XOR2_X1 U26330 ( .A1(n27763), .A2(n23346), .Z(n23498) );
  XOR2_X1 U26335 ( .A1(n24405), .A2(n24404), .Z(n31725) );
  INV_X2 U26337 ( .I(n8106), .ZN(n31730) );
  AOI21_X2 U26338 ( .A1(n31732), .A2(n21644), .B(n3418), .ZN(n22119) );
  NAND3_X2 U26339 ( .A1(n29389), .A2(n31893), .A3(n5424), .ZN(n5612) );
  AOI21_X2 U26345 ( .A1(n31736), .A2(n29158), .B(n3495), .ZN(n7905) );
  NAND2_X2 U26350 ( .A1(n31344), .A2(n9022), .ZN(n31736) );
  XOR2_X1 U26354 ( .A1(n31738), .A2(n31737), .Z(n31787) );
  XOR2_X1 U26355 ( .A1(n23277), .A2(n23234), .Z(n31738) );
  OR2_X1 U26356 ( .A1(n421), .A2(n6581), .Z(n26204) );
  XOR2_X1 U26373 ( .A1(n31739), .A2(n25908), .Z(Ciphertext[187]) );
  OAI22_X1 U26377 ( .A1(n7716), .A2(n25907), .B1(n25927), .B2(n690), .ZN(
        n31739) );
  OAI22_X1 U26378 ( .A1(n1094), .A2(n24044), .B1(n23602), .B2(n13412), .ZN(
        n26966) );
  AOI22_X2 U26388 ( .A1(n28491), .A2(n6453), .B1(n23111), .B2(n853), .ZN(n5893) );
  NAND2_X2 U26390 ( .A1(n28003), .A2(n9080), .ZN(n16429) );
  NOR2_X1 U26391 ( .A1(n11923), .A2(n6479), .ZN(n7444) );
  XNOR2_X1 U26392 ( .A1(n9185), .A2(n32861), .ZN(n16382) );
  AND2_X1 U26394 ( .A1(n5034), .A2(n28157), .Z(n19238) );
  NOR2_X1 U26399 ( .A1(n20052), .A2(n13327), .ZN(n31745) );
  XOR2_X1 U26403 ( .A1(n31747), .A2(n16125), .Z(n3339) );
  NOR2_X2 U26404 ( .A1(n31748), .A2(n15808), .ZN(n11744) );
  XOR2_X1 U26414 ( .A1(n8809), .A2(n31749), .Z(n8302) );
  XOR2_X1 U26416 ( .A1(n26230), .A2(n19755), .Z(n8809) );
  NAND2_X2 U26418 ( .A1(n20379), .A2(n6679), .ZN(n11303) );
  AND2_X1 U26424 ( .A1(n636), .A2(n1119), .Z(n28902) );
  XOR2_X1 U26426 ( .A1(n1590), .A2(n1587), .Z(n1589) );
  OAI21_X1 U26430 ( .A1(n31954), .A2(n2386), .B(n423), .ZN(n21644) );
  NAND2_X2 U26434 ( .A1(n6629), .A2(n12163), .ZN(n7555) );
  XOR2_X1 U26440 ( .A1(n17554), .A2(n20836), .Z(n20957) );
  OAI22_X2 U26442 ( .A1(n20048), .A2(n20047), .B1(n20546), .B2(n28904), .ZN(
        n20836) );
  XOR2_X1 U26443 ( .A1(n31751), .A2(n15470), .Z(n15092) );
  XOR2_X1 U26446 ( .A1(n22222), .A2(n22049), .Z(n9701) );
  XOR2_X1 U26447 ( .A1(n21913), .A2(n31457), .Z(n22049) );
  INV_X2 U26449 ( .I(n31753), .ZN(n26040) );
  XOR2_X1 U26450 ( .A1(Plaintext[25]), .A2(Key[25]), .Z(n31753) );
  XOR2_X1 U26451 ( .A1(n21481), .A2(n31105), .Z(n31754) );
  AOI21_X2 U26452 ( .A1(n26253), .A2(n13129), .B(n3659), .ZN(n3658) );
  XOR2_X1 U26454 ( .A1(n2384), .A2(n5647), .Z(n31756) );
  NAND2_X2 U26456 ( .A1(n18405), .A2(n3051), .ZN(n3060) );
  XOR2_X1 U26458 ( .A1(n16838), .A2(n31761), .Z(n188) );
  XOR2_X1 U26459 ( .A1(n31762), .A2(n28898), .Z(n31761) );
  NAND2_X1 U26460 ( .A1(n31763), .A2(n9558), .ZN(n26431) );
  NOR2_X1 U26461 ( .A1(n26142), .A2(n5395), .ZN(n31763) );
  XOR2_X1 U26462 ( .A1(n10789), .A2(n10788), .Z(n27732) );
  NAND2_X2 U26466 ( .A1(n5645), .A2(n31767), .ZN(n7345) );
  AOI22_X2 U26467 ( .A1(n5644), .A2(n18571), .B1(n953), .B2(n485), .ZN(n31767)
         );
  AOI22_X1 U26468 ( .A1(n1757), .A2(n1758), .B1(n1756), .B2(n13023), .ZN(
        n28116) );
  XOR2_X1 U26469 ( .A1(n21041), .A2(n4021), .Z(n31769) );
  XOR2_X1 U26470 ( .A1(n31770), .A2(n6940), .Z(n6938) );
  XOR2_X1 U26471 ( .A1(n24692), .A2(n24376), .Z(n31770) );
  XOR2_X1 U26472 ( .A1(n22171), .A2(n17258), .Z(n16861) );
  XOR2_X1 U26473 ( .A1(n31771), .A2(n8020), .Z(n17721) );
  NAND2_X1 U26475 ( .A1(n9249), .A2(n9248), .ZN(n9251) );
  XOR2_X1 U26479 ( .A1(n1851), .A2(n6574), .Z(n29228) );
  XOR2_X1 U26480 ( .A1(n18398), .A2(Key[184]), .Z(n31773) );
  NOR2_X2 U26484 ( .A1(n28836), .A2(n6530), .ZN(n31776) );
  NAND2_X2 U26486 ( .A1(n10656), .A2(n10655), .ZN(n9076) );
  OAI21_X2 U26490 ( .A1(n12029), .A2(n16484), .B(n4518), .ZN(n31777) );
  NOR2_X2 U26491 ( .A1(n18266), .A2(n18265), .ZN(n4858) );
  OAI22_X2 U26492 ( .A1(n20426), .A2(n12421), .B1(n20428), .B2(n32747), .ZN(
        n18265) );
  NAND2_X2 U26493 ( .A1(n31780), .A2(n31778), .ZN(n25136) );
  OAI21_X2 U26495 ( .A1(n7969), .A2(n196), .B(n31960), .ZN(n31781) );
  BUF_X2 U26496 ( .I(n16267), .Z(n31784) );
  INV_X2 U26497 ( .I(n4036), .ZN(n10579) );
  XOR2_X1 U26498 ( .A1(Plaintext[29]), .A2(Key[29]), .Z(n4036) );
  AOI21_X2 U26499 ( .A1(n25523), .A2(n27236), .B(n31786), .ZN(n25369) );
  INV_X2 U26500 ( .I(n13113), .ZN(n16386) );
  INV_X2 U26502 ( .I(n31787), .ZN(n23834) );
  OAI22_X1 U26503 ( .A1(n25380), .A2(n25379), .B1(n25377), .B2(n30302), .ZN(
        n27487) );
  AOI21_X1 U26504 ( .A1(n18459), .A2(n956), .B(n16854), .ZN(n7163) );
  INV_X2 U26505 ( .I(n17261), .ZN(n24265) );
  NAND2_X2 U26506 ( .A1(n12774), .A2(n26967), .ZN(n17261) );
  NOR2_X2 U26508 ( .A1(n28974), .A2(n31790), .ZN(n28782) );
  XOR2_X1 U26509 ( .A1(n19660), .A2(n29341), .Z(n26003) );
  INV_X2 U26512 ( .I(n22949), .ZN(n31795) );
  NAND2_X2 U26513 ( .A1(n6733), .A2(n19840), .ZN(n20431) );
  INV_X2 U26514 ( .I(n31797), .ZN(n26078) );
  NAND2_X1 U26515 ( .A1(n26817), .A2(n14625), .ZN(n31799) );
  XOR2_X1 U26516 ( .A1(n31800), .A2(n19443), .Z(n28216) );
  XOR2_X1 U26517 ( .A1(n27444), .A2(n7057), .Z(n31800) );
  XOR2_X1 U26521 ( .A1(n24602), .A2(n31803), .Z(n7535) );
  XOR2_X1 U26522 ( .A1(n25991), .A2(n7828), .Z(n31803) );
  NAND2_X2 U26526 ( .A1(n5418), .A2(n4191), .ZN(n26683) );
  XOR2_X1 U26529 ( .A1(n19543), .A2(n19702), .Z(n7375) );
  OAI22_X2 U26530 ( .A1(n229), .A2(n15920), .B1(n15919), .B2(n16724), .ZN(
        n31824) );
  OAI21_X2 U26534 ( .A1(n2744), .A2(n32298), .B(n14663), .ZN(n31813) );
  OAI21_X2 U26535 ( .A1(n18141), .A2(n20142), .B(n1458), .ZN(n31814) );
  INV_X2 U26543 ( .I(n31819), .ZN(n18960) );
  NOR2_X2 U26544 ( .A1(n4747), .A2(n12585), .ZN(n31819) );
  NAND2_X2 U26545 ( .A1(n6750), .A2(n6749), .ZN(n15829) );
  NOR2_X2 U26546 ( .A1(n31820), .A2(n29602), .ZN(n448) );
  INV_X2 U26547 ( .I(n25892), .ZN(n31822) );
  OAI21_X1 U26548 ( .A1(n773), .A2(n22945), .B(n31825), .ZN(n8923) );
  NOR2_X1 U26550 ( .A1(n16832), .A2(n18977), .ZN(n5842) );
  XOR2_X1 U26552 ( .A1(n19671), .A2(n17689), .Z(n26738) );
  AOI22_X2 U26553 ( .A1(n31827), .A2(n1055), .B1(n4749), .B2(n28478), .ZN(
        n11777) );
  OAI21_X2 U26554 ( .A1(n1175), .A2(n1051), .B(n25961), .ZN(n31827) );
  NOR2_X2 U26558 ( .A1(n31830), .A2(n29094), .ZN(n1474) );
  NOR2_X1 U26559 ( .A1(n19601), .A2(n10860), .ZN(n19614) );
  NAND2_X2 U26561 ( .A1(n28844), .A2(n20182), .ZN(n20775) );
  XOR2_X1 U26562 ( .A1(n9586), .A2(n17538), .Z(n3982) );
  XOR2_X1 U26564 ( .A1(n13586), .A2(n4329), .Z(n27152) );
  NOR2_X1 U26567 ( .A1(n5786), .A2(n12885), .ZN(n31833) );
  OAI21_X2 U26571 ( .A1(n31836), .A2(n16184), .B(n8539), .ZN(n21498) );
  NOR2_X2 U26572 ( .A1(n31030), .A2(n1333), .ZN(n31836) );
  NAND2_X2 U26573 ( .A1(n31923), .A2(n12610), .ZN(n5602) );
  XOR2_X1 U26575 ( .A1(n19409), .A2(n17551), .Z(n19732) );
  INV_X2 U26576 ( .I(n31839), .ZN(n9910) );
  AOI21_X2 U26579 ( .A1(n26591), .A2(n18729), .B(n31980), .ZN(n25971) );
  NOR2_X2 U26580 ( .A1(n13616), .A2(n13615), .ZN(n13614) );
  NOR2_X1 U26583 ( .A1(n17669), .A2(n23087), .ZN(n17668) );
  XOR2_X1 U26586 ( .A1(n9674), .A2(n31841), .Z(n28607) );
  XOR2_X1 U26587 ( .A1(n22171), .A2(n16027), .Z(n27312) );
  XOR2_X1 U26588 ( .A1(n6689), .A2(n6686), .Z(n10248) );
  XOR2_X1 U26590 ( .A1(n22113), .A2(n22196), .Z(n22289) );
  BUF_X2 U26591 ( .I(n3504), .Z(n31843) );
  XOR2_X1 U26592 ( .A1(n31844), .A2(n5846), .Z(n5844) );
  XOR2_X1 U26594 ( .A1(n19470), .A2(n27607), .Z(n5925) );
  XOR2_X1 U26599 ( .A1(n31849), .A2(n24539), .Z(n29277) );
  NAND2_X2 U26603 ( .A1(n3045), .A2(n3047), .ZN(n22227) );
  XOR2_X1 U26607 ( .A1(n3209), .A2(n2661), .Z(n31852) );
  NAND2_X2 U26608 ( .A1(n3211), .A2(n31853), .ZN(n21779) );
  AOI22_X2 U26612 ( .A1(n14828), .A2(n16915), .B1(n18464), .B2(n18489), .ZN(
        n31856) );
  NAND3_X2 U26613 ( .A1(n1772), .A2(n26979), .A3(n615), .ZN(n29137) );
  NAND2_X2 U26616 ( .A1(n13850), .A2(n12228), .ZN(n13041) );
  XOR2_X1 U26619 ( .A1(n23333), .A2(n1260), .Z(n23128) );
  OAI21_X1 U26620 ( .A1(n964), .A2(n713), .B(n7941), .ZN(n5903) );
  XOR2_X1 U26621 ( .A1(n12258), .A2(n29832), .Z(n26920) );
  OAI21_X2 U26622 ( .A1(n4497), .A2(n4496), .B(n26152), .ZN(n12211) );
  XOR2_X1 U26623 ( .A1(n14407), .A2(n13299), .Z(n4572) );
  NOR2_X2 U26624 ( .A1(n18699), .A2(n22), .ZN(n18833) );
  INV_X1 U26625 ( .I(n15139), .ZN(n18699) );
  XOR2_X1 U26626 ( .A1(n18388), .A2(Key[111]), .Z(n15139) );
  XOR2_X1 U26627 ( .A1(n22284), .A2(n22003), .Z(n1762) );
  BUF_X2 U26628 ( .I(n24616), .Z(n31866) );
  XOR2_X1 U26631 ( .A1(n9092), .A2(n9093), .Z(n31869) );
  NAND3_X2 U26632 ( .A1(n14838), .A2(n24344), .A3(n24342), .ZN(n24531) );
  NAND2_X2 U26636 ( .A1(n9561), .A2(n24084), .ZN(n24137) );
  NAND2_X2 U26637 ( .A1(n3170), .A2(n3172), .ZN(n7772) );
  NAND2_X1 U26638 ( .A1(n17535), .A2(n11957), .ZN(n24730) );
  AND2_X1 U26639 ( .A1(n23717), .A2(n10967), .Z(n23682) );
  NAND2_X2 U26640 ( .A1(n3845), .A2(n23999), .ZN(n24533) );
  XOR2_X1 U26642 ( .A1(n5194), .A2(n31875), .Z(n27883) );
  AOI21_X1 U26644 ( .A1(n25044), .A2(n31876), .B(n25062), .ZN(n8258) );
  NAND2_X1 U26645 ( .A1(n25058), .A2(n25057), .ZN(n31876) );
  OAI21_X1 U26646 ( .A1(n3229), .A2(n2983), .B(n14865), .ZN(n2264) );
  NOR2_X1 U26647 ( .A1(n20276), .A2(n14187), .ZN(n20277) );
  XOR2_X1 U26648 ( .A1(n6421), .A2(n31880), .Z(n25146) );
  XOR2_X1 U26649 ( .A1(n24840), .A2(n29417), .Z(n31880) );
  OAI21_X2 U26654 ( .A1(n11693), .A2(n17843), .B(n31885), .ZN(n18658) );
  NAND2_X2 U26655 ( .A1(n17843), .A2(n18446), .ZN(n31885) );
  XOR2_X1 U26657 ( .A1(n5184), .A2(n29412), .Z(n31887) );
  NAND2_X1 U26658 ( .A1(n31888), .A2(n16083), .ZN(n2729) );
  NOR2_X1 U26659 ( .A1(n23620), .A2(n30360), .ZN(n31888) );
  XOR2_X1 U26660 ( .A1(n20802), .A2(n25266), .Z(n7595) );
  OAI22_X2 U26661 ( .A1(n9587), .A2(n9588), .B1(n20075), .B2(n20360), .ZN(
        n20802) );
  BUF_X2 U26662 ( .I(n10312), .Z(n31891) );
  XOR2_X1 U26664 ( .A1(n28753), .A2(n23518), .Z(n31892) );
  NOR2_X1 U26665 ( .A1(n21848), .A2(n30291), .ZN(n12852) );
  AOI21_X2 U26666 ( .A1(n5611), .A2(n1216), .B(n31895), .ZN(n28304) );
  AOI21_X2 U26667 ( .A1(n8031), .A2(n7577), .B(n31898), .ZN(n7157) );
  XOR2_X1 U26669 ( .A1(n24573), .A2(n25991), .Z(n31899) );
  XOR2_X1 U26673 ( .A1(n26540), .A2(n24402), .Z(n31901) );
  NAND2_X1 U26677 ( .A1(n7334), .A2(n32859), .ZN(n31904) );
  XOR2_X1 U26680 ( .A1(n26075), .A2(n4771), .Z(n392) );
  XOR2_X1 U26681 ( .A1(n20849), .A2(n6857), .Z(n4771) );
  XOR2_X1 U26682 ( .A1(n19577), .A2(n19578), .Z(n4465) );
  INV_X2 U26683 ( .I(n19958), .ZN(n27808) );
  INV_X1 U26684 ( .I(n26088), .ZN(n20090) );
  INV_X2 U26686 ( .I(n26194), .ZN(n505) );
  NOR2_X2 U26688 ( .A1(n13314), .A2(n13310), .ZN(n21122) );
  NAND2_X2 U26689 ( .A1(n27249), .A2(n28549), .ZN(n28232) );
  XNOR2_X1 U26690 ( .A1(n22067), .A2(n16482), .ZN(n31912) );
  XNOR2_X1 U26691 ( .A1(n6771), .A2(n10935), .ZN(n31913) );
  INV_X2 U26692 ( .I(n3536), .ZN(n22491) );
  INV_X1 U26694 ( .I(n9953), .ZN(n11804) );
  INV_X1 U26695 ( .I(n6407), .ZN(n22362) );
  AND2_X1 U4340 ( .A1(n27077), .A2(n30010), .Z(n1490) );
  INV_X2 U1051 ( .I(n21704), .ZN(n26782) );
  NAND2_X2 U1695 ( .A1(n10323), .A2(n15434), .ZN(n7961) );
  AOI21_X2 U5747 ( .A1(n8022), .A2(n1271), .B(n12220), .ZN(n9918) );
  INV_X4 U14047 ( .I(n20052), .ZN(n19949) );
  BUF_X4 U3960 ( .I(n7251), .Z(n29223) );
  INV_X2 U1145 ( .I(n13712), .ZN(n26735) );
  INV_X2 U1873 ( .I(n26699), .ZN(n29200) );
  INV_X2 U5133 ( .I(n4289), .ZN(n20575) );
  INV_X2 U5403 ( .I(n17237), .ZN(n20570) );
  INV_X2 U1119 ( .I(n11063), .ZN(n15002) );
  NOR2_X2 U15357 ( .A1(n4665), .A2(n4664), .ZN(n4329) );
  INV_X2 U3390 ( .I(n18487), .ZN(n26520) );
  NAND3_X2 U15563 ( .A1(n23828), .A2(n23953), .A3(n13281), .ZN(n4824) );
  INV_X2 U7038 ( .I(n9871), .ZN(n22503) );
  NAND2_X2 U5912 ( .A1(n29365), .A2(n19826), .ZN(n30748) );
  NAND2_X2 U8233 ( .A1(n21107), .A2(n10546), .ZN(n21510) );
  NAND3_X2 U2384 ( .A1(n20949), .A2(n5822), .A3(n29062), .ZN(n20950) );
  BUF_X4 U867 ( .I(n17201), .Z(n29222) );
  OR2_X2 U14806 ( .A1(n6407), .A2(n11805), .Z(n12869) );
  NAND3_X2 U121 ( .A1(n11306), .A2(n25565), .A3(n11900), .ZN(n2018) );
  INV_X2 U54 ( .I(n25686), .ZN(n29243) );
  INV_X2 U2203 ( .I(n21761), .ZN(n21847) );
  NAND3_X2 U23123 ( .A1(n20178), .A2(n20179), .A3(n33301), .ZN(n20182) );
  INV_X2 U3531 ( .I(n10170), .ZN(n25695) );
  NAND2_X2 U1425 ( .A1(n18035), .A2(n10679), .ZN(n26848) );
  INV_X2 U10624 ( .I(n24235), .ZN(n10627) );
  INV_X4 U4438 ( .I(n561), .ZN(n1083) );
  OR2_X2 U11379 ( .A1(n21350), .A2(n30389), .Z(n21571) );
  AOI21_X2 U17315 ( .A1(n14473), .A2(n16943), .B(n4891), .ZN(n27446) );
  NAND2_X2 U21045 ( .A1(n981), .A2(n8217), .ZN(n16943) );
  NOR2_X2 U6595 ( .A1(n31108), .A2(n19052), .ZN(n3092) );
  BUF_X4 U1587 ( .I(n25185), .Z(n15641) );
  BUF_X4 U17991 ( .I(n10292), .Z(n30571) );
  NOR3_X2 U4868 ( .A1(n2296), .A2(n34046), .A3(n1322), .ZN(n2339) );
  INV_X2 U21491 ( .I(n19244), .ZN(n14698) );
  NAND2_X2 U3667 ( .A1(n30010), .A2(n4202), .ZN(n19244) );
  NAND2_X2 U4859 ( .A1(n1322), .A2(n34046), .ZN(n21830) );
  INV_X2 U14769 ( .I(n24147), .ZN(n24120) );
  NAND2_X2 U2978 ( .A1(n19234), .A2(n29003), .ZN(n8119) );
  OR2_X1 U5167 ( .A1(n8933), .A2(n4881), .Z(n11785) );
  NAND2_X2 U1690 ( .A1(n13920), .A2(n26881), .ZN(n9364) );
  INV_X4 U4967 ( .I(n19249), .ZN(n16274) );
  INV_X2 U6141 ( .I(n470), .ZN(n31670) );
  AND2_X2 U26023 ( .A1(n2207), .A2(n15411), .Z(n12316) );
  INV_X2 U1603 ( .I(n16122), .ZN(n27909) );
  NOR2_X2 U13418 ( .A1(n7673), .A2(n1333), .ZN(n26997) );
  NOR2_X2 U5917 ( .A1(n2606), .A2(n16630), .ZN(n20060) );
  BUF_X4 U15425 ( .I(n16453), .Z(n7557) );
  NAND2_X2 U14180 ( .A1(n16374), .A2(n9352), .ZN(n10231) );
  NOR2_X2 U23171 ( .A1(n9895), .A2(n8331), .ZN(n22048) );
  INV_X2 U3316 ( .I(n10285), .ZN(n25739) );
  INV_X4 U16585 ( .I(n13413), .ZN(n23756) );
  BUF_X2 U150 ( .I(n18242), .Z(n30512) );
  INV_X2 U3433 ( .I(n7280), .ZN(n7279) );
  NAND2_X2 U3187 ( .A1(n7195), .A2(n9663), .ZN(n9664) );
  NAND2_X2 U10260 ( .A1(n7044), .A2(n26777), .ZN(n21214) );
  NAND2_X2 U3464 ( .A1(n15179), .A2(n24254), .ZN(n13378) );
  AOI21_X2 U6410 ( .A1(n31765), .A2(n33139), .B(n17139), .ZN(n2741) );
  OAI21_X2 U2405 ( .A1(n12113), .A2(n10085), .B(n30512), .ZN(n14579) );
  NAND2_X2 U4135 ( .A1(n7486), .A2(n16374), .ZN(n28167) );
  NOR2_X2 U23081 ( .A1(n27336), .A2(n15026), .ZN(n21612) );
  INV_X4 U6334 ( .I(n22599), .ZN(n9580) );
  BUF_X2 U6036 ( .I(n27698), .Z(n29339) );
  NAND2_X2 U2902 ( .A1(n3077), .A2(n30191), .ZN(n24270) );
  INV_X2 U4665 ( .I(n25615), .ZN(n1202) );
  OAI22_X2 U12698 ( .A1(n3779), .A2(n18511), .B1(n12327), .B2(n11380), .ZN(
        n17130) );
  NOR2_X2 U7845 ( .A1(n29518), .A2(n12094), .ZN(n29138) );
  OAI21_X2 U3069 ( .A1(n22866), .A2(n23068), .B(n10641), .ZN(n12529) );
  NOR2_X2 U15717 ( .A1(n18791), .A2(n13548), .ZN(n9511) );
  NAND2_X2 U14677 ( .A1(n21702), .A2(n33833), .ZN(n6764) );
  AOI21_X2 U299 ( .A1(n11236), .A2(n32176), .B(n10381), .ZN(n3678) );
  NAND2_X2 U3269 ( .A1(n28338), .A2(n25756), .ZN(n25875) );
  BUF_X4 U3048 ( .I(n15715), .Z(n5471) );
  INV_X2 U44 ( .I(n32063), .ZN(n26198) );
  INV_X2 U2804 ( .I(n25897), .ZN(n27118) );
  AOI21_X2 U15211 ( .A1(n26185), .A2(n14463), .B(n33103), .ZN(n30625) );
  NOR2_X2 U9307 ( .A1(n22747), .A2(n1278), .ZN(n12220) );
  NAND2_X1 U11090 ( .A1(n15007), .A2(n1125), .ZN(n9451) );
  NOR2_X2 U7167 ( .A1(n1703), .A2(n32452), .ZN(n21161) );
  INV_X4 U2078 ( .I(n23085), .ZN(n17639) );
  INV_X4 U3302 ( .I(n25620), .ZN(n8186) );
  NAND2_X2 U14727 ( .A1(n28081), .A2(n32032), .ZN(n27113) );
  INV_X4 U18939 ( .I(n29200), .ZN(n30692) );
  BUF_X4 U1670 ( .I(n14564), .Z(n4468) );
  NAND2_X2 U1323 ( .A1(n19063), .A2(n19108), .ZN(n19365) );
  BUF_X2 U265 ( .I(n10170), .Z(n4146) );
  AOI22_X2 U1579 ( .A1(n9668), .A2(n9667), .B1(n11098), .B2(n1182), .ZN(n10481) );
  INV_X4 U8820 ( .I(n470), .ZN(n14213) );
  INV_X2 U807 ( .I(n7024), .ZN(n16225) );
  OAI21_X2 U5354 ( .A1(n13127), .A2(n31934), .B(n22444), .ZN(n17462) );
  INV_X2 U1040 ( .I(n156), .ZN(n13371) );
  AND2_X1 U4484 ( .A1(n18037), .A2(n8964), .Z(n22536) );
  INV_X2 U1800 ( .I(n19423), .ZN(n4942) );
  BUF_X2 U2549 ( .I(n24682), .Z(n27385) );
  BUF_X4 U1217 ( .I(n12211), .Z(n1008) );
  INV_X2 U5227 ( .I(n29272), .ZN(n980) );
  NAND3_X2 U800 ( .A1(n31506), .A2(n22488), .A3(n22489), .ZN(n10832) );
  INV_X2 U2279 ( .I(n713), .ZN(n314) );
  OAI21_X2 U639 ( .A1(n10895), .A2(n22900), .B(n3830), .ZN(n31758) );
  INV_X4 U4046 ( .I(n17184), .ZN(n957) );
  NOR2_X2 U14889 ( .A1(n23085), .A2(n23087), .ZN(n22967) );
  NAND2_X2 U5182 ( .A1(n16435), .A2(n18602), .ZN(n15909) );
  NOR2_X2 U17651 ( .A1(n10085), .A2(n7963), .ZN(n25839) );
  INV_X4 U4881 ( .I(n9220), .ZN(n12143) );
  AOI21_X2 U6555 ( .A1(n12912), .A2(n12911), .B(n810), .ZN(n26595) );
  NAND2_X2 U8503 ( .A1(n4639), .A2(n19883), .ZN(n4638) );
  NAND2_X2 U26384 ( .A1(n12257), .A2(n24873), .ZN(n8777) );
  NOR2_X2 U1360 ( .A1(n21839), .A2(n27937), .ZN(n13030) );
  BUF_X4 U4400 ( .I(n33146), .Z(n3468) );
  AND2_X1 U4761 ( .A1(n28329), .A2(n9430), .Z(n10045) );
  OAI21_X1 U21161 ( .A1(n12831), .A2(n12707), .B(n18922), .ZN(n12830) );
  AND2_X2 U1809 ( .A1(n2499), .A2(n12379), .Z(n20079) );
  INV_X2 U7587 ( .I(n15146), .ZN(n18892) );
  INV_X2 U20711 ( .I(n11677), .ZN(n12037) );
  NOR2_X2 U6718 ( .A1(n22666), .A2(n22664), .ZN(n26406) );
  INV_X2 U3993 ( .I(n12044), .ZN(n21406) );
  INV_X2 U2725 ( .I(n25295), .ZN(n25398) );
  INV_X2 U3686 ( .I(n25429), .ZN(n25453) );
  NAND2_X2 U2727 ( .A1(n25295), .A2(n25397), .ZN(n27586) );
  INV_X2 U3437 ( .I(n16534), .ZN(n842) );
  NAND3_X2 U10878 ( .A1(n13251), .A2(n1108), .A3(n1109), .ZN(n16928) );
  NAND2_X2 U943 ( .A1(n3567), .A2(n30529), .ZN(n11202) );
  INV_X2 U2930 ( .I(n31965), .ZN(n1017) );
  INV_X2 U24696 ( .I(n20614), .ZN(n20392) );
  INV_X2 U20610 ( .I(n18873), .ZN(n11460) );
  INV_X2 U207 ( .I(n6286), .ZN(n1239) );
  NAND2_X2 U11504 ( .A1(n28860), .A2(n28635), .ZN(n26682) );
  OAI22_X2 U6767 ( .A1(n27415), .A2(n16149), .B1(n22664), .B2(n16567), .ZN(
        n28860) );
  NOR2_X2 U5310 ( .A1(n23949), .A2(n11676), .ZN(n11708) );
  AND2_X1 U4052 ( .A1(n12211), .A2(n30690), .Z(n31335) );
  NAND2_X2 U8815 ( .A1(n15956), .A2(n13738), .ZN(n18463) );
  INV_X2 U5046 ( .I(n9375), .ZN(n23576) );
  NAND2_X2 U6079 ( .A1(n10126), .A2(n10127), .ZN(n6504) );
  NAND2_X2 U4373 ( .A1(n25142), .A2(n25184), .ZN(n25170) );
  INV_X4 U15083 ( .I(n13693), .ZN(n125) );
  NAND3_X2 U25336 ( .A1(n14973), .A2(n23785), .A3(n23903), .ZN(n23710) );
  AOI21_X2 U22375 ( .A1(n10700), .A2(n19115), .B(n25968), .ZN(n15143) );
  NAND2_X1 U12873 ( .A1(n16904), .A2(n17405), .ZN(n30064) );
  INV_X1 U12242 ( .I(n16904), .ZN(n29981) );
  NAND2_X2 U6760 ( .A1(n33761), .A2(n9427), .ZN(n9426) );
  NAND2_X2 U3799 ( .A1(n22364), .A2(n1125), .ZN(n3970) );
  NOR2_X2 U3349 ( .A1(n13796), .A2(n32253), .ZN(n29962) );
  INV_X2 U15551 ( .I(n17361), .ZN(n13950) );
  NOR2_X2 U10530 ( .A1(n10667), .A2(n10666), .ZN(n6490) );
  NOR2_X2 U7411 ( .A1(n29218), .A2(n30360), .ZN(n26241) );
  OAI22_X2 U16285 ( .A1(n5266), .A2(n18743), .B1(n18744), .B2(n18745), .ZN(
        n27261) );
  INV_X2 U869 ( .I(n575), .ZN(n1170) );
  NOR2_X2 U6762 ( .A1(n16432), .A2(n11930), .ZN(n1669) );
  INV_X2 U254 ( .I(n24308), .ZN(n27739) );
  AOI21_X2 U281 ( .A1(n24230), .A2(n24228), .B(n30696), .ZN(n30695) );
  INV_X2 U1191 ( .I(n21044), .ZN(n8284) );
  OAI21_X2 U10844 ( .A1(n6148), .A2(n26609), .B(n26608), .ZN(n26607) );
  AOI21_X2 U15376 ( .A1(n28900), .A2(n3487), .B(n28899), .ZN(n8285) );
  INV_X2 U3869 ( .I(n8084), .ZN(n27537) );
  NOR2_X2 U9191 ( .A1(n17288), .A2(n17287), .ZN(n17286) );
  INV_X2 U4878 ( .I(n32108), .ZN(n16403) );
  BUF_X4 U4448 ( .I(n25112), .Z(n25235) );
  INV_X2 U977 ( .I(n9737), .ZN(n31344) );
  INV_X4 U6479 ( .I(n12966), .ZN(n20427) );
  OAI21_X2 U1458 ( .A1(n11655), .A2(n27828), .B(n1331), .ZN(n30972) );
  INV_X4 U17361 ( .I(n11820), .ZN(n15964) );
  INV_X1 U48 ( .I(n10285), .ZN(n27164) );
  AOI21_X2 U12754 ( .A1(n6951), .A2(n32559), .B(n26827), .ZN(n6950) );
  INV_X2 U1904 ( .I(n19215), .ZN(n31503) );
  NAND2_X2 U1288 ( .A1(n15027), .A2(n20463), .ZN(n11035) );
  INV_X2 U19235 ( .I(n12866), .ZN(n21733) );
  NOR3_X2 U10119 ( .A1(n16358), .A2(n5269), .A3(n18705), .ZN(n10833) );
  NAND2_X2 U3671 ( .A1(n21579), .A2(n6669), .ZN(n21659) );
  INV_X1 U5990 ( .I(n16855), .ZN(n1183) );
  NAND2_X2 U7369 ( .A1(n17675), .A2(n9749), .ZN(n4639) );
  NOR2_X2 U8788 ( .A1(n5269), .A2(n18746), .ZN(n5266) );
  INV_X2 U6865 ( .I(n26415), .ZN(n23794) );
  NAND2_X1 U18021 ( .A1(n7067), .A2(n969), .ZN(n7069) );
  INV_X2 U6855 ( .I(n9153), .ZN(n10052) );
  INV_X4 U4808 ( .I(n11923), .ZN(n739) );
  NAND2_X2 U4669 ( .A1(n18983), .A2(n27021), .ZN(n18965) );
  INV_X2 U9972 ( .I(n19436), .ZN(n3417) );
  NOR2_X2 U15096 ( .A1(n7081), .A2(n25339), .ZN(n25233) );
  NAND2_X1 U12100 ( .A1(n18887), .A2(n10326), .ZN(n6362) );
  NAND2_X2 U11820 ( .A1(n12625), .A2(n31742), .ZN(n9728) );
  AOI21_X2 U5745 ( .A1(n7946), .A2(n29325), .B(n27589), .ZN(n7945) );
  OAI21_X2 U5909 ( .A1(n11832), .A2(n15052), .B(n14913), .ZN(n11831) );
  NAND2_X2 U1993 ( .A1(n19265), .A2(n18973), .ZN(n26469) );
  NAND2_X2 U2762 ( .A1(n24609), .A2(n28815), .ZN(n15232) );
  BUF_X2 U4982 ( .I(n19583), .Z(n27240) );
  BUF_X4 U2387 ( .I(n14002), .Z(n4135) );
  NAND3_X1 U2455 ( .A1(n16582), .A2(n16583), .A3(n7871), .ZN(n26877) );
  INV_X2 U2991 ( .I(n12561), .ZN(n919) );
  OR2_X1 U7098 ( .A1(n28904), .A2(n20545), .Z(n29356) );
  NOR2_X2 U3375 ( .A1(n23766), .A2(n23736), .ZN(n28637) );
  OR2_X2 U462 ( .A1(n5736), .A2(n9828), .Z(n29372) );
  NAND2_X2 U1104 ( .A1(n26573), .A2(n26513), .ZN(n31400) );
  OAI21_X1 U25118 ( .A1(n14251), .A2(n32830), .B(n22350), .ZN(n22650) );
  NAND2_X2 U6 ( .A1(n2962), .A2(n5839), .ZN(n25732) );
  AOI21_X2 U7766 ( .A1(n14491), .A2(n14703), .B(n28945), .ZN(n3257) );
  INV_X2 U3368 ( .I(n13862), .ZN(n1299) );
  INV_X1 U4430 ( .I(n18059), .ZN(n25227) );
  INV_X4 U6126 ( .I(n9561), .ZN(n14913) );
  BUF_X4 U6798 ( .I(n9107), .Z(n30365) );
  BUF_X2 U4281 ( .I(Key[157]), .Z(n16525) );
  BUF_X2 U4292 ( .I(Key[36]), .Z(n16497) );
  NAND2_X1 U18780 ( .A1(n16607), .A2(n25120), .ZN(n30673) );
  NAND2_X2 U370 ( .A1(n31531), .A2(n4124), .ZN(n2114) );
  INV_X4 U6558 ( .I(n15522), .ZN(n11745) );
  OAI21_X2 U3541 ( .A1(n14699), .A2(n14698), .B(n19245), .ZN(n14697) );
  NAND3_X2 U6203 ( .A1(n1057), .A2(n3928), .A3(n3927), .ZN(n5155) );
  INV_X2 U7331 ( .I(n20413), .ZN(n933) );
  INV_X2 U610 ( .I(n12878), .ZN(n13321) );
  INV_X2 U5973 ( .I(n18859), .ZN(n1057) );
  AOI21_X2 U2969 ( .A1(n16308), .A2(n14556), .B(n1022), .ZN(n20249) );
  NAND2_X2 U11643 ( .A1(n28899), .A2(n20362), .ZN(n20364) );
  INV_X2 U8355 ( .I(n599), .ZN(n21324) );
  OR2_X2 U15762 ( .A1(n23587), .A2(n23130), .Z(n8145) );
  AND2_X1 U4048 ( .A1(n17184), .A2(n17030), .Z(n18850) );
  NAND2_X2 U3258 ( .A1(n33909), .A2(n6961), .ZN(n9413) );
  NAND2_X2 U23948 ( .A1(n26573), .A2(n21687), .ZN(n12562) );
  NOR2_X2 U16155 ( .A1(n12320), .A2(n18581), .ZN(n30560) );
  INV_X4 U7043 ( .I(n7831), .ZN(n4525) );
  NOR2_X2 U8273 ( .A1(n8197), .A2(n154), .ZN(n15931) );
  OAI22_X2 U3438 ( .A1(n773), .A2(n9954), .B1(n22945), .B2(n850), .ZN(n26253)
         );
  NOR2_X1 U2133 ( .A1(n30619), .A2(n4220), .ZN(n12753) );
  INV_X2 U237 ( .I(n25890), .ZN(n7689) );
  NAND2_X2 U5090 ( .A1(n18078), .A2(n6679), .ZN(n1469) );
  INV_X2 U15596 ( .I(n21240), .ZN(n2239) );
  OAI21_X2 U25834 ( .A1(n17791), .A2(n20278), .B(n17790), .ZN(n28829) );
  NAND2_X2 U23973 ( .A1(n18169), .A2(n33312), .ZN(n18168) );
  NAND4_X2 U10497 ( .A1(n25768), .A2(n25770), .A3(n29168), .A4(n25769), .ZN(
        n26571) );
  NOR2_X2 U2442 ( .A1(n14752), .A2(n24915), .ZN(n24905) );
  INV_X4 U12077 ( .I(n8790), .ZN(n1009) );
  INV_X1 U15791 ( .I(n6969), .ZN(n6968) );
  BUF_X2 U3830 ( .I(n20423), .Z(n4647) );
  INV_X2 U11981 ( .I(n18960), .ZN(n18959) );
  INV_X2 U1121 ( .I(n32606), .ZN(n22608) );
  BUF_X2 U1989 ( .I(n2983), .Z(n42) );
  NOR2_X2 U5322 ( .A1(n9797), .A2(n11943), .ZN(n11078) );
  OAI21_X2 U1140 ( .A1(n27991), .A2(n21627), .B(n16601), .ZN(n28712) );
  NAND2_X2 U2964 ( .A1(n1287), .A2(n15644), .ZN(n30703) );
  OAI21_X2 U619 ( .A1(n17064), .A2(n11929), .B(n22830), .ZN(n18056) );
  NAND2_X2 U24244 ( .A1(n18472), .A2(n22), .ZN(n18389) );
  INV_X2 U2096 ( .I(n18696), .ZN(n12951) );
  INV_X2 U5806 ( .I(n10438), .ZN(n16306) );
  OAI21_X2 U24840 ( .A1(n21419), .A2(n4381), .B(n21117), .ZN(n21119) );
  BUF_X4 U3708 ( .I(n10974), .Z(n29047) );
  NAND2_X2 U21216 ( .A1(n14576), .A2(n14815), .ZN(n19966) );
  NAND2_X2 U7017 ( .A1(n680), .A2(n24610), .ZN(n3013) );
  INV_X2 U14 ( .I(n24927), .ZN(n24933) );
  INV_X2 U21764 ( .I(n18648), .ZN(n17114) );
  BUF_X2 U2366 ( .I(n18186), .Z(n10964) );
  NOR2_X2 U18311 ( .A1(n31428), .A2(n17477), .ZN(n18886) );
  OR2_X1 U4217 ( .A1(n6555), .A2(n14770), .Z(n9148) );
  INV_X2 U972 ( .I(n9789), .ZN(n10288) );
  NAND2_X2 U24634 ( .A1(n20025), .A2(n16461), .ZN(n20026) );
  OAI21_X2 U667 ( .A1(n22722), .A2(n22908), .B(n30447), .ZN(n22556) );
  INV_X2 U64 ( .I(n16751), .ZN(n16752) );
  INV_X2 U2273 ( .I(n4124), .ZN(n22720) );
  INV_X2 U4964 ( .I(n11900), .ZN(n25630) );
  NOR2_X2 U4755 ( .A1(n28704), .A2(n5433), .ZN(n19824) );
  AOI21_X2 U13447 ( .A1(n7767), .A2(n29819), .B(n30121), .ZN(n8114) );
  INV_X4 U2012 ( .I(n1060), .ZN(n31428) );
  INV_X2 U22052 ( .I(n19252), .ZN(n28276) );
  INV_X2 U23951 ( .I(n17559), .ZN(n19990) );
  INV_X2 U759 ( .I(n23086), .ZN(n28948) );
  NAND2_X1 U6654 ( .A1(n7319), .A2(n7318), .ZN(n2706) );
  INV_X4 U3382 ( .I(n8100), .ZN(n1172) );
  INV_X4 U5454 ( .I(n10845), .ZN(n1039) );
  INV_X2 U8396 ( .I(n10351), .ZN(n7719) );
  AOI21_X2 U8817 ( .A1(n18515), .A2(n11918), .B(n13663), .ZN(n9211) );
  OR2_X1 U4063 ( .A1(n22737), .A2(n2449), .Z(n23030) );
  NAND2_X2 U159 ( .A1(n9275), .A2(n24157), .ZN(n24206) );
  NAND3_X2 U3618 ( .A1(n32816), .A2(n21427), .A3(n33949), .ZN(n14618) );
  AOI21_X2 U5177 ( .A1(n19060), .A2(n9787), .B(n1374), .ZN(n2411) );
  NOR2_X2 U8730 ( .A1(n18363), .A2(n18161), .ZN(n18160) );
  NAND2_X2 U1741 ( .A1(n29208), .A2(n20043), .ZN(n11414) );
  NOR2_X2 U10126 ( .A1(n6470), .A2(n785), .ZN(n5122) );
  BUF_X4 U6257 ( .I(n6846), .Z(n5119) );
  OAI21_X1 U2188 ( .A1(n292), .A2(n12358), .B(n30019), .ZN(n24467) );
  NOR2_X2 U10177 ( .A1(n9305), .A2(n5225), .ZN(n9215) );
  INV_X2 U6340 ( .I(n8857), .ZN(n6748) );
  NOR2_X1 U14716 ( .A1(n6041), .A2(n6042), .ZN(n3996) );
  INV_X2 U13804 ( .I(n27007), .ZN(n22899) );
  OAI21_X2 U1725 ( .A1(n16675), .A2(n31745), .B(n29845), .ZN(n4209) );
  OR2_X2 U3435 ( .A1(n17306), .A2(n14911), .Z(n25887) );
  INV_X2 U4950 ( .I(n20630), .ZN(n20213) );
  OAI21_X2 U2625 ( .A1(n801), .A2(n31179), .B(n23640), .ZN(n29570) );
  NAND2_X2 U4224 ( .A1(n23956), .A2(n23824), .ZN(n18044) );
  NAND2_X2 U24872 ( .A1(n28869), .A2(n21430), .ZN(n21331) );
  NAND2_X2 U2072 ( .A1(n18618), .A2(n18779), .ZN(n30686) );
  BUF_X4 U15153 ( .I(n22871), .Z(n31861) );
  BUF_X2 U6098 ( .I(n18780), .Z(n31095) );
  NOR2_X2 U19953 ( .A1(n22339), .A2(n14145), .ZN(n22786) );
  OAI21_X2 U1477 ( .A1(n26554), .A2(n26553), .B(n25960), .ZN(n13705) );
  OAI22_X2 U8759 ( .A1(n18606), .A2(n18607), .B1(n18605), .B2(n18604), .ZN(
        n12768) );
  AOI21_X2 U10143 ( .A1(n18493), .A2(n5677), .B(n18324), .ZN(n15071) );
  AOI21_X2 U15790 ( .A1(n23082), .A2(n22885), .B(n13592), .ZN(n12450) );
  BUF_X2 U10828 ( .I(n23696), .Z(n8217) );
  NAND3_X2 U2484 ( .A1(n2715), .A2(n2716), .A3(n16473), .ZN(n2719) );
  NAND3_X2 U15767 ( .A1(n27103), .A2(n5757), .A3(n33571), .ZN(n21886) );
  INV_X4 U23588 ( .I(n17767), .ZN(n28502) );
  NAND2_X2 U5270 ( .A1(n29462), .A2(n12310), .ZN(n7839) );
  INV_X2 U3241 ( .I(n18983), .ZN(n17339) );
  OAI22_X2 U2798 ( .A1(n11299), .A2(n8453), .B1(n7430), .B2(n21328), .ZN(
        n21334) );
  NAND2_X2 U1681 ( .A1(n17688), .A2(n19901), .ZN(n20109) );
  NOR2_X2 U7614 ( .A1(n497), .A2(n18535), .ZN(n18704) );
  INV_X2 U8475 ( .I(n20633), .ZN(n2873) );
  NAND2_X1 U16674 ( .A1(n8955), .A2(n8958), .ZN(n27363) );
  NAND2_X2 U816 ( .A1(n6027), .A2(n20066), .ZN(n20094) );
  OAI22_X2 U4820 ( .A1(n25943), .A2(n11814), .B1(n12037), .B2(n21358), .ZN(
        n21359) );
  INV_X2 U19642 ( .I(n20120), .ZN(n20019) );
  INV_X1 U12950 ( .I(n7896), .ZN(n30075) );
  NOR2_X2 U7588 ( .A1(n1060), .A2(n18660), .ZN(n18887) );
  OAI21_X2 U15481 ( .A1(n1051), .A2(n18919), .B(n15534), .ZN(n4622) );
  NAND3_X2 U17232 ( .A1(n27814), .A2(n22981), .A3(n29329), .ZN(n30447) );
  BUF_X4 U1784 ( .I(n21006), .Z(n28262) );
  INV_X2 U175 ( .I(n9962), .ZN(n1246) );
  INV_X2 U20199 ( .I(n5226), .ZN(n24221) );
  NAND2_X2 U1227 ( .A1(n29676), .A2(n20392), .ZN(n28900) );
  INV_X4 U942 ( .I(n12585), .ZN(n1051) );
  OAI22_X2 U2833 ( .A1(n13913), .A2(n32951), .B1(n13219), .B2(n4210), .ZN(
        n13541) );
  NAND2_X1 U8138 ( .A1(n17734), .A2(n1132), .ZN(n11536) );
  OAI21_X2 U14017 ( .A1(n30181), .A2(n18292), .B(n18290), .ZN(n8482) );
  OAI21_X2 U12534 ( .A1(n30931), .A2(n17790), .B(n20562), .ZN(n3352) );
  INV_X2 U5649 ( .I(n17201), .ZN(n809) );
  INV_X2 U23 ( .I(n5942), .ZN(n6092) );
  NOR2_X2 U6646 ( .A1(n32005), .A2(n6597), .ZN(n6920) );
  INV_X2 U69 ( .I(n25437), .ZN(n11640) );
  OAI22_X2 U22948 ( .A1(n22817), .A2(n33968), .B1(n13597), .B2(n22818), .ZN(
        n22819) );
  OAI21_X2 U1537 ( .A1(n16011), .A2(n20359), .B(n30793), .ZN(n2319) );
  INV_X4 U6623 ( .I(n19220), .ZN(n9787) );
  NAND2_X2 U1868 ( .A1(n31161), .A2(n9563), .ZN(n11872) );
  INV_X2 U5709 ( .I(n548), .ZN(n15272) );
  INV_X2 U912 ( .I(n14760), .ZN(n1374) );
  NAND2_X2 U1069 ( .A1(n10456), .A2(n2300), .ZN(n2299) );
  INV_X2 U79 ( .I(n25378), .ZN(n750) );
  NOR2_X2 U20376 ( .A1(n8403), .A2(n8402), .ZN(n27972) );
  NAND2_X2 U6875 ( .A1(n6247), .A2(n893), .ZN(n11589) );
  OAI21_X2 U11866 ( .A1(n11971), .A2(n16307), .B(n8259), .ZN(n19929) );
  NAND2_X2 U1235 ( .A1(n1158), .A2(n20614), .ZN(n28603) );
  INV_X2 U2040 ( .I(n4734), .ZN(n22826) );
  OAI21_X2 U3448 ( .A1(n2923), .A2(n24057), .B(n27592), .ZN(n2922) );
  INV_X2 U2298 ( .I(n19849), .ZN(n9563) );
  INV_X2 U8584 ( .I(n11198), .ZN(n6970) );
  NOR2_X2 U6116 ( .A1(n33990), .A2(n2847), .ZN(n2851) );
  INV_X2 U9011 ( .I(n10183), .ZN(n10202) );
  INV_X4 U15564 ( .I(n23828), .ZN(n23669) );
  BUF_X2 U3188 ( .I(n7195), .Z(n31498) );
  OAI22_X2 U2858 ( .A1(n25113), .A2(n16632), .B1(n14895), .B2(n18132), .ZN(
        n27575) );
  INV_X2 U6285 ( .I(n22737), .ZN(n850) );
  INV_X1 U4835 ( .I(n21248), .ZN(n22521) );
  NAND2_X2 U5152 ( .A1(n12585), .A2(n25959), .ZN(n18958) );
  NOR2_X2 U14032 ( .A1(n32018), .A2(n28320), .ZN(n30182) );
  INV_X4 U2226 ( .I(n1931), .ZN(n16651) );
  INV_X2 U4378 ( .I(n14797), .ZN(n26608) );
  NOR2_X2 U660 ( .A1(n9377), .A2(n23017), .ZN(n14797) );
  NAND2_X2 U7461 ( .A1(n10453), .A2(n19050), .ZN(n10452) );
  INV_X2 U1050 ( .I(n21706), .ZN(n1316) );
  NAND2_X2 U25795 ( .A1(n28802), .A2(n3425), .ZN(n3424) );
  INV_X2 U8132 ( .I(n51), .ZN(n848) );
  INV_X2 U15119 ( .I(n9980), .ZN(n16933) );
  NOR2_X2 U4962 ( .A1(n13074), .A2(n34115), .ZN(n9615) );
  OAI22_X2 U10548 ( .A1(n4961), .A2(n26580), .B1(n4960), .B2(n15068), .ZN(
        n4959) );
  AOI21_X2 U15438 ( .A1(n7830), .A2(n33641), .B(n14563), .ZN(n7206) );
  NAND2_X2 U13433 ( .A1(n2514), .A2(n862), .ZN(n2513) );
  AOI21_X2 U16640 ( .A1(n18539), .A2(n18537), .B(n14651), .ZN(n5457) );
  NOR2_X2 U9115 ( .A1(n30724), .A2(n17604), .ZN(n30142) );
  INV_X2 U50 ( .I(n25901), .ZN(n7143) );
  NOR2_X2 U22526 ( .A1(n6298), .A2(n6666), .ZN(n31223) );
  INV_X2 U7000 ( .I(n17673), .ZN(n25403) );
  INV_X2 U5213 ( .I(n25479), .ZN(n25486) );
  NAND2_X2 U18060 ( .A1(n13407), .A2(n4381), .ZN(n7118) );
  NAND2_X2 U11455 ( .A1(n7206), .A2(n7205), .ZN(n7204) );
  INV_X2 U3329 ( .I(n10226), .ZN(n10513) );
  INV_X4 U13637 ( .I(n9133), .ZN(n10113) );
  AOI21_X2 U16375 ( .A1(n21580), .A2(n5795), .B(n3467), .ZN(n7349) );
  INV_X2 U880 ( .I(n17303), .ZN(n31506) );
  NAND2_X2 U8800 ( .A1(n34013), .A2(n4071), .ZN(n10105) );
  INV_X2 U687 ( .I(n6681), .ZN(n15874) );
  NAND2_X1 U10948 ( .A1(n24449), .A2(n1079), .ZN(n11696) );
  OAI21_X2 U8537 ( .A1(n8294), .A2(n8295), .B(n19863), .ZN(n2674) );
  NOR2_X2 U1297 ( .A1(n21705), .A2(n21704), .ZN(n21794) );
  INV_X4 U7188 ( .I(n21322), .ZN(n15015) );
  INV_X2 U582 ( .I(n28343), .ZN(n31810) );
  CLKBUF_X4 U9423 ( .I(n580), .Z(n29676) );
  INV_X2 U3544 ( .I(n31954), .ZN(n1007) );
  AOI21_X2 U324 ( .A1(n24263), .A2(n15974), .B(n1239), .ZN(n31785) );
  NOR2_X2 U7498 ( .A1(n10229), .A2(n33335), .ZN(n10857) );
  BUF_X4 U6299 ( .I(n20133), .Z(n16637) );
  AND2_X1 U4350 ( .A1(n29928), .A2(n11986), .Z(n7851) );
  NAND3_X2 U24657 ( .A1(n9688), .A2(n13920), .A3(n1154), .ZN(n20180) );
  INV_X2 U7025 ( .I(n25621), .ZN(n25752) );
  AOI22_X2 U11478 ( .A1(n1374), .A2(n29146), .B1(n31757), .B2(n16185), .ZN(
        n31213) );
  NAND2_X2 U20791 ( .A1(n22811), .A2(n22810), .ZN(n16028) );
  OAI21_X2 U6602 ( .A1(n11228), .A2(n7183), .B(n15595), .ZN(n31148) );
  INV_X2 U15127 ( .I(n19310), .ZN(n14178) );
  NAND2_X2 U10065 ( .A1(n10229), .A2(n25985), .ZN(n10352) );
  BUF_X2 U8016 ( .I(n15502), .Z(n31726) );
  NAND2_X2 U2408 ( .A1(n33146), .A2(n21721), .ZN(n21580) );
  INV_X2 U6571 ( .I(n17369), .ZN(n16081) );
  OAI22_X2 U1998 ( .A1(n18615), .A2(n31115), .B1(n18029), .B2(n16948), .ZN(
        n31459) );
  OAI22_X2 U13224 ( .A1(n1469), .A2(n20379), .B1(n2904), .B2(n2203), .ZN(
        n26907) );
  NAND2_X2 U1712 ( .A1(n2879), .A2(n868), .ZN(n31393) );
  NAND2_X2 U318 ( .A1(n10427), .A2(n9946), .ZN(n28488) );
  NOR2_X2 U3411 ( .A1(n27697), .A2(n20595), .ZN(n20258) );
  INV_X4 U10831 ( .I(n906), .ZN(n30641) );
  AOI22_X2 U26249 ( .A1(n4867), .A2(n24926), .B1(n24921), .B2(n15569), .ZN(
        n29127) );
  INV_X2 U4380 ( .I(n8622), .ZN(n13934) );
  OR2_X1 U11863 ( .A1(n8244), .A2(n2927), .Z(n2934) );
  NAND2_X2 U6249 ( .A1(n19267), .A2(n18974), .ZN(n13831) );
  NOR2_X2 U1977 ( .A1(n26417), .A2(n8141), .ZN(n19032) );
  NAND2_X2 U21417 ( .A1(n28130), .A2(n8137), .ZN(n29211) );
  INV_X2 U2050 ( .I(n27779), .ZN(n25169) );
  OAI21_X2 U2465 ( .A1(n3842), .A2(n1567), .B(n2909), .ZN(n27779) );
  NAND2_X2 U6787 ( .A1(n11268), .A2(n10031), .ZN(n27556) );
  AOI22_X2 U14331 ( .A1(n3407), .A2(n16694), .B1(n12061), .B2(n1360), .ZN(
        n15965) );
  NAND2_X2 U7360 ( .A1(n17456), .A2(n11350), .ZN(n11408) );
  AOI21_X2 U5993 ( .A1(n20125), .A2(n20124), .B(n20123), .ZN(n20126) );
  NAND2_X2 U6321 ( .A1(n1926), .A2(n17891), .ZN(n17890) );
  INV_X2 U21763 ( .I(n18392), .ZN(n15888) );
  BUF_X2 U24 ( .I(n17927), .Z(n29085) );
  OAI21_X1 U1762 ( .A1(n14426), .A2(n33069), .B(n8193), .ZN(n14425) );
  NAND2_X2 U7396 ( .A1(n19993), .A2(n1040), .ZN(n2288) );
  BUF_X2 U4161 ( .I(n17261), .Z(n28436) );
  NOR2_X2 U482 ( .A1(n4991), .A2(n23828), .ZN(n13196) );
  AOI21_X2 U20913 ( .A1(n14864), .A2(n21877), .B(n28059), .ZN(n15315) );
  INV_X4 U694 ( .I(n21070), .ZN(n21430) );
  NOR2_X2 U7543 ( .A1(n5456), .A2(n1185), .ZN(n6793) );
  NOR2_X2 U6567 ( .A1(n21583), .A2(n21781), .ZN(n8164) );
  AOI22_X2 U2089 ( .A1(n21711), .A2(n727), .B1(n862), .B2(n21710), .ZN(n6514)
         );
  NAND2_X2 U10422 ( .A1(n24224), .A2(n10687), .ZN(n28467) );
  INV_X2 U1511 ( .I(n3351), .ZN(n20789) );
  BUF_X4 U5430 ( .I(n2566), .Z(n2565) );
  NAND2_X2 U8407 ( .A1(n20486), .A2(n20485), .ZN(n20252) );
  OAI21_X2 U6476 ( .A1(n11445), .A2(n10848), .B(n10074), .ZN(n30552) );
  INV_X2 U14925 ( .I(n11676), .ZN(n30359) );
  NOR2_X2 U2368 ( .A1(n15371), .A2(n7868), .ZN(n17354) );
  CLKBUF_X4 U1495 ( .I(n16239), .Z(n5822) );
  NAND2_X2 U3041 ( .A1(n8219), .A2(n561), .ZN(n9612) );
  NAND3_X2 U6530 ( .A1(n27715), .A2(n17711), .A3(n11264), .ZN(n10152) );
  OAI21_X2 U1739 ( .A1(n27541), .A2(n27542), .B(n15110), .ZN(n31173) );
  NOR2_X2 U2002 ( .A1(n15789), .A2(n13554), .ZN(n30648) );
  NOR2_X2 U2505 ( .A1(n27), .A2(n23691), .ZN(n28688) );
  INV_X2 U5114 ( .I(n6556), .ZN(n17640) );
  NAND2_X2 U1369 ( .A1(n27715), .A2(n19947), .ZN(n27714) );
  INV_X2 U7427 ( .I(n5433), .ZN(n10444) );
  NAND2_X2 U3262 ( .A1(n26158), .A2(n26157), .ZN(n24063) );
  INV_X4 U4172 ( .I(n14849), .ZN(n1137) );
  AOI21_X2 U9497 ( .A1(n32079), .A2(n14848), .B(n33842), .ZN(n6698) );
  INV_X1 U15611 ( .I(n32647), .ZN(n21413) );
  BUF_X4 U5007 ( .I(n19122), .Z(n15534) );
  INV_X4 U45 ( .I(n25276), .ZN(n25278) );
  AOI22_X2 U2576 ( .A1(n22837), .A2(n10360), .B1(n22835), .B2(n22836), .ZN(
        n4231) );
  INV_X2 U18297 ( .I(n19484), .ZN(n27607) );
  INV_X4 U17842 ( .I(n3748), .ZN(n16443) );
  NOR2_X2 U2468 ( .A1(n3085), .A2(n384), .ZN(n11105) );
  INV_X2 U1723 ( .I(n20335), .ZN(n20546) );
  BUF_X2 U6943 ( .I(n5317), .Z(n29866) );
  AOI22_X2 U15945 ( .A1(n6770), .A2(n24191), .B1(n28726), .B2(n6769), .ZN(
        n6768) );
  AOI21_X2 U4557 ( .A1(n1155), .A2(n33721), .B(n32941), .ZN(n29692) );
  BUF_X4 U4261 ( .I(n13719), .Z(n13663) );
  OAI21_X2 U9493 ( .A1(n16953), .A2(n16952), .B(n18079), .ZN(n7703) );
  NAND2_X2 U10706 ( .A1(n15272), .A2(n23638), .ZN(n8799) );
  INV_X2 U1525 ( .I(n20670), .ZN(n21046) );
  INV_X4 U6500 ( .I(n20607), .ZN(n15217) );
  NAND3_X2 U17368 ( .A1(n17808), .A2(n29603), .A3(n17809), .ZN(n15745) );
  AOI21_X2 U1980 ( .A1(n16485), .A2(n13685), .B(n947), .ZN(n9078) );
  INV_X2 U1421 ( .I(n17711), .ZN(n942) );
  OAI21_X2 U2933 ( .A1(n33097), .A2(n1098), .B(n4538), .ZN(n17923) );
  AND2_X1 U7094 ( .A1(n13936), .A2(n31650), .Z(n29353) );
  BUF_X2 U5028 ( .I(n23683), .Z(n23864) );
  BUF_X4 U6974 ( .I(n24180), .Z(n5913) );
  NOR2_X1 U15167 ( .A1(n2069), .A2(n9788), .ZN(n28700) );
  BUF_X4 U12883 ( .I(n14339), .Z(n30065) );
  NAND2_X2 U15671 ( .A1(n6962), .A2(n4373), .ZN(n13583) );
  BUF_X4 U973 ( .I(n22411), .Z(n31551) );
  INV_X2 U502 ( .I(n23770), .ZN(n27910) );
  INV_X2 U599 ( .I(n23508), .ZN(n1259) );
  INV_X2 U871 ( .I(n9370), .ZN(n29232) );
  NOR2_X2 U19191 ( .A1(n14027), .A2(n8582), .ZN(n13572) );
  NAND2_X2 U425 ( .A1(n12817), .A2(n23752), .ZN(n12816) );
  BUF_X2 U74 ( .I(n25490), .Z(n4183) );
  OAI21_X2 U3547 ( .A1(n20594), .A2(n29603), .B(n20599), .ZN(n31401) );
  NAND2_X2 U6443 ( .A1(n27697), .A2(n27070), .ZN(n20599) );
  NAND2_X2 U1276 ( .A1(n28379), .A2(n744), .ZN(n19136) );
  INV_X2 U1103 ( .I(n30506), .ZN(n1326) );
  NOR2_X2 U14412 ( .A1(n19122), .A2(n30879), .ZN(n26550) );
  OAI21_X2 U224 ( .A1(n1634), .A2(n8004), .B(n4458), .ZN(n8003) );
  AOI22_X2 U15426 ( .A1(n1820), .A2(n992), .B1(n17394), .B2(n22583), .ZN(n1486) );
  NAND3_X2 U17000 ( .A1(n161), .A2(n1036), .A3(n27345), .ZN(n3272) );
  INV_X2 U5271 ( .I(n12310), .ZN(n5135) );
  NAND2_X2 U15075 ( .A1(n24057), .A2(n31918), .ZN(n24496) );
  AOI21_X2 U24626 ( .A1(n26567), .A2(n28471), .B(n741), .ZN(n20001) );
  NOR2_X2 U2425 ( .A1(n14384), .A2(n32384), .ZN(n11644) );
  NAND2_X2 U3175 ( .A1(n12715), .A2(n23318), .ZN(n3281) );
  INV_X4 U20445 ( .I(n29335), .ZN(n15322) );
  AND2_X1 U5109 ( .A1(n23692), .A2(n13147), .Z(n31239) );
  INV_X2 U5453 ( .I(n17405), .ZN(n19819) );
  NAND2_X1 U11065 ( .A1(n9030), .A2(n9032), .ZN(n30119) );
  OAI21_X2 U4623 ( .A1(n14461), .A2(n1316), .B(n21613), .ZN(n6253) );
  BUF_X2 U372 ( .I(n8178), .Z(n29977) );
  INV_X2 U9471 ( .I(n29854), .ZN(n26474) );
  INV_X1 U19205 ( .I(n30731), .ZN(n6257) );
  NAND2_X2 U15476 ( .A1(n786), .A2(n10858), .ZN(n10574) );
  NAND2_X2 U3150 ( .A1(n20155), .A2(n10059), .ZN(n2089) );
  NOR2_X2 U776 ( .A1(n28101), .A2(n29957), .ZN(n28035) );
  NOR2_X2 U8748 ( .A1(n15018), .A2(n1185), .ZN(n18161) );
  NAND2_X2 U2602 ( .A1(n15682), .A2(n23860), .ZN(n11158) );
  INV_X4 U19615 ( .I(n9390), .ZN(n15394) );
  NOR2_X2 U3695 ( .A1(n18617), .A2(n18616), .ZN(n16418) );
  INV_X2 U4377 ( .I(n25007), .ZN(n1205) );
  NAND2_X2 U12141 ( .A1(n11270), .A2(n33039), .ZN(n10247) );
  INV_X2 U26161 ( .I(n24785), .ZN(n1085) );
  NAND2_X2 U1479 ( .A1(n31004), .A2(n9439), .ZN(n31003) );
  INV_X1 U8086 ( .I(n16306), .ZN(n22621) );
  INV_X4 U13175 ( .I(n2256), .ZN(n22780) );
  NAND2_X2 U147 ( .A1(n18154), .A2(n25114), .ZN(n16024) );
  INV_X1 U480 ( .I(n2021), .ZN(n14497) );
  INV_X4 U2648 ( .I(n33069), .ZN(n19181) );
  INV_X2 U3895 ( .I(n27931), .ZN(n5335) );
  NAND3_X2 U8724 ( .A1(n22624), .A2(n22623), .A3(n2538), .ZN(n26393) );
  INV_X2 U5388 ( .I(n22098), .ZN(n22260) );
  INV_X2 U19442 ( .I(n22072), .ZN(n27837) );
  INV_X2 U8085 ( .I(n2547), .ZN(n994) );
  INV_X4 U439 ( .I(n22534), .ZN(n1120) );
  BUF_X4 U3579 ( .I(n5625), .Z(n4643) );
  INV_X2 U5524 ( .I(n7195), .ZN(n927) );
  BUF_X4 U3894 ( .I(n17967), .Z(n27345) );
  INV_X2 U1493 ( .I(n12804), .ZN(n21223) );
  INV_X2 U17223 ( .I(n16011), .ZN(n27426) );
  OAI21_X2 U10129 ( .A1(n9215), .A2(n18518), .B(n18672), .ZN(n9304) );
  INV_X2 U1419 ( .I(n21109), .ZN(n17438) );
  INV_X4 U5979 ( .I(n14454), .ZN(n3080) );
  BUF_X2 U1542 ( .I(n19289), .Z(n28528) );
  NOR2_X2 U6599 ( .A1(n19357), .A2(n19229), .ZN(n19354) );
  NOR2_X2 U5139 ( .A1(n5962), .A2(n28825), .ZN(n29928) );
  AOI21_X2 U8258 ( .A1(n15220), .A2(n15219), .B(n32799), .ZN(n15358) );
  AOI21_X2 U15782 ( .A1(n4371), .A2(n10947), .B(n13747), .ZN(n4370) );
  INV_X2 U4607 ( .I(n19947), .ZN(n11264) );
  BUF_X2 U2938 ( .I(n26363), .Z(n31072) );
  NAND2_X2 U13167 ( .A1(n28528), .A2(n10124), .ZN(n19076) );
  OAI21_X1 U3010 ( .A1(n23688), .A2(n17181), .B(n25987), .ZN(n23689) );
  BUF_X2 U1034 ( .I(n4034), .Z(n27850) );
  NAND2_X2 U834 ( .A1(n11161), .A2(n22669), .ZN(n2311) );
  OR2_X1 U4196 ( .A1(n24466), .A2(n292), .Z(n26281) );
  NOR2_X2 U15271 ( .A1(n776), .A2(n14686), .ZN(n28071) );
  NAND2_X2 U15622 ( .A1(n2577), .A2(n347), .ZN(n30291) );
  BUF_X4 U4752 ( .I(n596), .Z(n28287) );
  INV_X2 U21006 ( .I(n19637), .ZN(n15063) );
  INV_X4 U2639 ( .I(n17895), .ZN(n844) );
  NOR2_X2 U6995 ( .A1(n24973), .A2(n17118), .ZN(n17782) );
  AOI21_X2 U2513 ( .A1(n10589), .A2(n22919), .B(n10588), .ZN(n10760) );
  INV_X4 U7426 ( .I(n12168), .ZN(n8927) );
  NOR2_X2 U656 ( .A1(n28314), .A2(n3614), .ZN(n12728) );
  BUF_X2 U7069 ( .I(Key[177]), .Z(n25436) );
  INV_X2 U6929 ( .I(n23109), .ZN(n1264) );
  OR2_X1 U3623 ( .A1(n19915), .A2(n31671), .Z(n28208) );
  NOR2_X2 U22197 ( .A1(n818), .A2(n20411), .ZN(n28268) );
  OAI21_X2 U17087 ( .A1(n18953), .A2(n18952), .B(n28935), .ZN(n11336) );
  NAND2_X2 U4516 ( .A1(n20468), .A2(n14138), .ZN(n6536) );
  NAND2_X2 U8029 ( .A1(n27737), .A2(n30066), .ZN(n15919) );
  NAND2_X2 U6780 ( .A1(n12952), .A2(n16432), .ZN(n27737) );
  NAND2_X1 U10699 ( .A1(n14497), .A2(n14496), .ZN(n2036) );
  NAND2_X2 U18957 ( .A1(n19927), .A2(n30554), .ZN(n19928) );
  OAI21_X2 U9877 ( .A1(n6970), .A2(n19926), .B(n13591), .ZN(n19927) );
  BUF_X2 U4317 ( .I(Key[47]), .Z(n25195) );
  INV_X2 U6807 ( .I(n24243), .ZN(n24337) );
  CLKBUF_X2 U10231 ( .I(Key[159]), .Z(n25881) );
  NAND2_X1 U7842 ( .A1(n12020), .A2(n313), .ZN(n12858) );
  NAND2_X2 U2907 ( .A1(n20335), .A2(n30130), .ZN(n20411) );
  NAND2_X2 U2062 ( .A1(n489), .A2(n4194), .ZN(n17321) );
  NOR2_X2 U13793 ( .A1(n15434), .A2(n2843), .ZN(n17993) );
  INV_X4 U10085 ( .I(n29146), .ZN(n1179) );
  NAND2_X2 U4762 ( .A1(n24167), .A2(n24279), .ZN(n11121) );
  NOR2_X2 U7848 ( .A1(n23778), .A2(n23775), .ZN(n5438) );
  INV_X2 U6295 ( .I(n19406), .ZN(n31755) );
  INV_X2 U18497 ( .I(n14138), .ZN(n742) );
  NAND2_X2 U5298 ( .A1(n20059), .A2(n224), .ZN(n12696) );
  INV_X4 U21970 ( .I(n12707), .ZN(n13210) );
  NOR2_X1 U1238 ( .A1(n12354), .A2(n12394), .ZN(n30619) );
  INV_X2 U1157 ( .I(n21743), .ZN(n31654) );
  INV_X2 U689 ( .I(n16129), .ZN(n16906) );
  BUF_X2 U2145 ( .I(n12707), .Z(n12249) );
  AND2_X2 U3034 ( .A1(n26114), .A2(n10772), .Z(n23809) );
  OR2_X2 U2975 ( .A1(n5975), .A2(n625), .Z(n22364) );
  INV_X2 U14485 ( .I(n10390), .ZN(n4568) );
  AOI22_X2 U13486 ( .A1(n34005), .A2(n30932), .B1(n13475), .B2(n29715), .ZN(
        n15486) );
  NAND2_X2 U1558 ( .A1(n8689), .A2(n17234), .ZN(n32) );
  INV_X1 U1163 ( .I(n6842), .ZN(n21075) );
  OAI21_X2 U14037 ( .A1(n13428), .A2(n24780), .B(n3080), .ZN(n3079) );
  OAI21_X1 U9144 ( .A1(n29743), .A2(n12654), .B(n29742), .ZN(n7207) );
  NAND3_X2 U25183 ( .A1(n27589), .A2(n13778), .A3(n6149), .ZN(n23021) );
  OAI21_X2 U845 ( .A1(n28902), .A2(n22280), .B(n22379), .ZN(n261) );
  NAND2_X2 U6376 ( .A1(n20089), .A2(n2229), .ZN(n11120) );
  OR2_X1 U12927 ( .A1(n23805), .A2(n2752), .Z(n2004) );
  OAI21_X2 U2181 ( .A1(n2945), .A2(n13268), .B(n2943), .ZN(n15303) );
  INV_X4 U3750 ( .I(n14392), .ZN(n4113) );
  NAND3_X2 U5417 ( .A1(n33301), .A2(n13300), .A3(n20310), .ZN(n13563) );
  INV_X4 U6914 ( .I(n29785), .ZN(n24213) );
  OR2_X1 U4420 ( .A1(n32903), .A2(n16144), .Z(n2675) );
  INV_X2 U5718 ( .I(n10193), .ZN(n1098) );
  NAND3_X1 U15562 ( .A1(n23616), .A2(n33260), .A3(n23828), .ZN(n9998) );
  INV_X4 U13954 ( .I(n3601), .ZN(n18893) );
  INV_X2 U9950 ( .I(n17456), .ZN(n16579) );
  NOR2_X2 U2131 ( .A1(n15246), .A2(n15247), .ZN(n13302) );
  INV_X4 U2083 ( .I(n2019), .ZN(n29658) );
  BUF_X2 U7336 ( .I(n12375), .Z(n6553) );
  NOR2_X2 U2683 ( .A1(n10264), .A2(n959), .ZN(n8309) );
  INV_X2 U674 ( .I(n8490), .ZN(n11215) );
  NAND2_X2 U4586 ( .A1(n12836), .A2(n34054), .ZN(n6014) );
  BUF_X4 U2718 ( .I(n10657), .Z(n7007) );
  NAND3_X2 U1893 ( .A1(n26288), .A2(n29118), .A3(n19256), .ZN(n18526) );
  INV_X2 U755 ( .I(n33007), .ZN(n13474) );
  NAND3_X2 U14915 ( .A1(n14106), .A2(n14107), .A3(n9221), .ZN(n20503) );
  NAND2_X2 U18411 ( .A1(n19457), .A2(n33631), .ZN(n7708) );
  NAND2_X2 U3931 ( .A1(n33007), .A2(n33115), .ZN(n30364) );
  AOI21_X2 U15166 ( .A1(n24191), .A2(n795), .B(n28726), .ZN(n24172) );
  NOR2_X2 U2326 ( .A1(n27678), .A2(n1257), .ZN(n23308) );
  NOR2_X2 U6771 ( .A1(n22664), .A2(n22576), .ZN(n22454) );
  INV_X2 U10367 ( .I(n25513), .ZN(n1204) );
  INV_X4 U1532 ( .I(n13160), .ZN(n19137) );
  INV_X4 U974 ( .I(n22640), .ZN(n29626) );
  INV_X1 U4107 ( .I(n10673), .ZN(n23782) );
  INV_X4 U2350 ( .I(n12039), .ZN(n1213) );
  AOI21_X2 U15575 ( .A1(n16443), .A2(n24148), .B(n9946), .ZN(n8962) );
  NAND2_X2 U10964 ( .A1(n22843), .A2(n28330), .ZN(n5680) );
  INV_X2 U1833 ( .I(n31408), .ZN(n19969) );
  NOR2_X2 U25333 ( .A1(n1257), .A2(n10142), .ZN(n23698) );
  BUF_X2 U2610 ( .I(n25115), .Z(n14495) );
  INV_X2 U710 ( .I(n16315), .ZN(n15852) );
  NAND2_X2 U448 ( .A1(n18098), .A2(n27122), .ZN(n9620) );
  BUF_X4 U2775 ( .I(n24680), .Z(n25561) );
  INV_X2 U470 ( .I(n34125), .ZN(n1287) );
  AND2_X1 U16260 ( .A1(n5035), .A2(n987), .Z(n22509) );
  INV_X2 U854 ( .I(n502), .ZN(n13061) );
  NAND2_X2 U20478 ( .A1(n7792), .A2(n33403), .ZN(n30924) );
  OR2_X2 U13010 ( .A1(n18146), .A2(n24031), .Z(n24143) );
  OAI21_X2 U15492 ( .A1(n16443), .A2(n5335), .B(n29655), .ZN(n9521) );
  BUF_X4 U15043 ( .I(n25409), .Z(n419) );
  NAND2_X2 U289 ( .A1(n9824), .A2(n9823), .ZN(n9825) );
  NOR2_X2 U566 ( .A1(n8525), .A2(n23819), .ZN(n10749) );
  NOR2_X2 U20909 ( .A1(n21410), .A2(n16473), .ZN(n2941) );
  OAI21_X2 U2255 ( .A1(n24067), .A2(n32036), .B(n7503), .ZN(n10827) );
  BUF_X4 U248 ( .I(n6911), .Z(n27501) );
  AOI21_X2 U7250 ( .A1(n20566), .A2(n16515), .B(n12263), .ZN(n8941) );
  INV_X2 U7371 ( .I(n19601), .ZN(n13591) );
  INV_X2 U20282 ( .I(n27958), .ZN(n489) );
  INV_X2 U4181 ( .I(n16077), .ZN(n709) );
  OAI21_X2 U3851 ( .A1(n9261), .A2(n9262), .B(n29269), .ZN(n27756) );
  NAND2_X2 U25014 ( .A1(n621), .A2(n22557), .ZN(n22071) );
  BUF_X2 U4289 ( .I(Key[43]), .Z(n25190) );
  INV_X2 U16549 ( .I(n19969), .ZN(n30612) );
  INV_X2 U10864 ( .I(n13814), .ZN(n17188) );
  INV_X4 U12011 ( .I(n11940), .ZN(n29963) );
  AOI21_X2 U1909 ( .A1(n880), .A2(n879), .B(n15396), .ZN(n15395) );
  AND2_X2 U15465 ( .A1(n29124), .A2(n14587), .Z(n27159) );
  AOI21_X2 U2641 ( .A1(n22438), .A2(n12236), .B(n17007), .ZN(n17006) );
  NAND3_X2 U2616 ( .A1(n26459), .A2(n33544), .A3(n30459), .ZN(n14371) );
  INV_X2 U21563 ( .I(n19844), .ZN(n19923) );
  OR2_X2 U8316 ( .A1(n34151), .A2(n30387), .Z(n19888) );
  INV_X2 U5868 ( .I(n20519), .ZN(n20517) );
  NOR2_X2 U9048 ( .A1(n15665), .A2(n20056), .ZN(n17573) );
  NAND2_X2 U5448 ( .A1(n12398), .A2(n71), .ZN(n6405) );
  INV_X2 U14931 ( .I(n13040), .ZN(n28726) );
  INV_X2 U7640 ( .I(n14159), .ZN(n18853) );
  NAND3_X1 U2541 ( .A1(n5217), .A2(n26587), .A3(n14280), .ZN(n5216) );
  NOR2_X2 U3592 ( .A1(n7218), .A2(n8770), .ZN(n20304) );
  NAND2_X2 U4723 ( .A1(n20150), .A2(n20152), .ZN(n19915) );
  INV_X1 U5111 ( .I(n17590), .ZN(n21373) );
  INV_X2 U5914 ( .I(n29688), .ZN(n820) );
  NAND2_X2 U6151 ( .A1(n18496), .A2(n10043), .ZN(n8824) );
  INV_X1 U12195 ( .I(n24527), .ZN(n16253) );
  INV_X4 U1519 ( .I(n31970), .ZN(n763) );
  NOR2_X2 U2980 ( .A1(n25980), .A2(n397), .ZN(n8775) );
  NAND2_X1 U12914 ( .A1(n26858), .A2(n26856), .ZN(n21956) );
  BUF_X2 U6319 ( .I(n12452), .Z(n28923) );
  NAND2_X2 U2688 ( .A1(n18159), .A2(n29070), .ZN(n17873) );
  NAND2_X2 U18708 ( .A1(n10142), .A2(n33216), .ZN(n27679) );
  INV_X2 U14996 ( .I(n17717), .ZN(n11556) );
  INV_X2 U5754 ( .I(n23695), .ZN(n27163) );
  NAND2_X2 U16071 ( .A1(n26900), .A2(n27457), .ZN(n2221) );
  INV_X2 U3089 ( .I(n13670), .ZN(n28017) );
  OAI21_X2 U3844 ( .A1(n5745), .A2(n14119), .B(n8273), .ZN(n27377) );
  NOR2_X2 U7927 ( .A1(n17739), .A2(n32500), .ZN(n2222) );
  INV_X2 U274 ( .I(n29323), .ZN(n8273) );
  INV_X2 U7525 ( .I(n18988), .ZN(n19087) );
  NAND2_X2 U5617 ( .A1(n5135), .A2(n5380), .ZN(n30008) );
  INV_X1 U2086 ( .I(n18677), .ZN(n30558) );
  NAND2_X2 U2095 ( .A1(n15371), .A2(n31511), .ZN(n28973) );
  NAND2_X2 U12155 ( .A1(n18495), .A2(n28987), .ZN(n6026) );
  INV_X2 U5994 ( .I(n18847), .ZN(n18731) );
  OAI21_X2 U18265 ( .A1(n16461), .A2(n1042), .B(n6109), .ZN(n6108) );
  NAND2_X2 U4802 ( .A1(n2713), .A2(n7004), .ZN(n22838) );
  NOR2_X1 U535 ( .A1(n8082), .A2(n26780), .ZN(n8081) );
  NOR2_X2 U20256 ( .A1(n16189), .A2(n10686), .ZN(n15154) );
  INV_X4 U2818 ( .I(n563), .ZN(n11961) );
  BUF_X2 U5961 ( .I(n20445), .Z(n31768) );
  INV_X4 U2287 ( .I(n4373), .ZN(n5966) );
  NAND2_X2 U1669 ( .A1(n13341), .A2(n6098), .ZN(n13340) );
  NOR2_X2 U4976 ( .A1(n53), .A2(n7280), .ZN(n16882) );
  NAND3_X2 U17887 ( .A1(n26333), .A2(n9579), .A3(n16432), .ZN(n31689) );
  AOI22_X1 U7993 ( .A1(n17184), .A2(n18593), .B1(n18594), .B2(n18849), .ZN(
        n18598) );
  NAND2_X2 U25251 ( .A1(n9275), .A2(n32349), .ZN(n31543) );
  CLKBUF_X12 U2192 ( .I(n2956), .Z(n29011) );
  NOR2_X2 U3792 ( .A1(n23017), .A2(n23018), .ZN(n12416) );
  INV_X2 U16079 ( .I(n10420), .ZN(n25890) );
  INV_X4 U6200 ( .I(n23807), .ZN(n14664) );
  AOI22_X2 U5148 ( .A1(n10732), .A2(n16906), .B1(n21212), .B2(n21211), .ZN(
        n29503) );
  INV_X2 U7134 ( .I(n21721), .ZN(n1133) );
  NAND3_X2 U539 ( .A1(n187), .A2(n17773), .A3(n185), .ZN(n15677) );
  INV_X2 U11795 ( .I(n11408), .ZN(n3407) );
  NAND2_X2 U1524 ( .A1(n18913), .A2(n7995), .ZN(n19100) );
  BUF_X4 U5991 ( .I(n16855), .Z(n6597) );
  AOI21_X2 U22960 ( .A1(n16132), .A2(n1150), .B(n14710), .ZN(n20416) );
  OAI21_X2 U7550 ( .A1(n9090), .A2(n18633), .B(n18711), .ZN(n2987) );
  OAI21_X2 U5432 ( .A1(n215), .A2(n33763), .B(n214), .ZN(n23623) );
  NAND2_X1 U18436 ( .A1(n12391), .A2(n12392), .ZN(n30623) );
  CLKBUF_X4 U4855 ( .I(n20467), .Z(n26567) );
  INV_X2 U14940 ( .I(n11705), .ZN(n25348) );
  NAND2_X2 U10967 ( .A1(n22843), .A2(n33016), .ZN(n11467) );
  OAI21_X2 U15097 ( .A1(n1243), .A2(n23991), .B(n23990), .ZN(n23992) );
  AOI22_X2 U3338 ( .A1(n10853), .A2(n33822), .B1(n10857), .B2(n25985), .ZN(
        n31406) );
  INV_X4 U927 ( .I(n13295), .ZN(n19229) );
  NAND2_X2 U15784 ( .A1(n26544), .A2(n12143), .ZN(n31421) );
  OAI21_X2 U24134 ( .A1(n18226), .A2(n18848), .B(n18849), .ZN(n18224) );
  AOI21_X1 U3176 ( .A1(n12781), .A2(n12099), .B(n23318), .ZN(n12716) );
  NOR2_X1 U3419 ( .A1(n401), .A2(n8573), .ZN(n9123) );
  INV_X2 U1547 ( .I(n11103), .ZN(n30882) );
  INV_X2 U16111 ( .I(n10291), .ZN(n8270) );
  NOR2_X2 U11093 ( .A1(n30375), .A2(n19724), .ZN(n2927) );
  INV_X4 U6525 ( .I(n21237), .ZN(n21453) );
  NAND2_X1 U11283 ( .A1(n27317), .A2(n27316), .ZN(n30454) );
  NAND2_X2 U2807 ( .A1(n15833), .A2(n29938), .ZN(n15832) );
  NOR2_X2 U141 ( .A1(n10178), .A2(n10177), .ZN(n10176) );
  OAI22_X2 U26133 ( .A1(n29035), .A2(n29034), .B1(n6580), .B2(n729), .ZN(
        n11493) );
  NAND2_X2 U6393 ( .A1(n6611), .A2(n11624), .ZN(n13021) );
  NAND2_X2 U15117 ( .A1(n13037), .A2(n13035), .ZN(n19319) );
  OAI21_X2 U4376 ( .A1(n15189), .A2(n20155), .B(n11959), .ZN(n27111) );
  INV_X2 U2812 ( .I(n13510), .ZN(n16346) );
  NAND3_X2 U1665 ( .A1(n29365), .A2(n17672), .A3(n14731), .ZN(n30938) );
  NAND2_X2 U7114 ( .A1(n21632), .A2(n21871), .ZN(n4689) );
  INV_X4 U11935 ( .I(n6344), .ZN(n3989) );
  OR2_X2 U13567 ( .A1(n25695), .A2(n25628), .Z(n13641) );
  NOR2_X1 U21245 ( .A1(n28098), .A2(n18194), .ZN(n18192) );
  INV_X2 U598 ( .I(n21849), .ZN(n21763) );
  BUF_X4 U6353 ( .I(n31922), .Z(n16461) );
  INV_X1 U17036 ( .I(n2655), .ZN(n27378) );
  NAND2_X1 U2135 ( .A1(n12441), .A2(n7063), .ZN(n30562) );
  NAND2_X2 U21030 ( .A1(n32940), .A2(n295), .ZN(n15344) );
  OR2_X2 U12508 ( .A1(n13941), .A2(n1696), .Z(n19450) );
  OR2_X2 U17412 ( .A1(n30282), .A2(n6394), .Z(n4675) );
  AOI21_X2 U1752 ( .A1(n15383), .A2(n20066), .B(n30771), .ZN(n17346) );
  NOR2_X2 U2600 ( .A1(n15682), .A2(n23860), .ZN(n15681) );
  NOR2_X2 U17076 ( .A1(n27387), .A2(n13045), .ZN(n13043) );
  NOR2_X2 U17077 ( .A1(n15364), .A2(n3891), .ZN(n27387) );
  INV_X4 U11396 ( .I(n21630), .ZN(n2217) );
  NOR2_X2 U1956 ( .A1(n9345), .A2(n9344), .ZN(n9343) );
  NAND2_X2 U6237 ( .A1(n18767), .A2(n4624), .ZN(n17905) );
  NOR2_X1 U4616 ( .A1(n28494), .A2(n11938), .ZN(n12787) );
  NOR2_X1 U19587 ( .A1(n14264), .A2(n14261), .ZN(n30798) );
  NOR2_X2 U2617 ( .A1(n6599), .A2(n914), .ZN(n11797) );
  INV_X2 U1538 ( .I(n17586), .ZN(n17004) );
  INV_X2 U3754 ( .I(n18575), .ZN(n10043) );
  NOR2_X2 U25902 ( .A1(n19063), .A2(n19108), .ZN(n19110) );
  OR2_X1 U3779 ( .A1(n20219), .A2(n9014), .Z(n583) );
  INV_X4 U12728 ( .I(n1835), .ZN(n18633) );
  BUF_X2 U4883 ( .I(n9220), .Z(n7779) );
  NAND3_X2 U9693 ( .A1(n26499), .A2(n22828), .A3(n28327), .ZN(n26501) );
  NAND2_X2 U17097 ( .A1(n6082), .A2(n12654), .ZN(n14560) );
  INV_X2 U1324 ( .I(n18187), .ZN(n18185) );
  INV_X2 U13276 ( .I(n23057), .ZN(n31566) );
  NAND2_X2 U24688 ( .A1(n384), .A2(n20338), .ZN(n20340) );
  INV_X2 U6363 ( .I(n22119), .ZN(n22092) );
  OAI21_X2 U3859 ( .A1(n6285), .A2(n8290), .B(n14420), .ZN(n27695) );
  NAND2_X2 U10029 ( .A1(n18988), .A2(n6510), .ZN(n18899) );
  INV_X4 U7254 ( .I(n30879), .ZN(n18919) );
  NOR2_X2 U16238 ( .A1(n33022), .A2(n23034), .ZN(n16919) );
  AOI22_X2 U1411 ( .A1(n13680), .A2(n922), .B1(n28886), .B2(n13582), .ZN(
        n16085) );
  INV_X4 U6822 ( .I(n4568), .ZN(n26167) );
  INV_X4 U21313 ( .I(n24114), .ZN(n17068) );
  AOI22_X2 U4832 ( .A1(n18413), .A2(n18845), .B1(n18730), .B2(n18412), .ZN(
        n30336) );
  AOI21_X1 U23716 ( .A1(n20244), .A2(n20312), .B(n936), .ZN(n20245) );
  INV_X2 U7844 ( .I(n29303), .ZN(n21396) );
  AOI21_X1 U8726 ( .A1(n32009), .A2(n5677), .B(n5676), .ZN(n9840) );
  OAI22_X2 U4555 ( .A1(n1290), .A2(n6478), .B1(n33320), .B2(n22588), .ZN(
        n22438) );
  INV_X2 U11797 ( .I(n13610), .ZN(n13609) );
  INV_X2 U15013 ( .I(n7809), .ZN(n24260) );
  NAND2_X1 U14744 ( .A1(n16921), .A2(n28415), .ZN(n16920) );
  BUF_X2 U3129 ( .I(n13320), .Z(n25967) );
  NAND2_X2 U2660 ( .A1(n205), .A2(n204), .ZN(n20204) );
  NAND2_X2 U17965 ( .A1(n22478), .A2(n900), .ZN(n6956) );
  NOR3_X2 U1185 ( .A1(n31220), .A2(n517), .A3(n29084), .ZN(n15885) );
  NAND2_X1 U12980 ( .A1(n2070), .A2(n9146), .ZN(n2069) );
  NOR2_X1 U20432 ( .A1(n4067), .A2(n1281), .ZN(n11058) );
  OR2_X1 U3953 ( .A1(n8622), .A2(n3843), .Z(n29050) );
  NAND2_X2 U3877 ( .A1(n10031), .A2(n22876), .ZN(n14667) );
  NOR2_X2 U6166 ( .A1(n29239), .A2(n31428), .ZN(n28933) );
  INV_X2 U2621 ( .I(n19195), .ZN(n19606) );
  INV_X2 U5458 ( .I(n9759), .ZN(n16193) );
  INV_X4 U635 ( .I(n510), .ZN(n10686) );
  INV_X2 U6610 ( .I(n7680), .ZN(n1379) );
  AND2_X2 U13315 ( .A1(n20615), .A2(n9252), .Z(n20362) );
  OAI21_X2 U14493 ( .A1(n4339), .A2(n23103), .B(n3600), .ZN(n12790) );
  AOI21_X2 U21037 ( .A1(n905), .A2(n1116), .B(n12632), .ZN(n13104) );
  NAND3_X2 U8508 ( .A1(n7737), .A2(n11408), .A3(n32296), .ZN(n7736) );
  INV_X2 U16201 ( .I(n28697), .ZN(n3570) );
  INV_X2 U12957 ( .I(n11068), .ZN(n20008) );
  OAI21_X2 U2281 ( .A1(n17223), .A2(n12837), .B(n15108), .ZN(n8823) );
  NOR2_X2 U26328 ( .A1(n22396), .A2(n22398), .ZN(n5304) );
  NOR2_X2 U17397 ( .A1(n33915), .A2(n6345), .ZN(n11990) );
  NAND2_X2 U11903 ( .A1(n15267), .A2(n12168), .ZN(n3941) );
  INV_X2 U49 ( .I(n31407), .ZN(n27183) );
  NAND2_X2 U8786 ( .A1(n16538), .A2(n1189), .ZN(n14614) );
  NAND3_X1 U1410 ( .A1(n14943), .A2(n15400), .A3(n27455), .ZN(n14942) );
  INV_X4 U7641 ( .I(n24328), .ZN(n890) );
  NOR2_X2 U3095 ( .A1(n26912), .A2(n16648), .ZN(n15979) );
  AOI21_X2 U5470 ( .A1(n18953), .A2(n17445), .B(n18952), .ZN(n18924) );
  NAND2_X2 U14583 ( .A1(n14173), .A2(n19875), .ZN(n20290) );
  AOI21_X2 U5472 ( .A1(n19356), .A2(n6516), .B(n19359), .ZN(n14709) );
  NAND2_X1 U1748 ( .A1(n29202), .A2(n29201), .ZN(n20171) );
  NAND2_X2 U23504 ( .A1(n33659), .A2(n23559), .ZN(n16083) );
  INV_X4 U13400 ( .I(n27390), .ZN(n17185) );
  INV_X4 U1182 ( .I(n21259), .ZN(n28257) );
  OR2_X1 U20370 ( .A1(n30010), .A2(n27970), .Z(n7282) );
  INV_X4 U551 ( .I(n31220), .ZN(n17021) );
  OAI22_X1 U22594 ( .A1(n11156), .A2(n25916), .B1(n11155), .B2(n1206), .ZN(
        n28331) );
  OAI21_X2 U6751 ( .A1(n10310), .A2(n9958), .B(n22574), .ZN(n5453) );
  NAND2_X2 U15796 ( .A1(n4385), .A2(n28806), .ZN(n4384) );
  INV_X4 U10093 ( .I(n14812), .ZN(n16916) );
  OR3_X1 U3426 ( .A1(n1127), .A2(n9630), .A3(n3392), .Z(n2548) );
  INV_X2 U12826 ( .I(n7672), .ZN(n17341) );
  INV_X2 U16264 ( .I(n987), .ZN(n27298) );
  AOI21_X2 U6615 ( .A1(n29454), .A2(n1009), .B(n2339), .ZN(n2338) );
  INV_X2 U8489 ( .I(n20463), .ZN(n16518) );
  BUF_X2 U3147 ( .I(n21210), .Z(n16512) );
  INV_X2 U7738 ( .I(n5897), .ZN(n1081) );
  INV_X2 U4683 ( .I(n10775), .ZN(n26725) );
  NAND2_X2 U12040 ( .A1(n5033), .A2(n946), .ZN(n1767) );
  OR2_X1 U3643 ( .A1(n8444), .A2(n17117), .Z(n24878) );
  BUF_X2 U3812 ( .I(n8700), .Z(n8010) );
  NOR2_X2 U1664 ( .A1(n17263), .A2(n13154), .ZN(n26375) );
  NAND2_X2 U20496 ( .A1(n10389), .A2(n17186), .ZN(n27994) );
  NAND2_X2 U2421 ( .A1(n13884), .A2(n28203), .ZN(n31859) );
  CLKBUF_X4 U22350 ( .I(n24254), .Z(n28296) );
  NAND2_X2 U3488 ( .A1(n33889), .A2(n33147), .ZN(n2715) );
  NAND2_X2 U8457 ( .A1(n1150), .A2(n16684), .ZN(n1635) );
  AOI21_X2 U7602 ( .A1(n18633), .A2(n1439), .B(n17516), .ZN(n15811) );
  NAND2_X1 U10686 ( .A1(n16832), .A2(n1603), .ZN(n1602) );
  INV_X2 U16889 ( .I(n13147), .ZN(n23611) );
  INV_X2 U13694 ( .I(n19699), .ZN(n19619) );
  OAI21_X2 U14071 ( .A1(n732), .A2(n27228), .B(n16318), .ZN(n3112) );
  AOI21_X2 U14352 ( .A1(n21645), .A2(n861), .B(n27073), .ZN(n27754) );
  NAND2_X2 U290 ( .A1(n31419), .A2(n31421), .ZN(n30509) );
  NAND2_X1 U1826 ( .A1(n7462), .A2(n26320), .ZN(n26956) );
  NAND2_X2 U11035 ( .A1(n7066), .A2(n32678), .ZN(n27486) );
  INV_X4 U15623 ( .I(n16458), .ZN(n851) );
  NAND2_X2 U223 ( .A1(n16704), .A2(n25561), .ZN(n30561) );
  BUF_X4 U1492 ( .I(n34156), .Z(n31030) );
  BUF_X4 U7215 ( .I(n20882), .Z(n21163) );
  NOR2_X2 U633 ( .A1(n8967), .A2(n22956), .ZN(n28495) );
  OAI21_X2 U8970 ( .A1(n32911), .A2(n5202), .B(n25114), .ZN(n9050) );
  AOI21_X2 U4073 ( .A1(n24074), .A2(n24073), .B(n27038), .ZN(n9068) );
  INV_X2 U17337 ( .I(n27211), .ZN(n27458) );
  INV_X2 U6901 ( .I(n17150), .ZN(n893) );
  INV_X2 U1814 ( .I(n13327), .ZN(n29338) );
  NOR2_X2 U10582 ( .A1(n16443), .A2(n32178), .ZN(n10397) );
  OAI21_X2 U5496 ( .A1(n4518), .A2(n21078), .B(n28502), .ZN(n28501) );
  INV_X2 U20099 ( .I(n10337), .ZN(n11814) );
  NOR3_X1 U294 ( .A1(n30715), .A2(n1550), .A3(n28410), .ZN(n3214) );
  BUF_X4 U311 ( .I(n15227), .Z(n11200) );
  NAND3_X2 U24479 ( .A1(n19962), .A2(n28767), .A3(n6748), .ZN(n9978) );
  NAND2_X2 U2668 ( .A1(n8593), .A2(n22642), .ZN(n8332) );
  NOR2_X2 U1122 ( .A1(n9721), .A2(n17841), .ZN(n16189) );
  NAND2_X2 U10383 ( .A1(n9807), .A2(n1079), .ZN(n9806) );
  INV_X4 U3801 ( .I(n19332), .ZN(n7732) );
  INV_X1 U3181 ( .I(n23925), .ZN(n23763) );
  INV_X4 U20730 ( .I(n11744), .ZN(n18923) );
  OAI21_X2 U1085 ( .A1(n21187), .A2(n5239), .B(n5238), .ZN(n26413) );
  INV_X4 U14426 ( .I(n25889), .ZN(n14805) );
  INV_X1 U4980 ( .I(n25865), .ZN(n12266) );
  OAI22_X2 U8947 ( .A1(n12164), .A2(n32911), .B1(n9936), .B2(n12165), .ZN(
        n6629) );
  NAND2_X1 U15009 ( .A1(n30283), .A2(n14759), .ZN(n14758) );
  NOR2_X1 U15008 ( .A1(n16100), .A2(n7203), .ZN(n14759) );
  NAND3_X2 U3821 ( .A1(n20872), .A2(n12902), .A3(n20311), .ZN(n3402) );
  NAND2_X2 U853 ( .A1(n16009), .A2(n14281), .ZN(n14283) );
  INV_X4 U3540 ( .I(n19315), .ZN(n2081) );
  OAI21_X2 U3863 ( .A1(n7529), .A2(n7528), .B(n22986), .ZN(n29060) );
  NOR2_X2 U1720 ( .A1(n18137), .A2(n20910), .ZN(n18136) );
  OAI21_X1 U14880 ( .A1(n3862), .A2(n23608), .B(n3861), .ZN(n23610) );
  AOI22_X2 U16820 ( .A1(n7643), .A2(n10845), .B1(n19338), .B2(n5707), .ZN(
        n7327) );
  AOI21_X2 U4605 ( .A1(n25453), .A2(n17948), .B(n11640), .ZN(n25454) );
  INV_X2 U7255 ( .I(n18919), .ZN(n18621) );
  BUF_X4 U1083 ( .I(n7753), .Z(n230) );
  NAND2_X1 U440 ( .A1(n29360), .A2(n22636), .ZN(n15611) );
  AOI21_X2 U2435 ( .A1(n10113), .A2(n21149), .B(n2738), .ZN(n8727) );
  NAND2_X2 U748 ( .A1(n20200), .A2(n1789), .ZN(n205) );
  OR2_X2 U6915 ( .A1(n22591), .A2(n31549), .Z(n11873) );
  INV_X4 U5680 ( .I(n13343), .ZN(n794) );
  OR2_X2 U813 ( .A1(n22656), .A2(n17899), .Z(n13318) );
  CLKBUF_X4 U1611 ( .I(n18768), .Z(n28757) );
  INV_X4 U3809 ( .I(n1736), .ZN(n1329) );
  BUF_X2 U8606 ( .I(n9201), .Z(n2166) );
  NAND2_X2 U1589 ( .A1(n5535), .A2(n25337), .ZN(n5534) );
  BUF_X4 U1266 ( .I(n6255), .Z(n26471) );
  NAND2_X1 U17386 ( .A1(n12192), .A2(n12193), .ZN(n30469) );
  BUF_X2 U5010 ( .I(n12763), .Z(n29323) );
  NAND2_X2 U8011 ( .A1(n22522), .A2(n27638), .ZN(n10389) );
  INV_X1 U3055 ( .I(n17503), .ZN(n22752) );
  OAI22_X2 U1552 ( .A1(n3313), .A2(n18106), .B1(n9191), .B2(n10571), .ZN(n3312) );
  OAI22_X2 U11365 ( .A1(n26904), .A2(n8825), .B1(n11276), .B2(n21818), .ZN(
        n6699) );
  INV_X2 U7018 ( .I(n24874), .ZN(n17787) );
  INV_X1 U10749 ( .I(n17579), .ZN(n10498) );
  NAND2_X2 U15377 ( .A1(n11892), .A2(n10354), .ZN(n5140) );
  INV_X4 U592 ( .I(n21651), .ZN(n15371) );
  NOR2_X2 U8728 ( .A1(n22795), .A2(n33007), .ZN(n13120) );
  OAI22_X2 U8364 ( .A1(n18859), .A2(n18543), .B1(n18854), .B2(n18855), .ZN(
        n18417) );
  AOI21_X2 U3058 ( .A1(n14231), .A2(n1633), .B(n1887), .ZN(n1524) );
  BUF_X4 U5751 ( .I(n15329), .Z(n27875) );
  NAND3_X1 U3385 ( .A1(n13981), .A2(n11096), .A3(n13982), .ZN(n31090) );
  NAND2_X2 U166 ( .A1(n23982), .A2(n24246), .ZN(n13633) );
  NAND2_X2 U6968 ( .A1(n24325), .A2(n24328), .ZN(n24246) );
  NAND2_X2 U18955 ( .A1(n19844), .A2(n10086), .ZN(n7309) );
  NOR2_X2 U21506 ( .A1(n31097), .A2(n19923), .ZN(n4648) );
  OAI21_X2 U9883 ( .A1(n16029), .A2(n16346), .B(n940), .ZN(n2492) );
  NAND2_X2 U2675 ( .A1(n1874), .A2(n16323), .ZN(n9807) );
  INV_X2 U14139 ( .I(n21532), .ZN(n30678) );
  NAND2_X2 U4852 ( .A1(n27738), .A2(n12540), .ZN(n5059) );
  INV_X1 U261 ( .I(n29268), .ZN(n13291) );
  INV_X2 U23826 ( .I(n17143), .ZN(n18701) );
  NOR2_X1 U1397 ( .A1(n31906), .A2(n26774), .ZN(n5869) );
  NAND2_X1 U12156 ( .A1(n8860), .A2(n28056), .ZN(n12192) );
  NOR2_X2 U1899 ( .A1(n11075), .A2(n28345), .ZN(n30743) );
  NAND2_X1 U15092 ( .A1(n14209), .A2(n16231), .ZN(n8122) );
  NOR2_X2 U17244 ( .A1(n12221), .A2(n423), .ZN(n6447) );
  INV_X2 U10772 ( .I(n9328), .ZN(n3241) );
  NOR2_X2 U1897 ( .A1(n747), .A2(n30288), .ZN(n16973) );
  OAI21_X2 U11423 ( .A1(n18106), .A2(n18035), .B(n7723), .ZN(n7722) );
  OAI21_X1 U22287 ( .A1(n1132), .A2(n21811), .B(n31627), .ZN(n11167) );
  NAND3_X2 U2867 ( .A1(n434), .A2(n14449), .A3(n433), .ZN(n30199) );
  INV_X2 U8113 ( .I(n22225), .ZN(n10650) );
  NOR2_X1 U14089 ( .A1(n24329), .A2(n24328), .ZN(n30186) );
  NAND2_X1 U4930 ( .A1(n28261), .A2(n20546), .ZN(n20547) );
  AOI21_X2 U3145 ( .A1(n15611), .A2(n16240), .B(n15609), .ZN(n15608) );
  NAND2_X2 U2945 ( .A1(n2877), .A2(n23055), .ZN(n4845) );
  INV_X2 U16746 ( .I(n14619), .ZN(n14745) );
  AOI22_X2 U21720 ( .A1(n31120), .A2(n17483), .B1(n17482), .B2(n772), .ZN(
        n9747) );
  NOR2_X2 U19305 ( .A1(n31722), .A2(n28691), .ZN(n9973) );
  OAI21_X2 U10648 ( .A1(n13879), .A2(n17612), .B(n30980), .ZN(n13878) );
  NAND3_X2 U13153 ( .A1(n16261), .A2(n16262), .A3(n2229), .ZN(n16747) );
  BUF_X2 U4453 ( .I(n2256), .Z(n27694) );
  NAND2_X2 U4569 ( .A1(n28840), .A2(n15169), .ZN(n20430) );
  INV_X2 U1948 ( .I(n30663), .ZN(n30937) );
  AND2_X1 U4584 ( .A1(n15057), .A2(n10708), .Z(n14644) );
  INV_X4 U10286 ( .I(n6985), .ZN(n13592) );
  OR2_X2 U96 ( .A1(n8542), .A2(n13050), .Z(n25874) );
  BUF_X4 U17725 ( .I(n639), .Z(n30529) );
  INV_X2 U1115 ( .I(n14594), .ZN(n30115) );
  NAND2_X1 U18692 ( .A1(n30661), .A2(n30660), .ZN(n13707) );
  NOR2_X1 U11739 ( .A1(n7872), .A2(n20615), .ZN(n6797) );
  OAI22_X2 U2037 ( .A1(n8739), .A2(n18815), .B1(n18639), .B2(n9118), .ZN(n4843) );
  INV_X1 U5088 ( .I(n10757), .ZN(n12281) );
  NOR2_X2 U6796 ( .A1(n708), .A2(n28160), .ZN(n10138) );
  OAI21_X1 U15401 ( .A1(n23042), .A2(n17930), .B(n808), .ZN(n13121) );
  INV_X2 U11350 ( .I(n21496), .ZN(n21713) );
  INV_X1 U12524 ( .I(n11513), .ZN(n14483) );
  NAND2_X1 U14874 ( .A1(n21483), .A2(n1327), .ZN(n21484) );
  NAND2_X1 U20853 ( .A1(n21427), .A2(n33215), .ZN(n14598) );
  NAND3_X2 U3256 ( .A1(n1492), .A2(n1382), .A3(n19205), .ZN(n1491) );
  INV_X4 U9702 ( .I(n29314), .ZN(n22992) );
  NOR2_X1 U10870 ( .A1(n28141), .A2(n15885), .ZN(n31889) );
  CLKBUF_X4 U264 ( .I(n17037), .Z(n16957) );
  BUF_X4 U212 ( .I(n25382), .Z(n31149) );
  INV_X4 U71 ( .I(n25546), .ZN(n12864) );
  NAND2_X2 U2516 ( .A1(n11895), .A2(n22435), .ZN(n2522) );
  NOR2_X2 U18827 ( .A1(n6176), .A2(n2217), .ZN(n8274) );
  INV_X4 U17240 ( .I(n10724), .ZN(n30448) );
  INV_X4 U1636 ( .I(n14213), .ZN(n1182) );
  BUF_X4 U768 ( .I(n4084), .Z(n29648) );
  NAND2_X2 U345 ( .A1(n28745), .A2(n28744), .ZN(n4481) );
  INV_X1 U3612 ( .I(n7880), .ZN(n31509) );
  NAND2_X1 U1554 ( .A1(n30471), .A2(n15898), .ZN(n26720) );
  INV_X2 U3854 ( .I(n25), .ZN(n17955) );
  BUF_X2 U1688 ( .I(n20401), .Z(n27785) );
  BUF_X4 U1150 ( .I(n29258), .Z(n2551) );
  INV_X2 U14873 ( .I(n18198), .ZN(n12290) );
  OR2_X1 U5860 ( .A1(n26881), .A2(n13300), .Z(n13562) );
  INV_X4 U7184 ( .I(n505), .ZN(n5239) );
  INV_X4 U7900 ( .I(n7915), .ZN(n8547) );
  INV_X4 U8482 ( .I(n27504), .ZN(n29258) );
  OR2_X1 U7235 ( .A1(n8314), .A2(n17960), .Z(n29424) );
  INV_X2 U5312 ( .I(n31810), .ZN(n16271) );
  INV_X2 U8070 ( .I(n22589), .ZN(n22584) );
  INV_X4 U22583 ( .I(n28329), .ZN(n2023) );
  CLKBUF_X4 U1883 ( .I(n15960), .Z(n400) );
  NAND2_X1 U4772 ( .A1(n5494), .A2(n30832), .ZN(n12788) );
  NAND3_X1 U1526 ( .A1(n17270), .A2(n26800), .A3(n16762), .ZN(n29899) );
  NAND2_X2 U6189 ( .A1(n15211), .A2(n14159), .ZN(n28438) );
  NAND2_X2 U6230 ( .A1(n1057), .A2(n18721), .ZN(n6203) );
  INV_X2 U21203 ( .I(n16570), .ZN(n14034) );
  NOR2_X2 U10975 ( .A1(n16927), .A2(n22760), .ZN(n16926) );
  NAND2_X1 U5445 ( .A1(n9173), .A2(n20143), .ZN(n7820) );
  BUF_X2 U4186 ( .I(n8277), .Z(n28091) );
  AOI21_X2 U14680 ( .A1(n11013), .A2(n20052), .B(n3769), .ZN(n6931) );
  BUF_X4 U3287 ( .I(n18028), .Z(n27801) );
  INV_X4 U485 ( .I(n11895), .ZN(n1298) );
  NAND2_X2 U352 ( .A1(n8058), .A2(n18077), .ZN(n13109) );
  OR2_X1 U16168 ( .A1(n30988), .A2(n17271), .Z(n17272) );
  NOR2_X2 U10696 ( .A1(n8654), .A2(n11653), .ZN(n3983) );
  NAND3_X2 U7156 ( .A1(n21192), .A2(n26542), .A3(n33949), .ZN(n8046) );
  NAND2_X2 U2104 ( .A1(n20520), .A2(n5460), .ZN(n73) );
  NOR2_X2 U9351 ( .A1(n14157), .A2(n7179), .ZN(n14773) );
  NOR2_X1 U1659 ( .A1(n29409), .A2(n19792), .ZN(n30572) );
  NAND2_X2 U10000 ( .A1(n18667), .A2(n26518), .ZN(n8211) );
  AOI21_X2 U967 ( .A1(n909), .A2(n22427), .B(n22537), .ZN(n14388) );
  AOI22_X1 U4427 ( .A1(n17802), .A2(n6476), .B1(n17801), .B2(n16868), .ZN(
        n17800) );
  INV_X1 U8111 ( .I(n13553), .ZN(n1004) );
  INV_X4 U7434 ( .I(n12408), .ZN(n3790) );
  OAI21_X2 U5650 ( .A1(n22635), .A2(n22640), .B(n4511), .ZN(n4510) );
  NAND3_X2 U15070 ( .A1(n1243), .A2(n24193), .A3(n31918), .ZN(n23990) );
  AOI21_X2 U8769 ( .A1(n26036), .A2(n8273), .B(n26397), .ZN(n27391) );
  BUF_X2 U6984 ( .I(n8480), .Z(n27211) );
  NOR2_X1 U13505 ( .A1(n30124), .A2(n2764), .ZN(n31021) );
  NAND2_X2 U5753 ( .A1(n17568), .A2(n17567), .ZN(n22961) );
  INV_X1 U11507 ( .I(n29908), .ZN(n565) );
  NAND2_X2 U8612 ( .A1(n26751), .A2(n8237), .ZN(n8717) );
  NAND2_X2 U7441 ( .A1(n18668), .A2(n18669), .ZN(n8237) );
  INV_X2 U5080 ( .I(n3723), .ZN(n15798) );
  NAND2_X1 U16250 ( .A1(n31968), .A2(n17236), .ZN(n7035) );
  INV_X2 U516 ( .I(n22121), .ZN(n1305) );
  AOI21_X2 U6746 ( .A1(n26347), .A2(n22425), .B(n14728), .ZN(n22603) );
  NAND2_X2 U829 ( .A1(n16665), .A2(n28915), .ZN(n26347) );
  BUF_X2 U4041 ( .I(n10303), .Z(n22546) );
  NOR2_X1 U20479 ( .A1(n28614), .A2(n31174), .ZN(n7440) );
  NOR2_X2 U2413 ( .A1(n4318), .A2(n15550), .ZN(n13052) );
  INV_X2 U1813 ( .I(n871), .ZN(n7460) );
  NOR2_X2 U5023 ( .A1(n23930), .A2(n29269), .ZN(n23538) );
  NAND2_X2 U13660 ( .A1(n17726), .A2(n8834), .ZN(n31560) );
  AND2_X2 U19562 ( .A1(n8386), .A2(n32051), .Z(n18878) );
  INV_X2 U708 ( .I(n12315), .ZN(n22807) );
  NAND2_X2 U6636 ( .A1(n18760), .A2(n18759), .ZN(n15281) );
  NAND2_X2 U4085 ( .A1(n6249), .A2(n6248), .ZN(n23594) );
  NAND2_X2 U15979 ( .A1(n11232), .A2(n17832), .ZN(n7651) );
  INV_X2 U10893 ( .I(n8786), .ZN(n8415) );
  NAND2_X2 U8953 ( .A1(n16024), .A2(n32911), .ZN(n9936) );
  OR2_X2 U11201 ( .A1(n22599), .A2(n16432), .Z(n22510) );
  NOR2_X2 U23068 ( .A1(n4113), .A2(n27090), .ZN(n22775) );
  CLKBUF_X4 U1966 ( .I(n19206), .Z(n4202) );
  OAI21_X2 U6838 ( .A1(n22993), .A2(n22992), .B(n30388), .ZN(n22997) );
  BUF_X4 U5653 ( .I(n22978), .Z(n8990) );
  NAND3_X2 U8603 ( .A1(n26384), .A2(n17880), .A3(n26383), .ZN(n26589) );
  NAND2_X2 U25107 ( .A1(n22563), .A2(n14034), .ZN(n22564) );
  AOI21_X2 U15040 ( .A1(n27314), .A2(n15084), .B(n24983), .ZN(n15223) );
  NAND2_X2 U1848 ( .A1(n23940), .A2(n26965), .ZN(n13678) );
  INV_X2 U153 ( .I(n24436), .ZN(n718) );
  AOI22_X2 U1484 ( .A1(n1490), .A2(n27970), .B1(n19242), .B2(n1494), .ZN(
        n26293) );
  AND2_X1 U12836 ( .A1(n13354), .A2(n33789), .Z(n26836) );
  INV_X2 U15827 ( .I(n20310), .ZN(n1154) );
  INV_X4 U1004 ( .I(n22435), .ZN(n31636) );
  INV_X2 U16891 ( .I(n7463), .ZN(n11235) );
  INV_X1 U5715 ( .I(n522), .ZN(n29336) );
  NOR2_X2 U11050 ( .A1(n26628), .A2(n13677), .ZN(n27044) );
  INV_X2 U473 ( .I(n18098), .ZN(n22474) );
  BUF_X4 U4240 ( .I(n15411), .Z(n1883) );
  NAND3_X1 U15295 ( .A1(n17742), .A2(n17743), .A3(n17741), .ZN(n30583) );
  NOR3_X2 U18159 ( .A1(n31007), .A2(n21642), .A3(n32613), .ZN(n12274) );
  NAND2_X2 U14981 ( .A1(n25399), .A2(n1700), .ZN(n25402) );
  NOR2_X2 U24680 ( .A1(n20563), .A2(n17329), .ZN(n20285) );
  NOR2_X2 U14095 ( .A1(n32788), .A2(n15137), .ZN(n7437) );
  NOR2_X2 U53 ( .A1(n15531), .A2(n15530), .ZN(n15529) );
  NAND2_X2 U11126 ( .A1(n7398), .A2(n10630), .ZN(n6455) );
  NAND2_X1 U12629 ( .A1(n26808), .A2(n15971), .ZN(n9166) );
  INV_X2 U6549 ( .I(n20008), .ZN(n1359) );
  NAND2_X2 U6062 ( .A1(n10897), .A2(n14915), .ZN(n15546) );
  NAND2_X1 U23220 ( .A1(n15418), .A2(n15416), .ZN(n28444) );
  INV_X4 U655 ( .I(n758), .ZN(n23104) );
  OAI21_X2 U11520 ( .A1(n15632), .A2(n12027), .B(n31826), .ZN(n15631) );
  OAI22_X2 U14770 ( .A1(n25470), .A2(n25490), .B1(n25479), .B2(n25487), .ZN(
        n25492) );
  INV_X2 U3783 ( .I(n27741), .ZN(n7873) );
  INV_X2 U6286 ( .I(n18261), .ZN(n23100) );
  NAND2_X2 U14868 ( .A1(n25479), .A2(n25488), .ZN(n25463) );
  NOR2_X2 U1934 ( .A1(n19267), .A2(n19268), .ZN(n2098) );
  NAND2_X2 U417 ( .A1(n27163), .A2(n23872), .ZN(n31528) );
  BUF_X2 U1435 ( .I(n21442), .Z(n16180) );
  NAND2_X2 U9691 ( .A1(n17939), .A2(n32457), .ZN(n3211) );
  OAI21_X2 U8339 ( .A1(n31729), .A2(n29574), .B(n29573), .ZN(n17939) );
  OAI21_X1 U24760 ( .A1(n17200), .A2(n17199), .B(n25467), .ZN(n31492) );
  INV_X4 U4259 ( .I(n5225), .ZN(n16466) );
  NAND2_X1 U16121 ( .A1(n2052), .A2(n19782), .ZN(n19791) );
  INV_X2 U5460 ( .I(n20010), .ZN(n1167) );
  BUF_X4 U22924 ( .I(n14624), .Z(n28386) );
  INV_X2 U3604 ( .I(n23300), .ZN(n23414) );
  NAND2_X2 U6876 ( .A1(n4408), .A2(n976), .ZN(n5417) );
  NOR3_X2 U17074 ( .A1(n28625), .A2(n30793), .A3(n27386), .ZN(n4980) );
  NOR3_X2 U3281 ( .A1(n9817), .A2(n1019), .A3(n9816), .ZN(n29221) );
  INV_X2 U16610 ( .I(n14156), .ZN(n18637) );
  BUF_X2 U9000 ( .I(n15777), .Z(n11716) );
  NOR2_X2 U10988 ( .A1(n29242), .A2(n28680), .ZN(n22988) );
  NAND3_X2 U24731 ( .A1(n15468), .A2(n33154), .A3(n28899), .ZN(n20619) );
  INV_X2 U3090 ( .I(n15123), .ZN(n23033) );
  BUF_X4 U24127 ( .I(n20103), .Z(n28600) );
  CLKBUF_X4 U1505 ( .I(n19101), .Z(n6511) );
  AOI21_X2 U18259 ( .A1(n1246), .A2(n24311), .B(n7481), .ZN(n7480) );
  OAI22_X1 U10887 ( .A1(n6035), .A2(n3202), .B1(n3201), .B2(n1107), .ZN(n3200)
         );
  NAND3_X1 U10427 ( .A1(n29116), .A2(n30047), .A3(n25462), .ZN(n25458) );
  NAND2_X2 U14911 ( .A1(n31883), .A2(n24154), .ZN(n5367) );
  NOR2_X2 U857 ( .A1(n2471), .A2(n22926), .ZN(n9335) );
  INV_X4 U6707 ( .I(n16732), .ZN(n956) );
  INV_X4 U7652 ( .I(n18131), .ZN(n18815) );
  NAND2_X2 U20835 ( .A1(n15638), .A2(n33730), .ZN(n12847) );
  INV_X4 U846 ( .I(n19998), .ZN(n7609) );
  OAI22_X2 U26365 ( .A1(n19147), .A2(n15534), .B1(n1175), .B2(n1055), .ZN(
        n5654) );
  INV_X1 U1781 ( .I(n20886), .ZN(n29169) );
  INV_X2 U22629 ( .I(n19267), .ZN(n15869) );
  INV_X1 U6282 ( .I(n22848), .ZN(n15976) );
  BUF_X4 U3261 ( .I(n25894), .Z(n4993) );
  CLKBUF_X4 U2077 ( .I(n6039), .Z(n1125) );
  CLKBUF_X4 U4465 ( .I(n13232), .Z(n2744) );
  NAND2_X2 U6738 ( .A1(n23104), .A2(n23103), .ZN(n26161) );
  NAND2_X2 U4764 ( .A1(n24067), .A2(n10033), .ZN(n3216) );
  NAND3_X2 U21348 ( .A1(n28435), .A2(n27619), .A3(n27336), .ZN(n31886) );
  AOI21_X2 U17378 ( .A1(n17260), .A2(n71), .B(n12398), .ZN(n16977) );
  AND2_X2 U2697 ( .A1(n16275), .A2(n515), .Z(n21320) );
  INV_X2 U15270 ( .I(n32358), .ZN(n6119) );
  BUF_X4 U15544 ( .I(n11570), .Z(n15054) );
  BUF_X2 U8860 ( .I(Key[32]), .Z(n25428) );
  INV_X4 U3968 ( .I(n13905), .ZN(n23760) );
  BUF_X2 U4233 ( .I(n14255), .Z(n27577) );
  INV_X1 U4266 ( .I(n23827), .ZN(n26775) );
  NAND2_X1 U4706 ( .A1(n7756), .A2(n28257), .ZN(n27245) );
  INV_X2 U6077 ( .I(n18892), .ZN(n29683) );
  INV_X4 U22274 ( .I(n839), .ZN(n24154) );
  OAI21_X2 U3153 ( .A1(n19248), .A2(n3535), .B(n19247), .ZN(n19251) );
  NAND2_X2 U9823 ( .A1(n7307), .A2(n19844), .ZN(n3061) );
  NOR2_X1 U6180 ( .A1(n23712), .A2(n17234), .ZN(n14778) );
  BUF_X2 U3507 ( .I(n25696), .Z(n16609) );
  NAND3_X1 U15156 ( .A1(n1555), .A2(n9258), .A3(n27462), .ZN(n30779) );
  NAND3_X2 U16574 ( .A1(n22686), .A2(n33964), .A3(n22685), .ZN(n31902) );
  AOI21_X2 U1067 ( .A1(n11713), .A2(n17445), .B(n8192), .ZN(n11178) );
  NOR3_X2 U17214 ( .A1(n32831), .A2(n13703), .A3(n13525), .ZN(n6216) );
  NAND2_X2 U22560 ( .A1(n20484), .A2(n31009), .ZN(n28324) );
  AOI22_X2 U10139 ( .A1(n18470), .A2(n18007), .B1(n18469), .B2(n18006), .ZN(
        n18473) );
  AOI21_X2 U13278 ( .A1(n13730), .A2(n31826), .B(n6520), .ZN(n3888) );
  NOR2_X1 U12586 ( .A1(n15041), .A2(n12843), .ZN(n3035) );
  NAND2_X2 U84 ( .A1(n11696), .A2(n11697), .ZN(n11695) );
  OAI21_X2 U21458 ( .A1(n13036), .A2(n32143), .B(n29602), .ZN(n13035) );
  INV_X2 U14192 ( .I(n11516), .ZN(n13521) );
  NOR2_X2 U7833 ( .A1(n26282), .A2(n18033), .ZN(n18032) );
  NAND2_X2 U3594 ( .A1(n8770), .A2(n7218), .ZN(n20576) );
  NAND3_X2 U14799 ( .A1(n7803), .A2(n8033), .A3(n8107), .ZN(n7550) );
  INV_X2 U5904 ( .I(n31906), .ZN(n19960) );
  NAND2_X2 U14044 ( .A1(n16834), .A2(n26542), .ZN(n27016) );
  OAI21_X2 U11557 ( .A1(n21426), .A2(n13286), .B(n14168), .ZN(n16834) );
  INV_X2 U15050 ( .I(n26724), .ZN(n17828) );
  INV_X2 U8987 ( .I(n2023), .ZN(n26416) );
  OAI21_X2 U888 ( .A1(n25), .A2(n22621), .B(n995), .ZN(n22624) );
  OAI21_X2 U11040 ( .A1(n22024), .A2(n16170), .B(n2258), .ZN(n2257) );
  AOI22_X2 U4370 ( .A1(n11924), .A2(n29180), .B1(n21531), .B2(n8886), .ZN(
        n31244) );
  BUF_X2 U5894 ( .I(n19601), .Z(n19914) );
  BUF_X2 U5652 ( .I(n7012), .Z(n26884) );
  NOR2_X2 U4045 ( .A1(n18846), .A2(n17184), .ZN(n18413) );
  BUF_X4 U2215 ( .I(n16209), .Z(n100) );
  NAND2_X1 U6086 ( .A1(n6287), .A2(n10651), .ZN(n4520) );
  NAND2_X2 U1203 ( .A1(n8941), .A2(n28126), .ZN(n8940) );
  OAI21_X2 U542 ( .A1(n21794), .A2(n21792), .B(n30549), .ZN(n11560) );
  NAND3_X1 U25504 ( .A1(n24701), .A2(n11366), .A3(n25406), .ZN(n24704) );
  NAND2_X1 U10366 ( .A1(n6824), .A2(n6822), .ZN(n8743) );
  INV_X4 U3012 ( .I(n15278), .ZN(n8817) );
  CLKBUF_X4 U11232 ( .I(n19744), .Z(n29876) );
  OAI21_X2 U22907 ( .A1(n25160), .A2(n32553), .B(n25159), .ZN(n25163) );
  AOI22_X2 U18993 ( .A1(n25173), .A2(n7765), .B1(n8929), .B2(n25158), .ZN(
        n25159) );
  AOI22_X2 U1110 ( .A1(n19421), .A2(n29156), .B1(n19420), .B2(n19868), .ZN(
        n12705) );
  NAND2_X1 U11167 ( .A1(n29863), .A2(n5937), .ZN(n5935) );
  OAI22_X2 U15136 ( .A1(n11706), .A2(n22690), .B1(n8944), .B2(n32194), .ZN(
        n6943) );
  NAND2_X2 U16965 ( .A1(n355), .A2(n22690), .ZN(n8944) );
  NAND2_X2 U10991 ( .A1(n6371), .A2(n6370), .ZN(n6369) );
  AOI21_X2 U663 ( .A1(n26868), .A2(n14188), .B(n30904), .ZN(n6371) );
  INV_X2 U20735 ( .I(n11765), .ZN(n11923) );
  NOR2_X2 U9840 ( .A1(n29774), .A2(n20627), .ZN(n7836) );
  INV_X2 U5267 ( .I(n15063), .ZN(n27275) );
  OAI21_X2 U16179 ( .A1(n7765), .A2(n25175), .B(n25174), .ZN(n25177) );
  OAI21_X1 U10158 ( .A1(n882), .A2(n14213), .B(n12663), .ZN(n9046) );
  BUF_X4 U19699 ( .I(n27807), .Z(n30817) );
  NAND2_X2 U4071 ( .A1(n15068), .A2(n13601), .ZN(n23995) );
  NOR2_X2 U14839 ( .A1(n32890), .A2(n23807), .ZN(n13578) );
  AOI22_X2 U18599 ( .A1(n9316), .A2(n27077), .B1(n9315), .B2(n27818), .ZN(
        n9314) );
  BUF_X4 U359 ( .I(n13472), .Z(n7068) );
  NAND2_X2 U15977 ( .A1(n27367), .A2(n11232), .ZN(n26679) );
  NAND2_X2 U22597 ( .A1(n8862), .A2(n950), .ZN(n19329) );
  AOI22_X2 U24851 ( .A1(n21190), .A2(n21189), .B1(n33649), .B2(n21321), .ZN(
        n21191) );
  AOI21_X2 U17638 ( .A1(n18366), .A2(n18367), .B(n13254), .ZN(n27509) );
  BUF_X2 U5703 ( .I(n15617), .Z(n2471) );
  INV_X2 U22925 ( .I(n14605), .ZN(n17382) );
  BUF_X4 U3917 ( .I(n21693), .Z(n27635) );
  BUF_X4 U4904 ( .I(n18310), .Z(n14651) );
  OAI21_X2 U6391 ( .A1(n6954), .A2(n6953), .B(n1168), .ZN(n6952) );
  AND2_X2 U14473 ( .A1(n11707), .A2(n16462), .Z(n18634) );
  NOR2_X1 U9767 ( .A1(n16176), .A2(n782), .ZN(n5735) );
  NAND2_X2 U15621 ( .A1(n16611), .A2(n25149), .ZN(n6204) );
  NAND2_X2 U16070 ( .A1(n26900), .A2(n27457), .ZN(n30320) );
  OAI21_X1 U1388 ( .A1(n8348), .A2(n8349), .B(n9270), .ZN(n6945) );
  INV_X2 U2073 ( .I(n31773), .ZN(n8756) );
  NAND2_X1 U1620 ( .A1(n29995), .A2(n29994), .ZN(n29993) );
  NAND2_X1 U12381 ( .A1(n20259), .A2(n817), .ZN(n29995) );
  INV_X1 U541 ( .I(n4281), .ZN(n23593) );
  INV_X2 U11735 ( .I(n20328), .ZN(n11808) );
  NAND2_X2 U21396 ( .A1(n17993), .A2(n1350), .ZN(n17992) );
  BUF_X4 U6447 ( .I(n19260), .Z(n28379) );
  CLKBUF_X4 U11933 ( .I(n15476), .Z(n15381) );
  AOI21_X2 U16750 ( .A1(n13597), .A2(n30960), .B(n33675), .ZN(n5620) );
  INV_X2 U16956 ( .I(n21317), .ZN(n27367) );
  NOR2_X2 U7298 ( .A1(n33302), .A2(n32477), .ZN(n3240) );
  NAND2_X2 U4822 ( .A1(n17512), .A2(n28324), .ZN(n17511) );
  INV_X2 U21713 ( .I(n17916), .ZN(n22610) );
  NOR2_X1 U2353 ( .A1(n23058), .A2(n17462), .ZN(n28783) );
  NAND2_X1 U9126 ( .A1(n12568), .A2(n23896), .ZN(n3950) );
  NAND2_X1 U6990 ( .A1(n5140), .A2(n10216), .ZN(n10388) );
  INV_X2 U453 ( .I(n32926), .ZN(n15853) );
  NAND2_X1 U15964 ( .A1(n19803), .A2(n20006), .ZN(n27196) );
  NOR2_X2 U8995 ( .A1(n33120), .A2(n25697), .ZN(n3774) );
  NOR2_X2 U556 ( .A1(n13597), .A2(n15851), .ZN(n13619) );
  NOR2_X1 U5584 ( .A1(n23595), .A2(n11567), .ZN(n16969) );
  INV_X2 U5151 ( .I(n16625), .ZN(n941) );
  AOI22_X1 U22755 ( .A1(n17464), .A2(n30234), .B1(n22879), .B2(n22880), .ZN(
        n17463) );
  NAND2_X2 U17330 ( .A1(n2225), .A2(n7287), .ZN(n27457) );
  OR2_X2 U94 ( .A1(n1215), .A2(n25260), .Z(n6280) );
  NAND2_X1 U12095 ( .A1(n6207), .A2(n11122), .ZN(n8628) );
  NAND2_X2 U14752 ( .A1(n23791), .A2(n14460), .ZN(n9522) );
  OR2_X1 U3613 ( .A1(n13693), .A2(n20329), .Z(n20551) );
  NAND3_X1 U1338 ( .A1(n7386), .A2(n6309), .A3(n13291), .ZN(n6308) );
  OR2_X2 U184 ( .A1(n18151), .A2(n18150), .Z(n25591) );
  AOI21_X2 U122 ( .A1(n6551), .A2(n25332), .B(n15880), .ZN(n31786) );
  INV_X1 U198 ( .I(n15528), .ZN(n25411) );
  OAI21_X2 U4156 ( .A1(n13578), .A2(n6132), .B(n31208), .ZN(n6131) );
  INV_X1 U1874 ( .I(n16), .ZN(n29656) );
  OAI22_X2 U11432 ( .A1(n1785), .A2(n1329), .B1(n32248), .B2(n21061), .ZN(
        n1456) );
  NAND2_X1 U9703 ( .A1(n31350), .A2(n19291), .ZN(n31349) );
  NAND2_X1 U5752 ( .A1(n31871), .A2(n10344), .ZN(n10343) );
  INV_X2 U360 ( .I(n31437), .ZN(n1274) );
  OAI22_X2 U9347 ( .A1(n4812), .A2(n22467), .B1(n14376), .B2(n28865), .ZN(
        n4811) );
  NAND2_X1 U613 ( .A1(n13316), .A2(n13315), .ZN(n13314) );
  NOR2_X1 U19960 ( .A1(n30852), .A2(n12747), .ZN(n5248) );
  CLKBUF_X8 U15076 ( .I(n30978), .Z(n30769) );
  CLKBUF_X4 U8615 ( .I(n706), .Z(n25980) );
  CLKBUF_X4 U3155 ( .I(n16333), .Z(n9797) );
  BUF_X2 U7655 ( .I(Key[35]), .Z(n25131) );
  INV_X2 U22987 ( .I(n14798), .ZN(n17313) );
  INV_X4 U4239 ( .I(n1385), .ZN(n1047) );
  NOR2_X1 U11580 ( .A1(n28648), .A2(n986), .ZN(n26688) );
  NAND3_X2 U10973 ( .A1(n13597), .A2(n23093), .A3(n15039), .ZN(n23094) );
  INV_X4 U1530 ( .I(n9191), .ZN(n18106) );
  INV_X4 U5450 ( .I(n20100), .ZN(n937) );
  AOI21_X2 U1282 ( .A1(n15551), .A2(n16980), .B(n16979), .ZN(n16978) );
  NOR2_X2 U3177 ( .A1(n4205), .A2(n4204), .ZN(n5270) );
  BUF_X2 U2703 ( .I(n20939), .Z(n21357) );
  NOR2_X1 U17911 ( .A1(n5342), .A2(n27383), .ZN(n30984) );
  NAND2_X2 U7553 ( .A1(n18289), .A2(n18288), .ZN(n18290) );
  INV_X2 U8413 ( .I(n21085), .ZN(n11948) );
  NAND2_X2 U1614 ( .A1(n73), .A2(n14876), .ZN(n31878) );
  NAND2_X1 U19347 ( .A1(n23613), .A2(n29839), .ZN(n30754) );
  BUF_X2 U6874 ( .I(n29273), .Z(n31796) );
  NAND2_X2 U21118 ( .A1(n17466), .A2(n32242), .ZN(n12912) );
  NOR2_X2 U9500 ( .A1(n9206), .A2(n9204), .ZN(n5474) );
  BUF_X2 U11984 ( .I(n4314), .Z(n3727) );
  NAND2_X1 U21314 ( .A1(n17563), .A2(n17562), .ZN(n17561) );
  INV_X4 U10847 ( .I(n5381), .ZN(n9223) );
  NAND2_X2 U18711 ( .A1(n31007), .A2(n7553), .ZN(n21554) );
  INV_X2 U7148 ( .I(n17316), .ZN(n180) );
  OAI22_X2 U5636 ( .A1(n6225), .A2(n10529), .B1(n24216), .B2(n24109), .ZN(
        n10531) );
  NAND2_X1 U68 ( .A1(n27099), .A2(n9050), .ZN(n27731) );
  INV_X2 U5084 ( .I(n18539), .ZN(n14346) );
  NAND2_X2 U377 ( .A1(n26950), .A2(n8178), .ZN(n27826) );
  OAI21_X2 U3780 ( .A1(n20097), .A2(n1041), .B(n8182), .ZN(n8181) );
  INV_X2 U1295 ( .I(n26363), .ZN(n28471) );
  OR2_X2 U20140 ( .A1(n20208), .A2(n20207), .Z(n10460) );
  NAND3_X1 U21244 ( .A1(n19948), .A2(n20068), .A3(n20067), .ZN(n16084) );
  NOR2_X2 U7846 ( .A1(n23947), .A2(n29198), .ZN(n6272) );
  INV_X2 U10957 ( .I(n23088), .ZN(n14602) );
  NAND2_X1 U11700 ( .A1(n20159), .A2(n20333), .ZN(n12150) );
  OAI21_X1 U20901 ( .A1(n909), .A2(n5597), .B(n14388), .ZN(n14387) );
  AND3_X1 U4577 ( .A1(n10845), .A2(n34103), .A3(n6532), .Z(n10846) );
  NAND2_X2 U19901 ( .A1(n3180), .A2(n12886), .ZN(n9540) );
  NAND2_X2 U1638 ( .A1(n8454), .A2(n29867), .ZN(n11760) );
  NAND2_X2 U18580 ( .A1(n30640), .A2(n30639), .ZN(n22424) );
  OR2_X1 U10566 ( .A1(n9789), .A2(n11100), .Z(n17853) );
  INV_X2 U1183 ( .I(n20803), .ZN(n1343) );
  AOI21_X2 U21309 ( .A1(n22483), .A2(n9910), .B(n29158), .ZN(n15835) );
  INV_X2 U1880 ( .I(n19395), .ZN(n19740) );
  NOR3_X2 U20218 ( .A1(n15591), .A2(n15590), .A3(n20497), .ZN(n4061) );
  OAI21_X1 U11185 ( .A1(n22549), .A2(n27416), .B(n22315), .ZN(n22326) );
  INV_X4 U2948 ( .I(n11970), .ZN(n950) );
  NAND2_X2 U9365 ( .A1(n12334), .A2(n17960), .ZN(n12333) );
  INV_X1 U4083 ( .I(n24251), .ZN(n1092) );
  INV_X2 U3242 ( .I(n17439), .ZN(n21222) );
  BUF_X2 U20810 ( .I(n20657), .Z(n21079) );
  INV_X1 U3781 ( .I(n20097), .ZN(n20061) );
  NOR2_X1 U14397 ( .A1(n31514), .A2(n2906), .ZN(n30624) );
  INV_X1 U21302 ( .I(n18167), .ZN(n17730) );
  NOR2_X1 U14672 ( .A1(n2023), .A2(n23794), .ZN(n30251) );
  NAND3_X2 U14366 ( .A1(n31072), .A2(n28626), .A3(n28316), .ZN(n3465) );
  NOR2_X1 U14999 ( .A1(n25593), .A2(n13763), .ZN(n8246) );
  OAI21_X2 U10138 ( .A1(n18815), .A2(n18515), .B(n9211), .ZN(n8478) );
  INV_X4 U8776 ( .I(n18761), .ZN(n18288) );
  AOI22_X2 U24628 ( .A1(n20160), .A2(n20002), .B1(n742), .B2(n31072), .ZN(
        n20003) );
  NAND2_X1 U21284 ( .A1(n15490), .A2(n26965), .ZN(n13669) );
  NAND2_X2 U16414 ( .A1(n32012), .A2(n10629), .ZN(n27294) );
  NOR2_X1 U20599 ( .A1(n10381), .A2(n11435), .ZN(n11437) );
  NOR2_X2 U679 ( .A1(n22529), .A2(n28661), .ZN(n28660) );
  INV_X2 U11248 ( .I(n10946), .ZN(n4228) );
  NAND2_X2 U3102 ( .A1(n21378), .A2(n26798), .ZN(n13621) );
  NOR2_X2 U1618 ( .A1(n18805), .A2(n18806), .ZN(n18807) );
  NAND2_X2 U409 ( .A1(n23684), .A2(n28091), .ZN(n26529) );
  BUF_X2 U5882 ( .I(n9322), .Z(n30755) );
  NAND2_X2 U15593 ( .A1(n18383), .A2(n18515), .ZN(n4206) );
  AOI21_X2 U1251 ( .A1(n15053), .A2(n20243), .B(n26232), .ZN(n20246) );
  NAND2_X1 U18867 ( .A1(n10886), .A2(n8433), .ZN(n11179) );
  INV_X2 U25792 ( .I(n30231), .ZN(n28801) );
  NOR2_X2 U9903 ( .A1(n2391), .A2(n4215), .ZN(n10683) );
  INV_X1 U3114 ( .I(n23087), .ZN(n26243) );
  INV_X1 U3113 ( .I(n20037), .ZN(n28826) );
  INV_X4 U5143 ( .I(n14559), .ZN(n1358) );
  NAND2_X1 U10904 ( .A1(n13914), .A2(n3162), .ZN(n3161) );
  NOR2_X2 U20382 ( .A1(n10964), .A2(n10966), .ZN(n10965) );
  OAI22_X2 U3441 ( .A1(n19365), .A2(n27921), .B1(n19109), .B2(n5907), .ZN(
        n7185) );
  AND2_X2 U471 ( .A1(n13413), .A2(n27883), .Z(n23650) );
  NOR2_X2 U18475 ( .A1(n5248), .A2(n30627), .ZN(n28139) );
  NOR2_X1 U14398 ( .A1(n30318), .A2(n7272), .ZN(n7271) );
  INV_X1 U16031 ( .I(n34108), .ZN(n11182) );
  NAND2_X1 U14732 ( .A1(n27432), .A2(n27431), .ZN(n28652) );
  INV_X1 U11807 ( .I(n17494), .ZN(n24617) );
  NOR2_X2 U13772 ( .A1(n30155), .A2(n20141), .ZN(n15592) );
  OR2_X2 U17578 ( .A1(n6681), .A2(n16756), .Z(n21285) );
  INV_X1 U2069 ( .I(n34110), .ZN(n30697) );
  INV_X2 U22658 ( .I(n3503), .ZN(n28338) );
  NOR2_X1 U14407 ( .A1(n10651), .A2(n24061), .ZN(n10653) );
  NAND2_X1 U5330 ( .A1(n1890), .A2(n30867), .ZN(n4095) );
  INV_X2 U6243 ( .I(n26550), .ZN(n16592) );
  NOR2_X2 U9660 ( .A1(n833), .A2(n24667), .ZN(n28246) );
  INV_X1 U685 ( .I(n21253), .ZN(n17437) );
  INV_X1 U7283 ( .I(n17829), .ZN(n21252) );
  INV_X2 U17043 ( .I(n25582), .ZN(n27637) );
  BUF_X2 U3975 ( .I(n5306), .Z(n2539) );
  CLKBUF_X4 U4053 ( .I(n29470), .Z(n29305) );
  NOR2_X1 U14738 ( .A1(n29018), .A2(n2847), .ZN(n28281) );
  NAND2_X2 U16287 ( .A1(n19124), .A2(n27021), .ZN(n12270) );
  CLKBUF_X4 U4609 ( .I(n19796), .Z(n20052) );
  NAND3_X1 U13428 ( .A1(n15280), .A2(n22838), .A3(n13191), .ZN(n30853) );
  OAI21_X1 U1621 ( .A1(n13760), .A2(n33301), .B(n29983), .ZN(n4535) );
  NOR2_X1 U9597 ( .A1(n12372), .A2(n21121), .ZN(n12371) );
  INV_X2 U18197 ( .I(n31918), .ZN(n27592) );
  INV_X1 U15265 ( .I(n11707), .ZN(n27142) );
  INV_X1 U13160 ( .I(n1577), .ZN(n1581) );
  AOI22_X2 U7359 ( .A1(n870), .A2(n26368), .B1(n16811), .B2(n20044), .ZN(
        n15198) );
  NAND3_X2 U428 ( .A1(n17726), .A2(n16424), .A3(n11960), .ZN(n23835) );
  AOI21_X2 U650 ( .A1(n31712), .A2(n22701), .B(n23081), .ZN(n22704) );
  NAND3_X2 U16686 ( .A1(n30831), .A2(n25600), .A3(n25602), .ZN(n27308) );
  CLKBUF_X4 U4676 ( .I(n17431), .Z(n27560) );
  INV_X4 U23919 ( .I(n16933), .ZN(n21251) );
  INV_X2 U9290 ( .I(n6359), .ZN(n29659) );
  NOR2_X1 U12823 ( .A1(n15098), .A2(n23575), .ZN(n15097) );
  AOI21_X2 U4170 ( .A1(n21686), .A2(n21551), .B(n861), .ZN(n9493) );
  AOI21_X2 U1656 ( .A1(n12699), .A2(n11999), .B(n12651), .ZN(n12650) );
  NOR2_X2 U17431 ( .A1(n9549), .A2(n8422), .ZN(n18369) );
  NOR2_X2 U13658 ( .A1(n32087), .A2(n17132), .ZN(n27008) );
  CLKBUF_X4 U1176 ( .I(n12561), .Z(n26573) );
  NAND2_X1 U11634 ( .A1(n20223), .A2(n2203), .ZN(n2206) );
  NOR2_X1 U9612 ( .A1(n5332), .A2(n29768), .ZN(n30426) );
  INV_X2 U5420 ( .I(n12342), .ZN(n1024) );
  BUF_X2 U1196 ( .I(n7294), .Z(n28983) );
  NAND2_X2 U8576 ( .A1(n14589), .A2(n8611), .ZN(n13571) );
  INV_X1 U4099 ( .I(n7188), .ZN(n12932) );
  NAND2_X2 U930 ( .A1(n16570), .A2(n16556), .ZN(n22560) );
  INV_X2 U22823 ( .I(n34156), .ZN(n7673) );
  AOI21_X2 U21992 ( .A1(n32378), .A2(n22474), .B(n28225), .ZN(n17935) );
  INV_X2 U19914 ( .I(n11637), .ZN(n27901) );
  NOR2_X1 U12833 ( .A1(n26837), .A2(n26836), .ZN(n26835) );
  INV_X1 U19689 ( .I(n9549), .ZN(n18782) );
  NOR2_X1 U11867 ( .A1(n19897), .A2(n33743), .ZN(n15259) );
  BUF_X2 U2092 ( .I(n17405), .Z(n71) );
  INV_X2 U7868 ( .I(n23759), .ZN(n6662) );
  NOR2_X2 U10640 ( .A1(n22478), .A2(n32378), .ZN(n21968) );
  NOR2_X2 U9172 ( .A1(n7088), .A2(n2561), .ZN(n13402) );
  INV_X2 U22916 ( .I(n14572), .ZN(n16595) );
  NAND2_X1 U8533 ( .A1(n26376), .A2(n12892), .ZN(n12891) );
  AOI21_X1 U13509 ( .A1(n2766), .A2(n2767), .B(n31156), .ZN(n30124) );
  OAI21_X2 U14990 ( .A1(n10658), .A2(n17093), .B(n4041), .ZN(n21180) );
  INV_X1 U6361 ( .I(n6569), .ZN(n1131) );
  NAND2_X2 U25352 ( .A1(n23796), .A2(n14193), .ZN(n23803) );
  AOI21_X1 U3984 ( .A1(n19109), .A2(n6566), .B(n6565), .ZN(n6564) );
  NOR3_X2 U1074 ( .A1(n3168), .A2(n5017), .A3(n1325), .ZN(n29737) );
  NOR2_X2 U18582 ( .A1(n7990), .A2(n28701), .ZN(n9560) );
  BUF_X2 U4142 ( .I(n17204), .Z(n6297) );
  AOI22_X2 U7227 ( .A1(n20397), .A2(n7577), .B1(n20396), .B2(n20395), .ZN(
        n26216) );
  OR2_X1 U22434 ( .A1(n18187), .A2(n10080), .Z(n437) );
  AOI21_X1 U534 ( .A1(n12853), .A2(n13490), .B(n12852), .ZN(n12855) );
  NOR2_X2 U19905 ( .A1(n27899), .A2(n10117), .ZN(n10116) );
  OAI21_X2 U23534 ( .A1(n8824), .A2(n8948), .B(n8823), .ZN(n8822) );
  OAI21_X2 U886 ( .A1(n18985), .A2(n18984), .B(n15378), .ZN(n18986) );
  OAI21_X1 U14077 ( .A1(n14667), .A2(n802), .B(n22761), .ZN(n12907) );
  INV_X4 U7322 ( .I(n17157), .ZN(n23878) );
  INV_X4 U12897 ( .I(n15467), .ZN(n17394) );
  INV_X4 U4147 ( .I(n8965), .ZN(n909) );
  NAND2_X2 U24153 ( .A1(n179), .A2(n21438), .ZN(n20330) );
  NOR2_X1 U20022 ( .A1(n30858), .A2(n25084), .ZN(n25087) );
  INV_X2 U5343 ( .I(n13969), .ZN(n13157) );
  NOR2_X2 U23543 ( .A1(n28993), .A2(n31351), .ZN(n7403) );
  NAND2_X2 U3940 ( .A1(n7238), .A2(n349), .ZN(n11153) );
  BUF_X2 U4745 ( .I(n21428), .Z(n26542) );
  INV_X1 U25326 ( .I(n22143), .ZN(n3041) );
  INV_X2 U2613 ( .I(n23942), .ZN(n757) );
  NOR2_X1 U16233 ( .A1(n7344), .A2(n7343), .ZN(n29106) );
  INV_X2 U1518 ( .I(n16309), .ZN(n21867) );
  OAI21_X2 U8963 ( .A1(n5897), .A2(n17787), .B(n15084), .ZN(n16387) );
  NOR2_X1 U4730 ( .A1(n21415), .A2(n21416), .ZN(n27010) );
  NAND2_X2 U1969 ( .A1(n948), .A2(n19078), .ZN(n31539) );
  AOI22_X2 U17809 ( .A1(n18525), .A2(n19256), .B1(n26969), .B2(n33608), .ZN(
        n18527) );
  NAND2_X1 U14353 ( .A1(n4774), .A2(n3421), .ZN(n12576) );
  BUF_X2 U6009 ( .I(Key[115]), .Z(n16472) );
  BUF_X2 U4300 ( .I(Key[66]), .Z(n24623) );
  BUF_X2 U4311 ( .I(Key[145]), .Z(n16680) );
  BUF_X2 U7658 ( .I(Key[98]), .Z(n25208) );
  CLKBUF_X2 U7061 ( .I(Key[111]), .Z(n25610) );
  BUF_X2 U7671 ( .I(Key[97]), .Z(n24991) );
  BUF_X2 U10222 ( .I(Key[175]), .Z(n16381) );
  CLKBUF_X2 U4909 ( .I(Key[144]), .Z(n16575) );
  BUF_X2 U7663 ( .I(Key[106]), .Z(n16602) );
  BUF_X2 U10251 ( .I(Key[92]), .Z(n16671) );
  BUF_X2 U8861 ( .I(Key[19]), .Z(n25071) );
  CLKBUF_X2 U4280 ( .I(Key[33]), .Z(n25722) );
  CLKBUF_X2 U16647 ( .I(n494), .Z(n30371) );
  CLKBUF_X4 U6150 ( .I(n18429), .Z(n18510) );
  INV_X1 U10203 ( .I(n16561), .ZN(n1394) );
  INV_X1 U10198 ( .I(n24804), .ZN(n1410) );
  INV_X1 U508 ( .I(n25476), .ZN(n1404) );
  CLKBUF_X4 U5528 ( .I(n18357), .Z(n18797) );
  CLKBUF_X4 U3412 ( .I(n16596), .Z(n1430) );
  BUF_X2 U15934 ( .I(n18777), .Z(n12863) );
  INV_X1 U25448 ( .I(n31574), .ZN(n28231) );
  CLKBUF_X4 U21786 ( .I(n18392), .Z(n18711) );
  CLKBUF_X2 U12235 ( .I(n18498), .Z(n16435) );
  INV_X2 U8812 ( .I(n17813), .ZN(n5677) );
  CLKBUF_X2 U6094 ( .I(n16249), .Z(n29514) );
  CLKBUF_X4 U15066 ( .I(n17558), .Z(n5327) );
  OAI21_X1 U12168 ( .A1(n18428), .A2(n18832), .B(n18698), .ZN(n17254) );
  INV_X1 U3577 ( .I(n489), .ZN(n958) );
  INV_X1 U16380 ( .I(n19295), .ZN(n15859) );
  NAND2_X1 U12092 ( .A1(n10640), .A2(n10639), .ZN(n7285) );
  INV_X1 U12096 ( .I(n3986), .ZN(n3985) );
  CLKBUF_X4 U1568 ( .I(n2692), .Z(n26603) );
  INV_X2 U10044 ( .I(n31254), .ZN(n1376) );
  BUF_X2 U5168 ( .I(n9553), .Z(n3535) );
  INV_X2 U12701 ( .I(n30039), .ZN(n5610) );
  CLKBUF_X2 U1550 ( .I(n19149), .Z(n25961) );
  CLKBUF_X4 U15279 ( .I(n19335), .Z(n8212) );
  INV_X1 U10070 ( .I(n11477), .ZN(n19326) );
  CLKBUF_X2 U5014 ( .I(n4392), .Z(n29093) );
  BUF_X2 U3278 ( .I(n6763), .Z(n28157) );
  INV_X2 U24058 ( .I(n16801), .ZN(n11444) );
  NOR2_X1 U7775 ( .A1(n19228), .A2(n19357), .ZN(n13389) );
  OAI21_X1 U2698 ( .A1(n1049), .A2(n7687), .B(n11477), .ZN(n11113) );
  AOI21_X1 U23186 ( .A1(n2582), .A2(n30937), .B(n19053), .ZN(n8433) );
  INV_X1 U1912 ( .I(n19323), .ZN(n31618) );
  NOR2_X1 U17052 ( .A1(n18971), .A2(n1177), .ZN(n6024) );
  OAI21_X1 U17184 ( .A1(n27420), .A2(n29245), .B(n19263), .ZN(n9237) );
  AND2_X1 U15100 ( .A1(n18753), .A2(n17339), .Z(n12271) );
  INV_X1 U3417 ( .I(n19013), .ZN(n19010) );
  NOR2_X1 U25845 ( .A1(n19067), .A2(n31618), .ZN(n3133) );
  NAND2_X1 U8257 ( .A1(n30936), .A2(n9839), .ZN(n2583) );
  NAND2_X1 U3480 ( .A1(n4594), .A2(n34040), .ZN(n415) );
  NAND2_X1 U12847 ( .A1(n2598), .A2(n6795), .ZN(n30062) );
  NAND3_X1 U24473 ( .A1(n19352), .A2(n19351), .A3(n19350), .ZN(n19353) );
  CLKBUF_X4 U4969 ( .I(n253), .Z(n28601) );
  BUF_X2 U23579 ( .I(n19672), .Z(n31361) );
  CLKBUF_X4 U7818 ( .I(n30193), .Z(n29515) );
  INV_X1 U24480 ( .I(n19550), .ZN(n19379) );
  INV_X2 U4854 ( .I(n20064), .ZN(n20096) );
  BUF_X2 U5463 ( .I(n20098), .Z(n2606) );
  INV_X1 U22086 ( .I(n13941), .ZN(n19849) );
  BUF_X2 U19175 ( .I(n13922), .Z(n28704) );
  AND2_X1 U4520 ( .A1(n31951), .A2(n10860), .Z(n20153) );
  INV_X1 U841 ( .I(n8421), .ZN(n20032) );
  CLKBUF_X2 U26148 ( .I(n4577), .Z(n31684) );
  NOR2_X1 U1371 ( .A1(n33419), .A2(n16346), .ZN(n27787) );
  CLKBUF_X2 U4610 ( .I(n19419), .Z(n19886) );
  INV_X1 U5459 ( .I(n27748), .ZN(n4441) );
  CLKBUF_X4 U1803 ( .I(n26733), .Z(n30375) );
  CLKBUF_X4 U6430 ( .I(n27748), .Z(n26130) );
  INV_X2 U1417 ( .I(n26733), .ZN(n27938) );
  CLKBUF_X1 U6017 ( .I(n17559), .Z(n29944) );
  CLKBUF_X2 U3952 ( .I(n12241), .Z(n27624) );
  NAND2_X1 U9880 ( .A1(n9031), .A2(n27938), .ZN(n9030) );
  NOR2_X1 U9911 ( .A1(n9748), .A2(n4163), .ZN(n4162) );
  NAND2_X1 U7356 ( .A1(n12119), .A2(n18126), .ZN(n1681) );
  INV_X1 U19159 ( .I(n5470), .ZN(n27788) );
  NAND2_X1 U1347 ( .A1(n9149), .A2(n19840), .ZN(n27764) );
  BUF_X2 U6031 ( .I(n871), .Z(n31103) );
  NAND2_X1 U11817 ( .A1(n6223), .A2(n6221), .ZN(n19898) );
  INV_X1 U16217 ( .I(n570), .ZN(n20095) );
  INV_X1 U11898 ( .I(n19888), .ZN(n4972) );
  CLKBUF_X4 U25900 ( .I(n34153), .Z(n28876) );
  NAND2_X1 U11858 ( .A1(n19798), .A2(n29040), .ZN(n6645) );
  OAI21_X1 U9870 ( .A1(n19990), .A2(n1035), .B(n9661), .ZN(n9660) );
  NAND2_X1 U21584 ( .A1(n7461), .A2(n7460), .ZN(n28153) );
  NAND2_X1 U5977 ( .A1(n20094), .A2(n12669), .ZN(n10926) );
  NAND2_X1 U16811 ( .A1(n19828), .A2(n4587), .ZN(n28209) );
  CLKBUF_X4 U26295 ( .I(n7102), .Z(n31721) );
  NAND2_X1 U21600 ( .A1(n31106), .A2(n28767), .ZN(n27279) );
  OR2_X1 U15592 ( .A1(n4637), .A2(n4636), .Z(n4635) );
  INV_X2 U21598 ( .I(n6444), .ZN(n20078) );
  NAND2_X1 U21583 ( .A1(n28154), .A2(n28153), .ZN(n1976) );
  NAND2_X1 U24325 ( .A1(n31443), .A2(n20154), .ZN(n26543) );
  CLKBUF_X2 U24412 ( .I(n31668), .Z(n31454) );
  NOR2_X1 U5863 ( .A1(n17497), .A2(n26585), .ZN(n17693) );
  CLKBUF_X4 U6303 ( .I(n20560), .Z(n16684) );
  BUF_X1 U15346 ( .I(n9403), .Z(n31156) );
  INV_X1 U10545 ( .I(n28390), .ZN(n29792) );
  CLKBUF_X4 U4416 ( .I(n28064), .Z(n27755) );
  CLKBUF_X4 U8467 ( .I(n20371), .Z(n15898) );
  AOI21_X1 U4897 ( .A1(n27846), .A2(n12351), .B(n12832), .ZN(n2903) );
  CLKBUF_X4 U1706 ( .I(n17544), .Z(n28812) );
  CLKBUF_X4 U5436 ( .I(n16515), .Z(n28085) );
  AND2_X1 U13991 ( .A1(n20395), .A2(n7292), .Z(n7290) );
  NAND2_X1 U18155 ( .A1(n31811), .A2(n20606), .ZN(n20610) );
  OR2_X1 U8036 ( .A1(n15282), .A2(n3944), .Z(n17531) );
  CLKBUF_X2 U7187 ( .I(n12563), .Z(n26343) );
  INV_X2 U15776 ( .I(n9352), .ZN(n13768) );
  INV_X2 U8463 ( .I(n20529), .ZN(n1155) );
  INV_X1 U15811 ( .I(n20288), .ZN(n4964) );
  NOR2_X1 U22262 ( .A1(n17425), .A2(n266), .ZN(n17424) );
  INV_X1 U18863 ( .I(n14683), .ZN(n20251) );
  CLKBUF_X2 U8890 ( .I(n8903), .Z(n29628) );
  INV_X1 U1667 ( .I(n12227), .ZN(n12226) );
  INV_X1 U8452 ( .I(n20604), .ZN(n3751) );
  OAI21_X1 U22416 ( .A1(n1349), .A2(n1351), .B(n11312), .ZN(n31211) );
  NAND2_X1 U9805 ( .A1(n13537), .A2(n9688), .ZN(n13760) );
  NOR2_X1 U11638 ( .A1(n3746), .A2(n17322), .ZN(n4241) );
  OAI21_X1 U1206 ( .A1(n13090), .A2(n20494), .B(n20493), .ZN(n13089) );
  NOR2_X1 U11711 ( .A1(n27020), .A2(n6797), .ZN(n8325) );
  NAND2_X1 U2313 ( .A1(n120), .A2(n20199), .ZN(n1788) );
  NAND2_X1 U11725 ( .A1(n20321), .A2(n1032), .ZN(n10063) );
  INV_X1 U16452 ( .I(n4586), .ZN(n30340) );
  NAND2_X1 U21631 ( .A1(n31112), .A2(n31111), .ZN(n20177) );
  NAND2_X1 U5930 ( .A1(n30464), .A2(n15951), .ZN(n8959) );
  NAND2_X1 U11622 ( .A1(n2206), .A2(n2204), .ZN(n12479) );
  NAND2_X1 U1344 ( .A1(n15257), .A2(n15256), .ZN(n19910) );
  INV_X1 U11690 ( .I(n7978), .ZN(n20580) );
  OAI21_X1 U728 ( .A1(n20230), .A2(n20562), .B(n3352), .ZN(n20233) );
  AOI21_X1 U18510 ( .A1(n30632), .A2(n20493), .B(n17318), .ZN(n16858) );
  NAND2_X1 U9244 ( .A1(n29651), .A2(n26089), .ZN(n30446) );
  CLKBUF_X2 U22344 ( .I(n20900), .Z(n28295) );
  OAI21_X1 U17282 ( .A1(n16758), .A2(n20505), .B(n20504), .ZN(n13092) );
  CLKBUF_X4 U1852 ( .I(n6857), .Z(n15) );
  INV_X1 U11275 ( .I(n29652), .ZN(n20804) );
  CLKBUF_X2 U4201 ( .I(n20913), .Z(n3799) );
  CLKBUF_X4 U3140 ( .I(n7330), .Z(n25969) );
  CLKBUF_X2 U26653 ( .I(n20924), .Z(n31884) );
  INV_X1 U1192 ( .I(n4680), .ZN(n28897) );
  CLKBUF_X2 U22845 ( .I(n12748), .Z(n31277) );
  INV_X1 U4805 ( .I(n20648), .ZN(n26692) );
  INV_X1 U1184 ( .I(n12618), .ZN(n28584) );
  NAND2_X1 U1199 ( .A1(n2649), .A2(n17554), .ZN(n2648) );
  NAND2_X1 U22328 ( .A1(n31189), .A2(n31188), .ZN(n3403) );
  INV_X1 U23585 ( .I(n31423), .ZN(n20979) );
  NAND2_X1 U5883 ( .A1(n30083), .A2(n8579), .ZN(n8578) );
  INV_X2 U23503 ( .I(n17218), .ZN(n16072) );
  BUF_X2 U1481 ( .I(n11733), .Z(n29207) );
  CLKBUF_X2 U7072 ( .I(n21184), .Z(n17466) );
  CLKBUF_X4 U2723 ( .I(n21070), .Z(n164) );
  INV_X1 U5849 ( .I(n9351), .ZN(n9405) );
  CLKBUF_X2 U4792 ( .I(n21454), .Z(n27912) );
  CLKBUF_X4 U5879 ( .I(n4755), .Z(n30988) );
  CLKBUF_X2 U7286 ( .I(n17829), .Z(n28037) );
  CLKBUF_X4 U2502 ( .I(n21232), .Z(n16526) );
  CLKBUF_X4 U3387 ( .I(n11942), .Z(n7430) );
  INV_X2 U7214 ( .I(n16512), .ZN(n922) );
  CLKBUF_X4 U5499 ( .I(n21330), .Z(n8378) );
  INV_X2 U5146 ( .I(n16906), .ZN(n21209) );
  INV_X1 U7152 ( .I(n6192), .ZN(n11487) );
  INV_X1 U24777 ( .I(n21202), .ZN(n20791) );
  OR2_X1 U3996 ( .A1(n12044), .A2(n31114), .Z(n21114) );
  CLKBUF_X4 U7208 ( .I(n515), .Z(n4381) );
  INV_X2 U5529 ( .I(n13255), .ZN(n21211) );
  INV_X1 U21131 ( .I(n21297), .ZN(n15335) );
  NOR2_X1 U20884 ( .A1(n922), .A2(n13582), .ZN(n13581) );
  CLKBUF_X2 U26457 ( .I(n505), .Z(n31760) );
  CLKBUF_X4 U2195 ( .I(n10558), .Z(n4683) );
  NAND2_X1 U18974 ( .A1(n20705), .A2(n12756), .ZN(n30699) );
  INV_X1 U4716 ( .I(n3889), .ZN(n21077) );
  INV_X1 U8340 ( .I(n21398), .ZN(n16755) );
  CLKBUF_X2 U17350 ( .I(n21253), .Z(n27462) );
  CLKBUF_X4 U3043 ( .I(n11063), .Z(n9721) );
  INV_X1 U15576 ( .I(n8041), .ZN(n6826) );
  NAND2_X1 U11442 ( .A1(n6743), .A2(n13896), .ZN(n6501) );
  NAND2_X1 U16200 ( .A1(n7757), .A2(n21259), .ZN(n27246) );
  NAND2_X1 U1316 ( .A1(n30654), .A2(n21093), .ZN(n4919) );
  NOR2_X1 U15982 ( .A1(n12348), .A2(n12017), .ZN(n1687) );
  OR2_X1 U4701 ( .A1(n21176), .A2(n21175), .Z(n26468) );
  NOR2_X1 U9655 ( .A1(n12243), .A2(n1331), .ZN(n10093) );
  NAND2_X1 U7953 ( .A1(n12507), .A2(n10730), .ZN(n26302) );
  NAND2_X1 U18990 ( .A1(n8267), .A2(n21147), .ZN(n12018) );
  BUF_X2 U2874 ( .I(n9472), .Z(n28729) );
  NAND2_X1 U11368 ( .A1(n11152), .A2(n17217), .ZN(n11149) );
  CLKBUF_X2 U13769 ( .I(n21738), .Z(n30154) );
  INV_X1 U9586 ( .I(n2575), .ZN(n21848) );
  CLKBUF_X4 U2109 ( .I(n13113), .Z(n338) );
  NAND2_X1 U1152 ( .A1(n21315), .A2(n8011), .ZN(n9397) );
  INV_X2 U8317 ( .I(n21573), .ZN(n6660) );
  OR2_X1 U3669 ( .A1(n5795), .A2(n6669), .Z(n21660) );
  INV_X1 U5568 ( .I(n21235), .ZN(n4607) );
  CLKBUF_X2 U3915 ( .I(n8313), .Z(n28895) );
  INV_X1 U3037 ( .I(n7182), .ZN(n917) );
  INV_X2 U1764 ( .I(n16987), .ZN(n4234) );
  CLKBUF_X2 U1031 ( .I(n4356), .Z(n28387) );
  CLKBUF_X4 U3401 ( .I(n8790), .Z(n396) );
  BUF_X1 U6613 ( .I(n21761), .Z(n26443) );
  CLKBUF_X4 U4176 ( .I(n6669), .Z(n6483) );
  NAND4_X1 U22307 ( .A1(n13148), .A2(n13150), .A3(n13151), .A4(n13152), .ZN(
        n21786) );
  AND2_X1 U7247 ( .A1(n21779), .A2(n21743), .Z(n29434) );
  INV_X2 U608 ( .I(n21592), .ZN(n21793) );
  CLKBUF_X4 U2944 ( .I(n3539), .Z(n276) );
  INV_X2 U10651 ( .I(n31085), .ZN(n1136) );
  CLKBUF_X4 U15183 ( .I(n5016), .Z(n27619) );
  NAND2_X1 U6556 ( .A1(n1327), .A2(n21707), .ZN(n5788) );
  INV_X1 U3934 ( .I(n21649), .ZN(n16013) );
  NOR2_X1 U13927 ( .A1(n1535), .A2(n21749), .ZN(n1534) );
  AOI21_X1 U1211 ( .A1(n21649), .A2(n21648), .B(n31765), .ZN(n28432) );
  OAI21_X1 U21519 ( .A1(n21683), .A2(n26443), .B(n14870), .ZN(n14869) );
  NAND2_X1 U23265 ( .A1(n1316), .A2(n1319), .ZN(n15413) );
  NAND2_X1 U17466 ( .A1(n913), .A2(n9286), .ZN(n21125) );
  NAND2_X1 U2288 ( .A1(n14730), .A2(n16165), .ZN(n27759) );
  NOR2_X1 U14838 ( .A1(n3048), .A2(n31202), .ZN(n31201) );
  CLKBUF_X2 U10425 ( .I(n11458), .Z(n26562) );
  NAND2_X1 U21710 ( .A1(n12994), .A2(n12995), .ZN(n31118) );
  INV_X1 U1734 ( .I(n28432), .ZN(n28431) );
  NAND2_X1 U18387 ( .A1(n30616), .A2(n26163), .ZN(n275) );
  INV_X2 U893 ( .I(n21913), .ZN(n28162) );
  INV_X2 U12886 ( .I(n26875), .ZN(n8269) );
  CLKBUF_X2 U25966 ( .I(n22149), .Z(n28926) );
  INV_X2 U15748 ( .I(n16893), .ZN(n26957) );
  CLKBUF_X4 U889 ( .I(n22232), .Z(n28730) );
  INV_X1 U14920 ( .I(n7545), .ZN(n8359) );
  INV_X2 U4971 ( .I(n11166), .ZN(n22239) );
  INV_X1 U11220 ( .I(n22144), .ZN(n9311) );
  CLKBUF_X2 U14293 ( .I(n22367), .Z(n30205) );
  INV_X2 U22162 ( .I(n28263), .ZN(n629) );
  OR2_X1 U22049 ( .A1(n9757), .A2(n31692), .Z(n16986) );
  CLKBUF_X2 U3950 ( .I(n16710), .Z(n9022) );
  INV_X2 U6768 ( .I(n628), .ZN(n12496) );
  INV_X2 U6688 ( .I(n31914), .ZN(n22637) );
  CLKBUF_X2 U5804 ( .I(n9871), .Z(n8131) );
  BUF_X4 U5708 ( .I(n14514), .Z(n10354) );
  CLKBUF_X2 U11207 ( .I(n21971), .Z(n22489) );
  AND2_X1 U4474 ( .A1(n9064), .A2(n32055), .Z(n13079) );
  OR2_X1 U2471 ( .A1(n8505), .A2(n6955), .Z(n22475) );
  CLKBUF_X4 U5781 ( .I(n635), .Z(n22557) );
  INV_X1 U2839 ( .I(n16986), .ZN(n26367) );
  BUF_X2 U4568 ( .I(n5657), .Z(n27959) );
  NAND2_X1 U5645 ( .A1(n8912), .A2(n29903), .ZN(n8911) );
  INV_X1 U6343 ( .I(n22683), .ZN(n22686) );
  INV_X2 U13805 ( .I(n2858), .ZN(n22647) );
  NAND2_X1 U960 ( .A1(n22434), .A2(n701), .ZN(n10243) );
  AOI21_X1 U24655 ( .A1(n250), .A2(n5648), .B(n1292), .ZN(n31485) );
  INV_X1 U9812 ( .I(n22657), .ZN(n31267) );
  INV_X1 U2744 ( .I(n30529), .ZN(n11926) );
  AOI21_X1 U903 ( .A1(n32007), .A2(n26046), .B(n17394), .ZN(n29758) );
  INV_X2 U5669 ( .I(n16647), .ZN(n1001) );
  NAND2_X1 U24078 ( .A1(n28592), .A2(n22595), .ZN(n28681) );
  OAI21_X1 U14388 ( .A1(n32042), .A2(n4560), .B(n16334), .ZN(n30215) );
  NAND2_X1 U23023 ( .A1(n10654), .A2(n13525), .ZN(n18062) );
  NOR2_X1 U11051 ( .A1(n11615), .A2(n17631), .ZN(n11614) );
  OAI21_X1 U9960 ( .A1(n29736), .A2(n12840), .B(n22648), .ZN(n27307) );
  OAI21_X1 U19955 ( .A1(n15322), .A2(n11895), .B(n31636), .ZN(n10071) );
  NAND2_X1 U6952 ( .A1(n11243), .A2(n11245), .ZN(n26925) );
  NAND2_X1 U16957 ( .A1(n9108), .A2(n995), .ZN(n6685) );
  INV_X2 U4526 ( .I(n9224), .ZN(n13129) );
  INV_X1 U11672 ( .I(n31854), .ZN(n22849) );
  NAND2_X1 U19382 ( .A1(n22360), .A2(n1298), .ZN(n30762) );
  BUF_X2 U3088 ( .I(n15243), .Z(n27612) );
  BUF_X2 U4422 ( .I(n6798), .Z(n28853) );
  CLKBUF_X2 U5155 ( .I(n22909), .Z(n29328) );
  INV_X2 U22235 ( .I(n23053), .ZN(n28277) );
  NAND2_X1 U3436 ( .A1(n13129), .A2(n22945), .ZN(n31825) );
  INV_X2 U1750 ( .I(n13191), .ZN(n14420) );
  CLKBUF_X4 U777 ( .I(n5696), .Z(n3163) );
  CLKBUF_X4 U744 ( .I(n14126), .Z(n28680) );
  INV_X2 U5352 ( .I(n28942), .ZN(n773) );
  OAI21_X1 U6255 ( .A1(n6782), .A2(n26251), .B(n6942), .ZN(n10107) );
  NOR2_X1 U11027 ( .A1(n14977), .A2(n31867), .ZN(n7528) );
  CLKBUF_X2 U21941 ( .I(n22824), .Z(n28214) );
  BUF_X2 U4451 ( .I(n16297), .Z(n28330) );
  INV_X4 U6268 ( .I(n33675), .ZN(n15851) );
  CLKBUF_X4 U5013 ( .I(n31637), .Z(n29325) );
  OAI21_X1 U10956 ( .A1(n22813), .A2(n4937), .B(n17099), .ZN(n4936) );
  INV_X1 U18838 ( .I(n11383), .ZN(n22853) );
  NOR2_X1 U2506 ( .A1(n32091), .A2(n22919), .ZN(n2775) );
  NAND2_X1 U13339 ( .A1(n1746), .A2(n1745), .ZN(n4155) );
  NAND2_X1 U8039 ( .A1(n27263), .A2(n26312), .ZN(n26960) );
  INV_X1 U4374 ( .I(n27988), .ZN(n27987) );
  INV_X1 U2221 ( .I(n22792), .ZN(n29967) );
  NAND2_X1 U23505 ( .A1(n4487), .A2(n4486), .ZN(n28487) );
  NOR2_X1 U11882 ( .A1(n30968), .A2(n30967), .ZN(n30966) );
  NAND2_X1 U10907 ( .A1(n2078), .A2(n2076), .ZN(n5058) );
  NAND2_X1 U10889 ( .A1(n3778), .A2(n13778), .ZN(n13275) );
  CLKBUF_X2 U2119 ( .I(n5399), .Z(n26915) );
  INV_X1 U11644 ( .I(n23461), .ZN(n30274) );
  NAND2_X1 U4326 ( .A1(n26311), .A2(n26590), .ZN(n27701) );
  INV_X1 U596 ( .I(n23460), .ZN(n2862) );
  INV_X1 U10817 ( .I(n663), .ZN(n23853) );
  CLKBUF_X4 U469 ( .I(n22617), .Z(n27455) );
  CLKBUF_X4 U580 ( .I(n17015), .Z(n14974) );
  BUF_X4 U3504 ( .I(n22936), .Z(n23778) );
  CLKBUF_X4 U15236 ( .I(n665), .Z(n4069) );
  CLKBUF_X4 U2441 ( .I(n661), .Z(n6869) );
  BUF_X2 U15391 ( .I(n23025), .Z(n23775) );
  CLKBUF_X2 U3503 ( .I(n8838), .Z(n313) );
  INV_X2 U4810 ( .I(n23575), .ZN(n23939) );
  CLKBUF_X4 U17418 ( .I(n16534), .Z(n27474) );
  CLKBUF_X2 U483 ( .I(n23719), .Z(n16186) );
  INV_X2 U18798 ( .I(n8251), .ZN(n11240) );
  BUF_X4 U4234 ( .I(n15399), .Z(n1099) );
  NAND2_X1 U5276 ( .A1(n23575), .A2(n15722), .ZN(n12469) );
  INV_X1 U578 ( .I(n14133), .ZN(n1255) );
  NAND2_X1 U445 ( .A1(n23923), .A2(n11192), .ZN(n17543) );
  INV_X2 U262 ( .I(n8270), .ZN(n10145) );
  NAND2_X1 U16796 ( .A1(n979), .A2(n14473), .ZN(n17618) );
  CLKBUF_X4 U3684 ( .I(n15711), .Z(n25987) );
  NAND2_X1 U15843 ( .A1(n23653), .A2(n23746), .ZN(n23777) );
  NAND2_X1 U8874 ( .A1(n16186), .A2(n6869), .ZN(n8372) );
  INV_X2 U6879 ( .I(n11240), .ZN(n16388) );
  OR2_X1 U15293 ( .A1(n23899), .A2(n32711), .Z(n23704) );
  INV_X2 U22620 ( .I(n15623), .ZN(n16343) );
  CLKBUF_X4 U16075 ( .I(n23945), .Z(n27219) );
  NOR2_X1 U16018 ( .A1(n12848), .A2(n8045), .ZN(n27049) );
  NAND2_X1 U14330 ( .A1(n16212), .A2(n16211), .ZN(n28698) );
  NAND2_X1 U17524 ( .A1(n7141), .A2(n7139), .ZN(n23565) );
  NAND2_X1 U6846 ( .A1(n17950), .A2(n17949), .ZN(n3919) );
  AOI21_X1 U21070 ( .A1(n23955), .A2(n15616), .B(n23824), .ZN(n14014) );
  AOI21_X1 U6140 ( .A1(n18054), .A2(n9225), .B(n28855), .ZN(n24001) );
  AND2_X1 U13749 ( .A1(n23353), .A2(n17088), .Z(n29124) );
  OAI21_X1 U9132 ( .A1(n12433), .A2(n978), .B(n15351), .ZN(n17490) );
  NAND2_X1 U10764 ( .A1(n12592), .A2(n7781), .ZN(n7780) );
  AND2_X1 U6159 ( .A1(n16947), .A2(n7524), .Z(n14907) );
  NAND2_X1 U2325 ( .A1(n23308), .A2(n12603), .ZN(n12602) );
  INV_X2 U186 ( .I(n24201), .ZN(n738) );
  NOR2_X1 U15711 ( .A1(n12974), .A2(n5373), .ZN(n7407) );
  NAND2_X1 U21849 ( .A1(n845), .A2(n8914), .ZN(n3014) );
  INV_X1 U4094 ( .I(n10384), .ZN(n7169) );
  NAND2_X1 U10688 ( .A1(n13138), .A2(n13136), .ZN(n8380) );
  CLKBUF_X2 U5544 ( .I(n24240), .Z(n31862) );
  CLKBUF_X2 U2791 ( .I(n13623), .Z(n11255) );
  CLKBUF_X2 U12841 ( .I(n6286), .Z(n30061) );
  BUF_X2 U20942 ( .I(n3421), .Z(n31002) );
  BUF_X2 U3204 ( .I(n9919), .Z(n2444) );
  INV_X2 U246 ( .I(n24309), .ZN(n28040) );
  INV_X1 U3656 ( .I(n15227), .ZN(n24051) );
  NAND2_X1 U10587 ( .A1(n23608), .A2(n794), .ZN(n3861) );
  CLKBUF_X1 U5489 ( .I(n9146), .Z(n29819) );
  CLKBUF_X4 U15888 ( .I(n24053), .Z(n10381) );
  CLKBUF_X4 U258 ( .I(n11438), .Z(n28691) );
  NAND2_X1 U7758 ( .A1(n5914), .A2(n13260), .ZN(n3255) );
  CLKBUF_X4 U12931 ( .I(n16643), .Z(n8086) );
  AOI21_X1 U3549 ( .A1(n7099), .A2(n24246), .B(n28538), .ZN(n7098) );
  INV_X1 U10561 ( .I(n14052), .ZN(n8263) );
  NAND2_X1 U17209 ( .A1(n13239), .A2(n13109), .ZN(n13238) );
  AND3_X1 U15427 ( .A1(n6773), .A2(n7729), .A3(n7727), .Z(n27157) );
  OAI21_X1 U11409 ( .A1(n17566), .A2(n33182), .B(n305), .ZN(n5000) );
  NAND2_X1 U8546 ( .A1(n2398), .A2(n2400), .ZN(n29924) );
  CLKBUF_X4 U3025 ( .I(n9300), .Z(n4997) );
  NAND3_X1 U17062 ( .A1(n24502), .A2(n24500), .A3(n24501), .ZN(n30822) );
  CLKBUF_X4 U277 ( .I(n9708), .Z(n29320) );
  CLKBUF_X2 U13307 ( .I(n5762), .Z(n30104) );
  BUF_X2 U3379 ( .I(n24359), .Z(n13050) );
  INV_X1 U4059 ( .I(n9120), .ZN(n12676) );
  BUF_X2 U3645 ( .I(n17117), .Z(n15046) );
  BUF_X4 U15256 ( .I(n24368), .Z(n25707) );
  CLKBUF_X2 U4038 ( .I(n678), .Z(n28958) );
  BUF_X2 U4055 ( .I(n25188), .Z(n28591) );
  BUF_X2 U3221 ( .I(n25242), .Z(n25977) );
  CLKBUF_X2 U14574 ( .I(n29278), .Z(n30241) );
  INV_X2 U25820 ( .I(n24974), .ZN(n28815) );
  CLKBUF_X4 U23584 ( .I(n25150), .Z(n16293) );
  CLKBUF_X4 U5260 ( .I(n16659), .Z(n29334) );
  CLKBUF_X4 U156 ( .I(n13427), .Z(n1567) );
  CLKBUF_X2 U4037 ( .I(n25200), .Z(n26432) );
  INV_X2 U23995 ( .I(n32652), .ZN(n25025) );
  NOR2_X1 U1946 ( .A1(n32872), .A2(n2642), .ZN(n27757) );
  NAND2_X1 U8943 ( .A1(n25868), .A2(n11716), .ZN(n10066) );
  NOR2_X1 U14510 ( .A1(n10890), .A2(n32760), .ZN(n11082) );
  NAND2_X1 U3586 ( .A1(n836), .A2(n11045), .ZN(n24723) );
  NAND2_X1 U16312 ( .A1(n10454), .A2(n25566), .ZN(n27269) );
  NOR2_X1 U5320 ( .A1(n30877), .A2(n30876), .ZN(n31109) );
  NAND2_X1 U21630 ( .A1(n3955), .A2(n24413), .ZN(n31110) );
  CLKBUF_X4 U7042 ( .I(n17637), .Z(n30935) );
  BUF_X2 U4309 ( .I(Key[69]), .Z(n25911) );
  BUF_X2 U8859 ( .I(Key[183]), .Z(n16672) );
  BUF_X2 U7666 ( .I(Key[75]), .Z(n25364) );
  CLKBUF_X2 U4296 ( .I(Key[110]), .Z(n25274) );
  BUF_X2 U6005 ( .I(Key[121]), .Z(n25091) );
  CLKBUF_X2 U2282 ( .I(Key[51]), .Z(n23239) );
  CLKBUF_X2 U10244 ( .I(Key[18]), .Z(n16464) );
  BUF_X2 U4285 ( .I(Key[7]), .Z(n24999) );
  BUF_X2 U4649 ( .I(Key[72]), .Z(n24804) );
  CLKBUF_X2 U6122 ( .I(n18860), .Z(n31417) );
  INV_X1 U24564 ( .I(n19718), .ZN(n25104) );
  CLKBUF_X2 U12211 ( .I(n18773), .Z(n16522) );
  CLKBUF_X2 U2065 ( .I(n18228), .Z(n30472) );
  CLKBUF_X4 U1048 ( .I(n18884), .Z(n10669) );
  NOR2_X1 U10121 ( .A1(n18653), .A2(n31542), .ZN(n10640) );
  OAI21_X1 U10102 ( .A1(n18796), .A2(n18795), .B(n18799), .ZN(n3986) );
  NAND2_X1 U16024 ( .A1(n10220), .A2(n31972), .ZN(n8645) );
  BUF_X2 U6064 ( .I(n18257), .Z(n29715) );
  AND2_X1 U24266 ( .A1(n19322), .A2(n19274), .Z(n18415) );
  CLKBUF_X1 U21526 ( .I(n19224), .Z(n28147) );
  CLKBUF_X1 U6236 ( .I(n19053), .Z(n31108) );
  CLKBUF_X2 U3021 ( .I(n19149), .Z(n25960) );
  CLKBUF_X4 U20331 ( .I(n2971), .Z(n27965) );
  BUF_X2 U3969 ( .I(n27242), .Z(n26350) );
  CLKBUF_X2 U5004 ( .I(n18626), .Z(n28478) );
  OAI21_X1 U3133 ( .A1(n32790), .A2(n19137), .B(n744), .ZN(n4594) );
  NAND2_X1 U24444 ( .A1(n19189), .A2(n19257), .ZN(n19190) );
  NAND2_X1 U4992 ( .A1(n5082), .A2(n4405), .ZN(n5083) );
  CLKBUF_X2 U9910 ( .I(n18109), .Z(n29728) );
  NOR2_X1 U11956 ( .A1(n3073), .A2(n6575), .ZN(n3072) );
  CLKBUF_X2 U4957 ( .I(n29254), .Z(n29013) );
  BUF_X2 U6033 ( .I(n18199), .Z(n28183) );
  CLKBUF_X4 U1867 ( .I(n27808), .Z(n31823) );
  INV_X2 U4216 ( .I(n17495), .ZN(n939) );
  NOR2_X1 U19604 ( .A1(n8616), .A2(n19451), .ZN(n9379) );
  NAND2_X1 U24583 ( .A1(n1168), .A2(n10340), .ZN(n19823) );
  NAND2_X1 U17250 ( .A1(n27938), .A2(n13994), .ZN(n19805) );
  BUF_X2 U1831 ( .I(n20113), .Z(n31715) );
  INV_X2 U7390 ( .I(n15192), .ZN(n6644) );
  CLKBUF_X4 U5985 ( .I(n27070), .Z(n29603) );
  CLKBUF_X2 U3941 ( .I(n20614), .Z(n28527) );
  CLKBUF_X2 U5394 ( .I(n20634), .Z(n2203) );
  INV_X2 U3939 ( .I(n20634), .ZN(n20379) );
  CLKBUF_X2 U3492 ( .I(n816), .Z(n420) );
  NAND2_X1 U5936 ( .A1(n20258), .A2(n29603), .ZN(n29994) );
  CLKBUF_X4 U2847 ( .I(n10717), .Z(n1863) );
  BUF_X2 U5942 ( .I(n4460), .Z(n30793) );
  NOR2_X1 U1644 ( .A1(n20442), .A2(n1032), .ZN(n30952) );
  NAND2_X1 U4492 ( .A1(n1032), .A2(n18078), .ZN(n28135) );
  CLKBUF_X4 U1730 ( .I(n9831), .Z(n9688) );
  OAI21_X1 U26483 ( .A1(n4964), .A2(n31776), .B(n20174), .ZN(n27611) );
  BUF_X2 U4060 ( .I(n8625), .Z(n5141) );
  CLKBUF_X2 U2085 ( .I(n601), .Z(n67) );
  CLKBUF_X2 U5872 ( .I(n21168), .Z(n31874) );
  CLKBUF_X1 U1497 ( .I(n27503), .Z(n27773) );
  BUF_X4 U2729 ( .I(n16784), .Z(n28642) );
  CLKBUF_X4 U4190 ( .I(n18110), .Z(n6408) );
  NAND2_X2 U5856 ( .A1(n810), .A2(n27773), .ZN(n21366) );
  NOR2_X1 U1149 ( .A1(n21267), .A2(n31965), .ZN(n28922) );
  NOR2_X1 U8230 ( .A1(n12756), .A2(n810), .ZN(n12017) );
  OAI21_X1 U4734 ( .A1(n21138), .A2(n1553), .B(n9699), .ZN(n28754) );
  INV_X2 U1254 ( .I(n26622), .ZN(n21755) );
  INV_X1 U9651 ( .I(n26494), .ZN(n21153) );
  CLKBUF_X2 U4675 ( .I(n13442), .Z(n26163) );
  CLKBUF_X2 U14975 ( .I(n21849), .Z(n13490) );
  CLKBUF_X2 U5827 ( .I(n21573), .Z(n29552) );
  CLKBUF_X2 U4166 ( .I(n15863), .Z(n3821) );
  BUF_X2 U4171 ( .I(n12866), .Z(n15655) );
  NAND2_X1 U998 ( .A1(n5383), .A2(n5494), .ZN(n12391) );
  NAND2_X1 U22461 ( .A1(n7182), .A2(n196), .ZN(n5850) );
  INV_X2 U9582 ( .I(n4097), .ZN(n16165) );
  INV_X1 U5552 ( .I(n4356), .ZN(n21560) );
  NAND2_X1 U18339 ( .A1(n30978), .A2(n11301), .ZN(n3680) );
  NOR2_X1 U14323 ( .A1(n7476), .A2(n21854), .ZN(n27065) );
  BUF_X2 U21579 ( .I(n6442), .Z(n31102) );
  INV_X1 U15941 ( .I(n21749), .ZN(n1532) );
  OAI22_X1 U8120 ( .A1(n16723), .A2(n1134), .B1(n21283), .B2(n1312), .ZN(
        n16722) );
  NAND2_X1 U18390 ( .A1(n21839), .A2(n21685), .ZN(n30616) );
  NAND2_X1 U21177 ( .A1(n21591), .A2(n3756), .ZN(n15846) );
  INV_X1 U11964 ( .I(n21717), .ZN(n26732) );
  NAND2_X1 U21734 ( .A1(n21247), .A2(n31121), .ZN(n27753) );
  CLKBUF_X4 U3892 ( .I(n9129), .Z(n343) );
  INV_X1 U14540 ( .I(n12789), .ZN(n13146) );
  INV_X2 U5716 ( .I(n32753), .ZN(n29951) );
  CLKBUF_X2 U4547 ( .I(n17151), .Z(n27415) );
  INV_X2 U9436 ( .I(n16627), .ZN(n22434) );
  CLKBUF_X1 U16980 ( .I(n10183), .Z(n30405) );
  INV_X2 U2967 ( .I(n22926), .ZN(n22657) );
  BUF_X2 U762 ( .I(n29287), .Z(n16334) );
  INV_X2 U3173 ( .I(n4425), .ZN(n12043) );
  NAND2_X1 U4498 ( .A1(n33283), .A2(n994), .ZN(n27495) );
  OAI21_X1 U16505 ( .A1(n22434), .A2(n11895), .B(n28473), .ZN(n14329) );
  NOR2_X1 U25077 ( .A1(n22550), .A2(n15260), .ZN(n22392) );
  NAND3_X1 U6298 ( .A1(n15322), .A2(n11895), .A3(n22435), .ZN(n12688) );
  NAND3_X1 U4527 ( .A1(n22200), .A2(n8519), .A3(n31636), .ZN(n3384) );
  BUF_X4 U3565 ( .I(n15501), .Z(n29070) );
  BUF_X2 U7168 ( .I(n28942), .Z(n26251) );
  BUF_X2 U6955 ( .I(n6874), .Z(n3657) );
  BUF_X2 U697 ( .I(n23065), .Z(n4067) );
  BUF_X2 U6795 ( .I(n15123), .Z(n28313) );
  CLKBUF_X1 U20492 ( .I(n31854), .Z(n30925) );
  CLKBUF_X1 U4065 ( .I(n2449), .Z(n30455) );
  BUF_X2 U5644 ( .I(n15324), .Z(n26526) );
  OAI21_X1 U6837 ( .A1(n23096), .A2(n22786), .B(n18261), .ZN(n3297) );
  CLKBUF_X1 U2272 ( .I(n4124), .Z(n28849) );
  NOR2_X1 U10961 ( .A1(n22781), .A2(n29173), .ZN(n11741) );
  AOI21_X1 U2990 ( .A1(n28348), .A2(n28349), .B(n22720), .ZN(n5345) );
  NAND2_X1 U14187 ( .A1(n13004), .A2(n28853), .ZN(n13003) );
  BUF_X1 U24011 ( .I(n27175), .Z(n23238) );
  BUF_X2 U16177 ( .I(n23171), .Z(n27243) );
  CLKBUF_X4 U584 ( .I(n23916), .Z(n23721) );
  BUF_X2 U3223 ( .I(n29270), .Z(n354) );
  INV_X1 U6217 ( .I(n29271), .ZN(n895) );
  CLKBUF_X2 U4470 ( .I(n14031), .Z(n28273) );
  OAI21_X1 U6880 ( .A1(n11821), .A2(n8408), .B(n10142), .ZN(n13224) );
  BUF_X2 U410 ( .I(n17872), .Z(n6392) );
  OAI21_X1 U332 ( .A1(n31071), .A2(n13600), .B(n32520), .ZN(n31872) );
  CLKBUF_X1 U13696 ( .I(n24096), .Z(n30146) );
  OR2_X1 U9539 ( .A1(n24177), .A2(n15720), .Z(n14052) );
  NAND2_X1 U5520 ( .A1(n1092), .A2(n31342), .ZN(n31341) );
  AOI21_X1 U25164 ( .A1(n15537), .A2(n15899), .B(n28726), .ZN(n28725) );
  NAND2_X1 U5465 ( .A1(n31341), .A2(n29949), .ZN(n28522) );
  CLKBUF_X2 U2526 ( .I(n9353), .Z(n30358) );
  AND2_X1 U15900 ( .A1(n25628), .A2(n17523), .Z(n12926) );
  OR2_X1 U9006 ( .A1(n17641), .A2(n34169), .Z(n25566) );
  CLKBUF_X1 U2960 ( .I(n25277), .Z(n298) );
  AOI21_X1 U13184 ( .A1(n1205), .A2(n42), .B(n2264), .ZN(n2263) );
  NOR2_X1 U8145 ( .A1(n18034), .A2(n28923), .ZN(n18033) );
  INV_X2 U5395 ( .I(n20227), .ZN(n3972) );
  INV_X2 U20867 ( .I(n4119), .ZN(n21200) );
  INV_X2 U6301 ( .I(n19779), .ZN(n19434) );
  NOR2_X2 U105 ( .A1(n24725), .A2(n12699), .ZN(n12651) );
  OAI21_X2 U11678 ( .A1(n4468), .A2(n8998), .B(n12516), .ZN(n12515) );
  INV_X2 U6471 ( .I(n20385), .ZN(n12514) );
  BUF_X4 U15300 ( .I(n24823), .Z(n4240) );
  BUF_X4 U5953 ( .I(n17820), .Z(n3388) );
  INV_X4 U15203 ( .I(n5889), .ZN(n19063) );
  INV_X4 U8492 ( .I(n20384), .ZN(n8998) );
  AOI21_X2 U634 ( .A1(n21374), .A2(n4145), .B(n32452), .ZN(n21141) );
  AOI22_X2 U641 ( .A1(n27410), .A2(n27409), .B1(n17212), .B2(n29635), .ZN(
        n7584) );
  OAI21_X2 U9905 ( .A1(n939), .A2(n16489), .B(n4938), .ZN(n19438) );
  BUF_X4 U2684 ( .I(n25973), .Z(n25974) );
  BUF_X4 U16038 ( .I(n15212), .Z(n31263) );
  AOI21_X2 U3098 ( .A1(n24317), .A2(n14112), .B(n2913), .ZN(n9892) );
  NOR2_X2 U6590 ( .A1(n19259), .A2(n28379), .ZN(n6342) );
  BUF_X4 U594 ( .I(n17929), .Z(n26582) );
  NAND3_X2 U3414 ( .A1(n31381), .A2(n25821), .A3(n18246), .ZN(n8345) );
  NOR2_X2 U21542 ( .A1(n3183), .A2(n31824), .ZN(n22740) );
  NAND2_X1 U19079 ( .A1(n17578), .A2(n23874), .ZN(n23875) );
  NAND3_X2 U17316 ( .A1(n2128), .A2(n3006), .A3(n1934), .ZN(n30837) );
  INV_X4 U3866 ( .I(n31824), .ZN(n29173) );
  OAI21_X2 U21587 ( .A1(n831), .A2(n27262), .B(n25607), .ZN(n25600) );
  NOR2_X1 U6619 ( .A1(n4494), .A2(n27539), .ZN(n26152) );
  INV_X4 U8607 ( .I(n19926), .ZN(n20149) );
  OAI21_X2 U16275 ( .A1(n24152), .A2(n24154), .B(n27259), .ZN(n24066) );
  NOR2_X2 U8432 ( .A1(n29583), .A2(n6216), .ZN(n30122) );
  NOR2_X1 U4158 ( .A1(n300), .A2(n13263), .ZN(n13262) );
  INV_X2 U5519 ( .I(n29087), .ZN(n18571) );
  INV_X1 U17233 ( .I(n27428), .ZN(n12006) );
  NOR2_X1 U6147 ( .A1(n18639), .A2(n18815), .ZN(n18383) );
  NAND2_X1 U21163 ( .A1(n18633), .A2(n18710), .ZN(n16295) );
  INV_X1 U10456 ( .I(n29776), .ZN(n27958) );
  INV_X1 U22552 ( .I(n28321), .ZN(n14926) );
  INV_X2 U8805 ( .I(n18737), .ZN(n17360) );
  INV_X1 U984 ( .I(n18862), .ZN(n18738) );
  NOR2_X1 U26412 ( .A1(n15811), .A2(n27142), .ZN(n31748) );
  CLKBUF_X2 U3453 ( .I(n495), .Z(n46) );
  BUF_X2 U1639 ( .I(n18874), .Z(n16538) );
  NOR2_X1 U987 ( .A1(n1659), .A2(n5700), .ZN(n18400) );
  INV_X1 U7471 ( .I(n26249), .ZN(n18018) );
  INV_X1 U5185 ( .I(n962), .ZN(n6891) );
  INV_X1 U5120 ( .I(n18586), .ZN(n17166) );
  INV_X1 U6722 ( .I(n13719), .ZN(n8739) );
  BUF_X2 U7649 ( .I(n10664), .Z(n5269) );
  INV_X1 U6703 ( .I(n18756), .ZN(n18602) );
  INV_X1 U7650 ( .I(n18580), .ZN(n17419) );
  INV_X2 U6711 ( .I(n18722), .ZN(n18727) );
  OR2_X1 U12190 ( .A1(n490), .A2(n18723), .Z(n18584) );
  NOR2_X1 U975 ( .A1(n29182), .A2(n18727), .ZN(n11164) );
  INV_X1 U6701 ( .I(n7216), .ZN(n1853) );
  INV_X2 U6668 ( .I(n15873), .ZN(n1059) );
  NOR2_X1 U24350 ( .A1(n28675), .A2(n18687), .ZN(n18691) );
  INV_X1 U1009 ( .I(n15519), .ZN(n959) );
  NOR2_X1 U20742 ( .A1(n18559), .A2(n18623), .ZN(n18328) );
  NAND2_X1 U7624 ( .A1(n882), .A2(n11097), .ZN(n12876) );
  NOR2_X1 U23918 ( .A1(n882), .A2(n30472), .ZN(n17422) );
  NOR2_X1 U15509 ( .A1(n3954), .A2(n8386), .ZN(n18653) );
  NOR2_X1 U22518 ( .A1(n18815), .A2(n13663), .ZN(n18816) );
  INV_X2 U8806 ( .I(n15902), .ZN(n18875) );
  NAND2_X1 U10184 ( .A1(n18710), .A2(n18711), .ZN(n11270) );
  NOR2_X1 U10751 ( .A1(n15888), .A2(n32337), .ZN(n17190) );
  NAND2_X1 U12165 ( .A1(n16393), .A2(n13663), .ZN(n8735) );
  INV_X1 U10165 ( .I(n15211), .ZN(n18856) );
  INV_X2 U5522 ( .I(n18743), .ZN(n16358) );
  NAND2_X1 U24363 ( .A1(n18288), .A2(n27940), .ZN(n18760) );
  INV_X2 U7616 ( .I(n18774), .ZN(n18556) );
  INV_X1 U10208 ( .I(n16249), .ZN(n1186) );
  NAND2_X1 U8823 ( .A1(n18849), .A2(n18845), .ZN(n6312) );
  NOR2_X1 U5967 ( .A1(n5834), .A2(n18681), .ZN(n4926) );
  INV_X1 U14717 ( .I(n16915), .ZN(n6256) );
  INV_X1 U4901 ( .I(n490), .ZN(n11123) );
  INV_X1 U1608 ( .I(n488), .ZN(n1185) );
  NOR2_X1 U1822 ( .A1(n14651), .A2(n18638), .ZN(n14344) );
  INV_X1 U12151 ( .I(n9667), .ZN(n3018) );
  AND2_X1 U16367 ( .A1(n15966), .A2(n17030), .Z(n18733) );
  INV_X1 U2830 ( .I(n13445), .ZN(n18511) );
  INV_X1 U16157 ( .I(n18581), .ZN(n18726) );
  INV_X1 U3389 ( .I(n18487), .ZN(n18829) );
  OR2_X1 U2809 ( .A1(n15216), .A2(n15347), .Z(n18579) );
  NAND2_X1 U7551 ( .A1(n18288), .A2(n33472), .ZN(n18603) );
  NOR3_X1 U5029 ( .A1(n18881), .A2(n18880), .A3(n16588), .ZN(n10637) );
  NAND2_X1 U2836 ( .A1(n180), .A2(n18493), .ZN(n18326) );
  NAND2_X1 U8773 ( .A1(n5269), .A2(n18746), .ZN(n14705) );
  INV_X1 U6156 ( .I(n18579), .ZN(n6873) );
  NAND2_X1 U15658 ( .A1(n4259), .A2(n31579), .ZN(n18277) );
  NAND2_X1 U20416 ( .A1(n11164), .A2(n12320), .ZN(n11023) );
  NAND2_X1 U14039 ( .A1(n951), .A2(n8570), .ZN(n5646) );
  NOR2_X1 U12608 ( .A1(n15902), .A2(n10181), .ZN(n1710) );
  NOR2_X1 U26256 ( .A1(n16393), .A2(n18815), .ZN(n6393) );
  INV_X1 U1622 ( .I(n28438), .ZN(n18578) );
  INV_X1 U2006 ( .I(n18604), .ZN(n30181) );
  NOR2_X1 U19820 ( .A1(n10964), .A2(n12120), .ZN(n15136) );
  NOR2_X1 U7438 ( .A1(n31972), .A2(n28675), .ZN(n13860) );
  NAND2_X1 U14734 ( .A1(n1059), .A2(n9651), .ZN(n30255) );
  INV_X2 U7645 ( .I(n16474), .ZN(n17465) );
  NOR2_X1 U4891 ( .A1(n13014), .A2(n13013), .ZN(n18921) );
  INV_X1 U8781 ( .I(n18880), .ZN(n18112) );
  NOR2_X1 U10168 ( .A1(n16564), .A2(n18770), .ZN(n18495) );
  NAND2_X1 U3167 ( .A1(n18617), .A2(n16948), .ZN(n2042) );
  INV_X1 U4650 ( .I(n26040), .ZN(n732) );
  INV_X1 U24291 ( .I(n18563), .ZN(n18464) );
  AND2_X1 U12401 ( .A1(n18874), .A2(n27311), .Z(n14658) );
  INV_X1 U8813 ( .I(n34139), .ZN(n18566) );
  OAI21_X1 U23513 ( .A1(n18880), .A2(n16572), .B(n16588), .ZN(n16109) );
  NOR2_X1 U22172 ( .A1(n31972), .A2(n10283), .ZN(n18399) );
  AOI22_X1 U6168 ( .A1(n18543), .A2(n18854), .B1(n18307), .B2(n18853), .ZN(
        n18308) );
  NOR2_X1 U5971 ( .A1(n2042), .A2(n17224), .ZN(n6298) );
  OAI21_X1 U21153 ( .A1(n18553), .A2(n15694), .B(n28548), .ZN(n15693) );
  OAI22_X1 U992 ( .A1(n3436), .A2(n1853), .B1(n3437), .B2(n956), .ZN(n17131)
         );
  AOI21_X1 U20188 ( .A1(n31724), .A2(n6119), .B(n17843), .ZN(n18447) );
  NOR2_X1 U950 ( .A1(n13548), .A2(n26810), .ZN(n10125) );
  NOR2_X1 U6191 ( .A1(n18496), .A2(n10043), .ZN(n6666) );
  NOR2_X1 U18796 ( .A1(n18880), .A2(n16466), .ZN(n15984) );
  INV_X1 U1617 ( .I(n6138), .ZN(n26680) );
  NAND2_X1 U1596 ( .A1(n11097), .A2(n14213), .ZN(n26320) );
  NAND2_X1 U24225 ( .A1(n7454), .A2(n13514), .ZN(n18362) );
  NOR2_X1 U2049 ( .A1(n18643), .A2(n16766), .ZN(n31369) );
  NAND2_X1 U20825 ( .A1(n18817), .A2(n18714), .ZN(n16088) );
  NOR2_X1 U24326 ( .A1(n18584), .A2(n29602), .ZN(n18585) );
  NAND2_X1 U12130 ( .A1(n10565), .A2(n18574), .ZN(n10564) );
  AOI22_X1 U10120 ( .A1(n6393), .A2(n829), .B1(n18515), .B2(n7977), .ZN(n4114)
         );
  NOR3_X1 U20817 ( .A1(n13566), .A2(n18633), .A3(n1439), .ZN(n13565) );
  NAND2_X1 U14729 ( .A1(n16867), .A2(n30255), .ZN(n11470) );
  NAND2_X1 U24307 ( .A1(n33783), .A2(n18633), .ZN(n18508) );
  AOI22_X1 U6208 ( .A1(n10095), .A2(n18812), .B1(n18893), .B2(n27228), .ZN(
        n27618) );
  INV_X2 U3460 ( .I(n29223), .ZN(n1046) );
  NAND3_X1 U10132 ( .A1(n18516), .A2(n1572), .A3(n33548), .ZN(n14660) );
  INV_X1 U2007 ( .I(n18939), .ZN(n30958) );
  BUF_X2 U4241 ( .I(n16748), .Z(n13390) );
  INV_X2 U2535 ( .I(n16047), .ZN(n19088) );
  INV_X1 U5495 ( .I(n13673), .ZN(n19120) );
  INV_X1 U24384 ( .I(n19006), .ZN(n18876) );
  INV_X1 U4603 ( .I(n19325), .ZN(n19105) );
  NAND2_X1 U6184 ( .A1(n19267), .A2(n19265), .ZN(n19225) );
  NAND2_X1 U12364 ( .A1(n11477), .A2(n10714), .ZN(n19183) );
  INV_X1 U1986 ( .I(n8800), .ZN(n31152) );
  NAND2_X1 U6233 ( .A1(n5760), .A2(n18988), .ZN(n5761) );
  INV_X1 U8685 ( .I(n19089), .ZN(n6510) );
  INV_X1 U21808 ( .I(n19115), .ZN(n13329) );
  BUF_X2 U1147 ( .I(n14198), .Z(n6516) );
  INV_X2 U934 ( .I(n29757), .ZN(n1180) );
  INV_X2 U5009 ( .I(n19285), .ZN(n19078) );
  INV_X2 U5498 ( .I(n10974), .ZN(n10203) );
  INV_X1 U5479 ( .I(n19199), .ZN(n19093) );
  INV_X1 U15405 ( .I(n19049), .ZN(n949) );
  INV_X1 U3967 ( .I(n19167), .ZN(n824) );
  INV_X1 U14584 ( .I(n10714), .ZN(n1049) );
  INV_X1 U5955 ( .I(n2692), .ZN(n2901) );
  INV_X1 U21867 ( .I(n28197), .ZN(n15239) );
  INV_X1 U3180 ( .I(n19104), .ZN(n944) );
  INV_X1 U14351 ( .I(n8379), .ZN(n1054) );
  INV_X1 U920 ( .I(n8141), .ZN(n17386) );
  INV_X1 U8697 ( .I(n19265), .ZN(n2101) );
  INV_X2 U1938 ( .I(n29769), .ZN(n19179) );
  NAND2_X1 U15846 ( .A1(n25968), .A2(n8787), .ZN(n19114) );
  INV_X1 U12085 ( .I(n19274), .ZN(n19321) );
  NAND2_X1 U10014 ( .A1(n19248), .A2(n1050), .ZN(n5082) );
  NAND2_X1 U6229 ( .A1(n949), .A2(n19048), .ZN(n12708) );
  OAI21_X1 U21162 ( .A1(n27743), .A2(n29525), .B(n12500), .ZN(n12831) );
  NAND2_X1 U6620 ( .A1(n19158), .A2(n14811), .ZN(n19112) );
  NOR2_X1 U21465 ( .A1(n19357), .A2(n14624), .ZN(n16749) );
  NOR2_X1 U8681 ( .A1(n13390), .A2(n19228), .ZN(n18068) );
  NAND2_X1 U1950 ( .A1(n26891), .A2(n10700), .ZN(n13226) );
  INV_X1 U2999 ( .I(n19101), .ZN(n19009) );
  NOR2_X1 U9339 ( .A1(n880), .A2(n950), .ZN(n2039) );
  OR2_X1 U22149 ( .A1(n4747), .A2(n30879), .Z(n5653) );
  NOR2_X1 U7485 ( .A1(n17445), .A2(n7995), .ZN(n11714) );
  INV_X1 U12017 ( .I(n19100), .ZN(n11715) );
  OAI21_X1 U20393 ( .A1(n26830), .A2(n6516), .B(n19228), .ZN(n16768) );
  CLKBUF_X2 U21360 ( .I(n26969), .Z(n31074) );
  BUF_X2 U25977 ( .I(n19104), .Z(n28935) );
  NAND2_X1 U21560 ( .A1(n1380), .A2(n19222), .ZN(n12468) );
  NAND2_X1 U5238 ( .A1(n19318), .A2(n19319), .ZN(n19317) );
  NAND3_X1 U17411 ( .A1(n19040), .A2(n19049), .A3(n19042), .ZN(n18135) );
  INV_X1 U4999 ( .I(n1807), .ZN(n5656) );
  INV_X2 U7475 ( .I(n2935), .ZN(n1766) );
  INV_X2 U8673 ( .I(n19301), .ZN(n19291) );
  INV_X2 U26347 ( .I(n19180), .ZN(n784) );
  NOR2_X1 U21453 ( .A1(n18997), .A2(n18996), .ZN(n12937) );
  CLKBUF_X2 U1502 ( .I(n8024), .Z(n27818) );
  INV_X2 U12308 ( .I(n5491), .ZN(n17370) );
  NAND2_X1 U3709 ( .A1(n29047), .A2(n26417), .ZN(n5877) );
  NOR2_X1 U8708 ( .A1(n11940), .A2(n8379), .ZN(n1764) );
  INV_X1 U24129 ( .I(n19212), .ZN(n1373) );
  INV_X1 U5940 ( .I(n2799), .ZN(n3207) );
  INV_X1 U21428 ( .I(n19178), .ZN(n18957) );
  INV_X1 U6202 ( .I(n19156), .ZN(n27587) );
  INV_X1 U8712 ( .I(n15411), .ZN(n8742) );
  NAND2_X1 U8017 ( .A1(n31726), .A2(n19265), .ZN(n28447) );
  INV_X1 U4619 ( .I(n7197), .ZN(n19152) );
  INV_X1 U8627 ( .I(n8024), .ZN(n19242) );
  INV_X2 U1521 ( .I(n11203), .ZN(n827) );
  OR2_X1 U8252 ( .A1(n30879), .A2(n31746), .Z(n19148) );
  NAND2_X1 U8747 ( .A1(n19267), .A2(n19268), .ZN(n19270) );
  AOI21_X1 U16817 ( .A1(n19113), .A2(n19112), .B(n27587), .ZN(n27353) );
  CLKBUF_X2 U1804 ( .I(n19220), .Z(n4) );
  NAND2_X1 U3553 ( .A1(n1052), .A2(n26600), .ZN(n4658) );
  OAI21_X1 U26139 ( .A1(n19112), .A2(n12549), .B(n19113), .ZN(n26250) );
  NAND2_X1 U21716 ( .A1(n19179), .A2(n18957), .ZN(n11955) );
  AOI21_X1 U1469 ( .A1(n19103), .A2(n19100), .B(n17445), .ZN(n27076) );
  NOR2_X1 U4019 ( .A1(n4066), .A2(n19158), .ZN(n18970) );
  NAND2_X1 U1922 ( .A1(n4835), .A2(n30817), .ZN(n18967) );
  NAND2_X1 U10718 ( .A1(n19032), .A2(n10203), .ZN(n18788) );
  NAND3_X1 U5183 ( .A1(n19060), .A2(n9787), .A3(n1179), .ZN(n2410) );
  NOR2_X1 U12451 ( .A1(n19101), .A2(n11744), .ZN(n18952) );
  INV_X1 U12009 ( .I(n19085), .ZN(n18926) );
  NOR2_X1 U7454 ( .A1(n6343), .A2(n6342), .ZN(n9238) );
  NAND3_X1 U7463 ( .A1(n12468), .A2(n12505), .A3(n1378), .ZN(n12504) );
  INV_X1 U7497 ( .I(n9885), .ZN(n12815) );
  INV_X1 U8338 ( .I(n13219), .ZN(n26355) );
  AOI21_X1 U9980 ( .A1(n19217), .A2(n29), .B(n827), .ZN(n6578) );
  INV_X1 U5005 ( .I(n18958), .ZN(n4749) );
  NAND3_X1 U8641 ( .A1(n14148), .A2(n19088), .A3(n12807), .ZN(n18991) );
  NOR2_X1 U5933 ( .A1(n14233), .A2(n11203), .ZN(n18999) );
  OAI22_X1 U15432 ( .A1(n19090), .A2(n1047), .B1(n19091), .B2(n5760), .ZN(
        n17556) );
  OAI21_X1 U8878 ( .A1(n16768), .A2(n16769), .B(n18440), .ZN(n17997) );
  NAND2_X1 U9984 ( .A1(n9078), .A2(n2970), .ZN(n8828) );
  NAND2_X1 U22767 ( .A1(n8233), .A2(n19124), .ZN(n18955) );
  INV_X1 U7472 ( .I(n31658), .ZN(n15910) );
  INV_X1 U8706 ( .I(n18974), .ZN(n1048) );
  NAND2_X1 U938 ( .A1(n7134), .A2(n743), .ZN(n19039) );
  NAND2_X1 U5199 ( .A1(n947), .A2(n14312), .ZN(n6446) );
  NAND2_X1 U6587 ( .A1(n950), .A2(n7732), .ZN(n15396) );
  NAND2_X1 U3340 ( .A1(n1378), .A2(n16185), .ZN(n379) );
  INV_X1 U5487 ( .I(n19262), .ZN(n19140) );
  NOR2_X1 U4945 ( .A1(n5118), .A2(n7995), .ZN(n18953) );
  INV_X1 U901 ( .I(n27743), .ZN(n17238) );
  NAND2_X1 U1944 ( .A1(n1630), .A2(n33608), .ZN(n2703) );
  NAND2_X1 U8644 ( .A1(n2177), .A2(n19143), .ZN(n1631) );
  NOR2_X1 U1507 ( .A1(n15534), .A2(n4747), .ZN(n26553) );
  OAI22_X1 U9994 ( .A1(n19133), .A2(n15050), .B1(n19132), .B2(n1050), .ZN(
        n15126) );
  AOI21_X1 U22684 ( .A1(n7557), .A2(n12502), .B(n27941), .ZN(n13449) );
  AOI22_X1 U5467 ( .A1(n6142), .A2(n1054), .B1(n1373), .B2(n29963), .ZN(n4191)
         );
  OAI21_X1 U11316 ( .A1(n19179), .A2(n19181), .B(n13200), .ZN(n18917) );
  NOR2_X1 U6272 ( .A1(n11000), .A2(n19315), .ZN(n18230) );
  OAI21_X1 U15640 ( .A1(n32451), .A2(n19036), .B(n12850), .ZN(n12849) );
  NOR2_X1 U5214 ( .A1(n19038), .A2(n31139), .ZN(n7749) );
  NAND2_X1 U890 ( .A1(n29378), .A2(n827), .ZN(n18938) );
  OAI22_X1 U3160 ( .A1(n19154), .A2(n950), .B1(n8862), .B2(n879), .ZN(n13072)
         );
  NAND2_X1 U10027 ( .A1(n16068), .A2(n7968), .ZN(n17319) );
  NAND2_X1 U2534 ( .A1(n19309), .A2(n14178), .ZN(n2519) );
  AOI22_X1 U26143 ( .A1(n4102), .A2(n26417), .B1(n30412), .B2(n19032), .ZN(
        n29044) );
  NAND2_X1 U5244 ( .A1(n15845), .A2(n19281), .ZN(n15843) );
  OAI21_X1 U21190 ( .A1(n15628), .A2(n32908), .B(n28386), .ZN(n15627) );
  OAI21_X1 U8632 ( .A1(n7201), .A2(n7200), .B(n33581), .ZN(n7199) );
  OAI21_X1 U18140 ( .A1(n19291), .A2(n29223), .B(n13957), .ZN(n18927) );
  NOR2_X1 U21730 ( .A1(n11875), .A2(n28175), .ZN(n14355) );
  NOR2_X1 U8633 ( .A1(n14030), .A2(n5812), .ZN(n4386) );
  NAND2_X1 U7505 ( .A1(n19315), .A2(n31970), .ZN(n19151) );
  INV_X1 U8648 ( .I(n1494), .ZN(n1492) );
  NAND2_X1 U12420 ( .A1(n18477), .A2(n14760), .ZN(n18381) );
  NAND2_X1 U1512 ( .A1(n1883), .A2(n16699), .ZN(n12813) );
  NOR2_X1 U24469 ( .A1(n827), .A2(n7557), .ZN(n19349) );
  OAI21_X1 U12144 ( .A1(n19260), .A2(n744), .B(n16740), .ZN(n16741) );
  NAND2_X1 U8422 ( .A1(n19177), .A2(n19178), .ZN(n29580) );
  OAI21_X1 U21486 ( .A1(n1883), .A2(n12815), .B(n12813), .ZN(n18813) );
  OAI21_X1 U21017 ( .A1(n17527), .A2(n31029), .B(n26518), .ZN(n11295) );
  NAND2_X1 U1921 ( .A1(n10013), .A2(n2582), .ZN(n19056) );
  NAND3_X1 U1456 ( .A1(n9441), .A2(n9442), .A3(n1180), .ZN(n16797) );
  INV_X1 U5160 ( .I(n19676), .ZN(n1369) );
  BUF_X2 U10240 ( .I(Key[60]), .Z(n25598) );
  AOI22_X1 U15524 ( .A1(n19139), .A2(n28379), .B1(n19140), .B2(n16876), .ZN(
        n16875) );
  AOI21_X1 U6288 ( .A1(n18982), .A2(n13685), .B(n17508), .ZN(n17507) );
  NAND2_X1 U4983 ( .A1(n26289), .A2(n26288), .ZN(n8897) );
  NOR2_X1 U9970 ( .A1(n17528), .A2(n17526), .ZN(n13355) );
  CLKBUF_X2 U1451 ( .I(n19710), .Z(n25998) );
  NAND2_X1 U13057 ( .A1(n2126), .A2(n2125), .ZN(n16158) );
  INV_X1 U3091 ( .I(n19768), .ZN(n1363) );
  INV_X1 U24436 ( .I(n19136), .ZN(n19142) );
  INV_X1 U9765 ( .I(n9629), .ZN(n1368) );
  INV_X1 U18921 ( .I(n13480), .ZN(n7826) );
  INV_X1 U1885 ( .I(n31882), .ZN(n31057) );
  NOR3_X1 U4949 ( .A1(n1984), .A2(n5606), .A3(n5608), .ZN(n5605) );
  INV_X1 U20879 ( .I(n30411), .ZN(n19498) );
  INV_X1 U18294 ( .I(n14094), .ZN(n19566) );
  BUF_X2 U12519 ( .I(n14120), .Z(n26794) );
  CLKBUF_X2 U1891 ( .I(n6387), .Z(n30212) );
  INV_X1 U6569 ( .I(n14214), .ZN(n19375) );
  INV_X1 U2821 ( .I(n13645), .ZN(n19479) );
  INV_X1 U5273 ( .I(n19780), .ZN(n30712) );
  INV_X1 U6322 ( .I(n19568), .ZN(n2375) );
  INV_X1 U6269 ( .I(n12610), .ZN(n29046) );
  BUF_X2 U22847 ( .I(n29130), .Z(n31279) );
  INV_X1 U877 ( .I(n19378), .ZN(n1173) );
  BUF_X2 U15123 ( .I(Key[20]), .Z(n16581) );
  OAI22_X1 U3254 ( .A1(n7438), .A2(n12532), .B1(n7437), .B2(n7436), .ZN(n27144) );
  INV_X1 U1442 ( .I(n25266), .ZN(n26000) );
  CLKBUF_X2 U2103 ( .I(n16158), .Z(n29890) );
  INV_X1 U24031 ( .I(n31414), .ZN(n31908) );
  INV_X1 U16319 ( .I(n4883), .ZN(n14766) );
  INV_X1 U1881 ( .I(n24487), .ZN(n30993) );
  INV_X1 U10319 ( .I(n26551), .ZN(n219) );
  INV_X1 U11937 ( .I(n15189), .ZN(n2780) );
  INV_X1 U6314 ( .I(n11333), .ZN(n1040) );
  INV_X2 U8527 ( .I(n8443), .ZN(n6864) );
  INV_X1 U13579 ( .I(n568), .ZN(n1043) );
  INV_X1 U25215 ( .I(n31538), .ZN(n31906) );
  NAND2_X1 U7417 ( .A1(n1043), .A2(n16694), .ZN(n7923) );
  INV_X1 U9946 ( .I(n14576), .ZN(n20119) );
  NOR2_X1 U21561 ( .A1(n20099), .A2(n29216), .ZN(n13978) );
  INV_X1 U14087 ( .I(n9469), .ZN(n12045) );
  INV_X2 U11876 ( .I(n20113), .ZN(n20044) );
  NAND2_X1 U8517 ( .A1(n6611), .A2(n19991), .ZN(n17136) );
  INV_X2 U849 ( .I(n18089), .ZN(n8107) );
  BUF_X2 U2753 ( .I(n19857), .Z(n28645) );
  NAND2_X1 U12114 ( .A1(n8816), .A2(n29250), .ZN(n19933) );
  INV_X2 U2760 ( .I(n19857), .ZN(n20068) );
  INV_X1 U13413 ( .I(n2499), .ZN(n20076) );
  INV_X2 U862 ( .I(n11913), .ZN(n19986) );
  INV_X2 U14698 ( .I(n17575), .ZN(n20056) );
  INV_X1 U20330 ( .I(n10863), .ZN(n13327) );
  INV_X1 U19734 ( .I(n578), .ZN(n1165) );
  INV_X1 U7403 ( .I(n31453), .ZN(n20043) );
  INV_X1 U1438 ( .I(n1043), .ZN(n28684) );
  INV_X2 U19246 ( .I(n8684), .ZN(n17882) );
  BUF_X2 U2905 ( .I(n19885), .Z(n224) );
  INV_X2 U4606 ( .I(n14761), .ZN(n17260) );
  INV_X1 U820 ( .I(n19991), .ZN(n11624) );
  OAI22_X1 U1416 ( .A1(n11350), .A2(n28684), .B1(n7920), .B2(n1360), .ZN(
        n18003) );
  NAND2_X1 U5300 ( .A1(n19845), .A2(n16681), .ZN(n1878) );
  NAND2_X1 U11927 ( .A1(n29013), .A2(n502), .ZN(n15736) );
  OAI21_X1 U20999 ( .A1(n20136), .A2(n19834), .B(n15174), .ZN(n12634) );
  INV_X1 U10277 ( .I(n9201), .ZN(n26547) );
  NOR2_X1 U21536 ( .A1(n16092), .A2(n19966), .ZN(n15258) );
  NAND2_X1 U2685 ( .A1(n12682), .A2(n1169), .ZN(n28012) );
  NAND2_X1 U11036 ( .A1(n31468), .A2(n16154), .ZN(n29853) );
  NAND2_X1 U23549 ( .A1(n9876), .A2(n8301), .ZN(n20081) );
  NOR2_X1 U6408 ( .A1(n17260), .A2(n1699), .ZN(n15247) );
  INV_X1 U1832 ( .I(n20124), .ZN(n16155) );
  INV_X2 U19845 ( .I(n28704), .ZN(n10340) );
  INV_X2 U2866 ( .I(n20056), .ZN(n19883) );
  BUF_X2 U6375 ( .I(n8857), .Z(n431) );
  INV_X1 U836 ( .I(n20155), .ZN(n14747) );
  INV_X2 U9951 ( .I(n14457), .ZN(n5707) );
  INV_X1 U1776 ( .I(n32745), .ZN(n15551) );
  INV_X1 U8562 ( .I(n12045), .ZN(n19856) );
  NAND2_X1 U5286 ( .A1(n11521), .A2(n10947), .ZN(n28218) );
  INV_X1 U26411 ( .I(n29250), .ZN(n570) );
  OR2_X1 U3035 ( .A1(n10059), .A2(n9690), .Z(n19974) );
  INV_X2 U22765 ( .I(n20135), .ZN(n15286) );
  INV_X1 U4232 ( .I(n32807), .ZN(n19451) );
  INV_X1 U5456 ( .I(n11959), .ZN(n8611) );
  INV_X1 U1436 ( .I(n16595), .ZN(n20020) );
  INV_X2 U1828 ( .I(n27808), .ZN(n4142) );
  NAND2_X1 U11427 ( .A1(n16625), .A2(n29252), .ZN(n11593) );
  BUF_X2 U26138 ( .I(n19936), .Z(n29040) );
  INV_X2 U9916 ( .I(n15381), .ZN(n14976) );
  INV_X2 U7421 ( .I(n31448), .ZN(n20066) );
  NAND2_X1 U2520 ( .A1(n19724), .A2(n567), .ZN(n9031) );
  INV_X1 U14899 ( .I(n16298), .ZN(n31694) );
  AOI21_X1 U17922 ( .A1(n13327), .A2(n584), .B(n16489), .ZN(n14801) );
  NOR2_X1 U1847 ( .A1(n6532), .A2(n10845), .ZN(n19338) );
  OAI22_X1 U10882 ( .A1(n2089), .A2(n3486), .B1(n19974), .B2(n15189), .ZN(
        n27604) );
  NOR3_X1 U1797 ( .A1(n19808), .A2(n16491), .A3(n15278), .ZN(n11902) );
  OAI22_X1 U24641 ( .A1(n20085), .A2(n20084), .B1(n16664), .B2(n9876), .ZN(
        n20086) );
  AOI22_X1 U17717 ( .A1(n940), .A2(n4233), .B1(n4215), .B2(n20157), .ZN(n4230)
         );
  NOR2_X1 U10752 ( .A1(n20061), .A2(n27832), .ZN(n20062) );
  NOR2_X1 U20890 ( .A1(n20068), .A2(n20067), .ZN(n20069) );
  OAI22_X1 U12490 ( .A1(n19926), .A2(n13591), .B1(n19614), .B2(n27097), .ZN(
        n19623) );
  NAND3_X1 U17450 ( .A1(n9033), .A2(n19806), .A3(n30375), .ZN(n9032) );
  OAI21_X1 U1364 ( .A1(n16966), .A2(n28600), .B(n1699), .ZN(n20104) );
  NAND2_X1 U7368 ( .A1(n19951), .A2(n12045), .ZN(n2845) );
  NAND2_X1 U15514 ( .A1(n18003), .A2(n27624), .ZN(n4167) );
  AOI22_X1 U21123 ( .A1(n28852), .A2(n375), .B1(n15192), .B2(n19874), .ZN(
        n31048) );
  NOR2_X1 U1413 ( .A1(n27715), .A2(n28645), .ZN(n17712) );
  NAND2_X1 U19196 ( .A1(n33419), .A2(n20156), .ZN(n8591) );
  OAI21_X1 U20359 ( .A1(n17714), .A2(n17713), .B(n19451), .ZN(n10925) );
  NOR2_X1 U24643 ( .A1(n14083), .A2(n20120), .ZN(n20121) );
  NOR2_X1 U8563 ( .A1(n12657), .A2(n149), .ZN(n10768) );
  INV_X1 U3898 ( .I(n6027), .ZN(n30845) );
  AOI21_X1 U2122 ( .A1(n20056), .A2(n11958), .B(n15665), .ZN(n4637) );
  NOR2_X1 U1350 ( .A1(n19824), .A2(n15306), .ZN(n8431) );
  NAND2_X1 U1843 ( .A1(n14644), .A2(n20000), .ZN(n30790) );
  AND2_X1 U4518 ( .A1(n11198), .A2(n31951), .Z(n17156) );
  OAI21_X1 U21986 ( .A1(n11521), .A2(n28219), .B(n28218), .ZN(n19843) );
  NOR2_X1 U1390 ( .A1(n20099), .A2(n28087), .ZN(n9855) );
  NAND2_X1 U16569 ( .A1(n19969), .A2(n19970), .ZN(n2908) );
  NOR2_X1 U18847 ( .A1(n1164), .A2(n16694), .ZN(n8295) );
  INV_X1 U832 ( .I(n16154), .ZN(n19840) );
  OAI21_X1 U12300 ( .A1(n783), .A2(n20147), .B(n4602), .ZN(n4443) );
  NAND2_X1 U23500 ( .A1(n27597), .A2(n11961), .ZN(n17365) );
  NOR2_X1 U1395 ( .A1(n2694), .A2(n19995), .ZN(n26238) );
  INV_X1 U5156 ( .I(n3989), .ZN(n14927) );
  INV_X1 U10981 ( .I(n1358), .ZN(n29845) );
  NAND2_X1 U26176 ( .A1(n28208), .A2(n28209), .ZN(n5549) );
  AOI21_X1 U1787 ( .A1(n20081), .A2(n13585), .B(n32780), .ZN(n20087) );
  AOI22_X1 U8531 ( .A1(n9450), .A2(n33743), .B1(n16155), .B2(n20120), .ZN(
        n9449) );
  INV_X1 U14741 ( .I(n11872), .ZN(n27318) );
  NAND2_X1 U6527 ( .A1(n4233), .A2(n20043), .ZN(n13611) );
  NOR2_X1 U20260 ( .A1(n29208), .A2(n17389), .ZN(n10695) );
  NOR2_X1 U20064 ( .A1(n10272), .A2(n16694), .ZN(n10271) );
  NOR2_X1 U5889 ( .A1(n12337), .A2(n14210), .ZN(n20144) );
  INV_X1 U6554 ( .I(n17882), .ZN(n19943) );
  NOR2_X1 U2712 ( .A1(n31993), .A2(n8216), .ZN(n14134) );
  NOR2_X1 U15109 ( .A1(n1362), .A2(n18142), .ZN(n18141) );
  NAND2_X1 U21472 ( .A1(n14334), .A2(n16595), .ZN(n20125) );
  AND2_X1 U19704 ( .A1(n6275), .A2(n8933), .Z(n4855) );
  INV_X1 U21034 ( .I(n20076), .ZN(n16059) );
  NAND2_X1 U25903 ( .A1(n149), .A2(n29040), .ZN(n28880) );
  INV_X1 U7413 ( .I(n822), .ZN(n1438) );
  NOR2_X1 U5288 ( .A1(n4215), .A2(n940), .ZN(n10556) );
  INV_X1 U22551 ( .I(n33714), .ZN(n5598) );
  AOI21_X1 U6519 ( .A1(n20144), .A2(n20143), .B(n12851), .ZN(n2495) );
  NOR3_X1 U8265 ( .A1(n16059), .A2(n12379), .A3(n6444), .ZN(n12832) );
  OAI21_X1 U26088 ( .A1(n31697), .A2(n29284), .B(n31715), .ZN(n31676) );
  OAI21_X1 U24393 ( .A1(n20036), .A2(n8775), .B(n29187), .ZN(n28622) );
  OAI21_X1 U21275 ( .A1(n19932), .A2(n31103), .B(n579), .ZN(n14799) );
  AOI22_X1 U9887 ( .A1(n10465), .A2(n20077), .B1(n20079), .B2(n20078), .ZN(
        n12598) );
  OAI21_X1 U15158 ( .A1(n4972), .A2(n7014), .B(n19853), .ZN(n13283) );
  NAND3_X1 U17724 ( .A1(n6611), .A2(n28876), .A3(n30366), .ZN(n15850) );
  NAND2_X1 U6401 ( .A1(n19878), .A2(n20096), .ZN(n8183) );
  NAND3_X1 U6522 ( .A1(n13583), .A2(n6960), .A3(n12168), .ZN(n4498) );
  NAND2_X1 U1740 ( .A1(n20065), .A2(n2606), .ZN(n30922) );
  OAI22_X1 U11814 ( .A1(n12696), .A2(n821), .B1(n20059), .B2(n19886), .ZN(
        n2146) );
  NAND2_X1 U1351 ( .A1(n3366), .A2(n13585), .ZN(n13772) );
  NOR2_X1 U12313 ( .A1(n1458), .A2(n14210), .ZN(n2549) );
  OAI21_X1 U17681 ( .A1(n2933), .A2(n9875), .B(n1167), .ZN(n27517) );
  NAND2_X1 U1377 ( .A1(n10340), .A2(n17670), .ZN(n28912) );
  NAND2_X1 U22852 ( .A1(n31280), .A2(n15381), .ZN(n13397) );
  NAND2_X1 U1837 ( .A1(n19438), .A2(n1358), .ZN(n11) );
  NAND3_X1 U3893 ( .A1(n8783), .A2(n8782), .A3(n17967), .ZN(n20190) );
  OAI21_X1 U1335 ( .A1(n32000), .A2(n14622), .B(n29656), .ZN(n13955) );
  NAND2_X1 U6377 ( .A1(n20063), .A2(n20062), .ZN(n15310) );
  NAND3_X1 U6392 ( .A1(n27829), .A2(n27830), .A3(n20135), .ZN(n31585) );
  NAND2_X1 U2259 ( .A1(n18949), .A2(n7609), .ZN(n15436) );
  OAI21_X1 U5140 ( .A1(n2534), .A2(n8443), .B(n6200), .ZN(n16951) );
  NAND2_X1 U3360 ( .A1(n2845), .A2(n31080), .ZN(n13284) );
  NAND2_X1 U16560 ( .A1(n20026), .A2(n6109), .ZN(n30356) );
  NOR2_X1 U21215 ( .A1(n19867), .A2(n19868), .ZN(n12987) );
  OAI21_X1 U6420 ( .A1(n13157), .A2(n783), .B(n330), .ZN(n19832) );
  OAI22_X1 U1365 ( .A1(n3593), .A2(n20053), .B1(n11893), .B2(n15665), .ZN(
        n3592) );
  INV_X2 U1726 ( .I(n20560), .ZN(n20562) );
  INV_X2 U12098 ( .I(n20632), .ZN(n15162) );
  NAND2_X1 U24889 ( .A1(n3940), .A2(n3941), .ZN(n28696) );
  BUF_X2 U5429 ( .I(n14720), .Z(n11086) );
  INV_X2 U6486 ( .I(n31969), .ZN(n20360) );
  INV_X1 U18405 ( .I(n20404), .ZN(n2237) );
  INV_X1 U4204 ( .I(n20339), .ZN(n20590) );
  NAND2_X1 U20929 ( .A1(n20430), .A2(n20590), .ZN(n16133) );
  NAND2_X1 U2897 ( .A1(n20158), .A2(n30130), .ZN(n10614) );
  INV_X2 U9605 ( .I(n16606), .ZN(n20563) );
  INV_X1 U15862 ( .I(n29763), .ZN(n20524) );
  NOR2_X1 U3203 ( .A1(n11086), .A2(n12966), .ZN(n20263) );
  INV_X2 U12462 ( .I(n10847), .ZN(n10849) );
  NOR2_X1 U23084 ( .A1(n20371), .A2(n15027), .ZN(n20205) );
  NAND2_X1 U1280 ( .A1(n5471), .A2(n20374), .ZN(n1774) );
  INV_X2 U2166 ( .I(n2821), .ZN(n14731) );
  INV_X1 U20413 ( .I(n15169), .ZN(n20591) );
  INV_X2 U9827 ( .I(n20361), .ZN(n1789) );
  NAND2_X1 U1284 ( .A1(n1150), .A2(n20562), .ZN(n27316) );
  INV_X1 U7308 ( .I(n2843), .ZN(n16070) );
  NAND2_X1 U21108 ( .A1(n19864), .A2(n20360), .ZN(n13247) );
  CLKBUF_X2 U7348 ( .I(n20582), .Z(n26232) );
  INV_X2 U5103 ( .I(n6679), .ZN(n1032) );
  INV_X2 U4927 ( .I(n28261), .ZN(n818) );
  INV_X1 U7335 ( .I(n9025), .ZN(n935) );
  NAND2_X1 U21603 ( .A1(n20602), .A2(n6996), .ZN(n12184) );
  INV_X1 U7736 ( .I(n8870), .ZN(n11312) );
  INV_X1 U19661 ( .I(n14187), .ZN(n9484) );
  INV_X1 U1256 ( .I(n20329), .ZN(n1149) );
  INV_X2 U17294 ( .I(n20615), .ZN(n27741) );
  INV_X1 U11626 ( .I(n26881), .ZN(n13537) );
  INV_X1 U1265 ( .I(n9831), .ZN(n13538) );
  INV_X1 U15861 ( .I(n4460), .ZN(n20358) );
  INV_X1 U12773 ( .I(n20467), .ZN(n20160) );
  INV_X2 U3119 ( .I(n4254), .ZN(n20487) );
  INV_X1 U1294 ( .I(n7218), .ZN(n1034) );
  INV_X1 U10575 ( .I(n28390), .ZN(n6475) );
  INV_X2 U2899 ( .I(n30130), .ZN(n710) );
  AOI22_X1 U3587 ( .A1(n29453), .A2(n31504), .B1(n20524), .B2(n33222), .ZN(
        n8794) );
  INV_X2 U17626 ( .I(n32504), .ZN(n30987) );
  INV_X1 U4206 ( .I(n935), .ZN(n1030) );
  NAND2_X1 U17975 ( .A1(n20450), .A2(n14179), .ZN(n12227) );
  BUF_X4 U774 ( .I(n10847), .Z(n10848) );
  NOR2_X1 U2314 ( .A1(n20202), .A2(n20361), .ZN(n120) );
  NOR2_X1 U11738 ( .A1(n12169), .A2(n2879), .ZN(n20235) );
  INV_X1 U1705 ( .I(n14436), .ZN(n1151) );
  INV_X1 U783 ( .I(n33515), .ZN(n1152) );
  INV_X1 U9781 ( .I(n20327), .ZN(n11809) );
  INV_X1 U7285 ( .I(n3944), .ZN(n17866) );
  NAND2_X1 U11868 ( .A1(n1357), .A2(n20635), .ZN(n20442) );
  NAND2_X1 U21098 ( .A1(n16182), .A2(n15230), .ZN(n3644) );
  BUF_X2 U4886 ( .I(n20374), .Z(n27887) );
  INV_X1 U7317 ( .I(n17236), .ZN(n4807) );
  NOR2_X1 U24692 ( .A1(n20381), .A2(n30594), .ZN(n20382) );
  INV_X1 U6457 ( .I(n16452), .ZN(n20510) );
  NAND2_X1 U1241 ( .A1(n20428), .A2(n20427), .ZN(n4856) );
  NAND2_X1 U13218 ( .A1(n8870), .A2(n31668), .ZN(n26424) );
  BUF_X2 U7297 ( .I(n16606), .Z(n13589) );
  NOR2_X1 U22958 ( .A1(n1150), .A2(n20413), .ZN(n14710) );
  INV_X1 U4862 ( .I(n15230), .ZN(n20603) );
  NOR2_X1 U4263 ( .A1(n1349), .A2(n20447), .ZN(n30003) );
  NOR2_X1 U6498 ( .A1(n28812), .A2(n14049), .ZN(n20221) );
  INV_X1 U3773 ( .I(n12563), .ZN(n9854) );
  INV_X1 U1293 ( .I(n30763), .ZN(n28316) );
  INV_X1 U3410 ( .I(n27697), .ZN(n20497) );
  INV_X2 U8404 ( .I(n20489), .ZN(n20484) );
  INV_X2 U16246 ( .I(n31968), .ZN(n11637) );
  INV_X1 U2359 ( .I(n11303), .ZN(n12010) );
  INV_X1 U743 ( .I(n20401), .ZN(n20571) );
  NOR2_X1 U5440 ( .A1(n7577), .A2(n20395), .ZN(n20462) );
  INV_X1 U1698 ( .I(n20471), .ZN(n931) );
  NAND2_X1 U13916 ( .A1(n20317), .A2(n32504), .ZN(n2965) );
  INV_X1 U5442 ( .I(n20447), .ZN(n781) );
  NAND2_X1 U7391 ( .A1(n3944), .A2(n15282), .ZN(n1465) );
  NAND2_X1 U2555 ( .A1(n17866), .A2(n1355), .ZN(n15713) );
  NAND2_X1 U26568 ( .A1(n32033), .A2(n8031), .ZN(n31834) );
  NAND2_X1 U21395 ( .A1(n14369), .A2(n20507), .ZN(n17652) );
  INV_X1 U2126 ( .I(n30931), .ZN(n30413) );
  NOR2_X1 U17304 ( .A1(n5275), .A2(n10106), .ZN(n27442) );
  NOR2_X1 U7275 ( .A1(n1150), .A2(n20562), .ZN(n5952) );
  NAND2_X1 U14016 ( .A1(n20194), .A2(n27755), .ZN(n3065) );
  NAND3_X1 U23052 ( .A1(n28357), .A2(n31009), .A3(n20489), .ZN(n14945) );
  NAND2_X1 U735 ( .A1(n20412), .A2(n818), .ZN(n3137) );
  NOR2_X1 U13789 ( .A1(n14054), .A2(n2843), .ZN(n17043) );
  OAI22_X1 U7246 ( .A1(n19830), .A2(n20427), .B1(n28376), .B2(n14731), .ZN(
        n9725) );
  AOI21_X1 U1633 ( .A1(n20536), .A2(n20537), .B(n20541), .ZN(n11447) );
  NAND2_X1 U16846 ( .A1(n15045), .A2(n20563), .ZN(n16217) );
  NAND2_X1 U1564 ( .A1(n13353), .A2(n28288), .ZN(n5416) );
  NOR2_X1 U22977 ( .A1(n28527), .A2(n7873), .ZN(n14768) );
  NAND2_X1 U20838 ( .A1(n19930), .A2(n13589), .ZN(n16216) );
  NAND2_X1 U6296 ( .A1(n27697), .A2(n31804), .ZN(n26089) );
  NAND2_X1 U21531 ( .A1(n8998), .A2(n20630), .ZN(n14566) );
  AOI21_X1 U19868 ( .A1(n20538), .A2(n760), .B(n4071), .ZN(n11446) );
  NAND2_X1 U4843 ( .A1(n20382), .A2(n111), .ZN(n26987) );
  INV_X1 U11728 ( .I(n13253), .ZN(n8942) );
  OAI21_X1 U18289 ( .A1(n30603), .A2(n16123), .B(n16452), .ZN(n28752) );
  INV_X1 U5382 ( .I(n16144), .ZN(n930) );
  NOR2_X1 U11718 ( .A1(n13253), .A2(n28085), .ZN(n9776) );
  NAND2_X1 U13369 ( .A1(n20235), .A2(n33530), .ZN(n16488) );
  BUF_X2 U10454 ( .I(n29814), .Z(n29774) );
  INV_X1 U15324 ( .I(n5781), .ZN(n20493) );
  NAND2_X1 U11653 ( .A1(n16882), .A2(n9014), .ZN(n9288) );
  NAND2_X1 U11687 ( .A1(n8650), .A2(n2879), .ZN(n15954) );
  NOR2_X1 U7904 ( .A1(n29363), .A2(n29528), .ZN(n29527) );
  INV_X1 U19041 ( .I(n20224), .ZN(n11712) );
  NAND2_X1 U1549 ( .A1(n10848), .A2(n1349), .ZN(n10074) );
  NAND2_X1 U17889 ( .A1(n30553), .A2(n32061), .ZN(n31444) );
  NOR2_X1 U1841 ( .A1(n1151), .A2(n26587), .ZN(n7707) );
  NAND2_X1 U4856 ( .A1(n1149), .A2(n13693), .ZN(n13325) );
  NOR2_X1 U15901 ( .A1(n31072), .A2(n31961), .ZN(n20002) );
  INV_X1 U7556 ( .I(n13867), .ZN(n26257) );
  INV_X1 U15237 ( .I(n11453), .ZN(n27386) );
  AOI21_X1 U21606 ( .A1(n14368), .A2(n3944), .B(n14369), .ZN(n14367) );
  NAND3_X1 U9385 ( .A1(n10231), .A2(n20520), .A3(n16218), .ZN(n29672) );
  OAI21_X1 U24627 ( .A1(n28626), .A2(n26567), .B(n20001), .ZN(n20004) );
  AOI21_X1 U20924 ( .A1(n20325), .A2(n932), .B(n16174), .ZN(n16492) );
  OAI21_X1 U9776 ( .A1(n20405), .A2(n10848), .B(n11616), .ZN(n11618) );
  AOI22_X1 U12998 ( .A1(n3428), .A2(n29623), .B1(n1157), .B2(n17043), .ZN(
        n30079) );
  OAI22_X1 U21394 ( .A1(n17652), .A2(n20510), .B1(n20508), .B2(n20509), .ZN(
        n16774) );
  NAND3_X1 U1231 ( .A1(n28357), .A2(n20487), .A3(n20486), .ZN(n17513) );
  OAI21_X1 U8379 ( .A1(n12771), .A2(n12169), .B(n15954), .ZN(n8960) );
  NAND3_X1 U21604 ( .A1(n7116), .A2(n1160), .A3(n16182), .ZN(n14965) );
  AOI22_X1 U11380 ( .A1(n5950), .A2(n20562), .B1(n933), .B2(n16684), .ZN(n5949) );
  NAND2_X1 U9753 ( .A1(n13353), .A2(n30878), .ZN(n7054) );
  NAND3_X1 U23085 ( .A1(n20533), .A2(n1153), .A3(n15027), .ZN(n20353) );
  NOR2_X1 U9750 ( .A1(n20252), .A2(n20484), .ZN(n7479) );
  NAND3_X1 U17404 ( .A1(n14566), .A2(n20631), .A3(n111), .ZN(n14565) );
  AOI21_X1 U7622 ( .A1(n15045), .A2(n13589), .B(n9776), .ZN(n9775) );
  NAND3_X1 U1527 ( .A1(n30545), .A2(n30987), .A3(n7394), .ZN(n2770) );
  NOR2_X1 U20928 ( .A1(n20378), .A2(n5471), .ZN(n16139) );
  NAND3_X1 U20836 ( .A1(n20341), .A2(n20340), .A3(n26756), .ZN(n12846) );
  INV_X1 U1556 ( .I(n7397), .ZN(n20220) );
  NAND2_X1 U1205 ( .A1(n16787), .A2(n14177), .ZN(n14176) );
  OR2_X1 U9759 ( .A1(n20341), .A2(n1347), .Z(n14263) );
  OAI21_X1 U11645 ( .A1(n14571), .A2(n14005), .B(n15173), .ZN(n6311) );
  AOI21_X1 U23490 ( .A1(n31338), .A2(n3904), .B(n20238), .ZN(n9587) );
  AOI21_X1 U6481 ( .A1(n20358), .A2(n28625), .B(n31891), .ZN(n2320) );
  OAI21_X1 U7268 ( .A1(n3751), .A2(n3750), .B(n15217), .ZN(n20612) );
  NAND2_X1 U9796 ( .A1(n14051), .A2(n14050), .ZN(n31269) );
  NAND2_X1 U1544 ( .A1(n31422), .A2(n31210), .ZN(n30856) );
  NAND3_X1 U1565 ( .A1(n266), .A2(n20268), .A3(n20492), .ZN(n19954) );
  AOI21_X1 U6473 ( .A1(n20440), .A2(n2565), .B(n34155), .ZN(n20441) );
  NAND2_X1 U11747 ( .A1(n1159), .A2(n32201), .ZN(n2619) );
  INV_X1 U20528 ( .I(n30929), .ZN(n10489) );
  INV_X1 U17456 ( .I(n1344), .ZN(n20832) );
  INV_X1 U7239 ( .I(n20698), .ZN(n20783) );
  NAND2_X1 U734 ( .A1(n20899), .A2(n20954), .ZN(n4269) );
  NAND3_X1 U11677 ( .A1(n817), .A2(n20499), .A3(n33116), .ZN(n20500) );
  OAI21_X1 U8408 ( .A1(n20451), .A2(n16139), .B(n20452), .ZN(n2318) );
  AOI21_X1 U6497 ( .A1(n6530), .A2(n16174), .B(n29938), .ZN(n2250) );
  INV_X1 U1562 ( .I(n20963), .ZN(n30013) );
  INV_X1 U3813 ( .I(n20729), .ZN(n6548) );
  NOR2_X1 U12816 ( .A1(n30552), .A2(n1909), .ZN(n1908) );
  INV_X1 U6469 ( .I(n20849), .ZN(n13602) );
  INV_X1 U22770 ( .I(n29898), .ZN(n26255) );
  INV_X1 U7237 ( .I(n21043), .ZN(n20586) );
  INV_X1 U1187 ( .I(n2198), .ZN(n17659) );
  INV_X1 U3398 ( .I(n21016), .ZN(n26575) );
  INV_X1 U8368 ( .I(n17423), .ZN(n1341) );
  BUF_X2 U13935 ( .I(n1787), .Z(n30171) );
  BUF_X2 U1194 ( .I(n16173), .Z(n348) );
  BUF_X2 U1195 ( .I(n5572), .Z(n28864) );
  INV_X1 U8376 ( .I(n20954), .ZN(n4758) );
  INV_X1 U717 ( .I(n20961), .ZN(n20183) );
  INV_X1 U4200 ( .I(n20726), .ZN(n1338) );
  INV_X1 U723 ( .I(n20862), .ZN(n1342) );
  INV_X1 U11613 ( .I(n20905), .ZN(n5009) );
  CLKBUF_X2 U5895 ( .I(n20679), .Z(n28822) );
  INV_X1 U20594 ( .I(n519), .ZN(n924) );
  NAND2_X1 U5477 ( .A1(n16652), .A2(n14556), .ZN(n7756) );
  NAND2_X1 U2223 ( .A1(n17313), .A2(n28714), .ZN(n2230) );
  INV_X2 U8343 ( .I(n28642), .ZN(n16785) );
  INV_X2 U6459 ( .I(n1337), .ZN(n5883) );
  NAND2_X1 U14875 ( .A1(n29460), .A2(n26407), .ZN(n13130) );
  INV_X2 U13964 ( .I(n3193), .ZN(n11967) );
  INV_X1 U22158 ( .I(n28260), .ZN(n398) );
  INV_X1 U6451 ( .I(n15226), .ZN(n21267) );
  INV_X1 U24094 ( .I(n28594), .ZN(n21338) );
  INV_X2 U8203 ( .I(n17313), .ZN(n3673) );
  INV_X2 U7203 ( .I(n515), .ZN(n2822) );
  INV_X2 U7205 ( .I(n26712), .ZN(n21434) );
  INV_X1 U19491 ( .I(n26345), .ZN(n30783) );
  NAND2_X1 U20843 ( .A1(n33498), .A2(n29062), .ZN(n13101) );
  OR2_X1 U4947 ( .A1(n5392), .A2(n8074), .Z(n21402) );
  OAI21_X1 U17672 ( .A1(n11187), .A2(n21189), .B(n2822), .ZN(n27515) );
  NAND2_X1 U1663 ( .A1(n27939), .A2(n21328), .ZN(n26326) );
  INV_X1 U1133 ( .I(n21152), .ZN(n27689) );
  AOI21_X1 U5551 ( .A1(n4381), .A2(n21322), .B(n1145), .ZN(n7122) );
  CLKBUF_X2 U19988 ( .I(n6855), .Z(n30854) );
  INV_X2 U2831 ( .I(n14556), .ZN(n921) );
  INV_X2 U8602 ( .I(n21165), .ZN(n6075) );
  NAND2_X1 U3005 ( .A1(n21160), .A2(n17305), .ZN(n15428) );
  INV_X1 U13744 ( .I(n11272), .ZN(n7822) );
  INV_X1 U6462 ( .I(n21412), .ZN(n929) );
  INV_X1 U6536 ( .I(n34089), .ZN(n27382) );
  INV_X2 U12822 ( .I(n28668), .ZN(n18218) );
  INV_X2 U6465 ( .I(n27028), .ZN(n17699) );
  INV_X1 U5116 ( .I(n21221), .ZN(n6451) );
  INV_X2 U657 ( .I(n21403), .ZN(n1335) );
  INV_X1 U14559 ( .I(n26971), .ZN(n27842) );
  AND2_X1 U23300 ( .A1(n8681), .A2(n17829), .Z(n21138) );
  INV_X1 U4195 ( .I(n21233), .ZN(n9699) );
  INV_X1 U658 ( .I(n12037), .ZN(n1334) );
  INV_X1 U5842 ( .I(n16072), .ZN(n21115) );
  NAND2_X1 U15511 ( .A1(n14290), .A2(n21403), .ZN(n21404) );
  NOR2_X1 U3006 ( .A1(n34157), .A2(n31874), .ZN(n21212) );
  INV_X1 U690 ( .I(n601), .ZN(n925) );
  INV_X1 U18123 ( .I(n17271), .ZN(n21353) );
  NAND2_X1 U10925 ( .A1(n1018), .A2(n3193), .ZN(n21169) );
  NOR2_X1 U23460 ( .A1(n8490), .A2(n26407), .ZN(n15968) );
  AOI21_X1 U18565 ( .A1(n26014), .A2(n9699), .B(n21138), .ZN(n2464) );
  NAND2_X1 U8236 ( .A1(n8604), .A2(n5049), .ZN(n5048) );
  INV_X8 U6458 ( .I(n10533), .ZN(n926) );
  INV_X1 U8353 ( .I(n17985), .ZN(n21175) );
  NAND2_X1 U24823 ( .A1(n921), .A2(n16652), .ZN(n21052) );
  OAI21_X1 U13105 ( .A1(n27075), .A2(n21085), .B(n21173), .ZN(n2176) );
  NAND2_X1 U10182 ( .A1(n6075), .A2(n29750), .ZN(n31170) );
  NAND2_X1 U8298 ( .A1(n31909), .A2(n16072), .ZN(n15220) );
  INV_X1 U11569 ( .I(n6451), .ZN(n2574) );
  NOR2_X1 U24882 ( .A1(n6408), .A2(n34157), .ZN(n21383) );
  AND2_X1 U9773 ( .A1(n15559), .A2(n28594), .Z(n26829) );
  NAND2_X1 U2239 ( .A1(n7430), .A2(n164), .ZN(n21332) );
  INV_X1 U22578 ( .I(n29255), .ZN(n21325) );
  NOR2_X1 U22717 ( .A1(n21407), .A2(n4324), .ZN(n14098) );
  NAND2_X1 U17479 ( .A1(n30784), .A2(n27482), .ZN(n3696) );
  NOR2_X1 U628 ( .A1(n21163), .A2(n1148), .ZN(n20881) );
  INV_X1 U13168 ( .I(n10787), .ZN(n13194) );
  NOR2_X1 U21129 ( .A1(n11966), .A2(n21369), .ZN(n16313) );
  CLKBUF_X2 U4791 ( .I(n13255), .Z(n28886) );
  CLKBUF_X2 U5865 ( .I(n10533), .Z(n31826) );
  INV_X2 U6514 ( .I(n1146), .ZN(n8011) );
  NAND2_X1 U11523 ( .A1(n7122), .A2(n7121), .ZN(n7120) );
  NAND2_X1 U20944 ( .A1(n31003), .A2(n27912), .ZN(n1982) );
  INV_X2 U3146 ( .I(n17624), .ZN(n21192) );
  INV_X1 U2568 ( .I(n29460), .ZN(n20676) );
  INV_X1 U673 ( .I(n29256), .ZN(n779) );
  INV_X1 U11560 ( .I(n18035), .ZN(n3717) );
  INV_X2 U636 ( .I(n1145), .ZN(n21321) );
  INV_X1 U6518 ( .I(n17341), .ZN(n1019) );
  INV_X1 U6445 ( .I(n21241), .ZN(n8453) );
  NAND2_X1 U1423 ( .A1(n3673), .A2(n7007), .ZN(n3672) );
  NAND2_X1 U16731 ( .A1(n67), .A2(n1632), .ZN(n30379) );
  OR2_X1 U6134 ( .A1(n9663), .A2(n8243), .Z(n26021) );
  NOR2_X1 U620 ( .A1(n32347), .A2(n11912), .ZN(n21335) );
  INV_X1 U19504 ( .I(n9322), .ZN(n17455) );
  INV_X1 U3959 ( .I(n17305), .ZN(n12525) );
  INV_X1 U8341 ( .I(n21239), .ZN(n21448) );
  INV_X1 U8348 ( .I(n21306), .ZN(n29574) );
  NOR2_X1 U1433 ( .A1(n6075), .A2(n21085), .ZN(n31702) );
  NOR2_X1 U18947 ( .A1(n31498), .A2(n13730), .ZN(n30694) );
  OAI21_X1 U20953 ( .A1(n21353), .A2(n30784), .B(n27075), .ZN(n21082) );
  NAND2_X1 U8559 ( .A1(n21192), .A2(n21427), .ZN(n30889) );
  NAND3_X1 U15876 ( .A1(n13712), .A2(n21251), .A3(n20662), .ZN(n28340) );
  NOR2_X1 U2578 ( .A1(n9664), .A2(n926), .ZN(n10527) );
  AOI21_X1 U8303 ( .A1(n7690), .A2(n33745), .B(n28641), .ZN(n14722) );
  OAI21_X1 U1100 ( .A1(n4119), .A2(n30755), .B(n21408), .ZN(n14998) );
  NOR3_X1 U17655 ( .A1(n9518), .A2(n17699), .A3(n29062), .ZN(n1967) );
  AOI21_X1 U22732 ( .A1(n6584), .A2(n21408), .B(n510), .ZN(n31262) );
  NOR2_X1 U22240 ( .A1(n26861), .A2(n11948), .ZN(n21171) );
  OAI21_X1 U5567 ( .A1(n11457), .A2(n21335), .B(n21243), .ZN(n11456) );
  INV_X1 U1362 ( .I(n21354), .ZN(n2172) );
  NAND2_X1 U10435 ( .A1(n31170), .A2(n21173), .ZN(n27424) );
  NAND2_X1 U22023 ( .A1(n8197), .A2(n1337), .ZN(n9258) );
  NAND2_X1 U10968 ( .A1(n29122), .A2(n6908), .ZN(n6907) );
  NOR2_X1 U8334 ( .A1(n21099), .A2(n21252), .ZN(n7773) );
  OAI21_X1 U1234 ( .A1(n4569), .A2(n2676), .B(n33106), .ZN(n2834) );
  NAND3_X1 U14333 ( .A1(n15015), .A2(n599), .A3(n2822), .ZN(n7913) );
  NOR2_X1 U3588 ( .A1(n31909), .A2(n21406), .ZN(n21298) );
  NAND2_X1 U17293 ( .A1(n10148), .A2(n1020), .ZN(n27440) );
  NOR2_X1 U20402 ( .A1(n8011), .A2(n21434), .ZN(n30913) );
  INV_X1 U1132 ( .I(n6908), .ZN(n8957) );
  INV_X1 U10147 ( .I(n33641), .ZN(n27230) );
  NOR2_X1 U8282 ( .A1(n10730), .A2(n16459), .ZN(n21619) );
  NOR2_X1 U8240 ( .A1(n8378), .A2(n33882), .ZN(n13975) );
  INV_X1 U21409 ( .I(n29062), .ZN(n15444) );
  NOR2_X1 U15184 ( .A1(n7690), .A2(n21223), .ZN(n14273) );
  NOR2_X1 U13766 ( .A1(n21322), .A2(n2822), .ZN(n21323) );
  NAND2_X1 U6532 ( .A1(n21082), .A2(n26861), .ZN(n15961) );
  INV_X1 U7146 ( .I(n21619), .ZN(n11265) );
  NOR2_X1 U1285 ( .A1(n12746), .A2(n13921), .ZN(n28074) );
  OAI21_X1 U11471 ( .A1(n20795), .A2(n28287), .B(n33641), .ZN(n16046) );
  AOI22_X1 U2695 ( .A1(n21320), .A2(n28017), .B1(n21323), .B2(n11187), .ZN(
        n29799) );
  AOI21_X1 U616 ( .A1(n21054), .A2(n5111), .B(n14643), .ZN(n10980) );
  NAND2_X1 U1405 ( .A1(n5575), .A2(n21452), .ZN(n9392) );
  NAND2_X1 U9618 ( .A1(n21381), .A2(n21209), .ZN(n10733) );
  OAI21_X1 U8235 ( .A1(n13975), .A2(n21120), .B(n12363), .ZN(n12373) );
  NAND3_X1 U24931 ( .A1(n21411), .A2(n34037), .A3(n11315), .ZN(n28699) );
  NOR2_X1 U1327 ( .A1(n16180), .A2(n21443), .ZN(n31507) );
  AOI22_X1 U1381 ( .A1(n31673), .A2(n18218), .B1(n8539), .B2(n1911), .ZN(n1910) );
  NAND2_X1 U22915 ( .A1(n21169), .A2(n10092), .ZN(n28385) );
  AOI22_X1 U20869 ( .A1(n12324), .A2(n21398), .B1(n3933), .B2(n12325), .ZN(
        n21399) );
  OAI21_X1 U11459 ( .A1(n30727), .A2(n10113), .B(n8727), .ZN(n7543) );
  NAND2_X1 U4703 ( .A1(n26018), .A2(n20936), .ZN(n28299) );
  NOR2_X1 U9714 ( .A1(n8378), .A2(n7430), .ZN(n11480) );
  NOR2_X1 U9689 ( .A1(n7430), .A2(n12925), .ZN(n7446) );
  OAI21_X1 U9631 ( .A1(n14273), .A2(n21317), .B(n15261), .ZN(n14272) );
  NAND2_X1 U23659 ( .A1(n15622), .A2(n779), .ZN(n28526) );
  NOR2_X1 U14613 ( .A1(n17011), .A2(n10527), .ZN(n30246) );
  NAND3_X1 U26419 ( .A1(n11456), .A2(n21069), .A3(n17666), .ZN(n13442) );
  NAND2_X1 U3468 ( .A1(n21447), .A2(n31730), .ZN(n21824) );
  NAND2_X1 U14883 ( .A1(n21264), .A2(n11745), .ZN(n16851) );
  AOI21_X1 U1112 ( .A1(n1329), .A2(n21109), .B(n26167), .ZN(n26166) );
  INV_X1 U1300 ( .I(n21738), .ZN(n21864) );
  INV_X1 U5830 ( .I(n196), .ZN(n14397) );
  OAI21_X1 U17841 ( .A1(n29382), .A2(n30544), .B(n21443), .ZN(n31853) );
  OAI21_X1 U9650 ( .A1(n11979), .A2(n12521), .B(n32907), .ZN(n21089) );
  OAI21_X1 U9231 ( .A1(n28074), .A2(n25942), .B(n32347), .ZN(n6880) );
  NOR2_X1 U2590 ( .A1(n6879), .A2(n6881), .ZN(n6878) );
  AOI22_X1 U24887 ( .A1(n21420), .A2(n21419), .B1(n33649), .B2(n21418), .ZN(
        n21421) );
  NAND2_X1 U2304 ( .A1(n6212), .A2(n16553), .ZN(n21462) );
  NAND2_X1 U25924 ( .A1(n3973), .A2(n16046), .ZN(n8875) );
  INV_X2 U21957 ( .I(n15091), .ZN(n1312) );
  AOI21_X1 U20255 ( .A1(n21200), .A2(n10686), .B(n9721), .ZN(n16546) );
  INV_X1 U562 ( .I(n13652), .ZN(n21736) );
  INV_X1 U5402 ( .I(n8457), .ZN(n1016) );
  INV_X1 U1212 ( .I(n13884), .ZN(n16157) );
  INV_X1 U6383 ( .I(n17716), .ZN(n1321) );
  CLKBUF_X2 U5811 ( .I(n16222), .Z(n8079) );
  BUF_X2 U2582 ( .I(n9999), .Z(n2296) );
  INV_X2 U1255 ( .I(n31911), .ZN(n30440) );
  INV_X2 U5404 ( .I(n13114), .ZN(n1013) );
  INV_X2 U1215 ( .I(n10720), .ZN(n861) );
  INV_X1 U9305 ( .I(n27954), .ZN(n916) );
  INV_X1 U17120 ( .I(n27379), .ZN(n21672) );
  INV_X2 U4325 ( .I(n17888), .ZN(n11596) );
  AND2_X1 U15800 ( .A1(n18208), .A2(n18206), .Z(n27178) );
  INV_X1 U25923 ( .I(n8875), .ZN(n21858) );
  INV_X2 U1018 ( .I(n30769), .ZN(n11300) );
  INV_X1 U18795 ( .I(n30389), .ZN(n30677) );
  INV_X1 U1156 ( .I(n21816), .ZN(n912) );
  NOR2_X1 U3365 ( .A1(n16157), .A2(n21122), .ZN(n29784) );
  INV_X1 U1269 ( .I(n16023), .ZN(n10254) );
  NAND2_X1 U2573 ( .A1(n920), .A2(n21733), .ZN(n185) );
  NAND2_X1 U5558 ( .A1(n230), .A2(n21706), .ZN(n6351) );
  OAI21_X1 U10172 ( .A1(n11300), .A2(n17348), .B(n32252), .ZN(n4434) );
  NAND2_X1 U1159 ( .A1(n21518), .A2(n916), .ZN(n29690) );
  INV_X1 U1166 ( .I(n33766), .ZN(n11276) );
  INV_X2 U9550 ( .I(n21730), .ZN(n17773) );
  INV_X1 U13969 ( .I(n11756), .ZN(n12711) );
  NAND2_X1 U585 ( .A1(n1009), .A2(n21832), .ZN(n15813) );
  INV_X1 U1038 ( .I(n31102), .ZN(n26727) );
  AOI21_X1 U9503 ( .A1(n16864), .A2(n16863), .B(n31458), .ZN(n16445) );
  NAND2_X1 U8206 ( .A1(n31957), .A2(n2368), .ZN(n14848) );
  INV_X1 U11103 ( .I(n3379), .ZN(n10532) );
  NAND2_X1 U3802 ( .A1(n1321), .A2(n3420), .ZN(n31732) );
  INV_X1 U1197 ( .I(n21852), .ZN(n8706) );
  INV_X1 U15695 ( .I(n32904), .ZN(n862) );
  INV_X1 U11344 ( .I(n17274), .ZN(n21535) );
  NOR2_X1 U11872 ( .A1(n29947), .A2(n1008), .ZN(n5342) );
  NOR2_X1 U11831 ( .A1(n9590), .A2(n9591), .ZN(n9589) );
  CLKBUF_X2 U5589 ( .I(n13652), .Z(n28018) );
  NAND3_X1 U20806 ( .A1(n6231), .A2(n3250), .A3(n29180), .ZN(n31645) );
  INV_X1 U11405 ( .I(n32252), .ZN(n3140) );
  INV_X1 U8639 ( .I(n31859), .ZN(n31910) );
  OAI21_X1 U4629 ( .A1(n727), .A2(n7592), .B(n21496), .ZN(n2514) );
  INV_X1 U16512 ( .I(n14236), .ZN(n1138) );
  INV_X1 U4554 ( .I(n9999), .ZN(n11890) );
  AND2_X1 U18190 ( .A1(n12866), .A2(n17431), .Z(n21459) );
  AND2_X1 U1025 ( .A1(n15863), .A2(n28429), .Z(n534) );
  INV_X1 U4389 ( .I(n5170), .ZN(n21625) );
  INV_X1 U3675 ( .I(n31309), .ZN(n11499) );
  NAND2_X1 U24911 ( .A1(n30885), .A2(n27635), .ZN(n21529) );
  CLKBUF_X2 U4657 ( .I(n21767), .Z(n28395) );
  BUF_X8 U5399 ( .I(n4029), .Z(n3467) );
  OAI21_X1 U17971 ( .A1(n1009), .A2(n33981), .B(n11890), .ZN(n6969) );
  NOR2_X1 U1107 ( .A1(n432), .A2(n29302), .ZN(n12028) );
  NAND3_X1 U24859 ( .A1(n27560), .A2(n29854), .A3(n21730), .ZN(n21277) );
  NAND2_X1 U558 ( .A1(n10775), .A2(n21603), .ZN(n5851) );
  NOR3_X1 U4548 ( .A1(n11861), .A2(n31654), .A3(n21780), .ZN(n28141) );
  NOR2_X1 U1139 ( .A1(n5546), .A2(n6544), .ZN(n4311) );
  AND2_X1 U4774 ( .A1(n30832), .A2(n7811), .Z(n27466) );
  OAI22_X1 U4587 ( .A1(n28654), .A2(n1318), .B1(n21671), .B2(n918), .ZN(n14541) );
  NOR2_X1 U20737 ( .A1(n27596), .A2(n21632), .ZN(n30962) );
  NOR2_X1 U1013 ( .A1(n32519), .A2(n17887), .ZN(n8403) );
  NAND2_X1 U22943 ( .A1(n15838), .A2(n14681), .ZN(n15837) );
  NOR2_X1 U2580 ( .A1(n32865), .A2(n2296), .ZN(n2298) );
  NAND3_X1 U22469 ( .A1(n2217), .A2(n21628), .A3(n29322), .ZN(n21574) );
  NAND2_X1 U1127 ( .A1(n11861), .A2(n31317), .ZN(n4212) );
  AOI21_X1 U10778 ( .A1(n21535), .A2(n21566), .B(n21351), .ZN(n9884) );
  INV_X1 U1086 ( .I(n14595), .ZN(n30114) );
  NAND2_X1 U21522 ( .A1(n21581), .A2(n13133), .ZN(n16723) );
  NOR2_X1 U23870 ( .A1(n21571), .A2(n30678), .ZN(n21572) );
  OAI21_X1 U919 ( .A1(n17428), .A2(n21459), .B(n21730), .ZN(n13199) );
  NOR2_X1 U24909 ( .A1(n21781), .A2(n31220), .ZN(n21523) );
  NOR2_X1 U1747 ( .A1(n7326), .A2(n11797), .ZN(n7325) );
  INV_X1 U11335 ( .I(n11619), .ZN(n13248) );
  NOR2_X1 U532 ( .A1(n12275), .A2(n12274), .ZN(n12273) );
  NAND2_X1 U3901 ( .A1(n28824), .A2(n5309), .ZN(n14948) );
  NAND2_X1 U1124 ( .A1(n31711), .A2(n28018), .ZN(n28067) );
  BUF_X2 U1782 ( .I(n14691), .Z(n1) );
  NAND2_X1 U1931 ( .A1(n17406), .A2(n21830), .ZN(n21831) );
  NOR2_X1 U17012 ( .A1(n6544), .A2(n6489), .ZN(n4359) );
  NOR2_X1 U9575 ( .A1(n21777), .A2(n21743), .ZN(n21744) );
  AOI21_X1 U2585 ( .A1(n10699), .A2(n30441), .B(n30440), .ZN(n26671) );
  INV_X1 U1422 ( .I(n16147), .ZN(n21817) );
  INV_X1 U5124 ( .I(n26445), .ZN(n1014) );
  INV_X1 U6427 ( .I(n28450), .ZN(n864) );
  AND2_X1 U1063 ( .A1(n21573), .A2(n29322), .Z(n21607) );
  INV_X1 U23153 ( .I(n21832), .ZN(n15242) );
  NOR2_X1 U16913 ( .A1(n3539), .A2(n21781), .ZN(n17019) );
  NOR2_X1 U4390 ( .A1(n1135), .A2(n3468), .ZN(n8230) );
  NOR2_X1 U9583 ( .A1(n7553), .A2(n29234), .ZN(n13500) );
  INV_X1 U17358 ( .I(n32519), .ZN(n21701) );
  NOR2_X1 U17590 ( .A1(n29084), .A2(n11861), .ZN(n17018) );
  AOI22_X1 U5094 ( .A1(n21794), .A2(n15838), .B1(n21793), .B2(n21792), .ZN(
        n21795) );
  AOI21_X1 U7065 ( .A1(n21666), .A2(n1312), .B(n16577), .ZN(n2178) );
  NAND3_X1 U2935 ( .A1(n16194), .A2(n29302), .A3(n31458), .ZN(n21548) );
  OAI21_X1 U1054 ( .A1(n31335), .A2(n915), .B(n11499), .ZN(n11552) );
  OAI21_X1 U21991 ( .A1(n27704), .A2(n32865), .B(n1009), .ZN(n4131) );
  NOR2_X1 U14322 ( .A1(n27065), .A2(n1317), .ZN(n16163) );
  NAND2_X1 U8143 ( .A1(n5546), .A2(n1138), .ZN(n2709) );
  AOI22_X1 U2581 ( .A1(n2298), .A2(n21625), .B1(n2296), .B2(n396), .ZN(n2297)
         );
  NAND2_X1 U11391 ( .A1(n33146), .A2(n1133), .ZN(n4262) );
  NAND2_X1 U6381 ( .A1(n1647), .A2(n21520), .ZN(n1770) );
  NAND2_X1 U8142 ( .A1(n21852), .A2(n5546), .ZN(n2710) );
  NAND2_X1 U19647 ( .A1(n28729), .A2(n7813), .ZN(n12605) );
  NAND3_X1 U5817 ( .A1(n3467), .A2(n17077), .A3(n3468), .ZN(n3469) );
  NAND2_X1 U11298 ( .A1(n21701), .A2(n17887), .ZN(n15316) );
  INV_X1 U4658 ( .I(n27704), .ZN(n6967) );
  NAND2_X1 U19852 ( .A1(n12751), .A2(n32076), .ZN(n11448) );
  NAND2_X1 U9520 ( .A1(n21657), .A2(n8886), .ZN(n14829) );
  AOI21_X1 U5606 ( .A1(n21566), .A2(n3315), .B(n21570), .ZN(n3314) );
  OAI21_X1 U9543 ( .A1(n17019), .A2(n17018), .B(n31220), .ZN(n17017) );
  NAND2_X1 U1066 ( .A1(n30548), .A2(n3588), .ZN(n21525) );
  NAND2_X1 U7059 ( .A1(n7366), .A2(n7365), .ZN(n21680) );
  OAI22_X1 U1033 ( .A1(n32071), .A2(n30549), .B1(n21594), .B2(n21595), .ZN(
        n21597) );
  NAND2_X1 U7083 ( .A1(n1326), .A2(n15864), .ZN(n16012) );
  INV_X1 U26464 ( .I(n34084), .ZN(n1531) );
  OR2_X1 U519 ( .A1(n16796), .A2(n16192), .Z(n3722) );
  INV_X1 U3222 ( .I(n8269), .ZN(n1607) );
  OAI21_X1 U20926 ( .A1(n1531), .A2(n21804), .B(n11231), .ZN(n30999) );
  AOI22_X1 U9083 ( .A1(n29393), .A2(n3467), .B1(n1135), .B2(n4699), .ZN(n13540) );
  NOR2_X1 U22104 ( .A1(n21805), .A2(n3468), .ZN(n21722) );
  AOI22_X1 U15450 ( .A1(n26113), .A2(n16147), .B1(n6626), .B2(n1015), .ZN(
        n4880) );
  BUF_X2 U5093 ( .I(n17697), .Z(n4057) );
  NAND3_X1 U15766 ( .A1(n27103), .A2(n5757), .A3(n33571), .ZN(n30306) );
  BUF_X2 U15950 ( .I(n22249), .Z(n2353) );
  INV_X1 U11262 ( .I(n8392), .ZN(n1308) );
  INV_X1 U1042 ( .I(n22137), .ZN(n6812) );
  NAND2_X1 U11221 ( .A1(n910), .A2(n17362), .ZN(n6206) );
  INV_X1 U2271 ( .I(n34078), .ZN(n2308) );
  NAND2_X1 U1605 ( .A1(n26875), .A2(n22047), .ZN(n1609) );
  NAND2_X1 U13604 ( .A1(n21945), .A2(n12594), .ZN(n2777) );
  INV_X1 U7028 ( .I(n6771), .ZN(n22128) );
  INV_X1 U7618 ( .I(n27767), .ZN(n29501) );
  INV_X1 U13520 ( .I(n29693), .ZN(n26942) );
  INV_X1 U22737 ( .I(n22302), .ZN(n14125) );
  INV_X1 U1024 ( .I(n9809), .ZN(n21959) );
  INV_X1 U9481 ( .I(n22294), .ZN(n2554) );
  INV_X2 U26198 ( .I(n22681), .ZN(n31701) );
  INV_X1 U19066 ( .I(n8452), .ZN(n10680) );
  INV_X4 U13958 ( .I(n27004), .ZN(n22330) );
  INV_X2 U1253 ( .I(n5640), .ZN(n10724) );
  INV_X1 U3848 ( .I(n14307), .ZN(n22578) );
  INV_X1 U14614 ( .I(n32081), .ZN(n12530) );
  NAND2_X1 U16897 ( .A1(n33466), .A2(n22647), .ZN(n6187) );
  INV_X1 U5631 ( .I(n5657), .ZN(n12733) );
  BUF_X2 U4836 ( .I(n21941), .Z(n22645) );
  BUF_X2 U3296 ( .I(n22199), .Z(n11895) );
  INV_X1 U5800 ( .I(n34162), .ZN(n1119) );
  INV_X1 U3928 ( .I(n22332), .ZN(n2417) );
  INV_X1 U2741 ( .I(n22625), .ZN(n22497) );
  INV_X1 U18662 ( .I(n8099), .ZN(n22547) );
  INV_X2 U3076 ( .I(n16567), .ZN(n22666) );
  INV_X1 U20732 ( .I(n11749), .ZN(n16558) );
  INV_X1 U7048 ( .I(n27897), .ZN(n645) );
  INV_X1 U6713 ( .I(n10680), .ZN(n9456) );
  INV_X2 U1315 ( .I(n10568), .ZN(n14376) );
  INV_X2 U15233 ( .I(n22547), .ZN(n22550) );
  INV_X1 U8089 ( .I(n21869), .ZN(n22678) );
  INV_X1 U9468 ( .I(n8471), .ZN(n22398) );
  INV_X2 U13102 ( .I(n29304), .ZN(n905) );
  INV_X2 U3489 ( .I(n9515), .ZN(n22574) );
  NOR2_X1 U6687 ( .A1(n22681), .A2(n10354), .ZN(n9802) );
  CLKBUF_X2 U3705 ( .I(n22414), .Z(n137) );
  NOR2_X1 U5381 ( .A1(n16567), .A2(n16149), .ZN(n15805) );
  INV_X2 U19539 ( .I(n9234), .ZN(n9370) );
  BUF_X2 U4112 ( .I(n637), .Z(n14728) );
  INV_X2 U9463 ( .I(n9910), .ZN(n3495) );
  INV_X2 U23959 ( .I(n634), .ZN(n22626) );
  INV_X2 U456 ( .I(n12076), .ZN(n900) );
  INV_X1 U5798 ( .I(n22597), .ZN(n11930) );
  INV_X1 U1529 ( .I(n17879), .ZN(n22667) );
  INV_X2 U7757 ( .I(n9959), .ZN(n29508) );
  INV_X1 U11205 ( .I(n22452), .ZN(n6658) );
  INV_X1 U2047 ( .I(n22340), .ZN(n1300) );
  INV_X2 U4924 ( .I(n15089), .ZN(n11874) );
  NAND2_X1 U4369 ( .A1(n17147), .A2(n8965), .ZN(n18038) );
  OAI21_X1 U9399 ( .A1(n1290), .A2(n22588), .B(n22584), .ZN(n15007) );
  NAND3_X1 U5643 ( .A1(n2417), .A2(n16334), .A3(n12733), .ZN(n7053) );
  NAND2_X1 U22682 ( .A1(n14376), .A2(n29304), .ZN(n9751) );
  NOR3_X1 U6705 ( .A1(n29261), .A2(n900), .A3(n22394), .ZN(n13154) );
  NAND2_X1 U9430 ( .A1(n9578), .A2(n22599), .ZN(n9579) );
  OAI21_X1 U5373 ( .A1(n22401), .A2(n27390), .B(n32449), .ZN(n6749) );
  INV_X1 U4098 ( .I(n637), .ZN(n901) );
  NOR2_X1 U5670 ( .A1(n1116), .A2(n22672), .ZN(n12632) );
  NAND2_X1 U7637 ( .A1(n9022), .A2(n10612), .ZN(n11419) );
  NAND2_X1 U8014 ( .A1(n10206), .A2(n856), .ZN(n6709) );
  NAND2_X1 U421 ( .A1(n22389), .A2(n33966), .ZN(n17357) );
  INV_X2 U866 ( .I(n11932), .ZN(n26173) );
  INV_X1 U498 ( .I(n5379), .ZN(n904) );
  AOI21_X1 U5787 ( .A1(n22574), .A2(n16503), .B(n2471), .ZN(n12888) );
  INV_X1 U1443 ( .I(n2538), .ZN(n17123) );
  NAND2_X1 U926 ( .A1(n22549), .A2(n30668), .ZN(n25947) );
  INV_X2 U468 ( .I(n11920), .ZN(n22478) );
  BUF_X2 U21999 ( .I(n11916), .Z(n28669) );
  NAND2_X1 U13576 ( .A1(n468), .A2(n33964), .ZN(n22442) );
  INV_X1 U15542 ( .I(n33739), .ZN(n708) );
  INV_X2 U14853 ( .I(n28378), .ZN(n22483) );
  NAND2_X1 U3170 ( .A1(n4425), .A2(n22636), .ZN(n14478) );
  INV_X2 U5803 ( .I(n28825), .ZN(n4459) );
  AND2_X1 U21847 ( .A1(n22656), .A2(n17899), .Z(n22583) );
  INV_X1 U2749 ( .I(n1127), .ZN(n858) );
  NAND3_X1 U8208 ( .A1(n1125), .A2(n22584), .A3(n1290), .ZN(n29557) );
  BUF_X2 U4556 ( .I(n22580), .Z(n26878) );
  INV_X2 U826 ( .I(n17764), .ZN(n908) );
  INV_X1 U15795 ( .I(n9578), .ZN(n13078) );
  NOR3_X1 U19666 ( .A1(n16558), .A2(n31914), .A3(n22638), .ZN(n15609) );
  OAI21_X1 U7748 ( .A1(n15805), .A2(n22576), .B(n26453), .ZN(n27411) );
  AOI21_X1 U18298 ( .A1(n16531), .A2(n22612), .B(n855), .ZN(n7464) );
  INV_X1 U21751 ( .I(n468), .ZN(n22567) );
  NAND2_X1 U918 ( .A1(n22666), .A2(n22577), .ZN(n12439) );
  NAND2_X1 U13026 ( .A1(n1300), .A2(n22622), .ZN(n22623) );
  NAND3_X1 U3057 ( .A1(n1633), .A2(n2697), .A3(n28568), .ZN(n11376) );
  NOR2_X1 U18055 ( .A1(n22505), .A2(n14728), .ZN(n27574) );
  NOR2_X1 U11112 ( .A1(n22646), .A2(n4459), .ZN(n7850) );
  NAND2_X1 U1713 ( .A1(n22537), .A2(n17147), .ZN(n12698) );
  AOI21_X1 U6305 ( .A1(n1842), .A2(n30668), .B(n30669), .ZN(n22482) );
  NOR2_X1 U709 ( .A1(n16434), .A2(n8965), .ZN(n16549) );
  NOR2_X1 U11192 ( .A1(n22450), .A2(n17764), .ZN(n2657) );
  INV_X1 U7026 ( .I(n31931), .ZN(n22691) );
  NOR2_X1 U6715 ( .A1(n15752), .A2(n16483), .ZN(n14228) );
  NAND2_X1 U21038 ( .A1(n22475), .A2(n22474), .ZN(n17248) );
  AOI21_X1 U5377 ( .A1(n17185), .A2(n10862), .B(n8919), .ZN(n2486) );
  NAND2_X1 U20888 ( .A1(n8912), .A2(n17185), .ZN(n13874) );
  NOR2_X1 U9445 ( .A1(n16434), .A2(n22429), .ZN(n9425) );
  NOR3_X1 U835 ( .A1(n22330), .A2(n14376), .A3(n902), .ZN(n29957) );
  NOR2_X1 U8088 ( .A1(n1116), .A2(n905), .ZN(n29541) );
  NAND2_X1 U20828 ( .A1(n14231), .A2(n33966), .ZN(n15450) );
  OAI21_X1 U21257 ( .A1(n22576), .A2(n16567), .B(n6658), .ZN(n15379) );
  CLKBUF_X2 U12887 ( .I(n22599), .Z(n30066) );
  NOR2_X1 U874 ( .A1(n6401), .A2(n9653), .ZN(n6432) );
  AOI21_X1 U18640 ( .A1(n239), .A2(n7090), .B(n16137), .ZN(n2383) );
  NAND2_X1 U4829 ( .A1(n22402), .A2(n9739), .ZN(n13249) );
  INV_X1 U767 ( .I(n22634), .ZN(n1291) );
  NAND2_X1 U676 ( .A1(n5743), .A2(n9958), .ZN(n22924) );
  OAI21_X1 U8913 ( .A1(n17185), .A2(n26410), .B(n32449), .ZN(n26409) );
  INV_X1 U4346 ( .I(n29928), .ZN(n5960) );
  NAND2_X1 U2570 ( .A1(n2381), .A2(n7090), .ZN(n30510) );
  INV_X1 U7040 ( .I(n22486), .ZN(n1296) );
  INV_X1 U11166 ( .I(n7561), .ZN(n7560) );
  NAND2_X1 U25807 ( .A1(n1633), .A2(n17890), .ZN(n15448) );
  OAI22_X1 U848 ( .A1(n11928), .A2(n15379), .B1(n22454), .B2(n6658), .ZN(
        n26799) );
  NAND2_X1 U5683 ( .A1(n6956), .A2(n21963), .ZN(n29632) );
  AOI21_X1 U13557 ( .A1(n13525), .A2(n34058), .B(n22651), .ZN(n13524) );
  NAND2_X1 U9336 ( .A1(n11161), .A2(n22670), .ZN(n1579) );
  NAND3_X1 U5771 ( .A1(n10907), .A2(n28669), .A3(n8801), .ZN(n22459) );
  NAND2_X1 U3064 ( .A1(n22388), .A2(n1633), .ZN(n6063) );
  NAND2_X1 U2750 ( .A1(n7239), .A2(n6072), .ZN(n2408) );
  NAND3_X1 U18502 ( .A1(n13534), .A2(n12072), .A3(n22478), .ZN(n30631) );
  AOI21_X1 U8912 ( .A1(n17185), .A2(n8912), .B(n26409), .ZN(n26408) );
  OAI21_X1 U9341 ( .A1(n17960), .A2(n12335), .B(n12333), .ZN(n22011) );
  NOR2_X1 U18868 ( .A1(n7851), .A2(n7850), .ZN(n30688) );
  NAND2_X1 U12067 ( .A1(n26813), .A2(n1658), .ZN(n3670) );
  INV_X1 U11159 ( .I(n22633), .ZN(n7400) );
  NAND3_X1 U5372 ( .A1(n992), .A2(n1286), .A3(n10907), .ZN(n13895) );
  INV_X2 U15917 ( .I(n23056), .ZN(n31437) );
  NAND2_X1 U8430 ( .A1(n4100), .A2(n4459), .ZN(n5896) );
  INV_X1 U5654 ( .I(n22523), .ZN(n28938) );
  OAI21_X1 U12997 ( .A1(n29078), .A2(n17764), .B(n26867), .ZN(n4996) );
  NAND2_X1 U6276 ( .A1(n13895), .A2(n13892), .ZN(n4700) );
  NAND2_X1 U778 ( .A1(n7802), .A2(n22968), .ZN(n12471) );
  OAI21_X1 U9291 ( .A1(n32055), .A2(n12952), .B(n9580), .ZN(n229) );
  AOI22_X1 U792 ( .A1(n22594), .A2(n32831), .B1(n4918), .B2(n22651), .ZN(
        n29598) );
  OAI21_X1 U12930 ( .A1(n26065), .A2(n26862), .B(n1117), .ZN(n8667) );
  INV_X2 U773 ( .I(n22986), .ZN(n29242) );
  OAI21_X1 U11075 ( .A1(n5597), .A2(n1120), .B(n2253), .ZN(n2252) );
  NOR2_X1 U18443 ( .A1(n22471), .A2(n31019), .ZN(n17630) );
  NAND3_X1 U23174 ( .A1(n10282), .A2(n10354), .A3(n31701), .ZN(n22472) );
  BUF_X2 U12215 ( .I(n15299), .Z(n11268) );
  INV_X2 U21083 ( .I(n28077), .ZN(n641) );
  NAND2_X1 U1023 ( .A1(n16501), .A2(n16267), .ZN(n11018) );
  INV_X1 U2373 ( .I(n13129), .ZN(n6782) );
  INV_X2 U6924 ( .I(n22786), .ZN(n26667) );
  INV_X1 U18461 ( .I(n30868), .ZN(n1112) );
  INV_X1 U5065 ( .I(n17462), .ZN(n1269) );
  NOR2_X1 U6260 ( .A1(n26251), .A2(n23031), .ZN(n6876) );
  NAND2_X1 U2636 ( .A1(n15301), .A2(n17855), .ZN(n22761) );
  NOR2_X1 U21994 ( .A1(n26667), .A2(n32510), .ZN(n28648) );
  INV_X2 U15370 ( .I(n16280), .ZN(n16976) );
  NOR2_X1 U15232 ( .A1(n28313), .A2(n22894), .ZN(n12377) );
  INV_X2 U712 ( .I(n641), .ZN(n12259) );
  BUF_X2 U662 ( .I(n12701), .Z(n3891) );
  BUF_X2 U15662 ( .I(n13063), .Z(n28415) );
  CLKBUF_X2 U3498 ( .I(n22960), .Z(n8334) );
  INV_X2 U627 ( .I(n22951), .ZN(n28408) );
  INV_X2 U24869 ( .I(n31505), .ZN(n2635) );
  NAND2_X1 U17880 ( .A1(n28227), .A2(n31549), .ZN(n5205) );
  INV_X1 U12547 ( .I(n3670), .ZN(n22748) );
  INV_X2 U8649 ( .I(n29610), .ZN(n15718) );
  INV_X1 U4513 ( .I(n22950), .ZN(n2479) );
  INV_X1 U732 ( .I(n722), .ZN(n31358) );
  INV_X1 U17615 ( .I(n7802), .ZN(n22965) );
  INV_X1 U14395 ( .I(n23065), .ZN(n898) );
  INV_X1 U3479 ( .I(n22885), .ZN(n29958) );
  NAND2_X1 U699 ( .A1(n22983), .A2(n8040), .ZN(n28234) );
  NAND2_X1 U2728 ( .A1(n28974), .A2(n22933), .ZN(n2912) );
  NOR2_X1 U5679 ( .A1(n22780), .A2(n29175), .ZN(n29174) );
  NAND2_X1 U2128 ( .A1(n22473), .A2(n27589), .ZN(n7943) );
  BUF_X2 U10866 ( .I(n758), .Z(n26612) );
  AOI22_X1 U18597 ( .A1(n1278), .A2(n6975), .B1(n23010), .B2(n23014), .ZN(
        n23016) );
  OAI21_X1 U684 ( .A1(n27639), .A2(n23083), .B(n26243), .ZN(n30202) );
  NAND2_X1 U670 ( .A1(n13778), .A2(n27580), .ZN(n12417) );
  NAND2_X1 U9780 ( .A1(n28328), .A2(n29314), .ZN(n26499) );
  NAND2_X1 U678 ( .A1(n22946), .A2(n23034), .ZN(n5095) );
  AOI21_X1 U672 ( .A1(n897), .A2(n15704), .B(n10031), .ZN(n11084) );
  OAI21_X1 U6832 ( .A1(n23103), .A2(n23104), .B(n3600), .ZN(n5400) );
  NOR2_X1 U739 ( .A1(n23107), .A2(n23106), .ZN(n31455) );
  NAND2_X1 U6812 ( .A1(n17211), .A2(n27719), .ZN(n10895) );
  INV_X2 U560 ( .I(n10031), .ZN(n983) );
  NOR2_X1 U12893 ( .A1(n31358), .A2(n29384), .ZN(n26222) );
  AOI21_X1 U20900 ( .A1(n27798), .A2(n28680), .B(n22988), .ZN(n22993) );
  NOR2_X1 U528 ( .A1(n28867), .A2(n9213), .ZN(n15317) );
  NAND2_X1 U3557 ( .A1(n14129), .A2(n22968), .ZN(n23088) );
  NOR2_X1 U5704 ( .A1(n12259), .A2(n27556), .ZN(n27555) );
  INV_X1 U9289 ( .I(n22962), .ZN(n23081) );
  NAND2_X1 U2164 ( .A1(n22956), .A2(n987), .ZN(n6592) );
  NOR3_X1 U2816 ( .A1(n9293), .A2(n10031), .A3(n22876), .ZN(n10030) );
  INV_X1 U4115 ( .I(n22399), .ZN(n23043) );
  INV_X1 U361 ( .I(n22955), .ZN(n852) );
  NAND2_X1 U17164 ( .A1(n32119), .A2(n15851), .ZN(n5618) );
  INV_X1 U7917 ( .I(n31937), .ZN(n22866) );
  INV_X1 U4515 ( .I(n17161), .ZN(n1265) );
  INV_X1 U15674 ( .I(n22919), .ZN(n22880) );
  AND2_X1 U5336 ( .A1(n15324), .A2(n22856), .Z(n3296) );
  INV_X2 U741 ( .I(n28659), .ZN(n14188) );
  INV_X1 U3564 ( .I(n15501), .ZN(n989) );
  INV_X1 U5341 ( .I(n23070), .ZN(n1277) );
  AND2_X1 U4452 ( .A1(n6605), .A2(n22894), .Z(n22769) );
  CLKBUF_X2 U1181 ( .I(n14045), .Z(n16254) );
  NAND2_X1 U15665 ( .A1(n23034), .A2(n13063), .ZN(n22892) );
  NAND2_X1 U2611 ( .A1(n23033), .A2(n22894), .ZN(n23037) );
  INV_X1 U6965 ( .I(n23110), .ZN(n6453) );
  NOR2_X1 U14709 ( .A1(n6985), .A2(n23082), .ZN(n13396) );
  NAND3_X1 U546 ( .A1(n32868), .A2(n803), .A3(n14183), .ZN(n4710) );
  NAND3_X1 U23825 ( .A1(n1581), .A2(n22961), .A3(n8334), .ZN(n13365) );
  NAND3_X1 U14750 ( .A1(n18261), .A2(n986), .A3(n26667), .ZN(n22789) );
  OAI21_X1 U549 ( .A1(n4489), .A2(n23050), .B(n25994), .ZN(n4488) );
  NAND2_X1 U2318 ( .A1(n853), .A2(n23108), .ZN(n22614) );
  NAND2_X1 U9271 ( .A1(n14797), .A2(n33382), .ZN(n3851) );
  NAND3_X1 U2372 ( .A1(n28659), .A2(n22982), .A3(n22983), .ZN(n12702) );
  NAND3_X1 U355 ( .A1(n6800), .A2(n22655), .A3(n28408), .ZN(n22276) );
  AOI21_X1 U14942 ( .A1(n22876), .A2(n10031), .B(n11268), .ZN(n15298) );
  NAND2_X1 U15880 ( .A1(n898), .A2(n22826), .ZN(n22863) );
  NAND3_X1 U23053 ( .A1(n32868), .A2(n23158), .A3(n13751), .ZN(n4713) );
  NAND2_X1 U16748 ( .A1(n22738), .A2(n14610), .ZN(n8381) );
  NOR3_X1 U2583 ( .A1(n990), .A2(n1278), .A3(n4599), .ZN(n4652) );
  NOR2_X1 U21258 ( .A1(n13159), .A2(n16078), .ZN(n13635) );
  NOR2_X1 U4506 ( .A1(n23079), .A2(n22885), .ZN(n13411) );
  OAI21_X1 U11008 ( .A1(n29242), .A2(n31867), .B(n28328), .ZN(n7744) );
  NOR2_X1 U23542 ( .A1(n6592), .A2(n9778), .ZN(n6591) );
  NOR2_X1 U19423 ( .A1(n23111), .A2(n1264), .ZN(n27835) );
  NAND2_X1 U2269 ( .A1(n6012), .A2(n16022), .ZN(n22725) );
  NAND2_X1 U7928 ( .A1(n22760), .A2(n27612), .ZN(n22410) );
  NAND2_X1 U17430 ( .A1(n10360), .A2(n27389), .ZN(n6370) );
  NOR2_X1 U21543 ( .A1(n31854), .A2(n22780), .ZN(n22739) );
  NOR2_X1 U25150 ( .A1(n28867), .A2(n23101), .ZN(n22842) );
  NAND2_X1 U20488 ( .A1(n18240), .A2(n22774), .ZN(n11204) );
  OAI21_X1 U6919 ( .A1(n22762), .A2(n28314), .B(n12726), .ZN(n14680) );
  AOI21_X1 U10869 ( .A1(n22698), .A2(n30960), .B(n5689), .ZN(n22699) );
  NAND2_X1 U10953 ( .A1(n4805), .A2(n29648), .ZN(n4804) );
  NAND2_X1 U642 ( .A1(n28071), .A2(n22964), .ZN(n3692) );
  NOR2_X1 U13006 ( .A1(n28867), .A2(n985), .ZN(n30168) );
  NOR2_X1 U8698 ( .A1(n30488), .A2(n31455), .ZN(n4174) );
  NAND2_X1 U17761 ( .A1(n32088), .A2(n26526), .ZN(n14769) );
  OAI21_X1 U9446 ( .A1(n6149), .A2(n29325), .B(n33382), .ZN(n6148) );
  NOR2_X1 U3266 ( .A1(n16142), .A2(n16236), .ZN(n16993) );
  NOR2_X1 U2589 ( .A1(n27798), .A2(n22986), .ZN(n22864) );
  NAND2_X1 U12020 ( .A1(n27090), .A2(n29967), .ZN(n16514) );
  CLKBUF_X2 U625 ( .I(n31942), .Z(n3999) );
  INV_X1 U520 ( .I(n5620), .ZN(n5055) );
  NAND2_X1 U2342 ( .A1(n23045), .A2(n22795), .ZN(n15580) );
  NAND2_X1 U10913 ( .A1(n7047), .A2(n5178), .ZN(n5182) );
  OR2_X1 U17891 ( .A1(n4599), .A2(n14540), .Z(n14212) );
  OAI21_X1 U5749 ( .A1(n26507), .A2(n22901), .B(n15601), .ZN(n18177) );
  NAND3_X1 U9238 ( .A1(n802), .A2(n10031), .A3(n9293), .ZN(n11108) );
  OAI22_X1 U326 ( .A1(n12762), .A2(n32089), .B1(n22866), .B2(n1277), .ZN(n4268) );
  NAND2_X1 U9256 ( .A1(n22981), .A2(n2130), .ZN(n2111) );
  NOR2_X1 U6918 ( .A1(n30365), .A2(n28649), .ZN(n3174) );
  NAND2_X1 U16007 ( .A1(n4649), .A2(n990), .ZN(n4650) );
  OAI21_X1 U626 ( .A1(n29430), .A2(n29477), .B(n27589), .ZN(n7724) );
  NAND2_X1 U9252 ( .A1(n8084), .A2(n26373), .ZN(n7356) );
  AOI22_X1 U640 ( .A1(n23064), .A2(n30437), .B1(n10643), .B2(n1275), .ZN(
        n30080) );
  NAND3_X1 U20254 ( .A1(n13916), .A2(n22914), .A3(n12071), .ZN(n15341) );
  NOR2_X1 U18113 ( .A1(n8149), .A2(n8150), .ZN(n31394) );
  OAI21_X1 U7777 ( .A1(n17639), .A2(n28948), .B(n6236), .ZN(n26274) );
  BUF_X2 U26320 ( .I(n15341), .Z(n29190) );
  NAND2_X1 U5620 ( .A1(n14623), .A2(n11873), .ZN(n30741) );
  OAI21_X1 U7776 ( .A1(n14192), .A2(n6236), .B(n26274), .ZN(n11162) );
  BUF_X2 U1273 ( .I(n23453), .Z(n438) );
  INV_X1 U15079 ( .I(n30532), .ZN(n23461) );
  INV_X1 U22465 ( .I(n23273), .ZN(n23503) );
  INV_X1 U3603 ( .I(n23489), .ZN(n13216) );
  INV_X1 U4004 ( .I(n17871), .ZN(n23462) );
  NAND2_X1 U19931 ( .A1(n29160), .A2(n1260), .ZN(n3408) );
  NAND2_X1 U16062 ( .A1(n26900), .A2(n27457), .ZN(n30319) );
  CLKBUF_X2 U5750 ( .I(n6386), .Z(n3739) );
  INV_X1 U5049 ( .I(n23439), .ZN(n23413) );
  INV_X1 U600 ( .I(n13347), .ZN(n27220) );
  INV_X1 U589 ( .I(n23936), .ZN(n30949) );
  INV_X1 U24264 ( .I(n28611), .ZN(n14297) );
  INV_X1 U9219 ( .I(n17812), .ZN(n23951) );
  INV_X1 U9678 ( .I(n29704), .ZN(n28069) );
  INV_X1 U23439 ( .I(n15917), .ZN(n23578) );
  INV_X2 U3607 ( .I(n10213), .ZN(n801) );
  INV_X1 U11171 ( .I(n23765), .ZN(n29865) );
  INV_X1 U5696 ( .I(n30949), .ZN(n17181) );
  CLKBUF_X2 U4656 ( .I(n13361), .Z(n29185) );
  INV_X2 U13110 ( .I(n23735), .ZN(n1489) );
  INV_X1 U26258 ( .I(n29139), .ZN(n29271) );
  CLKBUF_X2 U5596 ( .I(n6474), .Z(n31179) );
  BUF_X2 U10829 ( .I(n23886), .Z(n17234) );
  INV_X1 U17601 ( .I(n9796), .ZN(n10279) );
  INV_X2 U2871 ( .I(n23201), .ZN(n4177) );
  INV_X1 U21008 ( .I(n28069), .ZN(n8045) );
  INV_X1 U14135 ( .I(n3169), .ZN(n8838) );
  INV_X1 U14960 ( .I(n23951), .ZN(n14473) );
  INV_X1 U19037 ( .I(n16563), .ZN(n23759) );
  OR2_X1 U4625 ( .A1(n17285), .A2(n17352), .Z(n23906) );
  INV_X1 U25858 ( .I(n28847), .ZN(n548) );
  INV_X1 U1857 ( .I(n23586), .ZN(n23910) );
  INV_X1 U9217 ( .I(n23754), .ZN(n12433) );
  INV_X1 U23116 ( .I(n16961), .ZN(n23945) );
  INV_X1 U309 ( .I(n29270), .ZN(n979) );
  INV_X1 U17142 ( .I(n14255), .ZN(n14164) );
  INV_X1 U282 ( .I(n23745), .ZN(n11567) );
  INV_X2 U19149 ( .I(n16333), .ZN(n8544) );
  AND2_X1 U5036 ( .A1(n2450), .A2(n23706), .Z(n2460) );
  INV_X1 U3606 ( .I(n499), .ZN(n10217) );
  NOR3_X1 U3536 ( .A1(n14473), .A2(n8217), .A3(n979), .ZN(n16862) );
  AOI21_X1 U23772 ( .A1(n981), .A2(n354), .B(n11888), .ZN(n17616) );
  NAND2_X1 U19360 ( .A1(n10213), .A2(n23871), .ZN(n23694) );
  NAND2_X1 U6850 ( .A1(n2460), .A2(n23782), .ZN(n9278) );
  NOR2_X1 U21773 ( .A1(n10217), .A2(n756), .ZN(n12094) );
  INV_X2 U6894 ( .I(n23786), .ZN(n23903) );
  AOI21_X1 U22127 ( .A1(n27678), .A2(n1257), .B(n844), .ZN(n31163) );
  INV_X1 U1916 ( .I(n23611), .ZN(n769) );
  BUF_X2 U5610 ( .I(n9430), .Z(n31890) );
  INV_X2 U400 ( .I(n6474), .ZN(n28367) );
  NAND2_X1 U16638 ( .A1(n23765), .A2(n23764), .ZN(n23923) );
  CLKBUF_X2 U5832 ( .I(n23755), .Z(n28222) );
  INV_X2 U15327 ( .I(n1099), .ZN(n978) );
  BUF_X2 U4222 ( .I(n23764), .Z(n28676) );
  INV_X2 U273 ( .I(n23756), .ZN(n23749) );
  INV_X2 U23685 ( .I(n28266), .ZN(n23891) );
  INV_X1 U5332 ( .I(n12974), .ZN(n17872) );
  INV_X1 U11142 ( .I(n26641), .ZN(n6394) );
  INV_X1 U292 ( .I(n23764), .ZN(n16337) );
  NAND2_X1 U16578 ( .A1(n5373), .A2(n299), .ZN(n5372) );
  INV_X1 U6176 ( .I(n23755), .ZN(n23726) );
  INV_X1 U7341 ( .I(n32711), .ZN(n23897) );
  INV_X1 U1464 ( .I(n27), .ZN(n23798) );
  INV_X1 U15458 ( .I(n31796), .ZN(n1254) );
  INV_X1 U4493 ( .I(n17245), .ZN(n7073) );
  NOR2_X1 U561 ( .A1(n27678), .A2(n8655), .ZN(n8654) );
  CLKBUF_X2 U13176 ( .I(n23742), .Z(n30089) );
  NOR2_X1 U3039 ( .A1(n31916), .A2(n29268), .ZN(n7140) );
  INV_X1 U464 ( .I(n9172), .ZN(n3687) );
  AOI21_X1 U9596 ( .A1(n29240), .A2(n33337), .B(n23841), .ZN(n17950) );
  INV_X1 U1595 ( .I(n30282), .ZN(n5163) );
  NOR2_X1 U23877 ( .A1(n893), .A2(n30059), .ZN(n23660) );
  NOR2_X1 U6177 ( .A1(n23778), .A2(n8547), .ZN(n15658) );
  NAND2_X1 U13682 ( .A1(n7005), .A2(n23910), .ZN(n1641) );
  OAI21_X1 U6897 ( .A1(n980), .A2(n23885), .B(n9278), .ZN(n9277) );
  NOR2_X1 U6193 ( .A1(n23855), .A2(n4177), .ZN(n2233) );
  NAND2_X1 U8486 ( .A1(n2023), .A2(n23793), .ZN(n23569) );
  INV_X1 U366 ( .I(n23753), .ZN(n26397) );
  NAND2_X1 U25144 ( .A1(n31938), .A2(n976), .ZN(n22833) );
  NAND2_X1 U386 ( .A1(n16343), .A2(n16496), .ZN(n26185) );
  NAND2_X1 U22389 ( .A1(n31435), .A2(n26114), .ZN(n31209) );
  NOR2_X1 U9389 ( .A1(n12722), .A2(n23611), .ZN(n26465) );
  INV_X1 U5031 ( .I(n11708), .ZN(n23811) );
  INV_X1 U18430 ( .I(n23877), .ZN(n30621) );
  BUF_X2 U550 ( .I(n14974), .Z(n28210) );
  NAND2_X1 U15352 ( .A1(n5372), .A2(n27474), .ZN(n4340) );
  NOR2_X1 U19677 ( .A1(n4319), .A2(n11968), .ZN(n17612) );
  INV_X1 U253 ( .I(n23672), .ZN(n144) );
  OAI21_X1 U6878 ( .A1(n11923), .A2(n23888), .B(n6479), .ZN(n11673) );
  AOI21_X1 U488 ( .A1(n30295), .A2(n30296), .B(n28676), .ZN(n30294) );
  NOR2_X1 U13380 ( .A1(n23704), .A2(n32308), .ZN(n17922) );
  NOR2_X1 U5714 ( .A1(n11050), .A2(n23708), .ZN(n23880) );
  NOR2_X1 U22780 ( .A1(n28266), .A2(n18133), .ZN(n23895) );
  AOI21_X1 U9156 ( .A1(n7073), .A2(n1256), .B(n1253), .ZN(n3371) );
  NAND2_X1 U20319 ( .A1(n29218), .A2(n10187), .ZN(n23558) );
  NOR2_X1 U484 ( .A1(n23891), .A2(n23892), .ZN(n30527) );
  INV_X1 U15323 ( .I(n23578), .ZN(n11096) );
  INV_X1 U3038 ( .I(n31916), .ZN(n3481) );
  INV_X1 U4242 ( .I(n10279), .ZN(n23787) );
  BUF_X2 U5608 ( .I(n17157), .Z(n14973) );
  INV_X1 U26617 ( .I(n23765), .ZN(n17087) );
  NAND2_X1 U6862 ( .A1(n14325), .A2(n23806), .ZN(n23805) );
  INV_X1 U2778 ( .I(n1098), .ZN(n27615) );
  CLKBUF_X2 U4793 ( .I(n893), .Z(n5357) );
  NAND2_X1 U16972 ( .A1(n23600), .A2(n6247), .ZN(n27369) );
  NAND2_X1 U26172 ( .A1(n11673), .A2(n23841), .ZN(n31690) );
  NAND2_X1 U13770 ( .A1(n10213), .A2(n6474), .ZN(n3401) );
  OAI21_X1 U25334 ( .A1(n6414), .A2(n16238), .B(n23906), .ZN(n23707) );
  INV_X1 U10760 ( .I(n23805), .ZN(n9900) );
  NOR2_X1 U16717 ( .A1(n23895), .A2(n29068), .ZN(n5555) );
  NOR2_X1 U446 ( .A1(n28855), .A2(n3687), .ZN(n9645) );
  OAI21_X1 U6909 ( .A1(n12528), .A2(n23782), .B(n11240), .ZN(n12527) );
  NAND3_X1 U25318 ( .A1(n23884), .A2(n756), .A3(n33936), .ZN(n23635) );
  NOR2_X1 U6890 ( .A1(n23953), .A2(n3481), .ZN(n7383) );
  NAND2_X1 U16991 ( .A1(n12658), .A2(n667), .ZN(n30409) );
  AOI22_X1 U449 ( .A1(n9002), .A2(n11621), .B1(n10753), .B2(n30359), .ZN(
        n30169) );
  OAI21_X1 U5297 ( .A1(n17750), .A2(n23773), .B(n23778), .ZN(n8719) );
  NOR2_X1 U5702 ( .A1(n23866), .A2(n843), .ZN(n24000) );
  NAND2_X1 U19527 ( .A1(n31179), .A2(n23871), .ZN(n28728) );
  NAND2_X1 U16718 ( .A1(n32434), .A2(n28266), .ZN(n5556) );
  OAI21_X1 U6911 ( .A1(n23953), .A2(n31601), .B(n29372), .ZN(n23564) );
  NAND2_X1 U25345 ( .A1(n23776), .A2(n8547), .ZN(n23747) );
  AOI21_X1 U13808 ( .A1(n3480), .A2(n16686), .B(n23953), .ZN(n28534) );
  INV_X1 U24612 ( .I(n14513), .ZN(n31479) );
  NOR2_X1 U6888 ( .A1(n29372), .A2(n4991), .ZN(n26837) );
  NAND2_X1 U415 ( .A1(n9382), .A2(n313), .ZN(n27811) );
  NAND2_X1 U25323 ( .A1(n23656), .A2(n23746), .ZN(n23657) );
  OAI21_X1 U420 ( .A1(n16969), .A2(n29474), .B(n23741), .ZN(n29795) );
  OAI21_X1 U6905 ( .A1(n15659), .A2(n15658), .B(n16271), .ZN(n31058) );
  OAI21_X1 U15194 ( .A1(n29269), .A2(n10993), .B(n23681), .ZN(n14124) );
  AOI22_X1 U3500 ( .A1(n15272), .A2(n10143), .B1(n4319), .B2(n23638), .ZN(
        n28850) );
  OAI21_X1 U14941 ( .A1(n23947), .A2(n13308), .B(n29294), .ZN(n1528) );
  AOI21_X1 U22047 ( .A1(n23493), .A2(n29240), .B(n31158), .ZN(n11492) );
  NAND2_X1 U23589 ( .A1(n28503), .A2(n23654), .ZN(n23658) );
  NAND2_X1 U21432 ( .A1(n8836), .A2(n5357), .ZN(n31082) );
  OAI21_X1 U12619 ( .A1(n23697), .A2(n11943), .B(n9772), .ZN(n30028) );
  NOR2_X1 U7816 ( .A1(n23896), .A2(n27615), .ZN(n10480) );
  OR2_X1 U15428 ( .A1(n23856), .A2(n25996), .Z(n9214) );
  NAND2_X1 U6854 ( .A1(n23704), .A2(n34008), .ZN(n4539) );
  NAND3_X1 U6861 ( .A1(n7073), .A2(n1253), .A3(n16677), .ZN(n7074) );
  AOI21_X1 U26068 ( .A1(n23593), .A2(n23891), .B(n23892), .ZN(n6723) );
  NAND2_X1 U12616 ( .A1(n30028), .A2(n33924), .ZN(n9770) );
  NOR2_X1 U3263 ( .A1(n10019), .A2(n10020), .ZN(n29699) );
  NAND2_X1 U340 ( .A1(n1920), .A2(n31890), .ZN(n14047) );
  NOR2_X1 U24501 ( .A1(n28637), .A2(n16118), .ZN(n4483) );
  NOR2_X1 U4089 ( .A1(n12722), .A2(n769), .ZN(n24331) );
  INV_X1 U18096 ( .I(n30505), .ZN(n1090) );
  INV_X1 U2017 ( .I(n24315), .ZN(n797) );
  INV_X2 U5280 ( .I(n24014), .ZN(n974) );
  INV_X1 U210 ( .I(n12374), .ZN(n1245) );
  NAND2_X1 U15615 ( .A1(n24159), .A2(n29157), .ZN(n9977) );
  BUF_X2 U3331 ( .I(n10226), .Z(n9275) );
  INV_X1 U21919 ( .I(n12356), .ZN(n23970) );
  NOR2_X1 U8247 ( .A1(n3667), .A2(n29561), .ZN(n5199) );
  INV_X2 U14704 ( .I(n3077), .ZN(n3148) );
  NAND2_X1 U283 ( .A1(n4655), .A2(n17261), .ZN(n24228) );
  INV_X2 U5877 ( .I(n26387), .ZN(n13343) );
  INV_X1 U8802 ( .I(n24207), .ZN(n24157) );
  INV_X2 U22219 ( .I(n13175), .ZN(n1244) );
  INV_X2 U8767 ( .I(n6713), .ZN(n737) );
  INV_X2 U6973 ( .I(n7465), .ZN(n793) );
  INV_X1 U6834 ( .I(n24164), .ZN(n14840) );
  NOR2_X1 U26170 ( .A1(n11503), .A2(n9616), .ZN(n1550) );
  INV_X1 U226 ( .I(n4655), .ZN(n16621) );
  INV_X1 U201 ( .I(n24087), .ZN(n24139) );
  INV_X2 U227 ( .I(n13223), .ZN(n24251) );
  INV_X1 U197 ( .I(n24141), .ZN(n7203) );
  INV_X1 U12982 ( .I(n6555), .ZN(n9146) );
  NAND2_X1 U7907 ( .A1(n24052), .A2(n24053), .ZN(n9976) );
  INV_X1 U301 ( .I(n24240), .ZN(n29043) );
  INV_X1 U200 ( .I(n24218), .ZN(n1240) );
  INV_X1 U12733 ( .I(n23748), .ZN(n15096) );
  INV_X1 U4781 ( .I(n24180), .ZN(n13260) );
  INV_X1 U22429 ( .I(n16215), .ZN(n796) );
  NAND2_X1 U13827 ( .A1(n33763), .A2(n24216), .ZN(n5098) );
  INV_X1 U3086 ( .I(n3421), .ZN(n24134) );
  INV_X1 U1970 ( .I(n6319), .ZN(n24013) );
  NOR2_X1 U3838 ( .A1(n24114), .A2(n24283), .ZN(n23961) );
  NAND2_X1 U21617 ( .A1(n16621), .A2(n28694), .ZN(n17940) );
  INV_X1 U220 ( .I(n16868), .ZN(n972) );
  NOR2_X1 U11016 ( .A1(n27104), .A2(n3077), .ZN(n29848) );
  NOR2_X1 U6940 ( .A1(n30289), .A2(n15068), .ZN(n31071) );
  NAND2_X1 U17734 ( .A1(n7546), .A2(n24221), .ZN(n11535) );
  NAND2_X1 U2068 ( .A1(n6003), .A2(n12356), .ZN(n5437) );
  NAND2_X1 U9138 ( .A1(n32917), .A2(n23970), .ZN(n26674) );
  BUF_X2 U4111 ( .I(n5199), .Z(n29141) );
  NAND2_X1 U6114 ( .A1(n9323), .A2(n8178), .ZN(n2247) );
  INV_X1 U14628 ( .I(n33832), .ZN(n14542) );
  BUF_X2 U1757 ( .I(n3718), .Z(n8) );
  CLKBUF_X2 U4215 ( .I(n17426), .Z(n8165) );
  NAND2_X1 U9102 ( .A1(n24052), .A2(n24185), .ZN(n24123) );
  INV_X2 U14723 ( .I(n24052), .ZN(n11463) );
  INV_X1 U271 ( .I(n29307), .ZN(n24272) );
  NAND2_X1 U6951 ( .A1(n24230), .A2(n31355), .ZN(n14861) );
  INV_X1 U2802 ( .I(n14195), .ZN(n14443) );
  INV_X1 U18877 ( .I(n2558), .ZN(n7150) );
  NOR2_X1 U6108 ( .A1(n2744), .A2(n31377), .ZN(n13170) );
  INV_X1 U374 ( .I(n1808), .ZN(n24237) );
  INV_X1 U10162 ( .I(n29157), .ZN(n29748) );
  INV_X1 U2784 ( .I(n9616), .ZN(n5308) );
  OAI21_X1 U13027 ( .A1(n4118), .A2(n4775), .B(n24134), .ZN(n17860) );
  NAND2_X1 U193 ( .A1(n10188), .A2(n13260), .ZN(n17943) );
  NAND3_X1 U25398 ( .A1(n24118), .A2(n24223), .A3(n24225), .ZN(n24119) );
  NAND2_X1 U15765 ( .A1(n792), .A2(n27104), .ZN(n2798) );
  NAND2_X1 U17015 ( .A1(n27661), .A2(n1240), .ZN(n6251) );
  NOR2_X1 U18960 ( .A1(n24092), .A2(n31096), .ZN(n30696) );
  NAND2_X1 U10574 ( .A1(n26027), .A2(n4024), .ZN(n3217) );
  NOR2_X1 U2115 ( .A1(n24292), .A2(n32936), .ZN(n24294) );
  INV_X1 U9057 ( .I(n13378), .ZN(n3603) );
  NOR2_X1 U12857 ( .A1(n891), .A2(n33597), .ZN(n23962) );
  INV_X1 U1991 ( .I(n24005), .ZN(n3903) );
  NOR2_X1 U2446 ( .A1(n32917), .A2(n17404), .ZN(n23701) );
  INV_X1 U152 ( .I(n24206), .ZN(n24009) );
  OAI21_X1 U11014 ( .A1(n10938), .A2(n29848), .B(n24268), .ZN(n31297) );
  NAND2_X1 U21830 ( .A1(n5631), .A2(n12143), .ZN(n24297) );
  INV_X1 U15608 ( .I(n24159), .ZN(n24124) );
  NAND2_X1 U20738 ( .A1(n9892), .A2(n14336), .ZN(n31868) );
  NOR2_X1 U327 ( .A1(n12862), .A2(n27661), .ZN(n27334) );
  NAND2_X1 U9711 ( .A1(n7779), .A2(n10104), .ZN(n28351) );
  NAND3_X1 U3078 ( .A1(n24027), .A2(n28040), .A3(n31002), .ZN(n24029) );
  NOR2_X1 U15567 ( .A1(n27436), .A2(n6476), .ZN(n11950) );
  OR2_X1 U5259 ( .A1(n11535), .A2(n3506), .Z(n11534) );
  NAND2_X1 U5474 ( .A1(n24182), .A2(n31722), .ZN(n17100) );
  NOR2_X1 U10590 ( .A1(n17232), .A2(n3506), .ZN(n17016) );
  NAND2_X1 U13737 ( .A1(n26459), .A2(n24093), .ZN(n29123) );
  INV_X1 U3611 ( .I(n24270), .ZN(n11721) );
  OAI22_X1 U9040 ( .A1(n7149), .A2(n15179), .B1(n14399), .B2(n29120), .ZN(
        n6877) );
  AOI21_X1 U10554 ( .A1(n11997), .A2(n12576), .B(n28040), .ZN(n10667) );
  NAND2_X1 U288 ( .A1(n30348), .A2(n24313), .ZN(n7483) );
  NAND2_X1 U15675 ( .A1(n14861), .A2(n11743), .ZN(n11742) );
  NAND2_X1 U17877 ( .A1(n27550), .A2(n32465), .ZN(n14724) );
  NAND3_X1 U18410 ( .A1(n24091), .A2(n16535), .A3(n24234), .ZN(n24655) );
  NAND2_X1 U9621 ( .A1(n24052), .A2(n24159), .ZN(n24183) );
  NAND2_X1 U20110 ( .A1(n33763), .A2(n31497), .ZN(n24109) );
  INV_X1 U6146 ( .I(n24220), .ZN(n1094) );
  NAND2_X1 U9079 ( .A1(n11463), .A2(n24053), .ZN(n30726) );
  INV_X1 U155 ( .I(n24216), .ZN(n24290) );
  INV_X1 U13048 ( .I(n11883), .ZN(n24233) );
  AND2_X1 U7357 ( .A1(n4286), .A2(n16052), .Z(n29473) );
  INV_X1 U214 ( .I(n28827), .ZN(n3219) );
  NAND2_X1 U308 ( .A1(n28300), .A2(n891), .ZN(n16683) );
  NOR2_X1 U19081 ( .A1(n3506), .A2(n7546), .ZN(n30715) );
  NAND3_X1 U7798 ( .A1(n24185), .A2(n11463), .A3(n1088), .ZN(n11461) );
  NOR2_X1 U1551 ( .A1(n24118), .A2(n10118), .ZN(n10117) );
  NAND3_X1 U7771 ( .A1(n2847), .A2(n24163), .A3(n24002), .ZN(n23988) );
  NAND2_X1 U20755 ( .A1(n23995), .A2(n24270), .ZN(n24385) );
  NAND3_X1 U189 ( .A1(n6001), .A2(n26516), .A3(n17404), .ZN(n17493) );
  OAI21_X1 U19785 ( .A1(n31113), .A2(n24290), .B(n11613), .ZN(n30826) );
  NAND3_X1 U5001 ( .A1(n33597), .A2(n7546), .A3(n24286), .ZN(n5307) );
  NAND2_X1 U18351 ( .A1(n24046), .A2(n13950), .ZN(n17233) );
  NAND2_X1 U23100 ( .A1(n24249), .A2(n24248), .ZN(n15085) );
  NAND2_X1 U284 ( .A1(n16683), .A2(n28409), .ZN(n30417) );
  NOR3_X1 U4996 ( .A1(n24202), .A2(n738), .A3(n27501), .ZN(n12262) );
  AOI21_X1 U8664 ( .A1(n31679), .A2(n23748), .B(n1499), .ZN(n1497) );
  NAND2_X1 U10635 ( .A1(n24273), .A2(n31918), .ZN(n11724) );
  NOR2_X1 U19113 ( .A1(n30726), .A2(n1088), .ZN(n26307) );
  OAI21_X1 U10571 ( .A1(n11950), .A2(n3632), .B(n28296), .ZN(n3631) );
  NOR2_X1 U291 ( .A1(n24107), .A2(n891), .ZN(n30096) );
  NAND3_X1 U9904 ( .A1(n2865), .A2(n27786), .A3(n31096), .ZN(n2186) );
  NAND2_X1 U5439 ( .A1(n31544), .A2(n31543), .ZN(n9367) );
  AOI21_X1 U6109 ( .A1(n12693), .A2(n12692), .B(n32917), .ZN(n12691) );
  NAND2_X1 U15924 ( .A1(n8142), .A2(n5490), .ZN(n24017) );
  AOI21_X1 U18278 ( .A1(n31002), .A2(n12982), .B(n28040), .ZN(n30598) );
  NAND2_X1 U11543 ( .A1(n5631), .A2(n24292), .ZN(n12429) );
  INV_X1 U5164 ( .I(n12868), .ZN(n2424) );
  NAND4_X1 U13150 ( .A1(n24343), .A2(n24342), .A3(n24344), .A4(n24341), .ZN(
        n31311) );
  NOR2_X1 U143 ( .A1(n28590), .A2(n9066), .ZN(n11042) );
  NAND2_X1 U279 ( .A1(n14445), .A2(n14444), .ZN(n31788) );
  BUF_X2 U3234 ( .I(n7679), .Z(n356) );
  CLKBUF_X2 U18973 ( .I(n24544), .Z(n27733) );
  INV_X2 U1275 ( .I(n5970), .ZN(n9907) );
  INV_X1 U10527 ( .I(n24393), .ZN(n8703) );
  BUF_X2 U5162 ( .I(n12868), .Z(n28977) );
  NOR2_X1 U13673 ( .A1(n16815), .A2(n26966), .ZN(n3295) );
  INV_X1 U2483 ( .I(n24805), .ZN(n14533) );
  NAND2_X1 U4747 ( .A1(n2421), .A2(n2420), .ZN(n17682) );
  CLKBUF_X2 U5418 ( .I(n24843), .Z(n10870) );
  INV_X1 U21378 ( .I(n28119), .ZN(n4886) );
  INV_X1 U4984 ( .I(n679), .ZN(n25397) );
  INV_X1 U19889 ( .I(n9932), .ZN(n10062) );
  INV_X1 U12755 ( .I(n25707), .ZN(n31570) );
  INV_X1 U2814 ( .I(n25394), .ZN(n13993) );
  BUF_X2 U15333 ( .I(n23668), .Z(n25871) );
  INV_X2 U5247 ( .I(n16957), .ZN(n9917) );
  INV_X1 U112 ( .I(n25536), .ZN(n833) );
  BUF_X2 U14756 ( .I(n25111), .Z(n25234) );
  INV_X1 U8982 ( .I(n25238), .ZN(n6910) );
  INV_X1 U115 ( .I(n5020), .ZN(n11987) );
  INV_X1 U14347 ( .I(n27072), .ZN(n17655) );
  INV_X1 U5957 ( .I(n25699), .ZN(n751) );
  INV_X1 U22211 ( .I(n24360), .ZN(n13042) );
  INV_X1 U235 ( .I(n680), .ZN(n24973) );
  INV_X1 U88 ( .I(n17240), .ZN(n885) );
  INV_X2 U2134 ( .I(n17655), .ZN(n25633) );
  NAND2_X1 U5956 ( .A1(n25867), .A2(n14111), .ZN(n10549) );
  INV_X1 U2638 ( .I(n10199), .ZN(n17839) );
  INV_X2 U5601 ( .I(n8219), .ZN(n1216) );
  NAND2_X1 U20653 ( .A1(n1567), .A2(n2092), .ZN(n30948) );
  INV_X1 U4981 ( .I(n15777), .ZN(n25870) );
  INV_X1 U4056 ( .I(n13993), .ZN(n11704) );
  NAND2_X1 U2860 ( .A1(n16632), .A2(n1786), .ZN(n27479) );
  INV_X1 U128 ( .I(n25766), .ZN(n27359) );
  CLKBUF_X2 U2509 ( .I(n25699), .Z(n28242) );
  INV_X1 U6777 ( .I(n15719), .ZN(n24983) );
  NAND2_X1 U8968 ( .A1(n11945), .A2(n15046), .ZN(n24609) );
  NOR2_X1 U188 ( .A1(n24361), .A2(n17118), .ZN(n30907) );
  BUF_X2 U2813 ( .I(n18156), .Z(n5202) );
  INV_X2 U5612 ( .I(n17963), .ZN(n25901) );
  INV_X2 U106 ( .I(n29629), .ZN(n14055) );
  INV_X1 U25721 ( .I(n25763), .ZN(n25704) );
  INV_X1 U80 ( .I(n11957), .ZN(n754) );
  INV_X1 U14968 ( .I(n18242), .ZN(n836) );
  NAND2_X1 U190 ( .A1(n25977), .A2(n11947), .ZN(n25239) );
  INV_X1 U13661 ( .I(n8892), .ZN(n25587) );
  INV_X1 U19564 ( .I(n28591), .ZN(n13709) );
  INV_X1 U3522 ( .I(n29334), .ZN(n8758) );
  INV_X1 U23355 ( .I(n14111), .ZN(n16835) );
  INV_X1 U2427 ( .I(n29279), .ZN(n717) );
  INV_X2 U91 ( .I(n25561), .ZN(n15880) );
  INV_X1 U4064 ( .I(n25885), .ZN(n884) );
  INV_X1 U9001 ( .I(n25760), .ZN(n1080) );
  NAND2_X1 U14842 ( .A1(n25013), .A2(n14020), .ZN(n4814) );
  OAI21_X1 U8487 ( .A1(n1221), .A2(n7689), .B(n25892), .ZN(n29594) );
  NAND2_X1 U13398 ( .A1(n27651), .A2(n25019), .ZN(n9402) );
  NOR2_X1 U2010 ( .A1(n25636), .A2(n25713), .ZN(n25639) );
  NOR2_X1 U109 ( .A1(n7413), .A2(n25900), .ZN(n10550) );
  OAI21_X1 U15038 ( .A1(n16528), .A2(n25412), .B(n419), .ZN(n28279) );
  NAND3_X1 U11003 ( .A1(n4968), .A2(n4967), .A3(n18264), .ZN(n29846) );
  NOR2_X1 U2004 ( .A1(n16850), .A2(n16957), .ZN(n26873) );
  NAND2_X1 U16046 ( .A1(n25398), .A2(n25397), .ZN(n25399) );
  OAI21_X1 U3747 ( .A1(n25900), .A2(n16835), .B(n790), .ZN(n15672) );
  NAND2_X1 U16628 ( .A1(n25205), .A2(n27376), .ZN(n27332) );
  NOR2_X1 U4733 ( .A1(n9127), .A2(n16113), .ZN(n11022) );
  INV_X1 U15520 ( .I(n5050), .ZN(n7317) );
  NOR2_X1 U20084 ( .A1(n31268), .A2(n25977), .ZN(n10314) );
  NAND2_X1 U15439 ( .A1(n17987), .A2(n25145), .ZN(n25184) );
  INV_X1 U162 ( .I(n32760), .ZN(n24873) );
  NAND2_X1 U10450 ( .A1(n3013), .A2(n28815), .ZN(n24877) );
  NAND2_X1 U23913 ( .A1(n11716), .A2(n4993), .ZN(n24310) );
  NAND2_X1 U26494 ( .A1(n25133), .A2(n31779), .ZN(n31778) );
  NOR2_X1 U20372 ( .A1(n17839), .A2(n30907), .ZN(n5115) );
  NOR2_X1 U3301 ( .A1(n25620), .A2(n25708), .ZN(n15354) );
  NOR2_X1 U2290 ( .A1(n13464), .A2(n9862), .ZN(n12522) );
  INV_X1 U25606 ( .I(n25339), .ZN(n25337) );
  NAND2_X1 U3293 ( .A1(n15255), .A2(n31945), .ZN(n25531) );
  INV_X1 U4433 ( .I(n6939), .ZN(n1082) );
  INV_X1 U10875 ( .I(n7350), .ZN(n6850) );
  INV_X1 U6999 ( .I(n12247), .ZN(n11106) );
  INV_X1 U7729 ( .I(n25587), .ZN(n25388) );
  INV_X1 U7022 ( .I(n25229), .ZN(n1215) );
  NOR2_X1 U25885 ( .A1(n25562), .A2(n16783), .ZN(n28866) );
  NOR2_X1 U2371 ( .A1(n15964), .A2(n25531), .ZN(n24633) );
  NOR2_X1 U10436 ( .A1(n15646), .A2(n27314), .ZN(n2999) );
  NAND3_X1 U78 ( .A1(n29976), .A2(n25183), .A3(n1218), .ZN(n14632) );
  NAND2_X1 U13514 ( .A1(n16609), .A2(n755), .ZN(n24430) );
  OAI21_X1 U2852 ( .A1(n25199), .A2(n1786), .B(n16632), .ZN(n27990) );
  NOR2_X1 U11238 ( .A1(n5791), .A2(n5793), .ZN(n5570) );
  NAND2_X1 U20208 ( .A1(n5387), .A2(n13349), .ZN(n4232) );
  NAND2_X1 U4016 ( .A1(n28564), .A2(n28562), .ZN(n15883) );
  AOI21_X1 U10297 ( .A1(n146), .A2(n9363), .B(n7064), .ZN(n25767) );
  NAND2_X1 U2333 ( .A1(n25396), .A2(n11556), .ZN(n25439) );
  NAND2_X1 U114 ( .A1(n15550), .A2(n4318), .ZN(n2182) );
  NOR2_X1 U75 ( .A1(n689), .A2(n15013), .ZN(n14539) );
  NOR2_X1 U13045 ( .A1(n15785), .A2(n26873), .ZN(n15783) );
  NOR2_X1 U4386 ( .A1(n10550), .A2(n8470), .ZN(n10547) );
  OAI22_X1 U2745 ( .A1(n2456), .A2(n25234), .B1(n25235), .B2(n25187), .ZN(
        n24570) );
  NAND2_X1 U17416 ( .A1(n25523), .A2(n25522), .ZN(n8442) );
  OAI21_X1 U67 ( .A1(n25896), .A2(n16113), .B(n13349), .ZN(n24708) );
  NAND3_X1 U15626 ( .A1(n17673), .A2(n14247), .A3(n25404), .ZN(n25441) );
  AOI21_X1 U9087 ( .A1(n11306), .A2(n25633), .B(n27637), .ZN(n12000) );
  OAI21_X1 U10381 ( .A1(n12025), .A2(n17367), .B(n25388), .ZN(n11823) );
  AOI21_X1 U23903 ( .A1(n24604), .A2(n15719), .B(n27314), .ZN(n17379) );
  OAI22_X1 U6028 ( .A1(n8186), .A2(n11944), .B1(n17092), .B2(n6939), .ZN(
        n15276) );
  NOR2_X1 U10372 ( .A1(n4095), .A2(n7041), .ZN(n11698) );
  NAND2_X1 U10428 ( .A1(n12058), .A2(n16752), .ZN(n11347) );
  AOI21_X1 U2719 ( .A1(n14484), .A2(n32761), .B(n11082), .ZN(n11429) );
  NAND2_X1 U12511 ( .A1(n1620), .A2(n25887), .ZN(n25914) );
  INV_X1 U7030 ( .I(n2270), .ZN(n15061) );
  INV_X1 U8008 ( .I(n10174), .ZN(n10504) );
  INV_X1 U15219 ( .I(n25376), .ZN(n25352) );
  INV_X2 U9998 ( .I(n1597), .ZN(n25738) );
  NAND2_X1 U14917 ( .A1(n25107), .A2(n11360), .ZN(n7862) );
  INV_X1 U4928 ( .I(n25478), .ZN(n25487) );
  CLKBUF_X2 U2934 ( .I(n7702), .Z(n7701) );
  INV_X1 U14791 ( .I(n25795), .ZN(n16111) );
  NAND2_X1 U57 ( .A1(n16494), .A2(n13640), .ZN(n13124) );
  INV_X2 U17512 ( .I(n16380), .ZN(n1951) );
  INV_X1 U1540 ( .I(n25154), .ZN(n25179) );
  INV_X1 U10377 ( .I(n25369), .ZN(n25367) );
  INV_X1 U24431 ( .I(n14915), .ZN(n25834) );
  OAI21_X1 U8903 ( .A1(n3489), .A2(n2536), .B(n32059), .ZN(n8951) );
  NOR2_X1 U1905 ( .A1(n30279), .A2(n25002), .ZN(n15078) );
  NAND2_X1 U15859 ( .A1(n25687), .A2(n25686), .ZN(n2016) );
  NOR2_X1 U7032 ( .A1(n5411), .A2(n7701), .ZN(n14434) );
  INV_X1 U23575 ( .I(n31360), .ZN(n25552) );
  NOR2_X1 U13124 ( .A1(n14199), .A2(n25863), .ZN(n13952) );
  NAND2_X1 U15732 ( .A1(n8202), .A2(n4525), .ZN(n4524) );
  INV_X1 U21482 ( .I(n25464), .ZN(n17200) );
  CLKBUF_X1 U4329 ( .I(n25557), .Z(n31647) );
  NAND2_X1 U25689 ( .A1(n29116), .A2(n25476), .ZN(n25474) );
  INV_X1 U10322 ( .I(n25738), .ZN(n25748) );
  INV_X1 U5548 ( .I(n25863), .ZN(n25854) );
  INV_X1 U19 ( .I(n24915), .ZN(n6154) );
  INV_X1 U7051 ( .I(n25724), .ZN(n25729) );
  INV_X1 U3985 ( .I(n13483), .ZN(n14944) );
  NAND4_X1 U4 ( .A1(n25914), .A2(n25922), .A3(n11019), .A4(n25913), .ZN(n25918) );
  NAND2_X1 U10329 ( .A1(n24351), .A2(n24927), .ZN(n24349) );
  NAND3_X1 U3 ( .A1(n25318), .A2(n17058), .A3(n17105), .ZN(n27063) );
  NOR2_X1 U7 ( .A1(n8639), .A2(n32398), .ZN(n32270) );
  INV_X1 U16 ( .I(n13960), .ZN(n25925) );
  INV_X1 U17 ( .I(n25106), .ZN(n32857) );
  BUF_X2 U18 ( .I(n25820), .Z(n11003) );
  NOR2_X1 U20 ( .A1(n16112), .A2(n12611), .ZN(n12395) );
  NOR2_X1 U21 ( .A1(n25788), .A2(n25796), .ZN(n25775) );
  NAND2_X1 U22 ( .A1(n7586), .A2(n11360), .ZN(n25093) );
  NAND2_X1 U25 ( .A1(n24925), .A2(n15799), .ZN(n24928) );
  NAND2_X1 U26 ( .A1(n34109), .A2(n25247), .ZN(n7924) );
  AND2_X1 U27 ( .A1(n25387), .A2(n33876), .Z(n32869) );
  INV_X1 U28 ( .I(n15323), .ZN(n712) );
  BUF_X2 U29 ( .I(n5578), .Z(n5043) );
  INV_X1 U30 ( .I(n24910), .ZN(n24902) );
  AOI21_X1 U31 ( .A1(n5810), .A2(n8186), .B(n32992), .ZN(n25731) );
  CLKBUF_X2 U32 ( .I(n25285), .Z(n28532) );
  INV_X1 U33 ( .I(n6595), .ZN(n33399) );
  INV_X1 U37 ( .I(n24955), .ZN(n1201) );
  INV_X1 U38 ( .I(n25820), .ZN(n17642) );
  NAND2_X1 U40 ( .A1(n32882), .A2(n10609), .ZN(n33900) );
  NOR2_X1 U42 ( .A1(n25818), .A2(n4450), .ZN(n9182) );
  OAI21_X2 U51 ( .A1(n32471), .A2(n32565), .B(n25010), .ZN(n25062) );
  OR2_X1 U55 ( .A1(n24572), .A2(n24570), .Z(n32882) );
  INV_X1 U56 ( .I(n24995), .ZN(n5072) );
  NAND2_X1 U59 ( .A1(n33632), .A2(n12968), .ZN(n25845) );
  NOR2_X1 U60 ( .A1(n32030), .A2(n14872), .ZN(n32311) );
  NAND3_X1 U61 ( .A1(n15051), .A2(n5659), .A3(n5755), .ZN(n30928) );
  AOI21_X1 U65 ( .A1(n25564), .A2(n3405), .B(n25582), .ZN(n32585) );
  NAND2_X1 U66 ( .A1(n32570), .A2(n5292), .ZN(n32135) );
  AND2_X1 U70 ( .A1(n13985), .A2(n25306), .Z(n32020) );
  NOR2_X1 U72 ( .A1(n33074), .A2(n16566), .ZN(n32626) );
  NAND3_X1 U73 ( .A1(n27119), .A2(n16339), .A3(n25412), .ZN(n33245) );
  NAND2_X1 U76 ( .A1(n33599), .A2(n33598), .ZN(n33632) );
  CLKBUF_X2 U77 ( .I(n7532), .Z(n31946) );
  NAND2_X1 U81 ( .A1(n6851), .A2(n12440), .ZN(n2000) );
  NAND2_X1 U82 ( .A1(n32828), .A2(n32761), .ZN(n8776) );
  NAND2_X1 U83 ( .A1(n11703), .A2(n25347), .ZN(n30930) );
  OAI21_X1 U85 ( .A1(n30372), .A2(n25329), .B(n28958), .ZN(n33880) );
  OAI21_X1 U86 ( .A1(n14991), .A2(n12093), .B(n30461), .ZN(n32205) );
  OAI21_X1 U87 ( .A1(n15555), .A2(n25893), .B(n9127), .ZN(n11020) );
  AOI21_X1 U89 ( .A1(n25711), .A2(n24729), .B(n4407), .ZN(n27208) );
  NOR2_X1 U92 ( .A1(n16783), .A2(n25561), .ZN(n30983) );
  NOR2_X1 U93 ( .A1(n1221), .A2(n547), .ZN(n12160) );
  NAND2_X1 U95 ( .A1(n25755), .A2(n28338), .ZN(n25876) );
  OR2_X1 U97 ( .A1(n28242), .A2(n25627), .Z(n32032) );
  AND2_X1 U98 ( .A1(n17240), .A2(n25012), .Z(n11977) );
  CLKBUF_X2 U99 ( .I(n25582), .Z(n27947) );
  NAND2_X1 U102 ( .A1(n28110), .A2(n1211), .ZN(n33002) );
  NOR2_X1 U104 ( .A1(n765), .A2(n25331), .ZN(n30522) );
  AND2_X1 U108 ( .A1(n9195), .A2(n25700), .Z(n32028) );
  OR2_X1 U110 ( .A1(n317), .A2(n16783), .Z(n32029) );
  INV_X1 U113 ( .I(n32878), .ZN(n32761) );
  AND2_X1 U116 ( .A1(n17240), .A2(n25014), .Z(n14991) );
  OR2_X1 U120 ( .A1(n24667), .A2(n16957), .Z(n33962) );
  INV_X1 U125 ( .I(n33067), .ZN(n33066) );
  NAND2_X1 U126 ( .A1(n16276), .A2(n25183), .ZN(n14630) );
  NAND2_X1 U140 ( .A1(n16751), .A2(n17987), .ZN(n14629) );
  NOR2_X1 U142 ( .A1(n1567), .A2(n25121), .ZN(n7771) );
  NAND2_X1 U144 ( .A1(n25891), .A2(n25890), .ZN(n30811) );
  INV_X2 U146 ( .I(n11045), .ZN(n25902) );
  BUF_X2 U148 ( .I(n25883), .Z(n15152) );
  INV_X2 U149 ( .I(n25409), .ZN(n752) );
  NOR2_X1 U154 ( .A1(n28338), .A2(n25755), .ZN(n28110) );
  NAND2_X1 U157 ( .A1(n25014), .A2(n11974), .ZN(n24977) );
  OR2_X1 U160 ( .A1(n10569), .A2(n4951), .Z(n25289) );
  INV_X1 U161 ( .I(n31945), .ZN(n16648) );
  AOI21_X1 U165 ( .A1(n15459), .A2(n25697), .B(n751), .ZN(n15458) );
  BUF_X2 U169 ( .I(n25238), .Z(n28136) );
  CLKBUF_X2 U172 ( .I(n17382), .Z(n27314) );
  CLKBUF_X1 U174 ( .I(n25334), .Z(n33460) );
  CLKBUF_X1 U177 ( .I(n16510), .Z(n32884) );
  AOI21_X1 U178 ( .A1(n31149), .A2(n16704), .B(n25561), .ZN(n33067) );
  BUF_X2 U179 ( .I(n25563), .Z(n317) );
  CLKBUF_X2 U180 ( .I(n24436), .Z(n33120) );
  OR2_X1 U183 ( .A1(n6725), .A2(n27181), .Z(n25584) );
  NAND2_X1 U185 ( .A1(n25295), .A2(n16650), .ZN(n25343) );
  INV_X1 U187 ( .I(n10569), .ZN(n5468) );
  BUF_X2 U191 ( .I(n25022), .Z(n25121) );
  BUF_X2 U199 ( .I(n14246), .Z(n33919) );
  INV_X1 U202 ( .I(n24692), .ZN(n14110) );
  INV_X1 U215 ( .I(n24547), .ZN(n32575) );
  BUF_X2 U216 ( .I(n3253), .Z(n30069) );
  INV_X1 U217 ( .I(n27115), .ZN(n32346) );
  OAI22_X1 U219 ( .A1(n17581), .A2(n3219), .B1(n15086), .B2(n15085), .ZN(
        n32871) );
  AOI21_X1 U221 ( .A1(n32470), .A2(n28827), .B(n25974), .ZN(n13217) );
  NAND2_X1 U222 ( .A1(n891), .A2(n33935), .ZN(n27397) );
  NAND2_X1 U228 ( .A1(n33123), .A2(n6978), .ZN(n6167) );
  NAND3_X1 U229 ( .A1(n16651), .A2(n30061), .A3(n29977), .ZN(n7729) );
  AOI22_X1 U233 ( .A1(n2853), .A2(n24163), .B1(n24002), .B2(n16552), .ZN(n2848) );
  OAI21_X1 U234 ( .A1(n13659), .A2(n29473), .B(n9219), .ZN(n29605) );
  AOI21_X1 U238 ( .A1(n24268), .A2(n11768), .B(n12644), .ZN(n11767) );
  OAI22_X1 U239 ( .A1(n24235), .A2(n24237), .B1(n11883), .B2(n24234), .ZN(
        n24239) );
  AOI21_X1 U242 ( .A1(n7150), .A2(n15179), .B(n9889), .ZN(n12341) );
  INV_X1 U243 ( .I(n32444), .ZN(n13659) );
  NAND2_X1 U244 ( .A1(n24052), .A2(n14123), .ZN(n24125) );
  NAND2_X1 U247 ( .A1(n14386), .A2(n7962), .ZN(n33951) );
  NAND2_X1 U249 ( .A1(n5132), .A2(n32228), .ZN(n5130) );
  NAND3_X1 U252 ( .A1(n890), .A2(n29141), .A3(n7361), .ZN(n7360) );
  OR2_X1 U255 ( .A1(n29634), .A2(n12374), .Z(n12054) );
  CLKBUF_X1 U256 ( .I(n10987), .Z(n28538) );
  OAI21_X1 U257 ( .A1(n32552), .A2(n32551), .B(n24213), .ZN(n24007) );
  NAND2_X1 U260 ( .A1(n10687), .A2(n13), .ZN(n13974) );
  NAND2_X1 U263 ( .A1(n24337), .A2(n33680), .ZN(n1998) );
  NOR2_X1 U266 ( .A1(n28300), .A2(n31985), .ZN(n6105) );
  NAND2_X1 U269 ( .A1(n24318), .A2(n2913), .ZN(n26488) );
  AOI21_X1 U270 ( .A1(n9946), .A2(n27931), .B(n4019), .ZN(n5708) );
  NAND2_X1 U272 ( .A1(n31377), .A2(n24317), .ZN(n32166) );
  NAND2_X1 U275 ( .A1(n24143), .A2(n27430), .ZN(n33653) );
  NOR2_X1 U280 ( .A1(n31355), .A2(n28694), .ZN(n33872) );
  OR2_X1 U286 ( .A1(n24141), .A2(n24084), .Z(n16017) );
  AOI22_X1 U293 ( .A1(n32062), .A2(n27739), .B1(n24133), .B2(n23714), .ZN(
        n2939) );
  NAND3_X1 U296 ( .A1(n32298), .A2(n14112), .A3(n2913), .ZN(n33912) );
  AOI21_X1 U298 ( .A1(n28410), .A2(n5308), .B(n3506), .ZN(n28409) );
  NAND3_X1 U300 ( .A1(n9066), .A2(n12982), .A3(n27739), .ZN(n16950) );
  NAND2_X1 U305 ( .A1(n24161), .A2(n24123), .ZN(n5969) );
  NAND2_X1 U306 ( .A1(n31342), .A2(n24249), .ZN(n32470) );
  INV_X2 U307 ( .I(n15179), .ZN(n15876) );
  NAND2_X1 U310 ( .A1(n24340), .A2(n24056), .ZN(n4049) );
  NOR2_X1 U314 ( .A1(n24309), .A2(n3421), .ZN(n24135) );
  INV_X1 U315 ( .I(n24248), .ZN(n31342) );
  INV_X2 U321 ( .I(n12143), .ZN(n33444) );
  BUF_X2 U331 ( .I(n24164), .Z(n2847) );
  NAND3_X1 U333 ( .A1(n13984), .A2(n5913), .A3(n31096), .ZN(n11743) );
  AND2_X1 U334 ( .A1(n2539), .A2(n11503), .Z(n31985) );
  NAND2_X1 U336 ( .A1(n31497), .A2(n10530), .ZN(n2529) );
  OR2_X1 U337 ( .A1(n24254), .A2(n33532), .Z(n7149) );
  INV_X1 U338 ( .I(n27430), .ZN(n33655) );
  NOR2_X1 U341 ( .A1(n24209), .A2(n24212), .ZN(n32551) );
  NAND2_X1 U343 ( .A1(n12644), .A2(n3148), .ZN(n4961) );
  NOR2_X1 U344 ( .A1(n24347), .A2(n3165), .ZN(n30121) );
  NAND2_X1 U346 ( .A1(n13334), .A2(n6713), .ZN(n1500) );
  INV_X2 U347 ( .I(n26120), .ZN(n2640) );
  INV_X1 U349 ( .I(n24053), .ZN(n24185) );
  INV_X2 U350 ( .I(n2826), .ZN(n24340) );
  BUF_X2 U351 ( .I(n6555), .Z(n6581) );
  OAI21_X1 U354 ( .A1(n24225), .A2(n10687), .B(n24223), .ZN(n32677) );
  NAND2_X1 U358 ( .A1(n7991), .A2(n26415), .ZN(n23997) );
  NAND2_X1 U362 ( .A1(n4024), .A2(n24312), .ZN(n29051) );
  INV_X1 U364 ( .I(n15720), .ZN(n14703) );
  NAND3_X1 U365 ( .A1(n15943), .A2(n23903), .A3(n15942), .ZN(n29575) );
  OAI21_X1 U367 ( .A1(n28688), .A2(n2233), .B(n23544), .ZN(n29052) );
  AOI22_X1 U368 ( .A1(n9768), .A2(n9797), .B1(n23787), .B2(n9769), .ZN(n32442)
         );
  AND2_X1 U378 ( .A1(n23867), .A2(n17895), .Z(n12090) );
  OAI21_X1 U379 ( .A1(n9736), .A2(n976), .B(n4408), .ZN(n6041) );
  NOR2_X1 U380 ( .A1(n29198), .A2(n33659), .ZN(n33055) );
  NOR2_X1 U381 ( .A1(n25987), .A2(n23575), .ZN(n27329) );
  NOR3_X1 U384 ( .A1(n2752), .A2(n23806), .A3(n28273), .ZN(n9899) );
  NOR2_X1 U385 ( .A1(n33828), .A2(n33827), .ZN(n4374) );
  NOR3_X1 U387 ( .A1(n32210), .A2(n7444), .A3(n32209), .ZN(n31084) );
  OAI21_X1 U392 ( .A1(n12070), .A2(n32522), .B(n23897), .ZN(n18117) );
  NAND3_X1 U396 ( .A1(n8835), .A2(n31560), .A3(n23600), .ZN(n6932) );
  OAI21_X1 U397 ( .A1(n30621), .A2(n30620), .B(n23878), .ZN(n33370) );
  AOI21_X1 U401 ( .A1(n30991), .A2(n23824), .B(n27893), .ZN(n24188) );
  NAND2_X1 U402 ( .A1(n28016), .A2(n32209), .ZN(n33043) );
  NAND2_X1 U405 ( .A1(n33340), .A2(n3371), .ZN(n32128) );
  NAND2_X1 U416 ( .A1(n33005), .A2(n23576), .ZN(n30803) );
  NOR2_X1 U418 ( .A1(n11904), .A2(n23860), .ZN(n12592) );
  NOR3_X1 U419 ( .A1(n6662), .A2(n23756), .A3(n23760), .ZN(n13903) );
  OAI21_X1 U422 ( .A1(n6661), .A2(n15600), .B(n17691), .ZN(n32607) );
  NAND2_X1 U423 ( .A1(n32986), .A2(n1920), .ZN(n7777) );
  AOI22_X1 U427 ( .A1(n15451), .A2(n33110), .B1(n2561), .B2(n2560), .ZN(n33071) );
  OAI21_X1 U431 ( .A1(n23634), .A2(n23633), .B(n11240), .ZN(n5227) );
  AOI22_X1 U432 ( .A1(n16224), .A2(n23754), .B1(n28297), .B2(n23726), .ZN(
        n33313) );
  OR2_X1 U433 ( .A1(n4281), .A2(n707), .Z(n31982) );
  INV_X1 U434 ( .I(n33867), .ZN(n32425) );
  AND2_X1 U435 ( .A1(n8270), .A2(n843), .Z(n10143) );
  INV_X1 U436 ( .I(n16320), .ZN(n23697) );
  CLKBUF_X2 U437 ( .I(n23588), .Z(n33103) );
  NOR2_X1 U443 ( .A1(n6414), .A2(n14975), .ZN(n32801) );
  INV_X1 U444 ( .I(n14335), .ZN(n23812) );
  NOR2_X1 U450 ( .A1(n756), .A2(n29272), .ZN(n10384) );
  AND2_X1 U454 ( .A1(n14975), .A2(n14974), .Z(n31981) );
  NOR2_X1 U459 ( .A1(n4069), .A2(n34009), .ZN(n32522) );
  NOR2_X1 U460 ( .A1(n32610), .A2(n11923), .ZN(n32609) );
  NAND2_X1 U467 ( .A1(n17777), .A2(n980), .ZN(n31759) );
  OAI21_X1 U472 ( .A1(n27678), .A2(n1257), .B(n32547), .ZN(n11654) );
  NOR2_X1 U474 ( .A1(n23897), .A2(n4069), .ZN(n33096) );
  NOR2_X1 U475 ( .A1(n32434), .A2(n32657), .ZN(n7262) );
  NAND2_X1 U478 ( .A1(n846), .A2(n13549), .ZN(n33340) );
  NAND2_X1 U481 ( .A1(n33670), .A2(n651), .ZN(n23881) );
  NOR2_X1 U486 ( .A1(n23775), .A2(n31810), .ZN(n17750) );
  NAND3_X1 U494 ( .A1(n26775), .A2(n16677), .A3(n17373), .ZN(n32354) );
  NAND2_X1 U495 ( .A1(n6247), .A2(n17726), .ZN(n8836) );
  OAI22_X1 U500 ( .A1(n8093), .A2(n33831), .B1(n23583), .B2(n27910), .ZN(
        n33018) );
  NOR2_X1 U501 ( .A1(n13905), .A2(n13413), .ZN(n15600) );
  NAND2_X1 U505 ( .A1(n23590), .A2(n6661), .ZN(n17691) );
  OR2_X1 U507 ( .A1(n23871), .A2(n6474), .Z(n32004) );
  BUF_X2 U509 ( .I(n11923), .Z(n33337) );
  INV_X1 U510 ( .I(n8838), .ZN(n6247) );
  INV_X1 U513 ( .I(n32999), .ZN(n2561) );
  NAND2_X1 U518 ( .A1(n10279), .A2(n9375), .ZN(n23882) );
  NAND2_X1 U522 ( .A1(n33354), .A2(n32711), .ZN(n5627) );
  CLKBUF_X2 U525 ( .I(n5736), .Z(n33260) );
  CLKBUF_X2 U526 ( .I(n15865), .Z(n14325) );
  INV_X1 U527 ( .I(n29472), .ZN(n23824) );
  BUF_X1 U530 ( .I(n9939), .Z(n33499) );
  INV_X2 U531 ( .I(n13998), .ZN(n33789) );
  NOR2_X1 U533 ( .A1(n14133), .A2(n32170), .ZN(n23825) );
  NAND2_X1 U536 ( .A1(n34036), .A2(n23767), .ZN(n1610) );
  NAND2_X1 U538 ( .A1(n13905), .A2(n26115), .ZN(n16292) );
  BUF_X2 U544 ( .I(n23156), .Z(n18204) );
  BUF_X2 U548 ( .I(n12974), .Z(n12658) );
  CLKBUF_X2 U555 ( .I(n17857), .Z(n25996) );
  CLKBUF_X2 U563 ( .I(n17812), .Z(n3760) );
  NAND2_X1 U567 ( .A1(n23867), .A2(n657), .ZN(n10140) );
  BUF_X2 U573 ( .I(n23202), .Z(n29217) );
  INV_X1 U574 ( .I(n23363), .ZN(n8915) );
  INV_X1 U575 ( .I(n23496), .ZN(n33111) );
  INV_X1 U576 ( .I(n23202), .ZN(n10625) );
  INV_X1 U579 ( .I(n11504), .ZN(n32214) );
  NAND2_X1 U581 ( .A1(n1565), .A2(n1564), .ZN(n27148) );
  NAND2_X1 U587 ( .A1(n11741), .A2(n11740), .ZN(n60) );
  NAND2_X1 U591 ( .A1(n32513), .A2(n22863), .ZN(n13918) );
  NAND2_X1 U593 ( .A1(n33640), .A2(n5182), .ZN(n33556) );
  OAI21_X1 U595 ( .A1(n22838), .A2(n33596), .B(n32827), .ZN(n4871) );
  NOR2_X1 U601 ( .A1(n6350), .A2(n29648), .ZN(n32324) );
  AND2_X1 U602 ( .A1(n5274), .A2(n10295), .Z(n11538) );
  NAND2_X1 U603 ( .A1(n2114), .A2(n8990), .ZN(n2113) );
  NOR2_X1 U604 ( .A1(n28689), .A2(n11059), .ZN(n32513) );
  NAND2_X1 U609 ( .A1(n29115), .A2(n17399), .ZN(n4649) );
  AOI22_X1 U611 ( .A1(n29329), .A2(n32935), .B1(n6433), .B2(n27814), .ZN(
        n22721) );
  CLKBUF_X2 U612 ( .I(n1266), .Z(n26373) );
  NAND2_X1 U614 ( .A1(n4845), .A2(n28974), .ZN(n4846) );
  OAI21_X1 U617 ( .A1(n27212), .A2(n31936), .B(n9293), .ZN(n16879) );
  NAND2_X1 U621 ( .A1(n32960), .A2(n32959), .ZN(n29401) );
  OAI21_X1 U623 ( .A1(n16975), .A2(n29391), .B(n23026), .ZN(n8853) );
  NAND2_X1 U624 ( .A1(n27798), .A2(n15349), .ZN(n33346) );
  NAND2_X1 U643 ( .A1(n23090), .A2(n33968), .ZN(n33932) );
  AOI21_X1 U644 ( .A1(n22720), .A2(n31531), .B(n32935), .ZN(n27775) );
  NAND2_X1 U645 ( .A1(n2712), .A2(n23106), .ZN(n32827) );
  OAI21_X1 U648 ( .A1(n11317), .A2(n33563), .B(n33562), .ZN(n22881) );
  INV_X1 U649 ( .I(n34017), .ZN(n29427) );
  OAI21_X1 U652 ( .A1(n33022), .A2(n30976), .B(n32258), .ZN(n22770) );
  NOR2_X1 U653 ( .A1(n12181), .A2(n15317), .ZN(n33510) );
  AOI21_X1 U654 ( .A1(n32307), .A2(n23079), .B(n6985), .ZN(n32318) );
  NAND2_X1 U665 ( .A1(n22769), .A2(n28415), .ZN(n32580) );
  OAI21_X1 U669 ( .A1(n4208), .A2(n23093), .B(n776), .ZN(n32964) );
  CLKBUF_X4 U671 ( .I(n23087), .Z(n6236) );
  NAND2_X1 U677 ( .A1(n6149), .A2(n22473), .ZN(n12418) );
  NOR2_X1 U681 ( .A1(n22832), .A2(n23000), .ZN(n22753) );
  AND2_X1 U682 ( .A1(n6835), .A2(n6836), .Z(n32868) );
  INV_X1 U686 ( .I(n22592), .ZN(n22900) );
  NOR2_X1 U688 ( .A1(n899), .A2(n30976), .ZN(n32959) );
  NAND2_X1 U691 ( .A1(n15935), .A2(n7047), .ZN(n23479) );
  CLKBUF_X2 U692 ( .I(n22848), .Z(n3184) );
  NOR2_X1 U701 ( .A1(n30909), .A2(n28313), .ZN(n15915) );
  NAND2_X1 U702 ( .A1(n14183), .A2(n5915), .ZN(n27296) );
  NAND2_X1 U705 ( .A1(n22792), .A2(n27090), .ZN(n32560) );
  NAND3_X1 U706 ( .A1(n15389), .A2(n27090), .A3(n4113), .ZN(n28178) );
  AOI21_X1 U707 ( .A1(n11495), .A2(n32820), .B(n1106), .ZN(n33179) );
  NOR2_X1 U711 ( .A1(n32842), .A2(n34017), .ZN(n15362) );
  INV_X1 U713 ( .I(n5682), .ZN(n30825) );
  NAND2_X1 U714 ( .A1(n22894), .A2(n30909), .ZN(n15190) );
  NOR2_X1 U720 ( .A1(n12586), .A2(n28697), .ZN(n22835) );
  AOI21_X1 U721 ( .A1(n23055), .A2(n3007), .B(n29107), .ZN(n14417) );
  NOR2_X1 U722 ( .A1(n32500), .A2(n23056), .ZN(n32424) );
  NAND3_X1 U726 ( .A1(n7181), .A2(n898), .A3(n4734), .ZN(n26312) );
  NAND2_X1 U727 ( .A1(n26526), .A2(n33132), .ZN(n22709) );
  INV_X1 U729 ( .I(n22832), .ZN(n79) );
  INV_X1 U731 ( .I(n22960), .ZN(n23082) );
  AND2_X1 U737 ( .A1(n9963), .A2(n30868), .Z(n32092) );
  INV_X1 U740 ( .I(n15456), .ZN(n12727) );
  INV_X2 U742 ( .I(n5274), .ZN(n11317) );
  AND2_X1 U745 ( .A1(n10528), .A2(n6975), .Z(n8022) );
  CLKBUF_X2 U746 ( .I(n27419), .Z(n32119) );
  INV_X2 U749 ( .I(n22795), .ZN(n23042) );
  INV_X2 U750 ( .I(n22798), .ZN(n772) );
  INV_X1 U753 ( .I(n22957), .ZN(n9778) );
  NOR2_X1 U756 ( .A1(n4580), .A2(n16486), .ZN(n13648) );
  CLKBUF_X2 U757 ( .I(n30293), .Z(n27798) );
  INV_X2 U758 ( .I(n31325), .ZN(n17211) );
  BUF_X2 U763 ( .I(n13762), .Z(n6800) );
  BUF_X2 U764 ( .I(n6605), .Z(n30909) );
  NOR2_X1 U765 ( .A1(n22885), .A2(n1577), .ZN(n22815) );
  INV_X1 U766 ( .I(n6799), .ZN(n22950) );
  INV_X2 U772 ( .I(n30297), .ZN(n1278) );
  NAND3_X1 U779 ( .A1(n32192), .A2(n32191), .A3(n5769), .ZN(n5573) );
  NAND2_X1 U781 ( .A1(n22530), .A2(n22531), .ZN(n12256) );
  AND2_X1 U784 ( .A1(n22442), .A2(n28692), .Z(n31934) );
  NAND2_X1 U785 ( .A1(n9425), .A2(n22539), .ZN(n4502) );
  NOR3_X1 U787 ( .A1(n5597), .A2(n22534), .A3(n16434), .ZN(n4503) );
  AOI22_X1 U794 ( .A1(n30065), .A2(n22570), .B1(n1297), .B2(n18073), .ZN(
        n33855) );
  NAND2_X1 U798 ( .A1(n32194), .A2(n32193), .ZN(n32192) );
  OAI21_X1 U801 ( .A1(n33061), .A2(n22407), .B(n32448), .ZN(n29982) );
  NAND2_X1 U805 ( .A1(n22530), .A2(n15643), .ZN(n6505) );
  INV_X1 U809 ( .I(n22612), .ZN(n32757) );
  AOI21_X1 U811 ( .A1(n22671), .A2(n29371), .B(n26098), .ZN(n33262) );
  NAND2_X1 U814 ( .A1(n2066), .A2(n22487), .ZN(n32680) );
  NOR2_X1 U817 ( .A1(n29078), .A2(n11917), .ZN(n33502) );
  AOI21_X1 U823 ( .A1(n11874), .A2(n16556), .B(n16570), .ZN(n33974) );
  OAI22_X1 U831 ( .A1(n14137), .A2(n5743), .B1(n22658), .B2(n22659), .ZN(
        n22366) );
  AOI21_X1 U838 ( .A1(n27959), .A2(n2418), .B(n11250), .ZN(n33463) );
  AND2_X1 U840 ( .A1(n22476), .A2(n22394), .Z(n15103) );
  INV_X1 U842 ( .I(n33227), .ZN(n3596) );
  NAND2_X1 U851 ( .A1(n12899), .A2(n22586), .ZN(n9452) );
  NAND2_X1 U856 ( .A1(n29261), .A2(n11920), .ZN(n21963) );
  NOR2_X1 U858 ( .A1(n34035), .A2(n5597), .ZN(n33061) );
  INV_X1 U861 ( .I(n15746), .ZN(n32193) );
  AOI21_X1 U864 ( .A1(n18038), .A2(n22427), .B(n28170), .ZN(n32446) );
  OR2_X1 U868 ( .A1(n22476), .A2(n29101), .Z(n12072) );
  OR2_X1 U870 ( .A1(n22474), .A2(n22476), .Z(n17247) );
  INV_X2 U872 ( .I(n29508), .ZN(n33455) );
  NOR2_X1 U881 ( .A1(n29078), .A2(n908), .ZN(n32823) );
  NOR3_X1 U883 ( .A1(n22636), .A2(n22640), .A3(n12043), .ZN(n22731) );
  NAND3_X1 U902 ( .A1(n16529), .A2(n22926), .A3(n22658), .ZN(n33368) );
  OAI21_X1 U905 ( .A1(n30334), .A2(n29461), .B(n30065), .ZN(n33982) );
  NOR2_X1 U906 ( .A1(n14728), .A2(n16375), .ZN(n12335) );
  INV_X1 U909 ( .I(n6976), .ZN(n22343) );
  BUF_X2 U910 ( .I(n6976), .Z(n239) );
  INV_X1 U913 ( .I(n26884), .ZN(n32831) );
  INV_X1 U936 ( .I(n29288), .ZN(n22558) );
  INV_X2 U948 ( .I(n22476), .ZN(n22377) );
  NAND2_X1 U952 ( .A1(n2858), .A2(n5961), .ZN(n7848) );
  INV_X1 U955 ( .I(n14227), .ZN(n32334) );
  NAND2_X1 U956 ( .A1(n22644), .A2(n22645), .ZN(n33026) );
  NAND2_X1 U965 ( .A1(n22330), .A2(n1116), .ZN(n11011) );
  NOR2_X1 U966 ( .A1(n14728), .A2(n12338), .ZN(n27878) );
  NAND3_X1 U968 ( .A1(n6242), .A2(n6244), .A3(n22639), .ZN(n32987) );
  NAND2_X1 U969 ( .A1(n22332), .A2(n28692), .ZN(n22569) );
  NAND2_X1 U971 ( .A1(n14251), .A2(n32830), .ZN(n12840) );
  NAND3_X1 U978 ( .A1(n33628), .A2(n6186), .A3(n6187), .ZN(n33619) );
  INV_X1 U980 ( .I(n9630), .ZN(n33281) );
  INV_X1 U981 ( .I(n22367), .ZN(n31964) );
  AND2_X1 U986 ( .A1(n27933), .A2(n26317), .Z(n22688) );
  CLKBUF_X2 U988 ( .I(n8420), .Z(n327) );
  BUF_X2 U993 ( .I(n9515), .Z(n5743) );
  BUF_X2 U996 ( .I(n22350), .Z(n1294) );
  NOR2_X1 U997 ( .A1(n33320), .A2(n8409), .ZN(n32569) );
  NAND2_X1 U999 ( .A1(n8131), .A2(n12496), .ZN(n9272) );
  INV_X1 U1002 ( .I(n4916), .ZN(n10654) );
  AOI21_X1 U1010 ( .A1(n32797), .A2(n17076), .B(n10354), .ZN(n13070) );
  NOR2_X1 U1012 ( .A1(n998), .A2(n1116), .ZN(n28019) );
  INV_X1 U1019 ( .I(n31692), .ZN(n10183) );
  INV_X1 U1021 ( .I(n5961), .ZN(n5991) );
  INV_X2 U1026 ( .I(n1926), .ZN(n16647) );
  INV_X1 U1028 ( .I(n22157), .ZN(n33593) );
  INV_X1 U1035 ( .I(n8617), .ZN(n22296) );
  BUF_X2 U1039 ( .I(n22160), .Z(n4295) );
  INV_X1 U1049 ( .I(n16237), .ZN(n1307) );
  INV_X1 U1055 ( .I(n22032), .ZN(n32714) );
  INV_X1 U1057 ( .I(n22211), .ZN(n33151) );
  INV_X1 U1062 ( .I(n29137), .ZN(n34063) );
  INV_X1 U1064 ( .I(n22113), .ZN(n31165) );
  INV_X1 U1072 ( .I(n22076), .ZN(n21892) );
  INV_X1 U1075 ( .I(n22283), .ZN(n1129) );
  NAND2_X1 U1076 ( .A1(n11727), .A2(n21964), .ZN(n11359) );
  INV_X1 U1079 ( .I(n22042), .ZN(n34014) );
  INV_X1 U1080 ( .I(n21945), .ZN(n32126) );
  NAND3_X1 U1081 ( .A1(n21933), .A2(n21932), .A3(n28895), .ZN(n6426) );
  NOR2_X1 U1082 ( .A1(n15639), .A2(n33298), .ZN(n10234) );
  NAND3_X1 U1087 ( .A1(n33481), .A2(n6238), .A3(n6237), .ZN(n33471) );
  NAND2_X1 U1089 ( .A1(n5228), .A2(n26671), .ZN(n31657) );
  NAND3_X1 U1090 ( .A1(n28895), .A2(n30440), .A3(n10699), .ZN(n32608) );
  NAND2_X1 U1091 ( .A1(n15465), .A2(n32833), .ZN(n32832) );
  AOI22_X1 U1092 ( .A1(n13248), .A2(n21546), .B1(n17429), .B2(n21730), .ZN(
        n7457) );
  AND2_X1 U1097 ( .A1(n2643), .A2(n21704), .Z(n32071) );
  OAI21_X1 U1099 ( .A1(n31260), .A2(n32384), .B(n8029), .ZN(n27631) );
  NOR2_X1 U1101 ( .A1(n21856), .A2(n13116), .ZN(n2352) );
  AOI22_X1 U1106 ( .A1(n16016), .A2(n276), .B1(n31220), .B2(n21778), .ZN(
        n33676) );
  OAI21_X1 U1108 ( .A1(n14641), .A2(n17078), .B(n32282), .ZN(n9686) );
  INV_X1 U1117 ( .I(n396), .ZN(n32321) );
  OAI21_X1 U1120 ( .A1(n17225), .A2(n17226), .B(n423), .ZN(n8077) );
  OAI21_X1 U1126 ( .A1(n11644), .A2(n29784), .B(n8029), .ZN(n11643) );
  OAI21_X1 U1128 ( .A1(n33520), .A2(n33519), .B(n4331), .ZN(n6766) );
  NOR2_X1 U1129 ( .A1(n14642), .A2(n914), .ZN(n28393) );
  AOI21_X1 U1142 ( .A1(n12626), .A2(n11619), .B(n26474), .ZN(n16192) );
  NOR2_X1 U1146 ( .A1(n915), .A2(n31911), .ZN(n32325) );
  NAND2_X1 U1151 ( .A1(n33242), .A2(n30769), .ZN(n32497) );
  NOR2_X1 U1153 ( .A1(n21652), .A2(n7553), .ZN(n33031) );
  OR2_X1 U1158 ( .A1(n21466), .A2(n31085), .Z(n32073) );
  INV_X1 U1160 ( .I(n32208), .ZN(n7366) );
  NAND2_X1 U1161 ( .A1(n21741), .A2(n423), .ZN(n33364) );
  NAND2_X1 U1165 ( .A1(n21625), .A2(n32865), .ZN(n32320) );
  NOR2_X1 U1168 ( .A1(n2643), .A2(n14681), .ZN(n21792) );
  INV_X1 U1171 ( .I(n32435), .ZN(n29286) );
  INV_X1 U1172 ( .I(n912), .ZN(n33842) );
  INV_X2 U1177 ( .I(n1013), .ZN(n32499) );
  OAI21_X1 U1180 ( .A1(n14384), .A2(n31042), .B(n32384), .ZN(n32208) );
  NAND2_X1 U1188 ( .A1(n21512), .A2(n26622), .ZN(n11719) );
  AND2_X1 U1190 ( .A1(n21860), .A2(n3286), .Z(n13116) );
  NOR2_X1 U1202 ( .A1(n11596), .A2(n11981), .ZN(n33520) );
  NAND2_X1 U1207 ( .A1(n13114), .A2(n30885), .ZN(n21586) );
  NAND2_X1 U1209 ( .A1(n12221), .A2(n21719), .ZN(n21490) );
  NAND3_X1 U1214 ( .A1(n33481), .A2(n21713), .A3(n5704), .ZN(n32994) );
  NAND2_X1 U1216 ( .A1(n12866), .A2(n13872), .ZN(n27023) );
  INV_X2 U1218 ( .I(n31956), .ZN(n1015) );
  INV_X1 U1219 ( .I(n2386), .ZN(n21489) );
  NOR2_X1 U1220 ( .A1(n30769), .A2(n32252), .ZN(n4432) );
  INV_X1 U1221 ( .I(n21604), .ZN(n1318) );
  INV_X1 U1222 ( .I(n21512), .ZN(n1327) );
  INV_X1 U1223 ( .I(n16954), .ZN(n21585) );
  INV_X2 U1225 ( .I(n1313), .ZN(n517) );
  INV_X1 U1228 ( .I(n33146), .ZN(n33731) );
  NAND2_X1 U1230 ( .A1(n2386), .A2(n31954), .ZN(n21717) );
  BUF_X2 U1239 ( .I(n7592), .Z(n33481) );
  INV_X1 U1245 ( .I(n31960), .ZN(n32643) );
  CLKBUF_X1 U1246 ( .I(n5086), .Z(n31953) );
  NAND2_X1 U1248 ( .A1(n32800), .A2(n15371), .ZN(n32372) );
  INV_X1 U1249 ( .I(n7592), .ZN(n16441) );
  INV_X1 U1250 ( .I(n12211), .ZN(n5228) );
  NAND2_X1 U1252 ( .A1(n21264), .A2(n21263), .ZN(n12640) );
  INV_X1 U1258 ( .I(n9472), .ZN(n5494) );
  INV_X1 U1260 ( .I(n3203), .ZN(n32505) );
  INV_X2 U1262 ( .I(n7868), .ZN(n27532) );
  AND2_X1 U1263 ( .A1(n21466), .A2(n1136), .Z(n4842) );
  OAI21_X1 U1264 ( .A1(n21222), .A2(n21109), .B(n26166), .ZN(n2570) );
  INV_X2 U1268 ( .I(n28099), .ZN(n777) );
  INV_X2 U1270 ( .I(n11755), .ZN(n7969) );
  NAND2_X1 U1271 ( .A1(n33802), .A2(n2834), .ZN(n5086) );
  NAND2_X1 U1272 ( .A1(n32455), .A2(n32454), .ZN(n21134) );
  NOR2_X1 U1277 ( .A1(n16204), .A2(n33167), .ZN(n17432) );
  NAND3_X1 U1281 ( .A1(n33926), .A2(n21336), .A3(n33925), .ZN(n5250) );
  NAND3_X1 U1286 ( .A1(n33755), .A2(n4988), .A3(n4324), .ZN(n4062) );
  NOR2_X1 U1291 ( .A1(n11138), .A2(n21411), .ZN(n2722) );
  OAI21_X1 U1296 ( .A1(n21403), .A2(n596), .B(n12654), .ZN(n29742) );
  OAI21_X1 U1301 ( .A1(n1867), .A2(n1868), .B(n21353), .ZN(n32330) );
  OR2_X1 U1309 ( .A1(n9191), .A2(n12323), .Z(n10573) );
  INV_X1 U1312 ( .I(n11299), .ZN(n31329) );
  AOI22_X1 U1313 ( .A1(n21099), .A2(n17437), .B1(n154), .B2(n21138), .ZN(
        n21067) );
  OAI22_X1 U1318 ( .A1(n29802), .A2(n21363), .B1(n21183), .B2(n21182), .ZN(
        n17685) );
  INV_X1 U1319 ( .I(n13593), .ZN(n8587) );
  NAND2_X1 U1321 ( .A1(n31730), .A2(n31728), .ZN(n18208) );
  AND2_X1 U1325 ( .A1(n2738), .A2(n9133), .Z(n29394) );
  INV_X1 U1328 ( .I(n32655), .ZN(n34081) );
  OR2_X1 U1329 ( .A1(n11967), .A2(n21358), .Z(n10092) );
  NOR2_X1 U1330 ( .A1(n4274), .A2(n17341), .ZN(n5039) );
  NOR2_X1 U1333 ( .A1(n32273), .A2(n8560), .ZN(n32407) );
  OAI21_X1 U1336 ( .A1(n31997), .A2(n5239), .B(n32203), .ZN(n32979) );
  NAND3_X1 U1342 ( .A1(n2831), .A2(n2833), .A3(n26167), .ZN(n33802) );
  NAND2_X1 U1343 ( .A1(n33972), .A2(n13073), .ZN(n13366) );
  NAND2_X1 U1345 ( .A1(n2370), .A2(n21441), .ZN(n32808) );
  OAI21_X1 U1358 ( .A1(n1020), .A2(n7007), .B(n3672), .ZN(n7051) );
  NOR2_X1 U1359 ( .A1(n26167), .A2(n1329), .ZN(n33113) );
  NOR3_X1 U1361 ( .A1(n31965), .A2(n28642), .A3(n29460), .ZN(n27608) );
  NAND2_X1 U1368 ( .A1(n5480), .A2(n32347), .ZN(n33925) );
  OAI21_X1 U1370 ( .A1(n922), .A2(n13255), .B(n6408), .ZN(n16640) );
  NOR2_X1 U1372 ( .A1(n32550), .A2(n1141), .ZN(n4497) );
  NAND2_X1 U1374 ( .A1(n32457), .A2(n32456), .ZN(n32455) );
  NAND2_X1 U1375 ( .A1(n5469), .A2(n26021), .ZN(n33523) );
  NOR2_X1 U1378 ( .A1(n4341), .A2(n30813), .ZN(n17011) );
  OAI22_X1 U1382 ( .A1(n810), .A2(n21365), .B1(n4076), .B2(n17466), .ZN(n29678) );
  NOR2_X1 U1383 ( .A1(n21251), .A2(n21078), .ZN(n30050) );
  NOR2_X1 U1385 ( .A1(n18106), .A2(n15522), .ZN(n33647) );
  INV_X1 U1386 ( .I(n21443), .ZN(n32457) );
  NAND2_X1 U1387 ( .A1(n32777), .A2(n32776), .ZN(n5018) );
  NAND2_X1 U1389 ( .A1(n2241), .A2(n2242), .ZN(n33735) );
  NAND2_X1 U1392 ( .A1(n16180), .A2(n16526), .ZN(n32456) );
  AND2_X1 U1394 ( .A1(n11967), .A2(n21358), .Z(n31674) );
  NAND2_X1 U1396 ( .A1(n21381), .A2(n16906), .ZN(n15985) );
  NAND2_X1 U1401 ( .A1(n21078), .A2(n4518), .ZN(n13401) );
  NAND2_X1 U1403 ( .A1(n14074), .A2(n21406), .ZN(n32322) );
  NAND2_X1 U1408 ( .A1(n33741), .A2(n4324), .ZN(n33171) );
  OR2_X1 U1418 ( .A1(n5395), .A2(n8028), .Z(n31997) );
  NAND2_X1 U1420 ( .A1(n21452), .A2(n780), .ZN(n29122) );
  BUF_X2 U1426 ( .I(n21438), .Z(n33745) );
  NOR2_X1 U1429 ( .A1(n21255), .A2(n28257), .ZN(n33137) );
  NAND2_X1 U1439 ( .A1(n33849), .A2(n32147), .ZN(n4076) );
  NOR2_X1 U1445 ( .A1(n33889), .A2(n33888), .ZN(n33887) );
  NOR2_X1 U1446 ( .A1(n17956), .A2(n349), .ZN(n32350) );
  NAND2_X1 U1447 ( .A1(n4337), .A2(n4971), .ZN(n32203) );
  NOR3_X1 U1448 ( .A1(n21163), .A2(n27170), .A3(n11734), .ZN(n33350) );
  NOR2_X1 U1450 ( .A1(n21219), .A2(n33496), .ZN(n32273) );
  NOR2_X1 U1455 ( .A1(n2738), .A2(n8924), .ZN(n8937) );
  NAND2_X1 U1457 ( .A1(n31909), .A2(n16668), .ZN(n21407) );
  INV_X2 U1459 ( .I(n16633), .ZN(n20949) );
  BUF_X2 U1460 ( .I(n3879), .Z(n30813) );
  BUF_X2 U1461 ( .I(n21395), .Z(n27955) );
  CLKBUF_X2 U1468 ( .I(n26677), .Z(n34131) );
  INV_X1 U1471 ( .I(n3193), .ZN(n32777) );
  BUF_X2 U1472 ( .I(n6493), .Z(n34054) );
  NAND2_X1 U1473 ( .A1(n6855), .A2(n32883), .ZN(n32239) );
  OAI21_X1 U1475 ( .A1(n349), .A2(n33496), .B(n33495), .ZN(n21146) );
  INV_X2 U1476 ( .I(n21452), .ZN(n1143) );
  OR2_X1 U1478 ( .A1(n34156), .A2(n28260), .Z(n31989) );
  INV_X1 U1487 ( .I(n4145), .ZN(n1703) );
  BUF_X2 U1488 ( .I(n9351), .Z(n9186) );
  CLKBUF_X2 U1489 ( .I(n13723), .Z(n32147) );
  NAND2_X1 U1490 ( .A1(n13692), .A2(n21357), .ZN(n33336) );
  INV_X1 U1509 ( .I(n29901), .ZN(n33496) );
  BUF_X2 U1510 ( .I(n10599), .Z(n33498) );
  BUF_X2 U1513 ( .I(n21258), .Z(n16652) );
  BUF_X2 U1516 ( .I(n13195), .Z(n10599) );
  OR2_X1 U1520 ( .A1(n31290), .A2(n31291), .Z(n32889) );
  INV_X1 U1523 ( .I(n20641), .ZN(n20920) );
  CLKBUF_X2 U1541 ( .I(n4680), .Z(n29918) );
  INV_X1 U1545 ( .I(n20970), .ZN(n29879) );
  INV_X1 U1546 ( .I(n20786), .ZN(n21024) );
  INV_X1 U1553 ( .I(n20928), .ZN(n12559) );
  NOR2_X1 U1555 ( .A1(n17317), .A2(n4980), .ZN(n32230) );
  NAND2_X1 U1570 ( .A1(n10105), .A2(n5735), .ZN(n5734) );
  OAI22_X1 U1572 ( .A1(n32033), .A2(n8031), .B1(n28799), .B2(n1356), .ZN(
        n32249) );
  NAND3_X1 U1573 ( .A1(n20302), .A2(n27600), .A3(n20360), .ZN(n12553) );
  OR2_X1 U1575 ( .A1(n14161), .A2(n20628), .Z(n20387) );
  NOR2_X1 U1576 ( .A1(n15898), .A2(n15027), .ZN(n11840) );
  AND2_X1 U1577 ( .A1(n20627), .A2(n9014), .Z(n14571) );
  OR2_X1 U1581 ( .A1(n20534), .A2(n28028), .Z(n30728) );
  AND2_X1 U1582 ( .A1(n33117), .A2(n14138), .Z(n2145) );
  AND2_X1 U1588 ( .A1(n33117), .A2(n20468), .Z(n3227) );
  AOI22_X1 U1591 ( .A1(n15638), .A2(n26756), .B1(n11017), .B2(n1347), .ZN(
        n33052) );
  CLKBUF_X2 U1593 ( .I(n28011), .Z(n34052) );
  NAND2_X1 U1594 ( .A1(n32765), .A2(n31891), .ZN(n32764) );
  NAND2_X1 U1597 ( .A1(n20607), .A2(n7577), .ZN(n33843) );
  NAND2_X1 U1601 ( .A1(n20551), .A2(n10834), .ZN(n12148) );
  NOR2_X1 U1602 ( .A1(n20243), .A2(n26471), .ZN(n32684) );
  NAND3_X1 U1604 ( .A1(n32941), .A2(n32940), .A3(n32939), .ZN(n29431) );
  NAND3_X1 U1606 ( .A1(n31969), .A2(n20072), .A3(n20073), .ZN(n3904) );
  NOR3_X1 U1610 ( .A1(n15898), .A2(n16518), .A3(n20534), .ZN(n184) );
  AND2_X1 U1615 ( .A1(n33117), .A2(n20467), .Z(n3463) );
  AND2_X1 U1619 ( .A1(n16144), .A2(n11984), .Z(n20194) );
  INV_X1 U1628 ( .I(n20608), .ZN(n33397) );
  INV_X1 U1641 ( .I(n10312), .ZN(n29553) );
  AND2_X1 U1643 ( .A1(n20515), .A2(n7242), .Z(n6121) );
  BUF_X2 U1649 ( .I(n30643), .Z(n4071) );
  CLKBUF_X2 U1653 ( .I(n20632), .Z(n111) );
  NAND2_X1 U1657 ( .A1(n12421), .A2(n14719), .ZN(n17672) );
  BUF_X2 U1660 ( .I(n30763), .Z(n31961) );
  CLKBUF_X1 U1662 ( .I(n14545), .Z(n29623) );
  INV_X1 U1666 ( .I(n31811), .ZN(n33398) );
  NAND2_X1 U1671 ( .A1(n28085), .A2(n20563), .ZN(n33194) );
  NAND2_X1 U1675 ( .A1(n20492), .A2(n26585), .ZN(n33944) );
  NAND2_X1 U1677 ( .A1(n3084), .A2(n20339), .ZN(n12244) );
  NOR2_X1 U1683 ( .A1(n25966), .A2(n20602), .ZN(n32341) );
  NAND2_X1 U1686 ( .A1(n9403), .A2(n20472), .ZN(n34113) );
  NOR2_X1 U1689 ( .A1(n12966), .A2(n12421), .ZN(n33734) );
  AND2_X1 U1692 ( .A1(n26566), .A2(n32989), .Z(n31975) );
  INV_X1 U1696 ( .I(n30643), .ZN(n10106) );
  INV_X1 U1697 ( .I(n3157), .ZN(n33091) );
  NOR2_X1 U1699 ( .A1(n16218), .A2(n7486), .ZN(n33776) );
  INV_X1 U1701 ( .I(n20549), .ZN(n31390) );
  BUF_X2 U1704 ( .I(n28840), .Z(n33730) );
  OR2_X1 U1707 ( .A1(n20613), .A2(n9252), .Z(n7872) );
  NAND2_X1 U1709 ( .A1(n28028), .A2(n32240), .ZN(n11036) );
  NAND2_X1 U1710 ( .A1(n20630), .A2(n31471), .ZN(n15225) );
  OAI21_X1 U1716 ( .A1(n939), .A2(n31442), .B(n19949), .ZN(n17496) );
  NAND2_X1 U1717 ( .A1(n30845), .A2(n149), .ZN(n34032) );
  NAND2_X1 U1718 ( .A1(n32377), .A2(n19820), .ZN(n11402) );
  NOR2_X1 U1719 ( .A1(n32197), .A2(n29187), .ZN(n2550) );
  OAI21_X1 U1721 ( .A1(n31993), .A2(n11142), .B(n29233), .ZN(n11141) );
  NAND2_X1 U1722 ( .A1(n11510), .A2(n12398), .ZN(n32956) );
  OAI21_X1 U1724 ( .A1(n31593), .A2(n16159), .B(n20033), .ZN(n33732) );
  NAND2_X1 U1728 ( .A1(n34006), .A2(n16489), .ZN(n3094) );
  OAI21_X1 U1732 ( .A1(n4215), .A2(n16346), .B(n34051), .ZN(n17242) );
  OAI21_X1 U1735 ( .A1(n19996), .A2(n19922), .B(n4674), .ZN(n4266) );
  NOR2_X1 U1737 ( .A1(n19932), .A2(n8817), .ZN(n10440) );
  NAND2_X1 U1738 ( .A1(n13569), .A2(n19925), .ZN(n32719) );
  AOI21_X1 U1743 ( .A1(n431), .A2(n19840), .B(n33504), .ZN(n16924) );
  NAND2_X1 U1746 ( .A1(n4215), .A2(n17243), .ZN(n34051) );
  INV_X1 U1751 ( .I(n6961), .ZN(n33148) );
  NOR3_X1 U1753 ( .A1(n20135), .A2(n32141), .A3(n12682), .ZN(n30155) );
  NAND2_X1 U1754 ( .A1(n9619), .A2(n1168), .ZN(n32674) );
  NOR2_X1 U1755 ( .A1(n4371), .A2(n19998), .ZN(n15366) );
  NOR2_X1 U1756 ( .A1(n19854), .A2(n19855), .ZN(n20070) );
  NAND2_X1 U1758 ( .A1(n7309), .A2(n3090), .ZN(n33439) );
  OAI21_X1 U1761 ( .A1(n3989), .A2(n11961), .B(n33627), .ZN(n28459) );
  NOR2_X1 U1763 ( .A1(n12075), .A2(n17495), .ZN(n34006) );
  NOR2_X1 U1765 ( .A1(n20020), .A2(n20120), .ZN(n19812) );
  NAND2_X1 U1768 ( .A1(n19898), .A2(n16092), .ZN(n14712) );
  NAND2_X1 U1769 ( .A1(n29853), .A2(n19961), .ZN(n33504) );
  NOR2_X1 U1770 ( .A1(n15192), .A2(n29040), .ZN(n15477) );
  NAND2_X1 U1773 ( .A1(n16977), .A2(n19920), .ZN(n32792) );
  AOI21_X1 U1775 ( .A1(n33264), .A2(n16848), .B(n13583), .ZN(n33553) );
  INV_X1 U1778 ( .I(n1826), .ZN(n33526) );
  NOR2_X1 U1785 ( .A1(n5966), .A2(n6962), .ZN(n32479) );
  NAND3_X1 U1786 ( .A1(n8259), .A2(n11199), .A3(n20154), .ZN(n19621) );
  INV_X1 U1789 ( .I(n10286), .ZN(n32197) );
  OAI21_X1 U1790 ( .A1(n13348), .A2(n6444), .B(n822), .ZN(n33769) );
  NAND3_X1 U1791 ( .A1(n7460), .A2(n16491), .A3(n7461), .ZN(n1814) );
  NOR3_X1 U1793 ( .A1(n19992), .A2(n19993), .A3(n1170), .ZN(n33271) );
  INV_X1 U1794 ( .I(n26237), .ZN(n33714) );
  OR2_X1 U1796 ( .A1(n16625), .A2(n17127), .Z(n8137) );
  AND2_X1 U1798 ( .A1(n16595), .A2(n14815), .Z(n9450) );
  AND2_X1 U1802 ( .A1(n28293), .A2(n17882), .Z(n31991) );
  NOR2_X1 U1805 ( .A1(n28293), .A2(n16681), .ZN(n19842) );
  AND2_X1 U1815 ( .A1(n27748), .A2(n26237), .Z(n11949) );
  OR2_X1 U1816 ( .A1(n11720), .A2(n10934), .Z(n14306) );
  NOR2_X1 U1819 ( .A1(n6344), .A2(n29446), .ZN(n19950) );
  CLKBUF_X2 U1824 ( .I(n6275), .Z(n26615) );
  INV_X1 U1825 ( .I(n19966), .ZN(n14575) );
  BUF_X2 U1827 ( .I(n19833), .Z(n20136) );
  BUF_X2 U1834 ( .I(n11720), .Z(n29187) );
  INV_X2 U1838 ( .I(n19938), .ZN(n1161) );
  INV_X1 U1840 ( .I(n32915), .ZN(n19885) );
  INV_X1 U1842 ( .I(n9161), .ZN(n19616) );
  NAND2_X1 U1846 ( .A1(n6022), .A2(n19056), .ZN(n11867) );
  CLKBUF_X2 U1850 ( .I(n19778), .Z(n28908) );
  INV_X1 U1853 ( .I(n24831), .ZN(n32981) );
  INV_X1 U1858 ( .I(n19778), .ZN(n33995) );
  OAI21_X1 U1859 ( .A1(n17677), .A2(n17678), .B(n31970), .ZN(n33088) );
  OAI21_X1 U1861 ( .A1(n28025), .A2(n18230), .B(n763), .ZN(n32431) );
  AOI22_X1 U1863 ( .A1(n19119), .A2(n19181), .B1(n29769), .B2(n14424), .ZN(
        n14423) );
  OR2_X1 U1866 ( .A1(n28949), .A2(n19080), .Z(n32057) );
  NOR2_X1 U1870 ( .A1(n27965), .A2(n25967), .ZN(n33825) );
  NAND2_X1 U1872 ( .A1(n19074), .A2(n30760), .ZN(n33852) );
  NAND2_X1 U1884 ( .A1(n19311), .A2(n19312), .ZN(n9683) );
  NOR2_X1 U1888 ( .A1(n1807), .A2(n4643), .ZN(n401) );
  NOR2_X1 U1889 ( .A1(n26518), .A2(n11085), .ZN(n11802) );
  CLKBUF_X1 U1892 ( .I(n29815), .Z(n33635) );
  CLKBUF_X1 U1894 ( .I(n30894), .Z(n33712) );
  AND2_X1 U1896 ( .A1(n10472), .A2(n31970), .Z(n32011) );
  NAND2_X1 U1900 ( .A1(n4714), .A2(n9646), .ZN(n16874) );
  AOI21_X1 U1902 ( .A1(n11074), .A2(n3093), .B(n2081), .ZN(n28345) );
  NAND2_X1 U1903 ( .A1(n33967), .A2(n4643), .ZN(n30661) );
  AOI21_X1 U1910 ( .A1(n826), .A2(n19290), .B(n19288), .ZN(n2717) );
  OAI21_X1 U1911 ( .A1(n33143), .A2(n19147), .B(n15534), .ZN(n32293) );
  AND2_X1 U1914 ( .A1(n7810), .A2(n19249), .Z(n9648) );
  OAI21_X1 U1915 ( .A1(n32653), .A2(n26037), .B(n17311), .ZN(n17819) );
  INV_X1 U1918 ( .I(n19348), .ZN(n33232) );
  INV_X1 U1919 ( .I(n9677), .ZN(n32219) );
  INV_X1 U1924 ( .I(n5625), .ZN(n18977) );
  NOR2_X1 U1925 ( .A1(n25960), .A2(n4747), .ZN(n33671) );
  INV_X1 U1927 ( .I(n19308), .ZN(n33718) );
  NOR2_X1 U1928 ( .A1(n19102), .A2(n944), .ZN(n8192) );
  INV_X1 U1937 ( .I(n18945), .ZN(n33967) );
  INV_X1 U1940 ( .I(n28379), .ZN(n32138) );
  NAND2_X1 U1941 ( .A1(n19078), .A2(n30501), .ZN(n30933) );
  INV_X1 U1942 ( .I(n19260), .ZN(n32790) );
  INV_X1 U1949 ( .I(n31947), .ZN(n27970) );
  BUF_X2 U1951 ( .I(n10228), .Z(n10227) );
  NOR2_X1 U1952 ( .A1(n18976), .A2(n14892), .ZN(n18945) );
  NAND2_X1 U1953 ( .A1(n764), .A2(n19167), .ZN(n10353) );
  AOI22_X1 U1958 ( .A1(n18641), .A2(n28238), .B1(n4259), .B2(n18642), .ZN(
        n32121) );
  NOR2_X1 U1959 ( .A1(n18974), .A2(n11322), .ZN(n34031) );
  CLKBUF_X2 U1963 ( .I(n30865), .Z(n31948) );
  INV_X2 U1965 ( .I(n18017), .ZN(n1384) );
  AOI22_X1 U1967 ( .A1(n18506), .A2(n9729), .B1(n18507), .B2(n1439), .ZN(
        n33396) );
  BUF_X4 U1973 ( .I(n10953), .Z(n2612) );
  NOR2_X1 U1974 ( .A1(n18866), .A2(n711), .ZN(n2507) );
  NOR2_X1 U1976 ( .A1(n33528), .A2(n33559), .ZN(n13112) );
  AND2_X1 U1979 ( .A1(n18566), .A2(n18324), .Z(n32009) );
  OAI21_X1 U1983 ( .A1(n18702), .A2(n16352), .B(n33736), .ZN(n18431) );
  OAI21_X1 U1984 ( .A1(n18866), .A2(n10283), .B(n18871), .ZN(n10220) );
  OAI21_X1 U1985 ( .A1(n18112), .A2(n18672), .B(n16572), .ZN(n33324) );
  NOR2_X1 U1988 ( .A1(n4259), .A2(n18768), .ZN(n33799) );
  NAND2_X1 U1992 ( .A1(n18510), .A2(n16352), .ZN(n33736) );
  NOR2_X1 U2009 ( .A1(n28009), .A2(n28010), .ZN(n33559) );
  NAND2_X1 U2013 ( .A1(n33997), .A2(n33999), .ZN(n32763) );
  NAND2_X1 U2015 ( .A1(n32411), .A2(n29309), .ZN(n32410) );
  NOR2_X1 U2016 ( .A1(n18603), .A2(n18602), .ZN(n32491) );
  NAND3_X1 U2019 ( .A1(n10043), .A2(n17255), .A3(n17223), .ZN(n32294) );
  NAND3_X1 U2021 ( .A1(n15108), .A2(n16881), .A3(n17255), .ZN(n10561) );
  NAND2_X1 U2022 ( .A1(n33999), .A2(n18672), .ZN(n9289) );
  NOR2_X1 U2023 ( .A1(n8400), .A2(n16614), .ZN(n18859) );
  INV_X1 U2027 ( .I(n18228), .ZN(n10903) );
  AND2_X1 U2032 ( .A1(n29315), .A2(n18397), .Z(n31986) );
  INV_X1 U2039 ( .I(n16995), .ZN(n15406) );
  INV_X2 U2046 ( .I(n6860), .ZN(n18854) );
  NOR2_X1 U2054 ( .A1(n18702), .A2(n18510), .ZN(n33792) );
  NOR2_X1 U2055 ( .A1(n10325), .A2(n18677), .ZN(n18679) );
  NAND2_X1 U2057 ( .A1(n18738), .A2(n17166), .ZN(n33207) );
  NAND2_X1 U2063 ( .A1(n16287), .A2(n31417), .ZN(n8860) );
  NAND2_X1 U2066 ( .A1(n16372), .A2(n12863), .ZN(n7497) );
  INV_X1 U2067 ( .I(n28245), .ZN(n6359) );
  BUF_X2 U2074 ( .I(n18295), .Z(n18324) );
  BUF_X2 U2079 ( .I(n18861), .Z(n16287) );
  BUF_X2 U2080 ( .I(n34110), .Z(n33093) );
  NAND2_X1 U2084 ( .A1(n18006), .A2(n30271), .ZN(n33040) );
  INV_X2 U2088 ( .I(n29309), .ZN(n33989) );
  BUF_X2 U2093 ( .I(n32096), .Z(n32798) );
  INV_X4 U2094 ( .I(n15716), .ZN(n727) );
  NAND3_X1 U2098 ( .A1(n18099), .A2(n15867), .A3(n6910), .ZN(n28217) );
  NAND2_X2 U2100 ( .A1(n22878), .A2(n23057), .ZN(n22933) );
  NAND2_X2 U2105 ( .A1(n27046), .A2(n25577), .ZN(n33305) );
  NOR2_X2 U2108 ( .A1(n123), .A2(n31327), .ZN(n2656) );
  NAND3_X2 U2112 ( .A1(n23177), .A2(n14350), .A3(n14756), .ZN(n23178) );
  INV_X2 U2118 ( .I(n8778), .ZN(n27150) );
  OAI22_X2 U2120 ( .A1(n15284), .A2(n10472), .B1(n11072), .B2(n2081), .ZN(
        n16909) );
  BUF_X4 U2130 ( .I(n24339), .Z(n16552) );
  NAND3_X2 U2132 ( .A1(n27833), .A2(n28917), .A3(n25609), .ZN(n28156) );
  NAND2_X2 U2136 ( .A1(n18261), .A2(n26739), .ZN(n22860) );
  INV_X2 U2137 ( .I(n23746), .ZN(n11392) );
  NOR2_X2 U2139 ( .A1(n32855), .A2(n25615), .ZN(n25607) );
  BUF_X2 U2141 ( .I(n23849), .Z(n31435) );
  NOR2_X1 U2144 ( .A1(n32301), .A2(n4607), .ZN(n8653) );
  NAND2_X2 U2147 ( .A1(n24262), .A2(n7809), .ZN(n15974) );
  NOR2_X2 U2152 ( .A1(n24104), .A2(n26750), .ZN(n24102) );
  NOR2_X2 U2153 ( .A1(n7093), .A2(n29566), .ZN(n2853) );
  BUF_X4 U2155 ( .I(n2860), .Z(n28957) );
  INV_X2 U2156 ( .I(n3181), .ZN(n32186) );
  NOR2_X2 U2158 ( .A1(n27651), .A2(n27461), .ZN(n33643) );
  NAND2_X2 U2159 ( .A1(n28181), .A2(n8140), .ZN(n21460) );
  OR2_X2 U2160 ( .A1(n4646), .A2(n31957), .Z(n32079) );
  NAND2_X2 U2163 ( .A1(n1015), .A2(n38), .ZN(n8825) );
  INV_X4 U2167 ( .I(n28840), .ZN(n26756) );
  INV_X2 U2169 ( .I(n25653), .ZN(n734) );
  AND2_X2 U2172 ( .A1(n30365), .A2(n22786), .Z(n32088) );
  NAND3_X2 U2173 ( .A1(n4436), .A2(n7810), .A3(n7680), .ZN(n4591) );
  NAND2_X2 U2175 ( .A1(n7093), .A2(n14839), .ZN(n24344) );
  BUF_X2 U2182 ( .I(n7293), .Z(n31957) );
  NAND2_X2 U2189 ( .A1(n29634), .A2(n14619), .ZN(n24153) );
  NAND2_X2 U2190 ( .A1(n25452), .A2(n15212), .ZN(n25430) );
  NAND2_X2 U2191 ( .A1(n5820), .A2(n28957), .ZN(n32712) );
  NAND3_X2 U2194 ( .A1(n15580), .A2(n6553), .A3(n30364), .ZN(n15579) );
  NOR2_X2 U2196 ( .A1(n7116), .A2(n12184), .ZN(n30148) );
  INV_X2 U2197 ( .I(n15051), .ZN(n15060) );
  INV_X2 U2199 ( .I(n22033), .ZN(n11727) );
  OAI22_X2 U2204 ( .A1(n30934), .A2(n18567), .B1(n17316), .B2(n17813), .ZN(
        n18423) );
  NAND2_X2 U2206 ( .A1(n18423), .A2(n18493), .ZN(n16806) );
  NAND2_X2 U2207 ( .A1(n9620), .A2(n22377), .ZN(n8176) );
  NAND2_X2 U2208 ( .A1(n24251), .A2(n3220), .ZN(n28827) );
  BUF_X4 U2209 ( .I(n23285), .Z(n3868) );
  BUF_X4 U2212 ( .I(n12617), .Z(n4774) );
  BUF_X2 U2213 ( .I(n15613), .Z(n32975) );
  AND2_X1 U2214 ( .A1(n9377), .A2(n23018), .Z(n33862) );
  BUF_X2 U2216 ( .I(n31453), .Z(n2391) );
  NOR2_X2 U2217 ( .A1(n13712), .A2(n21251), .ZN(n16204) );
  NAND2_X2 U2219 ( .A1(n16387), .A2(n4216), .ZN(n33044) );
  OAI21_X2 U2220 ( .A1(n3731), .A2(n3732), .B(n25236), .ZN(n3730) );
  BUF_X2 U2222 ( .I(n32051), .Z(n16389) );
  INV_X2 U2224 ( .I(n24269), .ZN(n33891) );
  BUF_X2 U2225 ( .I(n8808), .Z(n8301) );
  NOR2_X2 U2227 ( .A1(n14752), .A2(n10099), .ZN(n24904) );
  NAND2_X2 U2228 ( .A1(n30252), .A2(n28069), .ZN(n23750) );
  NAND2_X1 U2229 ( .A1(n11597), .A2(n11596), .ZN(n32739) );
  NOR3_X2 U2235 ( .A1(n14463), .A2(n16496), .A3(n29965), .ZN(n3445) );
  OAI21_X2 U2236 ( .A1(n19165), .A2(n11085), .B(n11444), .ZN(n11474) );
  NOR2_X1 U2238 ( .A1(n5304), .A2(n5305), .ZN(n33385) );
  INV_X2 U2240 ( .I(n6402), .ZN(n28200) );
  OAI21_X2 U2244 ( .A1(n21434), .A2(n5049), .B(n8010), .ZN(n21074) );
  INV_X2 U2248 ( .I(n16809), .ZN(n28658) );
  NOR2_X2 U2249 ( .A1(n28408), .A2(n13762), .ZN(n22861) );
  INV_X2 U2250 ( .I(n29213), .ZN(n584) );
  NAND3_X1 U2253 ( .A1(n32354), .A2(n7505), .A3(n7504), .ZN(n24314) );
  OR2_X1 U2257 ( .A1(n9159), .A2(n8602), .Z(n25944) );
  BUF_X2 U2258 ( .I(n22579), .Z(n16149) );
  AOI22_X2 U2260 ( .A1(n1315), .A2(n33857), .B1(n8569), .B2(n5078), .ZN(n5077)
         );
  NOR2_X2 U2262 ( .A1(n34009), .A2(n34008), .ZN(n6321) );
  OAI21_X2 U2263 ( .A1(n33808), .A2(n29965), .B(n28061), .ZN(n33759) );
  NAND2_X2 U2264 ( .A1(n1951), .A2(n25072), .ZN(n10301) );
  NOR3_X1 U2267 ( .A1(n33295), .A2(n30969), .A3(n24087), .ZN(n14197) );
  NAND3_X1 U2276 ( .A1(n2937), .A2(n8308), .A3(n23224), .ZN(n2803) );
  INV_X1 U2277 ( .I(n23224), .ZN(n26311) );
  CLKBUF_X4 U2278 ( .I(n20565), .Z(n17329) );
  NOR2_X1 U2280 ( .A1(n25681), .A2(n29243), .ZN(n25682) );
  NAND2_X1 U2289 ( .A1(n32879), .A2(n25675), .ZN(n25681) );
  NAND2_X1 U2296 ( .A1(n25002), .A2(n3229), .ZN(n2266) );
  AOI21_X1 U2297 ( .A1(n16127), .A2(n1134), .B(n6074), .ZN(n6678) );
  NAND2_X1 U2306 ( .A1(n15217), .A2(n20608), .ZN(n31714) );
  NOR2_X1 U2310 ( .A1(n7290), .A2(n20608), .ZN(n20186) );
  INV_X1 U2311 ( .I(n29815), .ZN(n32951) );
  NAND2_X1 U2312 ( .A1(n9646), .A2(n29815), .ZN(n7575) );
  BUF_X2 U2319 ( .I(n28714), .Z(n26133) );
  NOR2_X1 U2320 ( .A1(n4041), .A2(n17313), .ZN(n21158) );
  NAND2_X1 U2322 ( .A1(n13579), .A2(n22033), .ZN(n11728) );
  INV_X1 U2328 ( .I(n11205), .ZN(n29927) );
  INV_X2 U2332 ( .I(n6593), .ZN(n22956) );
  NOR2_X1 U2335 ( .A1(n6593), .A2(n15601), .ZN(n26047) );
  OAI21_X1 U2344 ( .A1(n4918), .A2(n1294), .B(n26884), .ZN(n10611) );
  NAND2_X1 U2346 ( .A1(n16964), .A2(n16963), .ZN(n16962) );
  CLKBUF_X1 U2347 ( .I(n10285), .Z(n28743) );
  AOI21_X1 U2349 ( .A1(n22379), .A2(n33966), .B(n636), .ZN(n22380) );
  CLKBUF_X1 U2351 ( .I(n21079), .Z(n32357) );
  NAND2_X1 U2354 ( .A1(n11652), .A2(n11651), .ZN(n8989) );
  NAND2_X1 U2355 ( .A1(n28568), .A2(n857), .ZN(n6062) );
  NAND2_X1 U2356 ( .A1(n9028), .A2(n32583), .ZN(n25176) );
  AOI21_X1 U2361 ( .A1(n20112), .A2(n20113), .B(n27808), .ZN(n20116) );
  AOI22_X1 U2362 ( .A1(n26787), .A2(n30230), .B1(n33624), .B2(n24337), .ZN(
        n2401) );
  NOR2_X1 U2365 ( .A1(n24244), .A2(n28374), .ZN(n26787) );
  AOI22_X1 U2369 ( .A1(n26367), .A2(n9370), .B1(n22503), .B2(n3332), .ZN(
        n31162) );
  NOR2_X1 U2375 ( .A1(n10202), .A2(n22503), .ZN(n22404) );
  INV_X1 U2376 ( .I(n11898), .ZN(n17781) );
  NOR3_X1 U2378 ( .A1(n10931), .A2(n28131), .A3(n137), .ZN(n2138) );
  AOI21_X1 U2380 ( .A1(n30205), .A2(n11629), .B(n28131), .ZN(n16964) );
  OAI22_X1 U2383 ( .A1(n14170), .A2(n25916), .B1(n25912), .B2(n25923), .ZN(
        n14067) );
  AOI21_X1 U2389 ( .A1(n1206), .A2(n25923), .B(n690), .ZN(n11156) );
  AOI21_X1 U2392 ( .A1(n25909), .A2(n1206), .B(n14067), .ZN(n8394) );
  NAND2_X1 U2393 ( .A1(n28743), .A2(n25743), .ZN(n25734) );
  OAI22_X1 U2398 ( .A1(n28743), .A2(n1597), .B1(n32863), .B2(n25746), .ZN(
        n25750) );
  NOR2_X1 U2399 ( .A1(n3019), .A2(n3229), .ZN(n25005) );
  NAND2_X1 U2400 ( .A1(n28639), .A2(n7862), .ZN(n3208) );
  NOR2_X1 U2401 ( .A1(n12861), .A2(n16688), .ZN(n27662) );
  INV_X2 U2402 ( .I(n16688), .ZN(n27661) );
  NAND2_X1 U2403 ( .A1(n18204), .A2(n29498), .ZN(n31266) );
  NAND2_X1 U2409 ( .A1(n1086), .A2(n24220), .ZN(n14445) );
  AOI21_X1 U2410 ( .A1(n1086), .A2(n24220), .B(n16688), .ZN(n14447) );
  NAND2_X1 U2411 ( .A1(n791), .A2(n24220), .ZN(n12862) );
  NAND3_X1 U2412 ( .A1(n25854), .A2(n14199), .A3(n10897), .ZN(n15544) );
  INV_X1 U2414 ( .I(n21530), .ZN(n33325) );
  OR2_X1 U2418 ( .A1(n21530), .A2(n29980), .Z(n31930) );
  NAND2_X1 U2420 ( .A1(n15456), .A2(n3614), .ZN(n22808) );
  NAND2_X1 U2422 ( .A1(n15456), .A2(n12315), .ZN(n15457) );
  NOR2_X1 U2423 ( .A1(n1997), .A2(n1995), .ZN(n24842) );
  INV_X2 U2430 ( .I(n700), .ZN(n1223) );
  OAI21_X1 U2433 ( .A1(n24249), .A2(n24248), .B(n24250), .ZN(n32976) );
  OAI22_X1 U2434 ( .A1(n4070), .A2(n1182), .B1(n10713), .B2(n30472), .ZN(n7493) );
  NAND2_X1 U2437 ( .A1(n30651), .A2(n24207), .ZN(n31160) );
  NAND2_X1 U2445 ( .A1(n2427), .A2(n24030), .ZN(n33963) );
  NAND2_X1 U2450 ( .A1(n5611), .A2(n25236), .ZN(n16400) );
  NAND2_X1 U2451 ( .A1(n25236), .A2(n25234), .ZN(n25133) );
  NOR2_X1 U2458 ( .A1(n25875), .A2(n717), .ZN(n13822) );
  CLKBUF_X1 U2461 ( .I(n7554), .Z(n33702) );
  INV_X2 U2466 ( .I(n24150), .ZN(n24317) );
  BUF_X1 U2469 ( .I(n25664), .Z(n3883) );
  INV_X2 U2470 ( .I(n8370), .ZN(n23892) );
  NOR2_X1 U2472 ( .A1(n8370), .A2(n28266), .ZN(n33827) );
  NAND2_X1 U2474 ( .A1(n8370), .A2(n23894), .ZN(n33829) );
  BUF_X2 U2475 ( .I(n8370), .Z(n32434) );
  OAI22_X1 U2476 ( .A1(n24737), .A2(n27162), .B1(n25836), .B2(n25860), .ZN(
        n28887) );
  INV_X2 U2477 ( .I(n24909), .ZN(n14752) );
  NAND2_X1 U2478 ( .A1(n24205), .A2(n24204), .ZN(n4519) );
  INV_X1 U2479 ( .I(n24205), .ZN(n33549) );
  NAND2_X1 U2481 ( .A1(n32328), .A2(n31160), .ZN(n24205) );
  NAND2_X1 U2486 ( .A1(n33543), .A2(n29056), .ZN(n29520) );
  OAI21_X1 U2487 ( .A1(n24260), .A2(n30280), .B(n8248), .ZN(n33543) );
  OAI21_X1 U2489 ( .A1(n32872), .A2(n15641), .B(n25184), .ZN(n9192) );
  CLKBUF_X1 U2490 ( .I(n24779), .Z(n32872) );
  NOR2_X1 U2492 ( .A1(n24994), .A2(n5072), .ZN(n26440) );
  NAND2_X1 U2494 ( .A1(n24902), .A2(n10755), .ZN(n24913) );
  INV_X1 U2499 ( .I(n10755), .ZN(n24903) );
  AOI21_X1 U2500 ( .A1(n16148), .A2(n22437), .B(n14219), .ZN(n4629) );
  INV_X1 U2501 ( .I(n3208), .ZN(n32100) );
  AOI21_X1 U2504 ( .A1(n26988), .A2(n6075), .B(n30783), .ZN(n2174) );
  NAND3_X1 U2507 ( .A1(n5411), .A2(n11019), .A3(n1206), .ZN(n25919) );
  OAI21_X1 U2508 ( .A1(n6154), .A2(n14075), .B(n24911), .ZN(n8980) );
  INV_X1 U2510 ( .I(n9247), .ZN(n25194) );
  NOR3_X1 U2514 ( .A1(n32577), .A2(n27062), .A3(n14837), .ZN(n8440) );
  NOR3_X1 U2515 ( .A1(n15078), .A2(n15079), .A3(n42), .ZN(n32577) );
  NAND2_X1 U2525 ( .A1(n32611), .A2(n32609), .ZN(n11670) );
  NAND2_X1 U2527 ( .A1(n32531), .A2(n22944), .ZN(n10108) );
  NOR2_X1 U2531 ( .A1(n22944), .A2(n3657), .ZN(n3659) );
  INV_X1 U2532 ( .I(n23171), .ZN(n8068) );
  NOR2_X1 U2533 ( .A1(n4193), .A2(n27668), .ZN(n25097) );
  NAND2_X1 U2536 ( .A1(n27668), .A2(n1203), .ZN(n25088) );
  CLKBUF_X1 U2539 ( .I(n11360), .Z(n27668) );
  NOR2_X1 U2542 ( .A1(n24984), .A2(n14454), .ZN(n16566) );
  OAI22_X1 U2543 ( .A1(n24984), .A2(n3080), .B1(n1081), .B2(n27926), .ZN(
        n17378) );
  NOR2_X1 U2550 ( .A1(n24213), .A2(n26914), .ZN(n342) );
  NAND2_X1 U2551 ( .A1(n3376), .A2(n7831), .ZN(n24988) );
  INV_X1 U2552 ( .I(n9963), .ZN(n10296) );
  BUF_X2 U2556 ( .I(n9963), .Z(n4750) );
  NAND3_X1 U2557 ( .A1(n6713), .A2(n7891), .A3(n793), .ZN(n24016) );
  NOR2_X1 U2559 ( .A1(n8835), .A2(n23750), .ZN(n23169) );
  NAND2_X1 U2560 ( .A1(n15059), .A2(n15062), .ZN(n15058) );
  AOI21_X1 U2561 ( .A1(n5178), .A2(n23482), .B(n22783), .ZN(n5681) );
  AOI21_X1 U2562 ( .A1(n25236), .A2(n25235), .B(n1216), .ZN(n4551) );
  NAND2_X1 U2563 ( .A1(n25128), .A2(n15323), .ZN(n25127) );
  AOI22_X1 U2569 ( .A1(n18497), .A2(n19087), .B1(n19088), .B2(n28171), .ZN(
        n18505) );
  NOR3_X1 U2577 ( .A1(n33093), .A2(n14248), .A3(n33101), .ZN(n29366) );
  BUF_X1 U2586 ( .I(n25228), .Z(n28388) );
  CLKBUF_X4 U2588 ( .I(n11887), .Z(n31807) );
  NOR3_X1 U2591 ( .A1(n33583), .A2(n11887), .A3(n23942), .ZN(n10020) );
  OR2_X1 U2592 ( .A1(n3103), .A2(n16022), .Z(n7626) );
  NAND2_X1 U2598 ( .A1(n6491), .A2(n20517), .ZN(n33240) );
  NAND2_X1 U2601 ( .A1(n27267), .A2(n6336), .ZN(n6334) );
  BUF_X2 U2603 ( .I(n3634), .Z(n28239) );
  AND2_X1 U2604 ( .A1(n15179), .A2(n2558), .Z(n6772) );
  OAI21_X1 U2605 ( .A1(n13560), .A2(n25587), .B(n15964), .ZN(n13559) );
  AOI21_X1 U2606 ( .A1(n24631), .A2(n25587), .B(n24633), .ZN(n11824) );
  CLKBUF_X2 U2612 ( .I(n17306), .Z(n31456) );
  NOR2_X1 U2614 ( .A1(n28329), .A2(n26415), .ZN(n2021) );
  NOR2_X1 U2619 ( .A1(n2141), .A2(n24335), .ZN(n33624) );
  INV_X1 U2622 ( .I(n16269), .ZN(n910) );
  BUF_X2 U2629 ( .I(n16269), .Z(n31105) );
  NAND3_X1 U2633 ( .A1(n16269), .A2(n21680), .A3(n21681), .ZN(n6570) );
  NAND2_X1 U2635 ( .A1(n25229), .A2(n28388), .ZN(n25261) );
  NOR3_X1 U2643 ( .A1(n25227), .A2(n15705), .A3(n15738), .ZN(n5532) );
  AOI21_X1 U2647 ( .A1(n33900), .A2(n10608), .B(n733), .ZN(n10606) );
  NAND3_X1 U2649 ( .A1(n733), .A2(n25278), .A3(n28532), .ZN(n24590) );
  NAND2_X1 U2652 ( .A1(n24262), .A2(n3205), .ZN(n8248) );
  NAND2_X1 U2654 ( .A1(n32859), .A2(n5713), .ZN(n28639) );
  CLKBUF_X2 U2656 ( .I(n20994), .Z(n28687) );
  INV_X1 U2657 ( .I(n20994), .ZN(n1339) );
  NAND2_X1 U2662 ( .A1(n28752), .A2(n17974), .ZN(n20994) );
  NOR2_X1 U2663 ( .A1(n14386), .A2(n24044), .ZN(n14249) );
  NAND3_X1 U2664 ( .A1(n25346), .A2(n24506), .A3(n753), .ZN(n10330) );
  AOI22_X1 U2665 ( .A1(n25732), .A2(n33386), .B1(n25730), .B2(n25731), .ZN(
        n32508) );
  NAND2_X1 U2667 ( .A1(n31941), .A2(n11704), .ZN(n24588) );
  OAI21_X1 U2680 ( .A1(n31941), .A2(n25392), .B(n13993), .ZN(n25442) );
  BUF_X2 U2686 ( .I(n28632), .Z(n31229) );
  NOR2_X1 U2689 ( .A1(n9181), .A2(n25820), .ZN(n25807) );
  NAND2_X1 U2691 ( .A1(n221), .A2(n13617), .ZN(n25569) );
  INV_X1 U2692 ( .I(n13617), .ZN(n6111) );
  NAND2_X1 U2693 ( .A1(n13617), .A2(n691), .ZN(n27046) );
  NAND2_X1 U2696 ( .A1(n13617), .A2(n8168), .ZN(n25568) );
  NAND2_X1 U2701 ( .A1(n33894), .A2(n6319), .ZN(n5089) );
  NOR2_X1 U2705 ( .A1(n33894), .A2(n6319), .ZN(n32526) );
  CLKBUF_X4 U2706 ( .I(n24471), .Z(n25013) );
  NOR2_X1 U2708 ( .A1(n419), .A2(n25405), .ZN(n25328) );
  NAND2_X1 U2710 ( .A1(n14810), .A2(n6402), .ZN(n25124) );
  NAND3_X1 U2711 ( .A1(n17872), .A2(n5373), .A3(n23901), .ZN(n17995) );
  NAND2_X1 U2713 ( .A1(n17149), .A2(n3898), .ZN(n5136) );
  CLKBUF_X2 U2721 ( .I(n25369), .Z(n30400) );
  NOR2_X1 U2722 ( .A1(n13883), .A2(n13811), .ZN(n25559) );
  BUF_X2 U2724 ( .I(n7925), .Z(n34109) );
  INV_X1 U2730 ( .I(n7925), .ZN(n3646) );
  OAI22_X1 U2731 ( .A1(n6061), .A2(n2697), .B1(n6062), .B2(n16647), .ZN(n33634) );
  NAND2_X1 U2736 ( .A1(n1805), .A2(n16647), .ZN(n6061) );
  NAND2_X1 U2739 ( .A1(n31155), .A2(n30505), .ZN(n31837) );
  NAND2_X1 U2742 ( .A1(n1090), .A2(n31155), .ZN(n10812) );
  BUF_X1 U2743 ( .I(n14531), .Z(n32553) );
  NOR2_X1 U2746 ( .A1(n25632), .A2(n29476), .ZN(n30423) );
  NOR3_X1 U2747 ( .A1(n30396), .A2(n10314), .A3(n14922), .ZN(n26528) );
  OAI21_X1 U2748 ( .A1(n33680), .A2(n33540), .B(n24243), .ZN(n23984) );
  NAND3_X1 U2752 ( .A1(n29495), .A2(n1127), .A3(n22670), .ZN(n33015) );
  INV_X1 U2757 ( .I(n23840), .ZN(n32611) );
  OAI21_X1 U2761 ( .A1(n13242), .A2(n23935), .B(n15097), .ZN(n14704) );
  NAND3_X1 U2763 ( .A1(n13242), .A2(n23575), .A3(n17181), .ZN(n33625) );
  OAI21_X1 U2764 ( .A1(n31959), .A2(n23935), .B(n13242), .ZN(n28530) );
  NAND2_X1 U2765 ( .A1(n31959), .A2(n13242), .ZN(n15803) );
  INV_X1 U2769 ( .I(n4034), .ZN(n1309) );
  NOR2_X1 U2773 ( .A1(n1500), .A2(n24072), .ZN(n1499) );
  BUF_X2 U2774 ( .I(n24072), .Z(n27038) );
  AOI21_X1 U2776 ( .A1(n25858), .A2(n14915), .B(n25854), .ZN(n24737) );
  NAND2_X1 U2777 ( .A1(n25858), .A2(n25859), .ZN(n25857) );
  NAND2_X1 U2779 ( .A1(n13947), .A2(n13946), .ZN(n13945) );
  INV_X1 U2781 ( .I(n11668), .ZN(n29660) );
  NAND3_X1 U2782 ( .A1(n23543), .A2(n23855), .A3(n14193), .ZN(n23547) );
  NAND2_X1 U2785 ( .A1(n5897), .A2(n17382), .ZN(n24984) );
  INV_X1 U2787 ( .I(n17382), .ZN(n13428) );
  NOR2_X1 U2788 ( .A1(n25460), .A2(n25475), .ZN(n32115) );
  CLKBUF_X2 U2789 ( .I(n25107), .Z(n4193) );
  NOR2_X1 U2792 ( .A1(n23857), .A2(n23201), .ZN(n25951) );
  NOR2_X1 U2795 ( .A1(n23201), .A2(n9152), .ZN(n29178) );
  CLKBUF_X2 U2797 ( .I(n25859), .Z(n13049) );
  AND2_X1 U2800 ( .A1(n25513), .A2(n25517), .Z(n25516) );
  OAI21_X1 U2806 ( .A1(n25081), .A2(n30330), .B(n32771), .ZN(n16104) );
  AOI22_X1 U2811 ( .A1(n1949), .A2(n30330), .B1(n1951), .B2(n16810), .ZN(
        n32771) );
  AOI21_X1 U2819 ( .A1(n25923), .A2(n25915), .B(n11019), .ZN(n14432) );
  CLKBUF_X4 U2820 ( .I(n13960), .Z(n11019) );
  NOR2_X1 U2828 ( .A1(n28694), .A2(n24004), .ZN(n5912) );
  OAI21_X1 U2829 ( .A1(n33871), .A2(n33872), .B(n24004), .ZN(n8001) );
  INV_X2 U2832 ( .I(n16273), .ZN(n8929) );
  AOI22_X1 U2834 ( .A1(n8207), .A2(n16273), .B1(n33851), .B2(n25174), .ZN(
        n25180) );
  INV_X1 U2835 ( .I(n3220), .ZN(n24069) );
  AOI21_X1 U2837 ( .A1(n24249), .A2(n24248), .B(n3220), .ZN(n29949) );
  NAND2_X1 U2843 ( .A1(n13223), .A2(n3220), .ZN(n1511) );
  INV_X1 U2844 ( .I(n5043), .ZN(n25211) );
  AOI21_X1 U2851 ( .A1(n1186), .A2(n18701), .B(n31012), .ZN(n13947) );
  NAND3_X1 U2854 ( .A1(n1186), .A2(n34110), .A3(n18701), .ZN(n33412) );
  INV_X2 U2861 ( .I(n18701), .ZN(n13554) );
  OAI22_X1 U2862 ( .A1(n32100), .A2(n25090), .B1(n25094), .B2(n25089), .ZN(
        n32529) );
  CLKBUF_X2 U2863 ( .I(n8678), .Z(n26753) );
  NOR2_X1 U2865 ( .A1(n8678), .A2(n25795), .ZN(n25797) );
  AND2_X1 U2875 ( .A1(n25317), .A2(n25313), .Z(n25320) );
  NAND4_X1 U2877 ( .A1(n693), .A2(n25070), .A3(n25069), .A4(n25068), .ZN(
        n29723) );
  INV_X1 U2878 ( .I(n7198), .ZN(n747) );
  OAI21_X1 U2881 ( .A1(n32270), .A2(n34170), .B(n24897), .ZN(n33081) );
  CLKBUF_X2 U2882 ( .I(n16940), .Z(n4024) );
  INV_X1 U2884 ( .I(n16940), .ZN(n24311) );
  NAND3_X1 U2886 ( .A1(n25744), .A2(n25739), .A3(n4415), .ZN(n32279) );
  INV_X1 U2887 ( .I(n1506), .ZN(n8235) );
  NAND2_X1 U2888 ( .A1(n4778), .A2(n4776), .ZN(n3589) );
  NOR3_X1 U2890 ( .A1(n8258), .A2(n16377), .A3(n8257), .ZN(n28486) );
  OR2_X1 U2891 ( .A1(n25473), .A2(n30047), .Z(n25460) );
  INV_X2 U2893 ( .I(n30584), .ZN(n16501) );
  NAND2_X1 U2895 ( .A1(n3909), .A2(n30584), .ZN(n22744) );
  NOR2_X1 U2904 ( .A1(n22953), .A2(n30584), .ZN(n22327) );
  NAND2_X1 U2911 ( .A1(n11105), .A2(n20591), .ZN(n11104) );
  NAND2_X1 U2912 ( .A1(n11255), .A2(n24327), .ZN(n9823) );
  NAND3_X1 U2913 ( .A1(n32510), .A2(n22855), .A3(n25979), .ZN(n22859) );
  NOR2_X1 U2914 ( .A1(n22709), .A2(n25979), .ZN(n14162) );
  NAND3_X1 U2927 ( .A1(n25979), .A2(n33132), .A3(n30365), .ZN(n22857) );
  AOI21_X1 U2931 ( .A1(n2480), .A2(n749), .B(n32177), .ZN(n25504) );
  CLKBUF_X2 U2932 ( .I(n6595), .Z(n2480) );
  NAND2_X1 U2937 ( .A1(n28427), .A2(n12471), .ZN(n10361) );
  NAND2_X1 U2940 ( .A1(n18084), .A2(n26390), .ZN(n24709) );
  NOR2_X1 U2941 ( .A1(n26390), .A2(n24310), .ZN(n9016) );
  NAND2_X1 U2942 ( .A1(n16609), .A2(n718), .ZN(n25583) );
  INV_X1 U2943 ( .I(n16609), .ZN(n13642) );
  NAND3_X1 U2946 ( .A1(n27113), .A2(n6092), .A3(n5926), .ZN(n36) );
  CLKBUF_X4 U2947 ( .I(n5492), .Z(n964) );
  NAND2_X1 U2949 ( .A1(n13488), .A2(n19867), .ZN(n28130) );
  NOR2_X1 U2952 ( .A1(n16271), .A2(n33679), .ZN(n33870) );
  NAND2_X1 U2956 ( .A1(n5091), .A2(n5292), .ZN(n24728) );
  INV_X1 U2957 ( .I(n10644), .ZN(n23064) );
  NOR2_X1 U2962 ( .A1(n714), .A2(n25006), .ZN(n15079) );
  NOR2_X1 U2963 ( .A1(n16519), .A2(n21662), .ZN(n13213) );
  NOR2_X1 U2966 ( .A1(n16519), .A2(n32898), .ZN(n14730) );
  NAND3_X1 U2968 ( .A1(n777), .A2(n21662), .A3(n16519), .ZN(n27760) );
  AOI21_X1 U2972 ( .A1(n7068), .A2(n24196), .B(n28784), .ZN(n2921) );
  NAND2_X1 U2973 ( .A1(n25724), .A2(n16494), .ZN(n25717) );
  OR2_X1 U2974 ( .A1(n675), .A2(n24779), .Z(n2727) );
  CLKBUF_X2 U2982 ( .I(n7940), .Z(n3376) );
  NAND2_X1 U2984 ( .A1(n25882), .A2(n5410), .ZN(n33176) );
  CLKBUF_X2 U2994 ( .I(n17824), .Z(n30396) );
  AOI21_X1 U2995 ( .A1(n14922), .A2(n17824), .B(n6034), .ZN(n16169) );
  NAND2_X1 U2997 ( .A1(n7515), .A2(n25221), .ZN(n15462) );
  INV_X1 U2998 ( .I(n25221), .ZN(n966) );
  NAND2_X1 U3000 ( .A1(n15421), .A2(n22832), .ZN(n23002) );
  OAI21_X1 U3001 ( .A1(n22752), .A2(n15421), .B(n16817), .ZN(n22618) );
  AND2_X1 U3003 ( .A1(n14873), .A2(n33155), .Z(n32030) );
  NOR2_X1 U3007 ( .A1(n13296), .A2(n13822), .ZN(n33516) );
  OAI21_X1 U3011 ( .A1(n10206), .A2(n28263), .B(n6709), .ZN(n6711) );
  OAI21_X1 U3014 ( .A1(n22583), .A2(n10206), .B(n28263), .ZN(n10796) );
  NAND2_X1 U3015 ( .A1(n33392), .A2(n6661), .ZN(n30185) );
  NAND2_X1 U3016 ( .A1(n16292), .A2(n23759), .ZN(n33392) );
  NAND2_X1 U3018 ( .A1(n31323), .A2(n32144), .ZN(n32272) );
  AOI22_X1 U3023 ( .A1(n25552), .A2(n13483), .B1(n33414), .B2(n13811), .ZN(
        n32144) );
  OAI21_X1 U3024 ( .A1(n16835), .A2(n700), .B(n25900), .ZN(n10756) );
  NAND3_X1 U3033 ( .A1(n13366), .A2(n8657), .A3(n13367), .ZN(n31734) );
  NAND2_X1 U3042 ( .A1(n7831), .A2(n24995), .ZN(n14208) );
  BUF_X2 U3046 ( .I(n14058), .Z(n27750) );
  NAND2_X1 U3047 ( .A1(n31907), .A2(n20507), .ZN(n14683) );
  AND2_X1 U3049 ( .A1(n3944), .A2(n31907), .Z(n16123) );
  INV_X1 U3051 ( .I(n31907), .ZN(n14369) );
  INV_X1 U3054 ( .I(n23456), .ZN(n30843) );
  BUF_X2 U3059 ( .I(n23456), .Z(n27481) );
  INV_X1 U3061 ( .I(n15425), .ZN(n25865) );
  INV_X1 U3062 ( .I(n21012), .ZN(n30487) );
  NAND2_X1 U3063 ( .A1(n22772), .A2(n1106), .ZN(n22773) );
  AND2_X1 U3066 ( .A1(n24171), .A2(n3483), .Z(n32041) );
  NAND2_X1 U3067 ( .A1(n34149), .A2(n834), .ZN(n12386) );
  INV_X1 U3068 ( .I(n834), .ZN(n32591) );
  CLKBUF_X2 U3070 ( .I(n18911), .Z(n33698) );
  NAND3_X1 U3071 ( .A1(n34074), .A2(n29395), .A3(n22682), .ZN(n3894) );
  NAND2_X1 U3072 ( .A1(n22772), .A2(n28957), .ZN(n22751) );
  NAND2_X1 U3073 ( .A1(n3300), .A2(n25375), .ZN(n25366) );
  NOR2_X1 U3074 ( .A1(n25376), .A2(n25375), .ZN(n14102) );
  NAND2_X1 U3075 ( .A1(n21840), .A2(n16987), .ZN(n21749) );
  NOR2_X1 U3080 ( .A1(n32063), .A2(n24955), .ZN(n24948) );
  CLKBUF_X4 U3081 ( .I(n24174), .Z(n25900) );
  NAND2_X1 U3084 ( .A1(n11899), .A2(n8307), .ZN(n24710) );
  OAI21_X1 U3085 ( .A1(n696), .A2(n1212), .B(n11899), .ZN(n4709) );
  NOR2_X1 U3092 ( .A1(n1202), .A2(n9982), .ZN(n12049) );
  INV_X1 U3093 ( .I(n32906), .ZN(n23152) );
  AOI22_X1 U3094 ( .A1(n33176), .A2(n14737), .B1(n5407), .B2(n32059), .ZN(
        n13902) );
  AND2_X1 U3096 ( .A1(n16033), .A2(n17661), .Z(n1933) );
  NAND2_X1 U3097 ( .A1(n1100), .A2(n16033), .ZN(n7781) );
  INV_X1 U3099 ( .I(n535), .ZN(n16033) );
  INV_X1 U3104 ( .I(n16853), .ZN(n28759) );
  NAND2_X1 U3106 ( .A1(n5259), .A2(n12450), .ZN(n12449) );
  INV_X1 U3107 ( .I(n23334), .ZN(n31567) );
  NAND2_X1 U3109 ( .A1(n30033), .A2(n8875), .ZN(n21740) );
  CLKBUF_X4 U3110 ( .I(n24408), .Z(n25756) );
  NOR2_X1 U3121 ( .A1(n22546), .A2(n22550), .ZN(n27406) );
  OAI21_X1 U3122 ( .A1(n22546), .A2(n27402), .B(n22550), .ZN(n26855) );
  NOR3_X1 U3123 ( .A1(n22546), .A2(n22549), .A3(n22547), .ZN(n32943) );
  INV_X1 U3128 ( .I(n24275), .ZN(n24196) );
  NOR2_X1 U3130 ( .A1(n30129), .A2(n33766), .ZN(n16229) );
  OAI21_X1 U3134 ( .A1(n912), .A2(n33766), .B(n1137), .ZN(n2718) );
  NAND2_X1 U3136 ( .A1(n33766), .A2(n2368), .ZN(n33841) );
  AOI21_X1 U3137 ( .A1(n912), .A2(n33766), .B(n38), .ZN(n16231) );
  NAND2_X1 U3142 ( .A1(n25141), .A2(n25145), .ZN(n2642) );
  CLKBUF_X2 U3143 ( .I(n25141), .Z(n16276) );
  INV_X1 U3151 ( .I(n25141), .ZN(n17987) );
  NAND2_X1 U3154 ( .A1(n31915), .A2(n11850), .ZN(n10470) );
  CLKBUF_X2 U3158 ( .I(n3874), .Z(n29839) );
  NAND2_X1 U3159 ( .A1(n27670), .A2(n22653), .ZN(n3951) );
  AOI22_X1 U3163 ( .A1(n16560), .A2(n22826), .B1(n23066), .B2(n7881), .ZN(
        n22653) );
  NAND2_X1 U3164 ( .A1(n23064), .A2(n28689), .ZN(n27670) );
  INV_X2 U3165 ( .I(n19907), .ZN(n20112) );
  NAND2_X1 U3166 ( .A1(n16058), .A2(n21396), .ZN(n27432) );
  NOR2_X1 U3168 ( .A1(n12325), .A2(n21396), .ZN(n12324) );
  NOR3_X1 U3171 ( .A1(n21396), .A2(n27955), .A3(n21400), .ZN(n32393) );
  NAND2_X1 U3174 ( .A1(n15746), .A2(n16205), .ZN(n3598) );
  NAND2_X1 U3185 ( .A1(n22690), .A2(n15746), .ZN(n32191) );
  NOR2_X1 U3194 ( .A1(n22690), .A2(n15746), .ZN(n30436) );
  NAND2_X1 U3201 ( .A1(n15746), .A2(n30333), .ZN(n31126) );
  NOR2_X1 U3202 ( .A1(n25967), .A2(n10700), .ZN(n15804) );
  NOR2_X1 U3205 ( .A1(n32186), .A2(n7188), .ZN(n9788) );
  NOR2_X1 U3206 ( .A1(n3165), .A2(n32186), .ZN(n34012) );
  INV_X1 U3207 ( .I(n12648), .ZN(n32785) );
  CLKBUF_X2 U3209 ( .I(n9107), .Z(n26739) );
  OR2_X1 U3211 ( .A1(n4184), .A2(n13191), .Z(n31052) );
  NAND2_X1 U3212 ( .A1(n4184), .A2(n13191), .ZN(n13995) );
  AND2_X1 U3213 ( .A1(n2635), .A2(n4184), .Z(n8290) );
  CLKBUF_X2 U3214 ( .I(n9708), .Z(n29318) );
  CLKBUF_X2 U3216 ( .I(n16331), .Z(n8347) );
  BUF_X2 U3217 ( .I(n21071), .Z(n21426) );
  OR2_X1 U3218 ( .A1(n17670), .A2(n5433), .Z(n29357) );
  NAND2_X1 U3219 ( .A1(n7081), .A2(n25232), .ZN(n10570) );
  OR2_X1 U3220 ( .A1(n339), .A2(n31217), .Z(n18344) );
  NOR2_X1 U3224 ( .A1(n32401), .A2(n339), .ZN(n9839) );
  INV_X2 U3228 ( .I(n339), .ZN(n19052) );
  AOI21_X1 U3229 ( .A1(n32401), .A2(n339), .B(n10015), .ZN(n2148) );
  OAI21_X1 U3230 ( .A1(n339), .A2(n10015), .B(n10017), .ZN(n31226) );
  OR3_X2 U3231 ( .A1(n989), .A2(n12578), .A3(n13648), .Z(n12577) );
  INV_X1 U3232 ( .I(n33857), .ZN(n33519) );
  NAND2_X1 U3236 ( .A1(n18830), .A2(n16915), .ZN(n3893) );
  AOI21_X1 U3239 ( .A1(n18830), .A2(n9), .B(n18829), .ZN(n29808) );
  INV_X1 U3244 ( .I(n3079), .ZN(n32565) );
  NAND2_X1 U3245 ( .A1(n10724), .A2(n906), .ZN(n4315) );
  AOI22_X1 U3246 ( .A1(n22643), .A2(n30448), .B1(n6297), .B2(n10724), .ZN(
        n13461) );
  INV_X1 U3247 ( .I(n19470), .ZN(n19561) );
  AND2_X1 U3249 ( .A1(n11515), .A2(n30713), .Z(n31180) );
  OAI21_X1 U3255 ( .A1(n867), .A2(n1469), .B(n20442), .ZN(n30929) );
  NAND2_X1 U3260 ( .A1(n19932), .A2(n8817), .ZN(n1812) );
  NAND2_X1 U3268 ( .A1(n11903), .A2(n2166), .ZN(n2167) );
  NAND2_X1 U3270 ( .A1(n2166), .A2(n28645), .ZN(n28022) );
  OAI21_X1 U3272 ( .A1(n2166), .A2(n20069), .B(n27715), .ZN(n6926) );
  INV_X1 U3276 ( .I(n32124), .ZN(n297) );
  BUF_X2 U3282 ( .I(Key[57]), .Z(n25856) );
  NOR2_X1 U3285 ( .A1(n5098), .A2(n24111), .ZN(n10178) );
  NAND2_X1 U3286 ( .A1(n13896), .A2(n16072), .ZN(n14074) );
  OAI22_X1 U3288 ( .A1(n4989), .A2(n4324), .B1(n13896), .B2(n32799), .ZN(
        n30654) );
  CLKBUF_X4 U3289 ( .I(n24866), .Z(n24667) );
  OAI22_X1 U3292 ( .A1(n803), .A2(n27450), .B1(n23158), .B2(n14183), .ZN(
        n27372) );
  OAI21_X1 U3295 ( .A1(n3379), .A2(n11756), .B(n31197), .ZN(n13034) );
  NAND2_X1 U3300 ( .A1(n31197), .A2(n28099), .ZN(n21664) );
  OAI21_X1 U3303 ( .A1(n15038), .A2(n16099), .B(n31479), .ZN(n5040) );
  BUF_X2 U3306 ( .I(n8926), .Z(n8207) );
  NOR2_X1 U3310 ( .A1(n25154), .A2(n8926), .ZN(n25158) );
  INV_X1 U3314 ( .I(n8926), .ZN(n25165) );
  NAND3_X1 U3317 ( .A1(n15423), .A2(n23848), .A3(n26114), .ZN(n6129) );
  INV_X1 U3318 ( .I(n30305), .ZN(n19416) );
  INV_X1 U3320 ( .I(n24573), .ZN(n11652) );
  NAND3_X1 U3323 ( .A1(n24573), .A2(n14410), .A3(n14412), .ZN(n8988) );
  CLKBUF_X2 U3324 ( .I(n21569), .Z(n29806) );
  INV_X1 U3327 ( .I(n21569), .ZN(n32506) );
  NAND2_X1 U3330 ( .A1(n3203), .A2(n21569), .ZN(n21491) );
  CLKBUF_X2 U3333 ( .I(n8622), .Z(n33434) );
  NAND3_X1 U3335 ( .A1(n21865), .A2(n30154), .A3(n28018), .ZN(n21739) );
  AOI22_X1 U3339 ( .A1(n26766), .A2(n8457), .B1(n21865), .B2(n21867), .ZN(
        n4516) );
  NAND2_X1 U3350 ( .A1(n21865), .A2(n21866), .ZN(n16241) );
  NAND2_X1 U3352 ( .A1(n32833), .A2(n21865), .ZN(n31711) );
  NOR2_X1 U3353 ( .A1(n21865), .A2(n21866), .ZN(n31334) );
  INV_X2 U3355 ( .I(n21865), .ZN(n15465) );
  CLKBUF_X2 U3356 ( .I(n22363), .Z(n6478) );
  CLKBUF_X4 U3357 ( .I(n16052), .Z(n5631) );
  INV_X2 U3358 ( .I(n16052), .ZN(n5632) );
  NAND3_X1 U3364 ( .A1(n4873), .A2(n23934), .A3(n11200), .ZN(n4872) );
  NOR3_X1 U3366 ( .A1(n33425), .A2(n28945), .A3(n11200), .ZN(n32929) );
  NAND3_X1 U3367 ( .A1(n27450), .A2(n32868), .A3(n803), .ZN(n13914) );
  NOR2_X1 U3372 ( .A1(n23051), .A2(n28277), .ZN(n17482) );
  NOR2_X1 U3378 ( .A1(n28277), .A2(n23051), .ZN(n16054) );
  CLKBUF_X4 U3381 ( .I(n19418), .Z(n19884) );
  NOR2_X1 U3383 ( .A1(n19418), .A2(n19885), .ZN(n13488) );
  CLKBUF_X4 U3384 ( .I(n2600), .Z(n29330) );
  INV_X1 U3388 ( .I(n5268), .ZN(n3146) );
  NOR3_X1 U3397 ( .A1(n29634), .A2(n14619), .A3(n24154), .ZN(n5613) );
  NOR2_X1 U3399 ( .A1(n9062), .A2(n31471), .ZN(n14568) );
  NAND2_X1 U3407 ( .A1(n9062), .A2(n20630), .ZN(n31469) );
  NOR3_X1 U3408 ( .A1(n5335), .A2(n24148), .A3(n3748), .ZN(n8543) );
  CLKBUF_X4 U3409 ( .I(n29279), .Z(n33585) );
  NAND2_X1 U3413 ( .A1(n25755), .A2(n29279), .ZN(n32343) );
  NAND2_X1 U3415 ( .A1(n31079), .A2(n30504), .ZN(n30503) );
  NAND2_X1 U3418 ( .A1(n15314), .A2(n15316), .ZN(n30284) );
  NOR2_X1 U3420 ( .A1(n23849), .A2(n26114), .ZN(n23808) );
  AOI22_X1 U3421 ( .A1(n12996), .A2(n100), .B1(n19057), .B2(n19058), .ZN(
        n19059) );
  NAND2_X1 U3425 ( .A1(n6718), .A2(n21719), .ZN(n14717) );
  NAND2_X1 U3427 ( .A1(n12221), .A2(n6718), .ZN(n21741) );
  INV_X1 U3429 ( .I(n6718), .ZN(n33083) );
  NAND2_X1 U3431 ( .A1(n17227), .A2(n6718), .ZN(n3420) );
  OR2_X1 U3444 ( .A1(n13913), .A2(n29815), .Z(n5223) );
  NAND2_X1 U3452 ( .A1(n24960), .A2(n24896), .ZN(n24939) );
  NOR2_X1 U3456 ( .A1(n8420), .A2(n29287), .ZN(n22683) );
  INV_X1 U3458 ( .I(n8420), .ZN(n2418) );
  NAND2_X1 U3459 ( .A1(n25012), .A2(n25015), .ZN(n24591) );
  NOR2_X1 U3466 ( .A1(n30145), .A2(n25015), .ZN(n33757) );
  NOR2_X1 U3469 ( .A1(n25015), .A2(n17240), .ZN(n12093) );
  INV_X2 U3471 ( .I(n24975), .ZN(n25015) );
  NOR2_X1 U3472 ( .A1(n33648), .A2(n29387), .ZN(n26389) );
  AOI21_X1 U3473 ( .A1(n12657), .A2(n20066), .B(n19874), .ZN(n19798) );
  AOI21_X1 U3476 ( .A1(n14976), .A2(n12657), .B(n20066), .ZN(n29905) );
  INV_X1 U3478 ( .I(n29258), .ZN(n17053) );
  INV_X1 U3482 ( .I(n3147), .ZN(n11768) );
  BUF_X2 U3484 ( .I(n3147), .Z(n31228) );
  NAND2_X1 U3491 ( .A1(n21072), .A2(n21428), .ZN(n2241) );
  NAND2_X1 U3495 ( .A1(n20009), .A2(n20008), .ZN(n20085) );
  NAND3_X1 U3496 ( .A1(n20009), .A2(n8301), .A3(n20008), .ZN(n9338) );
  OR3_X2 U3499 ( .A1(n20009), .A2(n20083), .A3(n11068), .Z(n9339) );
  CLKBUF_X2 U3501 ( .I(n22457), .Z(n16503) );
  INV_X2 U3505 ( .I(n12535), .ZN(n26513) );
  INV_X1 U3506 ( .I(n12548), .ZN(n18978) );
  NOR2_X1 U3511 ( .A1(n16916), .A2(n12548), .ZN(n6639) );
  NAND2_X1 U3516 ( .A1(n12548), .A2(n14812), .ZN(n19113) );
  CLKBUF_X1 U3521 ( .I(n17408), .Z(n27984) );
  CLKBUF_X2 U3523 ( .I(n13694), .Z(n27450) );
  NAND2_X1 U3524 ( .A1(n1177), .A2(n32332), .ZN(n32331) );
  INV_X2 U3530 ( .I(n1177), .ZN(n32671) );
  AOI21_X1 U3534 ( .A1(n19324), .A2(n19274), .B(n1177), .ZN(n19278) );
  OAI21_X1 U3537 ( .A1(n29965), .A2(n23912), .B(n23588), .ZN(n16539) );
  OAI21_X1 U3542 ( .A1(n16496), .A2(n34167), .B(n29965), .ZN(n28061) );
  NAND2_X1 U3545 ( .A1(n16496), .A2(n29965), .ZN(n26224) );
  INV_X2 U3546 ( .I(n20523), .ZN(n17790) );
  NAND2_X1 U3552 ( .A1(n30454), .A2(n20523), .ZN(n28484) );
  NOR2_X1 U3555 ( .A1(n16684), .A2(n20523), .ZN(n20280) );
  OAI21_X1 U3556 ( .A1(n16459), .A2(n31195), .B(n31498), .ZN(n2687) );
  OAI21_X1 U3558 ( .A1(n16459), .A2(n926), .B(n21077), .ZN(n12506) );
  NAND2_X1 U3561 ( .A1(n33523), .A2(n16459), .ZN(n2569) );
  BUF_X2 U3562 ( .I(n16248), .Z(n28904) );
  INV_X1 U3568 ( .I(n16248), .ZN(n26182) );
  BUF_X2 U3575 ( .I(n18064), .Z(n29216) );
  NAND2_X1 U3576 ( .A1(n18064), .A2(n34122), .ZN(n33570) );
  INV_X1 U3580 ( .I(n18064), .ZN(n1035) );
  OR2_X1 U3591 ( .A1(n10514), .A2(n18064), .Z(n29022) );
  CLKBUF_X1 U3595 ( .I(n16215), .Z(n10651) );
  INV_X1 U3596 ( .I(n16215), .ZN(n29883) );
  AND2_X1 U3599 ( .A1(n7935), .A2(n16215), .Z(n9368) );
  NOR2_X1 U3600 ( .A1(n16389), .A2(n28578), .ZN(n18671) );
  NOR3_X1 U3601 ( .A1(n16466), .A2(n16572), .A3(n16389), .ZN(n10638) );
  NAND2_X1 U3608 ( .A1(n31437), .A2(n23057), .ZN(n2877) );
  INV_X2 U3615 ( .I(n14359), .ZN(n1206) );
  NAND2_X1 U3619 ( .A1(n14359), .A2(n7702), .ZN(n25912) );
  CLKBUF_X2 U3621 ( .I(n24447), .Z(n16413) );
  NAND2_X1 U3622 ( .A1(n15116), .A2(n23742), .ZN(n23583) );
  OAI21_X1 U3630 ( .A1(n20460), .A2(n7852), .B(n7292), .ZN(n31898) );
  BUF_X2 U3631 ( .I(n7852), .Z(n8031) );
  INV_X1 U3636 ( .I(n16175), .ZN(n14968) );
  OAI21_X1 U3640 ( .A1(n34115), .A2(n1216), .B(n1083), .ZN(n8120) );
  NOR2_X1 U3653 ( .A1(n25234), .A2(n1083), .ZN(n3731) );
  INV_X2 U3655 ( .I(n34167), .ZN(n14463) );
  AOI21_X1 U3658 ( .A1(n2507), .A2(n10283), .B(n32409), .ZN(n32541) );
  INV_X1 U3664 ( .I(n19967), .ZN(n14334) );
  CLKBUF_X2 U3668 ( .I(n19967), .Z(n16092) );
  INV_X1 U3677 ( .I(n16562), .ZN(n32568) );
  NOR2_X1 U3690 ( .A1(n32483), .A2(n16562), .ZN(n2409) );
  INV_X1 U3691 ( .I(n16646), .ZN(n19834) );
  NAND2_X1 U3698 ( .A1(n19151), .A2(n11072), .ZN(n2152) );
  NOR2_X1 U3702 ( .A1(n6976), .A2(n5379), .ZN(n30718) );
  NAND2_X1 U3706 ( .A1(n6976), .A2(n5379), .ZN(n2381) );
  NOR3_X1 U3712 ( .A1(n2744), .A2(n24317), .A3(n26938), .ZN(n33512) );
  NAND2_X1 U3719 ( .A1(n26938), .A2(n13232), .ZN(n14663) );
  NAND2_X1 U3724 ( .A1(n26938), .A2(n32298), .ZN(n2993) );
  AOI22_X1 U3737 ( .A1(n24318), .A2(n26938), .B1(n2744), .B2(n24317), .ZN(
        n24319) );
  NAND2_X1 U3740 ( .A1(n6457), .A2(n11941), .ZN(n3113) );
  INV_X2 U3745 ( .I(n11941), .ZN(n16318) );
  NOR2_X1 U3748 ( .A1(n33834), .A2(n14419), .ZN(n29817) );
  INV_X1 U3749 ( .I(n7345), .ZN(n945) );
  NAND2_X1 U3751 ( .A1(n21627), .A2(n14095), .ZN(n14153) );
  NOR2_X1 U3752 ( .A1(n29322), .A2(n14095), .ZN(n33459) );
  NOR2_X1 U3756 ( .A1(n13773), .A2(n16333), .ZN(n9714) );
  OAI21_X1 U3757 ( .A1(n23881), .A2(n13773), .B(n23882), .ZN(n7170) );
  AOI22_X1 U3758 ( .A1(n9714), .A2(n23787), .B1(n10619), .B2(n13773), .ZN(
        n32942) );
  INV_X2 U3760 ( .I(n13773), .ZN(n16320) );
  NAND2_X1 U3763 ( .A1(n5915), .A2(n5696), .ZN(n28970) );
  INV_X2 U3765 ( .I(n14365), .ZN(n1355) );
  NOR2_X1 U3766 ( .A1(n14365), .A2(n31907), .ZN(n20435) );
  INV_X1 U3767 ( .I(n8625), .ZN(n13286) );
  INV_X1 U3770 ( .I(n20518), .ZN(n932) );
  CLKBUF_X2 U3774 ( .I(n20518), .Z(n6530) );
  BUF_X2 U3776 ( .I(n21198), .Z(n13896) );
  NOR2_X1 U3777 ( .A1(n31161), .A2(n8100), .ZN(n12297) );
  NOR2_X1 U3784 ( .A1(n4359), .A2(n4356), .ZN(n33746) );
  OAI21_X1 U3785 ( .A1(n21855), .A2(n12229), .B(n4356), .ZN(n33664) );
  NAND2_X1 U3786 ( .A1(n32642), .A2(n4356), .ZN(n21823) );
  OAI21_X1 U3788 ( .A1(n21853), .A2(n4356), .B(n5546), .ZN(n17748) );
  NAND2_X1 U3791 ( .A1(n4184), .A2(n13558), .ZN(n23107) );
  INV_X1 U3793 ( .I(n13558), .ZN(n2713) );
  NAND2_X1 U3796 ( .A1(n14131), .A2(n13558), .ZN(n13386) );
  CLKBUF_X2 U3798 ( .I(n22127), .Z(n28709) );
  INV_X1 U3808 ( .I(n22127), .ZN(n26193) );
  NAND2_X1 U3816 ( .A1(n16743), .A2(n16938), .ZN(n33423) );
  NAND2_X1 U3818 ( .A1(n10665), .A2(n18071), .ZN(n18254) );
  OAI21_X1 U3824 ( .A1(n17316), .A2(n34139), .B(n33687), .ZN(n12151) );
  AND2_X1 U3825 ( .A1(n23862), .A2(n26290), .Z(n9261) );
  NAND2_X1 U3829 ( .A1(n23862), .A2(n23864), .ZN(n33724) );
  INV_X1 U3831 ( .I(n15715), .ZN(n20377) );
  NOR2_X1 U3835 ( .A1(n14179), .A2(n15715), .ZN(n9719) );
  OAI21_X1 U3836 ( .A1(n1291), .A2(n26708), .B(n15853), .ZN(n7427) );
  OAI21_X1 U3842 ( .A1(n26173), .A2(n26708), .B(n29336), .ZN(n33105) );
  NOR2_X1 U3845 ( .A1(n26708), .A2(n26709), .ZN(n34002) );
  NAND2_X1 U3846 ( .A1(n22608), .A2(n26708), .ZN(n32450) );
  INV_X2 U3850 ( .I(n32605), .ZN(n26708) );
  BUF_X2 U3856 ( .I(n9292), .Z(n4975) );
  INV_X1 U3860 ( .I(n14821), .ZN(n20236) );
  BUF_X2 U3861 ( .I(n14821), .Z(n7486) );
  INV_X1 U3862 ( .I(n19679), .ZN(n17129) );
  NAND2_X1 U3868 ( .A1(n5318), .A2(n29634), .ZN(n16985) );
  CLKBUF_X2 U3870 ( .I(n5318), .Z(n28833) );
  CLKBUF_X4 U3871 ( .I(n20521), .Z(n16218) );
  NAND3_X1 U3873 ( .A1(n15096), .A2(n737), .A3(n27038), .ZN(n1837) );
  NAND2_X1 U3878 ( .A1(n33019), .A2(n15096), .ZN(n1496) );
  NAND3_X1 U3879 ( .A1(n15096), .A2(n13334), .A3(n27184), .ZN(n5129) );
  NAND2_X1 U3882 ( .A1(n25757), .A2(n26056), .ZN(n30259) );
  INV_X1 U3888 ( .I(n14682), .ZN(n2649) );
  INV_X1 U3896 ( .I(n9287), .ZN(n20628) );
  CLKBUF_X4 U3903 ( .I(n9287), .Z(n9014) );
  INV_X1 U3906 ( .I(n2859), .ZN(n31835) );
  BUF_X2 U3907 ( .I(n2859), .Z(n2738) );
  NAND3_X1 U3908 ( .A1(n5452), .A2(n4547), .A3(n16567), .ZN(n31418) );
  OAI22_X1 U3910 ( .A1(n5452), .A2(n6658), .B1(n22578), .B2(n29021), .ZN(n5449) );
  AOI21_X1 U3912 ( .A1(n5452), .A2(n22666), .B(n22576), .ZN(n5451) );
  CLKBUF_X4 U3916 ( .I(n22156), .Z(n22664) );
  INV_X1 U3920 ( .I(n23899), .ZN(n28914) );
  NAND2_X1 U3924 ( .A1(n6985), .A2(n1577), .ZN(n30945) );
  NOR2_X1 U3925 ( .A1(n12593), .A2(n7778), .ZN(n24293) );
  CLKBUF_X2 U3926 ( .I(n12593), .Z(n26544) );
  NAND2_X1 U3927 ( .A1(n12593), .A2(n7778), .ZN(n32444) );
  INV_X1 U3929 ( .I(n4897), .ZN(n15065) );
  NAND2_X1 U3930 ( .A1(n15720), .A2(n4897), .ZN(n15996) );
  NAND2_X1 U3932 ( .A1(n23738), .A2(n23737), .ZN(n23739) );
  INV_X1 U3936 ( .I(n21442), .ZN(n6277) );
  INV_X1 U3938 ( .I(n23429), .ZN(n29970) );
  NOR2_X1 U3943 ( .A1(n27726), .A2(n745), .ZN(n19287) );
  NAND2_X1 U3945 ( .A1(n19288), .A2(n745), .ZN(n9356) );
  INV_X1 U3951 ( .I(n19275), .ZN(n19320) );
  NAND2_X1 U3954 ( .A1(n19275), .A2(n19318), .ZN(n33108) );
  NAND2_X1 U3955 ( .A1(n27132), .A2(n19275), .ZN(n18419) );
  NAND3_X1 U3957 ( .A1(n808), .A2(n896), .A3(n22399), .ZN(n15578) );
  NAND2_X1 U3958 ( .A1(n32856), .A2(n25615), .ZN(n28791) );
  NOR2_X1 U3961 ( .A1(n5817), .A2(n30687), .ZN(n30990) );
  NAND2_X1 U3963 ( .A1(n2826), .A2(n24164), .ZN(n17280) );
  NOR2_X1 U3966 ( .A1(n14840), .A2(n2826), .ZN(n14839) );
  NAND2_X1 U3972 ( .A1(n4846), .A2(n4847), .ZN(n32480) );
  NAND2_X1 U3974 ( .A1(n12044), .A2(n27143), .ZN(n21297) );
  CLKBUF_X4 U3977 ( .I(n12044), .Z(n4324) );
  AND3_X1 U3979 ( .A1(n21115), .A2(n12044), .A3(n21405), .Z(n15466) );
  NOR2_X1 U3986 ( .A1(n24221), .A2(n5306), .ZN(n33935) );
  NOR3_X1 U3987 ( .A1(n27077), .A2(n30010), .A3(n5789), .ZN(n26164) );
  AND2_X1 U3991 ( .A1(n29763), .A2(n8374), .Z(n29453) );
  NOR2_X1 U3994 ( .A1(n8374), .A2(n29763), .ZN(n12541) );
  CLKBUF_X2 U3995 ( .I(n26724), .Z(n30573) );
  INV_X2 U3998 ( .I(n22816), .ZN(n23093) );
  NAND2_X1 U3999 ( .A1(n22816), .A2(n27419), .ZN(n12511) );
  NAND2_X1 U4000 ( .A1(n14686), .A2(n22816), .ZN(n22697) );
  INV_X1 U4002 ( .I(n14402), .ZN(n32500) );
  BUF_X2 U4003 ( .I(n14402), .Z(n29107) );
  INV_X2 U4007 ( .I(n22585), .ZN(n1290) );
  NAND2_X1 U4008 ( .A1(n6478), .A2(n22585), .ZN(n7239) );
  BUF_X2 U4009 ( .I(n22585), .Z(n32483) );
  CLKBUF_X2 U4010 ( .I(n7093), .Z(n33990) );
  CLKBUF_X1 U4011 ( .I(n13586), .Z(n33927) );
  NOR2_X1 U4013 ( .A1(n17872), .A2(n14756), .ZN(n7406) );
  INV_X2 U4017 ( .I(n20945), .ZN(n810) );
  NOR2_X1 U4018 ( .A1(n29240), .A2(n23713), .ZN(n32210) );
  NOR2_X1 U4026 ( .A1(n17234), .A2(n23713), .ZN(n31696) );
  NAND2_X1 U4027 ( .A1(n16615), .A2(n23735), .ZN(n23738) );
  OAI21_X1 U4028 ( .A1(n1489), .A2(n16121), .B(n16615), .ZN(n32931) );
  NOR2_X1 U4031 ( .A1(n16615), .A2(n23735), .ZN(n23351) );
  INV_X1 U4040 ( .I(n25119), .ZN(n24884) );
  OR3_X1 U4042 ( .A1(n25119), .A2(n18154), .A3(n27651), .Z(n25021) );
  NOR2_X1 U4047 ( .A1(n17879), .A2(n7965), .ZN(n13143) );
  NAND2_X1 U4054 ( .A1(n33032), .A2(n22791), .ZN(n15390) );
  NAND2_X1 U4057 ( .A1(n14770), .A2(n7188), .ZN(n2070) );
  AOI21_X1 U4061 ( .A1(n23621), .A2(n13176), .B(n15977), .ZN(n23622) );
  NOR2_X1 U4062 ( .A1(n13330), .A2(n947), .ZN(n14649) );
  NAND3_X1 U4067 ( .A1(n16485), .A2(n13330), .A3(n13328), .ZN(n13791) );
  INV_X1 U4068 ( .I(n13330), .ZN(n17508) );
  NOR2_X1 U4069 ( .A1(n13100), .A2(n17039), .ZN(n9967) );
  CLKBUF_X2 U4075 ( .I(n33986), .Z(n33822) );
  NOR2_X1 U4081 ( .A1(n1056), .A2(n33986), .ZN(n32218) );
  BUF_X2 U4082 ( .I(n1808), .Z(n1634) );
  CLKBUF_X2 U4084 ( .I(n1808), .Z(n32515) );
  OAI21_X1 U4086 ( .A1(n1808), .A2(n32102), .B(n16535), .ZN(n2427) );
  CLKBUF_X2 U4087 ( .I(n5863), .Z(n27596) );
  NOR2_X1 U4088 ( .A1(n26169), .A2(n30231), .ZN(n32233) );
  AND2_X1 U4091 ( .A1(n7463), .A2(n30231), .Z(n5821) );
  NOR2_X1 U4092 ( .A1(n30643), .A2(n27105), .ZN(n16176) );
  NAND2_X1 U4095 ( .A1(n24275), .A2(n2654), .ZN(n7067) );
  CLKBUF_X12 U4096 ( .I(n15077), .Z(n8576) );
  XOR2_X1 U4103 ( .A1(n10576), .A2(n17650), .Z(n31922) );
  OR2_X2 U4108 ( .A1(n12744), .A2(n17556), .Z(n31923) );
  INV_X2 U4110 ( .I(n33665), .ZN(n32930) );
  OR2_X1 U4114 ( .A1(n502), .A2(n5433), .Z(n31924) );
  INV_X2 U4116 ( .I(n20423), .ZN(n20566) );
  OAI21_X1 U4117 ( .A1(n28786), .A2(n1170), .B(n33241), .ZN(n32903) );
  OAI22_X2 U4118 ( .A1(n31444), .A2(n15714), .B1(n20224), .B2(n1030), .ZN(
        n1923) );
  AND2_X1 U4125 ( .A1(n21239), .A2(n5822), .Z(n31925) );
  AND2_X1 U4127 ( .A1(n30769), .A2(n26337), .Z(n31926) );
  OR2_X1 U4130 ( .A1(n8875), .A2(n30033), .Z(n31927) );
  INV_X1 U4131 ( .I(n21693), .ZN(n11301) );
  INV_X1 U4133 ( .I(n27635), .ZN(n33242) );
  INV_X2 U4138 ( .I(n7289), .ZN(n34050) );
  XNOR2_X1 U4143 ( .A1(n9536), .A2(n30018), .ZN(n31928) );
  XNOR2_X1 U4145 ( .A1(n14416), .A2(n15969), .ZN(n31929) );
  INV_X1 U4148 ( .I(n26317), .ZN(n11250) );
  INV_X4 U4150 ( .I(n28203), .ZN(n8029) );
  XNOR2_X1 U4151 ( .A1(n6543), .A2(n7152), .ZN(n31931) );
  XOR2_X1 U4153 ( .A1(n2309), .A2(n31303), .Z(n31932) );
  INV_X1 U4155 ( .I(n9535), .ZN(n22642) );
  CLKBUF_X4 U4157 ( .I(n9535), .Z(n33594) );
  OR2_X2 U4159 ( .A1(n22622), .A2(n22340), .Z(n31933) );
  NOR2_X2 U4162 ( .A1(n4396), .A2(n29288), .ZN(n33283) );
  BUF_X4 U4164 ( .I(n23005), .Z(n31942) );
  AND2_X1 U4167 ( .A1(n27752), .A2(n30293), .Z(n31935) );
  NAND2_X2 U4177 ( .A1(n33126), .A2(n11382), .ZN(n23391) );
  AND2_X1 U4180 ( .A1(n10031), .A2(n15301), .Z(n31936) );
  OR2_X2 U4183 ( .A1(n13894), .A2(n4700), .Z(n31937) );
  INV_X1 U4184 ( .I(n15722), .ZN(n23935) );
  INV_X1 U4191 ( .I(n10463), .ZN(n23918) );
  CLKBUF_X4 U4192 ( .I(n10463), .Z(n8760) );
  BUF_X4 U4198 ( .I(n23586), .Z(n16496) );
  AND2_X2 U4199 ( .A1(n31915), .A2(n26641), .Z(n31938) );
  INV_X2 U4203 ( .I(n24095), .ZN(n24097) );
  INV_X2 U4205 ( .I(n24171), .ZN(n24271) );
  INV_X4 U4208 ( .I(n29305), .ZN(n32308) );
  XOR2_X1 U4209 ( .A1(n27360), .A2(n24470), .Z(n31939) );
  INV_X2 U4212 ( .I(n25412), .ZN(n25406) );
  CLKBUF_X4 U4223 ( .I(n24511), .Z(n25412) );
  AND2_X1 U4228 ( .A1(n1080), .A2(n17120), .Z(n31940) );
  NOR2_X1 U4230 ( .A1(n16939), .A2(n25238), .ZN(n31941) );
  INV_X2 U4231 ( .I(n25044), .ZN(n27610) );
  NAND2_X1 U4246 ( .A1(n22744), .A2(n1266), .ZN(n9085) );
  OAI22_X1 U4248 ( .A1(n22744), .A2(n7310), .B1(n11018), .B2(n1266), .ZN(
        n30633) );
  NAND2_X1 U4250 ( .A1(n18681), .A2(n5700), .ZN(n19295) );
  OAI21_X1 U4251 ( .A1(n18681), .A2(n18683), .B(n29726), .ZN(n7320) );
  NAND2_X1 U4252 ( .A1(n25981), .A2(n18681), .ZN(n29726) );
  INV_X2 U4256 ( .I(n18681), .ZN(n15873) );
  OR2_X2 U4257 ( .A1(n14534), .A2(n32628), .Z(n6192) );
  AND2_X2 U4260 ( .A1(n20468), .A2(n28471), .Z(n17964) );
  BUF_X2 U4264 ( .I(n20468), .Z(n28626) );
  NOR2_X1 U4269 ( .A1(n12263), .A2(n17328), .ZN(n19930) );
  NOR2_X1 U4271 ( .A1(n13253), .A2(n17328), .ZN(n31398) );
  INV_X1 U4324 ( .I(n17328), .ZN(n3562) );
  NOR2_X1 U4327 ( .A1(n20566), .A2(n17328), .ZN(n28043) );
  AND2_X2 U4328 ( .A1(n6531), .A2(n17328), .Z(n15553) );
  AOI21_X1 U4330 ( .A1(n9285), .A2(n12827), .B(n31042), .ZN(n8651) );
  NOR2_X1 U4332 ( .A1(n9285), .A2(n12827), .ZN(n31484) );
  NAND2_X1 U4334 ( .A1(n21553), .A2(n12827), .ZN(n21235) );
  NAND2_X1 U4336 ( .A1(n9285), .A2(n12827), .ZN(n31041) );
  CLKBUF_X4 U4337 ( .I(n7463), .Z(n5820) );
  NOR2_X2 U4343 ( .A1(n13474), .A2(n6553), .ZN(n13142) );
  NAND2_X1 U4351 ( .A1(n32619), .A2(n2612), .ZN(n33795) );
  NAND2_X1 U4354 ( .A1(n30033), .A2(n29523), .ZN(n13115) );
  AOI21_X1 U4355 ( .A1(n21859), .A2(n30033), .B(n21858), .ZN(n2351) );
  INV_X2 U4358 ( .I(n10953), .ZN(n9646) );
  OR2_X2 U4360 ( .A1(n31787), .A2(n17150), .Z(n16091) );
  CLKBUF_X12 U4364 ( .I(n23005), .Z(n31943) );
  AND2_X2 U4368 ( .A1(n28014), .A2(n9753), .Z(n22674) );
  OR3_X2 U4375 ( .A1(n9737), .A2(n32078), .A3(n9910), .Z(n22421) );
  CLKBUF_X4 U4387 ( .I(n19456), .Z(n5825) );
  INV_X2 U4394 ( .I(n19456), .ZN(n19992) );
  AND2_X2 U4395 ( .A1(n17930), .A2(n12375), .Z(n9184) );
  OAI21_X1 U4396 ( .A1(n25306), .A2(n18059), .B(n1215), .ZN(n27443) );
  INV_X1 U4401 ( .I(n23454), .ZN(n23455) );
  AND3_X2 U4402 ( .A1(n21350), .A2(n32505), .A3(n14983), .Z(n3317) );
  NAND2_X1 U4405 ( .A1(n21350), .A2(n30389), .ZN(n16228) );
  NOR2_X1 U4406 ( .A1(n8140), .A2(n28181), .ZN(n2801) );
  INV_X2 U4410 ( .I(n5994), .ZN(n22114) );
  NOR2_X2 U4412 ( .A1(n30908), .A2(n10305), .ZN(n10307) );
  NAND2_X1 U4414 ( .A1(n31461), .A2(n24168), .ZN(n34136) );
  AND2_X2 U4417 ( .A1(n20561), .A2(n20413), .Z(n5953) );
  NOR2_X1 U4419 ( .A1(n33069), .A2(n784), .ZN(n18916) );
  NOR2_X1 U4421 ( .A1(n20119), .A2(n14815), .ZN(n20122) );
  INV_X2 U4425 ( .I(n14815), .ZN(n20021) );
  CLKBUF_X12 U4426 ( .I(n14815), .Z(n8371) );
  AND2_X2 U4428 ( .A1(n20561), .A2(n1636), .Z(n5950) );
  INV_X2 U4435 ( .I(n20561), .ZN(n30931) );
  INV_X1 U4436 ( .I(n30293), .ZN(n22828) );
  OR2_X2 U4437 ( .A1(n16603), .A2(n23144), .Z(n23712) );
  CLKBUF_X12 U4439 ( .I(n652), .Z(n27) );
  OR2_X2 U4440 ( .A1(n7463), .A2(n12055), .Z(n3901) );
  CLKBUF_X12 U4441 ( .I(n26317), .Z(n28692) );
  OAI21_X1 U4443 ( .A1(n9186), .A2(n424), .B(n780), .ZN(n9395) );
  NAND3_X1 U4444 ( .A1(n29088), .A2(n6493), .A3(n424), .ZN(n5687) );
  INV_X2 U4447 ( .I(n424), .ZN(n6908) );
  INV_X1 U4449 ( .I(n23230), .ZN(n12922) );
  NOR2_X1 U4454 ( .A1(n24060), .A2(n30191), .ZN(n26580) );
  NAND2_X1 U4456 ( .A1(n3147), .A2(n30191), .ZN(n14725) );
  AOI22_X1 U4457 ( .A1(n20524), .A2(n2958), .B1(n868), .B2(n31504), .ZN(n4398)
         );
  NAND2_X1 U4458 ( .A1(n2879), .A2(n2958), .ZN(n12771) );
  INV_X1 U4459 ( .I(n2958), .ZN(n33225) );
  OR2_X2 U4460 ( .A1(n28979), .A2(n26330), .Z(n26709) );
  INV_X1 U4461 ( .I(n13762), .ZN(n805) );
  AOI22_X1 U4464 ( .A1(n22950), .A2(n22949), .B1(n22951), .B2(n13762), .ZN(
        n17202) );
  CLKBUF_X12 U4467 ( .I(n13195), .Z(n27028) );
  INV_X1 U4469 ( .I(n3395), .ZN(n2763) );
  NAND2_X1 U4476 ( .A1(n2913), .A2(n24315), .ZN(n12005) );
  CLKBUF_X12 U4477 ( .I(n24315), .Z(n31377) );
  NOR2_X1 U4480 ( .A1(n31072), .A2(n33117), .ZN(n20308) );
  NOR2_X1 U4482 ( .A1(n742), .A2(n33117), .ZN(n3226) );
  AND2_X2 U4489 ( .A1(n33117), .A2(n26363), .Z(n29432) );
  INV_X1 U4490 ( .I(n24254), .ZN(n29120) );
  INV_X1 U4494 ( .I(n24747), .ZN(n33058) );
  CLKBUF_X12 U4495 ( .I(n22873), .Z(n18240) );
  NOR2_X1 U4496 ( .A1(n4135), .A2(n9377), .ZN(n33861) );
  BUF_X2 U4500 ( .I(n18575), .Z(n15108) );
  INV_X2 U4501 ( .I(n21579), .ZN(n21805) );
  OAI21_X1 U4503 ( .A1(n32634), .A2(n19093), .B(n8141), .ZN(n8013) );
  OR3_X2 U4507 ( .A1(n29047), .A2(n8141), .A3(n5813), .Z(n27930) );
  NAND2_X1 U4509 ( .A1(n8141), .A2(n19095), .ZN(n19097) );
  OAI22_X1 U4510 ( .A1(n19977), .A2(n14761), .B1(n1699), .B2(n32745), .ZN(
        n29548) );
  NAND2_X1 U4511 ( .A1(n28011), .A2(n20519), .ZN(n20288) );
  INV_X2 U4512 ( .I(n28011), .ZN(n16174) );
  OAI21_X1 U4519 ( .A1(n21466), .A2(n1134), .B(n6678), .ZN(n16889) );
  INV_X1 U4521 ( .I(n21466), .ZN(n16577) );
  NAND2_X1 U4524 ( .A1(n19165), .A2(n4835), .ZN(n19153) );
  CLKBUF_X4 U4530 ( .I(n8396), .Z(n7090) );
  INV_X1 U4533 ( .I(n8396), .ZN(n22460) );
  NAND2_X1 U4534 ( .A1(n17516), .A2(n1439), .ZN(n18316) );
  INV_X2 U4537 ( .I(n17516), .ZN(n18710) );
  BUF_X2 U4541 ( .I(n17516), .Z(n33783) );
  INV_X2 U4544 ( .I(n29634), .ZN(n24152) );
  AND2_X2 U4553 ( .A1(n31787), .A2(n23833), .Z(n29375) );
  OR2_X2 U4558 ( .A1(n23925), .A2(n14585), .Z(n11192) );
  BUF_X2 U4559 ( .I(n25589), .Z(n31945) );
  CLKBUF_X12 U4560 ( .I(n25703), .Z(n16323) );
  OR2_X2 U4561 ( .A1(n15057), .A2(n10708), .Z(n13650) );
  OAI21_X1 U4564 ( .A1(n6003), .A2(n24095), .B(n24015), .ZN(n4393) );
  AND3_X2 U4566 ( .A1(n14443), .A2(n6001), .A3(n24095), .Z(n29396) );
  NOR2_X1 U4567 ( .A1(n24095), .A2(n33868), .ZN(n12312) );
  AOI21_X1 U4571 ( .A1(n12452), .A2(n21463), .B(n26439), .ZN(n26325) );
  OAI21_X1 U4574 ( .A1(n33810), .A2(n21604), .B(n26439), .ZN(n27454) );
  INV_X2 U4588 ( .I(n30894), .ZN(n1177) );
  NAND2_X1 U4592 ( .A1(n30894), .A2(n19274), .ZN(n19323) );
  INV_X2 U4593 ( .I(n27419), .ZN(n776) );
  OR2_X2 U4596 ( .A1(n20148), .A2(n7865), .Z(n29422) );
  INV_X1 U4598 ( .I(n17098), .ZN(n16345) );
  NAND3_X1 U4602 ( .A1(n24325), .A2(n24328), .A3(n10987), .ZN(n26990) );
  NOR2_X1 U4617 ( .A1(n2302), .A2(n30219), .ZN(n2301) );
  NAND2_X1 U4618 ( .A1(n28429), .A2(n14691), .ZN(n21649) );
  NOR2_X1 U4620 ( .A1(n14691), .A2(n28429), .ZN(n2061) );
  CLKBUF_X12 U4621 ( .I(n28429), .Z(n33139) );
  CLKBUF_X12 U4622 ( .I(n17779), .Z(n17118) );
  INV_X1 U4626 ( .I(n17779), .ZN(n24974) );
  AND2_X2 U4628 ( .A1(n23746), .A2(n23603), .Z(n15659) );
  NOR2_X1 U4630 ( .A1(n11850), .A2(n31915), .ZN(n29590) );
  NOR2_X1 U4637 ( .A1(n6394), .A2(n11850), .ZN(n32574) );
  NAND2_X1 U4638 ( .A1(n4774), .A2(n12981), .ZN(n24027) );
  INV_X1 U4642 ( .I(n12981), .ZN(n12574) );
  CLKBUF_X12 U4660 ( .I(n12981), .Z(n4118) );
  OR2_X2 U4661 ( .A1(n23087), .A2(n23086), .Z(n26242) );
  NAND3_X2 U4663 ( .A1(n9915), .A2(n9916), .A3(n25390), .ZN(n33064) );
  CLKBUF_X4 U4666 ( .I(n23197), .Z(n23806) );
  CLKBUF_X12 U4671 ( .I(n30865), .Z(n31947) );
  CLKBUF_X12 U4672 ( .I(n30865), .Z(n31949) );
  INV_X1 U4674 ( .I(n13723), .ZN(n20945) );
  BUF_X4 U4678 ( .I(n25988), .Z(n31950) );
  INV_X1 U4679 ( .I(n11710), .ZN(n20332) );
  OAI21_X1 U4684 ( .A1(n6475), .A2(n31390), .B(n11710), .ZN(n8702) );
  NAND2_X1 U4686 ( .A1(n7873), .A2(n20613), .ZN(n28437) );
  NOR2_X1 U4690 ( .A1(n14129), .A2(n22968), .ZN(n22884) );
  INV_X1 U4692 ( .I(n14129), .ZN(n17084) );
  AND2_X2 U4693 ( .A1(n14129), .A2(n7802), .Z(n27639) );
  INV_X2 U4698 ( .I(n12323), .ZN(n28406) );
  AOI21_X1 U4712 ( .A1(n3717), .A2(n12323), .B(n30313), .ZN(n21176) );
  NAND2_X1 U4714 ( .A1(n12323), .A2(n595), .ZN(n21055) );
  AOI21_X1 U4717 ( .A1(n13386), .A2(n2638), .B(n4184), .ZN(n13384) );
  INV_X1 U4719 ( .I(n23741), .ZN(n23769) );
  NOR2_X1 U4721 ( .A1(n23741), .A2(n386), .ZN(n8093) );
  AOI21_X1 U4722 ( .A1(n23741), .A2(n17396), .B(n30895), .ZN(n33542) );
  AOI21_X1 U4727 ( .A1(n23741), .A2(n23597), .B(n23598), .ZN(n14551) );
  NAND2_X1 U4729 ( .A1(n23741), .A2(n30089), .ZN(n2878) );
  NAND2_X1 U4737 ( .A1(n27183), .A2(n25317), .ZN(n1803) );
  INV_X1 U4753 ( .I(n25317), .ZN(n31178) );
  AOI21_X1 U4757 ( .A1(n977), .A2(n13773), .B(n11943), .ZN(n4514) );
  OAI22_X1 U4759 ( .A1(n16320), .A2(n11943), .B1(n23882), .B2(n8544), .ZN(
        n33535) );
  NAND2_X1 U4765 ( .A1(n9714), .A2(n11943), .ZN(n7167) );
  AOI21_X1 U4770 ( .A1(n16320), .A2(n11943), .B(n8544), .ZN(n10620) );
  NAND2_X1 U4773 ( .A1(n15261), .A2(n21438), .ZN(n21440) );
  INV_X2 U4775 ( .I(n21438), .ZN(n15589) );
  OR2_X2 U4780 ( .A1(n29101), .A2(n15229), .Z(n17936) );
  AOI22_X1 U4785 ( .A1(n19030), .A2(n29223), .B1(n19300), .B2(n19029), .ZN(
        n31066) );
  AOI22_X1 U4786 ( .A1(n19085), .A2(n29223), .B1(n19084), .B2(n19300), .ZN(
        n28237) );
  AND3_X2 U4794 ( .A1(n20946), .A2(n10599), .A3(n10787), .Z(n34159) );
  OR2_X2 U4797 ( .A1(n20946), .A2(n13195), .Z(n21313) );
  NAND2_X1 U4801 ( .A1(n11086), .A2(n2821), .ZN(n20261) );
  NAND2_X1 U4809 ( .A1(n919), .A2(n28580), .ZN(n26527) );
  NOR2_X1 U4813 ( .A1(n28580), .A2(n12535), .ZN(n32148) );
  NAND2_X1 U4814 ( .A1(n28580), .A2(n10720), .ZN(n32435) );
  INV_X1 U4824 ( .I(n28580), .ZN(n21645) );
  INV_X1 U4825 ( .I(n12424), .ZN(n21777) );
  CLKBUF_X12 U4826 ( .I(n12424), .Z(n30940) );
  CLKBUF_X4 U4828 ( .I(n12424), .Z(n11861) );
  CLKBUF_X12 U4837 ( .I(n24372), .Z(n17833) );
  CLKBUF_X4 U4838 ( .I(n19829), .Z(n31951) );
  NAND2_X1 U4840 ( .A1(n23087), .A2(n4834), .ZN(n28427) );
  CLKBUF_X12 U4841 ( .I(n12804), .Z(n179) );
  INV_X1 U4851 ( .I(n20455), .ZN(n20457) );
  NAND2_X1 U4860 ( .A1(n20455), .A2(n15468), .ZN(n14767) );
  INV_X1 U4864 ( .I(n17517), .ZN(n33814) );
  NOR2_X1 U4866 ( .A1(n23110), .A2(n3103), .ZN(n22813) );
  NAND2_X1 U4870 ( .A1(n853), .A2(n3103), .ZN(n4935) );
  NAND2_X1 U4872 ( .A1(n16022), .A2(n3103), .ZN(n23108) );
  INV_X2 U4874 ( .I(n3103), .ZN(n6012) );
  OAI21_X1 U4875 ( .A1(n30168), .A2(n30167), .B(n22999), .ZN(n4305) );
  INV_X1 U4876 ( .I(n22999), .ZN(n7220) );
  OR2_X2 U4877 ( .A1(n9280), .A2(n22999), .Z(n9213) );
  OAI21_X2 U4880 ( .A1(n23101), .A2(n11956), .B(n22999), .ZN(n15935) );
  NAND2_X1 U4882 ( .A1(n29883), .A2(n7935), .ZN(n32328) );
  OR2_X2 U4884 ( .A1(n18039), .A2(n26699), .Z(n8182) );
  NAND2_X1 U4885 ( .A1(n31129), .A2(n23051), .ZN(n6102) );
  INV_X2 U4887 ( .I(n31129), .ZN(n1108) );
  NAND2_X1 U4888 ( .A1(n772), .A2(n31129), .ZN(n1746) );
  AND2_X2 U4889 ( .A1(n5962), .A2(n11986), .Z(n8846) );
  INV_X2 U4890 ( .I(n32253), .ZN(n14625) );
  NOR2_X1 U4892 ( .A1(n7279), .A2(n20627), .ZN(n8242) );
  OR2_X2 U4895 ( .A1(n20627), .A2(n7280), .Z(n17002) );
  BUF_X2 U4896 ( .I(n16954), .Z(n8886) );
  NAND2_X1 U4899 ( .A1(n16954), .A2(n15302), .ZN(n27338) );
  NOR2_X1 U4900 ( .A1(n28581), .A2(n16954), .ZN(n31231) );
  NOR2_X1 U4903 ( .A1(n14893), .A2(n5625), .ZN(n12996) );
  NAND2_X1 U4906 ( .A1(n19057), .A2(n5625), .ZN(n18944) );
  CLKBUF_X4 U4910 ( .I(n5086), .Z(n31954) );
  INV_X1 U4913 ( .I(n21891), .ZN(n2082) );
  OR2_X2 U4922 ( .A1(n31497), .A2(n24216), .Z(n215) );
  INV_X1 U4929 ( .I(n31497), .ZN(n24111) );
  NAND2_X1 U4932 ( .A1(n13175), .A2(n31497), .ZN(n13176) );
  NAND2_X1 U4937 ( .A1(n22791), .A2(n14392), .ZN(n31564) );
  NAND2_X1 U4939 ( .A1(n22871), .A2(n22791), .ZN(n22792) );
  INV_X1 U4940 ( .I(n7046), .ZN(n4063) );
  INV_X1 U4941 ( .I(n27880), .ZN(n621) );
  INV_X1 U4944 ( .I(n33288), .ZN(n30425) );
  OAI21_X1 U4946 ( .A1(n33288), .A2(n20317), .B(n20471), .ZN(n19402) );
  NAND3_X1 U4951 ( .A1(n34113), .A2(n20471), .A3(n33288), .ZN(n20248) );
  NAND2_X1 U4952 ( .A1(n16144), .A2(n28064), .ZN(n13599) );
  NAND3_X1 U4956 ( .A1(n16144), .A2(n20531), .A3(n20529), .ZN(n32840) );
  NOR2_X1 U4960 ( .A1(n5274), .A2(n32967), .ZN(n33344) );
  AOI21_X1 U4961 ( .A1(n1112), .A2(n5274), .B(n22931), .ZN(n30875) );
  OAI21_X1 U4966 ( .A1(n17297), .A2(n20324), .B(n20515), .ZN(n26576) );
  NAND2_X1 U4968 ( .A1(n16174), .A2(n20515), .ZN(n6491) );
  CLKBUF_X4 U4970 ( .I(n26750), .Z(n33544) );
  NAND2_X1 U4972 ( .A1(n1550), .A2(n24286), .ZN(n24047) );
  CLKBUF_X12 U4978 ( .I(n24286), .Z(n28300) );
  INV_X1 U4985 ( .I(n24286), .ZN(n17277) );
  INV_X2 U4993 ( .I(n1130), .ZN(n31706) );
  NAND2_X1 U5002 ( .A1(n879), .A2(n19330), .ZN(n19331) );
  INV_X1 U5003 ( .I(n17891), .ZN(n22379) );
  CLKBUF_X12 U5008 ( .I(n17891), .Z(n2697) );
  INV_X2 U5012 ( .I(n22361), .ZN(n6149) );
  NOR2_X1 U5015 ( .A1(n22361), .A2(n9575), .ZN(n27580) );
  NOR2_X1 U5018 ( .A1(n4135), .A2(n22361), .ZN(n32692) );
  NOR2_X1 U5019 ( .A1(n5119), .A2(n5118), .ZN(n19013) );
  OAI21_X1 U5021 ( .A1(n5118), .A2(n28929), .B(n6511), .ZN(n11489) );
  INV_X1 U5024 ( .I(n11720), .ZN(n11911) );
  NOR2_X1 U5025 ( .A1(n20507), .A2(n31907), .ZN(n16167) );
  NAND2_X1 U5026 ( .A1(n31907), .A2(n16452), .ZN(n33501) );
  AOI21_X1 U5027 ( .A1(n878), .A2(n5760), .B(n14498), .ZN(n18497) );
  NOR2_X1 U5032 ( .A1(n19089), .A2(n14498), .ZN(n15021) );
  INV_X2 U5038 ( .I(n14498), .ZN(n1385) );
  NOR2_X1 U5039 ( .A1(n26603), .A2(n32253), .ZN(n6142) );
  NAND2_X1 U5040 ( .A1(n15777), .A2(n9126), .ZN(n27272) );
  OAI21_X1 U5043 ( .A1(n16518), .A2(n28028), .B(n32240), .ZN(n20206) );
  NAND3_X1 U5044 ( .A1(n1153), .A2(n20534), .A3(n28028), .ZN(n18170) );
  INV_X2 U5051 ( .I(n28028), .ZN(n8206) );
  AOI22_X1 U5055 ( .A1(n17896), .A2(n31009), .B1(n28812), .B2(n4254), .ZN(
        n2609) );
  NOR2_X1 U5058 ( .A1(n19938), .A2(n16105), .ZN(n32109) );
  NOR2_X2 U5066 ( .A1(n28418), .A2(n28419), .ZN(n12599) );
  AOI21_X1 U5071 ( .A1(n16374), .A2(n16218), .B(n15893), .ZN(n13915) );
  NAND2_X1 U5072 ( .A1(n16374), .A2(n20236), .ZN(n14836) );
  NOR2_X1 U5073 ( .A1(n13768), .A2(n16374), .ZN(n15893) );
  OR2_X2 U5074 ( .A1(n16374), .A2(n20555), .Z(n32066) );
  INV_X1 U5075 ( .I(n9434), .ZN(n28647) );
  NAND2_X1 U5077 ( .A1(n9434), .A2(n29133), .ZN(n9637) );
  AND2_X2 U5081 ( .A1(n26848), .A2(n9744), .Z(n7723) );
  OR2_X2 U5085 ( .A1(n9744), .A2(n8899), .Z(n21263) );
  NAND2_X1 U5087 ( .A1(n34139), .A2(n18295), .ZN(n12154) );
  INV_X2 U5089 ( .I(n17817), .ZN(n19196) );
  NAND2_X1 U5099 ( .A1(n6290), .A2(n11085), .ZN(n19164) );
  NOR2_X1 U5100 ( .A1(n1165), .A2(n5433), .ZN(n11855) );
  BUF_X2 U5106 ( .I(n3007), .Z(n28974) );
  INV_X2 U5108 ( .I(n3007), .ZN(n17739) );
  OR2_X2 U5112 ( .A1(n7965), .A2(n2655), .Z(n26867) );
  CLKBUF_X12 U5118 ( .I(n7293), .Z(n31956) );
  CLKBUF_X12 U5119 ( .I(n7293), .Z(n31958) );
  NAND3_X1 U5126 ( .A1(n14161), .A2(n20628), .A3(n53), .ZN(n13172) );
  INV_X1 U5127 ( .I(n14161), .ZN(n20629) );
  NOR2_X1 U5132 ( .A1(n14005), .A2(n14161), .ZN(n30022) );
  NAND2_X1 U5136 ( .A1(n9616), .A2(n9625), .ZN(n8567) );
  CLKBUF_X4 U5138 ( .I(n9616), .Z(n891) );
  AOI21_X1 U5141 ( .A1(n25088), .A2(n25083), .B(n25082), .ZN(n30858) );
  BUF_X1 U5142 ( .I(n24960), .Z(n28662) );
  OAI21_X1 U5144 ( .A1(n13273), .A2(n30396), .B(n1213), .ZN(n6822) );
  BUF_X1 U5150 ( .I(n3565), .Z(n32678) );
  CLKBUF_X2 U5154 ( .I(n25188), .Z(n12476) );
  CLKBUF_X1 U5159 ( .I(n24646), .Z(n32759) );
  CLKBUF_X2 U5163 ( .I(n13695), .Z(n33699) );
  CLKBUF_X2 U5170 ( .I(n24618), .Z(n33348) );
  CLKBUF_X2 U5179 ( .I(n27922), .Z(n33492) );
  INV_X1 U5197 ( .I(n13458), .ZN(n32552) );
  CLKBUF_X2 U5201 ( .I(n24094), .Z(n32459) );
  NOR2_X1 U5205 ( .A1(n24263), .A2(n26950), .ZN(n5936) );
  INV_X2 U5207 ( .I(n24210), .ZN(n24322) );
  INV_X2 U5208 ( .I(n24008), .ZN(n9962) );
  NAND2_X1 U5209 ( .A1(n14038), .A2(n14039), .ZN(n14037) );
  INV_X1 U5210 ( .I(n5627), .ZN(n33104) );
  BUF_X2 U5211 ( .I(n23808), .Z(n32477) );
  CLKBUF_X2 U5212 ( .I(n8408), .Z(n33216) );
  INV_X1 U5215 ( .I(n23742), .ZN(n34036) );
  BUF_X2 U5216 ( .I(n23775), .Z(n33011) );
  CLKBUF_X2 U5218 ( .I(n29498), .Z(n32657) );
  CLKBUF_X1 U5219 ( .I(n10279), .Z(n33924) );
  INV_X2 U5220 ( .I(n662), .ZN(n31959) );
  CLKBUF_X2 U5225 ( .I(n23389), .Z(n32243) );
  NOR2_X1 U5226 ( .A1(n5983), .A2(n11308), .ZN(n26995) );
  BUF_X2 U5229 ( .I(n31937), .Z(n33522) );
  OAI22_X1 U5231 ( .A1(n3997), .A2(n7181), .B1(n22827), .B2(n11059), .ZN(n4476) );
  AOI21_X1 U5237 ( .A1(n28853), .A2(n28408), .B(n2479), .ZN(n32368) );
  BUF_X1 U5239 ( .I(n22880), .Z(n33395) );
  NAND2_X1 U5243 ( .A1(n22855), .A2(n28649), .ZN(n32509) );
  OR2_X1 U5246 ( .A1(n23057), .A2(n23056), .Z(n32086) );
  BUF_X1 U5248 ( .I(n11983), .Z(n34097) );
  NOR2_X1 U5250 ( .A1(n6782), .A2(n22945), .ZN(n33923) );
  NAND2_X1 U5251 ( .A1(n31636), .A2(n16627), .ZN(n31635) );
  NAND2_X1 U5253 ( .A1(n33056), .A2(n10796), .ZN(n29563) );
  INV_X1 U5254 ( .I(n22404), .ZN(n33402) );
  NAND2_X1 U5255 ( .A1(n16558), .A2(n22412), .ZN(n15119) );
  NOR2_X1 U5257 ( .A1(n22466), .A2(n998), .ZN(n28101) );
  CLKBUF_X2 U5258 ( .I(n27122), .Z(n32378) );
  CLKBUF_X2 U5262 ( .I(n7072), .Z(n33966) );
  OR2_X1 U5266 ( .A1(n14845), .A2(n16392), .Z(n32080) );
  CLKBUF_X2 U5269 ( .I(n22318), .Z(n32154) );
  CLKBUF_X4 U5274 ( .I(n7545), .Z(n32537) );
  CLKBUF_X4 U5275 ( .I(n14953), .Z(n2896) );
  INV_X1 U5279 ( .I(n33459), .ZN(n32314) );
  INV_X1 U5281 ( .I(n26206), .ZN(n32348) );
  NAND2_X1 U5285 ( .A1(n3472), .A2(n17077), .ZN(n34104) );
  CLKBUF_X1 U5287 ( .I(n914), .Z(n33322) );
  NAND2_X1 U5289 ( .A1(n31007), .A2(n32374), .ZN(n32373) );
  NOR2_X1 U5292 ( .A1(n21842), .A2(n30346), .ZN(n33907) );
  INV_X1 U5294 ( .I(n338), .ZN(n33908) );
  CLKBUF_X2 U5296 ( .I(n1652), .Z(n32282) );
  CLKBUF_X4 U5302 ( .I(n27379), .Z(n33810) );
  CLKBUF_X2 U5305 ( .I(n27336), .Z(n34098) );
  CLKBUF_X2 U5306 ( .I(n16278), .Z(n32642) );
  CLKBUF_X1 U5313 ( .I(n14864), .Z(n33833) );
  BUF_X4 U5314 ( .I(n5830), .Z(n31960) );
  AOI21_X1 U5318 ( .A1(n27689), .A2(n21151), .B(n27688), .ZN(n26494) );
  OAI21_X1 U5319 ( .A1(n21286), .A2(n32625), .B(n21285), .ZN(n32168) );
  CLKBUF_X2 U5321 ( .I(n21241), .Z(n33882) );
  CLKBUF_X2 U5323 ( .I(n16668), .Z(n33741) );
  NAND2_X1 U5333 ( .A1(n21400), .A2(n15874), .ZN(n32624) );
  CLKBUF_X2 U5344 ( .I(n4274), .Z(n34037) );
  NOR2_X1 U5345 ( .A1(n16473), .A2(n21152), .ZN(n33979) );
  BUF_X2 U5346 ( .I(n599), .Z(n33649) );
  CLKBUF_X2 U5349 ( .I(n8028), .Z(n16629) );
  NOR2_X1 U5350 ( .A1(n13573), .A2(n11635), .ZN(n30083) );
  BUF_X1 U5351 ( .I(n6431), .Z(n27375) );
  NOR2_X1 U5355 ( .A1(n20277), .A2(n29453), .ZN(n32304) );
  NAND2_X1 U5356 ( .A1(n20231), .A2(n20413), .ZN(n285) );
  OAI21_X1 U5359 ( .A1(n20492), .A2(n14863), .B(n33944), .ZN(n30632) );
  NAND2_X1 U5360 ( .A1(n26881), .A2(n20310), .ZN(n9832) );
  CLKBUF_X2 U5361 ( .I(n20472), .Z(n32201) );
  INV_X1 U5362 ( .I(n6536), .ZN(n33341) );
  CLKBUF_X2 U5363 ( .I(n1351), .Z(n32953) );
  CLKBUF_X2 U5364 ( .I(n20534), .Z(n32329) );
  NAND2_X1 U5365 ( .A1(n5781), .A2(n26585), .ZN(n17425) );
  CLKBUF_X4 U5366 ( .I(n30637), .Z(n33721) );
  CLKBUF_X2 U5367 ( .I(n20485), .Z(n31009) );
  NAND2_X1 U5368 ( .A1(n30017), .A2(n14281), .ZN(n33136) );
  CLKBUF_X2 U5371 ( .I(n20138), .Z(n32371) );
  CLKBUF_X2 U5376 ( .I(n17670), .Z(n32559) );
  CLKBUF_X2 U5379 ( .I(n34119), .Z(n33835) );
  NAND2_X1 U5380 ( .A1(n10192), .A2(n11798), .ZN(n33983) );
  BUF_X4 U5383 ( .I(n7492), .Z(n10472) );
  CLKBUF_X2 U5385 ( .I(n14194), .Z(n32485) );
  NAND2_X1 U5386 ( .A1(n27941), .A2(n32805), .ZN(n33230) );
  CLKBUF_X2 U5389 ( .I(n29781), .Z(n32401) );
  BUF_X1 U5391 ( .I(n25971), .Z(n34040) );
  BUF_X2 U5397 ( .I(n34107), .Z(n32908) );
  CLKBUF_X1 U5398 ( .I(n4016), .Z(n32805) );
  OAI22_X1 U5400 ( .A1(n27641), .A2(n18629), .B1(n18628), .B2(n18627), .ZN(
        n19149) );
  NOR2_X1 U5406 ( .A1(n18885), .A2(n10669), .ZN(n33255) );
  INV_X1 U5407 ( .I(n4733), .ZN(n18622) );
  NAND2_X1 U5408 ( .A1(n11123), .A2(n17419), .ZN(n33421) );
  INV_X1 U5409 ( .I(n29514), .ZN(n33101) );
  BUF_X2 U5410 ( .I(n18601), .Z(n33472) );
  NOR2_X1 U5414 ( .A1(n28686), .A2(n18228), .ZN(n33309) );
  CLKBUF_X2 U5416 ( .I(n26980), .Z(n32337) );
  NAND3_X1 U5421 ( .A1(n32724), .A2(n28516), .A3(n28517), .ZN(n32730) );
  AOI21_X1 U5424 ( .A1(n25683), .A2(n25684), .B(n25682), .ZN(n16541) );
  NAND2_X1 U5427 ( .A1(n14101), .A2(n16246), .ZN(n32724) );
  NOR2_X1 U5438 ( .A1(n33464), .A2(n25273), .ZN(n14070) );
  OAI22_X1 U5441 ( .A1(n25456), .A2(n33946), .B1(n25419), .B2(n25420), .ZN(
        n30746) );
  AOI22_X1 U5449 ( .A1(n25747), .A2(n25748), .B1(n25749), .B2(n25750), .ZN(
        n31599) );
  OAI22_X1 U5457 ( .A1(n10823), .A2(n1951), .B1(n10821), .B2(n1950), .ZN(
        n32190) );
  INV_X1 U5462 ( .I(n25857), .ZN(n406) );
  OAI22_X1 U5473 ( .A1(n33702), .A2(n788), .B1(n25128), .B2(n33138), .ZN(n6814) );
  NAND2_X1 U5475 ( .A1(n25412), .A2(n33921), .ZN(n9754) );
  CLKBUF_X2 U5478 ( .I(n31236), .Z(n33414) );
  BUF_X2 U5483 ( .I(n16509), .Z(n15359) );
  NOR2_X1 U5485 ( .A1(n25583), .A2(n28242), .ZN(n28098) );
  INV_X1 U5488 ( .I(n32427), .ZN(n7768) );
  NAND2_X1 U5494 ( .A1(n12386), .A2(n12369), .ZN(n32825) );
  NAND2_X1 U5497 ( .A1(n11994), .A2(n33199), .ZN(n26400) );
  BUF_X1 U5505 ( .I(n25403), .Z(n32920) );
  NOR2_X1 U5510 ( .A1(n24730), .A2(n17120), .ZN(n32556) );
  CLKBUF_X2 U5517 ( .I(n25865), .Z(n33196) );
  INV_X2 U5518 ( .I(n33919), .ZN(n31962) );
  CLKBUF_X2 U5527 ( .I(n17861), .Z(n32659) );
  CLKBUF_X4 U5530 ( .I(n11372), .Z(n33493) );
  BUF_X2 U5533 ( .I(n31783), .Z(n33761) );
  INV_X1 U5534 ( .I(n6863), .ZN(n32639) );
  CLKBUF_X2 U5539 ( .I(n14665), .Z(n33574) );
  INV_X1 U5541 ( .I(n16045), .ZN(n33375) );
  CLKBUF_X2 U5543 ( .I(n24760), .Z(n33447) );
  CLKBUF_X2 U5549 ( .I(n30323), .Z(n32660) );
  OAI21_X1 U5557 ( .A1(n23701), .A2(n6003), .B(n33727), .ZN(n23702) );
  INV_X1 U5560 ( .I(n32677), .ZN(n26851) );
  NAND2_X1 U5561 ( .A1(n1240), .A2(n24219), .ZN(n23625) );
  NAND2_X1 U5571 ( .A1(n29567), .A2(n29566), .ZN(n33853) );
  BUF_X1 U5574 ( .I(n14386), .Z(n33470) );
  NAND2_X1 U5575 ( .A1(n11200), .A2(n28945), .ZN(n9687) );
  CLKBUF_X2 U5577 ( .I(n24159), .Z(n32176) );
  CLKBUF_X2 U5579 ( .I(n15720), .Z(n33425) );
  CLKBUF_X2 U5585 ( .I(n4286), .Z(n32936) );
  CLKBUF_X2 U5590 ( .I(n33832), .Z(n32102) );
  CLKBUF_X4 U5593 ( .I(n11041), .Z(n9066) );
  INV_X1 U5597 ( .I(n2558), .ZN(n33532) );
  INV_X2 U5602 ( .I(n24106), .ZN(n24104) );
  INV_X2 U5603 ( .I(n8412), .ZN(n795) );
  BUF_X4 U5604 ( .I(n11789), .Z(n10687) );
  NAND2_X1 U5616 ( .A1(n32336), .A2(n23749), .ZN(n27340) );
  INV_X2 U5618 ( .I(n14080), .ZN(n23884) );
  CLKBUF_X4 U5622 ( .I(n386), .Z(n33867) );
  CLKBUF_X2 U5624 ( .I(n32711), .Z(n33097) );
  NOR2_X1 U5626 ( .A1(n23804), .A2(n14325), .ZN(n33595) );
  CLKBUF_X2 U5628 ( .I(n23822), .Z(n33110) );
  INV_X1 U5630 ( .I(n33679), .ZN(n32973) );
  OAI21_X1 U5635 ( .A1(n16496), .A2(n15623), .B(n8145), .ZN(n12777) );
  NOR2_X1 U5642 ( .A1(n6247), .A2(n33812), .ZN(n17563) );
  CLKBUF_X2 U5646 ( .I(n4892), .Z(n33221) );
  BUF_X1 U5648 ( .I(n10213), .Z(n26882) );
  CLKBUF_X2 U5651 ( .I(n23603), .Z(n33679) );
  INV_X2 U5655 ( .I(n29498), .ZN(n23894) );
  CLKBUF_X2 U5656 ( .I(n10673), .Z(n33936) );
  BUF_X2 U5658 ( .I(n23931), .Z(n10993) );
  CLKBUF_X2 U5660 ( .I(n7699), .Z(n33345) );
  CLKBUF_X2 U5661 ( .I(n9796), .Z(n33670) );
  INV_X1 U5662 ( .I(n23437), .ZN(n32640) );
  INV_X1 U5667 ( .I(n4273), .ZN(n32645) );
  INV_X1 U5671 ( .I(n23520), .ZN(n32922) );
  CLKBUF_X2 U5673 ( .I(n23292), .Z(n34047) );
  CLKBUF_X2 U5676 ( .I(n6373), .Z(n28927) );
  CLKBUF_X2 U5677 ( .I(n31727), .Z(n32516) );
  NAND3_X1 U5682 ( .A1(n22804), .A2(n33596), .A3(n22805), .ZN(n29818) );
  NAND2_X1 U5686 ( .A1(n22756), .A2(n14977), .ZN(n33347) );
  NAND2_X1 U5687 ( .A1(n12742), .A2(n32368), .ZN(n28846) );
  NAND2_X1 U5688 ( .A1(n31795), .A2(n22951), .ZN(n3201) );
  INV_X1 U5689 ( .I(n22694), .ZN(n33360) );
  OAI21_X1 U5691 ( .A1(n33923), .A2(n30455), .B(n6942), .ZN(n12443) );
  CLKBUF_X4 U5693 ( .I(n28934), .Z(n32935) );
  OR2_X1 U5694 ( .A1(n1577), .A2(n22885), .Z(n5259) );
  NAND2_X1 U5697 ( .A1(n22962), .A2(n29952), .ZN(n30946) );
  CLKBUF_X2 U5698 ( .I(n14686), .Z(n33968) );
  CLKBUF_X8 U5707 ( .I(n12619), .Z(n33675) );
  BUF_X2 U5721 ( .I(n22990), .Z(n31798) );
  BUF_X4 U5722 ( .I(n14201), .Z(n33132) );
  INV_X2 U5730 ( .I(n22971), .ZN(n23106) );
  AND2_X1 U5731 ( .A1(n22957), .A2(n5035), .Z(n32037) );
  CLKBUF_X4 U5736 ( .I(n28697), .Z(n30904) );
  NAND2_X1 U5737 ( .A1(n12097), .A2(n32080), .ZN(n32104) );
  AOI21_X1 U5738 ( .A1(n22571), .A2(n28473), .B(n31636), .ZN(n10904) );
  OAI21_X1 U5739 ( .A1(n4100), .A2(n4459), .B(n32344), .ZN(n13983) );
  NAND2_X1 U5744 ( .A1(n32406), .A2(n22663), .ZN(n26404) );
  INV_X1 U5755 ( .I(n22372), .ZN(n33180) );
  INV_X1 U5756 ( .I(n5766), .ZN(n33456) );
  NAND2_X1 U5762 ( .A1(n15812), .A2(n14228), .ZN(n33948) );
  NAND2_X1 U5765 ( .A1(n9546), .A2(n9547), .ZN(n9545) );
  NAND2_X1 U5769 ( .A1(n5960), .A2(n5963), .ZN(n22607) );
  INV_X1 U5770 ( .I(n7848), .ZN(n32344) );
  NAND2_X1 U5775 ( .A1(n22380), .A2(n22388), .ZN(n33753) );
  NOR2_X1 U5778 ( .A1(n32217), .A2(n32216), .ZN(n32215) );
  CLKBUF_X2 U5780 ( .I(n16558), .Z(n29597) );
  CLKBUF_X2 U5783 ( .I(n22491), .Z(n33750) );
  INV_X1 U5785 ( .I(n22600), .ZN(n7633) );
  AOI22_X1 U5786 ( .A1(n7490), .A2(n22359), .B1(n22551), .B2(n22391), .ZN(
        n30112) );
  INV_X2 U5790 ( .I(n11917), .ZN(n31963) );
  NAND2_X1 U5793 ( .A1(n16434), .A2(n22429), .ZN(n22408) );
  CLKBUF_X2 U5794 ( .I(n11892), .Z(n34074) );
  BUF_X2 U5799 ( .I(n622), .Z(n10282) );
  BUF_X2 U5807 ( .I(n11083), .Z(n10612) );
  CLKBUF_X2 U5812 ( .I(n25963), .Z(n34058) );
  INV_X1 U5813 ( .I(n30489), .ZN(n32114) );
  BUF_X2 U5818 ( .I(n6569), .Z(n32753) );
  CLKBUF_X4 U5823 ( .I(n22216), .Z(n34150) );
  INV_X1 U5826 ( .I(n34016), .ZN(n26351) );
  CLKBUF_X1 U5828 ( .I(n22145), .Z(n33072) );
  INV_X1 U5829 ( .I(n22133), .ZN(n32099) );
  INV_X1 U5833 ( .I(n10261), .ZN(n3797) );
  INV_X1 U5834 ( .I(n11458), .ZN(n33160) );
  NAND2_X1 U5835 ( .A1(n28665), .A2(n10689), .ZN(n33667) );
  NAND2_X1 U5839 ( .A1(n33459), .A2(n29552), .ZN(n607) );
  NAND2_X1 U5843 ( .A1(n7947), .A2(n7949), .ZN(n32149) );
  NAND2_X1 U5848 ( .A1(n33908), .A2(n33907), .ZN(n14738) );
  INV_X1 U5850 ( .I(n21622), .ZN(n21623) );
  NAND2_X1 U5855 ( .A1(n3048), .A2(n4097), .ZN(n31871) );
  INV_X1 U5861 ( .I(n26386), .ZN(n21683) );
  AND3_X1 U5864 ( .A1(n21872), .A2(n30832), .A3(n21870), .Z(n30963) );
  BUF_X2 U5867 ( .I(n13884), .Z(n32384) );
  CLKBUF_X2 U5869 ( .I(n1313), .Z(n31317) );
  CLKBUF_X4 U5876 ( .I(n11401), .Z(n7553) );
  NAND2_X1 U5878 ( .A1(n32223), .A2(n21188), .ZN(n10134) );
  INV_X1 U5881 ( .I(n8323), .ZN(n21663) );
  AOI22_X1 U5887 ( .A1(n6826), .A2(n21252), .B1(n9699), .B2(n11792), .ZN(n3924) );
  NAND2_X1 U5888 ( .A1(n21059), .A2(n17984), .ZN(n32521) );
  BUF_X4 U5893 ( .I(n29997), .Z(n32252) );
  NAND2_X1 U5900 ( .A1(n6198), .A2(n32001), .ZN(n33826) );
  NAND2_X1 U5902 ( .A1(n4341), .A2(n2689), .ZN(n34130) );
  CLKBUF_X1 U5905 ( .I(n26622), .Z(n32441) );
  OAI21_X1 U5906 ( .A1(n8393), .A2(n33889), .B(n33979), .ZN(n12690) );
  NAND2_X1 U5911 ( .A1(n32624), .A2(n12325), .ZN(n16198) );
  NAND2_X1 U5918 ( .A1(n31180), .A2(n17731), .ZN(n32815) );
  AND2_X1 U5921 ( .A1(n21253), .A2(n17829), .Z(n11792) );
  OAI21_X1 U5925 ( .A1(n32351), .A2(n32350), .B(n31614), .ZN(n17215) );
  NOR2_X1 U5927 ( .A1(n33684), .A2(n33683), .ZN(n33682) );
  NOR2_X1 U5928 ( .A1(n21284), .A2(n16473), .ZN(n7344) );
  NAND2_X1 U5939 ( .A1(n34121), .A2(n30755), .ZN(n27303) );
  BUF_X2 U5948 ( .I(n10787), .Z(n9518) );
  INV_X1 U5949 ( .I(n32239), .ZN(n13506) );
  BUF_X2 U5950 ( .I(n17144), .Z(n31614) );
  BUF_X2 U5954 ( .I(n8813), .Z(n7690) );
  CLKBUF_X2 U5960 ( .I(n21224), .Z(n5595) );
  OR2_X1 U5965 ( .A1(n15734), .A2(n15733), .Z(n21362) );
  INV_X1 U5966 ( .I(n602), .ZN(n33311) );
  CLKBUF_X4 U5968 ( .I(n8434), .Z(n32452) );
  BUF_X4 U5970 ( .I(n21266), .Z(n31965) );
  CLKBUF_X2 U5976 ( .I(n4858), .Z(n32310) );
  CLKBUF_X2 U5978 ( .I(n20766), .Z(n33969) );
  CLKBUF_X2 U5980 ( .I(n7653), .Z(n32581) );
  INV_X1 U5982 ( .I(n20742), .ZN(n20386) );
  CLKBUF_X2 U5984 ( .I(n20961), .Z(n32749) );
  INV_X1 U5986 ( .I(n7294), .ZN(n33234) );
  INV_X1 U5987 ( .I(n32996), .ZN(n7800) );
  INV_X2 U5989 ( .I(n20913), .ZN(n31966) );
  NOR2_X1 U6013 ( .A1(n33899), .A2(n30952), .ZN(n4909) );
  NOR2_X1 U6018 ( .A1(n28135), .A2(n2203), .ZN(n33899) );
  INV_X1 U6026 ( .I(n33944), .ZN(n34155) );
  NAND2_X1 U6032 ( .A1(n32277), .A2(n2237), .ZN(n32276) );
  NAND2_X1 U6034 ( .A1(n33341), .A2(n31961), .ZN(n19454) );
  INV_X1 U6037 ( .I(n33193), .ZN(n33192) );
  OAI21_X1 U6039 ( .A1(n20216), .A2(n8998), .B(n33639), .ZN(n20218) );
  INV_X1 U6040 ( .I(n9808), .ZN(n33307) );
  CLKBUF_X8 U6047 ( .I(n3086), .Z(n31967) );
  CLKBUF_X8 U6048 ( .I(n29337), .Z(n32504) );
  NOR2_X1 U6049 ( .A1(n20193), .A2(n20192), .ZN(n32939) );
  CLKBUF_X1 U6050 ( .I(n9352), .Z(n34132) );
  INV_X1 U6060 ( .I(n31863), .ZN(n33195) );
  INV_X4 U6066 ( .I(n30504), .ZN(n31968) );
  CLKBUF_X2 U6067 ( .I(n20344), .Z(n34013) );
  CLKBUF_X2 U6070 ( .I(n27697), .Z(n33116) );
  BUF_X2 U6072 ( .I(n7292), .Z(n31811) );
  NAND2_X1 U6073 ( .A1(n34105), .A2(n14479), .ZN(n29920) );
  AOI22_X1 U6074 ( .A1(n30404), .A2(n1035), .B1(n19562), .B2(n11624), .ZN(
        n33249) );
  CLKBUF_X2 U6078 ( .I(n20526), .Z(n33222) );
  AND2_X1 U6081 ( .A1(n29914), .A2(n17497), .Z(n20438) );
  NAND2_X1 U6084 ( .A1(n3790), .A2(n33769), .ZN(n33768) );
  OAI21_X1 U6089 ( .A1(n31988), .A2(n32371), .B(n32416), .ZN(n19839) );
  NAND2_X1 U6097 ( .A1(n19528), .A2(n1617), .ZN(n32740) );
  NAND2_X1 U6099 ( .A1(n6929), .A2(n6930), .ZN(n33896) );
  INV_X4 U6101 ( .I(n7762), .ZN(n31969) );
  NAND2_X1 U6106 ( .A1(n30614), .A2(n4201), .ZN(n33037) );
  NOR2_X1 U6111 ( .A1(n19939), .A2(n32109), .ZN(n5694) );
  BUF_X2 U6113 ( .I(n20110), .Z(n32408) );
  BUF_X1 U6115 ( .I(n13852), .Z(n29233) );
  CLKBUF_X2 U6118 ( .I(n12008), .Z(n34108) );
  BUF_X2 U6119 ( .I(n577), .Z(n27832) );
  CLKBUF_X1 U6131 ( .I(n10426), .Z(n32891) );
  BUF_X2 U6133 ( .I(n11630), .Z(n33419) );
  BUF_X2 U6152 ( .I(n20108), .Z(n16243) );
  CLKBUF_X2 U6157 ( .I(n7896), .Z(n32184) );
  CLKBUF_X2 U6161 ( .I(n33339), .Z(n32809) );
  INV_X1 U6167 ( .I(n19749), .ZN(n32206) );
  BUF_X2 U6170 ( .I(n19494), .Z(n207) );
  NAND2_X1 U6171 ( .A1(n32758), .A2(n13494), .ZN(n9080) );
  OAI21_X1 U6172 ( .A1(n33825), .A2(n26350), .B(n33824), .ZN(n17509) );
  NAND2_X1 U6174 ( .A1(n33231), .A2(n33230), .ZN(n10741) );
  NAND2_X1 U6175 ( .A1(n18360), .A2(n826), .ZN(n32675) );
  NAND2_X1 U6178 ( .A1(n32293), .A2(n32292), .ZN(n13706) );
  NAND2_X1 U6179 ( .A1(n29731), .A2(n29730), .ZN(n32676) );
  NAND2_X1 U6185 ( .A1(n27274), .A2(n27273), .ZN(n33229) );
  NAND2_X1 U6190 ( .A1(n17510), .A2(n26350), .ZN(n33824) );
  INV_X1 U6194 ( .I(n19363), .ZN(n32290) );
  CLKBUF_X2 U6199 ( .I(n30995), .Z(n32788) );
  CLKBUF_X2 U6206 ( .I(n19262), .Z(n33206) );
  OR2_X1 U6210 ( .A1(n1883), .A2(n16699), .Z(n9083) );
  NAND2_X1 U6242 ( .A1(n8662), .A2(n19178), .ZN(n33228) );
  AND2_X1 U6244 ( .A1(n8379), .A2(n2902), .Z(n32060) );
  CLKBUF_X2 U6248 ( .I(n19123), .Z(n27033) );
  CLKBUF_X8 U6252 ( .I(n19314), .Z(n31970) );
  INV_X2 U6254 ( .I(n19021), .ZN(n19288) );
  NAND2_X1 U6258 ( .A1(n15859), .A2(n30116), .ZN(n32720) );
  NAND2_X1 U6275 ( .A1(n18508), .A2(n18509), .ZN(n32439) );
  OR2_X1 U6278 ( .A1(n12648), .A2(n13016), .Z(n13014) );
  NAND2_X1 U6283 ( .A1(n33422), .A2(n33421), .ZN(n27253) );
  NAND2_X1 U6290 ( .A1(n29492), .A2(n18640), .ZN(n8736) );
  NOR2_X1 U6291 ( .A1(n9420), .A2(n14344), .ZN(n32097) );
  AND2_X1 U6292 ( .A1(n13554), .A2(n18510), .Z(n32003) );
  NAND2_X1 U6302 ( .A1(n13016), .A2(n32901), .ZN(n32786) );
  INV_X1 U6312 ( .I(n18726), .ZN(n33422) );
  INV_X1 U6315 ( .I(n17360), .ZN(n33208) );
  INV_X4 U6320 ( .I(n8756), .ZN(n31971) );
  INV_X1 U6332 ( .I(n14666), .ZN(n18516) );
  CLKBUF_X2 U6335 ( .I(n11460), .Z(n33548) );
  BUF_X2 U6338 ( .I(n18831), .Z(n13846) );
  INV_X4 U6342 ( .I(n29315), .ZN(n31972) );
  CLKBUF_X2 U6344 ( .I(n13445), .Z(n33941) );
  INV_X1 U6345 ( .I(n25570), .ZN(n32796) );
  INV_X1 U6346 ( .I(n25929), .ZN(n32130) );
  CLKBUF_X2 U6348 ( .I(n17168), .Z(n9) );
  CLKBUF_X1 U6349 ( .I(n493), .Z(n171) );
  CLKBUF_X2 U6360 ( .I(n18862), .Z(n33205) );
  INV_X1 U6362 ( .I(n24759), .ZN(n33693) );
  NAND2_X1 U6364 ( .A1(n10669), .A2(n18677), .ZN(n10670) );
  INV_X1 U6365 ( .I(n16572), .ZN(n33998) );
  CLKBUF_X2 U6366 ( .I(n18548), .Z(n16122) );
  INV_X1 U6367 ( .I(n18707), .ZN(n18535) );
  NAND2_X1 U6373 ( .A1(n11097), .A2(n882), .ZN(n4070) );
  INV_X2 U6378 ( .I(n12290), .ZN(n3218) );
  CLKBUF_X2 U6384 ( .I(n9930), .Z(n32358) );
  CLKBUF_X1 U6387 ( .I(n29182), .Z(n32143) );
  NOR2_X1 U6400 ( .A1(n8788), .A2(n18714), .ZN(n6590) );
  CLKBUF_X2 U6402 ( .I(n18588), .Z(n28056) );
  NAND2_X1 U6405 ( .A1(n5269), .A2(n18705), .ZN(n4043) );
  CLKBUF_X4 U6406 ( .I(n18373), .Z(n18805) );
  NOR2_X1 U6409 ( .A1(n18722), .A2(n18580), .ZN(n12190) );
  NOR2_X1 U6411 ( .A1(n33310), .A2(n33309), .ZN(n9668) );
  INV_X1 U6413 ( .I(n12074), .ZN(n18609) );
  NAND2_X1 U6415 ( .A1(n18633), .A2(n15888), .ZN(n15841) );
  NOR2_X1 U6416 ( .A1(n11390), .A2(n14926), .ZN(n18659) );
  CLKBUF_X1 U6417 ( .I(n18323), .Z(n18492) );
  NOR2_X1 U6424 ( .A1(n10844), .A2(n959), .ZN(n4267) );
  NAND2_X1 U6425 ( .A1(n9766), .A2(n18797), .ZN(n18796) );
  NAND2_X1 U6434 ( .A1(n13200), .A2(n19180), .ZN(n7751) );
  AOI21_X1 U6436 ( .A1(n31903), .A2(n18563), .B(n6256), .ZN(n18565) );
  AOI21_X1 U6439 ( .A1(n33040), .A2(n18695), .B(n16569), .ZN(n18391) );
  OAI21_X1 U6444 ( .A1(n18318), .A2(n18634), .B(n18711), .ZN(n30175) );
  NAND2_X1 U6449 ( .A1(n19057), .A2(n18994), .ZN(n32182) );
  NAND2_X1 U6460 ( .A1(n32219), .A2(n32218), .ZN(n10192) );
  NAND3_X1 U6461 ( .A1(n19181), .A2(n19178), .A3(n29769), .ZN(n13009) );
  NOR2_X1 U6464 ( .A1(n3784), .A2(n879), .ZN(n32758) );
  INV_X1 U6474 ( .I(n32622), .ZN(n8303) );
  INV_X1 U6477 ( .I(n30781), .ZN(n1056) );
  NAND2_X1 U6480 ( .A1(n28276), .A2(n1630), .ZN(n9442) );
  NAND2_X1 U6482 ( .A1(n19076), .A2(n19288), .ZN(n18360) );
  INV_X2 U6483 ( .I(n16093), .ZN(n1052) );
  INV_X1 U6484 ( .I(n14892), .ZN(n18995) );
  NOR2_X1 U6487 ( .A1(n19091), .A2(n19088), .ZN(n31174) );
  INV_X2 U6494 ( .I(n19258), .ZN(n744) );
  NOR2_X1 U6499 ( .A1(n19198), .A2(n26417), .ZN(n13891) );
  INV_X1 U6507 ( .I(n19103), .ZN(n11713) );
  NOR2_X1 U6511 ( .A1(n32932), .A2(n7492), .ZN(n17677) );
  AOI21_X1 U6512 ( .A1(n14625), .A2(n8379), .B(n2901), .ZN(n12850) );
  CLKBUF_X2 U6515 ( .I(n14812), .Z(n12549) );
  OAI21_X1 U6521 ( .A1(n19148), .A2(n19147), .B(n19150), .ZN(n18267) );
  OAI22_X1 U6526 ( .A1(n18475), .A2(n16185), .B1(n18901), .B2(n4), .ZN(n18476)
         );
  NAND2_X1 U6529 ( .A1(n6578), .A2(n6577), .ZN(n6576) );
  INV_X1 U6534 ( .I(n19520), .ZN(n10026) );
  INV_X1 U6538 ( .I(n6731), .ZN(n11320) );
  NAND2_X1 U6544 ( .A1(n14736), .A2(n14130), .ZN(n14735) );
  CLKBUF_X2 U6545 ( .I(n14094), .Z(n32286) );
  NOR2_X1 U6550 ( .A1(n33712), .A2(n33389), .ZN(n11581) );
  INV_X1 U6553 ( .I(n15787), .ZN(n29090) );
  CLKBUF_X1 U6557 ( .I(n5150), .Z(n32918) );
  INV_X1 U6560 ( .I(n26300), .ZN(n19722) );
  INV_X1 U6574 ( .I(n19466), .ZN(n17342) );
  INV_X1 U6577 ( .I(n19542), .ZN(n32231) );
  INV_X1 U6582 ( .I(n2362), .ZN(n12796) );
  INV_X1 U6583 ( .I(n31922), .ZN(n8292) );
  NOR2_X1 U6588 ( .A1(n13591), .A2(n11198), .ZN(n19828) );
  INV_X1 U6591 ( .I(n19746), .ZN(n30435) );
  INV_X1 U6592 ( .I(n11052), .ZN(n2679) );
  NAND2_X1 U6596 ( .A1(n34103), .A2(n6532), .ZN(n13657) );
  NAND2_X1 U6600 ( .A1(n20056), .A2(n32326), .ZN(n14099) );
  NAND2_X1 U6604 ( .A1(n32746), .A2(n32745), .ZN(n19977) );
  NAND2_X1 U6605 ( .A1(n19833), .A2(n1169), .ZN(n15174) );
  INV_X1 U6606 ( .I(n579), .ZN(n7461) );
  NOR2_X1 U6609 ( .A1(n27491), .A2(n19961), .ZN(n20128) );
  INV_X1 U6612 ( .I(n1361), .ZN(n9749) );
  INV_X1 U6614 ( .I(n1169), .ZN(n15593) );
  NOR2_X1 U6616 ( .A1(n27808), .A2(n20113), .ZN(n14729) );
  NOR2_X1 U6628 ( .A1(n29216), .A2(n19990), .ZN(n34106) );
  INV_X1 U6629 ( .I(n9106), .ZN(n31106) );
  CLKBUF_X2 U6631 ( .I(n20108), .Z(n33848) );
  NOR2_X1 U6638 ( .A1(n20097), .A2(n1041), .ZN(n30693) );
  INV_X1 U6639 ( .I(n20054), .ZN(n11893) );
  CLKBUF_X4 U6641 ( .I(n14458), .Z(n14281) );
  CLKBUF_X4 U6642 ( .I(n11333), .Z(n28293) );
  NAND2_X1 U6643 ( .A1(n20104), .A2(n873), .ZN(n15177) );
  NOR3_X1 U6649 ( .A1(n19724), .A2(n16461), .A3(n1042), .ZN(n30357) );
  INV_X1 U6652 ( .I(n19885), .ZN(n19799) );
  NAND2_X1 U6655 ( .A1(n29153), .A2(n576), .ZN(n9171) );
  CLKBUF_X4 U6656 ( .I(n16625), .Z(n29156) );
  INV_X2 U6659 ( .I(n16694), .ZN(n1360) );
  OAI21_X1 U6660 ( .A1(n4674), .A2(n6200), .B(n6263), .ZN(n3090) );
  CLKBUF_X4 U6678 ( .I(n18089), .Z(n161) );
  NAND2_X1 U6682 ( .A1(n33569), .A2(n17945), .ZN(n32673) );
  NAND2_X1 U6689 ( .A1(n9031), .A2(n1042), .ZN(n19941) );
  OAI21_X1 U6690 ( .A1(n27788), .A2(n27787), .B(n20157), .ZN(n30996) );
  NAND2_X1 U6691 ( .A1(n28685), .A2(n28684), .ZN(n28683) );
  AOI21_X1 U6692 ( .A1(n938), .A2(n20052), .B(n939), .ZN(n6929) );
  NAND2_X1 U6694 ( .A1(n8181), .A2(n16630), .ZN(n32775) );
  OAI21_X1 U6700 ( .A1(n20053), .A2(n1361), .B(n8616), .ZN(n15312) );
  INV_X1 U6709 ( .I(n10752), .ZN(n33525) );
  AOI21_X1 U6710 ( .A1(n27714), .A2(n27716), .B(n30355), .ZN(n26784) );
  OAI21_X1 U6731 ( .A1(n19950), .A2(n17363), .B(n729), .ZN(n14) );
  NAND2_X1 U6733 ( .A1(n295), .A2(n1155), .ZN(n20337) );
  INV_X1 U6734 ( .I(n20267), .ZN(n14863) );
  NAND2_X1 U6742 ( .A1(n31242), .A2(n15551), .ZN(n11505) );
  NOR2_X1 U6747 ( .A1(n20607), .A2(n20460), .ZN(n20396) );
  INV_X1 U6749 ( .I(n20410), .ZN(n28128) );
  NAND2_X1 U6754 ( .A1(n8903), .A2(n8870), .ZN(n4586) );
  NAND2_X1 U6755 ( .A1(n4807), .A2(n20571), .ZN(n29077) );
  NOR2_X1 U6756 ( .A1(n33091), .A2(n20545), .ZN(n13629) );
  CLKBUF_X4 U6757 ( .I(n20503), .Z(n28376) );
  NAND2_X1 U6761 ( .A1(n7242), .A2(n20228), .ZN(n20227) );
  INV_X1 U6764 ( .I(n19956), .ZN(n10380) );
  NOR2_X1 U6765 ( .A1(n20489), .A2(n33307), .ZN(n17897) );
  NAND3_X1 U6776 ( .A1(n26567), .A2(n3462), .A3(n741), .ZN(n19453) );
  CLKBUF_X2 U6778 ( .I(n7280), .Z(n32481) );
  AOI22_X1 U6779 ( .A1(n20251), .A2(n20510), .B1(n20509), .B2(n20435), .ZN(
        n17974) );
  NAND2_X1 U6782 ( .A1(n5471), .A2(n14179), .ZN(n20376) );
  INV_X1 U6785 ( .I(n9986), .ZN(n5589) );
  OAI21_X1 U6786 ( .A1(n20366), .A2(n7577), .B(n33843), .ZN(n20367) );
  NOR2_X1 U6788 ( .A1(n17329), .A2(n6531), .ZN(n9774) );
  INV_X2 U6789 ( .I(n15005), .ZN(n1352) );
  INV_X2 U6800 ( .I(n31533), .ZN(n30869) );
  NAND2_X1 U6805 ( .A1(n13629), .A2(n20335), .ZN(n13628) );
  NAND2_X1 U6806 ( .A1(n20297), .A2(n14836), .ZN(n14835) );
  NAND3_X1 U6810 ( .A1(n3944), .A2(n17975), .A3(n1355), .ZN(n14471) );
  NAND2_X1 U6813 ( .A1(n16004), .A2(n13786), .ZN(n13782) );
  INV_X1 U6814 ( .I(n20900), .ZN(n29167) );
  OAI21_X1 U6819 ( .A1(n11303), .A2(n1156), .B(n6616), .ZN(n20636) );
  NAND2_X1 U6823 ( .A1(n19454), .A2(n19453), .ZN(n3307) );
  INV_X1 U6825 ( .I(n12258), .ZN(n31860) );
  AOI21_X1 U6826 ( .A1(n29623), .A2(n1352), .B(n20419), .ZN(n20421) );
  NAND2_X1 U6828 ( .A1(n5781), .A2(n17497), .ZN(n19956) );
  CLKBUF_X1 U6839 ( .I(n21044), .Z(n30240) );
  INV_X1 U6840 ( .I(n20860), .ZN(n12671) );
  CLKBUF_X2 U6843 ( .I(n20680), .Z(n31233) );
  CLKBUF_X4 U6844 ( .I(n13864), .Z(n28315) );
  INV_X1 U6845 ( .I(n21025), .ZN(n8138) );
  INV_X1 U6849 ( .I(n17440), .ZN(n33085) );
  INV_X1 U6851 ( .I(n30492), .ZN(n20855) );
  INV_X1 U6853 ( .I(n28981), .ZN(n33892) );
  CLKBUF_X1 U6858 ( .I(n13189), .Z(n28400) );
  INV_X2 U6859 ( .I(n16526), .ZN(n31729) );
  NAND2_X1 U6860 ( .A1(n12037), .A2(n21270), .ZN(n27270) );
  NAND2_X1 U6872 ( .A1(n2738), .A2(n9133), .ZN(n8792) );
  INV_X2 U6881 ( .I(n28287), .ZN(n14563) );
  INV_X1 U6882 ( .I(n21210), .ZN(n16743) );
  NAND2_X1 U6889 ( .A1(n1022), .A2(n33684), .ZN(n7757) );
  NOR2_X1 U6902 ( .A1(n21085), .A2(n4755), .ZN(n29750) );
  CLKBUF_X2 U6904 ( .I(n13989), .Z(n32242) );
  INV_X2 U6913 ( .I(n11814), .ZN(n13692) );
  OAI21_X1 U6916 ( .A1(n33106), .A2(n21109), .B(n33705), .ZN(n10922) );
  NAND3_X1 U6920 ( .A1(n32357), .A2(n17767), .A3(n21078), .ZN(n26018) );
  NAND2_X1 U6921 ( .A1(n30646), .A2(n14721), .ZN(n17101) );
  NAND2_X1 U6922 ( .A1(n21379), .A2(n17313), .ZN(n2275) );
  NAND2_X1 U6925 ( .A1(n16668), .A2(n13896), .ZN(n15219) );
  NOR2_X1 U6927 ( .A1(n13896), .A2(n21115), .ZN(n29001) );
  NOR2_X1 U6930 ( .A1(n20879), .A2(n20880), .ZN(n29739) );
  INV_X1 U6933 ( .I(n929), .ZN(n33454) );
  INV_X1 U6939 ( .I(n11942), .ZN(n21431) );
  NOR2_X1 U6941 ( .A1(n20941), .A2(n16629), .ZN(n32980) );
  NAND2_X1 U6942 ( .A1(n13022), .A2(n32647), .ZN(n16117) );
  NAND2_X1 U6944 ( .A1(n20945), .A2(n27503), .ZN(n21183) );
  CLKBUF_X4 U6945 ( .I(n17731), .Z(n33972) );
  NAND2_X1 U6946 ( .A1(n21129), .A2(n21443), .ZN(n32454) );
  NOR2_X1 U6948 ( .A1(n21109), .A2(n1632), .ZN(n5488) );
  NAND2_X1 U6950 ( .A1(n14230), .A2(n21440), .ZN(n34083) );
  NAND2_X1 U6956 ( .A1(n27303), .A2(n27305), .ZN(n26903) );
  NOR2_X1 U6961 ( .A1(n6584), .A2(n9721), .ZN(n14997) );
  NAND2_X1 U6962 ( .A1(n7845), .A2(n1333), .ZN(n4179) );
  NOR2_X1 U6963 ( .A1(n27193), .A2(n32239), .ZN(n6879) );
  NOR2_X1 U6970 ( .A1(n11487), .A2(n33682), .ZN(n31848) );
  NOR2_X1 U6971 ( .A1(n11215), .A2(n28922), .ZN(n28921) );
  OAI22_X1 U6975 ( .A1(n10149), .A2(n3673), .B1(n2275), .B2(n7007), .ZN(n31215) );
  NAND2_X1 U6976 ( .A1(n21411), .A2(n5039), .ZN(n2721) );
  NOR2_X1 U6980 ( .A1(n33417), .A2(n33418), .ZN(n32116) );
  OR3_X1 U6983 ( .A1(n4683), .A2(n16639), .A3(n29255), .Z(n34158) );
  NOR2_X1 U6985 ( .A1(n4517), .A2(n21251), .ZN(n4284) );
  OAI21_X1 U6987 ( .A1(n21259), .A2(n16652), .B(n8757), .ZN(n6568) );
  INV_X2 U6989 ( .I(n16519), .ZN(n3048) );
  NOR2_X1 U6991 ( .A1(n17348), .A2(n32252), .ZN(n3703) );
  NOR2_X1 U6993 ( .A1(n15302), .A2(n15296), .ZN(n10875) );
  NOR2_X1 U6994 ( .A1(n338), .A2(n4234), .ZN(n4391) );
  INV_X2 U6996 ( .I(n16668), .ZN(n4989) );
  OAI22_X1 U6998 ( .A1(n21586), .A2(n32252), .B1(n3680), .B2(n26337), .ZN(
        n29595) );
  NOR2_X1 U7002 ( .A1(n21659), .A2(n8784), .ZN(n4117) );
  NAND2_X1 U7003 ( .A1(n29434), .A2(n517), .ZN(n21747) );
  NOR2_X1 U7004 ( .A1(n7969), .A2(n7182), .ZN(n7183) );
  INV_X1 U7008 ( .I(n21687), .ZN(n21514) );
  NOR2_X1 U7010 ( .A1(n5546), .A2(n4356), .ZN(n8705) );
  NAND2_X1 U7012 ( .A1(n5546), .A2(n14236), .ZN(n21622) );
  NAND3_X1 U7019 ( .A1(n30479), .A2(n21850), .A3(n21763), .ZN(n10968) );
  NAND2_X1 U7020 ( .A1(n21585), .A2(n15302), .ZN(n21234) );
  AOI21_X1 U7024 ( .A1(n4391), .A2(n13816), .B(n27816), .ZN(n6076) );
  INV_X1 U7035 ( .I(n8753), .ZN(n10456) );
  CLKBUF_X2 U7039 ( .I(n28762), .Z(n33468) );
  NAND3_X1 U7041 ( .A1(n32321), .A2(n21830), .A3(n32320), .ZN(n34001) );
  CLKBUF_X1 U7045 ( .I(n21789), .Z(n27543) );
  NOR2_X1 U7049 ( .A1(n16796), .A2(n16192), .ZN(n22126) );
  AOI21_X1 U7052 ( .A1(n2217), .A2(n16600), .B(n21772), .ZN(n12328) );
  NAND3_X1 U7055 ( .A1(n864), .A2(n15864), .A3(n12278), .ZN(n12277) );
  INV_X1 U7057 ( .I(n10205), .ZN(n30407) );
  CLKBUF_X2 U7058 ( .I(n22227), .Z(n33509) );
  NAND3_X1 U7063 ( .A1(n11657), .A2(n11656), .A3(n14829), .ZN(n17898) );
  AOI21_X1 U7068 ( .A1(n4311), .A2(n6489), .B(n4310), .ZN(n21624) );
  INV_X1 U7070 ( .I(n22000), .ZN(n21875) );
  INV_X1 U7073 ( .I(n6571), .ZN(n33707) );
  INV_X1 U7078 ( .I(n9267), .ZN(n11422) );
  INV_X1 U7079 ( .I(n9914), .ZN(n32696) );
  INV_X1 U7091 ( .I(n26933), .ZN(n32155) );
  NAND2_X1 U7097 ( .A1(n31701), .A2(n10282), .ZN(n32797) );
  INV_X1 U7099 ( .I(n15260), .ZN(n30669) );
  NOR2_X1 U7100 ( .A1(n31001), .A2(n26708), .ZN(n22342) );
  INV_X1 U7101 ( .I(n22487), .ZN(n1288) );
  INV_X1 U7104 ( .I(n17204), .ZN(n22644) );
  OAI21_X1 U7108 ( .A1(n9910), .A2(n29158), .B(n33237), .ZN(n31838) );
  CLKBUF_X2 U7110 ( .I(n29263), .Z(n355) );
  CLKBUF_X4 U7111 ( .I(n1805), .Z(n1633) );
  NOR2_X1 U7116 ( .A1(n1294), .A2(n14253), .ZN(n22594) );
  INV_X1 U7117 ( .I(n22622), .ZN(n995) );
  INV_X1 U7121 ( .I(n22491), .ZN(n17302) );
  AOI21_X1 U7125 ( .A1(n16745), .A2(n8919), .B(n32080), .ZN(n8918) );
  NOR2_X1 U7126 ( .A1(n22660), .A2(n809), .ZN(n30334) );
  CLKBUF_X1 U7127 ( .I(n17518), .Z(n14493) );
  CLKBUF_X2 U7130 ( .I(n22332), .Z(n33964) );
  CLKBUF_X4 U7131 ( .I(n8275), .Z(n1116) );
  NAND2_X1 U7133 ( .A1(n26098), .A2(n1127), .ZN(n13193) );
  NAND2_X1 U7137 ( .A1(n22460), .A2(n16137), .ZN(n22344) );
  NAND2_X1 U7138 ( .A1(n27880), .A2(n28312), .ZN(n33945) );
  INV_X1 U7145 ( .I(n12952), .ZN(n22511) );
  INV_X1 U7150 ( .I(n32448), .ZN(n1720) );
  NAND2_X1 U7151 ( .A1(n16884), .A2(n22336), .ZN(n26813) );
  OAI22_X1 U7158 ( .A1(n11419), .A2(n22420), .B1(n31345), .B2(n11420), .ZN(
        n3934) );
  NAND2_X1 U7164 ( .A1(n13524), .A2(n12840), .ZN(n32518) );
  CLKBUF_X2 U7169 ( .I(n16332), .Z(n27402) );
  OAI22_X1 U7173 ( .A1(n32680), .A2(n11629), .B1(n30205), .B2(n15581), .ZN(
        n2135) );
  INV_X1 U7175 ( .I(n10206), .ZN(n8801) );
  NAND2_X1 U7177 ( .A1(n32955), .A2(n29495), .ZN(n1580) );
  AOI22_X1 U7180 ( .A1(n22688), .A2(n22332), .B1(n2417), .B2(n12733), .ZN(
        n27034) );
  INV_X2 U7181 ( .I(n636), .ZN(n857) );
  NAND2_X1 U7189 ( .A1(n32823), .A2(n31963), .ZN(n27368) );
  NAND2_X1 U7193 ( .A1(n22475), .A2(n22377), .ZN(n31143) );
  INV_X2 U7198 ( .I(n10862), .ZN(n8912) );
  CLKBUF_X2 U7200 ( .I(n30868), .Z(n32967) );
  NAND3_X1 U7206 ( .A1(n903), .A2(n30564), .A3(n7848), .ZN(n29722) );
  INV_X1 U7209 ( .I(n2635), .ZN(n11298) );
  INV_X1 U7213 ( .I(n31566), .ZN(n33591) );
  OAI22_X1 U7216 ( .A1(n30455), .A2(n9954), .B1(n773), .B2(n6782), .ZN(n10280)
         );
  AOI22_X1 U7218 ( .A1(n22651), .A2(n4916), .B1(n22433), .B2(n14251), .ZN(
        n1661) );
  INV_X4 U7231 ( .I(n27090), .ZN(n22774) );
  INV_X2 U7232 ( .I(n17147), .ZN(n5597) );
  INV_X1 U7233 ( .I(n14978), .ZN(n22756) );
  INV_X1 U7236 ( .I(n3296), .ZN(n33388) );
  CLKBUF_X4 U7238 ( .I(n12729), .Z(n28314) );
  NAND2_X1 U7243 ( .A1(n32704), .A2(n15718), .ZN(n18239) );
  NOR2_X1 U7244 ( .A1(n4750), .A2(n30234), .ZN(n11540) );
  NAND2_X1 U7245 ( .A1(n31937), .A2(n15501), .ZN(n6350) );
  NAND2_X1 U7248 ( .A1(n7004), .A2(n22971), .ZN(n22805) );
  NOR2_X1 U7249 ( .A1(n23112), .A2(n23111), .ZN(n32525) );
  INV_X1 U7252 ( .I(n2449), .ZN(n23031) );
  NAND2_X1 U7253 ( .A1(n641), .A2(n22876), .ZN(n22766) );
  NAND2_X1 U7258 ( .A1(n6800), .A2(n1107), .ZN(n12742) );
  OAI21_X1 U7260 ( .A1(n28408), .A2(n6799), .B(n1107), .ZN(n6035) );
  NOR2_X1 U7262 ( .A1(n4750), .A2(n22919), .ZN(n10588) );
  INV_X1 U7266 ( .I(n28934), .ZN(n22908) );
  NAND2_X1 U7269 ( .A1(n6874), .A2(n2449), .ZN(n6942) );
  NAND2_X1 U7271 ( .A1(n31225), .A2(n15421), .ZN(n22383) );
  CLKBUF_X4 U7277 ( .I(n4208), .Z(n30960) );
  AOI21_X1 U7278 ( .A1(n30904), .A2(n28659), .B(n10360), .ZN(n5571) );
  INV_X1 U7279 ( .I(n23183), .ZN(n23241) );
  CLKBUF_X2 U7284 ( .I(n23209), .Z(n34100) );
  INV_X1 U7291 ( .I(n33971), .ZN(n1263) );
  OAI22_X1 U7292 ( .A1(n33996), .A2(n34097), .B1(n22938), .B2(n29173), .ZN(
        n16922) );
  INV_X1 U7296 ( .I(n16998), .ZN(n30362) );
  AOI22_X1 U7299 ( .A1(n26195), .A2(n10296), .B1(n32092), .B2(n30234), .ZN(
        n10759) );
  INV_X1 U7305 ( .I(n22867), .ZN(n33811) );
  CLKBUF_X2 U7307 ( .I(n5512), .Z(n33380) );
  NAND2_X1 U7311 ( .A1(n8381), .A2(n5211), .ZN(n10349) );
  OAI21_X1 U7312 ( .A1(n28970), .A2(n32868), .B(n3160), .ZN(n3159) );
  INV_X1 U7314 ( .I(n11249), .ZN(n32302) );
  INV_X1 U7315 ( .I(n4047), .ZN(n13888) );
  INV_X1 U7319 ( .I(n23153), .ZN(n33590) );
  NOR2_X1 U7326 ( .A1(n23938), .A2(n662), .ZN(n27266) );
  NOR2_X1 U7327 ( .A1(n23951), .A2(n16431), .ZN(n3759) );
  NOR2_X1 U7329 ( .A1(n23691), .A2(n23857), .ZN(n23570) );
  CLKBUF_X4 U7330 ( .I(n17285), .Z(n14975) );
  NAND2_X1 U7338 ( .A1(n27266), .A2(n23939), .ZN(n33626) );
  INV_X1 U7342 ( .I(n23706), .ZN(n33461) );
  INV_X1 U7343 ( .I(n10772), .ZN(n9328) );
  OAI21_X1 U7344 ( .A1(n23933), .A2(n29269), .B(n23527), .ZN(n13103) );
  BUF_X2 U7353 ( .I(n8270), .Z(n32602) );
  INV_X1 U7355 ( .I(n12104), .ZN(n33252) );
  NOR2_X1 U7358 ( .A1(n11392), .A2(n23653), .ZN(n6992) );
  NAND2_X1 U7362 ( .A1(n23777), .A2(n23778), .ZN(n32972) );
  NOR2_X1 U7367 ( .A1(n23858), .A2(n2023), .ZN(n1875) );
  INV_X1 U7370 ( .I(n651), .ZN(n977) );
  INV_X1 U7372 ( .I(n16686), .ZN(n1250) );
  NOR2_X1 U7374 ( .A1(n4743), .A2(n23638), .ZN(n18054) );
  INV_X2 U7375 ( .I(n18204), .ZN(n28265) );
  NAND2_X1 U7378 ( .A1(n23569), .A2(n23914), .ZN(n32843) );
  AOI21_X1 U7381 ( .A1(n13521), .A2(n29271), .B(n23795), .ZN(n16212) );
  INV_X1 U7382 ( .I(n32986), .ZN(n23915) );
  OAI21_X1 U7384 ( .A1(n23776), .A2(n31810), .B(n23775), .ZN(n23654) );
  NAND2_X1 U7392 ( .A1(n1099), .A2(n23755), .ZN(n14943) );
  NOR2_X1 U7393 ( .A1(n11589), .A2(n16424), .ZN(n33786) );
  CLKBUF_X1 U7402 ( .I(n666), .Z(n28365) );
  CLKBUF_X4 U7404 ( .I(n10187), .Z(n29198) );
  INV_X1 U7410 ( .I(n23867), .ZN(n23637) );
  INV_X1 U7412 ( .I(n23906), .ZN(n17288) );
  OAI22_X1 U7415 ( .A1(n10384), .A2(n16388), .B1(n2460), .B2(n11240), .ZN(
        n10382) );
  INV_X1 U7420 ( .I(n8547), .ZN(n1252) );
  NOR2_X1 U7428 ( .A1(n23826), .A2(n29839), .ZN(n8472) );
  NAND2_X1 U7431 ( .A1(n23939), .A2(n33499), .ZN(n30828) );
  NAND2_X1 U7433 ( .A1(n24095), .A2(n14195), .ZN(n1619) );
  OAI21_X1 U7442 ( .A1(n11708), .A2(n6272), .B(n4111), .ZN(n23671) );
  OAI22_X1 U7444 ( .A1(n23760), .A2(n26115), .B1(n23759), .B2(n13905), .ZN(
        n32336) );
  CLKBUF_X4 U7445 ( .I(n11516), .Z(n1920) );
  INV_X1 U7446 ( .I(n29370), .ZN(n33603) );
  NOR2_X1 U7449 ( .A1(n23773), .A2(n23775), .ZN(n16628) );
  NAND2_X1 U7451 ( .A1(n23961), .A2(n13343), .ZN(n6336) );
  CLKBUF_X4 U7453 ( .I(n10302), .Z(n6001) );
  NAND2_X1 U7456 ( .A1(n24204), .A2(n7935), .ZN(n9202) );
  NAND2_X1 U7459 ( .A1(n24114), .A2(n24283), .ZN(n23549) );
  CLKBUF_X1 U7466 ( .I(n30191), .Z(n32520) );
  NOR2_X1 U7467 ( .A1(n13378), .A2(n2558), .ZN(n4664) );
  INV_X2 U7469 ( .I(n6476), .ZN(n24253) );
  NAND3_X1 U7473 ( .A1(n8086), .A2(n24209), .A3(n8165), .ZN(n17676) );
  AOI21_X1 U7481 ( .A1(n24125), .A2(n24124), .B(n24182), .ZN(n24126) );
  OAI21_X1 U7484 ( .A1(n24176), .A2(n11200), .B(n17566), .ZN(n24179) );
  INV_X1 U7487 ( .I(n24568), .ZN(n30127) );
  NAND2_X1 U7491 ( .A1(n3549), .A2(n16573), .ZN(n2361) );
  NAND3_X1 U7492 ( .A1(n13660), .A2(n11937), .A3(n24198), .ZN(n32870) );
  NAND2_X1 U7494 ( .A1(n11439), .A2(n11440), .ZN(n24776) );
  INV_X1 U7500 ( .I(n18144), .ZN(n33028) );
  CLKBUF_X2 U7501 ( .I(n24811), .Z(n32814) );
  CLKBUF_X2 U7502 ( .I(n3694), .Z(n32623) );
  INV_X1 U7503 ( .I(n8152), .ZN(n24450) );
  INV_X1 U7513 ( .I(n24525), .ZN(n33090) );
  NAND2_X1 U7516 ( .A1(n4886), .A2(n32760), .ZN(n10629) );
  NAND2_X1 U7517 ( .A1(n5254), .A2(n11045), .ZN(n5273) );
  INV_X1 U7522 ( .I(n15318), .ZN(n29630) );
  INV_X1 U7527 ( .I(n25565), .ZN(n6071) );
  INV_X1 U7528 ( .I(n10248), .ZN(n13532) );
  NAND2_X1 U7529 ( .A1(n32878), .A2(n4885), .ZN(n10890) );
  INV_X1 U7530 ( .I(n25887), .ZN(n5553) );
  NOR2_X1 U7535 ( .A1(n25013), .A2(n24977), .ZN(n6364) );
  CLKBUF_X2 U7540 ( .I(n4885), .Z(n32106) );
  NAND2_X1 U7541 ( .A1(n25582), .A2(n11900), .ZN(n8712) );
  OAI22_X1 U7544 ( .A1(n25411), .A2(n752), .B1(n25412), .B2(n11366), .ZN(n1463) );
  CLKBUF_X2 U7545 ( .I(n11957), .Z(n33976) );
  CLKBUF_X4 U7546 ( .I(n24181), .Z(n25897) );
  NAND2_X1 U7547 ( .A1(n32590), .A2(n25889), .ZN(n32589) );
  INV_X1 U7548 ( .I(n24977), .ZN(n14993) );
  NAND2_X1 U7554 ( .A1(n25200), .A2(n12476), .ZN(n17928) );
  NAND3_X1 U7555 ( .A1(n1213), .A2(n25239), .A3(n14922), .ZN(n31545) );
  INV_X1 U7558 ( .I(n28096), .ZN(n25713) );
  INV_X1 U7560 ( .I(n17814), .ZN(n25904) );
  NOR2_X1 U7561 ( .A1(n25897), .A2(n9932), .ZN(n10136) );
  NAND2_X1 U7564 ( .A1(n27262), .A2(n10504), .ZN(n30656) );
  OAI21_X1 U7566 ( .A1(n32668), .A2(n32667), .B(n7081), .ZN(n28117) );
  AOI21_X1 U7568 ( .A1(n25866), .A2(n25889), .B(n1214), .ZN(n6851) );
  BUF_X1 U7571 ( .I(n12676), .Z(n33904) );
  NOR2_X1 U7572 ( .A1(n27757), .A2(n27758), .ZN(n33987) );
  CLKBUF_X2 U7574 ( .I(n25385), .Z(n6551) );
  NAND2_X1 U7578 ( .A1(n32825), .A2(n25866), .ZN(n32312) );
  NAND3_X1 U7580 ( .A1(n9495), .A2(n29331), .A3(n13640), .ZN(n26992) );
  INV_X2 U7591 ( .I(n7554), .ZN(n14810) );
  NAND2_X1 U7594 ( .A1(n12864), .A2(n13483), .ZN(n6391) );
  INV_X1 U7597 ( .I(n965), .ZN(n24946) );
  INV_X1 U7601 ( .I(n1209), .ZN(n33400) );
  NAND2_X1 U7604 ( .A1(n13124), .A2(n789), .ZN(n5786) );
  NOR2_X1 U7608 ( .A1(n25127), .A2(n1075), .ZN(n14638) );
  OAI22_X1 U7612 ( .A1(n25272), .A2(n28532), .B1(n25271), .B2(n30281), .ZN(
        n25273) );
  NAND2_X1 U7615 ( .A1(n25041), .A2(n25052), .ZN(n25048) );
  OAI21_X1 U7619 ( .A1(n25041), .A2(n25029), .B(n25060), .ZN(n25035) );
  BUF_X2 U7620 ( .I(Key[6]), .Z(n25832) );
  AOI21_X1 U7623 ( .A1(n5072), .A2(n24994), .B(n964), .ZN(n14318) );
  INV_X1 U7627 ( .I(n25418), .ZN(n33946) );
  INV_X1 U7629 ( .I(n13684), .ZN(n1076) );
  CLKBUF_X1 U7634 ( .I(Key[143]), .Z(n25801) );
  CLKBUF_X1 U7635 ( .I(Key[179]), .Z(n24937) );
  AOI21_X1 U7639 ( .A1(n2265), .A2(n714), .B(n2263), .ZN(n2262) );
  INV_X1 U7648 ( .I(n16525), .ZN(n17914) );
  AND2_X1 U7651 ( .A1(n15804), .A2(n13329), .Z(n31973) );
  AND2_X2 U7675 ( .A1(n11090), .A2(n11900), .Z(n31974) );
  AND2_X1 U7678 ( .A1(n32341), .A2(n20603), .Z(n31976) );
  OR2_X1 U7681 ( .A1(n24974), .A2(n11898), .Z(n31977) );
  AND2_X2 U7682 ( .A1(n29322), .A2(n14095), .Z(n31978) );
  AND3_X2 U7686 ( .A1(n32592), .A2(n32591), .A3(n32589), .Z(n31979) );
  AND2_X2 U7687 ( .A1(n29182), .A2(n18727), .Z(n31980) );
  OR3_X1 U7689 ( .A1(n9066), .A2(n12982), .A3(n24309), .Z(n31983) );
  AND2_X1 U7691 ( .A1(n1099), .A2(n27799), .Z(n31984) );
  AND2_X2 U7694 ( .A1(n29308), .A2(n29315), .Z(n31987) );
  AND2_X1 U7695 ( .A1(n20136), .A2(n19834), .Z(n31988) );
  AND2_X1 U7696 ( .A1(n3687), .A2(n32602), .Z(n31990) );
  AND2_X1 U7698 ( .A1(n19262), .A2(n19257), .Z(n31992) );
  AND2_X2 U7702 ( .A1(n16694), .A2(n19942), .Z(n31993) );
  AND2_X1 U7703 ( .A1(n25403), .A2(n16650), .Z(n31994) );
  AND2_X1 U7704 ( .A1(n6408), .A2(n16906), .Z(n31995) );
  AND2_X1 U7705 ( .A1(n7969), .A2(n31960), .Z(n31996) );
  OR2_X1 U7709 ( .A1(n14976), .A2(n149), .Z(n31998) );
  AND2_X1 U7713 ( .A1(n21251), .A2(n21249), .Z(n31999) );
  AND2_X1 U7715 ( .A1(n10947), .A2(n13747), .Z(n32000) );
  OR2_X1 U7716 ( .A1(n29574), .A2(n21303), .Z(n32001) );
  AND2_X1 U7718 ( .A1(n10295), .A2(n11317), .Z(n32002) );
  OR2_X2 U7719 ( .A1(n16732), .A2(n16854), .Z(n32005) );
  OR2_X1 U7720 ( .A1(n846), .A2(n16467), .Z(n32006) );
  OR2_X1 U7723 ( .A1(n28263), .A2(n907), .Z(n32007) );
  OR2_X1 U7724 ( .A1(n11392), .A2(n1252), .Z(n32008) );
  AND2_X1 U7726 ( .A1(n15421), .A2(n16078), .Z(n32010) );
  OR2_X2 U7732 ( .A1(n29334), .A2(n4886), .Z(n32012) );
  AND2_X1 U7734 ( .A1(n913), .A2(n13332), .Z(n32013) );
  OR2_X2 U7735 ( .A1(n3005), .A2(n8616), .Z(n32014) );
  XNOR2_X1 U7742 ( .A1(n23358), .A2(n25519), .ZN(n32015) );
  OR2_X1 U7746 ( .A1(n24125), .A2(n10381), .Z(n32016) );
  AND3_X1 U7747 ( .A1(n9934), .A2(n9962), .A3(n24201), .Z(n32017) );
  AND2_X1 U7750 ( .A1(n29314), .A2(n31867), .Z(n32018) );
  AND2_X1 U7751 ( .A1(n23881), .A2(n8544), .Z(n32019) );
  OR2_X2 U7752 ( .A1(n22491), .A2(n645), .Z(n32021) );
  XNOR2_X1 U7753 ( .A1(n33749), .A2(n1396), .ZN(n32022) );
  AND2_X1 U7754 ( .A1(n10252), .A2(n752), .Z(n32023) );
  XNOR2_X1 U7755 ( .A1(n14952), .A2(n24426), .ZN(n32024) );
  XNOR2_X1 U7768 ( .A1(n20786), .A2(n1393), .ZN(n32025) );
  XNOR2_X1 U7769 ( .A1(n14120), .A2(n16622), .ZN(n32026) );
  XOR2_X1 U7772 ( .A1(n29885), .A2(n16655), .Z(n32027) );
  OR2_X1 U7773 ( .A1(n2522), .A2(n15322), .Z(n32031) );
  OR2_X2 U7774 ( .A1(n7292), .A2(n20460), .Z(n32033) );
  XNOR2_X1 U7779 ( .A1(Plaintext[50]), .A2(Key[50]), .ZN(n32034) );
  AND2_X1 U7780 ( .A1(n25966), .A2(n9115), .Z(n32035) );
  AND2_X1 U7782 ( .A1(n24201), .A2(n6911), .Z(n32036) );
  AND2_X1 U7788 ( .A1(n1567), .A2(n8210), .Z(n32038) );
  OR2_X2 U7789 ( .A1(n21532), .A2(n30389), .Z(n32039) );
  OR2_X2 U7790 ( .A1(n18221), .A2(n14487), .Z(n32040) );
  INV_X2 U7794 ( .I(n9951), .ZN(n985) );
  NOR2_X1 U7797 ( .A1(n22332), .A2(n4330), .ZN(n32042) );
  AND2_X1 U7799 ( .A1(n30987), .A2(n32201), .Z(n32043) );
  XNOR2_X1 U7801 ( .A1(n19712), .A2(n25878), .ZN(n32044) );
  AND2_X2 U7802 ( .A1(n522), .A2(n7513), .Z(n32045) );
  XNOR2_X1 U7804 ( .A1(n19741), .A2(n24707), .ZN(n32046) );
  XNOR2_X1 U7807 ( .A1(n2073), .A2(n1393), .ZN(n32047) );
  OR2_X1 U7809 ( .A1(n22785), .A2(n3909), .Z(n32048) );
  CLKBUF_X4 U7814 ( .I(n564), .Z(n4215) );
  INV_X2 U7817 ( .I(n21812), .ZN(n1132) );
  AND2_X1 U7819 ( .A1(n24248), .A2(n28553), .Z(n32049) );
  INV_X1 U7822 ( .I(n7292), .ZN(n1356) );
  INV_X1 U7823 ( .I(n28945), .ZN(n33182) );
  OR2_X2 U7824 ( .A1(n30578), .A2(n33387), .Z(n32050) );
  INV_X1 U7826 ( .I(n17316), .ZN(n33688) );
  XOR2_X1 U7827 ( .A1(Plaintext[6]), .A2(Key[6]), .Z(n32051) );
  AND2_X2 U7830 ( .A1(n30572), .A2(n27585), .Z(n32052) );
  XNOR2_X1 U7834 ( .A1(n19744), .A2(n19743), .ZN(n32053) );
  OR2_X1 U7836 ( .A1(n8212), .A2(n2207), .Z(n32054) );
  CLKBUF_X4 U7838 ( .I(n18649), .Z(n16474) );
  XOR2_X1 U7840 ( .A1(n17284), .A2(n27268), .Z(n32055) );
  AND2_X1 U7843 ( .A1(n11444), .A2(n4835), .Z(n32056) );
  XOR2_X1 U7850 ( .A1(n11604), .A2(n1653), .Z(n32058) );
  AND2_X2 U7852 ( .A1(n2001), .A2(n2000), .Z(n32059) );
  CLKBUF_X2 U7853 ( .I(n9320), .Z(n26587) );
  INV_X1 U7855 ( .I(n19319), .ZN(n33432) );
  OR2_X1 U7857 ( .A1(n9025), .A2(n8870), .Z(n32061) );
  AND2_X2 U7858 ( .A1(n4775), .A2(n3421), .Z(n32062) );
  OR2_X2 U7860 ( .A1(n31656), .A2(n17295), .Z(n32063) );
  OR2_X1 U7863 ( .A1(n12548), .A2(n19156), .Z(n32064) );
  INV_X1 U7864 ( .I(n34010), .ZN(n29440) );
  NOR2_X1 U7866 ( .A1(n10714), .A2(n9319), .ZN(n34010) );
  XNOR2_X1 U7870 ( .A1(n9141), .A2(n20792), .ZN(n32065) );
  INV_X1 U7871 ( .I(n17144), .ZN(n21218) );
  XNOR2_X1 U7872 ( .A1(n20807), .A2(n20697), .ZN(n32067) );
  INV_X1 U7873 ( .I(n11630), .ZN(n17243) );
  NOR2_X1 U7874 ( .A1(n20208), .A2(n20207), .ZN(n32399) );
  INV_X1 U7875 ( .I(n16489), .ZN(n938) );
  INV_X1 U7881 ( .I(n33856), .ZN(n34154) );
  INV_X1 U7883 ( .I(n8813), .ZN(n14721) );
  AND2_X2 U7892 ( .A1(n12227), .A2(n20361), .Z(n32068) );
  XNOR2_X1 U7893 ( .A1(n20740), .A2(n20739), .ZN(n32069) );
  INV_X1 U7894 ( .I(n21952), .ZN(n32695) );
  XNOR2_X1 U7897 ( .A1(n20862), .A2(n13357), .ZN(n32070) );
  INV_X1 U7905 ( .I(n28254), .ZN(n21257) );
  CLKBUF_X2 U7909 ( .I(n28254), .Z(n33684) );
  INV_X1 U7912 ( .I(n21392), .ZN(n21368) );
  XNOR2_X1 U7918 ( .A1(n26785), .A2(n22220), .ZN(n32072) );
  XNOR2_X1 U7919 ( .A1(n13857), .A2(n13856), .ZN(n32074) );
  AND2_X1 U7924 ( .A1(n32815), .A2(n16117), .Z(n32075) );
  INV_X2 U7925 ( .I(n13382), .ZN(n1127) );
  OR2_X2 U7926 ( .A1(n6765), .A2(n17888), .Z(n32076) );
  XNOR2_X1 U7929 ( .A1(n623), .A2(n22022), .ZN(n32077) );
  XOR2_X1 U7930 ( .A1(n33202), .A2(n3353), .Z(n32078) );
  INV_X1 U7931 ( .I(n22148), .ZN(n22221) );
  XNOR2_X1 U7932 ( .A1(n6811), .A2(n6809), .ZN(n32081) );
  XNOR2_X1 U7933 ( .A1(n4589), .A2(n4590), .ZN(n32082) );
  XNOR2_X1 U7937 ( .A1(n22312), .A2(n21050), .ZN(n32083) );
  AND2_X2 U7938 ( .A1(n15314), .A2(n15316), .Z(n32084) );
  INV_X1 U7941 ( .I(n10402), .ZN(n28924) );
  INV_X1 U7946 ( .I(n26292), .ZN(n33237) );
  INV_X1 U7947 ( .I(n25963), .ZN(n32830) );
  XNOR2_X1 U7954 ( .A1(n7623), .A2(n7622), .ZN(n32085) );
  INV_X2 U7955 ( .I(n22425), .ZN(n1728) );
  AND2_X1 U7959 ( .A1(n28865), .A2(n22467), .Z(n32087) );
  INV_X1 U7961 ( .I(n622), .ZN(n11892) );
  AND2_X2 U7962 ( .A1(n15806), .A2(n4580), .Z(n32089) );
  NAND3_X1 U7963 ( .A1(n22398), .A2(n708), .A3(n17853), .ZN(n32090) );
  AND2_X1 U7964 ( .A1(n30234), .A2(n30868), .Z(n32091) );
  NAND2_X1 U7967 ( .A1(n9798), .A2(n28608), .ZN(n32093) );
  INV_X1 U7968 ( .I(n23886), .ZN(n23889) );
  INV_X2 U7969 ( .I(n14540), .ZN(n1271) );
  CLKBUF_X2 U7971 ( .I(n13704), .Z(n13525) );
  AND3_X2 U7973 ( .A1(n30651), .A2(n10226), .A3(n7935), .Z(n32094) );
  CLKBUF_X1 U7977 ( .I(n24870), .Z(n25152) );
  AND2_X1 U7978 ( .A1(n24143), .A2(n24142), .Z(n32095) );
  INV_X1 U7979 ( .I(n33235), .ZN(n736) );
  INV_X1 U7980 ( .I(n24242), .ZN(n33540) );
  XNOR2_X1 U7981 ( .A1(n6898), .A2(n33359), .ZN(n32096) );
  INV_X1 U7984 ( .I(n13232), .ZN(n14112) );
  INV_X1 U7985 ( .I(n24719), .ZN(n33155) );
  CLKBUF_X2 U7991 ( .I(n24719), .Z(n25866) );
  INV_X1 U7992 ( .I(n31783), .ZN(n25303) );
  XOR2_X1 U8000 ( .A1(n1994), .A2(n19627), .Z(n12413) );
  NAND2_X2 U8003 ( .A1(n5223), .A2(n33719), .ZN(n1994) );
  NAND2_X1 U8007 ( .A1(n7310), .A2(n3909), .ZN(n5832) );
  NAND2_X2 U8010 ( .A1(n28083), .A2(n4221), .ZN(n3909) );
  INV_X1 U8012 ( .I(n27728), .ZN(n19464) );
  XNOR2_X1 U8013 ( .A1(n3964), .A2(n19400), .ZN(n27728) );
  NOR2_X2 U8015 ( .A1(n14342), .A2(n32097), .ZN(n14624) );
  OAI21_X2 U8020 ( .A1(n32071), .A2(n30223), .B(n21653), .ZN(n30846) );
  XOR2_X1 U8021 ( .A1(n8583), .A2(n12539), .Z(n13455) );
  NAND2_X2 U8023 ( .A1(n21410), .A2(n10113), .ZN(n33886) );
  NAND2_X2 U8024 ( .A1(n33888), .A2(n31835), .ZN(n21410) );
  NAND3_X2 U8026 ( .A1(n32706), .A2(n28206), .A3(n22651), .ZN(n26568) );
  XOR2_X1 U8028 ( .A1(n22136), .A2(n32098), .Z(n32631) );
  XOR2_X1 U8031 ( .A1(n22134), .A2(n32099), .Z(n32098) );
  AOI21_X1 U8034 ( .A1(n31904), .A2(n32101), .B(n4193), .ZN(n31216) );
  OR2_X1 U8035 ( .A1(n7586), .A2(n5713), .Z(n32101) );
  NAND2_X2 U8037 ( .A1(n10922), .A2(n31677), .ZN(n1313) );
  NOR2_X1 U8042 ( .A1(n601), .A2(n1736), .ZN(n33705) );
  XOR2_X1 U8044 ( .A1(n3099), .A2(n32103), .Z(n7119) );
  XOR2_X1 U8045 ( .A1(n33892), .A2(n9464), .Z(n32103) );
  XOR2_X1 U8046 ( .A1(n9627), .A2(n20869), .Z(n28981) );
  NAND2_X2 U8050 ( .A1(n28733), .A2(n30197), .ZN(n9627) );
  OR2_X1 U8051 ( .A1(n20310), .A2(n7102), .Z(n16004) );
  NAND2_X2 U8052 ( .A1(n4079), .A2(n33724), .ZN(n23684) );
  NAND2_X2 U8053 ( .A1(n24292), .A2(n15520), .ZN(n24011) );
  NAND2_X2 U8054 ( .A1(n26529), .A2(n23685), .ZN(n9219) );
  AOI21_X2 U8058 ( .A1(n32104), .A2(n27094), .B(n22335), .ZN(n22999) );
  NOR2_X2 U8060 ( .A1(n20378), .A2(n27887), .ZN(n20323) );
  INV_X4 U8062 ( .I(n33817), .ZN(n22876) );
  NAND2_X2 U8068 ( .A1(n32105), .A2(n32090), .ZN(n33817) );
  INV_X2 U8071 ( .I(n8601), .ZN(n32105) );
  XOR2_X1 U8072 ( .A1(n27289), .A2(n7129), .Z(n9920) );
  INV_X2 U8080 ( .I(n32370), .ZN(n27390) );
  XOR2_X1 U8081 ( .A1(n5196), .A2(n31929), .Z(n32370) );
  NOR2_X2 U8082 ( .A1(n13903), .A2(n32107), .ZN(n32462) );
  NOR3_X2 U8087 ( .A1(n23749), .A2(n16781), .A3(n6661), .ZN(n32107) );
  AOI22_X2 U8094 ( .A1(n11022), .A2(n4993), .B1(n25896), .B2(n5387), .ZN(
        n32132) );
  NOR2_X2 U8099 ( .A1(n4993), .A2(n25870), .ZN(n25896) );
  NAND2_X2 U8100 ( .A1(n33044), .A2(n31946), .ZN(n32859) );
  BUF_X2 U8102 ( .I(n32787), .Z(n32108) );
  NAND2_X2 U8105 ( .A1(n33321), .A2(n4131), .ZN(n32255) );
  INV_X2 U8108 ( .I(n32109), .ZN(n2229) );
  NOR2_X2 U8109 ( .A1(n22557), .A2(n5379), .ZN(n32496) );
  AOI22_X2 U8114 ( .A1(n32110), .A2(n834), .B1(n1620), .B2(n12266), .ZN(n25790) );
  NAND2_X2 U8116 ( .A1(n12440), .A2(n25866), .ZN(n32110) );
  XOR2_X1 U8117 ( .A1(n14953), .A2(n14952), .Z(n32124) );
  XOR2_X1 U8118 ( .A1(n23469), .A2(n2854), .Z(n9200) );
  NAND2_X2 U8119 ( .A1(n30008), .A2(n7839), .ZN(n2854) );
  NOR2_X2 U8121 ( .A1(n927), .A2(n30813), .ZN(n2370) );
  XOR2_X1 U8122 ( .A1(n21023), .A2(n21025), .Z(n6792) );
  XOR2_X1 U8124 ( .A1(n13357), .A2(n5414), .Z(n21023) );
  OAI22_X2 U8125 ( .A1(n31964), .A2(n22487), .B1(n1289), .B2(n11629), .ZN(
        n16884) );
  INV_X2 U8127 ( .I(n9617), .ZN(n11629) );
  XOR2_X1 U8129 ( .A1(n2144), .A2(n5353), .Z(n9617) );
  XOR2_X1 U8131 ( .A1(n2267), .A2(n28998), .Z(n10657) );
  NAND3_X1 U8135 ( .A1(n25793), .A2(n25792), .A3(n25791), .ZN(n34070) );
  INV_X2 U8136 ( .I(n16486), .ZN(n22865) );
  NOR3_X1 U8137 ( .A1(n15382), .A2(n14905), .A3(n15476), .ZN(n30771) );
  XOR2_X1 U8139 ( .A1(n12972), .A2(n4992), .Z(n5487) );
  NOR2_X2 U8141 ( .A1(n1983), .A2(n5605), .ZN(n4992) );
  XOR2_X1 U8144 ( .A1(n4975), .A2(n12442), .Z(n13908) );
  BUF_X2 U8147 ( .I(n29898), .Z(n32111) );
  NOR2_X1 U8148 ( .A1(n10987), .A2(n24326), .ZN(n24329) );
  NAND2_X2 U8149 ( .A1(n29811), .A2(n31090), .ZN(n24326) );
  NAND2_X2 U8150 ( .A1(n22353), .A2(n27638), .ZN(n6750) );
  OAI22_X2 U8154 ( .A1(n26410), .A2(n27390), .B1(n29142), .B2(n8919), .ZN(
        n22353) );
  XOR2_X1 U8155 ( .A1(n30301), .A2(n5762), .Z(n24575) );
  NAND2_X1 U8156 ( .A1(n10231), .A2(n20236), .ZN(n13432) );
  XOR2_X1 U8157 ( .A1(n24643), .A2(n24753), .Z(n24419) );
  NAND2_X2 U8159 ( .A1(n24078), .A2(n24077), .ZN(n24643) );
  NAND2_X2 U8162 ( .A1(n33133), .A2(n31878), .ZN(n29898) );
  NOR3_X2 U8163 ( .A1(n32115), .A2(n32112), .A3(n17849), .ZN(n31571) );
  NOR3_X2 U8164 ( .A1(n4183), .A2(n25462), .A3(n29116), .ZN(n32112) );
  AOI21_X2 U8165 ( .A1(n14722), .A2(n14087), .B(n33352), .ZN(n5906) );
  NAND2_X2 U8166 ( .A1(n5820), .A2(n1106), .ZN(n23028) );
  AOI22_X2 U8167 ( .A1(n1232), .A2(n5079), .B1(n5080), .B2(n29985), .ZN(n5284)
         );
  NAND2_X2 U8170 ( .A1(n23981), .A2(n421), .ZN(n5080) );
  XOR2_X1 U8174 ( .A1(n6461), .A2(n14613), .Z(n32914) );
  XOR2_X1 U8177 ( .A1(n417), .A2(n32113), .Z(n7072) );
  XOR2_X1 U8179 ( .A1(n33840), .A2(n32114), .Z(n32113) );
  XOR2_X1 U8187 ( .A1(n22225), .A2(n34078), .Z(n16897) );
  XOR2_X1 U8190 ( .A1(n22190), .A2(n22191), .Z(n11358) );
  XOR2_X1 U8192 ( .A1(n7725), .A2(n21892), .Z(n22190) );
  AOI21_X2 U8197 ( .A1(n16001), .A2(n25753), .B(n1082), .ZN(n15709) );
  NAND2_X1 U8198 ( .A1(n25707), .A2(n25705), .ZN(n25753) );
  NAND3_X1 U8201 ( .A1(n11186), .A2(n25905), .A3(n25901), .ZN(n11185) );
  NAND2_X2 U8207 ( .A1(n21378), .A2(n15751), .ZN(n15728) );
  NAND2_X2 U8209 ( .A1(n21362), .A2(n2230), .ZN(n21378) );
  NOR2_X2 U8210 ( .A1(n33735), .A2(n32116), .ZN(n16987) );
  NOR2_X2 U8211 ( .A1(n1351), .A2(n20447), .ZN(n20405) );
  AOI21_X2 U8213 ( .A1(n32723), .A2(n28982), .B(n27373), .ZN(n20447) );
  XOR2_X1 U8214 ( .A1(n32117), .A2(n24740), .Z(n7759) );
  XOR2_X1 U8215 ( .A1(n33447), .A2(n705), .Z(n32117) );
  XOR2_X1 U8217 ( .A1(n33319), .A2(n32118), .Z(n11622) );
  XOR2_X1 U8219 ( .A1(n11782), .A2(n24803), .Z(n32118) );
  INV_X4 U8220 ( .I(n16305), .ZN(n32298) );
  AND2_X1 U8221 ( .A1(n9390), .A2(n13969), .Z(n5583) );
  XOR2_X1 U8222 ( .A1(n21891), .A2(n7289), .Z(n9193) );
  NAND2_X2 U8224 ( .A1(n1678), .A2(n1677), .ZN(n33117) );
  OAI21_X2 U8226 ( .A1(n21465), .A2(n11729), .B(n26728), .ZN(n16888) );
  XOR2_X1 U8229 ( .A1(n2956), .A2(n16520), .Z(n210) );
  NAND3_X2 U8234 ( .A1(n27759), .A2(n33372), .A3(n27760), .ZN(n2956) );
  XOR2_X1 U8238 ( .A1(n32120), .A2(n25783), .Z(Ciphertext[165]) );
  NAND3_X2 U8239 ( .A1(n28989), .A2(n17222), .A3(n26948), .ZN(n32120) );
  NAND2_X2 U8241 ( .A1(n28073), .A2(n32121), .ZN(n19314) );
  NAND2_X2 U8244 ( .A1(n32150), .A2(n32122), .ZN(n23928) );
  NAND3_X1 U8248 ( .A1(n16186), .A2(n4892), .A3(n23920), .ZN(n32122) );
  NAND2_X2 U8256 ( .A1(n7146), .A2(n32123), .ZN(n9159) );
  AOI22_X2 U8259 ( .A1(n21320), .A2(n11187), .B1(n21324), .B2(n28017), .ZN(
        n32123) );
  XOR2_X1 U8260 ( .A1(n23358), .A2(n23253), .Z(n23516) );
  NAND3_X2 U8261 ( .A1(n22751), .A2(n22750), .A3(n22749), .ZN(n23253) );
  NAND2_X2 U8264 ( .A1(n32126), .A2(n32125), .ZN(n26102) );
  INV_X2 U8266 ( .I(n12594), .ZN(n32125) );
  XOR2_X1 U8270 ( .A1(n13858), .A2(n7880), .Z(n32469) );
  XOR2_X1 U8272 ( .A1(n24545), .A2(n24544), .Z(n7880) );
  BUF_X2 U8275 ( .I(n16559), .Z(n32127) );
  NAND2_X2 U8281 ( .A1(n57), .A2(n32128), .ZN(n24254) );
  XOR2_X1 U8283 ( .A1(n19768), .A2(n19703), .Z(n19517) );
  AOI21_X2 U8288 ( .A1(n5654), .A2(n18621), .B(n31438), .ZN(n19768) );
  NAND2_X2 U8290 ( .A1(n10980), .A2(n32129), .ZN(n21767) );
  OR2_X1 U8291 ( .A1(n21051), .A2(n33684), .Z(n32129) );
  OAI21_X2 U8294 ( .A1(n6710), .A2(n6711), .B(n6712), .ZN(n6799) );
  NOR2_X2 U8295 ( .A1(n4207), .A2(n6877), .ZN(n7078) );
  AOI21_X2 U8296 ( .A1(n7151), .A2(n14995), .B(n972), .ZN(n4207) );
  XOR2_X1 U8297 ( .A1(n348), .A2(n32130), .Z(n12805) );
  NAND2_X1 U8299 ( .A1(n29981), .A2(n11507), .ZN(n19984) );
  NOR2_X2 U8300 ( .A1(n33720), .A2(n25784), .ZN(n32874) );
  NOR3_X2 U8301 ( .A1(n25757), .A2(n3275), .A3(n11899), .ZN(n33720) );
  OR2_X1 U8302 ( .A1(n8062), .A2(n4897), .Z(n4873) );
  INV_X2 U8304 ( .I(n25106), .ZN(n7334) );
  XOR2_X1 U8305 ( .A1(n5601), .A2(n33338), .Z(n8964) );
  XOR2_X1 U8309 ( .A1(n32131), .A2(n32895), .Z(n15731) );
  XOR2_X1 U8310 ( .A1(n32243), .A2(n33265), .Z(n32131) );
  OAI21_X2 U8311 ( .A1(n19051), .A2(n19000), .B(n27877), .ZN(n19423) );
  AOI22_X2 U8312 ( .A1(n18999), .A2(n19217), .B1(n19216), .B2(n31366), .ZN(
        n27877) );
  XOR2_X1 U8313 ( .A1(n23312), .A2(n23341), .Z(n11039) );
  NAND2_X1 U8314 ( .A1(n33235), .A2(n24866), .ZN(n16850) );
  XOR2_X1 U8315 ( .A1(n33161), .A2(n14065), .Z(n24866) );
  NOR2_X1 U8318 ( .A1(n25002), .A2(n3232), .ZN(n14609) );
  OAI21_X2 U8319 ( .A1(n15061), .A2(n15062), .B(n15059), .ZN(n25002) );
  XOR2_X1 U8320 ( .A1(n10631), .A2(n3935), .Z(n32417) );
  NOR2_X2 U8322 ( .A1(n14502), .A2(n4959), .ZN(n10631) );
  INV_X4 U8324 ( .I(n14001), .ZN(n24925) );
  NAND2_X2 U8325 ( .A1(n8776), .A2(n8777), .ZN(n14001) );
  AOI22_X2 U8330 ( .A1(n23912), .A2(n7005), .B1(n23910), .B2(n23588), .ZN(
        n33808) );
  INV_X2 U8333 ( .I(n16226), .ZN(n21078) );
  XOR2_X1 U8335 ( .A1(n26954), .A2(n13403), .Z(n16226) );
  NAND2_X2 U8336 ( .A1(n11020), .A2(n32132), .ZN(n13960) );
  XOR2_X1 U8346 ( .A1(n24513), .A2(n30323), .Z(n24788) );
  NAND3_X2 U8349 ( .A1(n4393), .A2(n17493), .A3(n17492), .ZN(n24513) );
  NOR2_X2 U8351 ( .A1(n12662), .A2(n34127), .ZN(n33306) );
  NAND2_X2 U8352 ( .A1(n7034), .A2(n32133), .ZN(n8238) );
  AOI22_X2 U8354 ( .A1(n7885), .A2(n33589), .B1(n23650), .B2(n28671), .ZN(
        n32133) );
  NAND2_X2 U8356 ( .A1(n22399), .A2(n17930), .ZN(n23046) );
  NAND2_X2 U8357 ( .A1(n21980), .A2(n21981), .ZN(n22399) );
  XOR2_X1 U8358 ( .A1(n32134), .A2(n19492), .Z(n706) );
  XOR2_X1 U8359 ( .A1(n27895), .A2(n19577), .Z(n32134) );
  OAI21_X2 U8361 ( .A1(n32135), .A2(n17762), .B(n8307), .ZN(n32731) );
  XOR2_X1 U8363 ( .A1(n32136), .A2(n1431), .Z(Ciphertext[163]) );
  NOR3_X1 U8366 ( .A1(n28854), .A2(n14615), .A3(n12395), .ZN(n32136) );
  XOR2_X1 U8369 ( .A1(n6466), .A2(n32137), .Z(n7) );
  XOR2_X1 U8371 ( .A1(n21893), .A2(n32072), .Z(n32137) );
  NOR2_X2 U8372 ( .A1(n30473), .A2(n24025), .ZN(n24936) );
  OAI22_X2 U8374 ( .A1(n13326), .A2(n14268), .B1(n14042), .B2(n1221), .ZN(
        n30473) );
  NAND2_X2 U8375 ( .A1(n32139), .A2(n32138), .ZN(n28539) );
  NOR2_X1 U8378 ( .A1(n31992), .A2(n13160), .ZN(n32139) );
  XOR2_X1 U8381 ( .A1(n32140), .A2(n24407), .Z(n17074) );
  XOR2_X1 U8387 ( .A1(n12422), .A2(n12512), .Z(n32140) );
  BUF_X2 U8388 ( .I(n1169), .Z(n32141) );
  NAND2_X2 U8389 ( .A1(n32142), .A2(n9085), .ZN(n5973) );
  NAND3_X2 U8394 ( .A1(n32048), .A2(n22953), .A3(n7544), .ZN(n32142) );
  XOR2_X1 U8395 ( .A1(n20789), .A2(n20787), .Z(n31070) );
  XOR2_X1 U8403 ( .A1(n10235), .A2(n1507), .Z(n28747) );
  XOR2_X1 U8405 ( .A1(n24842), .A2(n12720), .Z(n1507) );
  NAND2_X1 U8406 ( .A1(n18352), .A2(n9264), .ZN(n32769) );
  AOI22_X2 U8409 ( .A1(n16866), .A2(n22477), .B1(n27207), .B2(n18098), .ZN(
        n32482) );
  NAND3_X2 U8412 ( .A1(n3708), .A2(n8799), .A3(n32145), .ZN(n11754) );
  AOI22_X2 U8415 ( .A1(n4319), .A2(n17694), .B1(n29080), .B2(n30980), .ZN(
        n32145) );
  INV_X1 U8420 ( .I(n31185), .ZN(n20777) );
  NAND2_X2 U8423 ( .A1(n32288), .A2(n32146), .ZN(n1560) );
  NAND3_X2 U8425 ( .A1(n12429), .A2(n12430), .A3(n32936), .ZN(n32146) );
  XOR2_X1 U8426 ( .A1(n15517), .A2(n32870), .Z(n24746) );
  NAND2_X2 U8435 ( .A1(n15988), .A2(n13658), .ZN(n15517) );
  NAND2_X1 U8437 ( .A1(n2643), .A2(n14681), .ZN(n21469) );
  NAND2_X2 U8438 ( .A1(n8740), .A2(n21153), .ZN(n2643) );
  NOR2_X1 U8439 ( .A1(n25587), .A2(n25586), .ZN(n33500) );
  OAI21_X1 U8441 ( .A1(n13066), .A2(n9003), .B(n9954), .ZN(n30838) );
  XOR2_X1 U8443 ( .A1(n20861), .A2(n17423), .Z(n10169) );
  NAND2_X2 U8445 ( .A1(n14567), .A2(n14565), .ZN(n20861) );
  NOR2_X1 U8448 ( .A1(n32148), .A2(n861), .ZN(n29843) );
  NOR2_X2 U8451 ( .A1(n32149), .A2(n13212), .ZN(n6569) );
  NAND2_X1 U8454 ( .A1(n32151), .A2(n8760), .ZN(n32150) );
  NOR2_X1 U8461 ( .A1(n23920), .A2(n13361), .ZN(n32151) );
  XOR2_X1 U8462 ( .A1(n32733), .A2(n19679), .Z(n8637) );
  XOR2_X1 U8466 ( .A1(n30547), .A2(n32152), .Z(n23916) );
  XOR2_X1 U8473 ( .A1(n23334), .A2(n14527), .Z(n32152) );
  XOR2_X1 U8478 ( .A1(n20713), .A2(n32153), .Z(n21071) );
  XOR2_X1 U8479 ( .A1(n21020), .A2(n12618), .Z(n32153) );
  NOR2_X2 U8481 ( .A1(n8247), .A2(n8246), .ZN(n8245) );
  AOI22_X2 U8483 ( .A1(n6559), .A2(n20300), .B1(n20358), .B2(n16011), .ZN(
        n17177) );
  NOR2_X2 U8484 ( .A1(n20238), .A2(n11453), .ZN(n16011) );
  NOR2_X1 U8485 ( .A1(n33512), .A2(n16304), .ZN(n16410) );
  XOR2_X1 U8488 ( .A1(n32155), .A2(n32156), .Z(n33534) );
  XOR2_X1 U8490 ( .A1(n26462), .A2(n21944), .Z(n32156) );
  XOR2_X1 U8493 ( .A1(n32157), .A2(n25541), .Z(Ciphertext[120]) );
  NAND4_X2 U8499 ( .A1(n8805), .A2(n30134), .A3(n8804), .A4(n25555), .ZN(
        n32157) );
  NOR2_X1 U8500 ( .A1(n12302), .A2(n27925), .ZN(n32566) );
  AOI22_X2 U8501 ( .A1(n12482), .A2(n17005), .B1(n9294), .B2(n27990), .ZN(
        n16380) );
  OAI22_X2 U8502 ( .A1(n9294), .A2(n28591), .B1(n25199), .B2(n32873), .ZN(
        n12482) );
  INV_X2 U8507 ( .I(n23405), .ZN(n33476) );
  NAND2_X2 U8509 ( .A1(n30982), .A2(n16879), .ZN(n23405) );
  XOR2_X1 U8511 ( .A1(n19390), .A2(n19568), .Z(n2951) );
  XOR2_X1 U8512 ( .A1(n19629), .A2(n19389), .Z(n19568) );
  NAND3_X2 U8513 ( .A1(n20444), .A2(n30496), .A3(n20633), .ZN(n4469) );
  NAND2_X2 U8514 ( .A1(n30594), .A2(n15162), .ZN(n20444) );
  NOR2_X1 U8515 ( .A1(n31448), .A2(n19936), .ZN(n14905) );
  INV_X2 U8518 ( .I(n32158), .ZN(n11933) );
  XNOR2_X1 U8520 ( .A1(n284), .A2(n10051), .ZN(n32158) );
  NAND2_X2 U8521 ( .A1(n12214), .A2(n32159), .ZN(n16807) );
  NAND2_X2 U8522 ( .A1(n18324), .A2(n18567), .ZN(n32159) );
  INV_X2 U8534 ( .I(n29261), .ZN(n22477) );
  XOR2_X1 U8535 ( .A1(n32160), .A2(n24689), .Z(n24407) );
  XOR2_X1 U8538 ( .A1(n24785), .A2(n30327), .Z(n32160) );
  NAND2_X2 U8541 ( .A1(n17249), .A2(n32161), .ZN(n1266) );
  NAND3_X2 U8544 ( .A1(n17247), .A2(n17248), .A3(n9620), .ZN(n32161) );
  XOR2_X1 U8547 ( .A1(n15560), .A2(n22061), .Z(n14181) );
  NAND2_X2 U8548 ( .A1(n26102), .A2(n2777), .ZN(n15560) );
  XOR2_X1 U8549 ( .A1(n27175), .A2(n25783), .Z(n102) );
  NOR3_X2 U8551 ( .A1(n17740), .A2(n12445), .A3(n12444), .ZN(n27175) );
  NOR2_X2 U8552 ( .A1(n13319), .A2(n13255), .ZN(n21381) );
  AND2_X1 U8560 ( .A1(n17948), .A2(n15212), .Z(n29280) );
  XOR2_X1 U8561 ( .A1(n32162), .A2(n32467), .Z(n30492) );
  NAND2_X2 U8564 ( .A1(n3424), .A2(n30079), .ZN(n32467) );
  INV_X2 U8565 ( .I(n11665), .ZN(n32162) );
  XOR2_X1 U8567 ( .A1(n8070), .A2(n8069), .Z(n23587) );
  NOR2_X2 U8568 ( .A1(n23860), .A2(n23556), .ZN(n26955) );
  NAND2_X2 U8569 ( .A1(n28273), .A2(n17661), .ZN(n23556) );
  NAND2_X2 U8572 ( .A1(n18991), .A2(n18992), .ZN(n19400) );
  NOR2_X2 U8573 ( .A1(n13678), .A2(n33583), .ZN(n26628) );
  NAND2_X2 U8575 ( .A1(n206), .A2(n17375), .ZN(n30033) );
  NAND2_X2 U8577 ( .A1(n10939), .A2(n8268), .ZN(n20200) );
  NAND2_X2 U8580 ( .A1(n2495), .A2(n33003), .ZN(n10939) );
  NAND2_X2 U8581 ( .A1(n32163), .A2(n32289), .ZN(n31171) );
  NAND2_X1 U8586 ( .A1(n12208), .A2(n16305), .ZN(n32163) );
  INV_X2 U8592 ( .I(n26898), .ZN(n23034) );
  NAND3_X2 U8594 ( .A1(n33901), .A2(n1516), .A3(n30989), .ZN(n26898) );
  NAND2_X2 U8596 ( .A1(n22474), .A2(n29261), .ZN(n13185) );
  OAI21_X2 U8599 ( .A1(n8230), .A2(n32164), .B(n34104), .ZN(n26261) );
  NAND2_X1 U8600 ( .A1(n6483), .A2(n21580), .ZN(n32164) );
  NAND3_X1 U8601 ( .A1(n4086), .A2(n33097), .A3(n23628), .ZN(n33135) );
  BUF_X4 U8604 ( .I(n28374), .Z(n32323) );
  XOR2_X1 U8605 ( .A1(n4672), .A2(n32165), .Z(n5361) );
  XOR2_X1 U8611 ( .A1(n4671), .A2(n4771), .Z(n32165) );
  XOR2_X1 U8628 ( .A1(Plaintext[20]), .A2(Key[20]), .Z(n18655) );
  AOI22_X2 U8630 ( .A1(n4774), .A2(n11041), .B1(n12982), .B2(n24309), .ZN(
        n24199) );
  OAI22_X2 U8636 ( .A1(n4099), .A2(n6723), .B1(n31982), .B2(n18204), .ZN(
        n24309) );
  NOR3_X2 U8637 ( .A1(n33455), .A2(n9335), .A3(n5743), .ZN(n32636) );
  AOI21_X2 U8640 ( .A1(n32166), .A2(n2993), .B(n26545), .ZN(n2158) );
  XOR2_X1 U8642 ( .A1(n17519), .A2(n22275), .Z(n15618) );
  XOR2_X1 U8645 ( .A1(n14125), .A2(n7808), .Z(n17519) );
  NAND2_X1 U8650 ( .A1(n29614), .A2(n14418), .ZN(n32430) );
  NAND2_X1 U8651 ( .A1(n18133), .A2(n32309), .ZN(n23715) );
  XOR2_X1 U8652 ( .A1(n31237), .A2(n23537), .Z(n32309) );
  XOR2_X1 U8655 ( .A1(n20905), .A2(n27174), .Z(n20989) );
  NAND2_X2 U8658 ( .A1(n5951), .A2(n5949), .ZN(n20905) );
  XOR2_X1 U8666 ( .A1(n32167), .A2(n16775), .Z(n28179) );
  XOR2_X1 U8667 ( .A1(n27729), .A2(n20824), .Z(n32167) );
  XOR2_X1 U8668 ( .A1(n9207), .A2(n27693), .Z(n26317) );
  NOR2_X2 U8670 ( .A1(n29547), .A2(n32168), .ZN(n29523) );
  XOR2_X1 U8672 ( .A1(n26701), .A2(n23186), .Z(n23246) );
  NAND3_X2 U8675 ( .A1(n33777), .A2(n13365), .A3(n14516), .ZN(n26701) );
  INV_X2 U8677 ( .I(n21628), .ZN(n21772) );
  AOI22_X2 U8679 ( .A1(n31524), .A2(n23669), .B1(n23953), .B2(n33788), .ZN(
        n9995) );
  NAND2_X2 U8680 ( .A1(n12986), .A2(n32169), .ZN(n26585) );
  OAI21_X2 U8682 ( .A1(n19801), .A2(n19800), .B(n19867), .ZN(n32169) );
  XOR2_X1 U8688 ( .A1(n11218), .A2(n19529), .Z(n4578) );
  XOR2_X1 U8696 ( .A1(n30943), .A2(n19708), .Z(n19529) );
  XOR2_X1 U8700 ( .A1(n21014), .A2(n20718), .Z(n32379) );
  XOR2_X1 U8713 ( .A1(n2789), .A2(n2198), .Z(n20718) );
  OAI21_X1 U8714 ( .A1(n8334), .A2(n22962), .B(n22815), .ZN(n33049) );
  BUF_X2 U8716 ( .I(n15917), .Z(n32170) );
  XOR2_X1 U8719 ( .A1(n32171), .A2(n13863), .Z(n15205) );
  XOR2_X1 U8723 ( .A1(n32367), .A2(n27240), .Z(n32171) );
  BUF_X2 U8725 ( .I(n32081), .Z(n32172) );
  OAI21_X2 U8733 ( .A1(n30617), .A2(n19761), .B(n32173), .ZN(n20312) );
  AOI22_X2 U8734 ( .A1(n19759), .A2(n20045), .B1(n31715), .B2(n31823), .ZN(
        n32173) );
  NAND3_X2 U8736 ( .A1(n29668), .A2(n20414), .A3(n19908), .ZN(n29667) );
  XOR2_X1 U8741 ( .A1(n19626), .A2(n19624), .Z(n17541) );
  OAI22_X2 U8746 ( .A1(n12271), .A2(n12268), .B1(n7968), .B2(n18752), .ZN(
        n19626) );
  NAND2_X2 U8749 ( .A1(n33767), .A2(n32174), .ZN(n5211) );
  AOI22_X2 U8750 ( .A1(n32234), .A2(n32233), .B1(n5821), .B2(n16976), .ZN(
        n32174) );
  NAND2_X2 U8752 ( .A1(n31030), .A2(n1333), .ZN(n21411) );
  XOR2_X1 U8753 ( .A1(n14000), .A2(n5539), .Z(n24569) );
  NAND2_X2 U8754 ( .A1(n31039), .A2(n32836), .ZN(n5539) );
  NAND2_X2 U8756 ( .A1(n29502), .A2(n32175), .ZN(n11608) );
  NAND3_X1 U8757 ( .A1(n32917), .A2(n6003), .A3(n23970), .ZN(n32175) );
  NOR2_X2 U8758 ( .A1(n31979), .A2(n25843), .ZN(n25855) );
  OAI22_X2 U8763 ( .A1(n33196), .A2(n25887), .B1(n7350), .B2(n25866), .ZN(
        n25843) );
  OAI22_X2 U8770 ( .A1(n6553), .A2(n896), .B1(n23045), .B2(n23042), .ZN(n13341) );
  XOR2_X1 U8778 ( .A1(n18365), .A2(Key[49]), .Z(n32787) );
  OR2_X1 U8782 ( .A1(n8422), .A2(n9549), .Z(n10966) );
  OAI21_X2 U8791 ( .A1(n31925), .A2(n17039), .B(n15444), .ZN(n15443) );
  NOR2_X1 U8795 ( .A1(n10599), .A2(n10787), .ZN(n17039) );
  XOR2_X1 U8798 ( .A1(n6913), .A2(n19706), .Z(n32213) );
  XOR2_X1 U8803 ( .A1(n2920), .A2(n1944), .Z(n19706) );
  XOR2_X1 U8804 ( .A1(n7674), .A2(n7628), .Z(n5321) );
  XOR2_X1 U8807 ( .A1(n21040), .A2(n33814), .Z(n7674) );
  AOI21_X2 U8809 ( .A1(n11688), .A2(n1377), .B(n19309), .ZN(n19311) );
  XOR2_X1 U8811 ( .A1(n12738), .A2(n27673), .Z(n33354) );
  XOR2_X1 U8816 ( .A1(n20755), .A2(n21016), .Z(n20722) );
  NOR2_X2 U8819 ( .A1(n1929), .A2(n1930), .ZN(n21016) );
  NAND2_X2 U8824 ( .A1(n1472), .A2(n30935), .ZN(n32177) );
  XOR2_X1 U8825 ( .A1(n6373), .A2(n24991), .Z(n7211) );
  NAND2_X2 U8829 ( .A1(n30202), .A2(n33791), .ZN(n6373) );
  NOR2_X2 U8835 ( .A1(n14178), .A2(n19153), .ZN(n17528) );
  XOR2_X1 U8837 ( .A1(n1607), .A2(n28239), .Z(n17485) );
  XOR2_X1 U8838 ( .A1(n19517), .A2(n19518), .Z(n1615) );
  XOR2_X1 U8855 ( .A1(n5775), .A2(n14662), .Z(n8556) );
  XOR2_X1 U8858 ( .A1(n20803), .A2(n32894), .Z(n14662) );
  BUF_X2 U8871 ( .I(n26158), .Z(n32178) );
  XOR2_X1 U8879 ( .A1(n32179), .A2(n380), .Z(n33903) );
  XOR2_X1 U8882 ( .A1(n10649), .A2(n12627), .Z(n32179) );
  XOR2_X1 U8886 ( .A1(n20710), .A2(n14522), .Z(n26769) );
  XOR2_X1 U8887 ( .A1(n32180), .A2(n1196), .Z(Ciphertext[24]) );
  NOR2_X1 U8888 ( .A1(n32244), .A2(n24989), .ZN(n32180) );
  XOR2_X1 U8895 ( .A1(n15035), .A2(n15036), .Z(n15734) );
  INV_X2 U8896 ( .I(n32181), .ZN(n499) );
  XNOR2_X1 U8897 ( .A1(n31411), .A2(n10219), .ZN(n32181) );
  NAND2_X1 U8908 ( .A1(n4525), .A2(n24995), .ZN(n315) );
  NOR2_X1 U8916 ( .A1(n29361), .A2(n21373), .ZN(n8856) );
  XOR2_X1 U8917 ( .A1(n12720), .A2(n17912), .Z(n24749) );
  NAND2_X2 U8922 ( .A1(n16410), .A2(n16409), .ZN(n17912) );
  NOR2_X2 U8923 ( .A1(n32183), .A2(n32182), .ZN(n8091) );
  INV_X2 U8925 ( .I(n100), .ZN(n32183) );
  XOR2_X1 U8926 ( .A1(n22063), .A2(n16696), .Z(n22064) );
  NAND2_X2 U8929 ( .A1(n32204), .A2(n9961), .ZN(n22063) );
  XOR2_X1 U8932 ( .A1(n3030), .A2(n27767), .Z(n27601) );
  AND2_X1 U8933 ( .A1(n23082), .A2(n22962), .Z(n33294) );
  XOR2_X1 U8936 ( .A1(n5146), .A2(n139), .Z(n2345) );
  OAI22_X1 U8948 ( .A1(n22697), .A2(n33675), .B1(n22816), .B2(n27419), .ZN(
        n16463) );
  XOR2_X1 U8955 ( .A1(n23299), .A2(n12475), .Z(n12474) );
  XOR2_X1 U8957 ( .A1(n27174), .A2(n15877), .Z(n20778) );
  NAND2_X2 U8967 ( .A1(n32385), .A2(n20568), .ZN(n27174) );
  NAND2_X2 U8971 ( .A1(n14184), .A2(n14724), .ZN(n24837) );
  AOI22_X2 U8974 ( .A1(n31228), .A2(n33891), .B1(n3039), .B2(n3038), .ZN(
        n14184) );
  AOI21_X2 U8975 ( .A1(n32323), .A2(n33680), .B(n30230), .ZN(n26976) );
  NAND2_X1 U8977 ( .A1(n32976), .A2(n3220), .ZN(n1504) );
  OAI21_X2 U8981 ( .A1(n32185), .A2(n16367), .B(n16366), .ZN(n31282) );
  AOI22_X2 U8985 ( .A1(n239), .A2(n22557), .B1(n22343), .B2(n7090), .ZN(n32185) );
  AND2_X1 U8986 ( .A1(n33224), .A2(n2957), .Z(n12343) );
  AND2_X1 U8988 ( .A1(n18184), .A2(n32040), .Z(n17734) );
  NAND3_X2 U9005 ( .A1(n17415), .A2(n21345), .A3(n15422), .ZN(n18184) );
  AOI21_X2 U9007 ( .A1(n820), .A2(n33714), .B(n16568), .ZN(n4442) );
  INV_X1 U9010 ( .I(n13913), .ZN(n32952) );
  XNOR2_X1 U9022 ( .A1(n31477), .A2(n20754), .ZN(n31185) );
  XOR2_X1 U9023 ( .A1(n33369), .A2(n26140), .Z(n27736) );
  NAND2_X1 U9024 ( .A1(n23111), .A2(n3103), .ZN(n30476) );
  NAND2_X2 U9025 ( .A1(n29598), .A2(n32518), .ZN(n3103) );
  XOR2_X1 U9026 ( .A1(n13178), .A2(n8160), .Z(n13177) );
  NAND3_X2 U9028 ( .A1(n31998), .A2(n28880), .A3(n19874), .ZN(n27879) );
  OAI21_X2 U9031 ( .A1(n13950), .A2(n11503), .B(n24286), .ZN(n33184) );
  INV_X2 U9033 ( .I(n9624), .ZN(n11503) );
  NAND3_X2 U9034 ( .A1(n32), .A2(n25954), .A3(n6467), .ZN(n9624) );
  XOR2_X1 U9036 ( .A1(n20784), .A2(n20990), .Z(n20886) );
  NOR2_X2 U9041 ( .A1(n12479), .A2(n7033), .ZN(n20784) );
  OAI21_X2 U9044 ( .A1(n28406), .A2(n17985), .B(n32187), .ZN(n3313) );
  NAND2_X2 U9045 ( .A1(n28400), .A2(n17985), .ZN(n32187) );
  OAI21_X2 U9053 ( .A1(n9184), .A2(n32188), .B(n23043), .ZN(n23049) );
  NOR2_X2 U9056 ( .A1(n33007), .A2(n23042), .ZN(n32188) );
  XOR2_X1 U9059 ( .A1(n31769), .A2(n32189), .Z(n9626) );
  XOR2_X1 U9060 ( .A1(n28981), .A2(n10122), .Z(n32189) );
  XOR2_X1 U9062 ( .A1(n30482), .A2(n11326), .Z(n5509) );
  XOR2_X1 U9065 ( .A1(n32190), .A2(n25074), .Z(Ciphertext[44]) );
  INV_X2 U9068 ( .I(n22689), .ZN(n32194) );
  XOR2_X1 U9070 ( .A1(n9347), .A2(n32195), .Z(n29471) );
  XOR2_X1 U9072 ( .A1(n32715), .A2(n23384), .Z(n32195) );
  XOR2_X1 U9074 ( .A1(n33929), .A2(n32196), .Z(n29631) );
  XOR2_X1 U9076 ( .A1(n12659), .A2(n34112), .Z(n32196) );
  NAND2_X2 U9077 ( .A1(n25980), .A2(n397), .ZN(n10286) );
  NAND2_X2 U9078 ( .A1(n13139), .A2(n32198), .ZN(n12374) );
  AOI22_X2 U9080 ( .A1(n33870), .A2(n975), .B1(n23778), .B2(n6992), .ZN(n32198) );
  NAND2_X2 U9081 ( .A1(n6503), .A2(n32199), .ZN(n11897) );
  AOI21_X1 U9082 ( .A1(n22901), .A2(n852), .B(n26507), .ZN(n32199) );
  INV_X2 U9088 ( .I(n32200), .ZN(n27799) );
  XOR2_X1 U9089 ( .A1(n22518), .A2(n22517), .Z(n32200) );
  XOR2_X1 U9095 ( .A1(n7057), .A2(n11219), .Z(n11218) );
  NAND2_X2 U9097 ( .A1(n11178), .A2(n11177), .ZN(n7057) );
  XOR2_X1 U9098 ( .A1(n30041), .A2(n1417), .Z(n27349) );
  NAND2_X2 U9099 ( .A1(n30182), .A2(n29060), .ZN(n30041) );
  NAND2_X2 U9107 ( .A1(n31983), .A2(n6490), .ZN(n14058) );
  XOR2_X1 U9108 ( .A1(n13843), .A2(n19619), .Z(n13842) );
  NAND2_X2 U9109 ( .A1(n28821), .A2(n21437), .ZN(n6544) );
  NAND2_X2 U9110 ( .A1(n19961), .A2(n27491), .ZN(n19962) );
  XOR2_X1 U9111 ( .A1(n188), .A2(n32703), .Z(n11974) );
  XOR2_X1 U9114 ( .A1(n32124), .A2(n12614), .Z(n2900) );
  INV_X2 U9120 ( .I(n32202), .ZN(n8422) );
  XOR2_X1 U9121 ( .A1(Plaintext[61]), .A2(Key[61]), .Z(n32202) );
  XOR2_X1 U9122 ( .A1(n24469), .A2(n14762), .Z(n29809) );
  XOR2_X1 U9123 ( .A1(n2117), .A2(n24545), .Z(n24469) );
  NAND2_X2 U9130 ( .A1(n13340), .A2(n22758), .ZN(n31499) );
  OAI22_X1 U9131 ( .A1(n9792), .A2(n31231), .B1(n2202), .B2(n9793), .ZN(n32204) );
  XOR2_X1 U9133 ( .A1(n20906), .A2(n21003), .Z(n8026) );
  XOR2_X1 U9135 ( .A1(n20970), .A2(n21037), .Z(n20906) );
  AOI21_X1 U9140 ( .A1(n22999), .A2(n9280), .B(n32635), .ZN(n33640) );
  INV_X1 U9141 ( .I(n18269), .ZN(n33613) );
  NAND2_X2 U9146 ( .A1(n32637), .A2(n32205), .ZN(n7831) );
  XOR2_X1 U9147 ( .A1(n15978), .A2(n32206), .Z(n28978) );
  NOR2_X2 U9149 ( .A1(n27353), .A2(n6188), .ZN(n15978) );
  NAND2_X2 U9151 ( .A1(n11023), .A2(n32207), .ZN(n10943) );
  NOR2_X2 U9152 ( .A1(n448), .A2(n30560), .ZN(n32207) );
  NAND2_X2 U9155 ( .A1(n33551), .A2(n12913), .ZN(n32300) );
  NAND3_X2 U9158 ( .A1(n30587), .A2(n17884), .A3(n17883), .ZN(n32974) );
  INV_X2 U9170 ( .I(n23841), .ZN(n32209) );
  XOR2_X1 U9171 ( .A1(n3736), .A2(n32211), .Z(n28605) );
  XOR2_X1 U9173 ( .A1(n3735), .A2(n12618), .Z(n32211) );
  AOI22_X2 U9176 ( .A1(n32494), .A2(n32212), .B1(n6235), .B2(n10993), .ZN(
        n24147) );
  NAND2_X2 U9177 ( .A1(n13031), .A2(n23681), .ZN(n32212) );
  NAND2_X2 U9181 ( .A1(n14752), .A2(n10099), .ZN(n24908) );
  NAND2_X2 U9187 ( .A1(n6471), .A2(n18209), .ZN(n14957) );
  NAND2_X2 U9188 ( .A1(n31995), .A2(n21087), .ZN(n18209) );
  NAND2_X2 U9189 ( .A1(n21688), .A2(n12561), .ZN(n21551) );
  XOR2_X1 U9190 ( .A1(n11332), .A2(n3935), .Z(n10235) );
  NAND3_X2 U9194 ( .A1(n33689), .A2(n29584), .A3(n11331), .ZN(n11332) );
  NAND3_X2 U9196 ( .A1(n25853), .A2(n15546), .A3(n16673), .ZN(n30071) );
  NAND2_X2 U9211 ( .A1(n25834), .A2(n14199), .ZN(n25853) );
  XOR2_X1 U9212 ( .A1(n10582), .A2(n32511), .Z(n10679) );
  AOI21_X2 U9213 ( .A1(n22540), .A2(n22539), .B(n32448), .ZN(n32447) );
  NAND2_X2 U9214 ( .A1(n17147), .A2(n22427), .ZN(n22539) );
  NAND2_X2 U9218 ( .A1(n698), .A2(n29127), .ZN(n32443) );
  XOR2_X1 U9221 ( .A1(n6914), .A2(n32213), .Z(n15356) );
  INV_X2 U9223 ( .I(n2841), .ZN(n14841) );
  XOR2_X1 U9224 ( .A1(n23335), .A2(n32214), .Z(n2841) );
  INV_X1 U9225 ( .I(n6190), .ZN(n32820) );
  NAND2_X2 U9228 ( .A1(n14550), .A2(n14548), .ZN(n16554) );
  NAND2_X2 U9229 ( .A1(n12858), .A2(n27369), .ZN(n14550) );
  NOR2_X2 U9233 ( .A1(n31485), .A2(n32215), .ZN(n16280) );
  NOR2_X2 U9237 ( .A1(n30448), .A2(n33594), .ZN(n32216) );
  OAI21_X1 U9240 ( .A1(n10724), .A2(n22644), .B(n1292), .ZN(n32217) );
  XOR2_X1 U9251 ( .A1(n32220), .A2(n30049), .Z(n33487) );
  XOR2_X1 U9253 ( .A1(n32809), .A2(n32022), .Z(n32220) );
  NAND2_X1 U9254 ( .A1(n22789), .A2(n33388), .ZN(n33387) );
  XOR2_X1 U9258 ( .A1(n23341), .A2(n4564), .Z(n4563) );
  OAI22_X1 U9261 ( .A1(n32221), .A2(n5900), .B1(n5903), .B2(n17838), .ZN(
        n32235) );
  NOR2_X1 U9268 ( .A1(n24994), .A2(n7831), .ZN(n32221) );
  XOR2_X1 U9269 ( .A1(n22243), .A2(n22306), .Z(n21998) );
  NAND2_X2 U9273 ( .A1(n16163), .A2(n16164), .ZN(n22243) );
  XOR2_X1 U9275 ( .A1(n5767), .A2(n7605), .Z(n12871) );
  NAND2_X1 U9277 ( .A1(n32819), .A2(n12848), .ZN(n23170) );
  INV_X1 U9282 ( .I(n15324), .ZN(n32510) );
  XOR2_X1 U9283 ( .A1(n12659), .A2(n32222), .Z(n33662) );
  XOR2_X1 U9284 ( .A1(n2564), .A2(n14613), .Z(n32222) );
  INV_X2 U9285 ( .I(n16554), .ZN(n1086) );
  INV_X2 U9286 ( .I(n32550), .ZN(n32223) );
  NOR2_X2 U9288 ( .A1(n32957), .A2(n11513), .ZN(n32550) );
  NAND2_X2 U9299 ( .A1(n12900), .A2(n18026), .ZN(n31407) );
  NAND3_X1 U9304 ( .A1(n25296), .A2(n25344), .A3(n25397), .ZN(n18026) );
  NOR2_X2 U9306 ( .A1(n24200), .A2(n26027), .ZN(n28505) );
  AOI22_X2 U9309 ( .A1(n738), .A2(n24158), .B1(n7503), .B2(n24008), .ZN(n24200) );
  OAI21_X1 U9313 ( .A1(n14609), .A2(n25005), .B(n42), .ZN(n32227) );
  NAND3_X1 U9316 ( .A1(n32227), .A2(n14607), .A3(n25004), .ZN(n30063) );
  NAND3_X2 U9317 ( .A1(n30922), .A2(n30923), .A3(n6999), .ZN(n6997) );
  NAND2_X2 U9318 ( .A1(n7722), .A2(n32224), .ZN(n16954) );
  AOI22_X2 U9320 ( .A1(n21057), .A2(n11745), .B1(n7721), .B2(n28406), .ZN(
        n32224) );
  INV_X2 U9321 ( .I(n13970), .ZN(n28953) );
  OAI22_X2 U9324 ( .A1(n7157), .A2(n7154), .B1(n7291), .B2(n20604), .ZN(n13970) );
  NAND2_X1 U9329 ( .A1(n32225), .A2(n17383), .ZN(n16284) );
  NAND3_X1 U9334 ( .A1(n17089), .A2(n16661), .A3(n16660), .ZN(n32225) );
  NAND2_X2 U9337 ( .A1(n2529), .A2(n32226), .ZN(n8968) );
  NAND2_X2 U9342 ( .A1(n24289), .A2(n24110), .ZN(n32226) );
  XOR2_X1 U9344 ( .A1(n8761), .A2(n23330), .Z(n26279) );
  XOR2_X1 U9345 ( .A1(n23233), .A2(n23299), .Z(n8761) );
  XOR2_X1 U9346 ( .A1(n23454), .A2(n23474), .Z(n23324) );
  NOR2_X2 U9356 ( .A1(n17585), .A2(n12790), .ZN(n23454) );
  NAND2_X2 U9368 ( .A1(n10784), .A2(n10785), .ZN(n32253) );
  NAND2_X2 U9369 ( .A1(n816), .A2(n17237), .ZN(n9986) );
  NAND3_X2 U9370 ( .A1(n31805), .A2(n8589), .A3(n8592), .ZN(n17237) );
  CLKBUF_X4 U9372 ( .I(n14855), .Z(n4728) );
  AOI22_X2 U9379 ( .A1(n11317), .A2(n8365), .B1(n33563), .B2(n10296), .ZN(
        n32826) );
  XOR2_X1 U9384 ( .A1(n4680), .A2(n20835), .Z(n20993) );
  NOR2_X2 U9388 ( .A1(n4534), .A2(n4535), .ZN(n4680) );
  NOR2_X2 U9390 ( .A1(n33972), .A2(n21188), .ZN(n4494) );
  INV_X2 U9391 ( .I(n32229), .ZN(n32228) );
  OAI21_X2 U9393 ( .A1(n26120), .A2(n6713), .B(n27168), .ZN(n32229) );
  NOR2_X2 U9395 ( .A1(n4956), .A2(n28403), .ZN(n3935) );
  NAND2_X2 U9396 ( .A1(n18298), .A2(n18299), .ZN(n19445) );
  XOR2_X1 U9405 ( .A1(n12622), .A2(n30038), .Z(n625) );
  NAND2_X2 U9406 ( .A1(n32230), .A2(n16857), .ZN(n20733) );
  AOI21_X2 U9410 ( .A1(n22327), .A2(n722), .B(n22328), .ZN(n3512) );
  XOR2_X1 U9411 ( .A1(n19567), .A2(n32231), .Z(n2484) );
  XOR2_X1 U9412 ( .A1(n19386), .A2(n34119), .Z(n19567) );
  NOR2_X1 U9413 ( .A1(n19061), .A2(n19063), .ZN(n28498) );
  NOR2_X1 U9414 ( .A1(n19108), .A2(n5545), .ZN(n19061) );
  XOR2_X1 U9416 ( .A1(n32232), .A2(n1433), .Z(Ciphertext[35]) );
  AOI22_X1 U9417 ( .A1(n25007), .A2(n25008), .B1(n3155), .B2(n29110), .ZN(
        n32232) );
  INV_X2 U9419 ( .I(n5820), .ZN(n32234) );
  XOR2_X1 U9424 ( .A1(n32235), .A2(n1406), .Z(Ciphertext[26]) );
  NAND2_X2 U9429 ( .A1(n29904), .A2(n27840), .ZN(n32240) );
  XOR2_X1 U9432 ( .A1(n12972), .A2(n19529), .Z(n19533) );
  XOR2_X1 U9435 ( .A1(n30539), .A2(n5038), .Z(n11850) );
  XOR2_X1 U9437 ( .A1(n16200), .A2(n33274), .Z(n30539) );
  OAI22_X2 U9440 ( .A1(n14161), .A2(n10978), .B1(n7397), .B2(n32236), .ZN(
        n10159) );
  OAI21_X1 U9441 ( .A1(n1353), .A2(n20627), .B(n20628), .ZN(n32236) );
  AOI22_X2 U9444 ( .A1(n9014), .A2(n7552), .B1(n20627), .B2(n29814), .ZN(
        n10978) );
  XOR2_X1 U9447 ( .A1(n18929), .A2(n19538), .Z(n9636) );
  NAND2_X2 U9455 ( .A1(n28108), .A2(n9637), .ZN(n19538) );
  NAND2_X2 U9461 ( .A1(n2576), .A2(n16023), .ZN(n26386) );
  OAI21_X2 U9465 ( .A1(n14869), .A2(n14871), .B(n21684), .ZN(n22295) );
  NOR2_X2 U9466 ( .A1(n14292), .A2(n32237), .ZN(n2577) );
  NOR3_X2 U9467 ( .A1(n33641), .A2(n28287), .A3(n11915), .ZN(n32237) );
  XOR2_X1 U9469 ( .A1(n32238), .A2(n13886), .Z(n27503) );
  XOR2_X1 U9470 ( .A1(n21039), .A2(n20799), .Z(n32238) );
  XOR2_X1 U9472 ( .A1(n2920), .A2(n4362), .Z(n9161) );
  NOR2_X2 U9473 ( .A1(n5872), .A2(n4150), .ZN(n2920) );
  NOR2_X2 U9474 ( .A1(n12522), .A2(n11181), .ZN(n11180) );
  OR2_X2 U9477 ( .A1(n16), .A2(n11913), .Z(n4371) );
  XOR2_X1 U9478 ( .A1(n887), .A2(n5297), .Z(n5296) );
  XNOR2_X1 U9479 ( .A1(n5482), .A2(n34016), .ZN(n22164) );
  NOR2_X2 U9480 ( .A1(n27053), .A2(n21831), .ZN(n34016) );
  AOI22_X2 U9482 ( .A1(n32241), .A2(n21321), .B1(n4382), .B2(n21324), .ZN(
        n30745) );
  NOR2_X2 U9484 ( .A1(n15015), .A2(n28017), .ZN(n32241) );
  NAND2_X2 U9485 ( .A1(n21727), .A2(n21728), .ZN(n5482) );
  AOI21_X1 U9486 ( .A1(n5112), .A2(n315), .B(n314), .ZN(n32244) );
  NAND2_X2 U9487 ( .A1(n5789), .A2(n31948), .ZN(n19243) );
  NAND2_X2 U9488 ( .A1(n5155), .A2(n5154), .ZN(n5789) );
  NAND2_X1 U9492 ( .A1(n23826), .A2(n16467), .ZN(n27734) );
  AOI22_X1 U9496 ( .A1(n17760), .A2(n31907), .B1(n15282), .B2(n14365), .ZN(
        n14470) );
  NAND2_X2 U9499 ( .A1(n16804), .A2(n15198), .ZN(n31907) );
  OAI21_X2 U9506 ( .A1(n9652), .A2(n26081), .B(n26518), .ZN(n31036) );
  NOR2_X2 U9508 ( .A1(n33718), .A2(n6290), .ZN(n26081) );
  NAND2_X2 U9509 ( .A1(n27079), .A2(n6189), .ZN(n23474) );
  OAI22_X2 U9510 ( .A1(n23832), .A2(n7005), .B1(n15623), .B2(n34167), .ZN(
        n13936) );
  INV_X2 U9511 ( .I(n23587), .ZN(n7005) );
  AND2_X1 U9513 ( .A1(n22640), .A2(n11749), .Z(n14830) );
  XOR2_X1 U9514 ( .A1(n23280), .A2(n11326), .Z(n47) );
  XOR2_X1 U9517 ( .A1(n30315), .A2(n23405), .Z(n23280) );
  NAND2_X1 U9519 ( .A1(n22748), .A2(n30231), .ZN(n23027) );
  NOR2_X2 U9523 ( .A1(n22729), .A2(n22731), .ZN(n30231) );
  INV_X1 U9524 ( .I(n7052), .ZN(n33183) );
  OAI21_X2 U9526 ( .A1(n11280), .A2(n10828), .B(n11278), .ZN(n18669) );
  XNOR2_X1 U9527 ( .A1(n16641), .A2(n16472), .ZN(n32251) );
  XOR2_X1 U9528 ( .A1(n9877), .A2(n32245), .Z(n21330) );
  XOR2_X1 U9531 ( .A1(n32614), .A2(n30045), .Z(n32245) );
  NOR3_X2 U9535 ( .A1(n32246), .A2(n26465), .A3(n26464), .ZN(n11845) );
  NOR2_X1 U9538 ( .A1(n3289), .A2(n3288), .ZN(n32246) );
  XOR2_X1 U9548 ( .A1(n30997), .A2(n1396), .Z(n6852) );
  NOR2_X2 U9552 ( .A1(n31032), .A2(n34148), .ZN(n30997) );
  AOI21_X2 U9553 ( .A1(n32247), .A2(n33223), .B(n31293), .ZN(n24330) );
  AOI21_X1 U9554 ( .A1(n33144), .A2(n3860), .B(n14335), .ZN(n32247) );
  NAND2_X2 U9555 ( .A1(n23885), .A2(n15266), .ZN(n17777) );
  NAND2_X1 U9556 ( .A1(n17502), .A2(n32438), .ZN(n32338) );
  XOR2_X1 U9557 ( .A1(n22061), .A2(n22109), .Z(n5353) );
  XOR2_X1 U9561 ( .A1(n1310), .A2(n5476), .Z(n22109) );
  XOR2_X1 U9565 ( .A1(n5186), .A2(n28315), .Z(n20716) );
  XOR2_X1 U9566 ( .A1(n28953), .A2(n2356), .Z(n5186) );
  BUF_X2 U9569 ( .I(n17439), .Z(n32248) );
  AOI21_X2 U9571 ( .A1(n20186), .A2(n20187), .B(n32249), .ZN(n7889) );
  XOR2_X1 U9574 ( .A1(n28621), .A2(n32250), .Z(n26162) );
  XOR2_X1 U9580 ( .A1(n20806), .A2(n32251), .Z(n32250) );
  NAND2_X2 U9581 ( .A1(n13989), .A2(n32147), .ZN(n29802) );
  NAND2_X2 U9584 ( .A1(n11300), .A2(n32254), .ZN(n32535) );
  OAI22_X2 U9589 ( .A1(n31604), .A2(n11306), .B1(n12000), .B2(n32585), .ZN(
        n13483) );
  INV_X1 U9590 ( .I(n27152), .ZN(n33943) );
  OAI21_X2 U9594 ( .A1(n26337), .A2(n11301), .B(n29997), .ZN(n32254) );
  BUF_X4 U9598 ( .I(n28278), .Z(n33981) );
  OAI22_X2 U9599 ( .A1(n1125), .A2(n5440), .B1(n22588), .B2(n22589), .ZN(
        n12899) );
  XOR2_X1 U9600 ( .A1(n2653), .A2(n32906), .Z(n23290) );
  NAND2_X1 U9601 ( .A1(n8373), .A2(n16154), .ZN(n9151) );
  XOR2_X1 U9602 ( .A1(n28814), .A2(n32256), .Z(n4798) );
  XOR2_X1 U9603 ( .A1(n28354), .A2(n20974), .Z(n32256) );
  OAI22_X2 U9607 ( .A1(n5782), .A2(n27876), .B1(n266), .B2(n20495), .ZN(n5668)
         );
  NOR2_X2 U9608 ( .A1(n32257), .A2(n29354), .ZN(n28733) );
  NOR2_X2 U9609 ( .A1(n9364), .A2(n31721), .ZN(n32257) );
  INV_X2 U9613 ( .I(n8862), .ZN(n33884) );
  NAND2_X2 U9616 ( .A1(n33022), .A2(n17327), .ZN(n32258) );
  XOR2_X1 U9617 ( .A1(n32259), .A2(n4704), .Z(n7896) );
  OAI21_X2 U9619 ( .A1(n18959), .A2(n4622), .B(n4619), .ZN(n32259) );
  NOR2_X2 U9620 ( .A1(n4390), .A2(n32260), .ZN(n21842) );
  AOI21_X1 U9622 ( .A1(n3916), .A2(n14482), .B(n33454), .ZN(n32260) );
  NAND2_X2 U9623 ( .A1(n1965), .A2(n32261), .ZN(n6357) );
  NOR2_X2 U9627 ( .A1(n1968), .A2(n1967), .ZN(n32261) );
  XOR2_X1 U9629 ( .A1(n32262), .A2(n25993), .Z(n19565) );
  AOI21_X2 U9633 ( .A1(n31349), .A2(n14606), .B(n19303), .ZN(n25993) );
  INV_X2 U9638 ( .I(n19483), .ZN(n32262) );
  OAI21_X2 U9640 ( .A1(n13414), .A2(n1519), .B(n32754), .ZN(n28839) );
  OAI21_X2 U9643 ( .A1(n12312), .A2(n32263), .B(n6003), .ZN(n31718) );
  NOR2_X2 U9644 ( .A1(n32264), .A2(n24097), .ZN(n32263) );
  INV_X2 U9646 ( .I(n32917), .ZN(n32264) );
  NAND2_X2 U9647 ( .A1(n22765), .A2(n29795), .ZN(n29634) );
  NAND2_X2 U9649 ( .A1(n23631), .A2(n32265), .ZN(n24286) );
  NAND2_X2 U9652 ( .A1(n32426), .A2(n6392), .ZN(n32265) );
  OAI21_X2 U9654 ( .A1(n33470), .A2(n31788), .B(n32266), .ZN(n24761) );
  NAND2_X1 U9657 ( .A1(n1640), .A2(n14447), .ZN(n32266) );
  INV_X2 U9658 ( .I(n29540), .ZN(n15708) );
  XOR2_X1 U9662 ( .A1(n32267), .A2(n19368), .Z(n29540) );
  INV_X2 U9663 ( .I(n6387), .ZN(n32267) );
  INV_X2 U9665 ( .I(n24914), .ZN(n24911) );
  NAND2_X2 U9666 ( .A1(n29877), .A2(n17304), .ZN(n24914) );
  INV_X1 U9669 ( .I(n23729), .ZN(n30477) );
  NAND2_X1 U9670 ( .A1(n15722), .A2(n30949), .ZN(n23729) );
  AOI22_X2 U9671 ( .A1(n1219), .A2(n9862), .B1(n837), .B2(n9861), .ZN(n33737)
         );
  XOR2_X1 U9672 ( .A1(n7250), .A2(n22125), .Z(n3395) );
  NAND2_X2 U9673 ( .A1(n11585), .A2(n6076), .ZN(n7250) );
  XOR2_X1 U9676 ( .A1(n32268), .A2(n23375), .Z(n33710) );
  XOR2_X1 U9680 ( .A1(n23376), .A2(n23475), .Z(n32268) );
  NAND2_X2 U9681 ( .A1(n33239), .A2(n32269), .ZN(n24896) );
  NAND3_X1 U9685 ( .A1(n24477), .A2(n24591), .A3(n25013), .ZN(n32269) );
  BUF_X2 U9688 ( .I(n3964), .Z(n32271) );
  XOR2_X1 U9697 ( .A1(n32272), .A2(n25554), .Z(Ciphertext[123]) );
  INV_X1 U9699 ( .I(n31389), .ZN(n33357) );
  INV_X2 U9700 ( .I(n20581), .ZN(n936) );
  NAND2_X2 U9704 ( .A1(n9449), .A2(n19657), .ZN(n20581) );
  INV_X4 U9708 ( .I(n24326), .ZN(n24325) );
  NAND2_X2 U9710 ( .A1(n32274), .A2(n33335), .ZN(n33980) );
  NAND2_X2 U9713 ( .A1(n10353), .A2(n10352), .ZN(n32274) );
  NAND3_X2 U9715 ( .A1(n10261), .A2(n6599), .A3(n28395), .ZN(n33286) );
  NAND2_X2 U9716 ( .A1(n32275), .A2(n27269), .ZN(n17637) );
  AOI22_X2 U9717 ( .A1(n15979), .A2(n15964), .B1(n24865), .B2(n26912), .ZN(
        n32275) );
  NAND2_X2 U9720 ( .A1(n27856), .A2(n27916), .ZN(n27419) );
  INV_X1 U9721 ( .I(n20798), .ZN(n32392) );
  NAND2_X1 U9723 ( .A1(n32278), .A2(n32276), .ZN(n19457) );
  INV_X1 U9727 ( .I(n8770), .ZN(n32277) );
  NAND2_X1 U9728 ( .A1(n1034), .A2(n8770), .ZN(n32278) );
  NAND2_X2 U9732 ( .A1(n27337), .A2(n21394), .ZN(n14095) );
  OAI21_X1 U9735 ( .A1(n25740), .A2(n27189), .B(n32279), .ZN(n6524) );
  XOR2_X1 U9736 ( .A1(n5024), .A2(n20885), .Z(n15875) );
  NAND2_X2 U9738 ( .A1(n2292), .A2(n2293), .ZN(n20549) );
  AOI21_X2 U9739 ( .A1(n24269), .A2(n24268), .B(n11721), .ZN(n11723) );
  NAND2_X2 U9741 ( .A1(n32280), .A2(n33821), .ZN(n26445) );
  NAND2_X1 U9743 ( .A1(n30562), .A2(n14803), .ZN(n32280) );
  NOR2_X2 U9745 ( .A1(n15326), .A2(n15327), .ZN(n33646) );
  AOI22_X2 U9746 ( .A1(n26633), .A2(n20577), .B1(n20481), .B2(n20480), .ZN(
        n6228) );
  INV_X2 U9754 ( .I(n12008), .ZN(n4674) );
  NAND2_X1 U9757 ( .A1(n28645), .A2(n20067), .ZN(n26741) );
  NAND2_X2 U9763 ( .A1(n942), .A2(n19947), .ZN(n19948) );
  NAND2_X2 U9766 ( .A1(n7799), .A2(n32281), .ZN(n7798) );
  NAND2_X2 U9768 ( .A1(n20487), .A2(n9808), .ZN(n32281) );
  OR2_X1 U9769 ( .A1(n24153), .A2(n839), .Z(n32962) );
  NOR2_X1 U9770 ( .A1(n6326), .A2(n6325), .ZN(n6982) );
  XOR2_X1 U9774 ( .A1(n32283), .A2(n19412), .Z(n1694) );
  AOI21_X2 U9775 ( .A1(n18938), .A2(n29), .B(n18937), .ZN(n19412) );
  INV_X1 U9777 ( .I(n19400), .ZN(n32283) );
  NAND2_X2 U9778 ( .A1(n3983), .A2(n11654), .ZN(n31155) );
  XOR2_X1 U9784 ( .A1(n32284), .A2(n8487), .Z(Ciphertext[64]) );
  NAND3_X2 U9786 ( .A1(n8340), .A2(n8928), .A3(n8339), .ZN(n32284) );
  XOR2_X1 U9788 ( .A1(n32285), .A2(n7665), .Z(n7700) );
  XOR2_X1 U9791 ( .A1(n23424), .A2(n23307), .Z(n32285) );
  AOI22_X2 U9793 ( .A1(n7719), .A2(n16174), .B1(n34052), .B2(n20515), .ZN(
        n2251) );
  NAND2_X2 U9794 ( .A1(n3725), .A2(n3724), .ZN(n4782) );
  NOR2_X2 U9797 ( .A1(n9615), .A2(n9609), .ZN(n3725) );
  NAND2_X2 U9798 ( .A1(n31282), .A2(n22464), .ZN(n22962) );
  OAI21_X2 U9800 ( .A1(n16288), .A2(n25999), .B(n8233), .ZN(n16068) );
  XOR2_X1 U9802 ( .A1(n17004), .A2(n9440), .Z(n16689) );
  AND2_X1 U9811 ( .A1(n21357), .A2(n21358), .Z(n11655) );
  NAND2_X2 U9814 ( .A1(n32287), .A2(n3451), .ZN(n5915) );
  OAI21_X2 U9815 ( .A1(n3454), .A2(n3596), .B(n31931), .ZN(n32287) );
  INV_X4 U9816 ( .I(n29980), .ZN(n28581) );
  NAND2_X2 U9818 ( .A1(n30972), .A2(n28523), .ZN(n29980) );
  XOR2_X1 U9819 ( .A1(n4883), .A2(n19705), .Z(n3416) );
  XOR2_X1 U9820 ( .A1(n12779), .A2(n16150), .Z(n33804) );
  NAND2_X2 U9822 ( .A1(n8478), .A2(n4114), .ZN(n33069) );
  AOI22_X2 U9824 ( .A1(n31919), .A2(n24292), .B1(n7779), .B2(n26544), .ZN(
        n32288) );
  NAND2_X2 U9825 ( .A1(n14711), .A2(n14712), .ZN(n20414) );
  NOR2_X2 U9826 ( .A1(n5820), .A2(n16976), .ZN(n22772) );
  INV_X1 U9829 ( .I(n2913), .ZN(n32299) );
  NAND2_X2 U9830 ( .A1(n33458), .A2(n32298), .ZN(n32289) );
  NAND2_X2 U9831 ( .A1(n16787), .A2(n32329), .ZN(n26485) );
  NAND2_X2 U9833 ( .A1(n11035), .A2(n11036), .ZN(n16787) );
  INV_X4 U9835 ( .I(n33035), .ZN(n15027) );
  NAND2_X2 U9836 ( .A1(n18170), .A2(n18171), .ZN(n20208) );
  AOI21_X1 U9837 ( .A1(n16444), .A2(n19061), .B(n32290), .ZN(n7591) );
  NOR2_X1 U9839 ( .A1(n29213), .A2(n571), .ZN(n29423) );
  NOR2_X1 U9841 ( .A1(n26406), .A2(n16148), .ZN(n32406) );
  NAND2_X2 U9843 ( .A1(n32291), .A2(n20884), .ZN(n21693) );
  AOI22_X2 U9844 ( .A1(n812), .A2(n20881), .B1(n21163), .B2(n21367), .ZN(
        n32291) );
  OAI21_X2 U9845 ( .A1(n33488), .A2(n31239), .B(n29964), .ZN(n31497) );
  OR2_X1 U9846 ( .A1(n19122), .A2(n16361), .Z(n32292) );
  NAND2_X2 U9854 ( .A1(n10043), .A2(n18617), .ZN(n18615) );
  XOR2_X1 U9855 ( .A1(n8392), .A2(n22032), .Z(n22154) );
  NAND2_X2 U9856 ( .A1(n3702), .A2(n33315), .ZN(n8392) );
  XOR2_X1 U9858 ( .A1(n26272), .A2(n6031), .Z(n11006) );
  OAI21_X2 U9860 ( .A1(n14536), .A2(n31115), .B(n32294), .ZN(n10055) );
  XOR2_X1 U9863 ( .A1(n3267), .A2(n32295), .Z(n29470) );
  XOR2_X1 U9864 ( .A1(n17859), .A2(n23400), .Z(n32295) );
  BUF_X2 U9866 ( .I(n1164), .Z(n32296) );
  NAND2_X2 U9871 ( .A1(n32297), .A2(n4816), .ZN(n15275) );
  OAI22_X2 U9872 ( .A1(n20479), .A2(n20403), .B1(n20571), .B2(n31968), .ZN(
        n32297) );
  XOR2_X1 U9873 ( .A1(n31523), .A2(n16578), .Z(n2875) );
  NAND2_X2 U9875 ( .A1(n4846), .A2(n4847), .ZN(n31523) );
  NOR2_X2 U9882 ( .A1(n26595), .A2(n32300), .ZN(n13884) );
  NOR2_X2 U9884 ( .A1(n32384), .A2(n8029), .ZN(n32301) );
  NOR2_X2 U9885 ( .A1(n10862), .A2(n26410), .ZN(n22401) );
  XOR2_X1 U9889 ( .A1(n28315), .A2(n20873), .Z(n32726) );
  INV_X2 U9890 ( .I(n16805), .ZN(n18677) );
  XOR2_X1 U9892 ( .A1(Plaintext[2]), .A2(Key[2]), .Z(n16805) );
  XOR2_X1 U9897 ( .A1(n9018), .A2(n32302), .Z(n33331) );
  XOR2_X1 U9899 ( .A1(n23355), .A2(n23292), .Z(n11249) );
  XOR2_X1 U9900 ( .A1(n27423), .A2(n18028), .Z(n24561) );
  AOI21_X2 U9912 ( .A1(n342), .A2(n30579), .B(n33124), .ZN(n27423) );
  XOR2_X1 U9913 ( .A1(n32303), .A2(n16497), .Z(Ciphertext[108]) );
  NAND3_X1 U9918 ( .A1(n31492), .A2(n25482), .A3(n25458), .ZN(n32303) );
  NAND2_X2 U9920 ( .A1(n32304), .A2(n31078), .ZN(n20996) );
  NAND2_X2 U9921 ( .A1(n17496), .A2(n32305), .ZN(n17497) );
  AOI22_X2 U9932 ( .A1(n29338), .A2(n34152), .B1(n12075), .B2(n20052), .ZN(
        n32305) );
  XOR2_X1 U9938 ( .A1(n24691), .A2(n5762), .Z(n30563) );
  NAND2_X2 U9949 ( .A1(n32725), .A2(n31171), .ZN(n24691) );
  NAND3_X1 U9952 ( .A1(n25285), .A2(n16291), .A3(n25276), .ZN(n11257) );
  NAND2_X2 U9954 ( .A1(n10743), .A2(n33330), .ZN(n16291) );
  XOR2_X1 U9955 ( .A1(n32306), .A2(n16705), .Z(Ciphertext[134]) );
  NAND2_X1 U9957 ( .A1(n13996), .A2(n28775), .ZN(n32306) );
  NAND3_X2 U9961 ( .A1(n29741), .A2(n11109), .A3(n11108), .ZN(n23358) );
  NAND2_X1 U9962 ( .A1(n15241), .A2(n15242), .ZN(n34000) );
  OAI22_X2 U9967 ( .A1(n19329), .A2(n2040), .B1(n19328), .B2(n7732), .ZN(
        n18103) );
  INV_X1 U9969 ( .I(n20911), .ZN(n32342) );
  BUF_X4 U9971 ( .I(n28839), .Z(n33022) );
  NAND2_X1 U9973 ( .A1(n22885), .A2(n1577), .ZN(n32307) );
  NOR2_X2 U9975 ( .A1(n32308), .A2(n10193), .ZN(n6320) );
  NAND2_X2 U9976 ( .A1(n14412), .A2(n14410), .ZN(n11651) );
  NOR2_X2 U9977 ( .A1(n26079), .A2(n14249), .ZN(n14412) );
  AND2_X1 U9982 ( .A1(n28697), .A2(n22982), .Z(n22837) );
  NAND3_X1 U9985 ( .A1(n12293), .A2(n12295), .A3(n17928), .ZN(n32583) );
  XOR2_X1 U9987 ( .A1(n22075), .A2(n22141), .Z(n22267) );
  AOI22_X2 U9988 ( .A1(n6968), .A2(n15676), .B1(n12794), .B2(n6967), .ZN(
        n22141) );
  NOR2_X2 U9989 ( .A1(n27501), .A2(n24158), .ZN(n24067) );
  XOR2_X1 U9990 ( .A1(n13645), .A2(n19624), .Z(n16080) );
  AOI21_X2 U10002 ( .A1(n8906), .A2(n11955), .B(n30209), .ZN(n13645) );
  NAND2_X2 U10003 ( .A1(n32312), .A2(n32311), .ZN(n25816) );
  INV_X2 U10006 ( .I(n32313), .ZN(n14661) );
  XNOR2_X1 U10009 ( .A1(n6721), .A2(n6719), .ZN(n32313) );
  NAND3_X2 U10010 ( .A1(n32314), .A2(n6176), .A3(n16601), .ZN(n18163) );
  OR2_X2 U10012 ( .A1(n9717), .A2(n32315), .Z(n691) );
  OAI22_X1 U10015 ( .A1(n28283), .A2(n2378), .B1(n12230), .B2(n10497), .ZN(
        n32315) );
  AOI22_X2 U10017 ( .A1(n22780), .A2(n11983), .B1(n31824), .B2(n22848), .ZN(
        n22889) );
  OR2_X1 U10025 ( .A1(n7581), .A2(n1808), .Z(n33894) );
  NAND2_X2 U10033 ( .A1(n6581), .A2(n32317), .ZN(n23981) );
  XOR2_X1 U10035 ( .A1(n1991), .A2(n32316), .Z(n33082) );
  XOR2_X1 U10036 ( .A1(n1990), .A2(n31928), .Z(n32316) );
  INV_X2 U10037 ( .I(n7188), .ZN(n32317) );
  NAND2_X2 U10038 ( .A1(n32453), .A2(n3950), .ZN(n6555) );
  NAND4_X1 U10040 ( .A1(n6730), .A2(n4056), .A3(n25572), .A4(n25573), .ZN(
        n32702) );
  NAND2_X2 U10050 ( .A1(n15060), .A2(n11953), .ZN(n15059) );
  NOR2_X2 U10052 ( .A1(n22704), .A2(n32318), .ZN(n30532) );
  XOR2_X1 U10053 ( .A1(n32319), .A2(n3605), .Z(n11110) );
  XOR2_X1 U10056 ( .A1(n22000), .A2(n12882), .Z(n32319) );
  NAND2_X1 U10057 ( .A1(n17240), .A2(n11974), .ZN(n24484) );
  XOR2_X1 U10059 ( .A1(n24638), .A2(n24474), .Z(n24773) );
  AOI22_X2 U10061 ( .A1(n14847), .A2(n29566), .B1(n23781), .B2(n17280), .ZN(
        n24638) );
  NAND2_X2 U10062 ( .A1(n32322), .A2(n33171), .ZN(n3963) );
  NAND2_X2 U10066 ( .A1(n32877), .A2(n24060), .ZN(n12644) );
  AND2_X2 U10071 ( .A1(n652), .A2(n23201), .Z(n23796) );
  NAND2_X1 U10075 ( .A1(n15211), .A2(n28078), .ZN(n26068) );
  AOI21_X2 U10076 ( .A1(n29648), .A2(n32089), .B(n32324), .ZN(n16635) );
  XOR2_X1 U10079 ( .A1(n4314), .A2(n19370), .Z(n19742) );
  AOI21_X2 U10084 ( .A1(n7186), .A2(n7187), .B(n7185), .ZN(n4314) );
  XOR2_X1 U10088 ( .A1(n1085), .A2(n5539), .Z(n30917) );
  NOR2_X2 U10090 ( .A1(n17822), .A2(n32325), .ZN(n10735) );
  BUF_X2 U10091 ( .I(n32807), .Z(n32326) );
  AOI21_X2 U10092 ( .A1(n13227), .A2(n16485), .B(n32327), .ZN(n19583) );
  AOI21_X2 U10096 ( .A1(n19186), .A2(n13226), .B(n13685), .ZN(n32327) );
  NAND2_X2 U10103 ( .A1(n9995), .A2(n9998), .ZN(n24110) );
  NOR2_X2 U10107 ( .A1(n22483), .A2(n22372), .ZN(n33864) );
  INV_X8 U10110 ( .I(n18515), .ZN(n829) );
  AOI22_X2 U10112 ( .A1(n33240), .A2(n11666), .B1(n16492), .B2(n20227), .ZN(
        n11665) );
  NOR2_X2 U10113 ( .A1(n32326), .A2(n11364), .ZN(n1361) );
  XOR2_X1 U10114 ( .A1(n27192), .A2(n5322), .Z(n32807) );
  AOI22_X2 U10116 ( .A1(n30507), .A2(n1290), .B1(n22439), .B2(n12899), .ZN(
        n23018) );
  NAND2_X2 U10125 ( .A1(n12434), .A2(n27551), .ZN(n14619) );
  NOR2_X1 U10127 ( .A1(n8994), .A2(n20319), .ZN(n32440) );
  AOI21_X2 U10128 ( .A1(n19270), .A2(n19271), .B(n19269), .ZN(n19272) );
  NAND2_X2 U10130 ( .A1(n15961), .A2(n32330), .ZN(n21553) );
  NAND2_X2 U10133 ( .A1(n32670), .A2(n32331), .ZN(n9408) );
  OR2_X1 U10137 ( .A1(n27131), .A2(n19275), .Z(n32332) );
  INV_X4 U10141 ( .I(n31579), .ZN(n18643) );
  NOR2_X2 U10142 ( .A1(n1008), .A2(n32333), .ZN(n33298) );
  NAND2_X2 U10169 ( .A1(n10699), .A2(n915), .ZN(n32333) );
  OAI21_X1 U10170 ( .A1(n1581), .A2(n5260), .B(n5259), .ZN(n5261) );
  XOR2_X1 U10171 ( .A1(n11297), .A2(n24520), .Z(n24654) );
  NAND2_X2 U10173 ( .A1(n30732), .A2(n17233), .ZN(n11297) );
  NOR2_X1 U10176 ( .A1(n32335), .A2(n32334), .ZN(n8222) );
  NOR2_X1 U10178 ( .A1(n9456), .A2(n22660), .ZN(n32335) );
  XOR2_X1 U10179 ( .A1(n15606), .A2(n31457), .Z(n22182) );
  NAND2_X2 U10185 ( .A1(n12273), .A2(n9448), .ZN(n15606) );
  NAND3_X2 U10192 ( .A1(n20351), .A2(n28813), .A3(n20350), .ZN(n12364) );
  OAI22_X2 U10194 ( .A1(n25456), .A2(n32869), .B1(n25454), .B2(n25455), .ZN(
        n33248) );
  NOR2_X2 U10195 ( .A1(n408), .A2(n25433), .ZN(n25456) );
  XOR2_X1 U10202 ( .A1(n7889), .A2(n20961), .Z(n21025) );
  NAND3_X1 U10247 ( .A1(n891), .A2(n24221), .A3(n2539), .ZN(n9542) );
  INV_X1 U10254 ( .I(n8168), .ZN(n30285) );
  XOR2_X1 U10262 ( .A1(n6267), .A2(n12083), .Z(n17044) );
  AOI22_X2 U10264 ( .A1(n11566), .A2(n11565), .B1(n11564), .B2(n22705), .ZN(
        n32705) );
  NAND2_X2 U10265 ( .A1(n11132), .A2(n25289), .ZN(n25290) );
  NAND2_X2 U10270 ( .A1(n32338), .A2(n22755), .ZN(n12821) );
  OAI22_X2 U10271 ( .A1(n32339), .A2(n8614), .B1(n8613), .B2(n31271), .ZN(
        n12593) );
  NOR2_X2 U10272 ( .A1(n1978), .A2(n8615), .ZN(n32339) );
  INV_X1 U10276 ( .I(n23369), .ZN(n33929) );
  XOR2_X1 U10282 ( .A1(n24650), .A2(n32340), .Z(n28443) );
  XOR2_X1 U10283 ( .A1(n28579), .A2(n29589), .Z(n32340) );
  XOR2_X1 U10284 ( .A1(n6731), .A2(n19730), .Z(n26702) );
  XOR2_X1 U10288 ( .A1(n19558), .A2(n19474), .Z(n19730) );
  NAND2_X2 U10289 ( .A1(n27832), .A2(n29200), .ZN(n33875) );
  NAND2_X2 U10291 ( .A1(n9610), .A2(n2456), .ZN(n3724) );
  OR2_X2 U10293 ( .A1(n6359), .A2(n2019), .Z(n10844) );
  XOR2_X1 U10295 ( .A1(n1622), .A2(n1621), .Z(n11628) );
  XOR2_X1 U10300 ( .A1(n32342), .A2(n7630), .Z(n6159) );
  NAND2_X2 U10303 ( .A1(n6157), .A2(n4269), .ZN(n7630) );
  AND2_X1 U10305 ( .A1(n20097), .A2(n27832), .Z(n8146) );
  NAND2_X2 U10306 ( .A1(n4708), .A2(n32343), .ZN(n5091) );
  XOR2_X1 U10307 ( .A1(n24021), .A2(n32345), .Z(n26126) );
  XOR2_X1 U10308 ( .A1(n2278), .A2(n32346), .Z(n32345) );
  NAND3_X1 U10313 ( .A1(n5471), .A2(n20375), .A3(n10939), .ZN(n2317) );
  NAND2_X1 U10314 ( .A1(n9259), .A2(n30838), .ZN(n7278) );
  INV_X2 U10315 ( .I(n29215), .ZN(n6842) );
  NAND2_X1 U10316 ( .A1(n32347), .A2(n29215), .ZN(n30852) );
  XOR2_X1 U10337 ( .A1(n6843), .A2(n32464), .Z(n29215) );
  INV_X2 U10339 ( .I(n6855), .ZN(n32347) );
  NAND2_X1 U10345 ( .A1(n32617), .A2(n28554), .ZN(n22329) );
  NAND2_X2 U10346 ( .A1(n32348), .A2(n32039), .ZN(n21544) );
  NAND2_X2 U10347 ( .A1(n32506), .A2(n32505), .ZN(n26206) );
  BUF_X2 U10348 ( .I(n24207), .Z(n32349) );
  INV_X1 U10351 ( .I(n27842), .ZN(n32351) );
  AOI22_X2 U10353 ( .A1(n7262), .A2(n28265), .B1(n707), .B2(n7263), .ZN(n7261)
         );
  INV_X2 U10354 ( .I(n32352), .ZN(n29272) );
  XNOR2_X1 U10356 ( .A1(n7711), .A2(n33118), .ZN(n32352) );
  XOR2_X1 U10357 ( .A1(n32353), .A2(n3648), .Z(n28554) );
  XOR2_X1 U10375 ( .A1(n33408), .A2(n22070), .Z(n32353) );
  NOR2_X2 U10376 ( .A1(n5570), .A2(n32355), .ZN(n17273) );
  NOR3_X1 U10378 ( .A1(n26015), .A2(n15738), .A3(n25229), .ZN(n32355) );
  XOR2_X1 U10380 ( .A1(n18929), .A2(n30075), .Z(n30074) );
  XOR2_X1 U10384 ( .A1(n32356), .A2(n23311), .Z(n23827) );
  XOR2_X1 U10386 ( .A1(n33236), .A2(n14841), .Z(n32356) );
  XOR2_X1 U10387 ( .A1(n32722), .A2(n10236), .Z(n28514) );
  OR2_X1 U10388 ( .A1(n32919), .A2(n17439), .Z(n2831) );
  OAI21_X2 U10389 ( .A1(n11976), .A2(n883), .B(n32359), .ZN(n29754) );
  OAI21_X2 U10390 ( .A1(n4318), .A2(n15152), .B(n883), .ZN(n32359) );
  NAND3_X1 U10392 ( .A1(n26206), .A2(n26207), .A3(n1012), .ZN(n32688) );
  OAI21_X2 U10395 ( .A1(n29758), .A2(n29469), .B(n22459), .ZN(n14129) );
  XOR2_X1 U10405 ( .A1(n8018), .A2(n32360), .Z(n31771) );
  XOR2_X1 U10406 ( .A1(n34047), .A2(n7045), .Z(n32360) );
  INV_X1 U10409 ( .I(n21248), .ZN(n29142) );
  NAND2_X1 U10411 ( .A1(n13432), .A2(n13433), .ZN(n33133) );
  OR2_X1 U10412 ( .A1(n28308), .A2(n7368), .Z(n3889) );
  XOR2_X1 U10414 ( .A1(n32361), .A2(n25049), .Z(Ciphertext[39]) );
  NAND3_X2 U10418 ( .A1(n25048), .A2(n28220), .A3(n25046), .ZN(n32361) );
  NOR2_X1 U10419 ( .A1(n23793), .A2(n23794), .ZN(n1876) );
  XOR2_X1 U10421 ( .A1(n32362), .A2(n10951), .Z(n589) );
  XOR2_X1 U10424 ( .A1(n28295), .A2(n25578), .Z(n32362) );
  NAND2_X2 U10429 ( .A1(n27299), .A2(n4241), .ZN(n20900) );
  AOI21_X2 U10440 ( .A1(n23482), .A2(n7220), .B(n11956), .ZN(n9212) );
  AND2_X2 U10443 ( .A1(n15559), .A2(n21193), .Z(n21072) );
  XOR2_X1 U10444 ( .A1(n7880), .A2(n32363), .Z(n30173) );
  XOR2_X1 U10448 ( .A1(n6545), .A2(n2045), .Z(n32363) );
  NAND2_X1 U10449 ( .A1(n29753), .A2(n793), .ZN(n32369) );
  XOR2_X1 U10451 ( .A1(n32364), .A2(n23245), .Z(n22935) );
  XOR2_X1 U10452 ( .A1(n33380), .A2(n22932), .Z(n32364) );
  NOR2_X1 U10453 ( .A1(n4386), .A2(n4387), .ZN(n32612) );
  NOR2_X1 U10460 ( .A1(n22953), .A2(n7544), .ZN(n8082) );
  NAND2_X2 U10461 ( .A1(n16267), .A2(n30584), .ZN(n7544) );
  BUF_X4 U10463 ( .I(n3286), .Z(n21) );
  NAND2_X2 U10465 ( .A1(n11710), .A2(n20549), .ZN(n20327) );
  NAND2_X2 U10466 ( .A1(n2285), .A2(n26814), .ZN(n11710) );
  NAND2_X2 U10467 ( .A1(n3760), .A2(n981), .ZN(n23815) );
  AND2_X1 U10468 ( .A1(n11734), .A2(n17522), .Z(n2603) );
  XOR2_X1 U10470 ( .A1(n20803), .A2(n20802), .Z(n21012) );
  NAND2_X2 U10474 ( .A1(n20218), .A2(n20217), .ZN(n20803) );
  XOR2_X1 U10476 ( .A1(n33317), .A2(n26642), .Z(n17506) );
  XOR2_X1 U10477 ( .A1(n32365), .A2(n8464), .Z(n14934) );
  XOR2_X1 U10482 ( .A1(n21033), .A2(n15793), .Z(n32365) );
  XOR2_X1 U10483 ( .A1(n32366), .A2(n4610), .Z(n32489) );
  XOR2_X1 U10484 ( .A1(n27481), .A2(n7046), .Z(n32366) );
  BUF_X2 U10487 ( .I(n19749), .Z(n32367) );
  XOR2_X1 U10491 ( .A1(n9440), .A2(n22091), .Z(n30070) );
  XOR2_X1 U10493 ( .A1(n22031), .A2(n22243), .Z(n22091) );
  XOR2_X1 U10495 ( .A1(n24356), .A2(n24403), .Z(n17798) );
  NAND3_X2 U10502 ( .A1(n10176), .A2(n10179), .A3(n10175), .ZN(n24356) );
  NAND2_X2 U10504 ( .A1(n22737), .A2(n2449), .ZN(n22944) );
  OAI22_X2 U10505 ( .A1(n32369), .A2(n6654), .B1(n24073), .B2(n737), .ZN(n6651) );
  XOR2_X1 U10506 ( .A1(n23489), .A2(n23435), .Z(n30390) );
  OAI21_X2 U10509 ( .A1(n26526), .A2(n22710), .B(n8726), .ZN(n23435) );
  XOR2_X1 U10510 ( .A1(n18911), .A2(n19466), .Z(n10210) );
  NAND2_X2 U10514 ( .A1(n7420), .A2(n27553), .ZN(n18911) );
  OR2_X1 U10515 ( .A1(n10862), .A2(n17185), .Z(n12097) );
  XOR2_X1 U10517 ( .A1(n25993), .A2(n2388), .Z(n5861) );
  INV_X2 U10519 ( .I(n12934), .ZN(n23488) );
  NAND2_X2 U10520 ( .A1(n28401), .A2(n4305), .ZN(n12934) );
  NAND2_X1 U10521 ( .A1(n17134), .A2(n34165), .ZN(n15997) );
  NOR2_X1 U10535 ( .A1(n31033), .A2(n32929), .ZN(n30626) );
  NAND2_X1 U10537 ( .A1(n32373), .A2(n32372), .ZN(n9350) );
  INV_X1 U10538 ( .I(n32800), .ZN(n32374) );
  XOR2_X1 U10539 ( .A1(n30411), .A2(n19736), .Z(n19574) );
  OAI21_X2 U10540 ( .A1(n19142), .A2(n19141), .B(n16875), .ZN(n19736) );
  AOI22_X2 U10543 ( .A1(n28585), .A2(n33011), .B1(n23747), .B2(n16628), .ZN(
        n27168) );
  NAND2_X2 U10546 ( .A1(n11391), .A2(n11393), .ZN(n28585) );
  OAI21_X2 U10550 ( .A1(n20028), .A2(n1042), .B(n20025), .ZN(n8244) );
  INV_X2 U10553 ( .I(n14082), .ZN(n1042) );
  XOR2_X1 U10556 ( .A1(n7297), .A2(n7295), .Z(n14082) );
  NOR2_X2 U10558 ( .A1(n15358), .A2(n32375), .ZN(n11208) );
  OAI22_X2 U10562 ( .A1(n21114), .A2(n33741), .B1(n4989), .B2(n16072), .ZN(
        n32375) );
  NAND2_X2 U10563 ( .A1(n7974), .A2(n32376), .ZN(n25592) );
  NAND2_X1 U10564 ( .A1(n33095), .A2(n10248), .ZN(n32376) );
  INV_X2 U10565 ( .I(n19920), .ZN(n32377) );
  NAND2_X2 U10576 ( .A1(n32746), .A2(n14761), .ZN(n19920) );
  XOR2_X1 U10580 ( .A1(n32379), .A2(n26401), .Z(n13022) );
  XOR2_X1 U10585 ( .A1(n30058), .A2(n10915), .Z(n30057) );
  AOI22_X1 U10588 ( .A1(n15869), .A2(n19227), .B1(n18974), .B2(n19226), .ZN(
        n13939) );
  XOR2_X1 U10589 ( .A1(n20992), .A2(n1339), .Z(n20654) );
  XOR2_X1 U10592 ( .A1(n2953), .A2(n32380), .Z(n3392) );
  XOR2_X1 U10593 ( .A1(n3396), .A2(n3393), .Z(n32380) );
  XOR2_X1 U10595 ( .A1(n32381), .A2(n6175), .Z(n5962) );
  XOR2_X1 U10596 ( .A1(n21912), .A2(n297), .Z(n32381) );
  XOR2_X1 U10597 ( .A1(n28803), .A2(n20999), .Z(n17524) );
  XOR2_X1 U10600 ( .A1(n20839), .A2(n30543), .Z(n20999) );
  XOR2_X1 U10602 ( .A1(n23405), .A2(n1102), .Z(n23125) );
  NOR2_X2 U10603 ( .A1(n33585), .A2(n28338), .ZN(n25757) );
  NAND2_X1 U10604 ( .A1(n33610), .A2(n29597), .ZN(n22496) );
  XOR2_X1 U10605 ( .A1(n6502), .A2(n32382), .Z(n9796) );
  XOR2_X1 U10606 ( .A1(n23458), .A2(n11325), .Z(n32382) );
  AOI21_X2 U10611 ( .A1(n13860), .A2(n18687), .B(n32383), .ZN(n2593) );
  NOR3_X2 U10616 ( .A1(n18687), .A2(n18871), .A3(n29308), .ZN(n32383) );
  NAND2_X2 U10617 ( .A1(n14387), .A2(n18168), .ZN(n6593) );
  XOR2_X1 U10618 ( .A1(n23451), .A2(n23449), .Z(n9782) );
  XOR2_X1 U10621 ( .A1(n770), .A2(n31727), .Z(n23449) );
  NAND2_X2 U10622 ( .A1(n31759), .A2(n32656), .ZN(n33832) );
  XOR2_X1 U10625 ( .A1(n24788), .A2(n24746), .Z(n24024) );
  AOI22_X2 U10626 ( .A1(n28043), .A2(n28085), .B1(n26399), .B2(n31863), .ZN(
        n32385) );
  NAND2_X2 U10627 ( .A1(n8117), .A2(n8118), .ZN(n8130) );
  NAND2_X2 U10631 ( .A1(n5825), .A2(n31991), .ZN(n8117) );
  NAND2_X1 U10632 ( .A1(n23750), .A2(n12848), .ZN(n33165) );
  NOR2_X2 U10634 ( .A1(n29648), .A2(n23070), .ZN(n4803) );
  NOR3_X1 U10637 ( .A1(n31272), .A2(n16743), .A3(n32386), .ZN(n20879) );
  INV_X1 U10641 ( .I(n16938), .ZN(n32386) );
  OAI21_X2 U10644 ( .A1(n27535), .A2(n21778), .B(n276), .ZN(n12542) );
  XOR2_X1 U10647 ( .A1(n4741), .A2(n27000), .Z(n4740) );
  INV_X2 U10655 ( .I(n14545), .ZN(n1157) );
  NAND2_X2 U10656 ( .A1(n2674), .A2(n28285), .ZN(n14545) );
  XOR2_X1 U10657 ( .A1(n10320), .A2(n31828), .Z(n10708) );
  NAND2_X2 U10660 ( .A1(n32387), .A2(n23178), .ZN(n3147) );
  NAND2_X2 U10665 ( .A1(n31314), .A2(n30470), .ZN(n32387) );
  XOR2_X1 U10667 ( .A1(n31642), .A2(n30636), .Z(n30635) );
  INV_X2 U10669 ( .I(n14756), .ZN(n23902) );
  XOR2_X1 U10671 ( .A1(n15548), .A2(n27106), .Z(n4192) );
  XOR2_X1 U10674 ( .A1(n527), .A2(n9810), .Z(n31054) );
  XOR2_X1 U10675 ( .A1(n22030), .A2(n3550), .Z(n527) );
  XOR2_X1 U10676 ( .A1(n27052), .A2(n3126), .Z(n3169) );
  NOR2_X1 U10677 ( .A1(n1360), .A2(n17456), .ZN(n8294) );
  NAND3_X2 U10680 ( .A1(n32388), .A2(n11761), .A3(n11760), .ZN(n15877) );
  NAND2_X1 U10683 ( .A1(n30503), .A2(n7035), .ZN(n32388) );
  XOR2_X1 U10690 ( .A1(n1993), .A2(n17837), .Z(n20558) );
  NAND2_X2 U10697 ( .A1(n30450), .A2(n32418), .ZN(n1993) );
  AOI22_X2 U10698 ( .A1(n33522), .A2(n32389), .B1(n4803), .B2(n29070), .ZN(
        n4801) );
  NOR2_X2 U10701 ( .A1(n29070), .A2(n29648), .ZN(n32389) );
  NAND2_X2 U10702 ( .A1(n23987), .A2(n32390), .ZN(n33124) );
  NAND3_X2 U10711 ( .A1(n8), .A2(n13268), .A3(n8086), .ZN(n32390) );
  NAND2_X2 U10714 ( .A1(n25966), .A2(n819), .ZN(n10000) );
  NAND2_X1 U10716 ( .A1(n26806), .A2(n24335), .ZN(n29388) );
  XOR2_X1 U10717 ( .A1(n32391), .A2(n17440), .Z(n32919) );
  XOR2_X1 U10720 ( .A1(n27506), .A2(n32392), .Z(n32391) );
  AOI21_X2 U10721 ( .A1(n21206), .A2(n21289), .B(n32393), .ZN(n21207) );
  AOI22_X2 U10722 ( .A1(n20197), .A2(n20531), .B1(n13499), .B2(n27755), .ZN(
        n27646) );
  NOR2_X2 U10723 ( .A1(n1155), .A2(n32903), .ZN(n20197) );
  XOR2_X1 U10726 ( .A1(n31295), .A2(n21015), .Z(n2786) );
  XOR2_X1 U10727 ( .A1(n31704), .A2(n14918), .Z(n25110) );
  XOR2_X1 U10730 ( .A1(n1302), .A2(n17745), .Z(n9135) );
  XOR2_X1 U10732 ( .A1(n26863), .A2(n22013), .Z(n1302) );
  NOR2_X2 U10735 ( .A1(n11710), .A2(n28390), .ZN(n20550) );
  XOR2_X1 U10736 ( .A1(n17798), .A2(n24634), .Z(n16989) );
  XOR2_X1 U10739 ( .A1(n14499), .A2(n9943), .Z(n4222) );
  NAND2_X1 U10742 ( .A1(n32394), .A2(n16094), .ZN(n33991) );
  NAND2_X1 U10743 ( .A1(n28990), .A2(n33020), .ZN(n32394) );
  XOR2_X1 U10744 ( .A1(n32395), .A2(n527), .Z(n8154) );
  XOR2_X1 U10745 ( .A1(n13564), .A2(n33072), .Z(n32395) );
  OAI21_X1 U10746 ( .A1(n26471), .A2(n12872), .B(n33149), .ZN(n13000) );
  NAND2_X1 U10747 ( .A1(n13558), .A2(n7004), .ZN(n23105) );
  NAND3_X2 U10748 ( .A1(n14069), .A2(n22568), .A3(n22569), .ZN(n13558) );
  XOR2_X1 U10756 ( .A1(n32396), .A2(n24398), .Z(n16062) );
  XOR2_X1 U10758 ( .A1(n24395), .A2(n30607), .Z(n32396) );
  BUF_X2 U10759 ( .I(n10720), .Z(n32397) );
  OAI21_X2 U10761 ( .A1(n26198), .A2(n965), .B(n24947), .ZN(n32398) );
  AOI21_X2 U10766 ( .A1(n24161), .A2(n30595), .B(n3678), .ZN(n30307) );
  AND2_X1 U10768 ( .A1(n20584), .A2(n20583), .Z(n34045) );
  AOI22_X2 U10769 ( .A1(n17303), .A2(n17302), .B1(n14671), .B2(n22411), .ZN(
        n33299) );
  NOR2_X2 U10773 ( .A1(n26305), .A2(n7023), .ZN(n17303) );
  NAND3_X1 U10774 ( .A1(n16664), .A2(n12100), .A3(n20010), .ZN(n19782) );
  NOR2_X2 U10775 ( .A1(n1140), .A2(n5018), .ZN(n6219) );
  AOI22_X2 U10779 ( .A1(n27088), .A2(n17739), .B1(n23055), .B2(n2222), .ZN(
        n26900) );
  NAND2_X2 U10780 ( .A1(n32400), .A2(n18782), .ZN(n15166) );
  NAND2_X2 U10782 ( .A1(n18187), .A2(n30686), .ZN(n32400) );
  XOR2_X1 U10784 ( .A1(n33291), .A2(n27942), .Z(n4330) );
  XOR2_X1 U10786 ( .A1(n23371), .A2(n11504), .Z(n23473) );
  AOI22_X2 U10787 ( .A1(n3692), .A2(n32964), .B1(n3689), .B2(n13597), .ZN(
        n23371) );
  NOR2_X2 U10788 ( .A1(n12759), .A2(n12757), .ZN(n16641) );
  NOR2_X2 U10789 ( .A1(n30873), .A2(n32043), .ZN(n12759) );
  XOR2_X1 U10791 ( .A1(n16030), .A2(n33939), .Z(n13180) );
  XNOR2_X1 U10793 ( .A1(n14507), .A2(n8855), .ZN(n32502) );
  AOI22_X2 U10796 ( .A1(n21372), .A2(n21377), .B1(n33774), .B2(n32907), .ZN(
        n21573) );
  NOR2_X2 U10797 ( .A1(n21213), .A2(n12525), .ZN(n21372) );
  INV_X1 U10802 ( .I(n24787), .ZN(n26795) );
  NAND2_X2 U10803 ( .A1(n6741), .A2(n33489), .ZN(n24787) );
  NAND2_X2 U10805 ( .A1(n29256), .A2(n21079), .ZN(n13712) );
  NAND2_X2 U10807 ( .A1(n10361), .A2(n23086), .ZN(n33791) );
  XOR2_X1 U10809 ( .A1(n32402), .A2(n19766), .Z(n5856) );
  XOR2_X1 U10810 ( .A1(n32587), .A2(n13480), .Z(n32402) );
  XOR2_X1 U10812 ( .A1(n32403), .A2(n20823), .Z(n16770) );
  XOR2_X1 U10815 ( .A1(n16773), .A2(n17759), .Z(n32403) );
  BUF_X4 U10816 ( .I(n9172), .Z(n4319) );
  BUF_X2 U10818 ( .I(n33437), .Z(n32404) );
  NAND2_X2 U10820 ( .A1(n33784), .A2(n4206), .ZN(n5121) );
  OAI22_X1 U10822 ( .A1(n576), .A2(n5966), .B1(n29153), .B2(n4373), .ZN(n19924) );
  NOR2_X2 U10824 ( .A1(n32405), .A2(n30294), .ZN(n5317) );
  NOR3_X1 U10825 ( .A1(n17537), .A2(n16337), .A3(n23351), .ZN(n32405) );
  NAND2_X2 U10826 ( .A1(n32407), .A2(n12018), .ZN(n15863) );
  NAND3_X2 U10834 ( .A1(n16637), .A2(n27938), .A3(n8292), .ZN(n32528) );
  OR2_X2 U10839 ( .A1(n9920), .A2(n9490), .Z(n23933) );
  XOR2_X1 U10840 ( .A1(n20788), .A2(n21029), .Z(n20983) );
  NAND2_X2 U10841 ( .A1(n31269), .A2(n20612), .ZN(n20788) );
  NOR2_X1 U10845 ( .A1(n32410), .A2(n18687), .ZN(n32409) );
  INV_X2 U10846 ( .I(n18871), .ZN(n32411) );
  NOR2_X2 U10854 ( .A1(n5616), .A2(n5613), .ZN(n31893) );
  XOR2_X1 U10857 ( .A1(n12170), .A2(n12172), .Z(n20946) );
  XOR2_X1 U10862 ( .A1(n23137), .A2(n32975), .Z(n23168) );
  NOR2_X2 U10865 ( .A1(n32741), .A2(n29510), .ZN(n30824) );
  XOR2_X1 U10867 ( .A1(n32412), .A2(n22246), .Z(n26484) );
  XOR2_X1 U10871 ( .A1(n8475), .A2(n13651), .Z(n32412) );
  OAI21_X2 U10872 ( .A1(n7228), .A2(n31522), .B(n33820), .ZN(n33819) );
  AOI21_X1 U10873 ( .A1(n33530), .A2(n33225), .B(n33222), .ZN(n33224) );
  AOI21_X2 U10874 ( .A1(n24294), .A2(n24295), .B(n29352), .ZN(n32789) );
  XOR2_X1 U10876 ( .A1(n32413), .A2(n30514), .Z(n11877) );
  XOR2_X1 U10877 ( .A1(n28584), .A2(n20897), .Z(n32413) );
  BUF_X2 U10883 ( .I(n27021), .Z(n32414) );
  XOR2_X1 U10885 ( .A1(n13415), .A2(n23285), .Z(n31288) );
  NAND3_X2 U10886 ( .A1(n9791), .A2(n27544), .A3(n22441), .ZN(n23285) );
  NAND4_X1 U10890 ( .A1(n19235), .A2(n8119), .A3(n8118), .A4(n8117), .ZN(
        n19894) );
  OAI21_X2 U10897 ( .A1(n161), .A2(n27345), .B(n3310), .ZN(n19235) );
  XOR2_X1 U10898 ( .A1(n32415), .A2(n7257), .Z(n9126) );
  XOR2_X1 U10899 ( .A1(n24540), .A2(n17448), .Z(n32415) );
  XOR2_X1 U10901 ( .A1(n14337), .A2(n6974), .Z(n12972) );
  NAND2_X1 U10903 ( .A1(n19835), .A2(n32371), .ZN(n32416) );
  XOR2_X1 U10906 ( .A1(n32417), .A2(n1084), .Z(n10632) );
  NAND2_X1 U10914 ( .A1(n3558), .A2(n20404), .ZN(n32418) );
  OAI21_X2 U10918 ( .A1(n26078), .A2(n6581), .B(n32419), .ZN(n4956) );
  NAND3_X1 U10919 ( .A1(n14770), .A2(n6555), .A3(n7188), .ZN(n32419) );
  XOR2_X1 U10920 ( .A1(n32420), .A2(n27200), .Z(n27453) );
  XOR2_X1 U10922 ( .A1(n30706), .A2(n27778), .Z(n32420) );
  OR2_X1 U10927 ( .A1(n8965), .A2(n17140), .Z(n16412) );
  XOR2_X1 U10933 ( .A1(n9634), .A2(n9635), .Z(n10433) );
  NAND3_X1 U10936 ( .A1(n25045), .A2(n31640), .A3(n27610), .ZN(n25046) );
  NAND2_X1 U10937 ( .A1(n32422), .A2(n32421), .ZN(n24875) );
  NAND2_X1 U10939 ( .A1(n25015), .A2(n25012), .ZN(n32421) );
  NAND2_X1 U10941 ( .A1(n17240), .A2(n24975), .ZN(n32422) );
  OR2_X2 U10942 ( .A1(n23742), .A2(n15116), .Z(n27459) );
  AND2_X1 U10950 ( .A1(n21438), .A2(n8398), .Z(n30646) );
  XOR2_X1 U10954 ( .A1(n24691), .A2(n25064), .Z(n15792) );
  NOR2_X2 U10959 ( .A1(n7018), .A2(n14411), .ZN(n14410) );
  XOR2_X1 U10960 ( .A1(n91), .A2(n1416), .Z(n9308) );
  NAND2_X2 U10962 ( .A1(n31643), .A2(n29520), .ZN(n91) );
  AOI21_X2 U10966 ( .A1(n32423), .A2(n31483), .B(n29773), .ZN(n10710) );
  NOR2_X2 U10969 ( .A1(n23809), .A2(n14664), .ZN(n32423) );
  OR2_X1 U10972 ( .A1(n2643), .A2(n26782), .Z(n21470) );
  AOI22_X2 U10977 ( .A1(n32424), .A2(n33591), .B1(n2169), .B2(n17739), .ZN(
        n4847) );
  NAND3_X2 U10979 ( .A1(n32425), .A2(n27459), .A3(n23769), .ZN(n8286) );
  NOR3_X2 U10980 ( .A1(n4714), .A2(n32802), .A3(n1049), .ZN(n29768) );
  OAI22_X2 U10983 ( .A1(n23901), .A2(n5373), .B1(n1254), .B2(n667), .ZN(n32426) );
  AOI21_X2 U10985 ( .A1(n24888), .A2(n25149), .B(n16293), .ZN(n32427) );
  XOR2_X1 U10986 ( .A1(n2812), .A2(n32428), .Z(n13670) );
  XOR2_X1 U10987 ( .A1(n16178), .A2(n20974), .Z(n32428) );
  XOR2_X1 U10993 ( .A1(n19686), .A2(n19773), .Z(n9327) );
  NAND2_X2 U10995 ( .A1(n30426), .A2(n5329), .ZN(n19686) );
  NOR3_X1 U10996 ( .A1(n31216), .A2(n28270), .A3(n24857), .ZN(n33084) );
  INV_X2 U10999 ( .I(n32429), .ZN(n871) );
  XOR2_X1 U11001 ( .A1(n10722), .A2(n10723), .Z(n32429) );
  NAND2_X2 U11007 ( .A1(n32430), .A2(n23060), .ZN(n17775) );
  NAND2_X2 U11009 ( .A1(n32431), .A2(n33088), .ZN(n2073) );
  NAND2_X2 U11011 ( .A1(n26758), .A2(n32432), .ZN(n7287) );
  NAND2_X2 U11017 ( .A1(n2383), .A2(n22463), .ZN(n32432) );
  NAND2_X2 U11020 ( .A1(n23919), .A2(n6869), .ZN(n5759) );
  XOR2_X1 U11023 ( .A1(n9474), .A2(n10872), .Z(n14845) );
  NAND2_X2 U11025 ( .A1(n24148), .A2(n24147), .ZN(n11346) );
  NAND2_X2 U11028 ( .A1(n10500), .A2(n23574), .ZN(n24148) );
  XOR2_X1 U11032 ( .A1(n16283), .A2(n32433), .Z(n23719) );
  XOR2_X1 U11039 ( .A1(n23450), .A2(n23062), .Z(n32433) );
  XOR2_X1 U11041 ( .A1(n17504), .A2(n17505), .Z(n18075) );
  AND2_X1 U11042 ( .A1(n5466), .A2(n11571), .Z(n14510) );
  OAI22_X1 U11044 ( .A1(n21412), .A2(n14483), .B1(n13367), .B2(n11513), .ZN(
        n10135) );
  XOR2_X1 U11045 ( .A1(n20895), .A2(n14875), .Z(n3630) );
  OR2_X1 U11046 ( .A1(n21085), .A2(n14803), .Z(n26988) );
  NAND2_X2 U11048 ( .A1(n29754), .A2(n34069), .ZN(n14359) );
  NAND2_X2 U11052 ( .A1(n33379), .A2(n10003), .ZN(n22798) );
  OAI21_X2 U11056 ( .A1(n1047), .A2(n18988), .B(n5761), .ZN(n10373) );
  NAND2_X1 U11058 ( .A1(n30643), .A2(n5748), .ZN(n20537) );
  NOR2_X2 U11063 ( .A1(n30031), .A2(n9341), .ZN(n30643) );
  INV_X2 U11066 ( .I(n32436), .ZN(n24216) );
  NAND3_X2 U11073 ( .A1(n33431), .A2(n33457), .A3(n14166), .ZN(n32436) );
  BUF_X2 U11074 ( .I(n27921), .Z(n32437) );
  NAND2_X2 U11077 ( .A1(n10046), .A2(n23964), .ZN(n24676) );
  AOI22_X2 U11078 ( .A1(n29293), .A2(n31113), .B1(n10047), .B2(n10859), .ZN(
        n10046) );
  AOI22_X2 U11079 ( .A1(n8968), .A2(n24290), .B1(n32985), .B2(n2444), .ZN(
        n12454) );
  NAND2_X1 U11080 ( .A1(n12135), .A2(n17501), .ZN(n32438) );
  NAND2_X2 U11082 ( .A1(n25852), .A2(n25851), .ZN(n30805) );
  NOR2_X2 U11083 ( .A1(n10897), .A2(n16673), .ZN(n25852) );
  NAND2_X2 U11088 ( .A1(n32439), .A2(n33396), .ZN(n19180) );
  NAND2_X2 U11094 ( .A1(n11208), .A2(n21797), .ZN(n28824) );
  NOR2_X1 U11095 ( .A1(n33788), .A2(n31916), .ZN(n13354) );
  NOR2_X2 U11096 ( .A1(n14948), .A2(n29721), .ZN(n14952) );
  NOR2_X2 U11098 ( .A1(n32917), .A2(n12356), .ZN(n24015) );
  NAND2_X2 U11100 ( .A1(n21314), .A2(n28565), .ZN(n17698) );
  NOR2_X2 U11101 ( .A1(n32440), .A2(n29560), .ZN(n1344) );
  BUF_X4 U11102 ( .I(n14457), .Z(n34103) );
  OAI21_X2 U11105 ( .A1(n32437), .A2(n19111), .B(n28996), .ZN(n19629) );
  NOR3_X2 U11106 ( .A1(n10965), .A2(n18260), .A3(n18370), .ZN(n19360) );
  NAND2_X2 U11107 ( .A1(n33285), .A2(n1609), .ZN(n10087) );
  NAND2_X2 U11110 ( .A1(n9770), .A2(n32442), .ZN(n14123) );
  XOR2_X1 U11113 ( .A1(n32443), .A2(n31513), .Z(Ciphertext[8]) );
  XOR2_X1 U11115 ( .A1(n32445), .A2(n14899), .Z(n13716) );
  XOR2_X1 U11125 ( .A1(n21048), .A2(n5024), .Z(n32445) );
  NOR2_X2 U11127 ( .A1(n32447), .A2(n32446), .ZN(n16051) );
  INV_X2 U11128 ( .I(n22429), .ZN(n32448) );
  BUF_X2 U11129 ( .I(n22521), .Z(n32449) );
  NAND3_X2 U11132 ( .A1(n30071), .A2(n15544), .A3(n30805), .ZN(n32782) );
  AOI21_X2 U11135 ( .A1(n32450), .A2(n26173), .B(n31001), .ZN(n21929) );
  BUF_X2 U11136 ( .I(n14625), .Z(n32451) );
  OAI21_X2 U11138 ( .A1(n6320), .A2(n6321), .B(n28914), .ZN(n32453) );
  AOI21_X2 U11141 ( .A1(n27625), .A2(n5050), .B(n32911), .ZN(n32910) );
  NAND2_X2 U11143 ( .A1(n18154), .A2(n25019), .ZN(n5050) );
  XOR2_X1 U11144 ( .A1(n19558), .A2(n3131), .Z(n17840) );
  XOR2_X1 U11145 ( .A1(n32458), .A2(n25878), .Z(Ciphertext[180]) );
  NAND2_X1 U11147 ( .A1(n6047), .A2(n31075), .ZN(n32458) );
  XOR2_X1 U11148 ( .A1(n13471), .A2(n24621), .Z(n9467) );
  XOR2_X1 U11150 ( .A1(n11751), .A2(n3345), .Z(n24621) );
  NAND3_X1 U11151 ( .A1(n1081), .A2(n13428), .A3(n14454), .ZN(n7532) );
  NAND3_X1 U11153 ( .A1(n10862), .A2(n27390), .A3(n8919), .ZN(n17186) );
  XOR2_X1 U11154 ( .A1(n22313), .A2(n12980), .Z(n21885) );
  AOI21_X1 U11157 ( .A1(n10653), .A2(n24156), .B(n10652), .ZN(n6741) );
  NOR2_X2 U11162 ( .A1(n12043), .A2(n16240), .ZN(n15327) );
  AOI21_X2 U11165 ( .A1(n5160), .A2(n24093), .B(n888), .ZN(n5161) );
  NOR2_X1 U11179 ( .A1(n16408), .A2(n17601), .ZN(n33047) );
  AOI21_X2 U11182 ( .A1(n9105), .A2(n19814), .B(n32460), .ZN(n31533) );
  NOR2_X1 U11184 ( .A1(n19811), .A2(n19812), .ZN(n32460) );
  XOR2_X1 U11190 ( .A1(n11751), .A2(n16575), .Z(n5378) );
  NAND3_X2 U11191 ( .A1(n27397), .A2(n27396), .A3(n5307), .ZN(n11751) );
  XNOR2_X1 U11194 ( .A1(n20852), .A2(n20851), .ZN(n20930) );
  AOI22_X2 U11196 ( .A1(n10379), .A2(n20499), .B1(n10992), .B2(n20497), .ZN(
        n20851) );
  NOR2_X2 U11200 ( .A1(n11241), .A2(n12991), .ZN(n20852) );
  NAND2_X2 U11204 ( .A1(n29790), .A2(n28035), .ZN(n1577) );
  INV_X4 U11209 ( .I(n32461), .ZN(n20635) );
  AND3_X2 U11212 ( .A1(n1812), .A2(n1813), .A3(n1814), .Z(n32461) );
  NAND4_X2 U11214 ( .A1(n17480), .A2(n17479), .A3(n24353), .A4(n33343), .ZN(
        n32709) );
  NAND2_X2 U11215 ( .A1(n32462), .A2(n12237), .ZN(n13334) );
  NAND2_X2 U11216 ( .A1(n32463), .A2(n18142), .ZN(n30090) );
  OAI22_X2 U11219 ( .A1(n1362), .A2(n11911), .B1(n1458), .B2(n397), .ZN(n32463) );
  XOR2_X1 U11223 ( .A1(n31221), .A2(n22104), .Z(n29740) );
  NAND2_X2 U11228 ( .A1(n17124), .A2(n17122), .ZN(n22791) );
  NOR2_X1 U11229 ( .A1(n26013), .A2(n32778), .ZN(n29547) );
  XOR2_X1 U11234 ( .A1(n13395), .A2(n10628), .Z(n32464) );
  XOR2_X1 U11237 ( .A1(n19578), .A2(n19556), .Z(n5768) );
  BUF_X2 U11239 ( .I(n3148), .Z(n32465) );
  NOR2_X1 U11241 ( .A1(n21806), .A2(n21805), .ZN(n33985) );
  NAND2_X2 U11243 ( .A1(n1837), .A2(n1838), .ZN(n8636) );
  NAND2_X2 U11246 ( .A1(n32546), .A2(n337), .ZN(n16708) );
  NAND3_X2 U11247 ( .A1(n32466), .A2(n9232), .A3(n330), .ZN(n33140) );
  NAND2_X2 U11249 ( .A1(n15394), .A2(n26130), .ZN(n32466) );
  XOR2_X1 U11254 ( .A1(n16448), .A2(n20990), .Z(n34038) );
  NOR2_X2 U11256 ( .A1(n5059), .A2(n5061), .ZN(n16448) );
  NOR2_X2 U11258 ( .A1(n31220), .A2(n29084), .ZN(n27535) );
  NAND2_X2 U11259 ( .A1(n1508), .A2(n32468), .ZN(n24810) );
  AOI22_X2 U11261 ( .A1(n32049), .A2(n24251), .B1(n1511), .B2(n1513), .ZN(
        n32468) );
  OAI21_X1 U11264 ( .A1(n787), .A2(n5713), .B(n25106), .ZN(n18175) );
  INV_X2 U11265 ( .I(n11360), .ZN(n787) );
  NAND2_X2 U11266 ( .A1(n3223), .A2(n3225), .ZN(n11360) );
  OAI21_X2 U11269 ( .A1(n10645), .A2(n10646), .B(n7181), .ZN(n10329) );
  NAND3_X1 U11271 ( .A1(n8030), .A2(n16925), .A3(n16157), .ZN(n7324) );
  OR2_X1 U11277 ( .A1(n17637), .A2(n6595), .Z(n30523) );
  INV_X2 U11278 ( .I(n1026), .ZN(n33631) );
  NOR2_X2 U11286 ( .A1(n11187), .A2(n1145), .ZN(n11091) );
  INV_X2 U11287 ( .I(n10433), .ZN(n1145) );
  AND2_X1 U11289 ( .A1(n21604), .A2(n26439), .Z(n34028) );
  XOR2_X1 U11290 ( .A1(n31493), .A2(n22075), .Z(n16150) );
  XOR2_X1 U11291 ( .A1(n22105), .A2(n27633), .Z(n31649) );
  XOR2_X1 U11292 ( .A1(n17362), .A2(n22012), .Z(n22105) );
  XOR2_X1 U11297 ( .A1(n6771), .A2(n28762), .Z(n33203) );
  OAI21_X2 U11304 ( .A1(n34026), .A2(n21656), .B(n32535), .ZN(n28762) );
  XOR2_X1 U11309 ( .A1(n24618), .A2(n24393), .Z(n24504) );
  NOR2_X2 U11314 ( .A1(n28505), .A2(n12262), .ZN(n24618) );
  OAI22_X2 U11315 ( .A1(n28367), .A2(n10213), .B1(n23873), .B2(n17133), .ZN(
        n3571) );
  INV_X1 U11318 ( .I(n33996), .ZN(n22741) );
  NAND2_X1 U11320 ( .A1(n22848), .A2(n31854), .ZN(n33996) );
  XOR2_X1 U11321 ( .A1(n30029), .A2(n32469), .Z(n24565) );
  XOR2_X1 U11323 ( .A1(n9011), .A2(n9012), .Z(n9010) );
  NOR2_X2 U11324 ( .A1(n5741), .A2(n29306), .ZN(n6769) );
  INV_X1 U11325 ( .I(n18100), .ZN(n14593) );
  XNOR2_X1 U11326 ( .A1(n22137), .A2(n22158), .ZN(n18100) );
  XOR2_X1 U11330 ( .A1(n19565), .A2(n14146), .Z(n19429) );
  OR2_X2 U11331 ( .A1(n499), .A2(n33461), .Z(n17579) );
  NOR2_X2 U11332 ( .A1(n22563), .A2(n14034), .ZN(n32654) );
  NAND2_X2 U11333 ( .A1(n16447), .A2(n15089), .ZN(n22563) );
  XOR2_X1 U11334 ( .A1(n30380), .A2(n23488), .Z(n28587) );
  NOR2_X1 U11336 ( .A1(n15234), .A2(n3080), .ZN(n32471) );
  INV_X2 U11338 ( .I(n25444), .ZN(n25455) );
  NAND2_X2 U11339 ( .A1(n33245), .A2(n33258), .ZN(n25444) );
  NOR2_X2 U11345 ( .A1(n32472), .A2(n9725), .ZN(n32648) );
  AOI21_X2 U11351 ( .A1(n19826), .A2(n19827), .B(n29972), .ZN(n32472) );
  INV_X4 U11353 ( .I(n32635), .ZN(n11956) );
  INV_X2 U11354 ( .I(n18039), .ZN(n20097) );
  XOR2_X1 U11355 ( .A1(n17954), .A2(n17953), .Z(n18039) );
  AOI22_X2 U11357 ( .A1(n5080), .A2(n29985), .B1(n5079), .B2(n1232), .ZN(
        n30327) );
  AND3_X1 U11359 ( .A1(n11298), .A2(n14420), .A3(n4184), .Z(n33834) );
  NAND2_X2 U11361 ( .A1(n11823), .A2(n11824), .ZN(n30047) );
  XOR2_X1 U11362 ( .A1(n20716), .A2(n32473), .Z(n7918) );
  XOR2_X1 U11366 ( .A1(n7594), .A2(n20552), .Z(n32473) );
  XOR2_X1 U11369 ( .A1(n26920), .A2(n28134), .Z(n16275) );
  XOR2_X1 U11376 ( .A1(n61), .A2(n32474), .Z(n25963) );
  XOR2_X1 U11383 ( .A1(n21985), .A2(n15950), .Z(n32474) );
  XOR2_X1 U11385 ( .A1(n4583), .A2(n29458), .Z(n4581) );
  XOR2_X1 U11390 ( .A1(n5090), .A2(n24116), .Z(n24793) );
  NOR2_X2 U11393 ( .A1(n10531), .A2(n12002), .ZN(n5090) );
  XOR2_X1 U11403 ( .A1(n10235), .A2(n24685), .Z(n27290) );
  XOR2_X1 U11417 ( .A1(n24750), .A2(n5090), .Z(n24685) );
  INV_X2 U11422 ( .I(n14585), .ZN(n16615) );
  XOR2_X1 U11425 ( .A1(n14580), .A2(n14581), .Z(n14585) );
  NAND4_X2 U11431 ( .A1(n32475), .A2(n22857), .A3(n22859), .A4(n22860), .ZN(
        n23336) );
  NAND2_X2 U11434 ( .A1(n7797), .A2(n26667), .ZN(n32475) );
  AND2_X1 U11439 ( .A1(n20097), .A2(n20096), .Z(n7997) );
  AND2_X1 U11441 ( .A1(n25797), .A2(n16112), .Z(n14615) );
  NAND2_X2 U11443 ( .A1(n32476), .A2(n23479), .ZN(n29885) );
  OAI21_X2 U11444 ( .A1(n30825), .A2(n8415), .B(n33016), .ZN(n32476) );
  NOR2_X1 U11446 ( .A1(n28200), .A2(n15323), .ZN(n25129) );
  NAND3_X2 U11448 ( .A1(n14628), .A2(n14631), .A3(n14632), .ZN(n15323) );
  BUF_X2 U11453 ( .I(n13092), .Z(n32478) );
  NOR2_X2 U11461 ( .A1(n30832), .A2(n7811), .ZN(n5385) );
  OAI22_X2 U11468 ( .A1(n21196), .A2(n21195), .B1(n26542), .B2(n17624), .ZN(
        n30832) );
  OAI21_X2 U11473 ( .A1(n32479), .A2(n4855), .B(n33148), .ZN(n14106) );
  NAND2_X2 U11474 ( .A1(n2937), .A2(n8308), .ZN(n23511) );
  NAND2_X2 U11475 ( .A1(n33656), .A2(n2912), .ZN(n2937) );
  NAND2_X2 U11477 ( .A1(n11179), .A2(n19008), .ZN(n11219) );
  NAND2_X2 U11480 ( .A1(n32534), .A2(n27368), .ZN(n3007) );
  XOR2_X1 U11487 ( .A1(n32480), .A2(n23295), .Z(n81) );
  NAND2_X2 U11491 ( .A1(n33184), .A2(n2539), .ZN(n27396) );
  NAND3_X2 U11493 ( .A1(n983), .A2(n12259), .A3(n11268), .ZN(n11109) );
  XOR2_X1 U11496 ( .A1(n22169), .A2(n22168), .Z(n2162) );
  XOR2_X1 U11497 ( .A1(n1309), .A2(n16242), .Z(n22169) );
  INV_X2 U11498 ( .I(n4013), .ZN(n22132) );
  NAND2_X2 U11499 ( .A1(n3314), .A2(n3316), .ZN(n4013) );
  NAND2_X1 U11500 ( .A1(n33937), .A2(n28085), .ZN(n12808) );
  XOR2_X1 U11505 ( .A1(n7545), .A2(n22271), .Z(n22104) );
  NOR2_X2 U11508 ( .A1(n17418), .A2(n21347), .ZN(n22271) );
  NAND2_X2 U11510 ( .A1(n26375), .A2(n32482), .ZN(n17855) );
  NAND2_X1 U11514 ( .A1(n23708), .A2(n12680), .ZN(n15942) );
  AOI22_X2 U11515 ( .A1(n28428), .A2(n24134), .B1(n24135), .B2(n27739), .ZN(
        n27998) );
  XOR2_X1 U11526 ( .A1(n20918), .A2(n20834), .Z(n4949) );
  XOR2_X1 U11527 ( .A1(n20960), .A2(n1339), .Z(n20918) );
  AOI21_X2 U11528 ( .A1(n27150), .A2(n24925), .B(n24920), .ZN(n4867) );
  INV_X2 U11529 ( .I(n24936), .ZN(n24920) );
  NAND2_X2 U11531 ( .A1(n16216), .A2(n16217), .ZN(n13573) );
  INV_X2 U11532 ( .I(n6531), .ZN(n12263) );
  AOI22_X2 U11533 ( .A1(n19924), .A2(n26615), .B1(n8934), .B2(n33187), .ZN(
        n6531) );
  INV_X2 U11545 ( .I(n14737), .ZN(n963) );
  NOR2_X1 U11546 ( .A1(n8535), .A2(n10993), .ZN(n32494) );
  AND2_X1 U11548 ( .A1(n29203), .A2(n23578), .Z(n12326) );
  NOR2_X2 U11549 ( .A1(n13966), .A2(n13965), .ZN(n27066) );
  INV_X2 U11551 ( .I(n32484), .ZN(n29250) );
  XNOR2_X1 U11555 ( .A1(n4014), .A2(n4895), .ZN(n32484) );
  NAND3_X1 U11558 ( .A1(n26830), .A2(n13295), .A3(n13390), .ZN(n12114) );
  NOR2_X2 U11559 ( .A1(n9377), .A2(n23018), .ZN(n22473) );
  NAND2_X1 U11567 ( .A1(n28), .A2(n9793), .ZN(n9792) );
  NAND2_X2 U11572 ( .A1(n32978), .A2(n15925), .ZN(n9793) );
  NAND2_X1 U11577 ( .A1(n1207), .A2(n25277), .ZN(n27873) );
  NAND2_X2 U11579 ( .A1(n22277), .A2(n7), .ZN(n11033) );
  OAI22_X2 U11582 ( .A1(n22411), .A2(n7023), .B1(n645), .B2(n16225), .ZN(
        n22277) );
  INV_X2 U11584 ( .I(n32486), .ZN(n31448) );
  XNOR2_X1 U11587 ( .A1(n2952), .A2(n2951), .ZN(n32486) );
  NAND2_X2 U11588 ( .A1(n32528), .A2(n20134), .ZN(n31157) );
  INV_X2 U11590 ( .I(n32487), .ZN(n8028) );
  XNOR2_X1 U11591 ( .A1(n8026), .A2(n27091), .ZN(n32487) );
  AOI22_X2 U11600 ( .A1(n97), .A2(n98), .B1(n29708), .B2(n32488), .ZN(n18146)
         );
  NAND2_X2 U11604 ( .A1(n23823), .A2(n23672), .ZN(n32488) );
  XOR2_X1 U11606 ( .A1(n12539), .A2(n14875), .Z(n15353) );
  XOR2_X1 U11607 ( .A1(n32489), .A2(n647), .Z(n2200) );
  NAND2_X2 U11608 ( .A1(n32490), .A2(n29107), .ZN(n4542) );
  OAI22_X2 U11610 ( .A1(n23055), .A2(n17739), .B1(n22878), .B2(n31437), .ZN(
        n32490) );
  NAND2_X1 U11619 ( .A1(n29692), .A2(n10623), .ZN(n10369) );
  NOR2_X2 U11621 ( .A1(n32491), .A2(n12768), .ZN(n31746) );
  OAI21_X2 U11623 ( .A1(n12150), .A2(n20412), .B(n12149), .ZN(n30219) );
  XOR2_X1 U11624 ( .A1(n22285), .A2(n32492), .Z(n13382) );
  XOR2_X1 U11627 ( .A1(n2824), .A2(n5099), .Z(n32492) );
  AOI22_X2 U11631 ( .A1(n20308), .A2(n3462), .B1(n2145), .B2(n33691), .ZN(
        n20309) );
  BUF_X2 U11633 ( .I(n907), .Z(n32493) );
  XOR2_X1 U11635 ( .A1(n33160), .A2(n30495), .Z(n10482) );
  NOR2_X2 U11636 ( .A1(n33409), .A2(n13804), .ZN(n30495) );
  INV_X2 U11639 ( .I(n15064), .ZN(n19634) );
  OAI21_X2 U11647 ( .A1(n2411), .A2(n2412), .B(n2410), .ZN(n15064) );
  NAND2_X2 U11648 ( .A1(n19220), .A2(n5610), .ZN(n14760) );
  NAND2_X2 U11650 ( .A1(n18371), .A2(n18372), .ZN(n19220) );
  XOR2_X1 U11652 ( .A1(n4246), .A2(n5732), .Z(n9351) );
  XOR2_X1 U11654 ( .A1(n15161), .A2(n2117), .Z(n24674) );
  AOI21_X2 U11655 ( .A1(n24066), .A2(n14745), .B(n3918), .ZN(n15161) );
  XOR2_X1 U11656 ( .A1(n8328), .A2(n10888), .Z(n11620) );
  INV_X2 U11658 ( .I(n8306), .ZN(n30528) );
  NAND2_X2 U11659 ( .A1(n10510), .A2(n10511), .ZN(n8306) );
  AOI22_X2 U11660 ( .A1(n12987), .A2(n20059), .B1(n20058), .B2(n941), .ZN(
        n12986) );
  XOR2_X1 U11665 ( .A1(n11358), .A2(n11355), .Z(n16885) );
  NOR3_X2 U11666 ( .A1(n33911), .A2(n33919), .A3(n25295), .ZN(n11258) );
  NAND2_X2 U11667 ( .A1(n13197), .A2(n7957), .ZN(n22921) );
  NAND2_X2 U11669 ( .A1(n12869), .A2(n17853), .ZN(n13197) );
  NAND3_X2 U11670 ( .A1(n11584), .A2(n32495), .A3(n21667), .ZN(n22125) );
  OAI21_X2 U11671 ( .A1(n26175), .A2(n4842), .B(n28618), .ZN(n32495) );
  BUF_X2 U11679 ( .I(n15172), .Z(n13133) );
  NOR2_X1 U11682 ( .A1(n34012), .A2(n34011), .ZN(n3336) );
  NAND3_X2 U11683 ( .A1(n810), .A2(n21080), .A3(n21365), .ZN(n33551) );
  OAI22_X2 U11685 ( .A1(n32496), .A2(n30510), .B1(n6482), .B2(n7090), .ZN(
        n22974) );
  AOI21_X2 U11686 ( .A1(n32498), .A2(n32497), .B(n29595), .ZN(n3634) );
  NOR2_X2 U11688 ( .A1(n32588), .A2(n32499), .ZN(n32498) );
  XOR2_X1 U11691 ( .A1(n22085), .A2(n22173), .Z(n17207) );
  XOR2_X1 U11696 ( .A1(n32501), .A2(n29420), .Z(n4820) );
  XOR2_X1 U11699 ( .A1(n1865), .A2(n26646), .Z(n32501) );
  NAND2_X2 U11701 ( .A1(n789), .A2(n29331), .ZN(n5839) );
  XOR2_X1 U11702 ( .A1(n16617), .A2(n16618), .Z(n8452) );
  XOR2_X1 U11703 ( .A1(n2969), .A2(n2968), .Z(n3012) );
  NOR2_X2 U11705 ( .A1(n17590), .A2(n17305), .ZN(n21162) );
  XOR2_X1 U11706 ( .A1(n20786), .A2(n20960), .Z(n20688) );
  NOR2_X2 U11710 ( .A1(n14394), .A2(n8264), .ZN(n20786) );
  XOR2_X1 U11716 ( .A1(n32502), .A2(n3793), .Z(n33538) );
  XOR2_X1 U11719 ( .A1(n5356), .A2(n32077), .Z(n33934) );
  NAND2_X1 U11726 ( .A1(n32503), .A2(n14433), .ZN(n33873) );
  NAND2_X1 U11729 ( .A1(n27659), .A2(n14432), .ZN(n32503) );
  INV_X2 U11734 ( .I(n32507), .ZN(n24603) );
  XOR2_X1 U11736 ( .A1(n5790), .A2(n24652), .Z(n32507) );
  OAI21_X2 U11750 ( .A1(n2640), .A2(n737), .B(n7891), .ZN(n33019) );
  XOR2_X1 U11751 ( .A1(n32508), .A2(n12754), .Z(Ciphertext[155]) );
  NAND2_X2 U11757 ( .A1(n28526), .A2(n16934), .ZN(n28203) );
  NAND2_X2 U11759 ( .A1(n3163), .A2(n724), .ZN(n28831) );
  AOI21_X2 U11760 ( .A1(n26688), .A2(n32509), .B(n8876), .ZN(n31434) );
  XOR2_X1 U11761 ( .A1(n20895), .A2(n10581), .Z(n32511) );
  NAND3_X1 U11764 ( .A1(n30945), .A2(n30946), .A3(n23082), .ZN(n33777) );
  BUF_X2 U11766 ( .I(n32605), .Z(n32512) );
  NAND3_X2 U11771 ( .A1(n11814), .A2(n21358), .A3(n21357), .ZN(n33297) );
  NAND2_X2 U11772 ( .A1(n32514), .A2(n30084), .ZN(n2045) );
  AOI22_X2 U11773 ( .A1(n1634), .A2(n24233), .B1(n5066), .B2(n974), .ZN(n32514) );
  XOR2_X1 U11775 ( .A1(n32517), .A2(n25358), .Z(Ciphertext[98]) );
  NAND2_X1 U11776 ( .A1(n28469), .A2(n28470), .ZN(n32517) );
  OR2_X1 U11779 ( .A1(n13147), .A2(n13180), .Z(n11061) );
  NAND2_X2 U11782 ( .A1(n12452), .A2(n17098), .ZN(n21671) );
  NAND2_X2 U11785 ( .A1(n16851), .A2(n26468), .ZN(n12452) );
  XOR2_X1 U11787 ( .A1(n23371), .A2(n25040), .Z(n7411) );
  XOR2_X1 U11789 ( .A1(n22229), .A2(n8282), .Z(n5356) );
  OR2_X1 U11790 ( .A1(n33934), .A2(n33082), .Z(n22430) );
  NAND2_X2 U11793 ( .A1(n7144), .A2(n8602), .ZN(n32519) );
  NAND2_X1 U11794 ( .A1(n8926), .A2(n25176), .ZN(n11468) );
  NAND2_X2 U11798 ( .A1(n33620), .A2(n11111), .ZN(n8926) );
  XOR2_X1 U11803 ( .A1(n24358), .A2(n16416), .Z(n24719) );
  NAND2_X2 U11806 ( .A1(n14642), .A2(n17053), .ZN(n10261) );
  AND2_X1 U11808 ( .A1(n32926), .A2(n4862), .Z(n7429) );
  XOR2_X1 U11809 ( .A1(n22186), .A2(n9369), .Z(n5796) );
  XOR2_X1 U11813 ( .A1(n14639), .A2(n22080), .Z(n22186) );
  AOI22_X2 U11816 ( .A1(n32088), .A2(n33787), .B1(n7857), .B2(n28649), .ZN(
        n3170) );
  NOR2_X2 U11823 ( .A1(n33132), .A2(n25979), .ZN(n7857) );
  NAND2_X2 U11829 ( .A1(n32521), .A2(n17079), .ZN(n14640) );
  NAND2_X2 U11830 ( .A1(n33286), .A2(n9691), .ZN(n32881) );
  NAND3_X2 U11832 ( .A1(n11657), .A2(n14829), .A3(n11656), .ZN(n27130) );
  NOR2_X2 U11834 ( .A1(n11659), .A2(n11658), .ZN(n11657) );
  AOI21_X2 U11838 ( .A1(n5619), .A2(n5055), .B(n5054), .ZN(n12652) );
  OAI22_X2 U11839 ( .A1(n5618), .A2(n13597), .B1(n22886), .B2(n12511), .ZN(
        n5054) );
  XOR2_X1 U11842 ( .A1(n23261), .A2(n23237), .Z(n12573) );
  XOR2_X1 U11843 ( .A1(n7229), .A2(n23120), .Z(n23261) );
  NOR2_X2 U11844 ( .A1(n25446), .A2(n25444), .ZN(n25433) );
  NOR2_X2 U11845 ( .A1(n25058), .A2(n25062), .ZN(n17729) );
  NOR2_X2 U11854 ( .A1(n32523), .A2(n7649), .ZN(n6322) );
  NOR2_X1 U11857 ( .A1(n22596), .A2(n7633), .ZN(n32523) );
  INV_X2 U11859 ( .I(n10924), .ZN(n887) );
  NAND2_X2 U11861 ( .A1(n2153), .A2(n2154), .ZN(n10924) );
  XOR2_X1 U11864 ( .A1(n32524), .A2(n25436), .Z(Ciphertext[105]) );
  NAND2_X1 U11873 ( .A1(n25434), .A2(n33159), .ZN(n32524) );
  NOR2_X2 U11877 ( .A1(n29392), .A2(n32525), .ZN(n6400) );
  XOR2_X1 U11879 ( .A1(n33333), .A2(n22779), .Z(n11568) );
  XOR2_X1 U11886 ( .A1(n4047), .A2(n11668), .Z(n22779) );
  OAI21_X2 U11887 ( .A1(n33963), .A2(n32526), .B(n23699), .ZN(n5051) );
  AOI21_X2 U11890 ( .A1(n2949), .A2(n21771), .B(n2948), .ZN(n22173) );
  OAI22_X2 U11892 ( .A1(n1015), .A2(n38), .B1(n2368), .B2(n33766), .ZN(n21771)
         );
  XOR2_X1 U11893 ( .A1(n32527), .A2(n25728), .Z(Ciphertext[154]) );
  NAND4_X2 U11894 ( .A1(n25727), .A2(n25726), .A3(n34019), .A4(n25725), .ZN(
        n32527) );
  NAND2_X2 U11896 ( .A1(n31921), .A2(n13532), .ZN(n25593) );
  XOR2_X1 U11897 ( .A1(n27613), .A2(n1102), .Z(n23501) );
  NAND2_X2 U11901 ( .A1(n7217), .A2(n7724), .ZN(n27613) );
  XOR2_X1 U11905 ( .A1(n14058), .A2(n24819), .Z(n16838) );
  XOR2_X1 U11912 ( .A1(n32529), .A2(n25091), .Z(Ciphertext[49]) );
  NOR3_X1 U11913 ( .A1(n16226), .A2(n16933), .A3(n4518), .ZN(n33167) );
  BUF_X2 U11919 ( .I(n18254), .Z(n32530) );
  BUF_X2 U11926 ( .I(n22945), .Z(n32531) );
  NOR2_X2 U11928 ( .A1(n11259), .A2(n11258), .ZN(n32933) );
  BUF_X2 U11938 ( .I(n34161), .Z(n32532) );
  INV_X1 U11941 ( .I(n19167), .ZN(n33845) );
  AOI22_X2 U11946 ( .A1(n22839), .A2(n29329), .B1(n22840), .B2(n8990), .ZN(
        n33001) );
  OAI21_X1 U11955 ( .A1(n8923), .A2(n9954), .B(n32710), .ZN(n10495) );
  AOI22_X2 U11958 ( .A1(n17286), .A2(n23786), .B1(n17157), .B2(n15692), .ZN(
        n841) );
  NAND2_X2 U11960 ( .A1(n4110), .A2(n22832), .ZN(n17503) );
  NAND2_X2 U11971 ( .A1(n3520), .A2(n29349), .ZN(n4110) );
  XOR2_X1 U11974 ( .A1(n23533), .A2(n23529), .Z(n32841) );
  NAND2_X2 U11976 ( .A1(n4651), .A2(n4650), .ZN(n23529) );
  XOR2_X1 U11980 ( .A1(n32533), .A2(n24399), .Z(n34030) );
  XOR2_X1 U11982 ( .A1(n7574), .A2(n12493), .Z(n24399) );
  INV_X2 U11983 ( .I(n15588), .ZN(n32533) );
  NOR2_X2 U11985 ( .A1(n33132), .A2(n30365), .ZN(n7797) );
  NAND3_X2 U11987 ( .A1(n17773), .A2(n27024), .A3(n15655), .ZN(n21276) );
  NOR3_X2 U11989 ( .A1(n2657), .A2(n2656), .A3(n13143), .ZN(n32534) );
  NOR2_X1 U11992 ( .A1(n25784), .A2(n33720), .ZN(n25779) );
  NAND2_X1 U11994 ( .A1(n25779), .A2(n25790), .ZN(n25780) );
  NAND4_X2 U12002 ( .A1(n4899), .A2(n3820), .A3(n24365), .A4(n4898), .ZN(
        n32977) );
  NAND2_X2 U12003 ( .A1(n32536), .A2(n31531), .ZN(n32842) );
  NAND2_X2 U12006 ( .A1(n29329), .A2(n22978), .ZN(n32536) );
  XNOR2_X1 U12008 ( .A1(n21020), .A2(n20782), .ZN(n20168) );
  XOR2_X1 U12012 ( .A1(n20720), .A2(n10949), .Z(n20782) );
  INV_X2 U12013 ( .I(n7), .ZN(n630) );
  NOR2_X2 U12014 ( .A1(n75), .A2(n12929), .ZN(n9500) );
  AOI22_X2 U12016 ( .A1(n32658), .A2(n28314), .B1(n12728), .B2(n12727), .ZN(
        n30433) );
  AOI21_X2 U12022 ( .A1(n4375), .A2(n18204), .B(n4374), .ZN(n7188) );
  NAND2_X2 U12028 ( .A1(n25486), .A2(n25462), .ZN(n25482) );
  OR2_X1 U12030 ( .A1(n24335), .A2(n24242), .Z(n33669) );
  AOI21_X2 U12031 ( .A1(n22633), .A2(n11932), .B(n32512), .ZN(n7179) );
  INV_X2 U12046 ( .I(n32538), .ZN(n22633) );
  NOR2_X2 U12048 ( .A1(n522), .A2(n17916), .ZN(n32538) );
  NOR2_X1 U12049 ( .A1(n15882), .A2(n31994), .ZN(n32717) );
  NOR2_X2 U12054 ( .A1(n33533), .A2(n29830), .ZN(n646) );
  INV_X2 U12061 ( .I(n32539), .ZN(n10569) );
  XOR2_X1 U12062 ( .A1(n2210), .A2(n2211), .Z(n32539) );
  NOR2_X1 U12063 ( .A1(n22785), .A2(n30584), .ZN(n29384) );
  XOR2_X1 U12066 ( .A1(n3368), .A2(n32540), .Z(n22199) );
  XOR2_X1 U12068 ( .A1(n22186), .A2(n28005), .Z(n32540) );
  XOR2_X1 U12071 ( .A1(n23361), .A2(n32633), .Z(n29906) );
  XOR2_X1 U12072 ( .A1(n13216), .A2(n13814), .Z(n23361) );
  NAND2_X2 U12073 ( .A1(n32541), .A2(n2508), .ZN(n26969) );
  NOR2_X2 U12074 ( .A1(n16280), .A2(n7463), .ZN(n6190) );
  NAND2_X1 U12076 ( .A1(n4097), .A2(n28099), .ZN(n13828) );
  NAND2_X2 U12078 ( .A1(n26679), .A2(n34083), .ZN(n4097) );
  NOR2_X2 U12079 ( .A1(n32598), .A2(n32542), .ZN(n22249) );
  AOI21_X2 U12080 ( .A1(n21863), .A2(n21862), .B(n1016), .ZN(n32542) );
  NAND2_X2 U12083 ( .A1(n30649), .A2(n3840), .ZN(n11438) );
  NAND2_X2 U12088 ( .A1(n30448), .A2(n33026), .ZN(n9546) );
  XOR2_X1 U12091 ( .A1(n32543), .A2(n20668), .Z(n2881) );
  XOR2_X1 U12102 ( .A1(n2883), .A2(n31233), .Z(n32543) );
  XOR2_X1 U12103 ( .A1(n12652), .A2(n23200), .Z(n23343) );
  OR2_X1 U12106 ( .A1(n21395), .A2(n6681), .Z(n16058) );
  INV_X2 U12110 ( .I(n4862), .ZN(n32605) );
  OAI21_X2 U12112 ( .A1(n21414), .A2(n21413), .B(n1332), .ZN(n9905) );
  NOR2_X2 U12116 ( .A1(n29143), .A2(n28700), .ZN(n4287) );
  AOI22_X2 U12119 ( .A1(n32544), .A2(n21269), .B1(n28642), .B2(n29460), .ZN(
        n4082) );
  NOR2_X2 U12124 ( .A1(n28642), .A2(n21267), .ZN(n32544) );
  AND2_X2 U12126 ( .A1(n25198), .A2(n11985), .Z(n26015) );
  NAND2_X2 U12127 ( .A1(n32545), .A2(n7754), .ZN(n7753) );
  NAND2_X1 U12131 ( .A1(n27245), .A2(n27246), .ZN(n32545) );
  BUF_X4 U12133 ( .I(n22487), .Z(n33046) );
  NAND2_X2 U12134 ( .A1(n12443), .A2(n14617), .ZN(n23295) );
  NOR2_X1 U12137 ( .A1(n22592), .A2(n17408), .ZN(n17212) );
  AOI21_X2 U12139 ( .A1(n11246), .A2(n28131), .B(n26925), .ZN(n22592) );
  AOI22_X2 U12145 ( .A1(n28128), .A2(n9854), .B1(n20550), .B2(n125), .ZN(
        n32546) );
  AND2_X1 U12146 ( .A1(n4281), .A2(n18204), .Z(n7263) );
  AOI21_X2 U12148 ( .A1(n30219), .A2(n20955), .B(n2301), .ZN(n21020) );
  NAND2_X2 U12152 ( .A1(n32957), .A2(n34128), .ZN(n21188) );
  AOI21_X2 U12157 ( .A1(n1257), .A2(n844), .B(n23867), .ZN(n32547) );
  XOR2_X1 U12160 ( .A1(n28747), .A2(n32548), .Z(n7624) );
  XOR2_X1 U12161 ( .A1(n10869), .A2(n7450), .Z(n32548) );
  NOR2_X2 U12167 ( .A1(n21334), .A2(n32549), .ZN(n17416) );
  AOI21_X2 U12171 ( .A1(n21332), .A2(n21331), .B(n8378), .ZN(n32549) );
  XOR2_X1 U12173 ( .A1(n20904), .A2(n20754), .Z(n21034) );
  NAND2_X2 U12181 ( .A1(n162), .A2(n26478), .ZN(n20904) );
  NAND2_X2 U12183 ( .A1(n14805), .A2(n29278), .ZN(n12440) );
  XOR2_X1 U12184 ( .A1(n34160), .A2(n22098), .Z(n22229) );
  INV_X2 U12188 ( .I(n24810), .ZN(n9209) );
  XOR2_X1 U12200 ( .A1(n8754), .A2(n32554), .Z(n19899) );
  XOR2_X1 U12201 ( .A1(n7589), .A2(n7590), .Z(n32554) );
  OAI21_X1 U12202 ( .A1(n19322), .A2(n30894), .B(n19068), .ZN(n3132) );
  NAND2_X1 U12205 ( .A1(n21706), .A2(n15414), .ZN(n21754) );
  NAND3_X2 U12207 ( .A1(n15435), .A2(n15436), .A3(n32555), .ZN(n20305) );
  NAND2_X2 U12209 ( .A1(n29281), .A2(n19998), .ZN(n32555) );
  XOR2_X1 U12210 ( .A1(n22153), .A2(n22190), .Z(n5013) );
  NOR2_X2 U12213 ( .A1(n31940), .A2(n32556), .ZN(n33349) );
  XOR2_X1 U12214 ( .A1(n9914), .A2(n22161), .Z(n1938) );
  XOR2_X1 U12229 ( .A1(n8291), .A2(n3723), .Z(n22161) );
  XOR2_X1 U12231 ( .A1(n24602), .A2(n32557), .Z(n30220) );
  XOR2_X1 U12234 ( .A1(n15264), .A2(n4997), .Z(n32557) );
  OAI22_X2 U12236 ( .A1(n29630), .A2(n29629), .B1(n4886), .B2(n4885), .ZN(
        n12257) );
  INV_X2 U12261 ( .I(n11173), .ZN(n4885) );
  XOR2_X1 U12264 ( .A1(n10473), .A2(n10475), .Z(n11173) );
  XOR2_X1 U12267 ( .A1(n5253), .A2(n32558), .Z(n8939) );
  XNOR2_X1 U12290 ( .A1(n27114), .A2(n24522), .ZN(n5253) );
  INV_X2 U12291 ( .I(n24746), .ZN(n32558) );
  XOR2_X1 U12297 ( .A1(n14058), .A2(n25801), .Z(n13520) );
  OR2_X1 U12298 ( .A1(n10496), .A2(n22945), .Z(n32710) );
  AOI21_X2 U12302 ( .A1(n32560), .A2(n15718), .B(n22916), .ZN(n31399) );
  XOR2_X1 U12309 ( .A1(n5658), .A2(n10989), .Z(n5657) );
  AOI21_X2 U12312 ( .A1(n17860), .A2(n24029), .B(n32561), .ZN(n24847) );
  NOR3_X2 U12316 ( .A1(n28590), .A2(n9066), .A3(n4118), .ZN(n32561) );
  XOR2_X1 U12318 ( .A1(n32562), .A2(n31098), .Z(n26515) );
  XOR2_X1 U12319 ( .A1(n23459), .A2(n2862), .Z(n32562) );
  AOI21_X2 U12325 ( .A1(n31469), .A2(n31471), .B(n111), .ZN(n12991) );
  XOR2_X1 U12327 ( .A1(n32563), .A2(n17865), .Z(n31639) );
  XOR2_X1 U12328 ( .A1(n34088), .A2(n2278), .Z(n32563) );
  XOR2_X1 U12331 ( .A1(n14058), .A2(n24853), .Z(n24854) );
  NOR2_X2 U12333 ( .A1(n24238), .A2(n24239), .ZN(n24853) );
  INV_X2 U12335 ( .I(n23186), .ZN(n982) );
  OAI22_X2 U12342 ( .A1(n17083), .A2(n17639), .B1(n17085), .B2(n22884), .ZN(
        n23186) );
  XOR2_X1 U12345 ( .A1(n33606), .A2(n5215), .Z(n8251) );
  NAND2_X2 U12347 ( .A1(n14542), .A2(n32515), .ZN(n4458) );
  OAI22_X2 U12351 ( .A1(n21554), .A2(n32613), .B1(n21555), .B2(n21556), .ZN(
        n28413) );
  BUF_X2 U12353 ( .I(n22306), .Z(n32564) );
  NAND2_X2 U12354 ( .A1(n974), .A2(n33832), .ZN(n24235) );
  INV_X2 U12358 ( .I(n18665), .ZN(n2509) );
  NAND2_X2 U12360 ( .A1(n31972), .A2(n31971), .ZN(n18665) );
  XOR2_X1 U12363 ( .A1(n32566), .A2(n26001), .Z(Ciphertext[45]) );
  XOR2_X1 U12367 ( .A1(n12621), .A2(n12624), .Z(n30038) );
  XOR2_X1 U12369 ( .A1(n32567), .A2(n25040), .Z(Ciphertext[38]) );
  NAND2_X1 U12371 ( .A1(n6424), .A2(n33145), .ZN(n32567) );
  OAI21_X2 U12373 ( .A1(n32569), .A2(n32568), .B(n32483), .ZN(n17001) );
  NAND2_X2 U12374 ( .A1(n33585), .A2(n32571), .ZN(n32570) );
  INV_X2 U12375 ( .I(n28338), .ZN(n32571) );
  XOR2_X1 U12377 ( .A1(n14969), .A2(n32572), .Z(n32838) );
  XOR2_X1 U12380 ( .A1(n22198), .A2(n32573), .Z(n32572) );
  INV_X1 U12384 ( .I(n16697), .ZN(n32573) );
  NOR2_X2 U12385 ( .A1(n13696), .A2(n7953), .ZN(n20755) );
  NAND2_X2 U12386 ( .A1(n20459), .A2(n28899), .ZN(n162) );
  OAI22_X2 U12387 ( .A1(n32594), .A2(n27741), .B1(n1158), .B2(n20614), .ZN(
        n20459) );
  XOR2_X1 U12388 ( .A1(n4287), .A2(n31311), .Z(n6863) );
  NOR3_X2 U12389 ( .A1(n32574), .A2(n29037), .A3(n9736), .ZN(n33748) );
  NOR2_X1 U12390 ( .A1(n4423), .A2(n16313), .ZN(n4422) );
  XOR2_X1 U12392 ( .A1(n33267), .A2(n18107), .Z(n33391) );
  XOR2_X1 U12396 ( .A1(n32916), .A2(n32575), .Z(n15093) );
  XOR2_X1 U12397 ( .A1(n24475), .A2(n27115), .Z(n24547) );
  NOR2_X2 U12399 ( .A1(n32576), .A2(n7017), .ZN(n22302) );
  NAND2_X1 U12400 ( .A1(n8174), .A2(n11536), .ZN(n32576) );
  OAI21_X2 U12409 ( .A1(n14245), .A2(n14247), .B(n14243), .ZN(n25378) );
  OAI21_X2 U12410 ( .A1(n31962), .A2(n33915), .B(n33914), .ZN(n14245) );
  NAND2_X2 U12411 ( .A1(n30015), .A2(n12705), .ZN(n5003) );
  XOR2_X1 U12414 ( .A1(n19616), .A2(n19615), .Z(n19617) );
  OAI21_X2 U12416 ( .A1(n17453), .A2(n28120), .B(n15253), .ZN(n14288) );
  XOR2_X1 U12419 ( .A1(n6735), .A2(n32578), .Z(n9322) );
  XOR2_X1 U12425 ( .A1(n6739), .A2(n16178), .Z(n32578) );
  NAND2_X1 U12426 ( .A1(n3772), .A2(n3771), .ZN(n32615) );
  OAI22_X2 U12428 ( .A1(n32579), .A2(n25007), .B1(n3231), .B2(n3230), .ZN(
        n31182) );
  AOI21_X2 U12429 ( .A1(n3230), .A2(n25002), .B(n31122), .ZN(n32579) );
  NAND3_X2 U12430 ( .A1(n28776), .A2(n29401), .A3(n32580), .ZN(n23508) );
  NAND2_X2 U12433 ( .A1(n5091), .A2(n25709), .ZN(n4706) );
  NOR2_X1 U12434 ( .A1(n8086), .A2(n24212), .ZN(n26914) );
  INV_X4 U12435 ( .I(n21601), .ZN(n5704) );
  NAND2_X2 U12437 ( .A1(n7651), .A2(n329), .ZN(n21601) );
  XOR2_X1 U12444 ( .A1(n86), .A2(n85), .Z(n22656) );
  NOR2_X2 U12445 ( .A1(n3515), .A2(n6763), .ZN(n5032) );
  XOR2_X1 U12449 ( .A1(n28405), .A2(n32582), .Z(n13189) );
  XOR2_X1 U12459 ( .A1(n14968), .A2(n20640), .Z(n32582) );
  NAND2_X2 U12460 ( .A1(n12577), .A2(n23071), .ZN(n6676) );
  XOR2_X1 U12461 ( .A1(n21001), .A2(n20730), .Z(n16175) );
  OAI21_X2 U12464 ( .A1(n13783), .A2(n13784), .B(n13782), .ZN(n21001) );
  INV_X4 U12465 ( .I(n3515), .ZN(n2935) );
  XOR2_X1 U12466 ( .A1(n24807), .A2(n4329), .Z(n9571) );
  NAND2_X2 U12474 ( .A1(n27660), .A2(n27439), .ZN(n24807) );
  NAND2_X2 U12476 ( .A1(n11557), .A2(n12770), .ZN(n2958) );
  AOI22_X2 U12477 ( .A1(n20036), .A2(n2549), .B1(n14210), .B2(n12337), .ZN(
        n12770) );
  NAND2_X1 U12486 ( .A1(n13130), .A2(n21506), .ZN(n11687) );
  NAND2_X2 U12487 ( .A1(n33052), .A2(n28485), .ZN(n20670) );
  NAND2_X2 U12488 ( .A1(n8107), .A2(n11872), .ZN(n12296) );
  NAND2_X2 U12494 ( .A1(n20238), .A2(n11453), .ZN(n20075) );
  NOR2_X2 U12495 ( .A1(n11454), .A2(n2387), .ZN(n11453) );
  XOR2_X1 U12496 ( .A1(n7748), .A2(n25274), .Z(n4944) );
  NAND2_X2 U12500 ( .A1(n7108), .A2(n7109), .ZN(n7748) );
  OAI21_X2 U12502 ( .A1(n31507), .A2(n31730), .B(n21445), .ZN(n21827) );
  AOI22_X2 U12503 ( .A1(n21307), .A2(n21305), .B1(n16526), .B2(n21443), .ZN(
        n21445) );
  INV_X2 U12505 ( .I(n32584), .ZN(n29460) );
  XOR2_X1 U12507 ( .A1(n17281), .A2(n6205), .Z(n32584) );
  OAI21_X2 U12514 ( .A1(n33850), .A2(n9393), .B(n9392), .ZN(n32898) );
  NOR2_X2 U12516 ( .A1(n8380), .A2(n17805), .ZN(n24234) );
  NAND2_X1 U12518 ( .A1(n33383), .A2(n33382), .ZN(n7217) );
  NAND3_X2 U12531 ( .A1(n1873), .A2(n9339), .A3(n9338), .ZN(n30031) );
  XOR2_X1 U12533 ( .A1(n11490), .A2(n19531), .Z(n14316) );
  NAND2_X2 U12536 ( .A1(n18669), .A2(n18668), .ZN(n11490) );
  NAND2_X2 U12539 ( .A1(n33536), .A2(n31932), .ZN(n22455) );
  XOR2_X1 U12540 ( .A1(n2423), .A2(n32586), .Z(n8492) );
  XOR2_X1 U12541 ( .A1(n17682), .A2(n24752), .Z(n32586) );
  AOI21_X2 U12542 ( .A1(n4071), .A2(n20541), .B(n782), .ZN(n10718) );
  NAND2_X2 U12550 ( .A1(n7123), .A2(n7120), .ZN(n30346) );
  NAND2_X2 U12553 ( .A1(n7118), .A2(n27515), .ZN(n7123) );
  OAI21_X1 U12558 ( .A1(n1628), .A2(n4150), .B(n1627), .ZN(n32587) );
  NOR2_X2 U12564 ( .A1(n30769), .A2(n21697), .ZN(n32588) );
  NAND2_X2 U12570 ( .A1(n19198), .A2(n19200), .ZN(n28883) );
  NAND2_X2 U12573 ( .A1(n5813), .A2(n19199), .ZN(n19198) );
  XOR2_X1 U12574 ( .A1(n14855), .A2(n13470), .Z(n4729) );
  INV_X2 U12575 ( .I(n29278), .ZN(n32590) );
  NAND2_X2 U12580 ( .A1(n1214), .A2(n30241), .ZN(n32592) );
  INV_X2 U12581 ( .I(n28358), .ZN(n25210) );
  NAND2_X2 U12582 ( .A1(n4533), .A2(n33024), .ZN(n28358) );
  XOR2_X1 U12585 ( .A1(n4354), .A2(n32593), .Z(n14911) );
  XOR2_X1 U12587 ( .A1(n4352), .A2(n4353), .Z(n32593) );
  AND2_X2 U12588 ( .A1(n8838), .A2(n23834), .Z(n30060) );
  BUF_X2 U12589 ( .I(n17746), .Z(n32594) );
  NAND3_X1 U12593 ( .A1(n32596), .A2(n849), .A3(n32595), .ZN(n27263) );
  INV_X2 U12594 ( .I(n13807), .ZN(n32595) );
  INV_X1 U12595 ( .I(n23066), .ZN(n32596) );
  NAND2_X1 U12596 ( .A1(n18842), .A2(n33232), .ZN(n33231) );
  AOI21_X2 U12597 ( .A1(n3219), .A2(n25974), .B(n32597), .ZN(n3234) );
  AND2_X1 U12601 ( .A1(n3221), .A2(n3222), .Z(n32597) );
  NAND2_X2 U12603 ( .A1(n2727), .A2(n2642), .ZN(n25142) );
  XOR2_X1 U12604 ( .A1(n32111), .A2(n20992), .Z(n12330) );
  INV_X2 U12611 ( .I(n31017), .ZN(n16623) );
  XOR2_X1 U12612 ( .A1(n33604), .A2(n4840), .Z(n25894) );
  AOI21_X2 U12614 ( .A1(n30154), .A2(n16241), .B(n30152), .ZN(n32598) );
  XOR2_X1 U12615 ( .A1(n23145), .A2(n6348), .Z(n5194) );
  XOR2_X1 U12621 ( .A1(n23271), .A2(n33971), .Z(n6348) );
  OAI22_X2 U12624 ( .A1(n16623), .A2(n5707), .B1(n20000), .B2(n10845), .ZN(
        n7281) );
  INV_X2 U12631 ( .I(n10708), .ZN(n10845) );
  NAND2_X2 U12633 ( .A1(n25138), .A2(n32599), .ZN(n14189) );
  NAND2_X2 U12635 ( .A1(n32601), .A2(n32600), .ZN(n32599) );
  NOR2_X2 U12636 ( .A1(n11372), .A2(n9162), .ZN(n32600) );
  INV_X2 U12637 ( .I(n17824), .ZN(n32601) );
  XOR2_X1 U12638 ( .A1(n27121), .A2(n14613), .Z(n23521) );
  OAI21_X2 U12641 ( .A1(n32056), .A2(n32603), .B(n30817), .ZN(n10297) );
  NOR2_X1 U12642 ( .A1(n11444), .A2(n6290), .ZN(n32603) );
  BUF_X2 U12643 ( .I(n29693), .Z(n32604) );
  INV_X1 U12644 ( .I(n10630), .ZN(n22631) );
  NAND2_X2 U12646 ( .A1(n32606), .A2(n32605), .ZN(n10630) );
  INV_X2 U12647 ( .I(n7513), .ZN(n32606) );
  NOR2_X2 U12650 ( .A1(n29972), .A2(n20261), .ZN(n29528) );
  NAND2_X2 U12652 ( .A1(n32607), .A2(n27340), .ZN(n13412) );
  NAND2_X1 U12653 ( .A1(n14531), .A2(n7765), .ZN(n12458) );
  XOR2_X1 U12657 ( .A1(n11205), .A2(n15710), .Z(n32925) );
  OAI21_X2 U12659 ( .A1(n7626), .A2(n5895), .B(n5893), .ZN(n15710) );
  NAND3_X2 U12662 ( .A1(n31657), .A2(n14305), .A3(n32608), .ZN(n15825) );
  NAND3_X2 U12663 ( .A1(n32674), .A2(n8431), .A3(n19547), .ZN(n7102) );
  INV_X2 U12665 ( .I(n12758), .ZN(n9404) );
  NAND2_X2 U12666 ( .A1(n20471), .A2(n32504), .ZN(n12758) );
  NOR2_X1 U12667 ( .A1(n1597), .A2(n25746), .ZN(n24431) );
  NAND2_X2 U12671 ( .A1(n31591), .A2(n27486), .ZN(n1597) );
  AOI22_X2 U12672 ( .A1(n2873), .A2(n15162), .B1(n8998), .B2(n14568), .ZN(
        n14567) );
  XOR2_X1 U12673 ( .A1(n1173), .A2(n17091), .Z(n19662) );
  NAND2_X2 U12675 ( .A1(n33407), .A2(n13791), .ZN(n17091) );
  AND2_X1 U12677 ( .A1(n5673), .A2(n4286), .Z(n31419) );
  INV_X2 U12678 ( .I(n6479), .ZN(n32610) );
  OAI22_X2 U12684 ( .A1(n32612), .A2(n28806), .B1(n4384), .B2(n4387), .ZN(
        n10915) );
  XOR2_X1 U12688 ( .A1(n14206), .A2(n20652), .Z(n20710) );
  NAND2_X2 U12690 ( .A1(n20204), .A2(n20203), .ZN(n14206) );
  INV_X1 U12691 ( .I(n22426), .ZN(n32988) );
  INV_X2 U12692 ( .I(n7072), .ZN(n1805) );
  AND2_X1 U12699 ( .A1(n7868), .A2(n11401), .Z(n6807) );
  BUF_X2 U12703 ( .I(n32800), .Z(n32613) );
  XOR2_X1 U12707 ( .A1(n28897), .A2(n11691), .Z(n32614) );
  NOR2_X2 U12708 ( .A1(n18914), .A2(n27076), .ZN(n19483) );
  XOR2_X1 U12710 ( .A1(n10482), .A2(n1130), .Z(n417) );
  XOR2_X1 U12711 ( .A1(n22127), .A2(n8533), .Z(n1130) );
  XOR2_X1 U12715 ( .A1(n32615), .A2(n16619), .Z(Ciphertext[96]) );
  XOR2_X1 U12720 ( .A1(n24650), .A2(n24649), .Z(n33663) );
  XOR2_X1 U12722 ( .A1(n968), .A2(n24799), .Z(n24650) );
  XOR2_X1 U12724 ( .A1(n27516), .A2(n32616), .Z(n24511) );
  XOR2_X1 U12731 ( .A1(n24825), .A2(n24508), .Z(n32616) );
  INV_X2 U12734 ( .I(n32617), .ZN(n12488) );
  XNOR2_X1 U12737 ( .A1(n31054), .A2(n3120), .ZN(n32617) );
  NOR2_X1 U12739 ( .A1(n17030), .A2(n17029), .ZN(n18412) );
  NOR3_X2 U12740 ( .A1(n2137), .A2(n2138), .A3(n2135), .ZN(n12375) );
  OR2_X1 U12743 ( .A1(n27897), .A2(n3536), .Z(n22490) );
  XOR2_X1 U12746 ( .A1(n21907), .A2(n33300), .Z(n27897) );
  AND2_X1 U12747 ( .A1(n15964), .A2(n25586), .Z(n24631) );
  XOR2_X1 U12748 ( .A1(n32255), .A2(n3722), .Z(n22037) );
  BUF_X2 U12751 ( .I(n20043), .Z(n32618) );
  BUF_X2 U12752 ( .I(n10714), .Z(n32619) );
  XOR2_X1 U12756 ( .A1(n32620), .A2(n31852), .Z(n20483) );
  XOR2_X1 U12759 ( .A1(n20993), .A2(n20482), .Z(n32620) );
  XOR2_X1 U12760 ( .A1(n22251), .A2(n29693), .Z(n22150) );
  OAI22_X2 U12763 ( .A1(n12328), .A2(n6660), .B1(n21776), .B2(n21775), .ZN(
        n22251) );
  AND2_X1 U12764 ( .A1(n13667), .A2(n25123), .Z(n33413) );
  OAI21_X2 U12768 ( .A1(n32621), .A2(n4596), .B(n19140), .ZN(n4595) );
  INV_X2 U12771 ( .I(n19189), .ZN(n32621) );
  NAND2_X2 U12772 ( .A1(n744), .A2(n13160), .ZN(n19189) );
  INV_X1 U12777 ( .I(n31325), .ZN(n32837) );
  NAND3_X2 U12778 ( .A1(n880), .A2(n7732), .A3(n11970), .ZN(n32622) );
  BUF_X2 U12779 ( .I(n21203), .Z(n32625) );
  NAND2_X2 U12783 ( .A1(n17771), .A2(n32626), .ZN(n24996) );
  NAND2_X2 U12786 ( .A1(n34099), .A2(n1559), .ZN(n21532) );
  NOR2_X2 U12787 ( .A1(n22362), .A2(n8471), .ZN(n22542) );
  NAND2_X2 U12789 ( .A1(n10489), .A2(n10486), .ZN(n8568) );
  XOR2_X1 U12791 ( .A1(n32627), .A2(n6903), .Z(n7912) );
  XOR2_X1 U12802 ( .A1(n30482), .A2(n30362), .Z(n32627) );
  AOI22_X2 U12803 ( .A1(n10054), .A2(n19109), .B1(n19110), .B2(n27921), .ZN(
        n28996) );
  INV_X2 U12804 ( .I(n32628), .ZN(n26448) );
  XNOR2_X1 U12806 ( .A1(n9040), .A2(n9037), .ZN(n32628) );
  XOR2_X1 U12812 ( .A1(n29702), .A2(n19631), .Z(n14814) );
  NAND2_X1 U12818 ( .A1(n22745), .A2(n27166), .ZN(n33503) );
  XOR2_X1 U12821 ( .A1(n31639), .A2(n32629), .Z(n24779) );
  XOR2_X1 U12830 ( .A1(n24619), .A2(n33348), .Z(n32629) );
  AOI21_X1 U12840 ( .A1(n32630), .A2(n16273), .B(n12457), .ZN(n12456) );
  NAND2_X1 U12843 ( .A1(n12458), .A2(n16279), .ZN(n32630) );
  OR2_X1 U12845 ( .A1(n24027), .A2(n32934), .Z(n29292) );
  INV_X2 U12848 ( .I(n32631), .ZN(n22670) );
  XOR2_X1 U12853 ( .A1(n24825), .A2(n32632), .Z(n27946) );
  XOR2_X1 U12854 ( .A1(n4240), .A2(n12665), .Z(n32632) );
  XOR2_X1 U12855 ( .A1(n23174), .A2(n23189), .Z(n32633) );
  NAND2_X1 U12859 ( .A1(n4814), .A2(n24976), .ZN(n32735) );
  NAND2_X2 U12860 ( .A1(n12642), .A2(n11214), .ZN(n12866) );
  NOR2_X2 U12862 ( .A1(n29047), .A2(n29093), .ZN(n32634) );
  XOR2_X1 U12863 ( .A1(n19538), .A2(n32184), .Z(n14743) );
  NAND2_X2 U12866 ( .A1(n14749), .A2(n14750), .ZN(n32635) );
  AOI21_X2 U12875 ( .A1(n8499), .A2(n5690), .B(n27592), .ZN(n10793) );
  OAI22_X2 U12876 ( .A1(n9516), .A2(n9334), .B1(n32636), .B2(n9647), .ZN(
        n22949) );
  AOI22_X2 U12878 ( .A1(n14993), .A2(n25013), .B1(n24976), .B2(n14992), .ZN(
        n32637) );
  OAI22_X2 U12882 ( .A1(n5264), .A2(n1317), .B1(n21821), .B2(n5546), .ZN(
        n21562) );
  XOR2_X1 U12885 ( .A1(n29674), .A2(n26371), .Z(n30187) );
  XOR2_X1 U12890 ( .A1(n2809), .A2(n32638), .Z(n27894) );
  XOR2_X1 U12895 ( .A1(n33933), .A2(n32639), .Z(n32638) );
  XOR2_X1 U12898 ( .A1(n9983), .A2(n32640), .Z(n33253) );
  XOR2_X1 U12900 ( .A1(n23331), .A2(n23332), .Z(n23437) );
  NOR2_X2 U12901 ( .A1(n2086), .A2(n32641), .ZN(n10523) );
  AOI21_X2 U12902 ( .A1(n10524), .A2(n20338), .B(n20591), .ZN(n32641) );
  AND2_X1 U12904 ( .A1(n30233), .A2(n32643), .Z(n34148) );
  NOR2_X1 U12906 ( .A1(n33565), .A2(n26615), .ZN(n33187) );
  XOR2_X1 U12907 ( .A1(n19466), .A2(n16584), .Z(n19385) );
  OAI22_X2 U12912 ( .A1(n27420), .A2(n16741), .B1(n7419), .B2(n18751), .ZN(
        n19466) );
  BUF_X2 U12916 ( .I(n9678), .Z(n32644) );
  NAND2_X2 U12917 ( .A1(n792), .A2(n13601), .ZN(n24269) );
  XOR2_X1 U12919 ( .A1(n11736), .A2(n22227), .Z(n22143) );
  NAND2_X2 U12920 ( .A1(n13029), .A2(n3050), .ZN(n11736) );
  NAND2_X1 U12922 ( .A1(n32712), .A2(n16976), .ZN(n26858) );
  NAND2_X2 U12923 ( .A1(n33044), .A2(n31946), .ZN(n7586) );
  AOI22_X2 U12926 ( .A1(n16673), .A2(n25859), .B1(n14915), .B2(n25863), .ZN(
        n25836) );
  XOR2_X1 U12932 ( .A1(n32645), .A2(n23407), .Z(n236) );
  NOR2_X2 U12933 ( .A1(n9277), .A2(n29138), .ZN(n10226) );
  XOR2_X1 U12935 ( .A1(n32646), .A2(n29609), .Z(Ciphertext[50]) );
  OAI22_X1 U12936 ( .A1(n29076), .A2(n25097), .B1(n25095), .B2(n4193), .ZN(
        n32646) );
  NAND2_X2 U12938 ( .A1(n5897), .A2(n14454), .ZN(n15646) );
  NOR2_X2 U12939 ( .A1(n14281), .A2(n16009), .ZN(n7643) );
  AOI22_X2 U12940 ( .A1(n29180), .A2(n28581), .B1(n10875), .B2(n9793), .ZN(
        n29577) );
  OAI21_X1 U12941 ( .A1(n14117), .A2(n18460), .B(n15070), .ZN(n15069) );
  NOR2_X2 U12942 ( .A1(n33688), .A2(n33687), .ZN(n14117) );
  OAI21_X2 U12945 ( .A1(n1278), .A2(n6975), .B(n22747), .ZN(n22784) );
  NAND2_X2 U12946 ( .A1(n15633), .A2(n14540), .ZN(n22747) );
  NOR2_X1 U12954 ( .A1(n31967), .A2(n3084), .ZN(n3085) );
  NAND2_X2 U12966 ( .A1(n33439), .A2(n3061), .ZN(n3084) );
  NOR2_X1 U12967 ( .A1(n18715), .A2(n18716), .ZN(n18717) );
  INV_X1 U12970 ( .I(n33153), .ZN(n32647) );
  NAND2_X2 U12973 ( .A1(n7689), .A2(n25891), .ZN(n24985) );
  XOR2_X1 U12975 ( .A1(n24751), .A2(n7135), .Z(n2423) );
  NAND2_X2 U12979 ( .A1(n10848), .A2(n20405), .ZN(n5581) );
  NAND2_X2 U12985 ( .A1(n27965), .A2(n25968), .ZN(n8051) );
  OAI21_X2 U12986 ( .A1(n32649), .A2(n33974), .B(n12531), .ZN(n13679) );
  NOR2_X1 U12987 ( .A1(n12556), .A2(n15911), .ZN(n32649) );
  OR2_X2 U12988 ( .A1(n13427), .A2(n32652), .Z(n24888) );
  XOR2_X1 U12994 ( .A1(n19307), .A2(n14459), .Z(n30770) );
  XOR2_X1 U12995 ( .A1(n29856), .A2(n19403), .Z(n29661) );
  NOR2_X1 U13002 ( .A1(n10433), .A2(n7119), .ZN(n21117) );
  XOR2_X1 U13003 ( .A1(n19598), .A2(n10210), .Z(n10079) );
  XOR2_X1 U13004 ( .A1(n2611), .A2(n19470), .Z(n19598) );
  XOR2_X1 U13005 ( .A1(n32650), .A2(n33778), .Z(n11907) );
  XOR2_X1 U13008 ( .A1(n22166), .A2(n15367), .Z(n32650) );
  XOR2_X1 U13011 ( .A1(n29906), .A2(n13214), .Z(n28034) );
  NOR2_X2 U13013 ( .A1(n20751), .A2(n17341), .ZN(n28586) );
  NAND2_X2 U13019 ( .A1(n32651), .A2(n14019), .ZN(n26557) );
  NAND2_X2 U13020 ( .A1(n30366), .A2(n13077), .ZN(n32651) );
  XOR2_X1 U13025 ( .A1(n19649), .A2(n16349), .Z(n19497) );
  NAND2_X2 U13031 ( .A1(n18421), .A2(n18420), .ZN(n19649) );
  INV_X4 U13032 ( .I(n6765), .ZN(n11981) );
  NAND2_X2 U13034 ( .A1(n12506), .A2(n26302), .ZN(n6765) );
  NAND2_X2 U13037 ( .A1(n4800), .A2(n27811), .ZN(n7465) );
  NAND2_X2 U13039 ( .A1(n33165), .A2(n33166), .ZN(n4800) );
  XOR2_X1 U13044 ( .A1(n7808), .A2(n22231), .Z(n21993) );
  NOR2_X2 U13046 ( .A1(n11053), .A2(n30634), .ZN(n7808) );
  OAI21_X2 U13053 ( .A1(n12226), .A2(n12225), .B(n10939), .ZN(n12228) );
  INV_X2 U13056 ( .I(n8492), .ZN(n32652) );
  XOR2_X1 U13058 ( .A1(n20917), .A2(n29241), .Z(n21017) );
  OAI21_X2 U13060 ( .A1(n20177), .A2(n20176), .B(n20175), .ZN(n29241) );
  NOR2_X1 U13061 ( .A1(n11876), .A2(n28721), .ZN(n32653) );
  OAI21_X2 U13062 ( .A1(n655), .A2(n34166), .B(n23891), .ZN(n1818) );
  XOR2_X1 U13063 ( .A1(n30421), .A2(n30274), .Z(n33651) );
  XOR2_X1 U13065 ( .A1(n34062), .A2(n30229), .Z(n13922) );
  NOR2_X2 U13066 ( .A1(n24148), .A2(n1775), .ZN(n1973) );
  NOR2_X2 U13076 ( .A1(n14233), .A2(n32485), .ZN(n10740) );
  NOR2_X2 U13077 ( .A1(n32654), .A2(n16232), .ZN(n14749) );
  XNOR2_X1 U13085 ( .A1(n12459), .A2(n16708), .ZN(n20746) );
  OAI21_X2 U13086 ( .A1(n28641), .A2(n7690), .B(n15589), .ZN(n32655) );
  NAND2_X1 U13091 ( .A1(n28329), .A2(n7993), .ZN(n23914) );
  NAND2_X1 U13094 ( .A1(n20565), .A2(n16515), .ZN(n11368) );
  OAI21_X2 U13098 ( .A1(n7710), .A2(n33936), .B(n23884), .ZN(n32656) );
  XOR2_X1 U13103 ( .A1(n20641), .A2(n3350), .Z(n3351) );
  NAND3_X2 U13104 ( .A1(n12846), .A2(n12847), .A3(n14263), .ZN(n20641) );
  NAND2_X1 U13107 ( .A1(n19991), .A2(n937), .ZN(n17036) );
  INV_X2 U13109 ( .I(n22615), .ZN(n32658) );
  NAND2_X2 U13111 ( .A1(n851), .A2(n22810), .ZN(n22615) );
  XOR2_X1 U13113 ( .A1(n29810), .A2(n21000), .Z(n15817) );
  XOR2_X1 U13114 ( .A1(n51), .A2(n26656), .Z(n1793) );
  NOR2_X2 U13122 ( .A1(n3951), .A2(n22652), .ZN(n51) );
  OAI21_X2 U13126 ( .A1(n13230), .A2(n21234), .B(n29577), .ZN(n34078) );
  NAND3_X2 U13131 ( .A1(n1077), .A2(n4407), .A3(n24712), .ZN(n31372) );
  XOR2_X1 U13133 ( .A1(n9353), .A2(n8949), .Z(n24568) );
  NAND3_X2 U13148 ( .A1(n28703), .A2(n1504), .A3(n27735), .ZN(n9353) );
  XOR2_X1 U13163 ( .A1(n6904), .A2(n22267), .Z(n33214) );
  XOR2_X1 U13165 ( .A1(n4228), .A2(n7477), .Z(n6904) );
  NAND3_X2 U13166 ( .A1(n19120), .A2(n19181), .A3(n19180), .ZN(n8905) );
  XOR2_X1 U13171 ( .A1(n1003), .A2(n29121), .Z(n7288) );
  NAND2_X2 U13173 ( .A1(n4880), .A2(n8122), .ZN(n29121) );
  AND2_X2 U13174 ( .A1(n2234), .A2(n29052), .Z(n27117) );
  XOR2_X1 U13177 ( .A1(n32661), .A2(n20902), .Z(n5241) );
  XOR2_X1 U13179 ( .A1(n21046), .A2(n5024), .Z(n32661) );
  OAI21_X2 U13180 ( .A1(n4514), .A2(n23787), .B(n30803), .ZN(n7935) );
  NAND2_X2 U13183 ( .A1(n25210), .A2(n5578), .ZN(n7305) );
  OAI21_X2 U13187 ( .A1(n28688), .A2(n2233), .B(n23544), .ZN(n32866) );
  NAND2_X2 U13192 ( .A1(n32662), .A2(n31967), .ZN(n29780) );
  NAND2_X2 U13194 ( .A1(n26756), .A2(n3084), .ZN(n32662) );
  AOI22_X2 U13197 ( .A1(n1280), .A2(n22981), .B1(n34163), .B2(n28934), .ZN(
        n29791) );
  OAI21_X1 U13200 ( .A1(n33500), .A2(n29362), .B(n31945), .ZN(n33728) );
  XOR2_X1 U13204 ( .A1(n15948), .A2(n11995), .Z(n25589) );
  OAI21_X2 U13206 ( .A1(n32663), .A2(n32716), .B(n22726), .ZN(n31727) );
  NAND2_X1 U13208 ( .A1(n22725), .A2(n14555), .ZN(n32663) );
  XOR2_X1 U13212 ( .A1(n22037), .A2(n33217), .Z(n12622) );
  OAI22_X2 U13213 ( .A1(n1998), .A2(n1235), .B1(n1940), .B2(n24244), .ZN(n1997) );
  NAND2_X2 U13215 ( .A1(n1235), .A2(n28374), .ZN(n1940) );
  BUF_X4 U13216 ( .I(n5440), .Z(n33320) );
  XOR2_X1 U13219 ( .A1(n1713), .A2(n32664), .Z(n7012) );
  XOR2_X1 U13228 ( .A1(n34050), .A2(n1712), .Z(n32664) );
  INV_X2 U13230 ( .I(n32665), .ZN(n17289) );
  NAND2_X2 U13231 ( .A1(n31539), .A2(n28949), .ZN(n32665) );
  INV_X1 U13233 ( .I(n23464), .ZN(n33609) );
  XOR2_X1 U13234 ( .A1(n12796), .A2(n7387), .Z(n12795) );
  NAND2_X2 U13238 ( .A1(n32666), .A2(n31359), .ZN(n16060) );
  NOR2_X2 U13239 ( .A1(n30962), .A2(n30963), .ZN(n32666) );
  NAND2_X2 U13242 ( .A1(n9775), .A2(n9773), .ZN(n12478) );
  XOR2_X1 U13244 ( .A1(n9189), .A2(n30883), .Z(n24358) );
  NOR2_X2 U13254 ( .A1(n32829), .A2(n30000), .ZN(n2691) );
  XOR2_X1 U13258 ( .A1(n15666), .A2(n15669), .Z(n15226) );
  INV_X4 U13259 ( .I(n33616), .ZN(n26120) );
  XOR2_X1 U13260 ( .A1(n6758), .A2(n27174), .Z(n6757) );
  NAND2_X2 U13262 ( .A1(n13764), .A2(n25546), .ZN(n31360) );
  NAND3_X2 U13267 ( .A1(n33327), .A2(n25535), .A3(n25534), .ZN(n13764) );
  NOR3_X2 U13269 ( .A1(n8095), .A2(n30089), .A3(n33867), .ZN(n8094) );
  NOR2_X1 U13275 ( .A1(n7080), .A2(n4951), .ZN(n32667) );
  NOR2_X2 U13277 ( .A1(n17110), .A2(n32659), .ZN(n32668) );
  NAND2_X2 U13283 ( .A1(n9472), .A2(n21870), .ZN(n21632) );
  NAND2_X2 U13284 ( .A1(n33068), .A2(n33066), .ZN(n25387) );
  NAND2_X2 U13285 ( .A1(n32669), .A2(n4991), .ZN(n7384) );
  NAND2_X2 U13287 ( .A1(n33260), .A2(n33789), .ZN(n32669) );
  NAND2_X2 U13289 ( .A1(n118), .A2(n28058), .ZN(n22979) );
  XOR2_X1 U13293 ( .A1(n1228), .A2(n6168), .Z(n24800) );
  XOR2_X1 U13295 ( .A1(n21019), .A2(n20900), .Z(n20984) );
  NAND2_X2 U13299 ( .A1(n11104), .A2(n33815), .ZN(n21019) );
  NAND2_X2 U13300 ( .A1(n3844), .A2(n30336), .ZN(n19275) );
  XOR2_X1 U13301 ( .A1(n20649), .A2(n26691), .Z(n519) );
  NAND2_X2 U13302 ( .A1(n19232), .A2(n32671), .ZN(n32670) );
  OAI21_X2 U13303 ( .A1(n28856), .A2(n10478), .B(n19825), .ZN(n32747) );
  AOI21_X2 U13309 ( .A1(n1152), .A2(n13920), .B(n32672), .ZN(n4534) );
  OAI21_X2 U13310 ( .A1(n13920), .A2(n13538), .B(n13300), .ZN(n32672) );
  NAND2_X2 U13311 ( .A1(n18206), .A2(n18208), .ZN(n6718) );
  NOR2_X2 U13312 ( .A1(n18207), .A2(n21230), .ZN(n18206) );
  NAND2_X2 U13314 ( .A1(n32673), .A2(n17944), .ZN(n6899) );
  XOR2_X1 U13318 ( .A1(n24394), .A2(n13545), .Z(n24619) );
  BUF_X4 U13319 ( .I(n16451), .Z(n11703) );
  NAND2_X2 U13327 ( .A1(n22922), .A2(n22921), .ZN(n30868) );
  NAND2_X2 U13328 ( .A1(n33433), .A2(n252), .ZN(n22922) );
  AOI22_X2 U13329 ( .A1(n5598), .A2(n15394), .B1(n820), .B2(n26130), .ZN(n8406) );
  INV_X2 U13332 ( .I(n27781), .ZN(n19691) );
  NAND2_X2 U13333 ( .A1(n32676), .A2(n32675), .ZN(n27781) );
  NAND2_X1 U13335 ( .A1(n17716), .A2(n32679), .ZN(n6145) );
  OR2_X1 U13337 ( .A1(n2386), .A2(n16077), .Z(n32679) );
  XOR2_X1 U13341 ( .A1(n24805), .A2(n12800), .Z(n13471) );
  NAND2_X2 U13342 ( .A1(n18946), .A2(n18947), .ZN(n30443) );
  AOI22_X2 U13343 ( .A1(n13197), .A2(n22396), .B1(n10757), .B2(n1124), .ZN(
        n8601) );
  OAI21_X2 U13346 ( .A1(n7110), .A2(n31152), .B(n32681), .ZN(n3057) );
  NOR2_X2 U13355 ( .A1(n27617), .A2(n27616), .ZN(n32681) );
  NOR2_X2 U13363 ( .A1(n32790), .A2(n13160), .ZN(n27420) );
  NAND2_X2 U13364 ( .A1(n17446), .A2(n6203), .ZN(n19260) );
  AOI21_X2 U13365 ( .A1(n33116), .A2(n20595), .B(n817), .ZN(n20176) );
  XOR2_X1 U13366 ( .A1(n6812), .A2(n22075), .Z(n21912) );
  OAI21_X2 U13367 ( .A1(n32682), .A2(n27987), .B(n22959), .ZN(n23286) );
  NOR2_X1 U13373 ( .A1(n28877), .A2(n28878), .ZN(n32682) );
  NAND2_X2 U13374 ( .A1(n16607), .A2(n2092), .ZN(n3842) );
  XOR2_X1 U13377 ( .A1(n22192), .A2(n32683), .Z(n526) );
  INV_X1 U13384 ( .I(n25355), .ZN(n32683) );
  INV_X4 U13387 ( .I(n20613), .ZN(n1158) );
  NAND2_X2 U13390 ( .A1(n13954), .A2(n13955), .ZN(n20613) );
  NOR2_X2 U13395 ( .A1(n32684), .A2(n26633), .ZN(n26632) );
  OAI21_X2 U13396 ( .A1(n32671), .A2(n18415), .B(n32685), .ZN(n18421) );
  NAND2_X2 U13397 ( .A1(n33712), .A2(n18419), .ZN(n32685) );
  OAI21_X2 U13406 ( .A1(n32686), .A2(n3163), .B(n28970), .ZN(n30753) );
  INV_X1 U13407 ( .I(n32687), .ZN(n32686) );
  NOR2_X1 U13416 ( .A1(n724), .A2(n13694), .ZN(n32687) );
  INV_X2 U13421 ( .I(n10948), .ZN(n11931) );
  NAND3_X2 U13423 ( .A1(n15287), .A2(n25580), .A3(n25579), .ZN(n10948) );
  NOR2_X1 U13424 ( .A1(n30204), .A2(n11366), .ZN(n15531) );
  NAND2_X2 U13425 ( .A1(n32688), .A2(n9884), .ZN(n21925) );
  XOR2_X1 U13430 ( .A1(n32689), .A2(n17914), .Z(Ciphertext[85]) );
  AOI22_X1 U13431 ( .A1(n27680), .A2(n25268), .B1(n25286), .B2(n25280), .ZN(
        n32689) );
  NAND2_X2 U13434 ( .A1(n33238), .A2(n32690), .ZN(n4184) );
  AND2_X1 U13440 ( .A1(n29620), .A2(n13193), .Z(n32690) );
  INV_X2 U13443 ( .I(n24340), .ZN(n29567) );
  NAND2_X2 U13444 ( .A1(n4460), .A2(n20238), .ZN(n20302) );
  NOR2_X2 U13451 ( .A1(n19847), .A2(n31644), .ZN(n4460) );
  NAND2_X2 U13453 ( .A1(n1878), .A2(n32691), .ZN(n7232) );
  NAND2_X2 U13454 ( .A1(n2694), .A2(n15072), .ZN(n32691) );
  NAND2_X1 U13455 ( .A1(n2694), .A2(n19845), .ZN(n2693) );
  NAND2_X1 U13458 ( .A1(n14486), .A2(n14485), .ZN(n3788) );
  NAND2_X2 U13459 ( .A1(n29780), .A2(n16251), .ZN(n14486) );
  AND2_X1 U13462 ( .A1(n24308), .A2(n11041), .Z(n28428) );
  NAND2_X1 U13463 ( .A1(n32693), .A2(n32692), .ZN(n7942) );
  INV_X1 U13473 ( .I(n1279), .ZN(n32693) );
  NAND2_X2 U13475 ( .A1(n6512), .A2(n24430), .ZN(n25736) );
  NAND4_X2 U13476 ( .A1(n277), .A2(n25627), .A3(n25584), .A4(n17863), .ZN(
        n6512) );
  XOR2_X1 U13478 ( .A1(n32694), .A2(n17564), .Z(n8366) );
  XOR2_X1 U13481 ( .A1(n33509), .A2(n32695), .Z(n32694) );
  OAI21_X2 U13482 ( .A1(n17661), .A2(n11904), .B(n1100), .ZN(n155) );
  XOR2_X1 U13483 ( .A1(n32696), .A2(n22037), .Z(n32947) );
  XOR2_X1 U13484 ( .A1(n4219), .A2(n22283), .Z(n9914) );
  BUF_X2 U13485 ( .I(n31568), .Z(n32697) );
  XOR2_X1 U13492 ( .A1(n12785), .A2(n12789), .Z(n17745) );
  NAND2_X2 U13493 ( .A1(n12787), .A2(n12786), .ZN(n12789) );
  NAND2_X2 U13494 ( .A1(n30215), .A2(n27034), .ZN(n2449) );
  XOR2_X1 U13498 ( .A1(n20753), .A2(n20558), .Z(n11337) );
  XOR2_X1 U13510 ( .A1(n23194), .A2(n32698), .Z(n23197) );
  XOR2_X1 U13515 ( .A1(n23210), .A2(n29719), .Z(n32698) );
  AOI21_X2 U13516 ( .A1(n19236), .A2(n3515), .B(n31139), .ZN(n2280) );
  XOR2_X1 U13524 ( .A1(n32699), .A2(n18001), .Z(n30131) );
  XOR2_X1 U13525 ( .A1(n24427), .A2(n8050), .Z(n32699) );
  OAI22_X2 U13532 ( .A1(n30371), .A2(n18515), .B1(n1188), .B2(n13663), .ZN(
        n6470) );
  XOR2_X1 U13533 ( .A1(n31892), .A2(n32700), .Z(n26930) );
  XOR2_X1 U13534 ( .A1(n23240), .A2(n23238), .Z(n32700) );
  XOR2_X1 U13538 ( .A1(n23389), .A2(n31523), .Z(n23213) );
  OAI21_X2 U13540 ( .A1(n5681), .A2(n23485), .B(n5680), .ZN(n23389) );
  AOI21_X2 U13541 ( .A1(n22714), .A2(n14188), .B(n32701), .ZN(n16160) );
  OAI22_X2 U13542 ( .A1(n15364), .A2(n14188), .B1(n27389), .B2(n22836), .ZN(
        n32701) );
  NAND2_X1 U13548 ( .A1(n16197), .A2(n16198), .ZN(n30081) );
  NAND2_X2 U13549 ( .A1(n32995), .A2(n26501), .ZN(n33971) );
  OAI21_X2 U13550 ( .A1(n28414), .A2(n30869), .B(n20429), .ZN(n10992) );
  XOR2_X1 U13552 ( .A1(n32702), .A2(n16605), .Z(Ciphertext[130]) );
  XOR2_X1 U13553 ( .A1(n24481), .A2(n24482), .Z(n32703) );
  NAND2_X2 U13554 ( .A1(n29539), .A2(n30277), .ZN(n10097) );
  OAI21_X1 U13560 ( .A1(n14020), .A2(n25014), .B(n30461), .ZN(n34043) );
  NAND2_X2 U13561 ( .A1(n3247), .A2(n31645), .ZN(n30314) );
  AOI22_X2 U13562 ( .A1(n32949), .A2(n8886), .B1(n21585), .B2(n3248), .ZN(
        n3247) );
  NOR2_X1 U13566 ( .A1(n33032), .A2(n22873), .ZN(n32704) );
  OAI21_X2 U13569 ( .A1(n22956), .A2(n15601), .B(n22955), .ZN(n27988) );
  INV_X4 U13574 ( .I(n28714), .ZN(n1020) );
  OAI21_X2 U13577 ( .A1(n22825), .A2(n22823), .B(n32705), .ZN(n23467) );
  INV_X2 U13578 ( .I(n13334), .ZN(n719) );
  NAND2_X2 U13580 ( .A1(n15155), .A2(n2378), .ZN(n32950) );
  XOR2_X1 U13582 ( .A1(n7984), .A2(n28746), .Z(n15155) );
  AOI21_X2 U13584 ( .A1(n5555), .A2(n5556), .B(n4306), .ZN(n27104) );
  NAND2_X1 U13587 ( .A1(n13703), .A2(n34058), .ZN(n32706) );
  NAND2_X2 U13594 ( .A1(n23695), .A2(n14078), .ZN(n17578) );
  NAND3_X2 U13596 ( .A1(n17995), .A2(n29081), .A3(n8344), .ZN(n13530) );
  XOR2_X1 U13597 ( .A1(n31055), .A2(n23312), .Z(n6539) );
  XOR2_X1 U13601 ( .A1(n22288), .A2(n22266), .Z(n11816) );
  XOR2_X1 U13602 ( .A1(n33437), .A2(n22044), .Z(n22266) );
  XOR2_X1 U13605 ( .A1(n32707), .A2(n27699), .Z(n2455) );
  XOR2_X1 U13606 ( .A1(n22070), .A2(n457), .Z(n32707) );
  OAI21_X2 U13608 ( .A1(n5095), .A2(n5096), .B(n29621), .ZN(n30870) );
  NAND3_X1 U13613 ( .A1(n10010), .A2(n27092), .A3(n10007), .ZN(Ciphertext[126]) );
  XOR2_X1 U13618 ( .A1(n32708), .A2(n23311), .Z(n10937) );
  XOR2_X1 U13623 ( .A1(n28072), .A2(n15055), .Z(n32708) );
  INV_X2 U13624 ( .I(n25697), .ZN(n1718) );
  NAND2_X2 U13627 ( .A1(n33628), .A2(n33485), .ZN(n3711) );
  XOR2_X1 U13629 ( .A1(n32709), .A2(n16301), .Z(Ciphertext[9]) );
  AOI22_X2 U13632 ( .A1(n8780), .A2(n18219), .B1(n10136), .B2(n24607), .ZN(
        n29532) );
  AOI21_X2 U13633 ( .A1(n24161), .A2(n30595), .B(n3678), .ZN(n31416) );
  OAI21_X2 U13634 ( .A1(n16640), .A2(n12066), .B(n29739), .ZN(n29997) );
  INV_X2 U13639 ( .I(n26385), .ZN(n32711) );
  NAND2_X2 U13640 ( .A1(n33041), .A2(n3255), .ZN(n3253) );
  XOR2_X1 U13641 ( .A1(n32713), .A2(n16680), .Z(Ciphertext[73]) );
  OAI22_X1 U13642 ( .A1(n4613), .A2(n4188), .B1(n25207), .B2(n4614), .ZN(
        n32713) );
  XOR2_X1 U13645 ( .A1(n13480), .A2(n19749), .Z(n15297) );
  NAND2_X2 U13646 ( .A1(n7403), .A2(n7402), .ZN(n13480) );
  INV_X2 U13647 ( .I(n4735), .ZN(n22622) );
  XOR2_X1 U13650 ( .A1(n3812), .A2(n30901), .Z(n4735) );
  INV_X1 U13654 ( .I(n22015), .ZN(n11863) );
  XOR2_X1 U13655 ( .A1(n22015), .A2(n32714), .Z(n14796) );
  NOR2_X2 U13656 ( .A1(n28439), .A2(n9493), .ZN(n22015) );
  NAND2_X2 U13662 ( .A1(n34138), .A2(n32739), .ZN(n12376) );
  NOR2_X2 U13664 ( .A1(n15751), .A2(n4041), .ZN(n10973) );
  NAND2_X2 U13668 ( .A1(n1020), .A2(n17313), .ZN(n15751) );
  NOR2_X2 U13671 ( .A1(n5178), .A2(n11956), .ZN(n30167) );
  NOR2_X2 U13678 ( .A1(n5454), .A2(n24168), .ZN(n15253) );
  NAND2_X2 U13679 ( .A1(n13774), .A2(n8675), .ZN(n24168) );
  XOR2_X1 U13680 ( .A1(n23300), .A2(n23488), .Z(n32715) );
  XOR2_X1 U13681 ( .A1(n30303), .A2(n20924), .Z(n7031) );
  OAI22_X2 U13688 ( .A1(n17228), .A2(n10731), .B1(n15832), .B2(n20516), .ZN(
        n30303) );
  AOI21_X2 U13691 ( .A1(n5556), .A2(n5555), .B(n4306), .ZN(n32877) );
  OAI22_X2 U13692 ( .A1(n31266), .A2(n23892), .B1(n707), .B2(n23715), .ZN(
        n4306) );
  AOI21_X2 U13693 ( .A1(n23111), .A2(n1264), .B(n16254), .ZN(n32716) );
  OR2_X1 U13699 ( .A1(n13176), .A2(n24216), .Z(n10179) );
  INV_X2 U13700 ( .I(n24998), .ZN(n31122) );
  NAND2_X2 U13702 ( .A1(n25003), .A2(n2983), .ZN(n24998) );
  XOR2_X1 U13703 ( .A1(n29740), .A2(n22247), .Z(n22340) );
  NAND2_X2 U13704 ( .A1(n30745), .A2(n29799), .ZN(n28181) );
  AND2_X1 U13707 ( .A1(n15772), .A2(n8140), .Z(n4668) );
  NOR2_X2 U13708 ( .A1(n15883), .A2(n32717), .ZN(n25479) );
  INV_X2 U13712 ( .I(n24193), .ZN(n13040) );
  NAND2_X2 U13713 ( .A1(n3484), .A2(n31623), .ZN(n24193) );
  OAI21_X2 U13718 ( .A1(n22842), .A2(n22843), .B(n23482), .ZN(n22845) );
  NAND2_X1 U13724 ( .A1(n33938), .A2(n22626), .ZN(n6010) );
  NOR3_X1 U13725 ( .A1(n33102), .A2(n2480), .A3(n25509), .ZN(n25511) );
  NOR2_X2 U13727 ( .A1(n32719), .A2(n32718), .ZN(n17328) );
  NAND2_X2 U13730 ( .A1(n13570), .A2(n13571), .ZN(n32718) );
  NAND3_X2 U13732 ( .A1(n32720), .A2(n32849), .A3(n19294), .ZN(n7251) );
  NOR2_X2 U13733 ( .A1(n3181), .A2(n8125), .ZN(n31797) );
  NAND3_X2 U13734 ( .A1(n3166), .A2(n23835), .A3(n28497), .ZN(n8125) );
  XOR2_X1 U13735 ( .A1(n20852), .A2(n18102), .Z(n6758) );
  NOR2_X1 U13738 ( .A1(n11985), .A2(n11548), .ZN(n15738) );
  NAND2_X2 U13743 ( .A1(n17816), .A2(n32721), .ZN(n6911) );
  NOR2_X2 U13745 ( .A1(n16862), .A2(n10749), .ZN(n32721) );
  XOR2_X1 U13747 ( .A1(n26045), .A2(n24574), .Z(n32722) );
  NAND2_X1 U13750 ( .A1(n8200), .A2(n8201), .ZN(n22620) );
  NOR2_X2 U13753 ( .A1(n5451), .A2(n5449), .ZN(n33329) );
  XOR2_X1 U13757 ( .A1(n26084), .A2(n19556), .Z(n18065) );
  NAND3_X2 U13758 ( .A1(n2371), .A2(n2664), .A3(n32808), .ZN(n31197) );
  OR2_X1 U13768 ( .A1(n3860), .A2(n33722), .Z(n23566) );
  OAI22_X1 U13774 ( .A1(n5583), .A2(n33714), .B1(n26130), .B2(n13969), .ZN(
        n32723) );
  NAND3_X2 U13775 ( .A1(n25262), .A2(n25263), .A3(n6280), .ZN(n30281) );
  OAI22_X2 U13778 ( .A1(n1207), .A2(n12431), .B1(n16291), .B2(n25278), .ZN(
        n25286) );
  NOR2_X1 U13781 ( .A1(n13720), .A2(n29472), .ZN(n7475) );
  NOR2_X2 U13785 ( .A1(n10202), .A2(n11378), .ZN(n3186) );
  NAND2_X2 U13788 ( .A1(n31813), .A2(n24317), .ZN(n32725) );
  XOR2_X1 U13800 ( .A1(n32726), .A2(n6737), .Z(n6735) );
  XOR2_X1 U13801 ( .A1(n31900), .A2(n14060), .Z(n19967) );
  NAND4_X2 U13803 ( .A1(n30886), .A2(n12883), .A3(n12884), .A4(n13721), .ZN(
        n16940) );
  OAI21_X2 U13806 ( .A1(n10247), .A2(n11269), .B(n32727), .ZN(n10228) );
  AOI22_X2 U13807 ( .A1(n17190), .A2(n1439), .B1(n18634), .B2(n15888), .ZN(
        n32727) );
  XOR2_X1 U13809 ( .A1(n28640), .A2(n6420), .Z(n10954) );
  INV_X1 U13810 ( .I(n33846), .ZN(n29437) );
  OR2_X1 U13812 ( .A1(n33846), .A2(n19267), .Z(n15759) );
  XOR2_X1 U13813 ( .A1(n32728), .A2(n33699), .Z(n27790) );
  XOR2_X1 U13816 ( .A1(n27791), .A2(n12), .Z(n32728) );
  INV_X4 U13817 ( .I(n16966), .ZN(n32746) );
  NAND3_X2 U13818 ( .A1(n32729), .A2(n29431), .A3(n3065), .ZN(n12748) );
  NAND2_X1 U13820 ( .A1(n3069), .A2(n3068), .ZN(n32729) );
  XOR2_X1 U13832 ( .A1(n32730), .A2(n25364), .Z(Ciphertext[99]) );
  NAND2_X2 U13833 ( .A1(n34096), .A2(n14308), .ZN(n22127) );
  NAND2_X2 U13834 ( .A1(n21492), .A2(n21566), .ZN(n33644) );
  NAND2_X2 U13835 ( .A1(n987), .A2(n5035), .ZN(n16202) );
  NOR2_X1 U13840 ( .A1(n13295), .A2(n8606), .ZN(n15628) );
  NOR2_X2 U13841 ( .A1(n17515), .A2(n13565), .ZN(n13295) );
  XOR2_X1 U13843 ( .A1(n5884), .A2(n5885), .Z(n28545) );
  AND3_X1 U13844 ( .A1(n14255), .A2(n32170), .A3(n14133), .Z(n27893) );
  XOR2_X1 U13845 ( .A1(n11862), .A2(n14952), .Z(n22252) );
  NOR2_X2 U13850 ( .A1(n28413), .A2(n30374), .ZN(n11862) );
  XOR2_X1 U13851 ( .A1(n20688), .A2(n11512), .Z(n11514) );
  NAND3_X2 U13852 ( .A1(n24137), .A2(n15011), .A3(n6980), .ZN(n33123) );
  INV_X4 U13854 ( .I(n16286), .ZN(n9561) );
  OAI22_X2 U13856 ( .A1(n3825), .A2(n4308), .B1(n18236), .B2(n20111), .ZN(
        n20560) );
  NAND2_X2 U13857 ( .A1(n32731), .A2(n31146), .ZN(n3489) );
  XOR2_X1 U13861 ( .A1(n23145), .A2(n23280), .Z(n6388) );
  XOR2_X1 U13862 ( .A1(n2072), .A2(n32732), .Z(n2074) );
  XOR2_X1 U13866 ( .A1(n32733), .A2(n19470), .Z(n32732) );
  INV_X2 U13867 ( .I(n4321), .ZN(n32733) );
  XOR2_X1 U13869 ( .A1(n9848), .A2(n13745), .Z(n13743) );
  XOR2_X1 U13870 ( .A1(n24675), .A2(n3694), .Z(n9848) );
  BUF_X4 U13873 ( .I(n11676), .Z(n29218) );
  NAND2_X2 U13875 ( .A1(n28652), .A2(n32734), .ZN(n14681) );
  NAND2_X1 U13876 ( .A1(n15113), .A2(n15112), .ZN(n32734) );
  OAI21_X2 U13877 ( .A1(n32735), .A2(n14021), .B(n5624), .ZN(n2983) );
  AND2_X1 U13878 ( .A1(n16305), .A2(n11845), .Z(n24318) );
  INV_X4 U13880 ( .I(n5741), .ZN(n1243) );
  NAND2_X2 U13881 ( .A1(n33789), .A2(n33788), .ZN(n34164) );
  NAND2_X2 U13883 ( .A1(n21559), .A2(n6544), .ZN(n21852) );
  OR2_X1 U13884 ( .A1(n30832), .A2(n7811), .Z(n15494) );
  NOR3_X2 U13886 ( .A1(n33730), .A2(n1347), .A3(n3084), .ZN(n2086) );
  XOR2_X1 U13888 ( .A1(n13833), .A2(n22224), .Z(n13862) );
  NOR2_X2 U13889 ( .A1(n15458), .A2(n32736), .ZN(n28081) );
  NOR2_X1 U13895 ( .A1(n31490), .A2(n1718), .ZN(n32736) );
  AOI22_X2 U13897 ( .A1(n33779), .A2(n12452), .B1(n26439), .B2(n21672), .ZN(
        n11991) );
  NOR2_X1 U13900 ( .A1(n32888), .A2(n12040), .ZN(n12085) );
  XOR2_X1 U13901 ( .A1(n34126), .A2(n14985), .Z(n12040) );
  INV_X4 U13906 ( .I(n8057), .ZN(n20238) );
  NAND2_X2 U13908 ( .A1(n31062), .A2(n30790), .ZN(n8057) );
  NOR2_X1 U13913 ( .A1(n33031), .A2(n8733), .ZN(n30965) );
  NAND2_X2 U13917 ( .A1(n18976), .A2(n14892), .ZN(n1807) );
  NOR2_X2 U13918 ( .A1(n17131), .A2(n17130), .ZN(n14892) );
  OAI22_X2 U13919 ( .A1(n33748), .A2(n5040), .B1(n976), .B2(n4675), .ZN(n28945) );
  OAI22_X2 U13921 ( .A1(n20949), .A2(n5822), .B1(n16633), .B2(n21239), .ZN(
        n2888) );
  NAND2_X2 U13922 ( .A1(n2888), .A2(n17699), .ZN(n33859) );
  BUF_X2 U13923 ( .I(n24226), .Z(n32737) );
  NAND2_X2 U13924 ( .A1(n25187), .A2(n25234), .ZN(n13074) );
  INV_X2 U13925 ( .I(n32738), .ZN(n33621) );
  XNOR2_X1 U13932 ( .A1(n18364), .A2(Key[48]), .ZN(n32738) );
  NAND2_X1 U13947 ( .A1(n9876), .A2(n20010), .ZN(n19789) );
  INV_X2 U13948 ( .I(n10679), .ZN(n12323) );
  NOR2_X1 U13950 ( .A1(n3760), .A2(n33953), .ZN(n16430) );
  XOR2_X1 U13959 ( .A1(n9230), .A2(n14766), .Z(n27571) );
  XOR2_X1 U13960 ( .A1(n29262), .A2(n5875), .Z(n4087) );
  XOR2_X1 U13962 ( .A1(n22030), .A2(n27837), .Z(n29262) );
  NOR2_X1 U13963 ( .A1(n19907), .A2(n19958), .ZN(n29284) );
  AOI22_X2 U13965 ( .A1(n19996), .A2(n34108), .B1(n6263), .B2(n1957), .ZN(
        n1956) );
  INV_X2 U13966 ( .I(n17299), .ZN(n783) );
  XNOR2_X1 U13970 ( .A1(n17300), .A2(n19482), .ZN(n17299) );
  NAND2_X2 U13972 ( .A1(n32740), .A2(n19535), .ZN(n20401) );
  AOI21_X1 U13981 ( .A1(n14365), .A2(n3944), .B(n20509), .ZN(n19841) );
  INV_X2 U13986 ( .I(n15282), .ZN(n20509) );
  AOI21_X2 U13987 ( .A1(n19832), .A2(n8406), .B(n19831), .ZN(n15282) );
  AOI21_X2 U13988 ( .A1(n27501), .A2(n738), .B(n9934), .ZN(n14690) );
  NAND2_X2 U13989 ( .A1(n3748), .A2(n24120), .ZN(n10427) );
  OR2_X2 U13992 ( .A1(n2978), .A2(n33482), .Z(n9852) );
  XOR2_X1 U13994 ( .A1(n24492), .A2(n24693), .Z(n15862) );
  XOR2_X1 U14000 ( .A1(n15671), .A2(n15508), .Z(n24492) );
  INV_X2 U14003 ( .I(n27127), .ZN(n1079) );
  INV_X2 U14005 ( .I(n25277), .ZN(n25284) );
  NAND3_X2 U14007 ( .A1(n24588), .A2(n10330), .A3(n24585), .ZN(n25277) );
  NOR2_X1 U14009 ( .A1(n18874), .A2(n9909), .ZN(n14666) );
  NAND2_X1 U14010 ( .A1(n32938), .A2(n33803), .ZN(n23730) );
  NAND3_X2 U14012 ( .A1(n11629), .A2(n33046), .A3(n2066), .ZN(n22415) );
  OR2_X1 U14013 ( .A1(n9931), .A2(n7663), .Z(n33560) );
  NOR3_X1 U14019 ( .A1(n31702), .A2(n30783), .A3(n21086), .ZN(n32741) );
  NOR2_X2 U14026 ( .A1(n27687), .A2(n30271), .ZN(n18472) );
  NOR2_X2 U14027 ( .A1(n4225), .A2(n8285), .ZN(n21044) );
  XOR2_X1 U14034 ( .A1(n32742), .A2(n23213), .Z(n284) );
  XOR2_X1 U14036 ( .A1(n102), .A2(n27763), .Z(n32742) );
  AOI22_X2 U14041 ( .A1(n32743), .A2(n28867), .B1(n5178), .B2(n5177), .ZN(
        n26767) );
  NOR2_X2 U14042 ( .A1(n5178), .A2(n28330), .ZN(n32743) );
  NOR2_X2 U14046 ( .A1(n20038), .A2(n20135), .ZN(n19964) );
  NAND2_X2 U14048 ( .A1(n27911), .A2(n20037), .ZN(n20038) );
  XOR2_X1 U14049 ( .A1(n7636), .A2(n7634), .Z(n33856) );
  XOR2_X1 U14053 ( .A1(n19586), .A2(n11817), .Z(n7636) );
  NOR2_X2 U14055 ( .A1(n20453), .A2(n20454), .ZN(n16959) );
  NAND2_X2 U14056 ( .A1(n15176), .A2(n15177), .ZN(n20453) );
  XOR2_X1 U14057 ( .A1(n12376), .A2(n1917), .Z(n17128) );
  XOR2_X1 U14064 ( .A1(n8949), .A2(n24837), .Z(n15308) );
  NOR2_X2 U14066 ( .A1(n10793), .A2(n24172), .ZN(n8949) );
  XOR2_X1 U14067 ( .A1(n20983), .A2(n20686), .Z(n15526) );
  NAND2_X1 U14070 ( .A1(n8927), .A2(n15602), .ZN(n11770) );
  AND2_X1 U14072 ( .A1(n21253), .A2(n21233), .Z(n33263) );
  NAND2_X2 U14073 ( .A1(n12658), .A2(n23901), .ZN(n31275) );
  AOI22_X2 U14076 ( .A1(n26257), .A2(n16959), .B1(n28527), .B2(n20362), .ZN(
        n28332) );
  NAND2_X2 U14080 ( .A1(n31960), .A2(n11755), .ZN(n10775) );
  NAND2_X2 U14083 ( .A1(n22358), .A2(n22357), .ZN(n22986) );
  NAND2_X2 U14085 ( .A1(n22510), .A2(n8199), .ZN(n22358) );
  XOR2_X1 U14088 ( .A1(n32744), .A2(n1421), .Z(Ciphertext[150]) );
  AOI22_X1 U14090 ( .A1(n1076), .A2(n9552), .B1(n4253), .B2(n9495), .ZN(n32744) );
  INV_X2 U14099 ( .I(n245), .ZN(n32745) );
  NOR2_X1 U14100 ( .A1(n6118), .A2(n18795), .ZN(n8315) );
  XOR2_X1 U14101 ( .A1(n24455), .A2(n24788), .Z(n391) );
  XOR2_X1 U14103 ( .A1(n24790), .A2(n24512), .Z(n24455) );
  XOR2_X1 U14106 ( .A1(n23506), .A2(n23504), .Z(n2024) );
  XOR2_X1 U14110 ( .A1(n4400), .A2(n14293), .Z(n19537) );
  NOR2_X2 U14114 ( .A1(n19250), .A2(n19251), .ZN(n4400) );
  NAND2_X2 U14117 ( .A1(n32748), .A2(n5045), .ZN(n23792) );
  OAI21_X2 U14118 ( .A1(n1973), .A2(n3748), .B(n5335), .ZN(n32748) );
  BUF_X2 U14123 ( .I(n27931), .Z(n32750) );
  OAI21_X1 U14131 ( .A1(n21854), .A2(n21559), .B(n4356), .ZN(n5264) );
  NAND2_X2 U14132 ( .A1(n6878), .A2(n6880), .ZN(n4356) );
  NOR2_X2 U14134 ( .A1(n8671), .A2(n32751), .ZN(n14331) );
  NAND3_X2 U14136 ( .A1(n15696), .A2(n18074), .A3(n9512), .ZN(n32751) );
  NAND2_X2 U14142 ( .A1(n27139), .A2(n17746), .ZN(n3487) );
  AOI22_X2 U14144 ( .A1(n9660), .A2(n937), .B1(n13423), .B2(n29283), .ZN(
        n17746) );
  OAI21_X2 U14146 ( .A1(n32752), .A2(n31167), .B(n29738), .ZN(n19325) );
  NOR2_X2 U14148 ( .A1(n9289), .A2(n18671), .ZN(n32752) );
  XOR2_X1 U14150 ( .A1(n14645), .A2(n27167), .Z(n3235) );
  NOR2_X2 U14153 ( .A1(n1997), .A2(n1995), .ZN(n27167) );
  AOI22_X2 U14154 ( .A1(n26301), .A2(n9913), .B1(n13143), .B2(n11917), .ZN(
        n32754) );
  BUF_X4 U14156 ( .I(n21867), .Z(n30152) );
  XOR2_X1 U14158 ( .A1(n32755), .A2(n24503), .Z(n16659) );
  XOR2_X1 U14159 ( .A1(n10632), .A2(n24241), .Z(n32755) );
  NAND2_X2 U14160 ( .A1(n22613), .A2(n32756), .ZN(n16022) );
  AOI21_X2 U14165 ( .A1(n32045), .A2(n26173), .B(n32757), .ZN(n32756) );
  XOR2_X1 U14175 ( .A1(n13695), .A2(n24479), .Z(n14499) );
  NAND2_X2 U14176 ( .A1(n9398), .A2(n9933), .ZN(n13695) );
  NOR2_X2 U14178 ( .A1(n20312), .A2(n26566), .ZN(n20480) );
  XOR2_X1 U14182 ( .A1(n12972), .A2(n18929), .Z(n10861) );
  XOR2_X1 U14185 ( .A1(n2162), .A2(n2161), .Z(n2655) );
  XOR2_X1 U14186 ( .A1(n22220), .A2(n8617), .Z(n13020) );
  OAI21_X2 U14191 ( .A1(n16371), .A2(n8618), .B(n21739), .ZN(n22220) );
  NAND3_X2 U14193 ( .A1(n16962), .A2(n22415), .A3(n22416), .ZN(n15456) );
  NAND2_X2 U14197 ( .A1(n6380), .A2(n31428), .ZN(n34065) );
  XOR2_X1 U14198 ( .A1(n20869), .A2(n25457), .Z(n2055) );
  NAND2_X2 U14201 ( .A1(n26632), .A2(n13000), .ZN(n20869) );
  NAND2_X2 U14205 ( .A1(n20312), .A2(n20577), .ZN(n20243) );
  AOI22_X1 U14209 ( .A1(n6807), .A2(n29234), .B1(n32800), .B2(n27532), .ZN(
        n14308) );
  NOR2_X2 U14210 ( .A1(n21636), .A2(n21634), .ZN(n32800) );
  INV_X2 U14211 ( .I(n28950), .ZN(n32760) );
  NAND2_X2 U14215 ( .A1(n10), .A2(n32762), .ZN(n14342) );
  NAND3_X2 U14216 ( .A1(n14346), .A2(n18637), .A3(n14651), .ZN(n32762) );
  AOI21_X2 U14218 ( .A1(n28671), .A2(n23760), .B(n23756), .ZN(n4026) );
  NAND2_X2 U14221 ( .A1(n33837), .A2(n32763), .ZN(n18974) );
  XNOR2_X1 U14223 ( .A1(n29042), .A2(n20747), .ZN(n20958) );
  NAND2_X2 U14226 ( .A1(n183), .A2(n7956), .ZN(n20747) );
  AOI21_X2 U14227 ( .A1(n13104), .A2(n13105), .B(n22112), .ZN(n22894) );
  AOI22_X2 U14230 ( .A1(n32764), .A2(n27386), .B1(n13943), .B2(n20358), .ZN(
        n20963) );
  OR2_X1 U14234 ( .A1(n7762), .A2(n27600), .Z(n32765) );
  NAND2_X2 U14235 ( .A1(n8968), .A2(n24109), .ZN(n28253) );
  INV_X1 U14239 ( .I(n13063), .ZN(n32766) );
  NAND2_X1 U14240 ( .A1(n33023), .A2(n32766), .ZN(n5092) );
  XOR2_X1 U14246 ( .A1(n32767), .A2(n33877), .Z(n14439) );
  XOR2_X1 U14248 ( .A1(n6218), .A2(n6808), .Z(n32767) );
  NAND2_X1 U14250 ( .A1(n33657), .A2(n2911), .ZN(n33656) );
  OAI22_X2 U14258 ( .A1(n21453), .A2(n1143), .B1(n9186), .B2(n21237), .ZN(
        n33586) );
  INV_X2 U14259 ( .I(n32768), .ZN(n29882) );
  XOR2_X1 U14260 ( .A1(n2054), .A2(n2053), .Z(n32768) );
  AOI21_X2 U14261 ( .A1(n32769), .A2(n33324), .B(n15984), .ZN(n19021) );
  INV_X2 U14265 ( .I(n9810), .ZN(n9440) );
  XOR2_X1 U14267 ( .A1(n22306), .A2(n9809), .Z(n9810) );
  NOR2_X1 U14268 ( .A1(n10018), .A2(n3004), .ZN(n2560) );
  NAND2_X2 U14269 ( .A1(n5795), .A2(n21721), .ZN(n21806) );
  NAND3_X2 U14270 ( .A1(n3936), .A2(n10555), .A3(n4179), .ZN(n5795) );
  NOR2_X2 U14275 ( .A1(n16637), .A2(n1042), .ZN(n19903) );
  OR2_X1 U14277 ( .A1(n10312), .A2(n8057), .Z(n19864) );
  XOR2_X1 U14278 ( .A1(n24812), .A2(n32770), .Z(n26365) );
  XOR2_X1 U14281 ( .A1(n9650), .A2(n24811), .Z(n32770) );
  NAND3_X2 U14282 ( .A1(n21187), .A2(n17640), .A3(n34131), .ZN(n21083) );
  NAND2_X2 U14285 ( .A1(n5394), .A2(n5395), .ZN(n21187) );
  OAI21_X2 U14286 ( .A1(n33030), .A2(n14276), .B(n16728), .ZN(n14274) );
  OR2_X1 U14290 ( .A1(n31969), .A2(n10312), .Z(n31338) );
  XOR2_X1 U14295 ( .A1(n29624), .A2(n14340), .Z(n21232) );
  AOI21_X2 U14297 ( .A1(n29695), .A2(n20489), .B(n20487), .ZN(n17512) );
  NOR2_X2 U14301 ( .A1(n13015), .A2(n13845), .ZN(n12648) );
  XOR2_X1 U14303 ( .A1(n19642), .A2(n32058), .Z(n582) );
  XOR2_X1 U14308 ( .A1(n32772), .A2(n15679), .Z(n32915) );
  XOR2_X1 U14310 ( .A1(n17220), .A2(n32044), .Z(n32772) );
  XOR2_X1 U14311 ( .A1(n19710), .A2(n19408), .Z(n15913) );
  NOR2_X1 U14312 ( .A1(n12932), .A2(n9146), .ZN(n27309) );
  NOR2_X2 U14313 ( .A1(n17329), .A2(n4647), .ZN(n15045) );
  OAI21_X1 U14317 ( .A1(n22413), .A2(n14160), .B(n22486), .ZN(n14010) );
  XOR2_X1 U14320 ( .A1(n12934), .A2(n23435), .Z(n23155) );
  XOR2_X1 U14321 ( .A1(n24554), .A2(n24556), .Z(n1690) );
  XOR2_X1 U14334 ( .A1(n24846), .A2(n24741), .Z(n24554) );
  INV_X2 U14335 ( .I(n25345), .ZN(n14246) );
  NAND2_X2 U14339 ( .A1(n18958), .A2(n18621), .ZN(n18962) );
  XOR2_X1 U14343 ( .A1(n21012), .A2(n21011), .Z(n7015) );
  XOR2_X1 U14354 ( .A1(n15293), .A2(n13930), .Z(n30734) );
  NAND2_X2 U14359 ( .A1(n29464), .A2(n10349), .ZN(n15293) );
  NAND2_X2 U14360 ( .A1(n5428), .A2(n32773), .ZN(n8335) );
  OAI21_X2 U14361 ( .A1(n18750), .A2(n13243), .B(n959), .ZN(n32773) );
  NAND3_X2 U14362 ( .A1(n23002), .A2(n22831), .A3(n13159), .ZN(n12157) );
  XOR2_X1 U14368 ( .A1(n1994), .A2(n28601), .Z(n6913) );
  XOR2_X1 U14369 ( .A1(n32774), .A2(n590), .Z(n21053) );
  XOR2_X1 U14370 ( .A1(n21026), .A2(n20855), .Z(n32774) );
  AOI22_X2 U14375 ( .A1(n32775), .A2(n8183), .B1(n20060), .B2(n16789), .ZN(
        n29914) );
  INV_X1 U14378 ( .I(n4327), .ZN(n32776) );
  NAND2_X1 U14384 ( .A1(n27955), .A2(n21396), .ZN(n32778) );
  NAND2_X2 U14386 ( .A1(n9677), .A2(n10228), .ZN(n11798) );
  NAND2_X2 U14400 ( .A1(n30246), .A2(n32779), .ZN(n7182) );
  NAND2_X1 U14401 ( .A1(n3888), .A2(n3889), .ZN(n32779) );
  BUF_X2 U14402 ( .I(n20080), .Z(n32780) );
  OAI21_X2 U14405 ( .A1(n31463), .A2(n31464), .B(n25872), .ZN(n13053) );
  INV_X2 U14408 ( .I(n32781), .ZN(n29444) );
  NAND2_X2 U14413 ( .A1(n14054), .A2(n8130), .ZN(n32781) );
  XOR2_X1 U14416 ( .A1(n32782), .A2(n25856), .Z(Ciphertext[177]) );
  XOR2_X1 U14422 ( .A1(n32783), .A2(n465), .Z(n6420) );
  XOR2_X1 U14424 ( .A1(n30524), .A2(n16373), .Z(n32783) );
  INV_X2 U14427 ( .I(n28278), .ZN(n1322) );
  INV_X2 U14428 ( .I(n32784), .ZN(n18920) );
  NAND3_X2 U14430 ( .A1(n18833), .A2(n32786), .A3(n32785), .ZN(n32784) );
  NOR3_X1 U14434 ( .A1(n27262), .A2(n1202), .A3(n32856), .ZN(n27528) );
  OR2_X1 U14436 ( .A1(n16606), .A2(n20566), .Z(n33937) );
  OR3_X1 U14437 ( .A1(n28430), .A2(n20008), .A3(n29882), .Z(n1873) );
  XOR2_X1 U14443 ( .A1(n9507), .A2(n20976), .Z(n2812) );
  INV_X2 U14450 ( .I(n15516), .ZN(n9507) );
  XOR2_X1 U14453 ( .A1(n21009), .A2(n20873), .Z(n15516) );
  NAND2_X2 U14455 ( .A1(n32789), .A2(n3780), .ZN(n18028) );
  BUF_X2 U14461 ( .I(n33373), .Z(n32791) );
  NAND2_X2 U14463 ( .A1(n32792), .A2(n16978), .ZN(n20565) );
  NAND2_X2 U14472 ( .A1(n32793), .A2(n18270), .ZN(n21028) );
  OAI22_X2 U14474 ( .A1(n27901), .A2(n27902), .B1(n8819), .B2(n12999), .ZN(
        n32793) );
  NAND2_X2 U14476 ( .A1(n32794), .A2(n13106), .ZN(n3055) );
  NAND2_X2 U14477 ( .A1(n3057), .A2(n5139), .ZN(n13106) );
  OR2_X1 U14482 ( .A1(n3060), .A2(n3059), .Z(n32794) );
  XOR2_X1 U14486 ( .A1(n33427), .A2(n1540), .Z(n11720) );
  XOR2_X1 U14495 ( .A1(n20889), .A2(n32795), .Z(n27000) );
  XOR2_X1 U14496 ( .A1(n10159), .A2(n32796), .Z(n32795) );
  XOR2_X1 U14499 ( .A1(n28587), .A2(n15424), .Z(n27234) );
  NAND2_X2 U14501 ( .A1(n7881), .A2(n23065), .ZN(n22827) );
  NOR3_X2 U14503 ( .A1(n29455), .A2(n31073), .A3(n16722), .ZN(n21913) );
  NOR2_X1 U14505 ( .A1(n7993), .A2(n28329), .ZN(n5678) );
  NOR2_X1 U14506 ( .A1(n1773), .A2(n22551), .ZN(n22314) );
  NAND3_X2 U14509 ( .A1(n24233), .A2(n1634), .A3(n24236), .ZN(n23699) );
  XOR2_X1 U14512 ( .A1(n29137), .A2(n9412), .Z(n17395) );
  AOI22_X2 U14518 ( .A1(n1771), .A2(n1770), .B1(n1769), .B2(n2551), .ZN(n9412)
         );
  XOR2_X1 U14523 ( .A1(n20743), .A2(n1545), .Z(n7431) );
  XOR2_X1 U14524 ( .A1(n3009), .A2(n21047), .Z(n20743) );
  OAI22_X2 U14525 ( .A1(n20288), .A2(n10351), .B1(n20324), .B2(n20519), .ZN(
        n7255) );
  XOR2_X1 U14529 ( .A1(n9701), .A2(n33678), .Z(n22597) );
  BUF_X4 U14532 ( .I(n18655), .Z(n17843) );
  AND2_X1 U14538 ( .A1(n10847), .A2(n8870), .Z(n30004) );
  XOR2_X1 U14548 ( .A1(n18100), .A2(n22191), .Z(n6515) );
  NAND2_X2 U14551 ( .A1(n11359), .A2(n11728), .ZN(n22191) );
  BUF_X2 U14556 ( .I(n32069), .Z(n32799) );
  NAND2_X2 U14557 ( .A1(n22497), .A2(n16306), .ZN(n33010) );
  OAI22_X2 U14560 ( .A1(n22762), .A2(n22715), .B1(n22694), .B2(n851), .ZN(
        n33008) );
  XOR2_X1 U14565 ( .A1(n17369), .A2(n16429), .Z(n18929) );
  OR2_X1 U14566 ( .A1(n18098), .A2(n22476), .Z(n30384) );
  XOR2_X1 U14568 ( .A1(n14215), .A2(n19475), .Z(n11092) );
  XOR2_X1 U14570 ( .A1(n14214), .A2(n19367), .Z(n14215) );
  OAI22_X2 U14573 ( .A1(n12509), .A2(n32801), .B1(n23448), .B2(n28210), .ZN(
        n16215) );
  BUF_X2 U14575 ( .I(n19325), .Z(n32802) );
  INV_X2 U14581 ( .I(n32803), .ZN(n4145) );
  XOR2_X1 U14588 ( .A1(n33916), .A2(n1704), .Z(n32803) );
  XOR2_X1 U14589 ( .A1(n32804), .A2(n19575), .Z(n13305) );
  XOR2_X1 U14593 ( .A1(n26617), .A2(n8633), .Z(n32804) );
  XOR2_X1 U14602 ( .A1(n17351), .A2(n17350), .Z(n33152) );
  XOR2_X1 U14603 ( .A1(n4728), .A2(n31843), .Z(n5523) );
  NAND2_X2 U14604 ( .A1(n11266), .A2(n11265), .ZN(n21559) );
  NAND2_X2 U14605 ( .A1(n2355), .A2(n33664), .ZN(n22283) );
  OAI21_X2 U14606 ( .A1(n375), .A2(n29040), .B(n20092), .ZN(n31280) );
  NAND2_X2 U14608 ( .A1(n33286), .A2(n9691), .ZN(n14639) );
  XOR2_X1 U14610 ( .A1(n26255), .A2(n11636), .Z(n31575) );
  XOR2_X1 U14611 ( .A1(n33111), .A2(n23219), .Z(n15487) );
  XOR2_X1 U14612 ( .A1(n20912), .A2(n7458), .Z(n26954) );
  XOR2_X1 U14615 ( .A1(n8997), .A2(n20781), .Z(n7458) );
  NOR3_X2 U14616 ( .A1(n33985), .A2(n4117), .A3(n7349), .ZN(n7348) );
  XOR2_X1 U14622 ( .A1(n29936), .A2(n30676), .Z(n13427) );
  XOR2_X1 U14627 ( .A1(n21027), .A2(n21026), .Z(n12272) );
  NAND2_X2 U14632 ( .A1(n7007), .A2(n28190), .ZN(n10149) );
  AND2_X1 U14638 ( .A1(n25891), .A2(n25890), .Z(n33473) );
  NAND2_X2 U14640 ( .A1(n32806), .A2(n15631), .ZN(n7868) );
  OAI21_X2 U14642 ( .A1(n30694), .A2(n10483), .B(n926), .ZN(n32806) );
  NOR2_X2 U14644 ( .A1(n32108), .A2(n33621), .ZN(n18800) );
  OR2_X1 U14646 ( .A1(n17131), .A2(n17130), .Z(n28361) );
  OAI22_X2 U14648 ( .A1(n11049), .A2(n23608), .B1(n24285), .B2(n17068), .ZN(
        n27793) );
  XOR2_X1 U14649 ( .A1(n14762), .A2(n24826), .Z(n24808) );
  NAND2_X2 U14650 ( .A1(n29924), .A2(n2401), .ZN(n14762) );
  NAND2_X2 U14656 ( .A1(n2036), .A2(n32843), .ZN(n27931) );
  OAI22_X2 U14664 ( .A1(n33567), .A2(n33568), .B1(n9945), .B2(n10416), .ZN(
        n12720) );
  NAND2_X1 U14666 ( .A1(n11379), .A2(n14898), .ZN(n3436) );
  NAND2_X1 U14668 ( .A1(n26330), .A2(n22634), .ZN(n22612) );
  NOR2_X1 U14669 ( .A1(n33283), .A2(n858), .ZN(n33282) );
  NAND2_X1 U14675 ( .A1(n33282), .A2(n33280), .ZN(n33901) );
  NAND2_X2 U14681 ( .A1(n12358), .A2(n25890), .ZN(n30019) );
  XOR2_X1 U14684 ( .A1(n3576), .A2(n3574), .Z(n18182) );
  XOR2_X1 U14685 ( .A1(n32810), .A2(n24553), .Z(n9189) );
  OAI21_X2 U14688 ( .A1(n18127), .A2(n18128), .B(n24227), .ZN(n24553) );
  INV_X2 U14690 ( .I(n24847), .ZN(n32810) );
  BUF_X4 U14692 ( .I(n15296), .Z(n29180) );
  OAI22_X2 U14702 ( .A1(n32601), .A2(n25205), .B1(n13273), .B2(n25239), .ZN(
        n33494) );
  NAND2_X1 U14706 ( .A1(n10287), .A2(n33566), .ZN(n4341) );
  XOR2_X1 U14710 ( .A1(n12272), .A2(n21032), .Z(n33566) );
  NAND2_X2 U14711 ( .A1(n21674), .A2(n16345), .ZN(n28111) );
  NAND2_X2 U14713 ( .A1(n33810), .A2(n21604), .ZN(n21674) );
  XOR2_X1 U14719 ( .A1(n31486), .A2(n32811), .Z(n28107) );
  XOR2_X1 U14720 ( .A1(n30628), .A2(n21996), .Z(n32811) );
  XOR2_X1 U14724 ( .A1(n7107), .A2(n32812), .Z(n31737) );
  XOR2_X1 U14725 ( .A1(n34100), .A2(n32813), .Z(n32812) );
  INV_X1 U14728 ( .I(n25541), .ZN(n32813) );
  NOR2_X2 U14733 ( .A1(n25165), .A2(n25175), .ZN(n25173) );
  CLKBUF_X8 U14735 ( .I(n13473), .Z(n33007) );
  NAND2_X2 U14739 ( .A1(n29043), .A2(n8125), .ZN(n421) );
  XOR2_X1 U14740 ( .A1(n8067), .A2(n8065), .Z(n9490) );
  NAND3_X2 U14743 ( .A1(n31933), .A2(n1117), .A3(n7561), .ZN(n27856) );
  NAND3_X2 U14751 ( .A1(n17532), .A2(n20489), .A3(n4254), .ZN(n7799) );
  OR2_X1 U14753 ( .A1(n19101), .A2(n18923), .Z(n17444) );
  NOR2_X1 U14754 ( .A1(n10103), .A2(n10104), .ZN(n33601) );
  BUF_X2 U14763 ( .I(n13286), .Z(n32816) );
  NAND2_X2 U14768 ( .A1(n14959), .A2(n25013), .ZN(n14846) );
  NAND2_X2 U14774 ( .A1(n15277), .A2(n14799), .ZN(n33288) );
  XOR2_X1 U14776 ( .A1(n32817), .A2(n1198), .Z(Ciphertext[138]) );
  AOI22_X1 U14778 ( .A1(n28631), .A2(n11212), .B1(n9365), .B2(n734), .ZN(
        n32817) );
  NAND2_X2 U14782 ( .A1(n33304), .A2(n28194), .ZN(n16286) );
  XOR2_X1 U14792 ( .A1(n15691), .A2(n32818), .Z(n26630) );
  XOR2_X1 U14793 ( .A1(n23504), .A2(n15690), .Z(n32818) );
  NAND2_X2 U14795 ( .A1(n3379), .A2(n777), .ZN(n34084) );
  OAI22_X2 U14796 ( .A1(n21438), .A2(n21224), .B1(n21223), .B2(n8398), .ZN(
        n11232) );
  NAND3_X1 U14802 ( .A1(n16091), .A2(n8045), .A3(n30059), .ZN(n32819) );
  NOR2_X2 U14804 ( .A1(n8970), .A2(n279), .ZN(n32983) );
  NAND2_X2 U14807 ( .A1(n4289), .A2(n20401), .ZN(n31079) );
  XOR2_X1 U14808 ( .A1(n10758), .A2(n23164), .Z(n4446) );
  XOR2_X1 U14811 ( .A1(n23441), .A2(n23211), .Z(n23164) );
  INV_X2 U14812 ( .I(n28374), .ZN(n26806) );
  NAND2_X2 U14813 ( .A1(n32821), .A2(n23802), .ZN(n28374) );
  AND2_X1 U14818 ( .A1(n23803), .A2(n23801), .Z(n32821) );
  XOR2_X1 U14819 ( .A1(n19772), .A2(n19399), .Z(n19733) );
  NAND2_X2 U14821 ( .A1(n8576), .A2(n8857), .ZN(n9106) );
  OR2_X1 U14831 ( .A1(n26448), .A2(n21258), .Z(n33683) );
  NOR2_X2 U14832 ( .A1(n9195), .A2(n25701), .ZN(n25766) );
  NAND2_X1 U14833 ( .A1(n16170), .A2(n25), .ZN(n2258) );
  OR2_X1 U14841 ( .A1(n29342), .A2(n22398), .Z(n33190) );
  BUF_X2 U14844 ( .I(n2483), .Z(n32822) );
  XOR2_X1 U14846 ( .A1(n24528), .A2(n549), .Z(n28746) );
  XOR2_X1 U14847 ( .A1(n4662), .A2(n4661), .Z(n16536) );
  XOR2_X1 U14854 ( .A1(n32824), .A2(n23239), .Z(Ciphertext[75]) );
  NAND3_X2 U14857 ( .A1(n10942), .A2(n32990), .A3(n10940), .ZN(n32824) );
  XOR2_X1 U14858 ( .A1(n15877), .A2(n10159), .Z(n30985) );
  XOR2_X1 U14860 ( .A1(n31899), .A2(n10729), .Z(n5229) );
  INV_X4 U14862 ( .I(n25235), .ZN(n34115) );
  XOR2_X1 U14867 ( .A1(n23137), .A2(n23532), .Z(n23219) );
  OAI21_X2 U14870 ( .A1(n11064), .A2(n10687), .B(n28467), .ZN(n10811) );
  OAI22_X2 U14872 ( .A1(n32826), .A2(n2773), .B1(n2775), .B2(n11317), .ZN(
        n3519) );
  NAND2_X2 U14877 ( .A1(n4967), .A2(n14055), .ZN(n32828) );
  NAND2_X2 U14879 ( .A1(n29334), .A2(n15318), .ZN(n4967) );
  OAI21_X1 U14881 ( .A1(n5492), .A2(n24996), .B(n7940), .ZN(n9478) );
  NAND2_X2 U14882 ( .A1(n28647), .A2(n19530), .ZN(n28108) );
  NAND2_X2 U14884 ( .A1(n3266), .A2(n11967), .ZN(n28523) );
  NOR2_X2 U14885 ( .A1(n1940), .A2(n1233), .ZN(n32829) );
  NAND2_X2 U14886 ( .A1(n15253), .A2(n13472), .ZN(n6354) );
  XOR2_X1 U14888 ( .A1(n31727), .A2(n16705), .Z(n12924) );
  INV_X2 U14890 ( .I(n11845), .ZN(n24316) );
  OAI22_X1 U14891 ( .A1(n23946), .A2(n30359), .B1(n11676), .B2(n10187), .ZN(
        n8675) );
  OAI22_X2 U14892 ( .A1(n15225), .A2(n20381), .B1(n15162), .B2(n20633), .ZN(
        n11241) );
  NAND2_X2 U14898 ( .A1(n20445), .A2(n20384), .ZN(n20633) );
  BUF_X2 U14901 ( .I(n19901), .Z(n8421) );
  XOR2_X1 U14906 ( .A1(n20930), .A2(n20929), .Z(n33673) );
  NAND3_X2 U14908 ( .A1(n16235), .A2(n30152), .A3(n32832), .ZN(n21588) );
  INV_X2 U14909 ( .I(n21866), .ZN(n32833) );
  XOR2_X1 U14910 ( .A1(n32516), .A2(n25098), .Z(n23398) );
  OAI21_X2 U14916 ( .A1(n21254), .A2(n32644), .B(n32834), .ZN(n29854) );
  AOI22_X2 U14923 ( .A1(n15932), .A2(n9699), .B1(n15931), .B2(n27462), .ZN(
        n32834) );
  BUF_X2 U14926 ( .I(n22979), .Z(n27814) );
  BUF_X4 U14927 ( .I(n16568), .Z(n330) );
  XOR2_X1 U14934 ( .A1(n19637), .A2(n8633), .Z(n19433) );
  NAND2_X2 U14936 ( .A1(n14697), .A2(n19246), .ZN(n19637) );
  BUF_X4 U14937 ( .I(n23904), .Z(n6414) );
  XOR2_X1 U14938 ( .A1(n22171), .A2(n3781), .Z(n175) );
  XOR2_X1 U14939 ( .A1(n30999), .A2(n22211), .Z(n3781) );
  NAND2_X2 U14944 ( .A1(n16421), .A2(n8434), .ZN(n20780) );
  NAND3_X1 U14945 ( .A1(n31103), .A2(n29250), .A3(n19808), .ZN(n19809) );
  OAI22_X2 U14950 ( .A1(n14725), .A2(n27104), .B1(n31228), .B2(n2798), .ZN(
        n24383) );
  NAND2_X2 U14953 ( .A1(n31218), .A2(n7893), .ZN(n7892) );
  OAI21_X2 U14954 ( .A1(n3224), .A2(n1213), .B(n33493), .ZN(n3223) );
  XOR2_X1 U14967 ( .A1(n13455), .A2(n13456), .Z(n27257) );
  NAND2_X1 U14970 ( .A1(n28657), .A2(n28655), .ZN(n10823) );
  NAND2_X1 U14976 ( .A1(n4733), .A2(n14056), .ZN(n18625) );
  NAND2_X2 U14978 ( .A1(n26962), .A2(n16564), .ZN(n4733) );
  AND2_X1 U14984 ( .A1(n21426), .A2(n13286), .Z(n33418) );
  XOR2_X1 U14986 ( .A1(n7597), .A2(n7599), .Z(n22598) );
  XOR2_X1 U14987 ( .A1(n14277), .A2(n31552), .Z(n675) );
  XOR2_X1 U14988 ( .A1(n17798), .A2(n24494), .Z(n10685) );
  XOR2_X1 U14994 ( .A1(n24811), .A2(n24553), .Z(n24494) );
  NAND3_X2 U15001 ( .A1(n23711), .A2(n23709), .A3(n23710), .ZN(n12981) );
  BUF_X2 U15017 ( .I(n17338), .Z(n31850) );
  XOR2_X1 U15020 ( .A1(n32835), .A2(n13899), .Z(n21198) );
  XOR2_X1 U15022 ( .A1(n32892), .A2(n13898), .Z(n32835) );
  AOI22_X2 U15026 ( .A1(n17139), .A2(n28429), .B1(n30506), .B2(n28450), .ZN(
        n21488) );
  OAI21_X2 U15030 ( .A1(n5377), .A2(n5376), .B(n26516), .ZN(n32836) );
  NAND2_X2 U15031 ( .A1(n17561), .A2(n4349), .ZN(n24095) );
  AND2_X1 U15033 ( .A1(n25563), .A2(n28093), .Z(n25520) );
  INV_X1 U15034 ( .I(n30252), .ZN(n33813) );
  AND2_X1 U15039 ( .A1(n30252), .A2(n23833), .Z(n33812) );
  INV_X1 U15044 ( .I(n17280), .ZN(n31801) );
  NOR2_X2 U15057 ( .A1(n2209), .A2(n25686), .ZN(n14732) );
  NAND2_X2 U15059 ( .A1(n715), .A2(n28651), .ZN(n14795) );
  NOR2_X1 U15060 ( .A1(n32837), .A2(n27007), .ZN(n11566) );
  NAND2_X2 U15061 ( .A1(n13535), .A2(n30631), .ZN(n27007) );
  AOI21_X2 U15065 ( .A1(n23601), .A2(n5357), .B(n27049), .ZN(n14548) );
  XOR2_X1 U15077 ( .A1(n6329), .A2(n32838), .Z(n32924) );
  INV_X2 U15089 ( .I(n522), .ZN(n32926) );
  XOR2_X1 U15091 ( .A1(n19558), .A2(n19755), .Z(n19611) );
  NAND3_X2 U15094 ( .A1(n18526), .A2(n18527), .A3(n18528), .ZN(n19755) );
  NOR2_X2 U15095 ( .A1(n5704), .A2(n7592), .ZN(n21711) );
  XOR2_X1 U15098 ( .A1(n602), .A2(n2756), .Z(n4327) );
  XOR2_X1 U15099 ( .A1(n29832), .A2(n20684), .Z(n602) );
  XOR2_X1 U15101 ( .A1(n20956), .A2(n32839), .Z(n29303) );
  XOR2_X1 U15103 ( .A1(n27054), .A2(n20896), .Z(n32839) );
  NAND2_X2 U15110 ( .A1(n15344), .A2(n32840), .ZN(n34004) );
  NAND2_X2 U15111 ( .A1(n25592), .A2(n9862), .ZN(n388) );
  INV_X4 U15113 ( .I(n9219), .ZN(n24292) );
  OAI21_X2 U15118 ( .A1(n2325), .A2(n32323), .B(n24127), .ZN(n34093) );
  XOR2_X1 U15120 ( .A1(n32841), .A2(n23264), .Z(n27667) );
  NOR2_X2 U15122 ( .A1(n16922), .A2(n22743), .ZN(n23395) );
  BUF_X4 U15129 ( .I(n29321), .Z(n33992) );
  XOR2_X1 U15131 ( .A1(n19686), .A2(n32844), .Z(n19586) );
  INV_X2 U15132 ( .I(n19341), .ZN(n32844) );
  NAND2_X1 U15135 ( .A1(n33853), .A2(n29568), .ZN(n14838) );
  INV_X2 U15138 ( .I(n13073), .ZN(n21414) );
  NOR2_X1 U15139 ( .A1(n29322), .A2(n6176), .ZN(n2219) );
  INV_X2 U15141 ( .I(n6275), .ZN(n16848) );
  NAND2_X1 U15142 ( .A1(n12564), .A2(n33218), .ZN(n124) );
  NOR2_X1 U15143 ( .A1(n32852), .A2(n9480), .ZN(n27968) );
  NOR2_X1 U15154 ( .A1(n9052), .A2(n33643), .ZN(n27099) );
  OAI21_X1 U15172 ( .A1(n25053), .A2(n27610), .B(n32845), .ZN(n25055) );
  AOI22_X1 U15174 ( .A1(n17728), .A2(n25062), .B1(n17729), .B2(n27610), .ZN(
        n32845) );
  NAND2_X2 U15177 ( .A1(n27624), .A2(n1164), .ZN(n10272) );
  OAI21_X2 U15178 ( .A1(n31822), .A2(n25890), .B(n30811), .ZN(n31378) );
  NAND2_X2 U15182 ( .A1(n22655), .A2(n22951), .ZN(n22952) );
  NAND2_X2 U15185 ( .A1(n22258), .A2(n6540), .ZN(n22655) );
  OAI21_X2 U15187 ( .A1(n10221), .A2(n6981), .B(n1223), .ZN(n33197) );
  XOR2_X1 U15188 ( .A1(n32846), .A2(n30156), .Z(n31650) );
  XOR2_X1 U15190 ( .A1(n23123), .A2(n23124), .Z(n32846) );
  XOR2_X1 U15192 ( .A1(n21995), .A2(n22282), .Z(n15727) );
  XOR2_X1 U15193 ( .A1(n33150), .A2(n22255), .Z(n21995) );
  INV_X2 U15200 ( .I(n11805), .ZN(n33739) );
  AOI21_X2 U15205 ( .A1(n6802), .A2(n6675), .B(n6674), .ZN(n32860) );
  XOR2_X1 U15206 ( .A1(n32847), .A2(n25259), .Z(Ciphertext[83]) );
  AOI22_X1 U15210 ( .A1(n26497), .A2(n27429), .B1(n8035), .B2(n8036), .ZN(
        n32847) );
  NAND2_X2 U15215 ( .A1(n32848), .A2(n5888), .ZN(n17236) );
  NAND2_X1 U15221 ( .A1(n14988), .A2(n28912), .ZN(n32848) );
  NAND2_X1 U15223 ( .A1(n5789), .A2(n28885), .ZN(n19205) );
  OAI22_X2 U15224 ( .A1(n9645), .A2(n843), .B1(n5764), .B2(n548), .ZN(n9616)
         );
  AOI22_X2 U15226 ( .A1(n10145), .A2(n843), .B1(n9172), .B2(n11968), .ZN(n5764) );
  NAND3_X2 U15227 ( .A1(n29521), .A2(n15670), .A3(n10066), .ZN(n10469) );
  NAND2_X2 U15231 ( .A1(n11571), .A2(n15054), .ZN(n7871) );
  OR2_X1 U15234 ( .A1(n33189), .A2(n29230), .Z(n34121) );
  NAND2_X2 U15235 ( .A1(n26903), .A2(n28664), .ZN(n33146) );
  NOR2_X2 U15239 ( .A1(n11695), .A2(n11698), .ZN(n25670) );
  NAND3_X1 U15242 ( .A1(n19292), .A2(n18682), .A3(n746), .ZN(n32849) );
  XOR2_X1 U15247 ( .A1(n32850), .A2(n29550), .Z(n16401) );
  XOR2_X1 U15250 ( .A1(n572), .A2(n33742), .Z(n32850) );
  OR2_X1 U15252 ( .A1(n14780), .A2(n26447), .Z(n25684) );
  INV_X4 U15255 ( .I(n11956), .ZN(n28867) );
  INV_X2 U15257 ( .I(n32851), .ZN(n34167) );
  XOR2_X1 U15258 ( .A1(n6848), .A2(n28062), .Z(n32851) );
  XOR2_X1 U15260 ( .A1(n23506), .A2(n23126), .Z(n8071) );
  XOR2_X1 U15263 ( .A1(n29885), .A2(n23293), .Z(n23506) );
  NOR2_X1 U15264 ( .A1(n9479), .A2(n9478), .ZN(n32852) );
  NAND2_X1 U15272 ( .A1(n32853), .A2(n30740), .ZN(n7336) );
  NAND2_X1 U15274 ( .A1(n7341), .A2(n26744), .ZN(n32853) );
  AND3_X1 U15275 ( .A1(n15807), .A2(n21297), .A3(n4989), .Z(n26025) );
  XOR2_X1 U15280 ( .A1(n5149), .A2(n32854), .Z(n19527) );
  XOR2_X1 U15281 ( .A1(n8561), .A2(n26794), .Z(n32854) );
  BUF_X4 U15284 ( .I(n13670), .Z(n11187) );
  OR2_X1 U15285 ( .A1(n26374), .A2(n24340), .Z(n24343) );
  OAI21_X2 U15288 ( .A1(n11757), .A2(n11949), .B(n783), .ZN(n33323) );
  INV_X2 U15290 ( .I(n9958), .ZN(n14137) );
  BUF_X4 U15291 ( .I(n31721), .Z(n33301) );
  NAND2_X2 U15292 ( .A1(n24933), .A2(n24351), .ZN(n17479) );
  BUF_X4 U15296 ( .I(n25051), .Z(n31640) );
  NAND3_X1 U15301 ( .A1(n8766), .A2(n32897), .A3(n33399), .ZN(n4325) );
  INV_X1 U15302 ( .I(n888), .ZN(n24101) );
  NAND3_X1 U15305 ( .A1(n5160), .A2(n24104), .A3(n888), .ZN(n28524) );
  OAI21_X1 U15306 ( .A1(n24102), .A2(n12098), .B(n888), .ZN(n4928) );
  NAND2_X1 U15318 ( .A1(n24667), .A2(n25536), .ZN(n9915) );
  OAI21_X1 U15319 ( .A1(n24667), .A2(n25536), .B(n736), .ZN(n26921) );
  NOR2_X1 U15322 ( .A1(n8062), .A2(n11200), .ZN(n11201) );
  NAND2_X1 U15325 ( .A1(n3925), .A2(n20142), .ZN(n33003) );
  NAND3_X1 U15328 ( .A1(n10266), .A2(n10265), .A3(n10268), .ZN(n33513) );
  NOR2_X1 U15329 ( .A1(n26566), .A2(n20577), .ZN(n33149) );
  INV_X1 U15334 ( .I(n26566), .ZN(n8528) );
  NOR2_X1 U15336 ( .A1(n6230), .A2(n26566), .ZN(n27806) );
  OAI21_X1 U15338 ( .A1(n29271), .A2(n26415), .B(n30125), .ZN(n26221) );
  OAI21_X1 U15344 ( .A1(n33400), .A2(n33399), .B(n1204), .ZN(n33957) );
  NOR2_X2 U15345 ( .A1(n24888), .A2(n2092), .ZN(n28706) );
  NAND2_X1 U15350 ( .A1(n4243), .A2(n33480), .ZN(n24724) );
  INV_X2 U15358 ( .I(n10622), .ZN(n998) );
  NAND2_X1 U15359 ( .A1(n797), .A2(n24150), .ZN(n12208) );
  OAI21_X1 U15367 ( .A1(n797), .A2(n2744), .B(n26545), .ZN(n2746) );
  NOR2_X1 U15368 ( .A1(n10042), .A2(n12423), .ZN(n30569) );
  NAND2_X1 U15369 ( .A1(n1209), .A2(n16798), .ZN(n1472) );
  OR2_X1 U15381 ( .A1(n14490), .A2(n15065), .Z(n14491) );
  AOI22_X1 U15382 ( .A1(n8263), .A2(n14490), .B1(n15818), .B2(n15996), .ZN(
        n3845) );
  OAI22_X1 U15383 ( .A1(n24176), .A2(n15790), .B1(n14052), .B2(n14490), .ZN(
        n3256) );
  NAND2_X1 U15385 ( .A1(n1007), .A2(n2386), .ZN(n33367) );
  CLKBUF_X2 U15387 ( .I(n18818), .Z(n16393) );
  INV_X1 U15388 ( .I(n18818), .ZN(n18639) );
  NAND2_X1 U15392 ( .A1(n22883), .A2(n22882), .ZN(n33383) );
  NAND2_X1 U15393 ( .A1(n22883), .A2(n13274), .ZN(n3778) );
  AOI21_X1 U15400 ( .A1(n10045), .A2(n23795), .B(n5777), .ZN(n5776) );
  INV_X2 U15406 ( .I(n23795), .ZN(n845) );
  NAND2_X1 U15409 ( .A1(n13698), .A2(n25297), .ZN(n33956) );
  NOR2_X1 U15412 ( .A1(n6869), .A2(n23917), .ZN(n4197) );
  BUF_X1 U15413 ( .I(n25546), .Z(n8320) );
  NOR2_X1 U15414 ( .A1(n13334), .A2(n27168), .ZN(n6654) );
  INV_X1 U15415 ( .I(n5790), .ZN(n11868) );
  NAND2_X1 U15416 ( .A1(n7501), .A2(n6483), .ZN(n33955) );
  INV_X2 U15417 ( .I(n14650), .ZN(n25066) );
  INV_X1 U15421 ( .I(n30323), .ZN(n29670) );
  NAND2_X1 U15422 ( .A1(n25568), .A2(n3638), .ZN(n10959) );
  AOI21_X1 U15423 ( .A1(n9022), .A2(n33237), .B(n9910), .ZN(n7904) );
  NOR2_X1 U15429 ( .A1(n20575), .A2(n27785), .ZN(n27902) );
  NAND2_X1 U15430 ( .A1(n1463), .A2(n886), .ZN(n1462) );
  INV_X1 U15434 ( .I(n678), .ZN(n886) );
  CLKBUF_X4 U15444 ( .I(n18494), .Z(n16564) );
  NOR2_X2 U15445 ( .A1(n23539), .A2(n23538), .ZN(n12547) );
  BUF_X2 U15446 ( .I(n4287), .Z(n28579) );
  OAI21_X1 U15447 ( .A1(n23950), .A2(n30359), .B(n23620), .ZN(n13774) );
  AND2_X1 U15455 ( .A1(n13308), .A2(n23949), .Z(n23620) );
  NOR2_X1 U15456 ( .A1(n13698), .A2(n8105), .ZN(n15785) );
  NOR2_X1 U15459 ( .A1(n33460), .A2(n8105), .ZN(n15481) );
  OAI21_X1 U15463 ( .A1(n25537), .A2(n16826), .B(n8105), .ZN(n34033) );
  NOR2_X1 U15464 ( .A1(n33480), .A2(n18242), .ZN(n17815) );
  AOI21_X1 U15468 ( .A1(n17815), .A2(n25902), .B(n10792), .ZN(n12420) );
  INV_X1 U15469 ( .I(n17815), .ZN(n11186) );
  AOI22_X1 U15471 ( .A1(n10303), .A2(n22547), .B1(n22551), .B2(n27402), .ZN(
        n27416) );
  NAND2_X1 U15472 ( .A1(n25800), .A2(n25799), .ZN(n25802) );
  OR2_X2 U15475 ( .A1(n28557), .A2(n7806), .Z(n32855) );
  OR2_X2 U15477 ( .A1(n28557), .A2(n7806), .Z(n32856) );
  NAND2_X1 U15480 ( .A1(n22784), .A2(n3898), .ZN(n17900) );
  AND2_X1 U15482 ( .A1(n3515), .A2(n3340), .Z(n6780) );
  INV_X2 U15483 ( .I(n7555), .ZN(n788) );
  OAI21_X1 U15489 ( .A1(n8178), .A2(n1239), .B(n29056), .ZN(n29863) );
  NAND3_X1 U15495 ( .A1(n30280), .A2(n29056), .A3(n7809), .ZN(n7727) );
  CLKBUF_X8 U15496 ( .I(n8238), .Z(n32917) );
  OR2_X1 U15497 ( .A1(n7993), .A2(n2022), .Z(n23858) );
  INV_X2 U15499 ( .I(n7889), .ZN(n13457) );
  NOR2_X1 U15500 ( .A1(n34109), .A2(n5466), .ZN(n25237) );
  NAND2_X1 U15502 ( .A1(n6074), .A2(n21466), .ZN(n21283) );
  CLKBUF_X2 U15503 ( .I(n6074), .Z(n26728) );
  OAI21_X1 U15504 ( .A1(n27104), .A2(n24060), .B(n13601), .ZN(n3039) );
  INV_X1 U15506 ( .I(n16422), .ZN(n16112) );
  INV_X1 U15513 ( .I(n16529), .ZN(n1113) );
  OAI21_X1 U15516 ( .A1(n22567), .A2(n28692), .B(n22683), .ZN(n22568) );
  NOR2_X1 U15519 ( .A1(n9939), .A2(n23936), .ZN(n15098) );
  INV_X2 U15521 ( .I(n9939), .ZN(n13242) );
  AOI21_X1 U15529 ( .A1(n17166), .A2(n33205), .B(n16287), .ZN(n4505) );
  NOR2_X1 U15535 ( .A1(n16287), .A2(n31417), .ZN(n18864) );
  NAND2_X1 U15540 ( .A1(n14194), .A2(n11203), .ZN(n18842) );
  INV_X1 U15541 ( .I(n14194), .ZN(n19216) );
  NAND2_X1 U15543 ( .A1(n7557), .A2(n14194), .ZN(n16336) );
  OR2_X1 U15552 ( .A1(n13413), .A2(n16384), .Z(n23590) );
  INV_X1 U15565 ( .I(n25258), .ZN(n25250) );
  AND2_X1 U15566 ( .A1(n13532), .A2(n32875), .Z(n9861) );
  OAI22_X1 U15568 ( .A1(n28952), .A2(n16793), .B1(n25514), .B2(n2480), .ZN(
        n33401) );
  INV_X1 U15570 ( .I(n24643), .ZN(n242) );
  OAI21_X1 U15577 ( .A1(n13078), .A2(n9065), .B(n22595), .ZN(n22596) );
  NAND3_X1 U15584 ( .A1(n30708), .A2(n25102), .A3(n3824), .ZN(n32984) );
  NOR2_X1 U15588 ( .A1(n27233), .A2(n25951), .ZN(n27232) );
  NAND2_X1 U15589 ( .A1(n24232), .A2(n972), .ZN(n27381) );
  AOI22_X1 U15598 ( .A1(n6772), .A2(n29120), .B1(n24232), .B2(n14399), .ZN(
        n3633) );
  AOI22_X1 U15599 ( .A1(n2558), .A2(n24232), .B1(n6476), .B2(n14399), .ZN(
        n29836) );
  NAND2_X1 U15605 ( .A1(n25586), .A2(n34169), .ZN(n25530) );
  NOR2_X1 U15606 ( .A1(n25590), .A2(n25586), .ZN(n13560) );
  INV_X1 U15607 ( .I(n12042), .ZN(n967) );
  NAND2_X1 U15617 ( .A1(n1786), .A2(n12476), .ZN(n25113) );
  CLKBUF_X1 U15629 ( .I(n16380), .Z(n31207) );
  NAND2_X1 U15630 ( .A1(n25066), .A2(n31207), .ZN(n16836) );
  INV_X1 U15632 ( .I(n22832), .ZN(n806) );
  OR2_X2 U15635 ( .A1(n22832), .A2(n4110), .Z(n4731) );
  CLKBUF_X4 U15637 ( .I(n9301), .Z(n9195) );
  INV_X1 U15638 ( .I(n9870), .ZN(n22580) );
  INV_X1 U15642 ( .I(n25128), .ZN(n25130) );
  NAND2_X1 U15653 ( .A1(n25128), .A2(n1075), .ZN(n31617) );
  CLKBUF_X4 U15654 ( .I(n15012), .Z(n14454) );
  NAND2_X1 U15655 ( .A1(n4655), .A2(n14147), .ZN(n24092) );
  INV_X2 U15657 ( .I(n14147), .ZN(n28694) );
  OR3_X1 U15659 ( .A1(n7081), .A2(n25337), .A3(n11132), .Z(n25342) );
  INV_X1 U15660 ( .I(n30991), .ZN(n23955) );
  OAI21_X1 U15661 ( .A1(n15974), .A2(n29056), .B(n24263), .ZN(n13616) );
  NOR2_X2 U15666 ( .A1(n27854), .A2(n26949), .ZN(n13615) );
  NAND2_X1 U15667 ( .A1(n18143), .A2(n22499), .ZN(n32858) );
  NAND2_X2 U15669 ( .A1(n22500), .A2(n22691), .ZN(n18143) );
  OR2_X1 U15670 ( .A1(n25621), .A2(n25620), .Z(n16001) );
  NAND2_X1 U15673 ( .A1(n23026), .A2(n26169), .ZN(n11495) );
  CLKBUF_X4 U15677 ( .I(n23706), .Z(n14080) );
  INV_X1 U15679 ( .I(n25624), .ZN(n1219) );
  OAI21_X1 U15682 ( .A1(n24327), .A2(n24328), .B(n24326), .ZN(n28030) );
  INV_X1 U15684 ( .I(n12746), .ZN(n33926) );
  INV_X2 U15688 ( .I(n11912), .ZN(n12746) );
  BUF_X2 U15689 ( .I(n23834), .Z(n16424) );
  INV_X1 U15690 ( .I(n16424), .ZN(n33166) );
  NAND3_X1 U15691 ( .A1(n2640), .A2(n27038), .A3(n31615), .ZN(n668) );
  NOR3_X1 U15699 ( .A1(n793), .A2(n26120), .A3(n27038), .ZN(n17747) );
  NOR2_X1 U15700 ( .A1(n26120), .A2(n6713), .ZN(n8142) );
  NAND2_X1 U15702 ( .A1(n7753), .A2(n15414), .ZN(n21613) );
  OAI21_X1 U15710 ( .A1(n1316), .A2(n21752), .B(n15414), .ZN(n13662) );
  CLKBUF_X4 U15714 ( .I(n25654), .Z(n7083) );
  NAND2_X1 U15715 ( .A1(n8924), .A2(n31835), .ZN(n21151) );
  INV_X2 U15716 ( .I(n21395), .ZN(n12325) );
  INV_X4 U15718 ( .I(n23767), .ZN(n23770) );
  NOR2_X1 U15719 ( .A1(n9399), .A2(n22483), .ZN(n33021) );
  NAND3_X1 U15720 ( .A1(n9399), .A2(n22483), .A3(n8287), .ZN(n28463) );
  AOI21_X1 U15723 ( .A1(n12586), .A2(n22982), .B(n28234), .ZN(n8037) );
  NAND2_X1 U15728 ( .A1(n25760), .A2(n4407), .ZN(n30221) );
  OAI21_X1 U15733 ( .A1(n11898), .A2(n33278), .B(n24611), .ZN(n8648) );
  OAI21_X1 U15736 ( .A1(n1300), .A2(n22497), .B(n31933), .ZN(n22020) );
  NAND2_X1 U15740 ( .A1(n22628), .A2(n31933), .ZN(n33938) );
  AND3_X2 U15741 ( .A1(n32998), .A2(n3004), .A3(n23942), .Z(n10019) );
  CLKBUF_X2 U15742 ( .I(n2635), .Z(n33596) );
  NOR2_X1 U15744 ( .A1(n13995), .A2(n2635), .ZN(n30488) );
  NAND2_X1 U15750 ( .A1(n20429), .A2(n2928), .ZN(n31111) );
  NAND2_X1 U15753 ( .A1(n28414), .A2(n20429), .ZN(n17808) );
  INV_X1 U15754 ( .I(n20429), .ZN(n20498) );
  NOR2_X1 U15761 ( .A1(n20429), .A2(n2928), .ZN(n20259) );
  AND2_X2 U15764 ( .A1(n19901), .A2(n27655), .Z(n31593) );
  NOR2_X1 U15768 ( .A1(n6605), .A2(n30976), .ZN(n11925) );
  NAND2_X1 U15787 ( .A1(n25326), .A2(n16528), .ZN(n33921) );
  INV_X1 U15792 ( .I(n25796), .ZN(n25781) );
  OAI21_X1 U15798 ( .A1(n12395), .A2(n25797), .B(n25796), .ZN(n25800) );
  NOR2_X1 U15801 ( .A1(n19451), .A2(n16317), .ZN(n3591) );
  NAND2_X1 U15808 ( .A1(n7335), .A2(n32909), .ZN(n30708) );
  NAND2_X1 U15810 ( .A1(n1127), .A2(n2547), .ZN(n22669) );
  NOR2_X1 U15812 ( .A1(n2141), .A2(n24242), .ZN(n3947) );
  NAND2_X1 U15813 ( .A1(n5141), .A2(n21426), .ZN(n28342) );
  NAND2_X1 U15819 ( .A1(n21426), .A2(n17624), .ZN(n30091) );
  OAI22_X1 U15821 ( .A1(n30091), .A2(n28211), .B1(n21426), .B2(n28594), .ZN(
        n21195) );
  OAI21_X1 U15823 ( .A1(n17624), .A2(n21426), .B(n28342), .ZN(n21196) );
  INV_X1 U15824 ( .I(n15806), .ZN(n23069) );
  NAND2_X1 U15825 ( .A1(n23070), .A2(n15806), .ZN(n4806) );
  NAND2_X1 U15830 ( .A1(n22905), .A2(n15806), .ZN(n22907) );
  INV_X1 U15831 ( .I(n15296), .ZN(n18079) );
  AOI22_X1 U15835 ( .A1(n11058), .A2(n11059), .B1(n4067), .B2(n7181), .ZN(
        n11057) );
  OAI21_X1 U15837 ( .A1(n903), .A2(n4100), .B(n3810), .ZN(n9158) );
  NAND2_X2 U15838 ( .A1(n5741), .A2(n24193), .ZN(n5690) );
  NAND3_X1 U15844 ( .A1(n18220), .A2(n25697), .A3(n25695), .ZN(n33119) );
  AND3_X1 U15856 ( .A1(n25082), .A2(n25107), .A3(n787), .Z(n24857) );
  NAND2_X1 U15858 ( .A1(n33616), .A2(n27168), .ZN(n29753) );
  AOI22_X1 U15860 ( .A1(n8049), .A2(n719), .B1(n26120), .B2(n7891), .ZN(n11388) );
  OAI22_X1 U15863 ( .A1(n26120), .A2(n737), .B1(n793), .B2(n27168), .ZN(n8049)
         );
  NAND2_X1 U15866 ( .A1(n34009), .A2(n4069), .ZN(n17880) );
  AOI22_X1 U15873 ( .A1(n25013), .A2(n25014), .B1(n25015), .B2(n17240), .ZN(
        n6283) );
  INV_X2 U15879 ( .I(n11401), .ZN(n21642) );
  CLKBUF_X1 U15882 ( .I(n19938), .Z(n28644) );
  OR2_X1 U15886 ( .A1(n11548), .A2(n18075), .Z(n25260) );
  NAND3_X1 U15887 ( .A1(n16393), .A2(n18815), .A3(n18515), .ZN(n4645) );
  NOR2_X1 U15889 ( .A1(n15296), .A2(n9793), .ZN(n3248) );
  INV_X1 U15893 ( .I(n5708), .ZN(n33567) );
  NAND3_X2 U15895 ( .A1(n1243), .A2(n24272), .A3(n8412), .ZN(n24495) );
  NAND2_X2 U15896 ( .A1(n6400), .A2(n30123), .ZN(n32861) );
  XNOR2_X1 U15913 ( .A1(n24695), .A2(n24740), .ZN(n29545) );
  NAND2_X1 U15915 ( .A1(n6400), .A2(n30123), .ZN(n17052) );
  OAI21_X1 U15922 ( .A1(n25755), .A2(n717), .B(n11899), .ZN(n30877) );
  NAND2_X1 U15927 ( .A1(n13472), .A2(n2654), .ZN(n24279) );
  INV_X2 U15931 ( .I(n665), .ZN(n34008) );
  AOI22_X1 U15932 ( .A1(n20269), .A2(n5781), .B1(n17693), .B2(n20494), .ZN(
        n20650) );
  NAND2_X1 U15935 ( .A1(n15250), .A2(n15249), .ZN(n33958) );
  INV_X2 U15936 ( .I(n10281), .ZN(n32862) );
  NOR3_X1 U15939 ( .A1(n10606), .A2(n10605), .A3(n30018), .ZN(n27060) );
  INV_X1 U15940 ( .I(n4886), .ZN(n5755) );
  BUF_X2 U15948 ( .I(n28119), .Z(n32878) );
  INV_X1 U15953 ( .I(n23067), .ZN(n18159) );
  NOR2_X1 U15961 ( .A1(n23067), .A2(n23070), .ZN(n30967) );
  OAI22_X1 U15962 ( .A1(n12043), .A2(n31914), .B1(n29626), .B2(n22639), .ZN(
        n33610) );
  INV_X1 U15963 ( .I(n24829), .ZN(n11842) );
  NOR2_X1 U15968 ( .A1(n24250), .A2(n24248), .ZN(n31664) );
  NAND2_X1 U15972 ( .A1(n6512), .A2(n24430), .ZN(n32863) );
  AOI22_X1 U15973 ( .A1(n1219), .A2(n31921), .B1(n16397), .B2(n32896), .ZN(
        n33773) );
  NOR2_X1 U15981 ( .A1(n3487), .A2(n16959), .ZN(n27020) );
  INV_X2 U15985 ( .I(n16959), .ZN(n28899) );
  INV_X1 U15987 ( .I(n25014), .ZN(n24976) );
  AOI21_X1 U15990 ( .A1(n901), .A2(n8314), .B(n1728), .ZN(n26803) );
  NOR2_X1 U15998 ( .A1(n8766), .A2(n1209), .ZN(n33102) );
  INV_X1 U16001 ( .I(n25302), .ZN(n32864) );
  OAI21_X1 U16004 ( .A1(n11255), .A2(n24325), .B(n30186), .ZN(n9826) );
  NAND2_X1 U16005 ( .A1(n3729), .A2(n1083), .ZN(n3728) );
  CLKBUF_X1 U16008 ( .I(n19284), .Z(n30501) );
  CLKBUF_X12 U16009 ( .I(n20137), .Z(n27911) );
  AOI22_X1 U16010 ( .A1(n23957), .A2(n13720), .B1(n14232), .B2(n23825), .ZN(
        n29811) );
  NAND2_X1 U16019 ( .A1(n14133), .A2(n13720), .ZN(n13981) );
  AOI22_X1 U16022 ( .A1(n29541), .A2(n998), .B1(n905), .B2(n22467), .ZN(n29790) );
  NAND3_X1 U16023 ( .A1(n32868), .A2(n27622), .A3(n5915), .ZN(n12071) );
  OR2_X1 U16026 ( .A1(n17936), .A2(n11920), .Z(n18094) );
  NOR2_X1 U16027 ( .A1(n18098), .A2(n11920), .ZN(n16866) );
  INV_X2 U16030 ( .I(n7492), .ZN(n11000) );
  INV_X2 U16032 ( .I(n17273), .ZN(n11571) );
  CLKBUF_X1 U16034 ( .I(n28196), .Z(n33851) );
  INV_X2 U16036 ( .I(n11559), .ZN(n11904) );
  NOR3_X1 U16037 ( .A1(n23806), .A2(n11904), .A3(n1247), .ZN(n29705) );
  NAND2_X1 U16040 ( .A1(n1247), .A2(n11904), .ZN(n12248) );
  OAI21_X1 U16050 ( .A1(n1247), .A2(n11904), .B(n23806), .ZN(n15683) );
  AOI21_X1 U16051 ( .A1(n1100), .A2(n11904), .B(n28273), .ZN(n18167) );
  NAND2_X1 U16053 ( .A1(n1850), .A2(n12476), .ZN(n12295) );
  INV_X2 U16057 ( .I(n11987), .ZN(n25199) );
  CLKBUF_X4 U16061 ( .I(n25014), .Z(n14959) );
  INV_X1 U16072 ( .I(n386), .ZN(n17396) );
  NOR2_X1 U16074 ( .A1(n9778), .A2(n5035), .ZN(n28877) );
  INV_X1 U16076 ( .I(n3093), .ZN(n32932) );
  NAND2_X1 U16084 ( .A1(n3093), .A2(n5455), .ZN(n19313) );
  NAND2_X1 U16093 ( .A1(n10999), .A2(n3093), .ZN(n33261) );
  CLKBUF_X4 U16094 ( .I(n5612), .Z(n25991) );
  NAND2_X1 U16095 ( .A1(n25308), .A2(n32096), .ZN(n33169) );
  OAI21_X1 U16096 ( .A1(n25391), .A2(n17717), .B(n25962), .ZN(n9548) );
  NAND2_X1 U16098 ( .A1(n17717), .A2(n25962), .ZN(n18099) );
  NOR2_X1 U16099 ( .A1(n25487), .A2(n25462), .ZN(n17199) );
  NOR2_X1 U16100 ( .A1(n32750), .A2(n3748), .ZN(n33568) );
  INV_X1 U16101 ( .I(n13648), .ZN(n23068) );
  INV_X2 U16105 ( .I(n4580), .ZN(n23070) );
  NAND2_X1 U16107 ( .A1(n11754), .A2(n30505), .ZN(n14530) );
  CLKBUF_X4 U16108 ( .I(n8374), .Z(n2879) );
  NOR2_X1 U16109 ( .A1(n25296), .A2(n16650), .ZN(n28186) );
  AND2_X2 U16110 ( .A1(n2570), .A2(n30403), .Z(n32865) );
  NOR2_X1 U16114 ( .A1(n987), .A2(n22957), .ZN(n22901) );
  BUF_X2 U16115 ( .I(n17947), .Z(n29695) );
  AND2_X2 U16116 ( .A1(n25409), .A2(n15496), .Z(n25329) );
  NOR2_X1 U16117 ( .A1(n25995), .A2(n14737), .ZN(n7272) );
  NAND2_X1 U16120 ( .A1(n22886), .A2(n23093), .ZN(n13618) );
  NAND3_X1 U16123 ( .A1(n10376), .A2(n789), .A3(n13684), .ZN(n25727) );
  OAI21_X1 U16130 ( .A1(n25731), .A2(n16494), .B(n10376), .ZN(n1896) );
  CLKBUF_X4 U16140 ( .I(n25145), .Z(n29976) );
  NAND2_X1 U16141 ( .A1(n14972), .A2(n25973), .ZN(n28703) );
  NAND2_X1 U16144 ( .A1(n2456), .A2(n25234), .ZN(n8841) );
  NAND2_X1 U16145 ( .A1(n8784), .A2(n21579), .ZN(n3472) );
  OAI22_X1 U16146 ( .A1(n19010), .A2(n17445), .B1(n944), .B2(n17444), .ZN(
        n27460) );
  OR2_X2 U16164 ( .A1(n944), .A2(n18913), .Z(n5139) );
  OR2_X1 U16166 ( .A1(n8412), .A2(n29306), .Z(n15537) );
  AND3_X2 U16167 ( .A1(n30930), .A2(n30555), .A3(n28217), .Z(n32867) );
  NAND3_X1 U16173 ( .A1(n753), .A2(n17717), .A3(n28136), .ZN(n30555) );
  NAND3_X1 U16175 ( .A1(n29388), .A2(n33680), .A3(n33540), .ZN(n1475) );
  NAND2_X1 U16185 ( .A1(n25058), .A2(n25044), .ZN(n25059) );
  INV_X1 U16187 ( .I(n22856), .ZN(n986) );
  NAND2_X1 U16188 ( .A1(n13859), .A2(n6275), .ZN(n3940) );
  CLKBUF_X2 U16189 ( .I(n9133), .Z(n33147) );
  NOR2_X1 U16192 ( .A1(n19058), .A2(n945), .ZN(n5709) );
  AOI21_X1 U16193 ( .A1(n9982), .A2(n25615), .B(n10174), .ZN(n9981) );
  OAI21_X1 U16199 ( .A1(n21642), .A2(n21651), .B(n31511), .ZN(n21555) );
  INV_X1 U16202 ( .I(n24289), .ZN(n15977) );
  NOR2_X1 U16204 ( .A1(n21358), .A2(n5018), .ZN(n28882) );
  INV_X2 U16205 ( .I(n21358), .ZN(n1140) );
  AND3_X1 U16216 ( .A1(n16254), .A2(n23109), .A3(n23111), .Z(n78) );
  NOR2_X2 U16227 ( .A1(n31795), .A2(n28853), .ZN(n13006) );
  NAND2_X1 U16229 ( .A1(n23052), .A2(n23051), .ZN(n4006) );
  AOI21_X1 U16237 ( .A1(n1108), .A2(n23052), .B(n25994), .ZN(n4487) );
  NAND2_X1 U16239 ( .A1(n23052), .A2(n23053), .ZN(n1745) );
  OAI21_X1 U16244 ( .A1(n16054), .A2(n23052), .B(n31129), .ZN(n9949) );
  INV_X2 U16245 ( .I(n15038), .ZN(n9736) );
  INV_X2 U16256 ( .I(n16589), .ZN(n25187) );
  OAI21_X1 U16257 ( .A1(n25235), .A2(n8219), .B(n16589), .ZN(n3729) );
  INV_X2 U16258 ( .I(n25563), .ZN(n765) );
  INV_X1 U16261 ( .I(n25563), .ZN(n33394) );
  NAND2_X1 U16271 ( .A1(n25592), .A2(n25624), .ZN(n8854) );
  NOR2_X2 U16277 ( .A1(n25429), .A2(n11640), .ZN(n408) );
  NAND2_X1 U16278 ( .A1(n6662), .A2(n15600), .ZN(n7034) );
  NAND3_X1 U16279 ( .A1(n33078), .A2(n19180), .A3(n19178), .ZN(n13011) );
  AOI22_X1 U16281 ( .A1(n19177), .A2(n19180), .B1(n18114), .B2(n784), .ZN(
        n2126) );
  CLKBUF_X4 U16283 ( .I(n25903), .Z(n28455) );
  OAI21_X1 U16288 ( .A1(n25180), .A2(n25179), .B(n33428), .ZN(n25181) );
  OAI22_X1 U16289 ( .A1(n21159), .A2(n26133), .B1(n21158), .B2(n1020), .ZN(
        n28038) );
  OAI21_X1 U16294 ( .A1(n33507), .A2(n715), .B(n15462), .ZN(n7303) );
  NOR3_X1 U16302 ( .A1(n5926), .A2(n25571), .A3(n27113), .ZN(n30200) );
  NAND3_X1 U16303 ( .A1(n13660), .A2(n11937), .A3(n24198), .ZN(n17494) );
  CLKBUF_X12 U16305 ( .I(n22602), .Z(n16665) );
  NAND2_X1 U16310 ( .A1(n33107), .A2(n20419), .ZN(n10322) );
  NAND2_X1 U16315 ( .A1(n24056), .A2(n24002), .ZN(n24162) );
  INV_X2 U16318 ( .I(n24056), .ZN(n29566) );
  NAND2_X2 U16320 ( .A1(n21909), .A2(n32021), .ZN(n22730) );
  OR2_X2 U16323 ( .A1(n21688), .A2(n12561), .Z(n27073) );
  NAND2_X1 U16329 ( .A1(n28839), .A2(n13063), .ZN(n5374) );
  NAND2_X1 U16333 ( .A1(n12904), .A2(n18146), .ZN(n24144) );
  XNOR2_X1 U16334 ( .A1(n5023), .A2(n5022), .ZN(n32873) );
  OAI21_X1 U16338 ( .A1(n7334), .A2(n5713), .B(n25107), .ZN(n32909) );
  NAND2_X1 U16340 ( .A1(n8926), .A2(n25174), .ZN(n8925) );
  NAND3_X2 U16341 ( .A1(n1213), .A2(n9162), .A3(n6034), .ZN(n25138) );
  CLKBUF_X4 U16348 ( .I(n10943), .Z(n34005) );
  INV_X1 U16356 ( .I(n13349), .ZN(n33598) );
  OAI21_X1 U16360 ( .A1(n21162), .A2(n21161), .B(n21139), .ZN(n21140) );
  NAND2_X1 U16363 ( .A1(n21466), .A2(n31085), .ZN(n9666) );
  XNOR2_X1 U16365 ( .A1(n30749), .A2(n10332), .ZN(n20967) );
  INV_X1 U16366 ( .I(n10332), .ZN(n1345) );
  INV_X2 U16370 ( .I(n1294), .ZN(n13703) );
  AOI21_X1 U16371 ( .A1(n24718), .A2(n12266), .B(n11735), .ZN(n17304) );
  NAND2_X1 U16378 ( .A1(n20427), .A2(n12421), .ZN(n14620) );
  NAND2_X1 U16379 ( .A1(n28376), .A2(n12421), .ZN(n19827) );
  AOI21_X1 U16382 ( .A1(n12482), .A2(n12247), .B(n15274), .ZN(n11759) );
  XOR2_X1 U16390 ( .A1(n16989), .A2(n27896), .Z(n32875) );
  INV_X1 U16394 ( .I(n221), .ZN(n32876) );
  NOR2_X1 U16399 ( .A1(n24339), .A2(n24056), .ZN(n29018) );
  INV_X2 U16401 ( .I(n25176), .ZN(n16273) );
  NOR2_X1 U16402 ( .A1(n33353), .A2(n25257), .ZN(n32954) );
  XNOR2_X1 U16404 ( .A1(n24826), .A2(n24532), .ZN(n24673) );
  AND2_X2 U16416 ( .A1(n29681), .A2(n30802), .Z(n32879) );
  NAND2_X2 U16417 ( .A1(n33443), .A2(n33442), .ZN(n30802) );
  NAND2_X1 U16418 ( .A1(n33126), .A2(n11382), .ZN(n32880) );
  XOR2_X1 U16425 ( .A1(n13504), .A2(n12749), .Z(n32883) );
  INV_X1 U16426 ( .I(n5118), .ZN(n19011) );
  AOI21_X1 U16429 ( .A1(n22899), .A2(n22592), .B(n22705), .ZN(n10896) );
  INV_X1 U16430 ( .I(n12238), .ZN(n10126) );
  AOI21_X1 U16431 ( .A1(n32869), .A2(n25444), .B(n31263), .ZN(n15498) );
  NAND2_X2 U16435 ( .A1(n33243), .A2(n33644), .ZN(n32885) );
  XNOR2_X1 U16436 ( .A1(n32885), .A2(n10075), .ZN(n30671) );
  NAND2_X1 U16438 ( .A1(n33243), .A2(n33644), .ZN(n22059) );
  INV_X2 U16441 ( .I(n25175), .ZN(n14531) );
  INV_X1 U16450 ( .I(n19899), .ZN(n20033) );
  INV_X1 U16463 ( .I(n20577), .ZN(n32989) );
  NOR2_X1 U16464 ( .A1(n20312), .A2(n20577), .ZN(n17647) );
  NAND2_X1 U16470 ( .A1(n4396), .A2(n33281), .ZN(n33280) );
  OAI21_X1 U16474 ( .A1(n22558), .A2(n4396), .B(n9630), .ZN(n32955) );
  INV_X1 U16476 ( .I(n4396), .ZN(n22671) );
  OAI21_X1 U16484 ( .A1(n1140), .A2(n30267), .B(n11967), .ZN(n21273) );
  NOR2_X1 U16489 ( .A1(n12037), .A2(n11967), .ZN(n12492) );
  INV_X2 U16490 ( .I(n11967), .ZN(n1331) );
  INV_X1 U16491 ( .I(n7699), .ZN(n10142) );
  NAND2_X1 U16493 ( .A1(n20494), .A2(n17497), .ZN(n5779) );
  INV_X2 U16501 ( .I(n17497), .ZN(n20268) );
  NOR3_X1 U16502 ( .A1(n27752), .A2(n30293), .A3(n28680), .ZN(n13431) );
  OAI22_X1 U16506 ( .A1(n6074), .A2(n14012), .B1(n16127), .B2(n32073), .ZN(
        n21600) );
  OAI21_X1 U16510 ( .A1(n30318), .A2(n3489), .B(n747), .ZN(n7341) );
  AND2_X1 U16511 ( .A1(n26551), .A2(n3816), .Z(n19944) );
  INV_X1 U16514 ( .I(n22138), .ZN(n16210) );
  INV_X1 U16517 ( .I(n23813), .ZN(n23852) );
  CLKBUF_X12 U16521 ( .I(n11845), .Z(n26545) );
  NAND2_X1 U16524 ( .A1(n230), .A2(n21512), .ZN(n5787) );
  INV_X1 U16527 ( .I(n10219), .ZN(n33200) );
  NAND2_X1 U16528 ( .A1(n31566), .A2(n3007), .ZN(n23058) );
  NAND3_X1 U16530 ( .A1(n21392), .A2(n17522), .A3(n21163), .ZN(n4784) );
  AOI21_X1 U16535 ( .A1(n21163), .A2(n21392), .B(n17522), .ZN(n2604) );
  XNOR2_X1 U16538 ( .A1(Plaintext[31]), .A2(Key[31]), .ZN(n18139) );
  OAI21_X1 U16539 ( .A1(n20533), .A2(n20463), .B(n28028), .ZN(n4077) );
  XOR2_X1 U16540 ( .A1(n17498), .A2(n6397), .Z(n32886) );
  AOI21_X2 U16542 ( .A1(n5810), .A2(n8186), .B(n32992), .ZN(n32887) );
  INV_X1 U16544 ( .I(n24276), .ZN(n34137) );
  AOI21_X1 U16551 ( .A1(n3984), .A2(n24276), .B(n7068), .ZN(n24169) );
  AND2_X1 U16552 ( .A1(n31939), .A2(n9486), .Z(n7065) );
  AOI21_X1 U16557 ( .A1(n6662), .A2(n26115), .B(n5191), .ZN(n13906) );
  NAND2_X1 U16561 ( .A1(n24002), .A2(n2826), .ZN(n7171) );
  NOR2_X1 U16565 ( .A1(n25806), .A2(n25820), .ZN(n25817) );
  INV_X2 U16566 ( .I(n9126), .ZN(n16113) );
  NOR2_X1 U16572 ( .A1(n10967), .A2(n23862), .ZN(n30736) );
  INV_X1 U16575 ( .I(n23862), .ZN(n13031) );
  INV_X2 U16576 ( .I(n9252), .ZN(n580) );
  AND2_X1 U16577 ( .A1(n14600), .A2(n15299), .Z(n10405) );
  INV_X2 U16579 ( .I(n32096), .ZN(n25391) );
  AOI21_X1 U16581 ( .A1(n794), .A2(n4604), .B(n11049), .ZN(n13552) );
  NAND2_X1 U16593 ( .A1(n33857), .A2(n17888), .ZN(n27707) );
  NAND3_X1 U16594 ( .A1(n25043), .A2(n25062), .A3(n25042), .ZN(n28220) );
  NAND3_X1 U16595 ( .A1(n25731), .A2(n25724), .A3(n13640), .ZN(n25725) );
  INV_X2 U16596 ( .I(n23888), .ZN(n23887) );
  CLKBUF_X4 U16602 ( .I(n23888), .Z(n29240) );
  NOR2_X1 U16612 ( .A1(n9405), .A2(n21452), .ZN(n9324) );
  NOR2_X1 U16618 ( .A1(n7291), .A2(n7852), .ZN(n20397) );
  XOR2_X1 U16619 ( .A1(n27976), .A2(n30016), .Z(n32888) );
  AND3_X2 U16620 ( .A1(n7279), .A2(n14161), .A3(n20627), .Z(n31291) );
  AOI21_X1 U16624 ( .A1(n28736), .A2(n14810), .B(n788), .ZN(n8723) );
  INV_X2 U16629 ( .I(n16981), .ZN(n14232) );
  NAND2_X1 U16631 ( .A1(n16981), .A2(n11096), .ZN(n15616) );
  NOR2_X1 U16632 ( .A1(n30584), .A2(n3909), .ZN(n8083) );
  INV_X1 U16633 ( .I(n32452), .ZN(n7044) );
  OAI21_X1 U16637 ( .A1(n27685), .A2(n30832), .B(n9472), .ZN(n5495) );
  OAI21_X1 U16650 ( .A1(n5863), .A2(n7811), .B(n21872), .ZN(n12390) );
  NAND2_X1 U16655 ( .A1(n5863), .A2(n9472), .ZN(n12354) );
  NOR2_X1 U16660 ( .A1(n17720), .A2(n32858), .ZN(n12107) );
  INV_X2 U16661 ( .I(n17720), .ZN(n15601) );
  CLKBUF_X4 U16662 ( .I(n16798), .Z(n8766) );
  INV_X2 U16663 ( .I(n16798), .ZN(n749) );
  INV_X1 U16664 ( .I(n10858), .ZN(n25193) );
  NAND2_X1 U16665 ( .A1(n19320), .A2(n19274), .ZN(n33389) );
  NAND2_X1 U16666 ( .A1(n29317), .A2(n4908), .ZN(n8954) );
  NAND2_X1 U16667 ( .A1(n29317), .A2(n13694), .ZN(n23072) );
  AOI21_X1 U16669 ( .A1(n916), .A2(n196), .B(n11755), .ZN(n9898) );
  AOI21_X1 U16673 ( .A1(n5850), .A2(n27954), .B(n11755), .ZN(n5849) );
  INV_X1 U16676 ( .I(n17305), .ZN(n32907) );
  NAND2_X1 U16677 ( .A1(n21161), .A2(n17305), .ZN(n7050) );
  INV_X1 U16678 ( .I(n3286), .ZN(n17644) );
  INV_X2 U16679 ( .I(n12657), .ZN(n5371) );
  NAND2_X1 U16687 ( .A1(n13574), .A2(n29173), .ZN(n1561) );
  CLKBUF_X12 U16692 ( .I(n2655), .Z(n123) );
  AOI21_X1 U16694 ( .A1(n13059), .A2(n14811), .B(n12548), .ZN(n6188) );
  BUF_X2 U16695 ( .I(n18076), .Z(n11097) );
  INV_X1 U16700 ( .I(n18076), .ZN(n31669) );
  INV_X1 U16705 ( .I(n18861), .ZN(n18863) );
  XOR2_X1 U16706 ( .A1(n30767), .A2(n7071), .Z(n32890) );
  NAND3_X1 U16707 ( .A1(n14752), .A2(n10755), .A3(n27248), .ZN(n24365) );
  INV_X2 U16710 ( .I(n22979), .ZN(n31531) );
  NAND2_X1 U16712 ( .A1(n22978), .A2(n22979), .ZN(n28348) );
  OR2_X2 U16721 ( .A1(n29908), .A2(n11364), .Z(n3005) );
  NAND2_X1 U16722 ( .A1(n3169), .A2(n17150), .ZN(n12848) );
  OR2_X1 U16727 ( .A1(n28811), .A2(n16776), .Z(n23728) );
  OAI21_X1 U16729 ( .A1(n25987), .A2(n16776), .B(n23728), .ZN(n17134) );
  INV_X1 U16733 ( .I(n30045), .ZN(n32892) );
  OR2_X2 U16734 ( .A1(n32891), .A2(n8327), .Z(n6109) );
  OR2_X1 U16735 ( .A1(n31922), .A2(n32891), .Z(n9033) );
  NAND2_X1 U16736 ( .A1(n535), .A2(n23197), .ZN(n23804) );
  AOI21_X2 U16740 ( .A1(n23006), .A2(n3999), .B(n23004), .ZN(n32893) );
  AOI21_X2 U16741 ( .A1(n16883), .A2(n20220), .B(n30530), .ZN(n32894) );
  XOR2_X1 U16745 ( .A1(n22970), .A2(n23375), .Z(n32895) );
  NOR3_X1 U16749 ( .A1(n15139), .A2(n18006), .A3(n18007), .ZN(n18005) );
  INV_X1 U16757 ( .I(n14132), .ZN(n9568) );
  CLKBUF_X12 U16759 ( .I(n16309), .Z(n26766) );
  OAI21_X1 U16761 ( .A1(n14627), .A2(n17987), .B(n15641), .ZN(n15331) );
  NOR2_X1 U16764 ( .A1(n4897), .A2(n15227), .ZN(n27963) );
  AOI21_X1 U16766 ( .A1(n9687), .A2(n14490), .B(n4897), .ZN(n33390) );
  INV_X2 U16767 ( .I(n10612), .ZN(n31345) );
  INV_X1 U16772 ( .I(n837), .ZN(n32896) );
  NAND2_X2 U16774 ( .A1(n6656), .A2(n26614), .ZN(n32897) );
  NAND2_X1 U16776 ( .A1(n6656), .A2(n26614), .ZN(n25515) );
  NAND2_X2 U16778 ( .A1(n24864), .A2(n16397), .ZN(n6656) );
  NOR2_X2 U16780 ( .A1(n8149), .A2(n8150), .ZN(n32899) );
  OAI21_X1 U16782 ( .A1(n33850), .A2(n9393), .B(n9392), .ZN(n8323) );
  INV_X2 U16785 ( .I(n1877), .ZN(n31522) );
  BUF_X2 U16786 ( .I(n8088), .Z(n28737) );
  NOR2_X1 U16787 ( .A1(n723), .A2(n31325), .ZN(n11564) );
  NAND2_X1 U16789 ( .A1(n27719), .A2(n31325), .ZN(n10884) );
  NAND2_X1 U16799 ( .A1(n723), .A2(n31325), .ZN(n3830) );
  INV_X1 U16801 ( .I(n24803), .ZN(n33100) );
  NOR2_X1 U16803 ( .A1(n1269), .A2(n7287), .ZN(n2579) );
  AND2_X2 U16809 ( .A1(n27880), .A2(n1284), .Z(n27889) );
  CLKBUF_X12 U16815 ( .I(n7881), .Z(n28689) );
  NOR2_X1 U16816 ( .A1(n32595), .A2(n7881), .ZN(n16560) );
  NAND2_X1 U16830 ( .A1(n14133), .A2(n29472), .ZN(n23958) );
  INV_X1 U16831 ( .I(n25790), .ZN(n16422) );
  INV_X2 U16836 ( .I(n25790), .ZN(n25788) );
  NAND2_X1 U16838 ( .A1(n24062), .A2(n30651), .ZN(n6287) );
  NOR3_X1 U16841 ( .A1(n796), .A2(n30651), .A3(n24207), .ZN(n10652) );
  INV_X1 U16845 ( .I(n30651), .ZN(n970) );
  NAND2_X1 U16849 ( .A1(n7778), .A2(n9220), .ZN(n5673) );
  NAND2_X1 U16850 ( .A1(n25515), .A2(n6595), .ZN(n25510) );
  NOR2_X1 U16852 ( .A1(n22951), .A2(n13762), .ZN(n3202) );
  NOR2_X1 U16854 ( .A1(n2654), .A2(n5454), .ZN(n9581) );
  CLKBUF_X4 U16861 ( .I(n5454), .Z(n31461) );
  OR2_X2 U16863 ( .A1(n22565), .A2(n14676), .Z(n22680) );
  NAND3_X1 U16867 ( .A1(n25804), .A2(n25818), .A3(n11003), .ZN(n18246) );
  AOI22_X1 U16871 ( .A1(n25807), .A2(n25816), .B1(n25804), .B2(n25817), .ZN(
        n14009) );
  NAND2_X1 U16873 ( .A1(n15340), .A2(n28358), .ZN(n33507) );
  NOR2_X1 U16875 ( .A1(n28358), .A2(n15340), .ZN(n25207) );
  NAND2_X1 U16876 ( .A1(n3581), .A2(n30333), .ZN(n33227) );
  INV_X1 U16880 ( .I(n30333), .ZN(n34039) );
  NOR2_X1 U16892 ( .A1(n31263), .A2(n17948), .ZN(n25432) );
  NAND2_X1 U16894 ( .A1(n17948), .A2(n25437), .ZN(n25445) );
  INV_X1 U16902 ( .I(n17948), .ZN(n25425) );
  OAI21_X2 U16910 ( .A1(n6204), .A2(n28706), .B(n24889), .ZN(n32900) );
  INV_X1 U16914 ( .I(n9301), .ZN(n33681) );
  XOR2_X1 U16916 ( .A1(Plaintext[110]), .A2(Key[110]), .Z(n32901) );
  XOR2_X1 U16917 ( .A1(n10707), .A2(n27766), .Z(n32902) );
  OR2_X1 U16918 ( .A1(n23018), .A2(n9575), .Z(n13274) );
  NAND2_X1 U16927 ( .A1(n21811), .A2(n8140), .ZN(n15774) );
  OAI22_X2 U16928 ( .A1(n3866), .A2(n3867), .B1(n6568), .B2(n10096), .ZN(
        n32904) );
  OR2_X2 U16930 ( .A1(n32904), .A2(n21601), .Z(n6238) );
  CLKBUF_X12 U16931 ( .I(n31497), .Z(n31113) );
  AOI21_X1 U16932 ( .A1(n2444), .A2(n24216), .B(n31497), .ZN(n10047) );
  NOR2_X1 U16934 ( .A1(n889), .A2(n31497), .ZN(n6225) );
  AND3_X2 U16936 ( .A1(n25975), .A2(n21715), .A3(n5704), .Z(n9591) );
  NOR2_X1 U16937 ( .A1(n8270), .A2(n843), .ZN(n23788) );
  XOR2_X1 U16938 ( .A1(n17400), .A2(n32050), .Z(n32905) );
  AOI22_X2 U16941 ( .A1(n32010), .A2(n4110), .B1(n31942), .B2(n22383), .ZN(
        n8418) );
  XOR2_X1 U16942 ( .A1(n23475), .A2(n23417), .Z(n32906) );
  XOR2_X1 U16943 ( .A1(n22231), .A2(n22303), .Z(n30402) );
  NAND2_X2 U16949 ( .A1(n15847), .A2(n15846), .ZN(n22231) );
  XOR2_X1 U16951 ( .A1(n22240), .A2(n22197), .Z(n22167) );
  NOR2_X2 U16953 ( .A1(n21600), .A2(n21599), .ZN(n22240) );
  INV_X4 U16954 ( .I(n7892), .ZN(n20607) );
  XNOR2_X1 U16959 ( .A1(n33952), .A2(n31116), .ZN(n8434) );
  AOI22_X1 U16961 ( .A1(n25367), .A2(n30302), .B1(n3300), .B2(n25376), .ZN(
        n25380) );
  XOR2_X1 U16964 ( .A1(n19497), .A2(n17931), .Z(n12653) );
  NAND2_X2 U16967 ( .A1(n7647), .A2(n6494), .ZN(n5713) );
  NAND2_X2 U16969 ( .A1(n31309), .A2(n5228), .ZN(n21933) );
  NAND2_X1 U16971 ( .A1(n21213), .A2(n32907), .ZN(n17375) );
  NOR2_X2 U16974 ( .A1(n21160), .A2(n32902), .ZN(n21213) );
  INV_X2 U16975 ( .I(n20472), .ZN(n20317) );
  NAND2_X2 U16978 ( .A1(n19382), .A2(n27196), .ZN(n20472) );
  NOR2_X1 U16982 ( .A1(n1018), .A2(n21358), .ZN(n27828) );
  XOR2_X1 U16987 ( .A1(n29833), .A2(n33311), .Z(n1018) );
  XOR2_X1 U16999 ( .A1(n23367), .A2(n15941), .Z(n10758) );
  NOR2_X2 U17001 ( .A1(n31823), .A2(n16298), .ZN(n19759) );
  INV_X2 U17004 ( .I(n32910), .ZN(n28602) );
  INV_X2 U17006 ( .I(n560), .ZN(n32911) );
  XOR2_X1 U17007 ( .A1(n32912), .A2(n10064), .Z(n8277) );
  XOR2_X1 U17009 ( .A1(n27667), .A2(n10459), .Z(n32912) );
  NAND3_X2 U17011 ( .A1(n17108), .A2(n32913), .A3(n30151), .ZN(n25665) );
  NAND2_X2 U17014 ( .A1(n3774), .A2(n755), .ZN(n32913) );
  XOR2_X1 U17017 ( .A1(n32914), .A2(n14527), .Z(n15433) );
  NAND2_X1 U17023 ( .A1(n32086), .A2(n2226), .ZN(n2225) );
  INV_X1 U17025 ( .I(n13472), .ZN(n969) );
  NAND2_X2 U17028 ( .A1(n7613), .A2(n29788), .ZN(n13472) );
  XOR2_X1 U17029 ( .A1(n13794), .A2(n13792), .Z(n17037) );
  NAND2_X2 U17040 ( .A1(n17639), .A2(n22814), .ZN(n17085) );
  INV_X2 U17045 ( .I(n19908), .ZN(n870) );
  NAND2_X1 U17047 ( .A1(n6549), .A2(n3967), .ZN(n19908) );
  XOR2_X1 U17051 ( .A1(n33348), .A2(n33588), .Z(n32916) );
  INV_X2 U17061 ( .I(n32919), .ZN(n8469) );
  XOR2_X1 U17063 ( .A1(n32921), .A2(n2651), .Z(n28611) );
  XOR2_X1 U17065 ( .A1(n2653), .A2(n32922), .Z(n32921) );
  AOI21_X1 U17069 ( .A1(n28715), .A2(n24340), .B(n16552), .ZN(n14847) );
  INV_X1 U17071 ( .I(n2653), .ZN(n1865) );
  XOR2_X1 U17078 ( .A1(n31499), .A2(n29927), .Z(n2653) );
  NAND3_X2 U17082 ( .A1(n23772), .A2(n33668), .A3(n15402), .ZN(n7093) );
  XOR2_X1 U17084 ( .A1(n32923), .A2(n21014), .Z(n12557) );
  XOR2_X1 U17085 ( .A1(n13681), .A2(n12559), .Z(n32923) );
  NOR2_X1 U17086 ( .A1(n16868), .A2(n24254), .ZN(n17802) );
  XOR2_X1 U17093 ( .A1(n31133), .A2(n22250), .Z(n27693) );
  XOR2_X1 U17094 ( .A1(n31081), .A2(n23490), .Z(n28847) );
  INV_X2 U17095 ( .I(n32924), .ZN(n7513) );
  XOR2_X1 U17096 ( .A1(n32925), .A2(n10052), .Z(n31844) );
  NOR2_X2 U17104 ( .A1(n32045), .A2(n1291), .ZN(n7398) );
  XOR2_X1 U17105 ( .A1(n5703), .A2(n4173), .Z(n4718) );
  NAND2_X2 U17109 ( .A1(n24496), .A2(n24495), .ZN(n24498) );
  NAND2_X2 U17110 ( .A1(n12753), .A2(n32927), .ZN(n12785) );
  NAND3_X2 U17111 ( .A1(n15494), .A2(n12788), .A3(n7813), .ZN(n32927) );
  XOR2_X1 U17121 ( .A1(n12637), .A2(n32928), .Z(n17117) );
  XOR2_X1 U17124 ( .A1(n12636), .A2(n13309), .Z(n32928) );
  NOR2_X1 U17128 ( .A1(n1379), .A2(n19132), .ZN(n7418) );
  NAND2_X1 U17129 ( .A1(n4405), .A2(n19249), .ZN(n19132) );
  XOR2_X1 U17133 ( .A1(n10902), .A2(n32930), .Z(n33770) );
  XOR2_X1 U17135 ( .A1(n27098), .A2(n19654), .Z(n10902) );
  XOR2_X1 U17138 ( .A1(n10006), .A2(n22274), .Z(n22084) );
  INV_X2 U17140 ( .I(n21925), .ZN(n10006) );
  OAI21_X1 U17150 ( .A1(n28388), .A2(n10835), .B(n692), .ZN(n27342) );
  NAND2_X2 U17151 ( .A1(n33560), .A2(n27676), .ZN(n24008) );
  NAND2_X1 U17158 ( .A1(n32931), .A2(n17087), .ZN(n23927) );
  AOI22_X2 U17159 ( .A1(n11971), .A2(n20154), .B1(n20153), .B2(n8259), .ZN(
        n4420) );
  NOR2_X2 U17160 ( .A1(n19914), .A2(n31951), .ZN(n11971) );
  NOR2_X1 U17161 ( .A1(n31915), .A2(n26641), .ZN(n29037) );
  OAI21_X2 U17166 ( .A1(n31962), .A2(n24557), .B(n32933), .ZN(n25285) );
  AOI22_X1 U17168 ( .A1(n20076), .A2(n12408), .B1(n6444), .B2(n2499), .ZN(
        n3624) );
  NAND2_X1 U17169 ( .A1(n2654), .A2(n5454), .ZN(n8664) );
  OAI21_X1 U17171 ( .A1(n16474), .A2(n28344), .B(n18805), .ZN(n26909) );
  AOI22_X2 U17174 ( .A1(n32062), .A2(n32934), .B1(n24308), .B2(n24135), .ZN(
        n11830) );
  INV_X2 U17177 ( .I(n23714), .ZN(n32934) );
  XOR2_X1 U17181 ( .A1(n14781), .A2(n14783), .Z(n16603) );
  AND3_X1 U17182 ( .A1(n28641), .A2(n5595), .A3(n21223), .Z(n33352) );
  NAND2_X2 U17185 ( .A1(n1700), .A2(n32920), .ZN(n15768) );
  INV_X2 U17186 ( .I(n22108), .ZN(n7725) );
  NAND2_X2 U17187 ( .A1(n8078), .A2(n8077), .ZN(n22108) );
  XOR2_X1 U17188 ( .A1(n32937), .A2(n33017), .Z(n28615) );
  XOR2_X1 U17189 ( .A1(n23330), .A2(n23277), .Z(n32937) );
  INV_X2 U17198 ( .I(n32938), .ZN(n15722) );
  XNOR2_X1 U17202 ( .A1(n15507), .A2(n23377), .ZN(n32938) );
  INV_X2 U17205 ( .I(n20531), .ZN(n32940) );
  INV_X1 U17206 ( .I(n28064), .ZN(n32941) );
  OAI21_X2 U17208 ( .A1(n28786), .A2(n1170), .B(n33241), .ZN(n28064) );
  OAI21_X2 U17211 ( .A1(n10621), .A2(n10620), .B(n32942), .ZN(n10281) );
  AND2_X1 U17212 ( .A1(n5274), .A2(n8365), .Z(n26195) );
  NAND2_X2 U17215 ( .A1(n17008), .A2(n17006), .ZN(n5274) );
  NAND2_X2 U17217 ( .A1(n10760), .A2(n10759), .ZN(n15941) );
  NAND2_X2 U17218 ( .A1(n19310), .A2(n10828), .ZN(n18667) );
  AOI21_X2 U17221 ( .A1(n7662), .A2(n6366), .B(n32943), .ZN(n7660) );
  INV_X2 U17222 ( .I(n32945), .ZN(n3193) );
  XOR2_X1 U17224 ( .A1(n3298), .A2(n509), .Z(n32945) );
  XOR2_X1 U17225 ( .A1(n15360), .A2(n11193), .Z(n16998) );
  NOR2_X2 U17230 ( .A1(n22556), .A2(n15362), .ZN(n15360) );
  XOR2_X1 U17231 ( .A1(n10516), .A2(n2074), .Z(n10514) );
  NAND2_X1 U17235 ( .A1(n14633), .A2(n33701), .ZN(Ciphertext[57]) );
  NAND2_X2 U17242 ( .A1(n30870), .A2(n5092), .ZN(n13415) );
  XOR2_X1 U17248 ( .A1(n30284), .A2(n22123), .Z(n1971) );
  NAND2_X2 U17252 ( .A1(n12997), .A2(n14907), .ZN(n12982) );
  NAND2_X2 U17255 ( .A1(n29368), .A2(n30409), .ZN(n12997) );
  XOR2_X1 U17256 ( .A1(n15373), .A2(n17051), .Z(n33303) );
  NAND2_X2 U17257 ( .A1(n33987), .A2(n32946), .ZN(n25106) );
  NAND2_X1 U17260 ( .A1(n15331), .A2(n15332), .ZN(n32946) );
  XOR2_X1 U17261 ( .A1(n24674), .A2(n24673), .Z(n24679) );
  NAND2_X2 U17265 ( .A1(n1749), .A2(n29982), .ZN(n23052) );
  XOR2_X1 U17266 ( .A1(n32947), .A2(n22040), .Z(n22535) );
  INV_X2 U17267 ( .I(n13623), .ZN(n7361) );
  NAND4_X2 U17270 ( .A1(n3744), .A2(n7075), .A3(n7074), .A4(n7076), .ZN(n13623) );
  XOR2_X1 U17272 ( .A1(n23324), .A2(n32948), .Z(n11225) );
  XOR2_X1 U17274 ( .A1(n11227), .A2(n29082), .Z(n32948) );
  INV_X2 U17276 ( .I(n3250), .ZN(n32949) );
  NAND2_X2 U17280 ( .A1(n28581), .A2(n15302), .ZN(n3250) );
  OAI21_X2 U17281 ( .A1(n28096), .A2(n18151), .B(n32950), .ZN(n12856) );
  XOR2_X1 U17283 ( .A1(n5932), .A2(n6547), .Z(n15674) );
  NAND2_X2 U17290 ( .A1(n5933), .A2(n5935), .ZN(n5932) );
  XOR2_X1 U17291 ( .A1(n12310), .A2(n23388), .Z(n23220) );
  NAND3_X2 U17292 ( .A1(n12180), .A2(n5136), .A3(n9918), .ZN(n12310) );
  NAND2_X2 U17296 ( .A1(n4571), .A2(n9835), .ZN(n29781) );
  NOR2_X1 U17305 ( .A1(n16041), .A2(n25322), .ZN(n6234) );
  NAND3_X2 U17308 ( .A1(n30930), .A2(n30555), .A3(n28217), .ZN(n25322) );
  NAND2_X2 U17310 ( .A1(n23101), .A2(n11956), .ZN(n22783) );
  NAND2_X1 U17311 ( .A1(n32954), .A2(n11569), .ZN(n107) );
  OAI22_X2 U17319 ( .A1(n24149), .A2(n32750), .B1(n9946), .B2(n24063), .ZN(
        n24064) );
  INV_X4 U17320 ( .I(n1775), .ZN(n9946) );
  NAND2_X2 U17325 ( .A1(n27064), .A2(n1776), .ZN(n1775) );
  NAND2_X2 U17329 ( .A1(n32956), .A2(n11505), .ZN(n7552) );
  BUF_X2 U17333 ( .I(n33153), .Z(n32957) );
  OR2_X1 U17335 ( .A1(n33942), .A2(n30200), .Z(n31489) );
  XOR2_X1 U17336 ( .A1(n23296), .A2(n17766), .Z(n26371) );
  XOR2_X1 U17338 ( .A1(n19741), .A2(n19625), .Z(n19571) );
  NOR2_X2 U17339 ( .A1(n30670), .A2(n30768), .ZN(n19741) );
  XOR2_X1 U17340 ( .A1(n32958), .A2(n24918), .Z(Ciphertext[5]) );
  AOI22_X1 U17343 ( .A1(n8278), .A2(n10099), .B1(n24915), .B2(n24916), .ZN(
        n32958) );
  XOR2_X1 U17345 ( .A1(n24356), .A2(n24370), .Z(n24390) );
  INV_X2 U17346 ( .I(n28415), .ZN(n32960) );
  XOR2_X1 U17349 ( .A1(n2435), .A2(n32961), .Z(n22350) );
  XOR2_X1 U17357 ( .A1(n21984), .A2(n29418), .Z(n32961) );
  NOR2_X2 U17359 ( .A1(n745), .A2(n17817), .ZN(n19195) );
  NAND2_X2 U17363 ( .A1(n33122), .A2(n12826), .ZN(n17817) );
  NAND3_X2 U17377 ( .A1(n32963), .A2(n32962), .A3(n363), .ZN(n16045) );
  NAND3_X2 U17379 ( .A1(n5367), .A2(n5366), .A3(n28833), .ZN(n32963) );
  NAND2_X2 U17381 ( .A1(n5124), .A2(n32965), .ZN(n16960) );
  AOI22_X2 U17383 ( .A1(n18578), .A2(n18855), .B1(n6873), .B2(n18854), .ZN(
        n32965) );
  XOR2_X1 U17388 ( .A1(n29209), .A2(n11416), .Z(n16384) );
  XOR2_X1 U17401 ( .A1(n32966), .A2(n15338), .Z(n15153) );
  XOR2_X1 U17402 ( .A1(n15337), .A2(n20818), .Z(n32966) );
  NAND3_X2 U17405 ( .A1(n24079), .A2(n24080), .A3(n24081), .ZN(n24083) );
  NAND2_X2 U17407 ( .A1(n18754), .A2(n15193), .ZN(n19386) );
  AND2_X1 U17408 ( .A1(n18830), .A2(n6256), .Z(n17054) );
  XOR2_X1 U17414 ( .A1(n31092), .A2(n30126), .Z(n27435) );
  NOR2_X2 U17422 ( .A1(n22894), .A2(n6605), .ZN(n33023) );
  NAND2_X2 U17429 ( .A1(n29608), .A2(n33982), .ZN(n6605) );
  OAI22_X2 U17432 ( .A1(n18901), .A2(n9787), .B1(n30995), .B2(n1378), .ZN(
        n5872) );
  NAND2_X2 U17435 ( .A1(n1378), .A2(n29146), .ZN(n18901) );
  NAND2_X1 U17436 ( .A1(n16372), .A2(n12863), .ZN(n12875) );
  XOR2_X1 U17442 ( .A1(n32968), .A2(n17918), .Z(n16618) );
  XOR2_X1 U17443 ( .A1(n13651), .A2(n22048), .Z(n32968) );
  XOR2_X1 U17445 ( .A1(n24793), .A2(n11217), .Z(n30393) );
  AOI21_X2 U17446 ( .A1(n32969), .A2(n11381), .B(n32013), .ZN(n22085) );
  OR2_X1 U17451 ( .A1(n31859), .A2(n31484), .Z(n32969) );
  OAI21_X2 U17457 ( .A1(n8991), .A2(n10138), .B(n10137), .ZN(n22978) );
  XOR2_X1 U17458 ( .A1(n31901), .A2(n17904), .Z(n3503) );
  XOR2_X1 U17462 ( .A1(n22252), .A2(n14796), .Z(n8993) );
  XOR2_X1 U17464 ( .A1(n21769), .A2(n32970), .Z(n29287) );
  XOR2_X1 U17471 ( .A1(n21921), .A2(n22242), .Z(n32970) );
  NAND2_X2 U17476 ( .A1(n33516), .A2(n32971), .ZN(n25806) );
  NAND3_X1 U17477 ( .A1(n13819), .A2(n1211), .A3(n24710), .ZN(n32971) );
  OAI21_X2 U17478 ( .A1(n32973), .A2(n23778), .B(n32972), .ZN(n23354) );
  NOR2_X2 U17480 ( .A1(n9181), .A2(n17642), .ZN(n25812) );
  AOI22_X2 U17483 ( .A1(n24102), .A2(n24101), .B1(n14375), .B2(n24103), .ZN(
        n33505) );
  AOI22_X2 U17486 ( .A1(n11003), .A2(n9181), .B1(n25818), .B2(n25823), .ZN(
        n25825) );
  NAND2_X1 U17487 ( .A1(n28256), .A2(n28255), .ZN(n33450) );
  XOR2_X1 U17488 ( .A1(n32974), .A2(n16622), .Z(Ciphertext[3]) );
  NAND2_X2 U17492 ( .A1(n14828), .A2(n16782), .ZN(n18830) );
  AND2_X1 U17494 ( .A1(n29139), .A2(n33175), .Z(n32986) );
  XOR2_X1 U17495 ( .A1(n32977), .A2(n24748), .Z(Ciphertext[4]) );
  XOR2_X1 U17496 ( .A1(n10210), .A2(n19504), .Z(n5862) );
  NOR2_X1 U17499 ( .A1(n33155), .A2(n25889), .ZN(n11735) );
  NOR2_X2 U17500 ( .A1(n32980), .A2(n32979), .ZN(n32978) );
  OR2_X1 U17502 ( .A1(n8412), .A2(n24271), .Z(n8499) );
  XOR2_X1 U17503 ( .A1(n12494), .A2(n32981), .Z(n516) );
  NAND2_X2 U17504 ( .A1(n8940), .A2(n29835), .ZN(n12494) );
  XOR2_X1 U17506 ( .A1(n23140), .A2(n33073), .Z(n23144) );
  NAND2_X2 U17507 ( .A1(n32983), .A2(n33667), .ZN(n22197) );
  XOR2_X1 U17511 ( .A1(n32984), .A2(n25104), .Z(Ciphertext[51]) );
  OAI21_X2 U17522 ( .A1(n1244), .A2(n889), .B(n24289), .ZN(n32985) );
  NAND3_X1 U17523 ( .A1(n8614), .A2(n3860), .A3(n33722), .ZN(n29964) );
  NOR2_X2 U17528 ( .A1(n15718), .A2(n22873), .ZN(n9460) );
  INV_X4 U17532 ( .I(n865), .ZN(n33888) );
  OAI22_X1 U17533 ( .A1(n22952), .A2(n13762), .B1(n6801), .B2(n22951), .ZN(
        n6674) );
  NAND2_X2 U17536 ( .A1(n23915), .A2(n13521), .ZN(n7991) );
  BUF_X4 U17544 ( .I(n11676), .Z(n33659) );
  NAND2_X2 U17546 ( .A1(n32987), .A2(n11746), .ZN(n22729) );
  AOI21_X2 U17548 ( .A1(n30658), .A2(n1726), .B(n32988), .ZN(n29610) );
  CLKBUF_X4 U17555 ( .I(n14290), .Z(n33641) );
  NAND2_X2 U17557 ( .A1(n30119), .A2(n19735), .ZN(n26566) );
  NAND2_X2 U17558 ( .A1(n7204), .A2(n7207), .ZN(n21579) );
  XOR2_X1 U17559 ( .A1(n9369), .A2(n22150), .Z(n4589) );
  AOI22_X2 U17560 ( .A1(n5912), .A2(n17261), .B1(n10188), .B2(n5913), .ZN(
        n33041) );
  NOR2_X2 U17561 ( .A1(n24004), .A2(n841), .ZN(n10188) );
  NAND3_X1 U17562 ( .A1(n5043), .A2(n28358), .A3(n15340), .ZN(n32990) );
  NAND2_X1 U17564 ( .A1(n23092), .A2(n13597), .ZN(n33931) );
  NAND2_X2 U17565 ( .A1(n12147), .A2(n12148), .ZN(n20955) );
  NOR2_X1 U17566 ( .A1(n23942), .A2(n11933), .ZN(n15451) );
  XOR2_X1 U17567 ( .A1(n283), .A2(n24801), .Z(n24649) );
  NAND2_X2 U17574 ( .A1(n6165), .A2(n30509), .ZN(n24801) );
  XOR2_X1 U17577 ( .A1(n27145), .A2(n24478), .Z(n24551) );
  NAND2_X1 U17580 ( .A1(n14184), .A2(n14724), .ZN(n27145) );
  XOR2_X1 U17581 ( .A1(n32991), .A2(n2739), .Z(n2859) );
  XOR2_X1 U17582 ( .A1(n20777), .A2(n10412), .Z(n32991) );
  NAND3_X2 U17585 ( .A1(n11952), .A2(n20042), .A3(n410), .ZN(n16248) );
  NAND2_X1 U17586 ( .A1(n27110), .A2(n1169), .ZN(n20039) );
  XOR2_X1 U17588 ( .A1(n1615), .A2(n1616), .Z(n27110) );
  OAI22_X2 U17589 ( .A1(n14547), .A2(n25708), .B1(n17092), .B2(n25752), .ZN(
        n32992) );
  AOI22_X2 U17591 ( .A1(n8587), .A2(n29207), .B1(n34059), .B2(n32993), .ZN(
        n2790) );
  NAND2_X1 U17594 ( .A1(n17522), .A2(n28607), .ZN(n32993) );
  NAND3_X2 U17597 ( .A1(n7276), .A2(n28995), .A3(n32994), .ZN(n22274) );
  AOI22_X2 U17599 ( .A1(n31935), .A2(n29242), .B1(n11330), .B2(n29314), .ZN(
        n32995) );
  XOR2_X1 U17600 ( .A1(n6348), .A2(n33465), .Z(n5703) );
  XNOR2_X1 U17602 ( .A1(n20859), .A2(n10081), .ZN(n5518) );
  XOR2_X1 U17604 ( .A1(n33234), .A2(n9141), .Z(n10081) );
  AOI21_X2 U17607 ( .A1(n20327), .A2(n20328), .B(n1149), .ZN(n32996) );
  INV_X2 U17611 ( .I(n28975), .ZN(n32998) );
  NOR2_X2 U17619 ( .A1(n24925), .A2(n24936), .ZN(n24921) );
  AOI22_X2 U17620 ( .A1(n13258), .A2(n25712), .B1(n13924), .B2(n12314), .ZN(
        n33537) );
  XOR2_X1 U17623 ( .A1(n30104), .A2(n32997), .Z(n4682) );
  XOR2_X1 U17624 ( .A1(n15508), .A2(n7511), .Z(n32997) );
  OAI21_X1 U17627 ( .A1(n5867), .A2(n10822), .B(n25072), .ZN(n5866) );
  NOR2_X2 U17628 ( .A1(n13551), .A2(n13552), .ZN(n24394) );
  AOI22_X2 U17639 ( .A1(n5678), .A2(n1920), .B1(n2021), .B2(n845), .ZN(n33244)
         );
  NAND2_X2 U17642 ( .A1(n32999), .A2(n32998), .ZN(n23672) );
  INV_X2 U17644 ( .I(n23942), .ZN(n32999) );
  AOI22_X2 U17645 ( .A1(n30725), .A2(n26882), .B1(n23871), .B2(n3571), .ZN(
        n12841) );
  XOR2_X1 U17646 ( .A1(n11349), .A2(n16708), .Z(n5337) );
  OAI21_X2 U17647 ( .A1(n2251), .A2(n2250), .B(n12115), .ZN(n11349) );
  NAND2_X2 U17649 ( .A1(n33001), .A2(n34007), .ZN(n27252) );
  NAND2_X2 U17652 ( .A1(n8821), .A2(n8822), .ZN(n18017) );
  OAI21_X2 U17658 ( .A1(n8307), .A2(n5292), .B(n33002), .ZN(n25784) );
  XOR2_X1 U17659 ( .A1(n33004), .A2(n572), .Z(n10663) );
  XOR2_X1 U17661 ( .A1(n358), .A2(n14908), .Z(n33004) );
  INV_X1 U17662 ( .I(n33006), .ZN(n11077) );
  NAND2_X2 U17665 ( .A1(n32093), .A2(n33006), .ZN(n33005) );
  NAND2_X2 U17666 ( .A1(n33670), .A2(n16333), .ZN(n33006) );
  XOR2_X1 U17668 ( .A1(n20851), .A2(n20928), .Z(n33332) );
  AOI21_X2 U17670 ( .A1(n12782), .A2(n851), .B(n33008), .ZN(n23318) );
  OAI21_X2 U17671 ( .A1(n22908), .A2(n29329), .B(n22981), .ZN(n22910) );
  INV_X2 U17673 ( .I(n33009), .ZN(n17124) );
  AOI21_X2 U17674 ( .A1(n1300), .A2(n22626), .B(n33010), .ZN(n33009) );
  XOR2_X1 U17677 ( .A1(n13651), .A2(n16242), .Z(n22000) );
  NAND2_X2 U17678 ( .A1(n15698), .A2(n21873), .ZN(n16242) );
  AOI21_X1 U17682 ( .A1(n14524), .A2(n14525), .B(n17139), .ZN(n14151) );
  NAND2_X2 U17685 ( .A1(n6178), .A2(n6177), .ZN(n21626) );
  XOR2_X1 U17694 ( .A1(n15517), .A2(n24616), .Z(n24539) );
  NAND2_X2 U17695 ( .A1(n33012), .A2(n24208), .ZN(n24830) );
  OAI21_X2 U17698 ( .A1(n2463), .A2(n24206), .B(n33549), .ZN(n33012) );
  XOR2_X1 U17699 ( .A1(n27567), .A2(n33013), .Z(n9789) );
  XOR2_X1 U17705 ( .A1(n10519), .A2(n623), .Z(n33013) );
  OAI21_X1 U17709 ( .A1(n29335), .A2(n11895), .B(n22553), .ZN(n14776) );
  XOR2_X1 U17712 ( .A1(n33014), .A2(n24754), .Z(n7794) );
  XOR2_X1 U17713 ( .A1(n9281), .A2(n27852), .Z(n33014) );
  XNOR2_X1 U17715 ( .A1(n24516), .A2(n25598), .ZN(n33128) );
  NAND3_X2 U17718 ( .A1(n27495), .A2(n2548), .A3(n33015), .ZN(n2813) );
  XOR2_X1 U17720 ( .A1(n20835), .A2(n16641), .Z(n5630) );
  BUF_X2 U17726 ( .I(n31894), .Z(n33016) );
  XOR2_X1 U17732 ( .A1(n31860), .A2(n20765), .Z(n17804) );
  XOR2_X1 U17733 ( .A1(n28100), .A2(n532), .Z(n33017) );
  NOR2_X2 U17739 ( .A1(n8094), .A2(n33018), .ZN(n33616) );
  OR2_X2 U17743 ( .A1(n10327), .A2(n14238), .Z(n25905) );
  XOR2_X1 U17745 ( .A1(n33351), .A2(n28819), .Z(n10327) );
  XOR2_X1 U17749 ( .A1(n22148), .A2(n22318), .Z(n10598) );
  NAND2_X2 U17752 ( .A1(n21484), .A2(n21485), .ZN(n22148) );
  NAND2_X1 U17754 ( .A1(n28992), .A2(n25650), .ZN(n33020) );
  AOI22_X2 U17757 ( .A1(n29281), .A2(n7609), .B1(n10804), .B2(n10805), .ZN(
        n29615) );
  XOR2_X1 U17764 ( .A1(n24813), .A2(n7837), .Z(n7838) );
  NAND2_X2 U17766 ( .A1(n11388), .A2(n11387), .ZN(n24813) );
  XOR2_X1 U17768 ( .A1(n15384), .A2(n22036), .Z(n17918) );
  AOI21_X2 U17769 ( .A1(n21275), .A2(n21732), .B(n15385), .ZN(n15384) );
  XNOR2_X1 U17775 ( .A1(n25224), .A2(n28898), .ZN(n33579) );
  NOR3_X2 U17779 ( .A1(n30758), .A2(n33021), .A3(n3934), .ZN(n28077) );
  NAND3_X2 U17780 ( .A1(n4823), .A2(n4822), .A3(n4824), .ZN(n24257) );
  AOI22_X2 U17784 ( .A1(n23954), .A2(n4991), .B1(n7140), .B2(n13998), .ZN(
        n4822) );
  INV_X1 U17787 ( .I(n33023), .ZN(n9446) );
  NAND3_X2 U17791 ( .A1(n2348), .A2(n33945), .A3(n22344), .ZN(n23009) );
  NOR2_X2 U17794 ( .A1(n14594), .A2(n14595), .ZN(n21964) );
  NAND2_X1 U17797 ( .A1(n24162), .A2(n24340), .ZN(n23781) );
  AOI22_X1 U17803 ( .A1(n11069), .A2(n25292), .B1(n25196), .B2(n7081), .ZN(
        n33024) );
  NAND2_X2 U17804 ( .A1(n21680), .A2(n21681), .ZN(n17362) );
  NAND3_X1 U17805 ( .A1(n2342), .A2(n14540), .A3(n11626), .ZN(n33686) );
  XOR2_X1 U17808 ( .A1(n13041), .A2(n7653), .Z(n21033) );
  NAND2_X2 U17812 ( .A1(n13851), .A2(n30892), .ZN(n7653) );
  NOR2_X2 U17816 ( .A1(n33075), .A2(n29499), .ZN(n9890) );
  NAND2_X2 U17817 ( .A1(n9452), .A2(n9451), .ZN(n4834) );
  XOR2_X1 U17818 ( .A1(n33025), .A2(n10773), .Z(n23188) );
  XOR2_X1 U17821 ( .A1(n23368), .A2(n23247), .Z(n33025) );
  OAI21_X1 U17824 ( .A1(n14627), .A2(n1218), .B(n17987), .ZN(n33030) );
  XOR2_X1 U17827 ( .A1(n24536), .A2(n33027), .Z(n27490) );
  XOR2_X1 U17828 ( .A1(n8413), .A2(n33028), .Z(n33027) );
  NAND2_X2 U17835 ( .A1(n33029), .A2(n21104), .ZN(n15414) );
  OAI21_X2 U17843 ( .A1(n26735), .A2(n26736), .B(n21251), .ZN(n33029) );
  NOR2_X1 U17845 ( .A1(n22743), .A2(n16922), .ZN(n30315) );
  XOR2_X1 U17851 ( .A1(n29858), .A2(n17203), .Z(n17204) );
  AOI21_X2 U17856 ( .A1(n30050), .A2(n28502), .B(n31999), .ZN(n17079) );
  NAND2_X2 U17857 ( .A1(n15584), .A2(n33043), .ZN(n11041) );
  NOR2_X2 U17860 ( .A1(n23037), .A2(n28415), .ZN(n12444) );
  NAND2_X2 U17867 ( .A1(n13412), .A2(n9964), .ZN(n24044) );
  NAND2_X2 U17869 ( .A1(n9589), .A2(n21480), .ZN(n16269) );
  BUF_X2 U17873 ( .I(n16051), .Z(n33032) );
  NOR2_X2 U17874 ( .A1(n29246), .A2(n10955), .ZN(n28855) );
  INV_X2 U17881 ( .I(n18235), .ZN(n21692) );
  NAND2_X2 U17882 ( .A1(n5628), .A2(n3286), .ZN(n18235) );
  OAI21_X2 U17886 ( .A1(n33034), .A2(n33033), .B(n15149), .ZN(n29975) );
  NOR2_X2 U17900 ( .A1(n7238), .A2(n349), .ZN(n33033) );
  INV_X2 U17904 ( .I(n21219), .ZN(n33034) );
  NOR2_X2 U17905 ( .A1(n29305), .A2(n654), .ZN(n23705) );
  INV_X2 U17912 ( .I(n376), .ZN(n654) );
  XOR2_X1 U17913 ( .A1(n12579), .A2(n28031), .Z(n376) );
  AOI21_X2 U17916 ( .A1(n6704), .A2(n29905), .B(n31048), .ZN(n33035) );
  XOR2_X1 U17917 ( .A1(n27875), .A2(n33036), .Z(n11223) );
  XOR2_X1 U17919 ( .A1(n33823), .A2(n23391), .Z(n33036) );
  XOR2_X1 U17928 ( .A1(n10460), .A2(n20692), .Z(n20863) );
  NOR2_X2 U17930 ( .A1(n30612), .A2(n33037), .ZN(n16364) );
  NOR2_X1 U17932 ( .A1(n20206), .A2(n20464), .ZN(n20207) );
  INV_X2 U17933 ( .I(n33038), .ZN(n15438) );
  XOR2_X1 U17937 ( .A1(n3253), .A2(n12945), .Z(n33038) );
  NAND2_X1 U17941 ( .A1(n31522), .A2(n20257), .ZN(n33820) );
  BUF_X2 U17944 ( .I(n881), .Z(n33039) );
  XOR2_X1 U17951 ( .A1(n1307), .A2(n3704), .Z(n12627) );
  NOR2_X2 U17960 ( .A1(n9088), .A2(n33483), .ZN(n16237) );
  NAND2_X2 U17961 ( .A1(n6926), .A2(n29008), .ZN(n28028) );
  NAND2_X1 U17967 ( .A1(n19986), .A2(n16), .ZN(n19459) );
  XOR2_X1 U17968 ( .A1(n11580), .A2(n14621), .Z(n16) );
  XOR2_X1 U17969 ( .A1(n22143), .A2(n22144), .Z(n4627) );
  XNOR2_X1 U17978 ( .A1(n4529), .A2(n4530), .ZN(n33376) );
  OAI21_X2 U17979 ( .A1(n16372), .A2(n18554), .B(n9555), .ZN(n19249) );
  XOR2_X1 U17981 ( .A1(n22267), .A2(n22191), .Z(n30250) );
  NAND3_X2 U17982 ( .A1(n33228), .A2(n33229), .A3(n18956), .ZN(n19558) );
  AOI21_X1 U17983 ( .A1(n21228), .A2(n21305), .B(n21132), .ZN(n31728) );
  NAND2_X1 U17986 ( .A1(n4834), .A2(n23086), .ZN(n17669) );
  XOR2_X1 U17987 ( .A1(n29501), .A2(n22102), .Z(n22180) );
  NAND2_X2 U17989 ( .A1(n5289), .A2(n18218), .ZN(n13028) );
  NAND2_X2 U17996 ( .A1(n31989), .A2(n5836), .ZN(n5289) );
  XOR2_X1 U17998 ( .A1(n26889), .A2(n33042), .Z(n29075) );
  XOR2_X1 U18002 ( .A1(n11996), .A2(n23236), .Z(n33042) );
  NAND2_X2 U18006 ( .A1(n10149), .A2(n21379), .ZN(n10148) );
  OAI22_X2 U18007 ( .A1(n20458), .A2(n20459), .B1(n20457), .B2(n3487), .ZN(
        n21040) );
  NAND2_X2 U18009 ( .A1(n9976), .A2(n9977), .ZN(n24161) );
  NAND3_X2 U18011 ( .A1(n33045), .A2(n24295), .A3(n15520), .ZN(n6165) );
  NAND2_X2 U18015 ( .A1(n7779), .A2(n5631), .ZN(n33045) );
  NAND2_X2 U18016 ( .A1(n30185), .A2(n11418), .ZN(n2826) );
  OAI21_X2 U18019 ( .A1(n24009), .A2(n17602), .B(n33047), .ZN(n9708) );
  AOI22_X2 U18020 ( .A1(n22906), .A2(n33522), .B1(n989), .B2(n22907), .ZN(
        n5343) );
  NOR2_X2 U18025 ( .A1(n23069), .A2(n22865), .ZN(n22906) );
  XOR2_X1 U18033 ( .A1(n33048), .A2(n12717), .Z(n27042) );
  XOR2_X1 U18037 ( .A1(n23272), .A2(n15114), .Z(n33048) );
  NAND3_X2 U18039 ( .A1(n33049), .A2(n22701), .A3(n12646), .ZN(n23417) );
  INV_X1 U18041 ( .I(n22960), .ZN(n33050) );
  OR2_X1 U18043 ( .A1(n29952), .A2(n33050), .Z(n22701) );
  XOR2_X1 U18045 ( .A1(n22084), .A2(n27943), .Z(n27942) );
  AOI21_X1 U18051 ( .A1(n22332), .A2(n8420), .B(n28692), .ZN(n29823) );
  XOR2_X1 U18054 ( .A1(n33051), .A2(n23194), .Z(n27441) );
  XOR2_X1 U18058 ( .A1(n31567), .A2(n29012), .Z(n33051) );
  NAND2_X2 U18059 ( .A1(n10806), .A2(n33136), .ZN(n28840) );
  NOR2_X2 U18065 ( .A1(n16847), .A2(n19053), .ZN(n2584) );
  XOR2_X1 U18067 ( .A1(n27413), .A2(n27412), .Z(n28702) );
  BUF_X2 U18074 ( .I(n24610), .Z(n33053) );
  AND3_X1 U18077 ( .A1(n24243), .A2(n28374), .A3(n24242), .Z(n30000) );
  XOR2_X1 U18078 ( .A1(n33054), .A2(n25373), .Z(Ciphertext[100]) );
  NAND3_X2 U18081 ( .A1(n25372), .A2(n25371), .A3(n25370), .ZN(n33054) );
  OAI22_X2 U18083 ( .A1(n33055), .A2(n1528), .B1(n11708), .B2(n29294), .ZN(
        n31707) );
  INV_X4 U18086 ( .I(n6357), .ZN(n21832) );
  XOR2_X1 U18091 ( .A1(n23439), .A2(n10535), .Z(n23277) );
  NAND2_X2 U18093 ( .A1(n33728), .A2(n13559), .ZN(n15212) );
  OAI21_X2 U18094 ( .A1(n32493), .A2(n28669), .B(n629), .ZN(n33056) );
  XOR2_X1 U18095 ( .A1(n20664), .A2(n5647), .Z(n6701) );
  XOR2_X1 U18097 ( .A1(n20849), .A2(n20658), .Z(n20664) );
  XOR2_X1 U18098 ( .A1(n23790), .A2(n33057), .Z(n30398) );
  XOR2_X1 U18099 ( .A1(n9907), .A2(n33058), .Z(n33057) );
  XOR2_X1 U18100 ( .A1(n33059), .A2(n25355), .Z(Ciphertext[97]) );
  OAI22_X1 U18101 ( .A1(n25353), .A2(n25354), .B1(n25380), .B2(n25360), .ZN(
        n33059) );
  OAI22_X1 U18103 ( .A1(n24904), .A2(n24905), .B1(n24903), .B2(n10099), .ZN(
        n33717) );
  NAND2_X2 U18105 ( .A1(n33060), .A2(n23644), .ZN(n24226) );
  NAND2_X1 U18107 ( .A1(n3757), .A2(n34075), .ZN(n33060) );
  INV_X2 U18109 ( .I(n24219), .ZN(n1096) );
  OAI21_X2 U18110 ( .A1(n14037), .A2(n23604), .B(n32008), .ZN(n24219) );
  NOR2_X2 U18111 ( .A1(n23033), .A2(n6605), .ZN(n23035) );
  INV_X2 U18118 ( .I(n11933), .ZN(n33583) );
  XOR2_X1 U18124 ( .A1(n1988), .A2(n33062), .Z(n21455) );
  XOR2_X1 U18132 ( .A1(n21034), .A2(n1986), .Z(n33062) );
  XOR2_X1 U18137 ( .A1(n33063), .A2(n25428), .Z(Ciphertext[104]) );
  NAND2_X1 U18139 ( .A1(n33546), .A2(n25427), .ZN(n33063) );
  NAND2_X1 U18143 ( .A1(n25425), .A2(n25455), .ZN(n15500) );
  NAND2_X2 U18146 ( .A1(n15783), .A2(n33064), .ZN(n17948) );
  XOR2_X1 U18148 ( .A1(n12714), .A2(n23408), .Z(n3280) );
  NAND2_X2 U18151 ( .A1(n3282), .A2(n3281), .ZN(n12714) );
  OAI21_X2 U18152 ( .A1(n8279), .A2(n24118), .B(n33065), .ZN(n8502) );
  NAND2_X2 U18154 ( .A1(n24224), .A2(n24222), .ZN(n33065) );
  XOR2_X1 U18156 ( .A1(n8050), .A2(n24816), .Z(n24593) );
  NAND2_X2 U18162 ( .A1(n23610), .A2(n23609), .ZN(n8050) );
  NAND2_X1 U18164 ( .A1(n25383), .A2(n25561), .ZN(n33068) );
  NOR3_X2 U18167 ( .A1(n7776), .A2(n7775), .A3(n7232), .ZN(n1877) );
  AOI22_X2 U18174 ( .A1(n25925), .A2(n7701), .B1(n5411), .B2(n25923), .ZN(
        n25927) );
  NAND2_X2 U18177 ( .A1(n33071), .A2(n33070), .ZN(n2558) );
  OAI21_X2 U18189 ( .A1(n2563), .A2(n13402), .B(n26965), .ZN(n33070) );
  AND2_X1 U18193 ( .A1(n16625), .A2(n33430), .Z(n19801) );
  OAI21_X2 U18194 ( .A1(n15905), .A2(n1337), .B(n33209), .ZN(n12221) );
  XOR2_X1 U18195 ( .A1(n11324), .A2(n23165), .Z(n33073) );
  AND2_X1 U18202 ( .A1(n17770), .A2(n17787), .Z(n33074) );
  XOR2_X1 U18203 ( .A1(n19728), .A2(n32184), .Z(n17954) );
  XOR2_X1 U18209 ( .A1(n30943), .A2(n26751), .Z(n19728) );
  XOR2_X1 U18212 ( .A1(n20912), .A2(n20833), .Z(n30107) );
  XOR2_X1 U18213 ( .A1(n21040), .A2(n21018), .Z(n20912) );
  OAI22_X2 U18216 ( .A1(n17374), .A2(n2752), .B1(n1100), .B2(n23555), .ZN(
        n33075) );
  XOR2_X1 U18217 ( .A1(n23274), .A2(n1260), .Z(n23459) );
  NOR2_X2 U18220 ( .A1(n7921), .A2(n33076), .ZN(n7762) );
  OAI22_X2 U18228 ( .A1(n19862), .A2(n7920), .B1(n7922), .B2(n16694), .ZN(
        n33076) );
  NAND2_X2 U18233 ( .A1(n6123), .A2(n31148), .ZN(n14953) );
  NOR2_X2 U18234 ( .A1(n21719), .A2(n6718), .ZN(n17716) );
  NAND2_X2 U18236 ( .A1(n19249), .A2(n4436), .ZN(n19248) );
  XOR2_X1 U18239 ( .A1(n8921), .A2(n19585), .Z(n4169) );
  XOR2_X1 U18240 ( .A1(n1372), .A2(n19679), .Z(n19585) );
  XOR2_X1 U18243 ( .A1(n33077), .A2(n1402), .Z(Ciphertext[153]) );
  NOR2_X1 U18244 ( .A1(n31833), .A2(n5784), .ZN(n33077) );
  NOR2_X2 U18250 ( .A1(n18006), .A2(n13846), .ZN(n18470) );
  XOR2_X1 U18253 ( .A1(n12674), .A2(n32889), .Z(n10628) );
  NOR2_X2 U18254 ( .A1(n31290), .A2(n31291), .ZN(n20792) );
  NAND2_X2 U18263 ( .A1(n9966), .A2(n9965), .ZN(n27114) );
  XOR2_X1 U18266 ( .A1(Plaintext[110]), .A2(Key[110]), .Z(n33094) );
  NAND2_X1 U18268 ( .A1(n33069), .A2(n19120), .ZN(n18956) );
  INV_X2 U18273 ( .I(n19118), .ZN(n33078) );
  XOR2_X1 U18274 ( .A1(n33079), .A2(n19686), .Z(n17835) );
  XOR2_X1 U18276 ( .A1(n31731), .A2(n25578), .Z(n33079) );
  NAND2_X2 U18279 ( .A1(n33080), .A2(n33732), .ZN(n30130) );
  OAI22_X2 U18280 ( .A1(n20035), .A2(n20034), .B1(n16243), .B2(n2795), .ZN(
        n33080) );
  XOR2_X1 U18287 ( .A1(n33081), .A2(n16672), .Z(Ciphertext[15]) );
  INV_X2 U18288 ( .I(n33082), .ZN(n10438) );
  NAND2_X1 U18290 ( .A1(n17977), .A2(n17978), .ZN(n33431) );
  XOR2_X1 U18293 ( .A1(n705), .A2(n24813), .Z(n24797) );
  NOR2_X2 U18296 ( .A1(n13217), .A2(n8204), .ZN(n705) );
  AND2_X1 U18299 ( .A1(n12221), .A2(n33083), .Z(n17226) );
  XOR2_X1 U18300 ( .A1(n22183), .A2(n27190), .Z(n5976) );
  XOR2_X1 U18301 ( .A1(n33084), .A2(n28462), .Z(Ciphertext[52]) );
  INV_X2 U18302 ( .I(n34128), .ZN(n13073) );
  XOR2_X1 U18304 ( .A1(n33358), .A2(n33085), .Z(n34128) );
  XOR2_X1 U18305 ( .A1(n26530), .A2(n20860), .Z(n20668) );
  NOR2_X2 U18312 ( .A1(n8959), .A2(n8960), .ZN(n26530) );
  OAI21_X2 U18313 ( .A1(n22671), .A2(n27357), .B(n2311), .ZN(n30297) );
  NOR2_X2 U18315 ( .A1(n26663), .A2(n26784), .ZN(n4254) );
  NAND2_X2 U18316 ( .A1(n12496), .A2(n22503), .ZN(n22530) );
  NOR3_X1 U18319 ( .A1(n8902), .A2(n16798), .A3(n1204), .ZN(n16793) );
  OR2_X1 U18322 ( .A1(n3339), .A2(n25111), .Z(n33314) );
  XOR2_X1 U18323 ( .A1(n19409), .A2(n19398), .Z(n6731) );
  NAND2_X2 U18325 ( .A1(n10741), .A2(n10739), .ZN(n19409) );
  XOR2_X1 U18327 ( .A1(n15556), .A2(n29443), .Z(n30094) );
  XOR2_X1 U18342 ( .A1(n33086), .A2(n19496), .Z(n3283) );
  XOR2_X1 U18345 ( .A1(n29890), .A2(n1045), .Z(n33086) );
  XOR2_X1 U18349 ( .A1(n23459), .A2(n8974), .Z(n8973) );
  NAND2_X2 U18356 ( .A1(n25330), .A2(n6411), .ZN(n25375) );
  NAND2_X2 U18357 ( .A1(n33087), .A2(n25017), .ZN(n25058) );
  OAI21_X2 U18361 ( .A1(n11977), .A2(n14959), .B(n14846), .ZN(n33087) );
  NAND2_X2 U18364 ( .A1(n9826), .A2(n9825), .ZN(n24545) );
  XOR2_X1 U18365 ( .A1(n17095), .A2(n17096), .Z(n17094) );
  NAND3_X1 U18366 ( .A1(n14232), .A2(n27577), .A3(n13720), .ZN(n12883) );
  AOI21_X1 U18373 ( .A1(n33310), .A2(n18085), .B(n1182), .ZN(n15928) );
  OR2_X1 U18374 ( .A1(n1279), .A2(n4135), .Z(n7946) );
  NAND3_X2 U18375 ( .A1(n33089), .A2(n33750), .A3(n16225), .ZN(n21974) );
  NAND2_X2 U18376 ( .A1(n31551), .A2(n630), .ZN(n33089) );
  NAND2_X2 U18377 ( .A1(n263), .A2(n262), .ZN(n7293) );
  NOR2_X2 U18392 ( .A1(n1557), .A2(n26328), .ZN(n34099) );
  OAI21_X2 U18393 ( .A1(n33441), .A2(n13978), .B(n17136), .ZN(n33527) );
  XOR2_X1 U18395 ( .A1(n23375), .A2(n22970), .Z(n23517) );
  NOR2_X2 U18401 ( .A1(n27566), .A2(n7945), .ZN(n23375) );
  NAND2_X2 U18402 ( .A1(n21163), .A2(n11734), .ZN(n13593) );
  XOR2_X1 U18403 ( .A1(n33090), .A2(n24445), .Z(n27526) );
  XOR2_X1 U18412 ( .A1(n24691), .A2(n8050), .Z(n24525) );
  NAND3_X2 U18415 ( .A1(n11964), .A2(n13630), .A3(n13628), .ZN(n25988) );
  INV_X2 U18417 ( .I(n33092), .ZN(n9064) );
  XNOR2_X1 U18419 ( .A1(n33636), .A2(n7640), .ZN(n33092) );
  NOR2_X2 U18422 ( .A1(n29769), .A2(n19118), .ZN(n19119) );
  NAND2_X2 U18423 ( .A1(n926), .A2(n6520), .ZN(n10730) );
  XOR2_X1 U18428 ( .A1(n12454), .A2(n24836), .Z(n30493) );
  INV_X2 U18432 ( .I(n12748), .ZN(n26778) );
  NAND2_X2 U18439 ( .A1(n14501), .A2(n24059), .ZN(n13470) );
  NAND3_X2 U18444 ( .A1(n6354), .A2(n7069), .A3(n13306), .ZN(n14501) );
  XOR2_X1 U18446 ( .A1(n4312), .A2(n287), .Z(n9375) );
  OR2_X1 U18448 ( .A1(n12551), .A2(n3222), .Z(n24071) );
  XOR2_X1 U18459 ( .A1(n30131), .A2(n4682), .Z(n25696) );
  AOI22_X2 U18466 ( .A1(n28585), .A2(n33011), .B1(n23747), .B2(n16628), .ZN(
        n23748) );
  INV_X1 U18468 ( .I(n686), .ZN(n33095) );
  OR2_X1 U18469 ( .A1(n22999), .A2(n16297), .Z(n7219) );
  NOR2_X2 U18472 ( .A1(n17922), .A2(n33096), .ZN(n26883) );
  OR2_X1 U18474 ( .A1(n33766), .A2(n31958), .Z(n14209) );
  BUF_X2 U18479 ( .I(n16569), .Z(n33098) );
  XOR2_X1 U18480 ( .A1(n15297), .A2(n28710), .Z(n34118) );
  NOR2_X2 U18481 ( .A1(n20589), .A2(n31967), .ZN(n15638) );
  XOR2_X1 U18482 ( .A1(n33099), .A2(n6620), .Z(n33617) );
  XOR2_X1 U18483 ( .A1(n33100), .A2(n30917), .Z(n33099) );
  XOR2_X1 U18486 ( .A1(n3964), .A2(n19341), .Z(n31414) );
  NOR2_X2 U18489 ( .A1(n19162), .A2(n19161), .ZN(n19341) );
  NAND3_X2 U18490 ( .A1(n17692), .A2(n21747), .A3(n21746), .ZN(n4034) );
  AOI21_X2 U18493 ( .A1(n29632), .A2(n8176), .B(n21968), .ZN(n33115) );
  XOR2_X1 U18507 ( .A1(n20720), .A2(n31966), .Z(n20757) );
  NOR2_X2 U18511 ( .A1(n13597), .A2(n22964), .ZN(n12662) );
  XOR2_X1 U18512 ( .A1(n20558), .A2(n20718), .Z(n10391) );
  OAI22_X2 U18513 ( .A1(n7426), .A2(n33105), .B1(n7427), .B2(n15740), .ZN(
        n16315) );
  BUF_X2 U18514 ( .I(n4568), .Z(n33106) );
  INV_X4 U18516 ( .I(n8130), .ZN(n1350) );
  NAND2_X1 U18518 ( .A1(n14545), .A2(n8130), .ZN(n33107) );
  NOR2_X1 U18520 ( .A1(n15340), .A2(n5578), .ZN(n5173) );
  OAI21_X1 U18527 ( .A1(n33432), .A2(n19275), .B(n33108), .ZN(n18971) );
  XOR2_X1 U18536 ( .A1(n33109), .A2(n10332), .Z(n29828) );
  XOR2_X1 U18540 ( .A1(n20802), .A2(n25311), .Z(n33109) );
  XOR2_X1 U18541 ( .A1(n4321), .A2(n2388), .Z(n29028) );
  NOR3_X2 U18549 ( .A1(n6024), .A2(n11581), .A3(n6023), .ZN(n4321) );
  NAND2_X1 U18557 ( .A1(n21530), .A2(n29980), .ZN(n6231) );
  NOR2_X2 U18562 ( .A1(n28299), .A2(n28298), .ZN(n21530) );
  XOR2_X1 U18567 ( .A1(n2349), .A2(n1129), .Z(n22187) );
  OAI21_X2 U18578 ( .A1(n33113), .A2(n33112), .B(n2574), .ZN(n8391) );
  NOR2_X1 U18584 ( .A1(n1632), .A2(n17439), .ZN(n33112) );
  INV_X2 U18587 ( .I(n33114), .ZN(n23706) );
  XNOR2_X1 U18591 ( .A1(n17826), .A2(n33490), .ZN(n33114) );
  AND2_X1 U18594 ( .A1(n29980), .A2(n21530), .Z(n16952) );
  NAND2_X2 U18603 ( .A1(n14717), .A2(n12221), .ZN(n27595) );
  XOR2_X1 U18606 ( .A1(n24852), .A2(n8480), .Z(n24427) );
  NAND3_X2 U18608 ( .A1(n11962), .A2(n3021), .A3(n24071), .ZN(n24852) );
  NOR2_X1 U18610 ( .A1(n31664), .A2(n24069), .ZN(n31663) );
  XOR2_X1 U18612 ( .A1(n15588), .A2(n24600), .Z(n1441) );
  NAND2_X1 U18614 ( .A1(n28414), .A2(n27697), .ZN(n26800) );
  NAND2_X2 U18615 ( .A1(n2934), .A2(n19807), .ZN(n27697) );
  XOR2_X1 U18617 ( .A1(n23402), .A2(n27552), .Z(n33606) );
  NOR2_X2 U18621 ( .A1(n23052), .A2(n22798), .ZN(n6099) );
  XOR2_X1 U18623 ( .A1(n23415), .A2(n23414), .Z(n33118) );
  XOR2_X1 U18625 ( .A1(n24569), .A2(n15438), .Z(n10196) );
  OAI21_X2 U18627 ( .A1(n13642), .A2(n13641), .B(n33119), .ZN(n13637) );
  NOR2_X2 U18628 ( .A1(n33786), .A2(n4350), .ZN(n4349) );
  XOR2_X1 U18630 ( .A1(n5904), .A2(n23292), .Z(n33465) );
  OR2_X1 U18637 ( .A1(n17503), .A2(n31943), .Z(n13231) );
  XOR2_X1 U18639 ( .A1(n12252), .A2(n23196), .Z(n23451) );
  NAND2_X2 U18650 ( .A1(n22767), .A2(n22768), .ZN(n12252) );
  XOR2_X1 U18653 ( .A1(n33121), .A2(n11822), .Z(n27570) );
  XOR2_X1 U18660 ( .A1(n31611), .A2(n23296), .Z(n33121) );
  OAI21_X2 U18661 ( .A1(n8315), .A2(n14091), .B(n6119), .ZN(n33122) );
  NAND2_X2 U18663 ( .A1(n33708), .A2(n8463), .ZN(n22232) );
  XOR2_X1 U18664 ( .A1(n19625), .A2(n16429), .Z(n17540) );
  NOR2_X2 U18665 ( .A1(n27718), .A2(n19077), .ZN(n19625) );
  NAND2_X2 U18666 ( .A1(n21083), .A2(n7620), .ZN(n12827) );
  XOR2_X1 U18669 ( .A1(n5185), .A2(n31887), .Z(n33153) );
  NAND2_X2 U18670 ( .A1(n16297), .A2(n22999), .ZN(n5682) );
  XOR2_X1 U18672 ( .A1(n10005), .A2(n13873), .Z(n10004) );
  NAND2_X2 U18680 ( .A1(n33125), .A2(n33859), .ZN(n11755) );
  AOI21_X2 U18687 ( .A1(n21312), .A2(n13194), .B(n34159), .ZN(n33125) );
  NAND2_X1 U18688 ( .A1(n9917), .A2(n17044), .ZN(n9916) );
  NAND2_X2 U18690 ( .A1(n21390), .A2(n6179), .ZN(n6177) );
  NAND2_X1 U18691 ( .A1(n16716), .A2(n22889), .ZN(n33126) );
  XOR2_X1 U18693 ( .A1(n28448), .A2(n33127), .Z(n30526) );
  XOR2_X1 U18696 ( .A1(n24418), .A2(n33128), .Z(n33127) );
  AOI21_X2 U18701 ( .A1(n9689), .A2(n33515), .B(n33129), .ZN(n12902) );
  NOR3_X2 U18705 ( .A1(n33515), .A2(n13300), .A3(n1154), .ZN(n33129) );
  XOR2_X1 U18712 ( .A1(n15823), .A2(n33130), .Z(n10800) );
  XOR2_X1 U18714 ( .A1(n31584), .A2(n31884), .Z(n33130) );
  OAI21_X1 U18717 ( .A1(n33144), .A2(n14335), .B(n33722), .ZN(n3289) );
  INV_X2 U18720 ( .I(n8166), .ZN(n14335) );
  XOR2_X1 U18721 ( .A1(n33866), .A2(n1436), .Z(n8166) );
  NAND2_X2 U18722 ( .A1(n33131), .A2(n15624), .ZN(n31793) );
  NAND2_X2 U18723 ( .A1(n30561), .A2(n31149), .ZN(n33131) );
  NAND2_X2 U18724 ( .A1(n28253), .A2(n30826), .ZN(n13545) );
  AOI22_X2 U18726 ( .A1(n33180), .A2(n22483), .B1(n9022), .B2(n22297), .ZN(
        n4221) );
  OAI21_X1 U18728 ( .A1(n21705), .A2(n26782), .B(n2643), .ZN(n26479) );
  INV_X2 U18731 ( .I(n33134), .ZN(n10325) );
  XNOR2_X1 U18732 ( .A1(Plaintext[4]), .A2(Key[4]), .ZN(n33134) );
  NAND3_X1 U18734 ( .A1(n31977), .A2(n33277), .A3(n24611), .ZN(n24613) );
  OAI22_X2 U18739 ( .A1(n23811), .A2(n23559), .B1(n23558), .B2(n23947), .ZN(
        n23560) );
  NAND2_X2 U18743 ( .A1(n33135), .A2(n18117), .ZN(n5306) );
  NOR2_X2 U18745 ( .A1(n23007), .A2(n23013), .ZN(n10528) );
  OAI22_X2 U18754 ( .A1(n22348), .A2(n996), .B1(n7965), .B2(n22450), .ZN(
        n23013) );
  OAI21_X1 U18758 ( .A1(n8757), .A2(n21054), .B(n33137), .ZN(n33142) );
  NAND2_X1 U18759 ( .A1(n15323), .A2(n6402), .ZN(n33138) );
  XOR2_X1 U18761 ( .A1(n20690), .A2(n21047), .Z(n5775) );
  INV_X2 U18763 ( .I(n30191), .ZN(n24268) );
  NAND3_X2 U18768 ( .A1(n31691), .A2(n31690), .A3(n11670), .ZN(n30191) );
  NAND3_X2 U18769 ( .A1(n2167), .A2(n10152), .A3(n31173), .ZN(n26363) );
  NAND2_X2 U18771 ( .A1(n33797), .A2(n33694), .ZN(n10312) );
  XOR2_X1 U18775 ( .A1(n2820), .A2(n2819), .Z(n31101) );
  NOR2_X1 U18776 ( .A1(n23694), .A2(n28367), .ZN(n33226) );
  OAI21_X2 U18779 ( .A1(n9233), .A2(n18172), .B(n33140), .ZN(n29763) );
  AOI22_X2 U18781 ( .A1(n33141), .A2(n17238), .B1(n12249), .B2(n12497), .ZN(
        n19463) );
  OAI21_X2 U18782 ( .A1(n12249), .A2(n12500), .B(n18135), .ZN(n33141) );
  NAND2_X2 U18788 ( .A1(n33142), .A2(n31848), .ZN(n21719) );
  AOI22_X2 U18789 ( .A1(n21771), .A2(n26904), .B1(n2718), .B2(n38), .ZN(n4219)
         );
  BUF_X4 U18790 ( .I(n23499), .Z(n33293) );
  BUF_X2 U18802 ( .I(n18919), .Z(n33143) );
  BUF_X2 U18805 ( .I(n23813), .Z(n33144) );
  NAND2_X1 U18809 ( .A1(n11983), .A2(n31854), .ZN(n13575) );
  NAND2_X2 U18815 ( .A1(n22011), .A2(n26394), .ZN(n31854) );
  INV_X2 U18817 ( .I(n7515), .ZN(n715) );
  NAND2_X2 U18818 ( .A1(n26380), .A2(n1859), .ZN(n7515) );
  XOR2_X1 U18820 ( .A1(n4732), .A2(n32860), .Z(n23312) );
  OAI22_X2 U18822 ( .A1(n29789), .A2(n29922), .B1(n33690), .B2(n28263), .ZN(
        n14540) );
  XOR2_X1 U18829 ( .A1(n28323), .A2(n30041), .Z(n29643) );
  OAI21_X1 U18839 ( .A1(n31661), .A2(n31662), .B(n28070), .ZN(n33145) );
  NOR2_X1 U18848 ( .A1(n31932), .A2(n10197), .ZN(n12213) );
  NAND3_X1 U18852 ( .A1(n8206), .A2(n32240), .A3(n20534), .ZN(n20354) );
  XOR2_X1 U18856 ( .A1(n5472), .A2(n20813), .Z(n33508) );
  NAND2_X2 U18861 ( .A1(n2316), .A2(n2318), .ZN(n5472) );
  XNOR2_X1 U18865 ( .A1(n5742), .A2(n25054), .ZN(n33960) );
  NOR2_X2 U18871 ( .A1(n9201), .A2(n20067), .ZN(n11052) );
  NOR2_X1 U18874 ( .A1(n31263), .A2(n25452), .ZN(n25420) );
  XOR2_X1 U18875 ( .A1(n6863), .A2(n6862), .Z(n2557) );
  NOR2_X1 U18876 ( .A1(n28343), .A2(n31357), .ZN(n23773) );
  NAND2_X2 U18879 ( .A1(n30990), .A2(n26579), .ZN(n5454) );
  NOR2_X1 U18880 ( .A1(n8912), .A2(n16745), .ZN(n22335) );
  XOR2_X1 U18881 ( .A1(n13347), .A2(n23274), .Z(n17565) );
  NAND2_X2 U18883 ( .A1(n28355), .A2(n29114), .ZN(n23274) );
  NAND4_X2 U18884 ( .A1(n7091), .A2(n7094), .A3(n23988), .A4(n7095), .ZN(
        n10331) );
  OAI21_X1 U18886 ( .A1(n2066), .A2(n31964), .B(n1288), .ZN(n7819) );
  BUF_X2 U18888 ( .I(n30997), .Z(n33150) );
  XOR2_X1 U18889 ( .A1(n22173), .A2(n33151), .Z(n28000) );
  XOR2_X1 U18891 ( .A1(n33152), .A2(n23447), .Z(n17352) );
  OR2_X1 U18894 ( .A1(n18919), .A2(n18626), .Z(n33965) );
  BUF_X2 U18896 ( .I(n27741), .Z(n33154) );
  NAND2_X2 U18899 ( .A1(n33156), .A2(n28340), .ZN(n21569) );
  NOR2_X2 U18903 ( .A1(n4284), .A2(n4283), .ZN(n33156) );
  NAND2_X2 U18908 ( .A1(n14485), .A2(n14486), .ZN(n20992) );
  XOR2_X1 U18909 ( .A1(n12609), .A2(n33157), .Z(n7566) );
  XOR2_X1 U18914 ( .A1(n8284), .A2(n32889), .Z(n33157) );
  NOR2_X1 U18924 ( .A1(n25060), .A2(n25062), .ZN(n3122) );
  OAI21_X2 U18925 ( .A1(n20055), .A2(n8616), .B(n33158), .ZN(n17715) );
  NAND2_X2 U18927 ( .A1(n3005), .A2(n8616), .ZN(n33158) );
  XOR2_X1 U18930 ( .A1(n33756), .A2(n9464), .Z(n4727) );
  XOR2_X1 U18932 ( .A1(n29481), .A2(n31043), .Z(n9464) );
  OAI21_X1 U18937 ( .A1(n31142), .A2(n25444), .B(n31141), .ZN(n33159) );
  AND2_X1 U18942 ( .A1(n15623), .A2(n34167), .Z(n16540) );
  NAND3_X2 U18943 ( .A1(n7282), .A2(n7176), .A3(n19245), .ZN(n7109) );
  NAND2_X2 U18945 ( .A1(n3183), .A2(n22848), .ZN(n22937) );
  NAND2_X2 U18949 ( .A1(n3187), .A2(n2252), .ZN(n3183) );
  XOR2_X1 U18959 ( .A1(n15823), .A2(n29482), .Z(n27413) );
  XOR2_X1 U18964 ( .A1(n30749), .A2(n20670), .Z(n15823) );
  OAI22_X2 U18966 ( .A1(n4505), .A2(n4506), .B1(n18865), .B2(n18864), .ZN(
        n30865) );
  XOR2_X1 U18969 ( .A1(n14819), .A2(n23253), .Z(n23184) );
  NAND3_X2 U18971 ( .A1(n22943), .A2(n60), .A3(n22942), .ZN(n14819) );
  XOR2_X1 U18978 ( .A1(n14584), .A2(n23119), .Z(n6848) );
  XOR2_X1 U18991 ( .A1(n24651), .A2(n24653), .Z(n33161) );
  NOR3_X1 U18996 ( .A1(n25996), .A2(n652), .A3(n14193), .ZN(n27233) );
  NOR2_X2 U19005 ( .A1(n33162), .A2(n3947), .ZN(n1995) );
  NAND2_X1 U19007 ( .A1(n11563), .A2(n24244), .ZN(n33162) );
  XOR2_X1 U19013 ( .A1(n18125), .A2(n19783), .Z(n30757) );
  INV_X2 U19016 ( .I(n19708), .ZN(n18125) );
  NOR2_X2 U19024 ( .A1(n16907), .A2(n16909), .ZN(n19708) );
  INV_X1 U19027 ( .I(n33163), .ZN(n12201) );
  NOR2_X1 U19030 ( .A1(n24970), .A2(n3843), .ZN(n33163) );
  NAND2_X2 U19031 ( .A1(n33666), .A2(n30928), .ZN(n3843) );
  NOR2_X1 U19032 ( .A1(n4750), .A2(n8365), .ZN(n22879) );
  XOR2_X1 U19039 ( .A1(n23331), .A2(n23256), .Z(n30156) );
  XOR2_X1 U19040 ( .A1(n23438), .A2(n23534), .Z(n23256) );
  NAND2_X2 U19048 ( .A1(n28489), .A2(n33164), .ZN(n31129) );
  NAND2_X2 U19053 ( .A1(n5770), .A2(n5771), .ZN(n33164) );
  OAI21_X2 U19055 ( .A1(n19036), .A2(n26603), .B(n33168), .ZN(n5418) );
  NOR2_X2 U19056 ( .A1(n29962), .A2(n29963), .ZN(n33168) );
  OAI21_X2 U19057 ( .A1(n28136), .A2(n16451), .B(n33169), .ZN(n11705) );
  NAND2_X1 U19058 ( .A1(n28530), .A2(n26570), .ZN(n29934) );
  XOR2_X1 U19063 ( .A1(n33170), .A2(n5722), .Z(n6894) );
  XOR2_X1 U19067 ( .A1(n5724), .A2(n21045), .Z(n33170) );
  NAND2_X1 U19070 ( .A1(n24286), .A2(n17361), .ZN(n29576) );
  XOR2_X1 U19074 ( .A1(n16200), .A2(n23312), .Z(n11143) );
  AOI21_X2 U19087 ( .A1(n31978), .A2(n29552), .B(n33172), .ZN(n2215) );
  NOR3_X2 U19090 ( .A1(n2217), .A2(n21628), .A3(n33992), .ZN(n33172) );
  NAND2_X2 U19093 ( .A1(n16413), .A2(n6939), .ZN(n14547) );
  NAND2_X2 U19095 ( .A1(n33173), .A2(n28506), .ZN(n24084) );
  AOI21_X2 U19098 ( .A1(n14155), .A2(n28676), .B(n33174), .ZN(n33173) );
  INV_X1 U19119 ( .I(n23724), .ZN(n33174) );
  NAND2_X1 U19122 ( .A1(n14598), .A2(n21341), .ZN(n33417) );
  XOR2_X1 U19129 ( .A1(n23429), .A2(n16053), .Z(n4792) );
  NAND2_X2 U19130 ( .A1(n31365), .A2(n30433), .ZN(n16053) );
  INV_X2 U19131 ( .I(n33175), .ZN(n28329) );
  XNOR2_X1 U19138 ( .A1(n2024), .A2(n30190), .ZN(n33175) );
  XOR2_X1 U19139 ( .A1(n28999), .A2(n24388), .Z(n34073) );
  XOR2_X1 U19140 ( .A1(n24478), .A2(n24622), .Z(n24388) );
  NAND4_X1 U19143 ( .A1(n14637), .A2(n14763), .A3(n16578), .A4(n14635), .ZN(
        n33701) );
  AOI21_X2 U19144 ( .A1(n28330), .A2(n5178), .B(n7047), .ZN(n11466) );
  XOR2_X1 U19147 ( .A1(n10960), .A2(n30098), .Z(n21970) );
  INV_X1 U19152 ( .I(n15559), .ZN(n33215) );
  NOR2_X2 U19154 ( .A1(n22732), .A2(n22730), .ZN(n3668) );
  AOI21_X2 U19155 ( .A1(n21902), .A2(n22488), .B(n31551), .ZN(n22732) );
  NOR2_X2 U19156 ( .A1(n23326), .A2(n33177), .ZN(n31772) );
  OAI21_X2 U19163 ( .A1(n32006), .A2(n27219), .B(n33178), .ZN(n33177) );
  NAND2_X2 U19165 ( .A1(n23322), .A2(n27219), .ZN(n33178) );
  NOR2_X2 U19167 ( .A1(n33179), .A2(n4453), .ZN(n23143) );
  AOI22_X1 U19170 ( .A1(n25008), .A2(n24998), .B1(n15016), .B2(n15078), .ZN(
        n25000) );
  NAND2_X2 U19171 ( .A1(n10612), .A2(n9737), .ZN(n22372) );
  XOR2_X1 U19173 ( .A1(n2192), .A2(n1482), .Z(n1481) );
  XOR2_X1 U19178 ( .A1(n2198), .A2(n16331), .Z(n2192) );
  AOI21_X2 U19179 ( .A1(n16295), .A2(n2778), .B(n6295), .ZN(n15808) );
  NAND2_X2 U19180 ( .A1(n18711), .A2(n328), .ZN(n2778) );
  XOR2_X1 U19182 ( .A1(n11781), .A2(n33181), .Z(n11780) );
  XOR2_X1 U19183 ( .A1(n6454), .A2(n2896), .Z(n33181) );
  NOR2_X2 U19188 ( .A1(n15054), .A2(n25247), .ZN(n33353) );
  INV_X2 U19189 ( .I(n5544), .ZN(n25247) );
  NAND3_X2 U19193 ( .A1(n28117), .A2(n2214), .A3(n17925), .ZN(n5544) );
  OR2_X1 U19195 ( .A1(n15790), .A2(n33182), .Z(n23999) );
  OR2_X1 U19197 ( .A1(n33183), .A2(n22443), .Z(n6837) );
  XOR2_X1 U19203 ( .A1(n22282), .A2(n3395), .Z(n33202) );
  XOR2_X1 U19204 ( .A1(n22274), .A2(n22028), .Z(n22282) );
  NOR2_X2 U19207 ( .A1(n31640), .A2(n25062), .ZN(n25041) );
  XOR2_X1 U19210 ( .A1(n17552), .A2(n19536), .Z(n11251) );
  NAND2_X1 U19212 ( .A1(n25644), .A2(n34094), .ZN(n25646) );
  OAI22_X2 U19215 ( .A1(n33185), .A2(n1962), .B1(n20551), .B2(n26343), .ZN(
        n21009) );
  NOR3_X2 U19219 ( .A1(n20550), .A2(n31232), .A3(n125), .ZN(n33185) );
  OAI21_X2 U19221 ( .A1(n14437), .A2(n13796), .B(n33186), .ZN(n19241) );
  OAI21_X2 U19225 ( .A1(n1054), .A2(n26603), .B(n13796), .ZN(n33186) );
  AOI22_X1 U19227 ( .A1(n25432), .A2(n11640), .B1(n25453), .B2(n25433), .ZN(
        n25434) );
  XNOR2_X1 U19229 ( .A1(n231), .A2(n7619), .ZN(n33264) );
  NAND2_X2 U19230 ( .A1(n33980), .A2(n29801), .ZN(n5462) );
  NOR2_X2 U19231 ( .A1(n27973), .A2(n33188), .ZN(n27504) );
  OAI22_X2 U19241 ( .A1(n17438), .A2(n21060), .B1(n21222), .B2(n21061), .ZN(
        n33188) );
  INV_X2 U19244 ( .I(n33189), .ZN(n11063) );
  XNOR2_X1 U19248 ( .A1(n26769), .A2(n4263), .ZN(n33189) );
  NAND3_X2 U19254 ( .A1(n33191), .A2(n22299), .A3(n33190), .ZN(n13622) );
  NAND2_X1 U19257 ( .A1(n8136), .A2(n10757), .ZN(n33191) );
  NOR2_X2 U19258 ( .A1(n21566), .A2(n17274), .ZN(n33611) );
  NAND2_X2 U19260 ( .A1(n33192), .A2(n1788), .ZN(n1787) );
  AOI21_X2 U19265 ( .A1(n1774), .A2(n20200), .B(n1789), .ZN(n33193) );
  XOR2_X1 U19267 ( .A1(n8581), .A2(n11691), .Z(n20762) );
  NOR2_X2 U19275 ( .A1(n13573), .A2(n13572), .ZN(n8581) );
  AOI21_X1 U19280 ( .A1(n18737), .A2(n12166), .B(n16287), .ZN(n13026) );
  NAND2_X2 U19286 ( .A1(n33195), .A2(n33194), .ZN(n14027) );
  NOR2_X1 U19289 ( .A1(n17240), .A2(n24975), .ZN(n26020) );
  NOR2_X1 U19291 ( .A1(n14812), .A2(n14811), .ZN(n6637) );
  NAND2_X2 U19294 ( .A1(n17253), .A2(n17254), .ZN(n14812) );
  AND2_X2 U19301 ( .A1(n14001), .A2(n10371), .Z(n24351) );
  NOR2_X2 U19304 ( .A1(n23877), .A2(n23878), .ZN(n15245) );
  NOR2_X1 U19306 ( .A1(n3565), .A2(n25763), .ZN(n24448) );
  XOR2_X1 U19308 ( .A1(n24619), .A2(n5253), .Z(n8656) );
  NAND2_X2 U19309 ( .A1(n6982), .A2(n33197), .ZN(n7198) );
  INV_X2 U19310 ( .I(n31942), .ZN(n17501) );
  NAND2_X2 U19312 ( .A1(n33863), .A2(n92), .ZN(n23005) );
  XOR2_X1 U19319 ( .A1(n23454), .A2(n7520), .Z(n28493) );
  NAND2_X1 U19324 ( .A1(n33198), .A2(n14164), .ZN(n15207) );
  NAND2_X1 U19325 ( .A1(n23578), .A2(n16981), .ZN(n33198) );
  NAND2_X1 U19330 ( .A1(n11898), .A2(n24610), .ZN(n33199) );
  XOR2_X1 U19332 ( .A1(n1003), .A2(n22028), .Z(n22275) );
  XOR2_X1 U19336 ( .A1(n33201), .A2(n33200), .Z(n30042) );
  XOR2_X1 U19337 ( .A1(n14733), .A2(n6833), .Z(n33201) );
  AND2_X1 U19343 ( .A1(n29158), .A2(n28924), .Z(n33865) );
  NAND3_X1 U19349 ( .A1(n10295), .A2(n4750), .A3(n5274), .ZN(n27544) );
  XOR2_X1 U19353 ( .A1(n33203), .A2(n16060), .Z(n22285) );
  NAND2_X2 U19354 ( .A1(n1874), .A2(n11595), .ZN(n7066) );
  NAND2_X2 U19355 ( .A1(n5593), .A2(n7103), .ZN(n13347) );
  XOR2_X1 U19357 ( .A1(n26872), .A2(n34146), .Z(n9690) );
  XOR2_X1 U19361 ( .A1(n4285), .A2(n22138), .Z(n12980) );
  NOR2_X2 U19368 ( .A1(n3578), .A2(n3579), .ZN(n4285) );
  AOI22_X1 U19370 ( .A1(n6830), .A2(n6829), .B1(n6828), .B2(n1075), .ZN(n6827)
         );
  XOR2_X1 U19373 ( .A1(n8885), .A2(n32083), .Z(n21248) );
  XOR2_X1 U19374 ( .A1(n20837), .A2(n33204), .Z(n30778) );
  INV_X2 U19381 ( .I(n21007), .ZN(n33204) );
  NAND2_X2 U19390 ( .A1(n17431), .A2(n9076), .ZN(n11619) );
  NAND2_X2 U19404 ( .A1(n33262), .A2(n30105), .ZN(n15806) );
  OAI21_X1 U19405 ( .A1(n18738), .A2(n33208), .B(n33207), .ZN(n18736) );
  OAI21_X1 U19407 ( .A1(n26369), .A2(n11792), .B(n21233), .ZN(n33209) );
  XOR2_X1 U19410 ( .A1(n33210), .A2(n24798), .Z(n18155) );
  XOR2_X1 U19412 ( .A1(n24797), .A2(n31440), .Z(n33210) );
  NAND2_X2 U19415 ( .A1(n33212), .A2(n33211), .ZN(n15787) );
  AOI22_X1 U19419 ( .A1(n18907), .A2(n1056), .B1(n12128), .B2(n10227), .ZN(
        n33211) );
  NAND2_X1 U19430 ( .A1(n2517), .A2(n764), .ZN(n33212) );
  XOR2_X1 U19431 ( .A1(n33213), .A2(n32930), .Z(n31296) );
  XOR2_X1 U19439 ( .A1(n19487), .A2(n19737), .Z(n33213) );
  XOR2_X1 U19440 ( .A1(n33214), .A2(n30951), .Z(n29064) );
  INV_X4 U19451 ( .I(n9575), .ZN(n33382) );
  XOR2_X1 U19453 ( .A1(n15), .A2(n2989), .Z(n1986) );
  NAND2_X2 U19455 ( .A1(n21240), .A2(n11601), .ZN(n13152) );
  OAI22_X2 U19456 ( .A1(n21431), .A2(n21070), .B1(n21241), .B2(n606), .ZN(
        n21240) );
  NAND2_X2 U19457 ( .A1(n31418), .A2(n27411), .ZN(n4580) );
  INV_X1 U19461 ( .I(n28177), .ZN(n23424) );
  INV_X2 U19462 ( .I(n3260), .ZN(n10294) );
  OAI22_X2 U19466 ( .A1(n9711), .A2(n9677), .B1(n9710), .B2(n9709), .ZN(n3260)
         );
  NAND2_X2 U19471 ( .A1(n26404), .A2(n15019), .ZN(n23087) );
  NAND2_X2 U19475 ( .A1(n15831), .A2(n32002), .ZN(n17334) );
  NAND2_X2 U19481 ( .A1(n31264), .A2(n11954), .ZN(n12548) );
  NAND2_X2 U19484 ( .A1(n23998), .A2(n23997), .ZN(n14490) );
  NAND3_X2 U19486 ( .A1(n14047), .A2(n23914), .A3(n26221), .ZN(n23998) );
  XOR2_X1 U19488 ( .A1(n16060), .A2(n3682), .Z(n33217) );
  NAND3_X1 U19489 ( .A1(n11710), .A2(n13693), .A3(n28390), .ZN(n33218) );
  BUF_X2 U19493 ( .I(n16331), .Z(n33219) );
  XOR2_X1 U19494 ( .A1(n11124), .A2(n33220), .Z(n11175) );
  XOR2_X1 U19498 ( .A1(n30671), .A2(n11126), .Z(n33220) );
  XOR2_X1 U19505 ( .A1(n23324), .A2(n3322), .Z(n23041) );
  NAND2_X1 U19506 ( .A1(n25430), .A2(n25444), .ZN(n31141) );
  NOR2_X1 U19507 ( .A1(n8219), .A2(n3339), .ZN(n3732) );
  XOR2_X1 U19511 ( .A1(n24689), .A2(n27153), .Z(n24758) );
  NAND2_X2 U19516 ( .A1(n2691), .A2(n31553), .ZN(n24689) );
  INV_X4 U19519 ( .I(n10899), .ZN(n13349) );
  XOR2_X1 U19524 ( .A1(n12557), .A2(n33673), .Z(n14798) );
  INV_X1 U19532 ( .I(n1892), .ZN(n33223) );
  XOR2_X1 U19534 ( .A1(n22104), .A2(n28612), .Z(n6466) );
  NOR2_X2 U19537 ( .A1(n33226), .A2(n31396), .ZN(n33284) );
  NAND2_X1 U19541 ( .A1(n22500), .A2(n33227), .ZN(n26762) );
  XOR2_X1 U19544 ( .A1(n27792), .A2(n5126), .Z(n30333) );
  OAI21_X1 U19552 ( .A1(n16430), .A2(n3759), .B(n11888), .ZN(n34075) );
  XOR2_X1 U19554 ( .A1(n33233), .A2(n33975), .Z(n22367) );
  XOR2_X1 U19556 ( .A1(n12370), .A2(n22301), .Z(n33233) );
  NAND3_X1 U19563 ( .A1(n33962), .A2(n736), .A3(n33961), .ZN(n25336) );
  NAND2_X1 U19567 ( .A1(n4983), .A2(n2486), .ZN(n33379) );
  NAND2_X2 U19569 ( .A1(n8178), .A2(n1931), .ZN(n24263) );
  NAND2_X1 U19571 ( .A1(n24254), .A2(n2558), .ZN(n24255) );
  NAND2_X2 U19573 ( .A1(n16957), .A2(n25334), .ZN(n13698) );
  NAND2_X1 U19582 ( .A1(n17028), .A2(n66), .ZN(n28531) );
  NAND2_X2 U19583 ( .A1(n16041), .A2(n72), .ZN(n25316) );
  XOR2_X1 U19585 ( .A1(n2345), .A2(n17048), .Z(n33235) );
  XOR2_X1 U19586 ( .A1(n23310), .A2(n13888), .Z(n33236) );
  OR2_X1 U19590 ( .A1(n29494), .A2(n26098), .Z(n33238) );
  NAND2_X1 U19593 ( .A1(n31052), .A2(n7003), .ZN(n2636) );
  NOR2_X2 U19601 ( .A1(n6364), .A2(n6365), .ZN(n33239) );
  AOI22_X2 U19602 ( .A1(n19944), .A2(n2694), .B1(n17882), .B2(n16681), .ZN(
        n33241) );
  NAND3_X2 U19603 ( .A1(n22920), .A2(n12887), .A3(n22924), .ZN(n9963) );
  NAND2_X2 U19605 ( .A1(n29507), .A2(n12888), .ZN(n22920) );
  AOI22_X2 U19606 ( .A1(n22880), .A2(n33344), .B1(n32092), .B2(n8365), .ZN(
        n9791) );
  AND2_X1 U19608 ( .A1(n14335), .A2(n13147), .Z(n3288) );
  NOR2_X2 U19618 ( .A1(n33611), .A2(n29875), .ZN(n33243) );
  OAI21_X2 U19621 ( .A1(n5679), .A2(n5954), .B(n33244), .ZN(n4151) );
  XOR2_X1 U19622 ( .A1(n33892), .A2(n600), .Z(n6627) );
  NOR3_X1 U19629 ( .A1(n23841), .A2(n23840), .A3(n17234), .ZN(n31083) );
  INV_X2 U19630 ( .I(n33246), .ZN(n34156) );
  XOR2_X1 U19634 ( .A1(n5321), .A2(n30427), .Z(n33246) );
  INV_X2 U19635 ( .I(n33247), .ZN(n23767) );
  XOR2_X1 U19636 ( .A1(n10347), .A2(n12331), .Z(n33247) );
  XOR2_X1 U19637 ( .A1(n13496), .A2(n15438), .Z(n10200) );
  NAND3_X2 U19638 ( .A1(n17036), .A2(n19931), .A3(n17035), .ZN(n16515) );
  XOR2_X1 U19643 ( .A1(n7078), .A2(n27922), .Z(n26812) );
  XOR2_X1 U19644 ( .A1(n23291), .A2(n5512), .Z(n5511) );
  OAI22_X2 U19645 ( .A1(n27835), .A2(n27834), .B1(n22614), .B2(n22813), .ZN(
        n23291) );
  OAI21_X2 U19648 ( .A1(n2722), .A2(n5289), .B(n2721), .ZN(n33766) );
  XOR2_X1 U19649 ( .A1(n33248), .A2(n25457), .Z(Ciphertext[107]) );
  NAND2_X2 U19650 ( .A1(n29920), .A2(n33249), .ZN(n26881) );
  XOR2_X1 U19651 ( .A1(n22100), .A2(n22121), .Z(n17586) );
  NAND2_X2 U19653 ( .A1(n21725), .A2(n21724), .ZN(n22100) );
  XOR2_X1 U19654 ( .A1(n17797), .A2(n33250), .Z(n23944) );
  XOR2_X1 U19659 ( .A1(n33895), .A2(n23316), .Z(n33250) );
  NAND2_X2 U19669 ( .A1(n33251), .A2(n6311), .ZN(n17423) );
  AOI22_X2 U19683 ( .A1(n8242), .A2(n9014), .B1(n20629), .B2(n9255), .ZN(
        n33251) );
  NAND2_X2 U19693 ( .A1(n13196), .A2(n23953), .ZN(n4823) );
  XOR2_X1 U19695 ( .A1(n33253), .A2(n33252), .Z(n33269) );
  NAND2_X2 U19698 ( .A1(n25490), .A2(n25473), .ZN(n25464) );
  NOR2_X2 U19700 ( .A1(n84), .A2(n24672), .ZN(n25490) );
  AOI21_X1 U19703 ( .A1(n29748), .A2(n24052), .B(n24182), .ZN(n18179) );
  OAI21_X2 U19712 ( .A1(n33255), .A2(n33254), .B(n18889), .ZN(n11302) );
  NOR2_X2 U19713 ( .A1(n18886), .A2(n18887), .ZN(n33254) );
  NOR2_X2 U19714 ( .A1(n13349), .A2(n4993), .ZN(n15555) );
  INV_X2 U19722 ( .I(n33256), .ZN(n9630) );
  XOR2_X1 U19723 ( .A1(n4395), .A2(n22292), .Z(n33256) );
  OAI21_X1 U19731 ( .A1(n33257), .A2(n28246), .B(n16957), .ZN(n30025) );
  INV_X1 U19732 ( .I(n16850), .ZN(n33257) );
  OAI21_X2 U19739 ( .A1(n26038), .A2(n419), .B(n28279), .ZN(n33258) );
  XOR2_X1 U19741 ( .A1(n23361), .A2(n23362), .Z(n23366) );
  XOR2_X1 U19742 ( .A1(n23328), .A2(n7070), .Z(n23362) );
  NOR2_X2 U19744 ( .A1(n29328), .A2(n31531), .ZN(n2130) );
  OAI22_X2 U19748 ( .A1(n26422), .A2(n3999), .B1(n23002), .B2(n13159), .ZN(
        n23004) );
  XOR2_X1 U19764 ( .A1(n33259), .A2(n29108), .Z(n2108) );
  XOR2_X1 U19769 ( .A1(n33860), .A2(n24593), .Z(n33259) );
  OAI21_X2 U19770 ( .A1(n32011), .A2(n33261), .B(n17606), .ZN(n28674) );
  OAI22_X2 U19771 ( .A1(n1595), .A2(n21692), .B1(n21691), .B2(n2708), .ZN(
        n22113) );
  INV_X2 U19777 ( .I(n24031), .ZN(n1241) );
  OAI21_X2 U19778 ( .A1(n7384), .A2(n7383), .B(n6308), .ZN(n24031) );
  OAI22_X2 U19780 ( .A1(n34080), .A2(n17975), .B1(n19841), .B2(n10057), .ZN(
        n2198) );
  NOR2_X1 U19782 ( .A1(n28037), .A2(n33263), .ZN(n5858) );
  NAND2_X1 U19786 ( .A1(n32111), .A2(n26974), .ZN(n1734) );
  XOR2_X1 U19787 ( .A1(n24620), .A2(n12800), .Z(n24489) );
  NAND2_X2 U19796 ( .A1(n10777), .A2(n15570), .ZN(n24620) );
  XOR2_X1 U19797 ( .A1(n23291), .A2(n5212), .Z(n23403) );
  NAND2_X2 U19798 ( .A1(n9243), .A2(n9244), .ZN(n5212) );
  NOR2_X2 U19802 ( .A1(n31930), .A2(n18079), .ZN(n11659) );
  BUF_X2 U19804 ( .I(n15710), .Z(n33265) );
  OAI21_X2 U19806 ( .A1(n18970), .A2(n18600), .B(n33266), .ZN(n28806) );
  AOI22_X2 U19812 ( .A1(n6639), .A2(n19156), .B1(n6637), .B2(n6638), .ZN(
        n33266) );
  NAND2_X2 U19814 ( .A1(n5343), .A2(n17873), .ZN(n15114) );
  XOR2_X1 U19822 ( .A1(n22779), .A2(n23400), .Z(n33267) );
  XOR2_X1 U19829 ( .A1(n11514), .A2(n33268), .Z(n30570) );
  XOR2_X1 U19836 ( .A1(n30792), .A2(n1741), .Z(n33268) );
  INV_X2 U19839 ( .I(n33269), .ZN(n17157) );
  XOR2_X1 U19840 ( .A1(n3395), .A2(n27601), .Z(n2953) );
  NAND2_X2 U19842 ( .A1(n11904), .A2(n17661), .ZN(n17374) );
  XOR2_X1 U19843 ( .A1(n1923), .A2(n29167), .Z(n20870) );
  XOR2_X1 U19844 ( .A1(n5148), .A2(n101), .Z(n17380) );
  XOR2_X1 U19846 ( .A1(n5150), .A2(n29130), .Z(n5148) );
  INV_X2 U19847 ( .I(n33270), .ZN(n34157) );
  XOR2_X1 U19850 ( .A1(n14887), .A2(n17643), .Z(n33270) );
  XOR2_X1 U19851 ( .A1(n10780), .A2(n19486), .Z(n12145) );
  XOR2_X1 U19854 ( .A1(n26778), .A2(n11691), .Z(n20772) );
  AOI22_X2 U19861 ( .A1(n26466), .A2(n7041), .B1(n7064), .B2(n25704), .ZN(
        n9496) );
  NAND2_X2 U19863 ( .A1(n29503), .A2(n10733), .ZN(n28429) );
  NOR2_X2 U19864 ( .A1(n33272), .A2(n33271), .ZN(n26814) );
  NOR2_X2 U19871 ( .A1(n5825), .A2(n2288), .ZN(n33272) );
  NOR2_X2 U19873 ( .A1(n15150), .A2(n33273), .ZN(n24909) );
  AOI21_X2 U19876 ( .A1(n24362), .A2(n11945), .B(n33053), .ZN(n33273) );
  OR2_X1 U19877 ( .A1(n12290), .A2(n14926), .Z(n28383) );
  INV_X1 U19879 ( .I(n4790), .ZN(n33274) );
  XOR2_X1 U19881 ( .A1(n23388), .A2(n23499), .Z(n4790) );
  XOR2_X1 U19893 ( .A1(n17235), .A2(n33275), .Z(n23886) );
  XOR2_X1 U19896 ( .A1(n23460), .A2(n643), .Z(n33275) );
  XOR2_X1 U19897 ( .A1(n23469), .A2(n33276), .Z(n28031) );
  XOR2_X1 U19898 ( .A1(n31354), .A2(n23388), .Z(n33276) );
  NAND2_X1 U19904 ( .A1(n24974), .A2(n33278), .ZN(n33277) );
  INV_X2 U19911 ( .I(n24610), .ZN(n33278) );
  XOR2_X1 U19915 ( .A1(n24692), .A2(n29639), .Z(n29638) );
  XOR2_X1 U19919 ( .A1(n24533), .A2(n16141), .Z(n24692) );
  INV_X2 U19922 ( .I(n33279), .ZN(n7993) );
  XNOR2_X1 U19925 ( .A1(n5158), .A2(n5159), .ZN(n33279) );
  NAND2_X2 U19927 ( .A1(n33284), .A2(n5258), .ZN(n1808) );
  NAND2_X2 U19934 ( .A1(n21996), .A2(n8269), .ZN(n33285) );
  NAND3_X2 U19935 ( .A1(n22512), .A2(n22513), .A3(n22600), .ZN(n14044) );
  NAND2_X2 U19937 ( .A1(n6837), .A2(n33287), .ZN(n31894) );
  NAND4_X2 U19941 ( .A1(n22569), .A2(n7053), .A3(n22443), .A4(n22442), .ZN(
        n33287) );
  NOR2_X1 U19944 ( .A1(n9059), .A2(n7753), .ZN(n9058) );
  OAI22_X2 U19950 ( .A1(n21445), .A2(n6277), .B1(n21101), .B2(n16526), .ZN(
        n26622) );
  XOR2_X1 U19954 ( .A1(n23478), .A2(n12714), .Z(n27866) );
  XOR2_X1 U19956 ( .A1(n22157), .A2(n30275), .Z(n7911) );
  NAND2_X2 U19958 ( .A1(n115), .A2(n34084), .ZN(n30275) );
  NAND2_X1 U19966 ( .A1(n12006), .A2(n32901), .ZN(n18695) );
  XOR2_X1 U19970 ( .A1(n7045), .A2(n15183), .Z(n23145) );
  INV_X2 U19971 ( .I(n33289), .ZN(n26712) );
  XNOR2_X1 U19981 ( .A1(n13294), .A2(n13293), .ZN(n33289) );
  XOR2_X1 U19990 ( .A1(n6090), .A2(n33290), .Z(n31411) );
  XOR2_X1 U19991 ( .A1(n31499), .A2(n33823), .Z(n33290) );
  NAND2_X2 U19996 ( .A1(n7817), .A2(n135), .ZN(n22832) );
  AOI22_X2 U20001 ( .A1(n7169), .A2(n10498), .B1(n17580), .B2(n23885), .ZN(
        n24248) );
  XOR2_X1 U20007 ( .A1(n21891), .A2(n22256), .Z(n33291) );
  XOR2_X1 U20010 ( .A1(n5925), .A2(n19727), .Z(n29486) );
  XOR2_X1 U20011 ( .A1(n19386), .A2(n19403), .Z(n19727) );
  INV_X2 U20019 ( .I(n33292), .ZN(n4378) );
  XOR2_X1 U20023 ( .A1(n4379), .A2(n4380), .Z(n33292) );
  XOR2_X1 U20024 ( .A1(n12785), .A2(n16662), .Z(n14237) );
  NOR2_X2 U20025 ( .A1(n20636), .A2(n26907), .ZN(n20652) );
  AOI22_X2 U20026 ( .A1(n33294), .A2(n6985), .B1(n13411), .B2(n13592), .ZN(
        n3786) );
  XOR2_X1 U20030 ( .A1(n2894), .A2(n30331), .Z(n13198) );
  NAND2_X2 U20037 ( .A1(n26261), .A2(n3469), .ZN(n30331) );
  XOR2_X1 U20040 ( .A1(n10650), .A2(n33437), .Z(n22118) );
  NAND2_X2 U20045 ( .A1(n33676), .A2(n16014), .ZN(n33437) );
  BUF_X2 U20046 ( .I(n24138), .Z(n33295) );
  NAND3_X2 U20047 ( .A1(n31025), .A2(n8046), .A3(n14618), .ZN(n21738) );
  INV_X2 U20050 ( .I(n33296), .ZN(n26084) );
  XOR2_X1 U20055 ( .A1(n19395), .A2(n19230), .Z(n33296) );
  NAND2_X2 U20061 ( .A1(n31583), .A2(n33297), .ZN(n31473) );
  AOI21_X2 U20067 ( .A1(n8712), .A2(n8711), .B(n25633), .ZN(n31830) );
  NAND2_X2 U20073 ( .A1(n6835), .A2(n6836), .ZN(n29317) );
  OAI21_X2 U20076 ( .A1(n2986), .A2(n2987), .B(n29821), .ZN(n13320) );
  OR2_X1 U20089 ( .A1(n31034), .A2(n26170), .Z(n6309) );
  NAND2_X2 U20100 ( .A1(n10832), .A2(n33299), .ZN(n31325) );
  XOR2_X1 U20102 ( .A1(n21903), .A2(n31606), .Z(n33300) );
  NAND2_X2 U20106 ( .A1(n1567), .A2(n25152), .ZN(n30615) );
  NAND2_X2 U20107 ( .A1(n13028), .A2(n21498), .ZN(n13113) );
  BUF_X2 U20108 ( .I(n23807), .Z(n33302) );
  AND2_X1 U20109 ( .A1(n30282), .A2(n31915), .Z(n6042) );
  XOR2_X1 U20111 ( .A1(n33303), .A2(n3739), .Z(n15372) );
  NAND2_X1 U20114 ( .A1(n25177), .A2(n8929), .ZN(n33428) );
  OAI22_X2 U20115 ( .A1(n9404), .A2(n20165), .B1(n20164), .B2(n20476), .ZN(
        n33373) );
  NOR2_X2 U20116 ( .A1(n23966), .A2(n23967), .ZN(n29767) );
  NOR2_X2 U20122 ( .A1(n29834), .A2(n23771), .ZN(n23966) );
  AOI22_X2 U20128 ( .A1(n33221), .A2(n28306), .B1(n23722), .B2(n847), .ZN(
        n33304) );
  XOR2_X1 U20131 ( .A1(n16837), .A2(n536), .Z(n6175) );
  NAND2_X2 U20143 ( .A1(n33305), .A2(n5926), .ZN(n10385) );
  NAND2_X1 U20144 ( .A1(n9885), .A2(n15411), .ZN(n13252) );
  OAI22_X2 U20145 ( .A1(n1449), .A2(n34141), .B1(n26378), .B2(n1446), .ZN(
        n15411) );
  NAND2_X2 U20151 ( .A1(n33306), .A2(n22699), .ZN(n23282) );
  NOR2_X2 U20152 ( .A1(n33314), .A2(n34115), .ZN(n31895) );
  INV_X2 U20159 ( .I(n14612), .ZN(n12715) );
  NAND3_X2 U20160 ( .A1(n12418), .A2(n12781), .A3(n12417), .ZN(n14612) );
  NAND2_X1 U20166 ( .A1(n33308), .A2(n7023), .ZN(n11031) );
  OAI21_X1 U20170 ( .A1(n22491), .A2(n16225), .B(n27897), .ZN(n33308) );
  NOR2_X1 U20171 ( .A1(n29098), .A2(n29099), .ZN(n33569) );
  XOR2_X1 U20172 ( .A1(n28822), .A2(n29042), .Z(n20443) );
  INV_X2 U20175 ( .I(n11097), .ZN(n33310) );
  INV_X1 U20176 ( .I(n1018), .ZN(n30267) );
  INV_X4 U20194 ( .I(n21780), .ZN(n31220) );
  NAND2_X2 U20196 ( .A1(n15443), .A2(n33695), .ZN(n21780) );
  XOR2_X1 U20202 ( .A1(n3847), .A2(n12765), .Z(n12764) );
  BUF_X2 U20209 ( .I(n22537), .Z(n33312) );
  NAND2_X2 U20212 ( .A1(n33313), .A2(n23727), .ZN(n3880) );
  NAND3_X1 U20214 ( .A1(n7269), .A2(n7425), .A3(n7268), .ZN(n33318) );
  OAI21_X1 U20219 ( .A1(n996), .A2(n22667), .B(n22580), .ZN(n4994) );
  OAI21_X2 U20221 ( .A1(n31926), .A2(n32588), .B(n32499), .ZN(n33315) );
  INV_X2 U20223 ( .I(n11754), .ZN(n24118) );
  XOR2_X1 U20224 ( .A1(n12980), .A2(n33316), .Z(n8885) );
  XOR2_X1 U20226 ( .A1(n1308), .A2(n21892), .Z(n33316) );
  XOR2_X1 U20237 ( .A1(n9131), .A2(n23470), .Z(n33317) );
  INV_X4 U20238 ( .I(n654), .ZN(n34009) );
  OAI22_X2 U20242 ( .A1(n29342), .A2(n1124), .B1(n22542), .B2(n22397), .ZN(
        n8991) );
  NAND2_X2 U20247 ( .A1(n6257), .A2(n33739), .ZN(n29342) );
  NAND3_X1 U20248 ( .A1(n33318), .A2(n7265), .A3(n7266), .ZN(Ciphertext[181])
         );
  XOR2_X1 U20251 ( .A1(n14532), .A2(n24806), .Z(n33319) );
  AOI21_X2 U20252 ( .A1(n27947), .A2(n25630), .B(n31974), .ZN(n31604) );
  NAND2_X2 U20253 ( .A1(n26585), .A2(n17497), .ZN(n20495) );
  AOI22_X2 U20257 ( .A1(n12161), .A2(n34046), .B1(n396), .B2(n29454), .ZN(
        n33321) );
  INV_X1 U20258 ( .I(n2618), .ZN(n1348) );
  NAND2_X2 U20259 ( .A1(n9403), .A2(n33288), .ZN(n2618) );
  NAND2_X2 U20267 ( .A1(n33323), .A2(n30857), .ZN(n14720) );
  NAND2_X1 U20268 ( .A1(n29339), .A2(n29250), .ZN(n29872) );
  XOR2_X1 U20271 ( .A1(n8728), .A2(n13606), .Z(n20977) );
  NAND3_X2 U20281 ( .A1(n5734), .A2(n20408), .A3(n10290), .ZN(n13606) );
  AND2_X1 U20283 ( .A1(n33325), .A2(n15296), .Z(n21531) );
  NAND2_X2 U20286 ( .A1(n17715), .A2(n10925), .ZN(n29337) );
  XOR2_X1 U20287 ( .A1(Plaintext[10]), .A2(Key[10]), .Z(n8213) );
  XOR2_X1 U20290 ( .A1(n33326), .A2(n20916), .Z(n52) );
  XOR2_X1 U20293 ( .A1(n20792), .A2(n30163), .Z(n33326) );
  NAND2_X2 U20295 ( .A1(n7780), .A2(n29606), .ZN(n7778) );
  OR2_X1 U20297 ( .A1(n11820), .A2(n25531), .Z(n33327) );
  OR2_X1 U20299 ( .A1(n25724), .A2(n13640), .Z(n2962) );
  NOR2_X2 U20301 ( .A1(n11511), .A2(n14352), .ZN(n25724) );
  XOR2_X1 U20304 ( .A1(n33328), .A2(n19648), .Z(n31900) );
  XOR2_X1 U20305 ( .A1(n17129), .A2(n25993), .Z(n33328) );
  NAND3_X2 U20306 ( .A1(n33302), .A2(n23850), .A3(n3241), .ZN(n33457) );
  INV_X2 U20310 ( .I(n33329), .ZN(n758) );
  NAND2_X2 U20317 ( .A1(n22810), .A2(n12729), .ZN(n22694) );
  NAND2_X2 U20324 ( .A1(n13972), .A2(n22424), .ZN(n22810) );
  OAI21_X2 U20326 ( .A1(n10747), .A2(n25233), .B(n11132), .ZN(n33330) );
  XOR2_X1 U20327 ( .A1(n1707), .A2(n33331), .Z(n15865) );
  AND2_X1 U20328 ( .A1(n6118), .A2(n9766), .Z(n7726) );
  NAND2_X2 U20329 ( .A1(n16920), .A2(n16918), .ZN(n23355) );
  AOI22_X2 U20333 ( .A1(n30243), .A2(n29286), .B1(n15747), .B2(n21514), .ZN(
        n10233) );
  AOI21_X2 U20336 ( .A1(n23006), .A2(n3999), .B(n23004), .ZN(n7070) );
  XOR2_X1 U20338 ( .A1(n20987), .A2(n33332), .Z(n3298) );
  OAI22_X2 U20342 ( .A1(n14996), .A2(n14997), .B1(n14999), .B2(n14998), .ZN(
        n21761) );
  XOR2_X1 U20348 ( .A1(n32516), .A2(n29155), .Z(n33333) );
  XOR2_X1 U20349 ( .A1(n9464), .A2(n33334), .Z(n30214) );
  XOR2_X1 U20350 ( .A1(n26715), .A2(n28295), .Z(n33334) );
  BUF_X2 U20352 ( .I(n30781), .Z(n33335) );
  NAND2_X2 U20355 ( .A1(n1816), .A2(n1819), .ZN(n24220) );
  NAND2_X2 U20371 ( .A1(n30354), .A2(n14463), .ZN(n1816) );
  NAND2_X2 U20374 ( .A1(n33336), .A2(n27270), .ZN(n3266) );
  XOR2_X1 U20377 ( .A1(n5600), .A2(n22027), .Z(n33338) );
  XOR2_X1 U20381 ( .A1(n9904), .A2(n11102), .Z(n33339) );
  NAND2_X2 U20383 ( .A1(n11492), .A2(n11491), .ZN(n30651) );
  XOR2_X1 U20384 ( .A1(n15889), .A2(n15891), .Z(n14029) );
  XOR2_X1 U20387 ( .A1(n20848), .A2(n20729), .Z(n5724) );
  NAND2_X2 U20388 ( .A1(n26212), .A2(n29672), .ZN(n20848) );
  XOR2_X1 U20389 ( .A1(n5979), .A2(n3957), .Z(n9203) );
  NAND2_X2 U20401 ( .A1(n3440), .A2(n3439), .ZN(n13357) );
  NOR3_X2 U20403 ( .A1(n28276), .A2(n26969), .A3(n1180), .ZN(n31246) );
  OR2_X1 U20408 ( .A1(n3468), .A2(n8784), .Z(n26265) );
  NAND2_X2 U20414 ( .A1(n4878), .A2(n18897), .ZN(n29030) );
  NAND3_X2 U20419 ( .A1(n4611), .A2(n33686), .A3(n17774), .ZN(n15183) );
  NAND2_X1 U20420 ( .A1(n7751), .A2(n33069), .ZN(n8193) );
  NAND2_X2 U20421 ( .A1(n33342), .A2(n28888), .ZN(n3994) );
  NOR2_X2 U20424 ( .A1(n9016), .A2(n9017), .ZN(n33342) );
  NAND3_X1 U20426 ( .A1(n24924), .A2(n30328), .A3(n24925), .ZN(n33343) );
  XOR2_X1 U20428 ( .A1(n10196), .A2(n10194), .Z(n18220) );
  XOR2_X1 U20429 ( .A1(n22015), .A2(n4342), .Z(n12614) );
  NAND3_X1 U20430 ( .A1(n25449), .A2(n33658), .A3(n25447), .ZN(n33469) );
  NAND2_X2 U20436 ( .A1(n23864), .A2(n10993), .ZN(n23930) );
  XOR2_X1 U20438 ( .A1(n2917), .A2(n2918), .Z(n29288) );
  NOR2_X1 U20439 ( .A1(n25818), .A2(n25804), .ZN(n25811) );
  NAND2_X2 U20448 ( .A1(n11185), .A2(n12420), .ZN(n25804) );
  NAND3_X2 U20450 ( .A1(n22620), .A2(n33347), .A3(n33346), .ZN(n16073) );
  NAND2_X2 U20462 ( .A1(n33349), .A2(n31403), .ZN(n25863) );
  AOI21_X1 U20463 ( .A1(n21503), .A2(n13028), .B(n30346), .ZN(n21504) );
  NAND2_X2 U20465 ( .A1(n2570), .A2(n30403), .ZN(n34046) );
  XOR2_X1 U20469 ( .A1(n24801), .A2(n7603), .Z(n24567) );
  AOI21_X2 U20471 ( .A1(n4786), .A2(n11732), .B(n33350), .ZN(n4785) );
  XOR2_X1 U20486 ( .A1(n19728), .A2(n12223), .Z(n17193) );
  XOR2_X1 U20487 ( .A1(n19625), .A2(n19530), .Z(n12223) );
  XOR2_X1 U20499 ( .A1(n24388), .A2(n29140), .Z(n4418) );
  NAND3_X2 U20500 ( .A1(n12605), .A2(n12604), .A3(n5384), .ZN(n9536) );
  NOR2_X1 U20502 ( .A1(n34009), .A2(n32308), .ZN(n8849) );
  NAND2_X2 U20504 ( .A1(n8848), .A2(n8851), .ZN(n24159) );
  XOR2_X1 U20506 ( .A1(n17153), .A2(n8109), .Z(n33351) );
  XNOR2_X1 U20514 ( .A1(n16897), .A2(n21888), .ZN(n33975) );
  NAND2_X2 U20516 ( .A1(n1579), .A2(n1580), .ZN(n22960) );
  NAND2_X1 U20517 ( .A1(n28722), .A2(n7083), .ZN(n28990) );
  NAND2_X1 U20518 ( .A1(n25657), .A2(n25665), .ZN(n28722) );
  INV_X2 U20519 ( .I(n29042), .ZN(n30163) );
  NAND2_X2 U20522 ( .A1(n2620), .A2(n11412), .ZN(n29042) );
  INV_X2 U20525 ( .I(n24779), .ZN(n14627) );
  NAND2_X1 U20530 ( .A1(n13650), .A2(n13649), .ZN(n2293) );
  INV_X2 U20531 ( .I(n23385), .ZN(n26426) );
  NAND2_X2 U20537 ( .A1(n14466), .A2(n14465), .ZN(n23385) );
  INV_X2 U20540 ( .I(n33354), .ZN(n10193) );
  XOR2_X1 U20541 ( .A1(n7191), .A2(n33355), .Z(n15057) );
  XOR2_X1 U20545 ( .A1(n7193), .A2(n15157), .Z(n33355) );
  OAI22_X2 U20546 ( .A1(n33357), .A2(n33356), .B1(n13325), .B2(n26343), .ZN(
        n13696) );
  INV_X1 U20547 ( .I(n6475), .ZN(n33356) );
  XOR2_X1 U20554 ( .A1(n21027), .A2(n13338), .Z(n33358) );
  XOR2_X1 U20559 ( .A1(n24505), .A2(n6897), .Z(n33359) );
  AOI22_X2 U20564 ( .A1(n11705), .A2(n11704), .B1(n9548), .B2(n11703), .ZN(
        n16509) );
  NAND2_X2 U20567 ( .A1(n21087), .A2(n21209), .ZN(n21382) );
  OR2_X1 U20571 ( .A1(n18064), .A2(n12895), .Z(n9661) );
  NAND2_X2 U20573 ( .A1(n19910), .A2(n17633), .ZN(n20960) );
  NAND2_X1 U20577 ( .A1(n4066), .A2(n19158), .ZN(n13059) );
  NAND3_X1 U20578 ( .A1(n7968), .A2(n25999), .A3(n8233), .ZN(n19130) );
  NAND2_X1 U20579 ( .A1(n33360), .A2(n15456), .ZN(n26705) );
  NAND2_X2 U20582 ( .A1(n16134), .A2(n16133), .ZN(n14485) );
  XOR2_X1 U20584 ( .A1(n33361), .A2(n25929), .Z(Ciphertext[191]) );
  OAI22_X1 U20586 ( .A1(n25927), .A2(n25926), .B1(n25924), .B2(n25925), .ZN(
        n33361) );
  NAND2_X2 U20590 ( .A1(n20433), .A2(n20431), .ZN(n14365) );
  XOR2_X1 U20591 ( .A1(n33362), .A2(n14584), .Z(n5692) );
  XOR2_X1 U20593 ( .A1(n34120), .A2(n23533), .Z(n33362) );
  XOR2_X1 U20598 ( .A1(n5522), .A2(n5523), .Z(n29936) );
  INV_X2 U20605 ( .I(n33363), .ZN(n11784) );
  XOR2_X1 U20607 ( .A1(n22063), .A2(n9960), .Z(n33363) );
  NAND2_X2 U20621 ( .A1(n33365), .A2(n33364), .ZN(n21742) );
  NAND2_X2 U20625 ( .A1(n33367), .A2(n33366), .ZN(n33365) );
  INV_X2 U20628 ( .I(n423), .ZN(n33366) );
  NAND2_X2 U20633 ( .A1(n3854), .A2(n33368), .ZN(n33869) );
  XOR2_X1 U20634 ( .A1(n17765), .A2(n15821), .Z(n17879) );
  XOR2_X1 U20636 ( .A1(n23438), .A2(n23439), .Z(n3514) );
  NAND2_X2 U20637 ( .A1(n17460), .A2(n17458), .ZN(n23438) );
  INV_X2 U20644 ( .I(n2940), .ZN(n8924) );
  XOR2_X1 U20648 ( .A1(n2926), .A2(n2924), .Z(n2940) );
  XOR2_X1 U20649 ( .A1(n22229), .A2(n22230), .Z(n11282) );
  XOR2_X1 U20654 ( .A1(n22305), .A2(n22308), .Z(n22230) );
  XOR2_X1 U20656 ( .A1(n7057), .A2(n1984), .Z(n19578) );
  AOI21_X2 U20658 ( .A1(n33555), .A2(n19003), .B(n7749), .ZN(n1984) );
  XOR2_X1 U20663 ( .A1(n32478), .A2(n21028), .Z(n20787) );
  INV_X2 U20666 ( .I(n29296), .ZN(n30504) );
  OAI21_X2 U20669 ( .A1(n6631), .A2(n20144), .B(n6630), .ZN(n29296) );
  XNOR2_X1 U20671 ( .A1(n16303), .A2(n4028), .ZN(n33427) );
  NAND2_X2 U20672 ( .A1(n23556), .A2(n5685), .ZN(n29499) );
  XOR2_X1 U20674 ( .A1(n6348), .A2(n1708), .Z(n1707) );
  XOR2_X1 U20685 ( .A1(n20778), .A2(n31185), .Z(n33369) );
  NAND2_X2 U20694 ( .A1(n30222), .A2(n26576), .ZN(n31477) );
  NAND2_X2 U20696 ( .A1(n12315), .A2(n3614), .ZN(n22762) );
  NAND2_X2 U20700 ( .A1(n22418), .A2(n33582), .ZN(n12315) );
  OAI21_X2 U20701 ( .A1(n11714), .A2(n11715), .B(n19009), .ZN(n11177) );
  INV_X2 U20706 ( .I(n31511), .ZN(n31007) );
  NAND2_X2 U20708 ( .A1(n13292), .A2(n34158), .ZN(n31511) );
  NOR3_X1 U20717 ( .A1(n22634), .A2(n28979), .A3(n7513), .ZN(n18012) );
  NAND2_X2 U20718 ( .A1(n33370), .A2(n17387), .ZN(n24250) );
  OR2_X2 U20725 ( .A1(n8444), .A2(n9968), .Z(n24361) );
  NAND2_X2 U20728 ( .A1(n16639), .A2(n26712), .ZN(n21326) );
  XOR2_X1 U20729 ( .A1(n10758), .A2(n33371), .Z(n17014) );
  XOR2_X1 U20731 ( .A1(n23441), .A2(n23442), .Z(n33371) );
  NAND2_X1 U20734 ( .A1(n27594), .A2(n3016), .ZN(n33372) );
  NAND3_X1 U20748 ( .A1(n18752), .A2(n18753), .A3(n18983), .ZN(n18754) );
  NAND2_X2 U20753 ( .A1(n31850), .A2(n16288), .ZN(n18752) );
  XOR2_X1 U20754 ( .A1(n15093), .A2(n15934), .Z(n27182) );
  OAI21_X2 U20758 ( .A1(n15650), .A2(n4850), .B(n30106), .ZN(n30105) );
  XOR2_X1 U20760 ( .A1(n23363), .A2(n23385), .Z(n23463) );
  NAND2_X2 U20762 ( .A1(n29266), .A2(n16635), .ZN(n23363) );
  XOR2_X1 U20765 ( .A1(n33374), .A2(n19371), .Z(n19439) );
  INV_X2 U20766 ( .I(n19599), .ZN(n33374) );
  NAND2_X2 U20769 ( .A1(n7440), .A2(n7439), .ZN(n19371) );
  XOR2_X1 U20770 ( .A1(n33375), .A2(n24787), .Z(n8152) );
  NAND2_X2 U20771 ( .A1(n14309), .A2(n5115), .ZN(n24995) );
  XOR2_X1 U20776 ( .A1(n33377), .A2(n33376), .Z(n26284) );
  XOR2_X1 U20780 ( .A1(n9346), .A2(n31252), .Z(n33377) );
  NAND2_X2 U20784 ( .A1(n33832), .A2(n7581), .ZN(n24091) );
  XOR2_X1 U20795 ( .A1(n33378), .A2(n29447), .Z(n11248) );
  XOR2_X1 U20801 ( .A1(n19493), .A2(n34071), .Z(n33378) );
  INV_X1 U20803 ( .I(n25891), .ZN(n33474) );
  OAI21_X2 U20807 ( .A1(n10556), .A2(n16795), .B(n20043), .ZN(n17241) );
  XOR2_X1 U20808 ( .A1(n4020), .A2(n23537), .Z(n28407) );
  INV_X2 U20809 ( .I(n16310), .ZN(n33687) );
  XOR2_X1 U20811 ( .A1(n33381), .A2(n7572), .Z(n1942) );
  XOR2_X1 U20812 ( .A1(n5127), .A2(n31410), .Z(n33381) );
  OAI21_X2 U20813 ( .A1(n28543), .A2(n28544), .B(n33206), .ZN(n3900) );
  NOR2_X1 U20819 ( .A1(n4180), .A2(n29908), .ZN(n17714) );
  XOR2_X1 U20820 ( .A1(n22044), .A2(n9536), .Z(n8630) );
  NAND2_X2 U20822 ( .A1(n33384), .A2(n24613), .ZN(n8622) );
  OAI21_X2 U20829 ( .A1(n15231), .A2(n28815), .B(n15232), .ZN(n33384) );
  NAND2_X2 U20837 ( .A1(n33738), .A2(n33385), .ZN(n14002) );
  BUF_X2 U20841 ( .I(n13684), .Z(n33386) );
  AND2_X1 U20842 ( .A1(n25711), .A2(n4449), .Z(n13924) );
  NAND2_X2 U20845 ( .A1(n30044), .A2(n14856), .ZN(n14201) );
  AOI21_X1 U20846 ( .A1(n3717), .A2(n15522), .B(n12323), .ZN(n21058) );
  AOI22_X2 U20848 ( .A1(n13026), .A2(n17599), .B1(n13025), .B2(n13024), .ZN(
        n19274) );
  NAND2_X2 U20849 ( .A1(n28484), .A2(n28829), .ZN(n20990) );
  XNOR2_X1 U20856 ( .A1(n19389), .A2(n31882), .ZN(n26300) );
  OAI21_X1 U20857 ( .A1(n29432), .A2(n17964), .B(n742), .ZN(n15168) );
  NOR2_X2 U20859 ( .A1(n33390), .A2(n26874), .ZN(n16321) );
  INV_X2 U20862 ( .I(n33391), .ZN(n26641) );
  NAND2_X2 U20864 ( .A1(n25332), .A2(n16783), .ZN(n15624) );
  NAND2_X2 U20866 ( .A1(n33394), .A2(n33393), .ZN(n25332) );
  INV_X2 U20873 ( .I(n28093), .ZN(n33393) );
  NAND2_X2 U20876 ( .A1(n31886), .A2(n31572), .ZN(n34116) );
  OR2_X1 U20891 ( .A1(n26345), .A2(n4755), .Z(n12441) );
  OAI21_X2 U20893 ( .A1(n327), .A2(n17473), .B(n22443), .ZN(n13127) );
  NAND2_X2 U20894 ( .A1(n327), .A2(n27959), .ZN(n22443) );
  NOR2_X2 U20896 ( .A1(n11235), .A2(n22748), .ZN(n17707) );
  AOI22_X2 U20905 ( .A1(n33398), .A2(n33397), .B1(n7290), .B2(n15217), .ZN(
        n13547) );
  XOR2_X1 U20910 ( .A1(n33401), .A2(n16674), .Z(Ciphertext[118]) );
  XOR2_X1 U20911 ( .A1(n2854), .A2(n7832), .Z(n2857) );
  NAND2_X2 U20912 ( .A1(n6945), .A2(n33402), .ZN(n22945) );
  NAND2_X1 U20914 ( .A1(n9991), .A2(n10754), .ZN(n9990) );
  XOR2_X1 U20916 ( .A1(n14588), .A2(n1464), .Z(n9006) );
  NAND2_X2 U20921 ( .A1(n29581), .A2(n29580), .ZN(n1464) );
  AND3_X1 U20923 ( .A1(n20109), .A2(n33848), .A3(n8421), .Z(n2906) );
  BUF_X2 U20933 ( .I(n21755), .Z(n33403) );
  XOR2_X1 U20935 ( .A1(n31495), .A2(n33404), .Z(n31453) );
  XOR2_X1 U20949 ( .A1(n19541), .A2(n19471), .Z(n33404) );
  NOR2_X2 U20954 ( .A1(n33405), .A2(n13610), .ZN(n20545) );
  OAI21_X2 U20955 ( .A1(n11414), .A2(n33419), .B(n5470), .ZN(n13610) );
  INV_X1 U20956 ( .I(n33406), .ZN(n33405) );
  NAND2_X1 U20957 ( .A1(n13611), .A2(n12078), .ZN(n33406) );
  NOR2_X2 U20959 ( .A1(n14649), .A2(n26890), .ZN(n33407) );
  XOR2_X1 U20961 ( .A1(n23337), .A2(n23146), .Z(n2842) );
  XOR2_X1 U20962 ( .A1(n17775), .A2(n14077), .Z(n23337) );
  XOR2_X1 U20965 ( .A1(n1607), .A2(n30407), .Z(n33408) );
  XOR2_X1 U20968 ( .A1(n4728), .A2(n24839), .Z(n31340) );
  NAND2_X2 U20980 ( .A1(n3234), .A2(n28522), .ZN(n24839) );
  OAI22_X2 U20982 ( .A1(n21666), .A2(n1134), .B1(n31089), .B2(n1136), .ZN(
        n33409) );
  OAI21_X2 U20983 ( .A1(n33411), .A2(n33410), .B(n983), .ZN(n22768) );
  NOR2_X1 U20984 ( .A1(n33818), .A2(n641), .ZN(n33410) );
  INV_X1 U20985 ( .I(n6227), .ZN(n33411) );
  NOR2_X2 U20988 ( .A1(n24001), .A2(n24000), .ZN(n3220) );
  NAND3_X2 U20990 ( .A1(n15957), .A2(n18632), .A3(n33412), .ZN(n30781) );
  NAND2_X2 U20991 ( .A1(n33413), .A2(n33650), .ZN(n28736) );
  OR2_X1 U20992 ( .A1(n22491), .A2(n630), .Z(n21902) );
  INV_X2 U20994 ( .I(n33415), .ZN(n18496) );
  NOR2_X2 U20998 ( .A1(n17223), .A2(n17255), .ZN(n33415) );
  NOR3_X2 U21000 ( .A1(n5549), .A2(n5550), .A3(n33416), .ZN(n5548) );
  NOR3_X2 U21003 ( .A1(n30554), .A2(n19926), .A3(n4587), .ZN(n33416) );
  XOR2_X1 U21007 ( .A1(n14662), .A2(n8343), .Z(n28027) );
  AND2_X1 U21011 ( .A1(n386), .A2(n23745), .Z(n30895) );
  XOR2_X1 U21012 ( .A1(n2335), .A2(n28039), .Z(n13510) );
  OAI22_X2 U21016 ( .A1(n11538), .A2(n11539), .B1(n30875), .B2(n11540), .ZN(
        n23456) );
  XOR2_X1 U21020 ( .A1(n10758), .A2(n9671), .Z(n9670) );
  XOR2_X1 U21023 ( .A1(n23229), .A2(n26108), .Z(n28286) );
  XOR2_X1 U21024 ( .A1(n23419), .A2(n646), .Z(n23229) );
  NAND2_X2 U21028 ( .A1(n27272), .A2(n11752), .ZN(n18084) );
  INV_X4 U21035 ( .I(n33420), .ZN(n3944) );
  NOR2_X2 U21036 ( .A1(n3946), .A2(n3945), .ZN(n33420) );
  AND2_X1 U21043 ( .A1(n20375), .A2(n20374), .Z(n12225) );
  NAND2_X2 U21053 ( .A1(n30996), .A2(n2492), .ZN(n20375) );
  NAND2_X2 U21055 ( .A1(n33423), .A2(n27711), .ZN(n10732) );
  XOR2_X1 U21059 ( .A1(n20862), .A2(n16831), .Z(n21049) );
  NOR2_X2 U21060 ( .A1(n29993), .A2(n4061), .ZN(n20862) );
  XOR2_X1 U21062 ( .A1(n31200), .A2(n33424), .Z(n8694) );
  XOR2_X1 U21064 ( .A1(n16382), .A2(n23342), .Z(n33424) );
  INV_X1 U21071 ( .I(n33446), .ZN(n23851) );
  AND2_X1 U21072 ( .A1(n33446), .A2(n663), .Z(n5817) );
  NAND2_X2 U21078 ( .A1(n11385), .A2(n4760), .ZN(n2611) );
  XOR2_X1 U21080 ( .A1(n30535), .A2(n33426), .Z(n33803) );
  XOR2_X1 U21082 ( .A1(n23359), .A2(n32015), .Z(n33426) );
  XOR2_X1 U21086 ( .A1(n17307), .A2(n17308), .Z(n6434) );
  XOR2_X1 U21087 ( .A1(n12454), .A2(n12414), .Z(n24838) );
  XNOR2_X1 U21094 ( .A1(n7016), .A2(n21010), .ZN(n33521) );
  INV_X2 U21105 ( .I(n33429), .ZN(n34153) );
  XOR2_X1 U21107 ( .A1(n3070), .A2(n3074), .Z(n33429) );
  XOR2_X1 U21111 ( .A1(n8637), .A2(n2072), .Z(n31395) );
  INV_X2 U21113 ( .I(n33430), .ZN(n29252) );
  XOR2_X1 U21121 ( .A1(n19407), .A2(n8383), .Z(n33430) );
  NAND2_X2 U21124 ( .A1(n31970), .A2(n7197), .ZN(n11072) );
  NAND2_X1 U21126 ( .A1(n3979), .A2(n7502), .ZN(n33954) );
  OAI21_X2 U21127 ( .A1(n10757), .A2(n1124), .B(n10288), .ZN(n33433) );
  NOR2_X2 U21132 ( .A1(n26474), .A2(n17431), .ZN(n17428) );
  NAND2_X2 U21133 ( .A1(n27016), .A2(n33435), .ZN(n16278) );
  AOI22_X2 U21137 ( .A1(n7115), .A2(n21427), .B1(n21072), .B2(n21341), .ZN(
        n33435) );
  AOI21_X2 U21140 ( .A1(n20598), .A2(n5993), .B(n31401), .ZN(n20913) );
  XOR2_X1 U21142 ( .A1(n10026), .A2(n19627), .Z(n19723) );
  NAND2_X1 U21144 ( .A1(n33436), .A2(n8171), .ZN(n27585) );
  NOR2_X1 U21145 ( .A1(n27806), .A2(n20578), .ZN(n33436) );
  NOR2_X2 U21149 ( .A1(n10227), .A2(n764), .ZN(n18907) );
  NAND2_X1 U21150 ( .A1(n33586), .A2(n8957), .ZN(n8955) );
  OAI21_X2 U21156 ( .A1(n23112), .A2(n17099), .B(n33438), .ZN(n9041) );
  NAND3_X1 U21166 ( .A1(n6453), .A2(n23109), .A3(n16022), .ZN(n33438) );
  INV_X2 U21168 ( .I(n28702), .ZN(n4274) );
  XOR2_X1 U21173 ( .A1(n5138), .A2(n5137), .Z(n5188) );
  XOR2_X1 U21176 ( .A1(n2808), .A2(n33715), .Z(n17245) );
  XNOR2_X1 U21180 ( .A1(n23272), .A2(n23441), .ZN(n13190) );
  NAND2_X2 U21185 ( .A1(n4174), .A2(n5233), .ZN(n23272) );
  NAND2_X1 U21186 ( .A1(n7973), .A2(n33440), .ZN(n387) );
  AOI21_X1 U21192 ( .A1(n16397), .A2(n837), .B(n13763), .ZN(n33440) );
  INV_X2 U21197 ( .I(n19102), .ZN(n27617) );
  NAND2_X2 U21199 ( .A1(n18923), .A2(n19101), .ZN(n19102) );
  NAND2_X2 U21207 ( .A1(n28139), .A2(n5250), .ZN(n17888) );
  AND2_X1 U21208 ( .A1(n2697), .A2(n1119), .Z(n33854) );
  OR2_X1 U21210 ( .A1(n29944), .A2(n19991), .Z(n33441) );
  NOR2_X2 U21213 ( .A1(n30833), .A2(n12213), .ZN(n23007) );
  NAND2_X2 U21225 ( .A1(n18473), .A2(n15148), .ZN(n19057) );
  XOR2_X1 U21226 ( .A1(n3599), .A2(n19513), .Z(n19731) );
  NAND2_X2 U21247 ( .A1(n18928), .A2(n18927), .ZN(n19513) );
  NAND2_X1 U21249 ( .A1(n25621), .A2(n17499), .ZN(n33442) );
  INV_X1 U21251 ( .I(n31569), .ZN(n33443) );
  AOI22_X2 U21256 ( .A1(n18226), .A2(n18731), .B1(n18733), .B2(n18730), .ZN(
        n18225) );
  NOR2_X2 U21259 ( .A1(n957), .A2(n26155), .ZN(n18226) );
  INV_X2 U21268 ( .I(n33849), .ZN(n34089) );
  XOR2_X1 U21270 ( .A1(n13122), .A2(n32067), .Z(n33849) );
  NOR2_X2 U21272 ( .A1(n33444), .A2(n24012), .ZN(n31919) );
  NAND3_X2 U21273 ( .A1(n33445), .A2(n8591), .A3(n2391), .ZN(n31805) );
  NAND2_X2 U21303 ( .A1(n940), .A2(n4233), .ZN(n33445) );
  NOR2_X2 U21306 ( .A1(n13147), .A2(n17799), .ZN(n33446) );
  INV_X2 U21307 ( .I(n27894), .ZN(n10899) );
  XOR2_X1 U21310 ( .A1(n23476), .A2(n25881), .Z(n30955) );
  NAND2_X2 U21311 ( .A1(n2636), .A2(n2637), .ZN(n23476) );
  XOR2_X1 U21316 ( .A1(n19163), .A2(n19446), .Z(n4052) );
  XOR2_X1 U21323 ( .A1(n33448), .A2(n15117), .Z(n19163) );
  INV_X2 U21325 ( .I(n31731), .ZN(n33448) );
  XOR2_X1 U21327 ( .A1(n27362), .A2(n11483), .Z(n11548) );
  XOR2_X1 U21332 ( .A1(n19469), .A2(n33449), .Z(n10696) );
  XOR2_X1 U21334 ( .A1(n16792), .A2(n9503), .Z(n33449) );
  NAND2_X2 U21345 ( .A1(n4635), .A2(n4638), .ZN(n28011) );
  AOI22_X2 U21346 ( .A1(n7773), .A2(n8041), .B1(n5858), .B2(n5857), .ZN(n21512) );
  XOR2_X1 U21347 ( .A1(n26865), .A2(n7380), .Z(n2915) );
  XOR2_X1 U21349 ( .A1(n24450), .A2(n24409), .Z(n8691) );
  NAND2_X2 U21352 ( .A1(n1960), .A2(n1963), .ZN(n20873) );
  NOR2_X2 U21353 ( .A1(n1926), .A2(n1805), .ZN(n22280) );
  OAI22_X2 U21358 ( .A1(n33450), .A2(n20249), .B1(n16308), .B2(n28257), .ZN(
        n21743) );
  NOR2_X1 U21364 ( .A1(n15172), .A2(n21581), .ZN(n30652) );
  NAND2_X2 U21366 ( .A1(n14704), .A2(n15997), .ZN(n15720) );
  OAI21_X2 U21367 ( .A1(n4435), .A2(n4434), .B(n33451), .ZN(n22036) );
  AOI22_X2 U21377 ( .A1(n4432), .A2(n33242), .B1(n21697), .B2(n4433), .ZN(
        n33451) );
  XOR2_X1 U21383 ( .A1(n19598), .A2(n19647), .Z(n15776) );
  XOR2_X1 U21384 ( .A1(n4437), .A2(n33452), .Z(n16272) );
  XOR2_X1 U21389 ( .A1(n28441), .A2(n31754), .Z(n33452) );
  BUF_X2 U21392 ( .I(n24635), .Z(n33453) );
  AOI22_X2 U21393 ( .A1(n31080), .A2(n1681), .B1(n4301), .B2(n14927), .ZN(
        n1680) );
  OAI22_X2 U21401 ( .A1(n33456), .A2(n33455), .B1(n9647), .B2(n16529), .ZN(
        n4084) );
  OAI21_X1 U21416 ( .A1(n28240), .A2(n24031), .B(n24304), .ZN(n24033) );
  XOR2_X1 U21421 ( .A1(n30273), .A2(n29169), .Z(n31251) );
  XOR2_X1 U21423 ( .A1(n22005), .A2(n22067), .Z(n22288) );
  NAND2_X2 U21427 ( .A1(n2913), .A2(n24316), .ZN(n33458) );
  XOR2_X1 U21433 ( .A1(n23419), .A2(n4732), .Z(n4564) );
  NAND2_X2 U21435 ( .A1(n31434), .A2(n14769), .ZN(n23419) );
  NAND2_X2 U21442 ( .A1(n33462), .A2(n11340), .ZN(n30795) );
  NOR2_X2 U21444 ( .A1(n28391), .A2(n32094), .ZN(n33462) );
  AOI22_X2 U21466 ( .A1(n33463), .A2(n6649), .B1(n13369), .B2(n29823), .ZN(
        n29952) );
  NOR2_X1 U21467 ( .A1(n16290), .A2(n26061), .ZN(n33464) );
  XOR2_X1 U21469 ( .A1(n33465), .A2(n23501), .Z(n33550) );
  NAND2_X2 U21470 ( .A1(n26883), .A2(n17923), .ZN(n24207) );
  XOR2_X1 U21484 ( .A1(n24504), .A2(n24681), .Z(n6898) );
  XOR2_X1 U21489 ( .A1(n24830), .A2(n27114), .Z(n24681) );
  INV_X2 U21492 ( .I(n21326), .ZN(n1142) );
  XOR2_X1 U21493 ( .A1(n9218), .A2(n20964), .Z(n9217) );
  NAND2_X1 U21496 ( .A1(n5672), .A2(n5632), .ZN(n5671) );
  XOR2_X1 U21498 ( .A1(n17745), .A2(n22046), .Z(n3303) );
  OAI21_X1 U21499 ( .A1(n2858), .A2(n5961), .B(n33466), .ZN(n33485) );
  INV_X2 U21508 ( .I(n22606), .ZN(n33466) );
  NAND2_X2 U21517 ( .A1(n11402), .A2(n33467), .ZN(n12421) );
  OAI21_X2 U21518 ( .A1(n12397), .A2(n19819), .B(n12396), .ZN(n33467) );
  AOI22_X2 U21520 ( .A1(n22566), .A2(n13409), .B1(n22564), .B2(n16490), .ZN(
        n22971) );
  NAND2_X2 U21521 ( .A1(n11874), .A2(n12530), .ZN(n13409) );
  NOR2_X2 U21524 ( .A1(n28379), .A2(n19137), .ZN(n28543) );
  XOR2_X1 U21525 ( .A1(n23470), .A2(n33960), .Z(n33959) );
  NAND2_X2 U21538 ( .A1(n27701), .A2(n2803), .ZN(n23470) );
  AOI22_X2 U21539 ( .A1(n3494), .A2(n31345), .B1(n3911), .B2(n3495), .ZN(
        n28083) );
  NOR2_X2 U21547 ( .A1(n28378), .A2(n10612), .ZN(n3911) );
  NOR2_X1 U21548 ( .A1(n3348), .A2(n33503), .ZN(n28002) );
  XOR2_X1 U21550 ( .A1(n13802), .A2(n21898), .Z(n7114) );
  OAI22_X2 U21557 ( .A1(n12151), .A2(n28773), .B1(n12153), .B2(n33687), .ZN(
        n27021) );
  XOR2_X1 U21569 ( .A1(n33469), .A2(n25450), .Z(Ciphertext[106]) );
  NAND2_X2 U21573 ( .A1(n33471), .A2(n6514), .ZN(n22158) );
  INV_X2 U21574 ( .I(n4029), .ZN(n8784) );
  NAND2_X2 U21576 ( .A1(n29106), .A2(n7543), .ZN(n4029) );
  OAI21_X2 U21577 ( .A1(n33473), .A2(n31822), .B(n716), .ZN(n17022) );
  XOR2_X1 U21585 ( .A1(n31165), .A2(n22197), .Z(n14969) );
  NAND2_X2 U21586 ( .A1(n31037), .A2(n33475), .ZN(n24965) );
  NAND3_X1 U21591 ( .A1(n2886), .A2(n1221), .A3(n716), .ZN(n33475) );
  XOR2_X1 U21595 ( .A1(n33476), .A2(n34056), .Z(n33638) );
  OAI21_X2 U21597 ( .A1(n29570), .A2(n34168), .B(n32004), .ZN(n30394) );
  XOR2_X1 U21599 ( .A1(n33477), .A2(n20870), .Z(n14887) );
  XOR2_X1 U21601 ( .A1(n2055), .A2(n20955), .Z(n33477) );
  XOR2_X1 U21610 ( .A1(n3987), .A2(n33478), .Z(n29762) );
  XOR2_X1 U21612 ( .A1(n33574), .A2(n4997), .Z(n33478) );
  XOR2_X1 U21618 ( .A1(n33479), .A2(n12284), .Z(n31272) );
  XOR2_X1 U21623 ( .A1(n30492), .A2(n3617), .Z(n33479) );
  XOR2_X1 U21624 ( .A1(n14612), .A2(n23191), .Z(n23192) );
  INV_X2 U21626 ( .I(n6552), .ZN(n33480) );
  INV_X2 U21629 ( .I(n33482), .ZN(n10086) );
  XNOR2_X1 U21635 ( .A1(n2366), .A2(n2364), .ZN(n33482) );
  NOR2_X1 U21636 ( .A1(n15680), .A2(n21546), .ZN(n33483) );
  INV_X2 U21640 ( .I(n23150), .ZN(n1261) );
  NAND3_X2 U21641 ( .A1(n393), .A2(n18239), .A3(n28178), .ZN(n23150) );
  XOR2_X1 U21642 ( .A1(n10946), .A2(n11862), .Z(n12915) );
  XOR2_X1 U21647 ( .A1(n33484), .A2(n12896), .Z(n34122) );
  XOR2_X1 U21649 ( .A1(n19557), .A2(n27884), .Z(n33484) );
  XOR2_X1 U21670 ( .A1(n11781), .A2(n33486), .Z(n11641) );
  XOR2_X1 U21678 ( .A1(n10946), .A2(n22141), .Z(n33486) );
  XOR2_X1 U21692 ( .A1(n24810), .A2(n7879), .Z(n13858) );
  NAND2_X2 U21697 ( .A1(n6110), .A2(n5960), .ZN(n33760) );
  INV_X2 U21701 ( .I(n33487), .ZN(n29153) );
  NAND2_X2 U21705 ( .A1(n9171), .A2(n11785), .ZN(n33909) );
  AOI21_X2 U21712 ( .A1(n23812), .A2(n3860), .B(n11061), .ZN(n33488) );
  NOR2_X1 U21717 ( .A1(n33867), .A2(n23595), .ZN(n23584) );
  NAND2_X1 U21718 ( .A1(n9283), .A2(n9282), .ZN(n33489) );
  XOR2_X1 U21722 ( .A1(n23422), .A2(n23421), .Z(n33490) );
  NOR2_X2 U21736 ( .A1(n10973), .A2(n33491), .ZN(n10721) );
  NOR3_X1 U21744 ( .A1(n7007), .A2(n21379), .A3(n17313), .ZN(n33491) );
  XOR2_X1 U21745 ( .A1(n24562), .A2(n24563), .Z(n24564) );
  XOR2_X1 U21746 ( .A1(n26795), .A2(n24819), .Z(n24562) );
  NOR2_X2 U21748 ( .A1(n14189), .A2(n33494), .ZN(n25175) );
  XOR2_X1 U21749 ( .A1(n32648), .A2(n31950), .Z(n2785) );
  NAND2_X2 U21753 ( .A1(n349), .A2(n21218), .ZN(n33495) );
  OAI22_X2 U21754 ( .A1(n10871), .A2(n28825), .B1(n22606), .B2(n5961), .ZN(
        n6110) );
  XOR2_X1 U21755 ( .A1(n5186), .A2(n21011), .Z(n5185) );
  NOR2_X2 U21767 ( .A1(n33497), .A2(n31811), .ZN(n7154) );
  NOR2_X2 U21768 ( .A1(n20607), .A2(n7577), .ZN(n33497) );
  INV_X1 U21771 ( .I(n33501), .ZN(n17322) );
  AND2_X1 U21782 ( .A1(n1465), .A2(n33501), .Z(n34080) );
  INV_X2 U21783 ( .I(n13644), .ZN(n13681) );
  NAND2_X2 U21794 ( .A1(n7800), .A2(n31496), .ZN(n13644) );
  OR2_X1 U21796 ( .A1(n21392), .A2(n20882), .Z(n20883) );
  NOR2_X2 U21800 ( .A1(n20511), .A2(n16774), .ZN(n20730) );
  XOR2_X1 U21803 ( .A1(n33448), .A2(n19508), .Z(n19588) );
  NAND2_X2 U21807 ( .A1(n17507), .A2(n17509), .ZN(n19508) );
  NAND2_X2 U21812 ( .A1(n1684), .A2(n7392), .ZN(n20970) );
  OR2_X1 U21820 ( .A1(n18677), .A2(n18888), .Z(n10367) );
  NAND2_X2 U21825 ( .A1(n29089), .A2(n7316), .ZN(n5150) );
  OAI22_X2 U21831 ( .A1(n4994), .A2(n33502), .B1(n4996), .B2(n26878), .ZN(
        n15501) );
  XOR2_X1 U21832 ( .A1(n31597), .A2(n18189), .Z(n27633) );
  NAND2_X2 U21842 ( .A1(n10705), .A2(n14868), .ZN(n18189) );
  XOR2_X1 U21845 ( .A1(n8659), .A2(n23455), .Z(n7178) );
  NAND2_X2 U21848 ( .A1(n14371), .A2(n33505), .ZN(n17301) );
  NAND2_X2 U21851 ( .A1(n24189), .A2(n24186), .ZN(n8412) );
  XOR2_X1 U21856 ( .A1(n12653), .A2(n31638), .Z(n31468) );
  XOR2_X1 U21862 ( .A1(n33506), .A2(n16666), .Z(Ciphertext[81]) );
  NAND2_X1 U21863 ( .A1(n4226), .A2(n31281), .ZN(n33506) );
  INV_X2 U21865 ( .I(n33508), .ZN(n11869) );
  NOR2_X2 U21870 ( .A1(n5000), .A2(n5002), .ZN(n9300) );
  INV_X2 U21871 ( .I(n33510), .ZN(n29462) );
  XOR2_X1 U21900 ( .A1(n30747), .A2(n5482), .Z(n10519) );
  XOR2_X1 U21902 ( .A1(n33511), .A2(n4555), .Z(n17857) );
  XOR2_X1 U21903 ( .A1(n4554), .A2(n4559), .Z(n33511) );
  NOR2_X2 U21906 ( .A1(n5668), .A2(n5669), .ZN(n20690) );
  NAND2_X1 U21908 ( .A1(n33499), .A2(n17181), .ZN(n26570) );
  AND2_X1 U21909 ( .A1(n16809), .A2(n16380), .Z(n1949) );
  NAND2_X2 U21910 ( .A1(n24894), .A2(n14274), .ZN(n16809) );
  XOR2_X1 U21911 ( .A1(n33513), .A2(n16322), .Z(Ciphertext[136]) );
  XOR2_X1 U21912 ( .A1(n22141), .A2(n22055), .Z(n22206) );
  INV_X2 U21914 ( .I(n33514), .ZN(n12058) );
  NAND2_X2 U21923 ( .A1(n29976), .A2(n15641), .ZN(n33514) );
  NAND2_X1 U21926 ( .A1(n21427), .A2(n21338), .ZN(n21339) );
  NOR2_X2 U21935 ( .A1(n9994), .A2(n21826), .ZN(n28278) );
  NAND2_X2 U21938 ( .A1(n34015), .A2(n5687), .ZN(n21826) );
  BUF_X2 U21944 ( .I(n7102), .Z(n33515) );
  INV_X2 U21946 ( .I(n10001), .ZN(n819) );
  OAI22_X2 U21947 ( .A1(n1976), .A2(n16491), .B1(n1974), .B2(n10742), .ZN(
        n10001) );
  AND2_X1 U21948 ( .A1(n31437), .A2(n17462), .Z(n28777) );
  XOR2_X1 U21954 ( .A1(n2388), .A2(n19403), .Z(n19543) );
  OAI21_X2 U21955 ( .A1(n1871), .A2(n2390), .B(n16788), .ZN(n2388) );
  XOR2_X1 U21956 ( .A1(n33517), .A2(n24766), .Z(n15106) );
  XOR2_X1 U21960 ( .A1(n30358), .A2(n24764), .Z(n33517) );
  XOR2_X1 U21966 ( .A1(n30532), .A2(n23282), .Z(n23173) );
  XOR2_X1 U21971 ( .A1(n2072), .A2(n33518), .Z(n26854) );
  XOR2_X1 U21973 ( .A1(n8741), .A2(n29876), .Z(n33518) );
  NAND2_X2 U21974 ( .A1(n28463), .A2(n31006), .ZN(n3614) );
  XOR2_X1 U21975 ( .A1(Plaintext[168]), .A2(Key[168]), .Z(n17030) );
  XOR2_X1 U21978 ( .A1(n7015), .A2(n33521), .Z(n3879) );
  XOR2_X1 U21979 ( .A1(n10075), .A2(n10935), .Z(n12621) );
  NAND2_X2 U21981 ( .A1(n29729), .A2(n33524), .ZN(n6865) );
  NAND2_X2 U21993 ( .A1(n33526), .A2(n33525), .ZN(n33524) );
  NAND2_X2 U22001 ( .A1(n33527), .A2(n3087), .ZN(n3086) );
  NOR2_X2 U22003 ( .A1(n29659), .A2(n33558), .ZN(n33528) );
  NAND2_X2 U22004 ( .A1(n33529), .A2(n33730), .ZN(n3036) );
  INV_X2 U22005 ( .I(n10524), .ZN(n33529) );
  NAND2_X2 U22007 ( .A1(n31967), .A2(n3084), .ZN(n10524) );
  XOR2_X1 U22020 ( .A1(n1787), .A2(n14428), .Z(n11532) );
  AND2_X1 U22028 ( .A1(n24324), .A2(n30579), .Z(n2360) );
  NAND2_X2 U22031 ( .A1(n8), .A2(n8086), .ZN(n30579) );
  BUF_X2 U22032 ( .I(n29763), .Z(n33530) );
  XOR2_X1 U22037 ( .A1(n23529), .A2(n23287), .Z(n14584) );
  XOR2_X1 U22038 ( .A1(n4627), .A2(n15686), .Z(n17151) );
  INV_X2 U22044 ( .I(n33531), .ZN(n29688) );
  XOR2_X1 U22045 ( .A1(n5607), .A2(n5609), .Z(n33531) );
  XOR2_X1 U22053 ( .A1(n24760), .A2(n10084), .Z(n24743) );
  NAND3_X2 U22056 ( .A1(n8000), .A2(n8001), .A3(n24228), .ZN(n24760) );
  NAND3_X1 U22070 ( .A1(n4916), .A2(n34058), .A3(n14251), .ZN(n22351) );
  NOR2_X2 U22074 ( .A1(n16559), .A2(n12074), .ZN(n18641) );
  OR2_X1 U22077 ( .A1(n13431), .A2(n13430), .Z(n33533) );
  INV_X2 U22084 ( .I(n33534), .ZN(n4916) );
  NAND2_X2 U22091 ( .A1(n275), .A2(n9299), .ZN(n22318) );
  AOI21_X2 U22092 ( .A1(n11309), .A2(n23697), .B(n33535), .ZN(n11287) );
  XOR2_X1 U22099 ( .A1(n24422), .A2(n24423), .Z(n10172) );
  CLKBUF_X12 U22102 ( .I(n9870), .Z(n33536) );
  XOR2_X1 U22105 ( .A1(n21029), .A2(n12342), .Z(n20764) );
  NOR2_X2 U22110 ( .A1(n12343), .A2(n12344), .ZN(n12342) );
  NAND2_X2 U22113 ( .A1(n2961), .A2(n33537), .ZN(n13684) );
  INV_X2 U22114 ( .I(n33538), .ZN(n21160) );
  OAI22_X2 U22117 ( .A1(n18277), .A2(n18641), .B1(n18276), .B2(n4626), .ZN(
        n18279) );
  XOR2_X1 U22132 ( .A1(n14908), .A2(n16502), .Z(n15990) );
  NAND2_X2 U22140 ( .A1(n11070), .A2(n30743), .ZN(n14908) );
  AND2_X1 U22152 ( .A1(n17590), .A2(n21160), .Z(n12521) );
  XOR2_X1 U22155 ( .A1(n33539), .A2(n24798), .Z(n10209) );
  XOR2_X1 U22166 ( .A1(n24597), .A2(n27283), .Z(n33539) );
  NAND2_X1 U22183 ( .A1(n27514), .A2(n30673), .ZN(n33650) );
  OAI22_X2 U22185 ( .A1(n17767), .A2(n21078), .B1(n21079), .B2(n16933), .ZN(
        n15622) );
  NAND2_X2 U22189 ( .A1(n33541), .A2(n10928), .ZN(n23065) );
  NAND2_X1 U22190 ( .A1(n8427), .A2(n10654), .ZN(n33541) );
  AOI21_X2 U22218 ( .A1(n33542), .A2(n33830), .B(n23584), .ZN(n16643) );
  NOR2_X2 U22225 ( .A1(n6082), .A2(n21401), .ZN(n28426) );
  NAND2_X2 U22230 ( .A1(n21403), .A2(n596), .ZN(n21401) );
  NOR2_X2 U22231 ( .A1(n20070), .A2(n18036), .ZN(n27600) );
  XOR2_X1 U22236 ( .A1(n2520), .A2(n25879), .Z(n30421) );
  OAI22_X2 U22242 ( .A1(n2404), .A2(n2405), .B1(n17202), .B2(n22895), .ZN(
        n2520) );
  XOR2_X1 U22245 ( .A1(n2626), .A2(n33545), .Z(n18090) );
  XOR2_X1 U22247 ( .A1(n2628), .A2(n15188), .Z(n33545) );
  NAND2_X2 U22248 ( .A1(n18677), .A2(n10325), .ZN(n10364) );
  XOR2_X1 U22249 ( .A1(n23258), .A2(n23376), .Z(n23181) );
  OAI21_X2 U22254 ( .A1(n12529), .A2(n22906), .B(n14914), .ZN(n23258) );
  XOR2_X1 U22260 ( .A1(n32697), .A2(n19461), .Z(n5921) );
  NAND3_X2 U22261 ( .A1(n28372), .A2(n28371), .A3(n6193), .ZN(n31568) );
  INV_X1 U22264 ( .I(n1652), .ZN(n21461) );
  OAI22_X2 U22265 ( .A1(n28396), .A2(n21058), .B1(n21263), .B2(n11745), .ZN(
        n1652) );
  NAND2_X1 U22266 ( .A1(n15500), .A2(n15498), .ZN(n33546) );
  XOR2_X1 U22269 ( .A1(n18058), .A2(n22255), .Z(n17486) );
  XOR2_X1 U22270 ( .A1(n33547), .A2(n25567), .Z(Ciphertext[128]) );
  NAND4_X2 U22280 ( .A1(n10035), .A2(n37), .A3(n10039), .A4(n36), .ZN(n33547)
         );
  NOR2_X2 U22281 ( .A1(n12525), .A2(n20780), .ZN(n28420) );
  NAND2_X1 U22282 ( .A1(n10511), .A2(n10510), .ZN(n27282) );
  NAND3_X2 U22285 ( .A1(n10446), .A2(n10448), .A3(n10450), .ZN(n5762) );
  NAND3_X1 U22288 ( .A1(n22463), .A2(n22462), .A3(n22557), .ZN(n22464) );
  NAND2_X2 U22294 ( .A1(n22462), .A2(n22460), .ZN(n22463) );
  XOR2_X1 U22297 ( .A1(n31884), .A2(n16958), .Z(n2925) );
  NAND2_X2 U22302 ( .A1(n6775), .A2(n14366), .ZN(n16958) );
  NAND2_X2 U22303 ( .A1(n25025), .A2(n16293), .ZN(n25123) );
  OAI22_X2 U22305 ( .A1(n21571), .A2(n29806), .B1(n1012), .B2(n32039), .ZN(
        n3578) );
  XOR2_X1 U22310 ( .A1(n33550), .A2(n9550), .Z(n665) );
  XOR2_X1 U22313 ( .A1(n33552), .A2(n7596), .Z(n28236) );
  XOR2_X1 U22315 ( .A1(n30778), .A2(n3559), .Z(n33552) );
  XOR2_X1 U22316 ( .A1(n17301), .A2(n24442), .Z(n24825) );
  XOR2_X1 U22318 ( .A1(n7603), .A2(n24532), .Z(n7135) );
  NOR2_X2 U22326 ( .A1(n6334), .A2(n17067), .ZN(n24532) );
  AND2_X1 U22327 ( .A1(n18405), .A2(n5139), .Z(n3052) );
  OAI21_X2 U22335 ( .A1(n33553), .A2(n33909), .B(n5717), .ZN(n8087) );
  XOR2_X1 U22336 ( .A1(n24749), .A2(n33554), .Z(n7695) );
  XOR2_X1 U22337 ( .A1(n11651), .A2(n10070), .Z(n33554) );
  XOR2_X1 U22339 ( .A1(n16175), .A2(n20798), .Z(n9674) );
  XNOR2_X1 U22345 ( .A1(n31279), .A2(n25856), .ZN(n33838) );
  NAND3_X2 U22348 ( .A1(n5485), .A2(n2935), .A3(n19039), .ZN(n33555) );
  NAND2_X2 U22349 ( .A1(n33556), .A2(n26767), .ZN(n7045) );
  BUF_X2 U22352 ( .I(n24224), .Z(n33557) );
  NAND3_X1 U22354 ( .A1(n801), .A2(n28367), .A3(n23695), .ZN(n10160) );
  INV_X4 U22355 ( .I(n17930), .ZN(n896) );
  NAND2_X2 U22356 ( .A1(n3711), .A2(n34053), .ZN(n17930) );
  NOR2_X2 U22360 ( .A1(n33645), .A2(n7602), .ZN(n7604) );
  XOR2_X1 U22365 ( .A1(n20999), .A2(n21000), .Z(n21005) );
  INV_X2 U22366 ( .I(n28010), .ZN(n33558) );
  BUF_X2 U22378 ( .I(n578), .Z(n33561) );
  NOR2_X2 U22379 ( .A1(n33595), .A2(n29705), .ZN(n2005) );
  XOR2_X1 U22381 ( .A1(n1536), .A2(n1538), .Z(n7699) );
  XOR2_X1 U22385 ( .A1(n14181), .A2(n15561), .Z(n28312) );
  NAND2_X2 U22390 ( .A1(n11317), .A2(n4750), .ZN(n33562) );
  INV_X2 U22392 ( .I(n1112), .ZN(n33563) );
  XOR2_X1 U22394 ( .A1(n6746), .A2(n33575), .Z(n14398) );
  NAND2_X2 U22398 ( .A1(n7541), .A2(n33564), .ZN(n7802) );
  AOI22_X2 U22402 ( .A1(n13665), .A2(n13664), .B1(n26878), .B2(n908), .ZN(
        n33564) );
  NOR2_X2 U22422 ( .A1(n12168), .A2(n33264), .ZN(n33565) );
  NOR2_X2 U22431 ( .A1(n13541), .A2(n10398), .ZN(n19530) );
  XOR2_X1 U22438 ( .A1(n19672), .A2(n26683), .Z(n6156) );
  NAND2_X2 U22441 ( .A1(n28237), .A2(n14735), .ZN(n19672) );
  INV_X2 U22443 ( .I(n14321), .ZN(n24994) );
  NAND2_X2 U22445 ( .A1(n12679), .A2(n12678), .ZN(n14321) );
  AOI21_X2 U22454 ( .A1(n16873), .A2(n4210), .B(n16870), .ZN(n30411) );
  OR3_X1 U22456 ( .A1(n29695), .A2(n28812), .A3(n20489), .Z(n20254) );
  INV_X2 U22459 ( .I(n33570), .ZN(n27343) );
  BUF_X2 U22464 ( .I(n21820), .Z(n33571) );
  BUF_X2 U22466 ( .I(n22317), .Z(n33572) );
  NAND2_X2 U22468 ( .A1(n33573), .A2(n11008), .ZN(n13694) );
  NAND2_X1 U22472 ( .A1(n11010), .A2(n8252), .ZN(n33573) );
  NAND2_X1 U22473 ( .A1(n1619), .A2(n6003), .ZN(n33727) );
  XOR2_X1 U22478 ( .A1(n6745), .A2(n15424), .Z(n33575) );
  NAND2_X2 U22485 ( .A1(n33576), .A2(n9794), .ZN(n16147) );
  NOR2_X2 U22488 ( .A1(n2724), .A2(n2725), .ZN(n33576) );
  NAND2_X2 U22491 ( .A1(n384), .A2(n11103), .ZN(n16134) );
  NAND2_X2 U22492 ( .A1(n33577), .A2(n6663), .ZN(n7852) );
  AOI22_X2 U22503 ( .A1(n29284), .A2(n16298), .B1(n20116), .B2(n20118), .ZN(
        n33577) );
  XOR2_X1 U22505 ( .A1(n33578), .A2(n32074), .Z(n30445) );
  XOR2_X1 U22509 ( .A1(n6218), .A2(n20979), .Z(n33578) );
  XOR2_X1 U22513 ( .A1(n24419), .A2(n33579), .Z(n28819) );
  OAI21_X1 U22516 ( .A1(n9251), .A2(n786), .B(n33580), .ZN(n10587) );
  AOI22_X1 U22517 ( .A1(n3988), .A2(n4953), .B1(n4952), .B2(n27149), .ZN(
        n33580) );
  BUF_X2 U22520 ( .I(n946), .Z(n33581) );
  NAND2_X1 U22521 ( .A1(n30384), .A2(n30383), .ZN(n33582) );
  XOR2_X1 U22525 ( .A1(n12721), .A2(n20775), .Z(n20756) );
  NAND2_X2 U22527 ( .A1(n34045), .A2(n20585), .ZN(n12721) );
  XOR2_X1 U22528 ( .A1(n11897), .A2(n23519), .Z(n26338) );
  XOR2_X1 U22532 ( .A1(n12478), .A2(n20784), .Z(n20925) );
  XOR2_X1 U22533 ( .A1(n28968), .A2(n17869), .Z(n17867) );
  XOR2_X1 U22534 ( .A1(n27344), .A2(n33584), .Z(n28496) );
  XOR2_X1 U22535 ( .A1(n24800), .A2(n1227), .Z(n33584) );
  NOR3_X1 U22536 ( .A1(n15134), .A2(n13764), .A3(n31236), .ZN(n15133) );
  OAI22_X1 U22537 ( .A1(n8722), .A2(n25130), .B1(n8723), .B2(n712), .ZN(n27664) );
  XOR2_X1 U22540 ( .A1(n18042), .A2(n24647), .Z(n9868) );
  XOR2_X1 U22548 ( .A1(n6547), .A2(n24573), .Z(n24647) );
  AOI21_X2 U22549 ( .A1(n33615), .A2(n27443), .B(n32020), .ZN(n25317) );
  XOR2_X1 U22561 ( .A1(n11862), .A2(n33587), .Z(n21918) );
  INV_X1 U22564 ( .I(n24861), .ZN(n33587) );
  NAND3_X2 U22565 ( .A1(n9473), .A2(n12156), .A3(n12157), .ZN(n23271) );
  BUF_X2 U22567 ( .I(n12493), .Z(n33588) );
  NOR2_X2 U22570 ( .A1(n6661), .A2(n14092), .ZN(n33589) );
  XOR2_X1 U22582 ( .A1(n23518), .A2(n33590), .Z(n31751) );
  XOR2_X1 U22587 ( .A1(n8068), .A2(n16373), .Z(n23518) );
  XOR2_X1 U22598 ( .A1(n30528), .A2(n16693), .Z(n29772) );
  NOR2_X2 U22605 ( .A1(n28782), .A2(n28783), .ZN(n17460) );
  NAND3_X1 U22606 ( .A1(n22642), .A2(n6297), .A3(n22645), .ZN(n22337) );
  XOR2_X1 U22612 ( .A1(n32404), .A2(n33593), .Z(n31380) );
  NAND2_X2 U22626 ( .A1(n29605), .A2(n5671), .ZN(n12800) );
  AND2_X1 U22635 ( .A1(n10673), .A2(n23706), .Z(n23634) );
  BUF_X2 U22636 ( .I(n5226), .Z(n33597) );
  NAND2_X1 U22643 ( .A1(n26390), .A2(n9127), .ZN(n33599) );
  NAND2_X2 U22648 ( .A1(n10926), .A2(n27879), .ZN(n20471) );
  NAND2_X2 U22649 ( .A1(n695), .A2(n33600), .ZN(n2236) );
  NOR2_X2 U22653 ( .A1(n10251), .A2(n32023), .ZN(n33600) );
  NOR2_X2 U22657 ( .A1(n33602), .A2(n33601), .ZN(n5790) );
  NAND2_X2 U22661 ( .A1(n28351), .A2(n33603), .ZN(n33602) );
  NAND3_X2 U22663 ( .A1(n26667), .A2(n33132), .A3(n18261), .ZN(n1564) );
  NOR2_X1 U22669 ( .A1(n7868), .A2(n11401), .ZN(n21556) );
  NAND2_X2 U22672 ( .A1(n13152), .A2(n13150), .ZN(n11401) );
  NOR2_X1 U22676 ( .A1(n17956), .A2(n21220), .ZN(n10837) );
  XOR2_X1 U22677 ( .A1(n17400), .A2(n32050), .Z(n17766) );
  XOR2_X1 U22679 ( .A1(n31340), .A2(n24624), .Z(n33604) );
  XOR2_X1 U22681 ( .A1(n4790), .A2(n2142), .Z(n7665) );
  XOR2_X1 U22683 ( .A1(n20789), .A2(n20890), .Z(n28405) );
  NAND2_X2 U22685 ( .A1(n21545), .A2(n21544), .ZN(n22157) );
  NOR2_X2 U22686 ( .A1(n18672), .A2(n18881), .ZN(n18517) );
  INV_X2 U22687 ( .I(n18879), .ZN(n18672) );
  XOR2_X1 U22689 ( .A1(n18354), .A2(Key[8]), .Z(n18879) );
  NAND2_X2 U22690 ( .A1(n3137), .A2(n33605), .ZN(n3629) );
  NOR2_X2 U22692 ( .A1(n28269), .A2(n28268), .ZN(n33605) );
  XOR2_X1 U22694 ( .A1(n7705), .A2(n21028), .Z(n21031) );
  XOR2_X1 U22715 ( .A1(n33607), .A2(n10249), .Z(n10303) );
  XOR2_X1 U22716 ( .A1(n7288), .A2(n33747), .Z(n33607) );
  BUF_X2 U22724 ( .I(n29757), .Z(n33608) );
  AOI22_X1 U22726 ( .A1(n1830), .A2(n1832), .B1(n1833), .B2(n7555), .ZN(n33612) );
  NAND2_X2 U22731 ( .A1(n5075), .A2(n5077), .ZN(n8617) );
  XOR2_X1 U22736 ( .A1(n33609), .A2(n23315), .Z(n17797) );
  XOR2_X1 U22740 ( .A1(n29299), .A2(n23332), .Z(n23315) );
  XOR2_X1 U22743 ( .A1(n33612), .A2(n1390), .Z(Ciphertext[58]) );
  XOR2_X1 U22745 ( .A1(n33613), .A2(n33614), .Z(n29916) );
  XOR2_X1 U22747 ( .A1(n11062), .A2(n29955), .Z(n33614) );
  OAI21_X2 U22752 ( .A1(n33761), .A2(n13985), .B(n31060), .ZN(n33615) );
  INV_X2 U22757 ( .I(n33617), .ZN(n18156) );
  XOR2_X1 U22761 ( .A1(n33618), .A2(n20918), .Z(n28998) );
  XOR2_X1 U22763 ( .A1(n29918), .A2(n20652), .Z(n33618) );
  XOR2_X1 U22772 ( .A1(n8973), .A2(n8975), .Z(n27960) );
  NAND2_X1 U22784 ( .A1(n30888), .A2(n3901), .ZN(n33767) );
  NAND2_X2 U22791 ( .A1(n31629), .A2(n33619), .ZN(n2860) );
  AOI22_X2 U22793 ( .A1(n19188), .A2(n33672), .B1(n12316), .B2(n9538), .ZN(
        n31682) );
  NOR2_X2 U22794 ( .A1(n1883), .A2(n14597), .ZN(n19188) );
  OAI21_X2 U22796 ( .A1(n11112), .A2(n11409), .B(n25306), .ZN(n33620) );
  XOR2_X1 U22800 ( .A1(n24173), .A2(n33622), .Z(n24181) );
  XOR2_X1 U22801 ( .A1(n15368), .A2(n6050), .Z(n33622) );
  INV_X2 U22802 ( .I(n28181), .ZN(n15772) );
  OR2_X1 U22803 ( .A1(n28181), .A2(n17416), .Z(n21348) );
  INV_X1 U22805 ( .I(n22271), .ZN(n22218) );
  XOR2_X1 U22806 ( .A1(n22271), .A2(n24759), .Z(n29350) );
  XOR2_X1 U22810 ( .A1(n16073), .A2(n23336), .Z(n23496) );
  NAND2_X2 U22812 ( .A1(n20594), .A2(n20599), .ZN(n10379) );
  INV_X4 U22815 ( .I(n25806), .ZN(n9181) );
  NAND2_X2 U22819 ( .A1(n8759), .A2(n33623), .ZN(n20577) );
  AOI22_X2 U22821 ( .A1(n11587), .A2(n17696), .B1(n16243), .B2(n19971), .ZN(
        n33623) );
  XOR2_X1 U22828 ( .A1(n33905), .A2(n31725), .Z(n28142) );
  OAI21_X2 U22831 ( .A1(n31082), .A2(n30060), .B(n6932), .ZN(n29785) );
  NAND2_X2 U22836 ( .A1(n33626), .A2(n33625), .ZN(n33752) );
  BUF_X2 U22837 ( .I(n34151), .Z(n33627) );
  XOR2_X1 U22838 ( .A1(n24646), .A2(n15508), .Z(n24563) );
  NAND2_X2 U22841 ( .A1(n7884), .A2(n7883), .ZN(n24646) );
  AOI21_X2 U22846 ( .A1(n29849), .A2(n3236), .B(n7377), .ZN(n7620) );
  NOR2_X2 U22851 ( .A1(n5395), .A2(n505), .ZN(n7377) );
  BUF_X2 U22861 ( .I(n10871), .Z(n33628) );
  AOI22_X2 U22862 ( .A1(n24467), .A2(n27128), .B1(n31378), .B2(n1221), .ZN(
        n24947) );
  NOR2_X1 U22863 ( .A1(n29666), .A2(n19885), .ZN(n20058) );
  XOR2_X1 U22868 ( .A1(n392), .A2(n32085), .Z(n21356) );
  XOR2_X1 U22873 ( .A1(n33995), .A2(n28082), .Z(n13817) );
  NOR2_X2 U22874 ( .A1(n6590), .A2(n33629), .ZN(n2971) );
  OAI22_X2 U22876 ( .A1(n34066), .A2(n6587), .B1(n829), .B2(n785), .ZN(n33629)
         );
  AOI21_X2 U22878 ( .A1(n21558), .A2(n38), .B(n33630), .ZN(n22317) );
  OAI22_X2 U22881 ( .A1(n32079), .A2(n21817), .B1(n21820), .B2(n1015), .ZN(
        n33630) );
  XOR2_X1 U22883 ( .A1(n8761), .A2(n27548), .Z(n8765) );
  XOR2_X1 U22887 ( .A1(n20733), .A2(n20843), .Z(n21003) );
  NOR2_X2 U22889 ( .A1(n16858), .A2(n20496), .ZN(n20843) );
  OAI22_X2 U22892 ( .A1(n33631), .A2(n1028), .B1(n7228), .B2(n12917), .ZN(
        n7253) );
  NAND2_X2 U22899 ( .A1(n25845), .A2(n13944), .ZN(n25851) );
  NAND2_X2 U22908 ( .A1(n34044), .A2(n3447), .ZN(n3718) );
  BUF_X2 U22919 ( .I(n1944), .Z(n33633) );
  AOI21_X2 U22932 ( .A1(n6063), .A2(n6064), .B(n33634), .ZN(n22361) );
  INV_X4 U22938 ( .I(n28553), .ZN(n24249) );
  NAND2_X2 U22940 ( .A1(n7357), .A2(n7356), .ZN(n17400) );
  XOR2_X1 U22941 ( .A1(n6545), .A2(n24770), .Z(n2667) );
  NOR2_X2 U22942 ( .A1(n17747), .A2(n6651), .ZN(n6545) );
  XOR2_X1 U22949 ( .A1(n16917), .A2(n13299), .Z(n4291) );
  OAI21_X2 U22951 ( .A1(n3305), .A2(n2045), .B(n30248), .ZN(n16917) );
  XOR2_X1 U22952 ( .A1(n23391), .A2(n9153), .Z(n10289) );
  AND2_X1 U22953 ( .A1(n9578), .A2(n12952), .Z(n15920) );
  XOR2_X1 U22964 ( .A1(n27211), .A2(n24693), .Z(n27851) );
  XOR2_X1 U22971 ( .A1(n24753), .A2(n24853), .Z(n24693) );
  OR2_X1 U22972 ( .A1(n26120), .A2(n23748), .Z(n24074) );
  XOR2_X1 U22974 ( .A1(n7638), .A2(n7639), .Z(n33636) );
  XOR2_X1 U22983 ( .A1(n33637), .A2(n16738), .Z(n31655) );
  XOR2_X1 U22990 ( .A1(n27458), .A2(n7466), .Z(n33637) );
  XOR2_X1 U22994 ( .A1(n33638), .A2(n23314), .Z(n7616) );
  OAI21_X2 U23000 ( .A1(n31768), .A2(n111), .B(n8998), .ZN(n33639) );
  NOR2_X2 U23001 ( .A1(n21858), .A2(n29523), .ZN(n21856) );
  AOI21_X2 U23006 ( .A1(n30067), .A2(n29911), .B(n24099), .ZN(n24927) );
  XOR2_X1 U23008 ( .A1(n33642), .A2(n20711), .Z(n15047) );
  XOR2_X1 U23009 ( .A1(n2356), .A2(n1343), .Z(n33642) );
  AND2_X2 U23011 ( .A1(n4224), .A2(n33856), .Z(n13859) );
  OR2_X1 U23024 ( .A1(n22831), .A2(n4110), .Z(n9473) );
  NOR2_X1 U23025 ( .A1(n34064), .A2(n11215), .ZN(n1557) );
  XOR2_X1 U23037 ( .A1(n11665), .A2(n7705), .Z(n8189) );
  NOR2_X1 U23039 ( .A1(n15039), .A2(n32119), .ZN(n23092) );
  NAND3_X2 U23040 ( .A1(n23964), .A2(n10046), .A3(n18120), .ZN(n33645) );
  NOR2_X2 U23042 ( .A1(n33646), .A2(n15328), .ZN(n15324) );
  XOR2_X1 U23047 ( .A1(n20767), .A2(n20768), .Z(n10707) );
  XOR2_X1 U23054 ( .A1(n21009), .A2(n20715), .Z(n20768) );
  XOR2_X1 U23059 ( .A1(n19599), .A2(n2483), .Z(n19542) );
  NAND2_X1 U23062 ( .A1(n33647), .A2(n21175), .ZN(n13316) );
  NAND2_X1 U23064 ( .A1(n31894), .A2(n985), .ZN(n7221) );
  OR2_X1 U23066 ( .A1(n4327), .A2(n11677), .Z(n25943) );
  NOR2_X1 U23070 ( .A1(n1480), .A2(n1235), .ZN(n33648) );
  OAI21_X2 U23077 ( .A1(n25886), .A2(n4318), .B(n2182), .ZN(n34069) );
  XOR2_X1 U23080 ( .A1(n2592), .A2(n8138), .Z(n26511) );
  XOR2_X1 U23087 ( .A1(n9222), .A2(n23237), .Z(n26889) );
  XOR2_X1 U23093 ( .A1(n8695), .A2(n23430), .Z(n23237) );
  XOR2_X1 U23095 ( .A1(n27850), .A2(n22132), .Z(n22183) );
  XOR2_X1 U23096 ( .A1(n33651), .A2(n23505), .Z(n30964) );
  XOR2_X1 U23108 ( .A1(n31251), .A2(n33652), .Z(n9744) );
  XOR2_X1 U23120 ( .A1(n20711), .A2(n20642), .Z(n33652) );
  OR2_X2 U23121 ( .A1(n2655), .A2(n33536), .Z(n22450) );
  NAND2_X2 U23127 ( .A1(n33654), .A2(n33653), .ZN(n23679) );
  NAND2_X2 U23130 ( .A1(n24198), .A2(n33655), .ZN(n33654) );
  NAND2_X2 U23132 ( .A1(n1241), .A2(n24304), .ZN(n24198) );
  OR2_X1 U23133 ( .A1(n7287), .A2(n14402), .Z(n33657) );
  XOR2_X1 U23134 ( .A1(n19536), .A2(n400), .Z(n30016) );
  XOR2_X1 U23135 ( .A1(n19676), .A2(n19779), .Z(n19536) );
  XOR2_X1 U23144 ( .A1(n19409), .A2(n25598), .Z(n8055) );
  NAND2_X1 U23146 ( .A1(n27531), .A2(n25445), .ZN(n33658) );
  XOR2_X1 U23149 ( .A1(n27055), .A2(n11422), .Z(n8133) );
  NAND2_X2 U23152 ( .A1(n23354), .A2(n31058), .ZN(n24106) );
  NAND2_X2 U23157 ( .A1(n33660), .A2(n29575), .ZN(n17361) );
  NOR2_X2 U23165 ( .A1(n15245), .A2(n30717), .ZN(n33660) );
  NAND2_X2 U23168 ( .A1(n20309), .A2(n33661), .ZN(n30749) );
  AOI22_X2 U23176 ( .A1(n29432), .A2(n31961), .B1(n28626), .B2(n2134), .ZN(
        n33661) );
  XOR2_X1 U23184 ( .A1(n33662), .A2(n23188), .Z(n23025) );
  XOR2_X1 U23185 ( .A1(n9369), .A2(n30550), .Z(n9235) );
  XOR2_X1 U23194 ( .A1(n11481), .A2(n5476), .Z(n9369) );
  XOR2_X1 U23196 ( .A1(n15630), .A2(n17830), .Z(n8464) );
  XOR2_X1 U23198 ( .A1(n30013), .A2(n31477), .Z(n17830) );
  XOR2_X1 U23202 ( .A1(n33663), .A2(n15484), .Z(n17047) );
  NAND2_X2 U23205 ( .A1(n18379), .A2(n12534), .ZN(n29146) );
  OR2_X1 U23206 ( .A1(n25116), .A2(n18156), .Z(n25117) );
  XOR2_X1 U23209 ( .A1(n31568), .A2(n6488), .Z(n33665) );
  NAND2_X2 U23212 ( .A1(n11442), .A2(n31124), .ZN(n30234) );
  XOR2_X1 U23213 ( .A1(n9300), .A2(n13508), .Z(n24624) );
  NAND3_X2 U23215 ( .A1(n34079), .A2(n17943), .A3(n24266), .ZN(n13508) );
  XOR2_X1 U23217 ( .A1(n29652), .A2(n10332), .Z(n20711) );
  OAI22_X2 U23227 ( .A1(n10324), .A2(n11839), .B1(n11840), .B2(n4077), .ZN(
        n29652) );
  AOI22_X2 U23229 ( .A1(n1573), .A2(n24873), .B1(n5662), .B2(n8758), .ZN(
        n33666) );
  AOI21_X2 U23230 ( .A1(n1446), .A2(n8395), .B(n18800), .ZN(n1449) );
  NOR2_X1 U23231 ( .A1(n3790), .A2(n10465), .ZN(n19381) );
  OAI21_X2 U23234 ( .A1(n12322), .A2(n8611), .B(n5347), .ZN(n14179) );
  OAI21_X2 U23258 ( .A1(n15405), .A2(n15404), .B(n8095), .ZN(n33668) );
  NAND3_X2 U23262 ( .A1(n2004), .A2(n2003), .A3(n2005), .ZN(n2396) );
  NAND2_X1 U23282 ( .A1(n2141), .A2(n33669), .ZN(n2398) );
  XOR2_X1 U23283 ( .A1(n23535), .A2(n27708), .Z(n23234) );
  NAND2_X2 U23291 ( .A1(n3513), .A2(n3512), .ZN(n23535) );
  AOI22_X2 U23295 ( .A1(n33671), .A2(n18621), .B1(n18626), .B2(n26550), .ZN(
        n4619) );
  OAI21_X1 U23304 ( .A1(n15660), .A2(n14939), .B(n10470), .ZN(n23973) );
  NOR2_X2 U23306 ( .A1(n30282), .A2(n976), .ZN(n15660) );
  BUF_X2 U23308 ( .I(n9885), .Z(n33672) );
  XOR2_X1 U23309 ( .A1(n19632), .A2(n31415), .Z(n17552) );
  NAND2_X2 U23323 ( .A1(n33775), .A2(n33674), .ZN(n3181) );
  AOI22_X2 U23329 ( .A1(n7407), .A2(n23901), .B1(n7406), .B2(n1254), .ZN(
        n33674) );
  XOR2_X1 U23336 ( .A1(n19503), .A2(n9161), .Z(n9160) );
  XOR2_X1 U23349 ( .A1(n26623), .A2(n31057), .Z(n19503) );
  AOI22_X2 U23358 ( .A1(n18376), .A2(n4626), .B1(n32127), .B2(n18375), .ZN(
        n12534) );
  XOR2_X1 U23362 ( .A1(n33677), .A2(n1392), .Z(Ciphertext[54]) );
  NOR3_X2 U23364 ( .A1(n29227), .A2(n6814), .A3(n27518), .ZN(n33677) );
  XOR2_X1 U23366 ( .A1(n526), .A2(n6571), .Z(n33678) );
  OR3_X1 U23375 ( .A1(n12952), .A2(n22597), .A3(n4378), .Z(n22512) );
  AOI21_X1 U23376 ( .A1(n11113), .A2(n29815), .B(n15291), .ZN(n33719) );
  NOR2_X2 U23377 ( .A1(n7233), .A2(n12051), .ZN(n29815) );
  INV_X2 U23378 ( .I(n2396), .ZN(n33680) );
  NAND2_X2 U23379 ( .A1(n31707), .A2(n1525), .ZN(n24243) );
  NAND2_X2 U23380 ( .A1(n347), .A2(n2577), .ZN(n2576) );
  NAND3_X2 U23383 ( .A1(n4922), .A2(n4920), .A3(n14860), .ZN(n347) );
  NAND2_X2 U23384 ( .A1(n29681), .A2(n30802), .ZN(n2209) );
  NAND2_X2 U23388 ( .A1(n3592), .A2(n3590), .ZN(n30763) );
  INV_X1 U23389 ( .I(n25703), .ZN(n7041) );
  NAND2_X1 U23394 ( .A1(n25703), .A2(n33681), .ZN(n11595) );
  XOR2_X1 U23396 ( .A1(n17653), .A2(n24392), .Z(n25703) );
  XNOR2_X1 U23403 ( .A1(n3028), .A2(n3026), .ZN(n33950) );
  XOR2_X1 U23413 ( .A1(n21007), .A2(n25218), .Z(n15802) );
  NAND2_X2 U23416 ( .A1(n27611), .A2(n4965), .ZN(n21007) );
  XOR2_X1 U23417 ( .A1(n4701), .A2(n34118), .Z(n11364) );
  NAND2_X1 U23422 ( .A1(n4049), .A2(n28281), .ZN(n33689) );
  XOR2_X1 U23446 ( .A1(n33685), .A2(n23289), .Z(n27882) );
  XOR2_X1 U23465 ( .A1(n7011), .A2(n29082), .Z(n33685) );
  XNOR2_X1 U23484 ( .A1(n15801), .A2(n16803), .ZN(n28254) );
  NAND2_X1 U23486 ( .A1(n31561), .A2(n31467), .ZN(n29360) );
  NAND2_X2 U23502 ( .A1(n19290), .A2(n19021), .ZN(n2799) );
  AOI22_X2 U23506 ( .A1(n17394), .A2(n10206), .B1(n1286), .B2(n856), .ZN(
        n33690) );
  NOR2_X2 U23507 ( .A1(n7283), .A2(n26164), .ZN(n7108) );
  BUF_X2 U23511 ( .I(n28471), .Z(n33691) );
  NAND2_X2 U23514 ( .A1(n33692), .A2(n8391), .ZN(n21707) );
  NAND2_X1 U23515 ( .A1(n8468), .A2(n8466), .ZN(n33692) );
  XOR2_X1 U23517 ( .A1(n33698), .A2(n33693), .Z(n479) );
  NAND3_X2 U23520 ( .A1(n15109), .A2(n15111), .A3(n30355), .ZN(n33694) );
  NAND2_X1 U23522 ( .A1(n15441), .A2(n9518), .ZN(n33695) );
  OAI21_X1 U23529 ( .A1(n18537), .A2(n1184), .B(n18539), .ZN(n9420) );
  NOR2_X2 U23532 ( .A1(n14624), .A2(n14198), .ZN(n19359) );
  NAND2_X2 U23548 ( .A1(n33696), .A2(n13172), .ZN(n31290) );
  OAI21_X2 U23551 ( .A1(n29774), .A2(n30022), .B(n32481), .ZN(n33696) );
  OAI22_X2 U23554 ( .A1(n9176), .A2(n18969), .B1(n17593), .B2(n10472), .ZN(
        n33749) );
  XOR2_X1 U23567 ( .A1(n33697), .A2(n14701), .Z(n29642) );
  XOR2_X1 U23568 ( .A1(n30338), .A2(n32065), .Z(n33697) );
  XOR2_X1 U23570 ( .A1(n5051), .A2(n14665), .Z(n24473) );
  NAND2_X2 U23573 ( .A1(n23703), .A2(n23702), .ZN(n14665) );
  NAND3_X2 U23576 ( .A1(n34001), .A2(n21576), .A3(n34000), .ZN(n7545) );
  NAND2_X2 U23577 ( .A1(n33981), .A2(n5170), .ZN(n8753) );
  BUF_X2 U23580 ( .I(n3345), .Z(n33700) );
  NOR2_X2 U23587 ( .A1(n24218), .A2(n16554), .ZN(n14386) );
  NOR2_X2 U23594 ( .A1(n1355), .A2(n3944), .ZN(n30603) );
  NAND2_X2 U23595 ( .A1(n14974), .A2(n23786), .ZN(n23877) );
  NAND2_X1 U23596 ( .A1(n33703), .A2(n14443), .ZN(n23703) );
  NAND2_X1 U23598 ( .A1(n5437), .A2(n26674), .ZN(n33703) );
  NOR2_X2 U23599 ( .A1(n517), .A2(n21743), .ZN(n21778) );
  XOR2_X1 U23600 ( .A1(n33704), .A2(n1801), .Z(n26345) );
  XOR2_X1 U23601 ( .A1(n33984), .A2(n20887), .Z(n33704) );
  INV_X2 U23602 ( .I(n19950), .ZN(n6580) );
  XOR2_X1 U23606 ( .A1(n22324), .A2(n33706), .Z(n9168) );
  XOR2_X1 U23609 ( .A1(n22322), .A2(n33707), .Z(n33706) );
  XNOR2_X1 U23622 ( .A1(n27860), .A2(n721), .ZN(n33895) );
  AOI22_X2 U23629 ( .A1(n27595), .A2(n31954), .B1(n2386), .B2(n14794), .ZN(
        n33708) );
  NOR2_X1 U23636 ( .A1(n33709), .A2(n11902), .ZN(n15277) );
  NOR2_X1 U23639 ( .A1(n29872), .A2(n579), .ZN(n33709) );
  OAI21_X2 U23641 ( .A1(n30477), .A2(n27329), .B(n31959), .ZN(n15521) );
  XOR2_X1 U23646 ( .A1(n33710), .A2(n33711), .Z(n15507) );
  XOR2_X1 U23647 ( .A1(n2838), .A2(n29879), .Z(n27506) );
  AND2_X1 U23653 ( .A1(n9939), .A2(n15722), .Z(n23688) );
  NOR3_X1 U23658 ( .A1(n4286), .A2(n12593), .A3(n9220), .ZN(n29370) );
  INV_X2 U23663 ( .I(n21553), .ZN(n31042) );
  XOR2_X1 U23664 ( .A1(n31523), .A2(n24968), .Z(n33711) );
  AOI21_X2 U23666 ( .A1(n31861), .A2(n33713), .B(n12824), .ZN(n12823) );
  OAI22_X2 U23668 ( .A1(n22873), .A2(n18241), .B1(n27090), .B2(n4113), .ZN(
        n33713) );
  XOR2_X1 U23674 ( .A1(n33796), .A2(n19748), .Z(n29986) );
  XOR2_X1 U23675 ( .A1(n19436), .A2(n19583), .Z(n19748) );
  NAND2_X2 U23684 ( .A1(n29071), .A2(n11519), .ZN(n19040) );
  XOR2_X1 U23687 ( .A1(n15788), .A2(n19497), .Z(n11580) );
  NAND2_X2 U23688 ( .A1(n8645), .A2(n27628), .ZN(n30894) );
  XOR2_X1 U23690 ( .A1(n23173), .A2(n23247), .Z(n23369) );
  NAND2_X2 U23693 ( .A1(n33760), .A2(n13983), .ZN(n22816) );
  XOR2_X1 U23694 ( .A1(n23314), .A2(n26123), .Z(n33715) );
  NAND3_X2 U23696 ( .A1(n14708), .A2(n12114), .A3(n14709), .ZN(n8633) );
  XOR2_X1 U23697 ( .A1(n12750), .A2(n33716), .Z(n29908) );
  XOR2_X1 U23698 ( .A1(n30765), .A2(n32026), .Z(n33716) );
  NAND2_X2 U23705 ( .A1(n17756), .A2(n931), .ZN(n20247) );
  NAND2_X2 U23706 ( .A1(n32504), .A2(n5003), .ZN(n17756) );
  NAND2_X2 U23711 ( .A1(n3114), .A2(n3116), .ZN(n3964) );
  AND2_X1 U23712 ( .A1(n17245), .A2(n23944), .Z(n23322) );
  OAI21_X1 U23726 ( .A1(n10214), .A2(n24906), .B(n33717), .ZN(n9969) );
  NAND2_X1 U23729 ( .A1(n792), .A2(n30289), .ZN(n15175) );
  INV_X2 U23731 ( .I(n31650), .ZN(n23912) );
  NAND2_X1 U23740 ( .A1(n29965), .A2(n31650), .ZN(n31667) );
  XOR2_X1 U23743 ( .A1(n17889), .A2(n22223), .Z(n17891) );
  NAND2_X2 U23746 ( .A1(n4106), .A2(n29517), .ZN(n24262) );
  XOR2_X1 U23747 ( .A1(n23264), .A2(n6169), .Z(n9644) );
  AOI21_X2 U23749 ( .A1(n5261), .A2(n8127), .B(n8126), .ZN(n23264) );
  AOI21_X1 U23754 ( .A1(n19851), .A2(n19987), .B(n20000), .ZN(n34101) );
  XOR2_X1 U23763 ( .A1(n33959), .A2(n5445), .Z(n34134) );
  INV_X2 U23764 ( .I(n13180), .ZN(n33722) );
  NOR2_X2 U23771 ( .A1(n28002), .A2(n30633), .ZN(n23224) );
  XOR2_X1 U23775 ( .A1(n23266), .A2(n23267), .Z(n12538) );
  AOI22_X2 U23779 ( .A1(n22853), .A2(n22888), .B1(n22852), .B2(n22851), .ZN(
        n23266) );
  NAND3_X2 U23780 ( .A1(n15312), .A2(n15313), .A3(n32014), .ZN(n20371) );
  NAND3_X2 U23793 ( .A1(n9186), .A2(n21237), .A3(n780), .ZN(n34015) );
  XOR2_X1 U23794 ( .A1(n13545), .A2(n25567), .Z(n15986) );
  NAND2_X2 U23795 ( .A1(n14957), .A2(n29369), .ZN(n21688) );
  OAI21_X2 U23808 ( .A1(n2793), .A2(n16137), .B(n33723), .ZN(n2502) );
  NAND2_X2 U23809 ( .A1(n16137), .A2(n7090), .ZN(n33723) );
  NOR2_X2 U23813 ( .A1(n25234), .A2(n25235), .ZN(n5611) );
  XOR2_X1 U23815 ( .A1(n23534), .A2(n27860), .Z(n23411) );
  NOR2_X2 U23817 ( .A1(n33793), .A2(n34010), .ZN(n10398) );
  XOR2_X1 U23827 ( .A1(n2192), .A2(n20856), .Z(n12736) );
  XOR2_X1 U23855 ( .A1(n1993), .A2(n2989), .Z(n20856) );
  INV_X2 U23856 ( .I(n25517), .ZN(n1209) );
  NAND2_X2 U23862 ( .A1(n33956), .A2(n26277), .ZN(n25517) );
  OAI21_X2 U23874 ( .A1(n12992), .A2(n9879), .B(n4119), .ZN(n26524) );
  XOR2_X1 U23878 ( .A1(n30069), .A2(n30290), .Z(n29720) );
  XOR2_X1 U23879 ( .A1(n29241), .A2(n20775), .Z(n20723) );
  XOR2_X1 U23883 ( .A1(n33725), .A2(n25507), .Z(Ciphertext[116]) );
  NOR3_X2 U23884 ( .A1(n25504), .A2(n30165), .A3(n33772), .ZN(n33725) );
  XOR2_X1 U23889 ( .A1(n27790), .A2(n33726), .Z(n25228) );
  XOR2_X1 U23893 ( .A1(n24575), .A2(n28807), .Z(n33726) );
  XOR2_X1 U23898 ( .A1(n29912), .A2(n4302), .Z(n25111) );
  AND2_X1 U23901 ( .A1(n21218), .A2(n21220), .Z(n29900) );
  OAI21_X2 U23911 ( .A1(n3643), .A2(n32060), .B(n13796), .ZN(n30174) );
  NAND3_X2 U23912 ( .A1(n31868), .A2(n26488), .A3(n33912), .ZN(n3694) );
  NAND2_X2 U23914 ( .A1(n8905), .A2(n13647), .ZN(n30209) );
  NAND2_X1 U23917 ( .A1(n29690), .A2(n7182), .ZN(n10442) );
  NAND2_X2 U23922 ( .A1(n31960), .A2(n6442), .ZN(n21518) );
  NAND2_X1 U23929 ( .A1(n33729), .A2(n18631), .ZN(n3251) );
  XOR2_X1 U23930 ( .A1(n17622), .A2(Key[124]), .Z(n18631) );
  INV_X1 U23931 ( .I(n17143), .ZN(n33729) );
  OR2_X1 U23941 ( .A1(n33731), .A2(n5795), .Z(n3979) );
  NAND2_X2 U23945 ( .A1(n8442), .A2(n25521), .ZN(n31236) );
  XOR2_X1 U23950 ( .A1(Plaintext[185]), .A2(Key[185]), .Z(n18869) );
  OR2_X1 U23967 ( .A1(n22340), .A2(n16306), .Z(n22024) );
  OAI22_X2 U23969 ( .A1(n14690), .A2(n1246), .B1(n24200), .B2(n24311), .ZN(
        n3345) );
  NAND2_X2 U23970 ( .A1(n31619), .A2(n20780), .ZN(n33774) );
  NOR2_X1 U23974 ( .A1(n31504), .A2(n29763), .ZN(n8650) );
  AOI22_X2 U23975 ( .A1(n21652), .A2(n29234), .B1(n31511), .B2(n17354), .ZN(
        n34096) );
  NAND2_X2 U23980 ( .A1(n261), .A2(n28567), .ZN(n22951) );
  XOR2_X1 U23983 ( .A1(n33733), .A2(n25190), .Z(Ciphertext[67]) );
  NAND3_X2 U23987 ( .A1(n9705), .A2(n9704), .A3(n25189), .ZN(n33733) );
  XOR2_X1 U23991 ( .A1(n7348), .A2(n25252), .Z(n22208) );
  XOR2_X1 U23998 ( .A1(n24761), .A2(n24796), .Z(n24695) );
  INV_X2 U24002 ( .I(n33734), .ZN(n29365) );
  NAND2_X2 U24003 ( .A1(n9856), .A2(n33737), .ZN(n25557) );
  NOR2_X1 U24005 ( .A1(n7236), .A2(n7237), .ZN(n33738) );
  NAND2_X2 U24008 ( .A1(n25387), .A2(n33876), .ZN(n25452) );
  OR2_X2 U24021 ( .A1(n17405), .A2(n31248), .Z(n1699) );
  XNOR2_X1 U24022 ( .A1(n3781), .A2(n22166), .ZN(n2309) );
  NAND2_X2 U24024 ( .A1(n33906), .A2(n4498), .ZN(n9252) );
  INV_X2 U24028 ( .I(n30731), .ZN(n33740) );
  INV_X2 U24038 ( .I(n22978), .ZN(n6433) );
  NAND2_X2 U24039 ( .A1(n17432), .A2(n31777), .ZN(n17431) );
  XNOR2_X1 U24041 ( .A1(n10935), .A2(n5848), .ZN(n22061) );
  AOI22_X2 U24042 ( .A1(n3226), .A2(n33691), .B1(n3227), .B2(n26567), .ZN(
        n3439) );
  INV_X2 U24048 ( .I(n12478), .ZN(n21048) );
  INV_X1 U24059 ( .I(n6611), .ZN(n30404) );
  NAND2_X2 U24060 ( .A1(n28087), .A2(n34153), .ZN(n6611) );
  NAND2_X2 U24062 ( .A1(n27285), .A2(n31965), .ZN(n10546) );
  NAND2_X2 U24066 ( .A1(n19235), .A2(n8119), .ZN(n14054) );
  NAND2_X2 U24068 ( .A1(n3403), .A2(n3402), .ZN(n21045) );
  XOR2_X1 U24070 ( .A1(n19627), .A2(n28601), .Z(n33742) );
  XOR2_X1 U24077 ( .A1(n19642), .A2(n29988), .Z(n9103) );
  BUF_X2 U24079 ( .I(n14083), .Z(n33743) );
  XOR2_X1 U24081 ( .A1(n22149), .A2(n22192), .Z(n10703) );
  NAND3_X2 U24085 ( .A1(n6426), .A2(n21935), .A3(n21936), .ZN(n22192) );
  XOR2_X1 U24096 ( .A1(n28632), .A2(n25878), .Z(n26765) );
  NAND2_X2 U24098 ( .A1(n31889), .A2(n29878), .ZN(n28632) );
  NOR2_X2 U24099 ( .A1(n33744), .A2(n3798), .ZN(n10705) );
  NAND2_X2 U24100 ( .A1(n14153), .A2(n21574), .ZN(n33744) );
  INV_X2 U24101 ( .I(n22810), .ZN(n22715) );
  NOR2_X2 U24104 ( .A1(n9071), .A2(n29717), .ZN(n31309) );
  NAND2_X2 U24108 ( .A1(n18322), .A2(n18321), .ZN(n34082) );
  XOR2_X1 U24110 ( .A1(n17798), .A2(n24849), .Z(n5023) );
  NAND2_X2 U24114 ( .A1(n27589), .A2(n22882), .ZN(n27588) );
  AOI21_X2 U24123 ( .A1(n33746), .A2(n4358), .B(n8007), .ZN(n1544) );
  NAND2_X2 U24131 ( .A1(n936), .A2(n6255), .ZN(n15053) );
  XOR2_X1 U24136 ( .A1(n6852), .A2(n14125), .Z(n33747) );
  XOR2_X1 U24138 ( .A1(n9222), .A2(n7832), .Z(n2969) );
  XOR2_X1 U24144 ( .A1(n12821), .A2(n23253), .Z(n7832) );
  XOR2_X1 U24154 ( .A1(n33751), .A2(n20696), .Z(n21184) );
  XOR2_X1 U24157 ( .A1(n21042), .A2(n20796), .Z(n33751) );
  NOR2_X2 U24162 ( .A1(n31028), .A2(n33752), .ZN(n26157) );
  OAI21_X1 U24164 ( .A1(n33854), .A2(n22388), .B(n33753), .ZN(n22382) );
  NAND2_X2 U24165 ( .A1(n30467), .A2(n33754), .ZN(n12585) );
  AOI22_X1 U24179 ( .A1(n33799), .A2(n18767), .B1(n18768), .B2(n28238), .ZN(
        n33754) );
  NAND3_X2 U24184 ( .A1(n317), .A2(n31149), .A3(n25331), .ZN(n33874) );
  XOR2_X1 U24185 ( .A1(n22029), .A2(n22216), .Z(n22144) );
  AOI21_X2 U24188 ( .A1(n33954), .A2(n33955), .B(n21722), .ZN(n22029) );
  NAND2_X1 U24194 ( .A1(n31114), .A2(n16668), .ZN(n33755) );
  XOR2_X1 U24217 ( .A1(n20832), .A2(n31966), .Z(n33756) );
  AND2_X1 U24219 ( .A1(n8901), .A2(n11820), .Z(n10454) );
  NOR2_X2 U24221 ( .A1(n28227), .A2(n31549), .ZN(n5252) );
  AOI21_X2 U24229 ( .A1(n34043), .A2(n14964), .B(n33757), .ZN(n14960) );
  NOR2_X2 U24234 ( .A1(n29339), .A2(n16491), .ZN(n19932) );
  NAND2_X2 U24239 ( .A1(n33758), .A2(n14896), .ZN(n8790) );
  OAI21_X2 U24247 ( .A1(n34081), .A2(n21439), .B(n29933), .ZN(n33758) );
  XOR2_X1 U24248 ( .A1(n22107), .A2(n31649), .Z(n28014) );
  NAND2_X2 U24260 ( .A1(n23974), .A2(n23973), .ZN(n26750) );
  NAND2_X2 U24269 ( .A1(n33759), .A2(n23131), .ZN(n3077) );
  NAND2_X2 U24270 ( .A1(n9397), .A2(n9396), .ZN(n28099) );
  NAND2_X2 U24271 ( .A1(n33762), .A2(n11871), .ZN(n6610) );
  OAI21_X2 U24272 ( .A1(n17573), .A2(n17574), .B(n11958), .ZN(n33762) );
  BUF_X2 U24273 ( .I(n9919), .Z(n33763) );
  OR2_X1 U24286 ( .A1(n5032), .A2(n5034), .Z(n1768) );
  XOR2_X1 U24297 ( .A1(n23143), .A2(n6461), .Z(n22385) );
  XOR2_X1 U24309 ( .A1(n33764), .A2(n5145), .Z(n17476) );
  XOR2_X1 U24315 ( .A1(n29772), .A2(n24743), .Z(n33764) );
  XOR2_X1 U24318 ( .A1(n33765), .A2(n11784), .Z(n31346) );
  XOR2_X1 U24319 ( .A1(n28574), .A2(n28162), .Z(n33765) );
  XNOR2_X1 U24328 ( .A1(n23429), .A2(n1261), .ZN(n28177) );
  OAI21_X2 U24334 ( .A1(n9384), .A2(n5571), .B(n4231), .ZN(n23429) );
  NAND2_X1 U24352 ( .A1(n1106), .A2(n16280), .ZN(n14016) );
  XOR2_X1 U24353 ( .A1(n20690), .A2(n1394), .Z(n9274) );
  NAND2_X2 U24361 ( .A1(n21974), .A2(n21975), .ZN(n22795) );
  NAND2_X2 U24368 ( .A1(n26961), .A2(n33768), .ZN(n20492) );
  XOR2_X1 U24370 ( .A1(n33770), .A2(n30899), .Z(n30593) );
  INV_X4 U24377 ( .I(n6290), .ZN(n19165) );
  NAND2_X2 U24382 ( .A1(n7285), .A2(n7286), .ZN(n6290) );
  OAI21_X2 U24383 ( .A1(n29240), .A2(n739), .B(n33771), .ZN(n15585) );
  NAND2_X1 U24391 ( .A1(n23888), .A2(n23713), .ZN(n33771) );
  NOR2_X1 U24395 ( .A1(n25510), .A2(n8766), .ZN(n33772) );
  NAND2_X2 U24397 ( .A1(n11180), .A2(n33773), .ZN(n25657) );
  NOR3_X2 U24399 ( .A1(n330), .A2(n783), .A3(n26130), .ZN(n30546) );
  OAI21_X2 U24443 ( .A1(n9137), .A2(n27474), .B(n4340), .ZN(n33775) );
  AOI21_X2 U24447 ( .A1(n20296), .A2(n16218), .B(n33776), .ZN(n20299) );
  NAND2_X2 U24452 ( .A1(n24212), .A2(n3718), .ZN(n13458) );
  NAND2_X2 U24453 ( .A1(n9986), .A2(n27904), .ZN(n20479) );
  XOR2_X1 U24454 ( .A1(n13321), .A2(n23511), .Z(n13930) );
  NAND3_X1 U24458 ( .A1(n28167), .A2(n32066), .A3(n5460), .ZN(n26212) );
  NOR2_X1 U24490 ( .A1(n29539), .A2(n686), .ZN(n30998) );
  NAND2_X2 U24502 ( .A1(n4488), .A2(n28487), .ZN(n5512) );
  NAND2_X2 U24503 ( .A1(n3748), .A2(n1775), .ZN(n24149) );
  XOR2_X1 U24507 ( .A1(n31660), .A2(n4831), .Z(n33778) );
  AOI22_X2 U24513 ( .A1(n29407), .A2(n32499), .B1(n21696), .B2(n21697), .ZN(
        n21698) );
  NAND2_X1 U24518 ( .A1(n13654), .A2(n10845), .ZN(n34143) );
  INV_X2 U24525 ( .I(n17098), .ZN(n33779) );
  NOR2_X2 U24533 ( .A1(n26413), .A2(n5396), .ZN(n17098) );
  XOR2_X1 U24541 ( .A1(n3519), .A2(n23297), .Z(n17859) );
  NAND2_X2 U24542 ( .A1(n22618), .A2(n18056), .ZN(n23297) );
  NAND3_X1 U24547 ( .A1(n5239), .A2(n5395), .A3(n26677), .ZN(n5238) );
  XOR2_X1 U24551 ( .A1(n19557), .A2(n18072), .Z(n1698) );
  XOR2_X1 U24553 ( .A1(n33995), .A2(n8785), .Z(n19557) );
  NAND3_X1 U24565 ( .A1(n24340), .A2(n16552), .A3(n14840), .ZN(n24341) );
  OAI21_X2 U24567 ( .A1(n14314), .A2(n16395), .B(n33780), .ZN(n15144) );
  OAI21_X2 U24568 ( .A1(n15789), .A2(n17623), .B(n13554), .ZN(n33780) );
  OAI21_X2 U24571 ( .A1(n33781), .A2(n29282), .B(n27491), .ZN(n31218) );
  NOR2_X2 U24572 ( .A1(n431), .A2(n28767), .ZN(n33781) );
  XOR2_X1 U24579 ( .A1(n33782), .A2(n11834), .Z(n23899) );
  XOR2_X1 U24581 ( .A1(n23390), .A2(n26888), .Z(n33782) );
  XOR2_X1 U24586 ( .A1(n2415), .A2(n2414), .Z(n8398) );
  AOI21_X2 U24588 ( .A1(n18431), .A2(n13554), .B(n30001), .ZN(n34107) );
  NOR2_X1 U24590 ( .A1(n34101), .A2(n12300), .ZN(n31062) );
  NAND2_X2 U24592 ( .A1(n829), .A2(n33785), .ZN(n33784) );
  NOR2_X2 U24595 ( .A1(n13663), .A2(n11918), .ZN(n33785) );
  BUF_X2 U24613 ( .I(n25979), .Z(n33787) );
  OAI21_X2 U24614 ( .A1(n23828), .A2(n1250), .B(n34164), .ZN(n3482) );
  INV_X2 U24615 ( .I(n29268), .ZN(n33788) );
  INV_X2 U24616 ( .I(n33790), .ZN(n10181) );
  XOR2_X1 U24622 ( .A1(Plaintext[175]), .A2(Key[175]), .Z(n33790) );
  XOR2_X1 U24639 ( .A1(n11218), .A2(n11222), .Z(n11221) );
  OAI21_X2 U24642 ( .A1(n32003), .A2(n33792), .B(n33093), .ZN(n8550) );
  NAND2_X1 U24647 ( .A1(n33795), .A2(n33794), .ZN(n33793) );
  INV_X1 U24654 ( .I(n29815), .ZN(n33794) );
  XOR2_X1 U24662 ( .A1(n33633), .A2(n30435), .Z(n33796) );
  XOR2_X1 U24671 ( .A1(n24674), .A2(n17811), .Z(n5529) );
  INV_X2 U24674 ( .I(n9757), .ZN(n34125) );
  NAND2_X1 U24683 ( .A1(n28020), .A2(n28022), .ZN(n33797) );
  AOI21_X2 U24684 ( .A1(n33798), .A2(n1088), .B(n24126), .ZN(n10539) );
  NAND2_X2 U24689 ( .A1(n24123), .A2(n17100), .ZN(n33798) );
  OAI21_X2 U24693 ( .A1(n29553), .A2(n27600), .B(n20301), .ZN(n13943) );
  NAND3_X2 U24699 ( .A1(n32862), .A2(n974), .A3(n24234), .ZN(n24030) );
  XOR2_X1 U24700 ( .A1(n3416), .A2(n26456), .Z(n19455) );
  INV_X2 U24705 ( .I(n33800), .ZN(n29369) );
  NOR2_X2 U24722 ( .A1(n21087), .A2(n28886), .ZN(n33800) );
  XOR2_X1 U24723 ( .A1(n7931), .A2(n33801), .Z(n28608) );
  XOR2_X1 U24726 ( .A1(n7178), .A2(n23452), .Z(n33801) );
  AND2_X1 U24727 ( .A1(n13318), .A2(n15467), .Z(n29789) );
  INV_X2 U24728 ( .I(n33803), .ZN(n9939) );
  XOR2_X1 U24730 ( .A1(n9432), .A2(n26388), .Z(n17899) );
  XOR2_X1 U24733 ( .A1(n11667), .A2(n17775), .Z(n33806) );
  NAND2_X2 U24745 ( .A1(n2631), .A2(n2632), .ZN(n11667) );
  XOR2_X1 U24752 ( .A1(n33804), .A2(n11780), .Z(n11083) );
  OAI21_X2 U24756 ( .A1(n29355), .A2(n29626), .B(n33805), .ZN(n21981) );
  OAI21_X2 U24767 ( .A1(n29597), .A2(n16240), .B(n29626), .ZN(n33805) );
  AND2_X1 U24781 ( .A1(n5433), .A2(n33561), .Z(n6953) );
  XOR2_X1 U24786 ( .A1(n33806), .A2(n450), .Z(n1454) );
  XOR2_X1 U24788 ( .A1(n10585), .A2(n19518), .Z(n5436) );
  XOR2_X1 U24798 ( .A1(n10294), .A2(n19743), .Z(n10585) );
  NAND2_X2 U24799 ( .A1(n10383), .A2(n10382), .ZN(n24053) );
  XOR2_X1 U24809 ( .A1(n33807), .A2(n24968), .Z(Ciphertext[21]) );
  NAND3_X1 U24811 ( .A1(n17330), .A2(n699), .A3(n3846), .ZN(n33807) );
  NAND2_X2 U24816 ( .A1(n16121), .A2(n1489), .ZN(n23766) );
  INV_X2 U24836 ( .I(n33809), .ZN(n29282) );
  NAND2_X2 U24843 ( .A1(n16154), .A2(n8576), .ZN(n33809) );
  AOI22_X1 U24844 ( .A1(n22832), .A2(n17501), .B1(n22753), .B2(n15421), .ZN(
        n30207) );
  XOR2_X1 U24847 ( .A1(n23206), .A2(n33811), .Z(n16829) );
  XOR2_X1 U24853 ( .A1(n23262), .A2(n9153), .Z(n23206) );
  NAND2_X2 U24855 ( .A1(n24117), .A2(n24226), .ZN(n24224) );
  NAND2_X2 U24858 ( .A1(n18044), .A2(n15206), .ZN(n24117) );
  NAND2_X2 U24863 ( .A1(n7789), .A2(n30924), .ZN(n22075) );
  XOR2_X1 U24865 ( .A1(n20699), .A2(n1828), .Z(n20593) );
  XOR2_X1 U24868 ( .A1(Plaintext[76]), .A2(Key[76]), .Z(n31099) );
  OAI22_X2 U24871 ( .A1(n23903), .A2(n17157), .B1(n14975), .B2(n23786), .ZN(
        n23448) );
  XNOR2_X1 U24873 ( .A1(n22313), .A2(n7664), .ZN(n33816) );
  AOI21_X2 U24876 ( .A1(n20592), .A2(n1347), .B(n30882), .ZN(n33815) );
  NAND2_X1 U24878 ( .A1(n10248), .A2(n686), .ZN(n25624) );
  XOR2_X1 U24879 ( .A1(n21726), .A2(n22145), .Z(n21906) );
  NOR2_X2 U24881 ( .A1(n26690), .A2(n6253), .ZN(n22145) );
  XOR2_X1 U24894 ( .A1(n2104), .A2(n33816), .Z(n30994) );
  NAND2_X1 U24898 ( .A1(n33818), .A2(n33817), .ZN(n26109) );
  INV_X1 U24901 ( .I(n14600), .ZN(n33818) );
  NAND2_X2 U24906 ( .A1(n33819), .A2(n7698), .ZN(n7717) );
  XOR2_X1 U24908 ( .A1(n24473), .A2(n1507), .Z(n10277) );
  AOI22_X2 U24916 ( .A1(n2172), .A2(n30988), .B1(n2088), .B2(n2173), .ZN(
        n33821) );
  BUF_X2 U24923 ( .I(n23417), .Z(n33823) );
  NOR3_X2 U24934 ( .A1(n19992), .A2(n28293), .A3(n17882), .ZN(n7775) );
  XOR2_X1 U24935 ( .A1(n30449), .A2(n27669), .Z(n28109) );
  NAND3_X2 U24954 ( .A1(n19850), .A2(n4663), .A3(n27345), .ZN(n8016) );
  NAND2_X2 U24958 ( .A1(n21134), .A2(n33826), .ZN(n21715) );
  NAND2_X2 U24965 ( .A1(n33829), .A2(n28265), .ZN(n33828) );
  XOR2_X1 U24966 ( .A1(n9670), .A2(n9672), .Z(n11413) );
  NOR2_X1 U24967 ( .A1(n12336), .A2(n14523), .ZN(n33830) );
  OR2_X1 U24968 ( .A1(n30172), .A2(n23770), .Z(n33831) );
  NAND2_X2 U24971 ( .A1(n13934), .A2(n27134), .ZN(n3006) );
  AOI21_X2 U24972 ( .A1(n1120), .A2(n34035), .B(n28170), .ZN(n2253) );
  INV_X2 U24973 ( .I(n29687), .ZN(n21039) );
  XNOR2_X1 U24974 ( .A1(n20766), .A2(n32467), .ZN(n29687) );
  BUF_X2 U24986 ( .I(n8965), .Z(n34035) );
  AOI21_X2 U24987 ( .A1(n6138), .A2(n13788), .B(n15406), .ZN(n13202) );
  OAI21_X2 U24988 ( .A1(n8937), .A2(n30730), .B(n33888), .ZN(n6784) );
  XOR2_X1 U25003 ( .A1(n20993), .A2(n33836), .Z(n13504) );
  XOR2_X1 U25004 ( .A1(n8581), .A2(n29870), .Z(n33836) );
  AOI22_X2 U25008 ( .A1(n13448), .A2(n27941), .B1(n13450), .B2(n13449), .ZN(
        n34119) );
  NAND2_X2 U25018 ( .A1(n18443), .A2(n18881), .ZN(n33837) );
  XOR2_X1 U25029 ( .A1(n24372), .A2(n24829), .Z(n8791) );
  XOR2_X1 U25030 ( .A1(n24830), .A2(n24747), .Z(n24372) );
  NAND2_X1 U25032 ( .A1(n18537), .A2(n16042), .ZN(n18538) );
  XOR2_X1 U25033 ( .A1(n19579), .A2(n33838), .Z(n231) );
  XOR2_X1 U25040 ( .A1(n19658), .A2(n19698), .Z(n19579) );
  XOR2_X1 U25041 ( .A1(n23443), .A2(n32905), .Z(n3635) );
  XOR2_X1 U25043 ( .A1(n33839), .A2(n16355), .Z(Ciphertext[70]) );
  OAI22_X1 U25044 ( .A1(n9675), .A2(n9676), .B1(n11365), .B2(n12060), .ZN(
        n33839) );
  XOR2_X1 U25045 ( .A1(n32604), .A2(n22208), .Z(n33840) );
  XOR2_X1 U25057 ( .A1(n2989), .A2(n20801), .Z(n20987) );
  NAND2_X2 U25058 ( .A1(n3035), .A2(n3036), .ZN(n20801) );
  NAND2_X2 U25061 ( .A1(n9905), .A2(n9906), .ZN(n29937) );
  OAI21_X2 U25062 ( .A1(n2368), .A2(n33842), .B(n33841), .ZN(n21558) );
  AOI21_X2 U25063 ( .A1(n22910), .A2(n6433), .B(n5345), .ZN(n17871) );
  INV_X2 U25065 ( .I(n25571), .ZN(n25577) );
  OAI22_X2 U25066 ( .A1(n6640), .A2(n5929), .B1(n5930), .B2(n6641), .ZN(n25571) );
  XOR2_X1 U25069 ( .A1(n23271), .A2(n5904), .Z(n23458) );
  XOR2_X1 U25070 ( .A1(n17859), .A2(n23495), .Z(n3518) );
  OR2_X1 U25072 ( .A1(n25565), .A2(n25582), .Z(n1473) );
  NOR2_X2 U25073 ( .A1(n33844), .A2(n18907), .ZN(n29801) );
  NOR2_X2 U25080 ( .A1(n11798), .A2(n33845), .ZN(n33844) );
  NOR2_X2 U25087 ( .A1(n19268), .A2(n18974), .ZN(n33846) );
  XOR2_X1 U25091 ( .A1(n33847), .A2(n28896), .Z(n11089) );
  XOR2_X1 U25093 ( .A1(n24561), .A2(n24451), .Z(n33847) );
  XOR2_X1 U25096 ( .A1(n24756), .A2(n13496), .Z(n13163) );
  XOR2_X1 U25097 ( .A1(n3295), .A2(n13060), .Z(n24756) );
  XOR2_X1 U25098 ( .A1(n13724), .A2(n34111), .Z(n13723) );
  AOI21_X2 U25104 ( .A1(n8957), .A2(n34054), .B(n9395), .ZN(n33850) );
  NAND2_X2 U25108 ( .A1(n20010), .A2(n20008), .ZN(n13585) );
  XOR2_X1 U25112 ( .A1(n34024), .A2(n10985), .Z(n5675) );
  XOR2_X1 U25113 ( .A1(n3260), .A2(n19403), .Z(n19504) );
  OAI21_X2 U25115 ( .A1(n18789), .A2(n18790), .B(n18788), .ZN(n19403) );
  NOR2_X2 U25129 ( .A1(n6530), .A2(n20325), .ZN(n20324) );
  NAND2_X2 U25135 ( .A1(n5225), .A2(n32051), .ZN(n33999) );
  NAND2_X2 U25140 ( .A1(n33852), .A2(n30012), .ZN(n19520) );
  NAND2_X2 U25141 ( .A1(n23766), .A2(n28676), .ZN(n28745) );
  XOR2_X1 U25142 ( .A1(n24683), .A2(n24579), .Z(n17505) );
  XOR2_X1 U25151 ( .A1(n2278), .A2(n32871), .Z(n24579) );
  INV_X2 U25154 ( .I(n11576), .ZN(n865) );
  XOR2_X1 U25155 ( .A1(n5500), .A2(n11577), .Z(n11576) );
  NAND2_X2 U25160 ( .A1(n3501), .A2(n33855), .ZN(n13191) );
  INV_X2 U25163 ( .I(n21876), .ZN(n33857) );
  OR2_X1 U25170 ( .A1(n17888), .A2(n33857), .Z(n21590) );
  NAND2_X2 U25176 ( .A1(n30798), .A2(n14262), .ZN(n20892) );
  OAI22_X2 U25192 ( .A1(n29422), .A2(n33858), .B1(n4443), .B2(n4442), .ZN(
        n15715) );
  NOR2_X2 U25196 ( .A1(n330), .A2(n4441), .ZN(n33858) );
  XNOR2_X1 U25198 ( .A1(n10169), .A2(n26030), .ZN(n6604) );
  INV_X2 U25206 ( .I(n29322), .ZN(n21629) );
  XOR2_X1 U25208 ( .A1(n13520), .A2(n27950), .Z(n33860) );
  OAI21_X2 U25214 ( .A1(n33862), .A2(n33861), .B(n29325), .ZN(n3852) );
  AOI21_X2 U25219 ( .A1(n33865), .A2(n22483), .B(n33864), .ZN(n33863) );
  OR2_X1 U25220 ( .A1(n28723), .A2(n11089), .Z(n8711) );
  XOR2_X1 U25224 ( .A1(n16992), .A2(n23229), .Z(n33866) );
  BUF_X2 U25232 ( .I(n29767), .Z(n33868) );
  NAND3_X2 U25235 ( .A1(n23636), .A2(n5227), .A3(n23635), .ZN(n5226) );
  NOR2_X2 U25244 ( .A1(n33869), .A2(n22366), .ZN(n9377) );
  XOR2_X1 U25245 ( .A1(n23496), .A2(n23494), .Z(n3517) );
  NOR2_X2 U25246 ( .A1(n5913), .A2(n31096), .ZN(n33871) );
  XOR2_X1 U25255 ( .A1(n3504), .A2(n7679), .Z(n11217) );
  NAND3_X2 U25257 ( .A1(n7668), .A2(n3216), .A3(n3217), .ZN(n7679) );
  XOR2_X1 U25263 ( .A1(n33873), .A2(n25911), .Z(Ciphertext[189]) );
  NAND2_X2 U25268 ( .A1(n13979), .A2(n33874), .ZN(n30144) );
  XOR2_X1 U25270 ( .A1(n19400), .A2(n19399), .Z(n19546) );
  INV_X2 U25286 ( .I(n33875), .ZN(n20065) );
  NAND3_X2 U25292 ( .A1(n32029), .A2(n14139), .A3(n6551), .ZN(n33876) );
  XOR2_X1 U25296 ( .A1(n20588), .A2(n29850), .Z(n33877) );
  NOR2_X2 U25299 ( .A1(n30144), .A2(n33878), .ZN(n25488) );
  NOR3_X2 U25303 ( .A1(n28866), .A2(n25520), .A3(n25561), .ZN(n33878) );
  NAND3_X1 U25304 ( .A1(n14149), .A2(n25485), .A3(n33879), .ZN(Ciphertext[112]) );
  NAND3_X1 U25306 ( .A1(n25481), .A2(n30117), .A3(n30118), .ZN(n33879) );
  INV_X2 U25313 ( .I(n15212), .ZN(n25446) );
  NAND3_X2 U25314 ( .A1(n6818), .A2(n6817), .A3(n6990), .ZN(n12868) );
  NAND2_X2 U25316 ( .A1(n15529), .A2(n33880), .ZN(n25276) );
  XOR2_X1 U25321 ( .A1(n33881), .A2(n14526), .Z(Ciphertext[89]) );
  AOI22_X1 U25327 ( .A1(n16291), .A2(n11294), .B1(n25286), .B2(n28532), .ZN(
        n33881) );
  XOR2_X1 U25330 ( .A1(n11304), .A2(n20977), .Z(n6615) );
  XOR2_X1 U25335 ( .A1(n13844), .A2(n23368), .Z(n14527) );
  OAI21_X2 U25349 ( .A1(n26732), .A2(n26731), .B(n26710), .ZN(n8078) );
  NAND2_X2 U25355 ( .A1(n33883), .A2(n12527), .ZN(n12617) );
  NAND2_X2 U25359 ( .A1(n30720), .A2(n17580), .ZN(n33883) );
  AOI22_X2 U25362 ( .A1(n2039), .A2(n2040), .B1(n33885), .B2(n33884), .ZN(
        n2037) );
  NOR2_X2 U25368 ( .A1(n879), .A2(n880), .ZN(n33885) );
  XOR2_X1 U25369 ( .A1(n31234), .A2(n7137), .Z(n27012) );
  OR2_X1 U25371 ( .A1(n16987), .A2(n30346), .Z(n21843) );
  NOR2_X1 U25372 ( .A1(n8632), .A2(n31040), .ZN(n30730) );
  OAI21_X2 U25373 ( .A1(n33887), .A2(n10113), .B(n33886), .ZN(n8740) );
  INV_X2 U25376 ( .I(n21149), .ZN(n33889) );
  INV_X2 U25378 ( .I(n33890), .ZN(n17255) );
  XNOR2_X1 U25385 ( .A1(Plaintext[78]), .A2(Key[78]), .ZN(n33890) );
  XOR2_X1 U25386 ( .A1(n24675), .A2(n24487), .Z(n24488) );
  NAND3_X2 U25393 ( .A1(n12319), .A2(n10827), .A3(n12318), .ZN(n24675) );
  NOR2_X1 U25394 ( .A1(n11390), .A2(n18676), .ZN(n2105) );
  INV_X1 U25397 ( .I(n12282), .ZN(n18676) );
  XOR2_X1 U25400 ( .A1(Key[14]), .A2(Plaintext[14]), .Z(n12282) );
  NOR3_X1 U25410 ( .A1(n30935), .A2(n749), .A3(n1204), .ZN(n30165) );
  INV_X2 U25419 ( .I(n4782), .ZN(n4953) );
  XOR2_X1 U25422 ( .A1(n9218), .A2(n33893), .Z(n26236) );
  XOR2_X1 U25424 ( .A1(n21035), .A2(n5009), .Z(n33893) );
  NAND2_X1 U25428 ( .A1(n12900), .A2(n18026), .ZN(n72) );
  AOI21_X1 U25429 ( .A1(n27931), .A2(n26158), .B(n24120), .ZN(n10449) );
  OAI21_X2 U25434 ( .A1(n5952), .A2(n5953), .B(n15213), .ZN(n5951) );
  NAND2_X2 U25440 ( .A1(n33896), .A2(n6931), .ZN(n20534) );
  XOR2_X1 U25445 ( .A1(n16608), .A2(n32053), .Z(n34135) );
  XOR2_X1 U25450 ( .A1(n4321), .A2(n2611), .Z(n16608) );
  XOR2_X1 U25457 ( .A1(n33897), .A2(n15712), .Z(n15711) );
  XOR2_X1 U25463 ( .A1(n15293), .A2(n30565), .Z(n33897) );
  NAND2_X1 U25471 ( .A1(n33898), .A2(n19118), .ZN(n13647) );
  OAI21_X2 U25473 ( .A1(n3856), .A2(n18513), .B(n18512), .ZN(n19118) );
  NOR2_X1 U25474 ( .A1(n19120), .A2(n13646), .ZN(n33898) );
  NOR2_X1 U25480 ( .A1(n27060), .A2(n10603), .ZN(n33913) );
  NAND2_X2 U25481 ( .A1(n1982), .A2(n13151), .ZN(n21636) );
  NAND2_X2 U25483 ( .A1(n34054), .A2(n5575), .ZN(n13151) );
  INV_X1 U25484 ( .I(n16374), .ZN(n20298) );
  NAND2_X1 U25486 ( .A1(n33902), .A2(n16374), .ZN(n29201) );
  NAND2_X2 U25487 ( .A1(n34032), .A2(n17346), .ZN(n16374) );
  INV_X2 U25490 ( .I(n28166), .ZN(n33902) );
  INV_X2 U25493 ( .I(n33903), .ZN(n28263) );
  XOR2_X1 U25496 ( .A1(n16641), .A2(n13357), .Z(n3209) );
  NAND2_X2 U25498 ( .A1(n8502), .A2(n12629), .ZN(n24836) );
  NAND2_X1 U25508 ( .A1(n9058), .A2(n21509), .ZN(n9057) );
  XOR2_X1 U25513 ( .A1(n23246), .A2(n23244), .Z(n30912) );
  XOR2_X1 U25517 ( .A1(n15360), .A2(n13638), .Z(n23244) );
  AOI21_X1 U25519 ( .A1(n6475), .A2(n12563), .B(n13693), .ZN(n1962) );
  XOR2_X1 U25520 ( .A1(n1825), .A2(n23230), .Z(n23370) );
  NOR2_X2 U25543 ( .A1(n26607), .A2(n6150), .ZN(n1825) );
  XOR2_X1 U25555 ( .A1(n17811), .A2(n24439), .Z(n33905) );
  AOI22_X2 U25556 ( .A1(n6016), .A2(n34154), .B1(n4855), .B2(n6961), .ZN(
        n33906) );
  OAI21_X2 U25559 ( .A1(n8235), .A2(n12090), .B(n12602), .ZN(n24171) );
  XOR2_X1 U25563 ( .A1(n17973), .A2(n33910), .Z(n26846) );
  XOR2_X1 U25568 ( .A1(n17722), .A2(n32070), .Z(n33910) );
  BUF_X2 U25575 ( .I(n27182), .Z(n33911) );
  OAI22_X1 U25578 ( .A1(n33913), .A2(n10600), .B1(n10604), .B2(n16653), .ZN(
        Ciphertext[88]) );
  NAND2_X2 U25581 ( .A1(n33915), .A2(n33911), .ZN(n33914) );
  INV_X4 U25583 ( .I(n16650), .ZN(n33915) );
  AOI22_X2 U25589 ( .A1(n3596), .A2(n22691), .B1(n1122), .B2(n30436), .ZN(
        n28489) );
  XOR2_X1 U25594 ( .A1(n5501), .A2(n31576), .Z(n5504) );
  XOR2_X1 U25605 ( .A1(n3117), .A2(n3118), .Z(n33916) );
  NAND2_X2 U25618 ( .A1(n3247), .A2(n31645), .ZN(n27767) );
  XOR2_X1 U25623 ( .A1(n11651), .A2(n3544), .Z(n29538) );
  XOR2_X1 U25629 ( .A1(n16971), .A2(n33917), .Z(n27567) );
  XOR2_X1 U25630 ( .A1(n22243), .A2(n33918), .Z(n33917) );
  INV_X1 U25631 ( .I(n25364), .ZN(n33918) );
  NAND3_X2 U25632 ( .A1(n3310), .A2(n3309), .A3(n1036), .ZN(n1678) );
  NAND2_X1 U25633 ( .A1(n23771), .A2(n15116), .ZN(n23772) );
  NAND2_X2 U25635 ( .A1(n27459), .A2(n1610), .ZN(n23771) );
  XOR2_X1 U25638 ( .A1(n13727), .A2(n33920), .Z(n34111) );
  XOR2_X1 U25641 ( .A1(n31526), .A2(n1993), .Z(n33920) );
  XOR2_X1 U25642 ( .A1(n19378), .A2(n18102), .Z(n4986) );
  NOR2_X2 U25646 ( .A1(n26503), .A2(n18103), .ZN(n19378) );
  NAND2_X2 U25648 ( .A1(n26370), .A2(n7703), .ZN(n22076) );
  INV_X2 U25649 ( .I(n33922), .ZN(n14248) );
  XOR2_X1 U25650 ( .A1(Plaintext[122]), .A2(Key[122]), .Z(n33922) );
  NAND2_X2 U25652 ( .A1(n15303), .A2(n24007), .ZN(n24442) );
  AND2_X1 U25653 ( .A1(n10561), .A2(n18615), .Z(n26442) );
  NAND3_X2 U25655 ( .A1(n24867), .A2(n24667), .A3(n25536), .ZN(n26277) );
  NAND2_X2 U25657 ( .A1(n13693), .A2(n20329), .ZN(n20410) );
  NAND2_X2 U25661 ( .A1(n9413), .A2(n9097), .ZN(n13693) );
  NAND2_X2 U25663 ( .A1(n26012), .A2(n6131), .ZN(n7809) );
  INV_X2 U25665 ( .I(n33928), .ZN(n34163) );
  NAND3_X2 U25666 ( .A1(n17001), .A2(n22555), .A3(n413), .ZN(n33928) );
  XOR2_X1 U25673 ( .A1(n33930), .A2(n2015), .Z(n2013) );
  XOR2_X1 U25676 ( .A1(n24493), .A2(n705), .Z(n33930) );
  NAND4_X2 U25678 ( .A1(n13598), .A2(n33932), .A3(n23094), .A4(n33931), .ZN(
        n17278) );
  XOR2_X1 U25679 ( .A1(n15161), .A2(n24770), .Z(n33933) );
  INV_X2 U25680 ( .I(n33934), .ZN(n25) );
  OR2_X1 U25690 ( .A1(n31911), .A2(n21655), .Z(n29947) );
  XOR2_X1 U25694 ( .A1(n12923), .A2(n12921), .Z(n33939) );
  XOR2_X1 U25700 ( .A1(n22061), .A2(n33940), .Z(n21990) );
  XOR2_X1 U25703 ( .A1(n6771), .A2(n26942), .Z(n33940) );
  NAND2_X2 U25704 ( .A1(n27586), .A2(n25404), .ZN(n1700) );
  OAI21_X2 U25717 ( .A1(n16306), .A2(n22497), .B(n25), .ZN(n9108) );
  NAND2_X2 U25725 ( .A1(n3801), .A2(n6455), .ZN(n7881) );
  AND2_X1 U25726 ( .A1(n17143), .A2(n14248), .Z(n18821) );
  NAND3_X2 U25728 ( .A1(n6597), .A2(n1853), .A3(n18511), .ZN(n19042) );
  AOI21_X2 U25734 ( .A1(n11949), .A2(n20147), .B(n20148), .ZN(n28911) );
  NOR3_X1 U25741 ( .A1(n221), .A2(n25575), .A3(n5942), .ZN(n33942) );
  XOR2_X1 U25759 ( .A1(n33943), .A2(n24543), .Z(n6008) );
  XOR2_X1 U25762 ( .A1(n12313), .A2(n14762), .Z(n24543) );
  XOR2_X1 U25778 ( .A1(n28082), .A2(n19754), .Z(n19476) );
  NAND2_X2 U25781 ( .A1(n11801), .A2(n11800), .ZN(n28082) );
  NOR2_X1 U25783 ( .A1(n2613), .A2(n28344), .ZN(n11880) );
  NAND2_X2 U25788 ( .A1(n3124), .A2(n9801), .ZN(n4908) );
  NAND2_X2 U25789 ( .A1(n12891), .A2(n12894), .ZN(n14214) );
  OR2_X1 U25793 ( .A1(n32888), .A2(n14457), .Z(n19851) );
  XOR2_X1 U25801 ( .A1(n30258), .A2(n31857), .Z(n30257) );
  NAND3_X2 U25802 ( .A1(n15910), .A2(n29093), .A3(n19096), .ZN(n13889) );
  NAND2_X1 U25804 ( .A1(n15964), .A2(n25566), .ZN(n13421) );
  INV_X2 U25805 ( .I(n33945), .ZN(n6482) );
  XOR2_X1 U25809 ( .A1(n28709), .A2(n22078), .Z(n22079) );
  NAND2_X2 U25810 ( .A1(n31263), .A2(n25444), .ZN(n25418) );
  XOR2_X1 U25811 ( .A1(n23521), .A2(n23522), .Z(n23526) );
  AOI21_X2 U25812 ( .A1(n31981), .A2(n14973), .B(n23880), .ZN(n17387) );
  NAND3_X2 U25814 ( .A1(n33948), .A2(n14066), .A3(n33947), .ZN(n16486) );
  NAND2_X2 U25819 ( .A1(n29222), .A2(n30065), .ZN(n33947) );
  BUF_X2 U25825 ( .I(n16440), .Z(n33949) );
  INV_X2 U25829 ( .I(n8335), .ZN(n19154) );
  XNOR2_X1 U25830 ( .A1(n23404), .A2(n13638), .ZN(n23502) );
  NAND2_X2 U25832 ( .A1(n30853), .A2(n27695), .ZN(n23404) );
  NOR2_X2 U25833 ( .A1(n27814), .A2(n22981), .ZN(n22839) );
  XOR2_X1 U25836 ( .A1(n2143), .A2(n33950), .Z(n30125) );
  NAND3_X2 U25837 ( .A1(n24044), .A2(n24043), .A3(n33951), .ZN(n24522) );
  NAND3_X2 U25839 ( .A1(n4510), .A2(n34003), .A3(n13881), .ZN(n13807) );
  NAND2_X2 U25840 ( .A1(n25844), .A2(n25846), .ZN(n16673) );
  NAND2_X2 U25841 ( .A1(n25839), .A2(n25901), .ZN(n25844) );
  XOR2_X1 U25846 ( .A1(n12559), .A2(n20857), .Z(n31295) );
  XOR2_X1 U25848 ( .A1(n34067), .A2(n24751), .Z(n27523) );
  XOR2_X1 U25849 ( .A1(n24531), .A2(n2424), .Z(n24751) );
  AOI22_X2 U25851 ( .A1(n20093), .A2(n15192), .B1(n6027), .B2(n10768), .ZN(
        n4075) );
  NAND2_X1 U25852 ( .A1(n13242), .A2(n25987), .ZN(n27265) );
  XOR2_X1 U25853 ( .A1(n1848), .A2(n30664), .Z(n33952) );
  XOR2_X1 U25854 ( .A1(n30393), .A2(n29033), .Z(n25118) );
  INV_X2 U25856 ( .I(n33953), .ZN(n981) );
  XOR2_X1 U25859 ( .A1(n15731), .A2(n6485), .Z(n33953) );
  NOR2_X1 U25862 ( .A1(n23816), .A2(n6759), .ZN(n23817) );
  NAND2_X2 U25863 ( .A1(n15732), .A2(n16431), .ZN(n23816) );
  XOR2_X1 U25864 ( .A1(n24843), .A2(n14645), .Z(n10869) );
  NOR2_X2 U25865 ( .A1(n7358), .A2(n28029), .ZN(n14645) );
  XOR2_X1 U25867 ( .A1(n8993), .A2(n4251), .Z(n6407) );
  NAND2_X1 U25869 ( .A1(n23938), .A2(n9939), .ZN(n34165) );
  NOR2_X1 U25875 ( .A1(n386), .A2(n11567), .ZN(n10409) );
  INV_X2 U25879 ( .I(n2855), .ZN(n386) );
  XOR2_X1 U25880 ( .A1(n2857), .A2(n28286), .Z(n2855) );
  MUX2_X1 U25884 ( .I0(n24960), .I1(n24955), .S(n24947), .Z(n11428) );
  NAND2_X1 U25888 ( .A1(n33957), .A2(n30523), .ZN(n28952) );
  XOR2_X1 U25889 ( .A1(n33958), .A2(n24953), .Z(Ciphertext[14]) );
  NAND2_X1 U25896 ( .A1(n24667), .A2(n25390), .ZN(n33961) );
  NAND2_X1 U25897 ( .A1(n14763), .A2(n14635), .ZN(n14634) );
  NAND2_X1 U25899 ( .A1(n9227), .A2(n788), .ZN(n14635) );
  NOR2_X1 U25904 ( .A1(n14810), .A2(n28736), .ZN(n6831) );
  NOR2_X2 U25905 ( .A1(n27575), .A2(n34090), .ZN(n7554) );
  AOI22_X2 U25906 ( .A1(n18962), .A2(n16592), .B1(n31819), .B2(n33965), .ZN(
        n19711) );
  XOR2_X1 U25907 ( .A1(n24695), .A2(n24576), .Z(n27362) );
  XOR2_X1 U25908 ( .A1(n22075), .A2(n1433), .Z(n7685) );
  NAND4_X2 U25910 ( .A1(n26720), .A2(n20354), .A3(n26722), .A4(n20353), .ZN(
        n20766) );
  XOR2_X1 U25913 ( .A1(n26236), .A2(n33970), .Z(n5392) );
  XOR2_X1 U25916 ( .A1(n20785), .A2(n449), .Z(n33970) );
  NAND3_X2 U25919 ( .A1(n6865), .A2(n6866), .A3(n9015), .ZN(n9287) );
  NAND3_X2 U25926 ( .A1(n16514), .A2(n11204), .A3(n7625), .ZN(n11205) );
  XOR2_X1 U25928 ( .A1(n23344), .A2(n33973), .Z(n3576) );
  XOR2_X1 U25929 ( .A1(n1263), .A2(n23457), .Z(n33973) );
  OAI21_X1 U25930 ( .A1(n13032), .A2(n10497), .B(n28097), .ZN(n10393) );
  INV_X2 U25931 ( .I(n10392), .ZN(n10497) );
  XOR2_X1 U25932 ( .A1(n27526), .A2(n17159), .Z(n10392) );
  AOI21_X2 U25933 ( .A1(n16752), .A2(n25142), .B(n1547), .ZN(n25051) );
  INV_X2 U25937 ( .I(n14126), .ZN(n31867) );
  NAND3_X2 U25945 ( .A1(n29551), .A2(n22351), .A3(n10611), .ZN(n14126) );
  NAND2_X2 U25947 ( .A1(n8455), .A2(n26796), .ZN(n23499) );
  XOR2_X1 U25950 ( .A1(n22017), .A2(n31616), .Z(n27669) );
  NAND3_X2 U25959 ( .A1(n6145), .A2(n6146), .A3(n27529), .ZN(n22225) );
  XOR2_X1 U25960 ( .A1(n13067), .A2(n16584), .Z(n31590) );
  OAI21_X2 U25962 ( .A1(n29737), .A2(n16195), .B(n21564), .ZN(n13067) );
  NAND3_X2 U25963 ( .A1(n4715), .A2(n4716), .A3(n9646), .ZN(n4760) );
  INV_X2 U25965 ( .I(n33977), .ZN(n30282) );
  XOR2_X1 U25967 ( .A1(n30539), .A2(n5038), .Z(n33977) );
  XOR2_X1 U25968 ( .A1(n1762), .A2(n33978), .Z(n16124) );
  XOR2_X1 U25969 ( .A1(n26996), .A2(n22004), .Z(n33978) );
  XOR2_X1 U25970 ( .A1(n2117), .A2(n30795), .Z(n7562) );
  NAND3_X1 U25971 ( .A1(n785), .A2(n18515), .A3(n18639), .ZN(n29492) );
  NAND2_X2 U25978 ( .A1(n3919), .A2(n26391), .ZN(n4655) );
  XOR2_X1 U25979 ( .A1(n23343), .A2(n11249), .Z(n13375) );
  XOR2_X1 U25980 ( .A1(n34030), .A2(n30398), .Z(n25883) );
  XOR2_X1 U25981 ( .A1(n31288), .A2(n1980), .Z(n16992) );
  AND3_X1 U25988 ( .A1(n9328), .A2(n32890), .A3(n30820), .Z(n29773) );
  XOR2_X1 U25989 ( .A1(n7695), .A2(n29543), .Z(n10420) );
  AOI21_X2 U25990 ( .A1(n9177), .A2(n19146), .B(n33983), .ZN(n9904) );
  NAND2_X2 U25994 ( .A1(n13548), .A2(n15146), .ZN(n18546) );
  OAI22_X1 U25995 ( .A1(n29323), .A2(n11922), .B1(n23755), .B2(n15399), .ZN(
        n16224) );
  XOR2_X1 U25996 ( .A1(n26929), .A2(n20885), .Z(n33984) );
  NOR2_X2 U26000 ( .A1(n8736), .A2(n8734), .ZN(n33986) );
  NOR2_X1 U26004 ( .A1(n21463), .A2(n33810), .ZN(n26051) );
  XOR2_X1 U26007 ( .A1(n2667), .A2(n2666), .Z(n2665) );
  OR3_X1 U26008 ( .A1(n1358), .A2(n16489), .A3(n17495), .Z(n29844) );
  AOI21_X2 U26009 ( .A1(n18691), .A2(n33988), .B(n31987), .ZN(n18694) );
  NAND2_X2 U26011 ( .A1(n33989), .A2(n31971), .ZN(n33988) );
  XOR2_X1 U26014 ( .A1(n33991), .A2(n16604), .Z(Ciphertext[142]) );
  NOR2_X2 U26015 ( .A1(n29678), .A2(n15321), .ZN(n15302) );
  NOR2_X2 U26019 ( .A1(n33993), .A2(n27534), .ZN(n12983) );
  NOR2_X1 U26020 ( .A1(n14677), .A2(n9561), .ZN(n33993) );
  XOR2_X1 U26022 ( .A1(n24639), .A2(n33994), .Z(n11843) );
  XOR2_X1 U26026 ( .A1(n9145), .A2(n24638), .Z(n33994) );
  OAI22_X2 U26028 ( .A1(n7568), .A2(n7008), .B1(n19185), .B2(n29440), .ZN(
        n8785) );
  NOR2_X2 U26029 ( .A1(n8636), .A2(n9068), .ZN(n8480) );
  NOR2_X1 U26031 ( .A1(n34106), .A2(n27343), .ZN(n34105) );
  NAND2_X2 U26032 ( .A1(n2704), .A2(n9304), .ZN(n29757) );
  NOR2_X2 U26035 ( .A1(n9215), .A2(n33998), .ZN(n33997) );
  OAI21_X2 U26038 ( .A1(n7170), .A2(n32019), .B(n7167), .ZN(n28553) );
  XOR2_X1 U26039 ( .A1(n14422), .A2(n8358), .Z(n26934) );
  NOR2_X1 U26040 ( .A1(n3782), .A2(n15255), .ZN(n29362) );
  AOI21_X2 U26041 ( .A1(n7400), .A2(n1291), .B(n34002), .ZN(n3801) );
  NAND3_X1 U26042 ( .A1(n22637), .A2(n29626), .A3(n22636), .ZN(n34003) );
  NOR2_X2 U26045 ( .A1(n34004), .A2(n31022), .ZN(n20819) );
  XOR2_X1 U26049 ( .A1(n22067), .A2(n17555), .Z(n21946) );
  NAND2_X2 U26053 ( .A1(n2299), .A2(n2297), .ZN(n17555) );
  XOR2_X1 U26055 ( .A1(n10841), .A2(n6293), .Z(n28950) );
  XOR2_X1 U26058 ( .A1(n11102), .A2(n25500), .Z(n3131) );
  NAND2_X2 U26061 ( .A1(n3133), .A2(n3132), .ZN(n11102) );
  XOR2_X1 U26063 ( .A1(n16930), .A2(n14842), .Z(n29919) );
  AND2_X1 U26064 ( .A1(n20450), .A2(n20375), .Z(n20201) );
  XOR2_X1 U26065 ( .A1(n322), .A2(n24917), .Z(n16717) );
  NAND2_X2 U26077 ( .A1(n13834), .A2(n17411), .ZN(n23376) );
  XOR2_X1 U26081 ( .A1(n7469), .A2(n7472), .Z(n25185) );
  NAND3_X2 U26086 ( .A1(n16898), .A2(n27814), .A3(n29427), .ZN(n34007) );
  XOR2_X1 U26089 ( .A1(n4169), .A2(n8922), .Z(n8933) );
  XOR2_X1 U26093 ( .A1(n20888), .A2(n15268), .Z(n4741) );
  XOR2_X1 U26100 ( .A1(n20717), .A2(n30430), .Z(n15268) );
  NOR2_X1 U26104 ( .A1(n24347), .A2(n24346), .ZN(n34011) );
  XOR2_X1 U26105 ( .A1(n12494), .A2(n20825), .Z(n21026) );
  INV_X1 U26106 ( .I(n22164), .ZN(n1303) );
  XOR2_X1 U26108 ( .A1(n22164), .A2(n34014), .Z(n5884) );
  NOR2_X2 U26109 ( .A1(n4124), .A2(n22978), .ZN(n34017) );
  BUF_X2 U26111 ( .I(n19002), .Z(n34018) );
  NAND3_X1 U26123 ( .A1(n25729), .A2(n9495), .A3(n29331), .ZN(n34019) );
  AOI21_X2 U26127 ( .A1(n21367), .A2(n21369), .B(n21163), .ZN(n34059) );
  XOR2_X1 U26135 ( .A1(n34020), .A2(n22307), .Z(n2095) );
  XOR2_X1 U26140 ( .A1(n32564), .A2(n4057), .Z(n34020) );
  XOR2_X1 U26141 ( .A1(n29644), .A2(n19627), .Z(n19628) );
  NAND2_X2 U26144 ( .A1(n26987), .A2(n26986), .ZN(n20742) );
  INV_X2 U26145 ( .I(n11206), .ZN(n859) );
  XOR2_X1 U26150 ( .A1(n11206), .A2(n34021), .Z(n22177) );
  INV_X1 U26156 ( .I(n16672), .ZN(n34021) );
  NAND2_X2 U26158 ( .A1(n28431), .A2(n10874), .ZN(n11206) );
  NAND2_X1 U26164 ( .A1(n10470), .A2(n26641), .ZN(n2728) );
  XOR2_X1 U26165 ( .A1(n34022), .A2(n20866), .Z(n21210) );
  XOR2_X1 U26169 ( .A1(n29734), .A2(n6465), .Z(n34022) );
  NOR2_X2 U26173 ( .A1(n11990), .A2(n28186), .ZN(n12900) );
  NAND2_X2 U26178 ( .A1(n18551), .A2(n30192), .ZN(n4436) );
  XOR2_X1 U26179 ( .A1(n27152), .A2(n34023), .Z(n27360) );
  XOR2_X1 U26180 ( .A1(n9585), .A2(n24532), .Z(n34023) );
  XOR2_X1 U26181 ( .A1(n8637), .A2(n8504), .Z(n34024) );
  AOI21_X1 U26184 ( .A1(n32414), .A2(n25999), .B(n18983), .ZN(n5477) );
  XOR2_X1 U26188 ( .A1(n9006), .A2(n479), .Z(n9005) );
  XOR2_X1 U26189 ( .A1(n29709), .A2(n23119), .Z(n22969) );
  OAI21_X2 U26197 ( .A1(n32037), .A2(n32858), .B(n2002), .ZN(n22822) );
  NAND2_X2 U26203 ( .A1(n34025), .A2(n26682), .ZN(n13063) );
  NAND2_X1 U26204 ( .A1(n12439), .A2(n6657), .ZN(n34025) );
  AOI22_X2 U26206 ( .A1(n30769), .A2(n1013), .B1(n32252), .B2(n27635), .ZN(
        n34026) );
  AOI22_X2 U26209 ( .A1(n20278), .A2(n20562), .B1(n20280), .B2(n15213), .ZN(
        n17633) );
  XOR2_X1 U26210 ( .A1(n5253), .A2(n12011), .Z(n5256) );
  NAND2_X2 U26212 ( .A1(n10812), .A2(n9374), .ZN(n11064) );
  OAI21_X2 U26216 ( .A1(n34028), .A2(n34027), .B(n28923), .ZN(n17680) );
  NOR2_X1 U26217 ( .A1(n21604), .A2(n33810), .ZN(n34027) );
  XOR2_X1 U26218 ( .A1(n34029), .A2(n29007), .Z(n5187) );
  XOR2_X1 U26219 ( .A1(n19611), .A2(n5190), .Z(n34029) );
  NAND2_X2 U26223 ( .A1(n27440), .A2(n13621), .ZN(n29321) );
  INV_X2 U26224 ( .I(n34031), .ZN(n29398) );
  AOI21_X2 U26232 ( .A1(n24285), .A2(n794), .B(n24041), .ZN(n13551) );
  NAND2_X2 U26233 ( .A1(n26389), .A2(n1475), .ZN(n7574) );
  XOR2_X1 U26234 ( .A1(n20781), .A2(n20985), .Z(n7452) );
  NAND2_X2 U26237 ( .A1(n20287), .A2(n27478), .ZN(n20985) );
  NOR2_X1 U26239 ( .A1(n6831), .A2(n25129), .ZN(n6830) );
  NOR2_X2 U26242 ( .A1(n10699), .A2(n11499), .ZN(n17822) );
  NAND2_X2 U26245 ( .A1(n34033), .A2(n16827), .ZN(n25542) );
  XOR2_X1 U26246 ( .A1(n7828), .A2(n34034), .Z(n29000) );
  INV_X1 U26257 ( .I(n24843), .ZN(n34034) );
  NAND3_X2 U26260 ( .A1(n13205), .A2(n13204), .A3(n32016), .ZN(n24843) );
  XNOR2_X1 U26263 ( .A1(n7045), .A2(n7046), .ZN(n23344) );
  NOR2_X2 U26264 ( .A1(n3200), .A2(n4609), .ZN(n7046) );
  NAND3_X1 U26266 ( .A1(n767), .A2(n24340), .A3(n24163), .ZN(n11331) );
  OAI21_X2 U26270 ( .A1(n20283), .A2(n20282), .B(n20281), .ZN(n20781) );
  XOR2_X1 U26271 ( .A1(n34038), .A2(n21048), .Z(n14340) );
  INV_X2 U26273 ( .I(n9852), .ZN(n19996) );
  OAI22_X2 U26280 ( .A1(n13816), .A2(n21840), .B1(n16386), .B2(n30346), .ZN(
        n21748) );
  NAND2_X2 U26282 ( .A1(n21497), .A2(n21499), .ZN(n21840) );
  XOR2_X1 U26286 ( .A1(n15791), .A2(n14110), .Z(n34085) );
  NOR3_X1 U26290 ( .A1(n7935), .A2(n10513), .A3(n30651), .ZN(n16408) );
  NAND2_X2 U26296 ( .A1(n11033), .A2(n11031), .ZN(n30584) );
  XOR2_X1 U26298 ( .A1(n10585), .A2(n32047), .Z(n27717) );
  NAND2_X2 U26299 ( .A1(n13199), .A2(n15677), .ZN(n22055) );
  INV_X2 U26301 ( .I(n3581), .ZN(n6882) );
  NAND2_X1 U26307 ( .A1(n34039), .A2(n3581), .ZN(n31127) );
  XOR2_X1 U26308 ( .A1(n29260), .A2(n3584), .Z(n3581) );
  NAND3_X2 U26309 ( .A1(n21882), .A2(n21883), .A3(n12019), .ZN(n22737) );
  NAND2_X2 U26310 ( .A1(n9646), .A2(n19325), .ZN(n13913) );
  XOR2_X1 U26311 ( .A1(n34041), .A2(n30881), .Z(Ciphertext[20]) );
  AOI22_X1 U26315 ( .A1(n12203), .A2(n1208), .B1(n12201), .B2(n12202), .ZN(
        n34041) );
  XOR2_X1 U26316 ( .A1(n6020), .A2(n34042), .Z(n11986) );
  XOR2_X1 U26317 ( .A1(n6018), .A2(n31253), .Z(n34042) );
  XOR2_X1 U26322 ( .A1(n5067), .A2(n5068), .Z(n5070) );
  NAND2_X2 U26323 ( .A1(n1773), .A2(n15260), .ZN(n9411) );
  NOR2_X2 U26325 ( .A1(n3446), .A2(n3445), .ZN(n34044) );
  AOI21_X1 U26327 ( .A1(n3650), .A2(n33345), .B(n33216), .ZN(n3667) );
  XOR2_X1 U26331 ( .A1(n14742), .A2(n19722), .Z(n10024) );
  XOR2_X1 U26332 ( .A1(n5127), .A2(n1368), .Z(n14742) );
  NAND2_X1 U26333 ( .A1(n4908), .A2(n5696), .ZN(n22913) );
  XOR2_X1 U26336 ( .A1(Plaintext[157]), .A2(Key[157]), .Z(n16614) );
  INV_X2 U26342 ( .I(n10354), .ZN(n34048) );
  NAND2_X2 U26348 ( .A1(n639), .A2(n34048), .ZN(n29395) );
  NAND3_X2 U26353 ( .A1(n34049), .A2(n26176), .A3(n18341), .ZN(n10423) );
  NAND2_X2 U26360 ( .A1(n18185), .A2(n16426), .ZN(n34049) );
  XOR2_X1 U26361 ( .A1(n29589), .A2(n6545), .Z(n30807) );
  XOR2_X1 U26363 ( .A1(n31491), .A2(n12310), .Z(n30733) );
  NAND2_X2 U26364 ( .A1(n6110), .A2(n4100), .ZN(n34053) );
  XOR2_X1 U26367 ( .A1(n20727), .A2(n32162), .Z(n10164) );
  XOR2_X1 U26369 ( .A1(n6388), .A2(n6572), .Z(n13361) );
  NAND2_X2 U26370 ( .A1(n30846), .A2(n6619), .ZN(n6771) );
  NAND2_X2 U26371 ( .A1(n34055), .A2(n14561), .ZN(n16222) );
  NAND3_X2 U26372 ( .A1(n7205), .A2(n14560), .A3(n7830), .ZN(n34055) );
  BUF_X2 U26376 ( .I(n11193), .Z(n34056) );
  BUF_X2 U26379 ( .I(n16293), .Z(n34057) );
  NOR2_X2 U26383 ( .A1(n26387), .A2(n4151), .ZN(n11049) );
  NOR2_X2 U26386 ( .A1(n847), .A2(n23721), .ZN(n28306) );
  INV_X2 U26387 ( .I(n13361), .ZN(n847) );
  NOR2_X2 U26393 ( .A1(n23929), .A2(n23928), .ZN(n4897) );
  NOR3_X2 U26396 ( .A1(n4197), .A2(n11812), .A3(n847), .ZN(n23929) );
  NAND2_X2 U26397 ( .A1(n1601), .A2(n1600), .ZN(n27189) );
  NOR2_X2 U26398 ( .A1(n31245), .A2(n4531), .ZN(n1601) );
  XOR2_X1 U26402 ( .A1(n30273), .A2(n30487), .Z(n30486) );
  XOR2_X1 U26407 ( .A1(n16829), .A2(n34060), .Z(n23925) );
  XOR2_X1 U26408 ( .A1(n14733), .A2(n29194), .Z(n34060) );
  XOR2_X1 U26409 ( .A1(n22240), .A2(n22210), .Z(n21985) );
  XOR2_X1 U26410 ( .A1(n23261), .A2(n551), .Z(n5737) );
  XOR2_X1 U26422 ( .A1(n24579), .A2(n34061), .Z(n31132) );
  XOR2_X1 U26427 ( .A1(n11370), .A2(n7574), .Z(n34061) );
  NOR2_X1 U26429 ( .A1(n3646), .A2(n5466), .ZN(n25251) );
  XOR2_X1 U26432 ( .A1(n19552), .A2(n31908), .Z(n34062) );
  NAND2_X2 U26433 ( .A1(n5995), .A2(n5996), .ZN(n5994) );
  XOR2_X1 U26436 ( .A1(n34063), .A2(n22141), .Z(n30449) );
  NAND2_X1 U26437 ( .A1(n16034), .A2(n1017), .ZN(n34064) );
  NAND2_X2 U26439 ( .A1(n34065), .A2(n10829), .ZN(n16801) );
  NOR2_X2 U26445 ( .A1(n16393), .A2(n18515), .ZN(n34066) );
  XOR2_X1 U26448 ( .A1(n23143), .A2(n23273), .Z(n4554) );
  XOR2_X1 U26453 ( .A1(n20674), .A2(n20841), .Z(n17738) );
  XOR2_X1 U26455 ( .A1(n21037), .A2(n20892), .Z(n20841) );
  XOR2_X1 U26463 ( .A1(n4567), .A2(n4566), .Z(n34067) );
  NAND2_X2 U26465 ( .A1(n22382), .A2(n17357), .ZN(n15421) );
  INV_X4 U26474 ( .I(n8087), .ZN(n13920) );
  NAND2_X2 U26476 ( .A1(n34068), .A2(n26336), .ZN(n23536) );
  NAND2_X1 U26477 ( .A1(n2031), .A2(n2032), .ZN(n34068) );
  OAI21_X2 U26478 ( .A1(n18821), .A2(n12976), .B(n16352), .ZN(n12975) );
  XOR2_X1 U26481 ( .A1(n34070), .A2(n16530), .Z(Ciphertext[166]) );
  XOR2_X1 U26482 ( .A1(n11726), .A2(n19754), .Z(n34071) );
  OR2_X1 U26485 ( .A1(n16855), .A2(n6634), .Z(n6659) );
  NOR2_X1 U26487 ( .A1(n31783), .A2(n11985), .ZN(n7655) );
  INV_X2 U26488 ( .I(n11548), .ZN(n31783) );
  XOR2_X1 U26489 ( .A1(n24754), .A2(n34072), .Z(n24536) );
  XOR2_X1 U26501 ( .A1(n242), .A2(n27750), .Z(n34072) );
  XOR2_X1 U26507 ( .A1(n34073), .A2(n24369), .Z(n9125) );
  INV_X2 U26510 ( .I(n981), .ZN(n15732) );
  XOR2_X1 U26511 ( .A1(n19391), .A2(n34076), .Z(n29653) );
  XOR2_X1 U26518 ( .A1(n207), .A2(n34077), .Z(n34076) );
  INV_X2 U26519 ( .I(n19769), .ZN(n34077) );
  XOR2_X1 U26520 ( .A1(n26351), .A2(n22145), .Z(n22202) );
  NAND3_X2 U26523 ( .A1(n17941), .A2(n17940), .A3(n5913), .ZN(n34079) );
  XOR2_X1 U26524 ( .A1(n18028), .A2(n12797), .Z(n4332) );
  AOI21_X2 U26525 ( .A1(n18268), .A2(n19147), .B(n18267), .ZN(n19368) );
  XOR2_X1 U26527 ( .A1(n5737), .A2(n29807), .Z(n26170) );
  NAND2_X2 U26528 ( .A1(n26326), .A2(n2239), .ZN(n21497) );
  XOR2_X1 U26531 ( .A1(n9327), .A2(n29540), .Z(n5563) );
  XOR2_X1 U26532 ( .A1(n34085), .A2(n27851), .Z(n15235) );
  OR2_X1 U26533 ( .A1(n21862), .A2(n13652), .Z(n13653) );
  NAND2_X2 U26536 ( .A1(n21738), .A2(n21866), .ZN(n21862) );
  AOI21_X2 U26537 ( .A1(n21361), .A2(n15728), .B(n4906), .ZN(n29302) );
  XOR2_X1 U26538 ( .A1(n34086), .A2(n24435), .Z(Ciphertext[159]) );
  NOR2_X1 U26539 ( .A1(n24433), .A2(n24434), .ZN(n34086) );
  INV_X2 U26540 ( .I(n2132), .ZN(n13966) );
  NAND2_X1 U26541 ( .A1(n34162), .A2(n13862), .ZN(n2132) );
  XOR2_X1 U26542 ( .A1(n17040), .A2(n23121), .Z(n3081) );
  XOR2_X1 U26549 ( .A1(n23306), .A2(n23420), .Z(n23121) );
  OAI21_X2 U26551 ( .A1(n14767), .A2(n14768), .B(n8325), .ZN(n20961) );
  INV_X2 U26555 ( .I(n17426), .ZN(n24212) );
  OAI22_X2 U26556 ( .A1(n14746), .A2(n23651), .B1(n8330), .B2(n23650), .ZN(
        n17426) );
  BUF_X2 U26557 ( .I(n14236), .Z(n34087) );
  XOR2_X1 U26560 ( .A1(n11867), .A2(n27144), .Z(n19684) );
  XOR2_X1 U26563 ( .A1(n335), .A2(n14685), .Z(n22638) );
  XOR2_X1 U26565 ( .A1(n6607), .A2(n6608), .Z(n10675) );
  NOR2_X2 U26566 ( .A1(n29359), .A2(n5825), .ZN(n7776) );
  XOR2_X1 U26569 ( .A1(n11297), .A2(n25001), .Z(n34088) );
  NAND2_X2 U26570 ( .A1(n8418), .A2(n13231), .ZN(n23367) );
  NOR2_X2 U26574 ( .A1(n25968), .A2(n8787), .ZN(n13806) );
  NOR2_X2 U26577 ( .A1(n26432), .A2(n12247), .ZN(n34090) );
  XOR2_X1 U26578 ( .A1(n24854), .A2(n27423), .Z(n26435) );
  XOR2_X1 U26581 ( .A1(n24377), .A2(n34091), .Z(n10901) );
  XOR2_X1 U26582 ( .A1(n24559), .A2(n27750), .Z(n34091) );
  NAND2_X2 U26584 ( .A1(n28699), .A2(n34092), .ZN(n7811) );
  AOI22_X2 U26585 ( .A1(n1889), .A2(n17341), .B1(n5039), .B2(n18218), .ZN(
        n34092) );
  OR2_X1 U26589 ( .A1(n16042), .A2(n14156), .Z(n3344) );
  AOI21_X2 U26593 ( .A1(n2324), .A2(n26976), .B(n34093), .ZN(n16693) );
  BUF_X2 U26595 ( .I(n25665), .Z(n34094) );
  XOR2_X1 U26596 ( .A1(n23465), .A2(n34095), .Z(n4312) );
  XOR2_X1 U26597 ( .A1(n23488), .A2(n16548), .Z(n34095) );
  NAND2_X2 U26598 ( .A1(n3489), .A2(n2536), .ZN(n5410) );
  AND2_X1 U26600 ( .A1(n13525), .A2(n4916), .Z(n29736) );
  OR2_X1 U26601 ( .A1(n6286), .A2(n8178), .Z(n2245) );
  AOI22_X2 U26602 ( .A1(n5387), .A2(n25893), .B1(n16113), .B2(n28910), .ZN(
        n29521) );
  NAND2_X2 U26604 ( .A1(n19866), .A2(n17177), .ZN(n20692) );
  OAI21_X2 U26605 ( .A1(n3656), .A2(n32499), .B(n34102), .ZN(n10824) );
  NOR2_X2 U26606 ( .A1(n26913), .A2(n27836), .ZN(n34102) );
  NOR2_X2 U26609 ( .A1(n18510), .A2(n34110), .ZN(n15789) );
  INV_X2 U26610 ( .I(n18820), .ZN(n34110) );
  XOR2_X1 U26611 ( .A1(n18393), .A2(Key[120]), .Z(n18820) );
  XOR2_X1 U26614 ( .A1(n19764), .A2(n18453), .Z(n19620) );
  NAND2_X2 U26615 ( .A1(n17997), .A2(n17996), .ZN(n18453) );
  XNOR2_X1 U26618 ( .A1(n15419), .A2(n6867), .ZN(n12008) );
  XOR2_X1 U26629 ( .A1(n27349), .A2(n23274), .Z(n34112) );
  NAND3_X1 U26630 ( .A1(n27336), .A2(n26445), .A3(n31458), .ZN(n21564) );
  NAND2_X2 U26633 ( .A1(n1687), .A2(n1688), .ZN(n27336) );
  NAND2_X2 U26634 ( .A1(n34114), .A2(n15069), .ZN(n16209) );
  OR2_X1 U26635 ( .A1(n15071), .A2(n34139), .Z(n34114) );
  XOR2_X1 U26641 ( .A1(n8741), .A2(n19484), .Z(n19518) );
  OAI21_X2 U26643 ( .A1(n18459), .A2(n6597), .B(n956), .ZN(n11519) );
  OR3_X1 U26650 ( .A1(n25236), .A2(n8219), .A3(n34115), .Z(n16398) );
  XOR2_X1 U26651 ( .A1(n24489), .A2(n10474), .Z(n10473) );
  AOI21_X2 U26652 ( .A1(n2743), .A2(n12448), .B(n34116), .ZN(n21992) );
  XOR2_X1 U26656 ( .A1(n34117), .A2(n25815), .Z(Ciphertext[171]) );
  NAND2_X1 U26663 ( .A1(n25813), .A2(n25814), .ZN(n34117) );
  XOR2_X1 U26668 ( .A1(n11349), .A2(n7717), .Z(n2592) );
  XOR2_X1 U26670 ( .A1(n24407), .A2(n30986), .Z(n24408) );
  BUF_X2 U26671 ( .I(n16073), .Z(n34120) );
  INV_X2 U26672 ( .I(n34122), .ZN(n12895) );
  XOR2_X1 U26674 ( .A1(n9914), .A2(n3683), .Z(n6948) );
  OR2_X1 U26675 ( .A1(n7345), .A2(n19057), .Z(n16832) );
  INV_X2 U26676 ( .I(n34123), .ZN(n34169) );
  XOR2_X1 U26678 ( .A1(n8896), .A2(n8894), .Z(n34123) );
  XOR2_X1 U26679 ( .A1(n34124), .A2(n23411), .Z(n7711) );
  XOR2_X1 U26685 ( .A1(n23412), .A2(n32893), .Z(n34124) );
  NAND2_X1 U26687 ( .A1(n34125), .A2(n31692), .ZN(n9271) );
  XOR2_X1 U26693 ( .A1(n10184), .A2(n31100), .Z(n31692) );
  XOR2_X1 U26696 ( .A1(n17323), .A2(n15044), .Z(n34126) );
  OAI21_X2 U26697 ( .A1(n27520), .A2(n5089), .B(n24655), .ZN(n30323) );
  NOR2_X2 U26698 ( .A1(n12511), .A2(n15852), .ZN(n34127) );
  XOR2_X1 U26699 ( .A1(n236), .A2(n34129), .Z(n2312) );
  XOR2_X1 U26700 ( .A1(n23408), .A2(n32027), .Z(n34129) );
  OR2_X1 U26701 ( .A1(n29139), .A2(n27485), .Z(n23793) );
  NAND2_X2 U26702 ( .A1(n2687), .A2(n34130), .ZN(n11266) );
  XOR2_X1 U26703 ( .A1(n34133), .A2(n17793), .Z(n7987) );
  XOR2_X1 U26704 ( .A1(n32111), .A2(n16708), .Z(n34133) );
  XOR2_X1 U26705 ( .A1(n26214), .A2(n6395), .Z(n27933) );
  NOR2_X1 U26706 ( .A1(n8678), .A2(n32874), .ZN(n25789) );
  NOR2_X2 U26707 ( .A1(n15709), .A2(n15276), .ZN(n8678) );
  INV_X2 U26708 ( .I(n34134), .ZN(n13147) );
  INV_X2 U26709 ( .I(n6549), .ZN(n16811) );
  XOR2_X1 U26710 ( .A1(n34135), .A2(n8532), .Z(n6549) );
  OAI21_X2 U26711 ( .A1(n31461), .A2(n24195), .B(n34136), .ZN(n1857) );
  AOI22_X2 U26712 ( .A1(n1315), .A2(n11981), .B1(n4331), .B2(n21700), .ZN(
        n34138) );
  INV_X1 U26713 ( .I(n18295), .ZN(n30934) );
  XOR2_X1 U26714 ( .A1(Plaintext[84]), .A2(Key[84]), .Z(n18295) );
  INV_X2 U26715 ( .I(n15194), .ZN(n34139) );
  XOR2_X1 U26716 ( .A1(n20928), .A2(n15877), .Z(n20753) );
  AOI21_X2 U26717 ( .A1(n20557), .A2(n20556), .B(n15749), .ZN(n20928) );
  AOI22_X2 U26718 ( .A1(n21624), .A2(n17748), .B1(n21623), .B2(n28387), .ZN(
        n7477) );
  BUF_X2 U26719 ( .I(n12074), .Z(n34140) );
  BUF_X2 U26720 ( .I(n18801), .Z(n34141) );
  AOI22_X2 U26721 ( .A1(n34142), .A2(n28056), .B1(n18739), .B2(n16287), .ZN(
        n8203) );
  NOR2_X1 U26722 ( .A1(n18587), .A2(n18737), .ZN(n34142) );
  XOR2_X1 U26723 ( .A1(n23419), .A2(n27186), .Z(n23422) );
  NAND2_X2 U26724 ( .A1(n4776), .A2(n4778), .ZN(n27186) );
  XOR2_X1 U26725 ( .A1(n19556), .A2(n4992), .Z(n5607) );
  OAI21_X2 U26726 ( .A1(n13656), .A2(n13655), .B(n34143), .ZN(n10806) );
  NAND2_X2 U26727 ( .A1(n9508), .A2(n9512), .ZN(n4405) );
  XOR2_X1 U26728 ( .A1(n15028), .A2(n9434), .Z(n9586) );
  NAND2_X2 U26729 ( .A1(n8829), .A2(n8828), .ZN(n9434) );
  XOR2_X1 U26730 ( .A1(n10111), .A2(n12414), .Z(n29140) );
  NAND2_X2 U26731 ( .A1(n4520), .A2(n4519), .ZN(n10111) );
  INV_X2 U26732 ( .I(n34144), .ZN(n9663) );
  XOR2_X1 U26733 ( .A1(n10437), .A2(n10436), .Z(n34144) );
  XOR2_X1 U26734 ( .A1(n34145), .A2(n24619), .Z(n8845) );
  XOR2_X1 U26735 ( .A1(n24747), .A2(n31866), .Z(n34145) );
  NAND2_X1 U26736 ( .A1(n28414), .A2(n31533), .ZN(n31112) );
  AND2_X1 U26737 ( .A1(n651), .A2(n16333), .Z(n10619) );
  NAND3_X2 U26738 ( .A1(n8003), .A2(n8005), .A3(n24030), .ZN(n10084) );
  XOR2_X1 U26739 ( .A1(n1884), .A2(n31626), .Z(n8059) );
  OAI22_X2 U26740 ( .A1(n8653), .A2(n31260), .B1(n8651), .B2(n16157), .ZN(
        n29693) );
  XOR2_X1 U26741 ( .A1(n19543), .A2(n19542), .Z(n34146) );
  XOR2_X1 U26742 ( .A1(n21903), .A2(n21911), .Z(n14506) );
  XOR2_X1 U26743 ( .A1(n1305), .A2(n22291), .Z(n21911) );
  XOR2_X1 U26744 ( .A1(n9907), .A2(n24636), .Z(n24521) );
  OAI21_X2 U26745 ( .A1(n18179), .A2(n34147), .B(n11461), .ZN(n24826) );
  OAI22_X2 U26746 ( .A1(n24183), .A2(n28691), .B1(n10381), .B2(n24052), .ZN(
        n34147) );
  OR2_X1 U26747 ( .A1(n14080), .A2(n10217), .Z(n28507) );
  BUF_X2 U26748 ( .I(n25889), .Z(n34149) );
  XOR2_X1 U26749 ( .A1(n22222), .A2(n8324), .Z(n17889) );
  XOR2_X1 U26750 ( .A1(n26931), .A2(n22147), .Z(n22222) );
  XNOR2_X1 U26751 ( .A1(n3511), .A2(n27599), .ZN(n34151) );
  INV_X2 U26752 ( .I(n14456), .ZN(n31017) );
  NOR2_X1 U26753 ( .A1(n29213), .A2(n5837), .ZN(n34152) );
  INV_X2 U26754 ( .I(n27110), .ZN(n20037) );
  INV_X2 U26755 ( .I(n12670), .ZN(n17767) );
  INV_X4 U26756 ( .I(n8530), .ZN(n21865) );
  NAND2_X2 U26757 ( .A1(n8490), .A2(n31965), .ZN(n21506) );
  INV_X2 U26758 ( .I(n4274), .ZN(n8539) );
  AND2_X2 U26759 ( .A1(n30984), .A2(n31026), .Z(n34160) );
  INV_X2 U26760 ( .I(n11805), .ZN(n22397) );
  XOR2_X1 U26761 ( .A1(n14753), .A2(n11327), .Z(n34161) );
  XNOR2_X1 U26762 ( .A1(n6055), .A2(n28872), .ZN(n34162) );
  BUF_X2 U26763 ( .I(n22598), .Z(n16432) );
  INV_X2 U26764 ( .I(n8365), .ZN(n10295) );
  INV_X2 U26765 ( .I(n6093), .ZN(n28825) );
  NOR2_X2 U26766 ( .A1(n9041), .A2(n9042), .ZN(n30321) );
  INV_X2 U26767 ( .I(n17932), .ZN(n23786) );
  AND2_X1 U26768 ( .A1(n32309), .A2(n23894), .Z(n34166) );
  AND3_X1 U26769 ( .A1(n8694), .A2(n14078), .A3(n6474), .Z(n34168) );
  INV_X4 U26770 ( .I(n2967), .ZN(n11899) );
  AND2_X1 U26771 ( .A1(n24958), .A2(n24939), .Z(n34170) );
endmodule


module SPEEDY_Top ( clk, Plaintext, Key, Ciphertext );
  input [191:0] Plaintext;
  input [191:0] Key;
  output [191:0] Ciphertext;
  input clk;

  wire   [191:0] reg_in;
  wire   [191:0] reg_key;
  wire   [191:0] reg_out;

  DFFSNQ_X1 \reg_in_reg[191]  ( .D(Plaintext[191]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[191]) );
  DFFSNQ_X1 \reg_in_reg[190]  ( .D(Plaintext[190]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[190]) );
  DFFSNQ_X1 \reg_in_reg[189]  ( .D(Plaintext[189]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[189]) );
  DFFSNQ_X1 \reg_in_reg[188]  ( .D(Plaintext[188]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[188]) );
  DFFSNQ_X1 \reg_in_reg[187]  ( .D(Plaintext[187]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[187]) );
  DFFSNQ_X1 \reg_in_reg[186]  ( .D(Plaintext[186]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[186]) );
  DFFSNQ_X1 \reg_in_reg[184]  ( .D(Plaintext[184]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[184]) );
  DFFSNQ_X1 \reg_in_reg[183]  ( .D(Plaintext[183]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[183]) );
  DFFSNQ_X1 \reg_in_reg[182]  ( .D(Plaintext[182]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[182]) );
  DFFSNQ_X1 \reg_in_reg[181]  ( .D(Plaintext[181]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[181]) );
  DFFSNQ_X1 \reg_in_reg[180]  ( .D(Plaintext[180]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[180]) );
  DFFSNQ_X1 \reg_in_reg[179]  ( .D(Plaintext[179]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[179]) );
  DFFSNQ_X1 \reg_in_reg[178]  ( .D(Plaintext[178]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[178]) );
  DFFSNQ_X1 \reg_in_reg[177]  ( .D(Plaintext[177]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[177]) );
  DFFSNQ_X1 \reg_in_reg[176]  ( .D(Plaintext[176]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[176]) );
  DFFSNQ_X1 \reg_in_reg[175]  ( .D(Plaintext[175]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[175]) );
  DFFSNQ_X1 \reg_in_reg[174]  ( .D(Plaintext[174]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[174]) );
  DFFSNQ_X1 \reg_in_reg[173]  ( .D(Plaintext[173]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[173]) );
  DFFSNQ_X1 \reg_in_reg[172]  ( .D(Plaintext[172]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[172]) );
  DFFSNQ_X1 \reg_in_reg[171]  ( .D(Plaintext[171]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[171]) );
  DFFSNQ_X1 \reg_in_reg[170]  ( .D(Plaintext[170]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[170]) );
  DFFSNQ_X1 \reg_in_reg[169]  ( .D(Plaintext[169]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[169]) );
  DFFSNQ_X1 \reg_in_reg[168]  ( .D(Plaintext[168]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[168]) );
  DFFSNQ_X1 \reg_in_reg[167]  ( .D(Plaintext[167]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[167]) );
  DFFSNQ_X1 \reg_in_reg[166]  ( .D(Plaintext[166]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[166]) );
  DFFSNQ_X1 \reg_in_reg[165]  ( .D(Plaintext[165]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[165]) );
  DFFSNQ_X1 \reg_in_reg[164]  ( .D(Plaintext[164]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[164]) );
  DFFSNQ_X1 \reg_in_reg[163]  ( .D(Plaintext[163]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[163]) );
  DFFSNQ_X1 \reg_in_reg[162]  ( .D(Plaintext[162]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[162]) );
  DFFSNQ_X1 \reg_in_reg[161]  ( .D(Plaintext[161]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[161]) );
  DFFSNQ_X1 \reg_in_reg[160]  ( .D(Plaintext[160]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[160]) );
  DFFSNQ_X1 \reg_in_reg[159]  ( .D(Plaintext[159]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[159]) );
  DFFSNQ_X1 \reg_in_reg[158]  ( .D(Plaintext[158]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[158]) );
  DFFSNQ_X1 \reg_in_reg[157]  ( .D(Plaintext[157]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[157]) );
  DFFSNQ_X1 \reg_in_reg[156]  ( .D(Plaintext[156]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[156]) );
  DFFSNQ_X1 \reg_in_reg[155]  ( .D(Plaintext[155]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[155]) );
  DFFSNQ_X1 \reg_in_reg[154]  ( .D(Plaintext[154]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[154]) );
  DFFSNQ_X1 \reg_in_reg[153]  ( .D(Plaintext[153]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[153]) );
  DFFSNQ_X1 \reg_in_reg[152]  ( .D(Plaintext[152]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[152]) );
  DFFSNQ_X1 \reg_in_reg[151]  ( .D(Plaintext[151]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[151]) );
  DFFSNQ_X1 \reg_in_reg[150]  ( .D(Plaintext[150]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[150]) );
  DFFSNQ_X1 \reg_in_reg[149]  ( .D(Plaintext[149]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[149]) );
  DFFSNQ_X1 \reg_in_reg[148]  ( .D(Plaintext[148]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[148]) );
  DFFSNQ_X1 \reg_in_reg[147]  ( .D(Plaintext[147]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[147]) );
  DFFSNQ_X1 \reg_in_reg[146]  ( .D(Plaintext[146]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[146]) );
  DFFSNQ_X1 \reg_in_reg[145]  ( .D(Plaintext[145]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[145]) );
  DFFSNQ_X1 \reg_in_reg[144]  ( .D(Plaintext[144]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[144]) );
  DFFSNQ_X1 \reg_in_reg[143]  ( .D(Plaintext[143]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[143]) );
  DFFSNQ_X1 \reg_in_reg[142]  ( .D(Plaintext[142]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[142]) );
  DFFSNQ_X1 \reg_in_reg[141]  ( .D(Plaintext[141]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[141]) );
  DFFSNQ_X1 \reg_in_reg[140]  ( .D(Plaintext[140]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[140]) );
  DFFSNQ_X1 \reg_in_reg[139]  ( .D(Plaintext[139]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[139]) );
  DFFSNQ_X1 \reg_in_reg[138]  ( .D(Plaintext[138]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[138]) );
  DFFSNQ_X1 \reg_in_reg[137]  ( .D(Plaintext[137]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[137]) );
  DFFSNQ_X1 \reg_in_reg[136]  ( .D(Plaintext[136]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[136]) );
  DFFSNQ_X1 \reg_in_reg[135]  ( .D(Plaintext[135]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[135]) );
  DFFSNQ_X1 \reg_in_reg[134]  ( .D(Plaintext[134]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[134]) );
  DFFSNQ_X1 \reg_in_reg[133]  ( .D(Plaintext[133]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[133]) );
  DFFSNQ_X1 \reg_in_reg[132]  ( .D(Plaintext[132]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[132]) );
  DFFSNQ_X1 \reg_in_reg[131]  ( .D(Plaintext[131]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[131]) );
  DFFSNQ_X1 \reg_in_reg[130]  ( .D(Plaintext[130]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[130]) );
  DFFSNQ_X1 \reg_in_reg[129]  ( .D(Plaintext[129]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[129]) );
  DFFSNQ_X1 \reg_in_reg[128]  ( .D(Plaintext[128]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[128]) );
  DFFSNQ_X1 \reg_in_reg[127]  ( .D(Plaintext[127]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[127]) );
  DFFSNQ_X1 \reg_in_reg[126]  ( .D(Plaintext[126]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[126]) );
  DFFSNQ_X1 \reg_in_reg[125]  ( .D(Plaintext[125]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[125]) );
  DFFSNQ_X1 \reg_in_reg[124]  ( .D(Plaintext[124]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[124]) );
  DFFSNQ_X1 \reg_in_reg[123]  ( .D(Plaintext[123]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[123]) );
  DFFSNQ_X1 \reg_in_reg[122]  ( .D(Plaintext[122]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[122]) );
  DFFSNQ_X1 \reg_in_reg[121]  ( .D(Plaintext[121]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[121]) );
  DFFSNQ_X1 \reg_in_reg[120]  ( .D(Plaintext[120]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[120]) );
  DFFSNQ_X1 \reg_in_reg[119]  ( .D(Plaintext[119]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[119]) );
  DFFSNQ_X1 \reg_in_reg[118]  ( .D(Plaintext[118]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[118]) );
  DFFSNQ_X1 \reg_in_reg[117]  ( .D(Plaintext[117]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[117]) );
  DFFSNQ_X1 \reg_in_reg[116]  ( .D(Plaintext[116]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[116]) );
  DFFSNQ_X1 \reg_in_reg[115]  ( .D(Plaintext[115]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[115]) );
  DFFSNQ_X1 \reg_in_reg[114]  ( .D(Plaintext[114]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[114]) );
  DFFSNQ_X1 \reg_in_reg[113]  ( .D(Plaintext[113]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[113]) );
  DFFSNQ_X1 \reg_in_reg[112]  ( .D(Plaintext[112]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[112]) );
  DFFSNQ_X1 \reg_in_reg[110]  ( .D(Plaintext[110]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[110]) );
  DFFSNQ_X1 \reg_in_reg[109]  ( .D(Plaintext[109]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[109]) );
  DFFSNQ_X1 \reg_in_reg[108]  ( .D(Plaintext[108]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[108]) );
  DFFSNQ_X1 \reg_in_reg[107]  ( .D(Plaintext[107]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[107]) );
  DFFSNQ_X1 \reg_in_reg[106]  ( .D(Plaintext[106]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[106]) );
  DFFSNQ_X1 \reg_in_reg[105]  ( .D(Plaintext[105]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[105]) );
  DFFSNQ_X1 \reg_in_reg[104]  ( .D(Plaintext[104]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[104]) );
  DFFSNQ_X1 \reg_in_reg[103]  ( .D(Plaintext[103]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[103]) );
  DFFSNQ_X1 \reg_in_reg[102]  ( .D(Plaintext[102]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[102]) );
  DFFSNQ_X1 \reg_in_reg[100]  ( .D(Plaintext[100]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[100]) );
  DFFSNQ_X1 \reg_in_reg[99]  ( .D(Plaintext[99]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[99]) );
  DFFSNQ_X1 \reg_in_reg[98]  ( .D(Plaintext[98]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[98]) );
  DFFSNQ_X1 \reg_in_reg[97]  ( .D(Plaintext[97]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[97]) );
  DFFSNQ_X1 \reg_in_reg[96]  ( .D(Plaintext[96]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[96]) );
  DFFSNQ_X1 \reg_in_reg[95]  ( .D(Plaintext[95]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[95]) );
  DFFSNQ_X1 \reg_in_reg[94]  ( .D(Plaintext[94]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[94]) );
  DFFSNQ_X1 \reg_in_reg[93]  ( .D(Plaintext[93]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[93]) );
  DFFSNQ_X1 \reg_in_reg[92]  ( .D(Plaintext[92]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[92]) );
  DFFSNQ_X1 \reg_in_reg[91]  ( .D(Plaintext[91]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[91]) );
  DFFSNQ_X1 \reg_in_reg[90]  ( .D(Plaintext[90]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[90]) );
  DFFSNQ_X1 \reg_in_reg[89]  ( .D(Plaintext[89]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[89]) );
  DFFSNQ_X1 \reg_in_reg[88]  ( .D(Plaintext[88]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[88]) );
  DFFSNQ_X1 \reg_in_reg[87]  ( .D(Plaintext[87]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[87]) );
  DFFSNQ_X1 \reg_in_reg[86]  ( .D(Plaintext[86]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[86]) );
  DFFSNQ_X1 \reg_in_reg[85]  ( .D(Plaintext[85]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[85]) );
  DFFSNQ_X1 \reg_in_reg[84]  ( .D(Plaintext[84]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[84]) );
  DFFSNQ_X1 \reg_in_reg[82]  ( .D(Plaintext[82]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[82]) );
  DFFSNQ_X1 \reg_in_reg[81]  ( .D(Plaintext[81]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[81]) );
  DFFSNQ_X1 \reg_in_reg[79]  ( .D(Plaintext[79]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[79]) );
  DFFSNQ_X1 \reg_in_reg[78]  ( .D(Plaintext[78]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[78]) );
  DFFSNQ_X1 \reg_in_reg[77]  ( .D(Plaintext[77]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[77]) );
  DFFSNQ_X1 \reg_in_reg[76]  ( .D(Plaintext[76]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[76]) );
  DFFSNQ_X1 \reg_in_reg[75]  ( .D(Plaintext[75]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[75]) );
  DFFSNQ_X1 \reg_in_reg[74]  ( .D(Plaintext[74]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[74]) );
  DFFSNQ_X1 \reg_in_reg[73]  ( .D(Plaintext[73]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[73]) );
  DFFSNQ_X1 \reg_in_reg[72]  ( .D(Plaintext[72]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[72]) );
  DFFSNQ_X1 \reg_in_reg[71]  ( .D(Plaintext[71]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[71]) );
  DFFSNQ_X1 \reg_in_reg[70]  ( .D(Plaintext[70]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[70]) );
  DFFSNQ_X1 \reg_in_reg[69]  ( .D(Plaintext[69]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[69]) );
  DFFSNQ_X1 \reg_in_reg[68]  ( .D(Plaintext[68]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[68]) );
  DFFSNQ_X1 \reg_in_reg[67]  ( .D(Plaintext[67]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[67]) );
  DFFSNQ_X1 \reg_in_reg[66]  ( .D(Plaintext[66]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[66]) );
  DFFSNQ_X1 \reg_in_reg[65]  ( .D(Plaintext[65]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[65]) );
  DFFSNQ_X1 \reg_in_reg[64]  ( .D(Plaintext[64]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[64]) );
  DFFSNQ_X1 \reg_in_reg[63]  ( .D(Plaintext[63]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[63]) );
  DFFSNQ_X1 \reg_in_reg[62]  ( .D(Plaintext[62]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[62]) );
  DFFSNQ_X1 \reg_in_reg[61]  ( .D(Plaintext[61]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[61]) );
  DFFSNQ_X1 \reg_in_reg[60]  ( .D(Plaintext[60]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[60]) );
  DFFSNQ_X1 \reg_in_reg[58]  ( .D(Plaintext[58]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[58]) );
  DFFSNQ_X1 \reg_in_reg[57]  ( .D(Plaintext[57]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[57]) );
  DFFSNQ_X1 \reg_in_reg[56]  ( .D(Plaintext[56]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[56]) );
  DFFSNQ_X1 \reg_in_reg[55]  ( .D(Plaintext[55]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[55]) );
  DFFSNQ_X1 \reg_in_reg[54]  ( .D(Plaintext[54]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[54]) );
  DFFSNQ_X1 \reg_in_reg[53]  ( .D(Plaintext[53]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[53]) );
  DFFSNQ_X1 \reg_in_reg[52]  ( .D(Plaintext[52]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[52]) );
  DFFSNQ_X1 \reg_in_reg[51]  ( .D(Plaintext[51]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[51]) );
  DFFSNQ_X1 \reg_in_reg[50]  ( .D(Plaintext[50]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[50]) );
  DFFSNQ_X1 \reg_in_reg[49]  ( .D(Plaintext[49]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[49]) );
  DFFSNQ_X1 \reg_in_reg[48]  ( .D(Plaintext[48]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[48]) );
  DFFSNQ_X1 \reg_in_reg[47]  ( .D(Plaintext[47]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[47]) );
  DFFSNQ_X1 \reg_in_reg[46]  ( .D(Plaintext[46]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[46]) );
  DFFSNQ_X1 \reg_in_reg[45]  ( .D(Plaintext[45]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[45]) );
  DFFSNQ_X1 \reg_in_reg[44]  ( .D(Plaintext[44]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[44]) );
  DFFSNQ_X1 \reg_in_reg[43]  ( .D(Plaintext[43]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[43]) );
  DFFSNQ_X1 \reg_in_reg[42]  ( .D(Plaintext[42]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[42]) );
  DFFSNQ_X1 \reg_in_reg[41]  ( .D(Plaintext[41]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[41]) );
  DFFSNQ_X1 \reg_in_reg[40]  ( .D(Plaintext[40]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[40]) );
  DFFSNQ_X1 \reg_in_reg[39]  ( .D(Plaintext[39]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[39]) );
  DFFSNQ_X1 \reg_in_reg[38]  ( .D(Plaintext[38]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[38]) );
  DFFSNQ_X1 \reg_in_reg[37]  ( .D(Plaintext[37]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[37]) );
  DFFSNQ_X1 \reg_in_reg[36]  ( .D(Plaintext[36]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[36]) );
  DFFSNQ_X1 \reg_in_reg[35]  ( .D(Plaintext[35]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[35]) );
  DFFSNQ_X1 \reg_in_reg[34]  ( .D(Plaintext[34]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[34]) );
  DFFSNQ_X1 \reg_in_reg[33]  ( .D(Plaintext[33]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[33]) );
  DFFSNQ_X1 \reg_in_reg[32]  ( .D(Plaintext[32]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[32]) );
  DFFSNQ_X1 \reg_in_reg[31]  ( .D(Plaintext[31]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[31]) );
  DFFSNQ_X1 \reg_in_reg[30]  ( .D(Plaintext[30]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[30]) );
  DFFSNQ_X1 \reg_in_reg[29]  ( .D(Plaintext[29]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[29]) );
  DFFSNQ_X1 \reg_in_reg[28]  ( .D(Plaintext[28]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[28]) );
  DFFSNQ_X1 \reg_in_reg[27]  ( .D(Plaintext[27]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[27]) );
  DFFSNQ_X1 \reg_in_reg[26]  ( .D(Plaintext[26]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[26]) );
  DFFSNQ_X1 \reg_in_reg[25]  ( .D(Plaintext[25]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[25]) );
  DFFSNQ_X1 \reg_in_reg[24]  ( .D(Plaintext[24]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[24]) );
  DFFSNQ_X1 \reg_in_reg[23]  ( .D(Plaintext[23]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[23]) );
  DFFSNQ_X1 \reg_in_reg[22]  ( .D(Plaintext[22]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[22]) );
  DFFSNQ_X1 \reg_in_reg[21]  ( .D(Plaintext[21]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[21]) );
  DFFSNQ_X1 \reg_in_reg[20]  ( .D(Plaintext[20]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[20]) );
  DFFSNQ_X1 \reg_in_reg[19]  ( .D(Plaintext[19]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[19]) );
  DFFSNQ_X1 \reg_in_reg[18]  ( .D(Plaintext[18]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[18]) );
  DFFSNQ_X1 \reg_in_reg[17]  ( .D(Plaintext[17]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[17]) );
  DFFSNQ_X1 \reg_in_reg[16]  ( .D(Plaintext[16]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[16]) );
  DFFSNQ_X1 \reg_in_reg[15]  ( .D(Plaintext[15]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[15]) );
  DFFSNQ_X1 \reg_in_reg[14]  ( .D(Plaintext[14]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[14]) );
  DFFSNQ_X1 \reg_in_reg[13]  ( .D(Plaintext[13]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[13]) );
  DFFSNQ_X1 \reg_in_reg[12]  ( .D(Plaintext[12]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[12]) );
  DFFSNQ_X1 \reg_in_reg[11]  ( .D(Plaintext[11]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[11]) );
  DFFSNQ_X1 \reg_in_reg[10]  ( .D(Plaintext[10]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[10]) );
  DFFSNQ_X1 \reg_in_reg[9]  ( .D(Plaintext[9]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[9]) );
  DFFSNQ_X1 \reg_in_reg[8]  ( .D(Plaintext[8]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[8]) );
  DFFSNQ_X1 \reg_in_reg[7]  ( .D(Plaintext[7]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[7]) );
  DFFSNQ_X1 \reg_in_reg[6]  ( .D(Plaintext[6]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[6]) );
  DFFSNQ_X1 \reg_in_reg[5]  ( .D(Plaintext[5]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[5]) );
  DFFSNQ_X1 \reg_in_reg[4]  ( .D(Plaintext[4]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[4]) );
  DFFSNQ_X1 \reg_in_reg[3]  ( .D(Plaintext[3]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[3]) );
  DFFSNQ_X1 \reg_in_reg[2]  ( .D(Plaintext[2]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[2]) );
  DFFSNQ_X1 \reg_in_reg[1]  ( .D(Plaintext[1]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[1]) );
  DFFSNQ_X1 \reg_in_reg[0]  ( .D(Plaintext[0]), .CLK(clk), .SN(1'b1), .Q(
        reg_in[0]) );
  DFFSNQ_X1 \reg_key_reg[191]  ( .D(Key[191]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[191]) );
  DFFSNQ_X1 \reg_key_reg[190]  ( .D(Key[190]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[190]) );
  DFFSNQ_X1 \reg_key_reg[189]  ( .D(Key[189]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[189]) );
  DFFSNQ_X1 \reg_key_reg[188]  ( .D(Key[188]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[188]) );
  DFFSNQ_X1 \reg_key_reg[187]  ( .D(Key[187]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[187]) );
  DFFSNQ_X1 \reg_key_reg[186]  ( .D(Key[186]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[186]) );
  DFFSNQ_X1 \reg_key_reg[185]  ( .D(Key[185]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[185]) );
  DFFSNQ_X1 \reg_key_reg[184]  ( .D(Key[184]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[184]) );
  DFFSNQ_X1 \reg_key_reg[183]  ( .D(Key[183]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[183]) );
  DFFSNQ_X1 \reg_key_reg[182]  ( .D(Key[182]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[182]) );
  DFFSNQ_X1 \reg_key_reg[181]  ( .D(Key[181]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[181]) );
  DFFSNQ_X1 \reg_key_reg[180]  ( .D(Key[180]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[180]) );
  DFFSNQ_X1 \reg_key_reg[179]  ( .D(Key[179]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[179]) );
  DFFSNQ_X1 \reg_key_reg[178]  ( .D(Key[178]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[178]) );
  DFFSNQ_X1 \reg_key_reg[177]  ( .D(Key[177]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[177]) );
  DFFSNQ_X1 \reg_key_reg[176]  ( .D(Key[176]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[176]) );
  DFFSNQ_X1 \reg_key_reg[175]  ( .D(Key[175]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[175]) );
  DFFSNQ_X1 \reg_key_reg[174]  ( .D(Key[174]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[174]) );
  DFFSNQ_X1 \reg_key_reg[173]  ( .D(Key[173]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[173]) );
  DFFSNQ_X1 \reg_key_reg[172]  ( .D(Key[172]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[172]) );
  DFFSNQ_X1 \reg_key_reg[171]  ( .D(Key[171]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[171]) );
  DFFSNQ_X1 \reg_key_reg[170]  ( .D(Key[170]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[170]) );
  DFFSNQ_X1 \reg_key_reg[169]  ( .D(Key[169]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[169]) );
  DFFSNQ_X1 \reg_key_reg[168]  ( .D(Key[168]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[168]) );
  DFFSNQ_X1 \reg_key_reg[167]  ( .D(Key[167]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[167]) );
  DFFSNQ_X1 \reg_key_reg[166]  ( .D(Key[166]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[166]) );
  DFFSNQ_X1 \reg_key_reg[165]  ( .D(Key[165]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[165]) );
  DFFSNQ_X1 \reg_key_reg[164]  ( .D(Key[164]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[164]) );
  DFFSNQ_X1 \reg_key_reg[163]  ( .D(Key[163]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[163]) );
  DFFSNQ_X1 \reg_key_reg[162]  ( .D(Key[162]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[162]) );
  DFFSNQ_X1 \reg_key_reg[161]  ( .D(Key[161]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[161]) );
  DFFSNQ_X1 \reg_key_reg[160]  ( .D(Key[160]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[160]) );
  DFFSNQ_X1 \reg_key_reg[159]  ( .D(Key[159]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[159]) );
  DFFSNQ_X1 \reg_key_reg[158]  ( .D(Key[158]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[158]) );
  DFFSNQ_X1 \reg_key_reg[157]  ( .D(Key[157]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[157]) );
  DFFSNQ_X1 \reg_key_reg[156]  ( .D(Key[156]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[156]) );
  DFFSNQ_X1 \reg_key_reg[155]  ( .D(Key[155]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[155]) );
  DFFSNQ_X1 \reg_key_reg[154]  ( .D(Key[154]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[154]) );
  DFFSNQ_X1 \reg_key_reg[153]  ( .D(Key[153]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[153]) );
  DFFSNQ_X1 \reg_key_reg[152]  ( .D(Key[152]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[152]) );
  DFFSNQ_X1 \reg_key_reg[151]  ( .D(Key[151]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[151]) );
  DFFSNQ_X1 \reg_key_reg[150]  ( .D(Key[150]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[150]) );
  DFFSNQ_X1 \reg_key_reg[149]  ( .D(Key[149]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[149]) );
  DFFSNQ_X1 \reg_key_reg[148]  ( .D(Key[148]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[148]) );
  DFFSNQ_X1 \reg_key_reg[147]  ( .D(Key[147]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[147]) );
  DFFSNQ_X1 \reg_key_reg[146]  ( .D(Key[146]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[146]) );
  DFFSNQ_X1 \reg_key_reg[145]  ( .D(Key[145]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[145]) );
  DFFSNQ_X1 \reg_key_reg[144]  ( .D(Key[144]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[144]) );
  DFFSNQ_X1 \reg_key_reg[143]  ( .D(Key[143]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[143]) );
  DFFSNQ_X1 \reg_key_reg[142]  ( .D(Key[142]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[142]) );
  DFFSNQ_X1 \reg_key_reg[141]  ( .D(Key[141]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[141]) );
  DFFSNQ_X1 \reg_key_reg[140]  ( .D(Key[140]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[140]) );
  DFFSNQ_X1 \reg_key_reg[139]  ( .D(Key[139]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[139]) );
  DFFSNQ_X1 \reg_key_reg[138]  ( .D(Key[138]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[138]) );
  DFFSNQ_X1 \reg_key_reg[137]  ( .D(Key[137]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[137]) );
  DFFSNQ_X1 \reg_key_reg[136]  ( .D(Key[136]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[136]) );
  DFFSNQ_X1 \reg_key_reg[135]  ( .D(Key[135]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[135]) );
  DFFSNQ_X1 \reg_key_reg[134]  ( .D(Key[134]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[134]) );
  DFFSNQ_X1 \reg_key_reg[133]  ( .D(Key[133]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[133]) );
  DFFSNQ_X1 \reg_key_reg[132]  ( .D(Key[132]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[132]) );
  DFFSNQ_X1 \reg_key_reg[131]  ( .D(Key[131]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[131]) );
  DFFSNQ_X1 \reg_key_reg[130]  ( .D(Key[130]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[130]) );
  DFFSNQ_X1 \reg_key_reg[129]  ( .D(Key[129]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[129]) );
  DFFSNQ_X1 \reg_key_reg[128]  ( .D(Key[128]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[128]) );
  DFFSNQ_X1 \reg_key_reg[127]  ( .D(Key[127]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[127]) );
  DFFSNQ_X1 \reg_key_reg[126]  ( .D(Key[126]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[126]) );
  DFFSNQ_X1 \reg_key_reg[125]  ( .D(Key[125]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[125]) );
  DFFSNQ_X1 \reg_key_reg[124]  ( .D(Key[124]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[124]) );
  DFFSNQ_X1 \reg_key_reg[123]  ( .D(Key[123]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[123]) );
  DFFSNQ_X1 \reg_key_reg[122]  ( .D(Key[122]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[122]) );
  DFFSNQ_X1 \reg_key_reg[121]  ( .D(Key[121]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[121]) );
  DFFSNQ_X1 \reg_key_reg[120]  ( .D(Key[120]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[120]) );
  DFFSNQ_X1 \reg_key_reg[119]  ( .D(Key[119]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[119]) );
  DFFSNQ_X1 \reg_key_reg[118]  ( .D(Key[118]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[118]) );
  DFFSNQ_X1 \reg_key_reg[117]  ( .D(Key[117]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[117]) );
  DFFSNQ_X1 \reg_key_reg[116]  ( .D(Key[116]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[116]) );
  DFFSNQ_X1 \reg_key_reg[115]  ( .D(Key[115]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[115]) );
  DFFSNQ_X1 \reg_key_reg[114]  ( .D(Key[114]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[114]) );
  DFFSNQ_X1 \reg_key_reg[113]  ( .D(Key[113]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[113]) );
  DFFSNQ_X1 \reg_key_reg[112]  ( .D(Key[112]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[112]) );
  DFFSNQ_X1 \reg_key_reg[111]  ( .D(Key[111]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[111]) );
  DFFSNQ_X1 \reg_key_reg[110]  ( .D(Key[110]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[110]) );
  DFFSNQ_X1 \reg_key_reg[109]  ( .D(Key[109]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[109]) );
  DFFSNQ_X1 \reg_key_reg[108]  ( .D(Key[108]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[108]) );
  DFFSNQ_X1 \reg_key_reg[107]  ( .D(Key[107]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[107]) );
  DFFSNQ_X1 \reg_key_reg[106]  ( .D(Key[106]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[106]) );
  DFFSNQ_X1 \reg_key_reg[105]  ( .D(Key[105]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[105]) );
  DFFSNQ_X1 \reg_key_reg[104]  ( .D(Key[104]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[104]) );
  DFFSNQ_X1 \reg_key_reg[103]  ( .D(Key[103]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[103]) );
  DFFSNQ_X1 \reg_key_reg[102]  ( .D(Key[102]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[102]) );
  DFFSNQ_X1 \reg_key_reg[101]  ( .D(Key[101]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[101]) );
  DFFSNQ_X1 \reg_key_reg[100]  ( .D(Key[100]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[100]) );
  DFFSNQ_X1 \reg_key_reg[99]  ( .D(Key[99]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[99]) );
  DFFSNQ_X1 \reg_key_reg[98]  ( .D(Key[98]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[98]) );
  DFFSNQ_X1 \reg_key_reg[97]  ( .D(Key[97]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[97]) );
  DFFSNQ_X1 \reg_key_reg[96]  ( .D(Key[96]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[96]) );
  DFFSNQ_X1 \reg_key_reg[95]  ( .D(Key[95]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[95]) );
  DFFSNQ_X1 \reg_key_reg[94]  ( .D(Key[94]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[94]) );
  DFFSNQ_X1 \reg_key_reg[93]  ( .D(Key[93]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[93]) );
  DFFSNQ_X1 \reg_key_reg[92]  ( .D(Key[92]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[92]) );
  DFFSNQ_X1 \reg_key_reg[91]  ( .D(Key[91]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[91]) );
  DFFSNQ_X1 \reg_key_reg[90]  ( .D(Key[90]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[90]) );
  DFFSNQ_X1 \reg_key_reg[89]  ( .D(Key[89]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[89]) );
  DFFSNQ_X1 \reg_key_reg[88]  ( .D(Key[88]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[88]) );
  DFFSNQ_X1 \reg_key_reg[87]  ( .D(Key[87]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[87]) );
  DFFSNQ_X1 \reg_key_reg[86]  ( .D(Key[86]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[86]) );
  DFFSNQ_X1 \reg_key_reg[85]  ( .D(Key[85]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[85]) );
  DFFSNQ_X1 \reg_key_reg[84]  ( .D(Key[84]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[84]) );
  DFFSNQ_X1 \reg_key_reg[83]  ( .D(Key[83]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[83]) );
  DFFSNQ_X1 \reg_key_reg[82]  ( .D(Key[82]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[82]) );
  DFFSNQ_X1 \reg_key_reg[81]  ( .D(Key[81]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[81]) );
  DFFSNQ_X1 \reg_key_reg[80]  ( .D(Key[80]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[80]) );
  DFFSNQ_X1 \reg_key_reg[79]  ( .D(Key[79]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[79]) );
  DFFSNQ_X1 \reg_key_reg[78]  ( .D(Key[78]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[78]) );
  DFFSNQ_X1 \reg_key_reg[77]  ( .D(Key[77]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[77]) );
  DFFSNQ_X1 \reg_key_reg[76]  ( .D(Key[76]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[76]) );
  DFFSNQ_X1 \reg_key_reg[75]  ( .D(Key[75]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[75]) );
  DFFSNQ_X1 \reg_key_reg[74]  ( .D(Key[74]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[74]) );
  DFFSNQ_X1 \reg_key_reg[73]  ( .D(Key[73]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[73]) );
  DFFSNQ_X1 \reg_key_reg[72]  ( .D(Key[72]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[72]) );
  DFFSNQ_X1 \reg_key_reg[71]  ( .D(Key[71]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[71]) );
  DFFSNQ_X1 \reg_key_reg[70]  ( .D(Key[70]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[70]) );
  DFFSNQ_X1 \reg_key_reg[69]  ( .D(Key[69]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[69]) );
  DFFSNQ_X1 \reg_key_reg[68]  ( .D(Key[68]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[68]) );
  DFFSNQ_X1 \reg_key_reg[67]  ( .D(Key[67]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[67]) );
  DFFSNQ_X1 \reg_key_reg[66]  ( .D(Key[66]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[66]) );
  DFFSNQ_X1 \reg_key_reg[65]  ( .D(Key[65]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[65]) );
  DFFSNQ_X1 \reg_key_reg[64]  ( .D(Key[64]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[64]) );
  DFFSNQ_X1 \reg_key_reg[63]  ( .D(Key[63]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[63]) );
  DFFSNQ_X1 \reg_key_reg[62]  ( .D(Key[62]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[62]) );
  DFFSNQ_X1 \reg_key_reg[61]  ( .D(Key[61]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[61]) );
  DFFSNQ_X1 \reg_key_reg[60]  ( .D(Key[60]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[60]) );
  DFFSNQ_X1 \reg_key_reg[59]  ( .D(Key[59]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[59]) );
  DFFSNQ_X1 \reg_key_reg[58]  ( .D(Key[58]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[58]) );
  DFFSNQ_X1 \reg_key_reg[57]  ( .D(Key[57]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[57]) );
  DFFSNQ_X1 \reg_key_reg[56]  ( .D(Key[56]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[56]) );
  DFFSNQ_X1 \reg_key_reg[55]  ( .D(Key[55]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[55]) );
  DFFSNQ_X1 \reg_key_reg[54]  ( .D(Key[54]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[54]) );
  DFFSNQ_X1 \reg_key_reg[53]  ( .D(Key[53]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[53]) );
  DFFSNQ_X1 \reg_key_reg[52]  ( .D(Key[52]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[52]) );
  DFFSNQ_X1 \reg_key_reg[51]  ( .D(Key[51]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[51]) );
  DFFSNQ_X1 \reg_key_reg[50]  ( .D(Key[50]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[50]) );
  DFFSNQ_X1 \reg_key_reg[49]  ( .D(Key[49]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[49]) );
  DFFSNQ_X1 \reg_key_reg[48]  ( .D(Key[48]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[48]) );
  DFFSNQ_X1 \reg_key_reg[46]  ( .D(Key[46]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[46]) );
  DFFSNQ_X1 \reg_key_reg[45]  ( .D(Key[45]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[45]) );
  DFFSNQ_X1 \reg_key_reg[44]  ( .D(Key[44]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[44]) );
  DFFSNQ_X1 \reg_key_reg[43]  ( .D(Key[43]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[43]) );
  DFFSNQ_X1 \reg_key_reg[42]  ( .D(Key[42]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[42]) );
  DFFSNQ_X1 \reg_key_reg[41]  ( .D(Key[41]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[41]) );
  DFFSNQ_X1 \reg_key_reg[40]  ( .D(Key[40]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[40]) );
  DFFSNQ_X1 \reg_key_reg[39]  ( .D(Key[39]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[39]) );
  DFFSNQ_X1 \reg_key_reg[38]  ( .D(Key[38]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[38]) );
  DFFSNQ_X1 \reg_key_reg[37]  ( .D(Key[37]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[37]) );
  DFFSNQ_X1 \reg_key_reg[36]  ( .D(Key[36]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[36]) );
  DFFSNQ_X1 \reg_key_reg[35]  ( .D(Key[35]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[35]) );
  DFFSNQ_X1 \reg_key_reg[34]  ( .D(Key[34]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[34]) );
  DFFSNQ_X1 \reg_key_reg[33]  ( .D(Key[33]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[33]) );
  DFFSNQ_X1 \reg_key_reg[32]  ( .D(Key[32]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[32]) );
  DFFSNQ_X1 \reg_key_reg[31]  ( .D(Key[31]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[31]) );
  DFFSNQ_X1 \reg_key_reg[30]  ( .D(Key[30]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[30]) );
  DFFSNQ_X1 \reg_key_reg[29]  ( .D(Key[29]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[29]) );
  DFFSNQ_X1 \reg_key_reg[28]  ( .D(Key[28]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[28]) );
  DFFSNQ_X1 \reg_key_reg[27]  ( .D(Key[27]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[27]) );
  DFFSNQ_X1 \reg_key_reg[26]  ( .D(Key[26]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[26]) );
  DFFSNQ_X1 \reg_key_reg[25]  ( .D(Key[25]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[25]) );
  DFFSNQ_X1 \reg_key_reg[24]  ( .D(Key[24]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[24]) );
  DFFSNQ_X1 \reg_key_reg[23]  ( .D(Key[23]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[23]) );
  DFFSNQ_X1 \reg_key_reg[22]  ( .D(Key[22]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[22]) );
  DFFSNQ_X1 \reg_key_reg[21]  ( .D(Key[21]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[21]) );
  DFFSNQ_X1 \reg_key_reg[20]  ( .D(Key[20]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[20]) );
  DFFSNQ_X1 \reg_key_reg[19]  ( .D(Key[19]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[19]) );
  DFFSNQ_X1 \reg_key_reg[18]  ( .D(Key[18]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[18]) );
  DFFSNQ_X1 \reg_key_reg[17]  ( .D(Key[17]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[17]) );
  DFFSNQ_X1 \reg_key_reg[16]  ( .D(Key[16]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[16]) );
  DFFSNQ_X1 \reg_key_reg[15]  ( .D(Key[15]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[15]) );
  DFFSNQ_X1 \reg_key_reg[13]  ( .D(Key[13]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[13]) );
  DFFSNQ_X1 \reg_key_reg[12]  ( .D(Key[12]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[12]) );
  DFFSNQ_X1 \reg_key_reg[11]  ( .D(Key[11]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[11]) );
  DFFSNQ_X1 \reg_key_reg[10]  ( .D(Key[10]), .CLK(clk), .SN(1'b1), .Q(
        reg_key[10]) );
  DFFSNQ_X1 \reg_key_reg[9]  ( .D(Key[9]), .CLK(clk), .SN(1'b1), .Q(reg_key[9]) );
  DFFSNQ_X1 \reg_key_reg[7]  ( .D(Key[7]), .CLK(clk), .SN(1'b1), .Q(reg_key[7]) );
  DFFSNQ_X1 \reg_key_reg[6]  ( .D(Key[6]), .CLK(clk), .SN(1'b1), .Q(reg_key[6]) );
  DFFSNQ_X1 \reg_key_reg[5]  ( .D(Key[5]), .CLK(clk), .SN(1'b1), .Q(reg_key[5]) );
  DFFSNQ_X1 \reg_key_reg[4]  ( .D(Key[4]), .CLK(clk), .SN(1'b1), .Q(reg_key[4]) );
  DFFSNQ_X1 \reg_key_reg[3]  ( .D(Key[3]), .CLK(clk), .SN(1'b1), .Q(reg_key[3]) );
  DFFSNQ_X1 \reg_key_reg[2]  ( .D(Key[2]), .CLK(clk), .SN(1'b1), .Q(reg_key[2]) );
  DFFSNQ_X1 \reg_key_reg[1]  ( .D(Key[1]), .CLK(clk), .SN(1'b1), .Q(reg_key[1]) );
  DFFSNQ_X1 \reg_key_reg[0]  ( .D(Key[0]), .CLK(clk), .SN(1'b1), .Q(reg_key[0]) );
  DFFSNQ_X1 \Ciphertext_reg[190]  ( .D(reg_out[190]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[190]) );
  DFFSNQ_X1 \Ciphertext_reg[188]  ( .D(reg_out[188]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[188]) );
  DFFSNQ_X1 \Ciphertext_reg[184]  ( .D(reg_out[184]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[184]) );
  DFFSNQ_X1 \Ciphertext_reg[183]  ( .D(reg_out[183]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[183]) );
  DFFSNQ_X1 \Ciphertext_reg[172]  ( .D(reg_out[172]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[172]) );
  DFFSNQ_X1 \Ciphertext_reg[170]  ( .D(reg_out[170]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[170]) );
  DFFSNQ_X1 \Ciphertext_reg[169]  ( .D(reg_out[169]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[169]) );
  DFFSNQ_X1 \Ciphertext_reg[166]  ( .D(reg_out[166]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[166]) );
  DFFSNQ_X1 \Ciphertext_reg[165]  ( .D(reg_out[165]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[165]) );
  DFFSNQ_X1 \Ciphertext_reg[164]  ( .D(reg_out[164]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[164]) );
  DFFSNQ_X1 \Ciphertext_reg[163]  ( .D(reg_out[163]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[163]) );
  DFFSNQ_X1 \Ciphertext_reg[160]  ( .D(reg_out[160]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[160]) );
  DFFSNQ_X1 \Ciphertext_reg[156]  ( .D(reg_out[156]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[156]) );
  DFFSNQ_X1 \Ciphertext_reg[155]  ( .D(reg_out[155]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[155]) );
  DFFSNQ_X1 \Ciphertext_reg[154]  ( .D(reg_out[154]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[154]) );
  DFFSNQ_X1 \Ciphertext_reg[153]  ( .D(reg_out[153]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[153]) );
  DFFSNQ_X1 \Ciphertext_reg[150]  ( .D(reg_out[150]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[150]) );
  DFFSNQ_X1 \Ciphertext_reg[148]  ( .D(reg_out[148]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[148]) );
  DFFSNQ_X1 \Ciphertext_reg[144]  ( .D(reg_out[144]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[144]) );
  DFFSNQ_X1 \Ciphertext_reg[141]  ( .D(reg_out[141]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[141]) );
  DFFSNQ_X1 \Ciphertext_reg[140]  ( .D(reg_out[140]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[140]) );
  DFFSNQ_X1 \Ciphertext_reg[138]  ( .D(reg_out[138]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[138]) );
  DFFSNQ_X1 \Ciphertext_reg[136]  ( .D(reg_out[136]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[136]) );
  DFFSNQ_X1 \Ciphertext_reg[119]  ( .D(reg_out[119]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[119]) );
  DFFSNQ_X1 \Ciphertext_reg[118]  ( .D(reg_out[118]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[118]) );
  DFFSNQ_X1 \Ciphertext_reg[108]  ( .D(reg_out[108]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[108]) );
  DFFSNQ_X1 \Ciphertext_reg[107]  ( .D(reg_out[107]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[107]) );
  DFFSNQ_X1 \Ciphertext_reg[103]  ( .D(reg_out[103]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[103]) );
  DFFSNQ_X1 \Ciphertext_reg[99]  ( .D(reg_out[99]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[99]) );
  DFFSNQ_X1 \Ciphertext_reg[95]  ( .D(reg_out[95]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[95]) );
  DFFSNQ_X1 \Ciphertext_reg[94]  ( .D(reg_out[94]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[94]) );
  DFFSNQ_X1 \Ciphertext_reg[93]  ( .D(reg_out[93]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[93]) );
  DFFSNQ_X1 \Ciphertext_reg[92]  ( .D(reg_out[92]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[92]) );
  DFFSNQ_X1 \Ciphertext_reg[91]  ( .D(reg_out[91]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[91]) );
  DFFSNQ_X1 \Ciphertext_reg[89]  ( .D(reg_out[89]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[89]) );
  DFFSNQ_X1 \Ciphertext_reg[87]  ( .D(reg_out[87]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[87]) );
  DFFSNQ_X1 \Ciphertext_reg[85]  ( .D(reg_out[85]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[85]) );
  DFFSNQ_X1 \Ciphertext_reg[82]  ( .D(reg_out[82]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[82]) );
  DFFSNQ_X1 \Ciphertext_reg[81]  ( .D(reg_out[81]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[81]) );
  DFFSNQ_X1 \Ciphertext_reg[79]  ( .D(reg_out[79]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[79]) );
  DFFSNQ_X1 \Ciphertext_reg[76]  ( .D(reg_out[76]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[76]) );
  DFFSNQ_X1 \Ciphertext_reg[75]  ( .D(reg_out[75]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[75]) );
  DFFSNQ_X1 \Ciphertext_reg[72]  ( .D(reg_out[72]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[72]) );
  DFFSNQ_X1 \Ciphertext_reg[70]  ( .D(reg_out[70]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[70]) );
  DFFSNQ_X1 \Ciphertext_reg[69]  ( .D(reg_out[69]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[69]) );
  DFFSNQ_X1 \Ciphertext_reg[68]  ( .D(reg_out[68]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[68]) );
  DFFSNQ_X1 \Ciphertext_reg[65]  ( .D(reg_out[65]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[65]) );
  DFFSNQ_X1 \Ciphertext_reg[64]  ( .D(reg_out[64]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[64]) );
  DFFSNQ_X1 \Ciphertext_reg[63]  ( .D(reg_out[63]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[63]) );
  DFFSNQ_X1 \Ciphertext_reg[62]  ( .D(reg_out[62]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[62]) );
  DFFSNQ_X1 \Ciphertext_reg[58]  ( .D(reg_out[58]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[58]) );
  DFFSNQ_X1 \Ciphertext_reg[54]  ( .D(reg_out[54]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[54]) );
  DFFSNQ_X1 \Ciphertext_reg[53]  ( .D(reg_out[53]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[53]) );
  DFFSNQ_X1 \Ciphertext_reg[52]  ( .D(reg_out[52]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[52]) );
  DFFSNQ_X1 \Ciphertext_reg[50]  ( .D(reg_out[50]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[50]) );
  DFFSNQ_X1 \Ciphertext_reg[47]  ( .D(reg_out[47]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[47]) );
  DFFSNQ_X1 \Ciphertext_reg[45]  ( .D(reg_out[45]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[45]) );
  DFFSNQ_X1 \Ciphertext_reg[33]  ( .D(reg_out[33]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[33]) );
  DFFSNQ_X1 \Ciphertext_reg[32]  ( .D(reg_out[32]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[32]) );
  DFFSNQ_X1 \Ciphertext_reg[28]  ( .D(reg_out[28]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[28]) );
  DFFSNQ_X1 \Ciphertext_reg[26]  ( .D(reg_out[26]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[26]) );
  DFFSNQ_X1 \Ciphertext_reg[23]  ( .D(reg_out[23]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[23]) );
  DFFSNQ_X1 \Ciphertext_reg[20]  ( .D(reg_out[20]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[20]) );
  DFFSNQ_X1 \Ciphertext_reg[19]  ( .D(reg_out[19]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[19]) );
  DFFSNQ_X1 \Ciphertext_reg[18]  ( .D(reg_out[18]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[18]) );
  DFFSNQ_X1 \Ciphertext_reg[15]  ( .D(reg_out[15]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[15]) );
  DFFSNQ_X1 \Ciphertext_reg[11]  ( .D(reg_out[11]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[11]) );
  DFFSNQ_X1 \Ciphertext_reg[10]  ( .D(reg_out[10]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[10]) );
  DFFSNQ_X1 \Ciphertext_reg[9]  ( .D(reg_out[9]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[9]) );
  DFFSNQ_X1 \Ciphertext_reg[8]  ( .D(reg_out[8]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[8]) );
  DFFSNQ_X1 \Ciphertext_reg[4]  ( .D(reg_out[4]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[4]) );
  DFFRNQ_X1 \Ciphertext_reg[17]  ( .D(reg_out[17]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[17]) );
  DFFRNQ_X1 \Ciphertext_reg[112]  ( .D(reg_out[112]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[112]) );
  DFFRNQ_X1 \Ciphertext_reg[174]  ( .D(reg_out[174]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[174]) );
  DFFRNQ_X1 \Ciphertext_reg[105]  ( .D(reg_out[105]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[105]) );
  DFFRNQ_X1 \Ciphertext_reg[181]  ( .D(reg_out[181]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[181]) );
  DFFRNQ_X1 \Ciphertext_reg[36]  ( .D(reg_out[36]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[36]) );
  DFFRNQ_X1 \Ciphertext_reg[34]  ( .D(reg_out[34]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[34]) );
  DFFRNQ_X1 \Ciphertext_reg[106]  ( .D(reg_out[106]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[106]) );
  DFFRNQ_X1 \Ciphertext_reg[41]  ( .D(reg_out[41]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[41]) );
  DFFRNQ_X1 \Ciphertext_reg[157]  ( .D(reg_out[157]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[157]) );
  DFFRNQ_X1 \Ciphertext_reg[145]  ( .D(reg_out[145]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[145]) );
  DFFRNQ_X1 \Ciphertext_reg[114]  ( .D(reg_out[114]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[114]) );
  DFFRNQ_X1 \Ciphertext_reg[14]  ( .D(reg_out[14]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[14]) );
  DFFRNQ_X1 \Ciphertext_reg[122]  ( .D(reg_out[122]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[122]) );
  DFFRNQ_X1 \Ciphertext_reg[124]  ( .D(reg_out[124]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[124]) );
  DFFRNQ_X1 \Ciphertext_reg[88]  ( .D(reg_out[88]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[88]) );
  DFFRNQ_X1 \Ciphertext_reg[29]  ( .D(reg_out[29]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[29]) );
  DFFRNQ_X1 \Ciphertext_reg[42]  ( .D(reg_out[42]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[42]) );
  DFFRNQ_X1 \Ciphertext_reg[176]  ( .D(reg_out[176]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[176]) );
  DFFRNQ_X1 \Ciphertext_reg[98]  ( .D(reg_out[98]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[98]) );
  DFFRNQ_X1 \Ciphertext_reg[111]  ( .D(reg_out[111]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[111]) );
  DFFRNQ_X1 \Ciphertext_reg[37]  ( .D(reg_out[37]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[37]) );
  DFFRNQ_X1 \Ciphertext_reg[143]  ( .D(reg_out[143]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[143]) );
  DFFRNQ_X1 \Ciphertext_reg[130]  ( .D(reg_out[130]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[130]) );
  DFFRNQ_X1 \Ciphertext_reg[59]  ( .D(reg_out[59]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[59]) );
  DFFRNQ_X1 \Ciphertext_reg[129]  ( .D(reg_out[129]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[129]) );
  DFFRNQ_X1 \Ciphertext_reg[13]  ( .D(reg_out[13]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[13]) );
  DFFRNQ_X1 \Ciphertext_reg[115]  ( .D(reg_out[115]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[115]) );
  DFFRNQ_X1 \Ciphertext_reg[177]  ( .D(reg_out[177]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[177]) );
  DFFRNQ_X1 \Ciphertext_reg[44]  ( .D(reg_out[44]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[44]) );
  DFFRNQ_X1 \Ciphertext_reg[55]  ( .D(reg_out[55]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[55]) );
  DFFRNQ_X1 \Ciphertext_reg[116]  ( .D(reg_out[116]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[116]) );
  DFFRNQ_X1 \Ciphertext_reg[40]  ( .D(reg_out[40]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[40]) );
  DFFRNQ_X1 \Ciphertext_reg[25]  ( .D(reg_out[25]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[25]) );
  DFFRNQ_X1 \Ciphertext_reg[187]  ( .D(reg_out[187]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[187]) );
  DFFRNQ_X1 \Ciphertext_reg[38]  ( .D(reg_out[38]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[38]) );
  DFFRNQ_X1 \Ciphertext_reg[83]  ( .D(reg_out[83]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[83]) );
  DFFRNQ_X1 \Ciphertext_reg[30]  ( .D(reg_out[30]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[30]) );
  DFFRNQ_X1 \Ciphertext_reg[185]  ( .D(reg_out[185]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[185]) );
  DFFRNQ_X1 \Ciphertext_reg[178]  ( .D(reg_out[178]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[178]) );
  DFFRNQ_X1 \Ciphertext_reg[120]  ( .D(reg_out[120]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[120]) );
  DFFRNQ_X1 \Ciphertext_reg[133]  ( .D(reg_out[133]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[133]) );
  DFFRNQ_X1 \Ciphertext_reg[24]  ( .D(reg_out[24]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[24]) );
  DFFRNQ_X1 \Ciphertext_reg[123]  ( .D(reg_out[123]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[123]) );
  DFFRNQ_X1 \Ciphertext_reg[101]  ( .D(reg_out[101]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[101]) );
  DFFRNQ_X1 \Ciphertext_reg[167]  ( .D(reg_out[167]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[167]) );
  DFFRNQ_X1 \Ciphertext_reg[2]  ( .D(reg_out[2]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[2]) );
  DFFRNQ_X1 \Ciphertext_reg[158]  ( .D(reg_out[158]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[158]) );
  DFFRNQ_X1 \Ciphertext_reg[125]  ( .D(reg_out[125]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[125]) );
  DFFRNQ_X1 \Ciphertext_reg[121]  ( .D(reg_out[121]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[121]) );
  DFFRNQ_X1 \Ciphertext_reg[102]  ( .D(reg_out[102]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[102]) );
  DFFRNQ_X1 \Ciphertext_reg[131]  ( .D(reg_out[131]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[131]) );
  DFFRNQ_X1 \Ciphertext_reg[66]  ( .D(reg_out[66]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[66]) );
  DFFRNQ_X1 \Ciphertext_reg[22]  ( .D(reg_out[22]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[22]) );
  DFFRNQ_X1 \Ciphertext_reg[182]  ( .D(reg_out[182]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[182]) );
  DFFRNQ_X1 \Ciphertext_reg[97]  ( .D(reg_out[97]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[97]) );
  DFFRNQ_X1 \Ciphertext_reg[180]  ( .D(reg_out[180]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[180]) );
  DFFRNQ_X1 \Ciphertext_reg[73]  ( .D(reg_out[73]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[73]) );
  DFFRNQ_X1 \Ciphertext_reg[117]  ( .D(reg_out[117]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[117]) );
  DFFRNQ_X1 \Ciphertext_reg[78]  ( .D(reg_out[78]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[78]) );
  DFFRNQ_X1 \Ciphertext_reg[152]  ( .D(reg_out[152]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[152]) );
  DFFRNQ_X1 \Ciphertext_reg[39]  ( .D(reg_out[39]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[39]) );
  DFFRNQ_X1 \Ciphertext_reg[74]  ( .D(reg_out[74]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[74]) );
  DFFRNQ_X1 \Ciphertext_reg[179]  ( .D(reg_out[179]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[179]) );
  DFFRNQ_X1 \Ciphertext_reg[132]  ( .D(reg_out[132]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[132]) );
  DFFRNQ_X1 \Ciphertext_reg[109]  ( .D(reg_out[109]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[109]) );
  DFFRNQ_X1 \Ciphertext_reg[61]  ( .D(reg_out[61]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[61]) );
  DFFRNQ_X1 \Ciphertext_reg[16]  ( .D(reg_out[16]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[16]) );
  DFFRNQ_X1 \Ciphertext_reg[134]  ( .D(reg_out[134]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[134]) );
  DFFRNQ_X1 \Ciphertext_reg[80]  ( .D(reg_out[80]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[80]) );
  DFFRNQ_X1 \Ciphertext_reg[46]  ( .D(reg_out[46]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[46]) );
  DFFRNQ_X1 \Ciphertext_reg[43]  ( .D(reg_out[43]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[43]) );
  DFFRNQ_X1 \Ciphertext_reg[7]  ( .D(reg_out[7]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[7]) );
  DFFRNQ_X1 \Ciphertext_reg[110]  ( .D(reg_out[110]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[110]) );
  DFFRNQ_X1 \Ciphertext_reg[149]  ( .D(reg_out[149]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[149]) );
  DFFRNQ_X1 \Ciphertext_reg[175]  ( .D(reg_out[175]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[175]) );
  DFFRNQ_X1 \Ciphertext_reg[128]  ( .D(reg_out[128]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[128]) );
  DFFRNQ_X1 \Ciphertext_reg[127]  ( .D(reg_out[127]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[127]) );
  DFFRNQ_X1 \Ciphertext_reg[31]  ( .D(reg_out[31]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[31]) );
  DFFRNQ_X1 \Ciphertext_reg[96]  ( .D(reg_out[96]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[96]) );
  DFFRNQ_X1 \Ciphertext_reg[113]  ( .D(reg_out[113]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[113]) );
  DFFRNQ_X1 \Ciphertext_reg[6]  ( .D(reg_out[6]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[6]) );
  DFFRNQ_X1 \Ciphertext_reg[191]  ( .D(reg_out[191]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[191]) );
  DFFRNQ_X1 \Ciphertext_reg[77]  ( .D(reg_out[77]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[77]) );
  DFFRNQ_X1 \Ciphertext_reg[104]  ( .D(reg_out[104]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[104]) );
  DFFRNQ_X1 \Ciphertext_reg[71]  ( .D(reg_out[71]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[71]) );
  DFFRNQ_X1 \Ciphertext_reg[1]  ( .D(reg_out[1]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[1]) );
  DFFRNQ_X1 \Ciphertext_reg[60]  ( .D(reg_out[60]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[60]) );
  DFFRNQ_X1 \Ciphertext_reg[86]  ( .D(reg_out[86]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[86]) );
  DFFRNQ_X1 \Ciphertext_reg[139]  ( .D(reg_out[139]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[139]) );
  DFFRNQ_X1 \Ciphertext_reg[49]  ( .D(reg_out[49]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[49]) );
  DFFRNQ_X1 \Ciphertext_reg[173]  ( .D(reg_out[173]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[173]) );
  DFFRNQ_X1 \Ciphertext_reg[84]  ( .D(reg_out[84]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[84]) );
  DFFRNQ_X1 \Ciphertext_reg[35]  ( .D(reg_out[35]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[35]) );
  DFFRNQ_X1 \Ciphertext_reg[12]  ( .D(reg_out[12]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[12]) );
  DFFRNQ_X1 \Ciphertext_reg[146]  ( .D(reg_out[146]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[146]) );
  DFFRNQ_X1 \Ciphertext_reg[189]  ( .D(reg_out[189]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[189]) );
  DFFRNQ_X1 \Ciphertext_reg[137]  ( .D(reg_out[137]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[137]) );
  DFFRNQ_X1 \Ciphertext_reg[3]  ( .D(reg_out[3]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[3]) );
  DFFRNQ_X1 \Ciphertext_reg[142]  ( .D(reg_out[142]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[142]) );
  DFFRNQ_X1 \Ciphertext_reg[126]  ( .D(reg_out[126]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[126]) );
  DFFRNQ_X1 \Ciphertext_reg[162]  ( .D(reg_out[162]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[162]) );
  DFFRNQ_X1 \Ciphertext_reg[56]  ( .D(reg_out[56]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[56]) );
  DFFRNQ_X1 \Ciphertext_reg[5]  ( .D(reg_out[5]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[5]) );
  DFFRNQ_X1 \Ciphertext_reg[135]  ( .D(reg_out[135]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[135]) );
  DFFRNQ_X1 \Ciphertext_reg[57]  ( .D(reg_out[57]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[57]) );
  DFFRNQ_X1 \Ciphertext_reg[27]  ( .D(reg_out[27]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[27]) );
  DFFRNQ_X1 \Ciphertext_reg[90]  ( .D(reg_out[90]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[90]) );
  DFFRNQ_X1 \reg_key_reg[47]  ( .D(Key[47]), .CLK(clk), .RN(1'b1), .Q(
        reg_key[47]) );
  DFFRNQ_X1 \Ciphertext_reg[0]  ( .D(reg_out[0]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[0]) );
  DFFRNQ_X1 \Ciphertext_reg[151]  ( .D(reg_out[151]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[151]) );
  DFFRNQ_X1 \reg_in_reg[101]  ( .D(Plaintext[101]), .CLK(clk), .RN(1'b1), .Q(
        reg_in[101]) );
  DFFRNQ_X1 \reg_in_reg[59]  ( .D(Plaintext[59]), .CLK(clk), .RN(1'b1), .Q(
        reg_in[59]) );
  DFFSNQ_X1 \Ciphertext_reg[161]  ( .D(reg_out[161]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[161]) );
  DFFSNQ_X1 \Ciphertext_reg[67]  ( .D(reg_out[67]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[67]) );
  DFFSNQ_X1 \Ciphertext_reg[48]  ( .D(reg_out[48]), .CLK(clk), .SN(1'b1), .Q(
        Ciphertext[48]) );
  DFFRNQ_X1 \reg_in_reg[80]  ( .D(Plaintext[80]), .CLK(clk), .RN(1'b1), .Q(
        reg_in[80]) );
  DFFRNQ_X1 \reg_key_reg[14]  ( .D(Key[14]), .CLK(clk), .RN(1'b1), .Q(
        reg_key[14]) );
  DFFRNQ_X1 \reg_in_reg[185]  ( .D(Plaintext[185]), .CLK(clk), .RN(1'b1), .Q(
        reg_in[185]) );
  DFFRNQ_X1 \Ciphertext_reg[168]  ( .D(reg_out[168]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[168]) );
  SPEEDY_Rounds6_0 SPEEDY_instance ( .Plaintext(reg_in), .Key(reg_key), 
        .Ciphertext(reg_out) );
  DFFRNQ_X1 \Ciphertext_reg[186]  ( .D(reg_out[186]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[186]) );
  DFFRNQ_X1 \Ciphertext_reg[147]  ( .D(reg_out[147]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[147]) );
  DFFRNQ_X1 \Ciphertext_reg[21]  ( .D(reg_out[21]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[21]) );
  DFFSNQ_X1 \reg_key_reg[8]  ( .D(Key[8]), .CLK(clk), .SN(1'b1), .Q(reg_key[8]) );
  DFFRNQ_X1 \reg_in_reg[111]  ( .D(Plaintext[111]), .CLK(clk), .RN(1'b1), .Q(
        reg_in[111]) );
  DFFSNQ_X1 \Ciphertext_reg[100]  ( .D(reg_out[100]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[100]) );
  DFFRNQ_X1 \Ciphertext_reg[51]  ( .D(reg_out[51]), .CLK(clk), .RN(1'b1), .Q(
        Ciphertext[51]) );
  DFFSNQ_X1 \Ciphertext_reg[159]  ( .D(reg_out[159]), .CLK(clk), .SN(1'b1), 
        .Q(Ciphertext[159]) );
  DFFRNQ_X1 \Ciphertext_reg[171]  ( .D(reg_out[171]), .CLK(clk), .RN(1'b1), 
        .Q(Ciphertext[171]) );
  DFFRNQ_X1 \reg_in_reg[83]  ( .D(Plaintext[83]), .CLK(clk), .RN(1'b1), .Q(
        reg_in[83]) );
endmodule

